* File: sky130_fd_sc_hs__bufinv_8.pex.spice
* Created: Thu Aug 27 20:35:14 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HS__BUFINV_8%A 1 3 6 8 12
c30 6 0 7.51347e-20 $X=0.51 $Y=0.74
r31 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.385
+ $Y=1.515 $X2=0.385 $Y2=1.515
r32 8 12 4.06745 $w=4.23e-07 $l=1.5e-07 $layer=LI1_cond $X=0.337 $Y=1.665
+ $X2=0.337 $Y2=1.515
r33 4 11 38.6365 $w=3.35e-07 $l=2.10286e-07 $layer=POLY_cond $X=0.51 $Y=1.35
+ $X2=0.407 $Y2=1.515
r34 4 6 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=0.51 $Y=1.35 $X2=0.51
+ $Y2=0.74
r35 1 11 50.8664 $w=3.35e-07 $l=2.94958e-07 $layer=POLY_cond $X=0.505 $Y=1.765
+ $X2=0.407 $Y2=1.515
r36 1 3 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.505 $Y=1.765
+ $X2=0.505 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_HS__BUFINV_8%A_183_48# 1 2 3 4 15 17 19 22 24 26 27 29
+ 32 34 36 39 41 43 46 48 50 53 55 57 60 62 64 67 69 78 83 85 86 87 91 96 99 106
+ 107 108 125
c226 69 0 1.04254e-19 $X=4.65 $Y=1.465
c227 62 0 7.6204e-20 $X=4.285 $Y=1.765
c228 27 0 1.57415e-19 $X=1.905 $Y=1.765
c229 17 0 1.10108e-19 $X=1.005 $Y=1.765
r230 125 126 1.87306 $w=3.86e-07 $l=1.5e-08 $layer=POLY_cond $X=4.285 $Y=1.532
+ $X2=4.3 $Y2=1.532
r231 122 123 11.8627 $w=3.86e-07 $l=9.5e-08 $layer=POLY_cond $X=3.705 $Y=1.532
+ $X2=3.8 $Y2=1.532
r232 121 122 50.5725 $w=3.86e-07 $l=4.05e-07 $layer=POLY_cond $X=3.3 $Y=1.532
+ $X2=3.705 $Y2=1.532
r233 120 121 5.61917 $w=3.86e-07 $l=4.5e-08 $layer=POLY_cond $X=3.255 $Y=1.532
+ $X2=3.3 $Y2=1.532
r234 119 120 48.0751 $w=3.86e-07 $l=3.85e-07 $layer=POLY_cond $X=2.87 $Y=1.532
+ $X2=3.255 $Y2=1.532
r235 118 119 8.11658 $w=3.86e-07 $l=6.5e-08 $layer=POLY_cond $X=2.805 $Y=1.532
+ $X2=2.87 $Y2=1.532
r236 117 118 54.3187 $w=3.86e-07 $l=4.35e-07 $layer=POLY_cond $X=2.37 $Y=1.532
+ $X2=2.805 $Y2=1.532
r237 116 117 1.87306 $w=3.86e-07 $l=1.5e-08 $layer=POLY_cond $X=2.355 $Y=1.532
+ $X2=2.37 $Y2=1.532
r238 115 116 51.8212 $w=3.86e-07 $l=4.15e-07 $layer=POLY_cond $X=1.94 $Y=1.532
+ $X2=2.355 $Y2=1.532
r239 114 115 4.37047 $w=3.86e-07 $l=3.5e-08 $layer=POLY_cond $X=1.905 $Y=1.532
+ $X2=1.94 $Y2=1.532
r240 111 112 1.87306 $w=3.86e-07 $l=1.5e-08 $layer=POLY_cond $X=1.44 $Y=1.532
+ $X2=1.455 $Y2=1.532
r241 110 111 54.3187 $w=3.86e-07 $l=4.35e-07 $layer=POLY_cond $X=1.005 $Y=1.532
+ $X2=1.44 $Y2=1.532
r242 109 110 1.87306 $w=3.86e-07 $l=1.5e-08 $layer=POLY_cond $X=0.99 $Y=1.532
+ $X2=1.005 $Y2=1.532
r243 101 104 13.1378 $w=2.48e-07 $l=2.85e-07 $layer=LI1_cond $X=4.735 $Y=1.005
+ $X2=5.02 $Y2=1.005
r244 97 108 3.10218 $w=3.05e-07 $l=9.66954e-08 $layer=LI1_cond $X=5.985 $Y=2.31
+ $X2=5.96 $Y2=2.225
r245 97 99 3.70428 $w=2.78e-07 $l=9e-08 $layer=LI1_cond $X=5.985 $Y=2.31
+ $X2=5.985 $Y2=2.4
r246 94 108 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=5.96 $Y=2.14
+ $X2=5.96 $Y2=2.225
r247 94 96 5.41299 $w=3.28e-07 $l=1.55e-07 $layer=LI1_cond $X=5.96 $Y=2.14
+ $X2=5.96 $Y2=1.985
r248 93 107 4.07664 $w=3.3e-07 $l=1.25e-07 $layer=LI1_cond $X=5.96 $Y=1.13
+ $X2=5.96 $Y2=1.005
r249 93 96 29.8588 $w=3.28e-07 $l=8.55e-07 $layer=LI1_cond $X=5.96 $Y=1.13
+ $X2=5.96 $Y2=1.985
r250 89 107 4.07664 $w=3.3e-07 $l=1.25e-07 $layer=LI1_cond $X=5.96 $Y=0.88
+ $X2=5.96 $Y2=1.005
r251 89 91 12.7467 $w=3.28e-07 $l=3.65e-07 $layer=LI1_cond $X=5.96 $Y=0.88
+ $X2=5.96 $Y2=0.515
r252 88 106 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.175 $Y=2.225
+ $X2=5.01 $Y2=2.225
r253 87 108 3.51065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.795 $Y=2.225
+ $X2=5.96 $Y2=2.225
r254 87 88 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=5.795 $Y=2.225
+ $X2=5.175 $Y2=2.225
r255 86 104 4.84026 $w=2.48e-07 $l=1.05e-07 $layer=LI1_cond $X=5.125 $Y=1.005
+ $X2=5.02 $Y2=1.005
r256 85 107 2.3589 $w=2.5e-07 $l=1.65e-07 $layer=LI1_cond $X=5.795 $Y=1.005
+ $X2=5.96 $Y2=1.005
r257 85 86 30.8855 $w=2.48e-07 $l=6.7e-07 $layer=LI1_cond $X=5.795 $Y=1.005
+ $X2=5.125 $Y2=1.005
r258 81 104 1.92597 $w=2.05e-07 $l=1.25996e-07 $layer=LI1_cond $X=5.022 $Y=0.88
+ $X2=5.02 $Y2=1.005
r259 81 83 19.7472 $w=2.03e-07 $l=3.65e-07 $layer=LI1_cond $X=5.022 $Y=0.88
+ $X2=5.022 $Y2=0.515
r260 77 101 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.735 $Y=1.13
+ $X2=4.735 $Y2=1.005
r261 77 78 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=4.735 $Y=1.13
+ $X2=4.735 $Y2=1.3
r262 76 125 9.36528 $w=3.86e-07 $l=7.5e-08 $layer=POLY_cond $X=4.21 $Y=1.532
+ $X2=4.285 $Y2=1.532
r263 76 123 51.1969 $w=3.86e-07 $l=4.1e-07 $layer=POLY_cond $X=4.21 $Y=1.532
+ $X2=3.8 $Y2=1.532
r264 75 76 36.32 $w=1.7e-07 $l=6.8e-07 $layer=licon1_POLY $count=4 $X=4.21
+ $Y=1.465 $X2=4.21 $Y2=1.465
r265 72 114 9.36528 $w=3.86e-07 $l=7.5e-08 $layer=POLY_cond $X=1.83 $Y=1.532
+ $X2=1.905 $Y2=1.532
r266 72 112 46.8264 $w=3.86e-07 $l=3.75e-07 $layer=POLY_cond $X=1.83 $Y=1.532
+ $X2=1.455 $Y2=1.532
r267 71 75 83.1156 $w=3.28e-07 $l=2.38e-06 $layer=LI1_cond $X=1.83 $Y=1.465
+ $X2=4.21 $Y2=1.465
r268 71 72 36.32 $w=1.7e-07 $l=6.8e-07 $layer=licon1_POLY $count=4 $X=1.83
+ $Y=1.465 $X2=1.83 $Y2=1.465
r269 69 78 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.65 $Y=1.465
+ $X2=4.735 $Y2=1.3
r270 69 75 15.3659 $w=3.28e-07 $l=4.4e-07 $layer=LI1_cond $X=4.65 $Y=1.465
+ $X2=4.21 $Y2=1.465
r271 65 126 24.9932 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=4.3 $Y=1.3
+ $X2=4.3 $Y2=1.532
r272 65 67 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=4.3 $Y=1.3 $X2=4.3
+ $Y2=0.74
r273 62 125 24.9932 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=4.285 $Y=1.765
+ $X2=4.285 $Y2=1.532
r274 62 64 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=4.285 $Y=1.765
+ $X2=4.285 $Y2=2.4
r275 58 123 24.9932 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=3.8 $Y=1.3
+ $X2=3.8 $Y2=1.532
r276 58 60 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=3.8 $Y=1.3 $X2=3.8
+ $Y2=0.74
r277 55 122 24.9932 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=3.705 $Y=1.765
+ $X2=3.705 $Y2=1.532
r278 55 57 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.705 $Y=1.765
+ $X2=3.705 $Y2=2.4
r279 51 121 24.9932 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=3.3 $Y=1.3
+ $X2=3.3 $Y2=1.532
r280 51 53 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=3.3 $Y=1.3 $X2=3.3
+ $Y2=0.74
r281 48 120 24.9932 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=3.255 $Y=1.765
+ $X2=3.255 $Y2=1.532
r282 48 50 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.255 $Y=1.765
+ $X2=3.255 $Y2=2.4
r283 44 119 24.9932 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=2.87 $Y=1.3
+ $X2=2.87 $Y2=1.532
r284 44 46 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=2.87 $Y=1.3
+ $X2=2.87 $Y2=0.74
r285 41 118 24.9932 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=2.805 $Y=1.765
+ $X2=2.805 $Y2=1.532
r286 41 43 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.805 $Y=1.765
+ $X2=2.805 $Y2=2.4
r287 37 117 24.9932 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=2.37 $Y=1.3
+ $X2=2.37 $Y2=1.532
r288 37 39 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=2.37 $Y=1.3
+ $X2=2.37 $Y2=0.74
r289 34 116 24.9932 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=2.355 $Y=1.765
+ $X2=2.355 $Y2=1.532
r290 34 36 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.355 $Y=1.765
+ $X2=2.355 $Y2=2.4
r291 30 115 24.9932 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=1.94 $Y=1.3
+ $X2=1.94 $Y2=1.532
r292 30 32 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=1.94 $Y=1.3
+ $X2=1.94 $Y2=0.74
r293 27 114 24.9932 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=1.905 $Y=1.765
+ $X2=1.905 $Y2=1.532
r294 27 29 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.905 $Y=1.765
+ $X2=1.905 $Y2=2.4
r295 24 112 24.9932 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=1.455 $Y=1.765
+ $X2=1.455 $Y2=1.532
r296 24 26 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.455 $Y=1.765
+ $X2=1.455 $Y2=2.4
r297 20 111 24.9932 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=1.44 $Y=1.3
+ $X2=1.44 $Y2=1.532
r298 20 22 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=1.44 $Y=1.3
+ $X2=1.44 $Y2=0.74
r299 17 110 24.9932 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=1.005 $Y=1.765
+ $X2=1.005 $Y2=1.532
r300 17 19 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.005 $Y=1.765
+ $X2=1.005 $Y2=2.4
r301 13 109 24.9932 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=0.99 $Y=1.3
+ $X2=0.99 $Y2=1.532
r302 13 15 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=0.99 $Y=1.3
+ $X2=0.99 $Y2=0.74
r303 4 99 300 $w=1.7e-07 $l=6.30555e-07 $layer=licon1_PDIFF $count=2 $X=5.81
+ $Y=1.84 $X2=5.96 $Y2=2.4
r304 4 96 600 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=5.81
+ $Y=1.84 $X2=5.96 $Y2=1.985
r305 3 106 300 $w=1.7e-07 $l=5.34766e-07 $layer=licon1_PDIFF $count=2 $X=4.86
+ $Y=1.84 $X2=5.01 $Y2=2.305
r306 2 91 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=5.82
+ $Y=0.37 $X2=5.96 $Y2=0.515
r307 1 104 182 $w=1.7e-07 $l=6.63551e-07 $layer=licon1_NDIFF $count=1 $X=4.875
+ $Y=0.37 $X2=5.02 $Y2=0.965
r308 1 83 182 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=1 $X=4.875
+ $Y=0.37 $X2=5.02 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__BUFINV_8%A_27_368# 1 2 7 9 12 14 16 19 21 23 26 30
+ 34 36 37 38 41 42 45 46 47 49 52 54 64
c152 54 0 7.6204e-20 $X=5.475 $Y=1.485
c153 30 0 1.10108e-19 $X=0.28 $Y=2.815
c154 19 0 1.04254e-19 $X=5.245 $Y=0.74
c155 12 0 1.63832e-19 $X=4.8 $Y=0.74
c156 7 0 1.38632e-19 $X=4.785 $Y=1.765
r157 64 65 1.27177 $w=3.79e-07 $l=1e-08 $layer=POLY_cond $X=5.735 $Y=1.542
+ $X2=5.745 $Y2=1.542
r158 61 62 1.27177 $w=3.79e-07 $l=1e-08 $layer=POLY_cond $X=5.235 $Y=1.542
+ $X2=5.245 $Y2=1.542
r159 60 61 55.3219 $w=3.79e-07 $l=4.35e-07 $layer=POLY_cond $X=4.8 $Y=1.542
+ $X2=5.235 $Y2=1.542
r160 59 60 1.90765 $w=3.79e-07 $l=1.5e-08 $layer=POLY_cond $X=4.785 $Y=1.542
+ $X2=4.8 $Y2=1.542
r161 55 64 33.066 $w=3.79e-07 $l=2.6e-07 $layer=POLY_cond $X=5.475 $Y=1.542
+ $X2=5.735 $Y2=1.542
r162 55 62 29.2507 $w=3.79e-07 $l=2.3e-07 $layer=POLY_cond $X=5.475 $Y=1.542
+ $X2=5.245 $Y2=1.542
r163 54 55 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.475
+ $Y=1.485 $X2=5.475 $Y2=1.485
r164 49 51 7.33373 $w=3.28e-07 $l=2.1e-07 $layer=LI1_cond $X=0.28 $Y=2.115
+ $X2=0.28 $Y2=2.325
r165 46 54 7.77937 $w=6.13e-07 $l=4e-07 $layer=LI1_cond $X=5.297 $Y=1.885
+ $X2=5.297 $Y2=1.485
r166 46 47 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=4.99 $Y=1.885
+ $X2=4.565 $Y2=1.885
r167 44 47 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.48 $Y=1.97
+ $X2=4.565 $Y2=1.885
r168 44 45 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=4.48 $Y=1.97
+ $X2=4.48 $Y2=2.24
r169 43 52 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.89 $Y=2.325
+ $X2=0.805 $Y2=2.325
r170 42 45 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.395 $Y=2.325
+ $X2=4.48 $Y2=2.24
r171 42 43 228.668 $w=1.68e-07 $l=3.505e-06 $layer=LI1_cond $X=4.395 $Y=2.325
+ $X2=0.89 $Y2=2.325
r172 41 52 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.805 $Y=2.24
+ $X2=0.805 $Y2=2.325
r173 40 41 69.1551 $w=1.68e-07 $l=1.06e-06 $layer=LI1_cond $X=0.805 $Y=1.18
+ $X2=0.805 $Y2=2.24
r174 39 51 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.445 $Y=2.325
+ $X2=0.28 $Y2=2.325
r175 38 52 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.72 $Y=2.325
+ $X2=0.805 $Y2=2.325
r176 38 39 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=0.72 $Y=2.325
+ $X2=0.445 $Y2=2.325
r177 36 40 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.72 $Y=1.095
+ $X2=0.805 $Y2=1.18
r178 36 37 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=0.72 $Y=1.095
+ $X2=0.38 $Y2=1.095
r179 32 37 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.255 $Y=1.01
+ $X2=0.38 $Y2=1.095
r180 32 34 22.8184 $w=2.48e-07 $l=4.95e-07 $layer=LI1_cond $X=0.255 $Y=1.01
+ $X2=0.255 $Y2=0.515
r181 28 51 2.96841 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=0.28 $Y=2.41
+ $X2=0.28 $Y2=2.325
r182 28 30 14.1436 $w=3.28e-07 $l=4.05e-07 $layer=LI1_cond $X=0.28 $Y=2.41
+ $X2=0.28 $Y2=2.815
r183 24 65 24.5487 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=5.745 $Y=1.32
+ $X2=5.745 $Y2=1.542
r184 24 26 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=5.745 $Y=1.32
+ $X2=5.745 $Y2=0.74
r185 21 64 24.5487 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=5.735 $Y=1.765
+ $X2=5.735 $Y2=1.542
r186 21 23 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=5.735 $Y=1.765
+ $X2=5.735 $Y2=2.4
r187 17 62 24.5487 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=5.245 $Y=1.32
+ $X2=5.245 $Y2=1.542
r188 17 19 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=5.245 $Y=1.32
+ $X2=5.245 $Y2=0.74
r189 14 61 24.5487 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=5.235 $Y=1.765
+ $X2=5.235 $Y2=1.542
r190 14 16 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=5.235 $Y=1.765
+ $X2=5.235 $Y2=2.4
r191 10 60 24.5487 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=4.8 $Y=1.32
+ $X2=4.8 $Y2=1.542
r192 10 12 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=4.8 $Y=1.32 $X2=4.8
+ $Y2=0.74
r193 7 59 24.5487 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=4.785 $Y=1.765
+ $X2=4.785 $Y2=1.542
r194 7 9 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=4.785 $Y=1.765
+ $X2=4.785 $Y2=2.4
r195 2 49 400 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.115
r196 2 30 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.815
r197 1 34 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.15
+ $Y=0.37 $X2=0.295 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__BUFINV_8%VPWR 1 2 3 4 5 6 21 25 29 33 37 41 44 45 46
+ 48 53 58 67 71 78 79 82 85 88 91 94
r99 94 95 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r100 91 92 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r101 88 89 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r102 85 86 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r103 82 83 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r104 79 95 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=3.33 $X2=5.52
+ $Y2=3.33
r105 78 79 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r106 76 94 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.675 $Y=3.33
+ $X2=5.51 $Y2=3.33
r107 76 78 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=5.675 $Y=3.33
+ $X2=6 $Y2=3.33
r108 75 95 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=5.52 $Y2=3.33
r109 75 92 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=4.56 $Y2=3.33
r110 74 75 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r111 72 91 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.675 $Y=3.33
+ $X2=4.51 $Y2=3.33
r112 72 74 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=4.675 $Y=3.33
+ $X2=5.04 $Y2=3.33
r113 71 94 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.345 $Y=3.33
+ $X2=5.51 $Y2=3.33
r114 71 74 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=5.345 $Y=3.33
+ $X2=5.04 $Y2=3.33
r115 70 92 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=4.56 $Y2=3.33
r116 69 70 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r117 67 91 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.345 $Y=3.33
+ $X2=4.51 $Y2=3.33
r118 67 69 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=4.345 $Y=3.33
+ $X2=4.08 $Y2=3.33
r119 63 88 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.745 $Y=3.33
+ $X2=2.58 $Y2=3.33
r120 63 65 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=2.745 $Y=3.33
+ $X2=3.12 $Y2=3.33
r121 62 89 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r122 62 86 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.68 $Y2=3.33
r123 61 62 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r124 59 85 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.845 $Y=3.33
+ $X2=1.68 $Y2=3.33
r125 59 61 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=1.845 $Y=3.33
+ $X2=2.16 $Y2=3.33
r126 58 88 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.415 $Y=3.33
+ $X2=2.58 $Y2=3.33
r127 58 61 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=2.415 $Y=3.33
+ $X2=2.16 $Y2=3.33
r128 57 86 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=1.68 $Y2=3.33
r129 57 83 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r130 56 57 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r131 54 82 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.945 $Y=3.33
+ $X2=0.78 $Y2=3.33
r132 54 56 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.945 $Y=3.33
+ $X2=1.2 $Y2=3.33
r133 53 85 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.515 $Y=3.33
+ $X2=1.68 $Y2=3.33
r134 53 56 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=1.515 $Y=3.33
+ $X2=1.2 $Y2=3.33
r135 51 83 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r136 50 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r137 48 82 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.615 $Y=3.33
+ $X2=0.78 $Y2=3.33
r138 48 50 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=0.615 $Y=3.33
+ $X2=0.24 $Y2=3.33
r139 46 70 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=4.08 $Y2=3.33
r140 46 89 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=2.64 $Y2=3.33
r141 46 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r142 44 65 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=3.315 $Y=3.33
+ $X2=3.12 $Y2=3.33
r143 44 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.315 $Y=3.33
+ $X2=3.48 $Y2=3.33
r144 43 69 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=3.645 $Y=3.33
+ $X2=4.08 $Y2=3.33
r145 43 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.645 $Y=3.33
+ $X2=3.48 $Y2=3.33
r146 39 94 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.51 $Y=3.245
+ $X2=5.51 $Y2=3.33
r147 39 41 20.9535 $w=3.28e-07 $l=6e-07 $layer=LI1_cond $X=5.51 $Y=3.245
+ $X2=5.51 $Y2=2.645
r148 35 91 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.51 $Y=3.245
+ $X2=4.51 $Y2=3.33
r149 35 37 17.4613 $w=3.28e-07 $l=5e-07 $layer=LI1_cond $X=4.51 $Y=3.245
+ $X2=4.51 $Y2=2.745
r150 31 45 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.48 $Y=3.245
+ $X2=3.48 $Y2=3.33
r151 31 33 17.4613 $w=3.28e-07 $l=5e-07 $layer=LI1_cond $X=3.48 $Y=3.245
+ $X2=3.48 $Y2=2.745
r152 27 88 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.58 $Y=3.245
+ $X2=2.58 $Y2=3.33
r153 27 29 17.4613 $w=3.28e-07 $l=5e-07 $layer=LI1_cond $X=2.58 $Y=3.245
+ $X2=2.58 $Y2=2.745
r154 23 85 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.68 $Y=3.245
+ $X2=1.68 $Y2=3.33
r155 23 25 17.4613 $w=3.28e-07 $l=5e-07 $layer=LI1_cond $X=1.68 $Y=3.245
+ $X2=1.68 $Y2=2.745
r156 19 82 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.78 $Y=3.245
+ $X2=0.78 $Y2=3.33
r157 19 21 17.4613 $w=3.28e-07 $l=5e-07 $layer=LI1_cond $X=0.78 $Y=3.245
+ $X2=0.78 $Y2=2.745
r158 6 41 600 $w=1.7e-07 $l=8.99458e-07 $layer=licon1_PDIFF $count=1 $X=5.31
+ $Y=1.84 $X2=5.51 $Y2=2.645
r159 5 37 600 $w=1.7e-07 $l=9.77126e-07 $layer=licon1_PDIFF $count=1 $X=4.36
+ $Y=1.84 $X2=4.51 $Y2=2.745
r160 4 33 600 $w=1.7e-07 $l=9.77126e-07 $layer=licon1_PDIFF $count=1 $X=3.33
+ $Y=1.84 $X2=3.48 $Y2=2.745
r161 3 29 600 $w=1.7e-07 $l=9.77126e-07 $layer=licon1_PDIFF $count=1 $X=2.43
+ $Y=1.84 $X2=2.58 $Y2=2.745
r162 2 25 600 $w=1.7e-07 $l=9.77126e-07 $layer=licon1_PDIFF $count=1 $X=1.53
+ $Y=1.84 $X2=1.68 $Y2=2.745
r163 1 21 600 $w=1.7e-07 $l=1.00001e-06 $layer=licon1_PDIFF $count=1 $X=0.58
+ $Y=1.84 $X2=0.78 $Y2=2.745
.ends

.subckt PM_SKY130_FD_SC_HS__BUFINV_8%Y 1 2 3 4 5 6 7 8 25 33 37 39 43 45 49 51
+ 55 56 57 58 59 60
c102 59 0 2.3255e-19 $X=1.2 $Y=1.295
c103 45 0 1.63832e-19 $X=3.92 $Y=1.045
c104 33 0 1.38632e-19 $X=3.995 $Y=1.985
r105 59 60 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.225 $Y=1.295
+ $X2=1.225 $Y2=1.665
r106 59 72 5.76222 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=1.225 $Y=1.295
+ $X2=1.225 $Y2=1.13
r107 58 66 4.07664 $w=3.3e-07 $l=1.25e-07 $layer=LI1_cond $X=1.225 $Y=1.005
+ $X2=1.225 $Y2=0.88
r108 58 72 4.07664 $w=3.3e-07 $l=1.25e-07 $layer=LI1_cond $X=1.225 $Y=1.005
+ $X2=1.225 $Y2=1.13
r109 58 66 0.69845 $w=3.28e-07 $l=2e-08 $layer=LI1_cond $X=1.225 $Y=0.86
+ $X2=1.225 $Y2=0.88
r110 57 58 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=1.225 $Y=0.515
+ $X2=1.225 $Y2=0.86
r111 51 60 4.71454 $w=3.28e-07 $l=1.35e-07 $layer=LI1_cond $X=1.225 $Y=1.8
+ $X2=1.225 $Y2=1.665
r112 51 53 3.10749 $w=3.3e-07 $l=1.35e-07 $layer=LI1_cond $X=1.225 $Y=1.8
+ $X2=1.225 $Y2=1.935
r113 47 49 15.5405 $w=3.28e-07 $l=4.45e-07 $layer=LI1_cond $X=4.085 $Y=0.96
+ $X2=4.085 $Y2=0.515
r114 46 56 7.38875 $w=2.1e-07 $l=1.83916e-07 $layer=LI1_cond $X=3.25 $Y=1.045
+ $X2=3.085 $Y2=1.005
r115 45 47 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.92 $Y=1.045
+ $X2=4.085 $Y2=0.96
r116 45 46 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.92 $Y=1.045
+ $X2=3.25 $Y2=1.045
r117 41 56 0.221902 $w=3.3e-07 $l=1.25e-07 $layer=LI1_cond $X=3.085 $Y=0.88
+ $X2=3.085 $Y2=1.005
r118 41 43 12.7467 $w=3.28e-07 $l=3.65e-07 $layer=LI1_cond $X=3.085 $Y=0.88
+ $X2=3.085 $Y2=0.515
r119 40 55 4.08801 $w=2.5e-07 $l=9.5e-08 $layer=LI1_cond $X=2.25 $Y=1.005
+ $X2=2.155 $Y2=1.005
r120 39 56 7.38875 $w=2.1e-07 $l=1.65e-07 $layer=LI1_cond $X=2.92 $Y=1.005
+ $X2=3.085 $Y2=1.005
r121 39 40 30.8855 $w=2.48e-07 $l=6.7e-07 $layer=LI1_cond $X=2.92 $Y=1.005
+ $X2=2.25 $Y2=1.005
r122 35 55 2.34704 $w=1.9e-07 $l=1.25e-07 $layer=LI1_cond $X=2.155 $Y=0.88
+ $X2=2.155 $Y2=1.005
r123 35 37 21.3062 $w=1.88e-07 $l=3.65e-07 $layer=LI1_cond $X=2.155 $Y=0.88
+ $X2=2.155 $Y2=0.515
r124 31 33 41.1892 $w=2.68e-07 $l=9.65e-07 $layer=LI1_cond $X=3.03 $Y=1.935
+ $X2=3.995 $Y2=1.935
r125 29 31 38.4148 $w=2.68e-07 $l=9e-07 $layer=LI1_cond $X=2.13 $Y=1.935
+ $X2=3.03 $Y2=1.935
r126 27 53 3.79804 $w=2.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.39 $Y=1.935
+ $X2=1.225 $Y2=1.935
r127 27 29 31.5855 $w=2.68e-07 $l=7.4e-07 $layer=LI1_cond $X=1.39 $Y=1.935
+ $X2=2.13 $Y2=1.935
r128 26 58 2.3589 $w=2.5e-07 $l=1.65e-07 $layer=LI1_cond $X=1.39 $Y=1.005
+ $X2=1.225 $Y2=1.005
r129 25 55 4.08801 $w=2.5e-07 $l=9.5e-08 $layer=LI1_cond $X=2.06 $Y=1.005
+ $X2=2.155 $Y2=1.005
r130 25 26 30.8855 $w=2.48e-07 $l=6.7e-07 $layer=LI1_cond $X=2.06 $Y=1.005
+ $X2=1.39 $Y2=1.005
r131 8 33 600 $w=1.7e-07 $l=2.78209e-07 $layer=licon1_PDIFF $count=1 $X=3.78
+ $Y=1.84 $X2=3.995 $Y2=1.985
r132 7 31 600 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=2.88
+ $Y=1.84 $X2=3.03 $Y2=1.985
r133 6 29 600 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=1.98
+ $Y=1.84 $X2=2.13 $Y2=1.985
r134 5 53 600 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=1.08
+ $Y=1.84 $X2=1.23 $Y2=1.985
r135 4 49 91 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=2 $X=3.875
+ $Y=0.37 $X2=4.085 $Y2=0.515
r136 3 43 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.945
+ $Y=0.37 $X2=3.085 $Y2=0.515
r137 2 55 182 $w=1.7e-07 $l=6.61306e-07 $layer=licon1_NDIFF $count=1 $X=2.015
+ $Y=0.37 $X2=2.155 $Y2=0.965
r138 2 37 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=2.015
+ $Y=0.37 $X2=2.155 $Y2=0.515
r139 1 57 91 $w=1.7e-07 $l=2.20907e-07 $layer=licon1_NDIFF $count=2 $X=1.065
+ $Y=0.37 $X2=1.225 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__BUFINV_8%VGND 1 2 3 4 5 6 21 25 29 33 37 41 43 45 50
+ 55 60 65 70 77 78 81 84 87 90 93 96
r100 96 97 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r101 93 94 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r102 90 91 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r103 87 88 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r104 84 85 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r105 81 82 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r106 78 97 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=0 $X2=5.52
+ $Y2=0
r107 77 78 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=0 $X2=6 $Y2=0
r108 75 96 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.625 $Y=0 $X2=5.46
+ $Y2=0
r109 75 77 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=5.625 $Y=0 $X2=6
+ $Y2=0
r110 74 97 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=5.52
+ $Y2=0
r111 74 94 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=4.56
+ $Y2=0
r112 73 74 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r113 71 93 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.75 $Y=0 $X2=4.585
+ $Y2=0
r114 71 73 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=4.75 $Y=0 $X2=5.04
+ $Y2=0
r115 70 96 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.295 $Y=0 $X2=5.46
+ $Y2=0
r116 70 73 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=5.295 $Y=0
+ $X2=5.04 $Y2=0
r117 69 94 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=4.56
+ $Y2=0
r118 69 91 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=3.6
+ $Y2=0
r119 68 69 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r120 66 90 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.75 $Y=0 $X2=3.585
+ $Y2=0
r121 66 68 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=3.75 $Y=0 $X2=4.08
+ $Y2=0
r122 65 93 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.42 $Y=0 $X2=4.585
+ $Y2=0
r123 65 68 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=4.42 $Y=0 $X2=4.08
+ $Y2=0
r124 61 87 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.75 $Y=0 $X2=2.585
+ $Y2=0
r125 61 63 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=2.75 $Y=0 $X2=3.12
+ $Y2=0
r126 60 90 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.42 $Y=0 $X2=3.585
+ $Y2=0
r127 60 63 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=3.42 $Y=0 $X2=3.12
+ $Y2=0
r128 59 88 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r129 59 85 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.68
+ $Y2=0
r130 58 59 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r131 56 84 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.89 $Y=0 $X2=1.725
+ $Y2=0
r132 56 58 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=1.89 $Y=0 $X2=2.16
+ $Y2=0
r133 55 87 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.42 $Y=0 $X2=2.585
+ $Y2=0
r134 55 58 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=2.42 $Y=0 $X2=2.16
+ $Y2=0
r135 54 85 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=1.68
+ $Y2=0
r136 54 82 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r137 53 54 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r138 51 81 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.89 $Y=0 $X2=0.725
+ $Y2=0
r139 51 53 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=0.89 $Y=0 $X2=1.2
+ $Y2=0
r140 50 84 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.56 $Y=0 $X2=1.725
+ $Y2=0
r141 50 53 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=1.56 $Y=0 $X2=1.2
+ $Y2=0
r142 48 82 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r143 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r144 45 81 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.56 $Y=0 $X2=0.725
+ $Y2=0
r145 45 47 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=0.56 $Y=0 $X2=0.24
+ $Y2=0
r146 43 91 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=3.6
+ $Y2=0
r147 43 88 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=2.64
+ $Y2=0
r148 43 63 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r149 39 96 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.46 $Y=0.085
+ $X2=5.46 $Y2=0
r150 39 41 16.0644 $w=3.28e-07 $l=4.6e-07 $layer=LI1_cond $X=5.46 $Y=0.085
+ $X2=5.46 $Y2=0.545
r151 35 93 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.585 $Y=0.085
+ $X2=4.585 $Y2=0
r152 35 37 16.0644 $w=3.28e-07 $l=4.6e-07 $layer=LI1_cond $X=4.585 $Y=0.085
+ $X2=4.585 $Y2=0.545
r153 31 90 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.585 $Y=0.085
+ $X2=3.585 $Y2=0
r154 31 33 18.8582 $w=3.28e-07 $l=5.4e-07 $layer=LI1_cond $X=3.585 $Y=0.085
+ $X2=3.585 $Y2=0.625
r155 27 87 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.585 $Y=0.085
+ $X2=2.585 $Y2=0
r156 27 29 16.0644 $w=3.28e-07 $l=4.6e-07 $layer=LI1_cond $X=2.585 $Y=0.085
+ $X2=2.585 $Y2=0.545
r157 23 84 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.725 $Y=0.085
+ $X2=1.725 $Y2=0
r158 23 25 16.9374 $w=3.28e-07 $l=4.85e-07 $layer=LI1_cond $X=1.725 $Y=0.085
+ $X2=1.725 $Y2=0.57
r159 19 81 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.725 $Y=0.085
+ $X2=0.725 $Y2=0
r160 19 21 17.8105 $w=3.28e-07 $l=5.1e-07 $layer=LI1_cond $X=0.725 $Y=0.085
+ $X2=0.725 $Y2=0.595
r161 6 41 182 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_NDIFF $count=1 $X=5.32
+ $Y=0.37 $X2=5.46 $Y2=0.545
r162 5 37 182 $w=1.7e-07 $l=2.84341e-07 $layer=licon1_NDIFF $count=1 $X=4.375
+ $Y=0.37 $X2=4.585 $Y2=0.545
r163 4 33 182 $w=1.7e-07 $l=3.44347e-07 $layer=licon1_NDIFF $count=1 $X=3.375
+ $Y=0.37 $X2=3.585 $Y2=0.625
r164 3 29 182 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_NDIFF $count=1 $X=2.445
+ $Y=0.37 $X2=2.585 $Y2=0.545
r165 2 25 182 $w=1.7e-07 $l=2.93428e-07 $layer=licon1_NDIFF $count=1 $X=1.515
+ $Y=0.37 $X2=1.725 $Y2=0.57
r166 1 21 182 $w=1.7e-07 $l=2.86575e-07 $layer=licon1_NDIFF $count=1 $X=0.585
+ $Y=0.37 $X2=0.725 $Y2=0.595
.ends

