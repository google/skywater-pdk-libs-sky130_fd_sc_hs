* File: sky130_fd_sc_hs__and4b_1.pex.spice
* Created: Thu Aug 27 20:33:24 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HS__AND4B_1%A_N 3 5 7 10 11 14 15
r38 14 15 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.43
+ $Y=1.355 $X2=0.43 $Y2=1.355
r39 11 15 3.39186 $w=6.68e-07 $l=1.9e-07 $layer=LI1_cond $X=0.24 $Y=1.525
+ $X2=0.43 $Y2=1.525
r40 10 14 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=0.43 $Y=1.695
+ $X2=0.43 $Y2=1.355
r41 9 14 42.4377 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.43 $Y=1.19
+ $X2=0.43 $Y2=1.355
r42 5 10 67.48 $w=2.5e-07 $l=3.85681e-07 $layer=POLY_cond $X=0.505 $Y=2.045
+ $X2=0.43 $Y2=1.695
r43 5 7 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=0.505 $Y=2.045
+ $X2=0.505 $Y2=2.54
r44 3 9 279.457 $w=1.5e-07 $l=5.45e-07 $layer=POLY_cond $X=0.495 $Y=0.645
+ $X2=0.495 $Y2=1.19
.ends

.subckt PM_SKY130_FD_SC_HS__AND4B_1%A_27_74# 1 2 7 9 11 12 13 14 16 19 23 25 26
+ 27 28 30 32 36
r81 36 37 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.09
+ $Y=1.715 $X2=1.09 $Y2=1.715
r82 33 36 8.03218 $w=3.28e-07 $l=2.3e-07 $layer=LI1_cond $X=0.86 $Y=1.715
+ $X2=1.09 $Y2=1.715
r83 31 33 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.86 $Y=1.88
+ $X2=0.86 $Y2=1.715
r84 31 32 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=0.86 $Y=1.88 $X2=0.86
+ $Y2=2.03
r85 30 33 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.86 $Y=1.55
+ $X2=0.86 $Y2=1.715
r86 29 30 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=0.86 $Y=1.02
+ $X2=0.86 $Y2=1.55
r87 27 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.775 $Y=2.115
+ $X2=0.86 $Y2=2.03
r88 27 28 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=0.775 $Y=2.115
+ $X2=0.445 $Y2=2.115
r89 25 29 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.775 $Y=0.935
+ $X2=0.86 $Y2=1.02
r90 25 26 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.775 $Y=0.935
+ $X2=0.405 $Y2=0.935
r91 21 28 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.28 $Y=2.2
+ $X2=0.445 $Y2=2.115
r92 21 23 2.26996 $w=3.28e-07 $l=6.5e-08 $layer=LI1_cond $X=0.28 $Y=2.2 $X2=0.28
+ $Y2=2.265
r93 17 26 7.43784 $w=1.7e-07 $l=1.8262e-07 $layer=LI1_cond $X=0.26 $Y=0.85
+ $X2=0.405 $Y2=0.935
r94 17 19 8.14658 $w=2.88e-07 $l=2.05e-07 $layer=LI1_cond $X=0.26 $Y=0.85
+ $X2=0.26 $Y2=0.645
r95 14 16 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=1.69 $Y=0.545
+ $X2=1.69 $Y2=0.94
r96 12 14 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.615 $Y=0.47
+ $X2=1.69 $Y2=0.545
r97 12 13 184.596 $w=1.5e-07 $l=3.6e-07 $layer=POLY_cond $X=1.615 $Y=0.47
+ $X2=1.255 $Y2=0.47
r98 11 37 38.7299 $w=2.8e-07 $l=2.05122e-07 $layer=POLY_cond $X=1.18 $Y=1.55
+ $X2=1.09 $Y2=1.715
r99 10 13 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.18 $Y=0.545
+ $X2=1.255 $Y2=0.47
r100 10 11 515.33 $w=1.5e-07 $l=1.005e-06 $layer=POLY_cond $X=1.18 $Y=0.545
+ $X2=1.18 $Y2=1.55
r101 7 37 67.1335 $w=2.8e-07 $l=3.47059e-07 $layer=POLY_cond $X=1.055 $Y=2.045
+ $X2=1.09 $Y2=1.715
r102 7 9 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=1.055 $Y=2.045
+ $X2=1.055 $Y2=2.54
r103 2 23 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=2.12 $X2=0.28 $Y2=2.265
r104 1 19 182 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.645
.ends

.subckt PM_SKY130_FD_SC_HS__AND4B_1%B 1 3 6 8 9 10 11
c37 11 0 7.31803e-20 $X=2.16 $Y=1.665
c38 8 0 1.33203e-19 $X=1.675 $Y=1.795
r39 15 16 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.075
+ $Y=1.795 $X2=2.075 $Y2=1.795
r40 11 16 2.38921 $w=4.08e-07 $l=8.5e-08 $layer=LI1_cond $X=2.16 $Y=1.755
+ $X2=2.075 $Y2=1.755
r41 10 16 11.1028 $w=4.08e-07 $l=3.95e-07 $layer=LI1_cond $X=1.68 $Y=1.755
+ $X2=2.075 $Y2=1.755
r42 9 15 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=2.09 $Y=1.795
+ $X2=2.075 $Y2=1.795
r43 8 15 69.9445 $w=3.3e-07 $l=4e-07 $layer=POLY_cond $X=1.675 $Y=1.795
+ $X2=2.075 $Y2=1.795
r44 4 9 32.1775 $w=3.3e-07 $l=1.98997e-07 $layer=POLY_cond $X=2.165 $Y=1.63
+ $X2=2.09 $Y2=1.795
r45 4 6 315.351 $w=1.5e-07 $l=6.15e-07 $layer=POLY_cond $X=2.165 $Y=1.63
+ $X2=2.165 $Y2=1.015
r46 1 8 32.1775 $w=3.3e-07 $l=2.91548e-07 $layer=POLY_cond $X=1.585 $Y=2.045
+ $X2=1.675 $Y2=1.795
r47 1 3 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=1.585 $Y=2.045
+ $X2=1.585 $Y2=2.54
.ends

.subckt PM_SKY130_FD_SC_HS__AND4B_1%C 4 6 7 9 11 12 13 17 18
c47 11 0 7.31803e-20 $X=2.612 $Y=1.56
r48 17 20 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.645 $Y=0.42
+ $X2=2.645 $Y2=0.585
r49 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.645
+ $Y=0.42 $X2=2.645 $Y2=0.42
r50 13 18 0.138849 $w=4.13e-07 $l=5e-09 $layer=LI1_cond $X=2.64 $Y=0.462
+ $X2=2.645 $Y2=0.462
r51 12 13 13.3295 $w=4.13e-07 $l=4.8e-07 $layer=LI1_cond $X=2.16 $Y=0.462
+ $X2=2.64 $Y2=0.462
r52 10 11 60.4563 $w=1.8e-07 $l=1.5e-07 $layer=POLY_cond $X=2.612 $Y=1.41
+ $X2=2.612 $Y2=1.56
r53 7 9 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=2.655 $Y=2.045
+ $X2=2.655 $Y2=2.54
r54 6 7 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=2.655 $Y=1.955 $X2=2.655
+ $Y2=2.045
r55 6 11 153.54 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=2.655 $Y=1.955
+ $X2=2.655 $Y2=1.56
r56 4 10 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=2.555 $Y=1.015
+ $X2=2.555 $Y2=1.41
r57 4 20 220.489 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=2.555 $Y=1.015
+ $X2=2.555 $Y2=0.585
.ends

.subckt PM_SKY130_FD_SC_HS__AND4B_1%D 1 3 6 8
r37 8 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.15
+ $Y=1.715 $X2=3.15 $Y2=1.715
r38 4 11 38.6899 $w=2.83e-07 $l=2.06325e-07 $layer=POLY_cond $X=3.245 $Y=1.55
+ $X2=3.152 $Y2=1.715
r39 4 6 323.043 $w=1.5e-07 $l=6.3e-07 $layer=POLY_cond $X=3.245 $Y=1.55
+ $X2=3.245 $Y2=0.92
r40 1 11 66.7923 $w=2.83e-07 $l=3.31497e-07 $layer=POLY_cond $X=3.155 $Y=2.045
+ $X2=3.152 $Y2=1.715
r41 1 3 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=3.155 $Y=2.045
+ $X2=3.155 $Y2=2.54
.ends

.subckt PM_SKY130_FD_SC_HS__AND4B_1%A_226_424# 1 2 3 10 12 13 15 18 22 23 25 26
+ 30 35 36 38 40
c98 22 0 1.33203e-19 $X=2.595 $Y=1.295
r99 44 45 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.725
+ $Y=1.515 $X2=3.725 $Y2=1.515
r100 37 40 11.5244 $w=2.48e-07 $l=2.5e-07 $layer=LI1_cond $X=2.68 $Y=2.225
+ $X2=2.93 $Y2=2.225
r101 37 38 4.11343 $w=2.48e-07 $l=8.5e-08 $layer=LI1_cond $X=2.68 $Y=2.225
+ $X2=2.595 $Y2=2.225
r102 35 38 59.4556 $w=2.18e-07 $l=1.135e-06 $layer=LI1_cond $X=1.46 $Y=2.24
+ $X2=2.595 $Y2=2.24
r103 33 35 7.04571 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=1.295 $Y=2.295
+ $X2=1.46 $Y2=2.295
r104 30 40 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=2.93 $Y=2.815
+ $X2=2.93 $Y2=2.35
r105 27 36 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.765 $Y=1.295
+ $X2=2.68 $Y2=1.295
r106 26 44 8.97659 $w=2.99e-07 $l=2.95533e-07 $layer=LI1_cond $X=3.535 $Y=1.295
+ $X2=3.712 $Y2=1.515
r107 26 27 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=3.535 $Y=1.295
+ $X2=2.765 $Y2=1.295
r108 25 37 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.68 $Y=2.1
+ $X2=2.68 $Y2=2.225
r109 24 36 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.68 $Y=1.38
+ $X2=2.68 $Y2=1.295
r110 24 25 46.9733 $w=1.68e-07 $l=7.2e-07 $layer=LI1_cond $X=2.68 $Y=1.38
+ $X2=2.68 $Y2=2.1
r111 22 36 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.595 $Y=1.295
+ $X2=2.68 $Y2=1.295
r112 22 23 62.3048 $w=1.68e-07 $l=9.55e-07 $layer=LI1_cond $X=2.595 $Y=1.295
+ $X2=1.64 $Y2=1.295
r113 16 23 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.475 $Y=1.21
+ $X2=1.64 $Y2=1.295
r114 16 18 15.5405 $w=3.28e-07 $l=4.45e-07 $layer=LI1_cond $X=1.475 $Y=1.21
+ $X2=1.475 $Y2=0.765
r115 13 45 38.532 $w=3.11e-07 $l=2.06325e-07 $layer=POLY_cond $X=3.825 $Y=1.35
+ $X2=3.732 $Y2=1.515
r116 13 15 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=3.825 $Y=1.35
+ $X2=3.825 $Y2=0.87
r117 10 45 51.7056 $w=3.11e-07 $l=2.88531e-07 $layer=POLY_cond $X=3.815 $Y=1.765
+ $X2=3.732 $Y2=1.515
r118 10 12 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.815 $Y=1.765
+ $X2=3.815 $Y2=2.4
r119 3 40 600 $w=1.7e-07 $l=2.62678e-07 $layer=licon1_PDIFF $count=1 $X=2.73
+ $Y=2.12 $X2=2.93 $Y2=2.265
r120 3 30 600 $w=1.7e-07 $l=7.88686e-07 $layer=licon1_PDIFF $count=1 $X=2.73
+ $Y=2.12 $X2=2.93 $Y2=2.815
r121 2 33 600 $w=1.7e-07 $l=2.43926e-07 $layer=licon1_PDIFF $count=1 $X=1.13
+ $Y=2.12 $X2=1.295 $Y2=2.295
r122 1 18 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=1.33
+ $Y=0.62 $X2=1.475 $Y2=0.765
.ends

.subckt PM_SKY130_FD_SC_HS__AND4B_1%VPWR 1 2 3 12 18 21 22 23 25 35 36 39 44 50
r47 49 50 12.1537 $w=8.78e-07 $l=1.65e-07 $layer=LI1_cond $X=2.43 $Y=2.975
+ $X2=2.595 $Y2=2.975
r48 46 49 3.74318 $w=8.78e-07 $l=2.7e-07 $layer=LI1_cond $X=2.16 $Y=2.975
+ $X2=2.43 $Y2=2.975
r49 42 46 6.65455 $w=8.78e-07 $l=4.8e-07 $layer=LI1_cond $X=1.68 $Y=2.975
+ $X2=2.16 $Y2=2.975
r50 42 44 10.3515 $w=8.78e-07 $l=3.5e-08 $layer=LI1_cond $X=1.68 $Y=2.975
+ $X2=1.645 $Y2=2.975
r51 42 43 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r52 40 43 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.68 $Y2=3.33
r53 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r54 35 36 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r55 33 36 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=4.08 $Y2=3.33
r56 32 50 34.2513 $w=1.68e-07 $l=5.25e-07 $layer=LI1_cond $X=3.12 $Y=3.33
+ $X2=2.595 $Y2=3.33
r57 32 33 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r58 28 40 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r59 27 28 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r60 25 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.615 $Y=3.33
+ $X2=0.78 $Y2=3.33
r61 25 27 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=0.615 $Y=3.33
+ $X2=0.24 $Y2=3.33
r62 23 33 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=3.12 $Y2=3.33
r63 23 43 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.68 $Y2=3.33
r64 23 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r65 21 32 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=3.335 $Y=3.33
+ $X2=3.12 $Y2=3.33
r66 21 22 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.335 $Y=3.33
+ $X2=3.5 $Y2=3.33
r67 20 35 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=3.665 $Y=3.33
+ $X2=4.08 $Y2=3.33
r68 20 22 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.665 $Y=3.33
+ $X2=3.5 $Y2=3.33
r69 16 22 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.5 $Y=3.245 $X2=3.5
+ $Y2=3.33
r70 16 18 34.2241 $w=3.28e-07 $l=9.8e-07 $layer=LI1_cond $X=3.5 $Y=3.245 $X2=3.5
+ $Y2=2.265
r71 15 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.945 $Y=3.33
+ $X2=0.78 $Y2=3.33
r72 15 44 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=0.945 $Y=3.33
+ $X2=1.645 $Y2=3.33
r73 10 39 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.78 $Y=3.245
+ $X2=0.78 $Y2=3.33
r74 10 12 27.5888 $w=3.28e-07 $l=7.9e-07 $layer=LI1_cond $X=0.78 $Y=3.245
+ $X2=0.78 $Y2=2.455
r75 3 18 300 $w=1.7e-07 $l=3.34739e-07 $layer=licon1_PDIFF $count=2 $X=3.23
+ $Y=2.12 $X2=3.5 $Y2=2.265
r76 2 49 300 $w=1.7e-07 $l=1.01388e-06 $layer=licon1_PDIFF $count=2 $X=1.66
+ $Y=2.12 $X2=2.43 $Y2=2.685
r77 1 12 300 $w=1.7e-07 $l=4.2335e-07 $layer=licon1_PDIFF $count=2 $X=0.58
+ $Y=2.12 $X2=0.78 $Y2=2.455
.ends

.subckt PM_SKY130_FD_SC_HS__AND4B_1%X 1 2 9 13 14 15 16 23 32
r25 21 23 0.259705 $w=3.53e-07 $l=8e-09 $layer=LI1_cond $X=4.052 $Y=2.027
+ $X2=4.052 $Y2=2.035
r26 15 16 12.0114 $w=3.53e-07 $l=3.7e-07 $layer=LI1_cond $X=4.052 $Y=2.405
+ $X2=4.052 $Y2=2.775
r27 14 21 1.26606 $w=3.53e-07 $l=3.9e-08 $layer=LI1_cond $X=4.052 $Y=1.988
+ $X2=4.052 $Y2=2.027
r28 14 32 7.62255 $w=3.53e-07 $l=1.38e-07 $layer=LI1_cond $X=4.052 $Y=1.988
+ $X2=4.052 $Y2=1.85
r29 14 15 10.7778 $w=3.53e-07 $l=3.32e-07 $layer=LI1_cond $X=4.052 $Y=2.073
+ $X2=4.052 $Y2=2.405
r30 14 23 1.2336 $w=3.53e-07 $l=3.8e-08 $layer=LI1_cond $X=4.052 $Y=2.073
+ $X2=4.052 $Y2=2.035
r31 13 32 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.145 $Y=1.18
+ $X2=4.145 $Y2=1.85
r32 7 13 8.88861 $w=3.53e-07 $l=1.77e-07 $layer=LI1_cond $X=4.052 $Y=1.003
+ $X2=4.052 $Y2=1.18
r33 7 9 11.6218 $w=3.53e-07 $l=3.58e-07 $layer=LI1_cond $X=4.052 $Y=1.003
+ $X2=4.052 $Y2=0.645
r34 2 14 400 $w=1.7e-07 $l=2.38485e-07 $layer=licon1_PDIFF $count=1 $X=3.89
+ $Y=1.84 $X2=4.04 $Y2=2.015
r35 2 16 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=3.89
+ $Y=1.84 $X2=4.04 $Y2=2.815
r36 1 9 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.9 $Y=0.5
+ $X2=4.04 $Y2=0.645
.ends

.subckt PM_SKY130_FD_SC_HS__AND4B_1%VGND 1 2 9 13 15 17 22 32 33 36 39
r42 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r43 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r44 33 40 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=3.6
+ $Y2=0
r45 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r46 30 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.705 $Y=0 $X2=3.54
+ $Y2=0
r47 30 32 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=3.705 $Y=0 $X2=4.08
+ $Y2=0
r48 29 40 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=3.6
+ $Y2=0
r49 28 29 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r50 26 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r51 25 28 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=1.2 $Y=0 $X2=3.12
+ $Y2=0
r52 25 26 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r53 23 36 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=0.875 $Y=0 $X2=0.725
+ $Y2=0
r54 23 25 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.875 $Y=0 $X2=1.2
+ $Y2=0
r55 22 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.375 $Y=0 $X2=3.54
+ $Y2=0
r56 22 28 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=3.375 $Y=0 $X2=3.12
+ $Y2=0
r57 20 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r58 19 20 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r59 17 36 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=0.575 $Y=0 $X2=0.725
+ $Y2=0
r60 17 19 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=0.575 $Y=0 $X2=0.24
+ $Y2=0
r61 15 29 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=3.12
+ $Y2=0
r62 15 26 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.2
+ $Y2=0
r63 11 39 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.54 $Y=0.085
+ $X2=3.54 $Y2=0
r64 11 13 27.5888 $w=3.28e-07 $l=7.9e-07 $layer=LI1_cond $X=3.54 $Y=0.085
+ $X2=3.54 $Y2=0.875
r65 7 36 0.597483 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.725 $Y=0.085
+ $X2=0.725 $Y2=0
r66 7 9 16.5184 $w=2.98e-07 $l=4.3e-07 $layer=LI1_cond $X=0.725 $Y=0.085
+ $X2=0.725 $Y2=0.515
r67 2 13 182 $w=1.7e-07 $l=3.68951e-07 $layer=licon1_NDIFF $count=1 $X=3.32
+ $Y=0.6 $X2=3.54 $Y2=0.875
r68 1 9 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.37 $X2=0.71 $Y2=0.515
.ends

