* File: sky130_fd_sc_hs__a21o_2.pex.spice
* Created: Tue Sep  1 19:49:39 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HS__A21O_2%A_84_244# 1 2 7 9 10 12 13 15 16 18 19 22 26
+ 27 28 30 36 38 46
c87 22 0 1.09867e-19 $X=1.23 $Y=1.385
r88 45 46 17.088 $w=4.09e-07 $l=1.45e-07 $layer=POLY_cond $X=0.96 $Y=1.492
+ $X2=1.105 $Y2=1.492
r89 44 45 33.5868 $w=4.09e-07 $l=2.85e-07 $layer=POLY_cond $X=0.675 $Y=1.492
+ $X2=0.96 $Y2=1.492
r90 43 44 19.445 $w=4.09e-07 $l=1.65e-07 $layer=POLY_cond $X=0.51 $Y=1.492
+ $X2=0.675 $Y2=1.492
r91 34 36 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=2.13 $Y=0.84
+ $X2=2.13 $Y2=0.495
r92 30 32 32.7294 $w=2.48e-07 $l=7.1e-07 $layer=LI1_cond $X=1.665 $Y=2.105
+ $X2=1.665 $Y2=2.815
r93 28 30 10.6025 $w=2.48e-07 $l=2.3e-07 $layer=LI1_cond $X=1.665 $Y=1.875
+ $X2=1.665 $Y2=2.105
r94 26 34 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.965 $Y=0.925
+ $X2=2.13 $Y2=0.84
r95 26 27 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=1.965 $Y=0.925
+ $X2=1.395 $Y2=0.925
r96 24 27 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.31 $Y=1.01
+ $X2=1.395 $Y2=0.925
r97 24 38 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=1.31 $Y=1.01
+ $X2=1.31 $Y2=1.22
r98 23 46 14.7311 $w=4.09e-07 $l=1.25e-07 $layer=POLY_cond $X=1.23 $Y=1.492
+ $X2=1.105 $Y2=1.492
r99 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.23
+ $Y=1.385 $X2=1.23 $Y2=1.385
r100 20 28 28.2492 $w=1.68e-07 $l=4.33e-07 $layer=LI1_cond $X=1.232 $Y=1.79
+ $X2=1.665 $Y2=1.79
r101 20 22 11.3471 $w=3.23e-07 $l=3.2e-07 $layer=LI1_cond $X=1.232 $Y=1.705
+ $X2=1.232 $Y2=1.385
r102 19 38 8.35379 $w=3.23e-07 $l=1.62e-07 $layer=LI1_cond $X=1.232 $Y=1.382
+ $X2=1.232 $Y2=1.22
r103 19 22 0.106379 $w=3.23e-07 $l=3e-09 $layer=LI1_cond $X=1.232 $Y=1.382
+ $X2=1.232 $Y2=1.385
r104 16 46 26.4068 $w=1.5e-07 $l=2.72e-07 $layer=POLY_cond $X=1.105 $Y=1.22
+ $X2=1.105 $Y2=1.492
r105 16 18 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.105 $Y=1.22
+ $X2=1.105 $Y2=0.74
r106 13 45 26.4068 $w=1.5e-07 $l=2.73e-07 $layer=POLY_cond $X=0.96 $Y=1.765
+ $X2=0.96 $Y2=1.492
r107 13 15 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.96 $Y=1.765
+ $X2=0.96 $Y2=2.4
r108 10 44 26.4068 $w=1.5e-07 $l=2.72e-07 $layer=POLY_cond $X=0.675 $Y=1.22
+ $X2=0.675 $Y2=1.492
r109 10 12 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=0.675 $Y=1.22
+ $X2=0.675 $Y2=0.74
r110 7 43 26.4068 $w=1.5e-07 $l=2.73e-07 $layer=POLY_cond $X=0.51 $Y=1.765
+ $X2=0.51 $Y2=1.492
r111 7 9 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.51 $Y=1.765
+ $X2=0.51 $Y2=2.4
r112 2 32 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=1.58
+ $Y=1.96 $X2=1.705 $Y2=2.815
r113 2 30 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=1.58
+ $Y=1.96 $X2=1.705 $Y2=2.105
r114 1 36 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=1.99
+ $Y=0.37 $X2=2.13 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_HS__A21O_2%B1 3 8 9 10 11 14 15 16
c39 16 0 1.57121e-19 $X=1.825 $Y=1.22
c40 15 0 4.3623e-20 $X=1.825 $Y=1.385
c41 14 0 1.09867e-19 $X=1.825 $Y=1.385
r42 14 17 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.825 $Y=1.385
+ $X2=1.825 $Y2=1.55
r43 14 16 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.825 $Y=1.385
+ $X2=1.825 $Y2=1.22
r44 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.825
+ $Y=1.385 $X2=1.825 $Y2=1.385
r45 11 15 4.70716 $w=3.53e-07 $l=1.45e-07 $layer=LI1_cond $X=1.68 $Y=1.357
+ $X2=1.825 $Y2=1.357
r46 9 10 41.3838 $w=1.65e-07 $l=9.5e-08 $layer=POLY_cond $X=1.922 $Y=1.79
+ $X2=1.922 $Y2=1.885
r47 9 17 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=1.915 $Y=1.79
+ $X2=1.915 $Y2=1.55
r48 8 10 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=1.93 $Y=2.46
+ $X2=1.93 $Y2=1.885
r49 3 16 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.915 $Y=0.74
+ $X2=1.915 $Y2=1.22
.ends

.subckt PM_SKY130_FD_SC_HS__A21O_2%A1 3 5 6 8 9 12 14
c40 14 0 4.3623e-20 $X=2.365 $Y=1.22
c41 9 0 1.57121e-19 $X=2.64 $Y=1.295
r42 12 15 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.365 $Y=1.385
+ $X2=2.365 $Y2=1.55
r43 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.365 $Y=1.385
+ $X2=2.365 $Y2=1.22
r44 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.365
+ $Y=1.385 $X2=2.365 $Y2=1.385
r45 9 13 8.56545 $w=3.68e-07 $l=2.75e-07 $layer=LI1_cond $X=2.64 $Y=1.365
+ $X2=2.365 $Y2=1.365
r46 6 8 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=2.38 $Y=1.885
+ $X2=2.38 $Y2=2.46
r47 5 6 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=2.38 $Y=1.795 $X2=2.38
+ $Y2=1.885
r48 5 15 95.2339 $w=1.8e-07 $l=2.45e-07 $layer=POLY_cond $X=2.38 $Y=1.795
+ $X2=2.38 $Y2=1.55
r49 3 14 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=2.345 $Y=0.74
+ $X2=2.345 $Y2=1.22
.ends

.subckt PM_SKY130_FD_SC_HS__A21O_2%A2 1 3 6 9 10 11 17
r30 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.09
+ $Y=1.385 $X2=3.09 $Y2=1.385
r31 15 17 42.841 $w=3.3e-07 $l=2.45e-07 $layer=POLY_cond $X=2.845 $Y=1.385
+ $X2=3.09 $Y2=1.385
r32 13 15 5.24584 $w=3.3e-07 $l=3e-08 $layer=POLY_cond $X=2.815 $Y=1.385
+ $X2=2.845 $Y2=1.385
r33 11 18 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=3.09 $Y=1.295 $X2=3.09
+ $Y2=1.385
r34 9 10 41.3838 $w=1.65e-07 $l=9.5e-08 $layer=POLY_cond $X=2.837 $Y=1.79
+ $X2=2.837 $Y2=1.885
r35 7 15 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.845 $Y=1.55
+ $X2=2.845 $Y2=1.385
r36 7 9 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=2.845 $Y=1.55
+ $X2=2.845 $Y2=1.79
r37 6 10 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=2.83 $Y=2.46
+ $X2=2.83 $Y2=1.885
r38 1 13 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.815 $Y=1.22
+ $X2=2.815 $Y2=1.385
r39 1 3 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=2.815 $Y=1.22 $X2=2.815
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HS__A21O_2%VPWR 1 2 3 10 12 18 24 28 30 35 42 43 49 52
r44 52 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r45 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r46 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r47 43 53 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=2.64 $Y2=3.33
r48 42 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r49 40 52 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.77 $Y=3.33
+ $X2=2.605 $Y2=3.33
r50 40 42 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=2.77 $Y=3.33
+ $X2=3.12 $Y2=3.33
r51 39 53 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r52 38 39 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r53 36 49 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.35 $Y=3.33
+ $X2=1.185 $Y2=3.33
r54 36 38 52.8449 $w=1.68e-07 $l=8.1e-07 $layer=LI1_cond $X=1.35 $Y=3.33
+ $X2=2.16 $Y2=3.33
r55 35 52 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.44 $Y=3.33
+ $X2=2.605 $Y2=3.33
r56 35 38 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=2.44 $Y=3.33
+ $X2=2.16 $Y2=3.33
r57 34 50 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r58 34 47 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r59 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r60 31 46 4.0045 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=0.37 $Y=3.33
+ $X2=0.185 $Y2=3.33
r61 31 33 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=0.37 $Y=3.33
+ $X2=0.72 $Y2=3.33
r62 30 49 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.02 $Y=3.33
+ $X2=1.185 $Y2=3.33
r63 30 33 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=1.02 $Y=3.33 $X2=0.72
+ $Y2=3.33
r64 28 39 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r65 28 50 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r66 24 27 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=2.605 $Y=2.155
+ $X2=2.605 $Y2=2.835
r67 22 52 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.605 $Y=3.245
+ $X2=2.605 $Y2=3.33
r68 22 27 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=2.605 $Y=3.245
+ $X2=2.605 $Y2=2.835
r69 18 21 23.9219 $w=3.28e-07 $l=6.85e-07 $layer=LI1_cond $X=1.185 $Y=2.13
+ $X2=1.185 $Y2=2.815
r70 16 49 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.185 $Y=3.245
+ $X2=1.185 $Y2=3.33
r71 16 21 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=1.185 $Y=3.245
+ $X2=1.185 $Y2=2.815
r72 12 15 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=0.245 $Y=1.985
+ $X2=0.245 $Y2=2.815
r73 10 46 3.13866 $w=2.5e-07 $l=1.11018e-07 $layer=LI1_cond $X=0.245 $Y=3.245
+ $X2=0.185 $Y2=3.33
r74 10 15 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=0.245 $Y=3.245
+ $X2=0.245 $Y2=2.815
r75 3 27 400 $w=1.7e-07 $l=9.47035e-07 $layer=licon1_PDIFF $count=1 $X=2.455
+ $Y=1.96 $X2=2.605 $Y2=2.835
r76 3 24 400 $w=1.7e-07 $l=2.59374e-07 $layer=licon1_PDIFF $count=1 $X=2.455
+ $Y=1.96 $X2=2.605 $Y2=2.155
r77 2 21 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=1.035
+ $Y=1.84 $X2=1.185 $Y2=2.815
r78 2 18 400 $w=1.7e-07 $l=3.57211e-07 $layer=licon1_PDIFF $count=1 $X=1.035
+ $Y=1.84 $X2=1.185 $Y2=2.13
r79 1 15 400 $w=1.7e-07 $l=1.03562e-06 $layer=licon1_PDIFF $count=1 $X=0.16
+ $Y=1.84 $X2=0.285 $Y2=2.815
r80 1 12 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.16
+ $Y=1.84 $X2=0.285 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HS__A21O_2%X 1 2 9 13 14 15 16 17 33
r29 16 17 15.2287 $w=2.78e-07 $l=3.7e-07 $layer=LI1_cond $X=0.71 $Y=2.405
+ $X2=0.71 $Y2=2.775
r30 15 16 17.2866 $w=2.78e-07 $l=4.2e-07 $layer=LI1_cond $X=0.71 $Y=1.985
+ $X2=0.71 $Y2=2.405
r31 15 35 3.91007 $w=2.78e-07 $l=9.5e-08 $layer=LI1_cond $X=0.71 $Y=1.985
+ $X2=0.71 $Y2=1.89
r32 14 35 8.1553 $w=3.28e-07 $l=2.25e-07 $layer=LI1_cond $X=0.735 $Y=1.665
+ $X2=0.735 $Y2=1.89
r33 14 33 6.54453 $w=3.28e-07 $l=1.15e-07 $layer=LI1_cond $X=0.735 $Y=1.665
+ $X2=0.735 $Y2=1.55
r34 13 33 31.6883 $w=1.73e-07 $l=5e-07 $layer=LI1_cond $X=0.812 $Y=1.05
+ $X2=0.812 $Y2=1.55
r35 7 13 8.29065 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=0.89 $Y=0.885
+ $X2=0.89 $Y2=1.05
r36 7 9 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=0.89 $Y=0.885 $X2=0.89
+ $Y2=0.515
r37 2 17 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=1.84 $X2=0.735 $Y2=2.815
r38 2 15 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=1.84 $X2=0.735 $Y2=1.985
r39 1 9 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=0.75
+ $Y=0.37 $X2=0.89 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__A21O_2%A_401_392# 1 2 9 13 14 17
r29 17 19 32.7294 $w=2.48e-07 $l=7.1e-07 $layer=LI1_cond $X=3.095 $Y=2.105
+ $X2=3.095 $Y2=2.815
r30 15 17 9.91101 $w=2.48e-07 $l=2.15e-07 $layer=LI1_cond $X=3.095 $Y=1.89
+ $X2=3.095 $Y2=2.105
r31 13 15 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=2.97 $Y=1.805
+ $X2=3.095 $Y2=1.89
r32 13 14 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=2.97 $Y=1.805
+ $X2=2.24 $Y2=1.805
r33 9 11 32.7294 $w=2.48e-07 $l=7.1e-07 $layer=LI1_cond $X=2.115 $Y=2.105
+ $X2=2.115 $Y2=2.815
r34 7 14 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=2.115 $Y=1.89
+ $X2=2.24 $Y2=1.805
r35 7 9 9.91101 $w=2.48e-07 $l=2.15e-07 $layer=LI1_cond $X=2.115 $Y=1.89
+ $X2=2.115 $Y2=2.105
r36 2 19 400 $w=1.7e-07 $l=9.26971e-07 $layer=licon1_PDIFF $count=1 $X=2.905
+ $Y=1.96 $X2=3.055 $Y2=2.815
r37 2 17 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=2.905
+ $Y=1.96 $X2=3.055 $Y2=2.105
r38 1 11 400 $w=1.7e-07 $l=9.26971e-07 $layer=licon1_PDIFF $count=1 $X=2.005
+ $Y=1.96 $X2=2.155 $Y2=2.815
r39 1 9 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=2.005
+ $Y=1.96 $X2=2.155 $Y2=2.105
.ends

.subckt PM_SKY130_FD_SC_HS__A21O_2%VGND 1 2 3 12 16 18 20 23 24 25 30 34 40 44
r45 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r46 38 44 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r47 37 38 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r48 35 40 12.1981 $w=1.7e-07 $l=2.85e-07 $layer=LI1_cond $X=1.795 $Y=0 $X2=1.51
+ $Y2=0
r49 35 37 55.1283 $w=1.68e-07 $l=8.45e-07 $layer=LI1_cond $X=1.795 $Y=0 $X2=2.64
+ $Y2=0
r50 34 43 4.63344 $w=1.7e-07 $l=2.47e-07 $layer=LI1_cond $X=2.865 $Y=0 $X2=3.112
+ $Y2=0
r51 34 37 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=2.865 $Y=0 $X2=2.64
+ $Y2=0
r52 32 33 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r53 30 40 12.1981 $w=1.7e-07 $l=2.85e-07 $layer=LI1_cond $X=1.225 $Y=0 $X2=1.51
+ $Y2=0
r54 30 32 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=1.225 $Y=0 $X2=1.2
+ $Y2=0
r55 29 33 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=1.2
+ $Y2=0
r56 28 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r57 25 38 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.64
+ $Y2=0
r58 25 33 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r59 25 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r60 23 28 3.94706 $w=1.7e-07 $l=5.5e-08 $layer=LI1_cond $X=0.295 $Y=0 $X2=0.24
+ $Y2=0
r61 23 24 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.295 $Y=0 $X2=0.42
+ $Y2=0
r62 22 32 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=0.545 $Y=0 $X2=1.2
+ $Y2=0
r63 22 24 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.545 $Y=0 $X2=0.42
+ $Y2=0
r64 18 43 3.13273 $w=3.3e-07 $l=1.19143e-07 $layer=LI1_cond $X=3.03 $Y=0.085
+ $X2=3.112 $Y2=0
r65 18 20 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=3.03 $Y=0.085
+ $X2=3.03 $Y2=0.515
r66 14 40 2.39972 $w=5.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.51 $Y=0.085
+ $X2=1.51 $Y2=0
r67 14 16 8.81321 $w=5.68e-07 $l=4.2e-07 $layer=LI1_cond $X=1.51 $Y=0.085
+ $X2=1.51 $Y2=0.505
r68 10 24 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.42 $Y=0.085
+ $X2=0.42 $Y2=0
r69 10 12 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=0.42 $Y=0.085
+ $X2=0.42 $Y2=0.515
r70 3 20 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.89
+ $Y=0.37 $X2=3.03 $Y2=0.515
r71 2 16 91 $w=1.7e-07 $l=5.83609e-07 $layer=licon1_NDIFF $count=2 $X=1.18
+ $Y=0.37 $X2=1.7 $Y2=0.505
r72 1 12 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.335
+ $Y=0.37 $X2=0.46 $Y2=0.515
.ends

