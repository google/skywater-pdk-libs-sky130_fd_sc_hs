* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hs__einvp_1 A TE VGND VNB VPB VPWR Z
M1000 VPWR TE a_44_549# VPB pshort w=420000u l=150000u
+  ad=3.328e+11p pd=2.77e+06u as=2.646e+11p ps=2.1e+06u
M1001 a_318_74# TE VGND VNB nlowvt w=740000u l=150000u
+  ad=1.776e+11p pd=1.96e+06u as=2.276e+11p ps=2.16e+06u
M1002 Z A a_318_74# VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1003 VGND TE a_44_549# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=2.604e+11p ps=2.08e+06u
M1004 a_310_392# a_44_549# VPWR VPB pshort w=1e+06u l=150000u
+  ad=2.7e+11p pd=2.54e+06u as=0p ps=0u
M1005 Z A a_310_392# VPB pshort w=1e+06u l=150000u
+  ad=2.95e+11p pd=2.59e+06u as=0p ps=0u
.ends
