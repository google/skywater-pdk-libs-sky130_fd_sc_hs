# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_hs__o211a_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__o211a_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  6.720000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.075000 1.450000 6.595000 1.780000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.925000 1.450000 5.835000 1.780000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.444000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.505000 1.435000 2.835000 1.780000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.444000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.450000 1.450000 3.780000 1.780000 ;
    END
  END C1
  PIN X
    ANTENNADIFFAREA  1.086400 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 0.960000 1.760000 1.130000 ;
        RECT 0.125000 1.130000 0.355000 1.800000 ;
        RECT 0.125000 1.800000 1.945000 1.970000 ;
        RECT 0.580000 0.350000 0.830000 0.960000 ;
        RECT 0.615000 1.970000 0.945000 2.980000 ;
        RECT 1.510000 0.350000 1.760000 0.960000 ;
        RECT 1.615000 1.970000 1.945000 2.980000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 6.720000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 6.720000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 6.720000 0.085000 ;
      RECT 0.000000  3.245000 6.720000 3.415000 ;
      RECT 0.115000  2.140000 0.445000 3.245000 ;
      RECT 0.150000  0.085000 0.400000 0.790000 ;
      RECT 0.615000  1.300000 2.285000 1.630000 ;
      RECT 1.010000  0.085000 1.340000 0.790000 ;
      RECT 1.115000  2.140000 1.445000 3.245000 ;
      RECT 1.940000  0.085000 2.270000 1.130000 ;
      RECT 2.115000  1.630000 2.285000 1.950000 ;
      RECT 2.115000  1.950000 5.655000 2.120000 ;
      RECT 2.115000  2.290000 2.445000 3.245000 ;
      RECT 2.530000  0.255000 4.650000 0.425000 ;
      RECT 2.530000  0.425000 2.780000 1.265000 ;
      RECT 2.775000  2.120000 3.105000 2.815000 ;
      RECT 3.040000  0.595000 4.220000 0.765000 ;
      RECT 3.040000  0.765000 3.210000 1.285000 ;
      RECT 3.275000  2.290000 3.605000 3.245000 ;
      RECT 3.390000  0.935000 3.720000 1.110000 ;
      RECT 3.390000  1.110000 4.120000 1.280000 ;
      RECT 3.790000  2.120000 4.120000 2.815000 ;
      RECT 3.890000  0.765000 4.220000 0.940000 ;
      RECT 3.950000  1.280000 4.120000 1.950000 ;
      RECT 4.325000  2.290000 4.655000 3.245000 ;
      RECT 4.400000  0.425000 4.650000 1.110000 ;
      RECT 4.400000  1.110000 6.605000 1.280000 ;
      RECT 4.400000  1.280000 4.650000 1.285000 ;
      RECT 4.825000  2.290000 5.155000 2.905000 ;
      RECT 4.825000  2.905000 6.105000 3.075000 ;
      RECT 4.830000  0.085000 5.175000 0.935000 ;
      RECT 5.325000  2.120000 5.655000 2.735000 ;
      RECT 5.345000  0.605000 5.595000 1.110000 ;
      RECT 5.775000  0.085000 6.105000 0.940000 ;
      RECT 5.855000  1.950000 6.105000 2.905000 ;
      RECT 6.275000  0.605000 6.605000 1.110000 ;
      RECT 6.275000  1.950000 6.605000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
  END
END sky130_fd_sc_hs__o211a_4
END LIBRARY
