* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hs__sdfxtp_1 CLK D SCD SCE VGND VNB VPB VPWR Q
M1000 a_1520_74# a_828_74# a_1239_74# VNB nlowvt w=550000u l=150000u
+  ad=3.223e+11p pd=2.48e+06u as=1.5675e+11p ps=1.67e+06u
M1001 VPWR a_1736_74# a_1688_508# VPB pshort w=420000u l=150000u
+  ad=2.3028e+12p pd=1.727e+07u as=1.134e+11p ps=1.38e+06u
M1002 VPWR a_1239_74# a_1202_508# VPB pshort w=420000u l=150000u
+  ad=0p pd=0u as=1.05e+11p ps=1.34e+06u
M1003 a_630_74# CLK VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=1.52935e+12p ps=1.307e+07u
M1004 VGND a_1736_74# a_1688_100# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1005 a_301_74# D a_238_464# VPB pshort w=640000u l=150000u
+  ad=3.159e+11p pd=3.31e+06u as=1.728e+11p ps=1.82e+06u
M1006 VGND SCE a_35_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.197e+11p ps=1.41e+06u
M1007 a_1018_100# a_630_74# a_301_74# VNB nlowvt w=420000u l=150000u
+  ad=2.226e+11p pd=1.9e+06u as=3.612e+11p ps=3.4e+06u
M1008 a_1736_74# a_1520_74# VGND VNB nlowvt w=550000u l=150000u
+  ad=1.4575e+11p pd=1.63e+06u as=0p ps=0u
M1009 a_412_464# a_35_74# a_301_74# VPB pshort w=640000u l=150000u
+  ad=2.496e+11p pd=2.06e+06u as=0p ps=0u
M1010 a_1239_74# a_1018_100# VGND VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 Q a_1736_74# VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=3.248e+11p pd=2.82e+06u as=0p ps=0u
M1012 Q a_1736_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.035e+11p pd=2.03e+06u as=0p ps=0u
M1013 a_828_74# a_630_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=1.961e+11p pd=2.01e+06u as=0p ps=0u
M1014 a_223_74# a_35_74# VGND VNB nlowvt w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=0p ps=0u
M1015 a_301_74# D a_223_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_1688_508# a_828_74# a_1520_74# VPB pshort w=420000u l=150000u
+  ad=0p pd=0u as=3.927e+11p ps=2.79e+06u
M1017 a_1688_100# a_630_74# a_1520_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 VGND a_1239_74# a_1154_100# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.785e+11p ps=1.69e+06u
M1019 VPWR SCE a_35_74# VPB pshort w=640000u l=150000u
+  ad=0p pd=0u as=1.888e+11p ps=1.87e+06u
M1020 a_238_464# SCE VPWR VPB pshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_1736_74# a_1520_74# VPWR VPB pshort w=840000u l=150000u
+  ad=2.478e+11p pd=2.27e+06u as=0p ps=0u
M1022 VPWR SCD a_412_464# VPB pshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_1239_74# a_1018_100# VPWR VPB pshort w=840000u l=150000u
+  ad=4.662e+11p pd=2.79e+06u as=0p ps=0u
M1024 VGND SCD a_450_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1025 a_630_74# CLK VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=3.304e+11p pd=2.83e+06u as=0p ps=0u
M1026 a_450_74# SCE a_301_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 a_828_74# a_630_74# VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=3.304e+11p pd=2.83e+06u as=0p ps=0u
M1028 a_1154_100# a_828_74# a_1018_100# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1029 a_1202_508# a_630_74# a_1018_100# VPB pshort w=420000u l=150000u
+  ad=0p pd=0u as=1.47e+11p ps=1.54e+06u
M1030 a_1520_74# a_630_74# a_1239_74# VPB pshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1031 a_1018_100# a_828_74# a_301_74# VPB pshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
