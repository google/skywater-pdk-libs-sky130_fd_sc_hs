* File: sky130_fd_sc_hs__nor4bb_4.spice
* Created: Tue Sep  1 20:12:52 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hs__nor4bb_4.pex.spice"
.subckt sky130_fd_sc_hs__nor4bb_4  VNB VPB B A C_N D_N VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* D_N	D_N
* C_N	C_N
* A	A
* B	B
* VPB	VPB
* VNB	VNB
MM1001 N_Y_M1001_d N_B_M1001_g N_VGND_M1001_s VNB NLOWVT L=0.15 W=0.74 AD=0.1036
+ AS=0.2627 PD=1.02 PS=2.19 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75000.3 SB=75008.9
+ A=0.111 P=1.78 MULT=1
MM1011 N_VGND_M1011_d N_A_M1011_g N_Y_M1001_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.13875 AS=0.1036 PD=1.115 PS=1.02 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75000.7
+ SB=75008.4 A=0.111 P=1.78 MULT=1
MM1017 N_VGND_M1011_d N_A_M1017_g N_Y_M1017_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.13875 AS=0.12025 PD=1.115 PS=1.065 NRD=4.044 NRS=7.296 M=1 R=4.93333
+ SA=75001.2 SB=75007.9 A=0.111 P=1.78 MULT=1
MM1023 N_VGND_M1023_d N_A_M1023_g N_Y_M1017_s VNB NLOWVT L=0.15 W=0.74 AD=0.1443
+ AS=0.12025 PD=1.13 PS=1.065 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75001.7
+ SB=75007.4 A=0.111 P=1.78 MULT=1
MM1031 N_VGND_M1023_d N_A_M1031_g N_Y_M1031_s VNB NLOWVT L=0.15 W=0.74 AD=0.1443
+ AS=0.111 PD=1.13 PS=1.04 NRD=6.48 NRS=0 M=1 R=4.93333 SA=75002.2 SB=75006.9
+ A=0.111 P=1.78 MULT=1
MM1020 N_Y_M1031_s N_B_M1020_g N_VGND_M1020_s VNB NLOWVT L=0.15 W=0.74 AD=0.111
+ AS=0.1221 PD=1.04 PS=1.07 NRD=3.24 NRS=8.1 M=1 R=4.93333 SA=75002.7 SB=75006.4
+ A=0.111 P=1.78 MULT=1
MM1028 N_Y_M1028_d N_B_M1028_g N_VGND_M1020_s VNB NLOWVT L=0.15 W=0.74 AD=0.1295
+ AS=0.1221 PD=1.09 PS=1.07 NRD=0 NRS=0 M=1 R=4.93333 SA=75003.2 SB=75005.9
+ A=0.111 P=1.78 MULT=1
MM1034 N_Y_M1028_d N_B_M1034_g N_VGND_M1034_s VNB NLOWVT L=0.15 W=0.74 AD=0.1295
+ AS=0.1036 PD=1.09 PS=1.02 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75003.7 SB=75005.5
+ A=0.111 P=1.78 MULT=1
MM1009 N_VGND_M1034_s N_A_864_48#_M1009_g N_Y_M1009_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1295 PD=1.02 PS=1.09 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75004.1
+ SB=75005 A=0.111 P=1.78 MULT=1
MM1014 N_VGND_M1014_d N_A_864_48#_M1014_g N_Y_M1009_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1295 AS=0.1295 PD=1.09 PS=1.09 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75004.6
+ SB=75004.5 A=0.111 P=1.78 MULT=1
MM1035 N_VGND_M1014_d N_A_864_48#_M1035_g N_Y_M1035_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1295 AS=0.1258 PD=1.09 PS=1.08 NRD=0 NRS=0 M=1 R=4.93333 SA=75005.1
+ SB=75004 A=0.111 P=1.78 MULT=1
MM1004 N_VGND_M1004_d N_A_1162_48#_M1004_g N_Y_M1035_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1332 AS=0.1258 PD=1.1 PS=1.08 NRD=1.62 NRS=9.72 M=1 R=4.93333 SA=75005.6
+ SB=75003.5 A=0.111 P=1.78 MULT=1
MM1005 N_VGND_M1004_d N_A_1162_48#_M1005_g N_Y_M1005_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1332 AS=0.1036 PD=1.1 PS=1.02 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75006.1
+ SB=75003 A=0.111 P=1.78 MULT=1
MM1018 N_VGND_M1018_d N_A_1162_48#_M1018_g N_Y_M1005_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.2516 AS=0.1036 PD=1.42 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75006.5
+ SB=75002.6 A=0.111 P=1.78 MULT=1
MM1030 N_VGND_M1018_d N_A_1162_48#_M1030_g N_Y_M1030_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.2516 AS=0.11285 PD=1.42 PS=1.045 NRD=0 NRS=0 M=1 R=4.93333 SA=75007.4
+ SB=75001.8 A=0.111 P=1.78 MULT=1
MM1036 N_VGND_M1036_d N_A_864_48#_M1036_g N_Y_M1030_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.34965 AS=0.11285 PD=1.685 PS=1.045 NRD=0 NRS=4.044 M=1 R=4.93333
+ SA=75007.8 SB=75001.3 A=0.111 P=1.78 MULT=1
MM1025 N_A_864_48#_M1025_d N_C_N_M1025_g N_VGND_M1036_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.34965 PD=2.05 PS=1.685 NRD=0 NRS=52.692 M=1 R=4.93333
+ SA=75008.9 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1008 N_A_1162_48#_M1008_d N_D_N_M1008_g N_VGND_M1008_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.2109 AS=0.2627 PD=2.05 PS=2.19 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.3 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1010 N_A_27_368#_M1010_d N_B_M1010_g N_A_116_368#_M1010_s VPB PSHORT L=0.15
+ W=1.12 AD=0.3304 AS=0.196 PD=2.83 PS=1.47 NRD=1.7533 NRS=10.5395 M=1 R=7.46667
+ SA=75000.2 SB=75007.4 A=0.168 P=2.54 MULT=1
MM1021 N_VPWR_M1021_d N_A_M1021_g N_A_116_368#_M1010_s VPB PSHORT L=0.15 W=1.12
+ AD=0.196 AS=0.196 PD=1.47 PS=1.47 NRD=10.5395 NRS=1.7533 M=1 R=7.46667
+ SA=75000.7 SB=75006.9 A=0.168 P=2.54 MULT=1
MM1022 N_VPWR_M1021_d N_A_M1022_g N_A_116_368#_M1022_s VPB PSHORT L=0.15 W=1.12
+ AD=0.196 AS=0.168 PD=1.47 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.2 SB=75006.4 A=0.168 P=2.54 MULT=1
MM1024 N_VPWR_M1024_d N_A_M1024_g N_A_116_368#_M1022_s VPB PSHORT L=0.15 W=1.12
+ AD=0.2184 AS=0.168 PD=1.51 PS=1.42 NRD=14.0658 NRS=1.7533 M=1 R=7.46667
+ SA=75001.7 SB=75005.9 A=0.168 P=2.54 MULT=1
MM1033 N_VPWR_M1024_d N_A_M1033_g N_A_116_368#_M1033_s VPB PSHORT L=0.15 W=1.12
+ AD=0.2184 AS=0.207112 PD=1.51 PS=1.57 NRD=5.2599 NRS=1.7533 M=1 R=7.46667
+ SA=75002.2 SB=75005.4 A=0.168 P=2.54 MULT=1
MM1012 N_A_27_368#_M1012_d N_B_M1012_g N_A_116_368#_M1033_s VPB PSHORT L=0.15
+ W=1.12 AD=0.168 AS=0.207112 PD=1.42 PS=1.57 NRD=1.7533 NRS=11.426 M=1
+ R=7.46667 SA=75002.5 SB=75005.3 A=0.168 P=2.54 MULT=1
MM1015 N_A_27_368#_M1012_d N_B_M1015_g N_A_116_368#_M1015_s VPB PSHORT L=0.15
+ W=1.12 AD=0.168 AS=0.196 PD=1.42 PS=1.47 NRD=1.7533 NRS=10.5395 M=1 R=7.46667
+ SA=75003 SB=75004.9 A=0.168 P=2.54 MULT=1
MM1027 N_A_27_368#_M1027_d N_B_M1027_g N_A_116_368#_M1015_s VPB PSHORT L=0.15
+ W=1.12 AD=0.1736 AS=0.196 PD=1.43 PS=1.47 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75003.5 SB=75004.4 A=0.168 P=2.54 MULT=1
MM1007 N_A_27_368#_M1027_d N_A_864_48#_M1007_g N_A_897_349#_M1007_s VPB PSHORT
+ L=0.15 W=1.12 AD=0.1736 AS=0.168 PD=1.43 PS=1.42 NRD=3.5066 NRS=1.7533 M=1
+ R=7.46667 SA=75003.9 SB=75003.9 A=0.168 P=2.54 MULT=1
MM1013 N_A_27_368#_M1013_d N_A_864_48#_M1013_g N_A_897_349#_M1007_s VPB PSHORT
+ L=0.15 W=1.12 AD=0.30235 AS=0.168 PD=1.86 PS=1.42 NRD=37.8043 NRS=1.7533 M=1
+ R=7.46667 SA=75004.4 SB=75003.5 A=0.168 P=2.54 MULT=1
MM1032 N_A_27_368#_M1013_d N_A_864_48#_M1032_g N_A_897_349#_M1032_s VPB PSHORT
+ L=0.15 W=1.12 AD=0.30235 AS=0.168 PD=1.86 PS=1.42 NRD=37.8043 NRS=1.7533 M=1
+ R=7.46667 SA=75005 SB=75002.9 A=0.168 P=2.54 MULT=1
MM1002 N_Y_M1002_d N_A_1162_48#_M1002_g N_A_897_349#_M1032_s VPB PSHORT L=0.15
+ W=1.12 AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75005.4 SB=75002.4 A=0.168 P=2.54 MULT=1
MM1006 N_Y_M1002_d N_A_1162_48#_M1006_g N_A_897_349#_M1006_s VPB PSHORT L=0.15
+ W=1.12 AD=0.168 AS=0.1736 PD=1.42 PS=1.43 NRD=1.7533 NRS=2.6201 M=1 R=7.46667
+ SA=75005.9 SB=75002 A=0.168 P=2.54 MULT=1
MM1016 N_Y_M1016_d N_A_1162_48#_M1016_g N_A_897_349#_M1006_s VPB PSHORT L=0.15
+ W=1.12 AD=0.168 AS=0.1736 PD=1.42 PS=1.43 NRD=1.7533 NRS=2.6201 M=1 R=7.46667
+ SA=75006.3 SB=75001.5 A=0.168 P=2.54 MULT=1
MM1019 N_Y_M1016_d N_A_1162_48#_M1019_g N_A_897_349#_M1019_s VPB PSHORT L=0.15
+ W=1.12 AD=0.168 AS=0.3668 PD=1.42 PS=1.775 NRD=1.7533 NRS=32.9778 M=1
+ R=7.46667 SA=75006.8 SB=75001.1 A=0.168 P=2.54 MULT=1
MM1037 N_A_27_368#_M1037_d N_A_864_48#_M1037_g N_A_897_349#_M1019_s VPB PSHORT
+ L=0.15 W=1.12 AD=0.364 AS=0.3668 PD=2.89 PS=1.775 NRD=2.6201 NRS=1.7533 M=1
+ R=7.46667 SA=75007.6 SB=75000.2 A=0.168 P=2.54 MULT=1
MM1000 N_A_864_48#_M1000_d N_C_N_M1000_g N_VPWR_M1000_s VPB PSHORT L=0.15 W=0.84
+ AD=0.126 AS=0.2898 PD=1.14 PS=2.37 NRD=2.3443 NRS=3.5066 M=1 R=5.6 SA=75000.3
+ SB=75001.6 A=0.126 P=1.98 MULT=1
MM1003 N_A_864_48#_M1000_d N_C_N_M1003_g N_VPWR_M1003_s VPB PSHORT L=0.15 W=0.84
+ AD=0.126 AS=0.126 PD=1.14 PS=1.14 NRD=2.3443 NRS=2.3443 M=1 R=5.6 SA=75000.7
+ SB=75001.1 A=0.126 P=1.98 MULT=1
MM1026 N_A_1162_48#_M1026_d N_D_N_M1026_g N_VPWR_M1003_s VPB PSHORT L=0.15
+ W=0.84 AD=0.126 AS=0.126 PD=1.14 PS=1.14 NRD=2.3443 NRS=2.3443 M=1 R=5.6
+ SA=75001.2 SB=75000.7 A=0.126 P=1.98 MULT=1
MM1029 N_A_1162_48#_M1026_d N_D_N_M1029_g N_VPWR_M1029_s VPB PSHORT L=0.15
+ W=0.84 AD=0.126 AS=0.2478 PD=1.14 PS=2.27 NRD=2.3443 NRS=2.3443 M=1 R=5.6
+ SA=75001.6 SB=75000.2 A=0.126 P=1.98 MULT=1
DX38_noxref VNB VPB NWDIODE A=21.8297 P=26.75
*
.include "sky130_fd_sc_hs__nor4bb_4.pxi.spice"
*
.ends
*
*
