* File: sky130_fd_sc_hs__nand2_8.pex.spice
* Created: Tue Sep  1 20:08:48 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HS__NAND2_8%B 1 3 4 5 6 8 9 11 13 14 16 18 19 21 22 24
+ 25 27 30 34 38 40 41 42 44 45 47 49 50 51 52 53 54 55 56 57
c135 38 0 2.0568e-19 $X=3.855 $Y=0.74
r136 76 77 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.765
+ $Y=1.515 $X2=3.765 $Y2=1.515
r137 71 72 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.595
+ $Y=1.515 $X2=2.595 $Y2=1.515
r138 69 71 1.93834 $w=3.73e-07 $l=1.5e-08 $layer=POLY_cond $X=2.58 $Y=1.475
+ $X2=2.595 $Y2=1.475
r139 68 72 10.3184 $w=4.28e-07 $l=3.85e-07 $layer=LI1_cond $X=2.21 $Y=1.565
+ $X2=2.595 $Y2=1.565
r140 67 69 47.8123 $w=3.73e-07 $l=3.7e-07 $layer=POLY_cond $X=2.21 $Y=1.475
+ $X2=2.58 $Y2=1.475
r141 67 68 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.21
+ $Y=1.515 $X2=2.21 $Y2=1.515
r142 65 67 0.646113 $w=3.73e-07 $l=5e-09 $layer=POLY_cond $X=2.205 $Y=1.475
+ $X2=2.21 $Y2=1.475
r143 64 65 16.1528 $w=3.73e-07 $l=1.25e-07 $layer=POLY_cond $X=2.08 $Y=1.475
+ $X2=2.205 $Y2=1.475
r144 57 77 8.44232 $w=4.28e-07 $l=3.15e-07 $layer=LI1_cond $X=4.08 $Y=1.565
+ $X2=3.765 $Y2=1.565
r145 56 77 4.42216 $w=4.28e-07 $l=1.65e-07 $layer=LI1_cond $X=3.6 $Y=1.565
+ $X2=3.765 $Y2=1.565
r146 55 56 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=3.12 $Y=1.565
+ $X2=3.6 $Y2=1.565
r147 54 55 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=2.64 $Y=1.565
+ $X2=3.12 $Y2=1.565
r148 54 72 1.20605 $w=4.28e-07 $l=4.5e-08 $layer=LI1_cond $X=2.64 $Y=1.565
+ $X2=2.595 $Y2=1.565
r149 53 68 1.34005 $w=4.28e-07 $l=5e-08 $layer=LI1_cond $X=2.16 $Y=1.565
+ $X2=2.21 $Y2=1.565
r150 47 49 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=4.77 $Y=1.765
+ $X2=4.77 $Y2=2.4
r151 46 52 20.4101 $w=1.5e-07 $l=9.94987e-08 $layer=POLY_cond $X=4.41 $Y=1.65
+ $X2=4.32 $Y2=1.67
r152 45 47 26.9307 $w=1.5e-07 $l=1.53542e-07 $layer=POLY_cond $X=4.68 $Y=1.65
+ $X2=4.77 $Y2=1.765
r153 45 46 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=4.68 $Y=1.65
+ $X2=4.41 $Y2=1.65
r154 42 52 5.30422 $w=1.5e-07 $l=9.5e-08 $layer=POLY_cond $X=4.32 $Y=1.765
+ $X2=4.32 $Y2=1.67
r155 42 44 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=4.32 $Y=1.765
+ $X2=4.32 $Y2=2.4
r156 40 52 20.4101 $w=1.5e-07 $l=9.94987e-08 $layer=POLY_cond $X=4.23 $Y=1.65
+ $X2=4.32 $Y2=1.67
r157 40 41 153.83 $w=1.5e-07 $l=3e-07 $layer=POLY_cond $X=4.23 $Y=1.65 $X2=3.93
+ $Y2=1.65
r158 36 41 27.4728 $w=3.73e-07 $l=2.09165e-07 $layer=POLY_cond $X=3.855 $Y=1.475
+ $X2=3.93 $Y2=1.65
r159 36 76 11.63 $w=3.73e-07 $l=9e-08 $layer=POLY_cond $X=3.855 $Y=1.475
+ $X2=3.765 $Y2=1.475
r160 36 38 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=3.855 $Y=1.35
+ $X2=3.855 $Y2=0.74
r161 32 76 43.9357 $w=3.73e-07 $l=3.4e-07 $layer=POLY_cond $X=3.425 $Y=1.475
+ $X2=3.765 $Y2=1.475
r162 32 34 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=3.425 $Y=1.35
+ $X2=3.425 $Y2=0.74
r163 28 32 60.7346 $w=3.73e-07 $l=4.7e-07 $layer=POLY_cond $X=2.955 $Y=1.475
+ $X2=3.425 $Y2=1.475
r164 28 71 46.5201 $w=3.73e-07 $l=3.6e-07 $layer=POLY_cond $X=2.955 $Y=1.475
+ $X2=2.595 $Y2=1.475
r165 28 30 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.955 $Y=1.35
+ $X2=2.955 $Y2=0.74
r166 25 69 24.162 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=2.58 $Y=1.765
+ $X2=2.58 $Y2=1.475
r167 25 27 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.58 $Y=1.765
+ $X2=2.58 $Y2=2.4
r168 22 65 24.162 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=2.205 $Y=1.185
+ $X2=2.205 $Y2=1.475
r169 22 24 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=2.205 $Y=1.185
+ $X2=2.205 $Y2=0.74
r170 19 64 24.162 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=2.08 $Y=1.765
+ $X2=2.08 $Y2=1.475
r171 19 21 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.08 $Y=1.765
+ $X2=2.08 $Y2=2.4
r172 16 64 39.4129 $w=3.73e-07 $l=4.25999e-07 $layer=POLY_cond $X=1.775 $Y=1.185
+ $X2=2.08 $Y2=1.475
r173 16 18 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=1.775 $Y=1.185
+ $X2=1.775 $Y2=0.74
r174 15 51 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.42 $Y=1.26
+ $X2=1.345 $Y2=1.26
r175 14 16 27.4728 $w=3.73e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.7 $Y=1.26
+ $X2=1.775 $Y2=1.185
r176 14 15 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=1.7 $Y=1.26
+ $X2=1.42 $Y2=1.26
r177 11 51 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.345 $Y=1.185
+ $X2=1.345 $Y2=1.26
r178 11 13 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=1.345 $Y=1.185
+ $X2=1.345 $Y2=0.74
r179 10 50 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.99 $Y=1.26
+ $X2=0.915 $Y2=1.26
r180 9 51 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.27 $Y=1.26
+ $X2=1.345 $Y2=1.26
r181 9 10 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=1.27 $Y=1.26
+ $X2=0.99 $Y2=1.26
r182 6 50 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.915 $Y=1.185
+ $X2=0.915 $Y2=1.26
r183 6 8 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=0.915 $Y=1.185
+ $X2=0.915 $Y2=0.74
r184 4 50 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.84 $Y=1.26
+ $X2=0.915 $Y2=1.26
r185 4 5 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=0.84 $Y=1.26 $X2=0.56
+ $Y2=1.26
r186 1 5 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.485 $Y=1.185
+ $X2=0.56 $Y2=1.26
r187 1 3 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=0.485 $Y=1.185
+ $X2=0.485 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HS__NAND2_8%A 1 3 4 5 6 8 9 11 13 14 16 17 19 20 22 23
+ 25 26 28 29 31 32 34 35 37 38 40 41 47 48 49 54 55 77 79 89 93
c118 38 0 1.52276e-19 $X=7.66 $Y=1.765
c119 29 0 1.52276e-19 $X=7.21 $Y=1.765
r120 79 93 0.961134 $w=5.58e-07 $l=4.5e-08 $layer=LI1_cond $X=6.525 $Y=1.5
+ $X2=6.48 $Y2=1.5
r121 77 78 0.533186 $w=4.52e-07 $l=5e-09 $layer=POLY_cond $X=7.655 $Y=1.492
+ $X2=7.66 $Y2=1.492
r122 75 77 28.2589 $w=4.52e-07 $l=2.65e-07 $layer=POLY_cond $X=7.39 $Y=1.492
+ $X2=7.655 $Y2=1.492
r123 75 76 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.39
+ $Y=1.385 $X2=7.39 $Y2=1.385
r124 73 75 17.5951 $w=4.52e-07 $l=1.65e-07 $layer=POLY_cond $X=7.225 $Y=1.492
+ $X2=7.39 $Y2=1.492
r125 72 73 1.59956 $w=4.52e-07 $l=1.5e-08 $layer=POLY_cond $X=7.21 $Y=1.492
+ $X2=7.225 $Y2=1.492
r126 70 71 6.78005 $w=3.91e-07 $l=5.5e-08 $layer=POLY_cond $X=6.38 $Y=1.475
+ $X2=6.435 $Y2=1.475
r127 68 70 1.23274 $w=3.91e-07 $l=1e-08 $layer=POLY_cond $X=6.37 $Y=1.475
+ $X2=6.38 $Y2=1.475
r128 68 69 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.37
+ $Y=1.385 $X2=6.37 $Y2=1.385
r129 66 69 7.2619 $w=5.58e-07 $l=3.4e-07 $layer=LI1_cond $X=6.03 $Y=1.5 $X2=6.37
+ $Y2=1.5
r130 66 89 3.38932 $w=5.58e-07 $l=6.5e-08 $layer=LI1_cond $X=6.03 $Y=1.5
+ $X2=5.965 $Y2=1.5
r131 65 68 41.913 $w=3.91e-07 $l=3.4e-07 $layer=POLY_cond $X=6.03 $Y=1.475
+ $X2=6.37 $Y2=1.475
r132 65 66 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=6.03
+ $Y=1.385 $X2=6.03 $Y2=1.385
r133 63 65 3.08184 $w=3.91e-07 $l=2.5e-08 $layer=POLY_cond $X=6.005 $Y=1.475
+ $X2=6.03 $Y2=1.475
r134 62 63 15.4092 $w=3.91e-07 $l=1.25e-07 $layer=POLY_cond $X=5.88 $Y=1.475
+ $X2=6.005 $Y2=1.475
r135 61 62 37.5985 $w=3.91e-07 $l=3.05e-07 $layer=POLY_cond $X=5.575 $Y=1.475
+ $X2=5.88 $Y2=1.475
r136 58 76 7.2619 $w=5.58e-07 $l=3.4e-07 $layer=LI1_cond $X=7.05 $Y=1.5 $X2=7.39
+ $Y2=1.5
r137 57 58 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=7.05
+ $Y=1.385 $X2=7.05 $Y2=1.385
r138 55 71 10.5587 $w=3.91e-07 $l=1.21861e-07 $layer=POLY_cond $X=6.51 $Y=1.385
+ $X2=6.435 $Y2=1.475
r139 55 57 94.4251 $w=3.3e-07 $l=5.4e-07 $layer=POLY_cond $X=6.51 $Y=1.385
+ $X2=7.05 $Y2=1.385
r140 54 72 13.1977 $w=4.52e-07 $l=1.45186e-07 $layer=POLY_cond $X=7.12 $Y=1.385
+ $X2=7.21 $Y2=1.492
r141 54 57 12.2403 $w=3.3e-07 $l=7e-08 $layer=POLY_cond $X=7.12 $Y=1.385
+ $X2=7.05 $Y2=1.385
r142 49 76 1.06793 $w=5.58e-07 $l=5e-08 $layer=LI1_cond $X=7.44 $Y=1.5 $X2=7.39
+ $Y2=1.5
r143 48 58 1.92227 $w=5.58e-07 $l=9e-08 $layer=LI1_cond $X=6.96 $Y=1.5 $X2=7.05
+ $Y2=1.5
r144 47 93 0.427171 $w=5.58e-07 $l=2e-08 $layer=LI1_cond $X=6.46 $Y=1.5 $X2=6.48
+ $Y2=1.5
r145 47 69 1.92227 $w=5.58e-07 $l=9e-08 $layer=LI1_cond $X=6.46 $Y=1.5 $X2=6.37
+ $Y2=1.5
r146 47 48 8.8638 $w=5.58e-07 $l=4.15e-07 $layer=LI1_cond $X=6.545 $Y=1.5
+ $X2=6.96 $Y2=1.5
r147 47 79 0.427171 $w=5.58e-07 $l=2e-08 $layer=LI1_cond $X=6.545 $Y=1.5
+ $X2=6.525 $Y2=1.5
r148 45 61 27.7366 $w=3.91e-07 $l=2.25e-07 $layer=POLY_cond $X=5.35 $Y=1.475
+ $X2=5.575 $Y2=1.475
r149 44 89 21.4773 $w=3.28e-07 $l=6.15e-07 $layer=LI1_cond $X=5.35 $Y=1.385
+ $X2=5.965 $Y2=1.385
r150 44 45 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=5.35
+ $Y=1.385 $X2=5.35 $Y2=1.385
r151 38 78 28.877 $w=1.5e-07 $l=2.73e-07 $layer=POLY_cond $X=7.66 $Y=1.765
+ $X2=7.66 $Y2=1.492
r152 38 40 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=7.66 $Y=1.765
+ $X2=7.66 $Y2=2.4
r153 35 77 28.877 $w=1.5e-07 $l=2.72e-07 $layer=POLY_cond $X=7.655 $Y=1.22
+ $X2=7.655 $Y2=1.492
r154 35 37 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=7.655 $Y=1.22
+ $X2=7.655 $Y2=0.74
r155 32 73 28.877 $w=1.5e-07 $l=2.72e-07 $layer=POLY_cond $X=7.225 $Y=1.22
+ $X2=7.225 $Y2=1.492
r156 32 34 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=7.225 $Y=1.22
+ $X2=7.225 $Y2=0.74
r157 29 72 28.877 $w=1.5e-07 $l=2.73e-07 $layer=POLY_cond $X=7.21 $Y=1.765
+ $X2=7.21 $Y2=1.492
r158 29 31 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=7.21 $Y=1.765
+ $X2=7.21 $Y2=2.4
r159 26 71 25.3065 $w=1.5e-07 $l=2.55e-07 $layer=POLY_cond $X=6.435 $Y=1.22
+ $X2=6.435 $Y2=1.475
r160 26 28 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=6.435 $Y=1.22
+ $X2=6.435 $Y2=0.74
r161 23 70 25.3065 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=6.38 $Y=1.765
+ $X2=6.38 $Y2=1.475
r162 23 25 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=6.38 $Y=1.765
+ $X2=6.38 $Y2=2.4
r163 20 63 25.3065 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=6.005 $Y=1.185
+ $X2=6.005 $Y2=1.475
r164 20 22 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=6.005 $Y=1.185
+ $X2=6.005 $Y2=0.74
r165 17 62 25.3065 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=5.88 $Y=1.765
+ $X2=5.88 $Y2=1.475
r166 17 19 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=5.88 $Y=1.765
+ $X2=5.88 $Y2=2.4
r167 14 61 25.3065 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=5.575 $Y=1.185
+ $X2=5.575 $Y2=1.475
r168 14 16 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=5.575 $Y=1.185
+ $X2=5.575 $Y2=0.74
r169 11 45 25.2711 $w=3.91e-07 $l=3.7888e-07 $layer=POLY_cond $X=5.145 $Y=1.185
+ $X2=5.35 $Y2=1.475
r170 11 13 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=5.145 $Y=1.185
+ $X2=5.145 $Y2=0.74
r171 10 41 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.79 $Y=1.26
+ $X2=4.715 $Y2=1.26
r172 9 11 28.3191 $w=3.91e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.07 $Y=1.26
+ $X2=5.145 $Y2=1.185
r173 9 10 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=5.07 $Y=1.26
+ $X2=4.79 $Y2=1.26
r174 6 41 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.715 $Y=1.185
+ $X2=4.715 $Y2=1.26
r175 6 8 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=4.715 $Y=1.185
+ $X2=4.715 $Y2=0.74
r176 4 41 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.64 $Y=1.26
+ $X2=4.715 $Y2=1.26
r177 4 5 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=4.64 $Y=1.26 $X2=4.36
+ $Y2=1.26
r178 1 5 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.285 $Y=1.185
+ $X2=4.36 $Y2=1.26
r179 1 3 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=4.285 $Y=1.185
+ $X2=4.285 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HS__NAND2_8%VPWR 1 2 3 4 5 6 25 29 33 37 41 43 45 47 49
+ 54 60 68 76 87 89 92 95 101
r81 100 101 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r82 96 98 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=6.48 $Y2=3.33
r83 95 98 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r84 95 96 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r85 93 98 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=6.48 $Y2=3.33
r86 92 93 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r87 90 93 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=5.52 $Y2=3.33
r88 89 90 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r89 86 87 13.0375 $w=1.123e-06 $l=1.2e-07 $layer=LI1_cond $X=4.09 $Y=2.852
+ $X2=4.21 $Y2=2.852
r90 83 86 0.108444 $w=1.123e-06 $l=1e-08 $layer=LI1_cond $X=4.08 $Y=2.852
+ $X2=4.09 $Y2=2.852
r91 80 83 10.4107 $w=1.123e-06 $l=9.6e-07 $layer=LI1_cond $X=3.12 $Y=2.852
+ $X2=4.08 $Y2=2.852
r92 80 81 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r93 78 80 3.416 $w=1.123e-06 $l=3.15e-07 $layer=LI1_cond $X=2.805 $Y=2.852
+ $X2=3.12 $Y2=2.852
r94 75 81 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r95 74 78 1.78933 $w=1.123e-06 $l=1.65e-07 $layer=LI1_cond $X=2.64 $Y=2.852
+ $X2=2.805 $Y2=2.852
r96 74 76 11.7362 $w=1.123e-06 $l=3.8602e-08 $layer=LI1_cond $X=2.64 $Y=2.852
+ $X2=2.64 $Y2=2.852
r97 74 75 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r98 71 75 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.64 $Y2=3.33
r99 69 71 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.68 $Y2=3.33
r100 68 71 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r101 68 69 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r102 66 68 4.79618 $w=1.308e-06 $l=5.15e-07 $layer=LI1_cond $X=1.315 $Y=2.815
+ $X2=1.315 $Y2=3.33
r103 63 66 3.25954 $w=1.308e-06 $l=3.5e-07 $layer=LI1_cond $X=1.315 $Y=2.465
+ $X2=1.315 $Y2=2.815
r104 60 63 3.25954 $w=1.308e-06 $l=3.5e-07 $layer=LI1_cond $X=1.315 $Y=2.115
+ $X2=1.315 $Y2=2.465
r105 58 101 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=7.92 $Y2=3.33
r106 58 96 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=6.96 $Y2=3.33
r107 57 58 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r108 55 95 13.764 $w=1.7e-07 $l=3.55e-07 $layer=LI1_cond $X=7.15 $Y=3.33
+ $X2=6.795 $Y2=3.33
r109 55 57 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=7.15 $Y=3.33
+ $X2=7.44 $Y2=3.33
r110 54 100 4.746 $w=1.7e-07 $l=2.2e-07 $layer=LI1_cond $X=7.72 $Y=3.33 $X2=7.94
+ $Y2=3.33
r111 54 57 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=7.72 $Y=3.33
+ $X2=7.44 $Y2=3.33
r112 53 90 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=5.04 $Y2=3.33
r113 52 87 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=4.56 $Y=3.33
+ $X2=4.21 $Y2=3.33
r114 52 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r115 49 89 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.88 $Y=3.33
+ $X2=5.045 $Y2=3.33
r116 49 52 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=4.88 $Y=3.33
+ $X2=4.56 $Y2=3.33
r117 47 53 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=4.56 $Y2=3.33
r118 47 81 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=3.12 $Y2=3.33
r119 47 83 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r120 43 100 3.02018 $w=3.3e-07 $l=1.09087e-07 $layer=LI1_cond $X=7.885 $Y=3.245
+ $X2=7.94 $Y2=3.33
r121 43 45 30.3826 $w=3.28e-07 $l=8.7e-07 $layer=LI1_cond $X=7.885 $Y=3.245
+ $X2=7.885 $Y2=2.375
r122 39 95 2.89202 $w=7.1e-07 $l=8.5e-08 $layer=LI1_cond $X=6.795 $Y=3.245
+ $X2=6.795 $Y2=3.33
r123 39 41 14.6562 $w=7.08e-07 $l=8.7e-07 $layer=LI1_cond $X=6.795 $Y=3.245
+ $X2=6.795 $Y2=2.375
r124 38 92 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.77 $Y=3.33
+ $X2=5.605 $Y2=3.33
r125 37 95 13.764 $w=1.7e-07 $l=3.55e-07 $layer=LI1_cond $X=6.44 $Y=3.33
+ $X2=6.795 $Y2=3.33
r126 37 38 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=6.44 $Y=3.33
+ $X2=5.77 $Y2=3.33
r127 33 36 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=5.605 $Y=1.985
+ $X2=5.605 $Y2=2.815
r128 31 92 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.605 $Y=3.245
+ $X2=5.605 $Y2=3.33
r129 31 36 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=5.605 $Y=3.245
+ $X2=5.605 $Y2=2.815
r130 30 89 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.21 $Y=3.33
+ $X2=5.045 $Y2=3.33
r131 29 92 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.44 $Y=3.33
+ $X2=5.605 $Y2=3.33
r132 29 30 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=5.44 $Y=3.33
+ $X2=5.21 $Y2=3.33
r133 25 28 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=5.045 $Y=1.985
+ $X2=5.045 $Y2=2.815
r134 23 89 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.045 $Y=3.245
+ $X2=5.045 $Y2=3.33
r135 23 28 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=5.045 $Y=3.245
+ $X2=5.045 $Y2=2.815
r136 22 68 13.6074 $w=1.7e-07 $l=6.55e-07 $layer=LI1_cond $X=1.97 $Y=3.33
+ $X2=1.315 $Y2=3.33
r137 22 76 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.97 $Y=3.33
+ $X2=2.64 $Y2=3.33
r138 6 45 300 $w=1.7e-07 $l=6.05372e-07 $layer=licon1_PDIFF $count=2 $X=7.735
+ $Y=1.84 $X2=7.885 $Y2=2.375
r139 5 41 150 $w=1.7e-07 $l=7.54834e-07 $layer=licon1_PDIFF $count=4 $X=6.455
+ $Y=1.84 $X2=6.985 $Y2=2.375
r140 4 36 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=5.46
+ $Y=1.84 $X2=5.605 $Y2=2.815
r141 4 33 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=5.46
+ $Y=1.84 $X2=5.605 $Y2=1.985
r142 3 28 400 $w=1.7e-07 $l=1.07034e-06 $layer=licon1_PDIFF $count=1 $X=4.845
+ $Y=1.84 $X2=5.045 $Y2=2.815
r143 3 25 400 $w=1.7e-07 $l=2.62678e-07 $layer=licon1_PDIFF $count=1 $X=4.845
+ $Y=1.84 $X2=5.045 $Y2=1.985
r144 2 86 150 $w=1.7e-07 $l=1.71515e-06 $layer=licon1_PDIFF $count=4 $X=2.655
+ $Y=1.84 $X2=4.09 $Y2=2.455
r145 2 78 150 $w=1.7e-07 $l=6.85912e-07 $layer=licon1_PDIFF $count=4 $X=2.655
+ $Y=1.84 $X2=2.805 $Y2=2.455
r146 1 66 200 $w=1.7e-07 $l=1.19718e-06 $layer=licon1_PDIFF $count=3 $X=0.67
+ $Y=1.84 $X2=1.165 $Y2=2.815
r147 1 63 200 $w=1.7e-07 $l=1.45942e-06 $layer=licon1_PDIFF $count=3 $X=0.67
+ $Y=1.84 $X2=1.85 $Y2=2.465
r148 1 63 200 $w=1.7e-07 $l=6.98212e-07 $layer=licon1_PDIFF $count=3 $X=0.67
+ $Y=1.84 $X2=0.825 $Y2=2.465
r149 1 60 200 $w=1.7e-07 $l=6.17373e-07 $layer=licon1_PDIFF $count=3 $X=0.67
+ $Y=1.84 $X2=1.165 $Y2=2.115
.ends

.subckt PM_SKY130_FD_SC_HS__NAND2_8%Y 1 2 3 4 5 6 7 8 25 27 29 33 35 43 45 47 51
+ 53 56 59 64 68 69
c109 59 0 4.40404e-20 $X=4.545 $Y=1.13
c110 51 0 3.04552e-19 $X=7.435 $Y=2.425
r111 62 69 22.8742 $w=3.28e-07 $l=6.55e-07 $layer=LI1_cond $X=4.545 $Y=1.95
+ $X2=4.545 $Y2=1.295
r112 62 64 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.545 $Y=1.95
+ $X2=4.545 $Y2=2.035
r113 59 69 5.76222 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=4.545 $Y=1.13
+ $X2=4.545 $Y2=1.295
r114 59 61 3.23869 $w=3.3e-07 $l=1.91154e-07 $layer=LI1_cond $X=4.545 $Y=1.13
+ $X2=4.522 $Y2=0.95
r115 55 56 58.7166 $w=1.68e-07 $l=9e-07 $layer=LI1_cond $X=7.81 $Y=1.05 $X2=7.81
+ $Y2=1.95
r116 54 68 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=7.55 $Y=2.035
+ $X2=7.435 $Y2=2.035
r117 53 56 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.725 $Y=2.035
+ $X2=7.81 $Y2=1.95
r118 53 54 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=7.725 $Y=2.035
+ $X2=7.55 $Y2=2.035
r119 49 68 0.280307 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.435 $Y=2.12
+ $X2=7.435 $Y2=2.035
r120 49 51 15.2824 $w=2.28e-07 $l=3.05e-07 $layer=LI1_cond $X=7.435 $Y=2.12
+ $X2=7.435 $Y2=2.425
r121 48 66 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.27 $Y=2.035
+ $X2=6.105 $Y2=2.035
r122 47 68 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=7.32 $Y=2.035
+ $X2=7.435 $Y2=2.035
r123 47 48 68.5027 $w=1.68e-07 $l=1.05e-06 $layer=LI1_cond $X=7.32 $Y=2.035
+ $X2=6.27 $Y2=2.035
r124 43 66 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.105 $Y=2.12
+ $X2=6.105 $Y2=2.035
r125 43 45 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=6.105 $Y=2.12
+ $X2=6.105 $Y2=2.425
r126 40 42 50.2136 $w=2.78e-07 $l=1.22e-06 $layer=LI1_cond $X=6.22 $Y=0.91
+ $X2=7.44 $Y2=0.91
r127 38 40 35.3965 $w=2.78e-07 $l=8.6e-07 $layer=LI1_cond $X=5.36 $Y=0.91
+ $X2=6.22 $Y2=0.91
r128 36 61 3.63754 $w=2.8e-07 $l=2.07036e-07 $layer=LI1_cond $X=4.71 $Y=0.91
+ $X2=4.522 $Y2=0.95
r129 36 38 26.7531 $w=2.78e-07 $l=6.5e-07 $layer=LI1_cond $X=4.71 $Y=0.91
+ $X2=5.36 $Y2=0.91
r130 35 55 7.36005 $w=2.8e-07 $l=1.77482e-07 $layer=LI1_cond $X=7.725 $Y=0.91
+ $X2=7.81 $Y2=1.05
r131 35 42 11.7302 $w=2.78e-07 $l=2.85e-07 $layer=LI1_cond $X=7.725 $Y=0.91
+ $X2=7.44 $Y2=0.91
r132 31 64 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.545 $Y=2.12
+ $X2=4.545 $Y2=2.035
r133 31 33 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=4.545 $Y=2.12
+ $X2=4.545 $Y2=2.815
r134 30 58 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.47 $Y=2.035
+ $X2=2.305 $Y2=2.035
r135 29 64 3.80956 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.38 $Y=2.035
+ $X2=4.545 $Y2=2.035
r136 29 30 124.61 $w=1.68e-07 $l=1.91e-06 $layer=LI1_cond $X=4.38 $Y=2.035
+ $X2=2.47 $Y2=2.035
r137 25 58 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.305 $Y=2.12
+ $X2=2.305 $Y2=2.035
r138 25 27 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=2.305 $Y=2.12
+ $X2=2.305 $Y2=2.815
r139 8 68 600 $w=1.7e-07 $l=2.59374e-07 $layer=licon1_PDIFF $count=1 $X=7.285
+ $Y=1.84 $X2=7.435 $Y2=2.035
r140 8 51 300 $w=1.7e-07 $l=6.55725e-07 $layer=licon1_PDIFF $count=2 $X=7.285
+ $Y=1.84 $X2=7.435 $Y2=2.425
r141 7 66 600 $w=1.7e-07 $l=2.59374e-07 $layer=licon1_PDIFF $count=1 $X=5.955
+ $Y=1.84 $X2=6.105 $Y2=2.035
r142 7 45 300 $w=1.7e-07 $l=6.55725e-07 $layer=licon1_PDIFF $count=2 $X=5.955
+ $Y=1.84 $X2=6.105 $Y2=2.425
r143 6 64 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=4.395
+ $Y=1.84 $X2=4.545 $Y2=1.985
r144 6 33 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=4.395
+ $Y=1.84 $X2=4.545 $Y2=2.815
r145 5 58 400 $w=1.7e-07 $l=3.4187e-07 $layer=licon1_PDIFF $count=1 $X=2.155
+ $Y=1.84 $X2=2.305 $Y2=2.115
r146 5 27 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=2.155
+ $Y=1.84 $X2=2.305 $Y2=2.815
r147 4 42 182 $w=1.7e-07 $l=6.0597e-07 $layer=licon1_NDIFF $count=1 $X=7.3
+ $Y=0.37 $X2=7.44 $Y2=0.91
r148 3 40 182 $w=1.7e-07 $l=6.0597e-07 $layer=licon1_NDIFF $count=1 $X=6.08
+ $Y=0.37 $X2=6.22 $Y2=0.91
r149 2 38 182 $w=1.7e-07 $l=6.0597e-07 $layer=licon1_NDIFF $count=1 $X=5.22
+ $Y=0.37 $X2=5.36 $Y2=0.91
r150 1 61 182 $w=1.7e-07 $l=6.4622e-07 $layer=licon1_NDIFF $count=1 $X=4.36
+ $Y=0.37 $X2=4.5 $Y2=0.95
.ends

.subckt PM_SKY130_FD_SC_HS__NAND2_8%A_27_74# 1 2 3 4 5 6 7 8 9 30 32 33 36 38 42
+ 44 45 48 50 52 64 66 68
c104 52 0 1.6164e-19 $X=4.07 $Y=0.6
r105 62 64 39.8745 $w=2.48e-07 $l=8.65e-07 $layer=LI1_cond $X=7.01 $Y=0.475
+ $X2=7.875 $Y2=0.475
r106 60 62 56.2392 $w=2.48e-07 $l=1.22e-06 $layer=LI1_cond $X=5.79 $Y=0.475
+ $X2=7.01 $Y2=0.475
r107 58 60 39.644 $w=2.48e-07 $l=8.6e-07 $layer=LI1_cond $X=4.93 $Y=0.475
+ $X2=5.79 $Y2=0.475
r108 56 70 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.155 $Y=0.475
+ $X2=4.07 $Y2=0.475
r109 56 58 35.7257 $w=2.48e-07 $l=7.75e-07 $layer=LI1_cond $X=4.155 $Y=0.475
+ $X2=4.93 $Y2=0.475
r110 53 55 2.93583 $w=1.68e-07 $l=4.5e-08 $layer=LI1_cond $X=4.07 $Y=1.01
+ $X2=4.07 $Y2=0.965
r111 52 70 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.07 $Y=0.6
+ $X2=4.07 $Y2=0.475
r112 52 55 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=4.07 $Y=0.6
+ $X2=4.07 $Y2=0.965
r113 51 68 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=3.305 $Y=1.095
+ $X2=3.19 $Y2=1.095
r114 50 53 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.985 $Y=1.095
+ $X2=4.07 $Y2=1.01
r115 50 51 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=3.985 $Y=1.095
+ $X2=3.305 $Y2=1.095
r116 46 68 0.280307 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.19 $Y=1.01
+ $X2=3.19 $Y2=1.095
r117 46 48 24.8026 $w=2.28e-07 $l=4.95e-07 $layer=LI1_cond $X=3.19 $Y=1.01
+ $X2=3.19 $Y2=0.515
r118 45 67 7.71193 $w=2.34e-07 $l=1.67183e-07 $layer=LI1_cond $X=2.155 $Y=1.095
+ $X2=2.025 $Y2=1.18
r119 44 68 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=3.075 $Y=1.095
+ $X2=3.19 $Y2=1.095
r120 44 45 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=3.075 $Y=1.095
+ $X2=2.155 $Y2=1.095
r121 40 67 0.0633028 $w=2.6e-07 $l=1.7e-07 $layer=LI1_cond $X=2.025 $Y=1.01
+ $X2=2.025 $Y2=1.18
r122 40 42 21.9407 $w=2.58e-07 $l=4.95e-07 $layer=LI1_cond $X=2.025 $Y=1.01
+ $X2=2.025 $Y2=0.515
r123 39 66 3.85273 $w=2.67e-07 $l=9.5e-08 $layer=LI1_cond $X=1.225 $Y=1.182
+ $X2=1.13 $Y2=1.182
r124 38 67 13.1869 $w=3.45e-07 $l=3.37999e-07 $layer=LI1_cond $X=1.688 $Y=1.182
+ $X2=2.025 $Y2=1.18
r125 38 39 15.4661 $w=3.43e-07 $l=4.63e-07 $layer=LI1_cond $X=1.688 $Y=1.182
+ $X2=1.225 $Y2=1.182
r126 34 66 2.59883 $w=1.9e-07 $l=1.72e-07 $layer=LI1_cond $X=1.13 $Y=1.01
+ $X2=1.13 $Y2=1.182
r127 34 36 28.8947 $w=1.88e-07 $l=4.95e-07 $layer=LI1_cond $X=1.13 $Y=1.01
+ $X2=1.13 $Y2=0.515
r128 32 66 3.85273 $w=2.67e-07 $l=1.28199e-07 $layer=LI1_cond $X=1.035 $Y=1.26
+ $X2=1.13 $Y2=1.182
r129 32 33 39.6938 $w=1.88e-07 $l=6.8e-07 $layer=LI1_cond $X=1.035 $Y=1.26
+ $X2=0.355 $Y2=1.26
r130 28 33 6.98266 $w=1.9e-07 $l=1.65831e-07 $layer=LI1_cond $X=0.23 $Y=1.165
+ $X2=0.355 $Y2=1.26
r131 28 30 29.9635 $w=2.48e-07 $l=6.5e-07 $layer=LI1_cond $X=0.23 $Y=1.165
+ $X2=0.23 $Y2=0.515
r132 9 64 182 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=1 $X=7.73
+ $Y=0.37 $X2=7.875 $Y2=0.515
r133 8 62 91 $w=1.7e-07 $l=5.67891e-07 $layer=licon1_NDIFF $count=2 $X=6.51
+ $Y=0.37 $X2=7.01 $Y2=0.515
r134 7 60 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=5.65
+ $Y=0.37 $X2=5.79 $Y2=0.515
r135 6 58 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=4.79
+ $Y=0.37 $X2=4.93 $Y2=0.515
r136 5 70 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=3.93
+ $Y=0.37 $X2=4.07 $Y2=0.515
r137 5 55 182 $w=1.7e-07 $l=6.61306e-07 $layer=licon1_NDIFF $count=1 $X=3.93
+ $Y=0.37 $X2=4.07 $Y2=0.965
r138 4 48 91 $w=1.7e-07 $l=2.20907e-07 $layer=licon1_NDIFF $count=2 $X=3.03
+ $Y=0.37 $X2=3.19 $Y2=0.515
r139 3 42 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.85
+ $Y=0.37 $X2=1.99 $Y2=0.515
r140 2 36 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=0.99
+ $Y=0.37 $X2=1.13 $Y2=0.515
r141 1 30 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.37 $X2=0.27 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__NAND2_8%VGND 1 2 3 4 15 19 23 27 30 31 32 34 43 47
+ 57 58 61 64 67
r90 67 68 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r91 64 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r92 61 62 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r93 57 58 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=7.92 $Y=0
+ $X2=7.92 $Y2=0
r94 54 57 250.524 $w=1.68e-07 $l=3.84e-06 $layer=LI1_cond $X=4.08 $Y=0 $X2=7.92
+ $Y2=0
r95 52 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.805 $Y=0 $X2=3.64
+ $Y2=0
r96 52 54 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=3.805 $Y=0 $X2=4.08
+ $Y2=0
r97 51 68 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=3.6
+ $Y2=0
r98 51 65 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=2.64
+ $Y2=0
r99 50 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r100 48 64 12.3201 $w=1.7e-07 $l=2.9e-07 $layer=LI1_cond $X=2.905 $Y=0 $X2=2.615
+ $Y2=0
r101 48 50 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=2.905 $Y=0
+ $X2=3.12 $Y2=0
r102 47 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.475 $Y=0 $X2=3.64
+ $Y2=0
r103 47 50 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=3.475 $Y=0
+ $X2=3.12 $Y2=0
r104 46 65 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r105 45 46 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r106 43 64 12.3201 $w=1.7e-07 $l=2.9e-07 $layer=LI1_cond $X=2.325 $Y=0 $X2=2.615
+ $Y2=0
r107 43 45 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=2.325 $Y=0
+ $X2=2.16 $Y2=0
r108 42 46 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r109 42 62 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r110 41 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r111 39 61 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.865 $Y=0 $X2=0.7
+ $Y2=0
r112 39 41 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=0.865 $Y=0 $X2=1.2
+ $Y2=0
r113 37 62 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r114 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r115 34 61 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.535 $Y=0 $X2=0.7
+ $Y2=0
r116 34 36 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.535 $Y=0 $X2=0.24
+ $Y2=0
r117 32 58 1.07034 $w=4.9e-07 $l=3.84e-06 $layer=MET1_cond $X=4.08 $Y=0 $X2=7.92
+ $Y2=0
r118 32 68 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=3.6
+ $Y2=0
r119 32 54 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=4.08 $Y=0
+ $X2=4.08 $Y2=0
r120 30 41 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=1.395 $Y=0 $X2=1.2
+ $Y2=0
r121 30 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.395 $Y=0 $X2=1.56
+ $Y2=0
r122 29 45 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=1.725 $Y=0
+ $X2=2.16 $Y2=0
r123 29 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.725 $Y=0 $X2=1.56
+ $Y2=0
r124 25 67 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.64 $Y=0.085
+ $X2=3.64 $Y2=0
r125 25 27 19.2074 $w=3.28e-07 $l=5.5e-07 $layer=LI1_cond $X=3.64 $Y=0.085
+ $X2=3.64 $Y2=0.635
r126 21 64 2.44113 $w=5.8e-07 $l=8.5e-08 $layer=LI1_cond $X=2.615 $Y=0.085
+ $X2=2.615 $Y2=0
r127 21 23 8.45504 $w=5.78e-07 $l=4.1e-07 $layer=LI1_cond $X=2.615 $Y=0.085
+ $X2=2.615 $Y2=0.495
r128 17 31 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.56 $Y=0.085
+ $X2=1.56 $Y2=0
r129 17 19 20.6043 $w=3.28e-07 $l=5.9e-07 $layer=LI1_cond $X=1.56 $Y=0.085
+ $X2=1.56 $Y2=0.675
r130 13 61 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.7 $Y=0.085 $X2=0.7
+ $Y2=0
r131 13 15 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=0.7 $Y=0.085
+ $X2=0.7 $Y2=0.515
r132 4 27 182 $w=1.7e-07 $l=3.27605e-07 $layer=licon1_NDIFF $count=1 $X=3.5
+ $Y=0.37 $X2=3.64 $Y2=0.635
r133 3 23 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=2.28
+ $Y=0.37 $X2=2.42 $Y2=0.495
r134 2 19 182 $w=1.7e-07 $l=3.68409e-07 $layer=licon1_NDIFF $count=1 $X=1.42
+ $Y=0.37 $X2=1.56 $Y2=0.675
r135 1 15 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=0.56
+ $Y=0.37 $X2=0.7 $Y2=0.515
.ends

