* File: sky130_fd_sc_hs__a21bo_4.pex.spice
* Created: Thu Aug 27 20:24:16 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HS__A21BO_4%B1_N 2 3 5 9 12 14 20
c35 2 0 1.05294e-19 $X=0.495 $Y=1.795
r36 17 20 35.8466 $w=3.3e-07 $l=2.05e-07 $layer=POLY_cond $X=0.46 $Y=0.34
+ $X2=0.665 $Y2=0.34
r37 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.46
+ $Y=0.34 $X2=0.46 $Y2=0.34
r38 14 18 8.25846 $w=3.25e-07 $l=2.2e-07 $layer=LI1_cond $X=0.24 $Y=0.462
+ $X2=0.46 $Y2=0.462
r39 7 12 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.665 $Y=1.33
+ $X2=0.665 $Y2=1.405
r40 7 9 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=0.665 $Y=1.33
+ $X2=0.665 $Y2=0.935
r41 6 20 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.665 $Y=0.505
+ $X2=0.665 $Y2=0.34
r42 6 9 220.489 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=0.665 $Y=0.505
+ $X2=0.665 $Y2=0.935
r43 3 5 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=0.495 $Y=1.885
+ $X2=0.495 $Y2=2.46
r44 2 3 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=0.495 $Y=1.795 $X2=0.495
+ $Y2=1.885
r45 1 12 87.1702 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=0.495 $Y=1.405
+ $X2=0.665 $Y2=1.405
r46 1 2 122.444 $w=1.8e-07 $l=3.15e-07 $layer=POLY_cond $X=0.495 $Y=1.48
+ $X2=0.495 $Y2=1.795
.ends

.subckt PM_SKY130_FD_SC_HS__A21BO_4%A_187_338# 1 2 3 10 12 13 15 16 18 19 21 22
+ 24 25 27 28 30 31 33 34 41 42 46 50 52 53 56 58
c155 56 0 1.44963e-19 $X=4.95 $Y=0.76
c156 31 0 1.44963e-19 $X=2.545 $Y=1.35
c157 19 0 1.47805e-19 $X=1.685 $Y=1.35
r158 70 71 32.6215 $w=3.62e-07 $l=2.45e-07 $layer=POLY_cond $X=2.115 $Y=1.557
+ $X2=2.36 $Y2=1.557
r159 69 70 27.2956 $w=3.62e-07 $l=2.05e-07 $layer=POLY_cond $X=1.91 $Y=1.557
+ $X2=2.115 $Y2=1.557
r160 66 67 29.9586 $w=3.62e-07 $l=2.25e-07 $layer=POLY_cond $X=1.46 $Y=1.557
+ $X2=1.685 $Y2=1.557
r161 65 66 27.2956 $w=3.62e-07 $l=2.05e-07 $layer=POLY_cond $X=1.255 $Y=1.557
+ $X2=1.46 $Y2=1.557
r162 64 65 32.6215 $w=3.62e-07 $l=2.45e-07 $layer=POLY_cond $X=1.01 $Y=1.557
+ $X2=1.255 $Y2=1.557
r163 54 56 16.1342 $w=2.48e-07 $l=3.5e-07 $layer=LI1_cond $X=4.91 $Y=1.11
+ $X2=4.91 $Y2=0.76
r164 52 54 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=4.785 $Y=1.195
+ $X2=4.91 $Y2=1.11
r165 52 53 69.4813 $w=1.68e-07 $l=1.065e-06 $layer=LI1_cond $X=4.785 $Y=1.195
+ $X2=3.72 $Y2=1.195
r166 48 53 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=3.595 $Y=1.195
+ $X2=3.72 $Y2=1.195
r167 48 50 38.4916 $w=2.48e-07 $l=8.35e-07 $layer=LI1_cond $X=3.595 $Y=1.28
+ $X2=3.595 $Y2=2.115
r168 44 48 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=3.25 $Y=1.195
+ $X2=3.595 $Y2=1.195
r169 44 46 12.2229 $w=3.28e-07 $l=3.5e-07 $layer=LI1_cond $X=3.25 $Y=1.11
+ $X2=3.25 $Y2=0.76
r170 43 58 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.755 $Y=1.195
+ $X2=2.67 $Y2=1.195
r171 42 44 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=3.085 $Y=1.195
+ $X2=3.25 $Y2=1.195
r172 42 43 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=3.085 $Y=1.195
+ $X2=2.755 $Y2=1.195
r173 41 73 14.6464 $w=3.62e-07 $l=1.1e-07 $layer=POLY_cond $X=2.435 $Y=1.557
+ $X2=2.545 $Y2=1.557
r174 41 71 9.98619 $w=3.62e-07 $l=7.5e-08 $layer=POLY_cond $X=2.435 $Y=1.557
+ $X2=2.36 $Y2=1.557
r175 40 41 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=2.435
+ $Y=1.515 $X2=2.435 $Y2=1.515
r176 37 69 20.6381 $w=3.62e-07 $l=1.55e-07 $layer=POLY_cond $X=1.755 $Y=1.557
+ $X2=1.91 $Y2=1.557
r177 37 67 9.32044 $w=3.62e-07 $l=7e-08 $layer=POLY_cond $X=1.755 $Y=1.557
+ $X2=1.685 $Y2=1.557
r178 36 40 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=1.755 $Y=1.515
+ $X2=2.435 $Y2=1.515
r179 36 37 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.755
+ $Y=1.515 $X2=1.755 $Y2=1.515
r180 34 58 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=2.67 $Y=1.515
+ $X2=2.67 $Y2=1.195
r181 34 40 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=2.585 $Y=1.515
+ $X2=2.435 $Y2=1.515
r182 31 73 23.4391 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.545 $Y=1.35
+ $X2=2.545 $Y2=1.557
r183 31 33 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=2.545 $Y=1.35
+ $X2=2.545 $Y2=0.87
r184 28 71 23.4391 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=2.36 $Y=1.765
+ $X2=2.36 $Y2=1.557
r185 28 30 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.36 $Y=1.765
+ $X2=2.36 $Y2=2.4
r186 25 70 23.4391 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.115 $Y=1.35
+ $X2=2.115 $Y2=1.557
r187 25 27 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=2.115 $Y=1.35
+ $X2=2.115 $Y2=0.87
r188 22 69 23.4391 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=1.91 $Y=1.765
+ $X2=1.91 $Y2=1.557
r189 22 24 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.91 $Y=1.765
+ $X2=1.91 $Y2=2.4
r190 19 67 23.4391 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.685 $Y=1.35
+ $X2=1.685 $Y2=1.557
r191 19 21 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.685 $Y=1.35
+ $X2=1.685 $Y2=0.87
r192 16 66 23.4391 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=1.46 $Y=1.765
+ $X2=1.46 $Y2=1.557
r193 16 18 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.46 $Y=1.765
+ $X2=1.46 $Y2=2.4
r194 13 65 23.4391 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.255 $Y=1.35
+ $X2=1.255 $Y2=1.557
r195 13 15 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.255 $Y=1.35
+ $X2=1.255 $Y2=0.87
r196 10 64 23.4391 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=1.01 $Y=1.765
+ $X2=1.01 $Y2=1.557
r197 10 12 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.01 $Y=1.765
+ $X2=1.01 $Y2=2.4
r198 3 50 300 $w=1.7e-07 $l=2.17428e-07 $layer=licon1_PDIFF $count=2 $X=3.405
+ $Y=1.96 $X2=3.555 $Y2=2.115
r199 2 56 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=4.81
+ $Y=0.615 $X2=4.95 $Y2=0.76
r200 1 46 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.11
+ $Y=0.615 $X2=3.25 $Y2=0.76
.ends

.subckt PM_SKY130_FD_SC_HS__A21BO_4%A_29_392# 1 2 9 11 13 14 16 19 20 22 26 29
+ 31 34 35 36 39 45 47
c113 20 0 1.88367e-19 $X=3.78 $Y=1.885
r114 42 45 4.76873 $w=4.33e-07 $l=1.8e-07 $layer=LI1_cond $X=0.27 $Y=1.057
+ $X2=0.45 $Y2=1.057
r115 40 50 37.8582 $w=2.61e-07 $l=2.05e-07 $layer=POLY_cond $X=3.125 $Y=1.667
+ $X2=3.33 $Y2=1.667
r116 40 48 16.6207 $w=2.61e-07 $l=9e-08 $layer=POLY_cond $X=3.125 $Y=1.667
+ $X2=3.035 $Y2=1.667
r117 39 40 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.125
+ $Y=1.615 $X2=3.125 $Y2=1.615
r118 37 39 8.20679 $w=3.28e-07 $l=2.35e-07 $layer=LI1_cond $X=3.125 $Y=1.85
+ $X2=3.125 $Y2=1.615
r119 35 37 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.96 $Y=1.935
+ $X2=3.125 $Y2=1.85
r120 35 36 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=2.96 $Y=1.935
+ $X2=2.64 $Y2=1.935
r121 33 36 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.555 $Y=2.02
+ $X2=2.64 $Y2=1.935
r122 33 34 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=2.555 $Y=2.02
+ $X2=2.555 $Y2=2.27
r123 32 47 3.80956 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.435 $Y=2.355
+ $X2=0.27 $Y2=2.355
r124 31 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.47 $Y=2.355
+ $X2=2.555 $Y2=2.27
r125 31 32 132.765 $w=1.68e-07 $l=2.035e-06 $layer=LI1_cond $X=2.47 $Y=2.355
+ $X2=0.435 $Y2=2.355
r126 27 47 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.27 $Y=2.44
+ $X2=0.27 $Y2=2.355
r127 27 29 13.0959 $w=3.28e-07 $l=3.75e-07 $layer=LI1_cond $X=0.27 $Y=2.44
+ $X2=0.27 $Y2=2.815
r128 24 47 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.27 $Y=2.27
+ $X2=0.27 $Y2=2.355
r129 24 26 5.76222 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=0.27 $Y=2.27
+ $X2=0.27 $Y2=2.105
r130 23 42 2.35727 $w=3.3e-07 $l=2.18e-07 $layer=LI1_cond $X=0.27 $Y=1.275
+ $X2=0.27 $Y2=1.057
r131 23 26 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=0.27 $Y=1.275
+ $X2=0.27 $Y2=2.105
r132 20 22 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=3.78 $Y=1.885
+ $X2=3.78 $Y2=2.46
r133 19 20 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=3.78 $Y=1.795
+ $X2=3.78 $Y2=1.885
r134 18 19 75.7984 $w=1.8e-07 $l=1.95e-07 $layer=POLY_cond $X=3.78 $Y=1.6
+ $X2=3.78 $Y2=1.795
r135 14 18 58.1724 $w=2.61e-07 $l=3.82721e-07 $layer=POLY_cond $X=3.465 $Y=1.45
+ $X2=3.78 $Y2=1.6
r136 14 50 24.931 $w=2.61e-07 $l=2.76377e-07 $layer=POLY_cond $X=3.465 $Y=1.45
+ $X2=3.33 $Y2=1.667
r137 14 16 264.074 $w=1.5e-07 $l=5.15e-07 $layer=POLY_cond $X=3.465 $Y=1.45
+ $X2=3.465 $Y2=0.935
r138 11 50 15.717 $w=1.5e-07 $l=2.18e-07 $layer=POLY_cond $X=3.33 $Y=1.885
+ $X2=3.33 $Y2=1.667
r139 11 13 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=3.33 $Y=1.885
+ $X2=3.33 $Y2=2.46
r140 7 48 15.717 $w=1.5e-07 $l=2.17e-07 $layer=POLY_cond $X=3.035 $Y=1.45
+ $X2=3.035 $Y2=1.667
r141 7 9 264.074 $w=1.5e-07 $l=5.15e-07 $layer=POLY_cond $X=3.035 $Y=1.45
+ $X2=3.035 $Y2=0.935
r142 2 29 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=0.145
+ $Y=1.96 $X2=0.27 $Y2=2.815
r143 2 26 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.145
+ $Y=1.96 $X2=0.27 $Y2=2.105
r144 1 45 182 $w=1.7e-07 $l=4.98598e-07 $layer=licon1_NDIFF $count=1 $X=0.325
+ $Y=0.615 $X2=0.45 $Y2=1.055
.ends

.subckt PM_SKY130_FD_SC_HS__A21BO_4%A1 1 3 6 8 10 13 15 16 24
c47 13 0 1.44963e-19 $X=5.165 $Y=0.935
r48 24 25 4.41623 $w=3.82e-07 $l=3.5e-08 $layer=POLY_cond $X=5.13 $Y=1.667
+ $X2=5.165 $Y2=1.667
r49 22 24 47.3168 $w=3.82e-07 $l=3.75e-07 $layer=POLY_cond $X=4.755 $Y=1.667
+ $X2=5.13 $Y2=1.667
r50 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.755
+ $Y=1.615 $X2=4.755 $Y2=1.615
r51 20 22 2.52356 $w=3.82e-07 $l=2e-08 $layer=POLY_cond $X=4.735 $Y=1.667
+ $X2=4.755 $Y2=1.667
r52 19 20 6.93979 $w=3.82e-07 $l=5.5e-08 $layer=POLY_cond $X=4.68 $Y=1.667
+ $X2=4.735 $Y2=1.667
r53 16 23 9.95292 $w=3.28e-07 $l=2.85e-07 $layer=LI1_cond $X=5.04 $Y=1.615
+ $X2=4.755 $Y2=1.615
r54 15 23 6.80989 $w=3.28e-07 $l=1.95e-07 $layer=LI1_cond $X=4.56 $Y=1.615
+ $X2=4.755 $Y2=1.615
r55 11 25 24.74 $w=1.5e-07 $l=2.17e-07 $layer=POLY_cond $X=5.165 $Y=1.45
+ $X2=5.165 $Y2=1.667
r56 11 13 264.074 $w=1.5e-07 $l=5.15e-07 $layer=POLY_cond $X=5.165 $Y=1.45
+ $X2=5.165 $Y2=0.935
r57 8 24 24.74 $w=1.5e-07 $l=2.18e-07 $layer=POLY_cond $X=5.13 $Y=1.885 $X2=5.13
+ $Y2=1.667
r58 8 10 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=5.13 $Y=1.885
+ $X2=5.13 $Y2=2.46
r59 4 20 24.74 $w=1.5e-07 $l=2.17e-07 $layer=POLY_cond $X=4.735 $Y=1.45
+ $X2=4.735 $Y2=1.667
r60 4 6 264.074 $w=1.5e-07 $l=5.15e-07 $layer=POLY_cond $X=4.735 $Y=1.45
+ $X2=4.735 $Y2=0.935
r61 1 19 24.74 $w=1.5e-07 $l=2.18e-07 $layer=POLY_cond $X=4.68 $Y=1.885 $X2=4.68
+ $Y2=1.667
r62 1 3 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=4.68 $Y=1.885
+ $X2=4.68 $Y2=2.46
.ends

.subckt PM_SKY130_FD_SC_HS__A21BO_4%A2 1 2 3 5 9 10 12 13 14 16 20 23 25 29
r73 28 30 45.3519 $w=3.85e-07 $l=1.65e-07 $layer=POLY_cond $X=4.127 $Y=0.34
+ $X2=4.127 $Y2=0.505
r74 28 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.1
+ $Y=0.34 $X2=4.1 $Y2=0.34
r75 25 28 20.2238 $w=3.85e-07 $l=1.4e-07 $layer=POLY_cond $X=4.127 $Y=0.2
+ $X2=4.127 $Y2=0.34
r76 23 29 7.50834 $w=3.28e-07 $l=2.15e-07 $layer=LI1_cond $X=4.1 $Y=0.555
+ $X2=4.1 $Y2=0.34
r77 20 22 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=5.595 $Y=0.935
+ $X2=5.595 $Y2=1.33
r78 17 20 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=5.595 $Y=0.275
+ $X2=5.595 $Y2=0.935
r79 14 16 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=5.58 $Y=1.885
+ $X2=5.58 $Y2=2.46
r80 13 14 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=5.58 $Y=1.795 $X2=5.58
+ $Y2=1.885
r81 12 22 37.1337 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=5.58 $Y=1.42 $X2=5.58
+ $Y2=1.33
r82 12 13 145.766 $w=1.8e-07 $l=3.75e-07 $layer=POLY_cond $X=5.58 $Y=1.42
+ $X2=5.58 $Y2=1.795
r83 11 25 24.9301 $w=1.5e-07 $l=1.93e-07 $layer=POLY_cond $X=4.32 $Y=0.2
+ $X2=4.127 $Y2=0.2
r84 10 17 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.52 $Y=0.2
+ $X2=5.595 $Y2=0.275
r85 10 11 615.319 $w=1.5e-07 $l=1.2e-06 $layer=POLY_cond $X=5.52 $Y=0.2 $X2=4.32
+ $Y2=0.2
r86 9 21 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=4.245 $Y=0.935
+ $X2=4.245 $Y2=1.33
r87 9 30 220.489 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=4.245 $Y=0.935
+ $X2=4.245 $Y2=0.505
r88 3 5 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=4.23 $Y=1.885
+ $X2=4.23 $Y2=2.46
r89 2 3 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=4.23 $Y=1.795 $X2=4.23
+ $Y2=1.885
r90 1 21 37.1337 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=4.23 $Y=1.42 $X2=4.23
+ $Y2=1.33
r91 1 2 145.766 $w=1.8e-07 $l=3.75e-07 $layer=POLY_cond $X=4.23 $Y=1.42 $X2=4.23
+ $Y2=1.795
.ends

.subckt PM_SKY130_FD_SC_HS__A21BO_4%VPWR 1 2 3 4 5 18 22 26 30 34 37 38 40 41 42
+ 44 49 54 70 71 74 77 80
c88 30 0 1.88367e-19 $X=4.455 $Y=2.455
r89 80 81 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r90 77 78 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r91 74 75 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r92 70 71 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r93 68 71 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.04 $Y=3.33 $X2=6
+ $Y2=3.33
r94 67 68 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r95 65 68 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=5.04 $Y2=3.33
r96 64 65 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r97 61 64 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=3.12 $Y=3.33 $X2=4.08
+ $Y2=3.33
r98 59 80 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.75 $Y=3.33
+ $X2=2.585 $Y2=3.33
r99 59 61 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=2.75 $Y=3.33 $X2=3.12
+ $Y2=3.33
r100 58 81 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r101 58 78 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.68 $Y2=3.33
r102 57 58 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r103 55 77 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.85 $Y=3.33
+ $X2=1.685 $Y2=3.33
r104 55 57 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=1.85 $Y=3.33
+ $X2=2.16 $Y2=3.33
r105 54 80 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.42 $Y=3.33
+ $X2=2.585 $Y2=3.33
r106 54 57 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=2.42 $Y=3.33
+ $X2=2.16 $Y2=3.33
r107 53 78 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=1.68 $Y2=3.33
r108 53 75 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r109 52 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r110 50 74 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.95 $Y=3.33
+ $X2=0.785 $Y2=3.33
r111 50 52 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=0.95 $Y=3.33
+ $X2=1.2 $Y2=3.33
r112 49 77 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.52 $Y=3.33
+ $X2=1.685 $Y2=3.33
r113 49 52 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=1.52 $Y=3.33 $X2=1.2
+ $Y2=3.33
r114 47 75 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r115 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r116 44 74 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.62 $Y=3.33
+ $X2=0.785 $Y2=3.33
r117 44 46 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=0.62 $Y=3.33
+ $X2=0.24 $Y2=3.33
r118 42 65 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=4.08 $Y2=3.33
r119 42 81 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=2.64 $Y2=3.33
r120 42 61 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r121 40 67 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=5.27 $Y=3.33
+ $X2=5.04 $Y2=3.33
r122 40 41 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.27 $Y=3.33
+ $X2=5.395 $Y2=3.33
r123 39 70 31.3155 $w=1.68e-07 $l=4.8e-07 $layer=LI1_cond $X=5.52 $Y=3.33 $X2=6
+ $Y2=3.33
r124 39 41 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.52 $Y=3.33
+ $X2=5.395 $Y2=3.33
r125 37 64 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=4.29 $Y=3.33
+ $X2=4.08 $Y2=3.33
r126 37 38 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.29 $Y=3.33
+ $X2=4.415 $Y2=3.33
r127 36 67 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=4.54 $Y=3.33 $X2=5.04
+ $Y2=3.33
r128 36 38 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.54 $Y=3.33
+ $X2=4.415 $Y2=3.33
r129 32 41 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.395 $Y=3.245
+ $X2=5.395 $Y2=3.33
r130 32 34 36.4172 $w=2.48e-07 $l=7.9e-07 $layer=LI1_cond $X=5.395 $Y=3.245
+ $X2=5.395 $Y2=2.455
r131 28 38 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.415 $Y=3.245
+ $X2=4.415 $Y2=3.33
r132 28 30 36.4172 $w=2.48e-07 $l=7.9e-07 $layer=LI1_cond $X=4.415 $Y=3.245
+ $X2=4.415 $Y2=2.455
r133 24 80 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.585 $Y=3.245
+ $X2=2.585 $Y2=3.33
r134 24 26 16.4136 $w=3.28e-07 $l=4.7e-07 $layer=LI1_cond $X=2.585 $Y=3.245
+ $X2=2.585 $Y2=2.775
r135 20 77 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.685 $Y=3.245
+ $X2=1.685 $Y2=3.33
r136 20 22 16.4136 $w=3.28e-07 $l=4.7e-07 $layer=LI1_cond $X=1.685 $Y=3.245
+ $X2=1.685 $Y2=2.775
r137 16 74 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.785 $Y=3.245
+ $X2=0.785 $Y2=3.33
r138 16 18 16.4136 $w=3.28e-07 $l=4.7e-07 $layer=LI1_cond $X=0.785 $Y=3.245
+ $X2=0.785 $Y2=2.775
r139 5 34 300 $w=1.7e-07 $l=5.65044e-07 $layer=licon1_PDIFF $count=2 $X=5.205
+ $Y=1.96 $X2=5.355 $Y2=2.455
r140 4 30 300 $w=1.7e-07 $l=5.65044e-07 $layer=licon1_PDIFF $count=2 $X=4.305
+ $Y=1.96 $X2=4.455 $Y2=2.455
r141 3 26 600 $w=1.7e-07 $l=1.00721e-06 $layer=licon1_PDIFF $count=1 $X=2.435
+ $Y=1.84 $X2=2.585 $Y2=2.775
r142 2 22 600 $w=1.7e-07 $l=1.00721e-06 $layer=licon1_PDIFF $count=1 $X=1.535
+ $Y=1.84 $X2=1.685 $Y2=2.775
r143 1 18 600 $w=1.7e-07 $l=9.16215e-07 $layer=licon1_PDIFF $count=1 $X=0.57
+ $Y=1.96 $X2=0.785 $Y2=2.775
.ends

.subckt PM_SKY130_FD_SC_HS__A21BO_4%X 1 2 3 4 15 18 21 23 27 29 30 31 32
c55 27 0 1.44963e-19 $X=2.33 $Y=0.645
c56 18 0 1.05294e-19 $X=1.335 $Y=1.51
c57 15 0 1.47805e-19 $X=1.47 $Y=0.645
r58 32 38 10.4403 $w=5.88e-07 $l=5.15e-07 $layer=LI1_cond $X=0.72 $Y=1.805
+ $X2=1.235 $Y2=1.805
r59 30 38 0.304088 $w=5.88e-07 $l=1.5e-08 $layer=LI1_cond $X=1.25 $Y=1.805
+ $X2=1.235 $Y2=1.805
r60 30 31 2.31106 $w=4.2e-07 $l=8.5e-08 $layer=LI1_cond $X=1.25 $Y=1.805
+ $X2=1.335 $Y2=1.805
r61 25 27 16.8257 $w=2.48e-07 $l=3.65e-07 $layer=LI1_cond $X=2.29 $Y=1.01
+ $X2=2.29 $Y2=0.645
r62 24 29 2.57001 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=1.555 $Y=1.095
+ $X2=1.402 $Y2=1.095
r63 23 25 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=2.165 $Y=1.095
+ $X2=2.29 $Y2=1.01
r64 23 24 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=2.165 $Y=1.095
+ $X2=1.555 $Y2=1.095
r65 19 31 2.31106 $w=4.2e-07 $l=2.08207e-07 $layer=LI1_cond $X=1.42 $Y=1.975
+ $X2=1.335 $Y2=1.805
r66 19 21 32.9599 $w=2.48e-07 $l=7.15e-07 $layer=LI1_cond $X=1.42 $Y=1.975
+ $X2=2.135 $Y2=1.975
r67 18 31 4.73016 $w=1.7e-07 $l=2.95e-07 $layer=LI1_cond $X=1.335 $Y=1.51
+ $X2=1.335 $Y2=1.805
r68 17 29 3.87901 $w=2.37e-07 $l=1.13666e-07 $layer=LI1_cond $X=1.335 $Y=1.18
+ $X2=1.402 $Y2=1.095
r69 17 18 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=1.335 $Y=1.18
+ $X2=1.335 $Y2=1.51
r70 13 29 3.87901 $w=2.37e-07 $l=8.5e-08 $layer=LI1_cond $X=1.402 $Y=1.01
+ $X2=1.402 $Y2=1.095
r71 13 15 13.7915 $w=3.03e-07 $l=3.65e-07 $layer=LI1_cond $X=1.402 $Y=1.01
+ $X2=1.402 $Y2=0.645
r72 4 21 600 $w=1.7e-07 $l=2.38485e-07 $layer=licon1_PDIFF $count=1 $X=1.985
+ $Y=1.84 $X2=2.135 $Y2=2.015
r73 3 38 600 $w=1.7e-07 $l=2.22711e-07 $layer=licon1_PDIFF $count=1 $X=1.085
+ $Y=1.84 $X2=1.235 $Y2=2
r74 2 27 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.19
+ $Y=0.5 $X2=2.33 $Y2=0.645
r75 1 15 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.33
+ $Y=0.5 $X2=1.47 $Y2=0.645
.ends

.subckt PM_SKY130_FD_SC_HS__A21BO_4%A_596_392# 1 2 3 4 15 17 18 19 22 23 27 29
+ 31 33 38
r71 31 40 2.9222 $w=2.5e-07 $l=9e-08 $layer=LI1_cond $X=5.845 $Y=2.12 $X2=5.845
+ $Y2=2.03
r72 31 33 32.0379 $w=2.48e-07 $l=6.95e-07 $layer=LI1_cond $X=5.845 $Y=2.12
+ $X2=5.845 $Y2=2.815
r73 30 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.07 $Y=2.035
+ $X2=4.905 $Y2=2.035
r74 29 40 4.22096 $w=1.7e-07 $l=1.27475e-07 $layer=LI1_cond $X=5.72 $Y=2.035
+ $X2=5.845 $Y2=2.03
r75 29 30 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=5.72 $Y=2.035
+ $X2=5.07 $Y2=2.035
r76 25 38 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.905 $Y=2.12
+ $X2=4.905 $Y2=2.035
r77 25 27 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=4.905 $Y=2.12
+ $X2=4.905 $Y2=2.815
r78 24 36 3.40825 $w=1.7e-07 $l=8.74643e-08 $layer=LI1_cond $X=4.09 $Y=2.035
+ $X2=4.005 $Y2=2.03
r79 23 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.74 $Y=2.035
+ $X2=4.905 $Y2=2.035
r80 23 24 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=4.74 $Y=2.035
+ $X2=4.09 $Y2=2.035
r81 20 22 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=4.005 $Y=2.905
+ $X2=4.005 $Y2=2.815
r82 19 36 3.40825 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=4.005 $Y=2.12 $X2=4.005
+ $Y2=2.03
r83 19 22 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=4.005 $Y=2.12
+ $X2=4.005 $Y2=2.815
r84 17 20 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.92 $Y=2.99
+ $X2=4.005 $Y2=2.905
r85 17 18 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=3.92 $Y=2.99
+ $X2=3.27 $Y2=2.99
r86 13 18 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.105 $Y=2.905
+ $X2=3.27 $Y2=2.99
r87 13 15 19.2074 $w=3.28e-07 $l=5.5e-07 $layer=LI1_cond $X=3.105 $Y=2.905
+ $X2=3.105 $Y2=2.355
r88 4 40 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=5.655
+ $Y=1.96 $X2=5.805 $Y2=2.105
r89 4 33 400 $w=1.7e-07 $l=9.26971e-07 $layer=licon1_PDIFF $count=1 $X=5.655
+ $Y=1.96 $X2=5.805 $Y2=2.815
r90 3 38 400 $w=1.7e-07 $l=2.17428e-07 $layer=licon1_PDIFF $count=1 $X=4.755
+ $Y=1.96 $X2=4.905 $Y2=2.115
r91 3 27 400 $w=1.7e-07 $l=9.26971e-07 $layer=licon1_PDIFF $count=1 $X=4.755
+ $Y=1.96 $X2=4.905 $Y2=2.815
r92 2 36 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=3.855
+ $Y=1.96 $X2=4.005 $Y2=2.105
r93 2 22 400 $w=1.7e-07 $l=9.26971e-07 $layer=licon1_PDIFF $count=1 $X=3.855
+ $Y=1.96 $X2=4.005 $Y2=2.815
r94 1 15 300 $w=1.7e-07 $l=4.53211e-07 $layer=licon1_PDIFF $count=2 $X=2.98
+ $Y=1.96 $X2=3.105 $Y2=2.355
.ends

.subckt PM_SKY130_FD_SC_HS__A21BO_4%VGND 1 2 3 4 5 18 24 26 30 32 36 38 40 43 44
+ 45 46 47 56 65 68 72
r87 71 72 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=0 $X2=6 $Y2=0
r88 68 69 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r89 65 66 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r90 63 72 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=6
+ $Y2=0
r91 62 63 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r92 60 63 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=4.08 $Y=0 $X2=5.52
+ $Y2=0
r93 60 69 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=3.6
+ $Y2=0
r94 59 62 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=4.08 $Y=0 $X2=5.52
+ $Y2=0
r95 59 60 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r96 57 68 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.765 $Y=0 $X2=3.68
+ $Y2=0
r97 57 59 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=3.765 $Y=0 $X2=4.08
+ $Y2=0
r98 56 71 3.87298 $w=1.7e-07 $l=2.57e-07 $layer=LI1_cond $X=5.725 $Y=0 $X2=5.982
+ $Y2=0
r99 56 62 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=5.725 $Y=0 $X2=5.52
+ $Y2=0
r100 55 66 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.64
+ $Y2=0
r101 54 55 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r102 51 55 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r103 50 51 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r104 47 69 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=3.6
+ $Y2=0
r105 47 66 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=2.64
+ $Y2=0
r106 45 54 3.58824 $w=1.68e-07 $l=5.5e-08 $layer=LI1_cond $X=1.735 $Y=0 $X2=1.68
+ $Y2=0
r107 45 46 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.735 $Y=0 $X2=1.86
+ $Y2=0
r108 43 50 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=0.795 $Y=0 $X2=0.72
+ $Y2=0
r109 43 44 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.795 $Y=0 $X2=0.92
+ $Y2=0
r110 42 54 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=1.045 $Y=0
+ $X2=1.68 $Y2=0
r111 42 44 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.045 $Y=0 $X2=0.92
+ $Y2=0
r112 38 71 3.27018 $w=2.5e-07 $l=1.69245e-07 $layer=LI1_cond $X=5.85 $Y=0.085
+ $X2=5.982 $Y2=0
r113 38 40 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=5.85 $Y=0.085
+ $X2=5.85 $Y2=0.76
r114 34 68 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.68 $Y=0.085
+ $X2=3.68 $Y2=0
r115 34 36 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=3.68 $Y=0.085
+ $X2=3.68 $Y2=0.775
r116 33 65 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.845 $Y=0 $X2=2.72
+ $Y2=0
r117 32 68 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.595 $Y=0 $X2=3.68
+ $Y2=0
r118 32 33 48.9305 $w=1.68e-07 $l=7.5e-07 $layer=LI1_cond $X=3.595 $Y=0
+ $X2=2.845 $Y2=0
r119 28 65 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.72 $Y=0.085
+ $X2=2.72 $Y2=0
r120 28 30 31.8074 $w=2.48e-07 $l=6.9e-07 $layer=LI1_cond $X=2.72 $Y=0.085
+ $X2=2.72 $Y2=0.775
r121 27 46 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.985 $Y=0 $X2=1.86
+ $Y2=0
r122 26 65 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.595 $Y=0 $X2=2.72
+ $Y2=0
r123 26 27 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=2.595 $Y=0
+ $X2=1.985 $Y2=0
r124 22 46 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.86 $Y=0.085
+ $X2=1.86 $Y2=0
r125 22 24 26.5062 $w=2.48e-07 $l=5.75e-07 $layer=LI1_cond $X=1.86 $Y=0.085
+ $X2=1.86 $Y2=0.66
r126 18 20 21.4354 $w=2.48e-07 $l=4.65e-07 $layer=LI1_cond $X=0.92 $Y=0.645
+ $X2=0.92 $Y2=1.11
r127 16 44 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.92 $Y=0.085
+ $X2=0.92 $Y2=0
r128 16 18 25.8147 $w=2.48e-07 $l=5.6e-07 $layer=LI1_cond $X=0.92 $Y=0.085
+ $X2=0.92 $Y2=0.645
r129 5 40 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=5.67
+ $Y=0.615 $X2=5.81 $Y2=0.76
r130 4 36 182 $w=1.7e-07 $l=2.19089e-07 $layer=licon1_NDIFF $count=1 $X=3.54
+ $Y=0.615 $X2=3.68 $Y2=0.775
r131 3 30 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=2.62
+ $Y=0.5 $X2=2.76 $Y2=0.775
r132 2 24 182 $w=1.7e-07 $l=2.19089e-07 $layer=licon1_NDIFF $count=1 $X=1.76
+ $Y=0.5 $X2=1.9 $Y2=0.66
r133 1 20 182 $w=1.7e-07 $l=5.94916e-07 $layer=licon1_NDIFF $count=1 $X=0.74
+ $Y=0.615 $X2=0.96 $Y2=1.11
r134 1 18 182 $w=1.7e-07 $l=2.34521e-07 $layer=licon1_NDIFF $count=1 $X=0.74
+ $Y=0.615 $X2=0.96 $Y2=0.645
.ends

.subckt PM_SKY130_FD_SC_HS__A21BO_4%A_864_123# 1 2 9 11 12 15
r32 13 15 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=5.38 $Y=0.425
+ $X2=5.38 $Y2=0.76
r33 11 13 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=5.215 $Y=0.34
+ $X2=5.38 $Y2=0.425
r34 11 12 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=5.215 $Y=0.34
+ $X2=4.605 $Y2=0.34
r35 7 12 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.52 $Y=0.425
+ $X2=4.605 $Y2=0.34
r36 7 9 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=4.52 $Y=0.425 $X2=4.52
+ $Y2=0.765
r37 2 15 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=5.24
+ $Y=0.615 $X2=5.38 $Y2=0.76
r38 1 9 182 $w=1.7e-07 $l=2.64575e-07 $layer=licon1_NDIFF $count=1 $X=4.32
+ $Y=0.615 $X2=4.52 $Y2=0.765
.ends

