* File: sky130_fd_sc_hs__o31ai_2.pex.spice
* Created: Thu Aug 27 21:03:02 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HS__O31AI_2%A1 3 5 7 8 10 11 13 14 15 16 25
c49 16 0 1.44855e-19 $X=1.2 $Y=1.665
r50 23 25 47.0703 $w=3.84e-07 $l=3.75e-07 $layer=POLY_cond $X=0.585 $Y=1.475
+ $X2=0.96 $Y2=1.475
r51 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.585
+ $Y=1.515 $X2=0.585 $Y2=1.515
r52 21 23 9.41406 $w=3.84e-07 $l=7.5e-08 $layer=POLY_cond $X=0.51 $Y=1.475
+ $X2=0.585 $Y2=1.475
r53 15 16 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=0.72 $Y=1.565
+ $X2=1.2 $Y2=1.565
r54 15 24 3.61813 $w=4.28e-07 $l=1.35e-07 $layer=LI1_cond $X=0.72 $Y=1.565
+ $X2=0.585 $Y2=1.565
r55 14 24 9.24634 $w=4.28e-07 $l=3.45e-07 $layer=LI1_cond $X=0.24 $Y=1.565
+ $X2=0.585 $Y2=1.565
r56 11 25 13.1797 $w=3.84e-07 $l=3.38452e-07 $layer=POLY_cond $X=1.065 $Y=1.185
+ $X2=0.96 $Y2=1.475
r57 11 13 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=1.065 $Y=1.185
+ $X2=1.065 $Y2=0.74
r58 8 25 24.8669 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=0.96 $Y=1.765
+ $X2=0.96 $Y2=1.475
r59 8 10 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.96 $Y=1.765
+ $X2=0.96 $Y2=2.4
r60 5 21 24.8669 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=0.51 $Y=1.765
+ $X2=0.51 $Y2=1.475
r61 5 7 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.51 $Y=1.765
+ $X2=0.51 $Y2=2.4
r62 1 21 1.88281 $w=3.84e-07 $l=1.5e-08 $layer=POLY_cond $X=0.495 $Y=1.475
+ $X2=0.51 $Y2=1.475
r63 1 3 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=0.495 $Y=1.35
+ $X2=0.495 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HS__O31AI_2%A2 1 3 6 8 10 13 15 16 24
c55 24 0 1.15611e-19 $X=1.86 $Y=1.557
c56 16 0 7.40459e-20 $X=2.16 $Y=1.665
c57 13 0 3.67831e-20 $X=2.065 $Y=0.74
c58 1 0 1.44855e-19 $X=1.41 $Y=1.765
r59 22 24 20.0833 $w=3.12e-07 $l=1.3e-07 $layer=POLY_cond $X=1.73 $Y=1.557
+ $X2=1.86 $Y2=1.557
r60 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.73
+ $Y=1.515 $X2=1.73 $Y2=1.515
r61 20 22 36.3045 $w=3.12e-07 $l=2.35e-07 $layer=POLY_cond $X=1.495 $Y=1.557
+ $X2=1.73 $Y2=1.557
r62 16 23 11.5244 $w=4.28e-07 $l=4.3e-07 $layer=LI1_cond $X=2.16 $Y=1.565
+ $X2=1.73 $Y2=1.565
r63 15 23 1.34005 $w=4.28e-07 $l=5e-08 $layer=LI1_cond $X=1.68 $Y=1.565 $X2=1.73
+ $Y2=1.565
r64 11 24 31.6699 $w=3.12e-07 $l=2.92034e-07 $layer=POLY_cond $X=2.065 $Y=1.35
+ $X2=1.86 $Y2=1.557
r65 11 13 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.065 $Y=1.35
+ $X2=2.065 $Y2=0.74
r66 8 24 19.893 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=1.86 $Y=1.765
+ $X2=1.86 $Y2=1.557
r67 8 10 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.86 $Y=1.765
+ $X2=1.86 $Y2=2.4
r68 4 20 19.893 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.495 $Y=1.35
+ $X2=1.495 $Y2=1.557
r69 4 6 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.495 $Y=1.35
+ $X2=1.495 $Y2=0.74
r70 1 20 13.1314 $w=3.12e-07 $l=2.46868e-07 $layer=POLY_cond $X=1.41 $Y=1.765
+ $X2=1.495 $Y2=1.557
r71 1 3 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.41 $Y=1.765
+ $X2=1.41 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_HS__O31AI_2%A3 3 5 6 7 9 10 12 15 17 22 23
c66 10 0 7.53404e-20 $X=3.345 $Y=1.765
c67 7 0 7.40459e-20 $X=2.895 $Y=1.765
r68 23 24 3.19629 $w=3.77e-07 $l=2.5e-08 $layer=POLY_cond $X=3.345 $Y=1.557
+ $X2=3.37 $Y2=1.557
r69 21 23 8.31034 $w=3.77e-07 $l=6.5e-08 $layer=POLY_cond $X=3.28 $Y=1.557
+ $X2=3.345 $Y2=1.557
r70 21 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.28
+ $Y=1.515 $X2=3.28 $Y2=1.515
r71 19 21 49.2228 $w=3.77e-07 $l=3.85e-07 $layer=POLY_cond $X=2.895 $Y=1.557
+ $X2=3.28 $Y2=1.557
r72 17 22 4.28816 $w=4.28e-07 $l=1.6e-07 $layer=LI1_cond $X=3.12 $Y=1.565
+ $X2=3.28 $Y2=1.565
r73 13 24 24.4204 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.37 $Y=1.35
+ $X2=3.37 $Y2=1.557
r74 13 15 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=3.37 $Y=1.35
+ $X2=3.37 $Y2=0.74
r75 10 23 24.4204 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=3.345 $Y=1.765
+ $X2=3.345 $Y2=1.557
r76 10 12 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.345 $Y=1.765
+ $X2=3.345 $Y2=2.4
r77 7 19 24.4204 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=2.895 $Y=1.765
+ $X2=2.895 $Y2=1.557
r78 7 9 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.895 $Y=1.765
+ $X2=2.895 $Y2=2.4
r79 5 19 29.5789 $w=3.77e-07 $l=1.71184e-07 $layer=POLY_cond $X=2.805 $Y=1.425
+ $X2=2.895 $Y2=1.557
r80 5 6 120.5 $w=1.5e-07 $l=2.35e-07 $layer=POLY_cond $X=2.805 $Y=1.425 $X2=2.57
+ $Y2=1.425
r81 1 6 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.495 $Y=1.35
+ $X2=2.57 $Y2=1.425
r82 1 3 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.495 $Y=1.35
+ $X2=2.495 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HS__O31AI_2%B1 3 5 7 10 12 14 15 20 26
c56 15 0 1.34959e-19 $X=4.365 $Y=1.515
r57 29 34 1.74613 $w=3.28e-07 $l=5e-08 $layer=LI1_cond $X=4.53 $Y=1.465 $X2=4.53
+ $Y2=1.515
r58 28 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.53
+ $Y=1.465 $X2=4.53 $Y2=1.465
r59 26 28 28.7487 $w=3.94e-07 $l=2.35e-07 $layer=POLY_cond $X=4.295 $Y=1.532
+ $X2=4.53 $Y2=1.532
r60 25 26 1.83503 $w=3.94e-07 $l=1.5e-08 $layer=POLY_cond $X=4.28 $Y=1.532
+ $X2=4.295 $Y2=1.532
r61 22 23 5.50508 $w=3.94e-07 $l=4.5e-08 $layer=POLY_cond $X=3.8 $Y=1.532
+ $X2=3.845 $Y2=1.532
r62 20 29 5.93683 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=4.53 $Y=1.295
+ $X2=4.53 $Y2=1.465
r63 18 25 11.0102 $w=3.94e-07 $l=9e-08 $layer=POLY_cond $X=4.19 $Y=1.532
+ $X2=4.28 $Y2=1.532
r64 18 23 42.2056 $w=3.94e-07 $l=3.45e-07 $layer=POLY_cond $X=4.19 $Y=1.532
+ $X2=3.845 $Y2=1.532
r65 17 18 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.19
+ $Y=1.515 $X2=4.19 $Y2=1.515
r66 15 34 0.716491 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=4.365 $Y=1.515
+ $X2=4.53 $Y2=1.515
r67 15 17 6.11144 $w=3.28e-07 $l=1.75e-07 $layer=LI1_cond $X=4.365 $Y=1.515
+ $X2=4.19 $Y2=1.515
r68 12 26 25.4929 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=4.295 $Y=1.765
+ $X2=4.295 $Y2=1.532
r69 12 14 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=4.295 $Y=1.765
+ $X2=4.295 $Y2=2.4
r70 8 25 25.4929 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=4.28 $Y=1.3 $X2=4.28
+ $Y2=1.532
r71 8 10 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=4.28 $Y=1.3 $X2=4.28
+ $Y2=0.74
r72 5 23 25.4929 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=3.845 $Y=1.765
+ $X2=3.845 $Y2=1.532
r73 5 7 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.845 $Y=1.765
+ $X2=3.845 $Y2=2.4
r74 1 22 25.4929 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=3.8 $Y=1.3 $X2=3.8
+ $Y2=1.532
r75 1 3 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=3.8 $Y=1.3 $X2=3.8
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HS__O31AI_2%A_28_368# 1 2 3 10 12 14 18 20 27 29
r42 21 27 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.35 $Y=2.035
+ $X2=1.185 $Y2=2.035
r43 20 29 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.92 $Y=2.035
+ $X2=2.085 $Y2=2.035
r44 20 21 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=1.92 $Y=2.035
+ $X2=1.35 $Y2=2.035
r45 16 27 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.185 $Y=2.12
+ $X2=1.185 $Y2=2.035
r46 16 18 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=1.185 $Y=2.12
+ $X2=1.185 $Y2=2.815
r47 15 25 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.37 $Y=2.035
+ $X2=0.245 $Y2=2.035
r48 14 27 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.02 $Y=2.035
+ $X2=1.185 $Y2=2.035
r49 14 15 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=1.02 $Y=2.035
+ $X2=0.37 $Y2=2.035
r50 10 25 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.245 $Y=2.12
+ $X2=0.245 $Y2=2.035
r51 10 12 32.0379 $w=2.48e-07 $l=6.95e-07 $layer=LI1_cond $X=0.245 $Y=2.12
+ $X2=0.245 $Y2=2.815
r52 3 29 300 $w=1.7e-07 $l=3.4187e-07 $layer=licon1_PDIFF $count=2 $X=1.935
+ $Y=1.84 $X2=2.085 $Y2=2.115
r53 2 27 400 $w=1.7e-07 $l=3.4187e-07 $layer=licon1_PDIFF $count=1 $X=1.035
+ $Y=1.84 $X2=1.185 $Y2=2.115
r54 2 18 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=1.035
+ $Y=1.84 $X2=1.185 $Y2=2.815
r55 1 25 400 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_PDIFF $count=1 $X=0.14
+ $Y=1.84 $X2=0.285 $Y2=2.115
r56 1 12 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=0.14
+ $Y=1.84 $X2=0.285 $Y2=2.815
.ends

.subckt PM_SKY130_FD_SC_HS__O31AI_2%VPWR 1 2 9 13 16 17 18 20 33 34 37
r49 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r50 33 34 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r51 31 34 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.56 $Y2=3.33
r52 30 31 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r53 28 38 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r54 27 30 156.578 $w=1.68e-07 $l=2.4e-06 $layer=LI1_cond $X=1.2 $Y=3.33 $X2=3.6
+ $Y2=3.33
r55 27 28 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r56 25 37 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.82 $Y=3.33
+ $X2=0.695 $Y2=3.33
r57 25 27 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=0.82 $Y=3.33 $X2=1.2
+ $Y2=3.33
r58 23 38 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r59 22 23 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r60 20 37 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.57 $Y=3.33
+ $X2=0.695 $Y2=3.33
r61 20 22 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=0.57 $Y=3.33
+ $X2=0.24 $Y2=3.33
r62 18 31 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=2.4 $Y=3.33 $X2=3.6
+ $Y2=3.33
r63 18 28 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=2.4 $Y=3.33 $X2=1.2
+ $Y2=3.33
r64 16 30 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=3.985 $Y=3.33
+ $X2=3.6 $Y2=3.33
r65 16 17 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.985 $Y=3.33
+ $X2=4.07 $Y2=3.33
r66 15 33 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=4.155 $Y=3.33
+ $X2=4.56 $Y2=3.33
r67 15 17 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.155 $Y=3.33
+ $X2=4.07 $Y2=3.33
r68 11 17 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.07 $Y=3.245
+ $X2=4.07 $Y2=3.33
r69 11 13 58.0642 $w=1.68e-07 $l=8.9e-07 $layer=LI1_cond $X=4.07 $Y=3.245
+ $X2=4.07 $Y2=2.355
r70 7 37 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.695 $Y=3.245
+ $X2=0.695 $Y2=3.33
r71 7 9 36.4172 $w=2.48e-07 $l=7.9e-07 $layer=LI1_cond $X=0.695 $Y=3.245
+ $X2=0.695 $Y2=2.455
r72 2 13 300 $w=1.7e-07 $l=5.85214e-07 $layer=licon1_PDIFF $count=2 $X=3.92
+ $Y=1.84 $X2=4.07 $Y2=2.355
r73 1 9 300 $w=1.7e-07 $l=6.85912e-07 $layer=licon1_PDIFF $count=2 $X=0.585
+ $Y=1.84 $X2=0.735 $Y2=2.455
.ends

.subckt PM_SKY130_FD_SC_HS__O31AI_2%A_297_368# 1 2 9 11 12 15
r26 13 15 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=3.12 $Y=2.905
+ $X2=3.12 $Y2=2.455
r27 11 13 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.955 $Y=2.99
+ $X2=3.12 $Y2=2.905
r28 11 12 80.5722 $w=1.68e-07 $l=1.235e-06 $layer=LI1_cond $X=2.955 $Y=2.99
+ $X2=1.72 $Y2=2.99
r29 7 12 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.635 $Y=2.905
+ $X2=1.72 $Y2=2.99
r30 7 9 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=1.635 $Y=2.905
+ $X2=1.635 $Y2=2.455
r31 2 15 300 $w=1.7e-07 $l=6.85912e-07 $layer=licon1_PDIFF $count=2 $X=2.97
+ $Y=1.84 $X2=3.12 $Y2=2.455
r32 1 9 300 $w=1.7e-07 $l=6.85912e-07 $layer=licon1_PDIFF $count=2 $X=1.485
+ $Y=1.84 $X2=1.635 $Y2=2.455
.ends

.subckt PM_SKY130_FD_SC_HS__O31AI_2%Y 1 2 3 4 15 19 20 21 23 27 29 31 34 35 40
+ 43 44
c78 35 0 1.15611e-19 $X=2.67 $Y=1.82
c79 34 0 7.53404e-20 $X=2.67 $Y=1.985
r80 43 44 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=3.62 $Y=2.405
+ $X2=3.62 $Y2=2.775
r81 38 43 9.95292 $w=3.28e-07 $l=2.85e-07 $layer=LI1_cond $X=3.62 $Y=2.12
+ $X2=3.62 $Y2=2.405
r82 38 40 0.89609 $w=3.3e-07 $l=2.38642e-07 $layer=LI1_cond $X=3.62 $Y=2.12
+ $X2=3.455 $Y2=1.95
r83 36 37 3.67308 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=2.67 $Y=2.035
+ $X2=2.67 $Y2=2.12
r84 34 36 1.74613 $w=3.28e-07 $l=5e-08 $layer=LI1_cond $X=2.67 $Y=1.985 $X2=2.67
+ $Y2=2.035
r85 34 35 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=2.67 $Y=1.985
+ $X2=2.67 $Y2=1.82
r86 29 42 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.52 $Y=2.02 $X2=4.52
+ $Y2=1.935
r87 29 31 27.7634 $w=3.28e-07 $l=7.95e-07 $layer=LI1_cond $X=4.52 $Y=2.02
+ $X2=4.52 $Y2=2.815
r88 25 27 8.20679 $w=3.28e-07 $l=2.35e-07 $layer=LI1_cond $X=4.015 $Y=1.01
+ $X2=4.015 $Y2=0.775
r89 24 40 8.61065 $w=1.7e-07 $l=3.37417e-07 $layer=LI1_cond $X=3.785 $Y=1.935
+ $X2=3.455 $Y2=1.95
r90 23 42 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.355 $Y=1.935
+ $X2=4.52 $Y2=1.935
r91 23 24 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=4.355 $Y=1.935
+ $X2=3.785 $Y2=1.935
r92 22 36 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.835 $Y=2.035
+ $X2=2.67 $Y2=2.035
r93 21 40 8.61065 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.455 $Y=2.035
+ $X2=3.455 $Y2=1.95
r94 21 22 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=3.455 $Y=2.035
+ $X2=2.835 $Y2=2.035
r95 19 25 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.85 $Y=1.095
+ $X2=4.015 $Y2=1.01
r96 19 20 66.2193 $w=1.68e-07 $l=1.015e-06 $layer=LI1_cond $X=3.85 $Y=1.095
+ $X2=2.835 $Y2=1.095
r97 17 20 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.75 $Y=1.18
+ $X2=2.835 $Y2=1.095
r98 17 35 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=2.75 $Y=1.18 $X2=2.75
+ $Y2=1.82
r99 15 37 20.744 $w=2.48e-07 $l=4.5e-07 $layer=LI1_cond $X=2.63 $Y=2.57 $X2=2.63
+ $Y2=2.12
r100 4 42 400 $w=1.7e-07 $l=2.38485e-07 $layer=licon1_PDIFF $count=1 $X=4.37
+ $Y=1.84 $X2=4.52 $Y2=2.015
r101 4 31 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=4.37
+ $Y=1.84 $X2=4.52 $Y2=2.815
r102 3 44 400 $w=1.7e-07 $l=1.07034e-06 $layer=licon1_PDIFF $count=1 $X=3.42
+ $Y=1.84 $X2=3.62 $Y2=2.815
r103 3 40 400 $w=1.7e-07 $l=3.61421e-07 $layer=licon1_PDIFF $count=1 $X=3.42
+ $Y=1.84 $X2=3.62 $Y2=2.115
r104 2 34 600 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=2.525
+ $Y=1.84 $X2=2.67 $Y2=1.985
r105 2 15 600 $w=1.7e-07 $l=7.99218e-07 $layer=licon1_PDIFF $count=1 $X=2.525
+ $Y=1.84 $X2=2.67 $Y2=2.57
r106 1 27 182 $w=1.7e-07 $l=4.69814e-07 $layer=licon1_NDIFF $count=1 $X=3.875
+ $Y=0.37 $X2=4.015 $Y2=0.775
.ends

.subckt PM_SKY130_FD_SC_HS__O31AI_2%A_27_74# 1 2 3 4 5 18 20 21 24 26 29 30 35
+ 36 37 40 42 44
c81 30 0 3.67831e-20 $X=3.42 $Y=0.755
r82 44 46 8.3814 $w=3.28e-07 $l=2.4e-07 $layer=LI1_cond $X=2.28 $Y=0.515
+ $X2=2.28 $Y2=0.755
r83 38 40 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=4.515 $Y=0.425
+ $X2=4.515 $Y2=0.515
r84 36 38 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.35 $Y=0.34
+ $X2=4.515 $Y2=0.425
r85 36 37 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=4.35 $Y=0.34
+ $X2=3.67 $Y2=0.34
r86 33 35 3.45733 $w=2.48e-07 $l=7.5e-08 $layer=LI1_cond $X=3.545 $Y=0.67
+ $X2=3.545 $Y2=0.595
r87 32 37 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=3.545 $Y=0.425
+ $X2=3.67 $Y2=0.34
r88 32 35 7.83661 $w=2.48e-07 $l=1.7e-07 $layer=LI1_cond $X=3.545 $Y=0.425
+ $X2=3.545 $Y2=0.595
r89 31 46 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.445 $Y=0.755
+ $X2=2.28 $Y2=0.755
r90 30 33 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=3.42 $Y=0.755
+ $X2=3.545 $Y2=0.67
r91 30 31 63.6096 $w=1.68e-07 $l=9.75e-07 $layer=LI1_cond $X=3.42 $Y=0.755
+ $X2=2.445 $Y2=0.755
r92 28 46 2.96841 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=2.28 $Y=0.84
+ $X2=2.28 $Y2=0.755
r93 28 29 5.93683 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=2.28 $Y=0.84
+ $X2=2.28 $Y2=1.01
r94 27 42 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.445 $Y=1.095
+ $X2=1.28 $Y2=1.095
r95 26 29 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.115 $Y=1.095
+ $X2=2.28 $Y2=1.01
r96 26 27 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.115 $Y=1.095
+ $X2=1.445 $Y2=1.095
r97 22 42 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.28 $Y=1.01 $X2=1.28
+ $Y2=1.095
r98 22 24 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=1.28 $Y=1.01
+ $X2=1.28 $Y2=0.515
r99 20 42 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.115 $Y=1.095
+ $X2=1.28 $Y2=1.095
r100 20 21 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.115 $Y=1.095
+ $X2=0.445 $Y2=1.095
r101 16 21 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.28 $Y=1.01
+ $X2=0.445 $Y2=1.095
r102 16 18 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=0.28 $Y=1.01
+ $X2=0.28 $Y2=0.515
r103 5 40 91 $w=1.7e-07 $l=2.20907e-07 $layer=licon1_NDIFF $count=2 $X=4.355
+ $Y=0.37 $X2=4.515 $Y2=0.515
r104 4 35 182 $w=1.7e-07 $l=2.86575e-07 $layer=licon1_NDIFF $count=1 $X=3.445
+ $Y=0.37 $X2=3.585 $Y2=0.595
r105 3 44 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.14
+ $Y=0.37 $X2=2.28 $Y2=0.515
r106 2 24 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.14
+ $Y=0.37 $X2=1.28 $Y2=0.515
r107 1 18 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__O31AI_2%VGND 1 2 3 12 14 18 22 24 34 35 38 41 46 52
r59 50 52 9.13833 $w=5.83e-07 $l=1.2e-07 $layer=LI1_cond $X=3.12 $Y=0.207
+ $X2=3.24 $Y2=0.207
r60 50 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r61 48 50 3.8847 $w=5.83e-07 $l=1.9e-07 $layer=LI1_cond $X=2.93 $Y=0.207
+ $X2=3.12 $Y2=0.207
r62 45 51 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r63 44 48 5.92928 $w=5.83e-07 $l=2.9e-07 $layer=LI1_cond $X=2.64 $Y=0.207
+ $X2=2.93 $Y2=0.207
r64 44 46 6.99152 $w=5.83e-07 $l=1.5e-08 $layer=LI1_cond $X=2.64 $Y=0.207
+ $X2=2.625 $Y2=0.207
r65 44 45 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r66 41 42 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r67 39 42 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r68 38 39 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r69 34 35 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r70 32 35 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.56
+ $Y2=0
r71 32 51 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=3.12
+ $Y2=0
r72 31 34 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=3.6 $Y=0 $X2=4.56
+ $Y2=0
r73 31 52 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=3.6 $Y=0 $X2=3.24
+ $Y2=0
r74 31 32 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r75 27 39 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r76 26 27 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r77 24 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.615 $Y=0 $X2=0.78
+ $Y2=0
r78 24 26 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=0.615 $Y=0 $X2=0.24
+ $Y2=0
r79 22 45 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.4 $Y=0 $X2=2.64
+ $Y2=0
r80 22 42 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=2.4 $Y=0 $X2=1.68
+ $Y2=0
r81 21 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.945 $Y=0 $X2=1.78
+ $Y2=0
r82 21 46 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.945 $Y=0 $X2=2.625
+ $Y2=0
r83 16 41 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.78 $Y=0.085
+ $X2=1.78 $Y2=0
r84 16 18 20.0804 $w=3.28e-07 $l=5.75e-07 $layer=LI1_cond $X=1.78 $Y=0.085
+ $X2=1.78 $Y2=0.66
r85 15 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.945 $Y=0 $X2=0.78
+ $Y2=0
r86 14 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.615 $Y=0 $X2=1.78
+ $Y2=0
r87 14 15 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.615 $Y=0 $X2=0.945
+ $Y2=0
r88 10 38 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.78 $Y=0.085
+ $X2=0.78 $Y2=0
r89 10 12 20.0804 $w=3.28e-07 $l=5.75e-07 $layer=LI1_cond $X=0.78 $Y=0.085
+ $X2=0.78 $Y2=0.66
r90 3 48 182 $w=1.7e-07 $l=3.77094e-07 $layer=licon1_NDIFF $count=1 $X=2.57
+ $Y=0.37 $X2=2.93 $Y2=0.335
r91 2 18 182 $w=1.7e-07 $l=3.80789e-07 $layer=licon1_NDIFF $count=1 $X=1.57
+ $Y=0.37 $X2=1.78 $Y2=0.66
r92 1 12 182 $w=1.7e-07 $l=3.80789e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.37 $X2=0.78 $Y2=0.66
.ends

