* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hs__a211o_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
X0 a_600_392# C1 a_85_270# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=150000u
X1 a_85_270# B1 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X2 VGND C1 a_85_270# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X3 a_317_392# A2 VPWR VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=150000u
X4 X a_85_270# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X5 a_399_74# A1 a_85_270# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X6 VPWR A1 a_317_392# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=150000u
X7 VGND A2 a_399_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X8 VPWR a_85_270# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X9 X a_85_270# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X10 VGND a_85_270# X VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X11 a_317_392# B1 a_600_392# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=150000u
.ends
