* File: sky130_fd_sc_hs__or4_2.pex.spice
* Created: Thu Aug 27 21:06:44 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HS__OR4_2%D 3 5 7 8
r31 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.59
+ $Y=1.605 $X2=0.59 $Y2=1.605
r32 8 12 8.71359 $w=4.08e-07 $l=3.1e-07 $layer=LI1_cond $X=0.63 $Y=1.295
+ $X2=0.63 $Y2=1.605
r33 5 11 53.9634 $w=3.73e-07 $l=3.42929e-07 $layer=POLY_cond $X=0.795 $Y=1.885
+ $X2=0.655 $Y2=1.605
r34 5 7 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=0.795 $Y=1.885
+ $X2=0.795 $Y2=2.46
r35 1 11 39.1028 $w=3.73e-07 $l=1.72337e-07 $layer=POLY_cond $X=0.64 $Y=1.44
+ $X2=0.655 $Y2=1.605
r36 1 3 384.574 $w=1.5e-07 $l=7.5e-07 $layer=POLY_cond $X=0.64 $Y=1.44 $X2=0.64
+ $Y2=0.69
.ends

.subckt PM_SKY130_FD_SC_HS__OR4_2%C 3 6 7 9 10 11 12 13 19 20
c45 19 0 5.25652e-20 $X=1.17 $Y=1.33
c46 7 0 1.45554e-19 $X=1.215 $Y=1.885
r47 19 22 40.7132 $w=3.4e-07 $l=1.65e-07 $layer=POLY_cond $X=1.165 $Y=1.33
+ $X2=1.165 $Y2=1.495
r48 19 21 46.3065 $w=3.4e-07 $l=1.65e-07 $layer=POLY_cond $X=1.165 $Y=1.33
+ $X2=1.165 $Y2=1.165
r49 19 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.17
+ $Y=1.33 $X2=1.17 $Y2=1.33
r50 12 13 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.17 $Y=2.405
+ $X2=1.17 $Y2=2.775
r51 11 12 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.17 $Y=2.035
+ $X2=1.17 $Y2=2.405
r52 10 11 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.17 $Y=1.665
+ $X2=1.17 $Y2=2.035
r53 10 20 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=1.17 $Y=1.665
+ $X2=1.17 $Y2=1.33
r54 7 9 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=1.215 $Y=1.885
+ $X2=1.215 $Y2=2.46
r55 6 7 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=1.215 $Y=1.795 $X2=1.215
+ $Y2=1.885
r56 6 22 116.613 $w=1.8e-07 $l=3e-07 $layer=POLY_cond $X=1.215 $Y=1.795
+ $X2=1.215 $Y2=1.495
r57 3 21 243.564 $w=1.5e-07 $l=4.75e-07 $layer=POLY_cond $X=1.07 $Y=0.69
+ $X2=1.07 $Y2=1.165
.ends

.subckt PM_SKY130_FD_SC_HS__OR4_2%B 1 3 6 8 9 10 11 18
c36 6 0 1.02301e-19 $X=1.81 $Y=0.69
r37 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.71
+ $Y=1.515 $X2=1.71 $Y2=1.515
r38 10 11 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.71 $Y=2.405
+ $X2=1.71 $Y2=2.775
r39 9 10 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.71 $Y=2.035
+ $X2=1.71 $Y2=2.405
r40 8 9 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.71 $Y=1.665 $X2=1.71
+ $Y2=2.035
r41 8 18 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=1.71 $Y=1.665
+ $X2=1.71 $Y2=1.515
r42 4 17 38.7595 $w=2.78e-07 $l=2.07123e-07 $layer=POLY_cond $X=1.81 $Y=1.35
+ $X2=1.715 $Y2=1.515
r43 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.81 $Y=1.35 $X2=1.81
+ $Y2=0.69
r44 1 17 74.3026 $w=2.78e-07 $l=4.08044e-07 $layer=POLY_cond $X=1.635 $Y=1.885
+ $X2=1.715 $Y2=1.515
r45 1 3 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=1.635 $Y=1.885
+ $X2=1.635 $Y2=2.46
.ends

.subckt PM_SKY130_FD_SC_HS__OR4_2%A 1 3 6 8 12
r33 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.29
+ $Y=1.515 $X2=2.29 $Y2=1.515
r34 8 12 4.21625 $w=4.08e-07 $l=1.5e-07 $layer=LI1_cond $X=2.25 $Y=1.665
+ $X2=2.25 $Y2=1.515
r35 4 11 38.8629 $w=2.72e-07 $l=1.88348e-07 $layer=POLY_cond $X=2.24 $Y=1.35
+ $X2=2.29 $Y2=1.515
r36 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.24 $Y=1.35 $X2=2.24
+ $Y2=0.69
r37 1 11 75.1901 $w=2.72e-07 $l=4.05771e-07 $layer=POLY_cond $X=2.215 $Y=1.885
+ $X2=2.29 $Y2=1.515
r38 1 3 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=2.215 $Y=1.885
+ $X2=2.215 $Y2=2.46
.ends

.subckt PM_SKY130_FD_SC_HS__OR4_2%A_85_392# 1 2 3 10 12 15 17 19 22 25 26 27 30
+ 34 36 40 42 47 49 50 60
c111 50 0 5.25652e-20 $X=2.025 $Y=0.91
c112 47 0 1.45554e-19 $X=0.57 $Y=2.105
c113 42 0 1.02301e-19 $X=2.625 $Y=1.095
r114 59 60 42.7169 $w=3.78e-07 $l=3.35e-07 $layer=POLY_cond $X=2.915 $Y=1.532
+ $X2=3.25 $Y2=1.532
r115 56 59 5.10053 $w=3.78e-07 $l=4e-08 $layer=POLY_cond $X=2.875 $Y=1.532
+ $X2=2.915 $Y2=1.532
r116 56 57 9.56349 $w=3.78e-07 $l=7.5e-08 $layer=POLY_cond $X=2.875 $Y=1.532
+ $X2=2.8 $Y2=1.532
r117 55 56 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.875
+ $Y=1.465 $X2=2.875 $Y2=1.465
r118 50 51 6.46067 $w=3.28e-07 $l=1.85e-07 $layer=LI1_cond $X=2.025 $Y=0.91
+ $X2=2.025 $Y2=1.095
r119 44 47 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=0.17 $Y=2.025
+ $X2=0.57 $Y2=2.025
r120 43 51 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.19 $Y=1.095
+ $X2=2.025 $Y2=1.095
r121 42 55 15.0467 $w=3e-07 $l=4.6205e-07 $layer=LI1_cond $X=2.625 $Y=1.095
+ $X2=2.832 $Y2=1.465
r122 42 43 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=2.625 $Y=1.095
+ $X2=2.19 $Y2=1.095
r123 38 50 2.96841 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=2.025 $Y=0.825
+ $X2=2.025 $Y2=0.91
r124 38 40 10.826 $w=3.28e-07 $l=3.1e-07 $layer=LI1_cond $X=2.025 $Y=0.825
+ $X2=2.025 $Y2=0.515
r125 37 49 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.02 $Y=0.91
+ $X2=0.855 $Y2=0.91
r126 36 50 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.86 $Y=0.91
+ $X2=2.025 $Y2=0.91
r127 36 37 54.8021 $w=1.68e-07 $l=8.4e-07 $layer=LI1_cond $X=1.86 $Y=0.91
+ $X2=1.02 $Y2=0.91
r128 32 49 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.855 $Y=0.825
+ $X2=0.855 $Y2=0.91
r129 32 34 10.826 $w=3.28e-07 $l=3.1e-07 $layer=LI1_cond $X=0.855 $Y=0.825
+ $X2=0.855 $Y2=0.515
r130 30 47 24.6204 $w=3.28e-07 $l=7.05e-07 $layer=LI1_cond $X=0.57 $Y=2.815
+ $X2=0.57 $Y2=2.11
r131 26 49 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.69 $Y=0.91
+ $X2=0.855 $Y2=0.91
r132 26 27 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=0.69 $Y=0.91
+ $X2=0.255 $Y2=0.91
r133 25 44 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.17 $Y=1.94
+ $X2=0.17 $Y2=2.025
r134 24 27 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.17 $Y=0.995
+ $X2=0.255 $Y2=0.91
r135 24 25 61.6524 $w=1.68e-07 $l=9.45e-07 $layer=LI1_cond $X=0.17 $Y=0.995
+ $X2=0.17 $Y2=1.94
r136 20 60 12.1138 $w=3.78e-07 $l=2.75434e-07 $layer=POLY_cond $X=3.345 $Y=1.3
+ $X2=3.25 $Y2=1.532
r137 20 22 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=3.345 $Y=1.3
+ $X2=3.345 $Y2=0.74
r138 17 60 24.4846 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=3.25 $Y=1.765
+ $X2=3.25 $Y2=1.532
r139 17 19 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.25 $Y=1.765
+ $X2=3.25 $Y2=2.4
r140 13 59 24.4846 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=2.915 $Y=1.3
+ $X2=2.915 $Y2=1.532
r141 13 15 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=2.915 $Y=1.3
+ $X2=2.915 $Y2=0.74
r142 10 57 24.4846 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=2.8 $Y=1.765
+ $X2=2.8 $Y2=1.532
r143 10 12 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.8 $Y=1.765
+ $X2=2.8 $Y2=2.4
r144 3 47 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.425
+ $Y=1.96 $X2=0.57 $Y2=2.105
r145 3 30 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=0.425
+ $Y=1.96 $X2=0.57 $Y2=2.815
r146 2 40 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.885
+ $Y=0.37 $X2=2.025 $Y2=0.515
r147 1 34 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=0.715
+ $Y=0.37 $X2=0.855 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__OR4_2%VPWR 1 2 9 13 15 18 19 20 29 35
r38 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r39 32 35 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=3.6 $Y2=3.33
r40 31 32 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r41 29 34 4.65971 $w=1.7e-07 $l=2.4e-07 $layer=LI1_cond $X=3.36 $Y=3.33 $X2=3.6
+ $Y2=3.33
r42 29 31 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=3.36 $Y=3.33
+ $X2=3.12 $Y2=3.33
r43 28 32 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=3.12 $Y2=3.33
r44 27 28 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r45 23 27 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=0.24 $Y=3.33
+ $X2=2.16 $Y2=3.33
r46 23 24 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r47 20 28 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=2.16 $Y2=3.33
r48 20 24 0.468274 $w=4.9e-07 $l=1.68e-06 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=0.24 $Y2=3.33
r49 18 27 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=2.36 $Y=3.33 $X2=2.16
+ $Y2=3.33
r50 18 19 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.36 $Y=3.33
+ $X2=2.525 $Y2=3.33
r51 17 31 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=2.69 $Y=3.33
+ $X2=3.12 $Y2=3.33
r52 17 19 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.69 $Y=3.33
+ $X2=2.525 $Y2=3.33
r53 13 34 3.10647 $w=3.3e-07 $l=1.16619e-07 $layer=LI1_cond $X=3.525 $Y=3.245
+ $X2=3.6 $Y2=3.33
r54 13 15 35.621 $w=3.28e-07 $l=1.02e-06 $layer=LI1_cond $X=3.525 $Y=3.245
+ $X2=3.525 $Y2=2.225
r55 9 12 24.4458 $w=3.28e-07 $l=7e-07 $layer=LI1_cond $X=2.525 $Y=2.115
+ $X2=2.525 $Y2=2.815
r56 7 19 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.525 $Y=3.245
+ $X2=2.525 $Y2=3.33
r57 7 12 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=2.525 $Y=3.245
+ $X2=2.525 $Y2=2.815
r58 2 15 300 $w=1.7e-07 $l=4.74579e-07 $layer=licon1_PDIFF $count=2 $X=3.325
+ $Y=1.84 $X2=3.525 $Y2=2.225
r59 1 12 400 $w=1.7e-07 $l=9.65376e-07 $layer=licon1_PDIFF $count=1 $X=2.29
+ $Y=1.96 $X2=2.525 $Y2=2.815
r60 1 9 400 $w=1.7e-07 $l=3.02738e-07 $layer=licon1_PDIFF $count=1 $X=2.29
+ $Y=1.96 $X2=2.525 $Y2=2.115
.ends

.subckt PM_SKY130_FD_SC_HS__OR4_2%X 1 2 9 15 17 18 19 20 23 24
r41 23 24 18.5393 $w=2.28e-07 $l=3.7e-07 $layer=LI1_cond $X=3.6 $Y=1.295 $X2=3.6
+ $Y2=1.665
r42 22 24 6.76434 $w=2.28e-07 $l=1.35e-07 $layer=LI1_cond $X=3.6 $Y=1.8 $X2=3.6
+ $Y2=1.665
r43 21 23 8.26753 $w=2.28e-07 $l=1.65e-07 $layer=LI1_cond $X=3.6 $Y=1.13 $X2=3.6
+ $Y2=1.295
r44 19 21 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=3.485 $Y=1.045
+ $X2=3.6 $Y2=1.13
r45 19 20 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=3.485 $Y=1.045
+ $X2=3.215 $Y2=1.045
r46 17 22 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=3.485 $Y=1.885
+ $X2=3.6 $Y2=1.8
r47 17 18 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=3.485 $Y=1.885
+ $X2=3.19 $Y2=1.885
r48 13 20 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=3.09 $Y=0.96
+ $X2=3.215 $Y2=1.045
r49 13 15 20.5135 $w=2.48e-07 $l=4.45e-07 $layer=LI1_cond $X=3.09 $Y=0.96
+ $X2=3.09 $Y2=0.515
r50 9 11 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=3.025 $Y=1.985
+ $X2=3.025 $Y2=2.815
r51 7 18 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.025 $Y=1.97
+ $X2=3.19 $Y2=1.885
r52 7 9 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=3.025 $Y=1.97
+ $X2=3.025 $Y2=1.985
r53 2 11 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=2.875
+ $Y=1.84 $X2=3.025 $Y2=2.815
r54 2 9 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=2.875
+ $Y=1.84 $X2=3.025 $Y2=1.985
r55 1 15 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.99
+ $Y=0.37 $X2=3.13 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__OR4_2%VGND 1 2 3 4 13 15 17 21 25 27 29 31 33 38 47
+ 50 54
r58 53 54 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r59 50 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r60 47 48 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r61 45 48 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=1.2
+ $Y2=0
r62 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r63 42 54 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=3.6
+ $Y2=0
r64 42 51 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=2.64
+ $Y2=0
r65 41 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r66 39 50 10.3577 $w=1.7e-07 $l=2.18e-07 $layer=LI1_cond $X=2.795 $Y=0 $X2=2.577
+ $Y2=0
r67 39 41 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=2.795 $Y=0 $X2=3.12
+ $Y2=0
r68 38 53 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=3.395 $Y=0 $X2=3.617
+ $Y2=0
r69 38 41 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=3.395 $Y=0 $X2=3.12
+ $Y2=0
r70 37 51 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r71 36 37 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r72 34 47 11.015 $w=1.7e-07 $l=2.4e-07 $layer=LI1_cond $X=1.68 $Y=0 $X2=1.44
+ $Y2=0
r73 34 36 31.3155 $w=1.68e-07 $l=4.8e-07 $layer=LI1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r74 33 50 10.3577 $w=1.7e-07 $l=2.17e-07 $layer=LI1_cond $X=2.36 $Y=0 $X2=2.577
+ $Y2=0
r75 33 36 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=2.36 $Y=0 $X2=2.16
+ $Y2=0
r76 31 37 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=2.16
+ $Y2=0
r77 31 48 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=1.2
+ $Y2=0
r78 27 53 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=3.56 $Y=0.085
+ $X2=3.617 $Y2=0
r79 27 29 18.3343 $w=3.28e-07 $l=5.25e-07 $layer=LI1_cond $X=3.56 $Y=0.085
+ $X2=3.56 $Y2=0.61
r80 23 50 1.70358 $w=4.35e-07 $l=8.5e-08 $layer=LI1_cond $X=2.577 $Y=0.085
+ $X2=2.577 $Y2=0
r81 23 25 14.836 $w=4.33e-07 $l=5.6e-07 $layer=LI1_cond $X=2.577 $Y=0.085
+ $X2=2.577 $Y2=0.645
r82 19 47 1.96841 $w=4.8e-07 $l=8.5e-08 $layer=LI1_cond $X=1.44 $Y=0.085
+ $X2=1.44 $Y2=0
r83 19 21 10.0919 $w=4.78e-07 $l=4.05e-07 $layer=LI1_cond $X=1.44 $Y=0.085
+ $X2=1.44 $Y2=0.49
r84 18 44 5.3488 $w=1.7e-07 $l=2.55e-07 $layer=LI1_cond $X=0.51 $Y=0 $X2=0.255
+ $Y2=0
r85 17 47 11.015 $w=1.7e-07 $l=2.4e-07 $layer=LI1_cond $X=1.2 $Y=0 $X2=1.44
+ $Y2=0
r86 17 18 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.2 $Y=0 $X2=0.51
+ $Y2=0
r87 13 44 2.97855 $w=3.95e-07 $l=1.09864e-07 $layer=LI1_cond $X=0.312 $Y=0.085
+ $X2=0.255 $Y2=0
r88 13 15 11.8162 $w=3.93e-07 $l=4.05e-07 $layer=LI1_cond $X=0.312 $Y=0.085
+ $X2=0.312 $Y2=0.49
r89 4 29 182 $w=1.7e-07 $l=3.01993e-07 $layer=licon1_NDIFF $count=1 $X=3.42
+ $Y=0.37 $X2=3.56 $Y2=0.61
r90 3 25 182 $w=1.7e-07 $l=3.87137e-07 $layer=licon1_NDIFF $count=1 $X=2.315
+ $Y=0.37 $X2=2.585 $Y2=0.645
r91 2 21 182 $w=1.7e-07 $l=3.49893e-07 $layer=licon1_NDIFF $count=1 $X=1.145
+ $Y=0.37 $X2=1.44 $Y2=0.49
r92 1 15 182 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.345 $X2=0.31 $Y2=0.49
.ends

