* File: sky130_fd_sc_hs__a2bb2o_1.pex.spice
* Created: Tue Sep  1 19:51:40 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HS__A2BB2O_1%A_93_264# 1 2 7 9 12 15 16 17 19 20 22 23
+ 25 28 30 32 38 40
c101 40 0 7.12326e-20 $X=1.41 $Y=1.875
r102 35 38 6.46067 $w=3.28e-07 $l=1.85e-07 $layer=LI1_cond $X=0.63 $Y=1.485
+ $X2=0.815 $Y2=1.485
r103 35 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.63
+ $Y=1.485 $X2=0.63 $Y2=1.485
r104 30 32 33.5808 $w=1.78e-07 $l=5.45e-07 $layer=LI1_cond $X=2.19 $Y=1.12
+ $X2=2.735 $Y2=1.12
r105 26 28 9.42908 $w=3.28e-07 $l=2.7e-07 $layer=LI1_cond $X=2.35 $Y=2.905
+ $X2=2.35 $Y2=2.635
r106 24 30 6.82373 $w=1.8e-07 $l=1.25499e-07 $layer=LI1_cond $X=2.105 $Y=1.21
+ $X2=2.19 $Y2=1.12
r107 24 25 37.8396 $w=1.68e-07 $l=5.8e-07 $layer=LI1_cond $X=2.105 $Y=1.21
+ $X2=2.105 $Y2=1.79
r108 22 26 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.185 $Y=2.99
+ $X2=2.35 $Y2=2.905
r109 22 23 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=2.185 $Y=2.99
+ $X2=1.495 $Y2=2.99
r110 21 40 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.495 $Y=1.875
+ $X2=1.41 $Y2=1.875
r111 20 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.02 $Y=1.875
+ $X2=2.105 $Y2=1.79
r112 20 21 34.2513 $w=1.68e-07 $l=5.25e-07 $layer=LI1_cond $X=2.02 $Y=1.875
+ $X2=1.495 $Y2=1.875
r113 19 23 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.41 $Y=2.905
+ $X2=1.495 $Y2=2.99
r114 18 40 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.41 $Y=1.96
+ $X2=1.41 $Y2=1.875
r115 18 19 61.6524 $w=1.68e-07 $l=9.45e-07 $layer=LI1_cond $X=1.41 $Y=1.96
+ $X2=1.41 $Y2=2.905
r116 16 40 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.325 $Y=1.875
+ $X2=1.41 $Y2=1.875
r117 16 17 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=1.325 $Y=1.875
+ $X2=0.9 $Y2=1.875
r118 15 17 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.815 $Y=1.79
+ $X2=0.9 $Y2=1.875
r119 14 38 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.815 $Y=1.65
+ $X2=0.815 $Y2=1.485
r120 14 15 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=0.815 $Y=1.65
+ $X2=0.815 $Y2=1.79
r121 10 36 38.6072 $w=2.91e-07 $l=2.05122e-07 $layer=POLY_cond $X=0.72 $Y=1.32
+ $X2=0.63 $Y2=1.485
r122 10 12 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=0.72 $Y=1.32
+ $X2=0.72 $Y2=0.81
r123 7 36 57.6553 $w=2.91e-07 $l=3.1305e-07 $layer=POLY_cond $X=0.7 $Y=1.765
+ $X2=0.63 $Y2=1.485
r124 7 9 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.7 $Y=1.765 $X2=0.7
+ $Y2=2.4
r125 2 28 600 $w=1.7e-07 $l=7.34847e-07 $layer=licon1_PDIFF $count=1 $X=2.225
+ $Y=1.96 $X2=2.35 $Y2=2.635
r126 1 32 182 $w=1.7e-07 $l=5.55608e-07 $layer=licon1_NDIFF $count=1 $X=2.595
+ $Y=0.63 $X2=2.735 $Y2=1.12
.ends

.subckt PM_SKY130_FD_SC_HS__A2BB2O_1%A1_N 2 5 6 8 9 12 14
c42 14 0 1.8858e-19 $X=1.17 $Y=1.29
c43 12 0 7.12326e-20 $X=1.17 $Y=1.455
r44 12 15 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.17 $Y=1.455
+ $X2=1.17 $Y2=1.62
r45 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.17 $Y=1.455
+ $X2=1.17 $Y2=1.29
r46 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.17
+ $Y=1.455 $X2=1.17 $Y2=1.455
r47 9 13 6.95815 $w=2.63e-07 $l=1.6e-07 $layer=LI1_cond $X=1.202 $Y=1.295
+ $X2=1.202 $Y2=1.455
r48 6 8 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=1.215 $Y=1.885
+ $X2=1.215 $Y2=2.46
r49 5 14 123.713 $w=1.5e-07 $l=3.85e-07 $layer=POLY_cond $X=1.21 $Y=0.905
+ $X2=1.21 $Y2=1.29
r50 2 6 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=1.215 $Y=1.795 $X2=1.215
+ $Y2=1.885
r51 2 15 68.0242 $w=1.8e-07 $l=1.75e-07 $layer=POLY_cond $X=1.215 $Y=1.795
+ $X2=1.215 $Y2=1.62
.ends

.subckt PM_SKY130_FD_SC_HS__A2BB2O_1%A2_N 1 3 4 6 7
c39 7 0 1.96077e-19 $X=1.68 $Y=1.295
r40 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.71
+ $Y=1.455 $X2=1.71 $Y2=1.455
r41 7 11 6.0456 $w=3.03e-07 $l=1.6e-07 $layer=LI1_cond $X=1.697 $Y=1.295
+ $X2=1.697 $Y2=1.455
r42 4 10 39.2307 $w=2.57e-07 $l=1.90526e-07 $layer=POLY_cond $X=1.64 $Y=1.29
+ $X2=1.695 $Y2=1.455
r43 4 6 123.713 $w=1.5e-07 $l=3.85e-07 $layer=POLY_cond $X=1.64 $Y=1.29 $X2=1.64
+ $Y2=0.905
r44 1 10 88.9311 $w=2.57e-07 $l=4.72864e-07 $layer=POLY_cond $X=1.605 $Y=1.885
+ $X2=1.695 $Y2=1.455
r45 1 3 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=1.605 $Y=1.885
+ $X2=1.605 $Y2=2.46
.ends

.subckt PM_SKY130_FD_SC_HS__A2BB2O_1%A_257_126# 1 2 10 11 13 16 18 20 21 25 28
+ 30 32
c71 20 0 2.008e-20 $X=2.43 $Y=0.355
c72 18 0 1.8858e-19 $X=1.59 $Y=0.387
c73 10 0 1.96077e-19 $X=2.52 $Y=0.95
r74 32 35 8.47458 $w=3.03e-07 $l=1.65e-07 $layer=LI1_cond $X=2.512 $Y=1.615
+ $X2=2.512 $Y2=1.78
r75 32 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.5
+ $Y=1.615 $X2=2.5 $Y2=1.615
r76 28 35 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=2.445 $Y=2.13
+ $X2=2.445 $Y2=1.78
r77 26 30 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.995 $Y=2.215
+ $X2=1.83 $Y2=2.215
r78 25 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.36 $Y=2.215
+ $X2=2.445 $Y2=2.13
r79 25 26 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=2.36 $Y=2.215
+ $X2=1.995 $Y2=2.215
r80 21 38 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.43 $Y=0.355
+ $X2=2.43 $Y2=0.52
r81 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.43
+ $Y=0.355 $X2=2.43 $Y2=0.355
r82 18 20 36.5303 $w=2.63e-07 $l=8.4e-07 $layer=LI1_cond $X=1.59 $Y=0.387
+ $X2=2.43 $Y2=0.387
r83 14 18 6.86024 $w=2.65e-07 $l=2.09184e-07 $layer=LI1_cond $X=1.437 $Y=0.52
+ $X2=1.59 $Y2=0.387
r84 14 16 12.2801 $w=3.03e-07 $l=3.25e-07 $layer=LI1_cond $X=1.437 $Y=0.52
+ $X2=1.437 $Y2=0.845
r85 11 33 55.8646 $w=2.93e-07 $l=3.05205e-07 $layer=POLY_cond $X=2.575 $Y=1.885
+ $X2=2.5 $Y2=1.615
r86 11 13 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=2.575 $Y=1.885
+ $X2=2.575 $Y2=2.46
r87 10 38 220.489 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=2.52 $Y=0.95
+ $X2=2.52 $Y2=0.52
r88 8 33 38.5916 $w=2.93e-07 $l=1.74714e-07 $layer=POLY_cond $X=2.52 $Y=1.45
+ $X2=2.5 $Y2=1.615
r89 8 10 256.383 $w=1.5e-07 $l=5e-07 $layer=POLY_cond $X=2.52 $Y=1.45 $X2=2.52
+ $Y2=0.95
r90 2 30 300 $w=1.7e-07 $l=3.21364e-07 $layer=licon1_PDIFF $count=2 $X=1.68
+ $Y=1.96 $X2=1.83 $Y2=2.215
r91 1 16 182 $w=1.7e-07 $l=2.7627e-07 $layer=licon1_NDIFF $count=1 $X=1.285
+ $Y=0.63 $X2=1.425 $Y2=0.845
.ends

.subckt PM_SKY130_FD_SC_HS__A2BB2O_1%B2 3 5 7 8
c36 3 0 2.008e-20 $X=2.95 $Y=0.95
r37 8 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.04
+ $Y=1.615 $X2=3.04 $Y2=1.615
r38 5 11 55.8646 $w=2.93e-07 $l=2.77399e-07 $layer=POLY_cond $X=3.025 $Y=1.885
+ $X2=3.04 $Y2=1.615
r39 5 7 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=3.025 $Y=1.885
+ $X2=3.025 $Y2=2.46
r40 1 11 38.5916 $w=2.93e-07 $l=2.05122e-07 $layer=POLY_cond $X=2.95 $Y=1.45
+ $X2=3.04 $Y2=1.615
r41 1 3 256.383 $w=1.5e-07 $l=5e-07 $layer=POLY_cond $X=2.95 $Y=1.45 $X2=2.95
+ $Y2=0.95
.ends

.subckt PM_SKY130_FD_SC_HS__A2BB2O_1%B1 4 5 6 7 9 11 12 18
c31 4 0 5.93438e-20 $X=3.49 $Y=0.95
r32 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.65
+ $Y=0.355 $X2=3.65 $Y2=0.355
r33 15 18 27.9778 $w=3.3e-07 $l=1.6e-07 $layer=POLY_cond $X=3.49 $Y=0.355
+ $X2=3.65 $Y2=0.355
r34 12 19 11.941 $w=4.13e-07 $l=4.3e-07 $layer=LI1_cond $X=4.08 $Y=0.462
+ $X2=3.65 $Y2=0.462
r35 11 19 1.38849 $w=4.13e-07 $l=5e-08 $layer=LI1_cond $X=3.6 $Y=0.462 $X2=3.65
+ $Y2=0.462
r36 7 9 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=3.505 $Y=1.885
+ $X2=3.505 $Y2=2.46
r37 6 7 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=3.505 $Y=1.795 $X2=3.505
+ $Y2=1.885
r38 5 10 37.1337 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=3.505 $Y=1.435
+ $X2=3.505 $Y2=1.345
r39 5 6 139.935 $w=1.8e-07 $l=3.6e-07 $layer=POLY_cond $X=3.505 $Y=1.435
+ $X2=3.505 $Y2=1.795
r40 4 10 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=3.49 $Y=0.95
+ $X2=3.49 $Y2=1.345
r41 1 15 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.49 $Y=0.52
+ $X2=3.49 $Y2=0.355
r42 1 4 220.489 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=3.49 $Y=0.52 $X2=3.49
+ $Y2=0.95
.ends

.subckt PM_SKY130_FD_SC_HS__A2BB2O_1%X 1 2 9 13 14 15 16 31 32 35
r22 31 32 8.80985 $w=4.33e-07 $l=1.65e-07 $layer=LI1_cond $X=0.342 $Y=1.985
+ $X2=0.342 $Y2=1.82
r23 21 35 0.0529859 $w=4.33e-07 $l=2e-09 $layer=LI1_cond $X=0.342 $Y=2.037
+ $X2=0.342 $Y2=2.035
r24 16 28 1.05972 $w=4.33e-07 $l=4e-08 $layer=LI1_cond $X=0.342 $Y=2.775
+ $X2=0.342 $Y2=2.815
r25 15 16 9.80239 $w=4.33e-07 $l=3.7e-07 $layer=LI1_cond $X=0.342 $Y=2.405
+ $X2=0.342 $Y2=2.775
r26 14 35 1.1127 $w=4.33e-07 $l=4.2e-08 $layer=LI1_cond $X=0.342 $Y=1.993
+ $X2=0.342 $Y2=2.035
r27 14 31 0.211944 $w=4.33e-07 $l=8e-09 $layer=LI1_cond $X=0.342 $Y=1.993
+ $X2=0.342 $Y2=1.985
r28 14 15 8.66319 $w=4.33e-07 $l=3.27e-07 $layer=LI1_cond $X=0.342 $Y=2.078
+ $X2=0.342 $Y2=2.405
r29 14 21 1.08621 $w=4.33e-07 $l=4.1e-08 $layer=LI1_cond $X=0.342 $Y=2.078
+ $X2=0.342 $Y2=2.037
r30 13 32 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=0.21 $Y=1.15
+ $X2=0.21 $Y2=1.82
r31 7 13 11.032 $w=4.63e-07 $l=2.32e-07 $layer=LI1_cond $X=0.357 $Y=0.918
+ $X2=0.357 $Y2=1.15
r32 7 9 8.56546 $w=4.63e-07 $l=3.33e-07 $layer=LI1_cond $X=0.357 $Y=0.918
+ $X2=0.357 $Y2=0.585
r33 2 31 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.35
+ $Y=1.84 $X2=0.475 $Y2=1.985
r34 2 28 400 $w=1.7e-07 $l=1.03562e-06 $layer=licon1_PDIFF $count=1 $X=0.35
+ $Y=1.84 $X2=0.475 $Y2=2.815
r35 1 9 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.38
+ $Y=0.44 $X2=0.505 $Y2=0.585
.ends

.subckt PM_SKY130_FD_SC_HS__A2BB2O_1%VPWR 1 2 9 13 16 17 18 24 30 31 34
r47 34 35 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r48 31 35 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=3.12 $Y2=3.33
r49 30 31 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r50 28 34 9.14399 $w=1.7e-07 $l=1.8e-07 $layer=LI1_cond $X=3.445 $Y=3.33
+ $X2=3.265 $Y2=3.33
r51 28 30 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=3.445 $Y=3.33
+ $X2=4.08 $Y2=3.33
r52 26 27 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r53 24 34 9.14399 $w=1.7e-07 $l=1.8e-07 $layer=LI1_cond $X=3.085 $Y=3.33
+ $X2=3.265 $Y2=3.33
r54 24 26 122.979 $w=1.68e-07 $l=1.885e-06 $layer=LI1_cond $X=3.085 $Y=3.33
+ $X2=1.2 $Y2=3.33
r55 22 27 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r56 21 22 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r57 18 35 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=3.12 $Y2=3.33
r58 18 27 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.2 $Y2=3.33
r59 16 21 2.60963 $w=1.68e-07 $l=4e-08 $layer=LI1_cond $X=0.76 $Y=3.33 $X2=0.72
+ $Y2=3.33
r60 16 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.76 $Y=3.33
+ $X2=0.925 $Y2=3.33
r61 15 26 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=1.09 $Y=3.33 $X2=1.2
+ $Y2=3.33
r62 15 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.09 $Y=3.33
+ $X2=0.925 $Y2=3.33
r63 11 34 1.16013 $w=3.6e-07 $l=8.5e-08 $layer=LI1_cond $X=3.265 $Y=3.245
+ $X2=3.265 $Y2=3.33
r64 11 13 25.2897 $w=3.58e-07 $l=7.9e-07 $layer=LI1_cond $X=3.265 $Y=3.245
+ $X2=3.265 $Y2=2.455
r65 7 17 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.925 $Y=3.245
+ $X2=0.925 $Y2=3.33
r66 7 9 34.2241 $w=3.28e-07 $l=9.8e-07 $layer=LI1_cond $X=0.925 $Y=3.245
+ $X2=0.925 $Y2=2.265
r67 2 13 300 $w=1.7e-07 $l=5.71577e-07 $layer=licon1_PDIFF $count=2 $X=3.1
+ $Y=1.96 $X2=3.265 $Y2=2.455
r68 1 9 300 $w=1.7e-07 $l=4.94343e-07 $layer=licon1_PDIFF $count=2 $X=0.775
+ $Y=1.84 $X2=0.925 $Y2=2.265
.ends

.subckt PM_SKY130_FD_SC_HS__A2BB2O_1%A_530_392# 1 2 7 9 11 13 15
r30 13 20 2.9222 $w=2.5e-07 $l=9e-08 $layer=LI1_cond $X=3.77 $Y=2.12 $X2=3.77
+ $Y2=2.03
r31 13 15 32.0379 $w=2.48e-07 $l=6.95e-07 $layer=LI1_cond $X=3.77 $Y=2.12
+ $X2=3.77 $Y2=2.815
r32 12 18 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.885 $Y=2.035
+ $X2=2.8 $Y2=2.035
r33 11 20 4.22096 $w=1.7e-07 $l=1.27475e-07 $layer=LI1_cond $X=3.645 $Y=2.035
+ $X2=3.77 $Y2=2.03
r34 11 12 49.5829 $w=1.68e-07 $l=7.6e-07 $layer=LI1_cond $X=3.645 $Y=2.035
+ $X2=2.885 $Y2=2.035
r35 7 18 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.8 $Y=2.12 $X2=2.8
+ $Y2=2.035
r36 7 9 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=2.8 $Y=2.12 $X2=2.8
+ $Y2=2.815
r37 2 20 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=3.58
+ $Y=1.96 $X2=3.73 $Y2=2.105
r38 2 15 400 $w=1.7e-07 $l=9.26971e-07 $layer=licon1_PDIFF $count=1 $X=3.58
+ $Y=1.96 $X2=3.73 $Y2=2.815
r39 1 18 400 $w=1.7e-07 $l=2.17428e-07 $layer=licon1_PDIFF $count=1 $X=2.65
+ $Y=1.96 $X2=2.8 $Y2=2.115
r40 1 9 400 $w=1.7e-07 $l=9.26971e-07 $layer=licon1_PDIFF $count=1 $X=2.65
+ $Y=1.96 $X2=2.8 $Y2=2.815
.ends

.subckt PM_SKY130_FD_SC_HS__A2BB2O_1%VGND 1 2 3 12 14 19 21 22 23 25 26 28 29 31
+ 32 33 38 54 55
c77 14 0 5.93438e-20 $X=2.765 $Y=0.775
r78 54 55 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r79 52 55 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=4.08
+ $Y2=0
r80 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r81 49 52 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r82 48 49 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r83 45 48 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.2 $Y=0 $X2=2.64
+ $Y2=0
r84 45 46 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r85 42 46 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r86 41 42 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r87 38 49 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r88 38 46 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.2
+ $Y2=0
r89 33 36 4.88915 $w=3.28e-07 $l=1.4e-07 $layer=LI1_cond $X=3.705 $Y=0.925
+ $X2=3.705 $Y2=1.065
r90 31 51 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=3.145 $Y=0 $X2=3.12
+ $Y2=0
r91 31 32 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.145 $Y=0 $X2=3.23
+ $Y2=0
r92 30 54 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=3.315 $Y=0 $X2=4.08
+ $Y2=0
r93 30 32 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.315 $Y=0 $X2=3.23
+ $Y2=0
r94 28 48 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=2.765 $Y=0 $X2=2.64
+ $Y2=0
r95 28 29 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.765 $Y=0 $X2=2.85
+ $Y2=0
r96 27 51 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=2.935 $Y=0 $X2=3.12
+ $Y2=0
r97 27 29 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.935 $Y=0 $X2=2.85
+ $Y2=0
r98 25 41 3.26203 $w=1.68e-07 $l=5e-08 $layer=LI1_cond $X=0.77 $Y=0 $X2=0.72
+ $Y2=0
r99 25 26 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.77 $Y=0 $X2=0.935
+ $Y2=0
r100 24 45 6.52406 $w=1.68e-07 $l=1e-07 $layer=LI1_cond $X=1.1 $Y=0 $X2=1.2
+ $Y2=0
r101 24 26 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.1 $Y=0 $X2=0.935
+ $Y2=0
r102 22 33 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.54 $Y=0.925
+ $X2=3.705 $Y2=0.925
r103 22 23 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=3.54 $Y=0.925
+ $X2=3.315 $Y2=0.925
r104 21 23 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.23 $Y=0.84
+ $X2=3.315 $Y2=0.925
r105 20 32 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.23 $Y=0.085
+ $X2=3.23 $Y2=0
r106 20 21 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=3.23 $Y=0.085
+ $X2=3.23 $Y2=0.84
r107 18 29 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.85 $Y=0.085
+ $X2=2.85 $Y2=0
r108 18 19 39.4706 $w=1.68e-07 $l=6.05e-07 $layer=LI1_cond $X=2.85 $Y=0.085
+ $X2=2.85 $Y2=0.69
r109 14 19 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.765 $Y=0.775
+ $X2=2.85 $Y2=0.69
r110 14 16 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=2.765 $Y=0.775
+ $X2=2.305 $Y2=0.775
r111 10 26 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.935 $Y=0.085
+ $X2=0.935 $Y2=0
r112 10 12 17.4613 $w=3.28e-07 $l=5e-07 $layer=LI1_cond $X=0.935 $Y=0.085
+ $X2=0.935 $Y2=0.585
r113 3 36 182 $w=1.7e-07 $l=5.00125e-07 $layer=licon1_NDIFF $count=1 $X=3.565
+ $Y=0.63 $X2=3.705 $Y2=1.065
r114 2 16 91 $w=1.7e-07 $l=6.58521e-07 $layer=licon1_NDIFF $count=2 $X=1.715
+ $Y=0.63 $X2=2.305 $Y2=0.775
r115 1 12 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=0.795
+ $Y=0.44 $X2=0.935 $Y2=0.585
.ends

