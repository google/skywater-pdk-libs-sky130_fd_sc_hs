* File: sky130_fd_sc_hs__a221o_1.pex.spice
* Created: Tue Sep  1 19:50:08 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HS__A221O_1%A_148_260# 1 2 3 10 12 15 17 18 21 23 27 35
+ 37
r82 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.905
+ $Y=1.465 $X2=0.905 $Y2=1.465
r83 27 29 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=4.05 $Y=2.105
+ $X2=4.05 $Y2=2.815
r84 27 40 28.6365 $w=3.28e-07 $l=8.2e-07 $layer=LI1_cond $X=4.05 $Y=2.105
+ $X2=4.05 $Y2=1.285
r85 24 35 10.4332 $w=1.7e-07 $l=5.26498e-07 $layer=LI1_cond $X=2.86 $Y=1.2
+ $X2=2.42 $Y2=1.01
r86 23 40 2.83394 $w=3.53e-07 $l=8.5e-08 $layer=LI1_cond $X=4.037 $Y=1.2
+ $X2=4.037 $Y2=1.285
r87 23 37 6.33032 $w=3.53e-07 $l=1.95e-07 $layer=LI1_cond $X=4.037 $Y=1.2
+ $X2=4.037 $Y2=1.005
r88 23 24 65.2406 $w=1.68e-07 $l=1e-06 $layer=LI1_cond $X=3.86 $Y=1.2 $X2=2.86
+ $Y2=1.2
r89 19 35 1.73497 $w=4.4e-07 $l=2.2e-07 $layer=LI1_cond $X=2.64 $Y=1.01 $X2=2.42
+ $Y2=1.01
r90 19 21 12.834 $w=4.38e-07 $l=4.9e-07 $layer=LI1_cond $X=2.64 $Y=1.01 $X2=2.64
+ $Y2=0.52
r91 18 33 13.8043 $w=3.27e-07 $l=4.72345e-07 $layer=LI1_cond $X=1.205 $Y=1.095
+ $X2=0.972 $Y2=1.465
r92 17 35 10.4332 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.42 $Y=1.095
+ $X2=2.42 $Y2=1.01
r93 17 18 79.2674 $w=1.68e-07 $l=1.215e-06 $layer=LI1_cond $X=2.42 $Y=1.095
+ $X2=1.205 $Y2=1.095
r94 13 34 38.6549 $w=2.86e-07 $l=2.05122e-07 $layer=POLY_cond $X=0.995 $Y=1.3
+ $X2=0.905 $Y2=1.465
r95 13 15 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=0.995 $Y=1.3
+ $X2=0.995 $Y2=0.74
r96 10 34 61.4066 $w=2.86e-07 $l=3.26343e-07 $layer=POLY_cond $X=0.96 $Y=1.765
+ $X2=0.905 $Y2=1.465
r97 10 12 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.96 $Y=1.765
+ $X2=0.96 $Y2=2.4
r98 3 29 400 $w=1.7e-07 $l=9.26971e-07 $layer=licon1_PDIFF $count=1 $X=3.9
+ $Y=1.96 $X2=4.05 $Y2=2.815
r99 3 27 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=3.9
+ $Y=1.96 $X2=4.05 $Y2=2.105
r100 2 37 182 $w=1.7e-07 $l=4.54643e-07 $layer=licon1_NDIFF $count=1 $X=3.885
+ $Y=0.615 $X2=4.025 $Y2=1.005
r101 1 21 91 $w=1.7e-07 $l=2.498e-07 $layer=licon1_NDIFF $count=2 $X=2.445
+ $Y=0.395 $X2=2.64 $Y2=0.52
.ends

.subckt PM_SKY130_FD_SC_HS__A221O_1%A2 1 3 4 6 8 9
r39 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.46
+ $Y=1.515 $X2=1.46 $Y2=1.515
r40 9 14 5.89622 $w=4.28e-07 $l=2.2e-07 $layer=LI1_cond $X=1.68 $Y=1.565
+ $X2=1.46 $Y2=1.565
r41 6 8 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=2.01 $Y=1.11 $X2=2.01
+ $Y2=0.715
r42 5 13 62.3765 $w=2.55e-07 $l=4.04166e-07 $layer=POLY_cond $X=1.625 $Y=1.185
+ $X2=1.46 $Y2=1.515
r43 4 6 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.935 $Y=1.185
+ $X2=2.01 $Y2=1.11
r44 4 5 158.957 $w=1.5e-07 $l=3.1e-07 $layer=POLY_cond $X=1.935 $Y=1.185
+ $X2=1.625 $Y2=1.185
r45 1 13 78.0421 $w=2.55e-07 $l=3.77425e-07 $layer=POLY_cond $X=1.475 $Y=1.885
+ $X2=1.46 $Y2=1.515
r46 1 3 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=1.475 $Y=1.885
+ $X2=1.475 $Y2=2.46
.ends

.subckt PM_SKY130_FD_SC_HS__A221O_1%A1 1 3 6 8 12
r39 12 14 32.5859 $w=3.55e-07 $l=2.4e-07 $layer=POLY_cond $X=2.13 $Y=1.677
+ $X2=2.37 $Y2=1.677
r40 10 12 27.8338 $w=3.55e-07 $l=2.05e-07 $layer=POLY_cond $X=1.925 $Y=1.677
+ $X2=2.13 $Y2=1.677
r41 8 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.13
+ $Y=1.635 $X2=2.13 $Y2=1.635
r42 4 14 22.9692 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.37 $Y=1.47
+ $X2=2.37 $Y2=1.677
r43 4 6 387.138 $w=1.5e-07 $l=7.55e-07 $layer=POLY_cond $X=2.37 $Y=1.47 $X2=2.37
+ $Y2=0.715
r44 1 10 22.9692 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=1.925 $Y=1.885
+ $X2=1.925 $Y2=1.677
r45 1 3 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=1.925 $Y=1.885
+ $X2=1.925 $Y2=2.46
.ends

.subckt PM_SKY130_FD_SC_HS__A221O_1%B1 1 3 6 8 12
r33 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.82
+ $Y=1.615 $X2=2.82 $Y2=1.615
r34 8 12 6.38276 $w=3.23e-07 $l=1.8e-07 $layer=LI1_cond $X=2.64 $Y=1.617
+ $X2=2.82 $Y2=1.617
r35 4 11 38.5916 $w=2.93e-07 $l=2.05122e-07 $layer=POLY_cond $X=2.91 $Y=1.45
+ $X2=2.82 $Y2=1.615
r36 4 6 376.883 $w=1.5e-07 $l=7.35e-07 $layer=POLY_cond $X=2.91 $Y=1.45 $X2=2.91
+ $Y2=0.715
r37 1 11 55.8646 $w=2.93e-07 $l=3.05205e-07 $layer=POLY_cond $X=2.895 $Y=1.885
+ $X2=2.82 $Y2=1.615
r38 1 3 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=2.895 $Y=1.885
+ $X2=2.895 $Y2=2.46
.ends

.subckt PM_SKY130_FD_SC_HS__A221O_1%B2 3 5 7 8
c33 3 0 1.47272e-19 $X=3.27 $Y=0.715
r34 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.36
+ $Y=1.615 $X2=3.36 $Y2=1.615
r35 8 12 8.51035 $w=3.23e-07 $l=2.4e-07 $layer=LI1_cond $X=3.6 $Y=1.617 $X2=3.36
+ $Y2=1.617
r36 5 11 55.8646 $w=2.93e-07 $l=2.77399e-07 $layer=POLY_cond $X=3.345 $Y=1.885
+ $X2=3.36 $Y2=1.615
r37 5 7 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=3.345 $Y=1.885
+ $X2=3.345 $Y2=2.46
r38 1 11 38.5916 $w=2.93e-07 $l=2.05122e-07 $layer=POLY_cond $X=3.27 $Y=1.45
+ $X2=3.36 $Y2=1.615
r39 1 3 376.883 $w=1.5e-07 $l=7.35e-07 $layer=POLY_cond $X=3.27 $Y=1.45 $X2=3.27
+ $Y2=0.715
.ends

.subckt PM_SKY130_FD_SC_HS__A221O_1%C1 4 5 6 7 9 11 16 17
c30 17 0 1.47272e-19 $X=4.03 $Y=0.34
r31 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.03
+ $Y=0.34 $X2=4.03 $Y2=0.34
r32 13 16 38.4695 $w=3.3e-07 $l=2.2e-07 $layer=POLY_cond $X=3.81 $Y=0.34
+ $X2=4.03 $Y2=0.34
r33 11 17 7.50834 $w=3.28e-07 $l=2.15e-07 $layer=LI1_cond $X=4.03 $Y=0.555
+ $X2=4.03 $Y2=0.34
r34 7 9 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=3.825 $Y=1.885
+ $X2=3.825 $Y2=2.46
r35 6 7 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=3.825 $Y=1.795 $X2=3.825
+ $Y2=1.885
r36 5 10 37.1337 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=3.825 $Y=1.42 $X2=3.825
+ $Y2=1.33
r37 5 6 145.766 $w=1.8e-07 $l=3.75e-07 $layer=POLY_cond $X=3.825 $Y=1.42
+ $X2=3.825 $Y2=1.795
r38 4 10 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=3.81 $Y=0.935
+ $X2=3.81 $Y2=1.33
r39 1 13 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.81 $Y=0.505
+ $X2=3.81 $Y2=0.34
r40 1 4 220.489 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=3.81 $Y=0.505 $X2=3.81
+ $Y2=0.935
.ends

.subckt PM_SKY130_FD_SC_HS__A221O_1%X 1 2 12 14 15 16 27 28
r19 27 28 5.7419 $w=7.73e-07 $l=1.65e-07 $layer=LI1_cond $X=0.512 $Y=1.985
+ $X2=0.512 $Y2=1.82
r20 15 16 5.71031 $w=7.73e-07 $l=3.7e-07 $layer=LI1_cond $X=0.512 $Y=2.405
+ $X2=0.512 $Y2=2.775
r21 14 15 5.71031 $w=7.73e-07 $l=3.7e-07 $layer=LI1_cond $X=0.512 $Y=2.035
+ $X2=0.512 $Y2=2.405
r22 14 27 0.771663 $w=7.73e-07 $l=5e-08 $layer=LI1_cond $X=0.512 $Y=2.035
+ $X2=0.512 $Y2=1.985
r23 9 12 7.17647 $w=7.78e-07 $l=4.68e-07 $layer=LI1_cond $X=0.312 $Y=0.74
+ $X2=0.78 $Y2=0.74
r24 7 9 5.04298 $w=3.75e-07 $l=3.9e-07 $layer=LI1_cond $X=0.312 $Y=1.13
+ $X2=0.312 $Y2=0.74
r25 7 28 21.205 $w=3.73e-07 $l=6.9e-07 $layer=LI1_cond $X=0.312 $Y=1.13
+ $X2=0.312 $Y2=1.82
r26 2 16 400 $w=1.7e-07 $l=1.03562e-06 $layer=licon1_PDIFF $count=1 $X=0.61
+ $Y=1.84 $X2=0.735 $Y2=2.815
r27 2 27 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.61
+ $Y=1.84 $X2=0.735 $Y2=1.985
r28 1 12 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.655
+ $Y=0.37 $X2=0.78 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__A221O_1%VPWR 1 2 9 15 17 19 24 34 35 38 41
r45 38 39 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r46 34 35 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r47 32 35 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=4.08 $Y2=3.33
r48 31 34 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=2.64 $Y=3.33
+ $X2=4.08 $Y2=3.33
r49 31 32 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r50 29 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.315 $Y=3.33
+ $X2=2.15 $Y2=3.33
r51 29 31 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=2.315 $Y=3.33
+ $X2=2.64 $Y2=3.33
r52 28 39 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r53 27 28 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r54 25 38 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.35 $Y=3.33
+ $X2=1.225 $Y2=3.33
r55 25 27 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=1.35 $Y=3.33
+ $X2=1.68 $Y2=3.33
r56 24 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.985 $Y=3.33
+ $X2=2.15 $Y2=3.33
r57 24 27 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.985 $Y=3.33
+ $X2=1.68 $Y2=3.33
r58 22 39 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r59 21 22 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r60 19 38 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.1 $Y=3.33
+ $X2=1.225 $Y2=3.33
r61 19 21 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=1.1 $Y=3.33 $X2=0.72
+ $Y2=3.33
r62 17 32 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r63 17 28 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.68 $Y2=3.33
r64 17 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r65 13 41 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.15 $Y=3.245
+ $X2=2.15 $Y2=3.33
r66 13 15 26.8903 $w=3.28e-07 $l=7.7e-07 $layer=LI1_cond $X=2.15 $Y=3.245
+ $X2=2.15 $Y2=2.475
r67 9 12 32.2684 $w=2.48e-07 $l=7e-07 $layer=LI1_cond $X=1.225 $Y=2.115
+ $X2=1.225 $Y2=2.815
r68 7 38 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.225 $Y=3.245
+ $X2=1.225 $Y2=3.33
r69 7 12 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=1.225 $Y=3.245
+ $X2=1.225 $Y2=2.815
r70 2 15 300 $w=1.7e-07 $l=5.85214e-07 $layer=licon1_PDIFF $count=2 $X=2 $Y=1.96
+ $X2=2.15 $Y2=2.475
r71 1 12 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=1.035
+ $Y=1.84 $X2=1.185 $Y2=2.815
r72 1 9 400 $w=1.7e-07 $l=3.4187e-07 $layer=licon1_PDIFF $count=1 $X=1.035
+ $Y=1.84 $X2=1.185 $Y2=2.115
.ends

.subckt PM_SKY130_FD_SC_HS__A221O_1%A_310_392# 1 2 7 9 11 18
r32 12 16 4.19273 $w=1.7e-07 $l=1.29904e-07 $layer=LI1_cond $X=1.785 $Y=2.055
+ $X2=1.66 $Y2=2.045
r33 11 18 5.03363 $w=1.7e-07 $l=1.69926e-07 $layer=LI1_cond $X=2.955 $Y=2.055
+ $X2=3.12 $Y2=2.045
r34 11 12 76.3316 $w=1.68e-07 $l=1.17e-06 $layer=LI1_cond $X=2.955 $Y=2.055
+ $X2=1.785 $Y2=2.055
r35 7 16 2.95044 $w=2.5e-07 $l=9.5e-08 $layer=LI1_cond $X=1.66 $Y=2.14 $X2=1.66
+ $Y2=2.045
r36 7 9 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=1.66 $Y=2.14 $X2=1.66
+ $Y2=2.815
r37 2 18 300 $w=1.7e-07 $l=2.17428e-07 $layer=licon1_PDIFF $count=2 $X=2.97
+ $Y=1.96 $X2=3.12 $Y2=2.115
r38 1 16 400 $w=1.7e-07 $l=2.17428e-07 $layer=licon1_PDIFF $count=1 $X=1.55
+ $Y=1.96 $X2=1.7 $Y2=2.115
r39 1 9 400 $w=1.7e-07 $l=9.26971e-07 $layer=licon1_PDIFF $count=1 $X=1.55
+ $Y=1.96 $X2=1.7 $Y2=2.815
.ends

.subckt PM_SKY130_FD_SC_HS__A221O_1%A_509_392# 1 2 9 11 12 15
r24 15 18 38.8182 $w=1.98e-07 $l=7e-07 $layer=LI1_cond $X=3.585 $Y=2.115
+ $X2=3.585 $Y2=2.815
r25 13 18 4.99091 $w=1.98e-07 $l=9e-08 $layer=LI1_cond $X=3.585 $Y=2.905
+ $X2=3.585 $Y2=2.815
r26 11 13 6.87494 $w=1.7e-07 $l=1.36015e-07 $layer=LI1_cond $X=3.485 $Y=2.99
+ $X2=3.585 $Y2=2.905
r27 11 12 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=3.485 $Y=2.99
+ $X2=2.785 $Y2=2.99
r28 7 12 7.36005 $w=1.7e-07 $l=1.77482e-07 $layer=LI1_cond $X=2.645 $Y=2.905
+ $X2=2.785 $Y2=2.99
r29 7 9 17.6982 $w=2.78e-07 $l=4.3e-07 $layer=LI1_cond $X=2.645 $Y=2.905
+ $X2=2.645 $Y2=2.475
r30 2 18 400 $w=1.7e-07 $l=9.33863e-07 $layer=licon1_PDIFF $count=1 $X=3.42
+ $Y=1.96 $X2=3.585 $Y2=2.815
r31 2 15 400 $w=1.7e-07 $l=2.29783e-07 $layer=licon1_PDIFF $count=1 $X=3.42
+ $Y=1.96 $X2=3.585 $Y2=2.115
r32 1 9 300 $w=1.7e-07 $l=5.74108e-07 $layer=licon1_PDIFF $count=2 $X=2.545
+ $Y=1.96 $X2=2.67 $Y2=2.475
.ends

.subckt PM_SKY130_FD_SC_HS__A221O_1%VGND 1 2 9 11 18 28 29 34 42 44
r43 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r44 41 42 12.4865 $w=9.23e-07 $l=1.7e-07 $layer=LI1_cond $X=1.795 $Y=0.377
+ $X2=1.965 $Y2=0.377
r45 38 41 1.51676 $w=9.23e-07 $l=1.15e-07 $layer=LI1_cond $X=1.68 $Y=0.377
+ $X2=1.795 $Y2=0.377
r46 38 39 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r47 36 38 6.19892 $w=9.23e-07 $l=4.7e-07 $layer=LI1_cond $X=1.21 $Y=0.377
+ $X2=1.68 $Y2=0.377
r48 33 39 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=1.68
+ $Y2=0
r49 32 36 0.131892 $w=9.23e-07 $l=1e-08 $layer=LI1_cond $X=1.2 $Y=0.377 $X2=1.21
+ $Y2=0.377
r50 32 34 12.2887 $w=9.23e-07 $l=1.55e-07 $layer=LI1_cond $X=1.2 $Y=0.377
+ $X2=1.045 $Y2=0.377
r51 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r52 29 45 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=3.6
+ $Y2=0
r53 28 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r54 26 44 9.31531 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=3.69 $Y=0 $X2=3.505
+ $Y2=0
r55 26 28 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=3.69 $Y=0 $X2=4.08
+ $Y2=0
r56 25 45 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=3.6
+ $Y2=0
r57 24 25 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r58 21 24 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=2.16 $Y=0 $X2=3.12
+ $Y2=0
r59 21 42 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=2.16 $Y=0 $X2=1.965
+ $Y2=0
r60 18 44 9.31531 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=3.32 $Y=0 $X2=3.505
+ $Y2=0
r61 18 24 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=3.32 $Y=0 $X2=3.12
+ $Y2=0
r62 16 33 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r63 15 34 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.72 $Y=0 $X2=1.045
+ $Y2=0
r64 15 16 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r65 11 25 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=3.12
+ $Y2=0
r66 11 39 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.68
+ $Y2=0
r67 11 21 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r68 7 44 1.24149 $w=3.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.505 $Y=0.085
+ $X2=3.505 $Y2=0
r69 7 9 13.549 $w=3.68e-07 $l=4.35e-07 $layer=LI1_cond $X=3.505 $Y=0.085
+ $X2=3.505 $Y2=0.52
r70 2 9 91 $w=1.7e-07 $l=2.13542e-07 $layer=licon1_NDIFF $count=2 $X=3.345
+ $Y=0.395 $X2=3.505 $Y2=0.52
r71 1 41 182 $w=1.7e-07 $l=8.64147e-07 $layer=licon1_NDIFF $count=1 $X=1.07
+ $Y=0.37 $X2=1.795 $Y2=0.675
r72 1 36 182 $w=1.7e-07 $l=3.68409e-07 $layer=licon1_NDIFF $count=1 $X=1.07
+ $Y=0.37 $X2=1.21 $Y2=0.675
.ends

