# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_hs__einvn_4
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_hs__einvn_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.280000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  1.116000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.035000 1.180000 5.155000 1.550000 ;
    END
  END A
  PIN TE_B
    ANTENNAGATEAREA  0.951000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.300000 0.455000 1.780000 ;
    END
  END TE_B
  PIN Z
    ANTENNADIFFAREA  1.086400 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.485000 1.550000 3.815000 1.720000 ;
        RECT 3.485000 1.720000 4.715000 1.890000 ;
        RECT 3.485000 1.890000 3.815000 2.735000 ;
        RECT 3.615000 0.770000 4.655000 1.010000 ;
        RECT 3.615000 1.010000 3.865000 1.130000 ;
        RECT 3.615000 1.130000 3.815000 1.550000 ;
        RECT 4.385000 1.890000 4.715000 2.735000 ;
        RECT 4.485000 0.595000 4.655000 0.770000 ;
    END
  END Z
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 5.280000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 5.280000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.280000 0.085000 ;
      RECT 0.000000  3.245000 5.280000 3.415000 ;
      RECT 0.115000  0.085000 0.365000 1.130000 ;
      RECT 0.175000  1.950000 0.425000 3.245000 ;
      RECT 0.545000  0.300000 1.295000 1.130000 ;
      RECT 0.625000  1.130000 1.295000 1.310000 ;
      RECT 0.625000  1.310000 0.955000 2.980000 ;
      RECT 1.185000  1.480000 3.285000 1.650000 ;
      RECT 1.185000  1.650000 1.435000 2.980000 ;
      RECT 1.465000  0.350000 1.635000 1.140000 ;
      RECT 1.465000  1.140000 3.435000 1.310000 ;
      RECT 1.635000  1.820000 1.885000 3.245000 ;
      RECT 1.815000  0.085000 2.145000 0.970000 ;
      RECT 2.085000  1.650000 2.335000 2.980000 ;
      RECT 2.325000  0.350000 2.495000 1.140000 ;
      RECT 2.535000  1.820000 2.865000 3.245000 ;
      RECT 2.675000  0.085000 3.005000 0.970000 ;
      RECT 3.035000  1.650000 3.285000 2.905000 ;
      RECT 3.035000  2.905000 5.165000 3.075000 ;
      RECT 3.185000  0.255000 5.165000 0.425000 ;
      RECT 3.185000  0.425000 4.305000 0.600000 ;
      RECT 3.185000  0.600000 3.435000 1.140000 ;
      RECT 4.015000  2.060000 4.185000 2.905000 ;
      RECT 4.835000  0.425000 5.165000 1.010000 ;
      RECT 4.915000  1.820000 5.165000 2.905000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
  END
END sky130_fd_sc_hs__einvn_4
END LIBRARY
