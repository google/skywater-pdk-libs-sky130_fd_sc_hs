* File: sky130_fd_sc_hs__nand2_8.pxi.spice
* Created: Tue Sep  1 20:08:48 2020
* 
x_PM_SKY130_FD_SC_HS__NAND2_8%B N_B_c_108_n N_B_M1000_g N_B_c_109_n N_B_c_110_n
+ N_B_c_111_n N_B_M1001_g N_B_c_112_n N_B_c_113_n N_B_M1003_g N_B_c_114_n
+ N_B_c_115_n N_B_M1010_g N_B_c_127_n N_B_M1002_g N_B_c_116_n N_B_M1011_g
+ N_B_c_128_n N_B_M1007_g N_B_M1012_g N_B_M1016_g N_B_M1017_g N_B_c_120_n
+ N_B_c_121_n N_B_c_131_n N_B_M1008_g N_B_c_122_n N_B_c_133_n N_B_M1022_g
+ N_B_c_123_n N_B_c_124_n N_B_c_125_n B B B B B PM_SKY130_FD_SC_HS__NAND2_8%B
x_PM_SKY130_FD_SC_HS__NAND2_8%A N_A_c_243_n N_A_M1004_g N_A_c_244_n N_A_c_245_n
+ N_A_c_246_n N_A_M1005_g N_A_c_247_n N_A_c_248_n N_A_M1006_g N_A_c_249_n
+ N_A_M1009_g N_A_c_260_n N_A_M1015_g N_A_c_250_n N_A_M1013_g N_A_c_261_n
+ N_A_M1019_g N_A_c_251_n N_A_M1014_g N_A_c_262_n N_A_M1020_g N_A_c_252_n
+ N_A_M1018_g N_A_c_253_n N_A_M1023_g N_A_c_263_n N_A_M1021_g N_A_c_254_n A A A
+ N_A_c_256_n N_A_c_257_n N_A_c_258_n N_A_c_267_n N_A_c_259_n A
+ PM_SKY130_FD_SC_HS__NAND2_8%A
x_PM_SKY130_FD_SC_HS__NAND2_8%VPWR N_VPWR_M1002_d N_VPWR_M1007_d N_VPWR_M1022_d
+ N_VPWR_M1015_s N_VPWR_M1019_s N_VPWR_M1021_s N_VPWR_c_362_n N_VPWR_c_363_n
+ N_VPWR_c_364_n N_VPWR_c_365_n N_VPWR_c_366_n N_VPWR_c_367_n N_VPWR_c_368_n
+ VPWR N_VPWR_c_369_n N_VPWR_c_370_n N_VPWR_c_371_n N_VPWR_c_372_n
+ N_VPWR_c_373_n N_VPWR_c_374_n N_VPWR_c_375_n N_VPWR_c_376_n N_VPWR_c_377_n
+ N_VPWR_c_361_n PM_SKY130_FD_SC_HS__NAND2_8%VPWR
x_PM_SKY130_FD_SC_HS__NAND2_8%Y N_Y_M1004_s N_Y_M1006_s N_Y_M1013_s N_Y_M1018_s
+ N_Y_M1002_s N_Y_M1008_s N_Y_M1015_d N_Y_M1020_d N_Y_c_450_n N_Y_c_445_n
+ N_Y_c_455_n N_Y_c_446_n N_Y_c_461_n N_Y_c_485_n N_Y_c_447_n N_Y_c_491_n
+ N_Y_c_448_n N_Y_c_495_n N_Y_c_442_n N_Y_c_443_n N_Y_c_463_n N_Y_c_505_n Y
+ PM_SKY130_FD_SC_HS__NAND2_8%Y
x_PM_SKY130_FD_SC_HS__NAND2_8%A_27_74# N_A_27_74#_M1000_s N_A_27_74#_M1001_s
+ N_A_27_74#_M1010_s N_A_27_74#_M1012_s N_A_27_74#_M1017_s N_A_27_74#_M1005_d
+ N_A_27_74#_M1009_d N_A_27_74#_M1014_d N_A_27_74#_M1023_d N_A_27_74#_c_551_n
+ N_A_27_74#_c_552_n N_A_27_74#_c_553_n N_A_27_74#_c_554_n N_A_27_74#_c_555_n
+ N_A_27_74#_c_556_n N_A_27_74#_c_557_n N_A_27_74#_c_558_n N_A_27_74#_c_559_n
+ N_A_27_74#_c_560_n N_A_27_74#_c_561_n N_A_27_74#_c_562_n N_A_27_74#_c_563_n
+ N_A_27_74#_c_564_n PM_SKY130_FD_SC_HS__NAND2_8%A_27_74#
x_PM_SKY130_FD_SC_HS__NAND2_8%VGND N_VGND_M1000_d N_VGND_M1003_d N_VGND_M1011_d
+ N_VGND_M1016_d N_VGND_c_655_n N_VGND_c_656_n N_VGND_c_657_n N_VGND_c_658_n
+ N_VGND_c_659_n N_VGND_c_660_n VGND N_VGND_c_661_n N_VGND_c_662_n
+ N_VGND_c_663_n N_VGND_c_664_n N_VGND_c_665_n N_VGND_c_666_n N_VGND_c_667_n
+ N_VGND_c_668_n PM_SKY130_FD_SC_HS__NAND2_8%VGND
cc_1 VNB N_B_c_108_n 0.0183176f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=1.185
cc_2 VNB N_B_c_109_n 0.0152334f $X=-0.19 $Y=-0.245 $X2=0.84 $Y2=1.26
cc_3 VNB N_B_c_110_n 0.0109496f $X=-0.19 $Y=-0.245 $X2=0.56 $Y2=1.26
cc_4 VNB N_B_c_111_n 0.0145126f $X=-0.19 $Y=-0.245 $X2=0.915 $Y2=1.185
cc_5 VNB N_B_c_112_n 0.0151763f $X=-0.19 $Y=-0.245 $X2=1.27 $Y2=1.26
cc_6 VNB N_B_c_113_n 0.0140036f $X=-0.19 $Y=-0.245 $X2=1.345 $Y2=1.185
cc_7 VNB N_B_c_114_n 0.0152048f $X=-0.19 $Y=-0.245 $X2=1.7 $Y2=1.26
cc_8 VNB N_B_c_115_n 0.0140065f $X=-0.19 $Y=-0.245 $X2=1.775 $Y2=1.185
cc_9 VNB N_B_c_116_n 0.0165f $X=-0.19 $Y=-0.245 $X2=2.205 $Y2=1.185
cc_10 VNB N_B_M1012_g 0.0266771f $X=-0.19 $Y=-0.245 $X2=2.955 $Y2=0.74
cc_11 VNB N_B_M1016_g 0.0230786f $X=-0.19 $Y=-0.245 $X2=3.425 $Y2=0.74
cc_12 VNB N_B_M1017_g 0.0231092f $X=-0.19 $Y=-0.245 $X2=3.855 $Y2=0.74
cc_13 VNB N_B_c_120_n 0.0112897f $X=-0.19 $Y=-0.245 $X2=4.23 $Y2=1.65
cc_14 VNB N_B_c_121_n 0.129918f $X=-0.19 $Y=-0.245 $X2=3.93 $Y2=1.65
cc_15 VNB N_B_c_122_n 0.0149373f $X=-0.19 $Y=-0.245 $X2=4.68 $Y2=1.65
cc_16 VNB N_B_c_123_n 0.00666874f $X=-0.19 $Y=-0.245 $X2=0.915 $Y2=1.26
cc_17 VNB N_B_c_124_n 0.00666874f $X=-0.19 $Y=-0.245 $X2=1.345 $Y2=1.26
cc_18 VNB N_B_c_125_n 0.00470774f $X=-0.19 $Y=-0.245 $X2=4.32 $Y2=1.67
cc_19 VNB B 0.00594092f $X=-0.19 $Y=-0.245 $X2=3.995 $Y2=1.58
cc_20 VNB N_A_c_243_n 0.0153183f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=1.185
cc_21 VNB N_A_c_244_n 0.0106299f $X=-0.19 $Y=-0.245 $X2=0.84 $Y2=1.26
cc_22 VNB N_A_c_245_n 0.00815376f $X=-0.19 $Y=-0.245 $X2=0.56 $Y2=1.26
cc_23 VNB N_A_c_246_n 0.014839f $X=-0.19 $Y=-0.245 $X2=0.915 $Y2=1.185
cc_24 VNB N_A_c_247_n 0.0146698f $X=-0.19 $Y=-0.245 $X2=1.27 $Y2=1.26
cc_25 VNB N_A_c_248_n 0.0152285f $X=-0.19 $Y=-0.245 $X2=1.345 $Y2=1.185
cc_26 VNB N_A_c_249_n 0.0152356f $X=-0.19 $Y=-0.245 $X2=1.7 $Y2=1.26
cc_27 VNB N_A_c_250_n 0.0152356f $X=-0.19 $Y=-0.245 $X2=2.08 $Y2=2.4
cc_28 VNB N_A_c_251_n 0.0197869f $X=-0.19 $Y=-0.245 $X2=2.58 $Y2=2.4
cc_29 VNB N_A_c_252_n 0.0197799f $X=-0.19 $Y=-0.245 $X2=3.425 $Y2=1.35
cc_30 VNB N_A_c_253_n 0.0217216f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_c_254_n 0.00467678f $X=-0.19 $Y=-0.245 $X2=3.93 $Y2=1.65
cc_32 VNB A 6.48016e-19 $X=-0.19 $Y=-0.245 $X2=4.77 $Y2=2.4
cc_33 VNB N_A_c_256_n 0.0459053f $X=-0.19 $Y=-0.245 $X2=2.555 $Y2=1.58
cc_34 VNB N_A_c_257_n 0.112077f $X=-0.19 $Y=-0.245 $X2=3.035 $Y2=1.58
cc_35 VNB N_A_c_258_n 0.0502095f $X=-0.19 $Y=-0.245 $X2=3.765 $Y2=1.515
cc_36 VNB N_A_c_259_n 0.00311164f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_VPWR_c_361_n 0.342803f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_Y_c_442_n 0.0188945f $X=-0.19 $Y=-0.245 $X2=3.515 $Y2=1.58
cc_39 VNB N_Y_c_443_n 2.67464e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB Y 0.00540171f $X=-0.19 $Y=-0.245 $X2=2.58 $Y2=1.475
cc_41 VNB N_A_27_74#_c_551_n 0.033291f $X=-0.19 $Y=-0.245 $X2=2.955 $Y2=0.74
cc_42 VNB N_A_27_74#_c_552_n 0.0225159f $X=-0.19 $Y=-0.245 $X2=3.425 $Y2=1.35
cc_43 VNB N_A_27_74#_c_553_n 0.0187985f $X=-0.19 $Y=-0.245 $X2=3.425 $Y2=0.74
cc_44 VNB N_A_27_74#_c_554_n 0.00195975f $X=-0.19 $Y=-0.245 $X2=3.855 $Y2=1.35
cc_45 VNB N_A_27_74#_c_555_n 0.00740264f $X=-0.19 $Y=-0.245 $X2=3.855 $Y2=0.74
cc_46 VNB N_A_27_74#_c_556_n 0.00215184f $X=-0.19 $Y=-0.245 $X2=4.32 $Y2=1.765
cc_47 VNB N_A_27_74#_c_557_n 0.00512257f $X=-0.19 $Y=-0.245 $X2=4.32 $Y2=2.4
cc_48 VNB N_A_27_74#_c_558_n 0.00815104f $X=-0.19 $Y=-0.245 $X2=4.68 $Y2=1.65
cc_49 VNB N_A_27_74#_c_559_n 0.0023332f $X=-0.19 $Y=-0.245 $X2=4.77 $Y2=2.4
cc_50 VNB N_A_27_74#_c_560_n 0.00475718f $X=-0.19 $Y=-0.245 $X2=0.915 $Y2=1.26
cc_51 VNB N_A_27_74#_c_561_n 0.0016059f $X=-0.19 $Y=-0.245 $X2=4.32 $Y2=1.67
cc_52 VNB N_A_27_74#_c_562_n 0.0339639f $X=-0.19 $Y=-0.245 $X2=2.08 $Y2=1.475
cc_53 VNB N_A_27_74#_c_563_n 0.00367598f $X=-0.19 $Y=-0.245 $X2=2.21 $Y2=1.475
cc_54 VNB N_A_27_74#_c_564_n 0.00170472f $X=-0.19 $Y=-0.245 $X2=2.21 $Y2=1.515
cc_55 VNB N_VGND_c_655_n 0.00323505f $X=-0.19 $Y=-0.245 $X2=1.42 $Y2=1.26
cc_56 VNB N_VGND_c_656_n 0.002601f $X=-0.19 $Y=-0.245 $X2=2.08 $Y2=1.765
cc_57 VNB N_VGND_c_657_n 0.00753502f $X=-0.19 $Y=-0.245 $X2=2.205 $Y2=0.74
cc_58 VNB N_VGND_c_658_n 0.00329129f $X=-0.19 $Y=-0.245 $X2=2.58 $Y2=2.4
cc_59 VNB N_VGND_c_659_n 0.0150174f $X=-0.19 $Y=-0.245 $X2=2.955 $Y2=0.74
cc_60 VNB N_VGND_c_660_n 0.00604233f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_VGND_c_661_n 0.0170727f $X=-0.19 $Y=-0.245 $X2=3.425 $Y2=0.74
cc_62 VNB N_VGND_c_662_n 0.0168561f $X=-0.19 $Y=-0.245 $X2=4.32 $Y2=2.4
cc_63 VNB N_VGND_c_663_n 0.0159778f $X=-0.19 $Y=-0.245 $X2=4.77 $Y2=1.765
cc_64 VNB N_VGND_c_664_n 0.108913f $X=-0.19 $Y=-0.245 $X2=3.995 $Y2=1.58
cc_65 VNB N_VGND_c_665_n 0.432249f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_VGND_c_666_n 0.00604233f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_VGND_c_667_n 0.0109666f $X=-0.19 $Y=-0.245 $X2=2.08 $Y2=1.475
cc_68 VNB N_VGND_c_668_n 0.00604233f $X=-0.19 $Y=-0.245 $X2=2.21 $Y2=1.515
cc_69 VPB N_B_c_127_n 0.0185936f $X=-0.19 $Y=1.66 $X2=2.08 $Y2=1.765
cc_70 VPB N_B_c_128_n 0.0192409f $X=-0.19 $Y=1.66 $X2=2.58 $Y2=1.765
cc_71 VPB N_B_c_120_n 0.010401f $X=-0.19 $Y=1.66 $X2=4.23 $Y2=1.65
cc_72 VPB N_B_c_121_n 0.0699657f $X=-0.19 $Y=1.66 $X2=3.93 $Y2=1.65
cc_73 VPB N_B_c_131_n 0.017597f $X=-0.19 $Y=1.66 $X2=4.32 $Y2=1.765
cc_74 VPB N_B_c_122_n 0.0187089f $X=-0.19 $Y=1.66 $X2=4.68 $Y2=1.65
cc_75 VPB N_B_c_133_n 0.0174155f $X=-0.19 $Y=1.66 $X2=4.77 $Y2=1.765
cc_76 VPB N_B_c_125_n 0.00415909f $X=-0.19 $Y=1.66 $X2=4.32 $Y2=1.67
cc_77 VPB B 0.0179641f $X=-0.19 $Y=1.66 $X2=3.995 $Y2=1.58
cc_78 VPB N_A_c_260_n 0.0181247f $X=-0.19 $Y=1.66 $X2=1.775 $Y2=0.74
cc_79 VPB N_A_c_261_n 0.0174593f $X=-0.19 $Y=1.66 $X2=2.205 $Y2=0.74
cc_80 VPB N_A_c_262_n 0.0170613f $X=-0.19 $Y=1.66 $X2=2.955 $Y2=0.74
cc_81 VPB N_A_c_263_n 0.0177119f $X=-0.19 $Y=1.66 $X2=3.855 $Y2=0.74
cc_82 VPB A 0.00956512f $X=-0.19 $Y=1.66 $X2=4.77 $Y2=2.4
cc_83 VPB N_A_c_257_n 0.0166689f $X=-0.19 $Y=1.66 $X2=3.035 $Y2=1.58
cc_84 VPB N_A_c_258_n 0.0142296f $X=-0.19 $Y=1.66 $X2=3.765 $Y2=1.515
cc_85 VPB N_A_c_267_n 0.00398873f $X=-0.19 $Y=1.66 $X2=2.16 $Y2=1.565
cc_86 VPB N_VPWR_c_362_n 0.0203575f $X=-0.19 $Y=1.66 $X2=2.58 $Y2=1.765
cc_87 VPB N_VPWR_c_363_n 0.00725542f $X=-0.19 $Y=1.66 $X2=2.955 $Y2=0.74
cc_88 VPB N_VPWR_c_364_n 0.0181714f $X=-0.19 $Y=1.66 $X2=3.425 $Y2=0.74
cc_89 VPB N_VPWR_c_365_n 0.0185368f $X=-0.19 $Y=1.66 $X2=3.855 $Y2=0.74
cc_90 VPB N_VPWR_c_366_n 0.00610173f $X=-0.19 $Y=1.66 $X2=3.93 $Y2=1.65
cc_91 VPB N_VPWR_c_367_n 0.0118511f $X=-0.19 $Y=1.66 $X2=4.32 $Y2=2.4
cc_92 VPB N_VPWR_c_368_n 0.0359639f $X=-0.19 $Y=1.66 $X2=4.68 $Y2=1.65
cc_93 VPB N_VPWR_c_369_n 0.0186948f $X=-0.19 $Y=1.66 $X2=4.77 $Y2=2.4
cc_94 VPB N_VPWR_c_370_n 0.0159778f $X=-0.19 $Y=1.66 $X2=2.555 $Y2=1.58
cc_95 VPB N_VPWR_c_371_n 0.0901451f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_96 VPB N_VPWR_c_372_n 0.0231771f $X=-0.19 $Y=1.66 $X2=2.21 $Y2=1.515
cc_97 VPB N_VPWR_c_373_n 0.0185677f $X=-0.19 $Y=1.66 $X2=3.765 $Y2=1.515
cc_98 VPB N_VPWR_c_374_n 0.0483246f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_99 VPB N_VPWR_c_375_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_100 VPB N_VPWR_c_376_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_101 VPB N_VPWR_c_377_n 0.0132702f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_102 VPB N_VPWR_c_361_n 0.0975268f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_103 VPB N_Y_c_445_n 0.00289633f $X=-0.19 $Y=1.66 $X2=2.58 $Y2=2.4
cc_104 VPB N_Y_c_446_n 0.00257348f $X=-0.19 $Y=1.66 $X2=3.425 $Y2=0.74
cc_105 VPB N_Y_c_447_n 0.00289722f $X=-0.19 $Y=1.66 $X2=4.68 $Y2=1.65
cc_106 VPB N_Y_c_448_n 0.00233217f $X=-0.19 $Y=1.66 $X2=1.345 $Y2=1.26
cc_107 VPB N_Y_c_442_n 0.00618364f $X=-0.19 $Y=1.66 $X2=3.515 $Y2=1.58
cc_108 N_B_M1017_g N_A_c_243_n 0.0188633f $X=3.855 $Y=0.74 $X2=-0.19 $Y2=-0.245
cc_109 N_B_c_125_n N_A_c_244_n 0.0132758f $X=4.32 $Y=1.67 $X2=0 $Y2=0
cc_110 N_B_c_120_n N_A_c_245_n 0.0132758f $X=4.23 $Y=1.65 $X2=0 $Y2=0
cc_111 N_B_c_122_n N_A_c_254_n 0.0132758f $X=4.68 $Y=1.65 $X2=0 $Y2=0
cc_112 N_B_c_133_n N_VPWR_c_362_n 0.0261473f $X=4.77 $Y=1.765 $X2=0 $Y2=0
cc_113 N_B_c_131_n N_VPWR_c_369_n 0.00445602f $X=4.32 $Y=1.765 $X2=0 $Y2=0
cc_114 N_B_c_133_n N_VPWR_c_369_n 0.00445602f $X=4.77 $Y=1.765 $X2=0 $Y2=0
cc_115 N_B_c_109_n N_VPWR_c_371_n 0.00736641f $X=0.84 $Y=1.26 $X2=0 $Y2=0
cc_116 N_B_c_127_n N_VPWR_c_371_n 0.00399658f $X=2.08 $Y=1.765 $X2=0 $Y2=0
cc_117 N_B_c_121_n N_VPWR_c_371_n 0.00287171f $X=3.93 $Y=1.65 $X2=0 $Y2=0
cc_118 N_B_c_127_n N_VPWR_c_373_n 0.00445602f $X=2.08 $Y=1.765 $X2=0 $Y2=0
cc_119 N_B_c_128_n N_VPWR_c_373_n 0.00413917f $X=2.58 $Y=1.765 $X2=0 $Y2=0
cc_120 N_B_c_127_n N_VPWR_c_374_n 5.03529e-19 $X=2.08 $Y=1.765 $X2=0 $Y2=0
cc_121 N_B_c_128_n N_VPWR_c_374_n 0.0123325f $X=2.58 $Y=1.765 $X2=0 $Y2=0
cc_122 N_B_c_131_n N_VPWR_c_374_n 0.00400188f $X=4.32 $Y=1.765 $X2=0 $Y2=0
cc_123 N_B_c_127_n N_VPWR_c_361_n 0.0086218f $X=2.08 $Y=1.765 $X2=0 $Y2=0
cc_124 N_B_c_128_n N_VPWR_c_361_n 0.00813572f $X=2.58 $Y=1.765 $X2=0 $Y2=0
cc_125 N_B_c_131_n N_VPWR_c_361_n 0.00861697f $X=4.32 $Y=1.765 $X2=0 $Y2=0
cc_126 N_B_c_133_n N_VPWR_c_361_n 0.00861719f $X=4.77 $Y=1.765 $X2=0 $Y2=0
cc_127 N_B_c_127_n N_Y_c_450_n 0.0019041f $X=2.08 $Y=1.765 $X2=0 $Y2=0
cc_128 N_B_c_121_n N_Y_c_450_n 0.00186359f $X=3.93 $Y=1.65 $X2=0 $Y2=0
cc_129 B N_Y_c_450_n 0.0254779f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_130 N_B_c_127_n N_Y_c_445_n 0.00892941f $X=2.08 $Y=1.765 $X2=0 $Y2=0
cc_131 N_B_c_128_n N_Y_c_445_n 0.00464012f $X=2.58 $Y=1.765 $X2=0 $Y2=0
cc_132 N_B_c_128_n N_Y_c_455_n 0.0170494f $X=2.58 $Y=1.765 $X2=0 $Y2=0
cc_133 N_B_c_121_n N_Y_c_455_n 0.00911022f $X=3.93 $Y=1.65 $X2=0 $Y2=0
cc_134 N_B_c_131_n N_Y_c_455_n 0.0146467f $X=4.32 $Y=1.765 $X2=0 $Y2=0
cc_135 B N_Y_c_455_n 0.132799f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_136 N_B_c_131_n N_Y_c_446_n 0.0150947f $X=4.32 $Y=1.765 $X2=0 $Y2=0
cc_137 N_B_c_133_n N_Y_c_446_n 0.0095765f $X=4.77 $Y=1.765 $X2=0 $Y2=0
cc_138 N_B_c_122_n N_Y_c_461_n 6.66008e-19 $X=4.68 $Y=1.65 $X2=0 $Y2=0
cc_139 N_B_c_125_n N_Y_c_443_n 4.84695e-19 $X=4.32 $Y=1.67 $X2=0 $Y2=0
cc_140 N_B_c_131_n N_Y_c_463_n 2.24111e-19 $X=4.32 $Y=1.765 $X2=0 $Y2=0
cc_141 N_B_c_133_n N_Y_c_463_n 0.00170116f $X=4.77 $Y=1.765 $X2=0 $Y2=0
cc_142 N_B_M1017_g Y 0.00110836f $X=3.855 $Y=0.74 $X2=0 $Y2=0
cc_143 N_B_c_121_n Y 9.13145e-19 $X=3.93 $Y=1.65 $X2=0 $Y2=0
cc_144 N_B_c_131_n Y 0.00829499f $X=4.32 $Y=1.765 $X2=0 $Y2=0
cc_145 N_B_c_122_n Y 0.0224983f $X=4.68 $Y=1.65 $X2=0 $Y2=0
cc_146 N_B_c_133_n Y 0.0045128f $X=4.77 $Y=1.765 $X2=0 $Y2=0
cc_147 N_B_c_125_n Y 0.00422517f $X=4.32 $Y=1.67 $X2=0 $Y2=0
cc_148 B Y 0.0340849f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_149 N_B_c_108_n N_A_27_74#_c_551_n 0.00378532f $X=0.485 $Y=1.185 $X2=0 $Y2=0
cc_150 N_B_c_108_n N_A_27_74#_c_552_n 0.00680723f $X=0.485 $Y=1.185 $X2=0 $Y2=0
cc_151 N_B_c_109_n N_A_27_74#_c_552_n 0.00930473f $X=0.84 $Y=1.26 $X2=0 $Y2=0
cc_152 N_B_c_110_n N_A_27_74#_c_552_n 0.00728337f $X=0.56 $Y=1.26 $X2=0 $Y2=0
cc_153 N_B_c_111_n N_A_27_74#_c_552_n 0.00665856f $X=0.915 $Y=1.185 $X2=0 $Y2=0
cc_154 N_B_c_112_n N_A_27_74#_c_552_n 0.00121915f $X=1.27 $Y=1.26 $X2=0 $Y2=0
cc_155 N_B_c_123_n N_A_27_74#_c_552_n 0.00425286f $X=0.915 $Y=1.26 $X2=0 $Y2=0
cc_156 N_B_c_111_n N_A_27_74#_c_554_n 3.99083e-19 $X=0.915 $Y=1.185 $X2=0 $Y2=0
cc_157 N_B_c_113_n N_A_27_74#_c_554_n 3.99083e-19 $X=1.345 $Y=1.185 $X2=0 $Y2=0
cc_158 N_B_c_112_n N_A_27_74#_c_555_n 0.00121915f $X=1.27 $Y=1.26 $X2=0 $Y2=0
cc_159 N_B_c_113_n N_A_27_74#_c_555_n 0.0115179f $X=1.345 $Y=1.185 $X2=0 $Y2=0
cc_160 N_B_c_114_n N_A_27_74#_c_555_n 0.00932825f $X=1.7 $Y=1.26 $X2=0 $Y2=0
cc_161 N_B_c_124_n N_A_27_74#_c_555_n 0.00425286f $X=1.345 $Y=1.26 $X2=0 $Y2=0
cc_162 N_B_c_115_n N_A_27_74#_c_556_n 4.03226e-19 $X=1.775 $Y=1.185 $X2=0 $Y2=0
cc_163 N_B_c_116_n N_A_27_74#_c_556_n 0.0133277f $X=2.205 $Y=1.185 $X2=0 $Y2=0
cc_164 N_B_c_116_n N_A_27_74#_c_557_n 0.0124731f $X=2.205 $Y=1.185 $X2=0 $Y2=0
cc_165 N_B_M1012_g N_A_27_74#_c_557_n 0.0145095f $X=2.955 $Y=0.74 $X2=0 $Y2=0
cc_166 N_B_c_121_n N_A_27_74#_c_557_n 0.0101838f $X=3.93 $Y=1.65 $X2=0 $Y2=0
cc_167 B N_A_27_74#_c_557_n 0.0694732f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_168 N_B_c_114_n N_A_27_74#_c_558_n 3.12166e-19 $X=1.7 $Y=1.26 $X2=0 $Y2=0
cc_169 N_B_c_115_n N_A_27_74#_c_558_n 0.0116485f $X=1.775 $Y=1.185 $X2=0 $Y2=0
cc_170 N_B_c_116_n N_A_27_74#_c_558_n 0.00169705f $X=2.205 $Y=1.185 $X2=0 $Y2=0
cc_171 N_B_c_121_n N_A_27_74#_c_558_n 0.0180404f $X=3.93 $Y=1.65 $X2=0 $Y2=0
cc_172 B N_A_27_74#_c_558_n 0.00933702f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_173 N_B_M1012_g N_A_27_74#_c_559_n 4.44013e-19 $X=2.955 $Y=0.74 $X2=0 $Y2=0
cc_174 N_B_M1016_g N_A_27_74#_c_559_n 4.44013e-19 $X=3.425 $Y=0.74 $X2=0 $Y2=0
cc_175 N_B_M1016_g N_A_27_74#_c_560_n 0.0131399f $X=3.425 $Y=0.74 $X2=0 $Y2=0
cc_176 N_B_M1017_g N_A_27_74#_c_560_n 0.0128967f $X=3.855 $Y=0.74 $X2=0 $Y2=0
cc_177 N_B_c_120_n N_A_27_74#_c_560_n 0.00104959f $X=4.23 $Y=1.65 $X2=0 $Y2=0
cc_178 N_B_c_121_n N_A_27_74#_c_560_n 0.00230191f $X=3.93 $Y=1.65 $X2=0 $Y2=0
cc_179 B N_A_27_74#_c_560_n 0.0665294f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_180 N_B_c_111_n N_A_27_74#_c_563_n 0.00173424f $X=0.915 $Y=1.185 $X2=0 $Y2=0
cc_181 N_B_c_112_n N_A_27_74#_c_563_n 0.00780096f $X=1.27 $Y=1.26 $X2=0 $Y2=0
cc_182 N_B_c_121_n N_A_27_74#_c_564_n 0.00334528f $X=3.93 $Y=1.65 $X2=0 $Y2=0
cc_183 B N_A_27_74#_c_564_n 0.0197568f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_184 N_B_c_108_n N_VGND_c_655_n 0.0141343f $X=0.485 $Y=1.185 $X2=0 $Y2=0
cc_185 N_B_c_109_n N_VGND_c_655_n 7.59159e-19 $X=0.84 $Y=1.26 $X2=0 $Y2=0
cc_186 N_B_c_111_n N_VGND_c_655_n 0.0108532f $X=0.915 $Y=1.185 $X2=0 $Y2=0
cc_187 N_B_c_113_n N_VGND_c_655_n 5.07887e-19 $X=1.345 $Y=1.185 $X2=0 $Y2=0
cc_188 N_B_c_111_n N_VGND_c_656_n 4.64036e-19 $X=0.915 $Y=1.185 $X2=0 $Y2=0
cc_189 N_B_c_113_n N_VGND_c_656_n 0.010563f $X=1.345 $Y=1.185 $X2=0 $Y2=0
cc_190 N_B_c_114_n N_VGND_c_656_n 5.31749e-19 $X=1.7 $Y=1.26 $X2=0 $Y2=0
cc_191 N_B_c_115_n N_VGND_c_656_n 0.0106828f $X=1.775 $Y=1.185 $X2=0 $Y2=0
cc_192 N_B_c_116_n N_VGND_c_656_n 5.10222e-19 $X=2.205 $Y=1.185 $X2=0 $Y2=0
cc_193 N_B_c_116_n N_VGND_c_657_n 0.00351545f $X=2.205 $Y=1.185 $X2=0 $Y2=0
cc_194 N_B_M1012_g N_VGND_c_657_n 0.01382f $X=2.955 $Y=0.74 $X2=0 $Y2=0
cc_195 N_B_M1016_g N_VGND_c_657_n 4.5623e-19 $X=3.425 $Y=0.74 $X2=0 $Y2=0
cc_196 N_B_M1012_g N_VGND_c_658_n 4.58633e-19 $X=2.955 $Y=0.74 $X2=0 $Y2=0
cc_197 N_B_M1016_g N_VGND_c_658_n 0.010342f $X=3.425 $Y=0.74 $X2=0 $Y2=0
cc_198 N_B_M1017_g N_VGND_c_658_n 0.0104354f $X=3.855 $Y=0.74 $X2=0 $Y2=0
cc_199 N_B_c_111_n N_VGND_c_659_n 0.00383152f $X=0.915 $Y=1.185 $X2=0 $Y2=0
cc_200 N_B_c_113_n N_VGND_c_659_n 0.00383152f $X=1.345 $Y=1.185 $X2=0 $Y2=0
cc_201 N_B_c_108_n N_VGND_c_661_n 0.00383152f $X=0.485 $Y=1.185 $X2=0 $Y2=0
cc_202 N_B_c_115_n N_VGND_c_662_n 0.00383152f $X=1.775 $Y=1.185 $X2=0 $Y2=0
cc_203 N_B_c_116_n N_VGND_c_662_n 0.00434272f $X=2.205 $Y=1.185 $X2=0 $Y2=0
cc_204 N_B_M1012_g N_VGND_c_663_n 0.00383152f $X=2.955 $Y=0.74 $X2=0 $Y2=0
cc_205 N_B_M1016_g N_VGND_c_663_n 0.00383152f $X=3.425 $Y=0.74 $X2=0 $Y2=0
cc_206 N_B_M1017_g N_VGND_c_664_n 0.00383152f $X=3.855 $Y=0.74 $X2=0 $Y2=0
cc_207 N_B_c_108_n N_VGND_c_665_n 0.00761163f $X=0.485 $Y=1.185 $X2=0 $Y2=0
cc_208 N_B_c_111_n N_VGND_c_665_n 0.0075754f $X=0.915 $Y=1.185 $X2=0 $Y2=0
cc_209 N_B_c_113_n N_VGND_c_665_n 0.0075754f $X=1.345 $Y=1.185 $X2=0 $Y2=0
cc_210 N_B_c_115_n N_VGND_c_665_n 0.0075754f $X=1.775 $Y=1.185 $X2=0 $Y2=0
cc_211 N_B_c_116_n N_VGND_c_665_n 0.00822462f $X=2.205 $Y=1.185 $X2=0 $Y2=0
cc_212 N_B_M1012_g N_VGND_c_665_n 0.00757927f $X=2.955 $Y=0.74 $X2=0 $Y2=0
cc_213 N_B_M1016_g N_VGND_c_665_n 0.00757927f $X=3.425 $Y=0.74 $X2=0 $Y2=0
cc_214 N_B_M1017_g N_VGND_c_665_n 0.00757637f $X=3.855 $Y=0.74 $X2=0 $Y2=0
cc_215 N_A_c_247_n N_VPWR_c_362_n 0.010031f $X=5.07 $Y=1.26 $X2=0 $Y2=0
cc_216 N_A_c_257_n N_VPWR_c_362_n 6.1376e-19 $X=6.51 $Y=1.385 $X2=0 $Y2=0
cc_217 N_A_c_259_n N_VPWR_c_362_n 0.00143398f $X=5.965 $Y=1.5 $X2=0 $Y2=0
cc_218 N_A_c_260_n N_VPWR_c_364_n 0.0265292f $X=5.88 $Y=1.765 $X2=0 $Y2=0
cc_219 N_A_c_257_n N_VPWR_c_364_n 0.00829757f $X=6.51 $Y=1.385 $X2=0 $Y2=0
cc_220 N_A_c_259_n N_VPWR_c_364_n 0.0195977f $X=5.965 $Y=1.5 $X2=0 $Y2=0
cc_221 N_A_c_260_n N_VPWR_c_365_n 0.00445602f $X=5.88 $Y=1.765 $X2=0 $Y2=0
cc_222 N_A_c_261_n N_VPWR_c_365_n 0.00413917f $X=6.38 $Y=1.765 $X2=0 $Y2=0
cc_223 N_A_c_260_n N_VPWR_c_366_n 5.03756e-19 $X=5.88 $Y=1.765 $X2=0 $Y2=0
cc_224 N_A_c_261_n N_VPWR_c_366_n 0.0129143f $X=6.38 $Y=1.765 $X2=0 $Y2=0
cc_225 N_A_c_262_n N_VPWR_c_366_n 0.0126657f $X=7.21 $Y=1.765 $X2=0 $Y2=0
cc_226 N_A_c_263_n N_VPWR_c_366_n 5.02157e-19 $X=7.66 $Y=1.765 $X2=0 $Y2=0
cc_227 N_A_c_262_n N_VPWR_c_368_n 5.06484e-19 $X=7.21 $Y=1.765 $X2=0 $Y2=0
cc_228 N_A_c_263_n N_VPWR_c_368_n 0.0124858f $X=7.66 $Y=1.765 $X2=0 $Y2=0
cc_229 N_A_c_262_n N_VPWR_c_370_n 0.00413917f $X=7.21 $Y=1.765 $X2=0 $Y2=0
cc_230 N_A_c_263_n N_VPWR_c_370_n 0.00413917f $X=7.66 $Y=1.765 $X2=0 $Y2=0
cc_231 N_A_c_260_n N_VPWR_c_361_n 0.0086218f $X=5.88 $Y=1.765 $X2=0 $Y2=0
cc_232 N_A_c_261_n N_VPWR_c_361_n 0.00818187f $X=6.38 $Y=1.765 $X2=0 $Y2=0
cc_233 N_A_c_262_n N_VPWR_c_361_n 0.00817726f $X=7.21 $Y=1.765 $X2=0 $Y2=0
cc_234 N_A_c_263_n N_VPWR_c_361_n 0.00817726f $X=7.66 $Y=1.765 $X2=0 $Y2=0
cc_235 N_A_c_245_n N_Y_c_455_n 5.0821e-19 $X=4.36 $Y=1.26 $X2=0 $Y2=0
cc_236 N_A_c_246_n N_Y_c_461_n 0.00793829f $X=4.715 $Y=1.185 $X2=0 $Y2=0
cc_237 N_A_c_247_n N_Y_c_461_n 0.00377529f $X=5.07 $Y=1.26 $X2=0 $Y2=0
cc_238 N_A_c_248_n N_Y_c_461_n 0.0146292f $X=5.145 $Y=1.185 $X2=0 $Y2=0
cc_239 N_A_c_249_n N_Y_c_461_n 0.0113799f $X=5.575 $Y=1.185 $X2=0 $Y2=0
cc_240 N_A_c_250_n N_Y_c_461_n 0.0113799f $X=6.005 $Y=1.185 $X2=0 $Y2=0
cc_241 N_A_c_251_n N_Y_c_461_n 0.013733f $X=6.435 $Y=1.22 $X2=0 $Y2=0
cc_242 N_A_c_252_n N_Y_c_461_n 0.013733f $X=7.225 $Y=1.22 $X2=0 $Y2=0
cc_243 N_A_c_253_n N_Y_c_461_n 0.0175893f $X=7.655 $Y=1.22 $X2=0 $Y2=0
cc_244 N_A_c_256_n N_Y_c_461_n 0.0105545f $X=7.12 $Y=1.385 $X2=0 $Y2=0
cc_245 N_A_c_257_n N_Y_c_461_n 0.00753416f $X=6.51 $Y=1.385 $X2=0 $Y2=0
cc_246 N_A_c_258_n N_Y_c_461_n 0.00230817f $X=7.655 $Y=1.492 $X2=0 $Y2=0
cc_247 N_A_c_259_n N_Y_c_461_n 0.163412f $X=5.965 $Y=1.5 $X2=0 $Y2=0
cc_248 N_A_c_260_n N_Y_c_485_n 0.00202688f $X=5.88 $Y=1.765 $X2=0 $Y2=0
cc_249 N_A_c_257_n N_Y_c_485_n 6.5509e-19 $X=6.51 $Y=1.385 $X2=0 $Y2=0
cc_250 N_A_c_267_n N_Y_c_485_n 0.0244044f $X=6.525 $Y=1.5 $X2=0 $Y2=0
cc_251 N_A_c_259_n N_Y_c_485_n 7.48087e-19 $X=5.965 $Y=1.5 $X2=0 $Y2=0
cc_252 N_A_c_260_n N_Y_c_447_n 0.00892941f $X=5.88 $Y=1.765 $X2=0 $Y2=0
cc_253 N_A_c_261_n N_Y_c_447_n 0.00464047f $X=6.38 $Y=1.765 $X2=0 $Y2=0
cc_254 N_A_c_261_n N_Y_c_491_n 0.0165498f $X=6.38 $Y=1.765 $X2=0 $Y2=0
cc_255 N_A_c_262_n N_Y_c_491_n 0.0140762f $X=7.21 $Y=1.765 $X2=0 $Y2=0
cc_256 N_A_c_256_n N_Y_c_491_n 0.00195464f $X=7.12 $Y=1.385 $X2=0 $Y2=0
cc_257 N_A_c_267_n N_Y_c_491_n 0.0766712f $X=6.525 $Y=1.5 $X2=0 $Y2=0
cc_258 N_A_c_263_n N_Y_c_495_n 0.0176683f $X=7.66 $Y=1.765 $X2=0 $Y2=0
cc_259 N_A_c_262_n N_Y_c_442_n 5.80272e-19 $X=7.21 $Y=1.765 $X2=0 $Y2=0
cc_260 N_A_c_252_n N_Y_c_442_n 6.84216e-19 $X=7.225 $Y=1.22 $X2=0 $Y2=0
cc_261 N_A_c_253_n N_Y_c_442_n 0.00559507f $X=7.655 $Y=1.22 $X2=0 $Y2=0
cc_262 N_A_c_263_n N_Y_c_442_n 0.00610216f $X=7.66 $Y=1.765 $X2=0 $Y2=0
cc_263 A N_Y_c_442_n 0.043501f $X=7.355 $Y=1.58 $X2=0 $Y2=0
cc_264 N_A_c_258_n N_Y_c_442_n 0.0178746f $X=7.655 $Y=1.492 $X2=0 $Y2=0
cc_265 N_A_c_243_n N_Y_c_443_n 0.00472298f $X=4.285 $Y=1.185 $X2=0 $Y2=0
cc_266 N_A_c_246_n N_Y_c_443_n 0.00480024f $X=4.715 $Y=1.185 $X2=0 $Y2=0
cc_267 N_A_c_248_n N_Y_c_443_n 4.25175e-19 $X=5.145 $Y=1.185 $X2=0 $Y2=0
cc_268 A N_Y_c_505_n 0.0187638f $X=7.355 $Y=1.58 $X2=0 $Y2=0
cc_269 N_A_c_258_n N_Y_c_505_n 4.24887e-19 $X=7.655 $Y=1.492 $X2=0 $Y2=0
cc_270 N_A_c_243_n Y 5.82771e-19 $X=4.285 $Y=1.185 $X2=0 $Y2=0
cc_271 N_A_c_244_n Y 0.0110261f $X=4.64 $Y=1.26 $X2=0 $Y2=0
cc_272 N_A_c_246_n Y 0.00162787f $X=4.715 $Y=1.185 $X2=0 $Y2=0
cc_273 N_A_c_248_n Y 2.83995e-19 $X=5.145 $Y=1.185 $X2=0 $Y2=0
cc_274 N_A_c_254_n Y 0.00623952f $X=4.715 $Y=1.26 $X2=0 $Y2=0
cc_275 N_A_c_257_n Y 0.00128584f $X=6.51 $Y=1.385 $X2=0 $Y2=0
cc_276 N_A_c_259_n Y 0.0122173f $X=5.965 $Y=1.5 $X2=0 $Y2=0
cc_277 N_A_c_243_n N_A_27_74#_c_560_n 6.21217e-19 $X=4.285 $Y=1.185 $X2=0 $Y2=0
cc_278 N_A_c_243_n N_A_27_74#_c_562_n 0.0141739f $X=4.285 $Y=1.185 $X2=0 $Y2=0
cc_279 N_A_c_244_n N_A_27_74#_c_562_n 3.13775e-19 $X=4.64 $Y=1.26 $X2=0 $Y2=0
cc_280 N_A_c_246_n N_A_27_74#_c_562_n 0.0101463f $X=4.715 $Y=1.185 $X2=0 $Y2=0
cc_281 N_A_c_248_n N_A_27_74#_c_562_n 0.010218f $X=5.145 $Y=1.185 $X2=0 $Y2=0
cc_282 N_A_c_249_n N_A_27_74#_c_562_n 0.010218f $X=5.575 $Y=1.185 $X2=0 $Y2=0
cc_283 N_A_c_250_n N_A_27_74#_c_562_n 0.010218f $X=6.005 $Y=1.185 $X2=0 $Y2=0
cc_284 N_A_c_251_n N_A_27_74#_c_562_n 0.0103703f $X=6.435 $Y=1.22 $X2=0 $Y2=0
cc_285 N_A_c_252_n N_A_27_74#_c_562_n 0.0103703f $X=7.225 $Y=1.22 $X2=0 $Y2=0
cc_286 N_A_c_253_n N_A_27_74#_c_562_n 0.0103137f $X=7.655 $Y=1.22 $X2=0 $Y2=0
cc_287 N_A_c_243_n N_VGND_c_658_n 6.35276e-19 $X=4.285 $Y=1.185 $X2=0 $Y2=0
cc_288 N_A_c_243_n N_VGND_c_664_n 0.00291649f $X=4.285 $Y=1.185 $X2=0 $Y2=0
cc_289 N_A_c_246_n N_VGND_c_664_n 0.00291649f $X=4.715 $Y=1.185 $X2=0 $Y2=0
cc_290 N_A_c_248_n N_VGND_c_664_n 0.00291649f $X=5.145 $Y=1.185 $X2=0 $Y2=0
cc_291 N_A_c_249_n N_VGND_c_664_n 0.00291649f $X=5.575 $Y=1.185 $X2=0 $Y2=0
cc_292 N_A_c_250_n N_VGND_c_664_n 0.00291649f $X=6.005 $Y=1.185 $X2=0 $Y2=0
cc_293 N_A_c_251_n N_VGND_c_664_n 0.00291649f $X=6.435 $Y=1.22 $X2=0 $Y2=0
cc_294 N_A_c_252_n N_VGND_c_664_n 0.00291649f $X=7.225 $Y=1.22 $X2=0 $Y2=0
cc_295 N_A_c_253_n N_VGND_c_664_n 0.00291649f $X=7.655 $Y=1.22 $X2=0 $Y2=0
cc_296 N_A_c_243_n N_VGND_c_665_n 0.00359219f $X=4.285 $Y=1.185 $X2=0 $Y2=0
cc_297 N_A_c_246_n N_VGND_c_665_n 0.00359121f $X=4.715 $Y=1.185 $X2=0 $Y2=0
cc_298 N_A_c_248_n N_VGND_c_665_n 0.00359121f $X=5.145 $Y=1.185 $X2=0 $Y2=0
cc_299 N_A_c_249_n N_VGND_c_665_n 0.00359121f $X=5.575 $Y=1.185 $X2=0 $Y2=0
cc_300 N_A_c_250_n N_VGND_c_665_n 0.00359121f $X=6.005 $Y=1.185 $X2=0 $Y2=0
cc_301 N_A_c_251_n N_VGND_c_665_n 0.00361732f $X=6.435 $Y=1.22 $X2=0 $Y2=0
cc_302 N_A_c_252_n N_VGND_c_665_n 0.00361732f $X=7.225 $Y=1.22 $X2=0 $Y2=0
cc_303 N_A_c_253_n N_VGND_c_665_n 0.00362813f $X=7.655 $Y=1.22 $X2=0 $Y2=0
cc_304 N_VPWR_c_371_n N_Y_c_445_n 0.0331138f $X=1.165 $Y=2.115 $X2=0 $Y2=0
cc_305 N_VPWR_c_373_n N_Y_c_445_n 0.0145938f $X=2.64 $Y=2.852 $X2=0 $Y2=0
cc_306 N_VPWR_c_374_n N_Y_c_445_n 0.0298173f $X=4.21 $Y=2.852 $X2=0 $Y2=0
cc_307 N_VPWR_c_361_n N_Y_c_445_n 0.0120466f $X=7.92 $Y=3.33 $X2=0 $Y2=0
cc_308 N_VPWR_M1007_d N_Y_c_455_n 0.0397677f $X=2.655 $Y=1.84 $X2=0 $Y2=0
cc_309 N_VPWR_c_374_n N_Y_c_455_n 0.120654f $X=4.21 $Y=2.852 $X2=0 $Y2=0
cc_310 N_VPWR_c_362_n N_Y_c_446_n 0.0330222f $X=5.045 $Y=1.985 $X2=0 $Y2=0
cc_311 N_VPWR_c_369_n N_Y_c_446_n 0.014552f $X=4.88 $Y=3.33 $X2=0 $Y2=0
cc_312 N_VPWR_c_374_n N_Y_c_446_n 0.0268614f $X=4.21 $Y=2.852 $X2=0 $Y2=0
cc_313 N_VPWR_c_361_n N_Y_c_446_n 0.0119791f $X=7.92 $Y=3.33 $X2=0 $Y2=0
cc_314 N_VPWR_c_364_n N_Y_c_447_n 0.0330222f $X=5.605 $Y=1.985 $X2=0 $Y2=0
cc_315 N_VPWR_c_365_n N_Y_c_447_n 0.0145938f $X=6.44 $Y=3.33 $X2=0 $Y2=0
cc_316 N_VPWR_c_366_n N_Y_c_447_n 0.029897f $X=6.985 $Y=2.375 $X2=0 $Y2=0
cc_317 N_VPWR_c_361_n N_Y_c_447_n 0.0120466f $X=7.92 $Y=3.33 $X2=0 $Y2=0
cc_318 N_VPWR_M1019_s N_Y_c_491_n 0.014315f $X=6.455 $Y=1.84 $X2=0 $Y2=0
cc_319 N_VPWR_c_366_n N_Y_c_491_n 0.0480976f $X=6.985 $Y=2.375 $X2=0 $Y2=0
cc_320 N_VPWR_c_366_n N_Y_c_448_n 0.0298549f $X=6.985 $Y=2.375 $X2=0 $Y2=0
cc_321 N_VPWR_c_368_n N_Y_c_448_n 0.0266389f $X=7.885 $Y=2.375 $X2=0 $Y2=0
cc_322 N_VPWR_c_370_n N_Y_c_448_n 0.0101736f $X=7.72 $Y=3.33 $X2=0 $Y2=0
cc_323 N_VPWR_c_361_n N_Y_c_448_n 0.0084208f $X=7.92 $Y=3.33 $X2=0 $Y2=0
cc_324 N_VPWR_M1021_s N_Y_c_495_n 0.00879754f $X=7.735 $Y=1.84 $X2=0 $Y2=0
cc_325 N_VPWR_c_368_n N_Y_c_495_n 0.0100034f $X=7.885 $Y=2.375 $X2=0 $Y2=0
cc_326 N_VPWR_M1021_s N_Y_c_442_n 0.00415896f $X=7.735 $Y=1.84 $X2=0 $Y2=0
cc_327 N_VPWR_c_362_n Y 0.00563088f $X=5.045 $Y=1.985 $X2=0 $Y2=0
cc_328 N_VPWR_c_371_n N_A_27_74#_c_552_n 0.0125662f $X=1.165 $Y=2.115 $X2=0
+ $Y2=0
cc_329 N_VPWR_c_371_n N_A_27_74#_c_555_n 0.0162232f $X=1.165 $Y=2.115 $X2=0
+ $Y2=0
cc_330 N_VPWR_c_371_n N_A_27_74#_c_558_n 0.00605024f $X=1.165 $Y=2.115 $X2=0
+ $Y2=0
cc_331 N_VPWR_c_371_n N_A_27_74#_c_563_n 0.00704273f $X=1.165 $Y=2.115 $X2=0
+ $Y2=0
cc_332 N_Y_c_461_n N_A_27_74#_M1005_d 0.00533199f $X=7.725 $Y=0.91 $X2=0 $Y2=0
cc_333 N_Y_c_461_n N_A_27_74#_M1009_d 0.00331558f $X=7.725 $Y=0.91 $X2=0 $Y2=0
cc_334 N_Y_c_461_n N_A_27_74#_M1014_d 0.0143874f $X=7.725 $Y=0.91 $X2=0 $Y2=0
cc_335 N_Y_c_461_n N_A_27_74#_M1023_d 0.0138053f $X=7.725 $Y=0.91 $X2=0 $Y2=0
cc_336 N_Y_c_442_n N_A_27_74#_M1023_d 0.00225118f $X=7.81 $Y=1.95 $X2=0 $Y2=0
cc_337 N_Y_c_443_n N_A_27_74#_c_560_n 0.00542281f $X=4.545 $Y=1.13 $X2=0 $Y2=0
cc_338 Y N_A_27_74#_c_560_n 0.00359291f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_339 N_Y_M1004_s N_A_27_74#_c_562_n 0.00168993f $X=4.36 $Y=0.37 $X2=0 $Y2=0
cc_340 N_Y_M1006_s N_A_27_74#_c_562_n 0.00169393f $X=5.22 $Y=0.37 $X2=0 $Y2=0
cc_341 N_Y_M1013_s N_A_27_74#_c_562_n 0.00170263f $X=6.08 $Y=0.37 $X2=0 $Y2=0
cc_342 N_Y_M1018_s N_A_27_74#_c_562_n 0.00170263f $X=7.3 $Y=0.37 $X2=0 $Y2=0
cc_343 N_Y_c_461_n N_A_27_74#_c_562_n 0.178804f $X=7.725 $Y=0.91 $X2=0 $Y2=0
cc_344 N_Y_c_443_n N_A_27_74#_c_562_n 0.0204027f $X=4.545 $Y=1.13 $X2=0 $Y2=0
cc_345 N_A_27_74#_c_555_n N_VGND_M1003_d 0.00180346f $X=1.688 $Y=1.182 $X2=0
+ $Y2=0
cc_346 N_A_27_74#_c_557_n N_VGND_M1011_d 0.0064814f $X=3.075 $Y=1.095 $X2=0
+ $Y2=0
cc_347 N_A_27_74#_c_560_n N_VGND_M1016_d 0.00176461f $X=3.985 $Y=1.095 $X2=0
+ $Y2=0
cc_348 N_A_27_74#_c_551_n N_VGND_c_655_n 0.0238456f $X=0.27 $Y=0.515 $X2=0 $Y2=0
cc_349 N_A_27_74#_c_552_n N_VGND_c_655_n 0.0218173f $X=1.035 $Y=1.26 $X2=0 $Y2=0
cc_350 N_A_27_74#_c_554_n N_VGND_c_655_n 0.024929f $X=1.13 $Y=0.515 $X2=0 $Y2=0
cc_351 N_A_27_74#_c_554_n N_VGND_c_656_n 0.019113f $X=1.13 $Y=0.515 $X2=0 $Y2=0
cc_352 N_A_27_74#_c_555_n N_VGND_c_656_n 0.0160615f $X=1.688 $Y=1.182 $X2=0
+ $Y2=0
cc_353 N_A_27_74#_c_556_n N_VGND_c_656_n 0.0191484f $X=1.99 $Y=0.515 $X2=0 $Y2=0
cc_354 N_A_27_74#_c_558_n N_VGND_c_656_n 0.00188964f $X=2.155 $Y=1.095 $X2=0
+ $Y2=0
cc_355 N_A_27_74#_c_556_n N_VGND_c_657_n 0.0185872f $X=1.99 $Y=0.515 $X2=0 $Y2=0
cc_356 N_A_27_74#_c_557_n N_VGND_c_657_n 0.0413263f $X=3.075 $Y=1.095 $X2=0
+ $Y2=0
cc_357 N_A_27_74#_c_559_n N_VGND_c_657_n 0.0207899f $X=3.19 $Y=0.515 $X2=0 $Y2=0
cc_358 N_A_27_74#_c_559_n N_VGND_c_658_n 0.0191344f $X=3.19 $Y=0.515 $X2=0 $Y2=0
cc_359 N_A_27_74#_c_560_n N_VGND_c_658_n 0.0171619f $X=3.985 $Y=1.095 $X2=0
+ $Y2=0
cc_360 N_A_27_74#_c_561_n N_VGND_c_658_n 0.00985092f $X=4.07 $Y=0.6 $X2=0 $Y2=0
cc_361 N_A_27_74#_c_554_n N_VGND_c_659_n 0.00838873f $X=1.13 $Y=0.515 $X2=0
+ $Y2=0
cc_362 N_A_27_74#_c_551_n N_VGND_c_661_n 0.011066f $X=0.27 $Y=0.515 $X2=0 $Y2=0
cc_363 N_A_27_74#_c_556_n N_VGND_c_662_n 0.0114405f $X=1.99 $Y=0.515 $X2=0 $Y2=0
cc_364 N_A_27_74#_c_559_n N_VGND_c_663_n 0.0101736f $X=3.19 $Y=0.515 $X2=0 $Y2=0
cc_365 N_A_27_74#_c_561_n N_VGND_c_664_n 0.00758556f $X=4.07 $Y=0.6 $X2=0 $Y2=0
cc_366 N_A_27_74#_c_562_n N_VGND_c_664_n 0.157922f $X=7.875 $Y=0.515 $X2=0 $Y2=0
cc_367 N_A_27_74#_c_551_n N_VGND_c_665_n 0.00915947f $X=0.27 $Y=0.515 $X2=0
+ $Y2=0
cc_368 N_A_27_74#_c_554_n N_VGND_c_665_n 0.00694347f $X=1.13 $Y=0.515 $X2=0
+ $Y2=0
cc_369 N_A_27_74#_c_556_n N_VGND_c_665_n 0.00941304f $X=1.99 $Y=0.515 $X2=0
+ $Y2=0
cc_370 N_A_27_74#_c_559_n N_VGND_c_665_n 0.0084208f $X=3.19 $Y=0.515 $X2=0 $Y2=0
cc_371 N_A_27_74#_c_561_n N_VGND_c_665_n 0.00627867f $X=4.07 $Y=0.6 $X2=0 $Y2=0
cc_372 N_A_27_74#_c_562_n N_VGND_c_665_n 0.133324f $X=7.875 $Y=0.515 $X2=0 $Y2=0
