* File: sky130_fd_sc_hs__nor4b_2.pxi.spice
* Created: Tue Sep  1 20:12:27 2020
* 
x_PM_SKY130_FD_SC_HS__NOR4B_2%D_N N_D_N_c_95_n N_D_N_M1008_g N_D_N_M1002_g D_N
+ PM_SKY130_FD_SC_HS__NOR4B_2%D_N
x_PM_SKY130_FD_SC_HS__NOR4B_2%A_27_392# N_A_27_392#_M1002_s N_A_27_392#_M1008_s
+ N_A_27_392#_c_127_n N_A_27_392#_M1010_g N_A_27_392#_c_135_n
+ N_A_27_392#_M1001_g N_A_27_392#_c_128_n N_A_27_392#_M1011_g
+ N_A_27_392#_c_136_n N_A_27_392#_M1017_g N_A_27_392#_c_129_n
+ N_A_27_392#_c_130_n N_A_27_392#_c_131_n N_A_27_392#_c_132_n
+ N_A_27_392#_c_133_n N_A_27_392#_c_134_n PM_SKY130_FD_SC_HS__NOR4B_2%A_27_392#
x_PM_SKY130_FD_SC_HS__NOR4B_2%C N_C_M1012_g N_C_c_217_n N_C_M1004_g N_C_M1016_g
+ N_C_c_218_n N_C_M1006_g C C N_C_c_216_n PM_SKY130_FD_SC_HS__NOR4B_2%C
x_PM_SKY130_FD_SC_HS__NOR4B_2%B N_B_M1007_g N_B_c_270_n N_B_c_271_n N_B_c_279_n
+ N_B_M1000_g N_B_M1013_g N_B_c_273_n N_B_c_281_n N_B_M1003_g N_B_c_274_n B B
+ N_B_c_276_n PM_SKY130_FD_SC_HS__NOR4B_2%B
x_PM_SKY130_FD_SC_HS__NOR4B_2%A N_A_M1009_g N_A_c_336_n N_A_M1005_g N_A_c_337_n
+ N_A_M1015_g N_A_M1014_g A A A N_A_c_335_n PM_SKY130_FD_SC_HS__NOR4B_2%A
x_PM_SKY130_FD_SC_HS__NOR4B_2%VPWR N_VPWR_M1008_d N_VPWR_M1005_d N_VPWR_c_378_n
+ N_VPWR_c_379_n VPWR N_VPWR_c_380_n N_VPWR_c_381_n N_VPWR_c_382_n
+ N_VPWR_c_377_n N_VPWR_c_384_n N_VPWR_c_385_n PM_SKY130_FD_SC_HS__NOR4B_2%VPWR
x_PM_SKY130_FD_SC_HS__NOR4B_2%A_229_368# N_A_229_368#_M1001_d
+ N_A_229_368#_M1017_d N_A_229_368#_M1006_s N_A_229_368#_c_433_n
+ N_A_229_368#_c_434_n N_A_229_368#_c_435_n N_A_229_368#_c_447_n
+ N_A_229_368#_c_448_n N_A_229_368#_c_436_n N_A_229_368#_c_437_n
+ PM_SKY130_FD_SC_HS__NOR4B_2%A_229_368#
x_PM_SKY130_FD_SC_HS__NOR4B_2%Y N_Y_M1010_s N_Y_M1012_s N_Y_M1007_d N_Y_M1009_s
+ N_Y_M1001_s N_Y_c_481_n N_Y_c_494_n N_Y_c_497_n N_Y_c_490_n N_Y_c_504_n
+ N_Y_c_506_n N_Y_c_482_n N_Y_c_483_n N_Y_c_484_n N_Y_c_485_n N_Y_c_486_n
+ N_Y_c_487_n Y Y N_Y_c_489_n PM_SKY130_FD_SC_HS__NOR4B_2%Y
x_PM_SKY130_FD_SC_HS__NOR4B_2%A_498_368# N_A_498_368#_M1004_d
+ N_A_498_368#_M1000_d N_A_498_368#_c_587_n N_A_498_368#_c_594_n
+ N_A_498_368#_c_588_n PM_SKY130_FD_SC_HS__NOR4B_2%A_498_368#
x_PM_SKY130_FD_SC_HS__NOR4B_2%A_701_368# N_A_701_368#_M1000_s
+ N_A_701_368#_M1003_s N_A_701_368#_M1015_s N_A_701_368#_c_618_n
+ N_A_701_368#_c_619_n N_A_701_368#_c_628_n N_A_701_368#_c_620_n
+ N_A_701_368#_c_635_n N_A_701_368#_c_621_n N_A_701_368#_c_622_n
+ N_A_701_368#_c_641_n PM_SKY130_FD_SC_HS__NOR4B_2%A_701_368#
x_PM_SKY130_FD_SC_HS__NOR4B_2%VGND N_VGND_M1002_d N_VGND_M1011_d N_VGND_M1016_d
+ N_VGND_M1013_s N_VGND_M1014_d N_VGND_c_660_n N_VGND_c_661_n N_VGND_c_662_n
+ N_VGND_c_663_n N_VGND_c_664_n N_VGND_c_665_n VGND N_VGND_c_666_n
+ N_VGND_c_667_n N_VGND_c_668_n N_VGND_c_669_n N_VGND_c_670_n N_VGND_c_671_n
+ N_VGND_c_672_n PM_SKY130_FD_SC_HS__NOR4B_2%VGND
cc_1 VNB N_D_N_c_95_n 0.0264481f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.885
cc_2 VNB N_D_N_M1002_g 0.0450381f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=0.69
cc_3 VNB D_N 0.00165062f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_4 VNB N_A_27_392#_c_127_n 0.0182324f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_5 VNB N_A_27_392#_c_128_n 0.0183095f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_6 VNB N_A_27_392#_c_129_n 0.0390192f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_7 VNB N_A_27_392#_c_130_n 0.0189495f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_A_27_392#_c_131_n 0.0120801f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A_27_392#_c_132_n 0.0081778f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_27_392#_c_133_n 0.014353f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_27_392#_c_134_n 0.0808498f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_C_M1012_g 0.0257645f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.46
cc_13 VNB N_C_M1016_g 0.0249557f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.635
cc_14 VNB C 0.00340543f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_C_c_216_n 0.0337095f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_B_M1007_g 0.026244f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.46
cc_17 VNB N_B_c_270_n 0.0157093f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=0.69
cc_18 VNB N_B_c_271_n 0.00974905f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=0.69
cc_19 VNB N_B_M1013_g 0.0318253f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=1.635
cc_20 VNB N_B_c_273_n 0.0112417f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_B_c_274_n 0.0100834f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB B 0.00579351f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_B_c_276_n 0.0101463f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_M1009_g 0.0305489f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.46
cc_25 VNB N_A_M1014_g 0.0326296f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB A 0.0218856f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_c_335_n 0.0411845f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_VPWR_c_377_n 0.243291f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_Y_c_481_n 0.00291634f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_Y_c_482_n 0.00240191f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_Y_c_483_n 0.00517051f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_Y_c_484_n 0.00687852f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_Y_c_485_n 0.00263681f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_Y_c_486_n 0.0117419f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_Y_c_487_n 0.0028038f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB Y 0.00299091f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_Y_c_489_n 0.00245684f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_660_n 0.00894653f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_661_n 0.00830481f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_662_n 0.0120411f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_663_n 0.0421046f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_664_n 0.0223929f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_665_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_666_n 0.0184653f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_VGND_c_667_n 0.0187266f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_VGND_c_668_n 0.041024f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_VGND_c_669_n 0.0185686f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_VGND_c_670_n 0.0169675f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_VGND_c_671_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_VGND_c_672_n 0.313921f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VPB N_D_N_c_95_n 0.0504893f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.885
cc_52 VPB D_N 0.00249009f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_53 VPB N_A_27_392#_c_135_n 0.0177179f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.635
cc_54 VPB N_A_27_392#_c_136_n 0.0149021f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_55 VPB N_A_27_392#_c_130_n 0.0556875f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_56 VPB N_A_27_392#_c_134_n 0.0138781f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_57 VPB N_C_c_217_n 0.0154078f $X=-0.19 $Y=1.66 $X2=0.63 $Y2=0.69
cc_58 VPB N_C_c_218_n 0.0175567f $X=-0.19 $Y=1.66 $X2=0.7 $Y2=1.635
cc_59 VPB C 0.00596185f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_60 VPB N_C_c_216_n 0.0208819f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_61 VPB N_B_c_270_n 0.0103731f $X=-0.19 $Y=1.66 $X2=0.63 $Y2=0.69
cc_62 VPB N_B_c_271_n 0.00491078f $X=-0.19 $Y=1.66 $X2=0.63 $Y2=0.69
cc_63 VPB N_B_c_279_n 0.0186627f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_64 VPB N_B_c_273_n 0.00805595f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_65 VPB N_B_c_281_n 0.0155755f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_66 VPB N_B_c_274_n 0.00607543f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_67 VPB B 0.0140418f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_68 VPB N_B_c_276_n 0.00638865f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_69 VPB N_A_c_336_n 0.0153838f $X=-0.19 $Y=1.66 $X2=0.63 $Y2=0.69
cc_70 VPB N_A_c_337_n 0.0201619f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_71 VPB A 0.0149285f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_72 VPB N_A_c_335_n 0.0218327f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_73 VPB N_VPWR_c_378_n 0.0156399f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_74 VPB N_VPWR_c_379_n 0.00396467f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_75 VPB N_VPWR_c_380_n 0.0180274f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_76 VPB N_VPWR_c_381_n 0.0953726f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_77 VPB N_VPWR_c_382_n 0.018982f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_78 VPB N_VPWR_c_377_n 0.0917025f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_79 VPB N_VPWR_c_384_n 0.00614127f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_80 VPB N_VPWR_c_385_n 0.00601644f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_81 VPB N_A_229_368#_c_433_n 0.0130098f $X=-0.19 $Y=1.66 $X2=0.7 $Y2=1.635
cc_82 VPB N_A_229_368#_c_434_n 0.00479141f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_83 VPB N_A_229_368#_c_435_n 0.00431456f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_84 VPB N_A_229_368#_c_436_n 0.00226721f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_85 VPB N_A_229_368#_c_437_n 0.00257983f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_86 VPB N_Y_c_490_n 0.00314876f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_87 VPB N_Y_c_483_n 0.00305381f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_88 VPB N_A_498_368#_c_587_n 0.0192731f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_89 VPB N_A_498_368#_c_588_n 0.00216812f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_90 VPB N_A_701_368#_c_618_n 0.00198096f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.635
cc_91 VPB N_A_701_368#_c_619_n 0.00655998f $X=-0.19 $Y=1.66 $X2=0.7 $Y2=1.635
cc_92 VPB N_A_701_368#_c_620_n 0.00180901f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_93 VPB N_A_701_368#_c_621_n 0.00723723f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_94 VPB N_A_701_368#_c_622_n 0.0339676f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_95 N_D_N_M1002_g N_A_27_392#_c_127_n 0.0211411f $X=0.63 $Y=0.69 $X2=0 $Y2=0
cc_96 N_D_N_c_95_n N_A_27_392#_c_135_n 8.14646e-19 $X=0.505 $Y=1.885 $X2=0 $Y2=0
cc_97 N_D_N_M1002_g N_A_27_392#_c_129_n 0.0131116f $X=0.63 $Y=0.69 $X2=0 $Y2=0
cc_98 N_D_N_c_95_n N_A_27_392#_c_130_n 0.0197909f $X=0.505 $Y=1.885 $X2=0 $Y2=0
cc_99 N_D_N_M1002_g N_A_27_392#_c_130_n 0.00592896f $X=0.63 $Y=0.69 $X2=0 $Y2=0
cc_100 D_N N_A_27_392#_c_130_n 0.025547f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_101 N_D_N_c_95_n N_A_27_392#_c_131_n 0.00596036f $X=0.505 $Y=1.885 $X2=0
+ $Y2=0
cc_102 N_D_N_M1002_g N_A_27_392#_c_131_n 0.00449144f $X=0.63 $Y=0.69 $X2=0 $Y2=0
cc_103 D_N N_A_27_392#_c_131_n 0.00361618f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_104 N_D_N_c_95_n N_A_27_392#_c_132_n 3.08012e-19 $X=0.505 $Y=1.885 $X2=0
+ $Y2=0
cc_105 N_D_N_M1002_g N_A_27_392#_c_132_n 9.66795e-19 $X=0.63 $Y=0.69 $X2=0 $Y2=0
cc_106 D_N N_A_27_392#_c_132_n 0.00477495f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_107 N_D_N_c_95_n N_A_27_392#_c_133_n 0.00112087f $X=0.505 $Y=1.885 $X2=0
+ $Y2=0
cc_108 N_D_N_M1002_g N_A_27_392#_c_133_n 0.0117536f $X=0.63 $Y=0.69 $X2=0 $Y2=0
cc_109 D_N N_A_27_392#_c_133_n 0.0209481f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_110 N_D_N_c_95_n N_A_27_392#_c_134_n 0.0096455f $X=0.505 $Y=1.885 $X2=0 $Y2=0
cc_111 N_D_N_M1002_g N_A_27_392#_c_134_n 0.00670227f $X=0.63 $Y=0.69 $X2=0 $Y2=0
cc_112 D_N N_A_27_392#_c_134_n 0.00123122f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_113 N_D_N_c_95_n N_VPWR_c_378_n 0.0205212f $X=0.505 $Y=1.885 $X2=0 $Y2=0
cc_114 D_N N_VPWR_c_378_n 0.0220821f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_115 N_D_N_c_95_n N_VPWR_c_380_n 0.00413917f $X=0.505 $Y=1.885 $X2=0 $Y2=0
cc_116 N_D_N_c_95_n N_VPWR_c_377_n 0.00821221f $X=0.505 $Y=1.885 $X2=0 $Y2=0
cc_117 N_D_N_c_95_n N_A_229_368#_c_433_n 0.00369308f $X=0.505 $Y=1.885 $X2=0
+ $Y2=0
cc_118 N_D_N_c_95_n N_A_229_368#_c_435_n 5.94256e-19 $X=0.505 $Y=1.885 $X2=0
+ $Y2=0
cc_119 N_D_N_M1002_g N_VGND_c_660_n 0.00695483f $X=0.63 $Y=0.69 $X2=0 $Y2=0
cc_120 N_D_N_M1002_g N_VGND_c_664_n 0.00434272f $X=0.63 $Y=0.69 $X2=0 $Y2=0
cc_121 N_D_N_M1002_g N_VGND_c_672_n 0.0082535f $X=0.63 $Y=0.69 $X2=0 $Y2=0
cc_122 N_A_27_392#_c_128_n N_C_M1012_g 0.0180513f $X=1.7 $Y=1.22 $X2=0 $Y2=0
cc_123 N_A_27_392#_c_132_n N_C_M1012_g 8.7155e-19 $X=1.61 $Y=1.385 $X2=0 $Y2=0
cc_124 N_A_27_392#_c_134_n N_C_M1012_g 0.0240309f $X=1.7 $Y=1.492 $X2=0 $Y2=0
cc_125 N_A_27_392#_c_136_n N_C_c_217_n 0.0260422f $X=1.965 $Y=1.765 $X2=0 $Y2=0
cc_126 N_A_27_392#_c_136_n C 4.69145e-19 $X=1.965 $Y=1.765 $X2=0 $Y2=0
cc_127 N_A_27_392#_c_132_n C 0.0115655f $X=1.61 $Y=1.385 $X2=0 $Y2=0
cc_128 N_A_27_392#_c_134_n C 0.0139165f $X=1.7 $Y=1.492 $X2=0 $Y2=0
cc_129 N_A_27_392#_c_134_n N_C_c_216_n 0.00401348f $X=1.7 $Y=1.492 $X2=0 $Y2=0
cc_130 N_A_27_392#_c_135_n N_VPWR_c_378_n 0.00256389f $X=1.515 $Y=1.765 $X2=0
+ $Y2=0
cc_131 N_A_27_392#_c_130_n N_VPWR_c_378_n 0.0677511f $X=0.28 $Y=2.105 $X2=0
+ $Y2=0
cc_132 N_A_27_392#_c_133_n N_VPWR_c_378_n 9.48018e-19 $X=1.105 $Y=1.34 $X2=0
+ $Y2=0
cc_133 N_A_27_392#_c_130_n N_VPWR_c_380_n 0.011066f $X=0.28 $Y=2.105 $X2=0 $Y2=0
cc_134 N_A_27_392#_c_135_n N_VPWR_c_381_n 0.00278257f $X=1.515 $Y=1.765 $X2=0
+ $Y2=0
cc_135 N_A_27_392#_c_136_n N_VPWR_c_381_n 0.00278257f $X=1.965 $Y=1.765 $X2=0
+ $Y2=0
cc_136 N_A_27_392#_c_135_n N_VPWR_c_377_n 0.00358623f $X=1.515 $Y=1.765 $X2=0
+ $Y2=0
cc_137 N_A_27_392#_c_136_n N_VPWR_c_377_n 0.00353905f $X=1.965 $Y=1.765 $X2=0
+ $Y2=0
cc_138 N_A_27_392#_c_130_n N_VPWR_c_377_n 0.00915947f $X=0.28 $Y=2.105 $X2=0
+ $Y2=0
cc_139 N_A_27_392#_c_135_n N_A_229_368#_c_433_n 0.0139009f $X=1.515 $Y=1.765
+ $X2=0 $Y2=0
cc_140 N_A_27_392#_c_136_n N_A_229_368#_c_433_n 6.23098e-19 $X=1.965 $Y=1.765
+ $X2=0 $Y2=0
cc_141 N_A_27_392#_c_132_n N_A_229_368#_c_433_n 0.0198519f $X=1.61 $Y=1.385
+ $X2=0 $Y2=0
cc_142 N_A_27_392#_c_134_n N_A_229_368#_c_433_n 0.0079078f $X=1.7 $Y=1.492 $X2=0
+ $Y2=0
cc_143 N_A_27_392#_c_135_n N_A_229_368#_c_434_n 0.0107904f $X=1.515 $Y=1.765
+ $X2=0 $Y2=0
cc_144 N_A_27_392#_c_136_n N_A_229_368#_c_434_n 0.0122595f $X=1.965 $Y=1.765
+ $X2=0 $Y2=0
cc_145 N_A_27_392#_c_135_n N_A_229_368#_c_435_n 0.00262934f $X=1.515 $Y=1.765
+ $X2=0 $Y2=0
cc_146 N_A_27_392#_c_136_n N_A_229_368#_c_447_n 0.00193585f $X=1.965 $Y=1.765
+ $X2=0 $Y2=0
cc_147 N_A_27_392#_c_135_n N_A_229_368#_c_448_n 5.20641e-19 $X=1.515 $Y=1.765
+ $X2=0 $Y2=0
cc_148 N_A_27_392#_c_136_n N_A_229_368#_c_448_n 0.00574124f $X=1.965 $Y=1.765
+ $X2=0 $Y2=0
cc_149 N_A_27_392#_c_127_n N_Y_c_481_n 0.0054187f $X=1.2 $Y=1.22 $X2=0 $Y2=0
cc_150 N_A_27_392#_c_128_n N_Y_c_481_n 0.00252693f $X=1.7 $Y=1.22 $X2=0 $Y2=0
cc_151 N_A_27_392#_c_128_n N_Y_c_494_n 0.0130155f $X=1.7 $Y=1.22 $X2=0 $Y2=0
cc_152 N_A_27_392#_c_132_n N_Y_c_494_n 0.0128666f $X=1.61 $Y=1.385 $X2=0 $Y2=0
cc_153 N_A_27_392#_c_134_n N_Y_c_494_n 0.00946034f $X=1.7 $Y=1.492 $X2=0 $Y2=0
cc_154 N_A_27_392#_c_127_n N_Y_c_497_n 0.00209321f $X=1.2 $Y=1.22 $X2=0 $Y2=0
cc_155 N_A_27_392#_c_132_n N_Y_c_497_n 0.0256756f $X=1.61 $Y=1.385 $X2=0 $Y2=0
cc_156 N_A_27_392#_c_134_n N_Y_c_497_n 0.00105137f $X=1.7 $Y=1.492 $X2=0 $Y2=0
cc_157 N_A_27_392#_c_135_n N_Y_c_490_n 0.00124352f $X=1.515 $Y=1.765 $X2=0 $Y2=0
cc_158 N_A_27_392#_c_136_n N_Y_c_490_n 0.00262483f $X=1.965 $Y=1.765 $X2=0 $Y2=0
cc_159 N_A_27_392#_c_132_n N_Y_c_490_n 0.00728815f $X=1.61 $Y=1.385 $X2=0 $Y2=0
cc_160 N_A_27_392#_c_134_n N_Y_c_490_n 0.00244512f $X=1.7 $Y=1.492 $X2=0 $Y2=0
cc_161 N_A_27_392#_c_135_n N_Y_c_504_n 0.00279093f $X=1.515 $Y=1.765 $X2=0 $Y2=0
cc_162 N_A_27_392#_c_136_n N_Y_c_504_n 0.00554106f $X=1.965 $Y=1.765 $X2=0 $Y2=0
cc_163 N_A_27_392#_c_136_n N_Y_c_506_n 0.0171543f $X=1.965 $Y=1.765 $X2=0 $Y2=0
cc_164 N_A_27_392#_c_128_n N_Y_c_482_n 9.57264e-19 $X=1.7 $Y=1.22 $X2=0 $Y2=0
cc_165 N_A_27_392#_c_128_n N_Y_c_485_n 7.73117e-19 $X=1.7 $Y=1.22 $X2=0 $Y2=0
cc_166 N_A_27_392#_c_132_n N_Y_c_485_n 0.00131831f $X=1.61 $Y=1.385 $X2=0 $Y2=0
cc_167 N_A_27_392#_c_127_n N_VGND_c_660_n 0.0054296f $X=1.2 $Y=1.22 $X2=0 $Y2=0
cc_168 N_A_27_392#_c_129_n N_VGND_c_660_n 0.0249119f $X=0.415 $Y=0.515 $X2=0
+ $Y2=0
cc_169 N_A_27_392#_c_133_n N_VGND_c_660_n 0.0261348f $X=1.105 $Y=1.34 $X2=0
+ $Y2=0
cc_170 N_A_27_392#_c_129_n N_VGND_c_664_n 0.0205877f $X=0.415 $Y=0.515 $X2=0
+ $Y2=0
cc_171 N_A_27_392#_c_127_n N_VGND_c_666_n 0.00433834f $X=1.2 $Y=1.22 $X2=0 $Y2=0
cc_172 N_A_27_392#_c_128_n N_VGND_c_666_n 0.00384553f $X=1.7 $Y=1.22 $X2=0 $Y2=0
cc_173 N_A_27_392#_c_127_n N_VGND_c_670_n 3.64777e-19 $X=1.2 $Y=1.22 $X2=0 $Y2=0
cc_174 N_A_27_392#_c_128_n N_VGND_c_670_n 0.0117177f $X=1.7 $Y=1.22 $X2=0 $Y2=0
cc_175 N_A_27_392#_c_127_n N_VGND_c_672_n 0.00821665f $X=1.2 $Y=1.22 $X2=0 $Y2=0
cc_176 N_A_27_392#_c_128_n N_VGND_c_672_n 0.00374134f $X=1.7 $Y=1.22 $X2=0 $Y2=0
cc_177 N_A_27_392#_c_129_n N_VGND_c_672_n 0.0169844f $X=0.415 $Y=0.515 $X2=0
+ $Y2=0
cc_178 N_C_M1016_g N_B_M1007_g 0.0210645f $X=2.82 $Y=0.74 $X2=0 $Y2=0
cc_179 N_C_c_216_n N_B_c_271_n 0.0116958f $X=2.82 $Y=1.557 $X2=0 $Y2=0
cc_180 N_C_c_216_n B 8.19567e-19 $X=2.82 $Y=1.557 $X2=0 $Y2=0
cc_181 N_C_c_217_n N_VPWR_c_381_n 0.00444353f $X=2.415 $Y=1.765 $X2=0 $Y2=0
cc_182 N_C_c_218_n N_VPWR_c_381_n 0.00279479f $X=2.865 $Y=1.765 $X2=0 $Y2=0
cc_183 N_C_c_217_n N_VPWR_c_377_n 0.00857912f $X=2.415 $Y=1.765 $X2=0 $Y2=0
cc_184 N_C_c_218_n N_VPWR_c_377_n 0.00357714f $X=2.865 $Y=1.765 $X2=0 $Y2=0
cc_185 N_C_c_217_n N_A_229_368#_c_434_n 0.00125031f $X=2.415 $Y=1.765 $X2=0
+ $Y2=0
cc_186 N_C_c_217_n N_A_229_368#_c_436_n 0.0124723f $X=2.415 $Y=1.765 $X2=0 $Y2=0
cc_187 N_C_c_218_n N_A_229_368#_c_436_n 0.010317f $X=2.865 $Y=1.765 $X2=0 $Y2=0
cc_188 N_C_c_218_n N_A_229_368#_c_437_n 0.00452127f $X=2.865 $Y=1.765 $X2=0
+ $Y2=0
cc_189 N_C_M1012_g N_Y_c_494_n 0.0104376f $X=2.39 $Y=0.74 $X2=0 $Y2=0
cc_190 C N_Y_c_494_n 0.0154053f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_191 N_C_c_217_n N_Y_c_506_n 0.0106304f $X=2.415 $Y=1.765 $X2=0 $Y2=0
cc_192 N_C_c_218_n N_Y_c_506_n 0.015369f $X=2.865 $Y=1.765 $X2=0 $Y2=0
cc_193 C N_Y_c_506_n 0.0487216f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_194 N_C_c_216_n N_Y_c_506_n 0.00123707f $X=2.82 $Y=1.557 $X2=0 $Y2=0
cc_195 N_C_M1012_g N_Y_c_482_n 0.00798642f $X=2.39 $Y=0.74 $X2=0 $Y2=0
cc_196 N_C_M1016_g N_Y_c_482_n 0.00570416f $X=2.82 $Y=0.74 $X2=0 $Y2=0
cc_197 N_C_c_217_n N_Y_c_483_n 8.25832e-19 $X=2.415 $Y=1.765 $X2=0 $Y2=0
cc_198 N_C_M1016_g N_Y_c_483_n 0.00443118f $X=2.82 $Y=0.74 $X2=0 $Y2=0
cc_199 N_C_c_218_n N_Y_c_483_n 0.00615153f $X=2.865 $Y=1.765 $X2=0 $Y2=0
cc_200 C N_Y_c_483_n 0.0331353f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_201 N_C_c_216_n N_Y_c_483_n 0.0115413f $X=2.82 $Y=1.557 $X2=0 $Y2=0
cc_202 N_C_M1012_g N_Y_c_485_n 0.00661837f $X=2.39 $Y=0.74 $X2=0 $Y2=0
cc_203 N_C_M1016_g N_Y_c_485_n 0.0216954f $X=2.82 $Y=0.74 $X2=0 $Y2=0
cc_204 C N_Y_c_485_n 0.0269015f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_205 N_C_c_216_n N_Y_c_485_n 0.00357751f $X=2.82 $Y=1.557 $X2=0 $Y2=0
cc_206 N_C_M1016_g Y 6.11074e-19 $X=2.82 $Y=0.74 $X2=0 $Y2=0
cc_207 N_C_c_218_n N_A_498_368#_c_587_n 0.0109692f $X=2.865 $Y=1.765 $X2=0 $Y2=0
cc_208 N_C_c_217_n N_A_498_368#_c_588_n 0.00620718f $X=2.415 $Y=1.765 $X2=0
+ $Y2=0
cc_209 N_C_c_218_n N_A_498_368#_c_588_n 0.0108447f $X=2.865 $Y=1.765 $X2=0 $Y2=0
cc_210 N_C_c_218_n N_A_701_368#_c_618_n 9.2581e-19 $X=2.865 $Y=1.765 $X2=0 $Y2=0
cc_211 N_C_c_218_n N_A_701_368#_c_619_n 0.00443991f $X=2.865 $Y=1.765 $X2=0
+ $Y2=0
cc_212 N_C_M1016_g N_VGND_c_661_n 0.00470005f $X=2.82 $Y=0.74 $X2=0 $Y2=0
cc_213 N_C_M1012_g N_VGND_c_667_n 0.00434272f $X=2.39 $Y=0.74 $X2=0 $Y2=0
cc_214 N_C_M1016_g N_VGND_c_667_n 0.00434272f $X=2.82 $Y=0.74 $X2=0 $Y2=0
cc_215 N_C_M1012_g N_VGND_c_670_n 0.00400351f $X=2.39 $Y=0.74 $X2=0 $Y2=0
cc_216 N_C_M1012_g N_VGND_c_672_n 0.00436462f $X=2.39 $Y=0.74 $X2=0 $Y2=0
cc_217 N_C_M1016_g N_VGND_c_672_n 0.00821165f $X=2.82 $Y=0.74 $X2=0 $Y2=0
cc_218 N_B_c_281_n N_A_c_336_n 0.00823489f $X=4.325 $Y=1.765 $X2=0 $Y2=0
cc_219 N_B_c_274_n A 0.00256372f $X=4.325 $Y=1.605 $X2=0 $Y2=0
cc_220 B A 0.0298391f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_221 N_B_c_276_n A 5.80008e-19 $X=3.8 $Y=1.515 $X2=0 $Y2=0
cc_222 N_B_c_274_n N_A_c_335_n 0.0118804f $X=4.325 $Y=1.605 $X2=0 $Y2=0
cc_223 B N_A_c_335_n 7.03106e-19 $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_224 N_B_c_276_n N_A_c_335_n 0.0018393f $X=3.8 $Y=1.515 $X2=0 $Y2=0
cc_225 N_B_c_281_n N_VPWR_c_379_n 5.74542e-19 $X=4.325 $Y=1.765 $X2=0 $Y2=0
cc_226 N_B_c_279_n N_VPWR_c_381_n 0.00278257f $X=3.875 $Y=1.765 $X2=0 $Y2=0
cc_227 N_B_c_281_n N_VPWR_c_381_n 0.0044313f $X=4.325 $Y=1.765 $X2=0 $Y2=0
cc_228 N_B_c_279_n N_VPWR_c_377_n 0.00358623f $X=3.875 $Y=1.765 $X2=0 $Y2=0
cc_229 N_B_c_281_n N_VPWR_c_377_n 0.00854206f $X=4.325 $Y=1.765 $X2=0 $Y2=0
cc_230 N_B_M1007_g N_Y_c_483_n 0.00358729f $X=3.37 $Y=0.74 $X2=0 $Y2=0
cc_231 N_B_c_271_n N_Y_c_483_n 0.00111277f $X=3.445 $Y=1.515 $X2=0 $Y2=0
cc_232 B N_Y_c_483_n 0.0306983f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_233 N_B_c_276_n N_Y_c_483_n 2.30571e-19 $X=3.8 $Y=1.515 $X2=0 $Y2=0
cc_234 N_B_M1007_g N_Y_c_484_n 0.0131887f $X=3.37 $Y=0.74 $X2=0 $Y2=0
cc_235 B N_Y_c_484_n 0.0105458f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_236 N_B_M1007_g N_Y_c_485_n 4.69564e-19 $X=3.37 $Y=0.74 $X2=0 $Y2=0
cc_237 N_B_M1013_g N_Y_c_486_n 0.0169209f $X=3.89 $Y=0.74 $X2=0 $Y2=0
cc_238 N_B_c_273_n N_Y_c_486_n 0.00821843f $X=4.235 $Y=1.605 $X2=0 $Y2=0
cc_239 B N_Y_c_486_n 0.0329461f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_240 N_B_M1007_g Y 0.00856724f $X=3.37 $Y=0.74 $X2=0 $Y2=0
cc_241 N_B_M1013_g Y 0.00366931f $X=3.89 $Y=0.74 $X2=0 $Y2=0
cc_242 N_B_M1007_g N_Y_c_489_n 0.00116959f $X=3.37 $Y=0.74 $X2=0 $Y2=0
cc_243 N_B_c_270_n N_Y_c_489_n 0.00442617f $X=3.785 $Y=1.515 $X2=0 $Y2=0
cc_244 B N_Y_c_489_n 0.028285f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_245 N_B_c_279_n N_A_498_368#_c_587_n 0.0145139f $X=3.875 $Y=1.765 $X2=0 $Y2=0
cc_246 N_B_c_281_n N_A_498_368#_c_587_n 0.00396164f $X=4.325 $Y=1.765 $X2=0
+ $Y2=0
cc_247 N_B_c_279_n N_A_498_368#_c_594_n 0.0121561f $X=3.875 $Y=1.765 $X2=0 $Y2=0
cc_248 N_B_c_281_n N_A_498_368#_c_594_n 0.00641928f $X=4.325 $Y=1.765 $X2=0
+ $Y2=0
cc_249 N_B_c_270_n N_A_701_368#_c_618_n 0.0015368f $X=3.785 $Y=1.515 $X2=0 $Y2=0
cc_250 B N_A_701_368#_c_618_n 0.0221345f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_251 N_B_c_279_n N_A_701_368#_c_619_n 0.00787215f $X=3.875 $Y=1.765 $X2=0
+ $Y2=0
cc_252 N_B_c_279_n N_A_701_368#_c_628_n 0.0126853f $X=3.875 $Y=1.765 $X2=0 $Y2=0
cc_253 N_B_c_273_n N_A_701_368#_c_628_n 0.00118771f $X=4.235 $Y=1.605 $X2=0
+ $Y2=0
cc_254 N_B_c_281_n N_A_701_368#_c_628_n 0.0167755f $X=4.325 $Y=1.765 $X2=0 $Y2=0
cc_255 B N_A_701_368#_c_628_n 0.0313533f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_256 N_B_c_281_n N_A_701_368#_c_620_n 0.00554871f $X=4.325 $Y=1.765 $X2=0
+ $Y2=0
cc_257 N_B_M1007_g N_VGND_c_661_n 0.0027066f $X=3.37 $Y=0.74 $X2=0 $Y2=0
cc_258 N_B_M1007_g N_VGND_c_668_n 0.00504858f $X=3.37 $Y=0.74 $X2=0 $Y2=0
cc_259 N_B_M1013_g N_VGND_c_668_n 0.0159343f $X=3.89 $Y=0.74 $X2=0 $Y2=0
cc_260 N_B_M1007_g N_VGND_c_672_n 0.00891136f $X=3.37 $Y=0.74 $X2=0 $Y2=0
cc_261 N_B_M1013_g N_VGND_c_672_n 0.00758371f $X=3.89 $Y=0.74 $X2=0 $Y2=0
cc_262 N_A_c_336_n N_VPWR_c_379_n 0.0111113f $X=4.775 $Y=1.765 $X2=0 $Y2=0
cc_263 N_A_c_337_n N_VPWR_c_379_n 0.0132819f $X=5.235 $Y=1.765 $X2=0 $Y2=0
cc_264 N_A_c_336_n N_VPWR_c_381_n 0.00413917f $X=4.775 $Y=1.765 $X2=0 $Y2=0
cc_265 N_A_c_337_n N_VPWR_c_382_n 0.00444681f $X=5.235 $Y=1.765 $X2=0 $Y2=0
cc_266 N_A_c_336_n N_VPWR_c_377_n 0.0081781f $X=4.775 $Y=1.765 $X2=0 $Y2=0
cc_267 N_A_c_337_n N_VPWR_c_377_n 0.00881275f $X=5.235 $Y=1.765 $X2=0 $Y2=0
cc_268 N_A_M1009_g N_Y_c_486_n 0.0147517f $X=4.765 $Y=0.74 $X2=0 $Y2=0
cc_269 N_A_M1014_g N_Y_c_486_n 0.00185032f $X=5.25 $Y=0.74 $X2=0 $Y2=0
cc_270 A N_Y_c_486_n 0.0570125f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_271 N_A_c_335_n N_Y_c_486_n 0.00440097f $X=5.235 $Y=1.557 $X2=0 $Y2=0
cc_272 N_A_M1009_g N_Y_c_487_n 0.0153465f $X=4.765 $Y=0.74 $X2=0 $Y2=0
cc_273 N_A_M1014_g N_Y_c_487_n 4.79228e-19 $X=5.25 $Y=0.74 $X2=0 $Y2=0
cc_274 N_A_c_336_n N_A_498_368#_c_587_n 3.01915e-19 $X=4.775 $Y=1.765 $X2=0
+ $Y2=0
cc_275 A N_A_701_368#_c_628_n 0.00112091f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_276 N_A_c_336_n N_A_701_368#_c_620_n 0.00554978f $X=4.775 $Y=1.765 $X2=0
+ $Y2=0
cc_277 N_A_c_336_n N_A_701_368#_c_635_n 0.0127429f $X=4.775 $Y=1.765 $X2=0 $Y2=0
cc_278 N_A_c_337_n N_A_701_368#_c_635_n 0.0129941f $X=5.235 $Y=1.765 $X2=0 $Y2=0
cc_279 A N_A_701_368#_c_635_n 0.0485148f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_280 N_A_c_335_n N_A_701_368#_c_635_n 0.0013663f $X=5.235 $Y=1.557 $X2=0 $Y2=0
cc_281 A N_A_701_368#_c_621_n 0.0221348f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_282 N_A_c_337_n N_A_701_368#_c_622_n 0.00645576f $X=5.235 $Y=1.765 $X2=0
+ $Y2=0
cc_283 A N_A_701_368#_c_641_n 0.0150276f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_284 N_A_M1009_g N_VGND_c_663_n 5.65034e-19 $X=4.765 $Y=0.74 $X2=0 $Y2=0
cc_285 N_A_M1014_g N_VGND_c_663_n 0.0137863f $X=5.25 $Y=0.74 $X2=0 $Y2=0
cc_286 A N_VGND_c_663_n 0.023911f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_287 N_A_M1009_g N_VGND_c_668_n 0.00509578f $X=4.765 $Y=0.74 $X2=0 $Y2=0
cc_288 N_A_M1009_g N_VGND_c_669_n 0.00434272f $X=4.765 $Y=0.74 $X2=0 $Y2=0
cc_289 N_A_M1014_g N_VGND_c_669_n 0.00429299f $X=5.25 $Y=0.74 $X2=0 $Y2=0
cc_290 N_A_M1009_g N_VGND_c_672_n 0.00825583f $X=4.765 $Y=0.74 $X2=0 $Y2=0
cc_291 N_A_M1014_g N_VGND_c_672_n 0.00848048f $X=5.25 $Y=0.74 $X2=0 $Y2=0
cc_292 N_VPWR_c_378_n N_A_229_368#_c_433_n 0.0630028f $X=0.73 $Y=2.135 $X2=0
+ $Y2=0
cc_293 N_VPWR_c_381_n N_A_229_368#_c_434_n 0.053749f $X=4.835 $Y=3.33 $X2=0
+ $Y2=0
cc_294 N_VPWR_c_377_n N_A_229_368#_c_434_n 0.029846f $X=5.52 $Y=3.33 $X2=0 $Y2=0
cc_295 N_VPWR_c_378_n N_A_229_368#_c_435_n 0.0121617f $X=0.73 $Y=2.135 $X2=0
+ $Y2=0
cc_296 N_VPWR_c_381_n N_A_229_368#_c_435_n 0.0236039f $X=4.835 $Y=3.33 $X2=0
+ $Y2=0
cc_297 N_VPWR_c_377_n N_A_229_368#_c_435_n 0.012761f $X=5.52 $Y=3.33 $X2=0 $Y2=0
cc_298 N_VPWR_c_379_n N_A_498_368#_c_587_n 0.00279034f $X=5 $Y=2.455 $X2=0 $Y2=0
cc_299 N_VPWR_c_381_n N_A_498_368#_c_587_n 0.0955317f $X=4.835 $Y=3.33 $X2=0
+ $Y2=0
cc_300 N_VPWR_c_377_n N_A_498_368#_c_587_n 0.0539458f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_301 N_VPWR_c_381_n N_A_498_368#_c_588_n 0.0226868f $X=4.835 $Y=3.33 $X2=0
+ $Y2=0
cc_302 N_VPWR_c_377_n N_A_498_368#_c_588_n 0.0124868f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_303 N_VPWR_c_379_n N_A_701_368#_c_620_n 0.0449718f $X=5 $Y=2.455 $X2=0 $Y2=0
cc_304 N_VPWR_c_381_n N_A_701_368#_c_620_n 0.00749631f $X=4.835 $Y=3.33 $X2=0
+ $Y2=0
cc_305 N_VPWR_c_377_n N_A_701_368#_c_620_n 0.0062048f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_306 N_VPWR_M1005_d N_A_701_368#_c_635_n 0.00378686f $X=4.85 $Y=1.84 $X2=0
+ $Y2=0
cc_307 N_VPWR_c_379_n N_A_701_368#_c_635_n 0.0172332f $X=5 $Y=2.455 $X2=0 $Y2=0
cc_308 N_VPWR_c_379_n N_A_701_368#_c_622_n 0.0445954f $X=5 $Y=2.455 $X2=0 $Y2=0
cc_309 N_VPWR_c_382_n N_A_701_368#_c_622_n 0.011066f $X=5.52 $Y=3.33 $X2=0 $Y2=0
cc_310 N_VPWR_c_377_n N_A_701_368#_c_622_n 0.00915947f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_311 N_A_229_368#_c_434_n N_Y_M1001_s 0.00239636f $X=2.025 $Y=2.99 $X2=0 $Y2=0
cc_312 N_A_229_368#_c_433_n N_Y_c_490_n 0.020917f $X=1.29 $Y=1.985 $X2=0 $Y2=0
cc_313 N_A_229_368#_c_433_n N_Y_c_504_n 0.040027f $X=1.29 $Y=1.985 $X2=0 $Y2=0
cc_314 N_A_229_368#_c_434_n N_Y_c_504_n 0.012787f $X=2.025 $Y=2.99 $X2=0 $Y2=0
cc_315 N_A_229_368#_c_447_n N_Y_c_504_n 0.0117758f $X=2.15 $Y=2.46 $X2=0 $Y2=0
cc_316 N_A_229_368#_c_448_n N_Y_c_504_n 0.0175037f $X=2.15 $Y=2.905 $X2=0 $Y2=0
cc_317 N_A_229_368#_M1017_d N_Y_c_506_n 0.00395946f $X=2.04 $Y=1.84 $X2=0 $Y2=0
cc_318 N_A_229_368#_M1006_s N_Y_c_506_n 0.00388371f $X=2.94 $Y=1.84 $X2=0 $Y2=0
cc_319 N_A_229_368#_c_447_n N_Y_c_506_n 0.0155823f $X=2.15 $Y=2.46 $X2=0 $Y2=0
cc_320 N_A_229_368#_c_436_n N_Y_c_506_n 0.042844f $X=3.005 $Y=2.375 $X2=0 $Y2=0
cc_321 N_A_229_368#_M1006_s N_Y_c_483_n 0.00415896f $X=2.94 $Y=1.84 $X2=0 $Y2=0
cc_322 N_A_229_368#_c_436_n N_A_498_368#_M1004_d 0.00379409f $X=3.005 $Y=2.375
+ $X2=-0.19 $Y2=1.66
cc_323 N_A_229_368#_M1006_s N_A_498_368#_c_587_n 0.00291383f $X=2.94 $Y=1.84
+ $X2=0 $Y2=0
cc_324 N_A_229_368#_c_436_n N_A_498_368#_c_587_n 0.00445035f $X=3.005 $Y=2.375
+ $X2=0 $Y2=0
cc_325 N_A_229_368#_c_437_n N_A_498_368#_c_587_n 0.0183294f $X=3.13 $Y=2.46
+ $X2=0 $Y2=0
cc_326 N_A_229_368#_c_434_n N_A_498_368#_c_588_n 0.0125885f $X=2.025 $Y=2.99
+ $X2=0 $Y2=0
cc_327 N_A_229_368#_c_448_n N_A_498_368#_c_588_n 0.0184049f $X=2.15 $Y=2.905
+ $X2=0 $Y2=0
cc_328 N_A_229_368#_c_436_n N_A_498_368#_c_588_n 0.0166041f $X=3.005 $Y=2.375
+ $X2=0 $Y2=0
cc_329 N_A_229_368#_c_437_n N_A_498_368#_c_588_n 0.00704037f $X=3.13 $Y=2.46
+ $X2=0 $Y2=0
cc_330 N_A_229_368#_c_436_n N_A_701_368#_c_619_n 0.0119251f $X=3.005 $Y=2.375
+ $X2=0 $Y2=0
cc_331 N_A_229_368#_c_437_n N_A_701_368#_c_619_n 0.0177446f $X=3.13 $Y=2.46
+ $X2=0 $Y2=0
cc_332 N_Y_c_506_n N_A_498_368#_M1004_d 0.00359847f $X=2.925 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_333 N_Y_c_506_n N_A_701_368#_c_618_n 0.00860459f $X=2.925 $Y=2.035 $X2=0
+ $Y2=0
cc_334 N_Y_c_494_n N_VGND_M1011_d 0.0123139f $X=2.44 $Y=0.875 $X2=0 $Y2=0
cc_335 N_Y_c_484_n N_VGND_M1016_d 0.0016136f $X=3.44 $Y=1.095 $X2=0 $Y2=0
cc_336 N_Y_c_485_n N_VGND_M1016_d 0.00169317f $X=3.095 $Y=1.095 $X2=0 $Y2=0
cc_337 N_Y_c_486_n N_VGND_M1013_s 0.00926984f $X=4.815 $Y=1.095 $X2=0 $Y2=0
cc_338 N_Y_c_481_n N_VGND_c_660_n 0.0188454f $X=1.415 $Y=0.495 $X2=0 $Y2=0
cc_339 N_Y_c_482_n N_VGND_c_661_n 0.0172628f $X=2.605 $Y=0.515 $X2=0 $Y2=0
cc_340 N_Y_c_484_n N_VGND_c_661_n 0.0115978f $X=3.44 $Y=1.095 $X2=0 $Y2=0
cc_341 N_Y_c_485_n N_VGND_c_661_n 0.0128931f $X=3.095 $Y=1.095 $X2=0 $Y2=0
cc_342 Y N_VGND_c_661_n 0.0191764f $X=3.515 $Y=0.47 $X2=0 $Y2=0
cc_343 N_Y_c_486_n N_VGND_c_663_n 0.00540983f $X=4.815 $Y=1.095 $X2=0 $Y2=0
cc_344 N_Y_c_487_n N_VGND_c_663_n 0.0255552f $X=4.98 $Y=0.515 $X2=0 $Y2=0
cc_345 N_Y_c_481_n N_VGND_c_666_n 0.0157475f $X=1.415 $Y=0.495 $X2=0 $Y2=0
cc_346 N_Y_c_482_n N_VGND_c_667_n 0.0144922f $X=2.605 $Y=0.515 $X2=0 $Y2=0
cc_347 N_Y_c_486_n N_VGND_c_668_n 0.0424937f $X=4.815 $Y=1.095 $X2=0 $Y2=0
cc_348 N_Y_c_487_n N_VGND_c_668_n 0.0173963f $X=4.98 $Y=0.515 $X2=0 $Y2=0
cc_349 Y N_VGND_c_668_n 0.0339549f $X=3.515 $Y=0.47 $X2=0 $Y2=0
cc_350 N_Y_c_487_n N_VGND_c_669_n 0.0145639f $X=4.98 $Y=0.515 $X2=0 $Y2=0
cc_351 N_Y_c_481_n N_VGND_c_670_n 0.0124832f $X=1.415 $Y=0.495 $X2=0 $Y2=0
cc_352 N_Y_c_494_n N_VGND_c_670_n 0.0323939f $X=2.44 $Y=0.875 $X2=0 $Y2=0
cc_353 N_Y_c_482_n N_VGND_c_670_n 0.0102273f $X=2.605 $Y=0.515 $X2=0 $Y2=0
cc_354 N_Y_c_481_n N_VGND_c_672_n 0.0121127f $X=1.415 $Y=0.495 $X2=0 $Y2=0
cc_355 N_Y_c_494_n N_VGND_c_672_n 0.0123705f $X=2.44 $Y=0.875 $X2=0 $Y2=0
cc_356 N_Y_c_482_n N_VGND_c_672_n 0.0118826f $X=2.605 $Y=0.515 $X2=0 $Y2=0
cc_357 N_Y_c_487_n N_VGND_c_672_n 0.0119984f $X=4.98 $Y=0.515 $X2=0 $Y2=0
cc_358 Y N_VGND_c_672_n 0.0120948f $X=3.515 $Y=0.47 $X2=0 $Y2=0
cc_359 N_A_498_368#_c_587_n N_A_701_368#_M1000_s 0.00312144f $X=3.935 $Y=2.99
+ $X2=-0.19 $Y2=1.66
cc_360 N_A_498_368#_c_587_n N_A_701_368#_c_619_n 0.018931f $X=3.935 $Y=2.99
+ $X2=0 $Y2=0
cc_361 N_A_498_368#_c_594_n N_A_701_368#_c_619_n 0.0298377f $X=4.1 $Y=2.455
+ $X2=0 $Y2=0
cc_362 N_A_498_368#_M1000_d N_A_701_368#_c_628_n 0.00359365f $X=3.95 $Y=1.84
+ $X2=0 $Y2=0
cc_363 N_A_498_368#_c_594_n N_A_701_368#_c_628_n 0.0171813f $X=4.1 $Y=2.455
+ $X2=0 $Y2=0
cc_364 N_A_498_368#_c_587_n N_A_701_368#_c_620_n 0.00522251f $X=3.935 $Y=2.99
+ $X2=0 $Y2=0
cc_365 N_A_498_368#_c_594_n N_A_701_368#_c_620_n 0.0400262f $X=4.1 $Y=2.455
+ $X2=0 $Y2=0
