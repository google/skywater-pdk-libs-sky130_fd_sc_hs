* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hs__sdfsbp_1 CLK D SCD SCE SET_B VGND VNB VPB VPWR Q Q_N
X0 VPWR SET_B a_1762_74# VPB sky130_fd_pr__pfet_01v8 w=420000u l=150000u
X1 a_290_464# a_781_74# a_995_74# VPB sky130_fd_pr__pfet_01v8 w=420000u l=150000u
X2 a_206_464# D a_290_464# VPB sky130_fd_pr__pfet_01v8 w=640000u l=150000u
X3 a_2556_94# a_1762_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X4 a_1762_74# a_594_74# a_1600_347# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=150000u
X5 a_416_464# SCD VPWR VPB sky130_fd_pr__pfet_01v8 w=640000u l=150000u
X6 a_228_74# D a_290_464# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X7 a_1163_48# SET_B VPWR VPB sky130_fd_pr__pfet_01v8 w=420000u l=150000u
X8 VGND a_27_74# a_228_74# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X9 VPWR a_995_74# a_1600_347# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=150000u
X10 VPWR a_995_74# a_1163_48# VPB sky130_fd_pr__pfet_01v8 w=420000u l=150000u
X11 a_1954_74# SET_B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X12 VGND a_2556_94# Q VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X13 VPWR SCE a_206_464# VPB sky130_fd_pr__pfet_01v8 w=640000u l=150000u
X14 a_392_74# SCD VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X15 a_1411_74# SET_B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X16 a_1924_48# a_1762_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=420000u l=150000u
X17 a_290_464# SCE a_392_74# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X18 a_1712_374# a_1924_48# VPWR VPB sky130_fd_pr__pfet_01v8 w=420000u l=150000u
X19 a_290_464# a_27_74# a_416_464# VPB sky130_fd_pr__pfet_01v8 w=640000u l=150000u
X20 VPWR a_1762_74# Q_N VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X21 VPWR a_594_74# a_781_74# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X22 a_1684_74# a_781_74# a_1762_74# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X23 VGND a_1762_74# Q_N VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X24 a_995_74# a_594_74# a_1133_478# VPB sky130_fd_pr__pfet_01v8 w=420000u l=150000u
X25 VGND a_995_74# a_1684_74# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X26 VGND a_1762_74# a_1924_48# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X27 VGND a_594_74# a_781_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X28 a_290_464# a_594_74# a_995_74# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X29 a_2556_94# a_1762_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X30 a_1876_74# a_1924_48# a_1954_74# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X31 a_27_74# SCE VPWR VPB sky130_fd_pr__pfet_01v8 w=640000u l=150000u
X32 a_1163_48# a_995_74# a_1411_74# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X33 a_1762_74# a_594_74# a_1876_74# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X34 a_594_74# CLK VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X35 a_1712_374# a_781_74# a_1762_74# VPB sky130_fd_pr__pfet_01v8 w=420000u l=150000u
X36 a_1133_478# a_1163_48# VPWR VPB sky130_fd_pr__pfet_01v8 w=420000u l=150000u
X37 a_1115_74# a_1163_48# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X38 a_27_74# SCE VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X39 VPWR a_2556_94# Q VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X40 a_594_74# CLK VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X41 a_995_74# a_781_74# a_1115_74# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
.ends
