* File: sky130_fd_sc_hs__a31o_1.spice
* Created: Thu Aug 27 20:29:08 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hs__a31o_1.pex.spice"
.subckt sky130_fd_sc_hs__a31o_1  VNB VPB A3 A2 A1 B1 X VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* X	X
* B1	B1
* A1	A1
* A2	A2
* A3	A3
* VPB	VPB
* VNB	VNB
MM1007 N_VGND_M1007_d N_A_81_270#_M1007_g N_X_M1007_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.221517 AS=0.1961 PD=1.42638 PS=2.01 NRD=25.128 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75002.1 A=0.111 P=1.78 MULT=1
MM1008 A_265_120# N_A3_M1008_g N_VGND_M1007_d VNB NLOWVT L=0.15 W=0.64 AD=0.0672
+ AS=0.191583 PD=0.85 PS=1.23362 NRD=9.372 NRS=29.52 M=1 R=4.26667 SA=75000.9
+ SB=75001.7 A=0.096 P=1.58 MULT=1
MM1006 A_337_120# N_A2_M1006_g A_265_120# VNB NLOWVT L=0.15 W=0.64 AD=0.125625
+ AS=0.0672 PD=1.045 PS=0.85 NRD=26.484 NRS=9.372 M=1 R=4.26667 SA=75001.3
+ SB=75001.3 A=0.096 P=1.58 MULT=1
MM1009 N_A_81_270#_M1009_d N_A1_M1009_g A_337_120# VNB NLOWVT L=0.15 W=0.64
+ AD=0.1408 AS=0.125625 PD=1.08 PS=1.045 NRD=14.988 NRS=26.484 M=1 R=4.26667
+ SA=75001.8 SB=75000.8 A=0.096 P=1.58 MULT=1
MM1002 N_VGND_M1002_d N_B1_M1002_g N_A_81_270#_M1009_d VNB NLOWVT L=0.15 W=0.64
+ AD=0.1696 AS=0.1408 PD=1.81 PS=1.08 NRD=0 NRS=14.988 M=1 R=4.26667 SA=75002.4
+ SB=75000.2 A=0.096 P=1.58 MULT=1
MM1000 N_VPWR_M1000_d N_A_81_270#_M1000_g N_X_M1000_s VPB PSHORT L=0.15 W=1.12
+ AD=0.2968 AS=0.308 PD=1.7434 PS=2.79 NRD=21.9852 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75002.2 A=0.168 P=2.54 MULT=1
MM1001 N_A_250_392#_M1001_d N_A3_M1001_g N_VPWR_M1000_d VPB PSHORT L=0.15 W=1
+ AD=0.15 AS=0.265 PD=1.3 PS=1.5566 NRD=1.9503 NRS=24.6053 M=1 R=6.66667
+ SA=75000.9 SB=75001.7 A=0.15 P=2.3 MULT=1
MM1003 N_VPWR_M1003_d N_A2_M1003_g N_A_250_392#_M1001_d VPB PSHORT L=0.15 W=1
+ AD=0.24 AS=0.15 PD=1.48 PS=1.3 NRD=19.7 NRS=1.9503 M=1 R=6.66667 SA=75001.3
+ SB=75001.3 A=0.15 P=2.3 MULT=1
MM1004 N_A_250_392#_M1004_d N_A1_M1004_g N_VPWR_M1003_d VPB PSHORT L=0.15 W=1
+ AD=0.15 AS=0.24 PD=1.3 PS=1.48 NRD=1.9503 NRS=19.7 M=1 R=6.66667 SA=75002
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1005 N_A_81_270#_M1005_d N_B1_M1005_g N_A_250_392#_M1004_d VPB PSHORT L=0.15
+ W=1 AD=0.275 AS=0.15 PD=2.55 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=6.66667
+ SA=75002.4 SB=75000.2 A=0.15 P=2.3 MULT=1
DX10_noxref VNB VPB NWDIODE A=6.9564 P=11.2
*
.include "sky130_fd_sc_hs__a31o_1.pxi.spice"
*
.ends
*
*
