* File: sky130_fd_sc_hs__nand4_2.pex.spice
* Created: Thu Aug 27 20:51:51 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HS__NAND4_2%D 3 5 7 8 10 13 15 16 23 24
c42 23 0 9.82006e-20 $X=0.925 $Y=1.515
c43 13 0 8.01953e-20 $X=1.015 $Y=0.74
c44 8 0 1.84233e-19 $X=1 $Y=1.765
c45 5 0 1.64513e-19 $X=0.51 $Y=1.765
r46 24 25 1.928 $w=3.75e-07 $l=1.5e-08 $layer=POLY_cond $X=1 $Y=1.557 $X2=1.015
+ $Y2=1.557
r47 22 24 9.64 $w=3.75e-07 $l=7.5e-08 $layer=POLY_cond $X=0.925 $Y=1.557 $X2=1
+ $Y2=1.557
r48 22 23 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.925
+ $Y=1.515 $X2=0.925 $Y2=1.515
r49 20 22 53.3413 $w=3.75e-07 $l=4.15e-07 $layer=POLY_cond $X=0.51 $Y=1.557
+ $X2=0.925 $Y2=1.557
r50 19 20 1.928 $w=3.75e-07 $l=1.5e-08 $layer=POLY_cond $X=0.495 $Y=1.557
+ $X2=0.51 $Y2=1.557
r51 16 23 5.4942 $w=4.28e-07 $l=2.05e-07 $layer=LI1_cond $X=0.72 $Y=1.565
+ $X2=0.925 $Y2=1.565
r52 15 16 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=0.24 $Y=1.565
+ $X2=0.72 $Y2=1.565
r53 11 25 24.2915 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.015 $Y=1.35
+ $X2=1.015 $Y2=1.557
r54 11 13 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.015 $Y=1.35
+ $X2=1.015 $Y2=0.74
r55 8 24 24.2915 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=1 $Y=1.765 $X2=1
+ $Y2=1.557
r56 8 10 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1 $Y=1.765 $X2=1
+ $Y2=2.4
r57 5 20 24.2915 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=0.51 $Y=1.765
+ $X2=0.51 $Y2=1.557
r58 5 7 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.51 $Y=1.765
+ $X2=0.51 $Y2=2.4
r59 1 19 24.2915 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.495 $Y=1.35
+ $X2=0.495 $Y2=1.557
r60 1 3 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=0.495 $Y=1.35
+ $X2=0.495 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HS__NAND4_2%C 3 5 7 10 12 14 15 16 19 21 22
c54 22 0 8.45585e-20 $X=2.275 $Y=1.515
c55 19 0 6.47788e-20 $X=2.05 $Y=1.515
c56 12 0 3.22126e-20 $X=1.96 $Y=1.765
c57 5 0 2.97865e-19 $X=1.49 $Y=1.765
c58 3 0 1.87767e-19 $X=1.445 $Y=0.74
r59 28 30 3.28338 $w=3.67e-07 $l=2.5e-08 $layer=POLY_cond $X=1.935 $Y=1.557
+ $X2=1.96 $Y2=1.557
r60 28 29 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.935
+ $Y=1.515 $X2=1.935 $Y2=1.515
r61 26 28 7.88011 $w=3.67e-07 $l=6e-08 $layer=POLY_cond $X=1.875 $Y=1.557
+ $X2=1.935 $Y2=1.557
r62 25 26 50.564 $w=3.67e-07 $l=3.85e-07 $layer=POLY_cond $X=1.49 $Y=1.557
+ $X2=1.875 $Y2=1.557
r63 24 25 5.91008 $w=3.67e-07 $l=4.5e-08 $layer=POLY_cond $X=1.445 $Y=1.557
+ $X2=1.49 $Y2=1.557
r64 21 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.275
+ $Y=1.515 $X2=2.275 $Y2=1.515
r65 19 30 12.4159 $w=3.67e-07 $l=1.08995e-07 $layer=POLY_cond $X=2.05 $Y=1.515
+ $X2=1.96 $Y2=1.557
r66 19 21 39.3438 $w=3.3e-07 $l=2.25e-07 $layer=POLY_cond $X=2.05 $Y=1.515
+ $X2=2.275 $Y2=1.515
r67 16 22 3.08211 $w=4.28e-07 $l=1.15e-07 $layer=LI1_cond $X=2.16 $Y=1.565
+ $X2=2.275 $Y2=1.565
r68 16 29 6.03022 $w=4.28e-07 $l=2.25e-07 $layer=LI1_cond $X=2.16 $Y=1.565
+ $X2=1.935 $Y2=1.565
r69 15 29 6.83426 $w=4.28e-07 $l=2.55e-07 $layer=LI1_cond $X=1.68 $Y=1.565
+ $X2=1.935 $Y2=1.565
r70 12 30 23.77 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=1.96 $Y=1.765
+ $X2=1.96 $Y2=1.557
r71 12 14 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.96 $Y=1.765
+ $X2=1.96 $Y2=2.4
r72 8 26 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.875 $Y=1.35
+ $X2=1.875 $Y2=1.557
r73 8 10 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.875 $Y=1.35
+ $X2=1.875 $Y2=0.74
r74 5 25 23.77 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=1.49 $Y=1.765 $X2=1.49
+ $Y2=1.557
r75 5 7 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.49 $Y=1.765
+ $X2=1.49 $Y2=2.4
r76 1 24 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.445 $Y=1.35
+ $X2=1.445 $Y2=1.557
r77 1 3 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.445 $Y=1.35
+ $X2=1.445 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HS__NAND4_2%B 1 3 6 8 10 13 15 16 23
c54 16 0 1.06018e-19 $X=3.6 $Y=1.665
c55 13 0 1.79791e-19 $X=3.365 $Y=0.74
c56 8 0 1.34333e-19 $X=3.22 $Y=1.765
c57 1 0 6.86776e-20 $X=2.77 $Y=1.765
r58 23 25 11.7243 $w=3.7e-07 $l=9e-08 $layer=POLY_cond $X=3.275 $Y=1.557
+ $X2=3.365 $Y2=1.557
r59 23 24 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.275
+ $Y=1.515 $X2=3.275 $Y2=1.515
r60 21 23 7.16487 $w=3.7e-07 $l=5.5e-08 $layer=POLY_cond $X=3.22 $Y=1.557
+ $X2=3.275 $Y2=1.557
r61 20 21 37.127 $w=3.7e-07 $l=2.85e-07 $layer=POLY_cond $X=2.935 $Y=1.557
+ $X2=3.22 $Y2=1.557
r62 19 20 21.4946 $w=3.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.77 $Y=1.557
+ $X2=2.935 $Y2=1.557
r63 16 24 8.71033 $w=4.28e-07 $l=3.25e-07 $layer=LI1_cond $X=3.6 $Y=1.565
+ $X2=3.275 $Y2=1.565
r64 15 24 4.15415 $w=4.28e-07 $l=1.55e-07 $layer=LI1_cond $X=3.12 $Y=1.565
+ $X2=3.275 $Y2=1.565
r65 11 25 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.365 $Y=1.35
+ $X2=3.365 $Y2=1.557
r66 11 13 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=3.365 $Y=1.35
+ $X2=3.365 $Y2=0.74
r67 8 21 23.9667 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=3.22 $Y=1.765
+ $X2=3.22 $Y2=1.557
r68 8 10 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.22 $Y=1.765
+ $X2=3.22 $Y2=2.4
r69 4 20 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.935 $Y=1.35
+ $X2=2.935 $Y2=1.557
r70 4 6 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.935 $Y=1.35
+ $X2=2.935 $Y2=0.74
r71 1 19 23.9667 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=2.77 $Y=1.765
+ $X2=2.77 $Y2=1.557
r72 1 3 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.77 $Y=1.765
+ $X2=2.77 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_HS__NAND4_2%A 1 3 6 8 10 13 15 21 22
c48 8 0 1.89481e-19 $X=4.23 $Y=1.765
c49 6 0 1.79791e-19 $X=3.795 $Y=0.74
r50 22 23 1.95935 $w=3.69e-07 $l=1.5e-08 $layer=POLY_cond $X=4.23 $Y=1.557
+ $X2=4.245 $Y2=1.557
r51 20 22 23.5122 $w=3.69e-07 $l=1.8e-07 $layer=POLY_cond $X=4.05 $Y=1.557
+ $X2=4.23 $Y2=1.557
r52 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.05
+ $Y=1.515 $X2=4.05 $Y2=1.515
r53 18 20 33.3089 $w=3.69e-07 $l=2.55e-07 $layer=POLY_cond $X=3.795 $Y=1.557
+ $X2=4.05 $Y2=1.557
r54 17 18 1.95935 $w=3.69e-07 $l=1.5e-08 $layer=POLY_cond $X=3.78 $Y=1.557
+ $X2=3.795 $Y2=1.557
r55 15 21 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=4.05 $Y=1.665
+ $X2=4.05 $Y2=1.515
r56 11 23 23.9013 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.245 $Y=1.35
+ $X2=4.245 $Y2=1.557
r57 11 13 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=4.245 $Y=1.35
+ $X2=4.245 $Y2=0.74
r58 8 22 23.9013 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=4.23 $Y=1.765
+ $X2=4.23 $Y2=1.557
r59 8 10 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=4.23 $Y=1.765
+ $X2=4.23 $Y2=2.4
r60 4 18 23.9013 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.795 $Y=1.35
+ $X2=3.795 $Y2=1.557
r61 4 6 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=3.795 $Y=1.35
+ $X2=3.795 $Y2=0.74
r62 1 17 23.9013 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=3.78 $Y=1.765
+ $X2=3.78 $Y2=1.557
r63 1 3 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.78 $Y=1.765
+ $X2=3.78 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_HS__NAND4_2%VPWR 1 2 3 4 5 16 18 24 26 30 34 36 38 41 42
+ 43 45 54 62 65 69
r71 68 69 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r72 65 66 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r73 63 66 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.16 $Y2=3.33
r74 62 63 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r75 59 60 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r76 57 69 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=4.56 $Y2=3.33
r77 56 57 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r78 54 68 4.61575 $w=1.7e-07 $l=2.52e-07 $layer=LI1_cond $X=4.295 $Y=3.33
+ $X2=4.547 $Y2=3.33
r79 54 56 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=4.295 $Y=3.33
+ $X2=4.08 $Y2=3.33
r80 53 57 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=4.08 $Y2=3.33
r81 52 53 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r82 50 65 12.1981 $w=1.7e-07 $l=2.85e-07 $layer=LI1_cond $X=2.65 $Y=3.33
+ $X2=2.365 $Y2=3.33
r83 50 52 30.6631 $w=1.68e-07 $l=4.7e-07 $layer=LI1_cond $X=2.65 $Y=3.33
+ $X2=3.12 $Y2=3.33
r84 49 63 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r85 49 60 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r86 48 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r87 46 59 4.78727 $w=1.7e-07 $l=2.25e-07 $layer=LI1_cond $X=0.45 $Y=3.33
+ $X2=0.225 $Y2=3.33
r88 46 48 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=0.45 $Y=3.33 $X2=0.72
+ $Y2=3.33
r89 45 62 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.07 $Y=3.33
+ $X2=1.235 $Y2=3.33
r90 45 48 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=1.07 $Y=3.33
+ $X2=0.72 $Y2=3.33
r91 43 53 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=2.4 $Y=3.33
+ $X2=3.12 $Y2=3.33
r92 43 66 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.4 $Y=3.33
+ $X2=2.16 $Y2=3.33
r93 41 52 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=3.33 $Y=3.33
+ $X2=3.12 $Y2=3.33
r94 41 42 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.33 $Y=3.33
+ $X2=3.495 $Y2=3.33
r95 40 56 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=3.66 $Y=3.33
+ $X2=4.08 $Y2=3.33
r96 40 42 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.66 $Y=3.33
+ $X2=3.495 $Y2=3.33
r97 36 68 3.15043 $w=3.3e-07 $l=1.22327e-07 $layer=LI1_cond $X=4.46 $Y=3.245
+ $X2=4.547 $Y2=3.33
r98 36 38 29.1603 $w=3.28e-07 $l=8.35e-07 $layer=LI1_cond $X=4.46 $Y=3.245
+ $X2=4.46 $Y2=2.41
r99 32 42 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.495 $Y=3.245
+ $X2=3.495 $Y2=3.33
r100 32 34 29.1603 $w=3.28e-07 $l=8.35e-07 $layer=LI1_cond $X=3.495 $Y=3.245
+ $X2=3.495 $Y2=2.41
r101 28 65 2.39972 $w=5.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.365 $Y=3.245
+ $X2=2.365 $Y2=3.33
r102 28 30 16.5772 $w=5.68e-07 $l=7.9e-07 $layer=LI1_cond $X=2.365 $Y=3.245
+ $X2=2.365 $Y2=2.455
r103 27 62 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.4 $Y=3.33
+ $X2=1.235 $Y2=3.33
r104 26 65 12.1981 $w=1.7e-07 $l=2.85e-07 $layer=LI1_cond $X=2.08 $Y=3.33
+ $X2=2.365 $Y2=3.33
r105 26 27 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=2.08 $Y=3.33
+ $X2=1.4 $Y2=3.33
r106 22 62 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.235 $Y=3.245
+ $X2=1.235 $Y2=3.33
r107 22 24 29.1603 $w=3.28e-07 $l=8.35e-07 $layer=LI1_cond $X=1.235 $Y=3.245
+ $X2=1.235 $Y2=2.41
r108 18 21 26.833 $w=3.33e-07 $l=7.8e-07 $layer=LI1_cond $X=0.282 $Y=2.035
+ $X2=0.282 $Y2=2.815
r109 16 59 3.0213 $w=3.35e-07 $l=1.09864e-07 $layer=LI1_cond $X=0.282 $Y=3.245
+ $X2=0.225 $Y2=3.33
r110 16 21 14.7926 $w=3.33e-07 $l=4.3e-07 $layer=LI1_cond $X=0.282 $Y=3.245
+ $X2=0.282 $Y2=2.815
r111 5 38 300 $w=1.7e-07 $l=6.42845e-07 $layer=licon1_PDIFF $count=2 $X=4.305
+ $Y=1.84 $X2=4.46 $Y2=2.41
r112 4 34 300 $w=1.7e-07 $l=6.62495e-07 $layer=licon1_PDIFF $count=2 $X=3.295
+ $Y=1.84 $X2=3.495 $Y2=2.41
r113 3 30 150 $w=1.7e-07 $l=8.3179e-07 $layer=licon1_PDIFF $count=4 $X=2.035
+ $Y=1.84 $X2=2.545 $Y2=2.455
r114 2 24 300 $w=1.7e-07 $l=6.45058e-07 $layer=licon1_PDIFF $count=2 $X=1.075
+ $Y=1.84 $X2=1.235 $Y2=2.41
r115 1 21 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.815
r116 1 18 400 $w=1.7e-07 $l=2.57488e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.035
.ends

.subckt PM_SKY130_FD_SC_HS__NAND4_2%Y 1 2 3 4 5 16 18 20 24 26 30 32 36 40 42 44
+ 45 49 51 53 55 56 57
c87 53 0 1.34333e-19 $X=4.005 $Y=2.035
c88 45 0 1.79791e-19 $X=4.175 $Y=1.095
c89 36 0 1.80454e-19 $X=4.005 $Y=2.43
c90 24 0 1.99665e-19 $X=1.735 $Y=2.43
c91 18 0 3.32865e-19 $X=0.735 $Y=2.815
r92 56 57 10.2753 $w=3.98e-07 $l=2.85e-07 $layer=LI1_cond $X=4.56 $Y=1.665
+ $X2=4.56 $Y2=1.95
r93 55 56 18.5393 $w=2.28e-07 $l=3.7e-07 $layer=LI1_cond $X=4.56 $Y=1.295
+ $X2=4.56 $Y2=1.665
r94 54 55 5.76222 $w=2.28e-07 $l=1.15e-07 $layer=LI1_cond $X=4.56 $Y=1.18
+ $X2=4.56 $Y2=1.295
r95 44 54 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=4.445 $Y=1.095
+ $X2=4.56 $Y2=1.18
r96 44 45 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=4.445 $Y=1.095
+ $X2=4.175 $Y2=1.095
r97 43 53 7.27964 $w=1.85e-07 $l=1.43e-07 $layer=LI1_cond $X=4.125 $Y=2.05
+ $X2=3.982 $Y2=2.05
r98 42 57 3.66916 $w=2e-07 $l=1.15e-07 $layer=LI1_cond $X=4.445 $Y=2.05 $X2=4.56
+ $Y2=2.05
r99 42 43 17.7455 $w=1.98e-07 $l=3.2e-07 $layer=LI1_cond $X=4.445 $Y=2.05
+ $X2=4.125 $Y2=2.05
r100 38 45 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.01 $Y=1.01
+ $X2=4.175 $Y2=1.095
r101 38 40 6.9845 $w=3.28e-07 $l=2e-07 $layer=LI1_cond $X=4.01 $Y=1.01 $X2=4.01
+ $Y2=0.81
r102 34 53 0.156385 $w=2.85e-07 $l=1e-07 $layer=LI1_cond $X=3.982 $Y=2.15
+ $X2=3.982 $Y2=2.05
r103 34 36 11.3222 $w=2.83e-07 $l=2.8e-07 $layer=LI1_cond $X=3.982 $Y=2.15
+ $X2=3.982 $Y2=2.43
r104 33 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.16 $Y=2.035
+ $X2=2.995 $Y2=2.035
r105 32 53 7.27964 $w=1.85e-07 $l=1.49312e-07 $layer=LI1_cond $X=3.84 $Y=2.035
+ $X2=3.982 $Y2=2.05
r106 32 33 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=3.84 $Y=2.035
+ $X2=3.16 $Y2=2.035
r107 28 51 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.995 $Y=2.12
+ $X2=2.995 $Y2=2.035
r108 28 30 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=2.995 $Y=2.12
+ $X2=2.995 $Y2=2.815
r109 27 49 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.9 $Y=2.035
+ $X2=1.735 $Y2=2.035
r110 26 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.83 $Y=2.035
+ $X2=2.995 $Y2=2.035
r111 26 27 60.6738 $w=1.68e-07 $l=9.3e-07 $layer=LI1_cond $X=2.83 $Y=2.035
+ $X2=1.9 $Y2=2.035
r112 22 49 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.735 $Y=2.12
+ $X2=1.735 $Y2=2.035
r113 22 24 10.826 $w=3.28e-07 $l=3.1e-07 $layer=LI1_cond $X=1.735 $Y=2.12
+ $X2=1.735 $Y2=2.43
r114 21 47 4.42198 $w=1.7e-07 $l=1.33e-07 $layer=LI1_cond $X=0.9 $Y=2.035
+ $X2=0.767 $Y2=2.035
r115 20 49 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.57 $Y=2.035
+ $X2=1.735 $Y2=2.035
r116 20 21 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.57 $Y=2.035
+ $X2=0.9 $Y2=2.035
r117 16 47 2.82608 $w=2.65e-07 $l=8.5e-08 $layer=LI1_cond $X=0.767 $Y=2.12
+ $X2=0.767 $Y2=2.035
r118 16 18 30.2244 $w=2.63e-07 $l=6.95e-07 $layer=LI1_cond $X=0.767 $Y=2.12
+ $X2=0.767 $Y2=2.815
r119 5 53 600 $w=1.7e-07 $l=2.59374e-07 $layer=licon1_PDIFF $count=1 $X=3.855
+ $Y=1.84 $X2=4.005 $Y2=2.035
r120 5 36 300 $w=1.7e-07 $l=6.60757e-07 $layer=licon1_PDIFF $count=2 $X=3.855
+ $Y=1.84 $X2=4.005 $Y2=2.43
r121 4 51 400 $w=1.7e-07 $l=2.59374e-07 $layer=licon1_PDIFF $count=1 $X=2.845
+ $Y=1.84 $X2=2.995 $Y2=2.035
r122 4 30 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=2.845
+ $Y=1.84 $X2=2.995 $Y2=2.815
r123 3 49 600 $w=1.7e-07 $l=2.66786e-07 $layer=licon1_PDIFF $count=1 $X=1.565
+ $Y=1.84 $X2=1.735 $Y2=2.035
r124 3 24 300 $w=1.7e-07 $l=6.69627e-07 $layer=licon1_PDIFF $count=2 $X=1.565
+ $Y=1.84 $X2=1.735 $Y2=2.43
r125 2 47 400 $w=1.7e-07 $l=3.4187e-07 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=1.84 $X2=0.735 $Y2=2.115
r126 2 18 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=1.84 $X2=0.735 $Y2=2.815
r127 1 40 182 $w=1.7e-07 $l=5.05173e-07 $layer=licon1_NDIFF $count=1 $X=3.87
+ $Y=0.37 $X2=4.01 $Y2=0.81
.ends

.subckt PM_SKY130_FD_SC_HS__NAND4_2%A_27_74# 1 2 3 12 14 15 20 21 24
r37 22 24 5.93683 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=2.16 $Y=0.425
+ $X2=2.16 $Y2=0.595
r38 20 22 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.995 $Y=0.34
+ $X2=2.16 $Y2=0.425
r39 20 21 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.995 $Y=0.34
+ $X2=1.315 $Y2=0.34
r40 17 19 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=1.23 $Y=1.01
+ $X2=1.23 $Y2=0.515
r41 16 21 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.23 $Y=0.425
+ $X2=1.315 $Y2=0.34
r42 16 19 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=1.23 $Y=0.425 $X2=1.23
+ $Y2=0.515
r43 14 17 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.145 $Y=1.095
+ $X2=1.23 $Y2=1.01
r44 14 15 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=1.145 $Y=1.095
+ $X2=0.445 $Y2=1.095
r45 10 15 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.28 $Y=1.01
+ $X2=0.445 $Y2=1.095
r46 10 12 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=0.28 $Y=1.01
+ $X2=0.28 $Y2=0.515
r47 3 24 182 $w=1.7e-07 $l=3.1285e-07 $layer=licon1_NDIFF $count=1 $X=1.95
+ $Y=0.37 $X2=2.16 $Y2=0.595
r48 2 19 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.09
+ $Y=0.37 $X2=1.23 $Y2=0.515
r49 1 12 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__NAND4_2%VGND 1 6 8 10 20 21 24
c41 6 0 1.87767e-19 $X=0.78 $Y=0.635
r42 24 25 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r43 20 21 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r44 18 25 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r45 17 20 219.209 $w=1.68e-07 $l=3.36e-06 $layer=LI1_cond $X=1.2 $Y=0 $X2=4.56
+ $Y2=0
r46 17 18 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r47 15 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.945 $Y=0 $X2=0.78
+ $Y2=0
r48 15 17 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.945 $Y=0 $X2=1.2
+ $Y2=0
r49 13 25 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r50 12 13 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r51 10 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.615 $Y=0 $X2=0.78
+ $Y2=0
r52 10 12 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=0.615 $Y=0 $X2=0.24
+ $Y2=0
r53 8 21 0.602067 $w=4.9e-07 $l=2.16e-06 $layer=MET1_cond $X=2.4 $Y=0 $X2=4.56
+ $Y2=0
r54 8 18 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=2.4 $Y=0 $X2=1.2
+ $Y2=0
r55 4 24 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.78 $Y=0.085 $X2=0.78
+ $Y2=0
r56 4 6 19.2074 $w=3.28e-07 $l=5.5e-07 $layer=LI1_cond $X=0.78 $Y=0.085 $X2=0.78
+ $Y2=0.635
r57 1 6 182 $w=1.7e-07 $l=3.54789e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.37 $X2=0.78 $Y2=0.635
.ends

.subckt PM_SKY130_FD_SC_HS__NAND4_2%A_304_74# 1 2 9 11 12 15
c30 12 0 8.01953e-20 $X=1.825 $Y=1.095
c31 11 0 1.79791e-19 $X=2.985 $Y=1.095
r32 13 15 6.9845 $w=3.28e-07 $l=2e-07 $layer=LI1_cond $X=3.15 $Y=1.01 $X2=3.15
+ $Y2=0.81
r33 11 13 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.985 $Y=1.095
+ $X2=3.15 $Y2=1.01
r34 11 12 75.6791 $w=1.68e-07 $l=1.16e-06 $layer=LI1_cond $X=2.985 $Y=1.095
+ $X2=1.825 $Y2=1.095
r35 7 12 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.66 $Y=1.01
+ $X2=1.825 $Y2=1.095
r36 7 9 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=1.66 $Y=1.01 $X2=1.66
+ $Y2=0.86
r37 2 15 182 $w=1.7e-07 $l=5.05173e-07 $layer=licon1_NDIFF $count=1 $X=3.01
+ $Y=0.37 $X2=3.15 $Y2=0.81
r38 1 9 182 $w=1.7e-07 $l=5.55608e-07 $layer=licon1_NDIFF $count=1 $X=1.52
+ $Y=0.37 $X2=1.66 $Y2=0.86
.ends

.subckt PM_SKY130_FD_SC_HS__NAND4_2%A_515_74# 1 2 3 12 14 15 18 20 24 26
r37 22 24 5.93683 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=4.51 $Y=0.425
+ $X2=4.51 $Y2=0.595
r38 21 26 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=3.675 $Y=0.34
+ $X2=3.58 $Y2=0.34
r39 20 22 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.345 $Y=0.34
+ $X2=4.51 $Y2=0.425
r40 20 21 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.345 $Y=0.34
+ $X2=3.675 $Y2=0.34
r41 16 26 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=3.58 $Y=0.425
+ $X2=3.58 $Y2=0.34
r42 16 18 5.25359 $w=1.88e-07 $l=9e-08 $layer=LI1_cond $X=3.58 $Y=0.425 $X2=3.58
+ $Y2=0.515
r43 14 26 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=3.485 $Y=0.34
+ $X2=3.58 $Y2=0.34
r44 14 15 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.485 $Y=0.34
+ $X2=2.815 $Y2=0.34
r45 10 15 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=2.685 $Y=0.425
+ $X2=2.815 $Y2=0.34
r46 10 12 8.86495 $w=2.58e-07 $l=2e-07 $layer=LI1_cond $X=2.685 $Y=0.425
+ $X2=2.685 $Y2=0.625
r47 3 24 182 $w=1.7e-07 $l=3.05573e-07 $layer=licon1_NDIFF $count=1 $X=4.32
+ $Y=0.37 $X2=4.51 $Y2=0.595
r48 2 18 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.44
+ $Y=0.37 $X2=3.58 $Y2=0.515
r49 1 12 182 $w=1.7e-07 $l=3.19374e-07 $layer=licon1_NDIFF $count=1 $X=2.575
+ $Y=0.37 $X2=2.72 $Y2=0.625
.ends

