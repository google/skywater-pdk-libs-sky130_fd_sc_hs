* File: sky130_fd_sc_hs__or2_2.pxi.spice
* Created: Tue Sep  1 20:19:54 2020
* 
x_PM_SKY130_FD_SC_HS__OR2_2%B N_B_c_48_n N_B_M1004_g N_B_c_49_n N_B_M1001_g B
+ PM_SKY130_FD_SC_HS__OR2_2%B
x_PM_SKY130_FD_SC_HS__OR2_2%A N_A_c_71_n N_A_M1005_g N_A_M1006_g A A N_A_c_73_n
+ PM_SKY130_FD_SC_HS__OR2_2%A
x_PM_SKY130_FD_SC_HS__OR2_2%A_27_368# N_A_27_368#_M1004_d N_A_27_368#_M1001_s
+ N_A_27_368#_M1003_g N_A_27_368#_c_121_n N_A_27_368#_M1000_g
+ N_A_27_368#_M1007_g N_A_27_368#_c_122_n N_A_27_368#_M1002_g
+ N_A_27_368#_c_123_n N_A_27_368#_c_124_n N_A_27_368#_c_133_n
+ N_A_27_368#_c_114_n N_A_27_368#_c_115_n N_A_27_368#_c_116_n
+ N_A_27_368#_c_117_n N_A_27_368#_c_126_n N_A_27_368#_c_118_n
+ N_A_27_368#_c_128_n N_A_27_368#_c_160_p N_A_27_368#_c_119_n
+ N_A_27_368#_c_120_n PM_SKY130_FD_SC_HS__OR2_2%A_27_368#
x_PM_SKY130_FD_SC_HS__OR2_2%VPWR N_VPWR_M1005_d N_VPWR_M1002_s N_VPWR_c_212_n
+ N_VPWR_c_213_n N_VPWR_c_214_n VPWR N_VPWR_c_215_n N_VPWR_c_216_n
+ N_VPWR_c_217_n N_VPWR_c_211_n PM_SKY130_FD_SC_HS__OR2_2%VPWR
x_PM_SKY130_FD_SC_HS__OR2_2%X N_X_M1003_s N_X_M1000_d X X X X X
+ PM_SKY130_FD_SC_HS__OR2_2%X
x_PM_SKY130_FD_SC_HS__OR2_2%VGND N_VGND_M1004_s N_VGND_M1006_d N_VGND_M1007_d
+ N_VGND_c_268_n N_VGND_c_269_n N_VGND_c_270_n N_VGND_c_271_n N_VGND_c_272_n
+ VGND N_VGND_c_273_n N_VGND_c_274_n N_VGND_c_275_n N_VGND_c_276_n
+ PM_SKY130_FD_SC_HS__OR2_2%VGND
cc_1 VNB N_B_c_48_n 0.0205953f $X=-0.19 $Y=-0.245 $X2=0.49 $Y2=1.22
cc_2 VNB N_B_c_49_n 0.0677471f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.765
cc_3 VNB B 0.00785817f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_4 VNB N_A_c_71_n 0.0238748f $X=-0.19 $Y=-0.245 $X2=0.49 $Y2=1.22
cc_5 VNB N_A_M1006_g 0.0238971f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.34
cc_6 VNB N_A_c_73_n 0.00542652f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_7 VNB N_A_27_368#_M1003_g 0.0218443f $X=-0.19 $Y=-0.245 $X2=0.345 $Y2=1.385
cc_8 VNB N_A_27_368#_M1007_g 0.0260244f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A_27_368#_c_114_n 0.00241395f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_27_368#_c_115_n 0.00412876f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_27_368#_c_116_n 0.00278905f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_27_368#_c_117_n 0.00349145f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_27_368#_c_118_n 0.00121168f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_27_368#_c_119_n 0.00841735f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_27_368#_c_120_n 0.090597f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_VPWR_c_211_n 0.103974f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB X 0.00356546f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_18 VNB N_VGND_c_268_n 0.0120573f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.385
cc_19 VNB N_VGND_c_269_n 0.0358796f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.295
cc_20 VNB N_VGND_c_270_n 0.00647256f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_VGND_c_271_n 0.0117383f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_VGND_c_272_n 0.0441433f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_VGND_c_273_n 0.0175968f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_VGND_c_274_n 0.0168532f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_VGND_c_275_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_VGND_c_276_n 0.164475f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VPB N_B_c_49_n 0.0294453f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.765
cc_28 VPB N_A_c_71_n 0.0254102f $X=-0.19 $Y=1.66 $X2=0.49 $Y2=1.22
cc_29 VPB N_A_c_73_n 0.0027795f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_30 VPB N_A_27_368#_c_121_n 0.0169202f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.385
cc_31 VPB N_A_27_368#_c_122_n 0.0173077f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_32 VPB N_A_27_368#_c_123_n 0.0215662f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_33 VPB N_A_27_368#_c_124_n 0.017509f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_34 VPB N_A_27_368#_c_117_n 0.00111575f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_35 VPB N_A_27_368#_c_126_n 0.00748573f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_36 VPB N_A_27_368#_c_118_n 0.0246729f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_37 VPB N_A_27_368#_c_128_n 0.0071123f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_38 VPB N_A_27_368#_c_120_n 0.0134445f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_39 VPB N_VPWR_c_212_n 0.0104361f $X=-0.19 $Y=1.66 $X2=0.345 $Y2=1.385
cc_40 VPB N_VPWR_c_213_n 0.0120106f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.385
cc_41 VPB N_VPWR_c_214_n 0.0210177f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_42 VPB N_VPWR_c_215_n 0.033055f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_43 VPB N_VPWR_c_216_n 0.0183953f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_44 VPB N_VPWR_c_217_n 0.00614127f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_45 VPB N_VPWR_c_211_n 0.0602725f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_46 VPB X 0.00210362f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.21
cc_47 VPB X 4.20601e-19 $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.385
cc_48 N_B_c_49_n N_A_c_71_n 0.087086f $X=0.495 $Y=1.765 $X2=-0.19 $Y2=-0.245
cc_49 N_B_c_48_n N_A_M1006_g 0.00980177f $X=0.49 $Y=1.22 $X2=0 $Y2=0
cc_50 N_B_c_49_n N_A_M1006_g 0.00662485f $X=0.495 $Y=1.765 $X2=0 $Y2=0
cc_51 B N_A_M1006_g 7.98305e-19 $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_52 N_B_c_49_n N_A_c_73_n 0.0108231f $X=0.495 $Y=1.765 $X2=0 $Y2=0
cc_53 B N_A_c_73_n 0.0161951f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_54 N_B_c_49_n N_A_27_368#_c_123_n 0.0093155f $X=0.495 $Y=1.765 $X2=0 $Y2=0
cc_55 B N_A_27_368#_c_123_n 0.0197435f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_56 N_B_c_49_n N_A_27_368#_c_124_n 0.00695804f $X=0.495 $Y=1.765 $X2=0 $Y2=0
cc_57 N_B_c_49_n N_A_27_368#_c_133_n 0.0127906f $X=0.495 $Y=1.765 $X2=0 $Y2=0
cc_58 N_B_c_48_n N_A_27_368#_c_116_n 0.00218762f $X=0.49 $Y=1.22 $X2=0 $Y2=0
cc_59 N_B_c_49_n N_A_27_368#_c_128_n 2.24111e-19 $X=0.495 $Y=1.765 $X2=0 $Y2=0
cc_60 N_B_c_49_n N_VPWR_c_215_n 0.00481995f $X=0.495 $Y=1.765 $X2=0 $Y2=0
cc_61 N_B_c_49_n N_VPWR_c_211_n 0.00508379f $X=0.495 $Y=1.765 $X2=0 $Y2=0
cc_62 N_B_c_48_n N_VGND_c_269_n 0.0148675f $X=0.49 $Y=1.22 $X2=0 $Y2=0
cc_63 N_B_c_49_n N_VGND_c_269_n 0.00198489f $X=0.495 $Y=1.765 $X2=0 $Y2=0
cc_64 B N_VGND_c_269_n 0.0246129f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_65 N_B_c_48_n N_VGND_c_273_n 0.00421418f $X=0.49 $Y=1.22 $X2=0 $Y2=0
cc_66 N_B_c_48_n N_VGND_c_276_n 0.00432128f $X=0.49 $Y=1.22 $X2=0 $Y2=0
cc_67 N_A_M1006_g N_A_27_368#_M1003_g 0.0224491f $X=0.92 $Y=0.79 $X2=0 $Y2=0
cc_68 N_A_c_71_n N_A_27_368#_c_121_n 0.0287993f $X=0.885 $Y=1.765 $X2=0 $Y2=0
cc_69 N_A_c_73_n N_A_27_368#_c_121_n 0.00112187f $X=0.96 $Y=1.515 $X2=0 $Y2=0
cc_70 N_A_c_71_n N_A_27_368#_c_123_n 0.00106611f $X=0.885 $Y=1.765 $X2=0 $Y2=0
cc_71 N_A_c_73_n N_A_27_368#_c_123_n 0.013208f $X=0.96 $Y=1.515 $X2=0 $Y2=0
cc_72 N_A_c_71_n N_A_27_368#_c_124_n 0.00140708f $X=0.885 $Y=1.765 $X2=0 $Y2=0
cc_73 N_A_c_71_n N_A_27_368#_c_133_n 0.0140743f $X=0.885 $Y=1.765 $X2=0 $Y2=0
cc_74 N_A_c_73_n N_A_27_368#_c_133_n 0.0238741f $X=0.96 $Y=1.515 $X2=0 $Y2=0
cc_75 N_A_M1006_g N_A_27_368#_c_114_n 0.00781094f $X=0.92 $Y=0.79 $X2=0 $Y2=0
cc_76 N_A_c_71_n N_A_27_368#_c_115_n 0.00338829f $X=0.885 $Y=1.765 $X2=0 $Y2=0
cc_77 N_A_M1006_g N_A_27_368#_c_115_n 0.0113358f $X=0.92 $Y=0.79 $X2=0 $Y2=0
cc_78 N_A_c_73_n N_A_27_368#_c_115_n 0.0134037f $X=0.96 $Y=1.515 $X2=0 $Y2=0
cc_79 N_A_c_71_n N_A_27_368#_c_116_n 3.92011e-19 $X=0.885 $Y=1.765 $X2=0 $Y2=0
cc_80 N_A_M1006_g N_A_27_368#_c_116_n 0.00137818f $X=0.92 $Y=0.79 $X2=0 $Y2=0
cc_81 N_A_c_73_n N_A_27_368#_c_116_n 0.0229711f $X=0.96 $Y=1.515 $X2=0 $Y2=0
cc_82 N_A_c_71_n N_A_27_368#_c_117_n 0.00669135f $X=0.885 $Y=1.765 $X2=0 $Y2=0
cc_83 N_A_M1006_g N_A_27_368#_c_117_n 0.00340254f $X=0.92 $Y=0.79 $X2=0 $Y2=0
cc_84 N_A_c_73_n N_A_27_368#_c_117_n 0.0625707f $X=0.96 $Y=1.515 $X2=0 $Y2=0
cc_85 N_A_c_71_n N_A_27_368#_c_120_n 0.0232354f $X=0.885 $Y=1.765 $X2=0 $Y2=0
cc_86 N_A_M1006_g N_A_27_368#_c_120_n 0.00157274f $X=0.92 $Y=0.79 $X2=0 $Y2=0
cc_87 N_A_c_73_n N_A_27_368#_c_120_n 5.36155e-19 $X=0.96 $Y=1.515 $X2=0 $Y2=0
cc_88 N_A_c_73_n A_114_368# 0.00143032f $X=0.96 $Y=1.515 $X2=-0.19 $Y2=-0.245
cc_89 N_A_c_73_n N_VPWR_M1005_d 0.00311293f $X=0.96 $Y=1.515 $X2=-0.19
+ $Y2=-0.245
cc_90 N_A_c_71_n N_VPWR_c_212_n 0.00595217f $X=0.885 $Y=1.765 $X2=0 $Y2=0
cc_91 N_A_c_71_n N_VPWR_c_215_n 0.0049405f $X=0.885 $Y=1.765 $X2=0 $Y2=0
cc_92 N_A_c_71_n N_VPWR_c_211_n 0.00508379f $X=0.885 $Y=1.765 $X2=0 $Y2=0
cc_93 N_A_M1006_g N_VGND_c_269_n 5.06989e-19 $X=0.92 $Y=0.79 $X2=0 $Y2=0
cc_94 N_A_M1006_g N_VGND_c_270_n 0.00365474f $X=0.92 $Y=0.79 $X2=0 $Y2=0
cc_95 N_A_M1006_g N_VGND_c_273_n 0.00485498f $X=0.92 $Y=0.79 $X2=0 $Y2=0
cc_96 N_A_M1006_g N_VGND_c_276_n 0.00514438f $X=0.92 $Y=0.79 $X2=0 $Y2=0
cc_97 N_A_27_368#_c_133_n A_114_368# 0.00387262f $X=1.215 $Y=2.405 $X2=-0.19
+ $Y2=-0.245
cc_98 N_A_27_368#_c_133_n N_VPWR_M1005_d 0.00759042f $X=1.215 $Y=2.405 $X2=-0.19
+ $Y2=-0.245
cc_99 N_A_27_368#_c_117_n N_VPWR_M1005_d 0.00476863f $X=1.3 $Y=2.32 $X2=-0.19
+ $Y2=-0.245
cc_100 N_A_27_368#_c_160_p N_VPWR_M1005_d 8.40529e-19 $X=1.3 $Y=2.405 $X2=-0.19
+ $Y2=-0.245
cc_101 N_A_27_368#_c_126_n N_VPWR_M1002_s 0.00536103f $X=2.125 $Y=2.405 $X2=0
+ $Y2=0
cc_102 N_A_27_368#_c_118_n N_VPWR_M1002_s 0.00859407f $X=2.21 $Y=2.32 $X2=0
+ $Y2=0
cc_103 N_A_27_368#_c_121_n N_VPWR_c_212_n 0.0107345f $X=1.425 $Y=1.765 $X2=0
+ $Y2=0
cc_104 N_A_27_368#_c_122_n N_VPWR_c_212_n 0.00128695f $X=1.895 $Y=1.765 $X2=0
+ $Y2=0
cc_105 N_A_27_368#_c_124_n N_VPWR_c_212_n 0.00577095f $X=0.27 $Y=2.695 $X2=0
+ $Y2=0
cc_106 N_A_27_368#_c_133_n N_VPWR_c_212_n 0.0142094f $X=1.215 $Y=2.405 $X2=0
+ $Y2=0
cc_107 N_A_27_368#_c_160_p N_VPWR_c_212_n 0.00793448f $X=1.3 $Y=2.405 $X2=0
+ $Y2=0
cc_108 N_A_27_368#_c_121_n N_VPWR_c_214_n 0.00128695f $X=1.425 $Y=1.765 $X2=0
+ $Y2=0
cc_109 N_A_27_368#_c_122_n N_VPWR_c_214_n 0.0108017f $X=1.895 $Y=1.765 $X2=0
+ $Y2=0
cc_110 N_A_27_368#_c_126_n N_VPWR_c_214_n 0.0227777f $X=2.125 $Y=2.405 $X2=0
+ $Y2=0
cc_111 N_A_27_368#_c_124_n N_VPWR_c_215_n 0.0097982f $X=0.27 $Y=2.695 $X2=0
+ $Y2=0
cc_112 N_A_27_368#_c_121_n N_VPWR_c_216_n 0.00413917f $X=1.425 $Y=1.765 $X2=0
+ $Y2=0
cc_113 N_A_27_368#_c_122_n N_VPWR_c_216_n 0.00413917f $X=1.895 $Y=1.765 $X2=0
+ $Y2=0
cc_114 N_A_27_368#_c_121_n N_VPWR_c_211_n 0.0041466f $X=1.425 $Y=1.765 $X2=0
+ $Y2=0
cc_115 N_A_27_368#_c_122_n N_VPWR_c_211_n 0.00414695f $X=1.895 $Y=1.765 $X2=0
+ $Y2=0
cc_116 N_A_27_368#_c_124_n N_VPWR_c_211_n 0.0111907f $X=0.27 $Y=2.695 $X2=0
+ $Y2=0
cc_117 N_A_27_368#_c_133_n N_VPWR_c_211_n 0.0203661f $X=1.215 $Y=2.405 $X2=0
+ $Y2=0
cc_118 N_A_27_368#_c_126_n N_VPWR_c_211_n 0.0194473f $X=2.125 $Y=2.405 $X2=0
+ $Y2=0
cc_119 N_A_27_368#_c_160_p N_VPWR_c_211_n 0.00118533f $X=1.3 $Y=2.405 $X2=0
+ $Y2=0
cc_120 N_A_27_368#_c_126_n N_X_M1000_d 0.00618549f $X=2.125 $Y=2.405 $X2=0 $Y2=0
cc_121 N_A_27_368#_M1003_g X 0.00175981f $X=1.425 $Y=0.74 $X2=0 $Y2=0
cc_122 N_A_27_368#_c_121_n X 5.71627e-19 $X=1.425 $Y=1.765 $X2=0 $Y2=0
cc_123 N_A_27_368#_M1007_g X 0.0173853f $X=1.855 $Y=0.74 $X2=0 $Y2=0
cc_124 N_A_27_368#_c_122_n X 5.83312e-19 $X=1.895 $Y=1.765 $X2=0 $Y2=0
cc_125 N_A_27_368#_c_115_n X 0.0099082f $X=1.215 $Y=1.095 $X2=0 $Y2=0
cc_126 N_A_27_368#_c_117_n X 0.0575862f $X=1.3 $Y=2.32 $X2=0 $Y2=0
cc_127 N_A_27_368#_c_118_n X 0.0092052f $X=2.21 $Y=2.32 $X2=0 $Y2=0
cc_128 N_A_27_368#_c_119_n X 0.0241749f $X=2.13 $Y=1.465 $X2=0 $Y2=0
cc_129 N_A_27_368#_c_120_n X 0.0266948f $X=1.895 $Y=1.532 $X2=0 $Y2=0
cc_130 N_A_27_368#_c_122_n X 0.00537402f $X=1.895 $Y=1.765 $X2=0 $Y2=0
cc_131 N_A_27_368#_c_126_n X 0.0177271f $X=2.125 $Y=2.405 $X2=0 $Y2=0
cc_132 N_A_27_368#_c_118_n X 0.0159957f $X=2.21 $Y=2.32 $X2=0 $Y2=0
cc_133 N_A_27_368#_c_120_n X 0.00119064f $X=1.895 $Y=1.532 $X2=0 $Y2=0
cc_134 N_A_27_368#_c_115_n N_VGND_M1006_d 0.00267951f $X=1.215 $Y=1.095 $X2=0
+ $Y2=0
cc_135 N_A_27_368#_c_114_n N_VGND_c_269_n 0.0204407f $X=0.705 $Y=0.615 $X2=0
+ $Y2=0
cc_136 N_A_27_368#_M1003_g N_VGND_c_270_n 0.0111891f $X=1.425 $Y=0.74 $X2=0
+ $Y2=0
cc_137 N_A_27_368#_M1007_g N_VGND_c_270_n 5.12656e-19 $X=1.855 $Y=0.74 $X2=0
+ $Y2=0
cc_138 N_A_27_368#_c_114_n N_VGND_c_270_n 0.0139492f $X=0.705 $Y=0.615 $X2=0
+ $Y2=0
cc_139 N_A_27_368#_c_115_n N_VGND_c_270_n 0.0208721f $X=1.215 $Y=1.095 $X2=0
+ $Y2=0
cc_140 N_A_27_368#_M1007_g N_VGND_c_272_n 0.0185053f $X=1.855 $Y=0.74 $X2=0
+ $Y2=0
cc_141 N_A_27_368#_c_119_n N_VGND_c_272_n 0.0281178f $X=2.13 $Y=1.465 $X2=0
+ $Y2=0
cc_142 N_A_27_368#_c_120_n N_VGND_c_272_n 0.00255588f $X=1.895 $Y=1.532 $X2=0
+ $Y2=0
cc_143 N_A_27_368#_c_114_n N_VGND_c_273_n 0.0078096f $X=0.705 $Y=0.615 $X2=0
+ $Y2=0
cc_144 N_A_27_368#_M1003_g N_VGND_c_274_n 0.00383152f $X=1.425 $Y=0.74 $X2=0
+ $Y2=0
cc_145 N_A_27_368#_M1007_g N_VGND_c_274_n 0.00445602f $X=1.855 $Y=0.74 $X2=0
+ $Y2=0
cc_146 N_A_27_368#_M1003_g N_VGND_c_276_n 0.0075754f $X=1.425 $Y=0.74 $X2=0
+ $Y2=0
cc_147 N_A_27_368#_M1007_g N_VGND_c_276_n 0.00860452f $X=1.855 $Y=0.74 $X2=0
+ $Y2=0
cc_148 N_A_27_368#_c_114_n N_VGND_c_276_n 0.0085649f $X=0.705 $Y=0.615 $X2=0
+ $Y2=0
cc_149 X N_VGND_c_270_n 0.0177481f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_150 X N_VGND_c_272_n 0.0287813f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_151 X N_VGND_c_274_n 0.0105779f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_152 X N_VGND_c_276_n 0.00872261f $X=1.595 $Y=0.47 $X2=0 $Y2=0
