* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hs__fahcon_1 A B CI VGND VNB VPB VPWR COUT_N SUM
X0 a_369_365# B a_27_100# VPB sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X1 a_27_100# A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X2 a_1023_389# a_374_120# COUT_N VPB sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X3 a_369_365# B a_241_368# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X4 COUT_N a_369_365# a_1261_421# VPB sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X5 a_241_368# a_336_263# a_374_120# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X6 a_1719_368# a_369_365# a_1744_94# VPB sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X7 VPWR CI a_1606_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X8 VGND B a_1023_389# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X9 a_1261_421# CI VGND VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X10 VPWR B a_1023_389# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=150000u
X11 a_27_100# a_336_263# a_369_365# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X12 a_27_100# A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X13 a_1744_94# a_374_120# a_1719_368# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X14 a_241_368# a_336_263# a_369_365# VPB sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X15 a_336_263# B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X16 a_336_263# B VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X17 a_1261_421# CI VPWR VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=150000u
X18 VPWR a_1744_94# SUM VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X19 a_1606_368# a_369_365# a_1744_94# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X20 a_27_100# a_336_263# a_374_120# VPB sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X21 a_1744_94# a_374_120# a_1606_368# VPB sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X22 VGND CI a_1606_368# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X23 VGND a_1744_94# SUM VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X24 VPWR a_27_100# a_241_368# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=150000u
X25 a_374_120# B a_241_368# VPB sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X26 a_1719_368# a_1606_368# VPWR VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=150000u
X27 a_1719_368# a_1606_368# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X28 VGND a_27_100# a_241_368# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X29 a_1023_389# a_369_365# COUT_N VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X30 a_374_120# B a_27_100# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X31 COUT_N a_374_120# a_1261_421# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
.ends
