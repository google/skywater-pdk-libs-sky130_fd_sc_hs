* File: sky130_fd_sc_hs__dfsbp_2.spice
* Created: Thu Aug 27 20:39:11 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hs__dfsbp_2.pex.spice"
.subckt sky130_fd_sc_hs__dfsbp_2  VNB VPB D CLK SET_B VPWR Q_N Q VGND
* 
* VGND	VGND
* Q	Q
* Q_N	Q_N
* VPWR	VPWR
* SET_B	SET_B
* CLK	CLK
* D	D
* VPB	VPB
* VNB	VNB
MM1031 N_VGND_M1031_d N_D_M1031_g N_A_27_74#_M1031_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.1197 AS=0.1197 PD=1.41 PS=1.41 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1033 N_VGND_M1033_d N_CLK_M1033_g N_A_225_74#_M1033_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.2109 PD=1.02 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1018 N_A_398_74#_M1018_d N_A_225_74#_M1018_g N_VGND_M1033_d VNB NLOWVT L=0.15
+ W=0.74 AD=0.2072 AS=0.1036 PD=2.04 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.6 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1017 N_A_595_97#_M1017_d N_A_225_74#_M1017_g N_A_27_74#_M1017_s VNB NLOWVT
+ L=0.15 W=0.42 AD=0.1113 AS=0.1197 PD=0.95 PS=1.41 NRD=71.424 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75001.2 A=0.063 P=1.14 MULT=1
MM1036 A_731_97# N_A_398_74#_M1036_g N_A_595_97#_M1017_d VNB NLOWVT L=0.15
+ W=0.42 AD=0.0441 AS=0.1113 PD=0.63 PS=0.95 NRD=14.28 NRS=0 M=1 R=2.8
+ SA=75000.9 SB=75000.6 A=0.063 P=1.14 MULT=1
MM1024 N_VGND_M1024_d N_A_757_401#_M1024_g A_731_97# VNB NLOWVT L=0.15 W=0.42
+ AD=0.1197 AS=0.0441 PD=1.41 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75001.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1029 A_1001_74# N_A_595_97#_M1029_g N_A_757_401#_M1029_s VNB NLOWVT L=0.15
+ W=0.42 AD=0.0441 AS=0.1197 PD=0.63 PS=1.41 NRD=14.28 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75003 A=0.063 P=1.14 MULT=1
MM1026 N_VGND_M1026_d N_SET_B_M1026_g A_1001_74# VNB NLOWVT L=0.15 W=0.42
+ AD=0.15326 AS=0.0441 PD=1.13321 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75000.6
+ SB=75002.7 A=0.063 P=1.14 MULT=1
MM1012 A_1261_74# N_A_595_97#_M1012_g N_VGND_M1026_d VNB NLOWVT L=0.15 W=0.64
+ AD=0.0768 AS=0.23354 PD=0.88 PS=1.72679 NRD=12.18 NRS=3.744 M=1 R=4.26667
+ SA=75001.1 SB=75002.2 A=0.096 P=1.58 MULT=1
MM1020 N_A_1339_74#_M1020_d N_A_398_74#_M1020_g A_1261_74# VNB NLOWVT L=0.15
+ W=0.64 AD=0.139713 AS=0.0768 PD=1.28 PS=0.88 NRD=13.116 NRS=12.18 M=1
+ R=4.26667 SA=75001.4 SB=75001.8 A=0.096 P=1.58 MULT=1
MM1037 A_1453_118# N_A_225_74#_M1037_g N_A_1339_74#_M1020_d VNB NLOWVT L=0.15
+ W=0.42 AD=0.0504 AS=0.0916868 PD=0.66 PS=0.84 NRD=18.564 NRS=19.992 M=1 R=2.8
+ SA=75001.8 SB=75002.1 A=0.063 P=1.14 MULT=1
MM1021 A_1531_118# N_A_1501_92#_M1021_g A_1453_118# VNB NLOWVT L=0.15 W=0.42
+ AD=0.0504 AS=0.0504 PD=0.66 PS=0.66 NRD=18.564 NRS=18.564 M=1 R=2.8 SA=75002.2
+ SB=75001.7 A=0.063 P=1.14 MULT=1
MM1002 N_VGND_M1002_d N_SET_B_M1002_g A_1531_118# VNB NLOWVT L=0.15 W=0.42
+ AD=0.260625 AS=0.0504 PD=1.505 PS=0.66 NRD=161.58 NRS=18.564 M=1 R=2.8
+ SA=75002.6 SB=75001.3 A=0.063 P=1.14 MULT=1
MM1003 N_A_1501_92#_M1003_d N_A_1339_74#_M1003_g N_VGND_M1002_d VNB NLOWVT
+ L=0.15 W=0.42 AD=0.1533 AS=0.260625 PD=1.57 PS=1.505 NRD=22.848 NRS=161.58 M=1
+ R=2.8 SA=75003.6 SB=75000.3 A=0.063 P=1.14 MULT=1
MM1013 N_Q_N_M1013_d N_A_1339_74#_M1013_g N_VGND_M1013_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.2109 PD=1.02 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75000.6 A=0.111 P=1.78 MULT=1
MM1022 N_Q_N_M1013_d N_A_1339_74#_M1022_g N_VGND_M1022_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.2109 PD=1.02 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.6 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1008 N_VGND_M1008_d N_A_1339_74#_M1008_g N_A_2221_74#_M1008_s VNB NLOWVT
+ L=0.15 W=0.64 AD=0.136255 AS=0.1824 PD=1.07594 PS=1.85 NRD=13.116 NRS=0 M=1
+ R=4.26667 SA=75000.2 SB=75001.2 A=0.096 P=1.58 MULT=1
MM1004 N_VGND_M1008_d N_A_2221_74#_M1004_g N_Q_M1004_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.157545 AS=0.1036 PD=1.24406 PS=1.02 NRD=11.34 NRS=0 M=1 R=4.93333
+ SA=75000.7 SB=75000.6 A=0.111 P=1.78 MULT=1
MM1016 N_VGND_M1016_d N_A_2221_74#_M1016_g N_Q_M1004_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.1036 PD=2.05 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.1
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1000 N_VPWR_M1000_d N_D_M1000_g N_A_27_74#_M1000_s VPB PSHORT L=0.15 W=0.42
+ AD=0.1239 AS=0.1239 PD=1.43 PS=1.43 NRD=4.6886 NRS=4.6886 M=1 R=2.8 SA=75000.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1027 N_VPWR_M1027_d N_CLK_M1027_g N_A_225_74#_M1027_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.3304 PD=1.42 PS=2.83 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1030 N_A_398_74#_M1030_d N_A_225_74#_M1030_g N_VPWR_M1027_d VPB PSHORT L=0.15
+ W=1.12 AD=0.3304 AS=0.168 PD=2.83 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.7 SB=75000.2 A=0.168 P=2.54 MULT=1
MM1011 N_A_595_97#_M1011_d N_A_398_74#_M1011_g N_A_27_74#_M1011_s VPB PSHORT
+ L=0.15 W=0.42 AD=0.063 AS=0.1239 PD=0.72 PS=1.43 NRD=4.6886 NRS=4.6886 M=1
+ R=2.8 SA=75000.2 SB=75004.5 A=0.063 P=1.14 MULT=1
MM1014 A_706_463# N_A_225_74#_M1014_g N_A_595_97#_M1011_d VPB PSHORT L=0.15
+ W=0.42 AD=0.0567 AS=0.063 PD=0.69 PS=0.72 NRD=37.5088 NRS=4.6886 M=1 R=2.8
+ SA=75000.7 SB=75004.1 A=0.063 P=1.14 MULT=1
MM1032 N_VPWR_M1032_d N_A_757_401#_M1032_g A_706_463# VPB PSHORT L=0.15 W=0.42
+ AD=0.1961 AS=0.0567 PD=1.425 PS=0.69 NRD=193.198 NRS=37.5088 M=1 R=2.8
+ SA=75001.1 SB=75003.6 A=0.063 P=1.14 MULT=1
MM1028 N_A_757_401#_M1028_d N_A_595_97#_M1028_g N_VPWR_M1032_d VPB PSHORT L=0.15
+ W=0.42 AD=0.07665 AS=0.1961 PD=0.785 PS=1.425 NRD=4.6886 NRS=193.198 M=1 R=2.8
+ SA=75002 SB=75002.7 A=0.063 P=1.14 MULT=1
MM1009 N_VPWR_M1009_d N_SET_B_M1009_g N_A_757_401#_M1028_d VPB PSHORT L=0.15
+ W=0.42 AD=0.150431 AS=0.07665 PD=1.11507 PS=0.785 NRD=168.849 NRS=35.1645 M=1
+ R=2.8 SA=75002.5 SB=75002.2 A=0.063 P=1.14 MULT=1
MM1015 A_1258_341# N_A_595_97#_M1015_g N_VPWR_M1009_d VPB PSHORT L=0.15 W=1
+ AD=0.199812 AS=0.358169 PD=1.61 PS=2.65493 NRD=28.5256 NRS=23.6203 M=1
+ R=6.66667 SA=75001.5 SB=75000.9 A=0.15 P=2.3 MULT=1
MM1035 N_A_1339_74#_M1035_d N_A_225_74#_M1035_g A_1258_341# VPB PSHORT L=0.15
+ W=1 AD=0.315704 AS=0.199812 PD=2.33803 PS=1.61 NRD=1.9503 NRS=28.5256 M=1
+ R=6.66667 SA=75001.8 SB=75000.9 A=0.15 P=2.3 MULT=1
MM1034 A_1521_508# N_A_398_74#_M1034_g N_A_1339_74#_M1035_d VPB PSHORT L=0.15
+ W=0.42 AD=0.0567 AS=0.132596 PD=0.69 PS=0.981972 NRD=37.5088 NRS=90.2851 M=1
+ R=2.8 SA=75002.5 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1006 N_VPWR_M1006_d N_A_1501_92#_M1006_g A_1521_508# VPB PSHORT L=0.15 W=0.42
+ AD=0.063 AS=0.0567 PD=0.72 PS=0.69 NRD=4.6886 NRS=37.5088 M=1 R=2.8 SA=75002.9
+ SB=75000.7 A=0.063 P=1.14 MULT=1
MM1007 N_A_1339_74#_M1007_d N_SET_B_M1007_g N_VPWR_M1006_d VPB PSHORT L=0.15
+ W=0.42 AD=0.1218 AS=0.063 PD=1.42 PS=0.72 NRD=4.6886 NRS=4.6886 M=1 R=2.8
+ SA=75003.3 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1010 N_VPWR_M1010_d N_A_1339_74#_M1010_g N_A_1501_92#_M1010_s VPB PSHORT
+ L=0.15 W=0.42 AD=0.100418 AS=0.2544 PD=0.820909 PS=2.27 NRD=86.3451
+ NRS=258.306 M=1 R=2.8 SA=75000.3 SB=75001.2 A=0.063 P=1.14 MULT=1
MM1001 N_VPWR_M1010_d N_A_1339_74#_M1001_g N_Q_N_M1001_s VPB PSHORT L=0.15
+ W=1.12 AD=0.267782 AS=0.168 PD=2.18909 PS=1.42 NRD=1.7533 NRS=1.7533 M=1
+ R=7.46667 SA=75000.5 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1019 N_VPWR_M1019_d N_A_1339_74#_M1019_g N_Q_N_M1001_s VPB PSHORT L=0.15
+ W=1.12 AD=0.3248 AS=0.168 PD=2.82 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.9 SB=75000.2 A=0.168 P=2.54 MULT=1
MM1005 N_VPWR_M1005_d N_A_1339_74#_M1005_g N_A_2221_74#_M1005_s VPB PSHORT
+ L=0.15 W=1 AD=0.19566 AS=0.295 PD=1.41509 PS=2.59 NRD=17.73 NRS=1.9503 M=1
+ R=6.66667 SA=75000.2 SB=75001.2 A=0.15 P=2.3 MULT=1
MM1023 N_Q_M1023_d N_A_2221_74#_M1023_g N_VPWR_M1005_d VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.21914 PD=1.42 PS=1.58491 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.7 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1025 N_Q_M1023_d N_A_2221_74#_M1025_g N_VPWR_M1025_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.3304 PD=1.42 PS=2.83 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.1 SB=75000.2 A=0.168 P=2.54 MULT=1
DX38_noxref VNB VPB NWDIODE A=25.1893 P=30.67
c_136 VNB 0 1.55885e-19 $X=0 $Y=0
*
.include "sky130_fd_sc_hs__dfsbp_2.pxi.spice"
*
.ends
*
*
