# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_hs__a311oi_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  10.08000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  1.116000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.635000 1.350000 6.115000 1.780000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  1.116000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.045000 1.350000 3.715000 1.780000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  1.116000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.525000 1.350000 1.875000 1.780000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.894000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.775000 1.180000 7.555000 1.320000 ;
        RECT 6.775000 1.320000 7.785000 1.650000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.894000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.065000 1.220000 9.075000 1.550000 ;
        RECT 8.285000 1.180000 9.075000 1.220000 ;
    END
  END C1
  PIN Y
    ANTENNADIFFAREA  1.700600 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.330000 0.770000 4.660000 0.850000 ;
        RECT 4.330000 0.850000 9.425000 1.010000 ;
        RECT 4.330000 1.010000 6.380000 1.130000 ;
        RECT 6.130000 0.350000 6.380000 0.840000 ;
        RECT 6.130000 0.840000 9.425000 0.850000 ;
        RECT 7.760000 0.350000 8.010000 0.840000 ;
        RECT 7.760000 1.010000 8.010000 1.050000 ;
        RECT 8.355000 1.720000 9.425000 1.890000 ;
        RECT 8.355000 1.890000 8.525000 2.735000 ;
        RECT 8.700000 0.350000 9.955000 0.670000 ;
        RECT 8.700000 0.670000 9.425000 0.840000 ;
        RECT 9.255000 1.010000 9.425000 1.720000 ;
        RECT 9.255000 1.890000 9.425000 2.735000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 10.080000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 10.080000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 10.080000 0.085000 ;
      RECT 0.000000  3.245000 10.080000 3.415000 ;
      RECT 0.105000  1.820000  0.355000 3.245000 ;
      RECT 0.150000  0.350000  0.400000 1.010000 ;
      RECT 0.150000  1.010000  3.920000 1.180000 ;
      RECT 0.555000  1.950000  7.655000 2.120000 ;
      RECT 0.555000  2.120000  0.805000 2.980000 ;
      RECT 0.580000  0.085000  0.830000 0.840000 ;
      RECT 1.005000  2.290000  1.335000 3.245000 ;
      RECT 1.010000  0.350000  1.260000 1.010000 ;
      RECT 1.440000  0.085000  1.770000 0.840000 ;
      RECT 1.535000  2.120000  1.705000 2.980000 ;
      RECT 1.905000  2.290000  2.235000 3.245000 ;
      RECT 1.950000  0.350000  2.120000 0.975000 ;
      RECT 1.950000  0.975000  3.920000 1.010000 ;
      RECT 2.300000  0.350000  5.950000 0.600000 ;
      RECT 2.300000  0.600000  2.560000 0.680000 ;
      RECT 2.435000  2.120000  2.605000 2.980000 ;
      RECT 2.730000  0.770000  3.060000 0.975000 ;
      RECT 2.805000  2.290000  3.135000 3.245000 ;
      RECT 3.230000  0.600000  3.420000 0.680000 ;
      RECT 3.335000  2.120000  3.505000 2.980000 ;
      RECT 3.590000  0.770000  3.920000 0.975000 ;
      RECT 3.705000  2.290000  4.035000 3.245000 ;
      RECT 4.235000  1.820000  4.405000 1.950000 ;
      RECT 4.235000  2.120000  4.405000 2.980000 ;
      RECT 4.605000  2.290000  4.855000 3.245000 ;
      RECT 5.055000  2.120000  5.305000 2.980000 ;
      RECT 5.505000  2.290000  5.835000 3.245000 ;
      RECT 5.620000  0.600000  5.950000 0.680000 ;
      RECT 6.025000  2.320000  6.355000 2.905000 ;
      RECT 6.025000  2.905000  9.955000 3.075000 ;
      RECT 6.475000  1.820000  7.655000 1.950000 ;
      RECT 6.475000  2.120000  7.655000 2.150000 ;
      RECT 6.525000  2.150000  6.755000 2.735000 ;
      RECT 6.550000  0.085000  7.590000 0.670000 ;
      RECT 6.925000  2.320000  7.255000 2.905000 ;
      RECT 7.425000  2.150000  7.655000 2.735000 ;
      RECT 7.825000  1.820000  8.155000 2.905000 ;
      RECT 8.190000  0.085000  8.520000 0.670000 ;
      RECT 8.725000  2.060000  9.055000 2.905000 ;
      RECT 9.625000  1.820000  9.955000 2.905000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
      RECT 7.835000 -0.085000 8.005000 0.085000 ;
      RECT 7.835000  3.245000 8.005000 3.415000 ;
      RECT 8.315000 -0.085000 8.485000 0.085000 ;
      RECT 8.315000  3.245000 8.485000 3.415000 ;
      RECT 8.795000 -0.085000 8.965000 0.085000 ;
      RECT 8.795000  3.245000 8.965000 3.415000 ;
      RECT 9.275000 -0.085000 9.445000 0.085000 ;
      RECT 9.275000  3.245000 9.445000 3.415000 ;
      RECT 9.755000 -0.085000 9.925000 0.085000 ;
      RECT 9.755000  3.245000 9.925000 3.415000 ;
  END
END sky130_fd_sc_hs__a311oi_4
