* File: sky130_fd_sc_hs__a2111oi_1.pxi.spice
* Created: Tue Sep  1 19:48:06 2020
* 
x_PM_SKY130_FD_SC_HS__A2111OI_1%D1 N_D1_c_54_n N_D1_M1000_g N_D1_M1004_g D1
+ N_D1_c_56_n PM_SKY130_FD_SC_HS__A2111OI_1%D1
x_PM_SKY130_FD_SC_HS__A2111OI_1%C1 N_C1_c_78_n N_C1_M1007_g N_C1_M1008_g C1
+ N_C1_c_80_n PM_SKY130_FD_SC_HS__A2111OI_1%C1
x_PM_SKY130_FD_SC_HS__A2111OI_1%B1 N_B1_c_110_n N_B1_M1001_g N_B1_M1009_g B1
+ N_B1_c_112_n PM_SKY130_FD_SC_HS__A2111OI_1%B1
x_PM_SKY130_FD_SC_HS__A2111OI_1%A1 N_A1_c_140_n N_A1_M1005_g N_A1_M1003_g A1
+ N_A1_c_142_n PM_SKY130_FD_SC_HS__A2111OI_1%A1
x_PM_SKY130_FD_SC_HS__A2111OI_1%A2 N_A2_c_171_n N_A2_M1002_g N_A2_c_172_n
+ N_A2_M1006_g A2 PM_SKY130_FD_SC_HS__A2111OI_1%A2
x_PM_SKY130_FD_SC_HS__A2111OI_1%Y N_Y_M1004_d N_Y_M1009_d N_Y_M1000_s
+ N_Y_c_196_n N_Y_c_197_n N_Y_c_198_n N_Y_c_199_n N_Y_c_200_n N_Y_c_201_n
+ N_Y_c_202_n Y Y Y PM_SKY130_FD_SC_HS__A2111OI_1%Y
x_PM_SKY130_FD_SC_HS__A2111OI_1%A_342_368# N_A_342_368#_M1001_d
+ N_A_342_368#_M1006_d N_A_342_368#_c_260_n N_A_342_368#_c_256_n
+ N_A_342_368#_c_264_n N_A_342_368#_c_257_n N_A_342_368#_c_258_n
+ PM_SKY130_FD_SC_HS__A2111OI_1%A_342_368#
x_PM_SKY130_FD_SC_HS__A2111OI_1%VPWR N_VPWR_M1005_d N_VPWR_c_284_n
+ N_VPWR_c_285_n N_VPWR_c_286_n VPWR N_VPWR_c_287_n N_VPWR_c_283_n
+ PM_SKY130_FD_SC_HS__A2111OI_1%VPWR
x_PM_SKY130_FD_SC_HS__A2111OI_1%VGND N_VGND_M1004_s N_VGND_M1008_d
+ N_VGND_M1002_d N_VGND_c_312_n N_VGND_c_313_n N_VGND_c_314_n N_VGND_c_315_n
+ N_VGND_c_316_n N_VGND_c_317_n N_VGND_c_318_n N_VGND_c_319_n N_VGND_c_320_n
+ N_VGND_c_321_n VGND N_VGND_c_322_n PM_SKY130_FD_SC_HS__A2111OI_1%VGND
cc_1 VNB N_D1_c_54_n 0.0266193f $X=-0.19 $Y=-0.245 $X2=0.705 $Y2=1.765
cc_2 VNB N_D1_M1004_g 0.0273265f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=0.74
cc_3 VNB N_D1_c_56_n 0.00391874f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.515
cc_4 VNB N_C1_c_78_n 0.0262279f $X=-0.19 $Y=-0.245 $X2=0.705 $Y2=1.765
cc_5 VNB N_C1_M1008_g 0.0266005f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=0.74
cc_6 VNB N_C1_c_80_n 0.00165719f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.515
cc_7 VNB N_B1_c_110_n 0.0262515f $X=-0.19 $Y=-0.245 $X2=0.705 $Y2=1.765
cc_8 VNB N_B1_M1009_g 0.026609f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=0.74
cc_9 VNB N_B1_c_112_n 0.00166777f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.515
cc_10 VNB N_A1_c_140_n 0.0242864f $X=-0.19 $Y=-0.245 $X2=0.705 $Y2=1.765
cc_11 VNB N_A1_M1003_g 0.0250188f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=0.74
cc_12 VNB N_A1_c_142_n 0.00709957f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.515
cc_13 VNB N_A2_c_171_n 0.0215297f $X=-0.19 $Y=-0.245 $X2=0.705 $Y2=1.765
cc_14 VNB N_A2_c_172_n 0.0431106f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.35
cc_15 VNB A2 0.0349068f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_Y_c_196_n 0.0230393f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.515
cc_17 VNB N_Y_c_197_n 0.0103726f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.515
cc_18 VNB N_Y_c_198_n 0.0149129f $X=-0.19 $Y=-0.245 $X2=0.65 $Y2=1.515
cc_19 VNB N_Y_c_199_n 0.00206666f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_Y_c_200_n 0.0170798f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_Y_c_201_n 0.00240191f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_Y_c_202_n 0.00677638f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_VPWR_c_283_n 0.143779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_VGND_c_312_n 0.0279165f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.515
cc_25 VNB N_VGND_c_313_n 0.00974487f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_VGND_c_314_n 0.0344702f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_VGND_c_315_n 0.0129628f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_316_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_317_n 0.0169342f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_318_n 0.00788625f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_319_n 0.0110534f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_320_n 0.0312656f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_321_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_322_n 0.227536f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VPB N_D1_c_54_n 0.0306918f $X=-0.19 $Y=1.66 $X2=0.705 $Y2=1.765
cc_36 VPB N_D1_c_56_n 0.00369353f $X=-0.19 $Y=1.66 $X2=0.63 $Y2=1.515
cc_37 VPB N_C1_c_78_n 0.0270094f $X=-0.19 $Y=1.66 $X2=0.705 $Y2=1.765
cc_38 VPB N_C1_c_80_n 0.00296952f $X=-0.19 $Y=1.66 $X2=0.63 $Y2=1.515
cc_39 VPB N_B1_c_110_n 0.0287122f $X=-0.19 $Y=1.66 $X2=0.705 $Y2=1.765
cc_40 VPB N_B1_c_112_n 0.00279327f $X=-0.19 $Y=1.66 $X2=0.63 $Y2=1.515
cc_41 VPB N_A1_c_140_n 0.0274332f $X=-0.19 $Y=1.66 $X2=0.705 $Y2=1.765
cc_42 VPB N_A1_c_142_n 0.0039015f $X=-0.19 $Y=1.66 $X2=0.63 $Y2=1.515
cc_43 VPB N_A2_c_172_n 0.0316663f $X=-0.19 $Y=1.66 $X2=0.72 $Y2=1.35
cc_44 VPB N_Y_c_196_n 0.0148281f $X=-0.19 $Y=1.66 $X2=0.63 $Y2=1.515
cc_45 VPB Y 0.0614439f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_46 VPB N_A_342_368#_c_256_n 0.00327016f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_47 VPB N_A_342_368#_c_257_n 0.0151999f $X=-0.19 $Y=1.66 $X2=0.65 $Y2=1.515
cc_48 VPB N_A_342_368#_c_258_n 0.0360166f $X=-0.19 $Y=1.66 $X2=0.65 $Y2=1.665
cc_49 VPB N_VPWR_c_284_n 0.00695663f $X=-0.19 $Y=1.66 $X2=0.72 $Y2=0.74
cc_50 VPB N_VPWR_c_285_n 0.0609497f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_51 VPB N_VPWR_c_286_n 0.00691066f $X=-0.19 $Y=1.66 $X2=0.63 $Y2=1.515
cc_52 VPB N_VPWR_c_287_n 0.0236066f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_53 VPB N_VPWR_c_283_n 0.0765274f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_54 N_D1_c_54_n N_C1_c_78_n 0.099031f $X=0.705 $Y=1.765 $X2=-0.19 $Y2=-0.245
cc_55 N_D1_c_56_n N_C1_c_78_n 0.00238234f $X=0.63 $Y=1.515 $X2=-0.19 $Y2=-0.245
cc_56 N_D1_M1004_g N_C1_M1008_g 0.0195038f $X=0.72 $Y=0.74 $X2=0 $Y2=0
cc_57 N_D1_c_54_n N_C1_c_80_n 5.23576e-19 $X=0.705 $Y=1.765 $X2=0 $Y2=0
cc_58 N_D1_c_56_n N_C1_c_80_n 0.0344038f $X=0.63 $Y=1.515 $X2=0 $Y2=0
cc_59 N_D1_c_54_n N_Y_c_196_n 0.0112102f $X=0.705 $Y=1.765 $X2=0 $Y2=0
cc_60 N_D1_M1004_g N_Y_c_196_n 0.00477786f $X=0.72 $Y=0.74 $X2=0 $Y2=0
cc_61 N_D1_c_56_n N_Y_c_196_n 0.0330212f $X=0.63 $Y=1.515 $X2=0 $Y2=0
cc_62 N_D1_c_54_n N_Y_c_197_n 0.00126003f $X=0.705 $Y=1.765 $X2=0 $Y2=0
cc_63 N_D1_M1004_g N_Y_c_197_n 0.0148724f $X=0.72 $Y=0.74 $X2=0 $Y2=0
cc_64 N_D1_c_56_n N_Y_c_197_n 0.0279704f $X=0.63 $Y=1.515 $X2=0 $Y2=0
cc_65 N_D1_M1004_g N_Y_c_199_n 3.97481e-19 $X=0.72 $Y=0.74 $X2=0 $Y2=0
cc_66 N_D1_c_54_n Y 0.0298656f $X=0.705 $Y=1.765 $X2=0 $Y2=0
cc_67 N_D1_c_56_n Y 0.0264648f $X=0.63 $Y=1.515 $X2=0 $Y2=0
cc_68 N_D1_c_54_n N_VPWR_c_285_n 0.00291649f $X=0.705 $Y=1.765 $X2=0 $Y2=0
cc_69 N_D1_c_54_n N_VPWR_c_283_n 0.00363021f $X=0.705 $Y=1.765 $X2=0 $Y2=0
cc_70 N_D1_M1004_g N_VGND_c_312_n 0.0127749f $X=0.72 $Y=0.74 $X2=0 $Y2=0
cc_71 N_D1_M1004_g N_VGND_c_317_n 0.00383152f $X=0.72 $Y=0.74 $X2=0 $Y2=0
cc_72 N_D1_M1004_g N_VGND_c_322_n 0.00757637f $X=0.72 $Y=0.74 $X2=0 $Y2=0
cc_73 N_C1_c_78_n N_B1_c_110_n 0.0602631f $X=1.095 $Y=1.765 $X2=-0.19 $Y2=-0.245
cc_74 N_C1_c_80_n N_B1_c_110_n 0.00179181f $X=1.17 $Y=1.515 $X2=-0.19 $Y2=-0.245
cc_75 N_C1_M1008_g N_B1_M1009_g 0.0204655f $X=1.15 $Y=0.74 $X2=0 $Y2=0
cc_76 N_C1_c_78_n N_B1_c_112_n 0.00127792f $X=1.095 $Y=1.765 $X2=0 $Y2=0
cc_77 N_C1_c_80_n N_B1_c_112_n 0.0277337f $X=1.17 $Y=1.515 $X2=0 $Y2=0
cc_78 N_C1_M1008_g N_Y_c_199_n 0.00959601f $X=1.15 $Y=0.74 $X2=0 $Y2=0
cc_79 N_C1_c_78_n N_Y_c_200_n 7.68393e-19 $X=1.095 $Y=1.765 $X2=0 $Y2=0
cc_80 N_C1_M1008_g N_Y_c_200_n 0.01209f $X=1.15 $Y=0.74 $X2=0 $Y2=0
cc_81 N_C1_c_80_n N_Y_c_200_n 0.0175347f $X=1.17 $Y=1.515 $X2=0 $Y2=0
cc_82 N_C1_M1008_g N_Y_c_201_n 8.21695e-19 $X=1.15 $Y=0.74 $X2=0 $Y2=0
cc_83 N_C1_c_78_n N_Y_c_202_n 5.40529e-19 $X=1.095 $Y=1.765 $X2=0 $Y2=0
cc_84 N_C1_M1008_g N_Y_c_202_n 0.0015571f $X=1.15 $Y=0.74 $X2=0 $Y2=0
cc_85 N_C1_c_80_n N_Y_c_202_n 0.00799991f $X=1.17 $Y=1.515 $X2=0 $Y2=0
cc_86 N_C1_c_78_n Y 0.0392015f $X=1.095 $Y=1.765 $X2=0 $Y2=0
cc_87 N_C1_c_80_n Y 0.023085f $X=1.17 $Y=1.515 $X2=0 $Y2=0
cc_88 N_C1_c_78_n N_A_342_368#_c_256_n 7.61918e-19 $X=1.095 $Y=1.765 $X2=0 $Y2=0
cc_89 N_C1_c_78_n N_VPWR_c_285_n 0.00291649f $X=1.095 $Y=1.765 $X2=0 $Y2=0
cc_90 N_C1_c_78_n N_VPWR_c_283_n 0.0035986f $X=1.095 $Y=1.765 $X2=0 $Y2=0
cc_91 N_C1_M1008_g N_VGND_c_312_n 5.17822e-19 $X=1.15 $Y=0.74 $X2=0 $Y2=0
cc_92 N_C1_M1008_g N_VGND_c_313_n 0.0053617f $X=1.15 $Y=0.74 $X2=0 $Y2=0
cc_93 N_C1_M1008_g N_VGND_c_317_n 0.00434272f $X=1.15 $Y=0.74 $X2=0 $Y2=0
cc_94 N_C1_M1008_g N_VGND_c_322_n 0.00821949f $X=1.15 $Y=0.74 $X2=0 $Y2=0
cc_95 N_B1_c_110_n N_A1_c_140_n 0.043721f $X=1.635 $Y=1.765 $X2=-0.19 $Y2=-0.245
cc_96 N_B1_c_112_n N_A1_c_140_n 7.18891e-19 $X=1.71 $Y=1.515 $X2=-0.19
+ $Y2=-0.245
cc_97 N_B1_M1009_g N_A1_M1003_g 0.0204481f $X=1.8 $Y=0.74 $X2=0 $Y2=0
cc_98 N_B1_c_110_n N_A1_c_142_n 0.00214941f $X=1.635 $Y=1.765 $X2=0 $Y2=0
cc_99 N_B1_c_112_n N_A1_c_142_n 0.0347535f $X=1.71 $Y=1.515 $X2=0 $Y2=0
cc_100 N_B1_M1009_g N_Y_c_199_n 8.24465e-19 $X=1.8 $Y=0.74 $X2=0 $Y2=0
cc_101 N_B1_c_110_n N_Y_c_200_n 0.00124693f $X=1.635 $Y=1.765 $X2=0 $Y2=0
cc_102 N_B1_M1009_g N_Y_c_200_n 0.0136326f $X=1.8 $Y=0.74 $X2=0 $Y2=0
cc_103 N_B1_c_112_n N_Y_c_200_n 0.0248933f $X=1.71 $Y=1.515 $X2=0 $Y2=0
cc_104 N_B1_M1009_g N_Y_c_201_n 0.00990712f $X=1.8 $Y=0.74 $X2=0 $Y2=0
cc_105 N_B1_c_110_n Y 0.00958302f $X=1.635 $Y=1.765 $X2=0 $Y2=0
cc_106 N_B1_c_110_n N_A_342_368#_c_260_n 0.00344123f $X=1.635 $Y=1.765 $X2=0
+ $Y2=0
cc_107 N_B1_c_112_n N_A_342_368#_c_260_n 0.0131798f $X=1.71 $Y=1.515 $X2=0 $Y2=0
cc_108 N_B1_c_110_n N_A_342_368#_c_256_n 0.0128632f $X=1.635 $Y=1.765 $X2=0
+ $Y2=0
cc_109 N_B1_c_110_n N_VPWR_c_284_n 6.63234e-19 $X=1.635 $Y=1.765 $X2=0 $Y2=0
cc_110 N_B1_c_110_n N_VPWR_c_285_n 0.00445602f $X=1.635 $Y=1.765 $X2=0 $Y2=0
cc_111 N_B1_c_110_n N_VPWR_c_283_n 0.00860014f $X=1.635 $Y=1.765 $X2=0 $Y2=0
cc_112 N_B1_M1009_g N_VGND_c_313_n 0.00690689f $X=1.8 $Y=0.74 $X2=0 $Y2=0
cc_113 N_B1_M1009_g N_VGND_c_320_n 0.00434272f $X=1.8 $Y=0.74 $X2=0 $Y2=0
cc_114 N_B1_M1009_g N_VGND_c_322_n 0.00821949f $X=1.8 $Y=0.74 $X2=0 $Y2=0
cc_115 N_A1_M1003_g N_A2_c_171_n 0.039902f $X=2.23 $Y=0.74 $X2=-0.19 $Y2=-0.245
cc_116 N_A1_c_140_n N_A2_c_172_n 0.0488455f $X=2.175 $Y=1.765 $X2=0 $Y2=0
cc_117 N_A1_c_142_n N_A2_c_172_n 0.00351611f $X=2.25 $Y=1.515 $X2=0 $Y2=0
cc_118 N_A1_c_140_n A2 6.92182e-19 $X=2.175 $Y=1.765 $X2=0 $Y2=0
cc_119 N_A1_M1003_g A2 0.00101508f $X=2.23 $Y=0.74 $X2=0 $Y2=0
cc_120 N_A1_c_142_n A2 0.013398f $X=2.25 $Y=1.515 $X2=0 $Y2=0
cc_121 N_A1_c_140_n N_Y_c_200_n 5.48416e-19 $X=2.175 $Y=1.765 $X2=0 $Y2=0
cc_122 N_A1_M1003_g N_Y_c_200_n 0.00464229f $X=2.23 $Y=0.74 $X2=0 $Y2=0
cc_123 N_A1_c_142_n N_Y_c_200_n 0.0116188f $X=2.25 $Y=1.515 $X2=0 $Y2=0
cc_124 N_A1_M1003_g N_Y_c_201_n 0.0132273f $X=2.23 $Y=0.74 $X2=0 $Y2=0
cc_125 N_A1_c_140_n N_A_342_368#_c_256_n 0.00507867f $X=2.175 $Y=1.765 $X2=0
+ $Y2=0
cc_126 N_A1_c_140_n N_A_342_368#_c_264_n 0.0164123f $X=2.175 $Y=1.765 $X2=0
+ $Y2=0
cc_127 N_A1_c_142_n N_A_342_368#_c_264_n 0.0235693f $X=2.25 $Y=1.515 $X2=0 $Y2=0
cc_128 N_A1_c_140_n N_A_342_368#_c_257_n 5.93323e-19 $X=2.175 $Y=1.765 $X2=0
+ $Y2=0
cc_129 N_A1_c_140_n N_A_342_368#_c_258_n 7.54205e-19 $X=2.175 $Y=1.765 $X2=0
+ $Y2=0
cc_130 N_A1_c_140_n N_VPWR_c_284_n 0.0111932f $X=2.175 $Y=1.765 $X2=0 $Y2=0
cc_131 N_A1_c_140_n N_VPWR_c_285_n 0.00413917f $X=2.175 $Y=1.765 $X2=0 $Y2=0
cc_132 N_A1_c_140_n N_VPWR_c_283_n 0.00818558f $X=2.175 $Y=1.765 $X2=0 $Y2=0
cc_133 N_A1_M1003_g N_VGND_c_314_n 0.00253715f $X=2.23 $Y=0.74 $X2=0 $Y2=0
cc_134 N_A1_M1003_g N_VGND_c_320_n 0.00434272f $X=2.23 $Y=0.74 $X2=0 $Y2=0
cc_135 N_A1_M1003_g N_VGND_c_322_n 0.00821825f $X=2.23 $Y=0.74 $X2=0 $Y2=0
cc_136 N_A2_c_171_n N_Y_c_200_n 8.07707e-19 $X=2.7 $Y=1.22 $X2=0 $Y2=0
cc_137 N_A2_c_171_n N_Y_c_201_n 0.0019967f $X=2.7 $Y=1.22 $X2=0 $Y2=0
cc_138 N_A2_c_172_n N_A_342_368#_c_264_n 0.0135061f $X=2.715 $Y=1.765 $X2=0
+ $Y2=0
cc_139 A2 N_A_342_368#_c_264_n 0.00515375f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_140 N_A2_c_172_n N_A_342_368#_c_257_n 0.0071736f $X=2.715 $Y=1.765 $X2=0
+ $Y2=0
cc_141 A2 N_A_342_368#_c_257_n 0.0204504f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_142 N_A2_c_172_n N_A_342_368#_c_258_n 0.0114033f $X=2.715 $Y=1.765 $X2=0
+ $Y2=0
cc_143 N_A2_c_172_n N_VPWR_c_284_n 0.00734374f $X=2.715 $Y=1.765 $X2=0 $Y2=0
cc_144 N_A2_c_172_n N_VPWR_c_287_n 0.00445602f $X=2.715 $Y=1.765 $X2=0 $Y2=0
cc_145 N_A2_c_172_n N_VPWR_c_283_n 0.00861623f $X=2.715 $Y=1.765 $X2=0 $Y2=0
cc_146 N_A2_c_171_n N_VGND_c_314_n 0.0176088f $X=2.7 $Y=1.22 $X2=0 $Y2=0
cc_147 N_A2_c_172_n N_VGND_c_314_n 0.00111834f $X=2.715 $Y=1.765 $X2=0 $Y2=0
cc_148 A2 N_VGND_c_314_n 0.0259407f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_149 N_A2_c_171_n N_VGND_c_320_n 0.00383152f $X=2.7 $Y=1.22 $X2=0 $Y2=0
cc_150 N_A2_c_171_n N_VGND_c_322_n 0.00757998f $X=2.7 $Y=1.22 $X2=0 $Y2=0
cc_151 Y A_156_368# 0.00568393f $X=1.115 $Y=2.32 $X2=-0.19 $Y2=-0.245
cc_152 Y A_234_368# 0.013495f $X=1.115 $Y=2.32 $X2=-0.19 $Y2=-0.245
cc_153 Y N_A_342_368#_c_260_n 0.00791971f $X=1.115 $Y=2.32 $X2=0 $Y2=0
cc_154 Y N_A_342_368#_c_256_n 0.0385009f $X=1.115 $Y=2.32 $X2=0 $Y2=0
cc_155 Y N_VPWR_c_285_n 0.0519698f $X=1.115 $Y=2.32 $X2=0 $Y2=0
cc_156 Y N_VPWR_c_283_n 0.0424701f $X=1.115 $Y=2.32 $X2=0 $Y2=0
cc_157 N_Y_c_197_n N_VGND_M1004_s 0.00267685f $X=0.85 $Y=1.095 $X2=-0.19
+ $Y2=-0.245
cc_158 N_Y_c_200_n N_VGND_M1008_d 0.00487041f $X=1.85 $Y=1.095 $X2=0 $Y2=0
cc_159 N_Y_c_197_n N_VGND_c_312_n 0.0220026f $X=0.85 $Y=1.095 $X2=0 $Y2=0
cc_160 N_Y_c_199_n N_VGND_c_312_n 0.0182902f $X=0.935 $Y=0.515 $X2=0 $Y2=0
cc_161 N_Y_c_199_n N_VGND_c_313_n 0.018437f $X=0.935 $Y=0.515 $X2=0 $Y2=0
cc_162 N_Y_c_200_n N_VGND_c_313_n 0.0314044f $X=1.85 $Y=1.095 $X2=0 $Y2=0
cc_163 N_Y_c_201_n N_VGND_c_313_n 0.0192028f $X=2.015 $Y=0.515 $X2=0 $Y2=0
cc_164 N_Y_c_201_n N_VGND_c_314_n 0.018269f $X=2.015 $Y=0.515 $X2=0 $Y2=0
cc_165 N_Y_c_199_n N_VGND_c_317_n 0.0109942f $X=0.935 $Y=0.515 $X2=0 $Y2=0
cc_166 N_Y_c_201_n N_VGND_c_320_n 0.0144922f $X=2.015 $Y=0.515 $X2=0 $Y2=0
cc_167 N_Y_c_199_n N_VGND_c_322_n 0.00904371f $X=0.935 $Y=0.515 $X2=0 $Y2=0
cc_168 N_Y_c_201_n N_VGND_c_322_n 0.0118826f $X=2.015 $Y=0.515 $X2=0 $Y2=0
cc_169 N_A_342_368#_c_264_n N_VPWR_M1005_d 0.010589f $X=2.775 $Y=2.035 $X2=-0.19
+ $Y2=1.66
cc_170 N_A_342_368#_c_256_n N_VPWR_c_284_n 0.0271521f $X=1.88 $Y=2.435 $X2=0
+ $Y2=0
cc_171 N_A_342_368#_c_264_n N_VPWR_c_284_n 0.0234793f $X=2.775 $Y=2.035 $X2=0
+ $Y2=0
cc_172 N_A_342_368#_c_258_n N_VPWR_c_284_n 0.0266947f $X=2.94 $Y=2.815 $X2=0
+ $Y2=0
cc_173 N_A_342_368#_c_256_n N_VPWR_c_285_n 0.0163786f $X=1.88 $Y=2.435 $X2=0
+ $Y2=0
cc_174 N_A_342_368#_c_258_n N_VPWR_c_287_n 0.0145938f $X=2.94 $Y=2.815 $X2=0
+ $Y2=0
cc_175 N_A_342_368#_c_256_n N_VPWR_c_283_n 0.0135239f $X=1.88 $Y=2.435 $X2=0
+ $Y2=0
cc_176 N_A_342_368#_c_258_n N_VPWR_c_283_n 0.0120466f $X=2.94 $Y=2.815 $X2=0
+ $Y2=0
