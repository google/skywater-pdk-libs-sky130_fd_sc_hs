# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_hs__mux2i_4
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_hs__mux2i_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  10.08000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A0
    ANTENNAGATEAREA  1.116000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.225000 1.350000 3.235000 1.680000 ;
        RECT 2.525000 1.680000 3.235000 1.780000 ;
    END
  END A0
  PIN A1
    ANTENNAGATEAREA  1.116000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.535000 1.350000 1.885000 1.780000 ;
    END
  END A1
  PIN S
    ANTENNAGATEAREA  1.479000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.080000 1.180000 9.475000 1.540000 ;
    END
  END S
  PIN Y
    ANTENNADIFFAREA  2.868700 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.115000 0.405000 0.365000 1.010000 ;
        RECT 0.115000 1.010000 4.085000 1.180000 ;
        RECT 0.115000 1.180000 0.365000 1.185000 ;
        RECT 0.115000 1.820000 0.365000 1.950000 ;
        RECT 0.115000 1.950000 4.245000 2.120000 ;
        RECT 0.115000 2.120000 0.365000 2.980000 ;
        RECT 1.055000 0.595000 1.225000 1.010000 ;
        RECT 1.095000 2.120000 1.265000 2.735000 ;
        RECT 1.915000 2.120000 2.245000 2.735000 ;
        RECT 1.920000 0.595000 2.250000 0.935000 ;
        RECT 1.920000 0.935000 4.085000 1.010000 ;
        RECT 2.915000 2.120000 3.245000 2.395000 ;
        RECT 3.485000 1.550000 4.245000 1.950000 ;
        RECT 3.915000 1.180000 4.085000 1.550000 ;
        RECT 3.915000 2.120000 4.245000 2.395000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 10.080000 0.085000 ;
        RECT 4.935000  0.085000  5.185000 0.490000 ;
        RECT 5.875000  0.085000  6.205000 0.410000 ;
        RECT 6.895000  0.085000  7.225000 0.410000 ;
        RECT 7.905000  0.085000  8.325000 0.640000 ;
        RECT 8.995000  0.085000  9.325000 1.010000 ;
      LAYER mcon ;
        RECT 0.155000 -0.085000 0.325000 0.085000 ;
        RECT 0.635000 -0.085000 0.805000 0.085000 ;
        RECT 1.115000 -0.085000 1.285000 0.085000 ;
        RECT 1.595000 -0.085000 1.765000 0.085000 ;
        RECT 2.075000 -0.085000 2.245000 0.085000 ;
        RECT 2.555000 -0.085000 2.725000 0.085000 ;
        RECT 3.035000 -0.085000 3.205000 0.085000 ;
        RECT 3.515000 -0.085000 3.685000 0.085000 ;
        RECT 3.995000 -0.085000 4.165000 0.085000 ;
        RECT 4.475000 -0.085000 4.645000 0.085000 ;
        RECT 4.955000 -0.085000 5.125000 0.085000 ;
        RECT 5.435000 -0.085000 5.605000 0.085000 ;
        RECT 5.915000 -0.085000 6.085000 0.085000 ;
        RECT 6.395000 -0.085000 6.565000 0.085000 ;
        RECT 6.875000 -0.085000 7.045000 0.085000 ;
        RECT 7.355000 -0.085000 7.525000 0.085000 ;
        RECT 7.835000 -0.085000 8.005000 0.085000 ;
        RECT 8.315000 -0.085000 8.485000 0.085000 ;
        RECT 8.795000 -0.085000 8.965000 0.085000 ;
        RECT 9.275000 -0.085000 9.445000 0.085000 ;
        RECT 9.755000 -0.085000 9.925000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.245000 10.080000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 3.245000 10.080000 3.415000 ;
        RECT 4.475000 1.840000  6.080000 2.050000 ;
        RECT 4.475000 2.050000  9.010000 2.220000 ;
        RECT 6.730000 2.730000  7.060000 3.245000 ;
        RECT 7.730000 2.730000  8.060000 3.245000 ;
        RECT 8.760000 2.220000  9.010000 3.245000 ;
        RECT 9.635000 2.050000  9.965000 3.245000 ;
      LAYER mcon ;
        RECT 0.155000 3.245000 0.325000 3.415000 ;
        RECT 0.635000 3.245000 0.805000 3.415000 ;
        RECT 1.115000 3.245000 1.285000 3.415000 ;
        RECT 1.595000 3.245000 1.765000 3.415000 ;
        RECT 2.075000 3.245000 2.245000 3.415000 ;
        RECT 2.555000 3.245000 2.725000 3.415000 ;
        RECT 3.035000 3.245000 3.205000 3.415000 ;
        RECT 3.515000 3.245000 3.685000 3.415000 ;
        RECT 3.995000 3.245000 4.165000 3.415000 ;
        RECT 4.475000 3.245000 4.645000 3.415000 ;
        RECT 4.955000 3.245000 5.125000 3.415000 ;
        RECT 5.435000 3.245000 5.605000 3.415000 ;
        RECT 5.915000 3.245000 6.085000 3.415000 ;
        RECT 6.395000 3.245000 6.565000 3.415000 ;
        RECT 6.875000 3.245000 7.045000 3.415000 ;
        RECT 7.355000 3.245000 7.525000 3.415000 ;
        RECT 7.835000 3.245000 8.005000 3.415000 ;
        RECT 8.315000 3.245000 8.485000 3.415000 ;
        RECT 8.795000 3.245000 8.965000 3.415000 ;
        RECT 9.275000 3.245000 9.445000 3.415000 ;
        RECT 9.755000 3.245000 9.925000 3.415000 ;
      LAYER met1 ;
        RECT 0.000000 3.085000 10.080000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.545000 0.255000 4.765000 0.425000 ;
      RECT 0.545000 0.425000 0.875000 0.840000 ;
      RECT 0.565000 2.290000 0.895000 2.905000 ;
      RECT 0.565000 2.905000 6.560000 3.075000 ;
      RECT 1.405000 0.425000 1.735000 0.840000 ;
      RECT 1.465000 2.290000 1.715000 2.905000 ;
      RECT 2.415000 2.290000 2.745000 2.565000 ;
      RECT 2.415000 2.565000 5.130000 2.735000 ;
      RECT 2.420000 0.595000 4.425000 0.765000 ;
      RECT 3.415000 2.290000 3.745000 2.565000 ;
      RECT 4.255000 0.765000 4.425000 1.000000 ;
      RECT 4.255000 1.000000 6.715000 1.170000 ;
      RECT 4.595000 0.425000 4.765000 0.660000 ;
      RECT 4.595000 0.660000 7.735000 0.750000 ;
      RECT 4.595000 0.750000 5.525000 0.830000 ;
      RECT 4.960000 2.390000 8.560000 2.560000 ;
      RECT 4.960000 2.560000 5.130000 2.565000 ;
      RECT 5.150000 1.340000 6.840000 1.670000 ;
      RECT 5.300000 2.730000 6.560000 2.905000 ;
      RECT 5.355000 0.580000 7.735000 0.660000 ;
      RECT 6.385000 0.920000 6.715000 1.000000 ;
      RECT 6.670000 1.670000 6.840000 1.710000 ;
      RECT 6.670000 1.710000 9.825000 1.880000 ;
      RECT 7.230000 2.560000 7.560000 2.980000 ;
      RECT 7.405000 0.390000 7.735000 0.580000 ;
      RECT 7.405000 0.750000 7.735000 0.840000 ;
      RECT 7.405000 0.840000 8.825000 1.010000 ;
      RECT 8.230000 2.560000 8.560000 2.980000 ;
      RECT 8.495000 0.390000 8.825000 0.840000 ;
      RECT 9.185000 1.880000 9.455000 2.700000 ;
      RECT 9.495000 0.390000 9.825000 1.010000 ;
      RECT 9.655000 1.010000 9.825000 1.710000 ;
  END
END sky130_fd_sc_hs__mux2i_4
