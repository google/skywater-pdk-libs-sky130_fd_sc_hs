* File: sky130_fd_sc_hs__buf_1.pex.spice
* Created: Thu Aug 27 20:34:19 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HS__BUF_1%A 3 5 7 9 10 11
c34 5 0 8.14418e-20 $X=0.86 $Y=2.045
c35 3 0 1.25263e-20 $X=0.845 $Y=0.835
r36 11 15 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.745
+ $Y=1.615 $X2=0.745 $Y2=1.615
r37 10 11 16.7628 $w=3.28e-07 $l=4.8e-07 $layer=LI1_cond $X=0.24 $Y=1.615
+ $X2=0.72 $Y2=1.615
r38 9 15 4.37153 $w=3.3e-07 $l=2.5e-08 $layer=POLY_cond $X=0.77 $Y=1.615
+ $X2=0.745 $Y2=1.615
r39 5 9 131.349 $w=1.58e-07 $l=4.3e-07 $layer=POLY_cond $X=0.86 $Y=2.045
+ $X2=0.86 $Y2=1.615
r40 5 7 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=0.86 $Y=2.045 $X2=0.86
+ $Y2=2.54
r41 1 9 50.5074 $w=1.58e-07 $l=1.72337e-07 $layer=POLY_cond $X=0.845 $Y=1.45
+ $X2=0.86 $Y2=1.615
r42 1 3 315.351 $w=1.5e-07 $l=6.15e-07 $layer=POLY_cond $X=0.845 $Y=1.45
+ $X2=0.845 $Y2=0.835
.ends

.subckt PM_SKY130_FD_SC_HS__BUF_1%A_27_164# 1 2 7 9 12 16 18 20 21 22 23 29
c58 7 0 8.84994e-20 $X=1.41 $Y=1.765
r59 32 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.325
+ $Y=1.465 $X2=1.325 $Y2=1.465
r60 28 29 9.39634 $w=4.78e-07 $l=1.65e-07 $layer=LI1_cond $X=0.63 $Y=1.04
+ $X2=0.795 $Y2=1.04
r61 25 28 8.72141 $w=4.78e-07 $l=3.5e-07 $layer=LI1_cond $X=0.28 $Y=1.04
+ $X2=0.63 $Y2=1.04
r62 22 32 9.01297 $w=2.9e-07 $l=2.07123e-07 $layer=LI1_cond $X=1.215 $Y=1.63
+ $X2=1.31 $Y2=1.465
r63 22 23 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=1.215 $Y=1.63
+ $X2=1.215 $Y2=1.95
r64 20 23 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.13 $Y=2.035
+ $X2=1.215 $Y2=1.95
r65 20 21 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=1.13 $Y=2.035
+ $X2=0.8 $Y2=2.035
r66 18 32 11.3586 $w=2.9e-07 $l=3.48569e-07 $layer=LI1_cond $X=1.13 $Y=1.195
+ $X2=1.31 $Y2=1.465
r67 18 29 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=1.13 $Y=1.195
+ $X2=0.795 $Y2=1.195
r68 14 21 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.635 $Y=2.12
+ $X2=0.8 $Y2=2.035
r69 14 16 5.06376 $w=3.28e-07 $l=1.45e-07 $layer=LI1_cond $X=0.635 $Y=2.12
+ $X2=0.635 $Y2=2.265
r70 10 33 38.5916 $w=2.93e-07 $l=2.07123e-07 $layer=POLY_cond $X=1.425 $Y=1.3
+ $X2=1.33 $Y2=1.465
r71 10 12 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=1.425 $Y=1.3
+ $X2=1.425 $Y2=0.74
r72 7 33 60.7998 $w=2.93e-07 $l=3.37639e-07 $layer=POLY_cond $X=1.41 $Y=1.765
+ $X2=1.33 $Y2=1.465
r73 7 9 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.41 $Y=1.765
+ $X2=1.41 $Y2=2.4
r74 2 16 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=0.49
+ $Y=2.12 $X2=0.635 $Y2=2.265
r75 1 28 182 $w=1.7e-07 $l=5.6285e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.82 $X2=0.63 $Y2=0.965
r76 1 25 182 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.82 $X2=0.28 $Y2=0.965
.ends

.subckt PM_SKY130_FD_SC_HS__BUF_1%VPWR 1 6 8 10 17 18 21
r21 21 22 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r22 18 22 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r23 17 18 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r24 15 21 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.3 $Y=3.33
+ $X2=1.135 $Y2=3.33
r25 15 17 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=1.3 $Y=3.33 $X2=1.68
+ $Y2=3.33
r26 12 13 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r27 10 21 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.97 $Y=3.33
+ $X2=1.135 $Y2=3.33
r28 10 12 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=0.97 $Y=3.33
+ $X2=0.72 $Y2=3.33
r29 8 22 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=0.96 $Y=3.33
+ $X2=1.2 $Y2=3.33
r30 8 13 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=0.96 $Y=3.33
+ $X2=0.72 $Y2=3.33
r31 4 21 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.135 $Y=3.245
+ $X2=1.135 $Y2=3.33
r32 4 6 27.5888 $w=3.28e-07 $l=7.9e-07 $layer=LI1_cond $X=1.135 $Y=3.245
+ $X2=1.135 $Y2=2.455
r33 1 6 300 $w=1.7e-07 $l=4.2335e-07 $layer=licon1_PDIFF $count=2 $X=0.935
+ $Y=2.12 $X2=1.135 $Y2=2.455
.ends

.subckt PM_SKY130_FD_SC_HS__BUF_1%X 1 2 9 13 14 15 16 23 32
c25 32 0 8.84994e-20 $X=1.65 $Y=1.82
c26 14 0 8.14418e-20 $X=1.595 $Y=1.95
c27 13 0 1.25263e-20 $X=1.652 $Y=1.13
r28 21 23 1.12043 $w=3.58e-07 $l=3.5e-08 $layer=LI1_cond $X=1.65 $Y=2 $X2=1.65
+ $Y2=2.035
r29 15 16 11.8446 $w=3.58e-07 $l=3.7e-07 $layer=LI1_cond $X=1.65 $Y=2.405
+ $X2=1.65 $Y2=2.775
r30 14 21 0.800308 $w=3.58e-07 $l=2.5e-08 $layer=LI1_cond $X=1.65 $Y=1.975
+ $X2=1.65 $Y2=2
r31 14 32 8.1909 $w=3.58e-07 $l=1.55e-07 $layer=LI1_cond $X=1.65 $Y=1.975
+ $X2=1.65 $Y2=1.82
r32 14 15 11.0442 $w=3.58e-07 $l=3.45e-07 $layer=LI1_cond $X=1.65 $Y=2.06
+ $X2=1.65 $Y2=2.405
r33 14 23 0.800308 $w=3.58e-07 $l=2.5e-08 $layer=LI1_cond $X=1.65 $Y=2.06
+ $X2=1.65 $Y2=2.035
r34 13 32 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.745 $Y=1.13
+ $X2=1.745 $Y2=1.82
r35 7 13 8.88861 $w=3.53e-07 $l=1.77e-07 $layer=LI1_cond $X=1.652 $Y=0.953
+ $X2=1.652 $Y2=1.13
r36 7 9 14.2189 $w=3.53e-07 $l=4.38e-07 $layer=LI1_cond $X=1.652 $Y=0.953
+ $X2=1.652 $Y2=0.515
r37 2 14 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=1.485
+ $Y=1.84 $X2=1.635 $Y2=1.985
r38 2 16 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=1.485
+ $Y=1.84 $X2=1.635 $Y2=2.815
r39 1 9 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.5 $Y=0.37
+ $X2=1.64 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__BUF_1%VGND 1 6 8 10 17 18 21
r19 21 22 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r20 18 22 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r21 17 18 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r22 15 21 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.305 $Y=0 $X2=1.14
+ $Y2=0
r23 15 17 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=1.305 $Y=0 $X2=1.68
+ $Y2=0
r24 12 13 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r25 10 21 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.975 $Y=0 $X2=1.14
+ $Y2=0
r26 10 12 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.975 $Y=0 $X2=0.72
+ $Y2=0
r27 8 22 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=0.96 $Y=0 $X2=1.2
+ $Y2=0
r28 8 13 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=0.96 $Y=0 $X2=0.72
+ $Y2=0
r29 4 21 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.14 $Y=0.085 $X2=1.14
+ $Y2=0
r30 4 6 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=1.14 $Y=0.085 $X2=1.14
+ $Y2=0.515
r31 1 6 91 $w=1.7e-07 $l=2.41454e-07 $layer=licon1_NDIFF $count=2 $X=0.92
+ $Y=0.56 $X2=1.14 $Y2=0.515
.ends

