* File: sky130_fd_sc_hs__clkinv_1.pxi.spice
* Created: Thu Aug 27 20:36:57 2020
* 
x_PM_SKY130_FD_SC_HS__CLKINV_1%A N_A_c_31_n N_A_M1000_g N_A_M1002_g N_A_c_32_n
+ N_A_M1001_g A A N_A_c_28_n N_A_c_29_n N_A_c_30_n
+ PM_SKY130_FD_SC_HS__CLKINV_1%A
x_PM_SKY130_FD_SC_HS__CLKINV_1%VPWR N_VPWR_M1000_d N_VPWR_M1001_d N_VPWR_c_61_n
+ N_VPWR_c_62_n N_VPWR_c_63_n N_VPWR_c_64_n VPWR N_VPWR_c_65_n N_VPWR_c_60_n
+ PM_SKY130_FD_SC_HS__CLKINV_1%VPWR
x_PM_SKY130_FD_SC_HS__CLKINV_1%Y N_Y_M1002_d N_Y_M1000_s N_Y_c_86_n N_Y_c_81_n Y
+ Y Y Y Y N_Y_c_83_n Y N_Y_c_85_n PM_SKY130_FD_SC_HS__CLKINV_1%Y
x_PM_SKY130_FD_SC_HS__CLKINV_1%VGND N_VGND_M1002_s N_VGND_c_109_n N_VGND_c_110_n
+ VGND N_VGND_c_111_n N_VGND_c_112_n PM_SKY130_FD_SC_HS__CLKINV_1%VGND
cc_1 VNB N_A_M1002_g 0.027297f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=0.58
cc_2 VNB A 0.0282826f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_3 VNB N_A_c_28_n 0.0453666f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.425
cc_4 VNB N_A_c_29_n 0.0578814f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.085
cc_5 VNB N_A_c_30_n 0.00540078f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.765
cc_6 VNB N_VPWR_c_60_n 0.0641695f $X=-0.19 $Y=-0.245 $X2=0.44 $Y2=1.085
cc_7 VNB N_Y_c_81_n 0.00750462f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_8 VNB Y 0.0520536f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.615
cc_9 VNB N_Y_c_83_n 0.0160574f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.765
cc_10 VNB N_VGND_c_109_n 0.0122168f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=0.92
cc_11 VNB N_VGND_c_110_n 0.0282119f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=0.58
cc_12 VNB N_VGND_c_111_n 0.0282669f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_13 VNB N_VGND_c_112_n 0.11676f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VPB N_A_c_31_n 0.0177391f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=2.045
cc_15 VPB N_A_c_32_n 0.0171946f $X=-0.19 $Y=1.66 $X2=0.945 $Y2=2.045
cc_16 VPB A 0.0116764f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_17 VPB N_A_c_30_n 0.0620411f $X=-0.19 $Y=1.66 $X2=0.59 $Y2=1.765
cc_18 VPB N_VPWR_c_61_n 0.0103331f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_19 VPB N_VPWR_c_62_n 0.0473336f $X=-0.19 $Y=1.66 $X2=0.945 $Y2=2.54
cc_20 VPB N_VPWR_c_63_n 0.0116916f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.21
cc_21 VPB N_VPWR_c_64_n 0.0238695f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_22 VPB N_VPWR_c_65_n 0.0183948f $X=-0.19 $Y=1.66 $X2=0.72 $Y2=1.425
cc_23 VPB N_VPWR_c_60_n 0.0500475f $X=-0.19 $Y=1.66 $X2=0.44 $Y2=1.085
cc_24 VPB Y 0.0231436f $X=-0.19 $Y=1.66 $X2=0.72 $Y2=1.615
cc_25 VPB N_Y_c_85_n 0.0188872f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_26 N_A_c_31_n N_VPWR_c_62_n 0.0100772f $X=0.495 $Y=2.045 $X2=0 $Y2=0
cc_27 A N_VPWR_c_62_n 0.0136621f $X=0.155 $Y=1.58 $X2=0 $Y2=0
cc_28 N_A_c_31_n N_VPWR_c_64_n 4.01546e-19 $X=0.495 $Y=2.045 $X2=0 $Y2=0
cc_29 N_A_c_32_n N_VPWR_c_64_n 0.00896977f $X=0.945 $Y=2.045 $X2=0 $Y2=0
cc_30 N_A_c_31_n N_VPWR_c_65_n 0.00445915f $X=0.495 $Y=2.045 $X2=0 $Y2=0
cc_31 N_A_c_32_n N_VPWR_c_65_n 0.00413917f $X=0.945 $Y=2.045 $X2=0 $Y2=0
cc_32 N_A_c_31_n N_VPWR_c_60_n 0.0086132f $X=0.495 $Y=2.045 $X2=0 $Y2=0
cc_33 N_A_c_32_n N_VPWR_c_60_n 0.00817726f $X=0.945 $Y=2.045 $X2=0 $Y2=0
cc_34 N_A_c_31_n N_Y_c_86_n 0.00722275f $X=0.495 $Y=2.045 $X2=0 $Y2=0
cc_35 N_A_M1002_g N_Y_c_81_n 0.00458999f $X=0.565 $Y=0.58 $X2=0 $Y2=0
cc_36 A N_Y_c_81_n 0.00696579f $X=0.155 $Y=1.58 $X2=0 $Y2=0
cc_37 N_A_c_29_n N_Y_c_81_n 0.0121436f $X=0.59 $Y=1.085 $X2=0 $Y2=0
cc_38 N_A_M1002_g Y 0.00534936f $X=0.565 $Y=0.58 $X2=0 $Y2=0
cc_39 N_A_c_32_n Y 0.00218078f $X=0.945 $Y=2.045 $X2=0 $Y2=0
cc_40 A Y 0.0489624f $X=0.155 $Y=1.58 $X2=0 $Y2=0
cc_41 N_A_c_29_n Y 0.0372247f $X=0.59 $Y=1.085 $X2=0 $Y2=0
cc_42 N_A_c_31_n N_Y_c_85_n 0.00405592f $X=0.495 $Y=2.045 $X2=0 $Y2=0
cc_43 N_A_c_32_n N_Y_c_85_n 0.0250371f $X=0.945 $Y=2.045 $X2=0 $Y2=0
cc_44 A N_Y_c_85_n 0.0167215f $X=0.155 $Y=1.58 $X2=0 $Y2=0
cc_45 N_A_c_30_n N_Y_c_85_n 0.00764814f $X=0.59 $Y=1.765 $X2=0 $Y2=0
cc_46 N_A_M1002_g N_VGND_c_110_n 0.0124698f $X=0.565 $Y=0.58 $X2=0 $Y2=0
cc_47 A N_VGND_c_110_n 0.0151075f $X=0.155 $Y=1.58 $X2=0 $Y2=0
cc_48 N_A_c_29_n N_VGND_c_110_n 7.38054e-19 $X=0.59 $Y=1.085 $X2=0 $Y2=0
cc_49 N_A_M1002_g N_VGND_c_111_n 0.00433162f $X=0.565 $Y=0.58 $X2=0 $Y2=0
cc_50 N_A_M1002_g N_VGND_c_112_n 0.00825282f $X=0.565 $Y=0.58 $X2=0 $Y2=0
cc_51 N_VPWR_c_62_n N_Y_c_86_n 0.0347719f $X=0.27 $Y=2.265 $X2=0 $Y2=0
cc_52 N_VPWR_c_65_n N_Y_c_86_n 0.00933236f $X=1.005 $Y=3.33 $X2=0 $Y2=0
cc_53 N_VPWR_c_60_n N_Y_c_86_n 0.00993985f $X=1.2 $Y=3.33 $X2=0 $Y2=0
cc_54 N_VPWR_M1001_d N_Y_c_85_n 0.00426951f $X=1.02 $Y=2.12 $X2=0 $Y2=0
cc_55 N_VPWR_c_62_n N_Y_c_85_n 0.0233786f $X=0.27 $Y=2.265 $X2=0 $Y2=0
cc_56 N_VPWR_c_64_n N_Y_c_85_n 0.0222202f $X=1.17 $Y=2.79 $X2=0 $Y2=0
cc_57 N_Y_c_81_n N_VGND_c_110_n 0.0146598f $X=1.085 $Y=0.515 $X2=0 $Y2=0
cc_58 N_Y_c_81_n N_VGND_c_111_n 0.0197467f $X=1.085 $Y=0.515 $X2=0 $Y2=0
cc_59 N_Y_c_83_n N_VGND_c_111_n 0.010709f $X=1.205 $Y=0.68 $X2=0 $Y2=0
cc_60 N_Y_c_81_n N_VGND_c_112_n 0.0168182f $X=1.085 $Y=0.515 $X2=0 $Y2=0
cc_61 N_Y_c_83_n N_VGND_c_112_n 0.008864f $X=1.205 $Y=0.68 $X2=0 $Y2=0
