* File: sky130_fd_sc_hs__a221o_2.pxi.spice
* Created: Tue Sep  1 19:50:14 2020
* 
x_PM_SKY130_FD_SC_HS__A221O_2%A_89_260# N_A_89_260#_M1000_d N_A_89_260#_M1013_d
+ N_A_89_260#_M1012_d N_A_89_260#_c_95_n N_A_89_260#_M1003_g N_A_89_260#_M1001_g
+ N_A_89_260#_M1002_g N_A_89_260#_c_96_n N_A_89_260#_M1004_g N_A_89_260#_c_88_n
+ N_A_89_260#_c_89_n N_A_89_260#_c_107_p N_A_89_260#_c_191_p N_A_89_260#_c_90_n
+ N_A_89_260#_c_91_n N_A_89_260#_c_92_n N_A_89_260#_c_98_n N_A_89_260#_c_99_n
+ N_A_89_260#_c_100_n N_A_89_260#_c_93_n N_A_89_260#_c_94_n
+ PM_SKY130_FD_SC_HS__A221O_2%A_89_260#
x_PM_SKY130_FD_SC_HS__A221O_2%A2 N_A2_c_214_n N_A2_c_219_n N_A2_M1005_g
+ N_A2_M1007_g A2 N_A2_c_216_n N_A2_c_217_n PM_SKY130_FD_SC_HS__A221O_2%A2
x_PM_SKY130_FD_SC_HS__A221O_2%A1 N_A1_c_259_n N_A1_M1006_g N_A1_M1000_g A1
+ PM_SKY130_FD_SC_HS__A221O_2%A1
x_PM_SKY130_FD_SC_HS__A221O_2%B1 N_B1_c_296_n N_B1_M1010_g N_B1_M1008_g
+ N_B1_c_293_n N_B1_c_294_n B1 PM_SKY130_FD_SC_HS__A221O_2%B1
x_PM_SKY130_FD_SC_HS__A221O_2%B2 N_B2_M1009_g N_B2_c_336_n N_B2_c_341_n
+ N_B2_M1011_g B2 N_B2_c_338_n N_B2_c_339_n PM_SKY130_FD_SC_HS__A221O_2%B2
x_PM_SKY130_FD_SC_HS__A221O_2%C1 N_C1_M1012_g N_C1_c_376_n N_C1_M1013_g
+ N_C1_c_377_n N_C1_c_381_n C1 N_C1_c_379_n PM_SKY130_FD_SC_HS__A221O_2%C1
x_PM_SKY130_FD_SC_HS__A221O_2%VPWR N_VPWR_M1003_s N_VPWR_M1004_s N_VPWR_M1006_d
+ N_VPWR_c_407_n N_VPWR_c_408_n N_VPWR_c_409_n N_VPWR_c_410_n N_VPWR_c_411_n
+ VPWR N_VPWR_c_412_n N_VPWR_c_413_n N_VPWR_c_406_n N_VPWR_c_415_n
+ N_VPWR_c_416_n PM_SKY130_FD_SC_HS__A221O_2%VPWR
x_PM_SKY130_FD_SC_HS__A221O_2%X N_X_M1001_d N_X_M1003_d N_X_c_465_n N_X_c_466_n
+ N_X_c_467_n N_X_c_470_n N_X_c_471_n N_X_c_468_n X X X N_X_c_472_n X
+ PM_SKY130_FD_SC_HS__A221O_2%X
x_PM_SKY130_FD_SC_HS__A221O_2%A_316_392# N_A_316_392#_M1005_d
+ N_A_316_392#_M1010_d N_A_316_392#_c_511_n N_A_316_392#_c_512_n
+ N_A_316_392#_c_513_n N_A_316_392#_c_515_n N_A_316_392#_c_514_n
+ N_A_316_392#_c_516_n PM_SKY130_FD_SC_HS__A221O_2%A_316_392#
x_PM_SKY130_FD_SC_HS__A221O_2%A_515_392# N_A_515_392#_M1010_s
+ N_A_515_392#_M1011_d N_A_515_392#_c_553_n N_A_515_392#_c_554_n
+ N_A_515_392#_c_555_n N_A_515_392#_c_557_n
+ PM_SKY130_FD_SC_HS__A221O_2%A_515_392#
x_PM_SKY130_FD_SC_HS__A221O_2%VGND N_VGND_M1001_s N_VGND_M1002_s N_VGND_M1009_d
+ N_VGND_c_583_n N_VGND_c_584_n N_VGND_c_585_n N_VGND_c_586_n VGND
+ N_VGND_c_587_n N_VGND_c_588_n N_VGND_c_589_n N_VGND_c_590_n N_VGND_c_591_n
+ N_VGND_c_592_n PM_SKY130_FD_SC_HS__A221O_2%VGND
cc_1 VNB N_A_89_260#_M1001_g 0.0225612f $X=-0.19 $Y=-0.245 $X2=0.555 $Y2=0.74
cc_2 VNB N_A_89_260#_M1002_g 0.0215418f $X=-0.19 $Y=-0.245 $X2=0.985 $Y2=0.74
cc_3 VNB N_A_89_260#_c_88_n 0.00487008f $X=-0.19 $Y=-0.245 $X2=1.025 $Y2=1.465
cc_4 VNB N_A_89_260#_c_89_n 0.0018925f $X=-0.19 $Y=-0.245 $X2=1.11 $Y2=1.3
cc_5 VNB N_A_89_260#_c_90_n 0.00370085f $X=-0.19 $Y=-0.245 $X2=3.015 $Y2=1.72
cc_6 VNB N_A_89_260#_c_91_n 0.00827709f $X=-0.19 $Y=-0.245 $X2=3.89 $Y2=0.925
cc_7 VNB N_A_89_260#_c_92_n 0.0211949f $X=-0.19 $Y=-0.245 $X2=3.1 $Y2=0.925
cc_8 VNB N_A_89_260#_c_93_n 0.0215989f $X=-0.19 $Y=-0.245 $X2=4.055 $Y2=0.515
cc_9 VNB N_A_89_260#_c_94_n 0.0520328f $X=-0.19 $Y=-0.245 $X2=0.985 $Y2=1.532
cc_10 VNB N_A2_c_214_n 0.00331051f $X=-0.19 $Y=-0.245 $X2=3.915 $Y2=0.37
cc_11 VNB N_A2_M1007_g 0.0202188f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A2_c_216_n 0.0302333f $X=-0.19 $Y=-0.245 $X2=0.555 $Y2=1.3
cc_13 VNB N_A2_c_217_n 0.00614974f $X=-0.19 $Y=-0.245 $X2=0.555 $Y2=0.74
cc_14 VNB N_A1_c_259_n 0.0190052f $X=-0.19 $Y=-0.245 $X2=2.045 $Y2=0.37
cc_15 VNB N_A1_M1000_g 0.041392f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB A1 0.00165251f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_B1_M1008_g 0.0393008f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_B1_c_293_n 0.0226341f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_B1_c_294_n 0.00728357f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB B1 0.00359533f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=1.765
cc_21 VNB N_B2_c_336_n 0.00629801f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB B2 0.0064492f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_B2_c_338_n 0.0292541f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=2.4
cc_24 VNB N_B2_c_339_n 0.0171286f $X=-0.19 $Y=-0.245 $X2=0.555 $Y2=0.74
cc_25 VNB N_C1_c_376_n 0.024355f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_C1_c_377_n 0.00903766f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB C1 0.00666617f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=2.4
cc_28 VNB N_C1_c_379_n 0.0537945f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_VPWR_c_406_n 0.183584f $X=-0.19 $Y=-0.245 $X2=4.05 $Y2=1.89
cc_30 VNB N_X_c_465_n 0.0271257f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_X_c_466_n 0.00388534f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_X_c_467_n 0.0111704f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=1.765
cc_33 VNB N_X_c_468_n 0.00206666f $X=-0.19 $Y=-0.245 $X2=0.555 $Y2=0.74
cc_34 VNB N_VGND_c_583_n 0.0125919f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=1.765
cc_35 VNB N_VGND_c_584_n 0.0276293f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=2.4
cc_36 VNB N_VGND_c_585_n 0.00455857f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_586_n 0.00685406f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_587_n 0.0172524f $X=-0.19 $Y=-0.245 $X2=1.025 $Y2=1.465
cc_39 VNB N_VGND_c_588_n 0.0497854f $X=-0.19 $Y=-0.245 $X2=1.11 $Y2=1.09
cc_40 VNB N_VGND_c_589_n 0.0186742f $X=-0.19 $Y=-0.245 $X2=4.05 $Y2=1.89
cc_41 VNB N_VGND_c_590_n 0.257799f $X=-0.19 $Y=-0.245 $X2=4.05 $Y2=2.105
cc_42 VNB N_VGND_c_591_n 0.00971914f $X=-0.19 $Y=-0.245 $X2=4.055 $Y2=0.515
cc_43 VNB N_VGND_c_592_n 0.0069273f $X=-0.19 $Y=-0.245 $X2=2.725 $Y2=0.74
cc_44 VPB N_A_89_260#_c_95_n 0.0164244f $X=-0.19 $Y=1.66 $X2=0.54 $Y2=1.765
cc_45 VPB N_A_89_260#_c_96_n 0.0161704f $X=-0.19 $Y=1.66 $X2=0.99 $Y2=1.765
cc_46 VPB N_A_89_260#_c_90_n 5.72206e-19 $X=-0.19 $Y=1.66 $X2=3.015 $Y2=1.72
cc_47 VPB N_A_89_260#_c_98_n 0.0271121f $X=-0.19 $Y=1.66 $X2=3.885 $Y2=1.805
cc_48 VPB N_A_89_260#_c_99_n 9.2782e-19 $X=-0.19 $Y=1.66 $X2=3.1 $Y2=1.805
cc_49 VPB N_A_89_260#_c_100_n 0.0451244f $X=-0.19 $Y=1.66 $X2=4.05 $Y2=2.105
cc_50 VPB N_A_89_260#_c_94_n 0.0140194f $X=-0.19 $Y=1.66 $X2=0.985 $Y2=1.532
cc_51 VPB N_A2_c_214_n 0.00661751f $X=-0.19 $Y=1.66 $X2=3.915 $Y2=0.37
cc_52 VPB N_A2_c_219_n 0.0231724f $X=-0.19 $Y=1.66 $X2=3.9 $Y2=1.96
cc_53 VPB N_A2_c_217_n 0.00523119f $X=-0.19 $Y=1.66 $X2=0.555 $Y2=0.74
cc_54 VPB N_A1_c_259_n 0.0429114f $X=-0.19 $Y=1.66 $X2=2.045 $Y2=0.37
cc_55 VPB A1 0.00101673f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_56 VPB N_B1_c_296_n 0.0185476f $X=-0.19 $Y=1.66 $X2=2.045 $Y2=0.37
cc_57 VPB N_B1_c_293_n 0.0172704f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_58 VPB N_B1_c_294_n 0.0130302f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_59 VPB B1 0.00280744f $X=-0.19 $Y=1.66 $X2=0.54 $Y2=1.765
cc_60 VPB N_B2_c_336_n 0.00682148f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_61 VPB N_B2_c_341_n 0.0198828f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_62 VPB N_C1_c_377_n 0.00901237f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_63 VPB N_C1_c_381_n 0.0264129f $X=-0.19 $Y=1.66 $X2=0.54 $Y2=1.765
cc_64 VPB N_VPWR_c_407_n 0.0117686f $X=-0.19 $Y=1.66 $X2=0.54 $Y2=1.765
cc_65 VPB N_VPWR_c_408_n 0.0434034f $X=-0.19 $Y=1.66 $X2=0.54 $Y2=2.4
cc_66 VPB N_VPWR_c_409_n 0.0206041f $X=-0.19 $Y=1.66 $X2=0.555 $Y2=0.74
cc_67 VPB N_VPWR_c_410_n 0.00909434f $X=-0.19 $Y=1.66 $X2=0.985 $Y2=0.74
cc_68 VPB N_VPWR_c_411_n 0.0127089f $X=-0.19 $Y=1.66 $X2=1.025 $Y2=1.465
cc_69 VPB N_VPWR_c_412_n 0.018048f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_70 VPB N_VPWR_c_413_n 0.05134f $X=-0.19 $Y=1.66 $X2=3.1 $Y2=1.805
cc_71 VPB N_VPWR_c_406_n 0.0793798f $X=-0.19 $Y=1.66 $X2=4.05 $Y2=1.89
cc_72 VPB N_VPWR_c_415_n 0.0047828f $X=-0.19 $Y=1.66 $X2=4.055 $Y2=0.84
cc_73 VPB N_VPWR_c_416_n 0.00614127f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_74 VPB N_X_c_465_n 0.00726159f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_75 VPB N_X_c_470_n 0.00183065f $X=-0.19 $Y=1.66 $X2=0.54 $Y2=2.4
cc_76 VPB N_X_c_471_n 0.010032f $X=-0.19 $Y=1.66 $X2=0.54 $Y2=2.4
cc_77 VPB N_X_c_472_n 0.00183475f $X=-0.19 $Y=1.66 $X2=1.025 $Y2=1.465
cc_78 VPB X 0.00257348f $X=-0.19 $Y=1.66 $X2=0.95 $Y2=1.465
cc_79 VPB N_A_316_392#_c_511_n 0.00351688f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_80 VPB N_A_316_392#_c_512_n 0.00216998f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_81 VPB N_A_316_392#_c_513_n 0.0189278f $X=-0.19 $Y=1.66 $X2=0.54 $Y2=2.4
cc_82 VPB N_A_316_392#_c_514_n 0.00372599f $X=-0.19 $Y=1.66 $X2=0.985 $Y2=0.74
cc_83 VPB N_A_515_392#_c_553_n 0.0048276f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_84 VPB N_A_515_392#_c_554_n 0.00566895f $X=-0.19 $Y=1.66 $X2=0.54 $Y2=2.4
cc_85 VPB N_A_515_392#_c_555_n 0.00375341f $X=-0.19 $Y=1.66 $X2=0.54 $Y2=2.4
cc_86 N_A_89_260#_c_96_n N_A2_c_214_n 0.00439757f $X=0.99 $Y=1.765 $X2=0 $Y2=0
cc_87 N_A_89_260#_c_94_n N_A2_c_214_n 0.00610827f $X=0.985 $Y=1.532 $X2=0 $Y2=0
cc_88 N_A_89_260#_c_96_n N_A2_c_219_n 0.0167057f $X=0.99 $Y=1.765 $X2=0 $Y2=0
cc_89 N_A_89_260#_M1002_g N_A2_M1007_g 0.0222151f $X=0.985 $Y=0.74 $X2=0 $Y2=0
cc_90 N_A_89_260#_c_89_n N_A2_M1007_g 0.00309845f $X=1.11 $Y=1.3 $X2=0 $Y2=0
cc_91 N_A_89_260#_c_107_p N_A2_M1007_g 0.0146908f $X=2.02 $Y=1.005 $X2=0 $Y2=0
cc_92 N_A_89_260#_c_92_n N_A2_M1007_g 0.00212646f $X=3.1 $Y=0.925 $X2=0 $Y2=0
cc_93 N_A_89_260#_M1002_g N_A2_c_216_n 0.00157459f $X=0.985 $Y=0.74 $X2=0 $Y2=0
cc_94 N_A_89_260#_c_88_n N_A2_c_216_n 0.00191799f $X=1.025 $Y=1.465 $X2=0 $Y2=0
cc_95 N_A_89_260#_c_89_n N_A2_c_216_n 2.5812e-19 $X=1.11 $Y=1.3 $X2=0 $Y2=0
cc_96 N_A_89_260#_c_107_p N_A2_c_216_n 0.00146918f $X=2.02 $Y=1.005 $X2=0 $Y2=0
cc_97 N_A_89_260#_c_94_n N_A2_c_216_n 0.0153101f $X=0.985 $Y=1.532 $X2=0 $Y2=0
cc_98 N_A_89_260#_c_96_n N_A2_c_217_n 3.202e-19 $X=0.99 $Y=1.765 $X2=0 $Y2=0
cc_99 N_A_89_260#_c_88_n N_A2_c_217_n 0.0283357f $X=1.025 $Y=1.465 $X2=0 $Y2=0
cc_100 N_A_89_260#_c_89_n N_A2_c_217_n 0.00301343f $X=1.11 $Y=1.3 $X2=0 $Y2=0
cc_101 N_A_89_260#_c_107_p N_A2_c_217_n 0.0264353f $X=2.02 $Y=1.005 $X2=0 $Y2=0
cc_102 N_A_89_260#_c_94_n N_A2_c_217_n 0.00338938f $X=0.985 $Y=1.532 $X2=0 $Y2=0
cc_103 N_A_89_260#_c_92_n N_A1_c_259_n 0.00426639f $X=3.1 $Y=0.925 $X2=-0.19
+ $Y2=-0.245
cc_104 N_A_89_260#_c_107_p N_A1_M1000_g 0.012453f $X=2.02 $Y=1.005 $X2=0 $Y2=0
cc_105 N_A_89_260#_c_92_n N_A1_M1000_g 0.0138295f $X=3.1 $Y=0.925 $X2=0 $Y2=0
cc_106 N_A_89_260#_c_107_p A1 0.00330514f $X=2.02 $Y=1.005 $X2=0 $Y2=0
cc_107 N_A_89_260#_c_92_n A1 0.013448f $X=3.1 $Y=0.925 $X2=0 $Y2=0
cc_108 N_A_89_260#_c_99_n N_B1_c_296_n 0.00104043f $X=3.1 $Y=1.805 $X2=-0.19
+ $Y2=-0.245
cc_109 N_A_89_260#_c_90_n N_B1_M1008_g 0.0156215f $X=3.015 $Y=1.72 $X2=0 $Y2=0
cc_110 N_A_89_260#_c_92_n N_B1_M1008_g 0.0234179f $X=3.1 $Y=0.925 $X2=0 $Y2=0
cc_111 N_A_89_260#_c_92_n N_B1_c_293_n 0.00628063f $X=3.1 $Y=0.925 $X2=0 $Y2=0
cc_112 N_A_89_260#_c_90_n N_B1_c_294_n 0.00700708f $X=3.015 $Y=1.72 $X2=0 $Y2=0
cc_113 N_A_89_260#_c_99_n N_B1_c_294_n 0.00890858f $X=3.1 $Y=1.805 $X2=0 $Y2=0
cc_114 N_A_89_260#_c_90_n B1 0.019126f $X=3.015 $Y=1.72 $X2=0 $Y2=0
cc_115 N_A_89_260#_c_92_n B1 0.0160096f $X=3.1 $Y=0.925 $X2=0 $Y2=0
cc_116 N_A_89_260#_c_99_n B1 0.00476236f $X=3.1 $Y=1.805 $X2=0 $Y2=0
cc_117 N_A_89_260#_c_90_n N_B2_c_336_n 0.00343645f $X=3.015 $Y=1.72 $X2=0 $Y2=0
cc_118 N_A_89_260#_c_98_n N_B2_c_336_n 0.00538403f $X=3.885 $Y=1.805 $X2=0 $Y2=0
cc_119 N_A_89_260#_c_98_n N_B2_c_341_n 0.010248f $X=3.885 $Y=1.805 $X2=0 $Y2=0
cc_120 N_A_89_260#_c_100_n N_B2_c_341_n 0.00102747f $X=4.05 $Y=2.105 $X2=0 $Y2=0
cc_121 N_A_89_260#_c_90_n B2 0.0282982f $X=3.015 $Y=1.72 $X2=0 $Y2=0
cc_122 N_A_89_260#_c_91_n B2 0.0306748f $X=3.89 $Y=0.925 $X2=0 $Y2=0
cc_123 N_A_89_260#_c_98_n B2 0.0321363f $X=3.885 $Y=1.805 $X2=0 $Y2=0
cc_124 N_A_89_260#_c_91_n N_B2_c_338_n 0.00101381f $X=3.89 $Y=0.925 $X2=0 $Y2=0
cc_125 N_A_89_260#_c_98_n N_B2_c_338_n 0.00428104f $X=3.885 $Y=1.805 $X2=0 $Y2=0
cc_126 N_A_89_260#_c_90_n N_B2_c_339_n 0.0031703f $X=3.015 $Y=1.72 $X2=0 $Y2=0
cc_127 N_A_89_260#_c_91_n N_B2_c_339_n 0.0129716f $X=3.89 $Y=0.925 $X2=0 $Y2=0
cc_128 N_A_89_260#_c_92_n N_B2_c_339_n 0.00509793f $X=3.1 $Y=0.925 $X2=0 $Y2=0
cc_129 N_A_89_260#_c_93_n N_B2_c_339_n 6.8223e-19 $X=4.055 $Y=0.515 $X2=0 $Y2=0
cc_130 N_A_89_260#_c_91_n N_C1_c_376_n 0.0128498f $X=3.89 $Y=0.925 $X2=0 $Y2=0
cc_131 N_A_89_260#_c_93_n N_C1_c_376_n 0.00767918f $X=4.055 $Y=0.515 $X2=0 $Y2=0
cc_132 N_A_89_260#_c_98_n N_C1_c_377_n 0.0083321f $X=3.885 $Y=1.805 $X2=0 $Y2=0
cc_133 N_A_89_260#_c_98_n N_C1_c_381_n 0.01108f $X=3.885 $Y=1.805 $X2=0 $Y2=0
cc_134 N_A_89_260#_c_100_n N_C1_c_381_n 0.0142524f $X=4.05 $Y=2.105 $X2=0 $Y2=0
cc_135 N_A_89_260#_c_91_n C1 0.0255964f $X=3.89 $Y=0.925 $X2=0 $Y2=0
cc_136 N_A_89_260#_c_98_n C1 0.0275993f $X=3.885 $Y=1.805 $X2=0 $Y2=0
cc_137 N_A_89_260#_c_91_n N_C1_c_379_n 0.00180924f $X=3.89 $Y=0.925 $X2=0 $Y2=0
cc_138 N_A_89_260#_c_98_n N_C1_c_379_n 0.00220821f $X=3.885 $Y=1.805 $X2=0 $Y2=0
cc_139 N_A_89_260#_c_95_n N_VPWR_c_408_n 0.00993564f $X=0.54 $Y=1.765 $X2=0
+ $Y2=0
cc_140 N_A_89_260#_c_95_n N_VPWR_c_409_n 0.00445602f $X=0.54 $Y=1.765 $X2=0
+ $Y2=0
cc_141 N_A_89_260#_c_96_n N_VPWR_c_409_n 0.00445602f $X=0.99 $Y=1.765 $X2=0
+ $Y2=0
cc_142 N_A_89_260#_c_96_n N_VPWR_c_410_n 0.00653824f $X=0.99 $Y=1.765 $X2=0
+ $Y2=0
cc_143 N_A_89_260#_c_88_n N_VPWR_c_410_n 0.00374449f $X=1.025 $Y=1.465 $X2=0
+ $Y2=0
cc_144 N_A_89_260#_c_100_n N_VPWR_c_413_n 0.0145938f $X=4.05 $Y=2.105 $X2=0
+ $Y2=0
cc_145 N_A_89_260#_c_95_n N_VPWR_c_406_n 0.00861194f $X=0.54 $Y=1.765 $X2=0
+ $Y2=0
cc_146 N_A_89_260#_c_96_n N_VPWR_c_406_n 0.00858225f $X=0.99 $Y=1.765 $X2=0
+ $Y2=0
cc_147 N_A_89_260#_c_100_n N_VPWR_c_406_n 0.0120466f $X=4.05 $Y=2.105 $X2=0
+ $Y2=0
cc_148 N_A_89_260#_c_95_n N_X_c_465_n 0.00126333f $X=0.54 $Y=1.765 $X2=0 $Y2=0
cc_149 N_A_89_260#_M1001_g N_X_c_465_n 0.00617799f $X=0.555 $Y=0.74 $X2=0 $Y2=0
cc_150 N_A_89_260#_c_88_n N_X_c_465_n 0.024635f $X=1.025 $Y=1.465 $X2=0 $Y2=0
cc_151 N_A_89_260#_c_94_n N_X_c_465_n 0.0145794f $X=0.985 $Y=1.532 $X2=0 $Y2=0
cc_152 N_A_89_260#_M1001_g N_X_c_466_n 0.0142424f $X=0.555 $Y=0.74 $X2=0 $Y2=0
cc_153 N_A_89_260#_c_88_n N_X_c_466_n 0.0266522f $X=1.025 $Y=1.465 $X2=0 $Y2=0
cc_154 N_A_89_260#_c_89_n N_X_c_466_n 0.00221378f $X=1.11 $Y=1.3 $X2=0 $Y2=0
cc_155 N_A_89_260#_c_94_n N_X_c_466_n 0.00337043f $X=0.985 $Y=1.532 $X2=0 $Y2=0
cc_156 N_A_89_260#_c_95_n N_X_c_470_n 0.0142646f $X=0.54 $Y=1.765 $X2=0 $Y2=0
cc_157 N_A_89_260#_c_88_n N_X_c_470_n 0.00532205f $X=1.025 $Y=1.465 $X2=0 $Y2=0
cc_158 N_A_89_260#_c_94_n N_X_c_470_n 6.544e-19 $X=0.985 $Y=1.532 $X2=0 $Y2=0
cc_159 N_A_89_260#_M1001_g N_X_c_468_n 0.0128625f $X=0.555 $Y=0.74 $X2=0 $Y2=0
cc_160 N_A_89_260#_M1002_g N_X_c_468_n 3.97481e-19 $X=0.985 $Y=0.74 $X2=0 $Y2=0
cc_161 N_A_89_260#_c_95_n N_X_c_472_n 9.3899e-19 $X=0.54 $Y=1.765 $X2=0 $Y2=0
cc_162 N_A_89_260#_c_96_n N_X_c_472_n 0.00396299f $X=0.99 $Y=1.765 $X2=0 $Y2=0
cc_163 N_A_89_260#_c_88_n N_X_c_472_n 0.0276943f $X=1.025 $Y=1.465 $X2=0 $Y2=0
cc_164 N_A_89_260#_c_94_n N_X_c_472_n 0.00792231f $X=0.985 $Y=1.532 $X2=0 $Y2=0
cc_165 N_A_89_260#_c_95_n X 0.017229f $X=0.54 $Y=1.765 $X2=0 $Y2=0
cc_166 N_A_89_260#_c_96_n X 0.0113742f $X=0.99 $Y=1.765 $X2=0 $Y2=0
cc_167 N_A_89_260#_c_99_n N_A_316_392#_c_515_n 0.00415559f $X=3.1 $Y=1.805 $X2=0
+ $Y2=0
cc_168 N_A_89_260#_c_98_n N_A_316_392#_c_516_n 0.0150347f $X=3.885 $Y=1.805
+ $X2=0 $Y2=0
cc_169 N_A_89_260#_c_99_n N_A_316_392#_c_516_n 0.00780121f $X=3.1 $Y=1.805 $X2=0
+ $Y2=0
cc_170 N_A_89_260#_c_100_n N_A_515_392#_c_554_n 0.00549849f $X=4.05 $Y=2.105
+ $X2=0 $Y2=0
cc_171 N_A_89_260#_c_98_n N_A_515_392#_c_557_n 0.0138919f $X=3.885 $Y=1.805
+ $X2=0 $Y2=0
cc_172 N_A_89_260#_c_100_n N_A_515_392#_c_557_n 0.0550085f $X=4.05 $Y=2.105
+ $X2=0 $Y2=0
cc_173 N_A_89_260#_c_89_n N_VGND_M1002_s 2.53259e-19 $X=1.11 $Y=1.3 $X2=0 $Y2=0
cc_174 N_A_89_260#_c_107_p N_VGND_M1002_s 0.0111394f $X=2.02 $Y=1.005 $X2=0
+ $Y2=0
cc_175 N_A_89_260#_c_191_p N_VGND_M1002_s 8.64304e-19 $X=1.195 $Y=1.005 $X2=0
+ $Y2=0
cc_176 N_A_89_260#_c_91_n N_VGND_M1009_d 0.00620519f $X=3.89 $Y=0.925 $X2=0
+ $Y2=0
cc_177 N_A_89_260#_M1001_g N_VGND_c_584_n 0.00466772f $X=0.555 $Y=0.74 $X2=0
+ $Y2=0
cc_178 N_A_89_260#_M1001_g N_VGND_c_585_n 4.81239e-19 $X=0.555 $Y=0.74 $X2=0
+ $Y2=0
cc_179 N_A_89_260#_M1002_g N_VGND_c_585_n 0.0157538f $X=0.985 $Y=0.74 $X2=0
+ $Y2=0
cc_180 N_A_89_260#_c_107_p N_VGND_c_585_n 0.0248162f $X=2.02 $Y=1.005 $X2=0
+ $Y2=0
cc_181 N_A_89_260#_c_191_p N_VGND_c_585_n 0.00909352f $X=1.195 $Y=1.005 $X2=0
+ $Y2=0
cc_182 N_A_89_260#_c_92_n N_VGND_c_585_n 0.0146878f $X=3.1 $Y=0.925 $X2=0 $Y2=0
cc_183 N_A_89_260#_c_91_n N_VGND_c_586_n 0.0237091f $X=3.89 $Y=0.925 $X2=0 $Y2=0
cc_184 N_A_89_260#_c_92_n N_VGND_c_586_n 0.0114504f $X=3.1 $Y=0.925 $X2=0 $Y2=0
cc_185 N_A_89_260#_c_93_n N_VGND_c_586_n 0.0128115f $X=4.055 $Y=0.515 $X2=0
+ $Y2=0
cc_186 N_A_89_260#_M1001_g N_VGND_c_587_n 0.00434272f $X=0.555 $Y=0.74 $X2=0
+ $Y2=0
cc_187 N_A_89_260#_M1002_g N_VGND_c_587_n 0.00383152f $X=0.985 $Y=0.74 $X2=0
+ $Y2=0
cc_188 N_A_89_260#_c_92_n N_VGND_c_588_n 0.0386707f $X=3.1 $Y=0.925 $X2=0 $Y2=0
cc_189 N_A_89_260#_c_93_n N_VGND_c_589_n 0.0145323f $X=4.055 $Y=0.515 $X2=0
+ $Y2=0
cc_190 N_A_89_260#_M1001_g N_VGND_c_590_n 0.0082413f $X=0.555 $Y=0.74 $X2=0
+ $Y2=0
cc_191 N_A_89_260#_M1002_g N_VGND_c_590_n 0.0075754f $X=0.985 $Y=0.74 $X2=0
+ $Y2=0
cc_192 N_A_89_260#_c_91_n N_VGND_c_590_n 0.013929f $X=3.89 $Y=0.925 $X2=0 $Y2=0
cc_193 N_A_89_260#_c_92_n N_VGND_c_590_n 0.039097f $X=3.1 $Y=0.925 $X2=0 $Y2=0
cc_194 N_A_89_260#_c_93_n N_VGND_c_590_n 0.0119861f $X=4.055 $Y=0.515 $X2=0
+ $Y2=0
cc_195 N_A_89_260#_c_107_p A_337_74# 0.00672031f $X=2.02 $Y=1.005 $X2=-0.19
+ $Y2=-0.245
cc_196 N_A_89_260#_c_91_n A_603_74# 0.00390345f $X=3.89 $Y=0.925 $X2=-0.19
+ $Y2=-0.245
cc_197 N_A_89_260#_c_92_n A_603_74# 0.00199923f $X=3.1 $Y=0.925 $X2=-0.19
+ $Y2=-0.245
cc_198 N_A2_c_214_n N_A1_c_259_n 0.0133265f $X=1.505 $Y=1.795 $X2=-0.19
+ $Y2=-0.245
cc_199 N_A2_c_219_n N_A1_c_259_n 0.00842601f $X=1.505 $Y=1.885 $X2=-0.19
+ $Y2=-0.245
cc_200 N_A2_c_216_n N_A1_c_259_n 0.040834f $X=1.52 $Y=1.425 $X2=-0.19 $Y2=-0.245
cc_201 N_A2_c_217_n N_A1_c_259_n 4.02526e-19 $X=1.52 $Y=1.425 $X2=-0.19
+ $Y2=-0.245
cc_202 N_A2_M1007_g N_A1_M1000_g 0.040834f $X=1.61 $Y=0.74 $X2=0 $Y2=0
cc_203 N_A2_c_217_n N_A1_M1000_g 0.00666653f $X=1.52 $Y=1.425 $X2=0 $Y2=0
cc_204 N_A2_c_217_n A1 0.026544f $X=1.52 $Y=1.425 $X2=0 $Y2=0
cc_205 N_A2_c_219_n N_VPWR_c_410_n 0.00720533f $X=1.505 $Y=1.885 $X2=0 $Y2=0
cc_206 N_A2_c_216_n N_VPWR_c_410_n 4.65628e-19 $X=1.52 $Y=1.425 $X2=0 $Y2=0
cc_207 N_A2_c_217_n N_VPWR_c_410_n 0.00119394f $X=1.52 $Y=1.425 $X2=0 $Y2=0
cc_208 N_A2_c_219_n N_VPWR_c_411_n 5.53241e-19 $X=1.505 $Y=1.885 $X2=0 $Y2=0
cc_209 N_A2_c_219_n N_VPWR_c_412_n 0.00445602f $X=1.505 $Y=1.885 $X2=0 $Y2=0
cc_210 N_A2_c_219_n N_VPWR_c_406_n 0.00857973f $X=1.505 $Y=1.885 $X2=0 $Y2=0
cc_211 N_A2_c_219_n N_X_c_472_n 6.9999e-19 $X=1.505 $Y=1.885 $X2=0 $Y2=0
cc_212 N_A2_c_219_n N_A_316_392#_c_511_n 0.00248425f $X=1.505 $Y=1.885 $X2=0
+ $Y2=0
cc_213 N_A2_c_216_n N_A_316_392#_c_511_n 4.52853e-19 $X=1.52 $Y=1.425 $X2=0
+ $Y2=0
cc_214 N_A2_c_217_n N_A_316_392#_c_511_n 0.0180777f $X=1.52 $Y=1.425 $X2=0 $Y2=0
cc_215 N_A2_c_219_n N_A_316_392#_c_512_n 0.00883546f $X=1.505 $Y=1.885 $X2=0
+ $Y2=0
cc_216 N_A2_M1007_g N_VGND_c_585_n 0.017959f $X=1.61 $Y=0.74 $X2=0 $Y2=0
cc_217 N_A2_M1007_g N_VGND_c_588_n 0.00383152f $X=1.61 $Y=0.74 $X2=0 $Y2=0
cc_218 N_A2_M1007_g N_VGND_c_590_n 0.0075694f $X=1.61 $Y=0.74 $X2=0 $Y2=0
cc_219 N_A1_c_259_n N_B1_c_293_n 0.0215154f $X=1.955 $Y=1.885 $X2=0 $Y2=0
cc_220 A1 N_B1_c_293_n 0.00199005f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_221 N_A1_c_259_n B1 3.86748e-19 $X=1.955 $Y=1.885 $X2=0 $Y2=0
cc_222 A1 B1 0.0249007f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_223 N_A1_c_259_n N_VPWR_c_411_n 0.0131469f $X=1.955 $Y=1.885 $X2=0 $Y2=0
cc_224 N_A1_c_259_n N_VPWR_c_412_n 0.00413917f $X=1.955 $Y=1.885 $X2=0 $Y2=0
cc_225 N_A1_c_259_n N_VPWR_c_406_n 0.0081781f $X=1.955 $Y=1.885 $X2=0 $Y2=0
cc_226 N_A1_c_259_n N_A_316_392#_c_512_n 0.00605728f $X=1.955 $Y=1.885 $X2=0
+ $Y2=0
cc_227 N_A1_c_259_n N_A_316_392#_c_513_n 0.021584f $X=1.955 $Y=1.885 $X2=0 $Y2=0
cc_228 A1 N_A_316_392#_c_513_n 0.0253213f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_229 N_A1_c_259_n N_A_316_392#_c_514_n 0.00248989f $X=1.955 $Y=1.885 $X2=0
+ $Y2=0
cc_230 N_A1_c_259_n N_A_515_392#_c_553_n 8.38149e-19 $X=1.955 $Y=1.885 $X2=0
+ $Y2=0
cc_231 N_A1_c_259_n N_A_515_392#_c_555_n 5.75404e-19 $X=1.955 $Y=1.885 $X2=0
+ $Y2=0
cc_232 N_A1_M1000_g N_VGND_c_585_n 0.00165077f $X=1.97 $Y=0.74 $X2=0 $Y2=0
cc_233 N_A1_M1000_g N_VGND_c_588_n 0.00433139f $X=1.97 $Y=0.74 $X2=0 $Y2=0
cc_234 N_A1_M1000_g N_VGND_c_590_n 0.00822f $X=1.97 $Y=0.74 $X2=0 $Y2=0
cc_235 N_B1_c_294_n N_B2_c_336_n 0.0151757f $X=2.925 $Y=1.667 $X2=0 $Y2=0
cc_236 N_B1_c_296_n N_B2_c_341_n 0.0182718f $X=2.925 $Y=1.885 $X2=0 $Y2=0
cc_237 N_B1_M1008_g B2 3.61351e-19 $X=2.94 $Y=0.74 $X2=0 $Y2=0
cc_238 N_B1_c_294_n N_B2_c_338_n 0.039474f $X=2.925 $Y=1.667 $X2=0 $Y2=0
cc_239 N_B1_M1008_g N_B2_c_339_n 0.039474f $X=2.94 $Y=0.74 $X2=0 $Y2=0
cc_240 N_B1_c_296_n N_VPWR_c_411_n 0.00322745f $X=2.925 $Y=1.885 $X2=0 $Y2=0
cc_241 N_B1_c_296_n N_VPWR_c_413_n 0.00278271f $X=2.925 $Y=1.885 $X2=0 $Y2=0
cc_242 N_B1_c_296_n N_VPWR_c_406_n 0.00358708f $X=2.925 $Y=1.885 $X2=0 $Y2=0
cc_243 N_B1_c_293_n N_A_316_392#_c_513_n 5.92156e-19 $X=2.835 $Y=1.615 $X2=0
+ $Y2=0
cc_244 B1 N_A_316_392#_c_513_n 0.00634428f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_245 N_B1_c_296_n N_A_316_392#_c_515_n 0.0130599f $X=2.925 $Y=1.885 $X2=0
+ $Y2=0
cc_246 N_B1_c_293_n N_A_316_392#_c_515_n 0.00205663f $X=2.835 $Y=1.615 $X2=0
+ $Y2=0
cc_247 B1 N_A_316_392#_c_515_n 0.00146447f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_248 N_B1_c_296_n N_A_316_392#_c_514_n 0.00508098f $X=2.925 $Y=1.885 $X2=0
+ $Y2=0
cc_249 N_B1_c_293_n N_A_316_392#_c_514_n 0.00137755f $X=2.835 $Y=1.615 $X2=0
+ $Y2=0
cc_250 B1 N_A_316_392#_c_514_n 0.0148325f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_251 N_B1_c_296_n N_A_316_392#_c_516_n 0.0104527f $X=2.925 $Y=1.885 $X2=0
+ $Y2=0
cc_252 N_B1_c_296_n N_A_515_392#_c_553_n 0.00749293f $X=2.925 $Y=1.885 $X2=0
+ $Y2=0
cc_253 N_B1_c_293_n N_A_515_392#_c_553_n 3.17745e-19 $X=2.835 $Y=1.615 $X2=0
+ $Y2=0
cc_254 N_B1_c_296_n N_A_515_392#_c_554_n 0.0127203f $X=2.925 $Y=1.885 $X2=0
+ $Y2=0
cc_255 N_B1_M1008_g N_VGND_c_586_n 0.00143798f $X=2.94 $Y=0.74 $X2=0 $Y2=0
cc_256 N_B1_M1008_g N_VGND_c_588_n 0.00433139f $X=2.94 $Y=0.74 $X2=0 $Y2=0
cc_257 N_B1_M1008_g N_VGND_c_590_n 0.00451185f $X=2.94 $Y=0.74 $X2=0 $Y2=0
cc_258 B2 N_C1_c_376_n 0.00274822f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_259 N_B2_c_339_n N_C1_c_376_n 0.0225661f $X=3.39 $Y=1.22 $X2=0 $Y2=0
cc_260 N_B2_c_336_n N_C1_c_377_n 0.0105012f $X=3.375 $Y=1.795 $X2=0 $Y2=0
cc_261 N_B2_c_336_n N_C1_c_381_n 0.00416562f $X=3.375 $Y=1.795 $X2=0 $Y2=0
cc_262 N_B2_c_341_n N_C1_c_381_n 0.0173788f $X=3.375 $Y=1.885 $X2=0 $Y2=0
cc_263 B2 C1 0.0298222f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_264 N_B2_c_338_n C1 2.69235e-19 $X=3.39 $Y=1.385 $X2=0 $Y2=0
cc_265 N_B2_c_338_n N_C1_c_379_n 0.0207972f $X=3.39 $Y=1.385 $X2=0 $Y2=0
cc_266 N_B2_c_341_n N_VPWR_c_413_n 0.00278271f $X=3.375 $Y=1.885 $X2=0 $Y2=0
cc_267 N_B2_c_341_n N_VPWR_c_406_n 0.0035399f $X=3.375 $Y=1.885 $X2=0 $Y2=0
cc_268 N_B2_c_341_n N_A_316_392#_c_516_n 0.00863518f $X=3.375 $Y=1.885 $X2=0
+ $Y2=0
cc_269 N_B2_c_341_n N_A_515_392#_c_554_n 0.0124529f $X=3.375 $Y=1.885 $X2=0
+ $Y2=0
cc_270 N_B2_c_341_n N_A_515_392#_c_557_n 0.00628847f $X=3.375 $Y=1.885 $X2=0
+ $Y2=0
cc_271 N_B2_c_339_n N_VGND_c_586_n 0.00959637f $X=3.39 $Y=1.22 $X2=0 $Y2=0
cc_272 N_B2_c_339_n N_VGND_c_588_n 0.00383152f $X=3.39 $Y=1.22 $X2=0 $Y2=0
cc_273 N_B2_c_339_n N_VGND_c_590_n 0.00383367f $X=3.39 $Y=1.22 $X2=0 $Y2=0
cc_274 N_C1_c_381_n N_VPWR_c_413_n 0.00445602f $X=3.832 $Y=1.885 $X2=0 $Y2=0
cc_275 N_C1_c_381_n N_VPWR_c_406_n 0.00861895f $X=3.832 $Y=1.885 $X2=0 $Y2=0
cc_276 N_C1_c_381_n N_A_515_392#_c_554_n 0.00341066f $X=3.832 $Y=1.885 $X2=0
+ $Y2=0
cc_277 N_C1_c_381_n N_A_515_392#_c_557_n 0.00353834f $X=3.832 $Y=1.885 $X2=0
+ $Y2=0
cc_278 N_C1_c_376_n N_VGND_c_586_n 0.0051057f $X=3.84 $Y=1.22 $X2=0 $Y2=0
cc_279 N_C1_c_376_n N_VGND_c_589_n 0.00434272f $X=3.84 $Y=1.22 $X2=0 $Y2=0
cc_280 N_C1_c_376_n N_VGND_c_590_n 0.00449471f $X=3.84 $Y=1.22 $X2=0 $Y2=0
cc_281 N_VPWR_M1003_s N_X_c_470_n 0.0010131f $X=0.19 $Y=1.84 $X2=0 $Y2=0
cc_282 N_VPWR_c_408_n N_X_c_470_n 0.00517047f $X=0.315 $Y=2.305 $X2=0 $Y2=0
cc_283 N_VPWR_M1003_s N_X_c_471_n 0.00228818f $X=0.19 $Y=1.84 $X2=0 $Y2=0
cc_284 N_VPWR_c_408_n N_X_c_471_n 0.0167277f $X=0.315 $Y=2.305 $X2=0 $Y2=0
cc_285 N_VPWR_c_410_n N_X_c_472_n 0.00142382f $X=1.215 $Y=2.115 $X2=0 $Y2=0
cc_286 N_VPWR_c_408_n X 0.0563525f $X=0.315 $Y=2.305 $X2=0 $Y2=0
cc_287 N_VPWR_c_409_n X 0.014552f $X=1.13 $Y=3.33 $X2=0 $Y2=0
cc_288 N_VPWR_c_410_n X 0.0677182f $X=1.215 $Y=2.115 $X2=0 $Y2=0
cc_289 N_VPWR_c_406_n X 0.0119791f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_290 N_VPWR_c_410_n N_A_316_392#_c_511_n 0.00702872f $X=1.215 $Y=2.115 $X2=0
+ $Y2=0
cc_291 N_VPWR_c_410_n N_A_316_392#_c_512_n 0.0295792f $X=1.215 $Y=2.115 $X2=0
+ $Y2=0
cc_292 N_VPWR_c_411_n N_A_316_392#_c_512_n 0.0462948f $X=2.18 $Y=2.375 $X2=0
+ $Y2=0
cc_293 N_VPWR_c_412_n N_A_316_392#_c_512_n 0.0110241f $X=2.015 $Y=3.33 $X2=0
+ $Y2=0
cc_294 N_VPWR_c_406_n N_A_316_392#_c_512_n 0.00909194f $X=4.08 $Y=3.33 $X2=0
+ $Y2=0
cc_295 N_VPWR_M1006_d N_A_316_392#_c_513_n 0.00315345f $X=2.03 $Y=1.96 $X2=0
+ $Y2=0
cc_296 N_VPWR_c_411_n N_A_316_392#_c_513_n 0.0220544f $X=2.18 $Y=2.375 $X2=0
+ $Y2=0
cc_297 N_VPWR_c_411_n N_A_316_392#_c_516_n 0.00318324f $X=2.18 $Y=2.375 $X2=0
+ $Y2=0
cc_298 N_VPWR_c_411_n N_A_515_392#_c_553_n 0.038049f $X=2.18 $Y=2.375 $X2=0
+ $Y2=0
cc_299 N_VPWR_c_413_n N_A_515_392#_c_554_n 0.0582805f $X=4.08 $Y=3.33 $X2=0
+ $Y2=0
cc_300 N_VPWR_c_406_n N_A_515_392#_c_554_n 0.0326824f $X=4.08 $Y=3.33 $X2=0
+ $Y2=0
cc_301 N_VPWR_c_411_n N_A_515_392#_c_555_n 0.0139f $X=2.18 $Y=2.375 $X2=0 $Y2=0
cc_302 N_VPWR_c_413_n N_A_515_392#_c_555_n 0.0179117f $X=4.08 $Y=3.33 $X2=0
+ $Y2=0
cc_303 N_VPWR_c_406_n N_A_515_392#_c_555_n 0.00971754f $X=4.08 $Y=3.33 $X2=0
+ $Y2=0
cc_304 N_X_c_466_n N_VGND_M1001_s 9.24827e-19 $X=0.605 $Y=1.045 $X2=-0.19
+ $Y2=-0.245
cc_305 N_X_c_467_n N_VGND_M1001_s 0.00203367f $X=0.335 $Y=1.045 $X2=-0.19
+ $Y2=-0.245
cc_306 N_X_c_466_n N_VGND_c_584_n 0.00712308f $X=0.605 $Y=1.045 $X2=0 $Y2=0
cc_307 N_X_c_467_n N_VGND_c_584_n 0.0144736f $X=0.335 $Y=1.045 $X2=0 $Y2=0
cc_308 N_X_c_468_n N_VGND_c_584_n 0.0158413f $X=0.77 $Y=0.515 $X2=0 $Y2=0
cc_309 N_X_c_468_n N_VGND_c_585_n 0.0161194f $X=0.77 $Y=0.515 $X2=0 $Y2=0
cc_310 N_X_c_468_n N_VGND_c_587_n 0.0109942f $X=0.77 $Y=0.515 $X2=0 $Y2=0
cc_311 N_X_c_468_n N_VGND_c_590_n 0.00904371f $X=0.77 $Y=0.515 $X2=0 $Y2=0
cc_312 N_A_316_392#_c_515_n N_A_515_392#_M1010_s 0.00195543f $X=2.985 $Y=2.145
+ $X2=-0.19 $Y2=1.66
cc_313 N_A_316_392#_c_514_n N_A_515_392#_M1010_s 0.00462051f $X=2.635 $Y=2.035
+ $X2=-0.19 $Y2=1.66
cc_314 N_A_316_392#_c_515_n N_A_515_392#_c_553_n 0.00439071f $X=2.985 $Y=2.145
+ $X2=0 $Y2=0
cc_315 N_A_316_392#_c_514_n N_A_515_392#_c_553_n 0.0160063f $X=2.635 $Y=2.035
+ $X2=0 $Y2=0
cc_316 N_A_316_392#_c_516_n N_A_515_392#_c_553_n 0.0224621f $X=3.15 $Y=2.145
+ $X2=0 $Y2=0
cc_317 N_A_316_392#_M1010_d N_A_515_392#_c_554_n 0.00197722f $X=3 $Y=1.96 $X2=0
+ $Y2=0
cc_318 N_A_316_392#_c_515_n N_A_515_392#_c_554_n 0.00306905f $X=2.985 $Y=2.145
+ $X2=0 $Y2=0
cc_319 N_A_316_392#_c_516_n N_A_515_392#_c_554_n 0.0160685f $X=3.15 $Y=2.145
+ $X2=0 $Y2=0
cc_320 N_A_316_392#_c_516_n N_A_515_392#_c_557_n 0.0444964f $X=3.15 $Y=2.145
+ $X2=0 $Y2=0
