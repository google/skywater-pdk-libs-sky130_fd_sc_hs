* File: sky130_fd_sc_hs__fa_2.pxi.spice
* Created: Tue Sep  1 20:05:26 2020
* 
x_PM_SKY130_FD_SC_HS__FA_2%A N_A_M1017_g N_A_c_172_n N_A_M1019_g N_A_c_173_n
+ N_A_M1023_g N_A_c_174_n N_A_M1000_g N_A_c_175_n N_A_M1003_g N_A_c_176_n
+ N_A_M1015_g N_A_M1005_g N_A_c_178_n N_A_M1016_g N_A_c_179_n N_A_c_180_n
+ N_A_c_195_n N_A_c_181_n N_A_c_182_n N_A_c_183_n N_A_c_184_n N_A_c_185_n A
+ N_A_c_186_n N_A_c_187_n N_A_c_188_n PM_SKY130_FD_SC_HS__FA_2%A
x_PM_SKY130_FD_SC_HS__FA_2%CIN N_CIN_c_403_n N_CIN_M1027_g N_CIN_c_396_n
+ N_CIN_M1029_g N_CIN_c_397_n N_CIN_M1002_g N_CIN_c_398_n N_CIN_M1030_g
+ N_CIN_c_399_n N_CIN_M1024_g N_CIN_c_400_n N_CIN_M1021_g N_CIN_c_401_n
+ N_CIN_c_407_n N_CIN_c_425_n N_CIN_c_454_p N_CIN_c_408_n N_CIN_c_435_n
+ N_CIN_c_437_n N_CIN_c_409_n N_CIN_c_410_n CIN CIN N_CIN_c_402_n N_CIN_c_450_n
+ CIN CIN PM_SKY130_FD_SC_HS__FA_2%CIN
x_PM_SKY130_FD_SC_HS__FA_2%A_336_347# N_A_336_347#_M1029_d N_A_336_347#_M1027_d
+ N_A_336_347#_c_568_n N_A_336_347#_M1006_g N_A_336_347#_c_569_n
+ N_A_336_347#_M1001_g N_A_336_347#_c_570_n N_A_336_347#_M1020_g
+ N_A_336_347#_c_571_n N_A_336_347#_M1007_g N_A_336_347#_c_572_n
+ N_A_336_347#_c_573_n N_A_336_347#_c_584_n N_A_336_347#_M1031_g
+ N_A_336_347#_c_574_n N_A_336_347#_M1011_g N_A_336_347#_c_575_n
+ N_A_336_347#_c_576_n N_A_336_347#_c_598_n N_A_336_347#_c_665_p
+ N_A_336_347#_c_642_n N_A_336_347#_c_577_n N_A_336_347#_c_600_n
+ N_A_336_347#_c_578_n N_A_336_347#_c_615_n N_A_336_347#_c_579_n
+ N_A_336_347#_c_621_n N_A_336_347#_c_622_n N_A_336_347#_c_623_n
+ N_A_336_347#_c_759_p N_A_336_347#_c_580_n PM_SKY130_FD_SC_HS__FA_2%A_336_347#
x_PM_SKY130_FD_SC_HS__FA_2%B N_B_c_767_n N_B_M1008_g N_B_c_779_n N_B_c_780_n
+ N_B_c_768_n N_B_M1022_g N_B_c_783_n N_B_c_784_n N_B_c_769_n N_B_c_770_n
+ N_B_c_786_n N_B_c_787_n N_B_c_788_n N_B_M1028_g N_B_M1026_g N_B_c_790_n
+ N_B_c_771_n N_B_c_772_n N_B_c_792_n N_B_M1010_g N_B_M1014_g N_B_c_794_n
+ N_B_c_773_n N_B_c_774_n N_B_c_796_n N_B_M1012_g N_B_M1004_g N_B_c_775_n
+ N_B_c_798_n N_B_c_776_n N_B_c_799_n N_B_c_777_n N_B_c_800_n N_B_c_778_n B
+ N_B_c_802_n PM_SKY130_FD_SC_HS__FA_2%B
x_PM_SKY130_FD_SC_HS__FA_2%A_992_347# N_A_992_347#_M1001_d N_A_992_347#_M1006_d
+ N_A_992_347#_c_965_n N_A_992_347#_M1018_g N_A_992_347#_M1009_g
+ N_A_992_347#_c_967_n N_A_992_347#_c_968_n N_A_992_347#_c_976_n
+ N_A_992_347#_M1025_g N_A_992_347#_M1013_g N_A_992_347#_c_970_n
+ N_A_992_347#_c_980_n N_A_992_347#_c_984_n N_A_992_347#_c_977_n
+ N_A_992_347#_c_978_n N_A_992_347#_c_971_n N_A_992_347#_c_972_n
+ N_A_992_347#_c_973_n PM_SKY130_FD_SC_HS__FA_2%A_992_347#
x_PM_SKY130_FD_SC_HS__FA_2%A_27_378# N_A_27_378#_M1019_s N_A_27_378#_M1022_d
+ N_A_27_378#_c_1084_n N_A_27_378#_c_1092_n N_A_27_378#_c_1085_n
+ N_A_27_378#_c_1086_n PM_SKY130_FD_SC_HS__FA_2%A_27_378#
x_PM_SKY130_FD_SC_HS__FA_2%VPWR N_VPWR_M1019_d N_VPWR_M1000_d N_VPWR_M1010_d
+ N_VPWR_M1016_d N_VPWR_M1031_d N_VPWR_M1025_s N_VPWR_c_1119_n N_VPWR_c_1120_n
+ N_VPWR_c_1121_n N_VPWR_c_1122_n N_VPWR_c_1123_n N_VPWR_c_1124_n
+ N_VPWR_c_1125_n N_VPWR_c_1126_n N_VPWR_c_1127_n N_VPWR_c_1128_n VPWR
+ N_VPWR_c_1129_n N_VPWR_c_1130_n N_VPWR_c_1131_n N_VPWR_c_1132_n
+ N_VPWR_c_1133_n N_VPWR_c_1134_n N_VPWR_c_1135_n N_VPWR_c_1118_n
+ PM_SKY130_FD_SC_HS__FA_2%VPWR
x_PM_SKY130_FD_SC_HS__FA_2%A_683_347# N_A_683_347#_M1002_d N_A_683_347#_M1003_d
+ N_A_683_347#_c_1237_n N_A_683_347#_c_1238_n N_A_683_347#_c_1243_n
+ PM_SKY130_FD_SC_HS__FA_2%A_683_347#
x_PM_SKY130_FD_SC_HS__FA_2%COUT N_COUT_M1007_d N_COUT_M1020_s N_COUT_c_1280_n
+ N_COUT_c_1276_n COUT N_COUT_c_1278_n PM_SKY130_FD_SC_HS__FA_2%COUT
x_PM_SKY130_FD_SC_HS__FA_2%SUM N_SUM_M1009_d N_SUM_M1018_d N_SUM_c_1305_n
+ N_SUM_c_1306_n SUM SUM SUM SUM N_SUM_c_1307_n PM_SKY130_FD_SC_HS__FA_2%SUM
x_PM_SKY130_FD_SC_HS__FA_2%A_27_79# N_A_27_79#_M1017_s N_A_27_79#_M1008_d
+ N_A_27_79#_c_1345_n N_A_27_79#_c_1348_n N_A_27_79#_c_1346_n
+ N_A_27_79#_c_1355_n N_A_27_79#_c_1370_n N_A_27_79#_c_1356_n
+ PM_SKY130_FD_SC_HS__FA_2%A_27_79#
x_PM_SKY130_FD_SC_HS__FA_2%VGND N_VGND_M1017_d N_VGND_M1023_d N_VGND_M1014_d
+ N_VGND_M1005_d N_VGND_M1011_s N_VGND_M1013_s N_VGND_c_1381_n N_VGND_c_1382_n
+ N_VGND_c_1383_n N_VGND_c_1384_n VGND N_VGND_c_1385_n N_VGND_c_1386_n
+ N_VGND_c_1387_n N_VGND_c_1388_n N_VGND_c_1389_n N_VGND_c_1390_n
+ N_VGND_c_1391_n N_VGND_c_1392_n N_VGND_c_1393_n N_VGND_c_1394_n
+ N_VGND_c_1395_n PM_SKY130_FD_SC_HS__FA_2%VGND
x_PM_SKY130_FD_SC_HS__FA_2%A_701_79# N_A_701_79#_M1030_d N_A_701_79#_M1015_d
+ N_A_701_79#_c_1482_n N_A_701_79#_c_1485_n N_A_701_79#_c_1486_n
+ PM_SKY130_FD_SC_HS__FA_2%A_701_79#
cc_1 VNB N_A_M1017_g 0.0292213f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.765
cc_2 VNB N_A_c_172_n 0.059524f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.815
cc_3 VNB N_A_c_173_n 0.0176555f $X=-0.19 $Y=-0.245 $X2=2.75 $Y2=1.245
cc_4 VNB N_A_c_174_n 0.0221536f $X=-0.19 $Y=-0.245 $X2=2.765 $Y2=1.66
cc_5 VNB N_A_c_175_n 0.0228648f $X=-0.19 $Y=-0.245 $X2=4.435 $Y2=1.66
cc_6 VNB N_A_c_176_n 0.0192415f $X=-0.19 $Y=-0.245 $X2=4.45 $Y2=1.245
cc_7 VNB N_A_M1005_g 0.0244977f $X=-0.19 $Y=-0.245 $X2=6.34 $Y2=0.765
cc_8 VNB N_A_c_178_n 0.0260662f $X=-0.19 $Y=-0.245 $X2=6.355 $Y2=1.765
cc_9 VNB N_A_c_179_n 4.2027e-19 $X=-0.19 $Y=-0.245 $X2=2.495 $Y2=1.665
cc_10 VNB N_A_c_180_n 0.00472177f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.665
cc_11 VNB N_A_c_181_n 3.49925e-19 $X=-0.19 $Y=-0.245 $X2=2.785 $Y2=1.665
cc_12 VNB N_A_c_182_n 0.00247916f $X=-0.19 $Y=-0.245 $X2=6.335 $Y2=1.665
cc_13 VNB N_A_c_183_n 3.08548e-19 $X=-0.19 $Y=-0.245 $X2=4.225 $Y2=1.665
cc_14 VNB N_A_c_184_n 0.00715347f $X=-0.19 $Y=-0.245 $X2=4.08 $Y2=1.665
cc_15 VNB N_A_c_185_n 0.00176327f $X=-0.19 $Y=-0.245 $X2=6.48 $Y2=1.665
cc_16 VNB N_A_c_186_n 0.00357897f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.465
cc_17 VNB N_A_c_187_n 0.00546292f $X=-0.19 $Y=-0.245 $X2=2.84 $Y2=1.41
cc_18 VNB N_A_c_188_n 0.00195518f $X=-0.19 $Y=-0.245 $X2=6.43 $Y2=1.515
cc_19 VNB N_CIN_c_396_n 0.0195831f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_CIN_c_397_n 0.0256825f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.39
cc_21 VNB N_CIN_c_398_n 0.0185256f $X=-0.19 $Y=-0.245 $X2=2.75 $Y2=0.765
cc_22 VNB N_CIN_c_399_n 0.0257601f $X=-0.19 $Y=-0.245 $X2=2.765 $Y2=2.235
cc_23 VNB N_CIN_c_400_n 0.0173337f $X=-0.19 $Y=-0.245 $X2=4.435 $Y2=2.235
cc_24 VNB N_CIN_c_401_n 0.00375662f $X=-0.19 $Y=-0.245 $X2=4.45 $Y2=0.765
cc_25 VNB N_CIN_c_402_n 0.0345491f $X=-0.19 $Y=-0.245 $X2=2.84 $Y2=1.41
cc_26 VNB N_A_336_347#_c_568_n 0.0266503f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.39
cc_27 VNB N_A_336_347#_c_569_n 0.0179815f $X=-0.19 $Y=-0.245 $X2=2.75 $Y2=0.765
cc_28 VNB N_A_336_347#_c_570_n 0.030563f $X=-0.19 $Y=-0.245 $X2=2.765 $Y2=2.235
cc_29 VNB N_A_336_347#_c_571_n 0.0189208f $X=-0.19 $Y=-0.245 $X2=4.435 $Y2=2.235
cc_30 VNB N_A_336_347#_c_572_n 0.0117958f $X=-0.19 $Y=-0.245 $X2=4.45 $Y2=0.765
cc_31 VNB N_A_336_347#_c_573_n 0.0144982f $X=-0.19 $Y=-0.245 $X2=6.34 $Y2=0.765
cc_32 VNB N_A_336_347#_c_574_n 0.0184744f $X=-0.19 $Y=-0.245 $X2=6.355 $Y2=2.34
cc_33 VNB N_A_336_347#_c_575_n 0.00663775f $X=-0.19 $Y=-0.245 $X2=3.935
+ $Y2=1.665
cc_34 VNB N_A_336_347#_c_576_n 0.00414225f $X=-0.19 $Y=-0.245 $X2=6.335
+ $Y2=1.665
cc_35 VNB N_A_336_347#_c_577_n 0.00299485f $X=-0.19 $Y=-0.245 $X2=4.08 $Y2=1.665
cc_36 VNB N_A_336_347#_c_578_n 0.00120782f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_336_347#_c_579_n 0.0025057f $X=-0.19 $Y=-0.245 $X2=2.84 $Y2=1.41
cc_38 VNB N_A_336_347#_c_580_n 0.00656164f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_B_c_767_n 0.020601f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.3
cc_40 VNB N_B_c_768_n 0.028145f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.39
cc_41 VNB N_B_c_769_n 0.00567192f $X=-0.19 $Y=-0.245 $X2=2.765 $Y2=2.235
cc_42 VNB N_B_c_770_n 0.0134072f $X=-0.19 $Y=-0.245 $X2=2.765 $Y2=2.235
cc_43 VNB N_B_c_771_n 0.00588435f $X=-0.19 $Y=-0.245 $X2=6.355 $Y2=2.34
cc_44 VNB N_B_c_772_n 0.0135891f $X=-0.19 $Y=-0.245 $X2=6.355 $Y2=2.34
cc_45 VNB N_B_c_773_n 0.00559958f $X=-0.19 $Y=-0.245 $X2=4.08 $Y2=1.665
cc_46 VNB N_B_c_774_n 0.0161788f $X=-0.19 $Y=-0.245 $X2=4.08 $Y2=1.665
cc_47 VNB N_B_c_775_n 0.0150758f $X=-0.19 $Y=-0.245 $X2=0.35 $Y2=1.465
cc_48 VNB N_B_c_776_n 0.0158954f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.465
cc_49 VNB N_B_c_777_n 0.0146896f $X=-0.19 $Y=-0.245 $X2=2.84 $Y2=1.41
cc_50 VNB N_B_c_778_n 0.00380736f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_A_992_347#_c_965_n 0.0328658f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.39
cc_52 VNB N_A_992_347#_M1009_g 0.0226186f $X=-0.19 $Y=-0.245 $X2=2.765 $Y2=2.235
cc_53 VNB N_A_992_347#_c_967_n 0.0135027f $X=-0.19 $Y=-0.245 $X2=4.435 $Y2=1.66
cc_54 VNB N_A_992_347#_c_968_n 0.0149496f $X=-0.19 $Y=-0.245 $X2=4.45 $Y2=1.245
cc_55 VNB N_A_992_347#_M1013_g 0.0244428f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_A_992_347#_c_970_n 0.0111562f $X=-0.19 $Y=-0.245 $X2=6.355 $Y2=2.34
cc_57 VNB N_A_992_347#_c_971_n 0.00296222f $X=-0.19 $Y=-0.245 $X2=6.48 $Y2=1.665
cc_58 VNB N_A_992_347#_c_972_n 0.00607642f $X=-0.19 $Y=-0.245 $X2=0.35 $Y2=1.465
cc_59 VNB N_A_992_347#_c_973_n 0.0029615f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.465
cc_60 VNB N_VPWR_c_1118_n 0.382608f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_COUT_c_1276_n 0.00105681f $X=-0.19 $Y=-0.245 $X2=2.765 $Y2=2.235
cc_62 VNB N_SUM_c_1305_n 0.00250577f $X=-0.19 $Y=-0.245 $X2=2.75 $Y2=0.765
cc_63 VNB N_SUM_c_1306_n 0.00176823f $X=-0.19 $Y=-0.245 $X2=2.765 $Y2=2.235
cc_64 VNB N_SUM_c_1307_n 0.0020572f $X=-0.19 $Y=-0.245 $X2=4.225 $Y2=1.665
cc_65 VNB N_A_27_79#_c_1345_n 0.022885f $X=-0.19 $Y=-0.245 $X2=2.75 $Y2=0.765
cc_66 VNB N_A_27_79#_c_1346_n 0.00924515f $X=-0.19 $Y=-0.245 $X2=2.765 $Y2=2.235
cc_67 VNB N_VGND_c_1381_n 0.0107925f $X=-0.19 $Y=-0.245 $X2=6.34 $Y2=0.765
cc_68 VNB N_VGND_c_1382_n 0.0103473f $X=-0.19 $Y=-0.245 $X2=6.355 $Y2=2.34
cc_69 VNB N_VGND_c_1383_n 0.010678f $X=-0.19 $Y=-0.245 $X2=2.495 $Y2=1.665
cc_70 VNB N_VGND_c_1384_n 0.0467943f $X=-0.19 $Y=-0.245 $X2=3.935 $Y2=1.665
cc_71 VNB N_VGND_c_1385_n 0.0192741f $X=-0.19 $Y=-0.245 $X2=2.64 $Y2=1.665
cc_72 VNB N_VGND_c_1386_n 0.0538033f $X=-0.19 $Y=-0.245 $X2=4.08 $Y2=1.665
cc_73 VNB N_VGND_c_1387_n 0.0182626f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.465
cc_74 VNB N_VGND_c_1388_n 0.0758158f $X=-0.19 $Y=-0.245 $X2=4.36 $Y2=1.41
cc_75 VNB N_VGND_c_1389_n 0.0185038f $X=-0.19 $Y=-0.245 $X2=6.43 $Y2=1.515
cc_76 VNB N_VGND_c_1390_n 0.0194856f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.665
cc_77 VNB N_VGND_c_1391_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=2.64 $Y2=1.665
cc_78 VNB N_VGND_c_1392_n 0.00980973f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.665
cc_79 VNB N_VGND_c_1393_n 0.0158564f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_VGND_c_1394_n 0.0187415f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_81 VNB N_VGND_c_1395_n 0.522665f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_82 VNB N_A_701_79#_c_1482_n 0.00247806f $X=-0.19 $Y=-0.245 $X2=2.75 $Y2=0.765
cc_83 VPB N_A_c_172_n 0.0340295f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.815
cc_84 VPB N_A_c_174_n 0.0234011f $X=-0.19 $Y=1.66 $X2=2.765 $Y2=1.66
cc_85 VPB N_A_c_175_n 0.0248746f $X=-0.19 $Y=1.66 $X2=4.435 $Y2=1.66
cc_86 VPB N_A_c_178_n 0.0264704f $X=-0.19 $Y=1.66 $X2=6.355 $Y2=1.765
cc_87 VPB N_A_c_179_n 0.011005f $X=-0.19 $Y=1.66 $X2=2.495 $Y2=1.665
cc_88 VPB N_A_c_180_n 0.00683299f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.665
cc_89 VPB N_A_c_195_n 0.00671911f $X=-0.19 $Y=1.66 $X2=3.935 $Y2=1.665
cc_90 VPB N_A_c_181_n 3.31226e-19 $X=-0.19 $Y=1.66 $X2=2.785 $Y2=1.665
cc_91 VPB N_A_c_182_n 0.0126049f $X=-0.19 $Y=1.66 $X2=6.335 $Y2=1.665
cc_92 VPB N_A_c_183_n 0.0014314f $X=-0.19 $Y=1.66 $X2=4.225 $Y2=1.665
cc_93 VPB N_A_c_184_n 0.00579748f $X=-0.19 $Y=1.66 $X2=4.08 $Y2=1.665
cc_94 VPB N_A_c_185_n 0.00408517f $X=-0.19 $Y=1.66 $X2=6.48 $Y2=1.665
cc_95 VPB N_A_c_186_n 0.00277085f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.465
cc_96 VPB N_A_c_187_n 0.00253327f $X=-0.19 $Y=1.66 $X2=2.84 $Y2=1.41
cc_97 VPB N_A_c_188_n 0.00301871f $X=-0.19 $Y=1.66 $X2=6.43 $Y2=1.515
cc_98 VPB N_CIN_c_403_n 0.0147098f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.3
cc_99 VPB N_CIN_c_397_n 0.0251531f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.39
cc_100 VPB N_CIN_c_399_n 0.0248361f $X=-0.19 $Y=1.66 $X2=2.765 $Y2=2.235
cc_101 VPB N_CIN_c_401_n 2.09458e-19 $X=-0.19 $Y=1.66 $X2=4.45 $Y2=0.765
cc_102 VPB N_CIN_c_407_n 0.00218398f $X=-0.19 $Y=1.66 $X2=6.355 $Y2=2.34
cc_103 VPB N_CIN_c_408_n 0.00112438f $X=-0.19 $Y=1.66 $X2=3.935 $Y2=1.665
cc_104 VPB N_CIN_c_409_n 0.00242029f $X=-0.19 $Y=1.66 $X2=2.64 $Y2=1.665
cc_105 VPB N_CIN_c_410_n 2.62341e-19 $X=-0.19 $Y=1.66 $X2=4.08 $Y2=1.665
cc_106 VPB N_CIN_c_402_n 0.0179496f $X=-0.19 $Y=1.66 $X2=2.84 $Y2=1.41
cc_107 VPB N_A_336_347#_c_568_n 0.024396f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.39
cc_108 VPB N_A_336_347#_c_570_n 0.0252407f $X=-0.19 $Y=1.66 $X2=2.765 $Y2=2.235
cc_109 VPB N_A_336_347#_c_573_n 9.27735e-19 $X=-0.19 $Y=1.66 $X2=6.34 $Y2=0.765
cc_110 VPB N_A_336_347#_c_584_n 0.0233394f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_111 VPB N_A_336_347#_c_576_n 0.00145942f $X=-0.19 $Y=1.66 $X2=6.335 $Y2=1.665
cc_112 VPB N_A_336_347#_c_578_n 0.0010773f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_113 VPB N_B_c_779_n 0.00749723f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_114 VPB N_B_c_780_n 0.015767f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.815
cc_115 VPB N_B_c_768_n 0.0155687f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.39
cc_116 VPB N_B_M1022_g 0.00818226f $X=-0.19 $Y=1.66 $X2=2.75 $Y2=0.765
cc_117 VPB N_B_c_783_n 0.071366f $X=-0.19 $Y=1.66 $X2=2.75 $Y2=0.765
cc_118 VPB N_B_c_784_n 0.0139987f $X=-0.19 $Y=1.66 $X2=2.765 $Y2=1.66
cc_119 VPB N_B_c_770_n 7.3898e-19 $X=-0.19 $Y=1.66 $X2=2.765 $Y2=2.235
cc_120 VPB N_B_c_786_n 0.00796806f $X=-0.19 $Y=1.66 $X2=4.435 $Y2=1.66
cc_121 VPB N_B_c_787_n 0.0161956f $X=-0.19 $Y=1.66 $X2=4.435 $Y2=2.235
cc_122 VPB N_B_c_788_n 0.00604263f $X=-0.19 $Y=1.66 $X2=4.435 $Y2=2.235
cc_123 VPB N_B_M1028_g 0.00858468f $X=-0.19 $Y=1.66 $X2=4.45 $Y2=0.765
cc_124 VPB N_B_c_790_n 0.103205f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_125 VPB N_B_c_772_n 0.00904024f $X=-0.19 $Y=1.66 $X2=6.355 $Y2=2.34
cc_126 VPB N_B_c_792_n 0.00621372f $X=-0.19 $Y=1.66 $X2=2.495 $Y2=1.665
cc_127 VPB N_B_M1010_g 0.0101067f $X=-0.19 $Y=1.66 $X2=2.785 $Y2=1.665
cc_128 VPB N_B_c_794_n 0.14108f $X=-0.19 $Y=1.66 $X2=2.64 $Y2=1.665
cc_129 VPB N_B_c_774_n 0.00331323f $X=-0.19 $Y=1.66 $X2=4.08 $Y2=1.665
cc_130 VPB N_B_c_796_n 0.00570017f $X=-0.19 $Y=1.66 $X2=4.08 $Y2=1.665
cc_131 VPB N_B_M1012_g 0.00969195f $X=-0.19 $Y=1.66 $X2=6.48 $Y2=1.665
cc_132 VPB N_B_c_798_n 0.0089864f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.465
cc_133 VPB N_B_c_799_n 0.018297f $X=-0.19 $Y=1.66 $X2=2.84 $Y2=1.41
cc_134 VPB N_B_c_800_n 0.0297235f $X=-0.19 $Y=1.66 $X2=4.36 $Y2=1.41
cc_135 VPB N_B_c_778_n 4.92487e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_136 VPB N_B_c_802_n 0.00455707f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_137 VPB N_A_992_347#_c_965_n 0.024762f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.39
cc_138 VPB N_A_992_347#_c_968_n 0.00111912f $X=-0.19 $Y=1.66 $X2=4.45 $Y2=1.245
cc_139 VPB N_A_992_347#_c_976_n 0.0258095f $X=-0.19 $Y=1.66 $X2=4.45 $Y2=0.765
cc_140 VPB N_A_992_347#_c_977_n 0.00290363f $X=-0.19 $Y=1.66 $X2=2.64 $Y2=1.665
cc_141 VPB N_A_992_347#_c_978_n 0.00275916f $X=-0.19 $Y=1.66 $X2=2.64 $Y2=1.665
cc_142 VPB N_A_27_378#_c_1084_n 0.0145709f $X=-0.19 $Y=1.66 $X2=2.75 $Y2=0.765
cc_143 VPB N_A_27_378#_c_1085_n 0.0268148f $X=-0.19 $Y=1.66 $X2=4.435 $Y2=2.235
cc_144 VPB N_A_27_378#_c_1086_n 0.00279333f $X=-0.19 $Y=1.66 $X2=4.45 $Y2=0.765
cc_145 VPB N_VPWR_c_1119_n 0.0164359f $X=-0.19 $Y=1.66 $X2=6.34 $Y2=0.765
cc_146 VPB N_VPWR_c_1120_n 0.00837087f $X=-0.19 $Y=1.66 $X2=6.355 $Y2=2.34
cc_147 VPB N_VPWR_c_1121_n 0.00984397f $X=-0.19 $Y=1.66 $X2=3.935 $Y2=1.665
cc_148 VPB N_VPWR_c_1122_n 0.00788352f $X=-0.19 $Y=1.66 $X2=2.64 $Y2=1.665
cc_149 VPB N_VPWR_c_1123_n 0.0108116f $X=-0.19 $Y=1.66 $X2=2.64 $Y2=1.665
cc_150 VPB N_VPWR_c_1124_n 0.0588404f $X=-0.19 $Y=1.66 $X2=4.08 $Y2=1.665
cc_151 VPB N_VPWR_c_1125_n 0.0532034f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_152 VPB N_VPWR_c_1126_n 0.00436868f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_153 VPB N_VPWR_c_1127_n 0.0670335f $X=-0.19 $Y=1.66 $X2=0.35 $Y2=1.465
cc_154 VPB N_VPWR_c_1128_n 0.00614127f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.465
cc_155 VPB N_VPWR_c_1129_n 0.0193443f $X=-0.19 $Y=1.66 $X2=2.84 $Y2=1.41
cc_156 VPB N_VPWR_c_1130_n 0.0200644f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=1.665
cc_157 VPB N_VPWR_c_1131_n 0.0208129f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_158 VPB N_VPWR_c_1132_n 0.019486f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_159 VPB N_VPWR_c_1133_n 0.00757184f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_160 VPB N_VPWR_c_1134_n 0.00510111f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_161 VPB N_VPWR_c_1135_n 0.0178563f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_162 VPB N_VPWR_c_1118_n 0.0700796f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_163 VPB N_A_683_347#_c_1237_n 7.25211e-19 $X=-0.19 $Y=1.66 $X2=2.75 $Y2=0.765
cc_164 VPB N_A_683_347#_c_1238_n 0.00242661f $X=-0.19 $Y=1.66 $X2=4.435
+ $Y2=2.235
cc_165 VPB N_COUT_c_1276_n 0.00128407f $X=-0.19 $Y=1.66 $X2=2.765 $Y2=2.235
cc_166 VPB N_COUT_c_1278_n 0.00392752f $X=-0.19 $Y=1.66 $X2=4.435 $Y2=2.235
cc_167 VPB SUM 0.00164137f $X=-0.19 $Y=1.66 $X2=4.435 $Y2=1.66
cc_168 VPB SUM 0.00257348f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_169 VPB N_SUM_c_1307_n 8.45676e-19 $X=-0.19 $Y=1.66 $X2=4.225 $Y2=1.665
cc_170 N_A_c_179_n N_CIN_c_403_n 0.00201489f $X=2.495 $Y=1.665 $X2=-0.19
+ $Y2=-0.245
cc_171 N_A_c_174_n N_CIN_c_397_n 0.0498297f $X=2.765 $Y=1.66 $X2=0 $Y2=0
cc_172 N_A_c_195_n N_CIN_c_397_n 0.00344172f $X=3.935 $Y=1.665 $X2=0 $Y2=0
cc_173 N_A_c_181_n N_CIN_c_397_n 3.14434e-19 $X=2.785 $Y=1.665 $X2=0 $Y2=0
cc_174 N_A_c_187_n N_CIN_c_397_n 0.00181833f $X=2.84 $Y=1.41 $X2=0 $Y2=0
cc_175 N_A_c_173_n N_CIN_c_398_n 0.0198817f $X=2.75 $Y=1.245 $X2=0 $Y2=0
cc_176 N_A_c_182_n N_CIN_c_399_n 4.95816e-19 $X=6.335 $Y=1.665 $X2=0 $Y2=0
cc_177 N_A_c_179_n N_CIN_c_401_n 0.014025f $X=2.495 $Y=1.665 $X2=0 $Y2=0
cc_178 N_A_c_181_n N_CIN_c_401_n 7.08402e-19 $X=2.785 $Y=1.665 $X2=0 $Y2=0
cc_179 N_A_c_187_n N_CIN_c_401_n 0.0183851f $X=2.84 $Y=1.41 $X2=0 $Y2=0
cc_180 N_A_c_179_n N_CIN_c_407_n 0.0151462f $X=2.495 $Y=1.665 $X2=0 $Y2=0
cc_181 N_A_c_181_n N_CIN_c_407_n 0.00177234f $X=2.785 $Y=1.665 $X2=0 $Y2=0
cc_182 N_A_c_187_n N_CIN_c_407_n 0.0072747f $X=2.84 $Y=1.41 $X2=0 $Y2=0
cc_183 N_A_c_174_n N_CIN_c_425_n 0.0164464f $X=2.765 $Y=1.66 $X2=0 $Y2=0
cc_184 N_A_c_179_n N_CIN_c_425_n 0.0105527f $X=2.495 $Y=1.665 $X2=0 $Y2=0
cc_185 N_A_c_195_n N_CIN_c_425_n 0.0185306f $X=3.935 $Y=1.665 $X2=0 $Y2=0
cc_186 N_A_c_181_n N_CIN_c_425_n 0.00393208f $X=2.785 $Y=1.665 $X2=0 $Y2=0
cc_187 N_A_c_187_n N_CIN_c_425_n 0.0165874f $X=2.84 $Y=1.41 $X2=0 $Y2=0
cc_188 N_A_c_174_n N_CIN_c_408_n 0.00134925f $X=2.765 $Y=1.66 $X2=0 $Y2=0
cc_189 N_A_c_195_n N_CIN_c_408_n 0.0155819f $X=3.935 $Y=1.665 $X2=0 $Y2=0
cc_190 N_A_c_181_n N_CIN_c_408_n 0.00111887f $X=2.785 $Y=1.665 $X2=0 $Y2=0
cc_191 N_A_c_183_n N_CIN_c_408_n 0.00117756f $X=4.225 $Y=1.665 $X2=0 $Y2=0
cc_192 N_A_c_187_n N_CIN_c_408_n 0.0021498f $X=2.84 $Y=1.41 $X2=0 $Y2=0
cc_193 N_A_c_182_n N_CIN_c_435_n 0.0264144f $X=6.335 $Y=1.665 $X2=0 $Y2=0
cc_194 N_A_c_188_n N_CIN_c_435_n 0.00108359f $X=6.43 $Y=1.515 $X2=0 $Y2=0
cc_195 N_A_c_175_n N_CIN_c_437_n 0.0199556f $X=4.435 $Y=1.66 $X2=0 $Y2=0
cc_196 N_A_c_182_n N_CIN_c_437_n 0.00847825f $X=6.335 $Y=1.665 $X2=0 $Y2=0
cc_197 N_A_c_183_n N_CIN_c_437_n 0.00533814f $X=4.225 $Y=1.665 $X2=0 $Y2=0
cc_198 N_A_c_184_n N_CIN_c_437_n 0.0206888f $X=4.08 $Y=1.665 $X2=0 $Y2=0
cc_199 N_A_c_182_n N_CIN_c_409_n 0.0245402f $X=6.335 $Y=1.665 $X2=0 $Y2=0
cc_200 N_A_c_188_n N_CIN_c_409_n 0.00832169f $X=6.43 $Y=1.515 $X2=0 $Y2=0
cc_201 N_A_c_174_n N_CIN_c_410_n 3.97873e-19 $X=2.765 $Y=1.66 $X2=0 $Y2=0
cc_202 N_A_c_195_n N_CIN_c_410_n 0.00490934f $X=3.935 $Y=1.665 $X2=0 $Y2=0
cc_203 N_A_c_183_n N_CIN_c_410_n 9.52871e-19 $X=4.225 $Y=1.665 $X2=0 $Y2=0
cc_204 N_A_c_184_n N_CIN_c_410_n 0.0180651f $X=4.08 $Y=1.665 $X2=0 $Y2=0
cc_205 N_A_c_187_n N_CIN_c_410_n 0.0205242f $X=2.84 $Y=1.41 $X2=0 $Y2=0
cc_206 N_A_c_174_n CIN 2.08429e-19 $X=2.765 $Y=1.66 $X2=0 $Y2=0
cc_207 N_A_c_179_n N_CIN_c_402_n 0.0126f $X=2.495 $Y=1.665 $X2=0 $Y2=0
cc_208 N_A_c_195_n N_CIN_c_450_n 0.0163301f $X=3.935 $Y=1.665 $X2=0 $Y2=0
cc_209 N_A_c_183_n N_CIN_c_450_n 0.00493529f $X=4.225 $Y=1.665 $X2=0 $Y2=0
cc_210 N_A_c_184_n N_CIN_c_450_n 0.00787124f $X=4.08 $Y=1.665 $X2=0 $Y2=0
cc_211 N_A_c_179_n N_A_336_347#_M1027_d 0.00395264f $X=2.495 $Y=1.665 $X2=0
+ $Y2=0
cc_212 N_A_c_175_n N_A_336_347#_c_568_n 0.0558089f $X=4.435 $Y=1.66 $X2=0 $Y2=0
cc_213 N_A_c_182_n N_A_336_347#_c_568_n 0.00583338f $X=6.335 $Y=1.665 $X2=0
+ $Y2=0
cc_214 N_A_c_184_n N_A_336_347#_c_568_n 0.00115874f $X=4.08 $Y=1.665 $X2=0 $Y2=0
cc_215 N_A_c_176_n N_A_336_347#_c_569_n 0.0270001f $X=4.45 $Y=1.245 $X2=0 $Y2=0
cc_216 N_A_M1005_g N_A_336_347#_c_570_n 0.00229568f $X=6.34 $Y=0.765 $X2=0 $Y2=0
cc_217 N_A_c_178_n N_A_336_347#_c_570_n 0.0497937f $X=6.355 $Y=1.765 $X2=0 $Y2=0
cc_218 N_A_c_185_n N_A_336_347#_c_570_n 0.00354858f $X=6.48 $Y=1.665 $X2=0 $Y2=0
cc_219 N_A_c_188_n N_A_336_347#_c_570_n 0.00305605f $X=6.43 $Y=1.515 $X2=0 $Y2=0
cc_220 N_A_M1005_g N_A_336_347#_c_571_n 0.0178654f $X=6.34 $Y=0.765 $X2=0 $Y2=0
cc_221 N_A_c_179_n N_A_336_347#_c_576_n 0.0193041f $X=2.495 $Y=1.665 $X2=0 $Y2=0
cc_222 N_A_c_179_n N_A_336_347#_c_598_n 0.003536f $X=2.495 $Y=1.665 $X2=0 $Y2=0
cc_223 N_A_c_173_n N_A_336_347#_c_577_n 0.00199687f $X=2.75 $Y=1.245 $X2=0 $Y2=0
cc_224 N_A_c_173_n N_A_336_347#_c_600_n 0.0149278f $X=2.75 $Y=1.245 $X2=0 $Y2=0
cc_225 N_A_c_174_n N_A_336_347#_c_600_n 0.00405354f $X=2.765 $Y=1.66 $X2=0 $Y2=0
cc_226 N_A_c_175_n N_A_336_347#_c_600_n 0.00405354f $X=4.435 $Y=1.66 $X2=0 $Y2=0
cc_227 N_A_c_176_n N_A_336_347#_c_600_n 0.0118522f $X=4.45 $Y=1.245 $X2=0 $Y2=0
cc_228 N_A_c_179_n N_A_336_347#_c_600_n 0.00521189f $X=2.495 $Y=1.665 $X2=0
+ $Y2=0
cc_229 N_A_c_195_n N_A_336_347#_c_600_n 0.0199166f $X=3.935 $Y=1.665 $X2=0 $Y2=0
cc_230 N_A_c_181_n N_A_336_347#_c_600_n 0.00210494f $X=2.785 $Y=1.665 $X2=0
+ $Y2=0
cc_231 N_A_c_182_n N_A_336_347#_c_600_n 0.00561366f $X=6.335 $Y=1.665 $X2=0
+ $Y2=0
cc_232 N_A_c_183_n N_A_336_347#_c_600_n 0.00214331f $X=4.225 $Y=1.665 $X2=0
+ $Y2=0
cc_233 N_A_c_184_n N_A_336_347#_c_600_n 0.0383589f $X=4.08 $Y=1.665 $X2=0 $Y2=0
cc_234 N_A_c_187_n N_A_336_347#_c_600_n 0.0313356f $X=2.84 $Y=1.41 $X2=0 $Y2=0
cc_235 N_A_c_175_n N_A_336_347#_c_578_n 5.07555e-19 $X=4.435 $Y=1.66 $X2=0 $Y2=0
cc_236 N_A_c_176_n N_A_336_347#_c_578_n 0.0035272f $X=4.45 $Y=1.245 $X2=0 $Y2=0
cc_237 N_A_c_182_n N_A_336_347#_c_578_n 0.00935813f $X=6.335 $Y=1.665 $X2=0
+ $Y2=0
cc_238 N_A_c_184_n N_A_336_347#_c_578_n 0.0186719f $X=4.08 $Y=1.665 $X2=0 $Y2=0
cc_239 N_A_M1005_g N_A_336_347#_c_615_n 0.0117248f $X=6.34 $Y=0.765 $X2=0 $Y2=0
cc_240 N_A_c_178_n N_A_336_347#_c_615_n 9.98306e-19 $X=6.355 $Y=1.765 $X2=0
+ $Y2=0
cc_241 N_A_c_182_n N_A_336_347#_c_615_n 0.0257369f $X=6.335 $Y=1.665 $X2=0 $Y2=0
cc_242 N_A_c_185_n N_A_336_347#_c_615_n 0.00233398f $X=6.48 $Y=1.665 $X2=0 $Y2=0
cc_243 N_A_c_188_n N_A_336_347#_c_615_n 0.0147348f $X=6.43 $Y=1.515 $X2=0 $Y2=0
cc_244 N_A_M1005_g N_A_336_347#_c_579_n 0.00307272f $X=6.34 $Y=0.765 $X2=0 $Y2=0
cc_245 N_A_c_179_n N_A_336_347#_c_621_n 0.015434f $X=2.495 $Y=1.665 $X2=0 $Y2=0
cc_246 N_A_c_179_n N_A_336_347#_c_622_n 0.00625275f $X=2.495 $Y=1.665 $X2=0
+ $Y2=0
cc_247 N_A_c_179_n N_A_336_347#_c_623_n 0.00387496f $X=2.495 $Y=1.665 $X2=0
+ $Y2=0
cc_248 N_A_M1005_g N_A_336_347#_c_580_n 0.00196053f $X=6.34 $Y=0.765 $X2=0 $Y2=0
cc_249 N_A_c_178_n N_A_336_347#_c_580_n 0.00140769f $X=6.355 $Y=1.765 $X2=0
+ $Y2=0
cc_250 N_A_c_185_n N_A_336_347#_c_580_n 0.00102585f $X=6.48 $Y=1.665 $X2=0 $Y2=0
cc_251 N_A_c_188_n N_A_336_347#_c_580_n 0.0184416f $X=6.43 $Y=1.515 $X2=0 $Y2=0
cc_252 N_A_M1017_g N_B_c_767_n 0.0191562f $X=0.495 $Y=0.765 $X2=-0.19 $Y2=-0.245
cc_253 N_A_c_172_n N_B_c_779_n 0.00319861f $X=0.505 $Y=1.815 $X2=0 $Y2=0
cc_254 N_A_M1017_g N_B_c_768_n 0.0108341f $X=0.495 $Y=0.765 $X2=0 $Y2=0
cc_255 N_A_c_172_n N_B_c_768_n 0.00726414f $X=0.505 $Y=1.815 $X2=0 $Y2=0
cc_256 N_A_c_179_n N_B_c_768_n 0.0100044f $X=2.495 $Y=1.665 $X2=0 $Y2=0
cc_257 N_A_c_186_n N_B_c_768_n 2.17233e-19 $X=0.27 $Y=1.465 $X2=0 $Y2=0
cc_258 N_A_c_172_n N_B_M1022_g 0.0206901f $X=0.505 $Y=1.815 $X2=0 $Y2=0
cc_259 N_A_c_179_n N_B_M1022_g 0.00381423f $X=2.495 $Y=1.665 $X2=0 $Y2=0
cc_260 N_A_c_187_n N_B_c_769_n 0.00337199f $X=2.84 $Y=1.41 $X2=0 $Y2=0
cc_261 N_A_c_174_n N_B_c_770_n 0.0365084f $X=2.765 $Y=1.66 $X2=0 $Y2=0
cc_262 N_A_c_181_n N_B_c_770_n 7.31736e-19 $X=2.785 $Y=1.665 $X2=0 $Y2=0
cc_263 N_A_c_174_n N_B_c_786_n 0.00280186f $X=2.765 $Y=1.66 $X2=0 $Y2=0
cc_264 N_A_c_179_n N_B_c_788_n 0.00397396f $X=2.495 $Y=1.665 $X2=0 $Y2=0
cc_265 N_A_c_174_n N_B_M1028_g 0.0539834f $X=2.765 $Y=1.66 $X2=0 $Y2=0
cc_266 N_A_c_179_n N_B_M1028_g 0.00297635f $X=2.495 $Y=1.665 $X2=0 $Y2=0
cc_267 N_A_c_181_n N_B_M1028_g 7.31127e-19 $X=2.785 $Y=1.665 $X2=0 $Y2=0
cc_268 N_A_c_187_n N_B_M1028_g 8.20424e-19 $X=2.84 $Y=1.41 $X2=0 $Y2=0
cc_269 N_A_c_174_n N_B_c_790_n 0.0103562f $X=2.765 $Y=1.66 $X2=0 $Y2=0
cc_270 N_A_c_175_n N_B_c_771_n 0.015159f $X=4.435 $Y=1.66 $X2=0 $Y2=0
cc_271 N_A_c_184_n N_B_c_771_n 0.00612966f $X=4.08 $Y=1.665 $X2=0 $Y2=0
cc_272 N_A_c_175_n N_B_c_772_n 0.00718841f $X=4.435 $Y=1.66 $X2=0 $Y2=0
cc_273 N_A_c_195_n N_B_c_772_n 0.00392216f $X=3.935 $Y=1.665 $X2=0 $Y2=0
cc_274 N_A_c_183_n N_B_c_772_n 0.00191165f $X=4.225 $Y=1.665 $X2=0 $Y2=0
cc_275 N_A_c_195_n N_B_c_792_n 0.00174117f $X=3.935 $Y=1.665 $X2=0 $Y2=0
cc_276 N_A_c_183_n N_B_c_792_n 9.266e-19 $X=4.225 $Y=1.665 $X2=0 $Y2=0
cc_277 N_A_c_175_n N_B_M1010_g 0.0225413f $X=4.435 $Y=1.66 $X2=0 $Y2=0
cc_278 N_A_c_175_n N_B_c_794_n 0.0100145f $X=4.435 $Y=1.66 $X2=0 $Y2=0
cc_279 N_A_c_178_n N_B_c_774_n 0.0421668f $X=6.355 $Y=1.765 $X2=0 $Y2=0
cc_280 N_A_c_182_n N_B_c_774_n 0.00405176f $X=6.335 $Y=1.665 $X2=0 $Y2=0
cc_281 N_A_c_188_n N_B_c_774_n 0.00184828f $X=6.43 $Y=1.515 $X2=0 $Y2=0
cc_282 N_A_c_182_n N_B_c_796_n 0.00385187f $X=6.335 $Y=1.665 $X2=0 $Y2=0
cc_283 N_A_c_178_n N_B_M1012_g 0.0578524f $X=6.355 $Y=1.765 $X2=0 $Y2=0
cc_284 N_A_c_173_n N_B_c_775_n 0.0365084f $X=2.75 $Y=1.245 $X2=0 $Y2=0
cc_285 N_A_c_176_n N_B_c_776_n 0.0257242f $X=4.45 $Y=1.245 $X2=0 $Y2=0
cc_286 N_A_M1005_g N_B_c_777_n 0.0421668f $X=6.34 $Y=0.765 $X2=0 $Y2=0
cc_287 N_A_c_178_n N_B_c_800_n 0.00286536f $X=6.355 $Y=1.765 $X2=0 $Y2=0
cc_288 N_A_M1017_g N_B_c_778_n 0.00313715f $X=0.495 $Y=0.765 $X2=0 $Y2=0
cc_289 N_A_c_172_n N_B_c_778_n 8.64873e-19 $X=0.505 $Y=1.815 $X2=0 $Y2=0
cc_290 N_A_c_179_n N_B_c_778_n 0.0201027f $X=2.495 $Y=1.665 $X2=0 $Y2=0
cc_291 N_A_c_186_n N_B_c_778_n 0.017755f $X=0.27 $Y=1.465 $X2=0 $Y2=0
cc_292 N_A_c_179_n B 0.0027266f $X=2.495 $Y=1.665 $X2=0 $Y2=0
cc_293 N_A_c_172_n N_B_c_802_n 0.00549019f $X=0.505 $Y=1.815 $X2=0 $Y2=0
cc_294 N_A_c_179_n N_B_c_802_n 0.0125264f $X=2.495 $Y=1.665 $X2=0 $Y2=0
cc_295 N_A_c_180_n N_B_c_802_n 4.21253e-19 $X=0.385 $Y=1.665 $X2=0 $Y2=0
cc_296 N_A_c_186_n N_B_c_802_n 0.0103537f $X=0.27 $Y=1.465 $X2=0 $Y2=0
cc_297 N_A_c_182_n N_A_992_347#_M1006_d 0.00245688f $X=6.335 $Y=1.665 $X2=0
+ $Y2=0
cc_298 N_A_c_178_n N_A_992_347#_c_980_n 0.0146767f $X=6.355 $Y=1.765 $X2=0 $Y2=0
cc_299 N_A_c_182_n N_A_992_347#_c_980_n 0.0200918f $X=6.335 $Y=1.665 $X2=0 $Y2=0
cc_300 N_A_c_185_n N_A_992_347#_c_980_n 0.00261606f $X=6.48 $Y=1.665 $X2=0 $Y2=0
cc_301 N_A_c_188_n N_A_992_347#_c_980_n 0.0055978f $X=6.43 $Y=1.515 $X2=0 $Y2=0
cc_302 N_A_M1005_g N_A_992_347#_c_984_n 0.0121667f $X=6.34 $Y=0.765 $X2=0 $Y2=0
cc_303 N_A_c_179_n N_A_27_378#_M1022_d 0.00143238f $X=2.495 $Y=1.665 $X2=0 $Y2=0
cc_304 N_A_c_172_n N_A_27_378#_c_1084_n 0.00161023f $X=0.505 $Y=1.815 $X2=0
+ $Y2=0
cc_305 N_A_c_179_n N_A_27_378#_c_1084_n 2.96655e-19 $X=2.495 $Y=1.665 $X2=0
+ $Y2=0
cc_306 N_A_c_180_n N_A_27_378#_c_1084_n 0.00294111f $X=0.385 $Y=1.665 $X2=0
+ $Y2=0
cc_307 N_A_c_186_n N_A_27_378#_c_1084_n 0.0218249f $X=0.27 $Y=1.465 $X2=0 $Y2=0
cc_308 N_A_c_172_n N_A_27_378#_c_1092_n 0.0113294f $X=0.505 $Y=1.815 $X2=0 $Y2=0
cc_309 N_A_c_179_n N_A_27_378#_c_1092_n 0.0154426f $X=2.495 $Y=1.665 $X2=0 $Y2=0
cc_310 N_A_c_172_n N_A_27_378#_c_1085_n 0.00702625f $X=0.505 $Y=1.815 $X2=0
+ $Y2=0
cc_311 N_A_c_179_n N_A_27_378#_c_1085_n 3.53264e-19 $X=2.495 $Y=1.665 $X2=0
+ $Y2=0
cc_312 N_A_c_172_n N_A_27_378#_c_1086_n 0.00158491f $X=0.505 $Y=1.815 $X2=0
+ $Y2=0
cc_313 N_A_c_179_n N_A_27_378#_c_1086_n 0.0068788f $X=2.495 $Y=1.665 $X2=0 $Y2=0
cc_314 N_A_c_179_n N_VPWR_M1019_d 0.00317318f $X=2.495 $Y=1.665 $X2=-0.19
+ $Y2=-0.245
cc_315 N_A_c_195_n N_VPWR_M1000_d 0.00352864f $X=3.935 $Y=1.665 $X2=0 $Y2=0
cc_316 N_A_c_182_n N_VPWR_M1010_d 0.00109217f $X=6.335 $Y=1.665 $X2=0 $Y2=0
cc_317 N_A_c_183_n N_VPWR_M1010_d 0.00151528f $X=4.225 $Y=1.665 $X2=0 $Y2=0
cc_318 N_A_c_184_n N_VPWR_M1010_d 7.7392e-19 $X=4.08 $Y=1.665 $X2=0 $Y2=0
cc_319 N_A_c_172_n N_VPWR_c_1119_n 0.00528244f $X=0.505 $Y=1.815 $X2=0 $Y2=0
cc_320 N_A_c_174_n N_VPWR_c_1120_n 0.0135439f $X=2.765 $Y=1.66 $X2=0 $Y2=0
cc_321 N_A_c_175_n N_VPWR_c_1121_n 0.00418101f $X=4.435 $Y=1.66 $X2=0 $Y2=0
cc_322 N_A_c_178_n N_VPWR_c_1122_n 0.00839052f $X=6.355 $Y=1.765 $X2=0 $Y2=0
cc_323 N_A_c_178_n N_VPWR_c_1127_n 0.0049405f $X=6.355 $Y=1.765 $X2=0 $Y2=0
cc_324 N_A_c_172_n N_VPWR_c_1129_n 0.00513952f $X=0.505 $Y=1.815 $X2=0 $Y2=0
cc_325 N_A_c_172_n N_VPWR_c_1118_n 0.00523671f $X=0.505 $Y=1.815 $X2=0 $Y2=0
cc_326 N_A_c_174_n N_VPWR_c_1118_n 8.51577e-19 $X=2.765 $Y=1.66 $X2=0 $Y2=0
cc_327 N_A_c_175_n N_VPWR_c_1118_n 9.39239e-19 $X=4.435 $Y=1.66 $X2=0 $Y2=0
cc_328 N_A_c_178_n N_VPWR_c_1118_n 0.00508379f $X=6.355 $Y=1.765 $X2=0 $Y2=0
cc_329 N_A_c_179_n A_484_347# 6.14399e-19 $X=2.495 $Y=1.665 $X2=-0.19 $Y2=-0.245
cc_330 N_A_c_181_n A_484_347# 0.00157018f $X=2.785 $Y=1.665 $X2=-0.19 $Y2=-0.245
cc_331 N_A_c_187_n A_484_347# 8.66022e-19 $X=2.84 $Y=1.41 $X2=-0.19 $Y2=-0.245
cc_332 N_A_c_195_n N_A_683_347#_M1002_d 0.00110158f $X=3.935 $Y=1.665 $X2=-0.19
+ $Y2=-0.245
cc_333 N_A_c_182_n N_A_683_347#_M1003_d 0.00214261f $X=6.335 $Y=1.665 $X2=0
+ $Y2=0
cc_334 N_A_c_195_n N_A_683_347#_c_1237_n 8.4709e-19 $X=3.935 $Y=1.665 $X2=0
+ $Y2=0
cc_335 N_A_c_175_n N_A_683_347#_c_1238_n 0.00737612f $X=4.435 $Y=1.66 $X2=0
+ $Y2=0
cc_336 N_A_c_175_n N_A_683_347#_c_1243_n 0.00827287f $X=4.435 $Y=1.66 $X2=0
+ $Y2=0
cc_337 N_A_c_182_n A_1094_347# 0.00130281f $X=6.335 $Y=1.665 $X2=-0.19
+ $Y2=-0.245
cc_338 N_A_c_178_n N_COUT_c_1278_n 0.00146531f $X=6.355 $Y=1.765 $X2=0 $Y2=0
cc_339 N_A_M1017_g N_A_27_79#_c_1345_n 0.00837143f $X=0.495 $Y=0.765 $X2=0 $Y2=0
cc_340 N_A_M1017_g N_A_27_79#_c_1348_n 0.0129862f $X=0.495 $Y=0.765 $X2=0 $Y2=0
cc_341 N_A_c_179_n N_A_27_79#_c_1348_n 0.00766083f $X=2.495 $Y=1.665 $X2=0 $Y2=0
cc_342 N_A_M1017_g N_A_27_79#_c_1346_n 0.0020332f $X=0.495 $Y=0.765 $X2=0 $Y2=0
cc_343 N_A_c_172_n N_A_27_79#_c_1346_n 0.00224099f $X=0.505 $Y=1.815 $X2=0 $Y2=0
cc_344 N_A_c_179_n N_A_27_79#_c_1346_n 5.71069e-19 $X=2.495 $Y=1.665 $X2=0 $Y2=0
cc_345 N_A_c_180_n N_A_27_79#_c_1346_n 0.0013364f $X=0.385 $Y=1.665 $X2=0 $Y2=0
cc_346 N_A_c_186_n N_A_27_79#_c_1346_n 0.0235003f $X=0.27 $Y=1.465 $X2=0 $Y2=0
cc_347 N_A_M1017_g N_VGND_c_1381_n 0.00570879f $X=0.495 $Y=0.765 $X2=0 $Y2=0
cc_348 N_A_c_173_n N_VGND_c_1382_n 0.0160326f $X=2.75 $Y=1.245 $X2=0 $Y2=0
cc_349 N_A_M1017_g N_VGND_c_1385_n 0.00534051f $X=0.495 $Y=0.765 $X2=0 $Y2=0
cc_350 N_A_c_173_n N_VGND_c_1386_n 0.00465077f $X=2.75 $Y=1.245 $X2=0 $Y2=0
cc_351 N_A_c_176_n N_VGND_c_1388_n 0.00420132f $X=4.45 $Y=1.245 $X2=0 $Y2=0
cc_352 N_A_M1005_g N_VGND_c_1388_n 0.00846197f $X=6.34 $Y=0.765 $X2=0 $Y2=0
cc_353 N_A_c_176_n N_VGND_c_1393_n 0.00385053f $X=4.45 $Y=1.245 $X2=0 $Y2=0
cc_354 N_A_M1017_g N_VGND_c_1395_n 0.00537853f $X=0.495 $Y=0.765 $X2=0 $Y2=0
cc_355 N_A_c_173_n N_VGND_c_1395_n 0.00451796f $X=2.75 $Y=1.245 $X2=0 $Y2=0
cc_356 N_A_c_176_n N_VGND_c_1395_n 0.00537853f $X=4.45 $Y=1.245 $X2=0 $Y2=0
cc_357 N_A_M1005_g N_VGND_c_1395_n 0.00537853f $X=6.34 $Y=0.765 $X2=0 $Y2=0
cc_358 N_A_c_173_n N_A_701_79#_c_1482_n 3.90878e-19 $X=2.75 $Y=1.245 $X2=0 $Y2=0
cc_359 N_A_c_176_n N_A_701_79#_c_1482_n 8.56546e-19 $X=4.45 $Y=1.245 $X2=0 $Y2=0
cc_360 N_A_c_176_n N_A_701_79#_c_1485_n 0.00968656f $X=4.45 $Y=1.245 $X2=0 $Y2=0
cc_361 N_A_c_176_n N_A_701_79#_c_1486_n 0.00878341f $X=4.45 $Y=1.245 $X2=0 $Y2=0
cc_362 N_CIN_c_407_n N_A_336_347#_M1027_d 0.00245536f $X=2.14 $Y=1.95 $X2=0
+ $Y2=0
cc_363 N_CIN_c_454_p N_A_336_347#_M1027_d 0.0046269f $X=2.225 $Y=2.035 $X2=0
+ $Y2=0
cc_364 N_CIN_c_399_n N_A_336_347#_c_568_n 0.0501918f $X=5.395 $Y=1.66 $X2=0
+ $Y2=0
cc_365 N_CIN_c_435_n N_A_336_347#_c_568_n 0.015789f $X=5.305 $Y=1.83 $X2=0 $Y2=0
cc_366 N_CIN_c_409_n N_A_336_347#_c_568_n 0.0028202f $X=5.47 $Y=1.41 $X2=0 $Y2=0
cc_367 N_CIN_c_400_n N_A_336_347#_c_569_n 0.0277034f $X=5.52 $Y=1.245 $X2=0
+ $Y2=0
cc_368 N_CIN_c_403_n N_A_336_347#_c_576_n 0.00179211f $X=1.605 $Y=1.66 $X2=0
+ $Y2=0
cc_369 N_CIN_c_396_n N_A_336_347#_c_576_n 0.00330402f $X=1.86 $Y=1.245 $X2=0
+ $Y2=0
cc_370 N_CIN_c_401_n N_A_336_347#_c_576_n 0.0232781f $X=2.055 $Y=1.417 $X2=0
+ $Y2=0
cc_371 N_CIN_c_407_n N_A_336_347#_c_576_n 0.00347803f $X=2.14 $Y=1.95 $X2=0
+ $Y2=0
cc_372 N_CIN_c_402_n N_A_336_347#_c_576_n 0.0110899f $X=1.86 $Y=1.452 $X2=0
+ $Y2=0
cc_373 N_CIN_c_396_n N_A_336_347#_c_598_n 0.0152984f $X=1.86 $Y=1.245 $X2=0
+ $Y2=0
cc_374 N_CIN_c_401_n N_A_336_347#_c_598_n 0.0150423f $X=2.055 $Y=1.417 $X2=0
+ $Y2=0
cc_375 N_CIN_c_402_n N_A_336_347#_c_598_n 0.00673579f $X=1.86 $Y=1.452 $X2=0
+ $Y2=0
cc_376 N_CIN_c_407_n N_A_336_347#_c_642_n 0.00250584f $X=2.14 $Y=1.95 $X2=0
+ $Y2=0
cc_377 N_CIN_c_454_p N_A_336_347#_c_642_n 0.0138309f $X=2.225 $Y=2.035 $X2=0
+ $Y2=0
cc_378 N_CIN_c_396_n N_A_336_347#_c_577_n 0.00328097f $X=1.86 $Y=1.245 $X2=0
+ $Y2=0
cc_379 N_CIN_c_397_n N_A_336_347#_c_600_n 0.003457f $X=3.34 $Y=1.66 $X2=0 $Y2=0
cc_380 N_CIN_c_398_n N_A_336_347#_c_600_n 0.0151375f $X=3.43 $Y=1.245 $X2=0
+ $Y2=0
cc_381 N_CIN_c_435_n N_A_336_347#_c_600_n 0.00199472f $X=5.305 $Y=1.83 $X2=0
+ $Y2=0
cc_382 N_CIN_c_410_n N_A_336_347#_c_600_n 0.020621f $X=3.38 $Y=1.41 $X2=0 $Y2=0
cc_383 N_CIN_c_399_n N_A_336_347#_c_578_n 0.00120415f $X=5.395 $Y=1.66 $X2=0
+ $Y2=0
cc_384 N_CIN_c_400_n N_A_336_347#_c_578_n 9.1313e-19 $X=5.52 $Y=1.245 $X2=0
+ $Y2=0
cc_385 N_CIN_c_435_n N_A_336_347#_c_578_n 0.0168115f $X=5.305 $Y=1.83 $X2=0
+ $Y2=0
cc_386 N_CIN_c_409_n N_A_336_347#_c_578_n 0.0199626f $X=5.47 $Y=1.41 $X2=0 $Y2=0
cc_387 N_CIN_c_399_n N_A_336_347#_c_615_n 0.00359716f $X=5.395 $Y=1.66 $X2=0
+ $Y2=0
cc_388 N_CIN_c_400_n N_A_336_347#_c_615_n 0.0107724f $X=5.52 $Y=1.245 $X2=0
+ $Y2=0
cc_389 N_CIN_c_435_n N_A_336_347#_c_615_n 0.00172633f $X=5.305 $Y=1.83 $X2=0
+ $Y2=0
cc_390 N_CIN_c_409_n N_A_336_347#_c_615_n 0.0212826f $X=5.47 $Y=1.41 $X2=0 $Y2=0
cc_391 N_CIN_c_403_n N_A_336_347#_c_621_n 0.0152599f $X=1.605 $Y=1.66 $X2=0
+ $Y2=0
cc_392 N_CIN_c_401_n N_A_336_347#_c_621_n 0.0090667f $X=2.055 $Y=1.417 $X2=0
+ $Y2=0
cc_393 N_CIN_c_407_n N_A_336_347#_c_621_n 0.0132855f $X=2.14 $Y=1.95 $X2=0 $Y2=0
cc_394 N_CIN_c_402_n N_A_336_347#_c_621_n 0.00456175f $X=1.86 $Y=1.452 $X2=0
+ $Y2=0
cc_395 N_CIN_c_454_p N_A_336_347#_c_622_n 0.0107286f $X=2.225 $Y=2.035 $X2=0
+ $Y2=0
cc_396 N_CIN_c_401_n N_A_336_347#_c_623_n 0.020623f $X=2.055 $Y=1.417 $X2=0
+ $Y2=0
cc_397 N_CIN_c_402_n N_A_336_347#_c_623_n 0.00150385f $X=1.86 $Y=1.452 $X2=0
+ $Y2=0
cc_398 N_CIN_c_396_n N_B_c_767_n 0.01693f $X=1.86 $Y=1.245 $X2=-0.19 $Y2=-0.245
cc_399 N_CIN_c_403_n N_B_c_779_n 0.00255705f $X=1.605 $Y=1.66 $X2=0 $Y2=0
cc_400 N_CIN_c_402_n N_B_c_768_n 0.0169239f $X=1.86 $Y=1.452 $X2=0 $Y2=0
cc_401 N_CIN_c_403_n N_B_M1022_g 0.018678f $X=1.605 $Y=1.66 $X2=0 $Y2=0
cc_402 N_CIN_c_403_n N_B_c_783_n 0.0103487f $X=1.605 $Y=1.66 $X2=0 $Y2=0
cc_403 N_CIN_c_396_n N_B_c_769_n 0.00157551f $X=1.86 $Y=1.245 $X2=0 $Y2=0
cc_404 N_CIN_c_401_n N_B_c_769_n 0.00308749f $X=2.055 $Y=1.417 $X2=0 $Y2=0
cc_405 N_CIN_c_402_n N_B_c_769_n 0.0197345f $X=1.86 $Y=1.452 $X2=0 $Y2=0
cc_406 N_CIN_c_403_n N_B_c_786_n 0.0014644f $X=1.605 $Y=1.66 $X2=0 $Y2=0
cc_407 N_CIN_c_407_n N_B_c_788_n 9.85867e-19 $X=2.14 $Y=1.95 $X2=0 $Y2=0
cc_408 N_CIN_c_402_n N_B_c_788_n 0.00166586f $X=1.86 $Y=1.452 $X2=0 $Y2=0
cc_409 N_CIN_c_403_n N_B_M1028_g 0.0167295f $X=1.605 $Y=1.66 $X2=0 $Y2=0
cc_410 N_CIN_c_407_n N_B_M1028_g 0.00251859f $X=2.14 $Y=1.95 $X2=0 $Y2=0
cc_411 N_CIN_c_425_n N_B_M1028_g 0.0157453f $X=3.375 $Y=2.035 $X2=0 $Y2=0
cc_412 N_CIN_c_397_n N_B_c_790_n 0.0103728f $X=3.34 $Y=1.66 $X2=0 $Y2=0
cc_413 N_CIN_c_397_n N_B_c_771_n 0.0201396f $X=3.34 $Y=1.66 $X2=0 $Y2=0
cc_414 N_CIN_c_398_n N_B_c_771_n 0.00196948f $X=3.43 $Y=1.245 $X2=0 $Y2=0
cc_415 N_CIN_c_410_n N_B_c_771_n 0.00114716f $X=3.38 $Y=1.41 $X2=0 $Y2=0
cc_416 N_CIN_c_397_n N_B_c_772_n 0.00861901f $X=3.34 $Y=1.66 $X2=0 $Y2=0
cc_417 N_CIN_c_408_n N_B_c_772_n 0.00231522f $X=3.46 $Y=1.935 $X2=0 $Y2=0
cc_418 N_CIN_c_437_n N_B_c_792_n 2.72709e-19 $X=4.535 $Y=1.83 $X2=0 $Y2=0
cc_419 N_CIN_c_397_n N_B_M1010_g 0.0276136f $X=3.34 $Y=1.66 $X2=0 $Y2=0
cc_420 N_CIN_c_408_n N_B_M1010_g 0.00238604f $X=3.46 $Y=1.935 $X2=0 $Y2=0
cc_421 N_CIN_c_437_n N_B_M1010_g 6.5829e-19 $X=4.535 $Y=1.83 $X2=0 $Y2=0
cc_422 N_CIN_c_450_n N_B_M1010_g 0.01389f $X=4.088 $Y=2.042 $X2=0 $Y2=0
cc_423 N_CIN_c_399_n N_B_c_794_n 0.0100192f $X=5.395 $Y=1.66 $X2=0 $Y2=0
cc_424 N_CIN_c_399_n N_B_c_773_n 0.0209564f $X=5.395 $Y=1.66 $X2=0 $Y2=0
cc_425 N_CIN_c_400_n N_B_c_773_n 0.00196948f $X=5.52 $Y=1.245 $X2=0 $Y2=0
cc_426 N_CIN_c_409_n N_B_c_773_n 0.00153135f $X=5.47 $Y=1.41 $X2=0 $Y2=0
cc_427 N_CIN_c_399_n N_B_c_774_n 0.00617896f $X=5.395 $Y=1.66 $X2=0 $Y2=0
cc_428 N_CIN_c_409_n N_B_c_774_n 0.00150368f $X=5.47 $Y=1.41 $X2=0 $Y2=0
cc_429 N_CIN_c_435_n N_B_c_796_n 2.59657e-19 $X=5.305 $Y=1.83 $X2=0 $Y2=0
cc_430 N_CIN_c_399_n N_B_M1012_g 0.035569f $X=5.395 $Y=1.66 $X2=0 $Y2=0
cc_431 N_CIN_c_435_n N_B_M1012_g 0.00380739f $X=5.305 $Y=1.83 $X2=0 $Y2=0
cc_432 N_CIN_c_396_n N_B_c_775_n 0.018948f $X=1.86 $Y=1.245 $X2=0 $Y2=0
cc_433 N_CIN_c_398_n N_B_c_776_n 0.027619f $X=3.43 $Y=1.245 $X2=0 $Y2=0
cc_434 N_CIN_c_400_n N_B_c_777_n 0.0449656f $X=5.52 $Y=1.245 $X2=0 $Y2=0
cc_435 N_CIN_c_402_n N_B_c_778_n 3.09561e-19 $X=1.86 $Y=1.452 $X2=0 $Y2=0
cc_436 N_CIN_c_435_n N_A_992_347#_M1006_d 0.00592499f $X=5.305 $Y=1.83 $X2=0
+ $Y2=0
cc_437 N_CIN_c_399_n N_A_992_347#_c_980_n 0.0094745f $X=5.395 $Y=1.66 $X2=0
+ $Y2=0
cc_438 N_CIN_c_435_n N_A_992_347#_c_980_n 0.0084263f $X=5.305 $Y=1.83 $X2=0
+ $Y2=0
cc_439 N_CIN_c_400_n N_A_992_347#_c_984_n 0.0085641f $X=5.52 $Y=1.245 $X2=0
+ $Y2=0
cc_440 N_CIN_c_399_n N_A_992_347#_c_978_n 0.0109992f $X=5.395 $Y=1.66 $X2=0
+ $Y2=0
cc_441 N_CIN_c_435_n N_A_992_347#_c_978_n 0.0197772f $X=5.305 $Y=1.83 $X2=0
+ $Y2=0
cc_442 N_CIN_c_400_n N_A_992_347#_c_971_n 0.00545857f $X=5.52 $Y=1.245 $X2=0
+ $Y2=0
cc_443 N_CIN_c_403_n N_A_27_378#_c_1086_n 0.011693f $X=1.605 $Y=1.66 $X2=0 $Y2=0
cc_444 N_CIN_c_425_n N_VPWR_M1000_d 0.0093626f $X=3.375 $Y=2.035 $X2=0 $Y2=0
cc_445 N_CIN_c_437_n N_VPWR_M1010_d 0.00619008f $X=4.535 $Y=1.83 $X2=0 $Y2=0
cc_446 N_CIN_c_450_n N_VPWR_M1010_d 0.0022456f $X=4.088 $Y=2.042 $X2=0 $Y2=0
cc_447 N_CIN_c_397_n N_VPWR_c_1120_n 0.00789792f $X=3.34 $Y=1.66 $X2=0 $Y2=0
cc_448 N_CIN_c_425_n N_VPWR_c_1120_n 0.0212438f $X=3.375 $Y=2.035 $X2=0 $Y2=0
cc_449 N_CIN_c_397_n N_VPWR_c_1121_n 5.6418e-19 $X=3.34 $Y=1.66 $X2=0 $Y2=0
cc_450 N_CIN_c_403_n N_VPWR_c_1118_n 9.39239e-19 $X=1.605 $Y=1.66 $X2=0 $Y2=0
cc_451 N_CIN_c_397_n N_VPWR_c_1118_n 9.39239e-19 $X=3.34 $Y=1.66 $X2=0 $Y2=0
cc_452 N_CIN_c_399_n N_VPWR_c_1118_n 9.39239e-19 $X=5.395 $Y=1.66 $X2=0 $Y2=0
cc_453 N_CIN_c_425_n A_484_347# 0.00762779f $X=3.375 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_454 N_CIN_c_408_n N_A_683_347#_M1002_d 0.00227812f $X=3.46 $Y=1.935 $X2=-0.19
+ $Y2=-0.245
cc_455 CIN N_A_683_347#_M1002_d 7.96769e-19 $X=3.515 $Y=1.95 $X2=-0.19
+ $Y2=-0.245
cc_456 N_CIN_c_450_n N_A_683_347#_M1002_d 0.00408291f $X=4.088 $Y=2.042
+ $X2=-0.19 $Y2=-0.245
cc_457 N_CIN_c_435_n N_A_683_347#_M1003_d 0.00586137f $X=5.305 $Y=1.83 $X2=0
+ $Y2=0
cc_458 N_CIN_c_397_n N_A_683_347#_c_1237_n 0.00603929f $X=3.34 $Y=1.66 $X2=0
+ $Y2=0
cc_459 CIN N_A_683_347#_c_1237_n 0.00685294f $X=3.515 $Y=1.95 $X2=0 $Y2=0
cc_460 N_CIN_c_450_n N_A_683_347#_c_1237_n 0.013007f $X=4.088 $Y=2.042 $X2=0
+ $Y2=0
cc_461 N_CIN_c_435_n N_A_683_347#_c_1238_n 0.00773289f $X=5.305 $Y=1.83 $X2=0
+ $Y2=0
cc_462 N_CIN_c_437_n N_A_683_347#_c_1238_n 0.0010989f $X=4.535 $Y=1.83 $X2=0
+ $Y2=0
cc_463 N_CIN_c_437_n N_A_683_347#_c_1243_n 0.0216917f $X=4.535 $Y=1.83 $X2=0
+ $Y2=0
cc_464 N_CIN_c_450_n N_A_683_347#_c_1243_n 0.0180141f $X=4.088 $Y=2.042 $X2=0
+ $Y2=0
cc_465 N_CIN_c_435_n A_1094_347# 0.00427113f $X=5.305 $Y=1.83 $X2=-0.19
+ $Y2=-0.245
cc_466 N_CIN_c_396_n N_A_27_79#_c_1355_n 7.78141e-19 $X=1.86 $Y=1.245 $X2=0
+ $Y2=0
cc_467 N_CIN_c_396_n N_A_27_79#_c_1356_n 0.0102445f $X=1.86 $Y=1.245 $X2=0 $Y2=0
cc_468 N_CIN_c_402_n N_A_27_79#_c_1356_n 3.81313e-19 $X=1.86 $Y=1.452 $X2=0
+ $Y2=0
cc_469 N_CIN_c_398_n N_VGND_c_1382_n 0.00610458f $X=3.43 $Y=1.245 $X2=0 $Y2=0
cc_470 N_CIN_c_396_n N_VGND_c_1386_n 0.00533923f $X=1.86 $Y=1.245 $X2=0 $Y2=0
cc_471 N_CIN_c_398_n N_VGND_c_1387_n 0.00534051f $X=3.43 $Y=1.245 $X2=0 $Y2=0
cc_472 N_CIN_c_400_n N_VGND_c_1388_n 0.00419817f $X=5.52 $Y=1.245 $X2=0 $Y2=0
cc_473 N_CIN_c_396_n N_VGND_c_1395_n 0.00537853f $X=1.86 $Y=1.245 $X2=0 $Y2=0
cc_474 N_CIN_c_398_n N_VGND_c_1395_n 0.00537853f $X=3.43 $Y=1.245 $X2=0 $Y2=0
cc_475 N_CIN_c_400_n N_VGND_c_1395_n 0.00537853f $X=5.52 $Y=1.245 $X2=0 $Y2=0
cc_476 N_CIN_c_398_n N_A_701_79#_c_1482_n 0.00523166f $X=3.43 $Y=1.245 $X2=0
+ $Y2=0
cc_477 N_A_336_347#_c_576_n N_B_c_767_n 0.00605652f $X=1.46 $Y=1.745 $X2=-0.19
+ $Y2=-0.245
cc_478 N_A_336_347#_c_665_p N_B_c_767_n 0.00190527f $X=1.545 $Y=1.005 $X2=-0.19
+ $Y2=-0.245
cc_479 N_A_336_347#_c_576_n N_B_c_768_n 0.00141938f $X=1.46 $Y=1.745 $X2=0 $Y2=0
cc_480 N_A_336_347#_c_621_n N_B_M1022_g 0.0019933f $X=1.8 $Y=1.83 $X2=0 $Y2=0
cc_481 N_A_336_347#_c_622_n N_B_c_783_n 0.00768137f $X=2 $Y=2.455 $X2=0 $Y2=0
cc_482 N_A_336_347#_c_642_n N_B_M1028_g 0.00353603f $X=1.8 $Y=2.29 $X2=0 $Y2=0
cc_483 N_A_336_347#_c_622_n N_B_M1028_g 0.00576159f $X=2 $Y=2.455 $X2=0 $Y2=0
cc_484 N_A_336_347#_c_568_n N_B_c_794_n 0.010344f $X=4.885 $Y=1.66 $X2=0 $Y2=0
cc_485 N_A_336_347#_c_577_n N_B_c_775_n 0.00973989f $X=2.145 $Y=0.54 $X2=0 $Y2=0
cc_486 N_A_336_347#_c_600_n N_B_c_775_n 0.0117189f $X=4.765 $Y=1.005 $X2=0 $Y2=0
cc_487 N_A_336_347#_c_623_n N_B_c_775_n 9.8677e-19 $X=2.145 $Y=1.005 $X2=0 $Y2=0
cc_488 N_A_336_347#_c_600_n N_B_c_776_n 0.0124386f $X=4.765 $Y=1.005 $X2=0 $Y2=0
cc_489 N_A_336_347#_c_615_n N_B_c_777_n 0.0114492f $X=6.765 $Y=1.005 $X2=0 $Y2=0
cc_490 N_A_336_347#_c_576_n N_B_c_778_n 0.0218014f $X=1.46 $Y=1.745 $X2=0 $Y2=0
cc_491 N_A_336_347#_c_576_n N_B_c_802_n 0.0037895f $X=1.46 $Y=1.745 $X2=0 $Y2=0
cc_492 N_A_336_347#_c_621_n N_B_c_802_n 0.00561757f $X=1.8 $Y=1.83 $X2=0 $Y2=0
cc_493 N_A_336_347#_c_615_n N_A_992_347#_M1001_d 0.00615946f $X=6.765 $Y=1.005
+ $X2=-0.19 $Y2=-0.245
cc_494 N_A_336_347#_c_573_n N_A_992_347#_c_965_n 0.00175884f $X=7.47 $Y=1.675
+ $X2=0 $Y2=0
cc_495 N_A_336_347#_c_584_n N_A_992_347#_c_965_n 0.0213307f $X=7.47 $Y=1.765
+ $X2=0 $Y2=0
cc_496 N_A_336_347#_c_575_n N_A_992_347#_c_965_n 0.010916f $X=7.47 $Y=1.33 $X2=0
+ $Y2=0
cc_497 N_A_336_347#_c_574_n N_A_992_347#_M1009_g 0.0153227f $X=7.485 $Y=1.255
+ $X2=0 $Y2=0
cc_498 N_A_336_347#_c_570_n N_A_992_347#_c_980_n 0.0171525f $X=6.925 $Y=1.765
+ $X2=0 $Y2=0
cc_499 N_A_336_347#_c_584_n N_A_992_347#_c_980_n 0.0133594f $X=7.47 $Y=1.765
+ $X2=0 $Y2=0
cc_500 N_A_336_347#_c_570_n N_A_992_347#_c_984_n 3.23175e-19 $X=6.925 $Y=1.765
+ $X2=0 $Y2=0
cc_501 N_A_336_347#_c_571_n N_A_992_347#_c_984_n 0.0138642f $X=7.055 $Y=1.255
+ $X2=0 $Y2=0
cc_502 N_A_336_347#_c_574_n N_A_992_347#_c_984_n 0.0124144f $X=7.485 $Y=1.255
+ $X2=0 $Y2=0
cc_503 N_A_336_347#_c_615_n N_A_992_347#_c_984_n 0.081584f $X=6.765 $Y=1.005
+ $X2=0 $Y2=0
cc_504 N_A_336_347#_c_580_n N_A_992_347#_c_984_n 0.00436361f $X=7 $Y=1.42 $X2=0
+ $Y2=0
cc_505 N_A_336_347#_c_573_n N_A_992_347#_c_977_n 0.00320155f $X=7.47 $Y=1.675
+ $X2=0 $Y2=0
cc_506 N_A_336_347#_c_584_n N_A_992_347#_c_977_n 0.00468564f $X=7.47 $Y=1.765
+ $X2=0 $Y2=0
cc_507 N_A_336_347#_c_568_n N_A_992_347#_c_978_n 0.00366284f $X=4.885 $Y=1.66
+ $X2=0 $Y2=0
cc_508 N_A_336_347#_c_569_n N_A_992_347#_c_971_n 0.00239476f $X=5.02 $Y=1.245
+ $X2=0 $Y2=0
cc_509 N_A_336_347#_c_615_n N_A_992_347#_c_971_n 0.0200079f $X=6.765 $Y=1.005
+ $X2=0 $Y2=0
cc_510 N_A_336_347#_c_575_n N_A_992_347#_c_972_n 0.00320155f $X=7.47 $Y=1.33
+ $X2=0 $Y2=0
cc_511 N_A_336_347#_c_574_n N_A_992_347#_c_973_n 0.00320155f $X=7.485 $Y=1.255
+ $X2=0 $Y2=0
cc_512 N_A_336_347#_c_576_n N_A_27_378#_M1022_d 4.21214e-19 $X=1.46 $Y=1.745
+ $X2=0 $Y2=0
cc_513 N_A_336_347#_c_621_n N_A_27_378#_M1022_d 0.00363686f $X=1.8 $Y=1.83 $X2=0
+ $Y2=0
cc_514 N_A_336_347#_c_621_n N_A_27_378#_c_1086_n 0.00837331f $X=1.8 $Y=1.83
+ $X2=0 $Y2=0
cc_515 N_A_336_347#_c_622_n N_VPWR_c_1120_n 0.00916814f $X=2 $Y=2.455 $X2=0
+ $Y2=0
cc_516 N_A_336_347#_c_570_n N_VPWR_c_1122_n 0.0113821f $X=6.925 $Y=1.765 $X2=0
+ $Y2=0
cc_517 N_A_336_347#_c_584_n N_VPWR_c_1122_n 0.00142599f $X=7.47 $Y=1.765 $X2=0
+ $Y2=0
cc_518 N_A_336_347#_c_622_n N_VPWR_c_1125_n 0.00716517f $X=2 $Y=2.455 $X2=0
+ $Y2=0
cc_519 N_A_336_347#_c_570_n N_VPWR_c_1131_n 0.00413917f $X=6.925 $Y=1.765 $X2=0
+ $Y2=0
cc_520 N_A_336_347#_c_584_n N_VPWR_c_1131_n 0.00415318f $X=7.47 $Y=1.765 $X2=0
+ $Y2=0
cc_521 N_A_336_347#_c_570_n N_VPWR_c_1135_n 0.00110534f $X=6.925 $Y=1.765 $X2=0
+ $Y2=0
cc_522 N_A_336_347#_c_584_n N_VPWR_c_1135_n 0.0138746f $X=7.47 $Y=1.765 $X2=0
+ $Y2=0
cc_523 N_A_336_347#_c_568_n N_VPWR_c_1118_n 9.39239e-19 $X=4.885 $Y=1.66 $X2=0
+ $Y2=0
cc_524 N_A_336_347#_c_570_n N_VPWR_c_1118_n 0.00415345f $X=6.925 $Y=1.765 $X2=0
+ $Y2=0
cc_525 N_A_336_347#_c_584_n N_VPWR_c_1118_n 0.00415345f $X=7.47 $Y=1.765 $X2=0
+ $Y2=0
cc_526 N_A_336_347#_c_622_n N_VPWR_c_1118_n 0.0112052f $X=2 $Y=2.455 $X2=0 $Y2=0
cc_527 N_A_336_347#_c_568_n N_A_683_347#_c_1238_n 0.00665871f $X=4.885 $Y=1.66
+ $X2=0 $Y2=0
cc_528 N_A_336_347#_c_571_n N_COUT_c_1280_n 0.002376f $X=7.055 $Y=1.255 $X2=0
+ $Y2=0
cc_529 N_A_336_347#_c_572_n N_COUT_c_1280_n 0.00342367f $X=7.38 $Y=1.33 $X2=0
+ $Y2=0
cc_530 N_A_336_347#_c_574_n N_COUT_c_1280_n 0.00581486f $X=7.485 $Y=1.255 $X2=0
+ $Y2=0
cc_531 N_A_336_347#_c_580_n N_COUT_c_1280_n 0.00306471f $X=7 $Y=1.42 $X2=0 $Y2=0
cc_532 N_A_336_347#_c_570_n N_COUT_c_1276_n 0.00221371f $X=6.925 $Y=1.765 $X2=0
+ $Y2=0
cc_533 N_A_336_347#_c_571_n N_COUT_c_1276_n 8.6474e-19 $X=7.055 $Y=1.255 $X2=0
+ $Y2=0
cc_534 N_A_336_347#_c_573_n N_COUT_c_1276_n 0.00862707f $X=7.47 $Y=1.675 $X2=0
+ $Y2=0
cc_535 N_A_336_347#_c_584_n N_COUT_c_1276_n 0.0198732f $X=7.47 $Y=1.765 $X2=0
+ $Y2=0
cc_536 N_A_336_347#_c_574_n N_COUT_c_1276_n 0.00414001f $X=7.485 $Y=1.255 $X2=0
+ $Y2=0
cc_537 N_A_336_347#_c_575_n N_COUT_c_1276_n 0.00594554f $X=7.47 $Y=1.33 $X2=0
+ $Y2=0
cc_538 N_A_336_347#_c_579_n N_COUT_c_1276_n 0.00454656f $X=6.85 $Y=1.255 $X2=0
+ $Y2=0
cc_539 N_A_336_347#_c_580_n N_COUT_c_1276_n 0.0194098f $X=7 $Y=1.42 $X2=0 $Y2=0
cc_540 N_A_336_347#_c_570_n N_COUT_c_1278_n 0.0118952f $X=6.925 $Y=1.765 $X2=0
+ $Y2=0
cc_541 N_A_336_347#_c_572_n N_COUT_c_1278_n 0.00676361f $X=7.38 $Y=1.33 $X2=0
+ $Y2=0
cc_542 N_A_336_347#_c_584_n N_COUT_c_1278_n 2.28571e-19 $X=7.47 $Y=1.765 $X2=0
+ $Y2=0
cc_543 N_A_336_347#_c_580_n N_COUT_c_1278_n 0.011125f $X=7 $Y=1.42 $X2=0 $Y2=0
cc_544 N_A_336_347#_c_574_n N_SUM_c_1305_n 8.94563e-19 $X=7.485 $Y=1.255 $X2=0
+ $Y2=0
cc_545 N_A_336_347#_c_584_n SUM 0.00128072f $X=7.47 $Y=1.765 $X2=0 $Y2=0
cc_546 N_A_336_347#_c_576_n N_A_27_79#_M1008_d 0.00104465f $X=1.46 $Y=1.745
+ $X2=0 $Y2=0
cc_547 N_A_336_347#_c_598_n N_A_27_79#_M1008_d 0.00469593f $X=1.98 $Y=1.005
+ $X2=0 $Y2=0
cc_548 N_A_336_347#_c_665_p N_A_27_79#_M1008_d 0.00471217f $X=1.545 $Y=1.005
+ $X2=0 $Y2=0
cc_549 N_A_336_347#_c_665_p N_A_27_79#_c_1348_n 0.0135477f $X=1.545 $Y=1.005
+ $X2=0 $Y2=0
cc_550 N_A_336_347#_c_598_n N_A_27_79#_c_1356_n 0.0157342f $X=1.98 $Y=1.005
+ $X2=0 $Y2=0
cc_551 N_A_336_347#_c_665_p N_A_27_79#_c_1356_n 0.0144778f $X=1.545 $Y=1.005
+ $X2=0 $Y2=0
cc_552 N_A_336_347#_c_600_n N_VGND_M1023_d 0.0119522f $X=4.765 $Y=1.005 $X2=0
+ $Y2=0
cc_553 N_A_336_347#_c_600_n N_VGND_M1014_d 0.00727468f $X=4.765 $Y=1.005 $X2=0
+ $Y2=0
cc_554 N_A_336_347#_c_615_n N_VGND_M1005_d 0.0147652f $X=6.765 $Y=1.005 $X2=0
+ $Y2=0
cc_555 N_A_336_347#_c_579_n N_VGND_M1005_d 5.91846e-19 $X=6.85 $Y=1.255 $X2=0
+ $Y2=0
cc_556 N_A_336_347#_c_577_n N_VGND_c_1382_n 0.0108145f $X=2.145 $Y=0.54 $X2=0
+ $Y2=0
cc_557 N_A_336_347#_c_600_n N_VGND_c_1382_n 0.0299353f $X=4.765 $Y=1.005 $X2=0
+ $Y2=0
cc_558 N_A_336_347#_c_577_n N_VGND_c_1386_n 0.013278f $X=2.145 $Y=0.54 $X2=0
+ $Y2=0
cc_559 N_A_336_347#_c_569_n N_VGND_c_1388_n 0.00533923f $X=5.02 $Y=1.245 $X2=0
+ $Y2=0
cc_560 N_A_336_347#_c_571_n N_VGND_c_1388_n 0.00423577f $X=7.055 $Y=1.255 $X2=0
+ $Y2=0
cc_561 N_A_336_347#_c_571_n N_VGND_c_1389_n 0.0042262f $X=7.055 $Y=1.255 $X2=0
+ $Y2=0
cc_562 N_A_336_347#_c_574_n N_VGND_c_1389_n 0.0042262f $X=7.485 $Y=1.255 $X2=0
+ $Y2=0
cc_563 N_A_336_347#_c_574_n N_VGND_c_1394_n 0.00422051f $X=7.485 $Y=1.255 $X2=0
+ $Y2=0
cc_564 N_A_336_347#_c_569_n N_VGND_c_1395_n 0.00537853f $X=5.02 $Y=1.245 $X2=0
+ $Y2=0
cc_565 N_A_336_347#_c_571_n N_VGND_c_1395_n 0.00537853f $X=7.055 $Y=1.255 $X2=0
+ $Y2=0
cc_566 N_A_336_347#_c_574_n N_VGND_c_1395_n 0.00537853f $X=7.485 $Y=1.255 $X2=0
+ $Y2=0
cc_567 N_A_336_347#_c_577_n N_VGND_c_1395_n 0.0119308f $X=2.145 $Y=0.54 $X2=0
+ $Y2=0
cc_568 N_A_336_347#_c_600_n A_487_79# 0.00630082f $X=4.765 $Y=1.005 $X2=-0.19
+ $Y2=-0.245
cc_569 N_A_336_347#_c_600_n N_A_701_79#_M1030_d 0.0048411f $X=4.765 $Y=1.005
+ $X2=-0.19 $Y2=-0.245
cc_570 N_A_336_347#_c_600_n N_A_701_79#_M1015_d 0.00595956f $X=4.765 $Y=1.005
+ $X2=0 $Y2=0
cc_571 N_A_336_347#_c_578_n N_A_701_79#_M1015_d 5.82479e-19 $X=4.93 $Y=1.41
+ $X2=0 $Y2=0
cc_572 N_A_336_347#_c_759_p N_A_701_79#_M1015_d 0.00135186f $X=4.93 $Y=1.005
+ $X2=0 $Y2=0
cc_573 N_A_336_347#_c_600_n N_A_701_79#_c_1482_n 0.0162804f $X=4.765 $Y=1.005
+ $X2=0 $Y2=0
cc_574 N_A_336_347#_c_568_n N_A_701_79#_c_1485_n 5.7535e-19 $X=4.885 $Y=1.66
+ $X2=0 $Y2=0
cc_575 N_A_336_347#_c_569_n N_A_701_79#_c_1485_n 0.0092157f $X=5.02 $Y=1.245
+ $X2=0 $Y2=0
cc_576 N_A_336_347#_c_759_p N_A_701_79#_c_1485_n 0.0124344f $X=4.93 $Y=1.005
+ $X2=0 $Y2=0
cc_577 N_A_336_347#_c_600_n N_A_701_79#_c_1486_n 0.0563239f $X=4.765 $Y=1.005
+ $X2=0 $Y2=0
cc_578 N_A_336_347#_c_615_n A_1119_79# 0.00486686f $X=6.765 $Y=1.005 $X2=-0.19
+ $Y2=-0.245
cc_579 N_A_336_347#_c_615_n A_1205_79# 0.00369412f $X=6.765 $Y=1.005 $X2=-0.19
+ $Y2=-0.245
cc_580 N_B_c_794_n N_A_992_347#_c_980_n 0.00764906f $X=5.845 $Y=3.15 $X2=0 $Y2=0
cc_581 N_B_M1012_g N_A_992_347#_c_980_n 0.0139873f $X=5.935 $Y=2.34 $X2=0 $Y2=0
cc_582 N_B_c_777_n N_A_992_347#_c_984_n 0.0109897f $X=5.935 $Y=1.21 $X2=0 $Y2=0
cc_583 N_B_c_794_n N_A_992_347#_c_978_n 0.00638811f $X=5.845 $Y=3.15 $X2=0 $Y2=0
cc_584 N_B_M1012_g N_A_992_347#_c_978_n 0.00236384f $X=5.935 $Y=2.34 $X2=0 $Y2=0
cc_585 N_B_c_777_n N_A_992_347#_c_971_n 0.00108597f $X=5.935 $Y=1.21 $X2=0 $Y2=0
cc_586 N_B_M1022_g N_A_27_378#_c_1092_n 0.0120552f $X=1.155 $Y=2.235 $X2=0 $Y2=0
cc_587 B N_A_27_378#_c_1092_n 0.0152909f $X=0.635 $Y=1.95 $X2=0 $Y2=0
cc_588 N_B_M1022_g N_A_27_378#_c_1085_n 7.52797e-19 $X=1.155 $Y=2.235 $X2=0
+ $Y2=0
cc_589 N_B_c_779_n N_A_27_378#_c_1086_n 5.05692e-19 $X=1.155 $Y=2.9 $X2=0 $Y2=0
cc_590 N_B_M1022_g N_A_27_378#_c_1086_n 0.0106125f $X=1.155 $Y=2.235 $X2=0 $Y2=0
cc_591 N_B_c_783_n N_A_27_378#_c_1086_n 0.00398225f $X=2.255 $Y=3.15 $X2=0 $Y2=0
cc_592 B N_A_27_378#_c_1086_n 0.00264329f $X=0.635 $Y=1.95 $X2=0 $Y2=0
cc_593 B N_VPWR_M1019_d 0.00787393f $X=0.635 $Y=1.95 $X2=-0.19 $Y2=-0.245
cc_594 N_B_c_802_n N_VPWR_M1019_d 0.00328911f $X=0.72 $Y=1.92 $X2=-0.19
+ $Y2=-0.245
cc_595 N_B_c_779_n N_VPWR_c_1119_n 0.0147666f $X=1.155 $Y=2.9 $X2=0 $Y2=0
cc_596 N_B_M1022_g N_VPWR_c_1119_n 0.00265085f $X=1.155 $Y=2.235 $X2=0 $Y2=0
cc_597 N_B_c_786_n N_VPWR_c_1120_n 0.00653223f $X=2.345 $Y=2.9 $X2=0 $Y2=0
cc_598 N_B_M1028_g N_VPWR_c_1120_n 0.00190566f $X=2.345 $Y=2.235 $X2=0 $Y2=0
cc_599 N_B_c_790_n N_VPWR_c_1120_n 0.0259473f $X=3.755 $Y=3.15 $X2=0 $Y2=0
cc_600 N_B_M1010_g N_VPWR_c_1120_n 0.00253553f $X=3.845 $Y=2.39 $X2=0 $Y2=0
cc_601 N_B_c_799_n N_VPWR_c_1120_n 0.00266188f $X=3.845 $Y=3.15 $X2=0 $Y2=0
cc_602 N_B_M1010_g N_VPWR_c_1121_n 0.00901204f $X=3.845 $Y=2.39 $X2=0 $Y2=0
cc_603 N_B_c_794_n N_VPWR_c_1121_n 0.0228891f $X=5.845 $Y=3.15 $X2=0 $Y2=0
cc_604 N_B_c_799_n N_VPWR_c_1121_n 0.0123224f $X=3.845 $Y=3.15 $X2=0 $Y2=0
cc_605 N_B_c_800_n N_VPWR_c_1122_n 0.00558044f $X=5.935 $Y=3.15 $X2=0 $Y2=0
cc_606 N_B_c_784_n N_VPWR_c_1125_n 0.0555823f $X=1.245 $Y=3.15 $X2=0 $Y2=0
cc_607 N_B_c_794_n N_VPWR_c_1127_n 0.0543816f $X=5.845 $Y=3.15 $X2=0 $Y2=0
cc_608 N_B_c_790_n N_VPWR_c_1130_n 0.0232348f $X=3.755 $Y=3.15 $X2=0 $Y2=0
cc_609 N_B_c_783_n N_VPWR_c_1118_n 0.0315845f $X=2.255 $Y=3.15 $X2=0 $Y2=0
cc_610 N_B_c_784_n N_VPWR_c_1118_n 0.00780279f $X=1.245 $Y=3.15 $X2=0 $Y2=0
cc_611 N_B_c_790_n N_VPWR_c_1118_n 0.0374807f $X=3.755 $Y=3.15 $X2=0 $Y2=0
cc_612 N_B_c_794_n N_VPWR_c_1118_n 0.0448265f $X=5.845 $Y=3.15 $X2=0 $Y2=0
cc_613 N_B_c_798_n N_VPWR_c_1118_n 0.0109436f $X=2.345 $Y=3.15 $X2=0 $Y2=0
cc_614 N_B_c_799_n N_VPWR_c_1118_n 0.00453024f $X=3.845 $Y=3.15 $X2=0 $Y2=0
cc_615 N_B_c_800_n N_VPWR_c_1118_n 0.00805203f $X=5.935 $Y=3.15 $X2=0 $Y2=0
cc_616 N_B_c_790_n N_A_683_347#_c_1237_n 0.00619091f $X=3.755 $Y=3.15 $X2=0
+ $Y2=0
cc_617 N_B_M1010_g N_A_683_347#_c_1238_n 6.83896e-19 $X=3.845 $Y=2.39 $X2=0
+ $Y2=0
cc_618 N_B_c_794_n N_A_683_347#_c_1238_n 0.00601703f $X=5.845 $Y=3.15 $X2=0
+ $Y2=0
cc_619 N_B_M1010_g N_A_683_347#_c_1243_n 0.0115741f $X=3.845 $Y=2.39 $X2=0 $Y2=0
cc_620 N_B_c_794_n N_A_683_347#_c_1243_n 0.0024022f $X=5.845 $Y=3.15 $X2=0 $Y2=0
cc_621 N_B_c_767_n N_A_27_79#_c_1345_n 2.208e-19 $X=1.14 $Y=1.245 $X2=0 $Y2=0
cc_622 N_B_c_767_n N_A_27_79#_c_1348_n 0.00874326f $X=1.14 $Y=1.245 $X2=0 $Y2=0
cc_623 N_B_c_768_n N_A_27_79#_c_1348_n 0.00442488f $X=1.155 $Y=1.66 $X2=0 $Y2=0
cc_624 N_B_c_778_n N_A_27_79#_c_1348_n 0.0350363f $X=1 $Y=1.41 $X2=0 $Y2=0
cc_625 N_B_c_767_n N_A_27_79#_c_1346_n 2.41236e-19 $X=1.14 $Y=1.245 $X2=0 $Y2=0
cc_626 N_B_c_767_n N_A_27_79#_c_1355_n 0.00576482f $X=1.14 $Y=1.245 $X2=0 $Y2=0
cc_627 N_B_c_767_n N_A_27_79#_c_1370_n 0.00875087f $X=1.14 $Y=1.245 $X2=0 $Y2=0
cc_628 N_B_c_767_n N_A_27_79#_c_1356_n 0.00700064f $X=1.14 $Y=1.245 $X2=0 $Y2=0
cc_629 N_B_c_767_n N_VGND_c_1381_n 0.00479734f $X=1.14 $Y=1.245 $X2=0 $Y2=0
cc_630 N_B_c_775_n N_VGND_c_1382_n 0.00147287f $X=2.345 $Y=1.21 $X2=0 $Y2=0
cc_631 N_B_c_767_n N_VGND_c_1386_n 0.00404918f $X=1.14 $Y=1.245 $X2=0 $Y2=0
cc_632 N_B_c_775_n N_VGND_c_1386_n 0.00534051f $X=2.345 $Y=1.21 $X2=0 $Y2=0
cc_633 N_B_c_776_n N_VGND_c_1387_n 0.00420261f $X=3.845 $Y=1.21 $X2=0 $Y2=0
cc_634 N_B_c_777_n N_VGND_c_1388_n 0.0042262f $X=5.935 $Y=1.21 $X2=0 $Y2=0
cc_635 N_B_c_776_n N_VGND_c_1393_n 0.00348026f $X=3.845 $Y=1.21 $X2=0 $Y2=0
cc_636 N_B_c_767_n N_VGND_c_1395_n 0.00537853f $X=1.14 $Y=1.245 $X2=0 $Y2=0
cc_637 N_B_c_775_n N_VGND_c_1395_n 0.00537853f $X=2.345 $Y=1.21 $X2=0 $Y2=0
cc_638 N_B_c_776_n N_VGND_c_1395_n 0.00537853f $X=3.845 $Y=1.21 $X2=0 $Y2=0
cc_639 N_B_c_777_n N_VGND_c_1395_n 0.00537853f $X=5.935 $Y=1.21 $X2=0 $Y2=0
cc_640 N_B_c_776_n N_A_701_79#_c_1482_n 0.00558627f $X=3.845 $Y=1.21 $X2=0 $Y2=0
cc_641 N_B_c_776_n N_A_701_79#_c_1485_n 7.16157e-19 $X=3.845 $Y=1.21 $X2=0 $Y2=0
cc_642 N_B_c_776_n N_A_701_79#_c_1486_n 0.00933014f $X=3.845 $Y=1.21 $X2=0 $Y2=0
cc_643 N_A_992_347#_c_980_n N_VPWR_M1016_d 0.0129328f $X=7.88 $Y=2.405 $X2=0
+ $Y2=0
cc_644 N_A_992_347#_c_980_n N_VPWR_M1031_d 0.0186333f $X=7.88 $Y=2.405 $X2=0
+ $Y2=0
cc_645 N_A_992_347#_c_977_n N_VPWR_M1031_d 0.00976076f $X=7.965 $Y=2.32 $X2=0
+ $Y2=0
cc_646 N_A_992_347#_c_980_n N_VPWR_c_1122_n 0.0214521f $X=7.88 $Y=2.405 $X2=0
+ $Y2=0
cc_647 N_A_992_347#_c_976_n N_VPWR_c_1124_n 0.00963415f $X=8.61 $Y=1.765 $X2=0
+ $Y2=0
cc_648 N_A_992_347#_c_978_n N_VPWR_c_1127_n 0.00750989f $X=5.17 $Y=2.195 $X2=0
+ $Y2=0
cc_649 N_A_992_347#_c_965_n N_VPWR_c_1132_n 0.00445602f $X=8.16 $Y=1.765 $X2=0
+ $Y2=0
cc_650 N_A_992_347#_c_976_n N_VPWR_c_1132_n 0.00417277f $X=8.61 $Y=1.765 $X2=0
+ $Y2=0
cc_651 N_A_992_347#_c_965_n N_VPWR_c_1135_n 0.00562118f $X=8.16 $Y=1.765 $X2=0
+ $Y2=0
cc_652 N_A_992_347#_c_980_n N_VPWR_c_1135_n 0.0270364f $X=7.88 $Y=2.405 $X2=0
+ $Y2=0
cc_653 N_A_992_347#_c_965_n N_VPWR_c_1118_n 0.00858753f $X=8.16 $Y=1.765 $X2=0
+ $Y2=0
cc_654 N_A_992_347#_c_976_n N_VPWR_c_1118_n 0.00769383f $X=8.61 $Y=1.765 $X2=0
+ $Y2=0
cc_655 N_A_992_347#_c_980_n N_VPWR_c_1118_n 0.0615814f $X=7.88 $Y=2.405 $X2=0
+ $Y2=0
cc_656 N_A_992_347#_c_978_n N_VPWR_c_1118_n 0.00907713f $X=5.17 $Y=2.195 $X2=0
+ $Y2=0
cc_657 N_A_992_347#_c_978_n N_A_683_347#_c_1238_n 0.0186593f $X=5.17 $Y=2.195
+ $X2=0 $Y2=0
cc_658 N_A_992_347#_c_980_n A_1094_347# 0.00771309f $X=7.88 $Y=2.405 $X2=-0.19
+ $Y2=-0.245
cc_659 N_A_992_347#_c_980_n A_1202_368# 0.00624598f $X=7.88 $Y=2.405 $X2=-0.19
+ $Y2=-0.245
cc_660 N_A_992_347#_c_984_n N_COUT_M1007_d 0.00433887f $X=7.88 $Y=0.66 $X2=-0.19
+ $Y2=-0.245
cc_661 N_A_992_347#_c_980_n N_COUT_M1020_s 0.0089693f $X=7.88 $Y=2.405 $X2=0
+ $Y2=0
cc_662 N_A_992_347#_c_984_n N_COUT_c_1280_n 0.024721f $X=7.88 $Y=0.66 $X2=0
+ $Y2=0
cc_663 N_A_992_347#_c_973_n N_COUT_c_1280_n 0.00783929f $X=8.057 $Y=1.32 $X2=0
+ $Y2=0
cc_664 N_A_992_347#_c_965_n N_COUT_c_1276_n 4.03982e-19 $X=8.16 $Y=1.765 $X2=0
+ $Y2=0
cc_665 N_A_992_347#_c_980_n N_COUT_c_1276_n 0.0114263f $X=7.88 $Y=2.405 $X2=0
+ $Y2=0
cc_666 N_A_992_347#_c_977_n N_COUT_c_1276_n 0.0080394f $X=7.965 $Y=2.32 $X2=0
+ $Y2=0
cc_667 N_A_992_347#_c_973_n N_COUT_c_1276_n 0.0334028f $X=8.057 $Y=1.32 $X2=0
+ $Y2=0
cc_668 N_A_992_347#_c_980_n N_COUT_c_1278_n 0.0225082f $X=7.88 $Y=2.405 $X2=0
+ $Y2=0
cc_669 N_A_992_347#_M1009_g N_SUM_c_1305_n 0.00978782f $X=8.195 $Y=0.765 $X2=0
+ $Y2=0
cc_670 N_A_992_347#_M1013_g N_SUM_c_1305_n 0.00778673f $X=8.625 $Y=0.765 $X2=0
+ $Y2=0
cc_671 N_A_992_347#_c_984_n N_SUM_c_1305_n 0.0126255f $X=7.88 $Y=0.66 $X2=0
+ $Y2=0
cc_672 N_A_992_347#_c_973_n N_SUM_c_1305_n 0.0268531f $X=8.057 $Y=1.32 $X2=0
+ $Y2=0
cc_673 N_A_992_347#_M1009_g N_SUM_c_1306_n 0.00251262f $X=8.195 $Y=0.765 $X2=0
+ $Y2=0
cc_674 N_A_992_347#_c_967_n N_SUM_c_1306_n 0.00120743f $X=8.52 $Y=1.395 $X2=0
+ $Y2=0
cc_675 N_A_992_347#_M1013_g N_SUM_c_1306_n 0.00196897f $X=8.625 $Y=0.765 $X2=0
+ $Y2=0
cc_676 N_A_992_347#_c_965_n SUM 0.00360044f $X=8.16 $Y=1.765 $X2=0 $Y2=0
cc_677 N_A_992_347#_c_967_n SUM 0.00338114f $X=8.52 $Y=1.395 $X2=0 $Y2=0
cc_678 N_A_992_347#_c_976_n SUM 0.00233168f $X=8.61 $Y=1.765 $X2=0 $Y2=0
cc_679 N_A_992_347#_c_977_n SUM 0.019649f $X=7.965 $Y=2.32 $X2=0 $Y2=0
cc_680 N_A_992_347#_c_972_n SUM 0.00104314f $X=8.07 $Y=1.485 $X2=0 $Y2=0
cc_681 N_A_992_347#_c_965_n SUM 0.0134178f $X=8.16 $Y=1.765 $X2=0 $Y2=0
cc_682 N_A_992_347#_c_976_n SUM 0.0128557f $X=8.61 $Y=1.765 $X2=0 $Y2=0
cc_683 N_A_992_347#_c_965_n N_SUM_c_1307_n 0.00207353f $X=8.16 $Y=1.765 $X2=0
+ $Y2=0
cc_684 N_A_992_347#_M1009_g N_SUM_c_1307_n 9.71018e-19 $X=8.195 $Y=0.765 $X2=0
+ $Y2=0
cc_685 N_A_992_347#_c_967_n N_SUM_c_1307_n 0.00773415f $X=8.52 $Y=1.395 $X2=0
+ $Y2=0
cc_686 N_A_992_347#_c_968_n N_SUM_c_1307_n 0.00994975f $X=8.61 $Y=1.675 $X2=0
+ $Y2=0
cc_687 N_A_992_347#_c_976_n N_SUM_c_1307_n 0.00782818f $X=8.61 $Y=1.765 $X2=0
+ $Y2=0
cc_688 N_A_992_347#_M1013_g N_SUM_c_1307_n 0.008382f $X=8.625 $Y=0.765 $X2=0
+ $Y2=0
cc_689 N_A_992_347#_c_970_n N_SUM_c_1307_n 0.00647817f $X=8.61 $Y=1.395 $X2=0
+ $Y2=0
cc_690 N_A_992_347#_c_977_n N_SUM_c_1307_n 0.00538817f $X=7.965 $Y=2.32 $X2=0
+ $Y2=0
cc_691 N_A_992_347#_c_972_n N_SUM_c_1307_n 0.0243786f $X=8.07 $Y=1.485 $X2=0
+ $Y2=0
cc_692 N_A_992_347#_c_973_n N_SUM_c_1307_n 0.00538819f $X=8.057 $Y=1.32 $X2=0
+ $Y2=0
cc_693 N_A_992_347#_c_984_n N_VGND_M1005_d 0.0110898f $X=7.88 $Y=0.66 $X2=0
+ $Y2=0
cc_694 N_A_992_347#_c_984_n N_VGND_M1011_s 0.0188382f $X=7.88 $Y=0.66 $X2=0
+ $Y2=0
cc_695 N_A_992_347#_c_973_n N_VGND_M1011_s 0.0117254f $X=8.057 $Y=1.32 $X2=0
+ $Y2=0
cc_696 N_A_992_347#_M1013_g N_VGND_c_1384_n 0.00650727f $X=8.625 $Y=0.765 $X2=0
+ $Y2=0
cc_697 N_A_992_347#_c_984_n N_VGND_c_1388_n 0.0508119f $X=7.88 $Y=0.66 $X2=0
+ $Y2=0
cc_698 N_A_992_347#_c_971_n N_VGND_c_1388_n 0.0126849f $X=5.305 $Y=0.56 $X2=0
+ $Y2=0
cc_699 N_A_992_347#_c_984_n N_VGND_c_1389_n 0.0115584f $X=7.88 $Y=0.66 $X2=0
+ $Y2=0
cc_700 N_A_992_347#_M1009_g N_VGND_c_1390_n 0.00534051f $X=8.195 $Y=0.765 $X2=0
+ $Y2=0
cc_701 N_A_992_347#_M1013_g N_VGND_c_1390_n 0.00534051f $X=8.625 $Y=0.765 $X2=0
+ $Y2=0
cc_702 N_A_992_347#_M1009_g N_VGND_c_1394_n 0.00382295f $X=8.195 $Y=0.765 $X2=0
+ $Y2=0
cc_703 N_A_992_347#_c_984_n N_VGND_c_1394_n 0.0336382f $X=7.88 $Y=0.66 $X2=0
+ $Y2=0
cc_704 N_A_992_347#_M1009_g N_VGND_c_1395_n 0.00537853f $X=8.195 $Y=0.765 $X2=0
+ $Y2=0
cc_705 N_A_992_347#_M1013_g N_VGND_c_1395_n 0.00537853f $X=8.625 $Y=0.765 $X2=0
+ $Y2=0
cc_706 N_A_992_347#_c_984_n N_VGND_c_1395_n 0.0545367f $X=7.88 $Y=0.66 $X2=0
+ $Y2=0
cc_707 N_A_992_347#_c_971_n N_VGND_c_1395_n 0.0116693f $X=5.305 $Y=0.56 $X2=0
+ $Y2=0
cc_708 N_A_992_347#_c_984_n A_1119_79# 0.00447592f $X=7.88 $Y=0.66 $X2=-0.19
+ $Y2=-0.245
cc_709 N_A_992_347#_c_984_n A_1205_79# 0.00339738f $X=7.88 $Y=0.66 $X2=-0.19
+ $Y2=-0.245
cc_710 N_A_27_378#_c_1092_n N_VPWR_M1019_d 0.0113157f $X=1.215 $Y=2.405
+ $X2=-0.19 $Y2=1.66
cc_711 N_A_27_378#_c_1092_n N_VPWR_c_1119_n 0.0296023f $X=1.215 $Y=2.405 $X2=0
+ $Y2=0
cc_712 N_A_27_378#_c_1085_n N_VPWR_c_1119_n 0.0102777f $X=0.28 $Y=2.405 $X2=0
+ $Y2=0
cc_713 N_A_27_378#_c_1086_n N_VPWR_c_1119_n 0.00650757f $X=1.38 $Y=2.25 $X2=0
+ $Y2=0
cc_714 N_A_27_378#_c_1086_n N_VPWR_c_1125_n 0.00747926f $X=1.38 $Y=2.25 $X2=0
+ $Y2=0
cc_715 N_A_27_378#_c_1085_n N_VPWR_c_1129_n 0.0120606f $X=0.28 $Y=2.405 $X2=0
+ $Y2=0
cc_716 N_A_27_378#_c_1092_n N_VPWR_c_1118_n 0.0127953f $X=1.215 $Y=2.405 $X2=0
+ $Y2=0
cc_717 N_A_27_378#_c_1085_n N_VPWR_c_1118_n 0.0122796f $X=0.28 $Y=2.405 $X2=0
+ $Y2=0
cc_718 N_A_27_378#_c_1086_n N_VPWR_c_1118_n 0.00904062f $X=1.38 $Y=2.25 $X2=0
+ $Y2=0
cc_719 N_VPWR_c_1120_n N_A_683_347#_c_1237_n 0.0251519f $X=2.99 $Y=2.455 $X2=0
+ $Y2=0
cc_720 N_VPWR_c_1130_n N_A_683_347#_c_1237_n 0.00687345f $X=3.905 $Y=3.33 $X2=0
+ $Y2=0
cc_721 N_VPWR_c_1118_n N_A_683_347#_c_1237_n 0.00888901f $X=8.88 $Y=3.33 $X2=0
+ $Y2=0
cc_722 N_VPWR_c_1121_n N_A_683_347#_c_1238_n 0.00645158f $X=4.095 $Y=2.745 $X2=0
+ $Y2=0
cc_723 N_VPWR_c_1127_n N_A_683_347#_c_1238_n 0.00731715f $X=6.535 $Y=3.33 $X2=0
+ $Y2=0
cc_724 N_VPWR_c_1118_n N_A_683_347#_c_1238_n 0.00895337f $X=8.88 $Y=3.33 $X2=0
+ $Y2=0
cc_725 N_VPWR_M1010_d N_A_683_347#_c_1243_n 0.00737327f $X=3.92 $Y=1.89 $X2=0
+ $Y2=0
cc_726 N_VPWR_c_1121_n N_A_683_347#_c_1243_n 0.0258287f $X=4.095 $Y=2.745 $X2=0
+ $Y2=0
cc_727 N_VPWR_c_1118_n N_A_683_347#_c_1243_n 0.0118804f $X=8.88 $Y=3.33 $X2=0
+ $Y2=0
cc_728 N_VPWR_c_1124_n SUM 0.0866997f $X=8.835 $Y=1.985 $X2=0 $Y2=0
cc_729 N_VPWR_c_1132_n SUM 0.0155928f $X=8.75 $Y=3.33 $X2=0 $Y2=0
cc_730 N_VPWR_c_1135_n SUM 0.0103327f $X=7.79 $Y=2.815 $X2=0 $Y2=0
cc_731 N_VPWR_c_1118_n SUM 0.0127818f $X=8.88 $Y=3.33 $X2=0 $Y2=0
cc_732 N_VPWR_c_1124_n N_VGND_c_1384_n 0.00873044f $X=8.835 $Y=1.985 $X2=0 $Y2=0
cc_733 N_SUM_c_1305_n N_VGND_c_1384_n 0.0293573f $X=8.41 $Y=0.54 $X2=0 $Y2=0
cc_734 N_SUM_c_1305_n N_VGND_c_1390_n 0.0131608f $X=8.41 $Y=0.54 $X2=0 $Y2=0
cc_735 N_SUM_c_1305_n N_VGND_c_1394_n 0.0018709f $X=8.41 $Y=0.54 $X2=0 $Y2=0
cc_736 N_SUM_c_1305_n N_VGND_c_1395_n 0.0118885f $X=8.41 $Y=0.54 $X2=0 $Y2=0
cc_737 N_A_27_79#_c_1348_n N_VGND_M1017_d 0.013096f $X=1.035 $Y=0.99 $X2=-0.19
+ $Y2=-0.245
cc_738 N_A_27_79#_c_1345_n N_VGND_c_1381_n 0.014266f $X=0.28 $Y=0.54 $X2=0 $Y2=0
cc_739 N_A_27_79#_c_1348_n N_VGND_c_1381_n 0.019282f $X=1.035 $Y=0.99 $X2=0
+ $Y2=0
cc_740 N_A_27_79#_c_1345_n N_VGND_c_1385_n 0.0132298f $X=0.28 $Y=0.54 $X2=0
+ $Y2=0
cc_741 N_A_27_79#_c_1370_n N_VGND_c_1386_n 0.00502025f $X=1.205 $Y=0.585 $X2=0
+ $Y2=0
cc_742 N_A_27_79#_c_1356_n N_VGND_c_1386_n 0.0176852f $X=1.5 $Y=0.585 $X2=0
+ $Y2=0
cc_743 N_A_27_79#_c_1345_n N_VGND_c_1395_n 0.0119092f $X=0.28 $Y=0.54 $X2=0
+ $Y2=0
cc_744 N_A_27_79#_c_1370_n N_VGND_c_1395_n 0.00586634f $X=1.205 $Y=0.585 $X2=0
+ $Y2=0
cc_745 N_A_27_79#_c_1356_n N_VGND_c_1395_n 0.0207666f $X=1.5 $Y=0.585 $X2=0
+ $Y2=0
cc_746 N_VGND_c_1382_n N_A_701_79#_c_1482_n 0.0132266f $X=3.055 $Y=0.54 $X2=0
+ $Y2=0
cc_747 N_VGND_c_1387_n N_A_701_79#_c_1482_n 0.0126214f $X=3.99 $Y=0 $X2=0 $Y2=0
cc_748 N_VGND_c_1393_n N_A_701_79#_c_1482_n 0.00201367f $X=4.08 $Y=0 $X2=0 $Y2=0
cc_749 N_VGND_c_1395_n N_A_701_79#_c_1482_n 0.0116492f $X=8.88 $Y=0 $X2=0 $Y2=0
cc_750 N_VGND_c_1388_n N_A_701_79#_c_1485_n 0.0133589f $X=6.47 $Y=0 $X2=0 $Y2=0
cc_751 N_VGND_c_1395_n N_A_701_79#_c_1485_n 0.0161161f $X=8.88 $Y=0 $X2=0 $Y2=0
cc_752 N_VGND_M1014_d N_A_701_79#_c_1486_n 0.00736239f $X=3.935 $Y=0.395 $X2=0
+ $Y2=0
cc_753 N_VGND_c_1387_n N_A_701_79#_c_1486_n 0.0029521f $X=3.99 $Y=0 $X2=0 $Y2=0
cc_754 N_VGND_c_1388_n N_A_701_79#_c_1486_n 0.00294479f $X=6.47 $Y=0 $X2=0 $Y2=0
cc_755 N_VGND_c_1393_n N_A_701_79#_c_1486_n 0.0243979f $X=4.08 $Y=0 $X2=0 $Y2=0
cc_756 N_VGND_c_1395_n N_A_701_79#_c_1486_n 0.0121896f $X=8.88 $Y=0 $X2=0 $Y2=0
