* File: sky130_fd_sc_hs__or2b_2.pxi.spice
* Created: Tue Sep  1 20:20:13 2020
* 
x_PM_SKY130_FD_SC_HS__OR2B_2%B_N N_B_N_M1002_g N_B_N_c_64_n N_B_N_M1007_g B_N
+ N_B_N_c_65_n PM_SKY130_FD_SC_HS__OR2B_2%B_N
x_PM_SKY130_FD_SC_HS__OR2B_2%A_187_48# N_A_187_48#_M1003_d N_A_187_48#_M1004_d
+ N_A_187_48#_M1005_g N_A_187_48#_c_101_n N_A_187_48#_M1000_g
+ N_A_187_48#_M1006_g N_A_187_48#_c_102_n N_A_187_48#_M1009_g N_A_187_48#_c_92_n
+ N_A_187_48#_c_93_n N_A_187_48#_c_94_n N_A_187_48#_c_95_n N_A_187_48#_c_103_n
+ N_A_187_48#_c_96_n N_A_187_48#_c_97_n N_A_187_48#_c_98_n N_A_187_48#_c_99_n
+ N_A_187_48#_c_105_n N_A_187_48#_c_100_n PM_SKY130_FD_SC_HS__OR2B_2%A_187_48#
x_PM_SKY130_FD_SC_HS__OR2B_2%A N_A_c_195_n N_A_M1001_g N_A_M1003_g A N_A_c_197_n
+ PM_SKY130_FD_SC_HS__OR2B_2%A
x_PM_SKY130_FD_SC_HS__OR2B_2%A_27_368# N_A_27_368#_M1002_s N_A_27_368#_M1007_s
+ N_A_27_368#_c_231_n N_A_27_368#_M1004_g N_A_27_368#_M1008_g
+ N_A_27_368#_c_233_n N_A_27_368#_c_234_n N_A_27_368#_c_235_n
+ N_A_27_368#_c_236_n N_A_27_368#_c_268_n N_A_27_368#_c_241_n
+ N_A_27_368#_c_237_n N_A_27_368#_c_238_n PM_SKY130_FD_SC_HS__OR2B_2%A_27_368#
x_PM_SKY130_FD_SC_HS__OR2B_2%VPWR N_VPWR_M1007_d N_VPWR_M1009_s N_VPWR_c_321_n
+ N_VPWR_c_322_n N_VPWR_c_323_n N_VPWR_c_324_n VPWR N_VPWR_c_325_n
+ N_VPWR_c_320_n N_VPWR_c_327_n PM_SKY130_FD_SC_HS__OR2B_2%VPWR
x_PM_SKY130_FD_SC_HS__OR2B_2%X N_X_M1005_d N_X_M1000_d N_X_c_355_n N_X_c_369_n
+ N_X_c_359_n X X X PM_SKY130_FD_SC_HS__OR2B_2%X
x_PM_SKY130_FD_SC_HS__OR2B_2%VGND N_VGND_M1002_d N_VGND_M1006_s N_VGND_M1008_d
+ N_VGND_c_394_n N_VGND_c_395_n N_VGND_c_396_n N_VGND_c_397_n VGND
+ N_VGND_c_398_n N_VGND_c_399_n N_VGND_c_400_n N_VGND_c_401_n N_VGND_c_402_n
+ N_VGND_c_403_n PM_SKY130_FD_SC_HS__OR2B_2%VGND
cc_1 VNB N_B_N_M1002_g 0.0335026f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=0.835
cc_2 VNB N_B_N_c_64_n 0.034329f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.765
cc_3 VNB N_B_N_c_65_n 0.0146969f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.515
cc_4 VNB N_A_187_48#_M1005_g 0.0217666f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_5 VNB N_A_187_48#_M1006_g 0.024884f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_6 VNB N_A_187_48#_c_92_n 0.0117673f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_7 VNB N_A_187_48#_c_93_n 4.49632e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_A_187_48#_c_94_n 0.00280429f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A_187_48#_c_95_n 0.0126244f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_187_48#_c_96_n 0.00389497f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_187_48#_c_97_n 0.0716833f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_187_48#_c_98_n 0.00292651f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_187_48#_c_99_n 0.00658719f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_187_48#_c_100_n 0.0242522f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_c_195_n 0.0270095f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=1.35
cc_16 VNB N_A_M1003_g 0.0336313f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.26
cc_17 VNB N_A_c_197_n 0.00176544f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.515
cc_18 VNB N_A_27_368#_c_231_n 0.0362251f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.26
cc_19 VNB N_A_27_368#_M1008_g 0.0312833f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.515
cc_20 VNB N_A_27_368#_c_233_n 0.0214174f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_27_368#_c_234_n 0.00518554f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_27_368#_c_235_n 0.00961237f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_27_368#_c_236_n 0.00871721f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_27_368#_c_237_n 2.57084e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_27_368#_c_238_n 0.00602679f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_VPWR_c_320_n 0.143779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_X_c_355_n 0.00169063f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_28 VNB X 0.0024448f $X=-0.19 $Y=-0.245 $X2=0.337 $Y2=1.515
cc_29 VNB X 0.00423402f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_394_n 0.0157594f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.515
cc_31 VNB N_VGND_c_395_n 0.0102093f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_396_n 0.0122168f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_397_n 0.0302304f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_398_n 0.0204283f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_399_n 0.019013f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_400_n 0.018855f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_401_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_402_n 0.0127985f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_403_n 0.20914f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VPB N_B_N_c_64_n 0.0355634f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.765
cc_41 VPB N_B_N_c_65_n 0.00743971f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.515
cc_42 VPB N_A_187_48#_c_101_n 0.0183785f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.515
cc_43 VPB N_A_187_48#_c_102_n 0.018677f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_44 VPB N_A_187_48#_c_103_n 0.0393709f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_45 VPB N_A_187_48#_c_97_n 0.0149615f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_46 VPB N_A_187_48#_c_105_n 0.0114988f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_47 VPB N_A_187_48#_c_100_n 0.00780236f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_48 VPB N_A_c_195_n 0.0270058f $X=-0.19 $Y=1.66 $X2=0.5 $Y2=1.35
cc_49 VPB N_A_c_197_n 0.00371807f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.515
cc_50 VPB N_A_27_368#_c_231_n 0.0253489f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.26
cc_51 VPB N_A_27_368#_c_236_n 0.00324248f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_52 VPB N_A_27_368#_c_241_n 0.0348664f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_53 VPB N_A_27_368#_c_237_n 0.00130347f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_54 VPB N_VPWR_c_321_n 0.0170949f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.515
cc_55 VPB N_VPWR_c_322_n 0.0111109f $X=-0.19 $Y=1.66 $X2=0.337 $Y2=1.665
cc_56 VPB N_VPWR_c_323_n 0.0246006f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_57 VPB N_VPWR_c_324_n 0.00614127f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_58 VPB N_VPWR_c_325_n 0.0399421f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_59 VPB N_VPWR_c_320_n 0.103022f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_60 VPB N_VPWR_c_327_n 0.0274851f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_61 VPB N_X_c_355_n 0.00184297f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_62 VPB N_X_c_359_n 0.00352644f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.515
cc_63 N_B_N_M1002_g N_A_187_48#_M1005_g 0.0192799f $X=0.5 $Y=0.835 $X2=0 $Y2=0
cc_64 N_B_N_c_64_n N_A_187_48#_c_101_n 0.0246567f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_65 N_B_N_c_64_n N_A_187_48#_c_97_n 0.0121446f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_66 N_B_N_M1002_g N_A_27_368#_c_233_n 0.00874924f $X=0.5 $Y=0.835 $X2=0 $Y2=0
cc_67 N_B_N_M1002_g N_A_27_368#_c_234_n 0.0117776f $X=0.5 $Y=0.835 $X2=0 $Y2=0
cc_68 N_B_N_c_64_n N_A_27_368#_c_234_n 7.87309e-19 $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_69 N_B_N_c_65_n N_A_27_368#_c_234_n 0.00722636f $X=0.385 $Y=1.515 $X2=0 $Y2=0
cc_70 N_B_N_M1002_g N_A_27_368#_c_235_n 0.00377477f $X=0.5 $Y=0.835 $X2=0 $Y2=0
cc_71 N_B_N_c_64_n N_A_27_368#_c_235_n 0.00160577f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_72 N_B_N_c_65_n N_A_27_368#_c_235_n 0.0281151f $X=0.385 $Y=1.515 $X2=0 $Y2=0
cc_73 N_B_N_M1002_g N_A_27_368#_c_236_n 0.00374987f $X=0.5 $Y=0.835 $X2=0 $Y2=0
cc_74 N_B_N_c_64_n N_A_27_368#_c_236_n 0.00712517f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_75 N_B_N_c_65_n N_A_27_368#_c_236_n 0.0329132f $X=0.385 $Y=1.515 $X2=0 $Y2=0
cc_76 N_B_N_c_64_n N_A_27_368#_c_241_n 0.0289543f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_77 N_B_N_c_65_n N_A_27_368#_c_241_n 0.0338821f $X=0.385 $Y=1.515 $X2=0 $Y2=0
cc_78 N_B_N_c_64_n N_VPWR_c_321_n 0.00415725f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_79 N_B_N_c_64_n N_VPWR_c_320_n 0.00462577f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_80 N_B_N_c_64_n N_VPWR_c_327_n 0.00393265f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_81 N_B_N_M1002_g X 6.25529e-19 $X=0.5 $Y=0.835 $X2=0 $Y2=0
cc_82 N_B_N_M1002_g N_VGND_c_394_n 0.00456881f $X=0.5 $Y=0.835 $X2=0 $Y2=0
cc_83 N_B_N_M1002_g N_VGND_c_398_n 0.0043356f $X=0.5 $Y=0.835 $X2=0 $Y2=0
cc_84 N_B_N_M1002_g N_VGND_c_403_n 0.00487769f $X=0.5 $Y=0.835 $X2=0 $Y2=0
cc_85 N_A_187_48#_c_102_n N_A_c_195_n 0.0295781f $X=1.705 $Y=1.765 $X2=-0.19
+ $Y2=-0.245
cc_86 N_A_187_48#_c_92_n N_A_c_195_n 0.001217f $X=2.405 $Y=1.065 $X2=-0.19
+ $Y2=-0.245
cc_87 N_A_187_48#_c_96_n N_A_c_195_n 0.00103081f $X=1.63 $Y=1.465 $X2=-0.19
+ $Y2=-0.245
cc_88 N_A_187_48#_c_97_n N_A_c_195_n 0.0204599f $X=1.63 $Y=1.465 $X2=-0.19
+ $Y2=-0.245
cc_89 N_A_187_48#_M1006_g N_A_M1003_g 0.00791742f $X=1.445 $Y=0.74 $X2=0 $Y2=0
cc_90 N_A_187_48#_c_92_n N_A_M1003_g 0.0163044f $X=2.405 $Y=1.065 $X2=0 $Y2=0
cc_91 N_A_187_48#_c_94_n N_A_M1003_g 0.00334116f $X=2.57 $Y=0.515 $X2=0 $Y2=0
cc_92 N_A_187_48#_c_96_n N_A_M1003_g 2.80126e-19 $X=1.63 $Y=1.465 $X2=0 $Y2=0
cc_93 N_A_187_48#_c_97_n N_A_M1003_g 0.00168337f $X=1.63 $Y=1.465 $X2=0 $Y2=0
cc_94 N_A_187_48#_c_98_n N_A_M1003_g 0.00266234f $X=1.63 $Y=1.3 $X2=0 $Y2=0
cc_95 N_A_187_48#_c_102_n N_A_c_197_n 3.33341e-19 $X=1.705 $Y=1.765 $X2=0 $Y2=0
cc_96 N_A_187_48#_c_92_n N_A_c_197_n 0.021788f $X=2.405 $Y=1.065 $X2=0 $Y2=0
cc_97 N_A_187_48#_c_96_n N_A_c_197_n 0.0159518f $X=1.63 $Y=1.465 $X2=0 $Y2=0
cc_98 N_A_187_48#_c_97_n N_A_c_197_n 0.00346501f $X=1.63 $Y=1.465 $X2=0 $Y2=0
cc_99 N_A_187_48#_c_95_n N_A_27_368#_c_231_n 0.00168154f $X=3.105 $Y=1.065 $X2=0
+ $Y2=0
cc_100 N_A_187_48#_c_99_n N_A_27_368#_c_231_n 0.00282246f $X=2.57 $Y=1.065 $X2=0
+ $Y2=0
cc_101 N_A_187_48#_c_105_n N_A_27_368#_c_231_n 0.0322195f $X=3.04 $Y=1.985 $X2=0
+ $Y2=0
cc_102 N_A_187_48#_c_100_n N_A_27_368#_c_231_n 0.00540056f $X=3.075 $Y=1.82
+ $X2=0 $Y2=0
cc_103 N_A_187_48#_c_94_n N_A_27_368#_M1008_g 0.0128081f $X=2.57 $Y=0.515 $X2=0
+ $Y2=0
cc_104 N_A_187_48#_c_95_n N_A_27_368#_M1008_g 0.0127833f $X=3.105 $Y=1.065 $X2=0
+ $Y2=0
cc_105 N_A_187_48#_c_99_n N_A_27_368#_M1008_g 0.00267461f $X=2.57 $Y=1.065 $X2=0
+ $Y2=0
cc_106 N_A_187_48#_c_100_n N_A_27_368#_M1008_g 0.00533837f $X=3.075 $Y=1.82
+ $X2=0 $Y2=0
cc_107 N_A_187_48#_M1005_g N_A_27_368#_c_233_n 5.25364e-19 $X=1.01 $Y=0.74 $X2=0
+ $Y2=0
cc_108 N_A_187_48#_M1005_g N_A_27_368#_c_234_n 0.00118159f $X=1.01 $Y=0.74 $X2=0
+ $Y2=0
cc_109 N_A_187_48#_M1005_g N_A_27_368#_c_236_n 0.00250805f $X=1.01 $Y=0.74 $X2=0
+ $Y2=0
cc_110 N_A_187_48#_c_101_n N_A_27_368#_c_236_n 0.00146678f $X=1.04 $Y=1.765
+ $X2=0 $Y2=0
cc_111 N_A_187_48#_c_97_n N_A_27_368#_c_236_n 0.00290361f $X=1.63 $Y=1.465 $X2=0
+ $Y2=0
cc_112 N_A_187_48#_c_101_n N_A_27_368#_c_268_n 0.0191027f $X=1.04 $Y=1.765 $X2=0
+ $Y2=0
cc_113 N_A_187_48#_c_102_n N_A_27_368#_c_268_n 0.0182331f $X=1.705 $Y=1.765
+ $X2=0 $Y2=0
cc_114 N_A_187_48#_c_103_n N_A_27_368#_c_268_n 0.0142079f $X=3.04 $Y=2.695 $X2=0
+ $Y2=0
cc_115 N_A_187_48#_c_96_n N_A_27_368#_c_268_n 0.00374667f $X=1.63 $Y=1.465 $X2=0
+ $Y2=0
cc_116 N_A_187_48#_c_97_n N_A_27_368#_c_268_n 4.90248e-19 $X=1.63 $Y=1.465 $X2=0
+ $Y2=0
cc_117 N_A_187_48#_c_101_n N_A_27_368#_c_241_n 0.00735817f $X=1.04 $Y=1.765
+ $X2=0 $Y2=0
cc_118 N_A_187_48#_c_105_n N_A_27_368#_c_237_n 0.0315234f $X=3.04 $Y=1.985 $X2=0
+ $Y2=0
cc_119 N_A_187_48#_c_100_n N_A_27_368#_c_237_n 0.00639198f $X=3.075 $Y=1.82
+ $X2=0 $Y2=0
cc_120 N_A_187_48#_c_95_n N_A_27_368#_c_238_n 0.0145294f $X=3.105 $Y=1.065 $X2=0
+ $Y2=0
cc_121 N_A_187_48#_c_99_n N_A_27_368#_c_238_n 0.0170429f $X=2.57 $Y=1.065 $X2=0
+ $Y2=0
cc_122 N_A_187_48#_c_105_n N_A_27_368#_c_238_n 0.00497567f $X=3.04 $Y=1.985
+ $X2=0 $Y2=0
cc_123 N_A_187_48#_c_100_n N_A_27_368#_c_238_n 0.0251406f $X=3.075 $Y=1.82 $X2=0
+ $Y2=0
cc_124 N_A_187_48#_c_101_n N_VPWR_c_321_n 0.0139308f $X=1.04 $Y=1.765 $X2=0
+ $Y2=0
cc_125 N_A_187_48#_c_102_n N_VPWR_c_321_n 0.00217981f $X=1.705 $Y=1.765 $X2=0
+ $Y2=0
cc_126 N_A_187_48#_c_101_n N_VPWR_c_322_n 0.00217981f $X=1.04 $Y=1.765 $X2=0
+ $Y2=0
cc_127 N_A_187_48#_c_102_n N_VPWR_c_322_n 0.0138722f $X=1.705 $Y=1.765 $X2=0
+ $Y2=0
cc_128 N_A_187_48#_c_101_n N_VPWR_c_323_n 0.00413917f $X=1.04 $Y=1.765 $X2=0
+ $Y2=0
cc_129 N_A_187_48#_c_102_n N_VPWR_c_323_n 0.00413917f $X=1.705 $Y=1.765 $X2=0
+ $Y2=0
cc_130 N_A_187_48#_c_103_n N_VPWR_c_325_n 0.011933f $X=3.04 $Y=2.695 $X2=0 $Y2=0
cc_131 N_A_187_48#_c_101_n N_VPWR_c_320_n 0.0081943f $X=1.04 $Y=1.765 $X2=0
+ $Y2=0
cc_132 N_A_187_48#_c_102_n N_VPWR_c_320_n 0.0081943f $X=1.705 $Y=1.765 $X2=0
+ $Y2=0
cc_133 N_A_187_48#_c_103_n N_VPWR_c_320_n 0.0135963f $X=3.04 $Y=2.695 $X2=0
+ $Y2=0
cc_134 N_A_187_48#_M1005_g N_X_c_355_n 0.00296721f $X=1.01 $Y=0.74 $X2=0 $Y2=0
cc_135 N_A_187_48#_c_101_n N_X_c_355_n 0.00123216f $X=1.04 $Y=1.765 $X2=0 $Y2=0
cc_136 N_A_187_48#_M1006_g N_X_c_355_n 0.0014407f $X=1.445 $Y=0.74 $X2=0 $Y2=0
cc_137 N_A_187_48#_c_102_n N_X_c_355_n 9.35381e-19 $X=1.705 $Y=1.765 $X2=0 $Y2=0
cc_138 N_A_187_48#_c_93_n N_X_c_355_n 9.15778e-19 $X=1.795 $Y=1.065 $X2=0 $Y2=0
cc_139 N_A_187_48#_c_96_n N_X_c_355_n 0.0181937f $X=1.63 $Y=1.465 $X2=0 $Y2=0
cc_140 N_A_187_48#_c_97_n N_X_c_355_n 0.0226131f $X=1.63 $Y=1.465 $X2=0 $Y2=0
cc_141 N_A_187_48#_c_98_n N_X_c_355_n 0.0062371f $X=1.63 $Y=1.3 $X2=0 $Y2=0
cc_142 N_A_187_48#_c_101_n N_X_c_369_n 0.00845785f $X=1.04 $Y=1.765 $X2=0 $Y2=0
cc_143 N_A_187_48#_c_102_n N_X_c_359_n 0.0102028f $X=1.705 $Y=1.765 $X2=0 $Y2=0
cc_144 N_A_187_48#_c_96_n N_X_c_359_n 0.0128197f $X=1.63 $Y=1.465 $X2=0 $Y2=0
cc_145 N_A_187_48#_c_97_n N_X_c_359_n 0.0112221f $X=1.63 $Y=1.465 $X2=0 $Y2=0
cc_146 N_A_187_48#_M1005_g X 0.00874049f $X=1.01 $Y=0.74 $X2=0 $Y2=0
cc_147 N_A_187_48#_M1006_g X 0.0125066f $X=1.445 $Y=0.74 $X2=0 $Y2=0
cc_148 N_A_187_48#_M1005_g X 0.00231072f $X=1.01 $Y=0.74 $X2=0 $Y2=0
cc_149 N_A_187_48#_M1006_g X 0.00360017f $X=1.445 $Y=0.74 $X2=0 $Y2=0
cc_150 N_A_187_48#_c_93_n X 0.00969017f $X=1.795 $Y=1.065 $X2=0 $Y2=0
cc_151 N_A_187_48#_c_97_n X 0.00222206f $X=1.63 $Y=1.465 $X2=0 $Y2=0
cc_152 N_A_187_48#_c_92_n N_VGND_M1006_s 0.00423176f $X=2.405 $Y=1.065 $X2=0
+ $Y2=0
cc_153 N_A_187_48#_c_93_n N_VGND_M1006_s 0.00421622f $X=1.795 $Y=1.065 $X2=0
+ $Y2=0
cc_154 N_A_187_48#_c_95_n N_VGND_M1008_d 0.00361779f $X=3.105 $Y=1.065 $X2=0
+ $Y2=0
cc_155 N_A_187_48#_M1005_g N_VGND_c_394_n 0.0062918f $X=1.01 $Y=0.74 $X2=0 $Y2=0
cc_156 N_A_187_48#_M1006_g N_VGND_c_395_n 0.00495353f $X=1.445 $Y=0.74 $X2=0
+ $Y2=0
cc_157 N_A_187_48#_c_92_n N_VGND_c_395_n 0.0309019f $X=2.405 $Y=1.065 $X2=0
+ $Y2=0
cc_158 N_A_187_48#_c_93_n N_VGND_c_395_n 0.0152767f $X=1.795 $Y=1.065 $X2=0
+ $Y2=0
cc_159 N_A_187_48#_c_94_n N_VGND_c_395_n 0.0200457f $X=2.57 $Y=0.515 $X2=0 $Y2=0
cc_160 N_A_187_48#_c_96_n N_VGND_c_395_n 0.00200141f $X=1.63 $Y=1.465 $X2=0
+ $Y2=0
cc_161 N_A_187_48#_c_97_n N_VGND_c_395_n 0.00102847f $X=1.63 $Y=1.465 $X2=0
+ $Y2=0
cc_162 N_A_187_48#_c_94_n N_VGND_c_397_n 0.0172462f $X=2.57 $Y=0.515 $X2=0 $Y2=0
cc_163 N_A_187_48#_c_95_n N_VGND_c_397_n 0.0278586f $X=3.105 $Y=1.065 $X2=0
+ $Y2=0
cc_164 N_A_187_48#_M1005_g N_VGND_c_399_n 0.00434272f $X=1.01 $Y=0.74 $X2=0
+ $Y2=0
cc_165 N_A_187_48#_M1006_g N_VGND_c_399_n 0.00439937f $X=1.445 $Y=0.74 $X2=0
+ $Y2=0
cc_166 N_A_187_48#_c_94_n N_VGND_c_400_n 0.0145639f $X=2.57 $Y=0.515 $X2=0 $Y2=0
cc_167 N_A_187_48#_M1005_g N_VGND_c_403_n 0.00825333f $X=1.01 $Y=0.74 $X2=0
+ $Y2=0
cc_168 N_A_187_48#_M1006_g N_VGND_c_403_n 0.0084116f $X=1.445 $Y=0.74 $X2=0
+ $Y2=0
cc_169 N_A_187_48#_c_94_n N_VGND_c_403_n 0.0119984f $X=2.57 $Y=0.515 $X2=0 $Y2=0
cc_170 N_A_c_195_n N_A_27_368#_c_231_n 0.0543908f $X=2.275 $Y=1.765 $X2=0 $Y2=0
cc_171 N_A_M1003_g N_A_27_368#_c_231_n 0.0231545f $X=2.29 $Y=0.69 $X2=0 $Y2=0
cc_172 N_A_c_197_n N_A_27_368#_c_231_n 5.00732e-19 $X=2.2 $Y=1.515 $X2=0 $Y2=0
cc_173 N_A_M1003_g N_A_27_368#_M1008_g 0.0244563f $X=2.29 $Y=0.69 $X2=0 $Y2=0
cc_174 N_A_c_195_n N_A_27_368#_c_268_n 0.0173941f $X=2.275 $Y=1.765 $X2=0 $Y2=0
cc_175 N_A_c_197_n N_A_27_368#_c_268_n 0.0106437f $X=2.2 $Y=1.515 $X2=0 $Y2=0
cc_176 N_A_c_195_n N_A_27_368#_c_237_n 0.00993389f $X=2.275 $Y=1.765 $X2=0 $Y2=0
cc_177 N_A_c_197_n N_A_27_368#_c_237_n 0.00983193f $X=2.2 $Y=1.515 $X2=0 $Y2=0
cc_178 N_A_M1003_g N_A_27_368#_c_238_n 0.00253418f $X=2.29 $Y=0.69 $X2=0 $Y2=0
cc_179 N_A_c_197_n N_A_27_368#_c_238_n 0.0241464f $X=2.2 $Y=1.515 $X2=0 $Y2=0
cc_180 N_A_c_195_n N_VPWR_c_322_n 0.0105558f $X=2.275 $Y=1.765 $X2=0 $Y2=0
cc_181 N_A_c_195_n N_VPWR_c_325_n 0.0049405f $X=2.275 $Y=1.765 $X2=0 $Y2=0
cc_182 N_A_c_195_n N_VPWR_c_320_n 0.00508379f $X=2.275 $Y=1.765 $X2=0 $Y2=0
cc_183 N_A_c_195_n N_X_c_359_n 0.00110758f $X=2.275 $Y=1.765 $X2=0 $Y2=0
cc_184 N_A_M1003_g N_VGND_c_395_n 0.011727f $X=2.29 $Y=0.69 $X2=0 $Y2=0
cc_185 N_A_M1003_g N_VGND_c_400_n 0.00398535f $X=2.29 $Y=0.69 $X2=0 $Y2=0
cc_186 N_A_M1003_g N_VGND_c_403_n 0.00788205f $X=2.29 $Y=0.69 $X2=0 $Y2=0
cc_187 N_A_27_368#_c_236_n N_VPWR_M1007_d 0.00285261f $X=0.805 $Y=1.95 $X2=-0.19
+ $Y2=-0.245
cc_188 N_A_27_368#_c_268_n N_VPWR_M1007_d 8.29358e-19 $X=2.535 $Y=2.325
+ $X2=-0.19 $Y2=-0.245
cc_189 N_A_27_368#_c_241_n N_VPWR_M1007_d 0.0112471f $X=0.89 $Y=2.325 $X2=-0.19
+ $Y2=-0.245
cc_190 N_A_27_368#_c_268_n N_VPWR_M1009_s 0.0143552f $X=2.535 $Y=2.325 $X2=0
+ $Y2=0
cc_191 N_A_27_368#_c_268_n N_VPWR_c_321_n 0.00249443f $X=2.535 $Y=2.325 $X2=0
+ $Y2=0
cc_192 N_A_27_368#_c_241_n N_VPWR_c_321_n 0.0294588f $X=0.89 $Y=2.325 $X2=0
+ $Y2=0
cc_193 N_A_27_368#_c_268_n N_VPWR_c_322_n 0.0219756f $X=2.535 $Y=2.325 $X2=0
+ $Y2=0
cc_194 N_A_27_368#_c_231_n N_VPWR_c_325_n 0.0049405f $X=2.695 $Y=1.765 $X2=0
+ $Y2=0
cc_195 N_A_27_368#_c_231_n N_VPWR_c_320_n 0.00508379f $X=2.695 $Y=1.765 $X2=0
+ $Y2=0
cc_196 N_A_27_368#_c_241_n N_VPWR_c_320_n 0.0100331f $X=0.89 $Y=2.325 $X2=0
+ $Y2=0
cc_197 N_A_27_368#_c_241_n N_VPWR_c_327_n 0.00671799f $X=0.89 $Y=2.325 $X2=0
+ $Y2=0
cc_198 N_A_27_368#_c_268_n N_X_M1000_d 0.0206477f $X=2.535 $Y=2.325 $X2=0 $Y2=0
cc_199 N_A_27_368#_c_236_n N_X_c_355_n 0.0456299f $X=0.805 $Y=1.95 $X2=0 $Y2=0
cc_200 N_A_27_368#_c_236_n N_X_c_369_n 0.0100844f $X=0.805 $Y=1.95 $X2=0 $Y2=0
cc_201 N_A_27_368#_c_268_n N_X_c_369_n 0.00886631f $X=2.535 $Y=2.325 $X2=0 $Y2=0
cc_202 N_A_27_368#_c_241_n N_X_c_369_n 0.0103743f $X=0.89 $Y=2.325 $X2=0 $Y2=0
cc_203 N_A_27_368#_c_268_n N_X_c_359_n 0.0266632f $X=2.535 $Y=2.325 $X2=0 $Y2=0
cc_204 N_A_27_368#_c_233_n X 0.00439955f $X=0.285 $Y=0.835 $X2=0 $Y2=0
cc_205 N_A_27_368#_c_234_n X 0.00940933f $X=0.72 $Y=1.095 $X2=0 $Y2=0
cc_206 N_A_27_368#_c_268_n A_470_368# 0.0109095f $X=2.535 $Y=2.325 $X2=-0.19
+ $Y2=-0.245
cc_207 N_A_27_368#_c_237_n A_470_368# 0.00467536f $X=2.62 $Y=2.24 $X2=-0.19
+ $Y2=-0.245
cc_208 N_A_27_368#_c_234_n N_VGND_M1002_d 0.0033541f $X=0.72 $Y=1.095 $X2=-0.19
+ $Y2=-0.245
cc_209 N_A_27_368#_c_233_n N_VGND_c_394_n 0.0114804f $X=0.285 $Y=0.835 $X2=0
+ $Y2=0
cc_210 N_A_27_368#_c_234_n N_VGND_c_394_n 0.0213686f $X=0.72 $Y=1.095 $X2=0
+ $Y2=0
cc_211 N_A_27_368#_M1008_g N_VGND_c_395_n 6.4117e-19 $X=2.785 $Y=0.69 $X2=0
+ $Y2=0
cc_212 N_A_27_368#_M1008_g N_VGND_c_397_n 0.00656895f $X=2.785 $Y=0.69 $X2=0
+ $Y2=0
cc_213 N_A_27_368#_c_233_n N_VGND_c_398_n 0.00811255f $X=0.285 $Y=0.835 $X2=0
+ $Y2=0
cc_214 N_A_27_368#_M1008_g N_VGND_c_400_n 0.00434272f $X=2.785 $Y=0.69 $X2=0
+ $Y2=0
cc_215 N_A_27_368#_M1008_g N_VGND_c_403_n 0.00824856f $X=2.785 $Y=0.69 $X2=0
+ $Y2=0
cc_216 N_A_27_368#_c_233_n N_VGND_c_403_n 0.0106114f $X=0.285 $Y=0.835 $X2=0
+ $Y2=0
cc_217 X N_VGND_c_394_n 0.0182902f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_218 X N_VGND_c_395_n 0.018141f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_219 X N_VGND_c_399_n 0.0145071f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_220 X N_VGND_c_403_n 0.0119067f $X=1.115 $Y=0.47 $X2=0 $Y2=0
