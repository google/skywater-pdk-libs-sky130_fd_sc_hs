* File: sky130_fd_sc_hs__a2bb2oi_2.pex.spice
* Created: Tue Sep  1 19:52:03 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HS__A2BB2OI_2%A1_N 1 3 4 5 7 11 13 15 19
r29 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.27
+ $Y=0.45 $X2=0.27 $Y2=0.45
r30 15 18 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=0.27 $Y=0.36 $X2=0.27
+ $Y2=0.45
r31 13 19 3.66686 $w=3.28e-07 $l=1.05e-07 $layer=LI1_cond $X=0.27 $Y=0.555
+ $X2=0.27 $Y2=0.45
r32 11 12 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=0.985 $Y=0.83
+ $X2=0.985 $Y2=1.225
r33 8 11 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=0.985 $Y=0.435
+ $X2=0.985 $Y2=0.83
r34 5 7 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=0.97 $Y=1.885
+ $X2=0.97 $Y2=2.46
r35 4 5 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=0.97 $Y=1.795 $X2=0.97
+ $Y2=1.885
r36 3 12 37.1337 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=0.97 $Y=1.315 $X2=0.97
+ $Y2=1.225
r37 3 4 186.581 $w=1.8e-07 $l=4.8e-07 $layer=POLY_cond $X=0.97 $Y=1.315 $X2=0.97
+ $Y2=1.795
r38 2 15 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.435 $Y=0.36
+ $X2=0.27 $Y2=0.36
r39 1 8 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.91 $Y=0.36
+ $X2=0.985 $Y2=0.435
r40 1 2 243.564 $w=1.5e-07 $l=4.75e-07 $layer=POLY_cond $X=0.91 $Y=0.36
+ $X2=0.435 $Y2=0.36
.ends

.subckt PM_SKY130_FD_SC_HS__A2BB2OI_2%A2_N 1 3 6 8 12
c33 12 0 1.88217e-19 $X=1.435 $Y=1.615
c34 6 0 1.77687e-19 $X=1.46 $Y=0.83
r35 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.435
+ $Y=1.615 $X2=1.435 $Y2=1.615
r36 8 12 8.20679 $w=3.28e-07 $l=2.35e-07 $layer=LI1_cond $X=1.2 $Y=1.615
+ $X2=1.435 $Y2=1.615
r37 4 11 38.5916 $w=2.93e-07 $l=1.77059e-07 $layer=POLY_cond $X=1.46 $Y=1.45
+ $X2=1.435 $Y2=1.615
r38 4 6 317.915 $w=1.5e-07 $l=6.2e-07 $layer=POLY_cond $X=1.46 $Y=1.45 $X2=1.46
+ $Y2=0.83
r39 1 11 55.8646 $w=2.93e-07 $l=3.05205e-07 $layer=POLY_cond $X=1.36 $Y=1.885
+ $X2=1.435 $Y2=1.615
r40 1 3 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=1.36 $Y=1.885
+ $X2=1.36 $Y2=2.46
.ends

.subckt PM_SKY130_FD_SC_HS__A2BB2OI_2%A_212_102# 1 2 9 13 15 17 18 19 20 22 23
+ 27 29 30 33 35 38 39
c92 39 0 1.56524e-19 $X=1.665 $Y=1.95
c93 27 0 1.77687e-19 $X=1.22 $Y=0.655
c94 20 0 4.43259e-20 $X=2.92 $Y=1.765
c95 19 0 1.88217e-19 $X=2.56 $Y=1.575
c96 15 0 9.92294e-20 $X=2.47 $Y=1.765
r97 46 47 13.0663 $w=3.32e-07 $l=9e-08 $layer=POLY_cond $X=2.38 $Y=1.542
+ $X2=2.47 $Y2=1.542
r98 43 46 49.3614 $w=3.32e-07 $l=3.4e-07 $layer=POLY_cond $X=2.04 $Y=1.542
+ $X2=2.38 $Y2=1.542
r99 43 44 13.0663 $w=3.32e-07 $l=9e-08 $layer=POLY_cond $X=2.04 $Y=1.542
+ $X2=1.95 $Y2=1.542
r100 42 43 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.04
+ $Y=1.485 $X2=2.04 $Y2=1.485
r101 38 39 9.45624 $w=4.88e-07 $l=1.65e-07 $layer=LI1_cond $X=1.665 $Y=2.115
+ $X2=1.665 $Y2=1.95
r102 35 42 8.98608 $w=3.5e-07 $l=2.26892e-07 $layer=LI1_cond $X=1.825 $Y=1.65
+ $X2=1.972 $Y2=1.485
r103 35 39 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=1.825 $Y=1.65
+ $X2=1.825 $Y2=1.95
r104 31 38 1.95278 $w=4.88e-07 $l=8e-08 $layer=LI1_cond $X=1.665 $Y=2.195
+ $X2=1.665 $Y2=2.115
r105 31 33 15.1341 $w=4.88e-07 $l=6.2e-07 $layer=LI1_cond $X=1.665 $Y=2.195
+ $X2=1.665 $Y2=2.815
r106 29 42 10.1086 $w=3.5e-07 $l=3.89076e-07 $layer=LI1_cond $X=1.74 $Y=1.195
+ $X2=1.972 $Y2=1.485
r107 29 30 26.7487 $w=1.68e-07 $l=4.1e-07 $layer=LI1_cond $X=1.74 $Y=1.195
+ $X2=1.33 $Y2=1.195
r108 25 30 7.47753 $w=1.7e-07 $l=1.85699e-07 $layer=LI1_cond $X=1.182 $Y=1.11
+ $X2=1.33 $Y2=1.195
r109 25 27 17.775 $w=2.93e-07 $l=4.55e-07 $layer=LI1_cond $X=1.182 $Y=1.11
+ $X2=1.182 $Y2=0.655
r110 20 23 76.0046 $w=1.8e-07 $l=1.9e-07 $layer=POLY_cond $X=2.92 $Y=1.765
+ $X2=2.92 $Y2=1.575
r111 20 22 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.92 $Y=1.765
+ $X2=2.92 $Y2=2.4
r112 19 47 27.7253 $w=3.32e-07 $l=1.05214e-07 $layer=POLY_cond $X=2.56 $Y=1.575
+ $X2=2.47 $Y2=1.542
r113 18 23 7.1379 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=2.83 $Y=1.575 $X2=2.92
+ $Y2=1.575
r114 18 19 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=2.83 $Y=1.575
+ $X2=2.56 $Y2=1.575
r115 15 47 21.3668 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=2.47 $Y=1.765
+ $X2=2.47 $Y2=1.542
r116 15 17 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.47 $Y=1.765
+ $X2=2.47 $Y2=2.4
r117 11 46 21.3668 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=2.38 $Y=1.32
+ $X2=2.38 $Y2=1.542
r118 11 13 276.894 $w=1.5e-07 $l=5.4e-07 $layer=POLY_cond $X=2.38 $Y=1.32
+ $X2=2.38 $Y2=0.78
r119 7 44 21.3668 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=1.95 $Y=1.32
+ $X2=1.95 $Y2=1.542
r120 7 9 276.894 $w=1.5e-07 $l=5.4e-07 $layer=POLY_cond $X=1.95 $Y=1.32 $X2=1.95
+ $Y2=0.78
r121 2 38 400 $w=1.7e-07 $l=2.17428e-07 $layer=licon1_PDIFF $count=1 $X=1.435
+ $Y=1.96 $X2=1.585 $Y2=2.115
r122 2 33 400 $w=1.7e-07 $l=9.26971e-07 $layer=licon1_PDIFF $count=1 $X=1.435
+ $Y=1.96 $X2=1.585 $Y2=2.815
r123 1 27 91 $w=1.7e-07 $l=2.20907e-07 $layer=licon1_NDIFF $count=2 $X=1.06
+ $Y=0.51 $X2=1.22 $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_HS__A2BB2OI_2%B2 1 3 6 8 10 13 15 21 22
c53 21 0 1.73551e-19 $X=3.57 $Y=1.485
c54 13 0 2.40437e-20 $X=3.845 $Y=0.74
c55 8 0 1.25206e-19 $X=3.82 $Y=1.765
r56 22 23 3.08184 $w=3.91e-07 $l=2.5e-08 $layer=POLY_cond $X=3.82 $Y=1.542
+ $X2=3.845 $Y2=1.542
r57 20 22 30.8184 $w=3.91e-07 $l=2.5e-07 $layer=POLY_cond $X=3.57 $Y=1.542
+ $X2=3.82 $Y2=1.542
r58 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.57
+ $Y=1.485 $X2=3.57 $Y2=1.485
r59 18 20 19.1074 $w=3.91e-07 $l=1.55e-07 $layer=POLY_cond $X=3.415 $Y=1.542
+ $X2=3.57 $Y2=1.542
r60 17 18 5.54731 $w=3.91e-07 $l=4.5e-08 $layer=POLY_cond $X=3.37 $Y=1.542
+ $X2=3.415 $Y2=1.542
r61 15 21 6.28605 $w=3.28e-07 $l=1.8e-07 $layer=LI1_cond $X=3.57 $Y=1.665
+ $X2=3.57 $Y2=1.485
r62 11 23 25.3065 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=3.845 $Y=1.32
+ $X2=3.845 $Y2=1.542
r63 11 13 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=3.845 $Y=1.32
+ $X2=3.845 $Y2=0.74
r64 8 22 25.3065 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=3.82 $Y=1.765
+ $X2=3.82 $Y2=1.542
r65 8 10 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.82 $Y=1.765
+ $X2=3.82 $Y2=2.4
r66 4 18 25.3065 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=3.415 $Y=1.32
+ $X2=3.415 $Y2=1.542
r67 4 6 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=3.415 $Y=1.32
+ $X2=3.415 $Y2=0.74
r68 1 17 25.3065 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=3.37 $Y=1.765
+ $X2=3.37 $Y2=1.542
r69 1 3 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.37 $Y=1.765
+ $X2=3.37 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_HS__A2BB2OI_2%B1 1 3 6 10 12 14 15 16 24
c42 16 0 1.25206e-19 $X=4.56 $Y=1.665
c43 6 0 3.50294e-19 $X=4.275 $Y=0.74
r44 24 25 1.9127 $w=3.78e-07 $l=1.5e-08 $layer=POLY_cond $X=4.705 $Y=1.557
+ $X2=4.72 $Y2=1.557
r45 22 24 45.9048 $w=3.78e-07 $l=3.6e-07 $layer=POLY_cond $X=4.345 $Y=1.557
+ $X2=4.705 $Y2=1.557
r46 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.345
+ $Y=1.515 $X2=4.345 $Y2=1.515
r47 20 22 8.92593 $w=3.78e-07 $l=7e-08 $layer=POLY_cond $X=4.275 $Y=1.557
+ $X2=4.345 $Y2=1.557
r48 19 20 0.637566 $w=3.78e-07 $l=5e-09 $layer=POLY_cond $X=4.27 $Y=1.557
+ $X2=4.275 $Y2=1.557
r49 16 23 5.76222 $w=4.28e-07 $l=2.15e-07 $layer=LI1_cond $X=4.56 $Y=1.565
+ $X2=4.345 $Y2=1.565
r50 15 23 7.10226 $w=4.28e-07 $l=2.65e-07 $layer=LI1_cond $X=4.08 $Y=1.565
+ $X2=4.345 $Y2=1.565
r51 12 25 24.4846 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=4.72 $Y=1.765
+ $X2=4.72 $Y2=1.557
r52 12 14 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=4.72 $Y=1.765
+ $X2=4.72 $Y2=2.4
r53 8 24 24.4846 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.705 $Y=1.35
+ $X2=4.705 $Y2=1.557
r54 8 10 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=4.705 $Y=1.35
+ $X2=4.705 $Y2=0.74
r55 4 20 24.4846 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.275 $Y=1.35
+ $X2=4.275 $Y2=1.557
r56 4 6 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=4.275 $Y=1.35
+ $X2=4.275 $Y2=0.74
r57 1 19 24.4846 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=4.27 $Y=1.765
+ $X2=4.27 $Y2=1.557
r58 1 3 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=4.27 $Y=1.765
+ $X2=4.27 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_HS__A2BB2OI_2%VPWR 1 2 3 12 18 22 24 26 31 39 46 47 50
+ 53 56
r57 56 57 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r58 53 54 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r59 50 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r60 47 57 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=4.56 $Y2=3.33
r61 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r62 44 56 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.66 $Y=3.33
+ $X2=4.495 $Y2=3.33
r63 44 46 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=4.66 $Y=3.33
+ $X2=5.04 $Y2=3.33
r64 43 57 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=4.56 $Y2=3.33
r65 43 54 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=3.6 $Y2=3.33
r66 42 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r67 40 53 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.76 $Y=3.33
+ $X2=3.595 $Y2=3.33
r68 40 42 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=3.76 $Y=3.33 $X2=4.08
+ $Y2=3.33
r69 39 56 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.33 $Y=3.33
+ $X2=4.495 $Y2=3.33
r70 39 42 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=4.33 $Y=3.33
+ $X2=4.08 $Y2=3.33
r71 38 54 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=3.6 $Y2=3.33
r72 37 38 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r73 35 51 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r74 34 37 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=1.2 $Y=3.33
+ $X2=3.12 $Y2=3.33
r75 34 35 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r76 32 50 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.91 $Y=3.33
+ $X2=0.745 $Y2=3.33
r77 32 34 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=0.91 $Y=3.33 $X2=1.2
+ $Y2=3.33
r78 31 53 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.43 $Y=3.33
+ $X2=3.595 $Y2=3.33
r79 31 37 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=3.43 $Y=3.33
+ $X2=3.12 $Y2=3.33
r80 29 51 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r81 28 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r82 26 50 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.58 $Y=3.33
+ $X2=0.745 $Y2=3.33
r83 26 28 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=0.58 $Y=3.33
+ $X2=0.24 $Y2=3.33
r84 24 38 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r85 24 35 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=1.2 $Y2=3.33
r86 20 56 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.495 $Y=3.245
+ $X2=4.495 $Y2=3.33
r87 20 22 27.5888 $w=3.28e-07 $l=7.9e-07 $layer=LI1_cond $X=4.495 $Y=3.245
+ $X2=4.495 $Y2=2.455
r88 16 53 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.595 $Y=3.245
+ $X2=3.595 $Y2=3.33
r89 16 18 27.5888 $w=3.28e-07 $l=7.9e-07 $layer=LI1_cond $X=3.595 $Y=3.245
+ $X2=3.595 $Y2=2.455
r90 12 15 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=0.745 $Y=2.105
+ $X2=0.745 $Y2=2.815
r91 10 50 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.745 $Y=3.245
+ $X2=0.745 $Y2=3.33
r92 10 15 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=0.745 $Y=3.245
+ $X2=0.745 $Y2=2.815
r93 3 22 300 $w=1.7e-07 $l=6.85912e-07 $layer=licon1_PDIFF $count=2 $X=4.345
+ $Y=1.84 $X2=4.495 $Y2=2.455
r94 2 18 300 $w=1.7e-07 $l=6.85912e-07 $layer=licon1_PDIFF $count=2 $X=3.445
+ $Y=1.84 $X2=3.595 $Y2=2.455
r95 1 15 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=0.62
+ $Y=1.96 $X2=0.745 $Y2=2.815
r96 1 12 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.62
+ $Y=1.96 $X2=0.745 $Y2=2.105
.ends

.subckt PM_SKY130_FD_SC_HS__A2BB2OI_2%A_424_368# 1 2 3 4 15 19 20 21 24 25 29 31
+ 33 35 40
c62 25 0 1.58807e-19 $X=3.96 $Y=2.035
c63 21 0 9.92294e-20 $X=3.105 $Y=2.12
r64 33 42 3.1514 $w=2.5e-07 $l=1.5e-07 $layer=LI1_cond $X=4.985 $Y=2.12
+ $X2=4.985 $Y2=1.97
r65 33 35 12.9074 $w=2.48e-07 $l=2.8e-07 $layer=LI1_cond $X=4.985 $Y=2.12
+ $X2=4.985 $Y2=2.4
r66 32 40 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.13 $Y=2.035
+ $X2=4.045 $Y2=2.035
r67 31 42 3.99177 $w=1.7e-07 $l=1.5411e-07 $layer=LI1_cond $X=4.86 $Y=2.035
+ $X2=4.985 $Y2=1.97
r68 31 32 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=4.86 $Y=2.035
+ $X2=4.13 $Y2=2.035
r69 27 40 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.045 $Y=2.12
+ $X2=4.045 $Y2=2.035
r70 27 29 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=4.045 $Y=2.12
+ $X2=4.045 $Y2=2.815
r71 26 38 3.99177 $w=1.7e-07 $l=1.5411e-07 $layer=LI1_cond $X=3.23 $Y=2.035
+ $X2=3.105 $Y2=1.97
r72 25 40 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.96 $Y=2.035
+ $X2=4.045 $Y2=2.035
r73 25 26 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=3.96 $Y=2.035
+ $X2=3.23 $Y2=2.035
r74 22 24 23.2793 $w=2.48e-07 $l=5.05e-07 $layer=LI1_cond $X=3.105 $Y=2.905
+ $X2=3.105 $Y2=2.4
r75 21 38 3.1514 $w=2.5e-07 $l=1.5e-07 $layer=LI1_cond $X=3.105 $Y=2.12
+ $X2=3.105 $Y2=1.97
r76 21 24 12.9074 $w=2.48e-07 $l=2.8e-07 $layer=LI1_cond $X=3.105 $Y=2.12
+ $X2=3.105 $Y2=2.4
r77 19 22 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=2.98 $Y=2.99
+ $X2=3.105 $Y2=2.905
r78 19 20 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=2.98 $Y=2.99
+ $X2=2.33 $Y2=2.99
r79 15 18 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=2.205 $Y=1.985
+ $X2=2.205 $Y2=2.815
r80 13 20 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=2.205 $Y=2.905
+ $X2=2.33 $Y2=2.99
r81 13 18 4.14879 $w=2.48e-07 $l=9e-08 $layer=LI1_cond $X=2.205 $Y=2.905
+ $X2=2.205 $Y2=2.815
r82 4 42 600 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=4.795
+ $Y=1.84 $X2=4.945 $Y2=1.985
r83 4 35 300 $w=1.7e-07 $l=6.30555e-07 $layer=licon1_PDIFF $count=2 $X=4.795
+ $Y=1.84 $X2=4.945 $Y2=2.4
r84 3 40 400 $w=1.7e-07 $l=3.4187e-07 $layer=licon1_PDIFF $count=1 $X=3.895
+ $Y=1.84 $X2=4.045 $Y2=2.115
r85 3 29 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=3.895
+ $Y=1.84 $X2=4.045 $Y2=2.815
r86 2 38 600 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=2.995
+ $Y=1.84 $X2=3.145 $Y2=1.985
r87 2 24 300 $w=1.7e-07 $l=6.30555e-07 $layer=licon1_PDIFF $count=2 $X=2.995
+ $Y=1.84 $X2=3.145 $Y2=2.4
r88 1 18 400 $w=1.7e-07 $l=1.03562e-06 $layer=licon1_PDIFF $count=1 $X=2.12
+ $Y=1.84 $X2=2.245 $Y2=2.815
r89 1 15 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=2.12
+ $Y=1.84 $X2=2.245 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HS__A2BB2OI_2%Y 1 2 3 12 14 15 18 20 22 25 29 30 37
c59 37 0 1.58807e-19 $X=3.235 $Y=1.195
c60 25 0 5.94286e-20 $X=3.63 $Y=0.95
c61 22 0 2.40437e-20 $X=3.465 $Y=1.065
r62 30 37 7.44484 $w=4.28e-07 $l=1.15e-07 $layer=LI1_cond $X=3.12 $Y=1.195
+ $X2=3.235 $Y2=1.195
r63 25 27 4.01609 $w=3.28e-07 $l=1.15e-07 $layer=LI1_cond $X=3.63 $Y=0.95
+ $X2=3.63 $Y2=1.065
r64 22 27 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.465 $Y=1.065
+ $X2=3.63 $Y2=1.065
r65 22 37 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=3.465 $Y=1.065
+ $X2=3.235 $Y2=1.065
r66 21 29 4.50329 $w=3e-07 $l=1.28e-07 $layer=LI1_cond $X=2.78 $Y=1.195
+ $X2=2.652 $Y2=1.195
r67 20 30 2.6801 $w=4.28e-07 $l=1e-07 $layer=LI1_cond $X=3.02 $Y=1.195 $X2=3.12
+ $Y2=1.195
r68 20 21 6.43224 $w=4.28e-07 $l=2.4e-07 $layer=LI1_cond $X=3.02 $Y=1.195
+ $X2=2.78 $Y2=1.195
r69 16 29 1.93381 $w=2.55e-07 $l=2.15e-07 $layer=LI1_cond $X=2.652 $Y=1.41
+ $X2=2.652 $Y2=1.195
r70 16 18 25.9865 $w=2.53e-07 $l=5.75e-07 $layer=LI1_cond $X=2.652 $Y=1.41
+ $X2=2.652 $Y2=1.985
r71 14 29 4.50329 $w=3e-07 $l=1.82784e-07 $layer=LI1_cond $X=2.525 $Y=1.065
+ $X2=2.652 $Y2=1.195
r72 14 15 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=2.525 $Y=1.065
+ $X2=2.25 $Y2=1.065
r73 10 15 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.165 $Y=0.98
+ $X2=2.25 $Y2=1.065
r74 10 12 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=2.165 $Y=0.98
+ $X2=2.165 $Y2=0.555
r75 3 18 300 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=2 $X=2.545
+ $Y=1.84 $X2=2.695 $Y2=1.985
r76 2 25 182 $w=1.7e-07 $l=6.4622e-07 $layer=licon1_NDIFF $count=1 $X=3.49
+ $Y=0.37 $X2=3.63 $Y2=0.95
r77 1 12 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.025
+ $Y=0.41 $X2=2.165 $Y2=0.555
.ends

.subckt PM_SKY130_FD_SC_HS__A2BB2OI_2%VGND 1 2 3 4 15 19 23 27 30 31 32 34 39 44
+ 57 58 61 64 67
r77 64 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r78 61 62 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r79 57 58 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r80 55 58 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=5.04
+ $Y2=0
r81 54 55 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r82 52 55 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=4.08
+ $Y2=0
r83 51 54 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=3.12 $Y=0 $X2=4.08
+ $Y2=0
r84 51 52 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r85 49 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.76 $Y=0 $X2=2.595
+ $Y2=0
r86 49 51 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=2.76 $Y=0 $X2=3.12
+ $Y2=0
r87 48 65 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.68
+ $Y2=0
r88 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r89 45 64 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.9 $Y=0 $X2=1.735
+ $Y2=0
r90 45 47 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=1.9 $Y=0 $X2=2.16
+ $Y2=0
r91 44 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.43 $Y=0 $X2=2.595
+ $Y2=0
r92 44 47 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=2.43 $Y=0 $X2=2.16
+ $Y2=0
r93 43 65 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=1.68
+ $Y2=0
r94 43 62 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r95 42 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r96 40 61 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.855 $Y=0 $X2=0.73
+ $Y2=0
r97 40 42 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.855 $Y=0 $X2=1.2
+ $Y2=0
r98 39 64 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.57 $Y=0 $X2=1.735
+ $Y2=0
r99 39 42 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=1.57 $Y=0 $X2=1.2
+ $Y2=0
r100 37 62 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r101 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r102 34 61 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.605 $Y=0 $X2=0.73
+ $Y2=0
r103 34 36 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=0.605 $Y=0
+ $X2=0.24 $Y2=0
r104 32 52 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r105 32 48 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=2.16
+ $Y2=0
r106 32 67 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r107 30 54 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=4.325 $Y=0 $X2=4.08
+ $Y2=0
r108 30 31 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.325 $Y=0 $X2=4.45
+ $Y2=0
r109 29 57 30.3369 $w=1.68e-07 $l=4.65e-07 $layer=LI1_cond $X=4.575 $Y=0
+ $X2=5.04 $Y2=0
r110 29 31 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.575 $Y=0 $X2=4.45
+ $Y2=0
r111 25 31 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.45 $Y=0.085
+ $X2=4.45 $Y2=0
r112 25 27 23.5098 $w=2.48e-07 $l=5.1e-07 $layer=LI1_cond $X=4.45 $Y=0.085
+ $X2=4.45 $Y2=0.595
r113 21 67 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.595 $Y=0.085
+ $X2=2.595 $Y2=0
r114 21 23 19.5566 $w=3.28e-07 $l=5.6e-07 $layer=LI1_cond $X=2.595 $Y=0.085
+ $X2=2.595 $Y2=0.645
r115 17 64 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.735 $Y=0.085
+ $X2=1.735 $Y2=0
r116 17 19 23.0489 $w=3.28e-07 $l=6.6e-07 $layer=LI1_cond $X=1.735 $Y=0.085
+ $X2=1.735 $Y2=0.745
r117 13 61 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.73 $Y=0.085
+ $X2=0.73 $Y2=0
r118 13 15 26.7367 $w=2.48e-07 $l=5.8e-07 $layer=LI1_cond $X=0.73 $Y=0.085
+ $X2=0.73 $Y2=0.665
r119 4 27 182 $w=1.7e-07 $l=2.86575e-07 $layer=licon1_NDIFF $count=1 $X=4.35
+ $Y=0.37 $X2=4.49 $Y2=0.595
r120 3 23 182 $w=1.7e-07 $l=2.96859e-07 $layer=licon1_NDIFF $count=1 $X=2.455
+ $Y=0.41 $X2=2.595 $Y2=0.645
r121 2 19 182 $w=1.7e-07 $l=3.19726e-07 $layer=licon1_NDIFF $count=1 $X=1.535
+ $Y=0.51 $X2=1.735 $Y2=0.745
r122 1 15 91 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_NDIFF $count=2 $X=0.645
+ $Y=0.51 $X2=0.77 $Y2=0.665
.ends

.subckt PM_SKY130_FD_SC_HS__A2BB2OI_2%A_615_74# 1 2 3 10 14 18 19 22
c34 14 0 1.6164e-19 $X=4.06 $Y=0.6
r35 20 22 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=4.92 $Y=1.01
+ $X2=4.92 $Y2=0.515
r36 18 20 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.755 $Y=1.095
+ $X2=4.92 $Y2=1.01
r37 18 19 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=4.755 $Y=1.095
+ $X2=4.145 $Y2=1.095
r38 15 19 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.06 $Y=1.01
+ $X2=4.145 $Y2=1.095
r39 15 17 2.93583 $w=1.68e-07 $l=4.5e-08 $layer=LI1_cond $X=4.06 $Y=1.01
+ $X2=4.06 $Y2=0.965
r40 14 25 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.06 $Y=0.6 $X2=4.06
+ $Y2=0.475
r41 14 17 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=4.06 $Y=0.6
+ $X2=4.06 $Y2=0.965
r42 10 25 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.975 $Y=0.475
+ $X2=4.06 $Y2=0.475
r43 10 12 35.7257 $w=2.48e-07 $l=7.75e-07 $layer=LI1_cond $X=3.975 $Y=0.475
+ $X2=3.2 $Y2=0.475
r44 3 22 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=4.78
+ $Y=0.37 $X2=4.92 $Y2=0.515
r45 2 25 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=3.92
+ $Y=0.37 $X2=4.06 $Y2=0.515
r46 2 17 182 $w=1.7e-07 $l=6.61306e-07 $layer=licon1_NDIFF $count=1 $X=3.92
+ $Y=0.37 $X2=4.06 $Y2=0.965
r47 1 12 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=3.075
+ $Y=0.37 $X2=3.2 $Y2=0.515
.ends

