# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_hs__a221oi_2
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_hs__a221oi_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.760000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.558000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.405000 1.430000 3.735000 1.950000 ;
        RECT 3.405000 1.950000 5.065000 2.120000 ;
        RECT 4.895000 1.430000 5.635000 1.780000 ;
        RECT 4.895000 1.780000 5.065000 1.950000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.558000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.965000 1.430000 4.675000 1.780000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.558000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.245000 1.430000 1.595000 1.680000 ;
        RECT 1.425000 1.680000 1.595000 1.950000 ;
        RECT 1.425000 1.950000 3.235000 2.120000 ;
        RECT 2.525000 1.550000 3.235000 1.950000 ;
        RECT 2.685000 1.430000 3.015000 1.550000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.558000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.945000 1.430000 2.275000 1.780000 ;
    END
  END B2
  PIN C1
    ANTENNAGATEAREA  0.558000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.585000 1.350000 0.915000 1.780000 ;
    END
  END C1
  PIN Y
    ANTENNADIFFAREA  1.172200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 0.350000 0.380000 1.010000 ;
        RECT 0.125000 1.010000 1.260000 1.090000 ;
        RECT 0.125000 1.090000 5.430000 1.180000 ;
        RECT 0.125000 1.180000 0.380000 1.950000 ;
        RECT 0.125000 1.950000 0.885000 2.120000 ;
        RECT 0.555000 2.120000 0.885000 2.735000 ;
        RECT 1.090000 0.350000 1.260000 1.010000 ;
        RECT 1.090000 1.180000 5.430000 1.260000 ;
        RECT 2.950000 0.350000 3.180000 1.090000 ;
        RECT 5.180000 0.350000 5.430000 1.090000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 5.760000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 5.760000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.760000 0.085000 ;
      RECT 0.000000  3.245000 5.760000 3.415000 ;
      RECT 0.105000  2.290000 0.355000 2.905000 ;
      RECT 0.105000  2.905000 3.165000 2.980000 ;
      RECT 0.105000  2.980000 2.265000 3.075000 ;
      RECT 0.560000  0.085000 0.910000 0.840000 ;
      RECT 1.085000  1.850000 1.255000 2.905000 ;
      RECT 1.440000  0.350000 1.770000 0.750000 ;
      RECT 1.440000  0.750000 2.780000 0.920000 ;
      RECT 1.455000  2.290000 5.035000 2.460000 ;
      RECT 1.455000  2.460000 1.815000 2.735000 ;
      RECT 1.940000  0.085000 2.280000 0.580000 ;
      RECT 2.015000  2.630000 3.165000 2.905000 ;
      RECT 2.450000  0.330000 2.780000 0.750000 ;
      RECT 3.350000  0.330000 4.030000 0.750000 ;
      RECT 3.350000  0.750000 5.000000 0.920000 ;
      RECT 3.355000  2.630000 3.605000 3.245000 ;
      RECT 3.805000  2.460000 4.135000 2.980000 ;
      RECT 4.200000  0.085000 4.530000 0.580000 ;
      RECT 4.335000  2.630000 4.505000 3.245000 ;
      RECT 4.700000  0.330000 5.000000 0.750000 ;
      RECT 4.705000  2.460000 5.035000 2.980000 ;
      RECT 5.235000  1.950000 5.485000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
  END
END sky130_fd_sc_hs__a221oi_2
