* File: sky130_fd_sc_hs__dfrbp_1.spice
* Created: Tue Sep  1 19:59:39 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hs__dfrbp_1.pex.spice"
.subckt sky130_fd_sc_hs__dfrbp_1  VNB VPB D RESET_B CLK VPWR Q_N Q VGND
* 
* VGND	VGND
* Q	Q
* Q_N	Q_N
* VPWR	VPWR
* CLK	CLK
* RESET_B	RESET_B
* D	D
* VPB	VPB
* VNB	VNB
MM1011 A_125_78# N_D_M1011_g N_A_38_78#_M1011_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.0504 AS=0.1197 PD=0.66 PS=1.41 NRD=18.564 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1033 N_VGND_M1033_d N_RESET_B_M1033_g A_125_78# VNB NLOWVT L=0.15 W=0.42
+ AD=0.1365 AS=0.0504 PD=1.49 PS=0.66 NRD=11.424 NRS=18.564 M=1 R=2.8 SA=75000.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1002 N_VGND_M1002_d N_CLK_M1002_g N_A_319_360#_M1002_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1554 AS=0.2109 PD=1.16 PS=2.05 NRD=11.34 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75000.8 A=0.111 P=1.78 MULT=1
MM1013 N_A_498_360#_M1013_d N_A_319_360#_M1013_g N_VGND_M1002_d VNB NLOWVT
+ L=0.15 W=0.74 AD=0.2109 AS=0.1554 PD=2.05 PS=1.16 NRD=0 NRS=11.34 M=1
+ R=4.93333 SA=75000.8 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1020 N_A_706_463#_M1020_d N_A_319_360#_M1020_g N_A_38_78#_M1020_s VNB NLOWVT
+ L=0.15 W=0.42 AD=0.0735 AS=0.1197 PD=0.77 PS=1.41 NRD=19.992 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75003.8 A=0.063 P=1.14 MULT=1
MM1018 A_832_118# N_A_498_360#_M1018_g N_A_706_463#_M1020_d VNB NLOWVT L=0.15
+ W=0.42 AD=0.0504 AS=0.0735 PD=0.66 PS=0.77 NRD=18.564 NRS=0 M=1 R=2.8
+ SA=75000.7 SB=75003.3 A=0.063 P=1.14 MULT=1
MM1006 A_910_118# N_A_841_401#_M1006_g A_832_118# VNB NLOWVT L=0.15 W=0.42
+ AD=0.0504 AS=0.0504 PD=0.66 PS=0.66 NRD=18.564 NRS=18.564 M=1 R=2.8 SA=75001.1
+ SB=75002.9 A=0.063 P=1.14 MULT=1
MM1022 N_VGND_M1022_d N_RESET_B_M1022_g A_910_118# VNB NLOWVT L=0.15 W=0.42
+ AD=0.126872 AS=0.0504 PD=1.00642 PS=0.66 NRD=70.584 NRS=18.564 M=1 R=2.8
+ SA=75001.5 SB=75002.5 A=0.063 P=1.14 MULT=1
MM1004 N_A_841_401#_M1004_d N_A_706_463#_M1004_g N_VGND_M1022_d VNB NLOWVT
+ L=0.15 W=0.64 AD=0.1611 AS=0.193328 PD=1.22 PS=1.53358 NRD=15.936 NRS=15.936
+ M=1 R=4.26667 SA=75001.5 SB=75002.4 A=0.096 P=1.58 MULT=1
MM1007 N_A_1224_74#_M1007_d N_A_498_360#_M1007_g N_A_841_401#_M1004_d VNB NLOWVT
+ L=0.15 W=0.64 AD=0.261434 AS=0.1611 PD=1.85962 PS=1.22 NRD=81.552 NRS=15.936
+ M=1 R=4.26667 SA=75002.1 SB=75001.8 A=0.096 P=1.58 MULT=1
MM1003 A_1434_74# N_A_319_360#_M1003_g N_A_1224_74#_M1007_d VNB NLOWVT L=0.15
+ W=0.42 AD=0.0504 AS=0.171566 PD=0.66 PS=1.22038 NRD=18.564 NRS=52.848 M=1
+ R=2.8 SA=75002.8 SB=75001.6 A=0.063 P=1.14 MULT=1
MM1029 N_VGND_M1029_d N_A_1482_48#_M1029_g A_1434_74# VNB NLOWVT L=0.15 W=0.42
+ AD=0.0861 AS=0.0504 PD=0.83 PS=0.66 NRD=18.564 NRS=18.564 M=1 R=2.8 SA=75003.2
+ SB=75001.2 A=0.063 P=1.14 MULT=1
MM1030 A_1624_74# N_RESET_B_M1030_g N_VGND_M1029_d VNB NLOWVT L=0.15 W=0.42
+ AD=0.0504 AS=0.0861 PD=0.66 PS=0.83 NRD=18.564 NRS=18.564 M=1 R=2.8 SA=75003.7
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1031 N_A_1482_48#_M1031_d N_A_1224_74#_M1031_g A_1624_74# VNB NLOWVT L=0.15
+ W=0.42 AD=0.1197 AS=0.0504 PD=1.41 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8
+ SA=75004.1 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1014 N_Q_N_M1014_d N_A_1224_74#_M1014_g N_VGND_M1014_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.2627 AS=0.2109 PD=2.19 PS=2.05 NRD=11.34 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75000.3 A=0.111 P=1.78 MULT=1
MM1012 N_VGND_M1012_d N_A_1224_74#_M1012_g N_A_2026_424#_M1012_s VNB NLOWVT
+ L=0.15 W=0.55 AD=0.104351 AS=0.15675 PD=0.929457 PS=1.67 NRD=13.632 NRS=0 M=1
+ R=3.66667 SA=75000.2 SB=75000.7 A=0.0825 P=1.4 MULT=1
MM1009 N_Q_M1009_d N_A_2026_424#_M1009_g N_VGND_M1012_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.140399 PD=2.05 PS=1.25054 NRD=0 NRS=1.62 M=1 R=4.93333
+ SA=75000.6 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1000 N_A_38_78#_M1000_d N_D_M1000_g N_VPWR_M1000_s VPB PSHORT L=0.15 W=0.42
+ AD=0.063 AS=0.1239 PD=0.72 PS=1.43 NRD=4.6886 NRS=4.6886 M=1 R=2.8 SA=75000.2
+ SB=75000.7 A=0.063 P=1.14 MULT=1
MM1001 N_VPWR_M1001_d N_RESET_B_M1001_g N_A_38_78#_M1000_d VPB PSHORT L=0.15
+ W=0.42 AD=0.1239 AS=0.063 PD=1.43 PS=0.72 NRD=4.6886 NRS=4.6886 M=1 R=2.8
+ SA=75000.7 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1017 N_VPWR_M1017_d N_CLK_M1017_g N_A_319_360#_M1017_s VPB PSHORT L=0.15
+ W=1.12 AD=0.168 AS=0.3304 PD=1.42 PS=2.83 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1023 N_A_498_360#_M1023_d N_A_319_360#_M1023_g N_VPWR_M1017_d VPB PSHORT
+ L=0.15 W=1.12 AD=0.3304 AS=0.168 PD=2.83 PS=1.42 NRD=1.7533 NRS=1.7533 M=1
+ R=7.46667 SA=75000.7 SB=75000.2 A=0.168 P=2.54 MULT=1
MM1021 N_A_706_463#_M1021_d N_A_498_360#_M1021_g N_A_38_78#_M1021_s VPB PSHORT
+ L=0.15 W=0.42 AD=0.063 AS=0.1239 PD=0.72 PS=1.43 NRD=4.6886 NRS=4.6886 M=1
+ R=2.8 SA=75000.2 SB=75001.7 A=0.063 P=1.14 MULT=1
MM1025 A_796_463# N_A_319_360#_M1025_g N_A_706_463#_M1021_d VPB PSHORT L=0.15
+ W=0.42 AD=0.0504 AS=0.063 PD=0.66 PS=0.72 NRD=30.4759 NRS=4.6886 M=1 R=2.8
+ SA=75000.7 SB=75001.2 A=0.063 P=1.14 MULT=1
MM1005 N_VPWR_M1005_d N_A_841_401#_M1005_g A_796_463# VPB PSHORT L=0.15 W=0.42
+ AD=0.139975 AS=0.0504 PD=1.155 PS=0.66 NRD=130.512 NRS=30.4759 M=1 R=2.8
+ SA=75001.1 SB=75000.8 A=0.063 P=1.14 MULT=1
MM1027 N_A_706_463#_M1027_d N_RESET_B_M1027_g N_VPWR_M1005_d VPB PSHORT L=0.15
+ W=0.42 AD=0.1176 AS=0.139975 PD=1.4 PS=1.155 NRD=7.0329 NRS=130.512 M=1 R=2.8
+ SA=75001.7 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1028 N_A_841_401#_M1028_d N_A_706_463#_M1028_g N_VPWR_M1028_s VPB PSHORT
+ L=0.15 W=1 AD=0.15 AS=0.295 PD=1.3 PS=2.59 NRD=1.9503 NRS=1.9503 M=1 R=6.66667
+ SA=75000.2 SB=75001.8 A=0.15 P=2.3 MULT=1
MM1032 N_A_1224_74#_M1032_d N_A_319_360#_M1032_g N_A_841_401#_M1028_d VPB PSHORT
+ L=0.15 W=1 AD=0.273028 AS=0.15 PD=2.25352 PS=1.3 NRD=26.5753 NRS=1.9503 M=1
+ R=6.66667 SA=75000.7 SB=75001.3 A=0.15 P=2.3 MULT=1
MM1015 A_1465_471# N_A_498_360#_M1015_g N_A_1224_74#_M1032_d VPB PSHORT L=0.15
+ W=0.42 AD=0.0567 AS=0.114672 PD=0.69 PS=0.946479 NRD=37.5088 NRS=68.0044 M=1
+ R=2.8 SA=75001.3 SB=75002.4 A=0.063 P=1.14 MULT=1
MM1026 N_VPWR_M1026_d N_A_1482_48#_M1026_g A_1465_471# VPB PSHORT L=0.15 W=0.42
+ AD=0.0756 AS=0.0567 PD=0.78 PS=0.69 NRD=16.4101 NRS=37.5088 M=1 R=2.8
+ SA=75001.7 SB=75002 A=0.063 P=1.14 MULT=1
MM1016 N_A_1482_48#_M1016_d N_RESET_B_M1016_g N_VPWR_M1026_d VPB PSHORT L=0.15
+ W=0.42 AD=0.063 AS=0.0756 PD=0.72 PS=0.78 NRD=4.6886 NRS=21.0987 M=1 R=2.8
+ SA=75002.2 SB=75001.5 A=0.063 P=1.14 MULT=1
MM1019 N_VPWR_M1019_d N_A_1224_74#_M1019_g N_A_1482_48#_M1016_d VPB PSHORT
+ L=0.15 W=0.42 AD=0.0943091 AS=0.063 PD=0.81 PS=0.72 NRD=37.5088 NRS=4.6886 M=1
+ R=2.8 SA=75002.6 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1024 N_Q_N_M1024_d N_A_1224_74#_M1024_g N_VPWR_M1019_d VPB PSHORT L=0.15
+ W=1.12 AD=0.6888 AS=0.251491 PD=3.47 PS=2.16 NRD=1.7533 NRS=1.7533 M=1
+ R=7.46667 SA=75001.3 SB=75000.5 A=0.168 P=2.54 MULT=1
MM1008 N_VPWR_M1008_d N_A_1224_74#_M1008_g N_A_2026_424#_M1008_s VPB PSHORT
+ L=0.15 W=0.84 AD=0.1644 AS=0.2478 PD=1.27286 PS=2.27 NRD=10.5395 NRS=2.3443
+ M=1 R=5.6 SA=75000.2 SB=75000.7 A=0.126 P=1.98 MULT=1
MM1010 N_Q_M1010_d N_A_2026_424#_M1010_g N_VPWR_M1008_d VPB PSHORT L=0.15 W=1.12
+ AD=0.3304 AS=0.2192 PD=2.83 PS=1.69714 NRD=1.7533 NRS=5.2599 M=1 R=7.46667
+ SA=75000.6 SB=75000.2 A=0.168 P=2.54 MULT=1
DX34_noxref VNB VPB NWDIODE A=22.4586 P=27.73
c_122 VNB 0 1.03779e-19 $X=0 $Y=0
c_236 VPB 0 1.13494e-19 $X=0 $Y=3.085
c_1690 A_1465_471# 0 1.04385e-19 $X=7.325 $Y=2.355
*
.include "sky130_fd_sc_hs__dfrbp_1.pxi.spice"
*
.ends
*
*
