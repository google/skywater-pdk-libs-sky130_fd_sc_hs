* File: sky130_fd_sc_hs__fah_2.pex.spice
* Created: Tue Sep  1 20:05:45 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HS__FAH_2%A_81_260# 1 2 7 9 12 18 23 26 29 32
c58 29 0 1.98792e-19 $X=1.31 $Y=1.465
c59 7 0 1.11723e-19 $X=0.495 $Y=1.765
r60 32 34 16.3735 $w=4.78e-07 $l=4.45e-07 $layer=LI1_cond $X=1.465 $Y=0.675
+ $X2=1.465 $Y2=1.12
r61 28 29 3.31764 $w=3.28e-07 $l=9.5e-08 $layer=LI1_cond $X=1.215 $Y=1.465
+ $X2=1.31 $Y2=1.465
r62 25 28 8.03218 $w=3.28e-07 $l=2.3e-07 $layer=LI1_cond $X=0.985 $Y=1.465
+ $X2=1.215 $Y2=1.465
r63 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.985
+ $Y=1.465 $X2=0.985 $Y2=1.465
r64 23 29 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.31 $Y=1.3 $X2=1.31
+ $Y2=1.465
r65 23 34 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=1.31 $Y=1.3 $X2=1.31
+ $Y2=1.12
r66 18 20 32.7294 $w=2.48e-07 $l=7.1e-07 $layer=LI1_cond $X=1.215 $Y=2.105
+ $X2=1.215 $Y2=2.815
r67 16 28 2.36532 $w=2.5e-07 $l=1.65e-07 $layer=LI1_cond $X=1.215 $Y=1.63
+ $X2=1.215 $Y2=1.465
r68 16 18 21.8964 $w=2.48e-07 $l=4.75e-07 $layer=LI1_cond $X=1.215 $Y=1.63
+ $X2=1.215 $Y2=2.105
r69 15 26 56.8299 $w=3.3e-07 $l=3.25e-07 $layer=POLY_cond $X=0.66 $Y=1.465
+ $X2=0.985 $Y2=1.465
r70 10 15 40.2336 $w=2.33e-07 $l=1.89658e-07 $layer=POLY_cond $X=0.585 $Y=1.3
+ $X2=0.532 $Y2=1.465
r71 10 12 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=0.585 $Y=1.3
+ $X2=0.585 $Y2=0.74
r72 7 15 68.1606 $w=2.33e-07 $l=3.17962e-07 $layer=POLY_cond $X=0.495 $Y=1.765
+ $X2=0.532 $Y2=1.465
r73 7 9 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.495 $Y=1.765
+ $X2=0.495 $Y2=2.4
r74 2 20 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=1.12
+ $Y=1.96 $X2=1.255 $Y2=2.815
r75 2 18 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=1.12
+ $Y=1.96 $X2=1.255 $Y2=2.105
r76 1 32 91 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_NDIFF $count=2 $X=1.395
+ $Y=0.525 $X2=1.54 $Y2=0.675
.ends

.subckt PM_SKY130_FD_SC_HS__FAH_2%A 2 3 5 6 8 10 11 13 14 16 17 24 26
c65 11 0 2.00363e-19 $X=1.99 $Y=1.885
c66 10 0 4.97865e-21 $X=1.99 $Y=1.795
c67 6 0 2.24154e-20 $X=1.825 $Y=1.29
c68 3 0 8.47849e-20 $X=1.48 $Y=1.885
r69 25 26 46.3382 $w=3.3e-07 $l=2.65e-07 $layer=POLY_cond $X=1.99 $Y=1.455
+ $X2=2.255 $Y2=1.455
r70 23 25 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=1.915 $Y=1.455
+ $X2=1.99 $Y2=1.455
r71 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.915
+ $Y=1.455 $X2=1.915 $Y2=1.455
r72 21 23 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=1.825 $Y=1.455
+ $X2=1.915 $Y2=1.455
r73 19 21 60.3271 $w=3.3e-07 $l=3.45e-07 $layer=POLY_cond $X=1.48 $Y=1.455
+ $X2=1.825 $Y2=1.455
r74 17 24 5.73629 $w=4.88e-07 $l=2.35e-07 $layer=LI1_cond $X=1.68 $Y=1.535
+ $X2=1.915 $Y2=1.535
r75 14 26 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.255 $Y=1.29
+ $X2=2.255 $Y2=1.455
r76 14 16 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=2.255 $Y=1.29
+ $X2=2.255 $Y2=0.845
r77 11 13 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=1.99 $Y=1.885
+ $X2=1.99 $Y2=2.46
r78 10 11 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=1.99 $Y=1.795 $X2=1.99
+ $Y2=1.885
r79 9 25 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.99 $Y=1.62
+ $X2=1.99 $Y2=1.455
r80 9 10 68.0242 $w=1.8e-07 $l=1.75e-07 $layer=POLY_cond $X=1.99 $Y=1.62
+ $X2=1.99 $Y2=1.795
r81 6 21 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.825 $Y=1.29
+ $X2=1.825 $Y2=1.455
r82 6 8 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=1.825 $Y=1.29
+ $X2=1.825 $Y2=0.845
r83 3 5 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=1.48 $Y=1.885
+ $X2=1.48 $Y2=2.46
r84 2 3 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=1.48 $Y=1.795 $X2=1.48
+ $Y2=1.885
r85 1 19 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.48 $Y=1.62
+ $X2=1.48 $Y2=1.455
r86 1 2 68.0242 $w=1.8e-07 $l=1.75e-07 $layer=POLY_cond $X=1.48 $Y=1.62 $X2=1.48
+ $Y2=1.795
.ends

.subckt PM_SKY130_FD_SC_HS__FAH_2%B 3 5 7 10 11 13 14 16 17 18 21 25 26 29 33 34
+ 36 39 40 41 44 45 46 48 50 52 53 54 60 61 69
c210 60 0 4.57584e-20 $X=2.64 $Y=1.665
c211 53 0 1.90307e-19 $X=4.5 $Y=0.68
c212 41 0 1.42825e-19 $X=5.435 $Y=1.005
c213 40 0 5.25489e-20 $X=5.875 $Y=1.005
c214 33 0 3.17652e-19 $X=4.505 $Y=1.44
c215 21 0 9.95712e-20 $X=7.125 $Y=0.74
c216 18 0 9.54589e-20 $X=6.745 $Y=1.315
c217 17 0 1.97436e-19 $X=7.05 $Y=1.315
c218 14 0 1.04626e-19 $X=6.655 $Y=1.765
c219 5 0 1.75179e-20 $X=3.56 $Y=2.045
r220 60 61 12.5413 $w=3.38e-07 $l=3.7e-07 $layer=LI1_cond $X=2.725 $Y=1.665
+ $X2=2.725 $Y2=2.035
r221 58 73 53.1237 $w=5.58e-07 $l=6.15e-07 $layer=POLY_cond $X=6.04 $Y=1.482
+ $X2=6.655 $Y2=1.482
r222 57 58 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.04
+ $Y=1.085 $X2=6.04 $Y2=1.085
r223 54 57 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=6.04 $Y=1.005 $X2=6.04
+ $Y2=1.085
r224 48 50 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=3.605 $Y=1.795
+ $X2=3.605 $Y2=1.63
r225 48 49 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.605
+ $Y=1.795 $X2=3.605 $Y2=1.795
r226 45 65 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.705 $Y=1.52
+ $X2=2.705 $Y2=1.355
r227 44 46 8.47192 $w=3.38e-07 $l=1.65e-07 $layer=LI1_cond $X=2.725 $Y=1.52
+ $X2=2.725 $Y2=1.355
r228 44 45 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.705
+ $Y=1.52 $X2=2.705 $Y2=1.52
r229 42 60 4.74535 $w=3.38e-07 $l=1.4e-07 $layer=LI1_cond $X=2.725 $Y=1.525
+ $X2=2.725 $Y2=1.665
r230 42 44 0.169477 $w=3.38e-07 $l=5e-09 $layer=LI1_cond $X=2.725 $Y=1.525
+ $X2=2.725 $Y2=1.52
r231 40 54 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.875 $Y=1.005
+ $X2=6.04 $Y2=1.005
r232 40 41 28.7059 $w=1.68e-07 $l=4.4e-07 $layer=LI1_cond $X=5.875 $Y=1.005
+ $X2=5.435 $Y2=1.005
r233 39 41 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.35 $Y=0.92
+ $X2=5.435 $Y2=1.005
r234 38 39 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=5.35 $Y=0.765
+ $X2=5.35 $Y2=0.92
r235 37 53 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=4.595 $Y=0.68
+ $X2=4.5 $Y2=0.68
r236 36 38 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.265 $Y=0.68
+ $X2=5.35 $Y2=0.765
r237 36 37 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.265 $Y=0.68
+ $X2=4.595 $Y2=0.68
r238 34 69 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.505 $Y=1.44
+ $X2=4.505 $Y2=1.275
r239 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.505
+ $Y=1.44 $X2=4.505 $Y2=1.44
r240 31 53 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=4.5 $Y=0.765
+ $X2=4.5 $Y2=0.68
r241 31 33 39.4019 $w=1.88e-07 $l=6.75e-07 $layer=LI1_cond $X=4.5 $Y=0.765
+ $X2=4.5 $Y2=1.44
r242 30 52 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.735 $Y=0.68
+ $X2=3.65 $Y2=0.68
r243 29 53 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=4.405 $Y=0.68
+ $X2=4.5 $Y2=0.68
r244 29 30 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.405 $Y=0.68
+ $X2=3.735 $Y2=0.68
r245 27 52 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.65 $Y=0.765
+ $X2=3.65 $Y2=0.68
r246 27 50 56.4332 $w=1.68e-07 $l=8.65e-07 $layer=LI1_cond $X=3.65 $Y=0.765
+ $X2=3.65 $Y2=1.63
r247 25 52 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.565 $Y=0.68
+ $X2=3.65 $Y2=0.68
r248 25 26 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.565 $Y=0.68
+ $X2=2.895 $Y2=0.68
r249 23 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.81 $Y=0.765
+ $X2=2.895 $Y2=0.68
r250 23 46 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=2.81 $Y=0.765
+ $X2=2.81 $Y2=1.355
r251 19 21 256.383 $w=1.5e-07 $l=5e-07 $layer=POLY_cond $X=7.125 $Y=1.24
+ $X2=7.125 $Y2=0.74
r252 18 73 36.977 $w=5.58e-07 $l=2.07169e-07 $layer=POLY_cond $X=6.745 $Y=1.315
+ $X2=6.655 $Y2=1.482
r253 17 19 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=7.05 $Y=1.315
+ $X2=7.125 $Y2=1.24
r254 17 18 156.394 $w=1.5e-07 $l=3.05e-07 $layer=POLY_cond $X=7.05 $Y=1.315
+ $X2=6.745 $Y2=1.315
r255 14 73 34.2028 $w=1.5e-07 $l=2.83e-07 $layer=POLY_cond $X=6.655 $Y=1.765
+ $X2=6.655 $Y2=1.482
r256 14 16 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=6.655 $Y=1.765
+ $X2=6.655 $Y2=2.4
r257 11 58 32.3925 $w=5.58e-07 $l=7.26701e-07 $layer=POLY_cond $X=5.665 $Y=2.045
+ $X2=6.04 $Y2=1.482
r258 11 13 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=5.665 $Y=2.045
+ $X2=5.665 $Y2=2.54
r259 10 69 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=4.445 $Y=0.845
+ $X2=4.445 $Y2=1.275
r260 5 49 52.2586 $w=2.99e-07 $l=2.7157e-07 $layer=POLY_cond $X=3.56 $Y=2.045
+ $X2=3.605 $Y2=1.795
r261 5 7 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=3.56 $Y=2.045
+ $X2=3.56 $Y2=2.54
r262 3 65 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=2.685 $Y=0.845
+ $X2=2.685 $Y2=1.355
.ends

.subckt PM_SKY130_FD_SC_HS__FAH_2%A_481_379# 1 2 7 9 10 11 13 14 16 17 18 20 21
+ 23 24 25 28 34 35 37 40 41 43 46 47 55
c167 37 0 8.21497e-20 $X=6.715 $Y=1.845
c168 34 0 1.61089e-19 $X=5.2 $Y=1.42
c169 24 0 1.90025e-19 $X=5.035 $Y=1.92
c170 17 0 1.56563e-19 $X=3.98 $Y=1.315
r171 55 57 4.88915 $w=3.28e-07 $l=1.4e-07 $layer=LI1_cond $X=6.88 $Y=1.845
+ $X2=6.88 $Y2=1.985
r172 46 49 3.54598 $w=2.58e-07 $l=8e-08 $layer=LI1_cond $X=5.235 $Y=1.765
+ $X2=5.235 $Y2=1.845
r173 46 47 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.2
+ $Y=1.765 $X2=5.2 $Y2=1.765
r174 41 43 13.7944 $w=3.28e-07 $l=3.95e-07 $layer=LI1_cond $X=7.34 $Y=1.19
+ $X2=7.34 $Y2=0.795
r175 40 55 2.96841 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=6.88 $Y=1.76
+ $X2=6.88 $Y2=1.845
r176 39 41 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=6.88 $Y=1.275
+ $X2=7.34 $Y2=1.275
r177 39 40 13.969 $w=3.28e-07 $l=4e-07 $layer=LI1_cond $X=6.88 $Y=1.36 $X2=6.88
+ $Y2=1.76
r178 38 49 3.22376 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=5.365 $Y=1.845
+ $X2=5.235 $Y2=1.845
r179 37 55 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.715 $Y=1.845
+ $X2=6.88 $Y2=1.845
r180 37 38 88.0749 $w=1.68e-07 $l=1.35e-06 $layer=LI1_cond $X=6.715 $Y=1.845
+ $X2=5.365 $Y2=1.845
r181 36 47 13.9889 $w=3.3e-07 $l=8e-08 $layer=POLY_cond $X=5.2 $Y=1.845 $X2=5.2
+ $Y2=1.765
r182 34 47 60.3271 $w=3.3e-07 $l=3.45e-07 $layer=POLY_cond $X=5.2 $Y=1.42
+ $X2=5.2 $Y2=1.765
r183 34 35 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.2 $Y=1.42
+ $X2=5.2 $Y2=1.255
r184 32 33 30.456 $w=1.82e-07 $l=1.15e-07 $layer=POLY_cond $X=4.055 $Y=1.945
+ $X2=4.17 $Y2=1.945
r185 29 31 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=3.155 $Y=1.315
+ $X2=3.445 $Y2=1.315
r186 28 35 131.747 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=5.29 $Y=0.845
+ $X2=5.29 $Y2=1.255
r187 25 33 25.4679 $w=1.82e-07 $l=1.01735e-07 $layer=POLY_cond $X=4.26 $Y=1.92
+ $X2=4.17 $Y2=1.945
r188 24 36 32.1775 $w=1.5e-07 $l=1.98997e-07 $layer=POLY_cond $X=5.035 $Y=1.92
+ $X2=5.2 $Y2=1.845
r189 24 25 397.394 $w=1.5e-07 $l=7.75e-07 $layer=POLY_cond $X=5.035 $Y=1.92
+ $X2=4.26 $Y2=1.92
r190 21 33 7.39479 $w=1.5e-07 $l=1e-07 $layer=POLY_cond $X=4.17 $Y=2.045
+ $X2=4.17 $Y2=1.945
r191 21 23 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=4.17 $Y=2.045
+ $X2=4.17 $Y2=2.54
r192 20 32 7.39479 $w=1.5e-07 $l=1e-07 $layer=POLY_cond $X=4.055 $Y=1.845
+ $X2=4.055 $Y2=1.945
r193 19 20 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=4.055 $Y=1.39
+ $X2=4.055 $Y2=1.845
r194 18 31 38.4574 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.52 $Y=1.315
+ $X2=3.445 $Y2=1.315
r195 17 19 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.98 $Y=1.315
+ $X2=4.055 $Y2=1.39
r196 17 18 235.872 $w=1.5e-07 $l=4.6e-07 $layer=POLY_cond $X=3.98 $Y=1.315
+ $X2=3.52 $Y2=1.315
r197 14 31 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.445 $Y=1.24
+ $X2=3.445 $Y2=1.315
r198 14 16 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=3.445 $Y=1.24
+ $X2=3.445 $Y2=0.845
r199 12 29 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.155 $Y=1.39
+ $X2=3.155 $Y2=1.315
r200 12 13 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=3.155 $Y=1.39
+ $X2=3.155 $Y2=1.895
r201 10 13 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.08 $Y=1.97
+ $X2=3.155 $Y2=1.895
r202 10 11 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=3.08 $Y=1.97
+ $X2=2.57 $Y2=1.97
r203 7 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.495 $Y=2.045
+ $X2=2.57 $Y2=1.97
r204 7 9 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=2.495 $Y=2.045
+ $X2=2.495 $Y2=2.54
r205 2 57 600 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=6.73
+ $Y=1.84 $X2=6.88 $Y2=1.985
r206 1 43 182 $w=1.7e-07 $l=4.90026e-07 $layer=licon1_NDIFF $count=1 $X=7.2
+ $Y=0.37 $X2=7.34 $Y2=0.795
.ends

.subckt PM_SKY130_FD_SC_HS__FAH_2%A_514_424# 1 2 7 9 12 14 16 19 21 26 27 30 31
+ 32 33 36 38 39 40 43 44 46 51 52 53 55 57 63 64 69 73 74 76 78 83 84
c246 69 0 2.00084e-19 $X=7.34 $Y=1.795
c247 44 0 3.062e-19 $X=8.575 $Y=1.39
c248 21 0 1.54605e-19 $X=3.065 $Y=2.555
c249 19 0 1.00227e-19 $X=10.285 $Y=0.715
r250 84 92 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=10.375 $Y=1.52
+ $X2=10.375 $Y2=1.355
r251 83 84 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.375
+ $Y=1.52 $X2=10.375 $Y2=1.52
r252 80 83 7.15912 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=10.17 $Y=1.52
+ $X2=10.375 $Y2=1.52
r253 76 79 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=9.41 $Y=1.795
+ $X2=9.41 $Y2=1.96
r254 76 78 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=9.41 $Y=1.795
+ $X2=9.41 $Y2=1.63
r255 76 77 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.475
+ $Y=1.795 $X2=9.475 $Y2=1.795
r256 69 72 8.51388 $w=2.88e-07 $l=1.65e-07 $layer=LI1_cond $X=7.36 $Y=1.795
+ $X2=7.36 $Y2=1.96
r257 69 70 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.34
+ $Y=1.795 $X2=7.34 $Y2=1.795
r258 64 66 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=6.31 $Y=2.185
+ $X2=6.31 $Y2=2.325
r259 62 63 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=3.285 $Y=2.555
+ $X2=3.45 $Y2=2.555
r260 60 62 4.71454 $w=3.28e-07 $l=1.35e-07 $layer=LI1_cond $X=3.15 $Y=2.555
+ $X2=3.285 $Y2=2.555
r261 57 59 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=3.23 $Y=1.02
+ $X2=3.23 $Y2=1.185
r262 55 80 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.17 $Y=1.355
+ $X2=10.17 $Y2=1.52
r263 54 55 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=10.17 $Y=0.765
+ $X2=10.17 $Y2=1.355
r264 52 54 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=10.085 $Y=0.68
+ $X2=10.17 $Y2=0.765
r265 52 53 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=10.085 $Y=0.68
+ $X2=9.415 $Y2=0.68
r266 51 79 61.6524 $w=1.68e-07 $l=9.45e-07 $layer=LI1_cond $X=9.49 $Y=2.905
+ $X2=9.49 $Y2=1.96
r267 48 53 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.33 $Y=0.765
+ $X2=9.415 $Y2=0.68
r268 48 78 56.4332 $w=1.68e-07 $l=8.65e-07 $layer=LI1_cond $X=9.33 $Y=0.765
+ $X2=9.33 $Y2=1.63
r269 47 74 7.13466 $w=1.7e-07 $l=1.28e-07 $layer=LI1_cond $X=8.735 $Y=2.99
+ $X2=8.607 $Y2=2.99
r270 46 51 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.405 $Y=2.99
+ $X2=9.49 $Y2=2.905
r271 46 47 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=9.405 $Y=2.99
+ $X2=8.735 $Y2=2.99
r272 44 88 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=8.575 $Y=1.39
+ $X2=8.575 $Y2=1.225
r273 43 44 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.575
+ $Y=1.39 $X2=8.575 $Y2=1.39
r274 41 74 0.067832 $w=2.55e-07 $l=8.5e-08 $layer=LI1_cond $X=8.607 $Y=2.905
+ $X2=8.607 $Y2=2.99
r275 41 43 68.4687 $w=2.53e-07 $l=1.515e-06 $layer=LI1_cond $X=8.607 $Y=2.905
+ $X2=8.607 $Y2=1.39
r276 39 74 7.13466 $w=1.7e-07 $l=1.27e-07 $layer=LI1_cond $X=8.48 $Y=2.99
+ $X2=8.607 $Y2=2.99
r277 39 40 71.4385 $w=1.68e-07 $l=1.095e-06 $layer=LI1_cond $X=8.48 $Y=2.99
+ $X2=7.385 $Y2=2.99
r278 38 40 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.3 $Y=2.905
+ $X2=7.385 $Y2=2.99
r279 37 73 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.3 $Y=2.41 $X2=7.3
+ $Y2=2.325
r280 37 38 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=7.3 $Y=2.41
+ $X2=7.3 $Y2=2.905
r281 36 73 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.3 $Y=2.24 $X2=7.3
+ $Y2=2.325
r282 36 72 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=7.3 $Y=2.24 $X2=7.3
+ $Y2=1.96
r283 34 66 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.395 $Y=2.325
+ $X2=6.31 $Y2=2.325
r284 33 73 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.215 $Y=2.325
+ $X2=7.3 $Y2=2.325
r285 33 34 53.4973 $w=1.68e-07 $l=8.2e-07 $layer=LI1_cond $X=7.215 $Y=2.325
+ $X2=6.395 $Y2=2.325
r286 31 64 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.225 $Y=2.185
+ $X2=6.31 $Y2=2.185
r287 31 32 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=6.225 $Y=2.185
+ $X2=5.555 $Y2=2.185
r288 29 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.47 $Y=2.27
+ $X2=5.555 $Y2=2.185
r289 29 30 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=5.47 $Y=2.27
+ $X2=5.47 $Y2=2.55
r290 27 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.385 $Y=2.635
+ $X2=5.47 $Y2=2.55
r291 27 63 126.241 $w=1.68e-07 $l=1.935e-06 $layer=LI1_cond $X=5.385 $Y=2.635
+ $X2=3.45 $Y2=2.635
r292 26 60 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.15 $Y=2.39
+ $X2=3.15 $Y2=2.555
r293 26 59 78.615 $w=1.68e-07 $l=1.205e-06 $layer=LI1_cond $X=3.15 $Y=2.39
+ $X2=3.15 $Y2=1.185
r294 21 60 2.96841 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=3.065 $Y=2.555
+ $X2=3.15 $Y2=2.555
r295 21 23 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=3.065 $Y=2.555
+ $X2=2.72 $Y2=2.555
r296 19 92 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=10.285 $Y=0.715
+ $X2=10.285 $Y2=1.355
r297 14 77 52.2586 $w=2.99e-07 $l=2.85044e-07 $layer=POLY_cond $X=9.4 $Y=2.045
+ $X2=9.475 $Y2=1.795
r298 14 16 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=9.4 $Y=2.045
+ $X2=9.4 $Y2=2.54
r299 12 88 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=8.625 $Y=0.715
+ $X2=8.625 $Y2=1.225
r300 7 70 50.1894 $w=3.66e-07 $l=3.02903e-07 $layer=POLY_cond $X=7.18 $Y=2.045
+ $X2=7.297 $Y2=1.795
r301 7 9 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=7.18 $Y=2.045
+ $X2=7.18 $Y2=2.54
r302 2 62 600 $w=1.7e-07 $l=9.0678e-07 $layer=licon1_PDIFF $count=1 $X=2.57
+ $Y=2.12 $X2=3.285 $Y2=2.555
r303 2 23 600 $w=1.7e-07 $l=5.04455e-07 $layer=licon1_PDIFF $count=1 $X=2.57
+ $Y=2.12 $X2=2.72 $Y2=2.555
r304 1 57 182 $w=1.7e-07 $l=6.9114e-07 $layer=licon1_NDIFF $count=1 $X=2.76
+ $Y=0.525 $X2=3.23 $Y2=1.02
.ends

.subckt PM_SKY130_FD_SC_HS__FAH_2%A_849_424# 1 2 7 9 10 11 12 14 15 18 19 20 23
+ 25 28 29 31 35 36 38 41 46 49 51 53 56 57 58 60 61 62 65 67 71 75 76 80
c209 80 0 2.97007e-19 $X=7.822 $Y=1.275
c210 71 0 1.90025e-19 $X=4.93 $Y=1.02
c211 53 0 2.83882e-20 $X=6.375 $Y=1.44
c212 23 0 1.66419e-19 $X=9.455 $Y=0.715
c213 7 0 1.77494e-19 $X=7.6 $Y=1.11
c214 1 0 1.90307e-19 $X=4.52 $Y=0.525
r215 76 78 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=5.62 $Y=1.345
+ $X2=5.62 $Y2=1.44
r216 73 74 5.66838 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=4.93 $Y=1.345
+ $X2=4.93 $Y2=1.43
r217 71 73 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=4.93 $Y=1.02
+ $X2=4.93 $Y2=1.345
r218 67 68 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=7.88
+ $Y=1.44 $X2=7.88 $Y2=1.44
r219 65 80 7.79447 $w=2.93e-07 $l=1.47e-07 $layer=LI1_cond $X=7.822 $Y=1.422
+ $X2=7.822 $Y2=1.275
r220 65 67 0.703186 $w=2.93e-07 $l=1.8e-08 $layer=LI1_cond $X=7.822 $Y=1.422
+ $X2=7.822 $Y2=1.44
r221 63 80 55.4545 $w=1.68e-07 $l=8.5e-07 $layer=LI1_cond $X=7.76 $Y=0.425
+ $X2=7.76 $Y2=1.275
r222 61 63 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.675 $Y=0.34
+ $X2=7.76 $Y2=0.425
r223 61 62 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=7.675 $Y=0.34
+ $X2=7.005 $Y2=0.34
r224 59 62 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.92 $Y=0.425
+ $X2=7.005 $Y2=0.34
r225 59 60 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=6.92 $Y=0.425
+ $X2=6.92 $Y2=0.85
r226 57 60 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.835 $Y=0.935
+ $X2=6.92 $Y2=0.85
r227 57 58 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=6.835 $Y=0.935
+ $X2=6.545 $Y2=0.935
r228 55 58 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.46 $Y=1.02
+ $X2=6.545 $Y2=0.935
r229 55 56 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=6.46 $Y=1.02
+ $X2=6.46 $Y2=1.355
r230 54 78 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.705 $Y=1.44
+ $X2=5.62 $Y2=1.44
r231 53 56 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.375 $Y=1.44
+ $X2=6.46 $Y2=1.355
r232 53 54 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=6.375 $Y=1.44
+ $X2=5.705 $Y2=1.44
r233 52 73 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.095 $Y=1.345
+ $X2=4.93 $Y2=1.345
r234 51 76 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.535 $Y=1.345
+ $X2=5.62 $Y2=1.345
r235 51 52 28.7059 $w=1.68e-07 $l=4.4e-07 $layer=LI1_cond $X=5.535 $Y=1.345
+ $X2=5.095 $Y2=1.345
r236 47 75 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.935 $Y=2.225
+ $X2=4.85 $Y2=2.225
r237 47 49 5.30124 $w=2.48e-07 $l=1.15e-07 $layer=LI1_cond $X=4.935 $Y=2.225
+ $X2=5.05 $Y2=2.225
r238 46 75 2.76166 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.85 $Y=2.1
+ $X2=4.85 $Y2=2.225
r239 46 74 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.85 $Y=2.1
+ $X2=4.85 $Y2=1.43
r240 39 41 133.319 $w=1.5e-07 $l=2.6e-07 $layer=POLY_cond $X=9.925 $Y=1.97
+ $X2=10.185 $Y2=1.97
r241 35 68 62.0758 $w=3.3e-07 $l=3.55e-07 $layer=POLY_cond $X=7.88 $Y=1.795
+ $X2=7.88 $Y2=1.44
r242 29 41 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=10.185 $Y=2.045
+ $X2=10.185 $Y2=1.97
r243 29 31 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=10.185 $Y=2.045
+ $X2=10.185 $Y2=2.54
r244 28 39 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=9.925 $Y=1.895
+ $X2=9.925 $Y2=1.97
r245 27 28 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=9.925 $Y=1.39
+ $X2=9.925 $Y2=1.895
r246 26 38 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=9.53 $Y=1.315
+ $X2=9.455 $Y2=1.315
r247 25 27 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=9.85 $Y=1.315
+ $X2=9.925 $Y2=1.39
r248 25 26 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=9.85 $Y=1.315
+ $X2=9.53 $Y2=1.315
r249 21 38 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=9.455 $Y=1.24
+ $X2=9.455 $Y2=1.315
r250 21 23 269.202 $w=1.5e-07 $l=5.25e-07 $layer=POLY_cond $X=9.455 $Y=1.24
+ $X2=9.455 $Y2=0.715
r251 19 38 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=9.38 $Y=1.315
+ $X2=9.455 $Y2=1.315
r252 19 20 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=9.38 $Y=1.315
+ $X2=9.1 $Y2=1.315
r253 17 20 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=9.025 $Y=1.39
+ $X2=9.1 $Y2=1.315
r254 17 18 207.67 $w=1.5e-07 $l=4.05e-07 $layer=POLY_cond $X=9.025 $Y=1.39
+ $X2=9.025 $Y2=1.795
r255 16 36 7.1379 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=8.46 $Y=1.87 $X2=8.37
+ $Y2=1.87
r256 15 18 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=8.95 $Y=1.87
+ $X2=9.025 $Y2=1.795
r257 15 16 251.255 $w=1.5e-07 $l=4.9e-07 $layer=POLY_cond $X=8.95 $Y=1.87
+ $X2=8.46 $Y2=1.87
r258 12 36 70.174 $w=1.8e-07 $l=1.75e-07 $layer=POLY_cond $X=8.37 $Y=2.045
+ $X2=8.37 $Y2=1.87
r259 12 14 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=8.37 $Y=2.045
+ $X2=8.37 $Y2=2.54
r260 11 35 32.1775 $w=1.5e-07 $l=1.98997e-07 $layer=POLY_cond $X=8.045 $Y=1.87
+ $X2=7.88 $Y2=1.795
r261 10 36 7.1379 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=8.28 $Y=1.87 $X2=8.37
+ $Y2=1.87
r262 10 11 120.5 $w=1.5e-07 $l=2.35e-07 $layer=POLY_cond $X=8.28 $Y=1.87
+ $X2=8.045 $Y2=1.87
r263 7 68 65.1981 $w=2.07e-07 $l=3.52987e-07 $layer=POLY_cond $X=7.6 $Y=1.11
+ $X2=7.88 $Y2=1.275
r264 7 9 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=7.6 $Y=1.11 $X2=7.6
+ $Y2=0.715
r265 2 49 300 $w=1.7e-07 $l=8.745e-07 $layer=licon1_PDIFF $count=2 $X=4.245
+ $Y=2.12 $X2=5.05 $Y2=2.265
r266 1 71 182 $w=1.7e-07 $l=6.69309e-07 $layer=licon1_NDIFF $count=1 $X=4.52
+ $Y=0.525 $X2=4.93 $Y2=1.02
.ends

.subckt PM_SKY130_FD_SC_HS__FAH_2%A_1689_424# 1 2 3 4 15 17 19 23 28 29 35 37 39
+ 41 43 44 46
c116 37 0 5.31033e-20 $X=11.24 $Y=2.075
r117 46 48 16.8178 $w=4.28e-07 $l=5.9e-07 $layer=LI1_cond $X=11.11 $Y=0.715
+ $X2=11.7 $Y2=0.715
r118 43 44 6.71605 $w=3.28e-07 $l=1.15e-07 $layer=LI1_cond $X=9.07 $Y=2.245
+ $X2=9.07 $Y2=2.13
r119 41 44 70.1337 $w=1.68e-07 $l=1.075e-06 $layer=LI1_cond $X=8.99 $Y=1.055
+ $X2=8.99 $Y2=2.13
r120 37 39 24.2013 $w=2.48e-07 $l=5.25e-07 $layer=LI1_cond $X=11.24 $Y=2.075
+ $X2=11.765 $Y2=2.075
r121 35 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=11.075
+ $Y=1.635 $X2=11.075 $Y2=1.635
r122 33 37 6.8199 $w=2.5e-07 $l=1.82071e-07 $layer=LI1_cond $X=11.11 $Y=1.95
+ $X2=11.24 $Y2=2.075
r123 33 35 13.9623 $w=2.58e-07 $l=3.15e-07 $layer=LI1_cond $X=11.11 $Y=1.95
+ $X2=11.11 $Y2=1.635
r124 32 46 3.65327 $w=2.6e-07 $l=3.4e-07 $layer=LI1_cond $X=11.11 $Y=1.055
+ $X2=11.11 $Y2=0.715
r125 32 35 25.7083 $w=2.58e-07 $l=5.8e-07 $layer=LI1_cond $X=11.11 $Y=1.055
+ $X2=11.11 $Y2=1.635
r126 31 46 7.41121 $w=4.28e-07 $l=2.6e-07 $layer=LI1_cond $X=10.85 $Y=0.715
+ $X2=11.11 $Y2=0.715
r127 30 31 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=10.85 $Y=0.425
+ $X2=10.85 $Y2=0.675
r128 28 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=10.765 $Y=0.34
+ $X2=10.85 $Y2=0.425
r129 28 29 110.257 $w=1.68e-07 $l=1.69e-06 $layer=LI1_cond $X=10.765 $Y=0.34
+ $X2=9.075 $Y2=0.34
r130 21 41 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=8.91 $Y=0.89
+ $X2=8.91 $Y2=1.055
r131 21 23 12.2229 $w=3.28e-07 $l=3.5e-07 $layer=LI1_cond $X=8.91 $Y=0.89
+ $X2=8.91 $Y2=0.54
r132 20 29 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=8.91 $Y=0.425
+ $X2=9.075 $Y2=0.34
r133 20 23 4.01609 $w=3.28e-07 $l=1.15e-07 $layer=LI1_cond $X=8.91 $Y=0.425
+ $X2=8.91 $Y2=0.54
r134 17 36 49.8163 $w=4.02e-07 $l=3.1225e-07 $layer=POLY_cond $X=10.87 $Y=1.885
+ $X2=11.01 $Y2=1.635
r135 17 19 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=10.87 $Y=1.885
+ $X2=10.87 $Y2=2.46
r136 13 36 39.6247 $w=4.02e-07 $l=2.29783e-07 $layer=POLY_cond $X=10.855 $Y=1.47
+ $X2=11.01 $Y2=1.635
r137 13 15 387.138 $w=1.5e-07 $l=7.55e-07 $layer=POLY_cond $X=10.855 $Y=1.47
+ $X2=10.855 $Y2=0.715
r138 4 39 600 $w=1.7e-07 $l=2.17428e-07 $layer=licon1_PDIFF $count=1 $X=11.615
+ $Y=1.96 $X2=11.765 $Y2=2.115
r139 3 43 300 $w=1.7e-07 $l=6.84653e-07 $layer=licon1_PDIFF $count=2 $X=8.445
+ $Y=2.12 $X2=9.07 $Y2=2.245
r140 2 48 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=11.56
+ $Y=0.395 $X2=11.7 $Y2=0.54
r141 1 23 91 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=2 $X=8.7
+ $Y=0.395 $X2=8.91 $Y2=0.54
.ends

.subckt PM_SKY130_FD_SC_HS__FAH_2%CI 3 5 6 8 9 10 11
c43 9 0 2.46841e-20 $X=11.505 $Y=1.11
c44 6 0 4.06256e-19 $X=11.54 $Y=1.885
r45 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=11.615
+ $Y=1.615 $X2=11.615 $Y2=1.615
r46 11 15 5.06376 $w=3.28e-07 $l=1.45e-07 $layer=LI1_cond $X=11.76 $Y=1.615
+ $X2=11.615 $Y2=1.615
r47 9 10 53.9552 $w=1.9e-07 $l=1.5e-07 $layer=POLY_cond $X=11.505 $Y=1.11
+ $X2=11.505 $Y2=1.26
r48 6 14 55.8646 $w=2.93e-07 $l=3.05205e-07 $layer=POLY_cond $X=11.54 $Y=1.885
+ $X2=11.615 $Y2=1.615
r49 6 8 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=11.54 $Y=1.885
+ $X2=11.54 $Y2=2.46
r50 5 14 38.5916 $w=2.93e-07 $l=2.05122e-07 $layer=POLY_cond $X=11.525 $Y=1.45
+ $X2=11.615 $Y2=1.615
r51 5 10 97.4255 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=11.525 $Y=1.45
+ $X2=11.525 $Y2=1.26
r52 3 9 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=11.485 $Y=0.715
+ $X2=11.485 $Y2=1.11
.ends

.subckt PM_SKY130_FD_SC_HS__FAH_2%A_1451_424# 1 2 7 9 10 12 13 15 16 18 19 22 24
+ 25 31 32 38 39
c132 39 0 1.08693e-19 $X=12.24 $Y=0.925
c133 38 0 7.1893e-20 $X=12.24 $Y=0.925
c134 31 0 1.39782e-19 $X=12.095 $Y=0.925
c135 24 0 1.77494e-19 $X=8.225 $Y=1.04
c136 22 0 5.88905e-20 $X=12.965 $Y=1.492
c137 13 0 2.25411e-19 $X=12.965 $Y=1.22
c138 7 0 1.78707e-19 $X=12.53 $Y=1.765
r139 42 43 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=12.25
+ $Y=1.385 $X2=12.25 $Y2=1.385
r140 39 43 16.0644 $w=3.28e-07 $l=4.6e-07 $layer=LI1_cond $X=12.25 $Y=0.925
+ $X2=12.25 $Y2=1.385
r141 38 39 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.24 $Y=0.925
+ $X2=12.24 $Y2=0.925
r142 35 50 10.6717 $w=4.63e-07 $l=4.05e-07 $layer=LI1_cond $X=8.285 $Y=0.925
+ $X2=8.285 $Y2=0.52
r143 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=0.925
+ $X2=8.4 $Y2=0.925
r144 32 34 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=8.545 $Y=0.925
+ $X2=8.4 $Y2=0.925
r145 31 38 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=12.095 $Y=0.925
+ $X2=12.24 $Y2=0.925
r146 31 32 4.39356 $w=1.4e-07 $l=3.55e-06 $layer=MET1_cond $X=12.095 $Y=0.925
+ $X2=8.545 $Y2=0.925
r147 25 27 1.58159 $w=6.03e-07 $l=8e-08 $layer=LI1_cond $X=8.225 $Y=2.432
+ $X2=8.145 $Y2=2.432
r148 24 35 8.16564 $w=4.63e-07 $l=1.41863e-07 $layer=LI1_cond $X=8.225 $Y=1.04
+ $X2=8.285 $Y2=0.925
r149 24 25 71.1123 $w=1.68e-07 $l=1.09e-06 $layer=LI1_cond $X=8.225 $Y=1.04
+ $X2=8.225 $Y2=2.13
r150 22 23 1.59956 $w=4.52e-07 $l=1.5e-08 $layer=POLY_cond $X=12.965 $Y=1.492
+ $X2=12.98 $Y2=1.492
r151 21 22 45.854 $w=4.52e-07 $l=4.3e-07 $layer=POLY_cond $X=12.535 $Y=1.492
+ $X2=12.965 $Y2=1.492
r152 20 21 0.533186 $w=4.52e-07 $l=5e-09 $layer=POLY_cond $X=12.53 $Y=1.492
+ $X2=12.535 $Y2=1.492
r153 19 42 33.2236 $w=3.3e-07 $l=1.9e-07 $layer=POLY_cond $X=12.44 $Y=1.385
+ $X2=12.25 $Y2=1.385
r154 19 20 13.1977 $w=4.52e-07 $l=1.45186e-07 $layer=POLY_cond $X=12.44 $Y=1.385
+ $X2=12.53 $Y2=1.492
r155 16 23 28.877 $w=1.5e-07 $l=2.73e-07 $layer=POLY_cond $X=12.98 $Y=1.765
+ $X2=12.98 $Y2=1.492
r156 16 18 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=12.98 $Y=1.765
+ $X2=12.98 $Y2=2.4
r157 13 22 28.877 $w=1.5e-07 $l=2.72e-07 $layer=POLY_cond $X=12.965 $Y=1.22
+ $X2=12.965 $Y2=1.492
r158 13 15 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=12.965 $Y=1.22
+ $X2=12.965 $Y2=0.74
r159 10 21 28.877 $w=1.5e-07 $l=2.72e-07 $layer=POLY_cond $X=12.535 $Y=1.22
+ $X2=12.535 $Y2=1.492
r160 10 12 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=12.535 $Y=1.22
+ $X2=12.535 $Y2=0.74
r161 7 20 28.877 $w=1.5e-07 $l=2.73e-07 $layer=POLY_cond $X=12.53 $Y=1.765
+ $X2=12.53 $Y2=1.492
r162 7 9 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=12.53 $Y=1.765
+ $X2=12.53 $Y2=2.4
r163 2 27 150 $w=1.7e-07 $l=9.50447e-07 $layer=licon1_PDIFF $count=4 $X=7.255
+ $Y=2.12 $X2=8.145 $Y2=2.245
r164 1 50 91 $w=1.7e-07 $l=5.64048e-07 $layer=licon1_NDIFF $count=2 $X=7.675
+ $Y=0.395 $X2=8.18 $Y2=0.52
.ends

.subckt PM_SKY130_FD_SC_HS__FAH_2%A_1895_424# 1 2 7 9 12 14 16 19 24 26 27 29 32
+ 34 37 38 42 49 55
c123 55 0 1.93712e-19 $X=13.89 $Y=1.532
c124 37 0 1.00227e-19 $X=9.91 $Y=2.1
r125 55 56 1.81203 $w=3.99e-07 $l=1.5e-08 $layer=POLY_cond $X=13.89 $Y=1.532
+ $X2=13.905 $Y2=1.532
r126 54 55 51.3409 $w=3.99e-07 $l=4.25e-07 $layer=POLY_cond $X=13.465 $Y=1.532
+ $X2=13.89 $Y2=1.532
r127 50 54 2.41604 $w=3.99e-07 $l=2e-08 $layer=POLY_cond $X=13.445 $Y=1.532
+ $X2=13.465 $Y2=1.532
r128 50 52 1.81203 $w=3.99e-07 $l=1.5e-08 $layer=POLY_cond $X=13.445 $Y=1.532
+ $X2=13.43 $Y2=1.532
r129 49 50 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=13.445
+ $Y=1.465 $X2=13.445 $Y2=1.465
r130 46 49 4.53993 $w=3.28e-07 $l=1.3e-07 $layer=LI1_cond $X=13.315 $Y=1.465
+ $X2=13.445 $Y2=1.465
r131 42 44 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=11.885 $Y=2.455
+ $X2=11.885 $Y2=2.685
r132 38 40 4.53993 $w=3.28e-07 $l=1.3e-07 $layer=LI1_cond $X=9.91 $Y=2.685
+ $X2=9.91 $Y2=2.815
r133 36 37 59.6952 $w=1.68e-07 $l=9.15e-07 $layer=LI1_cond $X=9.83 $Y=1.185
+ $X2=9.83 $Y2=2.1
r134 34 36 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=9.75 $Y=1.02
+ $X2=9.75 $Y2=1.185
r135 31 46 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=13.315 $Y=1.63
+ $X2=13.315 $Y2=1.465
r136 31 32 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=13.315 $Y=1.63
+ $X2=13.315 $Y2=2.37
r137 30 42 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=11.97 $Y=2.455
+ $X2=11.885 $Y2=2.455
r138 29 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=13.23 $Y=2.455
+ $X2=13.315 $Y2=2.37
r139 29 30 82.2032 $w=1.68e-07 $l=1.26e-06 $layer=LI1_cond $X=13.23 $Y=2.455
+ $X2=11.97 $Y2=2.455
r140 28 38 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.075 $Y=2.685
+ $X2=9.91 $Y2=2.685
r141 27 44 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=11.8 $Y=2.685
+ $X2=11.885 $Y2=2.685
r142 27 28 112.54 $w=1.68e-07 $l=1.725e-06 $layer=LI1_cond $X=11.8 $Y=2.685
+ $X2=10.075 $Y2=2.685
r143 26 37 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=9.91 $Y=2.265
+ $X2=9.91 $Y2=2.1
r144 24 38 2.96841 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=9.91 $Y=2.6
+ $X2=9.91 $Y2=2.685
r145 24 26 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=9.91 $Y=2.6
+ $X2=9.91 $Y2=2.265
r146 17 56 25.8008 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=13.905 $Y=1.3
+ $X2=13.905 $Y2=1.532
r147 17 19 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=13.905 $Y=1.3
+ $X2=13.905 $Y2=0.74
r148 14 55 25.8008 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=13.89 $Y=1.765
+ $X2=13.89 $Y2=1.532
r149 14 16 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=13.89 $Y=1.765
+ $X2=13.89 $Y2=2.4
r150 10 54 25.8008 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=13.465 $Y=1.3
+ $X2=13.465 $Y2=1.532
r151 10 12 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=13.465 $Y=1.3
+ $X2=13.465 $Y2=0.74
r152 7 52 25.8008 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=13.43 $Y=1.765
+ $X2=13.43 $Y2=1.532
r153 7 9 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=13.43 $Y=1.765
+ $X2=13.43 $Y2=2.4
r154 2 40 600 $w=1.7e-07 $l=8.862e-07 $layer=licon1_PDIFF $count=1 $X=9.475
+ $Y=2.12 $X2=9.91 $Y2=2.815
r155 2 26 600 $w=1.7e-07 $l=5.02295e-07 $layer=licon1_PDIFF $count=1 $X=9.475
+ $Y=2.12 $X2=9.91 $Y2=2.265
r156 1 34 182 $w=1.7e-07 $l=7.26722e-07 $layer=licon1_NDIFF $count=1 $X=9.53
+ $Y=0.395 $X2=9.75 $Y2=1.02
.ends

.subckt PM_SKY130_FD_SC_HS__FAH_2%VPWR 1 2 3 4 5 6 7 22 24 28 34 38 42 44 46 50
+ 52 57 65 73 78 83 92 95 98 105 108 112
c130 34 0 2.96008e-20 $X=6.43 $Y=2.745
r131 111 112 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=14.16 $Y=3.33
+ $X2=14.16 $Y2=3.33
r132 108 109 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.2 $Y=3.33
+ $X2=13.2 $Y2=3.33
r133 105 106 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.24 $Y=3.33
+ $X2=12.24 $Y2=3.33
r134 101 102 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.28 $Y=3.33
+ $X2=11.28 $Y2=3.33
r135 98 101 9.24987 $w=3.78e-07 $l=3.05e-07 $layer=LI1_cond $X=11.205 $Y=3.025
+ $X2=11.205 $Y2=3.33
r136 95 96 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r137 92 93 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r138 89 90 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r139 87 112 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=13.68 $Y=3.33
+ $X2=14.16 $Y2=3.33
r140 87 109 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=13.68 $Y=3.33
+ $X2=13.2 $Y2=3.33
r141 86 87 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.68 $Y=3.33
+ $X2=13.68 $Y2=3.33
r142 84 108 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=13.37 $Y=3.33
+ $X2=13.205 $Y2=3.33
r143 84 86 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=13.37 $Y=3.33
+ $X2=13.68 $Y2=3.33
r144 83 111 4.02656 $w=1.7e-07 $l=1.77e-07 $layer=LI1_cond $X=14.045 $Y=3.33
+ $X2=14.222 $Y2=3.33
r145 83 86 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=14.045 $Y=3.33
+ $X2=13.68 $Y2=3.33
r146 82 109 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.72 $Y=3.33
+ $X2=13.2 $Y2=3.33
r147 82 106 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.72 $Y=3.33
+ $X2=12.24 $Y2=3.33
r148 81 82 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.72 $Y=3.33
+ $X2=12.72 $Y2=3.33
r149 79 105 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12.47 $Y=3.33
+ $X2=12.305 $Y2=3.33
r150 79 81 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=12.47 $Y=3.33
+ $X2=12.72 $Y2=3.33
r151 78 108 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=13.04 $Y=3.33
+ $X2=13.205 $Y2=3.33
r152 78 81 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=13.04 $Y=3.33
+ $X2=12.72 $Y2=3.33
r153 77 106 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.76 $Y=3.33
+ $X2=12.24 $Y2=3.33
r154 77 102 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.76 $Y=3.33
+ $X2=11.28 $Y2=3.33
r155 76 77 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.76 $Y=3.33
+ $X2=11.76 $Y2=3.33
r156 74 101 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=11.395 $Y=3.33
+ $X2=11.205 $Y2=3.33
r157 74 76 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=11.395 $Y=3.33
+ $X2=11.76 $Y2=3.33
r158 73 105 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12.14 $Y=3.33
+ $X2=12.305 $Y2=3.33
r159 73 76 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=12.14 $Y=3.33
+ $X2=11.76 $Y2=3.33
r160 72 102 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.8 $Y=3.33
+ $X2=11.28 $Y2=3.33
r161 71 72 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=10.8 $Y=3.33
+ $X2=10.8 $Y2=3.33
r162 69 96 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=6.48 $Y2=3.33
r163 68 71 250.524 $w=1.68e-07 $l=3.84e-06 $layer=LI1_cond $X=6.96 $Y=3.33
+ $X2=10.8 $Y2=3.33
r164 68 69 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r165 66 95 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.595 $Y=3.33
+ $X2=6.43 $Y2=3.33
r166 66 68 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=6.595 $Y=3.33
+ $X2=6.96 $Y2=3.33
r167 65 101 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=11.015 $Y=3.33
+ $X2=11.205 $Y2=3.33
r168 65 71 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=11.015 $Y=3.33
+ $X2=10.8 $Y2=3.33
r169 64 96 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=3.33 $X2=6.48
+ $Y2=3.33
r170 63 64 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=6 $Y=3.33
+ $X2=6 $Y2=3.33
r171 61 64 1.07034 $w=4.9e-07 $l=3.84e-06 $layer=MET1_cond $X=2.16 $Y=3.33 $X2=6
+ $Y2=3.33
r172 61 93 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.68 $Y2=3.33
r173 60 63 250.524 $w=1.68e-07 $l=3.84e-06 $layer=LI1_cond $X=2.16 $Y=3.33 $X2=6
+ $Y2=3.33
r174 60 61 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r175 58 92 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.87 $Y=3.33
+ $X2=1.705 $Y2=3.33
r176 58 60 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=1.87 $Y=3.33
+ $X2=2.16 $Y2=3.33
r177 57 95 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.265 $Y=3.33
+ $X2=6.43 $Y2=3.33
r178 57 63 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=6.265 $Y=3.33
+ $X2=6 $Y2=3.33
r179 56 93 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=1.68 $Y2=3.33
r180 56 90 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.24 $Y2=3.33
r181 55 56 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r182 53 89 4.0754 $w=1.7e-07 $l=1.8e-07 $layer=LI1_cond $X=0.36 $Y=3.33 $X2=0.18
+ $Y2=3.33
r183 53 55 54.8021 $w=1.68e-07 $l=8.4e-07 $layer=LI1_cond $X=0.36 $Y=3.33
+ $X2=1.2 $Y2=3.33
r184 52 92 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.54 $Y=3.33
+ $X2=1.705 $Y2=3.33
r185 52 55 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=1.54 $Y=3.33
+ $X2=1.2 $Y2=3.33
r186 50 72 1.00344 $w=4.9e-07 $l=3.6e-06 $layer=MET1_cond $X=7.2 $Y=3.33
+ $X2=10.8 $Y2=3.33
r187 50 69 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=7.2 $Y=3.33
+ $X2=6.96 $Y2=3.33
r188 46 49 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=14.17 $Y=1.985
+ $X2=14.17 $Y2=2.815
r189 44 111 3.1166 $w=2.5e-07 $l=1.07912e-07 $layer=LI1_cond $X=14.17 $Y=3.245
+ $X2=14.222 $Y2=3.33
r190 44 49 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=14.17 $Y=3.245
+ $X2=14.17 $Y2=2.815
r191 40 108 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=13.205 $Y=3.245
+ $X2=13.205 $Y2=3.33
r192 40 42 15.3659 $w=3.28e-07 $l=4.4e-07 $layer=LI1_cond $X=13.205 $Y=3.245
+ $X2=13.205 $Y2=2.805
r193 36 105 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=12.305 $Y=3.245
+ $X2=12.305 $Y2=3.33
r194 36 38 15.3659 $w=3.28e-07 $l=4.4e-07 $layer=LI1_cond $X=12.305 $Y=3.245
+ $X2=12.305 $Y2=2.805
r195 32 95 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.43 $Y=3.245
+ $X2=6.43 $Y2=3.33
r196 32 34 17.4613 $w=3.28e-07 $l=5e-07 $layer=LI1_cond $X=6.43 $Y=3.245
+ $X2=6.43 $Y2=2.745
r197 28 31 24.4458 $w=3.28e-07 $l=7e-07 $layer=LI1_cond $X=1.705 $Y=2.115
+ $X2=1.705 $Y2=2.815
r198 26 92 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.705 $Y=3.245
+ $X2=1.705 $Y2=3.33
r199 26 31 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=1.705 $Y=3.245
+ $X2=1.705 $Y2=2.815
r200 22 89 3.10183 $w=2.55e-07 $l=1.07912e-07 $layer=LI1_cond $X=0.232 $Y=3.245
+ $X2=0.18 $Y2=3.33
r201 22 24 41.5783 $w=2.53e-07 $l=9.2e-07 $layer=LI1_cond $X=0.232 $Y=3.245
+ $X2=0.232 $Y2=2.325
r202 7 49 400 $w=1.7e-07 $l=1.05428e-06 $layer=licon1_PDIFF $count=1 $X=13.965
+ $Y=1.84 $X2=14.13 $Y2=2.815
r203 7 46 400 $w=1.7e-07 $l=2.26164e-07 $layer=licon1_PDIFF $count=1 $X=13.965
+ $Y=1.84 $X2=14.13 $Y2=1.985
r204 6 42 600 $w=1.7e-07 $l=1.03729e-06 $layer=licon1_PDIFF $count=1 $X=13.055
+ $Y=1.84 $X2=13.205 $Y2=2.805
r205 5 38 600 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_PDIFF $count=1 $X=12.17
+ $Y=2.65 $X2=12.305 $Y2=2.805
r206 4 98 600 $w=1.7e-07 $l=1.18791e-06 $layer=licon1_PDIFF $count=1 $X=10.945
+ $Y=1.96 $X2=11.205 $Y2=3.025
r207 3 34 600 $w=1.7e-07 $l=9.70155e-07 $layer=licon1_PDIFF $count=1 $X=6.295
+ $Y=1.84 $X2=6.43 $Y2=2.745
r208 2 31 400 $w=1.7e-07 $l=9.26971e-07 $layer=licon1_PDIFF $count=1 $X=1.555
+ $Y=1.96 $X2=1.705 $Y2=2.815
r209 2 28 400 $w=1.7e-07 $l=2.17428e-07 $layer=licon1_PDIFF $count=1 $X=1.555
+ $Y=1.96 $X2=1.705 $Y2=2.115
r210 1 24 300 $w=1.7e-07 $l=5.48361e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.84 $X2=0.27 $Y2=2.325
.ends

.subckt PM_SKY130_FD_SC_HS__FAH_2%A_114_368# 1 2 3 4 14 17 21 23 27 28 32 34 35
+ 41 45
c101 35 0 1.93813e-19 $X=0.385 $Y=1.295
c102 34 0 1.29241e-19 $X=3.935 $Y=1.295
r103 42 48 10.7189 $w=3.13e-07 $l=2.75e-07 $layer=LI1_cond $X=4.07 $Y=1.295
+ $X2=4.07 $Y2=1.02
r104 41 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=1.295
+ $X2=4.08 $Y2=1.295
r105 38 45 10.6381 $w=2.89e-07 $l=2.52e-07 $layer=LI1_cond $X=0.24 $Y=1.215
+ $X2=0.492 $Y2=1.215
r106 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=1.295
+ $X2=0.24 $Y2=1.295
r107 35 37 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=0.385 $Y=1.295
+ $X2=0.24 $Y2=1.295
r108 34 41 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.935 $Y=1.295
+ $X2=4.08 $Y2=1.295
r109 34 35 4.39356 $w=1.4e-07 $l=3.55e-06 $layer=MET1_cond $X=3.935 $Y=1.295
+ $X2=0.385 $Y2=1.295
r110 27 42 7.01145 $w=3.13e-07 $l=1.35647e-07 $layer=LI1_cond $X=4.025 $Y=1.41
+ $X2=4.07 $Y2=1.295
r111 27 28 46.9733 $w=1.68e-07 $l=7.2e-07 $layer=LI1_cond $X=4.025 $Y=1.41
+ $X2=4.025 $Y2=2.13
r112 23 28 7.14316 $w=2.5e-07 $l=1.62019e-07 $layer=LI1_cond $X=3.94 $Y=2.255
+ $X2=4.025 $Y2=2.13
r113 23 25 3.45733 $w=2.48e-07 $l=7.5e-08 $layer=LI1_cond $X=3.94 $Y=2.255
+ $X2=3.865 $Y2=2.255
r114 19 45 14.4796 $w=2.89e-07 $l=4.52895e-07 $layer=LI1_cond $X=0.835 $Y=0.96
+ $X2=0.492 $Y2=1.215
r115 19 21 19.7245 $w=2.58e-07 $l=4.45e-07 $layer=LI1_cond $X=0.835 $Y=0.96
+ $X2=0.835 $Y2=0.515
r116 17 32 28.8111 $w=3.28e-07 $l=8.25e-07 $layer=LI1_cond $X=0.72 $Y=2.815
+ $X2=0.72 $Y2=1.99
r117 14 32 14.8749 $w=1.68e-07 $l=2.28e-07 $layer=LI1_cond $X=0.492 $Y=1.905
+ $X2=0.72 $Y2=1.905
r118 13 45 0.205252 $w=3.15e-07 $l=2.55e-07 $layer=LI1_cond $X=0.492 $Y=1.47
+ $X2=0.492 $Y2=1.215
r119 13 14 12.8049 $w=3.13e-07 $l=3.5e-07 $layer=LI1_cond $X=0.492 $Y=1.47
+ $X2=0.492 $Y2=1.82
r120 4 25 600 $w=1.7e-07 $l=3.05205e-07 $layer=licon1_PDIFF $count=1 $X=3.635
+ $Y=2.12 $X2=3.865 $Y2=2.295
r121 3 32 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=0.57
+ $Y=1.84 $X2=0.72 $Y2=1.985
r122 3 17 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=0.57
+ $Y=1.84 $X2=0.72 $Y2=2.815
r123 2 48 182 $w=1.7e-07 $l=7.58123e-07 $layer=licon1_NDIFF $count=1 $X=3.52
+ $Y=0.525 $X2=4.07 $Y2=1.02
r124 1 21 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=0.66
+ $Y=0.37 $X2=0.8 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__FAH_2%A_413_392# 1 2 3 4 13 16 22 23 24 25 26 29 31
+ 33 34
c88 34 0 2.83882e-20 $X=5.77 $Y=0.34
c89 26 0 2.24154e-20 $X=2.555 $Y=0.34
c90 24 0 8.47849e-20 $X=2.385 $Y=2.975
c91 2 0 1.42825e-19 $X=5.365 $Y=0.525
r92 34 37 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=5.77 $Y=0.34
+ $X2=5.77 $Y2=0.665
r93 32 33 9.02376 $w=2.48e-07 $l=1.7e-07 $layer=LI1_cond $X=2.385 $Y=1.015
+ $X2=2.385 $Y2=1.185
r94 31 33 54.1497 $w=1.68e-07 $l=8.3e-07 $layer=LI1_cond $X=2.3 $Y=2.015 $X2=2.3
+ $Y2=1.185
r95 27 29 9.95292 $w=3.28e-07 $l=2.85e-07 $layer=LI1_cond $X=5.89 $Y=2.89
+ $X2=5.89 $Y2=2.605
r96 25 34 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.605 $Y=0.34
+ $X2=5.77 $Y2=0.34
r97 25 26 198.984 $w=1.68e-07 $l=3.05e-06 $layer=LI1_cond $X=5.605 $Y=0.34
+ $X2=2.555 $Y2=0.34
r98 23 27 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=5.725 $Y=2.975
+ $X2=5.89 $Y2=2.89
r99 23 24 217.904 $w=1.68e-07 $l=3.34e-06 $layer=LI1_cond $X=5.725 $Y=2.975
+ $X2=2.385 $Y2=2.975
r100 22 32 15.9037 $w=2.48e-07 $l=3.45e-07 $layer=LI1_cond $X=2.43 $Y=0.67
+ $X2=2.43 $Y2=1.015
r101 19 26 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=2.43 $Y=0.425
+ $X2=2.555 $Y2=0.34
r102 19 22 11.2939 $w=2.48e-07 $l=2.45e-07 $layer=LI1_cond $X=2.43 $Y=0.425
+ $X2=2.43 $Y2=0.67
r103 14 24 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.22 $Y=2.89
+ $X2=2.385 $Y2=2.975
r104 14 16 22.525 $w=3.28e-07 $l=6.45e-07 $layer=LI1_cond $X=2.22 $Y=2.89
+ $X2=2.22 $Y2=2.245
r105 13 31 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=2.22 $Y=2.18
+ $X2=2.22 $Y2=2.015
r106 13 16 2.26996 $w=3.28e-07 $l=6.5e-08 $layer=LI1_cond $X=2.22 $Y=2.18
+ $X2=2.22 $Y2=2.245
r107 4 29 600 $w=1.7e-07 $l=5.54955e-07 $layer=licon1_PDIFF $count=1 $X=5.74
+ $Y=2.12 $X2=5.89 $Y2=2.605
r108 3 16 300 $w=1.7e-07 $l=3.54119e-07 $layer=licon1_PDIFF $count=2 $X=2.065
+ $Y=1.96 $X2=2.22 $Y2=2.245
r109 2 37 182 $w=1.7e-07 $l=4.69814e-07 $layer=licon1_NDIFF $count=1 $X=5.365
+ $Y=0.525 $X2=5.77 $Y2=0.665
r110 1 22 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.33
+ $Y=0.525 $X2=2.47 $Y2=0.67
.ends

.subckt PM_SKY130_FD_SC_HS__FAH_2%A_2052_424# 1 2 7 13 16 19
c39 19 0 2.46841e-20 $X=10.725 $Y=1.1
c40 16 0 1.18856e-19 $X=10.725 $Y=2.13
r41 17 19 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=10.51 $Y=1.1
+ $X2=10.725 $Y2=1.1
r42 15 19 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.725 $Y=1.185
+ $X2=10.725 $Y2=1.1
r43 15 16 61.6524 $w=1.68e-07 $l=9.45e-07 $layer=LI1_cond $X=10.725 $Y=1.185
+ $X2=10.725 $Y2=2.13
r44 11 17 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.51 $Y=1.015
+ $X2=10.51 $Y2=1.1
r45 11 13 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=10.51 $Y=1.015
+ $X2=10.51 $Y2=0.825
r46 7 16 7.51767 $w=3e-07 $l=1.8775e-07 $layer=LI1_cond $X=10.64 $Y=2.28
+ $X2=10.725 $Y2=2.13
r47 7 9 5.57014 $w=2.98e-07 $l=1.45e-07 $layer=LI1_cond $X=10.64 $Y=2.28
+ $X2=10.495 $Y2=2.28
r48 2 9 600 $w=1.7e-07 $l=3.10403e-07 $layer=licon1_PDIFF $count=1 $X=10.26
+ $Y=2.12 $X2=10.495 $Y2=2.295
r49 1 13 182 $w=1.7e-07 $l=4.994e-07 $layer=licon1_NDIFF $count=1 $X=10.36
+ $Y=0.395 $X2=10.51 $Y2=0.825
.ends

.subckt PM_SKY130_FD_SC_HS__FAH_2%COUT 1 2 9 11 12 25
c22 11 0 1.93712e-19 $X=12.635 $Y=1.58
r23 16 25 1.78887 $w=3.33e-07 $l=5.2e-08 $layer=LI1_cond $X=12.752 $Y=1.717
+ $X2=12.752 $Y2=1.665
r24 11 25 0.584822 $w=3.33e-07 $l=1.7e-08 $layer=LI1_cond $X=12.752 $Y=1.648
+ $X2=12.752 $Y2=1.665
r25 11 23 4.13832 $w=3.33e-07 $l=9.8e-08 $layer=LI1_cond $X=12.752 $Y=1.648
+ $X2=12.752 $Y2=1.55
r26 11 12 9.52916 $w=3.33e-07 $l=2.77e-07 $layer=LI1_cond $X=12.752 $Y=1.733
+ $X2=12.752 $Y2=2.01
r27 11 16 0.550421 $w=3.33e-07 $l=1.6e-08 $layer=LI1_cond $X=12.752 $Y=1.733
+ $X2=12.752 $Y2=1.717
r28 9 23 47.7111 $w=2.48e-07 $l=1.035e-06 $layer=LI1_cond $X=12.71 $Y=0.515
+ $X2=12.71 $Y2=1.55
r29 2 12 600 $w=1.7e-07 $l=2.33238e-07 $layer=licon1_PDIFF $count=1 $X=12.605
+ $Y=1.84 $X2=12.755 $Y2=2.01
r30 1 9 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=12.61
+ $Y=0.37 $X2=12.75 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__FAH_2%SUM 1 2 9 11 13 19 20
c36 20 0 1.21085e-19 $X=14.16 $Y=1.295
c37 19 0 2.31759e-20 $X=13.722 $Y=1.82
c38 9 0 1.4004e-19 $X=13.685 $Y=0.52
r39 26 27 2.09656 $w=6.11e-07 $l=2.33675e-07 $layer=LI1_cond $X=13.685 $Y=0.965
+ $X2=13.79 $Y2=1.152
r40 20 27 7.38789 $w=6.11e-07 $l=3.7e-07 $layer=LI1_cond $X=14.16 $Y=1.152
+ $X2=13.79 $Y2=1.152
r41 17 27 8.43407 $w=1.7e-07 $l=3.53e-07 $layer=LI1_cond $X=13.79 $Y=1.505
+ $X2=13.79 $Y2=1.152
r42 17 19 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=13.79 $Y=1.505
+ $X2=13.79 $Y2=1.82
r43 13 15 31.3616 $w=3.03e-07 $l=8.3e-07 $layer=LI1_cond $X=13.722 $Y=1.985
+ $X2=13.722 $Y2=2.815
r44 11 19 7.98337 $w=3.03e-07 $l=1.52e-07 $layer=LI1_cond $X=13.722 $Y=1.972
+ $X2=13.722 $Y2=1.82
r45 11 13 0.491205 $w=3.03e-07 $l=1.3e-08 $layer=LI1_cond $X=13.722 $Y=1.972
+ $X2=13.722 $Y2=1.985
r46 7 26 0.698854 $w=6.11e-07 $l=1.81659e-07 $layer=LI1_cond $X=13.65 $Y=0.8
+ $X2=13.685 $Y2=0.965
r47 7 9 11.9513 $w=2.68e-07 $l=2.8e-07 $layer=LI1_cond $X=13.65 $Y=0.8 $X2=13.65
+ $Y2=0.52
r48 2 15 400 $w=1.7e-07 $l=1.04964e-06 $layer=licon1_PDIFF $count=1 $X=13.505
+ $Y=1.84 $X2=13.66 $Y2=2.815
r49 2 13 400 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_PDIFF $count=1 $X=13.505
+ $Y=1.84 $X2=13.66 $Y2=1.985
r50 1 26 182 $w=1.7e-07 $l=6.63551e-07 $layer=licon1_NDIFF $count=1 $X=13.54
+ $Y=0.37 $X2=13.685 $Y2=0.965
r51 1 9 182 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_NDIFF $count=1 $X=13.54
+ $Y=0.37 $X2=13.685 $Y2=0.52
.ends

.subckt PM_SKY130_FD_SC_HS__FAH_2%VGND 1 2 3 4 5 6 7 22 24 28 32 36 40 44 46 48
+ 51 52 54 55 56 65 79 83 88 97 100 103 107
r136 106 107 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=14.16 $Y=0
+ $X2=14.16 $Y2=0
r137 103 104 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.2 $Y=0
+ $X2=13.2 $Y2=0
r138 100 101 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.24 $Y=0
+ $X2=12.24 $Y2=0
r139 97 98 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=0 $X2=6.48
+ $Y2=0
r140 94 95 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r141 92 107 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=13.68 $Y=0
+ $X2=14.16 $Y2=0
r142 92 104 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=13.68 $Y=0
+ $X2=13.2 $Y2=0
r143 91 92 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.68 $Y=0
+ $X2=13.68 $Y2=0
r144 89 103 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=13.345 $Y=0
+ $X2=13.18 $Y2=0
r145 89 91 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=13.345 $Y=0
+ $X2=13.68 $Y2=0
r146 88 106 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=13.955 $Y=0
+ $X2=14.177 $Y2=0
r147 88 91 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=13.955 $Y=0
+ $X2=13.68 $Y2=0
r148 87 104 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.72 $Y=0
+ $X2=13.2 $Y2=0
r149 87 101 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.72 $Y=0
+ $X2=12.24 $Y2=0
r150 86 87 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.72 $Y=0
+ $X2=12.72 $Y2=0
r151 84 100 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12.405 $Y=0
+ $X2=12.24 $Y2=0
r152 84 86 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=12.405 $Y=0
+ $X2=12.72 $Y2=0
r153 83 103 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=13.015 $Y=0
+ $X2=13.18 $Y2=0
r154 83 86 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=13.015 $Y=0
+ $X2=12.72 $Y2=0
r155 82 101 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.76 $Y=0
+ $X2=12.24 $Y2=0
r156 81 82 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=11.76 $Y=0
+ $X2=11.76 $Y2=0
r157 79 100 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12.075 $Y=0
+ $X2=12.24 $Y2=0
r158 79 81 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=12.075 $Y=0
+ $X2=11.76 $Y2=0
r159 78 82 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=10.8 $Y=0
+ $X2=11.76 $Y2=0
r160 77 78 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=10.8 $Y=0
+ $X2=10.8 $Y2=0
r161 75 98 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=0 $X2=6.48
+ $Y2=0
r162 74 77 250.524 $w=1.68e-07 $l=3.84e-06 $layer=LI1_cond $X=6.96 $Y=0 $X2=10.8
+ $Y2=0
r163 74 75 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=6.96 $Y=0
+ $X2=6.96 $Y2=0
r164 72 97 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.665 $Y=0 $X2=6.5
+ $Y2=0
r165 72 74 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=6.665 $Y=0 $X2=6.96
+ $Y2=0
r166 71 98 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=0 $X2=6.48
+ $Y2=0
r167 70 71 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=6 $Y=0 $X2=6
+ $Y2=0
r168 68 71 1.07034 $w=4.9e-07 $l=3.84e-06 $layer=MET1_cond $X=2.16 $Y=0 $X2=6
+ $Y2=0
r169 67 70 250.524 $w=1.68e-07 $l=3.84e-06 $layer=LI1_cond $X=2.16 $Y=0 $X2=6
+ $Y2=0
r170 67 68 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=2.16 $Y=0
+ $X2=2.16 $Y2=0
r171 65 97 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.335 $Y=0 $X2=6.5
+ $Y2=0
r172 65 70 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=6.335 $Y=0 $X2=6
+ $Y2=0
r173 64 68 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r174 63 64 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r175 61 64 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r176 61 95 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r177 60 63 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r178 60 61 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r179 58 94 4.9356 $w=1.7e-07 $l=2.68e-07 $layer=LI1_cond $X=0.535 $Y=0 $X2=0.267
+ $Y2=0
r180 58 60 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=0.535 $Y=0
+ $X2=0.72 $Y2=0
r181 56 78 1.00344 $w=4.9e-07 $l=3.6e-06 $layer=MET1_cond $X=7.2 $Y=0 $X2=10.8
+ $Y2=0
r182 56 75 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=7.2 $Y=0 $X2=6.96
+ $Y2=0
r183 54 77 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=11.105 $Y=0
+ $X2=10.8 $Y2=0
r184 54 55 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=11.105 $Y=0
+ $X2=11.23 $Y2=0
r185 53 81 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=11.355 $Y=0
+ $X2=11.76 $Y2=0
r186 53 55 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=11.355 $Y=0
+ $X2=11.23 $Y2=0
r187 51 63 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=1.875 $Y=0
+ $X2=1.68 $Y2=0
r188 51 52 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.875 $Y=0 $X2=2
+ $Y2=0
r189 50 67 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=2.125 $Y=0 $X2=2.16
+ $Y2=0
r190 50 52 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.125 $Y=0 $X2=2
+ $Y2=0
r191 46 106 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=14.12 $Y=0.085
+ $X2=14.177 $Y2=0
r192 46 48 15.5405 $w=3.28e-07 $l=4.45e-07 $layer=LI1_cond $X=14.12 $Y=0.085
+ $X2=14.12 $Y2=0.53
r193 42 103 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=13.18 $Y=0.085
+ $X2=13.18 $Y2=0
r194 42 44 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=13.18 $Y=0.085
+ $X2=13.18 $Y2=0.515
r195 38 100 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=12.24 $Y=0.085
+ $X2=12.24 $Y2=0
r196 38 40 13.6198 $w=3.28e-07 $l=3.9e-07 $layer=LI1_cond $X=12.24 $Y=0.085
+ $X2=12.24 $Y2=0.475
r197 34 55 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=11.23 $Y=0.085
+ $X2=11.23 $Y2=0
r198 34 36 11.7549 $w=2.48e-07 $l=2.55e-07 $layer=LI1_cond $X=11.23 $Y=0.085
+ $X2=11.23 $Y2=0.34
r199 30 97 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.5 $Y=0.085 $X2=6.5
+ $Y2=0
r200 30 32 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=6.5 $Y=0.085
+ $X2=6.5 $Y2=0.515
r201 26 52 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2 $Y=0.085 $X2=2
+ $Y2=0
r202 26 28 27.1977 $w=2.48e-07 $l=5.9e-07 $layer=LI1_cond $X=2 $Y=0.085 $X2=2
+ $Y2=0.675
r203 22 94 3.13079 $w=3.65e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.352 $Y=0.085
+ $X2=0.267 $Y2=0
r204 22 24 18.1549 $w=3.63e-07 $l=5.75e-07 $layer=LI1_cond $X=0.352 $Y=0.085
+ $X2=0.352 $Y2=0.66
r205 7 48 182 $w=1.7e-07 $l=2.19089e-07 $layer=licon1_NDIFF $count=1 $X=13.98
+ $Y=0.37 $X2=14.12 $Y2=0.53
r206 6 44 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=13.04
+ $Y=0.37 $X2=13.18 $Y2=0.515
r207 5 40 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=12.105
+ $Y=0.33 $X2=12.24 $Y2=0.475
r208 4 36 182 $w=1.7e-07 $l=2.86182e-07 $layer=licon1_NDIFF $count=1 $X=10.93
+ $Y=0.395 $X2=11.19 $Y2=0.34
r209 3 32 182 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=1 $X=6.355
+ $Y=0.37 $X2=6.5 $Y2=0.515
r210 2 28 182 $w=1.7e-07 $l=2.08567e-07 $layer=licon1_NDIFF $count=1 $X=1.9
+ $Y=0.525 $X2=2.04 $Y2=0.675
r211 1 24 182 $w=1.7e-07 $l=3.61248e-07 $layer=licon1_NDIFF $count=1 $X=0.21
+ $Y=0.37 $X2=0.37 $Y2=0.66
.ends

