* File: sky130_fd_sc_hs__or4b_2.pex.spice
* Created: Tue Sep  1 20:21:28 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HS__OR4B_2%D_N 1 3 6 8 12
c26 6 0 2.621e-19 $X=0.51 $Y=0.835
c27 1 0 1.46046e-19 $X=0.505 $Y=1.765
r28 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.385
+ $Y=1.515 $X2=0.385 $Y2=1.515
r29 8 12 4.06745 $w=4.23e-07 $l=1.5e-07 $layer=LI1_cond $X=0.337 $Y=1.665
+ $X2=0.337 $Y2=1.515
r30 4 11 38.571 $w=3.25e-07 $l=2.12238e-07 $layer=POLY_cond $X=0.51 $Y=1.35
+ $X2=0.402 $Y2=1.515
r31 4 6 264.074 $w=1.5e-07 $l=5.15e-07 $layer=POLY_cond $X=0.51 $Y=1.35 $X2=0.51
+ $Y2=0.835
r32 1 11 51.1772 $w=3.25e-07 $l=2.97069e-07 $layer=POLY_cond $X=0.505 $Y=1.765
+ $X2=0.402 $Y2=1.515
r33 1 3 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=0.505 $Y=1.765
+ $X2=0.505 $Y2=2.26
.ends

.subckt PM_SKY130_FD_SC_HS__OR4B_2%A_190_48# 1 2 3 12 15 16 18 19 23 25 27 28 30
+ 31 32 35 41 43 47 55 57 59 60 62 63
c121 57 0 1.3676e-19 $X=2.34 $Y=1.045
c122 41 0 1.69342e-19 $X=3.54 $Y=0.615
c123 32 0 1.7764e-19 $X=1.745 $Y=1.045
r124 62 63 8.53881 $w=3.68e-07 $l=1.65e-07 $layer=LI1_cond $X=4.05 $Y=2.105
+ $X2=4.05 $Y2=1.94
r125 58 60 8.46729 $w=3.08e-07 $l=1.65e-07 $layer=LI1_cond $X=3.54 $Y=1.115
+ $X2=3.705 $Y2=1.115
r126 58 59 8.46729 $w=3.08e-07 $l=1.65e-07 $layer=LI1_cond $X=3.54 $Y=1.115
+ $X2=3.375 $Y2=1.115
r127 53 64 14.46 $w=3e-07 $l=9e-08 $layer=POLY_cond $X=1.555 $Y=1.465 $X2=1.555
+ $Y2=1.375
r128 52 55 3.31764 $w=3.28e-07 $l=9.5e-08 $layer=LI1_cond $X=1.565 $Y=1.465
+ $X2=1.66 $Y2=1.465
r129 52 53 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.565
+ $Y=1.465 $X2=1.565 $Y2=1.465
r130 49 63 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.15 $Y=1.27
+ $X2=4.15 $Y2=1.94
r131 45 62 0.622942 $w=3.68e-07 $l=2e-08 $layer=LI1_cond $X=4.05 $Y=2.125
+ $X2=4.05 $Y2=2.105
r132 45 47 21.4915 $w=3.68e-07 $l=6.9e-07 $layer=LI1_cond $X=4.05 $Y=2.125
+ $X2=4.05 $Y2=2.815
r133 43 49 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.065 $Y=1.185
+ $X2=4.15 $Y2=1.27
r134 43 60 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=4.065 $Y=1.185
+ $X2=3.705 $Y2=1.185
r135 39 58 0.331605 $w=3.3e-07 $l=1.55e-07 $layer=LI1_cond $X=3.54 $Y=0.96
+ $X2=3.54 $Y2=1.115
r136 39 41 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=3.54 $Y=0.96
+ $X2=3.54 $Y2=0.615
r137 38 57 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.505 $Y=1.045
+ $X2=2.34 $Y2=1.045
r138 38 59 56.7594 $w=1.68e-07 $l=8.7e-07 $layer=LI1_cond $X=2.505 $Y=1.045
+ $X2=3.375 $Y2=1.045
r139 33 57 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.34 $Y=0.96
+ $X2=2.34 $Y2=1.045
r140 33 35 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=2.34 $Y=0.96
+ $X2=2.34 $Y2=0.615
r141 31 57 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.175 $Y=1.045
+ $X2=2.34 $Y2=1.045
r142 31 32 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=2.175 $Y=1.045
+ $X2=1.745 $Y2=1.045
r143 30 55 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.66 $Y=1.3
+ $X2=1.66 $Y2=1.465
r144 29 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.66 $Y=1.13
+ $X2=1.745 $Y2=1.045
r145 29 30 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=1.66 $Y=1.13
+ $X2=1.66 $Y2=1.3
r146 25 53 60.2419 $w=3e-07 $l=3.30908e-07 $layer=POLY_cond $X=1.49 $Y=1.765
+ $X2=1.555 $Y2=1.465
r147 25 27 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.49 $Y=1.765
+ $X2=1.49 $Y2=2.4
r148 21 64 24.0919 $w=3e-07 $l=1.32288e-07 $layer=POLY_cond $X=1.455 $Y=1.3
+ $X2=1.555 $Y2=1.375
r149 21 23 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=1.455 $Y=1.3
+ $X2=1.455 $Y2=0.74
r150 20 28 6.66866 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=1.13 $Y=1.375
+ $X2=1.04 $Y2=1.375
r151 19 64 18.9685 $w=1.5e-07 $l=1.75e-07 $layer=POLY_cond $X=1.38 $Y=1.375
+ $X2=1.555 $Y2=1.375
r152 19 20 128.191 $w=1.5e-07 $l=2.5e-07 $layer=POLY_cond $X=1.38 $Y=1.375
+ $X2=1.13 $Y2=1.375
r153 16 18 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.04 $Y=1.765
+ $X2=1.04 $Y2=2.4
r154 15 16 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=1.04 $Y=1.675
+ $X2=1.04 $Y2=1.765
r155 14 28 18.8402 $w=1.65e-07 $l=7.5e-08 $layer=POLY_cond $X=1.04 $Y=1.45
+ $X2=1.04 $Y2=1.375
r156 14 15 87.4597 $w=1.8e-07 $l=2.25e-07 $layer=POLY_cond $X=1.04 $Y=1.45
+ $X2=1.04 $Y2=1.675
r157 10 28 18.8402 $w=1.65e-07 $l=8.21584e-08 $layer=POLY_cond $X=1.025 $Y=1.3
+ $X2=1.04 $Y2=1.375
r158 10 12 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=1.025 $Y=1.3
+ $X2=1.025 $Y2=0.74
r159 3 62 400 $w=1.7e-07 $l=3.65377e-07 $layer=licon1_PDIFF $count=1 $X=3.73
+ $Y=1.96 $X2=4.03 $Y2=2.105
r160 3 47 400 $w=1.7e-07 $l=9.93743e-07 $layer=licon1_PDIFF $count=1 $X=3.73
+ $Y=1.96 $X2=4.03 $Y2=2.815
r161 2 41 91 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=2 $X=3.355
+ $Y=0.47 $X2=3.54 $Y2=0.615
r162 1 35 91 $w=1.7e-07 $l=2.83373e-07 $layer=licon1_NDIFF $count=2 $X=2.12
+ $Y=0.47 $X2=2.34 $Y2=0.615
.ends

.subckt PM_SKY130_FD_SC_HS__OR4B_2%A 3 5 7 8 9 14
c39 3 0 1.08939e-19 $X=2.045 $Y=0.79
r40 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.11
+ $Y=1.515 $X2=2.11 $Y2=1.515
r41 8 9 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=2.11 $Y=1.665 $X2=2.11
+ $Y2=2.035
r42 8 14 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=2.11 $Y=1.665
+ $X2=2.11 $Y2=1.515
r43 5 13 75.1901 $w=2.72e-07 $l=4.05771e-07 $layer=POLY_cond $X=2.185 $Y=1.885
+ $X2=2.11 $Y2=1.515
r44 5 7 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=2.185 $Y=1.885
+ $X2=2.185 $Y2=2.46
r45 1 13 38.8629 $w=2.72e-07 $l=1.94808e-07 $layer=POLY_cond $X=2.045 $Y=1.35
+ $X2=2.11 $Y2=1.515
r46 1 3 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=2.045 $Y=1.35
+ $X2=2.045 $Y2=0.79
.ends

.subckt PM_SKY130_FD_SC_HS__OR4B_2%B 1 3 6 8 9
c34 1 0 1.3676e-19 $X=2.605 $Y=1.885
r35 8 9 13.969 $w=3.28e-07 $l=4e-07 $layer=LI1_cond $X=2.65 $Y=1.635 $X2=2.65
+ $Y2=2.035
r36 8 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.65
+ $Y=1.635 $X2=2.65 $Y2=1.635
r37 4 13 38.5562 $w=2.99e-07 $l=1.72337e-07 $layer=POLY_cond $X=2.635 $Y=1.47
+ $X2=2.65 $Y2=1.635
r38 4 6 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=2.635 $Y=1.47
+ $X2=2.635 $Y2=0.79
r39 1 13 52.2586 $w=2.99e-07 $l=2.7157e-07 $layer=POLY_cond $X=2.605 $Y=1.885
+ $X2=2.65 $Y2=1.635
r40 1 3 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=2.605 $Y=1.885
+ $X2=2.605 $Y2=2.46
.ends

.subckt PM_SKY130_FD_SC_HS__OR4B_2%C 1 3 6 8 9 10
c30 6 0 1.69342e-19 $X=3.28 $Y=0.79
r31 9 10 12.183 $w=3.48e-07 $l=3.7e-07 $layer=LI1_cond $X=3.18 $Y=2.035 $X2=3.18
+ $Y2=2.405
r32 8 9 13.1708 $w=3.48e-07 $l=4e-07 $layer=LI1_cond $X=3.18 $Y=1.635 $X2=3.18
+ $Y2=2.035
r33 8 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.19
+ $Y=1.635 $X2=3.19 $Y2=1.635
r34 4 15 38.5562 $w=2.99e-07 $l=2.05122e-07 $layer=POLY_cond $X=3.28 $Y=1.47
+ $X2=3.19 $Y2=1.635
r35 4 6 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=3.28 $Y=1.47 $X2=3.28
+ $Y2=0.79
r36 1 15 52.2586 $w=2.99e-07 $l=2.85044e-07 $layer=POLY_cond $X=3.115 $Y=1.885
+ $X2=3.19 $Y2=1.635
r37 1 3 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=3.115 $Y=1.885
+ $X2=3.115 $Y2=2.46
.ends

.subckt PM_SKY130_FD_SC_HS__OR4B_2%A_27_368# 1 2 7 9 12 16 18 19 21 22 23 25 26
+ 27 29 36
r96 36 37 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.73
+ $Y=1.605 $X2=3.73 $Y2=1.605
r97 33 36 4.1907 $w=3.28e-07 $l=1.2e-07 $layer=LI1_cond $X=3.61 $Y=1.605
+ $X2=3.73 $Y2=1.605
r98 31 32 10.1828 $w=6.29e-07 $l=5.25e-07 $layer=LI1_cond $X=0.28 $Y=2.325
+ $X2=0.805 $Y2=2.325
r99 28 33 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.61 $Y=1.77
+ $X2=3.61 $Y2=1.605
r100 28 29 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=3.61 $Y=1.77
+ $X2=3.61 $Y2=2.69
r101 26 29 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.525 $Y=2.775
+ $X2=3.61 $Y2=2.69
r102 26 27 69.1551 $w=1.68e-07 $l=1.06e-06 $layer=LI1_cond $X=3.525 $Y=2.775
+ $X2=2.465 $Y2=2.775
r103 25 27 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.38 $Y=2.69
+ $X2=2.465 $Y2=2.775
r104 24 25 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=2.38 $Y=2.49 $X2=2.38
+ $Y2=2.69
r105 23 32 9.00042 $w=6.29e-07 $l=1.18427e-07 $layer=LI1_cond $X=0.89 $Y=2.405
+ $X2=0.805 $Y2=2.325
r106 22 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.295 $Y=2.405
+ $X2=2.38 $Y2=2.49
r107 22 23 91.6631 $w=1.68e-07 $l=1.405e-06 $layer=LI1_cond $X=2.295 $Y=2.405
+ $X2=0.89 $Y2=2.405
r108 21 32 8.62214 $w=1.7e-07 $l=3.75e-07 $layer=LI1_cond $X=0.805 $Y=1.95
+ $X2=0.805 $Y2=2.325
r109 20 21 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=0.805 $Y=1.18
+ $X2=0.805 $Y2=1.95
r110 18 20 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.72 $Y=1.095
+ $X2=0.805 $Y2=1.18
r111 18 19 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=0.72 $Y=1.095
+ $X2=0.46 $Y2=1.095
r112 14 19 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.295 $Y=1.01
+ $X2=0.46 $Y2=1.095
r113 14 16 6.11144 $w=3.28e-07 $l=1.75e-07 $layer=LI1_cond $X=0.295 $Y=1.01
+ $X2=0.295 $Y2=0.835
r114 10 37 38.6072 $w=2.91e-07 $l=1.77059e-07 $layer=POLY_cond $X=3.755 $Y=1.44
+ $X2=3.73 $Y2=1.605
r115 10 12 333.298 $w=1.5e-07 $l=6.5e-07 $layer=POLY_cond $X=3.755 $Y=1.44
+ $X2=3.755 $Y2=0.79
r116 7 37 57.6553 $w=2.91e-07 $l=3.15278e-07 $layer=POLY_cond $X=3.655 $Y=1.885
+ $X2=3.73 $Y2=1.605
r117 7 9 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=3.655 $Y=1.885
+ $X2=3.655 $Y2=2.46
r118 2 31 300 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.115
r119 1 16 182 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_NDIFF $count=1 $X=0.15
+ $Y=0.56 $X2=0.295 $Y2=0.835
.ends

.subckt PM_SKY130_FD_SC_HS__OR4B_2%VPWR 1 2 11 13 15 25 26 29 32
r45 29 30 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r46 25 26 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r47 22 25 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=2.16 $Y=3.33
+ $X2=4.08 $Y2=3.33
r48 20 22 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=2.125 $Y=3.33
+ $X2=2.16 $Y2=3.33
r49 19 36 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=1.68 $Y2=3.33
r50 19 30 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r51 18 19 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r52 16 29 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.98 $Y=3.33
+ $X2=0.815 $Y2=3.33
r53 16 18 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=0.98 $Y=3.33 $X2=1.2
+ $Y2=3.33
r54 15 20 8.04321 $w=1.7e-07 $l=2.88e-07 $layer=LI1_cond $X=1.837 $Y=3.33
+ $X2=2.125 $Y2=3.33
r55 15 36 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r56 15 32 10.7127 $w=5.73e-07 $l=5.15e-07 $layer=LI1_cond $X=1.837 $Y=3.33
+ $X2=1.837 $Y2=2.815
r57 15 18 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=1.55 $Y=3.33 $X2=1.2
+ $Y2=3.33
r58 13 26 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=4.08 $Y2=3.33
r59 13 36 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.68 $Y2=3.33
r60 13 22 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r61 9 29 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.815 $Y=3.245
+ $X2=0.815 $Y2=3.33
r62 9 11 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=0.815 $Y=3.245
+ $X2=0.815 $Y2=2.78
r63 2 32 600 $w=1.7e-07 $l=1.10176e-06 $layer=licon1_PDIFF $count=1 $X=1.565
+ $Y=1.84 $X2=1.835 $Y2=2.815
r64 1 11 600 $w=1.7e-07 $l=1.05095e-06 $layer=licon1_PDIFF $count=1 $X=0.58
+ $Y=1.84 $X2=0.815 $Y2=2.78
.ends

.subckt PM_SKY130_FD_SC_HS__OR4B_2%X 1 2 9 13 14 18
c38 18 0 1.42209e-19 $X=1.245 $Y=1.82
c39 14 0 1.46046e-19 $X=1.2 $Y=2.035
c40 13 0 2.2883e-19 $X=1.232 $Y=1.13
r41 14 18 8.53881 $w=3.68e-07 $l=1.65e-07 $layer=LI1_cond $X=1.245 $Y=1.985
+ $X2=1.245 $Y2=1.82
r42 13 18 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.145 $Y=1.13
+ $X2=1.145 $Y2=1.82
r43 7 13 8.71323 $w=3.43e-07 $l=1.72e-07 $layer=LI1_cond $X=1.232 $Y=0.958
+ $X2=1.232 $Y2=1.13
r44 7 9 14.798 $w=3.43e-07 $l=4.43e-07 $layer=LI1_cond $X=1.232 $Y=0.958
+ $X2=1.232 $Y2=0.515
r45 2 14 600 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=1.115
+ $Y=1.84 $X2=1.265 $Y2=1.985
r46 1 9 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.1 $Y=0.37
+ $X2=1.24 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__OR4B_2%VGND 1 2 3 4 17 21 25 27 29 31 33 38 43 49 52
+ 55 59
r61 58 59 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r62 55 56 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r63 52 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r64 49 50 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r65 47 59 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.08
+ $Y2=0
r66 47 56 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=3.12
+ $Y2=0
r67 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r68 44 55 11.5608 $w=1.7e-07 $l=2.6e-07 $layer=LI1_cond $X=3.205 $Y=0 $X2=2.945
+ $Y2=0
r69 44 46 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=3.205 $Y=0 $X2=3.6
+ $Y2=0
r70 43 58 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=3.875 $Y=0 $X2=4.097
+ $Y2=0
r71 43 46 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=3.875 $Y=0 $X2=3.6
+ $Y2=0
r72 42 56 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r73 41 42 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r74 39 52 10.1275 $w=1.7e-07 $l=2.1e-07 $layer=LI1_cond $X=1.995 $Y=0 $X2=1.785
+ $Y2=0
r75 39 41 42.0802 $w=1.68e-07 $l=6.45e-07 $layer=LI1_cond $X=1.995 $Y=0 $X2=2.64
+ $Y2=0
r76 38 55 11.5608 $w=1.7e-07 $l=2.6e-07 $layer=LI1_cond $X=2.685 $Y=0 $X2=2.945
+ $Y2=0
r77 38 41 2.93583 $w=1.68e-07 $l=4.5e-08 $layer=LI1_cond $X=2.685 $Y=0 $X2=2.64
+ $Y2=0
r78 37 53 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=1.68
+ $Y2=0
r79 37 50 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r80 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r81 34 49 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.89 $Y=0 $X2=0.765
+ $Y2=0
r82 34 36 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=0.89 $Y=0 $X2=1.2
+ $Y2=0
r83 33 52 10.1275 $w=1.7e-07 $l=2.1e-07 $layer=LI1_cond $X=1.575 $Y=0 $X2=1.785
+ $Y2=0
r84 33 36 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=1.575 $Y=0 $X2=1.2
+ $Y2=0
r85 31 42 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r86 31 53 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.68
+ $Y2=0
r87 27 58 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=4.04 $Y=0.085
+ $X2=4.097 $Y2=0
r88 27 29 21.1281 $w=3.28e-07 $l=6.05e-07 $layer=LI1_cond $X=4.04 $Y=0.085
+ $X2=4.04 $Y2=0.69
r89 23 55 2.17428 $w=5.2e-07 $l=8.5e-08 $layer=LI1_cond $X=2.945 $Y=0.085
+ $X2=2.945 $Y2=0
r90 23 25 12.1908 $w=5.18e-07 $l=5.3e-07 $layer=LI1_cond $X=2.945 $Y=0.085
+ $X2=2.945 $Y2=0.615
r91 19 52 1.60615 $w=4.2e-07 $l=8.5e-08 $layer=LI1_cond $X=1.785 $Y=0.085
+ $X2=1.785 $Y2=0
r92 19 21 14.5427 $w=4.18e-07 $l=5.3e-07 $layer=LI1_cond $X=1.785 $Y=0.085
+ $X2=1.785 $Y2=0.615
r93 15 49 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.765 $Y=0.085
+ $X2=0.765 $Y2=0
r94 15 17 23.5098 $w=2.48e-07 $l=5.1e-07 $layer=LI1_cond $X=0.765 $Y=0.085
+ $X2=0.765 $Y2=0.595
r95 4 29 182 $w=1.7e-07 $l=3.07571e-07 $layer=licon1_NDIFF $count=1 $X=3.83
+ $Y=0.47 $X2=4.04 $Y2=0.69
r96 3 25 182 $w=1.7e-07 $l=2.98831e-07 $layer=licon1_NDIFF $count=1 $X=2.71
+ $Y=0.47 $X2=2.945 $Y2=0.615
r97 2 21 182 $w=1.7e-07 $l=3.57071e-07 $layer=licon1_NDIFF $count=1 $X=1.53
+ $Y=0.37 $X2=1.785 $Y2=0.615
r98 1 17 182 $w=1.7e-07 $l=2.36854e-07 $layer=licon1_NDIFF $count=1 $X=0.585
+ $Y=0.56 $X2=0.805 $Y2=0.595
.ends

