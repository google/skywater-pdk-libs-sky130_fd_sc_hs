# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_hs__nor3b_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__nor3b_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.800000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.558000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.485000 1.350000 4.675000 1.780000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.558000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.605000 1.350000 3.275000 1.780000 ;
    END
  END B
  PIN C_N
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425000 1.450000 0.835000 1.780000 ;
    END
  END C_N
  PIN Y
    ANTENNADIFFAREA  1.005700 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.120000 0.350000 1.395000 0.770000 ;
        RECT 1.120000 0.770000 2.695000 0.940000 ;
        RECT 1.565000 0.940000 2.695000 0.960000 ;
        RECT 1.565000 0.960000 4.185000 1.130000 ;
        RECT 1.640000 1.130000 1.810000 2.735000 ;
        RECT 2.505000 0.350000 2.695000 0.770000 ;
        RECT 3.925000 0.350000 4.185000 0.960000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 4.800000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 4.800000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.800000 0.085000 ;
      RECT 0.000000  3.245000 4.800000 3.415000 ;
      RECT 0.085000  0.350000 0.450000 1.110000 ;
      RECT 0.085000  1.110000 1.335000 1.280000 ;
      RECT 0.085000  1.280000 0.255000 1.950000 ;
      RECT 0.085000  1.950000 0.360000 2.980000 ;
      RECT 0.560000  1.950000 0.890000 3.245000 ;
      RECT 0.620000  0.085000 0.950000 0.940000 ;
      RECT 1.005000  1.280000 1.335000 1.550000 ;
      RECT 1.110000  1.820000 1.440000 2.905000 ;
      RECT 1.110000  2.905000 3.240000 3.075000 ;
      RECT 1.565000  0.085000 2.335000 0.600000 ;
      RECT 2.010000  1.820000 2.290000 2.905000 ;
      RECT 2.460000  1.950000 4.240000 2.120000 ;
      RECT 2.460000  2.120000 2.790000 2.735000 ;
      RECT 2.865000  0.085000 3.755000 0.770000 ;
      RECT 2.970000  2.290000 3.240000 2.905000 ;
      RECT 3.460000  2.290000 3.790000 3.245000 ;
      RECT 3.990000  2.120000 4.240000 2.980000 ;
      RECT 4.355000  0.085000 4.685000 1.130000 ;
      RECT 4.425000  1.950000 4.690000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
  END
END sky130_fd_sc_hs__nor3b_2
END LIBRARY
