# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_hs__sdfrtp_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  14.88000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.565000 0.810000 2.100000 1.265000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  1.086400 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 12.535000 0.350000 12.865000 0.930000 ;
        RECT 12.535000 0.930000 14.255000 1.100000 ;
        RECT 13.085000 1.770000 14.755000 1.940000 ;
        RECT 13.085000 1.940000 13.415000 2.980000 ;
        RECT 14.065000 1.940000 14.280000 2.980000 ;
        RECT 14.085000 0.350000 14.255000 0.930000 ;
        RECT 14.085000 1.100000 14.255000 1.300000 ;
        RECT 14.085000 1.300000 14.755000 1.770000 ;
    END
  END Q
  PIN RESET_B
    ANTENNAGATEAREA  0.411000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT  3.935000 1.920000  4.225000 1.965000 ;
        RECT  3.935000 1.965000 10.945000 2.105000 ;
        RECT  3.935000 2.105000  4.225000 2.150000 ;
        RECT  7.775000 1.920000  8.065000 1.965000 ;
        RECT  7.775000 2.105000  8.065000 2.150000 ;
        RECT 10.655000 1.920000 10.945000 1.965000 ;
        RECT 10.655000 2.105000 10.945000 2.150000 ;
    END
  END RESET_B
  PIN SCD
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.945000 1.440000 3.275000 2.150000 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605000 1.490000 2.735000 1.660000 ;
        RECT 0.605000 1.660000 1.795000 1.835000 ;
        RECT 2.405000 1.260000 2.735000 1.490000 ;
    END
  END SCE
  PIN CLK
    ANTENNAGATEAREA  0.261000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 3.840000 1.180000 4.195000 1.260000 ;
        RECT 3.840000 1.260000 4.635000 1.590000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 14.880000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 14.880000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 14.880000 0.085000 ;
      RECT  0.000000  3.245000 14.880000 3.415000 ;
      RECT  0.115000  0.350000  0.365000 0.935000 ;
      RECT  0.115000  0.935000  1.140000 1.265000 ;
      RECT  0.115000  1.265000  0.285000 2.005000 ;
      RECT  0.115000  2.005000  2.705000 2.175000 ;
      RECT  0.115000  2.175000  0.445000 2.980000 ;
      RECT  0.545000  0.085000  0.875000 0.765000 ;
      RECT  0.615000  2.345000  1.565000 3.245000 ;
      RECT  1.105000  0.255000  3.500000 0.425000 ;
      RECT  1.105000  0.425000  1.435000 0.640000 ;
      RECT  2.105000  2.345000  3.995000 2.420000 ;
      RECT  2.105000  2.420000  6.075000 2.515000 ;
      RECT  2.105000  2.515000  2.435000 2.980000 ;
      RECT  2.270000  0.595000  2.735000 0.845000 ;
      RECT  2.375000  1.830000  2.705000 2.005000 ;
      RECT  2.565000  0.845000  2.735000 0.920000 ;
      RECT  2.565000  0.920000  3.615000 1.090000 ;
      RECT  3.095000  2.685000  3.425000 3.245000 ;
      RECT  3.225000  0.425000  3.500000 0.750000 ;
      RECT  3.445000  1.090000  3.615000 2.330000 ;
      RECT  3.445000  2.330000  3.995000 2.345000 ;
      RECT  3.615000  2.515000  6.075000 2.580000 ;
      RECT  3.615000  2.580000  4.645000 2.590000 ;
      RECT  3.615000  2.590000  3.995000 2.980000 ;
      RECT  3.670000  0.085000  3.995000 0.750000 ;
      RECT  3.785000  1.830000  4.165000 2.160000 ;
      RECT  4.165000  0.550000  4.535000 0.750000 ;
      RECT  4.335000  1.820000  4.975000 1.990000 ;
      RECT  4.335000  1.990000  4.515000 2.250000 ;
      RECT  4.365000  0.750000  4.535000 0.920000 ;
      RECT  4.365000  0.920000  4.975000 1.090000 ;
      RECT  4.580000  2.410000  6.075000 2.420000 ;
      RECT  4.705000  2.750000  5.035000 3.245000 ;
      RECT  4.715000  0.085000  5.045000 0.750000 ;
      RECT  4.805000  1.090000  4.975000 1.410000 ;
      RECT  4.805000  1.410000  5.280000 1.740000 ;
      RECT  4.805000  1.740000  4.975000 1.820000 ;
      RECT  5.155000  1.910000  6.205000 1.915000 ;
      RECT  5.155000  1.915000  5.655000 2.240000 ;
      RECT  5.195000  0.920000  5.620000 1.240000 ;
      RECT  5.215000  0.330000  7.225000 0.500000 ;
      RECT  5.215000  0.500000  5.620000 0.920000 ;
      RECT  5.450000  1.240000  5.620000 1.585000 ;
      RECT  5.450000  1.585000  6.205000 1.910000 ;
      RECT  5.745000  2.580000  6.075000 2.755000 ;
      RECT  5.790000  0.670000  5.990000 1.245000 ;
      RECT  5.790000  1.245000  6.545000 1.415000 ;
      RECT  5.825000  2.085000  6.545000 2.255000 ;
      RECT  5.825000  2.255000  6.075000 2.410000 ;
      RECT  6.160000  0.670000  6.470000 0.905000 ;
      RECT  6.160000  0.905000  6.885000 1.075000 ;
      RECT  6.245000  2.425000  8.055000 2.490000 ;
      RECT  6.245000  2.490000  6.885000 2.755000 ;
      RECT  6.375000  1.415000  6.545000 2.085000 ;
      RECT  6.715000  1.075000  6.885000 2.320000 ;
      RECT  6.715000  2.320000  8.055000 2.425000 ;
      RECT  7.055000  0.500000  7.225000 0.580000 ;
      RECT  7.055000  0.580000  8.100000 0.750000 ;
      RECT  7.055000  0.920000  8.655000 1.090000 ;
      RECT  7.055000  1.090000  7.325000 1.945000 ;
      RECT  7.170000  2.660000  7.520000 3.245000 ;
      RECT  7.430000  0.085000  7.760000 0.410000 ;
      RECT  7.495000  1.260000  8.315000 1.575000 ;
      RECT  7.495000  1.575000  7.665000 2.320000 ;
      RECT  7.725000  2.490000  8.055000 2.755000 ;
      RECT  7.835000  1.820000  8.145000 2.150000 ;
      RECT  7.930000  0.255000  8.995000 0.425000 ;
      RECT  7.930000  0.425000  8.100000 0.580000 ;
      RECT  8.270000  0.595000  8.655000 0.920000 ;
      RECT  8.365000  1.745000  8.535000 3.245000 ;
      RECT  8.485000  1.090000  8.655000 1.405000 ;
      RECT  8.485000  1.405000  9.065000 1.575000 ;
      RECT  8.735000  1.575000  9.065000 2.755000 ;
      RECT  8.825000  0.425000  8.995000 0.905000 ;
      RECT  8.825000  0.905000  9.415000 1.235000 ;
      RECT  9.165000  0.405000  9.755000 0.735000 ;
      RECT  9.245000  1.235000  9.415000 2.065000 ;
      RECT  9.245000  2.065000  9.955000 2.380000 ;
      RECT  9.270000  2.550000 10.295000 2.880000 ;
      RECT  9.585000  0.735000  9.755000 0.885000 ;
      RECT  9.585000  0.885000 11.245000 1.055000 ;
      RECT  9.585000  1.055000  9.755000 1.725000 ;
      RECT  9.585000  1.725000 10.295000 1.895000 ;
      RECT 10.015000  1.225000 10.345000 1.385000 ;
      RECT 10.015000  1.385000 11.585000 1.555000 ;
      RECT 10.125000  1.895000 10.295000 2.550000 ;
      RECT 10.140000  0.085000 10.580000 0.680000 ;
      RECT 10.465000  2.520000 10.795000 3.245000 ;
      RECT 10.585000  1.820000 10.915000 2.150000 ;
      RECT 10.915000  1.055000 11.245000 1.215000 ;
      RECT 11.000000  2.520000 11.330000 2.980000 ;
      RECT 11.040000  0.385000 11.585000 0.715000 ;
      RECT 11.160000  1.555000 11.330000 2.520000 ;
      RECT 11.415000  0.715000 11.585000 1.385000 ;
      RECT 11.650000  1.820000 11.900000 3.245000 ;
      RECT 11.755000  0.350000 11.925000 1.270000 ;
      RECT 11.755000  1.270000 13.850000 1.600000 ;
      RECT 12.100000  1.600000 12.430000 2.700000 ;
      RECT 12.105000  0.085000 12.365000 1.100000 ;
      RECT 12.635000  1.820000 12.885000 3.245000 ;
      RECT 13.035000  0.085000 13.905000 0.760000 ;
      RECT 13.615000  2.110000 13.865000 3.245000 ;
      RECT 14.435000  0.085000 14.765000 1.130000 ;
      RECT 14.470000  2.110000 14.765000 3.245000 ;
    LAYER mcon ;
      RECT  0.155000 -0.085000  0.325000 0.085000 ;
      RECT  0.155000  3.245000  0.325000 3.415000 ;
      RECT  0.635000 -0.085000  0.805000 0.085000 ;
      RECT  0.635000  3.245000  0.805000 3.415000 ;
      RECT  1.115000 -0.085000  1.285000 0.085000 ;
      RECT  1.115000  3.245000  1.285000 3.415000 ;
      RECT  1.595000 -0.085000  1.765000 0.085000 ;
      RECT  1.595000  3.245000  1.765000 3.415000 ;
      RECT  2.075000 -0.085000  2.245000 0.085000 ;
      RECT  2.075000  3.245000  2.245000 3.415000 ;
      RECT  2.555000 -0.085000  2.725000 0.085000 ;
      RECT  2.555000  3.245000  2.725000 3.415000 ;
      RECT  3.035000 -0.085000  3.205000 0.085000 ;
      RECT  3.035000  3.245000  3.205000 3.415000 ;
      RECT  3.515000 -0.085000  3.685000 0.085000 ;
      RECT  3.515000  3.245000  3.685000 3.415000 ;
      RECT  3.995000 -0.085000  4.165000 0.085000 ;
      RECT  3.995000  1.950000  4.165000 2.120000 ;
      RECT  3.995000  3.245000  4.165000 3.415000 ;
      RECT  4.475000 -0.085000  4.645000 0.085000 ;
      RECT  4.475000  3.245000  4.645000 3.415000 ;
      RECT  4.955000 -0.085000  5.125000 0.085000 ;
      RECT  4.955000  3.245000  5.125000 3.415000 ;
      RECT  5.435000 -0.085000  5.605000 0.085000 ;
      RECT  5.435000  3.245000  5.605000 3.415000 ;
      RECT  5.915000 -0.085000  6.085000 0.085000 ;
      RECT  5.915000  3.245000  6.085000 3.415000 ;
      RECT  6.395000 -0.085000  6.565000 0.085000 ;
      RECT  6.395000  3.245000  6.565000 3.415000 ;
      RECT  6.875000 -0.085000  7.045000 0.085000 ;
      RECT  6.875000  3.245000  7.045000 3.415000 ;
      RECT  7.355000 -0.085000  7.525000 0.085000 ;
      RECT  7.355000  3.245000  7.525000 3.415000 ;
      RECT  7.835000 -0.085000  8.005000 0.085000 ;
      RECT  7.835000  1.950000  8.005000 2.120000 ;
      RECT  7.835000  3.245000  8.005000 3.415000 ;
      RECT  8.315000 -0.085000  8.485000 0.085000 ;
      RECT  8.315000  3.245000  8.485000 3.415000 ;
      RECT  8.795000 -0.085000  8.965000 0.085000 ;
      RECT  8.795000  3.245000  8.965000 3.415000 ;
      RECT  9.275000 -0.085000  9.445000 0.085000 ;
      RECT  9.275000  3.245000  9.445000 3.415000 ;
      RECT  9.755000 -0.085000  9.925000 0.085000 ;
      RECT  9.755000  3.245000  9.925000 3.415000 ;
      RECT 10.235000 -0.085000 10.405000 0.085000 ;
      RECT 10.235000  3.245000 10.405000 3.415000 ;
      RECT 10.715000 -0.085000 10.885000 0.085000 ;
      RECT 10.715000  1.950000 10.885000 2.120000 ;
      RECT 10.715000  3.245000 10.885000 3.415000 ;
      RECT 11.195000 -0.085000 11.365000 0.085000 ;
      RECT 11.195000  3.245000 11.365000 3.415000 ;
      RECT 11.675000 -0.085000 11.845000 0.085000 ;
      RECT 11.675000  3.245000 11.845000 3.415000 ;
      RECT 12.155000 -0.085000 12.325000 0.085000 ;
      RECT 12.155000  3.245000 12.325000 3.415000 ;
      RECT 12.635000 -0.085000 12.805000 0.085000 ;
      RECT 12.635000  3.245000 12.805000 3.415000 ;
      RECT 13.115000 -0.085000 13.285000 0.085000 ;
      RECT 13.115000  3.245000 13.285000 3.415000 ;
      RECT 13.595000 -0.085000 13.765000 0.085000 ;
      RECT 13.595000  3.245000 13.765000 3.415000 ;
      RECT 14.075000 -0.085000 14.245000 0.085000 ;
      RECT 14.075000  3.245000 14.245000 3.415000 ;
      RECT 14.555000 -0.085000 14.725000 0.085000 ;
      RECT 14.555000  3.245000 14.725000 3.415000 ;
  END
END sky130_fd_sc_hs__sdfrtp_4
