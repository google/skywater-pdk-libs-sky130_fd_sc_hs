# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_sc_hs__a31oi_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__a31oi_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.320000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.558000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.505000 1.430000 4.195000 1.780000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.558000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605000 1.430000 1.545000 1.780000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.558000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105000 1.090000 2.115000 1.260000 ;
        RECT 0.105000 1.260000 0.435000 1.550000 ;
        RECT 1.785000 1.260000 2.115000 1.550000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.447000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.325000 1.180000 2.995000 1.550000 ;
    END
  END B1
  PIN Y
    ANTENNADIFFAREA  1.090800 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.475000 1.720000 3.335000 1.890000 ;
        RECT 2.475000 1.890000 2.805000 2.735000 ;
        RECT 2.545000 0.255000 4.205000 0.425000 ;
        RECT 2.545000 0.425000 3.260000 0.580000 ;
        RECT 3.165000 1.090000 4.205000 1.260000 ;
        RECT 3.165000 1.260000 3.335000 1.720000 ;
        RECT 3.875000 0.425000 4.205000 1.090000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 4.320000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.000000 0.000000 4.320000 0.245000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.660000 4.510000 3.520000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 4.320000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.320000 0.085000 ;
      RECT 0.000000  3.245000 4.320000 3.415000 ;
      RECT 0.115000  0.085000 0.365000 0.920000 ;
      RECT 0.115000  1.820000 0.365000 1.950000 ;
      RECT 0.115000  1.950000 2.275000 2.120000 ;
      RECT 0.115000  2.120000 0.365000 2.980000 ;
      RECT 0.545000  0.255000 1.875000 0.425000 ;
      RECT 0.545000  0.425000 0.875000 0.920000 ;
      RECT 0.565000  2.290000 0.895000 3.245000 ;
      RECT 1.045000  0.595000 1.375000 0.750000 ;
      RECT 1.045000  0.750000 3.705000 0.920000 ;
      RECT 1.065000  2.120000 1.395000 2.980000 ;
      RECT 1.545000  0.425000 1.875000 0.580000 ;
      RECT 1.595000  2.290000 1.845000 3.245000 ;
      RECT 2.015000  2.120000 2.275000 2.905000 ;
      RECT 2.015000  2.905000 3.255000 3.075000 ;
      RECT 2.045000  0.085000 2.375000 0.580000 ;
      RECT 2.975000  2.060000 4.205000 2.230000 ;
      RECT 2.975000  2.230000 3.255000 2.905000 ;
      RECT 3.425000  2.400000 3.755000 3.245000 ;
      RECT 3.430000  0.670000 3.705000 0.750000 ;
      RECT 3.875000  1.950000 4.205000 2.060000 ;
      RECT 3.925000  2.230000 4.205000 2.980000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
  END
END sky130_fd_sc_hs__a31oi_2
END LIBRARY
