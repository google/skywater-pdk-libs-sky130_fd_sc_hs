* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hs__a2bb2o_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
X0 VPWR a_221_74# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X1 a_293_333# A2_N a_546_378# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=150000u
X2 a_149_74# B2 a_221_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X3 VPWR B2 a_61_392# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=150000u
X4 VGND A2_N a_293_333# VNB sky130_fd_pr__nfet_01v8_lvt w=550000u l=150000u
X5 a_61_392# a_293_333# a_221_74# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=150000u
X6 X a_221_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X7 a_293_333# A1_N VGND VNB sky130_fd_pr__nfet_01v8_lvt w=550000u l=150000u
X8 X a_221_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X9 VGND B1 a_149_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X10 VGND a_221_74# X VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X11 a_61_392# B1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=150000u
X12 a_546_378# A1_N VPWR VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=150000u
X13 a_221_74# a_293_333# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
.ends
