* File: sky130_fd_sc_hs__o221a_2.pex.spice
* Created: Tue Sep  1 20:15:32 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HS__O221A_2%C1 1 3 4 6 7 12
r28 12 13 30.8329 $w=3.83e-07 $l=2.45e-07 $layer=POLY_cond $X=0.505 $Y=1.492
+ $X2=0.75 $Y2=1.492
r29 10 12 29.5744 $w=3.83e-07 $l=2.35e-07 $layer=POLY_cond $X=0.27 $Y=1.492
+ $X2=0.505 $Y2=1.492
r30 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.27
+ $Y=1.385 $X2=0.27 $Y2=1.385
r31 7 11 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=0.27 $Y=1.295 $X2=0.27
+ $Y2=1.385
r32 4 13 24.8035 $w=1.5e-07 $l=2.72e-07 $layer=POLY_cond $X=0.75 $Y=1.22
+ $X2=0.75 $Y2=1.492
r33 4 6 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=0.75 $Y=1.22 $X2=0.75
+ $Y2=0.74
r34 1 12 24.8035 $w=1.5e-07 $l=2.73e-07 $layer=POLY_cond $X=0.505 $Y=1.765
+ $X2=0.505 $Y2=1.492
r35 1 3 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=0.505 $Y=1.765
+ $X2=0.505 $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_HS__O221A_2%B1 3 5 7 8 12 13
c39 3 0 5.3557e-20 $X=1.245 $Y=0.74
r40 11 13 2.55477 $w=2.83e-07 $l=1.5e-08 $layer=POLY_cond $X=1.23 $Y=1.557
+ $X2=1.245 $Y2=1.557
r41 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.23
+ $Y=1.515 $X2=1.23 $Y2=1.515
r42 8 12 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=1.23 $Y=1.665
+ $X2=1.23 $Y2=1.515
r43 5 13 57.9081 $w=2.83e-07 $l=4.31648e-07 $layer=POLY_cond $X=1.585 $Y=1.765
+ $X2=1.245 $Y2=1.557
r44 5 7 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=1.585 $Y=1.765
+ $X2=1.585 $Y2=2.34
r45 1 13 17.601 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.245 $Y=1.35
+ $X2=1.245 $Y2=1.557
r46 1 3 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.245 $Y=1.35
+ $X2=1.245 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HS__O221A_2%B2 1 3 4 5 6 8 13 14
c39 6 0 1.20527e-19 $X=2.005 $Y=1.765
c40 1 0 1.67816e-19 $X=1.75 $Y=1.185
r41 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.08
+ $Y=1.515 $X2=2.08 $Y2=1.515
r42 14 19 2.14408 $w=4.28e-07 $l=8e-08 $layer=LI1_cond $X=2.16 $Y=1.565 $X2=2.08
+ $Y2=1.565
r43 13 19 10.7204 $w=4.28e-07 $l=4e-07 $layer=LI1_cond $X=1.68 $Y=1.565 $X2=2.08
+ $Y2=1.565
r44 6 18 53.429 $w=2.79e-07 $l=2.85044e-07 $layer=POLY_cond $X=2.005 $Y=1.765
+ $X2=2.08 $Y2=1.515
r45 6 8 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=2.005 $Y=1.765
+ $X2=2.005 $Y2=2.34
r46 5 18 1.29086 $w=3.3e-07 $l=8.75758e-08 $layer=POLY_cond $X=2.08 $Y=1.515
+ $X2=2.08 $Y2=1.515
r47 4 9 169.213 $w=1.5e-07 $l=3.3e-07 $layer=POLY_cond $X=2.08 $Y=1.26 $X2=1.75
+ $Y2=1.26
r48 4 5 31.475 $w=3.3e-07 $l=1.8e-07 $layer=POLY_cond $X=2.08 $Y=1.335 $X2=2.08
+ $Y2=1.515
r49 1 9 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.75 $Y=1.185 $X2=1.75
+ $Y2=1.26
r50 1 3 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=1.75 $Y=1.185
+ $X2=1.75 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HS__O221A_2%A2 1 3 6 8 12
c29 12 0 1.20527e-19 $X=2.65 $Y=1.515
r30 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.65
+ $Y=1.515 $X2=2.65 $Y2=1.515
r31 8 12 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=2.65 $Y=1.665
+ $X2=2.65 $Y2=1.515
r32 4 11 38.5562 $w=2.99e-07 $l=2.05122e-07 $layer=POLY_cond $X=2.74 $Y=1.35
+ $X2=2.65 $Y2=1.515
r33 4 6 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.74 $Y=1.35 $X2=2.74
+ $Y2=0.74
r34 1 11 52.2586 $w=2.99e-07 $l=2.85044e-07 $layer=POLY_cond $X=2.575 $Y=1.765
+ $X2=2.65 $Y2=1.515
r35 1 3 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=2.575 $Y=1.765
+ $X2=2.575 $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_HS__O221A_2%A1 1 3 6 8 12
c35 1 0 1.17931e-19 $X=3.145 $Y=1.765
r36 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.22
+ $Y=1.515 $X2=3.22 $Y2=1.515
r37 8 12 4.54912 $w=3.78e-07 $l=1.5e-07 $layer=LI1_cond $X=3.195 $Y=1.665
+ $X2=3.195 $Y2=1.515
r38 4 11 38.5562 $w=2.99e-07 $l=1.88348e-07 $layer=POLY_cond $X=3.17 $Y=1.35
+ $X2=3.22 $Y2=1.515
r39 4 6 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=3.17 $Y=1.35 $X2=3.17
+ $Y2=0.74
r40 1 11 52.2586 $w=2.99e-07 $l=2.85044e-07 $layer=POLY_cond $X=3.145 $Y=1.765
+ $X2=3.22 $Y2=1.515
r41 1 3 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=3.145 $Y=1.765
+ $X2=3.145 $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_HS__O221A_2%A_27_368# 1 2 3 12 14 16 17 21 24 25 27 28
+ 31 35 38 39 43 45 48 53 54 56 60
r112 61 63 14.557 $w=2.98e-07 $l=9e-08 $layer=POLY_cond $X=3.765 $Y=1.485
+ $X2=3.765 $Y2=1.395
r113 60 61 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.76
+ $Y=1.485 $X2=3.76 $Y2=1.485
r114 57 60 3.84148 $w=3.28e-07 $l=1.1e-07 $layer=LI1_cond $X=3.65 $Y=1.485
+ $X2=3.76 $Y2=1.485
r115 52 53 5.41145 $w=2.98e-07 $l=8.5e-08 $layer=LI1_cond $X=0.69 $Y=1.97
+ $X2=0.775 $Y2=1.97
r116 50 52 15.7501 $w=2.98e-07 $l=4.1e-07 $layer=LI1_cond $X=0.28 $Y=1.97
+ $X2=0.69 $Y2=1.97
r117 47 57 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.65 $Y=1.65
+ $X2=3.65 $Y2=1.485
r118 47 48 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=3.65 $Y=1.65 $X2=3.65
+ $Y2=1.95
r119 46 56 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.395 $Y=2.035
+ $X2=2.23 $Y2=2.035
r120 45 48 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.565 $Y=2.035
+ $X2=3.65 $Y2=1.95
r121 45 46 76.3316 $w=1.68e-07 $l=1.17e-06 $layer=LI1_cond $X=3.565 $Y=2.035
+ $X2=2.395 $Y2=2.035
r122 41 56 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.23 $Y=2.12
+ $X2=2.23 $Y2=2.035
r123 41 43 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=2.23 $Y=2.12
+ $X2=2.23 $Y2=2.375
r124 39 56 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.065 $Y=2.035
+ $X2=2.23 $Y2=2.035
r125 39 53 84.1604 $w=1.68e-07 $l=1.29e-06 $layer=LI1_cond $X=2.065 $Y=2.035
+ $X2=0.775 $Y2=2.035
r126 38 52 4.061 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=0.69 $Y=1.82 $X2=0.69
+ $Y2=1.97
r127 38 54 52.8449 $w=1.68e-07 $l=8.1e-07 $layer=LI1_cond $X=0.69 $Y=1.82
+ $X2=0.69 $Y2=1.01
r128 33 54 9.72165 $w=4.03e-07 $l=2.02e-07 $layer=LI1_cond $X=0.572 $Y=0.808
+ $X2=0.572 $Y2=1.01
r129 33 35 8.33743 $w=4.03e-07 $l=2.93e-07 $layer=LI1_cond $X=0.572 $Y=0.808
+ $X2=0.572 $Y2=0.515
r130 29 50 0.126616 $w=3.3e-07 $l=1.5e-07 $layer=LI1_cond $X=0.28 $Y=2.12
+ $X2=0.28 $Y2=1.97
r131 29 31 20.0804 $w=3.28e-07 $l=5.75e-07 $layer=LI1_cond $X=0.28 $Y=2.12
+ $X2=0.28 $Y2=2.695
r132 25 27 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=4.295 $Y=1.765
+ $X2=4.295 $Y2=2.4
r133 24 25 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=4.295 $Y=1.675
+ $X2=4.295 $Y2=1.765
r134 23 28 18.8402 $w=1.65e-07 $l=9.87421e-08 $layer=POLY_cond $X=4.295 $Y=1.47
+ $X2=4.24 $Y2=1.395
r135 23 24 79.6855 $w=1.8e-07 $l=2.05e-07 $layer=POLY_cond $X=4.295 $Y=1.47
+ $X2=4.295 $Y2=1.675
r136 19 28 18.8402 $w=1.65e-07 $l=1.04283e-07 $layer=POLY_cond $X=4.17 $Y=1.32
+ $X2=4.24 $Y2=1.395
r137 19 21 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=4.17 $Y=1.32
+ $X2=4.17 $Y2=0.74
r138 18 63 18.8112 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=3.935 $Y=1.395
+ $X2=3.765 $Y2=1.395
r139 17 28 6.66866 $w=1.5e-07 $l=1.45e-07 $layer=POLY_cond $X=4.095 $Y=1.395
+ $X2=4.24 $Y2=1.395
r140 17 18 82.0426 $w=1.5e-07 $l=1.6e-07 $layer=POLY_cond $X=4.095 $Y=1.395
+ $X2=3.935 $Y2=1.395
r141 14 61 57.1617 $w=2.98e-07 $l=3.1749e-07 $layer=POLY_cond $X=3.845 $Y=1.765
+ $X2=3.765 $Y2=1.485
r142 14 16 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.845 $Y=1.765
+ $X2=3.845 $Y2=2.4
r143 10 63 24.0039 $w=2.98e-07 $l=8.66025e-08 $layer=POLY_cond $X=3.74 $Y=1.32
+ $X2=3.765 $Y2=1.395
r144 10 12 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=3.74 $Y=1.32
+ $X2=3.74 $Y2=0.74
r145 3 56 600 $w=1.7e-07 $l=2.59374e-07 $layer=licon1_PDIFF $count=1 $X=2.08
+ $Y=1.84 $X2=2.23 $Y2=2.035
r146 3 43 300 $w=1.7e-07 $l=6.05372e-07 $layer=licon1_PDIFF $count=2 $X=2.08
+ $Y=1.84 $X2=2.23 $Y2=2.375
r147 2 50 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=1.985
r148 2 31 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.695
r149 1 35 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.39
+ $Y=0.37 $X2=0.535 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__O221A_2%VPWR 1 2 3 12 16 20 22 26 28 33 41 47 50 54
r47 53 54 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r48 50 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r49 47 48 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r50 45 54 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=4.56 $Y2=3.33
r51 45 51 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=3.6 $Y2=3.33
r52 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r53 42 50 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.735 $Y=3.33
+ $X2=3.57 $Y2=3.33
r54 42 44 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=3.735 $Y=3.33
+ $X2=4.08 $Y2=3.33
r55 41 53 4.01252 $w=1.7e-07 $l=1.82e-07 $layer=LI1_cond $X=4.435 $Y=3.33
+ $X2=4.617 $Y2=3.33
r56 41 44 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=4.435 $Y=3.33
+ $X2=4.08 $Y2=3.33
r57 40 51 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=3.6 $Y2=3.33
r58 39 40 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r59 37 48 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r60 36 39 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.68 $Y=3.33
+ $X2=3.12 $Y2=3.33
r61 36 37 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r62 34 47 15.5867 $w=1.7e-07 $l=4.55e-07 $layer=LI1_cond $X=1.525 $Y=3.33
+ $X2=1.07 $Y2=3.33
r63 34 36 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=1.525 $Y=3.33
+ $X2=1.68 $Y2=3.33
r64 33 50 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.405 $Y=3.33
+ $X2=3.57 $Y2=3.33
r65 33 39 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=3.405 $Y=3.33
+ $X2=3.12 $Y2=3.33
r66 31 48 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=1.2 $Y2=3.33
r67 30 31 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r68 28 47 15.5867 $w=1.7e-07 $l=4.55e-07 $layer=LI1_cond $X=0.615 $Y=3.33
+ $X2=1.07 $Y2=3.33
r69 28 30 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=0.615 $Y=3.33
+ $X2=0.24 $Y2=3.33
r70 26 40 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=2.4 $Y=3.33
+ $X2=3.12 $Y2=3.33
r71 26 37 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=2.4 $Y=3.33
+ $X2=1.68 $Y2=3.33
r72 22 25 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=4.56 $Y=1.985
+ $X2=4.56 $Y2=2.815
r73 20 53 3.13065 $w=2.5e-07 $l=1.09864e-07 $layer=LI1_cond $X=4.56 $Y=3.245
+ $X2=4.617 $Y2=3.33
r74 20 25 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=4.56 $Y=3.245
+ $X2=4.56 $Y2=2.815
r75 16 19 12.5721 $w=3.28e-07 $l=3.6e-07 $layer=LI1_cond $X=3.57 $Y=2.455
+ $X2=3.57 $Y2=2.815
r76 14 50 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.57 $Y=3.245
+ $X2=3.57 $Y2=3.33
r77 14 19 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=3.57 $Y=3.245
+ $X2=3.57 $Y2=2.815
r78 10 47 3.36946 $w=9.1e-07 $l=8.5e-08 $layer=LI1_cond $X=1.07 $Y=3.245
+ $X2=1.07 $Y2=3.33
r79 10 12 11.6637 $w=9.08e-07 $l=8.7e-07 $layer=LI1_cond $X=1.07 $Y=3.245
+ $X2=1.07 $Y2=2.375
r80 3 25 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=4.37
+ $Y=1.84 $X2=4.52 $Y2=2.815
r81 3 22 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=4.37
+ $Y=1.84 $X2=4.52 $Y2=1.985
r82 2 19 600 $w=1.7e-07 $l=1.13661e-06 $layer=licon1_PDIFF $count=1 $X=3.22
+ $Y=1.84 $X2=3.57 $Y2=2.815
r83 2 16 600 $w=1.7e-07 $l=7.70373e-07 $layer=licon1_PDIFF $count=1 $X=3.22
+ $Y=1.84 $X2=3.57 $Y2=2.455
r84 1 12 150 $w=1.7e-07 $l=1.01277e-06 $layer=licon1_PDIFF $count=4 $X=0.58
+ $Y=1.84 $X2=1.36 $Y2=2.375
.ends

.subckt PM_SKY130_FD_SC_HS__O221A_2%X 1 2 9 14 15 16 17 23 29
c36 14 0 1.17931e-19 $X=4.07 $Y=1.985
r37 21 29 0.805779 $w=4.73e-07 $l=3.2e-08 $layer=LI1_cond $X=4.027 $Y=0.893
+ $X2=4.027 $Y2=0.925
r38 17 31 9.71933 $w=4.73e-07 $l=1.79e-07 $layer=LI1_cond $X=4.027 $Y=0.951
+ $X2=4.027 $Y2=1.13
r39 17 29 0.654696 $w=4.73e-07 $l=2.6e-08 $layer=LI1_cond $X=4.027 $Y=0.951
+ $X2=4.027 $Y2=0.925
r40 17 21 0.679876 $w=4.73e-07 $l=2.7e-08 $layer=LI1_cond $X=4.027 $Y=0.866
+ $X2=4.027 $Y2=0.893
r41 16 17 7.83117 $w=4.73e-07 $l=3.11e-07 $layer=LI1_cond $X=4.027 $Y=0.555
+ $X2=4.027 $Y2=0.866
r42 16 23 1.00722 $w=4.73e-07 $l=4e-08 $layer=LI1_cond $X=4.027 $Y=0.555
+ $X2=4.027 $Y2=0.515
r43 15 31 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=4.18 $Y=1.82 $X2=4.18
+ $Y2=1.13
r44 14 15 8.51103 $w=3.58e-07 $l=1.65e-07 $layer=LI1_cond $X=4.085 $Y=1.985
+ $X2=4.085 $Y2=1.82
r45 7 14 0.480185 $w=3.58e-07 $l=1.5e-08 $layer=LI1_cond $X=4.085 $Y=2 $X2=4.085
+ $Y2=1.985
r46 7 9 26.09 $w=3.58e-07 $l=8.15e-07 $layer=LI1_cond $X=4.085 $Y=2 $X2=4.085
+ $Y2=2.815
r47 2 14 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=3.92
+ $Y=1.84 $X2=4.07 $Y2=1.985
r48 2 9 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=3.92
+ $Y=1.84 $X2=4.07 $Y2=2.815
r49 1 23 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.815
+ $Y=0.37 $X2=3.955 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__O221A_2%A_165_74# 1 2 9 12 13
r26 13 16 8.03218 $w=3.28e-07 $l=2.3e-07 $layer=LI1_cond $X=1.965 $Y=0.435
+ $X2=1.965 $Y2=0.665
r27 10 12 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.115 $Y=0.435
+ $X2=1.03 $Y2=0.435
r28 9 13 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.8 $Y=0.435
+ $X2=1.965 $Y2=0.435
r29 9 10 44.6898 $w=1.68e-07 $l=6.85e-07 $layer=LI1_cond $X=1.8 $Y=0.435
+ $X2=1.115 $Y2=0.435
r30 2 16 182 $w=1.7e-07 $l=3.58225e-07 $layer=licon1_NDIFF $count=1 $X=1.825
+ $Y=0.37 $X2=1.965 $Y2=0.665
r31 1 12 91 $w=1.7e-07 $l=2.67862e-07 $layer=licon1_NDIFF $count=2 $X=0.825
+ $Y=0.37 $X2=1.03 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__O221A_2%A_264_74# 1 2 7 11 14
c35 14 0 1.67816e-19 $X=1.495 $Y=0.965
c36 7 0 5.3557e-20 $X=2.87 $Y=1.095
r37 14 16 4.60977 $w=3.23e-07 $l=1.3e-07 $layer=LI1_cond $X=1.457 $Y=0.965
+ $X2=1.457 $Y2=1.095
r38 9 11 22.8184 $w=2.48e-07 $l=4.95e-07 $layer=LI1_cond $X=2.995 $Y=1.01
+ $X2=2.995 $Y2=0.515
r39 8 16 4.53325 $w=1.7e-07 $l=1.63e-07 $layer=LI1_cond $X=1.62 $Y=1.095
+ $X2=1.457 $Y2=1.095
r40 7 9 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=2.87 $Y=1.095
+ $X2=2.995 $Y2=1.01
r41 7 8 81.5508 $w=1.68e-07 $l=1.25e-06 $layer=LI1_cond $X=2.87 $Y=1.095
+ $X2=1.62 $Y2=1.095
r42 2 11 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.815
+ $Y=0.37 $X2=2.955 $Y2=0.515
r43 1 14 182 $w=1.7e-07 $l=6.76868e-07 $layer=licon1_NDIFF $count=1 $X=1.32
+ $Y=0.37 $X2=1.495 $Y2=0.965
.ends

.subckt PM_SKY130_FD_SC_HS__O221A_2%VGND 1 2 3 12 16 18 20 23 24 26 27 28 40 46
r54 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r55 43 46 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=4.56
+ $Y2=0
r56 42 43 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r57 40 45 4.01252 $w=1.7e-07 $l=1.82e-07 $layer=LI1_cond $X=4.435 $Y=0 $X2=4.617
+ $Y2=0
r58 40 42 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=4.435 $Y=0 $X2=4.08
+ $Y2=0
r59 39 43 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=4.08
+ $Y2=0
r60 38 39 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r61 35 36 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r62 32 36 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=0.24 $Y=0 $X2=2.16
+ $Y2=0
r63 31 35 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=0.24 $Y=0 $X2=2.16
+ $Y2=0
r64 31 32 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r65 28 39 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=2.4 $Y=0 $X2=3.12
+ $Y2=0
r66 28 36 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.4 $Y=0 $X2=2.16
+ $Y2=0
r67 26 38 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=3.29 $Y=0 $X2=3.12
+ $Y2=0
r68 26 27 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.29 $Y=0 $X2=3.455
+ $Y2=0
r69 25 42 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=3.62 $Y=0 $X2=4.08
+ $Y2=0
r70 25 27 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.62 $Y=0 $X2=3.455
+ $Y2=0
r71 23 35 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=2.36 $Y=0 $X2=2.16
+ $Y2=0
r72 23 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.36 $Y=0 $X2=2.525
+ $Y2=0
r73 22 38 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=2.69 $Y=0 $X2=3.12
+ $Y2=0
r74 22 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.69 $Y=0 $X2=2.525
+ $Y2=0
r75 18 45 3.13065 $w=2.5e-07 $l=1.09864e-07 $layer=LI1_cond $X=4.56 $Y=0.085
+ $X2=4.617 $Y2=0
r76 18 20 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=4.56 $Y=0.085
+ $X2=4.56 $Y2=0.515
r77 14 27 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.455 $Y=0.085
+ $X2=3.455 $Y2=0
r78 14 16 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=3.455 $Y=0.085
+ $X2=3.455 $Y2=0.515
r79 10 24 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.525 $Y=0.085
+ $X2=2.525 $Y2=0
r80 10 12 20.2551 $w=3.28e-07 $l=5.8e-07 $layer=LI1_cond $X=2.525 $Y=0.085
+ $X2=2.525 $Y2=0.665
r81 3 20 91 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_NDIFF $count=2 $X=4.245
+ $Y=0.37 $X2=4.52 $Y2=0.515
r82 2 16 91 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=2 $X=3.245
+ $Y=0.37 $X2=3.455 $Y2=0.515
r83 1 12 182 $w=1.7e-07 $l=3.60278e-07 $layer=licon1_NDIFF $count=1 $X=2.38
+ $Y=0.37 $X2=2.525 $Y2=0.665
.ends

