* NGSPICE file created from sky130_fd_sc_hs__a311oi_1.ext - technology: sky130A

.subckt sky130_fd_sc_hs__a311oi_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
M1000 a_156_368# A3 VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=6.72e+11p pd=5.68e+06u as=8.456e+11p ps=5.99e+06u
M1001 VPWR A2 a_156_368# VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1002 a_231_74# A2 a_159_74# VNB nlowvt w=740000u l=150000u
+  ad=2.886e+11p pd=2.26e+06u as=1.554e+11p ps=1.9e+06u
M1003 Y C1 VGND VNB nlowvt w=740000u l=150000u
+  ad=4.847e+11p pd=4.27e+06u as=4.847e+11p ps=4.27e+06u
M1004 a_159_74# A3 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 Y C1 a_462_368# VPB pshort w=1.12e+06u l=150000u
+  ad=3.08e+11p pd=2.79e+06u as=3.696e+11p ps=2.9e+06u
M1006 Y A1 a_231_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_156_368# A1 VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_462_368# B1 a_156_368# VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VGND B1 Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

