* File: sky130_fd_sc_hs__dlrtn_2.pex.spice
* Created: Thu Aug 27 20:41:32 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HS__DLRTN_2%D 3 5 7 8
r27 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.6
+ $Y=1.615 $X2=0.6 $Y2=1.615
r28 8 12 4.1907 $w=3.28e-07 $l=1.2e-07 $layer=LI1_cond $X=0.72 $Y=1.615 $X2=0.6
+ $Y2=1.615
r29 5 11 56.8989 $w=3.02e-07 $l=3.1881e-07 $layer=POLY_cond $X=0.675 $Y=1.895
+ $X2=0.592 $Y2=1.615
r30 5 7 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=0.675 $Y=1.895
+ $X2=0.675 $Y2=2.39
r31 1 11 38.5446 $w=3.02e-07 $l=2.07918e-07 $layer=POLY_cond $X=0.495 $Y=1.45
+ $X2=0.592 $Y2=1.615
r32 1 3 253.819 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=0.495 $Y=1.45
+ $X2=0.495 $Y2=0.955
.ends

.subckt PM_SKY130_FD_SC_HS__DLRTN_2%GATE_N 3 5 7 8
r35 8 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.17
+ $Y=1.615 $X2=1.17 $Y2=1.615
r36 5 11 57.6553 $w=2.91e-07 $l=3.06268e-07 $layer=POLY_cond $X=1.225 $Y=1.895
+ $X2=1.17 $Y2=1.615
r37 5 7 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=1.225 $Y=1.895
+ $X2=1.225 $Y2=2.39
r38 1 11 38.6072 $w=2.91e-07 $l=2.03101e-07 $layer=POLY_cond $X=1.085 $Y=1.45
+ $X2=1.17 $Y2=1.615
r39 1 3 302.532 $w=1.5e-07 $l=5.9e-07 $layer=POLY_cond $X=1.085 $Y=1.45
+ $X2=1.085 $Y2=0.86
.ends

.subckt PM_SKY130_FD_SC_HS__DLRTN_2%A_232_98# 1 2 7 10 11 13 16 20 22 24 25 26
+ 31 32 34 35 38 42 43 48 53
r120 52 53 2.03662 $w=3.55e-07 $l=1.5e-08 $layer=POLY_cond $X=3.8 $Y=2.237
+ $X2=3.815 $Y2=2.237
r121 47 48 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=1.74 $Y=1.505
+ $X2=1.74 $Y2=1.415
r122 46 47 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.74
+ $Y=1.505 $X2=1.74 $Y2=1.505
r123 42 43 8.60763 $w=3.88e-07 $l=1.65e-07 $layer=LI1_cond $X=1.48 $Y=2.115
+ $X2=1.48 $Y2=1.95
r124 39 53 46.8423 $w=3.55e-07 $l=3.45e-07 $layer=POLY_cond $X=4.16 $Y=2.237
+ $X2=3.815 $Y2=2.237
r125 38 39 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.16
+ $Y=2.195 $X2=4.16 $Y2=2.195
r126 36 38 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=4.16 $Y=2.52
+ $X2=4.16 $Y2=2.195
r127 34 36 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.995 $Y=2.605
+ $X2=4.16 $Y2=2.52
r128 34 35 151.358 $w=1.68e-07 $l=2.32e-06 $layer=LI1_cond $X=3.995 $Y=2.605
+ $X2=1.675 $Y2=2.605
r129 32 46 9.11389 $w=2.71e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.59 $Y=1.67
+ $X2=1.675 $Y2=1.505
r130 32 43 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=1.59 $Y=1.67
+ $X2=1.59 $Y2=1.95
r131 31 35 8.28377 $w=1.7e-07 $l=2.33666e-07 $layer=LI1_cond $X=1.48 $Y=2.52
+ $X2=1.675 $Y2=2.605
r132 30 42 0.886495 $w=3.88e-07 $l=3e-08 $layer=LI1_cond $X=1.48 $Y=2.145
+ $X2=1.48 $Y2=2.115
r133 30 31 11.0812 $w=3.88e-07 $l=3.75e-07 $layer=LI1_cond $X=1.48 $Y=2.145
+ $X2=1.48 $Y2=2.52
r134 26 46 18.9077 $w=2.71e-07 $l=4.2e-07 $layer=LI1_cond $X=1.675 $Y=1.085
+ $X2=1.675 $Y2=1.505
r135 26 28 7.15912 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=1.505 $Y=1.085
+ $X2=1.3 $Y2=1.085
r136 22 53 22.9692 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=3.815 $Y=2.445
+ $X2=3.815 $Y2=2.237
r137 22 24 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=3.815 $Y=2.445
+ $X2=3.815 $Y2=2.73
r138 18 52 22.9692 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.8 $Y=2.03
+ $X2=3.8 $Y2=2.237
r139 18 20 687.106 $w=1.5e-07 $l=1.34e-06 $layer=POLY_cond $X=3.8 $Y=2.03
+ $X2=3.8 $Y2=0.69
r140 14 25 18.8402 $w=1.65e-07 $l=8.21584e-08 $layer=POLY_cond $X=2.25 $Y=1.34
+ $X2=2.235 $Y2=1.415
r141 14 16 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=2.25 $Y=1.34
+ $X2=2.25 $Y2=0.78
r142 11 13 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=2.235 $Y=1.885
+ $X2=2.235 $Y2=2.38
r143 10 11 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=2.235 $Y=1.795
+ $X2=2.235 $Y2=1.885
r144 9 25 18.8402 $w=1.65e-07 $l=7.5e-08 $layer=POLY_cond $X=2.235 $Y=1.49
+ $X2=2.235 $Y2=1.415
r145 9 10 118.556 $w=1.8e-07 $l=3.05e-07 $layer=POLY_cond $X=2.235 $Y=1.49
+ $X2=2.235 $Y2=1.795
r146 8 48 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.905 $Y=1.415
+ $X2=1.74 $Y2=1.415
r147 7 25 6.66866 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=2.145 $Y=1.415
+ $X2=2.235 $Y2=1.415
r148 7 8 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=2.145 $Y=1.415
+ $X2=1.905 $Y2=1.415
r149 2 42 300 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=2 $X=1.3
+ $Y=1.97 $X2=1.45 $Y2=2.115
r150 1 28 182 $w=1.7e-07 $l=6.16036e-07 $layer=licon1_NDIFF $count=1 $X=1.16
+ $Y=0.49 $X2=1.3 $Y2=1.04
.ends

.subckt PM_SKY130_FD_SC_HS__DLRTN_2%A_27_136# 1 2 7 8 9 11 12 14 16 20 25 26 29
+ 32 34 35
c78 7 0 5.22992e-20 $X=2.855 $Y=1.59
r79 34 35 9.6413 $w=5.18e-07 $l=1.65e-07 $layer=LI1_cond $X=0.355 $Y=2.115
+ $X2=0.355 $Y2=1.95
r80 32 35 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=0.18 $Y=1.25 $X2=0.18
+ $Y2=1.95
r81 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.78
+ $Y=1.425 $X2=2.78 $Y2=1.425
r82 27 29 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=2.78 $Y=0.75
+ $X2=2.78 $Y2=1.425
r83 25 27 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.615 $Y=0.665
+ $X2=2.78 $Y2=0.75
r84 25 26 141.572 $w=1.68e-07 $l=2.17e-06 $layer=LI1_cond $X=2.615 $Y=0.665
+ $X2=0.445 $Y2=0.665
r85 18 32 8.81775 $w=3.48e-07 $l=1.75e-07 $layer=LI1_cond $X=0.27 $Y=1.075
+ $X2=0.27 $Y2=1.25
r86 18 20 3.95123 $w=3.48e-07 $l=1.2e-07 $layer=LI1_cond $X=0.27 $Y=1.075
+ $X2=0.27 $Y2=0.955
r87 17 26 7.93686 $w=1.7e-07 $l=2.13307e-07 $layer=LI1_cond $X=0.27 $Y=0.75
+ $X2=0.445 $Y2=0.665
r88 17 20 6.75002 $w=3.48e-07 $l=2.05e-07 $layer=LI1_cond $X=0.27 $Y=0.75
+ $X2=0.27 $Y2=0.955
r89 14 16 134.96 $w=1.5e-07 $l=4.2e-07 $layer=POLY_cond $X=3.41 $Y=1.11 $X2=3.41
+ $Y2=0.69
r90 13 30 42.3736 $w=2.73e-07 $l=3.11769e-07 $layer=POLY_cond $X=2.945 $Y=1.185
+ $X2=2.78 $Y2=1.425
r91 12 14 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.335 $Y=1.185
+ $X2=3.41 $Y2=1.11
r92 12 13 199.979 $w=1.5e-07 $l=3.9e-07 $layer=POLY_cond $X=3.335 $Y=1.185
+ $X2=2.945 $Y2=1.185
r93 9 11 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=2.855 $Y=1.885
+ $X2=2.855 $Y2=2.46
r94 8 9 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=2.855 $Y=1.795 $X2=2.855
+ $Y2=1.885
r95 7 30 34.7287 $w=2.73e-07 $l=1.98997e-07 $layer=POLY_cond $X=2.855 $Y=1.59
+ $X2=2.78 $Y2=1.425
r96 7 8 79.6855 $w=1.8e-07 $l=2.05e-07 $layer=POLY_cond $X=2.855 $Y=1.59
+ $X2=2.855 $Y2=1.795
r97 2 34 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=0.305
+ $Y=1.97 $X2=0.45 $Y2=2.115
r98 1 20 182 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.68 $X2=0.28 $Y2=0.955
.ends

.subckt PM_SKY130_FD_SC_HS__DLRTN_2%A_373_82# 1 2 7 9 12 16 21 23 25 26 31 33 34
c94 31 0 5.22992e-20 $X=2.16 $Y=1.045
r95 33 36 6.33844 $w=3.98e-07 $l=2.2e-07 $layer=LI1_cond $X=2.045 $Y=1.925
+ $X2=2.045 $Y2=2.145
r96 33 34 6.34273 $w=3.98e-07 $l=8.5e-08 $layer=LI1_cond $X=2.045 $Y=1.925
+ $X2=2.045 $Y2=1.84
r97 29 31 6.45368 $w=2.48e-07 $l=1.4e-07 $layer=LI1_cond $X=2.02 $Y=1.045
+ $X2=2.16 $Y2=1.045
r98 26 40 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.25 $Y=1.355
+ $X2=4.25 $Y2=1.19
r99 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.25
+ $Y=1.355 $X2=4.25 $Y2=1.355
r100 23 25 26.7157 $w=3.28e-07 $l=7.65e-07 $layer=LI1_cond $X=3.485 $Y=1.355
+ $X2=4.25 $Y2=1.355
r101 21 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.32
+ $Y=1.635 $X2=3.32 $Y2=1.635
r102 19 21 7.15912 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=3.32 $Y=1.84
+ $X2=3.32 $Y2=1.635
r103 18 23 6.81649 $w=3.3e-07 $l=2.33345e-07 $layer=LI1_cond $X=3.32 $Y=1.52
+ $X2=3.485 $Y2=1.355
r104 18 21 4.01609 $w=3.28e-07 $l=1.15e-07 $layer=LI1_cond $X=3.32 $Y=1.52
+ $X2=3.32 $Y2=1.635
r105 17 33 5.77842 $w=1.7e-07 $l=2e-07 $layer=LI1_cond $X=2.245 $Y=1.925
+ $X2=2.045 $Y2=1.925
r106 16 19 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.155 $Y=1.925
+ $X2=3.32 $Y2=1.84
r107 16 17 59.369 $w=1.68e-07 $l=9.1e-07 $layer=LI1_cond $X=3.155 $Y=1.925
+ $X2=2.245 $Y2=1.925
r108 14 31 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.16 $Y=1.17
+ $X2=2.16 $Y2=1.045
r109 14 34 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.16 $Y=1.17
+ $X2=2.16 $Y2=1.84
r110 12 40 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=4.275 $Y=0.58
+ $X2=4.275 $Y2=1.19
r111 7 22 52.2586 $w=2.99e-07 $l=2.7157e-07 $layer=POLY_cond $X=3.275 $Y=1.885
+ $X2=3.32 $Y2=1.635
r112 7 9 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=3.275 $Y=1.885
+ $X2=3.275 $Y2=2.46
r113 2 36 600 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_PDIFF $count=1 $X=1.865
+ $Y=1.96 $X2=2.01 $Y2=2.145
r114 1 29 182 $w=1.7e-07 $l=6.68019e-07 $layer=licon1_NDIFF $count=1 $X=1.865
+ $Y=0.41 $X2=2.02 $Y2=1.005
.ends

.subckt PM_SKY130_FD_SC_HS__DLRTN_2%A_913_406# 1 2 7 9 12 14 15 16 19 20 22 25
+ 27 30 33 35 37 39 40 41 48 54 56 58 59 60 66 70
c130 60 0 3.65537e-20 $X=5.795 $Y=1.72
c131 56 0 7.28369e-20 $X=6.505 $Y=1.805
c132 20 0 1.03995e-19 $X=7.145 $Y=1.765
r133 67 70 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=6.68 $Y=1.485
+ $X2=6.68 $Y2=1.395
r134 66 68 14.5672 $w=2.68e-07 $l=3.2e-07 $layer=LI1_cond $X=6.675 $Y=1.485
+ $X2=6.675 $Y2=1.805
r135 66 67 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.68
+ $Y=1.485 $X2=6.68 $Y2=1.485
r136 63 64 5.33075 $w=4.98e-07 $l=1.65e-07 $layer=LI1_cond $X=5.795 $Y=2.195
+ $X2=5.795 $Y2=2.36
r137 62 63 5.02353 $w=4.98e-07 $l=2.1e-07 $layer=LI1_cond $X=5.795 $Y=1.985
+ $X2=5.795 $Y2=2.195
r138 59 62 4.30588 $w=4.98e-07 $l=1.8e-07 $layer=LI1_cond $X=5.795 $Y=1.805
+ $X2=5.795 $Y2=1.985
r139 59 60 7.60339 $w=4.98e-07 $l=8.5e-08 $layer=LI1_cond $X=5.795 $Y=1.805
+ $X2=5.795 $Y2=1.72
r140 58 60 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=5.63 $Y=1.13
+ $X2=5.63 $Y2=1.72
r141 57 59 7.15667 $w=1.7e-07 $l=2.5e-07 $layer=LI1_cond $X=6.045 $Y=1.805
+ $X2=5.795 $Y2=1.805
r142 56 68 3.40055 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=6.505 $Y=1.805
+ $X2=6.675 $Y2=1.805
r143 56 57 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=6.505 $Y=1.805
+ $X2=6.045 $Y2=1.805
r144 54 64 15.8897 $w=3.28e-07 $l=4.55e-07 $layer=LI1_cond $X=5.88 $Y=2.815
+ $X2=5.88 $Y2=2.36
r145 46 58 9.72165 $w=4.03e-07 $l=2.02e-07 $layer=LI1_cond $X=5.512 $Y=0.928
+ $X2=5.512 $Y2=1.13
r146 46 48 11.7521 $w=4.03e-07 $l=4.13e-07 $layer=LI1_cond $X=5.512 $Y=0.928
+ $X2=5.512 $Y2=0.515
r147 43 44 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.73
+ $Y=2.195 $X2=4.73 $Y2=2.195
r148 41 63 3.16914 $w=3.3e-07 $l=2.5e-07 $layer=LI1_cond $X=5.545 $Y=2.195
+ $X2=5.795 $Y2=2.195
r149 41 43 28.4618 $w=3.28e-07 $l=8.15e-07 $layer=LI1_cond $X=5.545 $Y=2.195
+ $X2=4.73 $Y2=2.195
r150 35 37 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=7.595 $Y=1.765
+ $X2=7.595 $Y2=2.4
r151 31 40 18.8402 $w=1.65e-07 $l=7.98436e-08 $layer=POLY_cond $X=7.585 $Y=1.32
+ $X2=7.595 $Y2=1.395
r152 31 33 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=7.585 $Y=1.32
+ $X2=7.585 $Y2=0.74
r153 30 35 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=7.595 $Y=1.675
+ $X2=7.595 $Y2=1.765
r154 29 40 18.8402 $w=1.65e-07 $l=7.5e-08 $layer=POLY_cond $X=7.595 $Y=1.47
+ $X2=7.595 $Y2=1.395
r155 29 30 79.6855 $w=1.8e-07 $l=2.05e-07 $layer=POLY_cond $X=7.595 $Y=1.47
+ $X2=7.595 $Y2=1.675
r156 28 39 13.2179 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=7.235 $Y=1.395
+ $X2=7.145 $Y2=1.395
r157 27 40 6.66866 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=7.505 $Y=1.395
+ $X2=7.595 $Y2=1.395
r158 27 28 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=7.505 $Y=1.395
+ $X2=7.235 $Y2=1.395
r159 23 39 10.9219 $w=1.5e-07 $l=7.98436e-08 $layer=POLY_cond $X=7.155 $Y=1.32
+ $X2=7.145 $Y2=1.395
r160 23 25 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=7.155 $Y=1.32
+ $X2=7.155 $Y2=0.74
r161 20 22 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=7.145 $Y=1.765
+ $X2=7.145 $Y2=2.4
r162 19 20 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=7.145 $Y=1.675
+ $X2=7.145 $Y2=1.765
r163 18 39 10.9219 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=7.145 $Y=1.47
+ $X2=7.145 $Y2=1.395
r164 18 19 79.6855 $w=1.8e-07 $l=2.05e-07 $layer=POLY_cond $X=7.145 $Y=1.47
+ $X2=7.145 $Y2=1.675
r165 17 70 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.845 $Y=1.395
+ $X2=6.68 $Y2=1.395
r166 16 39 13.2179 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=7.055 $Y=1.395
+ $X2=7.145 $Y2=1.395
r167 16 17 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=7.055 $Y=1.395
+ $X2=6.845 $Y2=1.395
r168 15 44 34.1752 $w=2.99e-07 $l=1.72337e-07 $layer=POLY_cond $X=4.715 $Y=2.03
+ $X2=4.73 $Y2=2.195
r169 14 38 37.1337 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=4.715 $Y=1.77
+ $X2=4.715 $Y2=1.68
r170 14 15 101.065 $w=1.8e-07 $l=2.6e-07 $layer=POLY_cond $X=4.715 $Y=1.77
+ $X2=4.715 $Y2=2.03
r171 12 38 564.043 $w=1.5e-07 $l=1.1e-06 $layer=POLY_cond $X=4.7 $Y=0.58 $X2=4.7
+ $Y2=1.68
r172 7 44 52.2586 $w=2.99e-07 $l=2.85044e-07 $layer=POLY_cond $X=4.655 $Y=2.445
+ $X2=4.73 $Y2=2.195
r173 7 9 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=4.655 $Y=2.445
+ $X2=4.655 $Y2=2.73
r174 2 62 400 $w=1.7e-07 $l=2.20907e-07 $layer=licon1_PDIFF $count=1 $X=5.72
+ $Y=1.84 $X2=5.88 $Y2=1.985
r175 2 54 400 $w=1.7e-07 $l=1.05196e-06 $layer=licon1_PDIFF $count=1 $X=5.72
+ $Y=1.84 $X2=5.88 $Y2=2.815
r176 1 48 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=5.33
+ $Y=0.37 $X2=5.475 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__DLRTN_2%A_670_392# 1 2 7 9 12 15 16 21 22 23 26 28
+ 29 33 35
c95 15 0 1.01066e-19 $X=5.555 $Y=1.515
c96 7 0 7.28369e-20 $X=5.645 $Y=1.765
r97 33 35 8.6688 $w=4.03e-07 $l=1.65e-07 $layer=LI1_cond $X=5.172 $Y=1.515
+ $X2=5.172 $Y2=1.35
r98 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.21
+ $Y=1.515 $X2=5.21 $Y2=1.515
r99 30 35 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=5.055 $Y=1.02
+ $X2=5.055 $Y2=1.35
r100 28 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.97 $Y=0.935
+ $X2=5.055 $Y2=1.02
r101 28 29 48.6043 $w=1.68e-07 $l=7.45e-07 $layer=LI1_cond $X=4.97 $Y=0.935
+ $X2=4.225 $Y2=0.935
r102 24 29 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.06 $Y=0.85
+ $X2=4.225 $Y2=0.935
r103 24 26 9.42908 $w=3.28e-07 $l=2.7e-07 $layer=LI1_cond $X=4.06 $Y=0.85
+ $X2=4.06 $Y2=0.58
r104 22 33 7.3984 $w=4.03e-07 $l=2.6e-07 $layer=LI1_cond $X=5.172 $Y=1.775
+ $X2=5.172 $Y2=1.515
r105 22 23 74.7005 $w=1.68e-07 $l=1.145e-06 $layer=LI1_cond $X=4.97 $Y=1.775
+ $X2=3.825 $Y2=1.775
r106 20 23 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.74 $Y=1.86
+ $X2=3.825 $Y2=1.775
r107 20 21 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=3.74 $Y=1.86
+ $X2=3.74 $Y2=2.18
r108 16 21 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.655 $Y=2.265
+ $X2=3.74 $Y2=2.18
r109 16 18 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=3.655 $Y=2.265
+ $X2=3.5 $Y2=2.265
r110 15 34 60.3271 $w=3.3e-07 $l=3.45e-07 $layer=POLY_cond $X=5.555 $Y=1.515
+ $X2=5.21 $Y2=1.515
r111 10 15 44.1289 $w=1.9e-07 $l=1.79374e-07 $layer=POLY_cond $X=5.69 $Y=1.35
+ $X2=5.66 $Y2=1.515
r112 10 12 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=5.69 $Y=1.35
+ $X2=5.69 $Y2=0.74
r113 7 15 65.692 $w=1.9e-07 $l=2.57391e-07 $layer=POLY_cond $X=5.645 $Y=1.765
+ $X2=5.66 $Y2=1.515
r114 7 9 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=5.645 $Y=1.765
+ $X2=5.645 $Y2=2.4
r115 2 18 600 $w=1.7e-07 $l=3.72525e-07 $layer=licon1_PDIFF $count=1 $X=3.35
+ $Y=1.96 $X2=3.5 $Y2=2.265
r116 1 26 182 $w=1.7e-07 $l=2.8801e-07 $layer=licon1_NDIFF $count=1 $X=3.875
+ $Y=0.37 $X2=4.06 $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_HS__DLRTN_2%RESET_B 1 3 4 6 7 11
c30 1 0 3.65537e-20 $X=6.08 $Y=1.22
r31 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.14
+ $Y=1.385 $X2=6.14 $Y2=1.385
r32 7 11 4.3606 $w=3.68e-07 $l=1.4e-07 $layer=LI1_cond $X=6 $Y=1.365 $X2=6.14
+ $Y2=1.365
r33 4 10 77.2841 $w=2.7e-07 $l=3.97115e-07 $layer=POLY_cond $X=6.105 $Y=1.765
+ $X2=6.14 $Y2=1.385
r34 4 6 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=6.105 $Y=1.765
+ $X2=6.105 $Y2=2.4
r35 1 10 38.9026 $w=2.7e-07 $l=1.92678e-07 $layer=POLY_cond $X=6.08 $Y=1.22
+ $X2=6.14 $Y2=1.385
r36 1 3 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=6.08 $Y=1.22 $X2=6.08
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HS__DLRTN_2%VPWR 1 2 3 4 5 18 22 26 28 30 35 36 37 43 55
+ 60 66 71 74 76 80
r81 79 80 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r82 76 77 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r83 73 74 11.3415 $w=7.83e-07 $l=1.65e-07 $layer=LI1_cond $X=5.38 $Y=3.022
+ $X2=5.545 $Y2=3.022
r84 69 73 5.18047 $w=7.83e-07 $l=3.4e-07 $layer=LI1_cond $X=5.04 $Y=3.022
+ $X2=5.38 $Y2=3.022
r85 69 71 13.7794 $w=7.83e-07 $l=3.25e-07 $layer=LI1_cond $X=5.04 $Y=3.022
+ $X2=4.715 $Y2=3.022
r86 69 70 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r87 66 67 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r88 64 80 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=7.92 $Y2=3.33
r89 64 77 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=6.48 $Y2=3.33
r90 63 64 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r91 61 76 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.65 $Y=3.33
+ $X2=6.485 $Y2=3.33
r92 61 63 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=6.65 $Y=3.33
+ $X2=7.44 $Y2=3.33
r93 60 79 4.82984 $w=1.7e-07 $l=2.27e-07 $layer=LI1_cond $X=7.705 $Y=3.33
+ $X2=7.932 $Y2=3.33
r94 60 63 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=7.705 $Y=3.33
+ $X2=7.44 $Y2=3.33
r95 59 77 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=3.33 $X2=6.48
+ $Y2=3.33
r96 59 70 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6 $Y=3.33 $X2=5.04
+ $Y2=3.33
r97 58 74 29.6845 $w=1.68e-07 $l=4.55e-07 $layer=LI1_cond $X=6 $Y=3.33 $X2=5.545
+ $Y2=3.33
r98 58 59 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r99 55 76 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.32 $Y=3.33
+ $X2=6.485 $Y2=3.33
r100 55 58 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=6.32 $Y=3.33 $X2=6
+ $Y2=3.33
r101 54 70 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=5.04 $Y2=3.33
r102 53 71 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=4.56 $Y=3.33
+ $X2=4.715 $Y2=3.33
r103 53 54 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r104 51 66 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.71 $Y=3.33
+ $X2=2.545 $Y2=3.33
r105 51 53 120.695 $w=1.68e-07 $l=1.85e-06 $layer=LI1_cond $X=2.71 $Y=3.33
+ $X2=4.56 $Y2=3.33
r106 49 67 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r107 48 49 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r108 46 49 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.16 $Y2=3.33
r109 45 48 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.2 $Y=3.33 $X2=2.16
+ $Y2=3.33
r110 45 46 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r111 43 66 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.38 $Y=3.33
+ $X2=2.545 $Y2=3.33
r112 43 48 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=2.38 $Y=3.33
+ $X2=2.16 $Y2=3.33
r113 41 46 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r114 40 41 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r115 37 54 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=4.56 $Y2=3.33
r116 37 67 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=2.64 $Y2=3.33
r117 35 40 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=0.785 $Y=3.33
+ $X2=0.72 $Y2=3.33
r118 35 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.785 $Y=3.33
+ $X2=0.95 $Y2=3.33
r119 34 45 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=1.115 $Y=3.33
+ $X2=1.2 $Y2=3.33
r120 34 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.115 $Y=3.33
+ $X2=0.95 $Y2=3.33
r121 30 33 28.1332 $w=3.38e-07 $l=8.3e-07 $layer=LI1_cond $X=7.875 $Y=1.985
+ $X2=7.875 $Y2=2.815
r122 28 79 3.02131 $w=3.4e-07 $l=1.09864e-07 $layer=LI1_cond $X=7.875 $Y=3.245
+ $X2=7.932 $Y2=3.33
r123 28 33 14.575 $w=3.38e-07 $l=4.3e-07 $layer=LI1_cond $X=7.875 $Y=3.245
+ $X2=7.875 $Y2=2.815
r124 24 76 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.485 $Y=3.245
+ $X2=6.485 $Y2=3.33
r125 24 26 35.621 $w=3.28e-07 $l=1.02e-06 $layer=LI1_cond $X=6.485 $Y=3.245
+ $X2=6.485 $Y2=2.225
r126 20 66 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.545 $Y=3.245
+ $X2=2.545 $Y2=3.33
r127 20 22 7.68295 $w=3.28e-07 $l=2.2e-07 $layer=LI1_cond $X=2.545 $Y=3.245
+ $X2=2.545 $Y2=3.025
r128 16 36 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.95 $Y=3.245
+ $X2=0.95 $Y2=3.33
r129 16 18 39.4624 $w=3.28e-07 $l=1.13e-06 $layer=LI1_cond $X=0.95 $Y=3.245
+ $X2=0.95 $Y2=2.115
r130 5 33 400 $w=1.7e-07 $l=1.07261e-06 $layer=licon1_PDIFF $count=1 $X=7.67
+ $Y=1.84 $X2=7.875 $Y2=2.815
r131 5 30 400 $w=1.7e-07 $l=2.67862e-07 $layer=licon1_PDIFF $count=1 $X=7.67
+ $Y=1.84 $X2=7.875 $Y2=1.985
r132 4 26 300 $w=1.7e-07 $l=5.15412e-07 $layer=licon1_PDIFF $count=2 $X=6.18
+ $Y=1.84 $X2=6.485 $Y2=2.225
r133 3 73 300 $w=1.7e-07 $l=7.75403e-07 $layer=licon1_PDIFF $count=2 $X=4.73
+ $Y=2.52 $X2=5.38 $Y2=2.795
r134 2 22 600 $w=1.7e-07 $l=1.17665e-06 $layer=licon1_PDIFF $count=1 $X=2.31
+ $Y=1.96 $X2=2.545 $Y2=3.025
r135 1 18 300 $w=1.7e-07 $l=2.62678e-07 $layer=licon1_PDIFF $count=2 $X=0.75
+ $Y=1.97 $X2=0.95 $Y2=2.115
.ends

.subckt PM_SKY130_FD_SC_HS__DLRTN_2%Q 1 2 9 13 14 15 16 29 30
c36 30 0 1.03995e-19 $X=7.19 $Y=1.82
r37 29 30 10.7408 $w=6.88e-07 $l=1.65e-07 $layer=LI1_cond $X=7.19 $Y=1.985
+ $X2=7.19 $Y2=1.82
r38 16 26 0.693379 $w=6.88e-07 $l=4e-08 $layer=LI1_cond $X=7.19 $Y=2.775
+ $X2=7.19 $Y2=2.815
r39 15 16 6.41375 $w=6.88e-07 $l=3.7e-07 $layer=LI1_cond $X=7.19 $Y=2.405
+ $X2=7.19 $Y2=2.775
r40 15 20 4.16027 $w=6.88e-07 $l=2.4e-07 $layer=LI1_cond $X=7.19 $Y=2.405
+ $X2=7.19 $Y2=2.165
r41 14 20 2.25348 $w=6.88e-07 $l=1.3e-07 $layer=LI1_cond $X=7.19 $Y=2.035
+ $X2=7.19 $Y2=2.165
r42 14 29 0.866723 $w=6.88e-07 $l=5e-08 $layer=LI1_cond $X=7.19 $Y=2.035
+ $X2=7.19 $Y2=1.985
r43 13 30 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=7.45 $Y=1.47
+ $X2=7.45 $Y2=1.82
r44 7 13 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=7.37 $Y=1.305
+ $X2=7.37 $Y2=1.47
r45 7 9 27.5888 $w=3.28e-07 $l=7.9e-07 $layer=LI1_cond $X=7.37 $Y=1.305 $X2=7.37
+ $Y2=0.515
r46 2 29 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=7.22
+ $Y=1.84 $X2=7.37 $Y2=1.985
r47 2 26 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=7.22
+ $Y=1.84 $X2=7.37 $Y2=2.815
r48 1 9 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=7.23
+ $Y=0.37 $X2=7.37 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__DLRTN_2%VGND 1 2 3 4 5 18 22 24 26 28 30 43 51 56 63
+ 70 74 76 79 83
c75 18 0 1.01066e-19 $X=4.915 $Y=0.515
r76 82 83 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=0 $X2=7.92
+ $Y2=0
r77 79 80 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=0 $X2=6.48
+ $Y2=0
r78 76 77 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r79 72 74 9.36575 $w=4.93e-07 $l=1.6e-07 $layer=LI1_cond $X=3.12 $Y=0.162
+ $X2=3.28 $Y2=0.162
r80 72 73 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r81 69 72 0.120816 $w=4.93e-07 $l=5e-09 $layer=LI1_cond $X=3.115 $Y=0.162
+ $X2=3.12 $Y2=0.162
r82 69 70 23.2596 $w=4.93e-07 $l=7.35e-07 $layer=LI1_cond $X=3.115 $Y=0.162
+ $X2=2.38 $Y2=0.162
r83 63 66 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=0.79 $Y=0 $X2=0.79
+ $Y2=0.325
r84 63 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r85 60 83 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=0 $X2=7.92
+ $Y2=0
r86 60 80 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=7.44 $Y=0 $X2=6.48
+ $Y2=0
r87 59 60 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.44 $Y=0 $X2=7.44
+ $Y2=0
r88 57 79 15.5458 $w=1.7e-07 $l=4.53e-07 $layer=LI1_cond $X=7.035 $Y=0 $X2=6.582
+ $Y2=0
r89 57 59 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=7.035 $Y=0 $X2=7.44
+ $Y2=0
r90 56 82 4.71369 $w=1.7e-07 $l=2.27e-07 $layer=LI1_cond $X=7.705 $Y=0 $X2=7.932
+ $Y2=0
r91 56 59 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=7.705 $Y=0 $X2=7.44
+ $Y2=0
r92 55 80 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=0 $X2=6.48
+ $Y2=0
r93 55 77 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6 $Y=0 $X2=5.04
+ $Y2=0
r94 54 55 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6 $Y=0 $X2=6 $Y2=0
r95 52 76 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.08 $Y=0 $X2=4.915
+ $Y2=0
r96 52 54 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=5.08 $Y=0 $X2=6
+ $Y2=0
r97 51 79 15.5458 $w=1.7e-07 $l=4.52e-07 $layer=LI1_cond $X=6.13 $Y=0 $X2=6.582
+ $Y2=0
r98 51 54 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=6.13 $Y=0 $X2=6
+ $Y2=0
r99 50 77 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=5.04
+ $Y2=0
r100 49 50 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r101 47 73 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=3.12
+ $Y2=0
r102 46 49 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=3.6 $Y=0 $X2=4.56
+ $Y2=0
r103 46 74 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=3.6 $Y=0 $X2=3.28
+ $Y2=0
r104 46 47 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r105 43 76 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.75 $Y=0 $X2=4.915
+ $Y2=0
r106 43 49 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=4.75 $Y=0 $X2=4.56
+ $Y2=0
r107 42 73 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=3.12
+ $Y2=0
r108 41 70 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=2.16 $Y=0 $X2=2.38
+ $Y2=0
r109 41 42 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r110 39 42 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r111 39 64 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r112 38 41 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r113 38 39 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r114 36 63 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.955 $Y=0 $X2=0.79
+ $Y2=0
r115 36 38 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=0.955 $Y=0 $X2=1.2
+ $Y2=0
r116 33 64 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r117 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r118 30 63 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.625 $Y=0 $X2=0.79
+ $Y2=0
r119 30 32 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=0.625 $Y=0
+ $X2=0.24 $Y2=0
r120 28 50 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=4.56
+ $Y2=0
r121 28 47 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=3.6
+ $Y2=0
r122 24 82 3.05248 $w=3.3e-07 $l=1.11781e-07 $layer=LI1_cond $X=7.87 $Y=0.085
+ $X2=7.932 $Y2=0
r123 24 26 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=7.87 $Y=0.085
+ $X2=7.87 $Y2=0.515
r124 20 79 3.35974 $w=9.05e-07 $l=8.5e-08 $layer=LI1_cond $X=6.582 $Y=0.085
+ $X2=6.582 $Y2=0
r125 20 22 5.79669 $w=9.03e-07 $l=4.3e-07 $layer=LI1_cond $X=6.582 $Y=0.085
+ $X2=6.582 $Y2=0.515
r126 16 76 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.915 $Y=0.085
+ $X2=4.915 $Y2=0
r127 16 18 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=4.915 $Y=0.085
+ $X2=4.915 $Y2=0.515
r128 5 26 91 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=2 $X=7.66
+ $Y=0.37 $X2=7.87 $Y2=0.515
r129 4 22 45.5 $w=1.7e-07 $l=7.84156e-07 $layer=licon1_NDIFF $count=4 $X=6.155
+ $Y=0.37 $X2=6.87 $Y2=0.515
r130 3 18 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=4.775
+ $Y=0.37 $X2=4.915 $Y2=0.515
r131 2 69 91 $w=1.7e-07 $l=8.31414e-07 $layer=licon1_NDIFF $count=2 $X=2.325
+ $Y=0.41 $X2=3.115 $Y2=0.325
r132 1 66 182 $w=1.7e-07 $l=4.51802e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.68 $X2=0.79 $Y2=0.325
.ends

