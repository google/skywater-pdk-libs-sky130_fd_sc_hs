# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_hs__bufbuf_16
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_hs__bufbuf_16 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  12.96000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.300000 0.505000 1.780000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  4.401600 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT  5.635000 0.350000  5.885000 1.900000 ;
        RECT  5.660000 1.900000  5.885000 1.920000 ;
        RECT  5.660000 1.920000  5.990000 2.980000 ;
        RECT  6.535000 0.350000  6.780000 1.650000 ;
        RECT  6.610000 1.650000  6.780000 1.920000 ;
        RECT  6.610000 1.920000  6.940000 2.980000 ;
        RECT  7.385000 0.350000  7.680000 1.650000 ;
        RECT  7.510000 1.650000  7.680000 1.920000 ;
        RECT  7.510000 1.920000  7.840000 2.980000 ;
        RECT  8.285000 0.350000  8.580000 1.650000 ;
        RECT  8.410000 1.650000  8.580000 1.920000 ;
        RECT  8.410000 1.920000  8.740000 2.980000 ;
        RECT  9.215000 0.350000  9.480000 1.650000 ;
        RECT  9.310000 1.650000  9.480000 1.920000 ;
        RECT  9.310000 1.920000  9.640000 2.980000 ;
        RECT 10.145000 0.350000 10.395000 1.650000 ;
        RECT 10.210000 1.650000 10.395000 1.920000 ;
        RECT 10.210000 1.920000 10.540000 2.980000 ;
        RECT 11.110000 0.350000 11.325000 1.920000 ;
        RECT 11.110000 1.920000 11.440000 2.980000 ;
        RECT 12.015000 0.350000 12.345000 1.150000 ;
        RECT 12.060000 1.150000 12.345000 2.020000 ;
        RECT 12.060000 2.020000 12.390000 2.980000 ;
      LAYER mcon ;
        RECT  5.760000 1.950000  5.930000 2.120000 ;
        RECT  6.675000 1.950000  6.845000 2.120000 ;
        RECT  7.595000 1.950000  7.765000 2.120000 ;
        RECT  8.485000 1.950000  8.655000 2.120000 ;
        RECT  9.405000 1.950000  9.575000 2.120000 ;
        RECT 10.295000 1.950000 10.465000 2.120000 ;
        RECT 11.195000 1.950000 11.365000 2.120000 ;
        RECT 12.115000 1.950000 12.285000 2.120000 ;
      LAYER met1 ;
        RECT 5.700000 1.920000 12.380000 2.150000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT  0.000000 -0.085000 12.960000 0.085000 ;
        RECT  0.560000  0.085000  0.890000 0.790000 ;
        RECT  1.420000  0.085000  1.670000 0.790000 ;
        RECT  2.415000  0.085000  2.745000 1.130000 ;
        RECT  3.345000  0.085000  3.675000 0.810000 ;
        RECT  4.275000  0.085000  4.605000 0.810000 ;
        RECT  5.275000  0.085000  5.455000 1.130000 ;
        RECT  6.065000  0.085000  6.315000 1.130000 ;
        RECT  6.960000  0.085000  7.175000 1.130000 ;
        RECT  7.850000  0.085000  8.115000 1.130000 ;
        RECT  8.750000  0.085000  9.045000 1.130000 ;
        RECT  9.665000  0.085000  9.975000 1.130000 ;
        RECT 10.575000  0.085000 10.905000 1.130000 ;
        RECT 11.505000  0.085000 11.835000 1.130000 ;
        RECT 12.515000  0.085000 12.845000 1.130000 ;
      LAYER mcon ;
        RECT  0.155000 -0.085000  0.325000 0.085000 ;
        RECT  0.635000 -0.085000  0.805000 0.085000 ;
        RECT  1.115000 -0.085000  1.285000 0.085000 ;
        RECT  1.595000 -0.085000  1.765000 0.085000 ;
        RECT  2.075000 -0.085000  2.245000 0.085000 ;
        RECT  2.555000 -0.085000  2.725000 0.085000 ;
        RECT  3.035000 -0.085000  3.205000 0.085000 ;
        RECT  3.515000 -0.085000  3.685000 0.085000 ;
        RECT  3.995000 -0.085000  4.165000 0.085000 ;
        RECT  4.475000 -0.085000  4.645000 0.085000 ;
        RECT  4.955000 -0.085000  5.125000 0.085000 ;
        RECT  5.435000 -0.085000  5.605000 0.085000 ;
        RECT  5.915000 -0.085000  6.085000 0.085000 ;
        RECT  6.395000 -0.085000  6.565000 0.085000 ;
        RECT  6.875000 -0.085000  7.045000 0.085000 ;
        RECT  7.355000 -0.085000  7.525000 0.085000 ;
        RECT  7.835000 -0.085000  8.005000 0.085000 ;
        RECT  8.315000 -0.085000  8.485000 0.085000 ;
        RECT  8.795000 -0.085000  8.965000 0.085000 ;
        RECT  9.275000 -0.085000  9.445000 0.085000 ;
        RECT  9.755000 -0.085000  9.925000 0.085000 ;
        RECT 10.235000 -0.085000 10.405000 0.085000 ;
        RECT 10.715000 -0.085000 10.885000 0.085000 ;
        RECT 11.195000 -0.085000 11.365000 0.085000 ;
        RECT 11.675000 -0.085000 11.845000 0.085000 ;
        RECT 12.155000 -0.085000 12.325000 0.085000 ;
        RECT 12.635000 -0.085000 12.805000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.245000 12.960000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT  0.000000 3.245000 12.960000 3.415000 ;
        RECT  0.645000 2.290000  0.815000 3.245000 ;
        RECT  1.545000 2.140000  1.715000 3.245000 ;
        RECT  2.490000 1.820000  2.740000 3.245000 ;
        RECT  3.470000 2.160000  3.640000 3.245000 ;
        RECT  4.370000 2.160000  4.540000 3.245000 ;
        RECT  5.280000 1.925000  5.450000 3.245000 ;
        RECT  6.160000 1.925000  6.410000 3.245000 ;
        RECT  7.140000 1.925000  7.310000 3.245000 ;
        RECT  8.040000 1.925000  8.210000 3.245000 ;
        RECT  8.940000 1.925000  9.110000 3.245000 ;
        RECT  9.840000 1.925000 10.010000 3.245000 ;
        RECT 10.740000 1.925000 10.910000 3.245000 ;
        RECT 11.640000 1.925000 11.890000 3.245000 ;
        RECT 12.590000 1.820000 12.840000 3.245000 ;
      LAYER mcon ;
        RECT  0.155000 3.245000  0.325000 3.415000 ;
        RECT  0.635000 3.245000  0.805000 3.415000 ;
        RECT  1.115000 3.245000  1.285000 3.415000 ;
        RECT  1.595000 3.245000  1.765000 3.415000 ;
        RECT  2.075000 3.245000  2.245000 3.415000 ;
        RECT  2.555000 3.245000  2.725000 3.415000 ;
        RECT  3.035000 3.245000  3.205000 3.415000 ;
        RECT  3.515000 3.245000  3.685000 3.415000 ;
        RECT  3.995000 3.245000  4.165000 3.415000 ;
        RECT  4.475000 3.245000  4.645000 3.415000 ;
        RECT  4.955000 3.245000  5.125000 3.415000 ;
        RECT  5.435000 3.245000  5.605000 3.415000 ;
        RECT  5.915000 3.245000  6.085000 3.415000 ;
        RECT  6.395000 3.245000  6.565000 3.415000 ;
        RECT  6.875000 3.245000  7.045000 3.415000 ;
        RECT  7.355000 3.245000  7.525000 3.415000 ;
        RECT  7.835000 3.245000  8.005000 3.415000 ;
        RECT  8.315000 3.245000  8.485000 3.415000 ;
        RECT  8.795000 3.245000  8.965000 3.415000 ;
        RECT  9.275000 3.245000  9.445000 3.415000 ;
        RECT  9.755000 3.245000  9.925000 3.415000 ;
        RECT 10.235000 3.245000 10.405000 3.415000 ;
        RECT 10.715000 3.245000 10.885000 3.415000 ;
        RECT 11.195000 3.245000 11.365000 3.415000 ;
        RECT 11.675000 3.245000 11.845000 3.415000 ;
        RECT 12.155000 3.245000 12.325000 3.415000 ;
        RECT 12.635000 3.245000 12.805000 3.415000 ;
      LAYER met1 ;
        RECT 0.000000 3.085000 12.960000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.115000 1.950000  0.845000 2.120000 ;
      RECT  0.115000 2.120000  0.445000 2.980000 ;
      RECT  0.130000 0.350000  0.380000 0.960000 ;
      RECT  0.130000 0.960000  0.845000 1.130000 ;
      RECT  0.675000 1.130000  0.845000 1.300000 ;
      RECT  0.675000 1.300000  1.875000 1.630000 ;
      RECT  0.675000 1.630000  0.845000 1.950000 ;
      RECT  1.015000 1.800000  2.245000 1.970000 ;
      RECT  1.015000 1.970000  1.345000 2.980000 ;
      RECT  1.070000 0.350000  1.240000 0.960000 ;
      RECT  1.070000 0.960000  2.215000 1.130000 ;
      RECT  1.855000 0.350000  2.215000 0.960000 ;
      RECT  1.915000 1.970000  2.245000 2.980000 ;
      RECT  2.045000 1.130000  2.215000 1.320000 ;
      RECT  2.045000 1.320000  4.480000 1.650000 ;
      RECT  2.045000 1.650000  2.245000 1.800000 ;
      RECT  2.915000 0.350000  3.165000 0.980000 ;
      RECT  2.915000 0.980000  5.105000 1.150000 ;
      RECT  2.940000 1.820000  5.080000 1.990000 ;
      RECT  2.940000 1.990000  3.270000 2.980000 ;
      RECT  3.840000 1.990000  4.170000 2.980000 ;
      RECT  3.845000 0.350000  4.095000 0.980000 ;
      RECT  4.750000 1.990000  5.080000 2.980000 ;
      RECT  4.775000 0.350000  5.025000 0.980000 ;
      RECT  4.845000 1.150000  5.105000 1.320000 ;
      RECT  4.845000 1.320000  5.405000 1.755000 ;
      RECT  4.845000 1.755000  5.080000 1.820000 ;
      RECT  6.055000 1.320000  6.365000 1.750000 ;
      RECT  6.950000 1.320000  7.215000 1.750000 ;
      RECT  7.850000 1.320000  8.115000 1.750000 ;
      RECT  8.750000 1.320000  9.045000 1.750000 ;
      RECT  9.650000 1.320000  9.975000 1.750000 ;
      RECT 10.565000 1.320000 10.940000 1.750000 ;
      RECT 11.495000 1.320000 11.890000 1.750000 ;
    LAYER mcon ;
      RECT  5.180000 1.580000  5.350000 1.750000 ;
      RECT  6.125000 1.580000  6.295000 1.750000 ;
      RECT  7.000000 1.580000  7.170000 1.750000 ;
      RECT  7.900000 1.580000  8.070000 1.750000 ;
      RECT  8.820000 1.580000  8.990000 1.750000 ;
      RECT  9.730000 1.580000  9.900000 1.750000 ;
      RECT 10.675000 1.580000 10.845000 1.750000 ;
      RECT 11.600000 1.580000 11.770000 1.750000 ;
    LAYER met1 ;
      RECT 5.110000 1.550000 11.830000 1.780000 ;
  END
END sky130_fd_sc_hs__bufbuf_16
