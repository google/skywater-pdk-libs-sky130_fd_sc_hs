* File: sky130_fd_sc_hs__nand3_4.pex.spice
* Created: Tue Sep  1 20:09:24 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HS__NAND3_4%A 1 3 4 6 7 9 10 12 13 15 16 18 19 20 32 33
c62 32 0 7.45181e-20 $X=1.37 $Y=1.515
r63 31 33 12.1952 $w=4.15e-07 $l=1.05e-07 $layer=POLY_cond $X=1.37 $Y=1.495
+ $X2=1.475 $Y2=1.495
r64 31 32 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.37
+ $Y=1.515 $X2=1.37 $Y2=1.515
r65 29 31 2.90361 $w=4.15e-07 $l=2.5e-08 $layer=POLY_cond $X=1.345 $Y=1.495
+ $X2=1.37 $Y2=1.495
r66 28 29 49.9422 $w=4.15e-07 $l=4.3e-07 $layer=POLY_cond $X=0.915 $Y=1.495
+ $X2=1.345 $Y2=1.495
r67 26 28 26.1325 $w=4.15e-07 $l=2.25e-07 $layer=POLY_cond $X=0.69 $Y=1.495
+ $X2=0.915 $Y2=1.495
r68 26 27 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=0.69
+ $Y=1.515 $X2=0.69 $Y2=1.515
r69 24 26 21.4867 $w=4.15e-07 $l=1.85e-07 $layer=POLY_cond $X=0.505 $Y=1.495
+ $X2=0.69 $Y2=1.495
r70 23 24 2.32289 $w=4.15e-07 $l=2e-08 $layer=POLY_cond $X=0.485 $Y=1.495
+ $X2=0.505 $Y2=1.495
r71 20 32 4.55617 $w=4.28e-07 $l=1.7e-07 $layer=LI1_cond $X=1.2 $Y=1.565
+ $X2=1.37 $Y2=1.565
r72 19 20 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=0.72 $Y=1.565
+ $X2=1.2 $Y2=1.565
r73 19 27 0.80403 $w=4.28e-07 $l=3e-08 $layer=LI1_cond $X=0.72 $Y=1.565 $X2=0.69
+ $Y2=1.565
r74 16 33 34.8434 $w=4.15e-07 $l=4.13521e-07 $layer=POLY_cond $X=1.775 $Y=1.225
+ $X2=1.475 $Y2=1.495
r75 16 18 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=1.775 $Y=1.225
+ $X2=1.775 $Y2=0.78
r76 13 33 26.7644 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=1.475 $Y=1.765
+ $X2=1.475 $Y2=1.495
r77 13 15 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.475 $Y=1.765
+ $X2=1.475 $Y2=2.4
r78 10 29 26.7644 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=1.345 $Y=1.225
+ $X2=1.345 $Y2=1.495
r79 10 12 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=1.345 $Y=1.225
+ $X2=1.345 $Y2=0.78
r80 7 28 26.7644 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=0.915 $Y=1.225
+ $X2=0.915 $Y2=1.495
r81 7 9 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=0.915 $Y=1.225
+ $X2=0.915 $Y2=0.78
r82 4 24 26.7644 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=0.505 $Y=1.765
+ $X2=0.505 $Y2=1.495
r83 4 6 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.505 $Y=1.765
+ $X2=0.505 $Y2=2.4
r84 1 23 26.7644 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=0.485 $Y=1.225
+ $X2=0.485 $Y2=1.495
r85 1 3 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=0.485 $Y=1.225
+ $X2=0.485 $Y2=0.78
.ends

.subckt PM_SKY130_FD_SC_HS__NAND3_4%B 1 3 6 8 10 13 17 21 28 32 33 34 45
c66 45 0 1.88335e-19 $X=3.405 $Y=1.515
c67 21 0 4.53359e-20 $X=3.495 $Y=0.78
c68 17 0 1.20944e-20 $X=3.065 $Y=0.78
c69 6 0 1.07122e-19 $X=2.205 $Y=0.78
c70 1 0 7.45181e-20 $X=1.975 $Y=1.765
r71 45 47 11.5372 $w=3.76e-07 $l=9e-08 $layer=POLY_cond $X=3.405 $Y=1.557
+ $X2=3.495 $Y2=1.557
r72 45 46 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.405
+ $Y=1.515 $X2=3.405 $Y2=1.515
r73 43 45 43.5851 $w=3.76e-07 $l=3.4e-07 $layer=POLY_cond $X=3.065 $Y=1.557
+ $X2=3.405 $Y2=1.557
r74 40 41 26.9202 $w=3.76e-07 $l=2.1e-07 $layer=POLY_cond $X=2.425 $Y=1.557
+ $X2=2.635 $Y2=1.557
r75 34 46 5.22619 $w=4.28e-07 $l=1.95e-07 $layer=LI1_cond $X=3.6 $Y=1.565
+ $X2=3.405 $Y2=1.565
r76 33 46 7.63829 $w=4.28e-07 $l=2.85e-07 $layer=LI1_cond $X=3.12 $Y=1.565
+ $X2=3.405 $Y2=1.565
r77 31 43 43.5851 $w=3.76e-07 $l=3.4e-07 $layer=POLY_cond $X=2.725 $Y=1.557
+ $X2=3.065 $Y2=1.557
r78 31 41 11.5372 $w=3.76e-07 $l=9e-08 $layer=POLY_cond $X=2.725 $Y=1.557
+ $X2=2.635 $Y2=1.557
r79 30 32 5.82291 $w=4.28e-07 $l=1.65e-07 $layer=LI1_cond $X=2.725 $Y=1.565
+ $X2=2.56 $Y2=1.565
r80 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.725
+ $Y=1.515 $X2=2.725 $Y2=1.515
r81 28 33 3.48413 $w=4.28e-07 $l=1.3e-07 $layer=LI1_cond $X=2.99 $Y=1.565
+ $X2=3.12 $Y2=1.565
r82 28 30 7.10226 $w=4.28e-07 $l=2.65e-07 $layer=LI1_cond $X=2.99 $Y=1.565
+ $X2=2.725 $Y2=1.565
r83 26 40 16.6649 $w=3.76e-07 $l=1.3e-07 $layer=POLY_cond $X=2.295 $Y=1.557
+ $X2=2.425 $Y2=1.557
r84 26 38 11.5372 $w=3.76e-07 $l=9e-08 $layer=POLY_cond $X=2.295 $Y=1.557
+ $X2=2.205 $Y2=1.557
r85 25 32 10.9071 $w=2.78e-07 $l=2.65e-07 $layer=LI1_cond $X=2.295 $Y=1.49
+ $X2=2.56 $Y2=1.49
r86 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.295
+ $Y=1.515 $X2=2.295 $Y2=1.515
r87 19 47 24.356 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.495 $Y=1.35
+ $X2=3.495 $Y2=1.557
r88 19 21 292.277 $w=1.5e-07 $l=5.7e-07 $layer=POLY_cond $X=3.495 $Y=1.35
+ $X2=3.495 $Y2=0.78
r89 15 43 24.356 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.065 $Y=1.35
+ $X2=3.065 $Y2=1.557
r90 15 17 292.277 $w=1.5e-07 $l=5.7e-07 $layer=POLY_cond $X=3.065 $Y=1.35
+ $X2=3.065 $Y2=0.78
r91 11 41 24.356 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.635 $Y=1.35
+ $X2=2.635 $Y2=1.557
r92 11 13 292.277 $w=1.5e-07 $l=5.7e-07 $layer=POLY_cond $X=2.635 $Y=1.35
+ $X2=2.635 $Y2=0.78
r93 8 40 24.356 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=2.425 $Y=1.765
+ $X2=2.425 $Y2=1.557
r94 8 10 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.425 $Y=1.765
+ $X2=2.425 $Y2=2.4
r95 4 38 24.356 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.205 $Y=1.35
+ $X2=2.205 $Y2=1.557
r96 4 6 292.277 $w=1.5e-07 $l=5.7e-07 $layer=POLY_cond $X=2.205 $Y=1.35
+ $X2=2.205 $Y2=0.78
r97 1 38 29.484 $w=3.76e-07 $l=3.17396e-07 $layer=POLY_cond $X=1.975 $Y=1.765
+ $X2=2.205 $Y2=1.557
r98 1 3 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.975 $Y=1.765
+ $X2=1.975 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_HS__NAND3_4%C 1 3 4 6 9 13 17 21 28 32 33 34 35 50
c64 32 0 2.21572e-19 $X=4.495 $Y=1.56
c65 21 0 1.6164e-19 $X=5.755 $Y=0.78
r66 50 52 12.5376 $w=3.46e-07 $l=9e-08 $layer=POLY_cond $X=5.665 $Y=1.552
+ $X2=5.755 $Y2=1.552
r67 50 51 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=5.665
+ $Y=1.505 $X2=5.665 $Y2=1.505
r68 48 50 47.3642 $w=3.46e-07 $l=3.4e-07 $layer=POLY_cond $X=5.325 $Y=1.552
+ $X2=5.665 $Y2=1.552
r69 46 48 47.3642 $w=3.46e-07 $l=3.4e-07 $layer=POLY_cond $X=4.985 $Y=1.552
+ $X2=5.325 $Y2=1.552
r70 46 47 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=4.985
+ $Y=1.505 $X2=4.985 $Y2=1.505
r71 44 46 12.5376 $w=3.46e-07 $l=9e-08 $layer=POLY_cond $X=4.895 $Y=1.552
+ $X2=4.985 $Y2=1.552
r72 41 42 16.0202 $w=3.46e-07 $l=1.15e-07 $layer=POLY_cond $X=4.35 $Y=1.552
+ $X2=4.465 $Y2=1.552
r73 35 51 8.77428 $w=4.38e-07 $l=3.35e-07 $layer=LI1_cond $X=6 $Y=1.56 $X2=5.665
+ $Y2=1.56
r74 34 51 3.79782 $w=4.38e-07 $l=1.45e-07 $layer=LI1_cond $X=5.52 $Y=1.56
+ $X2=5.665 $Y2=1.56
r75 33 34 12.5721 $w=4.38e-07 $l=4.8e-07 $layer=LI1_cond $X=5.04 $Y=1.56
+ $X2=5.52 $Y2=1.56
r76 33 47 1.44055 $w=4.38e-07 $l=5.5e-08 $layer=LI1_cond $X=5.04 $Y=1.56
+ $X2=4.985 $Y2=1.56
r77 31 44 34.8266 $w=3.46e-07 $l=2.5e-07 $layer=POLY_cond $X=4.645 $Y=1.552
+ $X2=4.895 $Y2=1.552
r78 31 42 25.0751 $w=3.46e-07 $l=1.8e-07 $layer=POLY_cond $X=4.645 $Y=1.552
+ $X2=4.465 $Y2=1.552
r79 30 32 5.26886 $w=4.38e-07 $l=1.5e-07 $layer=LI1_cond $X=4.645 $Y=1.56
+ $X2=4.495 $Y2=1.56
r80 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.645
+ $Y=1.505 $X2=4.645 $Y2=1.505
r81 28 47 1.30959 $w=4.38e-07 $l=5e-08 $layer=LI1_cond $X=4.935 $Y=1.56
+ $X2=4.985 $Y2=1.56
r82 28 30 7.59565 $w=4.38e-07 $l=2.9e-07 $layer=LI1_cond $X=4.935 $Y=1.56
+ $X2=4.645 $Y2=1.56
r83 26 41 6.26879 $w=3.46e-07 $l=4.5e-08 $layer=POLY_cond $X=4.305 $Y=1.552
+ $X2=4.35 $Y2=1.552
r84 26 39 56.4191 $w=3.46e-07 $l=4.05e-07 $layer=POLY_cond $X=4.305 $Y=1.552
+ $X2=3.9 $Y2=1.552
r85 25 32 7.55049 $w=2.88e-07 $l=1.9e-07 $layer=LI1_cond $X=4.305 $Y=1.485
+ $X2=4.495 $Y2=1.485
r86 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.305
+ $Y=1.505 $X2=4.305 $Y2=1.505
r87 19 52 22.3532 $w=1.5e-07 $l=2.12e-07 $layer=POLY_cond $X=5.755 $Y=1.34
+ $X2=5.755 $Y2=1.552
r88 19 21 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=5.755 $Y=1.34
+ $X2=5.755 $Y2=0.78
r89 15 48 22.3532 $w=1.5e-07 $l=2.12e-07 $layer=POLY_cond $X=5.325 $Y=1.34
+ $X2=5.325 $Y2=1.552
r90 15 17 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=5.325 $Y=1.34
+ $X2=5.325 $Y2=0.78
r91 11 44 22.3532 $w=1.5e-07 $l=2.12e-07 $layer=POLY_cond $X=4.895 $Y=1.34
+ $X2=4.895 $Y2=1.552
r92 11 13 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=4.895 $Y=1.34
+ $X2=4.895 $Y2=0.78
r93 7 42 22.3532 $w=1.5e-07 $l=2.12e-07 $layer=POLY_cond $X=4.465 $Y=1.34
+ $X2=4.465 $Y2=1.552
r94 7 9 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=4.465 $Y=1.34
+ $X2=4.465 $Y2=0.78
r95 4 41 22.3532 $w=1.5e-07 $l=2.13e-07 $layer=POLY_cond $X=4.35 $Y=1.765
+ $X2=4.35 $Y2=1.552
r96 4 6 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=4.35 $Y=1.765
+ $X2=4.35 $Y2=2.4
r97 1 39 22.3532 $w=1.5e-07 $l=2.13e-07 $layer=POLY_cond $X=3.9 $Y=1.765 $X2=3.9
+ $Y2=1.552
r98 1 3 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.9 $Y=1.765 $X2=3.9
+ $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_HS__NAND3_4%VPWR 1 2 3 4 13 15 19 21 23 33 40 41 47 52
+ 60 62
r54 71 73 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=5.52 $Y2=3.33
r55 65 68 3.36552 $w=1.303e-06 $l=3.6e-07 $layer=LI1_cond $X=5.112 $Y=2.455
+ $X2=5.112 $Y2=2.815
r56 62 65 3.17854 $w=1.303e-06 $l=3.4e-07 $layer=LI1_cond $X=5.112 $Y=2.115
+ $X2=5.112 $Y2=2.455
r57 59 60 13.0375 $w=1.123e-06 $l=1.2e-07 $layer=LI1_cond $X=3.67 $Y=2.852
+ $X2=3.79 $Y2=2.852
r58 56 59 0.759111 $w=1.123e-06 $l=7e-08 $layer=LI1_cond $X=3.6 $Y=2.852
+ $X2=3.67 $Y2=2.852
r59 56 57 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r60 54 56 10.248 $w=1.123e-06 $l=9.45e-07 $layer=LI1_cond $X=2.655 $Y=2.852
+ $X2=3.6 $Y2=2.852
r61 50 54 0.162667 $w=1.123e-06 $l=1.5e-08 $layer=LI1_cond $X=2.64 $Y=2.852
+ $X2=2.655 $Y2=2.852
r62 50 52 12.8748 $w=1.123e-06 $l=1.05e-07 $layer=LI1_cond $X=2.64 $Y=2.852
+ $X2=2.535 $Y2=2.852
r63 50 51 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r64 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r65 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r66 41 73 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=3.33 $X2=5.52
+ $Y2=3.33
r67 40 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r68 38 40 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=5.765 $Y=3.33 $X2=6
+ $Y2=3.33
r69 37 71 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=4.56 $Y2=3.33
r70 37 57 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=3.6 $Y2=3.33
r71 36 60 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=4.08 $Y=3.33
+ $X2=3.79 $Y2=3.33
r72 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r73 33 38 13.5804 $w=1.7e-07 $l=6.53e-07 $layer=LI1_cond $X=5.112 $Y=3.33
+ $X2=5.765 $Y2=3.33
r74 33 73 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r75 33 71 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r76 33 68 4.81456 $w=1.303e-06 $l=5.15e-07 $layer=LI1_cond $X=5.112 $Y=3.33
+ $X2=5.112 $Y2=2.815
r77 33 36 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=4.46 $Y=3.33
+ $X2=4.08 $Y2=3.33
r78 32 51 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r79 32 48 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.68 $Y2=3.33
r80 31 52 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=2.16 $Y=3.33
+ $X2=2.535 $Y2=3.33
r81 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r82 29 47 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.865 $Y=3.33
+ $X2=1.7 $Y2=3.33
r83 29 31 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=1.865 $Y=3.33
+ $X2=2.16 $Y2=3.33
r84 27 48 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=1.68 $Y2=3.33
r85 27 45 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.24 $Y2=3.33
r86 26 27 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r87 24 44 4.73185 $w=1.7e-07 $l=2.23e-07 $layer=LI1_cond $X=0.445 $Y=3.33
+ $X2=0.222 $Y2=3.33
r88 24 26 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=0.445 $Y=3.33
+ $X2=1.2 $Y2=3.33
r89 23 47 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.535 $Y=3.33
+ $X2=1.7 $Y2=3.33
r90 23 26 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=1.535 $Y=3.33
+ $X2=1.2 $Y2=3.33
r91 21 57 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=3.6 $Y2=3.33
r92 21 51 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=2.64 $Y2=3.33
r93 17 47 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.7 $Y=3.245 $X2=1.7
+ $Y2=3.33
r94 17 19 27.5888 $w=3.28e-07 $l=7.9e-07 $layer=LI1_cond $X=1.7 $Y=3.245 $X2=1.7
+ $Y2=2.455
r95 13 44 3.03433 $w=3.3e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.28 $Y=3.245
+ $X2=0.222 $Y2=3.33
r96 13 15 29.6841 $w=3.28e-07 $l=8.5e-07 $layer=LI1_cond $X=0.28 $Y=3.245
+ $X2=0.28 $Y2=2.395
r97 4 68 200 $w=1.7e-07 $l=1.19718e-06 $layer=licon1_PDIFF $count=3 $X=4.425
+ $Y=1.84 $X2=4.92 $Y2=2.815
r98 4 65 200 $w=1.7e-07 $l=1.45026e-06 $layer=licon1_PDIFF $count=3 $X=4.425
+ $Y=1.84 $X2=5.6 $Y2=2.455
r99 4 65 200 $w=1.7e-07 $l=6.8815e-07 $layer=licon1_PDIFF $count=3 $X=4.425
+ $Y=1.84 $X2=4.58 $Y2=2.455
r100 4 62 200 $w=1.7e-07 $l=6.17373e-07 $layer=licon1_PDIFF $count=3 $X=4.425
+ $Y=1.84 $X2=4.92 $Y2=2.115
r101 3 59 200 $w=1.7e-07 $l=1.44515e-06 $layer=licon1_PDIFF $count=3 $X=2.5
+ $Y=1.84 $X2=3.67 $Y2=2.455
r102 3 54 200 $w=1.7e-07 $l=6.8815e-07 $layer=licon1_PDIFF $count=3 $X=2.5
+ $Y=1.84 $X2=2.655 $Y2=2.455
r103 2 19 300 $w=1.7e-07 $l=6.85912e-07 $layer=licon1_PDIFF $count=2 $X=1.55
+ $Y=1.84 $X2=1.7 $Y2=2.455
r104 1 15 300 $w=1.7e-07 $l=6.23298e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.395
.ends

.subckt PM_SKY130_FD_SC_HS__NAND3_4%Y 1 2 3 4 5 16 17 18 19 22 26 28 30 34 38 40
+ 42 44 48 50 52 55 56
c97 28 0 9.50231e-20 $X=1.395 $Y=1.095
r98 55 56 18.5393 $w=2.28e-07 $l=3.7e-07 $layer=LI1_cond $X=0.24 $Y=1.295
+ $X2=0.24 $Y2=1.665
r99 47 56 14.2803 $w=2.28e-07 $l=2.85e-07 $layer=LI1_cond $X=0.24 $Y=1.95
+ $X2=0.24 $Y2=1.665
r100 46 55 5.76222 $w=2.28e-07 $l=1.15e-07 $layer=LI1_cond $X=0.24 $Y=1.18
+ $X2=0.24 $Y2=1.295
r101 42 54 3.0656 $w=3.3e-07 $l=1.5e-07 $layer=LI1_cond $X=4.125 $Y=2.12
+ $X2=4.125 $Y2=1.97
r102 42 44 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=4.125 $Y=2.12
+ $X2=4.125 $Y2=2.815
r103 41 52 8.61065 $w=1.7e-07 $l=1.94808e-07 $layer=LI1_cond $X=2.365 $Y=2.035
+ $X2=2.2 $Y2=1.97
r104 40 54 4.70058 $w=1.7e-07 $l=1.94808e-07 $layer=LI1_cond $X=3.96 $Y=2.035
+ $X2=4.125 $Y2=1.97
r105 40 41 104.059 $w=1.68e-07 $l=1.595e-06 $layer=LI1_cond $X=3.96 $Y=2.035
+ $X2=2.365 $Y2=2.035
r106 36 52 0.89609 $w=3.3e-07 $l=1.5e-07 $layer=LI1_cond $X=2.2 $Y=2.12 $X2=2.2
+ $Y2=1.97
r107 36 38 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=2.2 $Y=2.12
+ $X2=2.2 $Y2=2.815
r108 32 34 11.5244 $w=3.28e-07 $l=3.3e-07 $layer=LI1_cond $X=1.56 $Y=1.01
+ $X2=1.56 $Y2=0.68
r109 31 50 14.1623 $w=1.7e-07 $l=3.75e-07 $layer=LI1_cond $X=1.365 $Y=2.035
+ $X2=0.99 $Y2=2.035
r110 30 52 8.61065 $w=1.7e-07 $l=1.94808e-07 $layer=LI1_cond $X=2.035 $Y=2.035
+ $X2=2.2 $Y2=1.97
r111 30 31 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.035 $Y=2.035
+ $X2=1.365 $Y2=2.035
r112 29 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.865 $Y=1.095
+ $X2=0.7 $Y2=1.095
r113 28 32 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.395 $Y=1.095
+ $X2=1.56 $Y2=1.01
r114 28 29 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=1.395 $Y=1.095
+ $X2=0.865 $Y2=1.095
r115 24 50 3.00456 $w=7.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.99 $Y=2.12
+ $X2=0.99 $Y2=2.035
r116 24 26 11.0837 $w=7.48e-07 $l=6.95e-07 $layer=LI1_cond $X=0.99 $Y=2.12
+ $X2=0.99 $Y2=2.815
r117 20 48 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.7 $Y=1.01 $X2=0.7
+ $Y2=1.095
r118 20 22 11.5244 $w=3.28e-07 $l=3.3e-07 $layer=LI1_cond $X=0.7 $Y=1.01 $X2=0.7
+ $Y2=0.68
r119 19 47 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=0.355 $Y=2.035
+ $X2=0.24 $Y2=1.95
r120 18 50 14.1623 $w=1.7e-07 $l=3.75e-07 $layer=LI1_cond $X=0.615 $Y=2.035
+ $X2=0.99 $Y2=2.035
r121 18 19 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=0.615 $Y=2.035
+ $X2=0.355 $Y2=2.035
r122 17 46 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=0.355 $Y=1.095
+ $X2=0.24 $Y2=1.18
r123 16 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.535 $Y=1.095
+ $X2=0.7 $Y2=1.095
r124 16 17 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=0.535 $Y=1.095
+ $X2=0.355 $Y2=1.095
r125 5 54 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=3.975
+ $Y=1.84 $X2=4.125 $Y2=1.985
r126 5 44 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=3.975
+ $Y=1.84 $X2=4.125 $Y2=2.815
r127 4 52 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=2.05
+ $Y=1.84 $X2=2.2 $Y2=1.985
r128 4 38 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=2.05
+ $Y=1.84 $X2=2.2 $Y2=2.815
r129 3 50 200 $w=1.7e-07 $l=3.43875e-07 $layer=licon1_PDIFF $count=3 $X=0.58
+ $Y=1.84 $X2=0.735 $Y2=2.115
r130 3 26 200 $w=1.7e-07 $l=1.04964e-06 $layer=licon1_PDIFF $count=3 $X=0.58
+ $Y=1.84 $X2=0.735 $Y2=2.815
r131 2 34 91 $w=1.7e-07 $l=3.32716e-07 $layer=licon1_NDIFF $count=2 $X=1.42
+ $Y=0.41 $X2=1.56 $Y2=0.68
r132 1 22 91 $w=1.7e-07 $l=3.32716e-07 $layer=licon1_NDIFF $count=2 $X=0.56
+ $Y=0.41 $X2=0.7 $Y2=0.68
.ends

.subckt PM_SKY130_FD_SC_HS__NAND3_4%A_27_82# 1 2 3 4 5 18 20 21 24 26 30 32 36
+ 38 42 44 45 46
r66 40 42 6.42709 $w=2.58e-07 $l=1.45e-07 $layer=LI1_cond $X=3.745 $Y=0.425
+ $X2=3.745 $Y2=0.57
r67 39 46 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=2.945 $Y=0.34
+ $X2=2.85 $Y2=0.34
r68 38 40 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=3.615 $Y=0.34
+ $X2=3.745 $Y2=0.425
r69 38 39 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.615 $Y=0.34
+ $X2=2.945 $Y2=0.34
r70 34 46 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=2.85 $Y=0.425
+ $X2=2.85 $Y2=0.34
r71 34 36 8.46412 $w=1.88e-07 $l=1.45e-07 $layer=LI1_cond $X=2.85 $Y=0.425
+ $X2=2.85 $Y2=0.57
r72 33 45 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.075 $Y=0.34
+ $X2=1.99 $Y2=0.34
r73 32 46 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=2.755 $Y=0.34
+ $X2=2.85 $Y2=0.34
r74 32 33 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=2.755 $Y=0.34
+ $X2=2.075 $Y2=0.34
r75 28 45 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.99 $Y=0.425
+ $X2=1.99 $Y2=0.34
r76 28 30 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=1.99 $Y=0.425
+ $X2=1.99 $Y2=0.555
r77 27 44 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.215 $Y=0.34
+ $X2=1.13 $Y2=0.34
r78 26 45 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.905 $Y=0.34
+ $X2=1.99 $Y2=0.34
r79 26 27 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.905 $Y=0.34
+ $X2=1.215 $Y2=0.34
r80 22 44 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.13 $Y=0.425
+ $X2=1.13 $Y2=0.34
r81 22 24 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=1.13 $Y=0.425
+ $X2=1.13 $Y2=0.615
r82 20 44 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.045 $Y=0.34
+ $X2=1.13 $Y2=0.34
r83 20 21 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.045 $Y=0.34
+ $X2=0.355 $Y2=0.34
r84 16 21 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.23 $Y=0.425
+ $X2=0.355 $Y2=0.34
r85 16 18 8.75857 $w=2.48e-07 $l=1.9e-07 $layer=LI1_cond $X=0.23 $Y=0.425
+ $X2=0.23 $Y2=0.615
r86 5 42 182 $w=1.7e-07 $l=2.19089e-07 $layer=licon1_NDIFF $count=1 $X=3.57
+ $Y=0.41 $X2=3.71 $Y2=0.57
r87 4 36 182 $w=1.7e-07 $l=2.19089e-07 $layer=licon1_NDIFF $count=1 $X=2.71
+ $Y=0.41 $X2=2.85 $Y2=0.57
r88 3 30 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.85
+ $Y=0.41 $X2=1.99 $Y2=0.555
r89 2 24 182 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_NDIFF $count=1 $X=0.99
+ $Y=0.41 $X2=1.13 $Y2=0.615
r90 1 18 182 $w=1.7e-07 $l=2.64008e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.41 $X2=0.27 $Y2=0.615
.ends

.subckt PM_SKY130_FD_SC_HS__NAND3_4%A_456_82# 1 2 3 4 13 15 19 21 23 25 28 33 38
c66 23 0 1.6164e-19 $X=5.54 $Y=0.92
c67 15 0 1.20944e-20 $X=4.585 $Y=1.045
c68 13 0 2.41975e-20 $X=3.115 $Y=1.045
r69 33 35 12.7467 $w=3.28e-07 $l=3.65e-07 $layer=LI1_cond $X=3.28 $Y=0.68
+ $X2=3.28 $Y2=1.045
r70 28 30 12.7467 $w=3.28e-07 $l=3.65e-07 $layer=LI1_cond $X=2.42 $Y=0.68
+ $X2=2.42 $Y2=1.045
r71 23 40 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.54 $Y=0.92
+ $X2=5.54 $Y2=1.045
r72 23 25 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=5.54 $Y=0.92
+ $X2=5.54 $Y2=0.555
r73 22 38 4.08801 $w=2.5e-07 $l=9.5e-08 $layer=LI1_cond $X=4.775 $Y=1.045
+ $X2=4.68 $Y2=1.045
r74 21 40 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.455 $Y=1.045
+ $X2=5.54 $Y2=1.045
r75 21 22 31.3464 $w=2.48e-07 $l=6.8e-07 $layer=LI1_cond $X=5.455 $Y=1.045
+ $X2=4.775 $Y2=1.045
r76 17 38 2.34704 $w=1.9e-07 $l=1.25e-07 $layer=LI1_cond $X=4.68 $Y=0.92
+ $X2=4.68 $Y2=1.045
r77 17 19 21.3062 $w=1.88e-07 $l=3.65e-07 $layer=LI1_cond $X=4.68 $Y=0.92
+ $X2=4.68 $Y2=0.555
r78 16 35 2.36532 $w=2.5e-07 $l=1.65e-07 $layer=LI1_cond $X=3.445 $Y=1.045
+ $X2=3.28 $Y2=1.045
r79 15 38 4.08801 $w=2.5e-07 $l=9.5e-08 $layer=LI1_cond $X=4.585 $Y=1.045
+ $X2=4.68 $Y2=1.045
r80 15 16 52.5514 $w=2.48e-07 $l=1.14e-06 $layer=LI1_cond $X=4.585 $Y=1.045
+ $X2=3.445 $Y2=1.045
r81 14 30 2.36532 $w=2.5e-07 $l=1.65e-07 $layer=LI1_cond $X=2.585 $Y=1.045
+ $X2=2.42 $Y2=1.045
r82 13 35 2.36532 $w=2.5e-07 $l=1.65e-07 $layer=LI1_cond $X=3.115 $Y=1.045
+ $X2=3.28 $Y2=1.045
r83 13 14 24.4318 $w=2.48e-07 $l=5.3e-07 $layer=LI1_cond $X=3.115 $Y=1.045
+ $X2=2.585 $Y2=1.045
r84 4 40 182 $w=1.7e-07 $l=6.61306e-07 $layer=licon1_NDIFF $count=1 $X=5.4
+ $Y=0.41 $X2=5.54 $Y2=1.005
r85 4 25 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=5.4
+ $Y=0.41 $X2=5.54 $Y2=0.555
r86 3 38 182 $w=1.7e-07 $l=6.61306e-07 $layer=licon1_NDIFF $count=1 $X=4.54
+ $Y=0.41 $X2=4.68 $Y2=1.005
r87 3 19 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=4.54
+ $Y=0.41 $X2=4.68 $Y2=0.555
r88 2 33 91 $w=1.7e-07 $l=3.32716e-07 $layer=licon1_NDIFF $count=2 $X=3.14
+ $Y=0.41 $X2=3.28 $Y2=0.68
r89 1 28 91 $w=1.7e-07 $l=3.32716e-07 $layer=licon1_NDIFF $count=2 $X=2.28
+ $Y=0.41 $X2=2.42 $Y2=0.68
.ends

.subckt PM_SKY130_FD_SC_HS__NAND3_4%VGND 1 2 3 12 16 18 20 23 24 25 34 38 44 48
r67 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=0 $X2=6 $Y2=0
r68 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r69 42 48 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=6
+ $Y2=0
r70 42 45 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=5.04
+ $Y2=0
r71 41 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r72 39 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.275 $Y=0 $X2=5.11
+ $Y2=0
r73 39 41 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=5.275 $Y=0 $X2=5.52
+ $Y2=0
r74 38 47 4.76062 $w=1.7e-07 $l=2.17e-07 $layer=LI1_cond $X=5.805 $Y=0 $X2=6.022
+ $Y2=0
r75 38 41 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=5.805 $Y=0 $X2=5.52
+ $Y2=0
r76 37 45 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=5.04
+ $Y2=0
r77 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r78 34 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.945 $Y=0 $X2=5.11
+ $Y2=0
r79 34 36 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=4.945 $Y=0 $X2=4.56
+ $Y2=0
r80 33 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=4.56
+ $Y2=0
r81 32 33 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=4.08 $Y=0
+ $X2=4.08 $Y2=0
r82 28 32 250.524 $w=1.68e-07 $l=3.84e-06 $layer=LI1_cond $X=0.24 $Y=0 $X2=4.08
+ $Y2=0
r83 28 29 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=0.24 $Y=0
+ $X2=0.24 $Y2=0
r84 25 33 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=4.08
+ $Y2=0
r85 25 29 0.802756 $w=4.9e-07 $l=2.88e-06 $layer=MET1_cond $X=3.12 $Y=0 $X2=0.24
+ $Y2=0
r86 23 32 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=4.085 $Y=0 $X2=4.08
+ $Y2=0
r87 23 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.085 $Y=0 $X2=4.25
+ $Y2=0
r88 22 36 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=4.415 $Y=0 $X2=4.56
+ $Y2=0
r89 22 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.415 $Y=0 $X2=4.25
+ $Y2=0
r90 18 47 3.00555 $w=3.3e-07 $l=1.07912e-07 $layer=LI1_cond $X=5.97 $Y=0.085
+ $X2=6.022 $Y2=0
r91 18 20 16.4136 $w=3.28e-07 $l=4.7e-07 $layer=LI1_cond $X=5.97 $Y=0.085
+ $X2=5.97 $Y2=0.555
r92 14 44 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.11 $Y=0.085
+ $X2=5.11 $Y2=0
r93 14 16 17.4613 $w=3.28e-07 $l=5e-07 $layer=LI1_cond $X=5.11 $Y=0.085 $X2=5.11
+ $Y2=0.585
r94 10 24 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.25 $Y=0.085
+ $X2=4.25 $Y2=0
r95 10 12 17.4613 $w=3.28e-07 $l=5e-07 $layer=LI1_cond $X=4.25 $Y=0.085 $X2=4.25
+ $Y2=0.585
r96 3 20 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=5.83
+ $Y=0.41 $X2=5.97 $Y2=0.555
r97 2 16 182 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_NDIFF $count=1 $X=4.97
+ $Y=0.41 $X2=5.11 $Y2=0.585
r98 1 12 182 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_NDIFF $count=1 $X=4.115
+ $Y=0.41 $X2=4.25 $Y2=0.585
.ends

