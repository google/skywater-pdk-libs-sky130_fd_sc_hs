* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hs__and2_4 A B VGND VNB VPB VPWR X
M1000 a_83_269# B VPWR VPB pshort w=840000u l=150000u
+  ad=5.25e+11p pd=4.61e+06u as=1.58705e+12p ps=1.328e+07u
M1001 a_83_269# A VPWR VPB pshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1002 VGND a_83_269# X VNB nlowvt w=740000u l=150000u
+  ad=8.594e+11p pd=8.14e+06u as=5.254e+11p ps=4.38e+06u
M1003 VPWR a_83_269# X VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=6.944e+11p ps=5.72e+06u
M1004 X a_83_269# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_83_269# A a_504_119# VNB nlowvt w=640000u l=150000u
+  ad=2.08e+11p pd=1.93e+06u as=3.872e+11p ps=3.77e+06u
M1006 VPWR B a_83_269# VPB pshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VPWR A a_83_269# VPB pshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VGND a_83_269# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_504_119# B VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_504_119# A a_83_269# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VGND B a_504_119# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VPWR a_83_269# X VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 X a_83_269# VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 X a_83_269# VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 X a_83_269# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
