* File: sky130_fd_sc_hs__a2111oi_4.pex.spice
* Created: Thu Aug 27 20:23:07 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HS__A2111OI_4%D1 1 3 4 6 7 9 10 12 13 15 16 18 19 20 21
+ 36 37
c70 16 0 4.80185e-20 $X=1.845 $Y=1.765
r71 37 38 1.69321 $w=4.27e-07 $l=1.5e-08 $layer=POLY_cond $X=1.83 $Y=1.492
+ $X2=1.845 $Y2=1.492
r72 35 37 10.1593 $w=4.27e-07 $l=9e-08 $layer=POLY_cond $X=1.74 $Y=1.492
+ $X2=1.83 $Y2=1.492
r73 35 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.74
+ $Y=1.385 $X2=1.74 $Y2=1.385
r74 32 35 38.3794 $w=4.27e-07 $l=3.4e-07 $layer=POLY_cond $X=1.4 $Y=1.492
+ $X2=1.74 $Y2=1.492
r75 32 33 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.4
+ $Y=1.385 $X2=1.4 $Y2=1.385
r76 30 32 0.564403 $w=4.27e-07 $l=5e-09 $layer=POLY_cond $X=1.395 $Y=1.492
+ $X2=1.4 $Y2=1.492
r77 29 30 50.7963 $w=4.27e-07 $l=4.5e-07 $layer=POLY_cond $X=0.945 $Y=1.492
+ $X2=1.395 $Y2=1.492
r78 27 29 25.3981 $w=4.27e-07 $l=2.25e-07 $layer=POLY_cond $X=0.72 $Y=1.492
+ $X2=0.945 $Y2=1.492
r79 25 27 25.3981 $w=4.27e-07 $l=2.25e-07 $layer=POLY_cond $X=0.495 $Y=1.492
+ $X2=0.72 $Y2=1.492
r80 21 36 1.86883 $w=3.68e-07 $l=6e-08 $layer=LI1_cond $X=1.68 $Y=1.365 $X2=1.74
+ $Y2=1.365
r81 21 33 8.72119 $w=3.68e-07 $l=2.8e-07 $layer=LI1_cond $X=1.68 $Y=1.365
+ $X2=1.4 $Y2=1.365
r82 20 33 6.22942 $w=3.68e-07 $l=2e-07 $layer=LI1_cond $X=1.2 $Y=1.365 $X2=1.4
+ $Y2=1.365
r83 19 20 14.9506 $w=3.68e-07 $l=4.8e-07 $layer=LI1_cond $X=0.72 $Y=1.365
+ $X2=1.2 $Y2=1.365
r84 19 27 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=0.72
+ $Y=1.385 $X2=0.72 $Y2=1.385
r85 16 38 27.4666 $w=1.5e-07 $l=2.73e-07 $layer=POLY_cond $X=1.845 $Y=1.765
+ $X2=1.845 $Y2=1.492
r86 16 18 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.845 $Y=1.765
+ $X2=1.845 $Y2=2.4
r87 13 37 27.4666 $w=1.5e-07 $l=2.72e-07 $layer=POLY_cond $X=1.83 $Y=1.22
+ $X2=1.83 $Y2=1.492
r88 13 15 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.83 $Y=1.22 $X2=1.83
+ $Y2=0.74
r89 10 32 27.4666 $w=1.5e-07 $l=2.72e-07 $layer=POLY_cond $X=1.4 $Y=1.22 $X2=1.4
+ $Y2=1.492
r90 10 12 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.4 $Y=1.22 $X2=1.4
+ $Y2=0.74
r91 7 30 27.4666 $w=1.5e-07 $l=2.73e-07 $layer=POLY_cond $X=1.395 $Y=1.765
+ $X2=1.395 $Y2=1.492
r92 7 9 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.395 $Y=1.765
+ $X2=1.395 $Y2=2.4
r93 4 29 27.4666 $w=1.5e-07 $l=2.73e-07 $layer=POLY_cond $X=0.945 $Y=1.765
+ $X2=0.945 $Y2=1.492
r94 4 6 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.945 $Y=1.765
+ $X2=0.945 $Y2=2.4
r95 1 25 27.4666 $w=1.5e-07 $l=2.73e-07 $layer=POLY_cond $X=0.495 $Y=1.765
+ $X2=0.495 $Y2=1.492
r96 1 3 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.495 $Y=1.765
+ $X2=0.495 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_HS__A2111OI_4%C1 3 5 7 10 12 14 15 17 18 20 21 22 34 35
c78 35 0 4.80185e-20 $X=3.42 $Y=1.515
c79 34 0 1.12785e-19 $X=3.42 $Y=1.515
c80 12 0 1.0185e-19 $X=2.745 $Y=1.765
r81 34 36 27.3174 $w=3.97e-07 $l=2.25e-07 $layer=POLY_cond $X=3.42 $Y=1.542
+ $X2=3.645 $Y2=1.542
r82 34 35 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.42
+ $Y=1.515 $X2=3.42 $Y2=1.515
r83 32 34 27.3174 $w=3.97e-07 $l=2.25e-07 $layer=POLY_cond $X=3.195 $Y=1.542
+ $X2=3.42 $Y2=1.542
r84 31 32 54.6348 $w=3.97e-07 $l=4.5e-07 $layer=POLY_cond $X=2.745 $Y=1.542
+ $X2=3.195 $Y2=1.542
r85 30 31 6.67758 $w=3.97e-07 $l=5.5e-08 $layer=POLY_cond $X=2.69 $Y=1.542
+ $X2=2.745 $Y2=1.542
r86 28 30 35.2091 $w=3.97e-07 $l=2.9e-07 $layer=POLY_cond $X=2.4 $Y=1.542
+ $X2=2.69 $Y2=1.542
r87 28 29 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.4
+ $Y=1.515 $X2=2.4 $Y2=1.515
r88 26 28 12.7481 $w=3.97e-07 $l=1.05e-07 $layer=POLY_cond $X=2.295 $Y=1.542
+ $X2=2.4 $Y2=1.542
r89 25 26 4.24937 $w=3.97e-07 $l=3.5e-08 $layer=POLY_cond $X=2.26 $Y=1.542
+ $X2=2.295 $Y2=1.542
r90 22 35 8.0403 $w=4.28e-07 $l=3e-07 $layer=LI1_cond $X=3.12 $Y=1.565 $X2=3.42
+ $Y2=1.565
r91 21 22 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=2.64 $Y=1.565
+ $X2=3.12 $Y2=1.565
r92 21 29 6.43224 $w=4.28e-07 $l=2.4e-07 $layer=LI1_cond $X=2.64 $Y=1.565
+ $X2=2.4 $Y2=1.565
r93 18 36 25.678 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=3.645 $Y=1.765
+ $X2=3.645 $Y2=1.542
r94 18 20 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.645 $Y=1.765
+ $X2=3.645 $Y2=2.4
r95 15 32 25.678 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=3.195 $Y=1.765
+ $X2=3.195 $Y2=1.542
r96 15 17 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.195 $Y=1.765
+ $X2=3.195 $Y2=2.4
r97 12 31 25.678 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=2.745 $Y=1.765
+ $X2=2.745 $Y2=1.542
r98 12 14 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.745 $Y=1.765
+ $X2=2.745 $Y2=2.4
r99 8 30 25.678 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=2.69 $Y=1.32 $X2=2.69
+ $Y2=1.542
r100 8 10 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=2.69 $Y=1.32
+ $X2=2.69 $Y2=0.74
r101 5 26 25.678 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=2.295 $Y=1.765
+ $X2=2.295 $Y2=1.542
r102 5 7 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.295 $Y=1.765
+ $X2=2.295 $Y2=2.4
r103 1 25 25.678 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=2.26 $Y=1.32
+ $X2=2.26 $Y2=1.542
r104 1 3 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=2.26 $Y=1.32 $X2=2.26
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HS__A2111OI_4%B1 3 7 9 11 12 14 15 17 18 20 21 22 23 36
+ 37
c72 37 0 1.06992e-19 $X=5.91 $Y=1.515
c73 18 0 1.42688e-20 $X=5.985 $Y=1.765
r74 36 38 10.3879 $w=3.48e-07 $l=7.5e-08 $layer=POLY_cond $X=5.91 $Y=1.557
+ $X2=5.985 $Y2=1.557
r75 36 37 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=5.91
+ $Y=1.515 $X2=5.91 $Y2=1.515
r76 34 36 51.9397 $w=3.48e-07 $l=3.75e-07 $layer=POLY_cond $X=5.535 $Y=1.557
+ $X2=5.91 $Y2=1.557
r77 33 34 62.3276 $w=3.48e-07 $l=4.5e-07 $layer=POLY_cond $X=5.085 $Y=1.557
+ $X2=5.535 $Y2=1.557
r78 32 33 62.3276 $w=3.48e-07 $l=4.5e-07 $layer=POLY_cond $X=4.635 $Y=1.557
+ $X2=5.085 $Y2=1.557
r79 31 32 25.6236 $w=3.48e-07 $l=1.85e-07 $layer=POLY_cond $X=4.45 $Y=1.557
+ $X2=4.635 $Y2=1.557
r80 29 31 1.38506 $w=3.48e-07 $l=1e-08 $layer=POLY_cond $X=4.44 $Y=1.557
+ $X2=4.45 $Y2=1.557
r81 29 30 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=4.44
+ $Y=1.515 $X2=4.44 $Y2=1.515
r82 23 37 10.4524 $w=4.28e-07 $l=3.9e-07 $layer=LI1_cond $X=5.52 $Y=1.565
+ $X2=5.91 $Y2=1.565
r83 22 23 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=5.04 $Y=1.565
+ $X2=5.52 $Y2=1.565
r84 21 22 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=4.56 $Y=1.565
+ $X2=5.04 $Y2=1.565
r85 21 30 3.21612 $w=4.28e-07 $l=1.2e-07 $layer=LI1_cond $X=4.56 $Y=1.565
+ $X2=4.44 $Y2=1.565
r86 18 38 22.4912 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=5.985 $Y=1.765
+ $X2=5.985 $Y2=1.557
r87 18 20 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=5.985 $Y=1.765
+ $X2=5.985 $Y2=2.4
r88 15 34 22.4912 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=5.535 $Y=1.765
+ $X2=5.535 $Y2=1.557
r89 15 17 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=5.535 $Y=1.765
+ $X2=5.535 $Y2=2.4
r90 12 33 22.4912 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=5.085 $Y=1.765
+ $X2=5.085 $Y2=1.557
r91 12 14 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=5.085 $Y=1.765
+ $X2=5.085 $Y2=2.4
r92 9 32 22.4912 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=4.635 $Y=1.765
+ $X2=4.635 $Y2=1.557
r93 9 11 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=4.635 $Y=1.765
+ $X2=4.635 $Y2=2.4
r94 5 31 22.4912 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.45 $Y=1.35
+ $X2=4.45 $Y2=1.557
r95 5 7 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=4.45 $Y=1.35 $X2=4.45
+ $Y2=0.74
r96 1 29 58.1724 $w=3.48e-07 $l=5.13167e-07 $layer=POLY_cond $X=4.02 $Y=1.35
+ $X2=4.44 $Y2=1.557
r97 1 3 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=4.02 $Y=1.35 $X2=4.02
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HS__A2111OI_4%A1 1 3 6 8 10 13 15 17 20 22 24 27 29 30
+ 31 47
c85 31 0 1.11272e-19 $X=7.92 $Y=1.665
c86 27 0 1.20142e-20 $X=7.79 $Y=0.74
c87 22 0 1.16815e-20 $X=7.785 $Y=1.765
c88 1 0 1.06992e-19 $X=6.435 $Y=1.765
r89 47 48 0.651351 $w=3.7e-07 $l=5e-09 $layer=POLY_cond $X=7.785 $Y=1.557
+ $X2=7.79 $Y2=1.557
r90 45 47 9.77027 $w=3.7e-07 $l=7.5e-08 $layer=POLY_cond $X=7.71 $Y=1.557
+ $X2=7.785 $Y2=1.557
r91 45 46 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=7.71
+ $Y=1.515 $X2=7.71 $Y2=1.515
r92 43 45 45.5946 $w=3.7e-07 $l=3.5e-07 $layer=POLY_cond $X=7.36 $Y=1.557
+ $X2=7.71 $Y2=1.557
r93 42 43 3.25676 $w=3.7e-07 $l=2.5e-08 $layer=POLY_cond $X=7.335 $Y=1.557
+ $X2=7.36 $Y2=1.557
r94 41 42 52.7595 $w=3.7e-07 $l=4.05e-07 $layer=POLY_cond $X=6.93 $Y=1.557
+ $X2=7.335 $Y2=1.557
r95 40 41 5.86216 $w=3.7e-07 $l=4.5e-08 $layer=POLY_cond $X=6.885 $Y=1.557
+ $X2=6.93 $Y2=1.557
r96 38 40 25.4027 $w=3.7e-07 $l=1.95e-07 $layer=POLY_cond $X=6.69 $Y=1.557
+ $X2=6.885 $Y2=1.557
r97 38 39 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.69
+ $Y=1.515 $X2=6.69 $Y2=1.515
r98 36 38 24.7514 $w=3.7e-07 $l=1.9e-07 $layer=POLY_cond $X=6.5 $Y=1.557
+ $X2=6.69 $Y2=1.557
r99 35 36 8.46757 $w=3.7e-07 $l=6.5e-08 $layer=POLY_cond $X=6.435 $Y=1.557
+ $X2=6.5 $Y2=1.557
r100 31 46 5.62821 $w=4.28e-07 $l=2.1e-07 $layer=LI1_cond $X=7.92 $Y=1.565
+ $X2=7.71 $Y2=1.565
r101 30 46 7.23627 $w=4.28e-07 $l=2.7e-07 $layer=LI1_cond $X=7.44 $Y=1.565
+ $X2=7.71 $Y2=1.565
r102 29 30 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=6.96 $Y=1.565
+ $X2=7.44 $Y2=1.565
r103 29 39 7.23627 $w=4.28e-07 $l=2.7e-07 $layer=LI1_cond $X=6.96 $Y=1.565
+ $X2=6.69 $Y2=1.565
r104 25 48 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=7.79 $Y=1.35
+ $X2=7.79 $Y2=1.557
r105 25 27 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=7.79 $Y=1.35
+ $X2=7.79 $Y2=0.74
r106 22 47 23.9667 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=7.785 $Y=1.765
+ $X2=7.785 $Y2=1.557
r107 22 24 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=7.785 $Y=1.765
+ $X2=7.785 $Y2=2.4
r108 18 43 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=7.36 $Y=1.35
+ $X2=7.36 $Y2=1.557
r109 18 20 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=7.36 $Y=1.35
+ $X2=7.36 $Y2=0.74
r110 15 42 23.9667 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=7.335 $Y=1.765
+ $X2=7.335 $Y2=1.557
r111 15 17 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=7.335 $Y=1.765
+ $X2=7.335 $Y2=2.4
r112 11 41 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=6.93 $Y=1.35
+ $X2=6.93 $Y2=1.557
r113 11 13 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=6.93 $Y=1.35
+ $X2=6.93 $Y2=0.74
r114 8 40 23.9667 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=6.885 $Y=1.765
+ $X2=6.885 $Y2=1.557
r115 8 10 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=6.885 $Y=1.765
+ $X2=6.885 $Y2=2.4
r116 4 36 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=6.5 $Y=1.35 $X2=6.5
+ $Y2=1.557
r117 4 6 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=6.5 $Y=1.35 $X2=6.5
+ $Y2=0.74
r118 1 35 23.9667 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=6.435 $Y=1.765
+ $X2=6.435 $Y2=1.557
r119 1 3 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=6.435 $Y=1.765
+ $X2=6.435 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_HS__A2111OI_4%A2 3 5 7 10 12 14 17 19 21 24 26 28 29 30
+ 31 46 47
c76 46 0 1.16815e-20 $X=9.39 $Y=1.515
c77 5 0 9.70031e-20 $X=8.235 $Y=1.765
c78 3 0 2.06049e-19 $X=8.22 $Y=0.74
r79 47 48 9.77027 $w=3.7e-07 $l=7.5e-08 $layer=POLY_cond $X=9.51 $Y=1.557
+ $X2=9.585 $Y2=1.557
r80 45 47 15.6324 $w=3.7e-07 $l=1.2e-07 $layer=POLY_cond $X=9.39 $Y=1.557
+ $X2=9.51 $Y2=1.557
r81 45 46 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=9.39
+ $Y=1.515 $X2=9.39 $Y2=1.515
r82 43 45 33.2189 $w=3.7e-07 $l=2.55e-07 $layer=POLY_cond $X=9.135 $Y=1.557
+ $X2=9.39 $Y2=1.557
r83 42 43 7.16487 $w=3.7e-07 $l=5.5e-08 $layer=POLY_cond $X=9.08 $Y=1.557
+ $X2=9.135 $Y2=1.557
r84 41 42 51.4568 $w=3.7e-07 $l=3.95e-07 $layer=POLY_cond $X=8.685 $Y=1.557
+ $X2=9.08 $Y2=1.557
r85 40 41 4.55946 $w=3.7e-07 $l=3.5e-08 $layer=POLY_cond $X=8.65 $Y=1.557
+ $X2=8.685 $Y2=1.557
r86 38 40 36.4757 $w=3.7e-07 $l=2.8e-07 $layer=POLY_cond $X=8.37 $Y=1.557
+ $X2=8.65 $Y2=1.557
r87 38 39 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=8.37
+ $Y=1.515 $X2=8.37 $Y2=1.515
r88 36 38 17.5865 $w=3.7e-07 $l=1.35e-07 $layer=POLY_cond $X=8.235 $Y=1.557
+ $X2=8.37 $Y2=1.557
r89 35 36 1.95405 $w=3.7e-07 $l=1.5e-08 $layer=POLY_cond $X=8.22 $Y=1.557
+ $X2=8.235 $Y2=1.557
r90 31 46 0.80403 $w=4.28e-07 $l=3e-08 $layer=LI1_cond $X=9.36 $Y=1.565 $X2=9.39
+ $Y2=1.565
r91 30 31 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=8.88 $Y=1.565
+ $X2=9.36 $Y2=1.565
r92 29 30 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=8.4 $Y=1.565
+ $X2=8.88 $Y2=1.565
r93 29 39 0.80403 $w=4.28e-07 $l=3e-08 $layer=LI1_cond $X=8.4 $Y=1.565 $X2=8.37
+ $Y2=1.565
r94 26 48 23.9667 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=9.585 $Y=1.765
+ $X2=9.585 $Y2=1.557
r95 26 28 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=9.585 $Y=1.765
+ $X2=9.585 $Y2=2.4
r96 22 47 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=9.51 $Y=1.35
+ $X2=9.51 $Y2=1.557
r97 22 24 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=9.51 $Y=1.35
+ $X2=9.51 $Y2=0.74
r98 19 43 23.9667 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=9.135 $Y=1.765
+ $X2=9.135 $Y2=1.557
r99 19 21 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=9.135 $Y=1.765
+ $X2=9.135 $Y2=2.4
r100 15 42 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=9.08 $Y=1.35
+ $X2=9.08 $Y2=1.557
r101 15 17 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=9.08 $Y=1.35
+ $X2=9.08 $Y2=0.74
r102 12 41 23.9667 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=8.685 $Y=1.765
+ $X2=8.685 $Y2=1.557
r103 12 14 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=8.685 $Y=1.765
+ $X2=8.685 $Y2=2.4
r104 8 40 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=8.65 $Y=1.35
+ $X2=8.65 $Y2=1.557
r105 8 10 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=8.65 $Y=1.35
+ $X2=8.65 $Y2=0.74
r106 5 36 23.9667 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=8.235 $Y=1.765
+ $X2=8.235 $Y2=1.557
r107 5 7 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=8.235 $Y=1.765
+ $X2=8.235 $Y2=2.4
r108 1 35 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=8.22 $Y=1.35
+ $X2=8.22 $Y2=1.557
r109 1 3 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=8.22 $Y=1.35 $X2=8.22
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HS__A2111OI_4%A_29_368# 1 2 3 4 5 18 20 21 24 26 28 31
+ 32 36 38 42 46 48
c70 28 0 6.36857e-20 $X=2.07 $Y=2.12
c71 26 0 1.0185e-19 $X=1.905 $Y=2.99
r72 39 46 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=3.085 $Y=2.035
+ $X2=2.97 $Y2=2.035
r73 38 48 4.17978 $w=1.7e-07 $l=1.94808e-07 $layer=LI1_cond $X=3.705 $Y=2.035
+ $X2=3.87 $Y2=1.97
r74 38 39 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=3.705 $Y=2.035
+ $X2=3.085 $Y2=2.035
r75 34 46 0.280307 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.97 $Y=2.12
+ $X2=2.97 $Y2=2.035
r76 34 36 22.5478 $w=2.28e-07 $l=4.5e-07 $layer=LI1_cond $X=2.97 $Y=2.12
+ $X2=2.97 $Y2=2.57
r77 33 44 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.235 $Y=2.035
+ $X2=2.07 $Y2=2.035
r78 32 46 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=2.855 $Y=2.035
+ $X2=2.97 $Y2=2.035
r79 32 33 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=2.855 $Y=2.035
+ $X2=2.235 $Y2=2.035
r80 29 31 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=2.07 $Y=2.905 $X2=2.07
+ $Y2=2.815
r81 28 44 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.07 $Y=2.12 $X2=2.07
+ $Y2=2.035
r82 28 31 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=2.07 $Y=2.12
+ $X2=2.07 $Y2=2.815
r83 27 42 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.255 $Y=2.99
+ $X2=1.17 $Y2=2.99
r84 26 29 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.905 $Y=2.99
+ $X2=2.07 $Y2=2.905
r85 26 27 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=1.905 $Y=2.99
+ $X2=1.255 $Y2=2.99
r86 22 42 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.17 $Y=2.905
+ $X2=1.17 $Y2=2.99
r87 22 24 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.17 $Y=2.905
+ $X2=1.17 $Y2=2.225
r88 20 42 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.085 $Y=2.99
+ $X2=1.17 $Y2=2.99
r89 20 21 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=1.085 $Y=2.99
+ $X2=0.355 $Y2=2.99
r90 16 21 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.23 $Y=2.905
+ $X2=0.355 $Y2=2.99
r91 16 18 31.3464 $w=2.48e-07 $l=6.8e-07 $layer=LI1_cond $X=0.23 $Y=2.905
+ $X2=0.23 $Y2=2.225
r92 5 48 300 $w=1.7e-07 $l=2.74955e-07 $layer=licon1_PDIFF $count=2 $X=3.72
+ $Y=1.84 $X2=3.87 $Y2=2.05
r93 4 46 600 $w=1.7e-07 $l=2.59374e-07 $layer=licon1_PDIFF $count=1 $X=2.82
+ $Y=1.84 $X2=2.97 $Y2=2.035
r94 4 36 600 $w=1.7e-07 $l=8.01499e-07 $layer=licon1_PDIFF $count=1 $X=2.82
+ $Y=1.84 $X2=2.97 $Y2=2.57
r95 3 44 400 $w=1.7e-07 $l=2.59374e-07 $layer=licon1_PDIFF $count=1 $X=1.92
+ $Y=1.84 $X2=2.07 $Y2=2.035
r96 3 31 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=1.92
+ $Y=1.84 $X2=2.07 $Y2=2.815
r97 2 24 300 $w=1.7e-07 $l=4.53845e-07 $layer=licon1_PDIFF $count=2 $X=1.02
+ $Y=1.84 $X2=1.17 $Y2=2.225
r98 1 18 300 $w=1.7e-07 $l=4.43114e-07 $layer=licon1_PDIFF $count=2 $X=0.145
+ $Y=1.84 $X2=0.27 $Y2=2.225
.ends

.subckt PM_SKY130_FD_SC_HS__A2111OI_4%Y 1 2 3 4 5 6 7 22 23 24 28 30 34 38 40 44
+ 46 50 54 57 59 61 64 67 68 70 74 75 79 84
c133 70 0 4.44094e-20 $X=7.575 $Y=0.95
c134 54 0 1.20142e-20 $X=7.41 $Y=1.022
c135 40 0 4.90994e-20 $X=2.39 $Y=0.925
r136 79 84 2.75584 $w=2.28e-07 $l=5.5e-08 $layer=LI1_cond $X=0.24 $Y=1.72
+ $X2=0.24 $Y2=1.665
r137 75 79 2.9826 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.24 $Y=1.805
+ $X2=0.24 $Y2=1.72
r138 75 84 0.751593 $w=2.28e-07 $l=1.5e-08 $layer=LI1_cond $X=0.24 $Y=1.65
+ $X2=0.24 $Y2=1.665
r139 74 75 17.7877 $w=2.28e-07 $l=3.55e-07 $layer=LI1_cond $X=0.24 $Y=1.295
+ $X2=0.24 $Y2=1.65
r140 70 72 2.51442 $w=3.28e-07 $l=7.2e-08 $layer=LI1_cond $X=7.575 $Y=0.95
+ $X2=7.575 $Y2=1.022
r141 66 68 7.23236 $w=4.08e-07 $l=1.65e-07 $layer=LI1_cond $X=6.715 $Y=0.975
+ $X2=6.88 $Y2=0.975
r142 66 67 7.51706 $w=4.08e-07 $l=1.65e-07 $layer=LI1_cond $X=6.715 $Y=0.975
+ $X2=6.55 $Y2=0.975
r143 61 62 7.83661 $w=2.48e-07 $l=1.7e-07 $layer=LI1_cond $X=2.515 $Y=0.925
+ $X2=2.515 $Y2=1.095
r144 56 74 14.2803 $w=2.28e-07 $l=2.85e-07 $layer=LI1_cond $X=0.24 $Y=1.01
+ $X2=0.24 $Y2=1.295
r145 54 72 3.26307 $w=2.15e-07 $l=1.65e-07 $layer=LI1_cond $X=7.41 $Y=1.022
+ $X2=7.575 $Y2=1.022
r146 54 68 28.4091 $w=2.13e-07 $l=5.3e-07 $layer=LI1_cond $X=7.41 $Y=1.022
+ $X2=6.88 $Y2=1.022
r147 53 64 6.51676 $w=1.87e-07 $l=1.25e-07 $layer=LI1_cond $X=4.32 $Y=1.077
+ $X2=4.195 $Y2=1.077
r148 53 67 120.647 $w=2.03e-07 $l=2.23e-06 $layer=LI1_cond $X=4.32 $Y=1.077
+ $X2=6.55 $Y2=1.077
r149 48 64 0.330231 $w=2.5e-07 $l=1.02e-07 $layer=LI1_cond $X=4.195 $Y=0.975
+ $X2=4.195 $Y2=1.077
r150 48 50 21.205 $w=2.48e-07 $l=4.6e-07 $layer=LI1_cond $X=4.195 $Y=0.975
+ $X2=4.195 $Y2=0.515
r151 47 62 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.64 $Y=1.095
+ $X2=2.515 $Y2=1.095
r152 46 64 6.51676 $w=1.87e-07 $l=1.33697e-07 $layer=LI1_cond $X=4.07 $Y=1.095
+ $X2=4.195 $Y2=1.077
r153 46 47 93.2941 $w=1.68e-07 $l=1.43e-06 $layer=LI1_cond $X=4.07 $Y=1.095
+ $X2=2.64 $Y2=1.095
r154 42 61 3.91831 $w=2.48e-07 $l=8.5e-08 $layer=LI1_cond $X=2.515 $Y=0.84
+ $X2=2.515 $Y2=0.925
r155 42 44 14.9818 $w=2.48e-07 $l=3.25e-07 $layer=LI1_cond $X=2.515 $Y=0.84
+ $X2=2.515 $Y2=0.515
r156 41 59 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.7 $Y=0.925
+ $X2=1.615 $Y2=0.925
r157 40 61 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.39 $Y=0.925
+ $X2=2.515 $Y2=0.925
r158 40 41 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=2.39 $Y=0.925
+ $X2=1.7 $Y2=0.925
r159 36 59 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.615 $Y=0.84
+ $X2=1.615 $Y2=0.925
r160 36 38 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.615 $Y=0.84
+ $X2=1.615 $Y2=0.495
r161 32 34 4.37928 $w=2.48e-07 $l=9.5e-08 $layer=LI1_cond $X=1.58 $Y=1.89
+ $X2=1.58 $Y2=1.985
r162 31 57 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.885 $Y=1.805
+ $X2=0.72 $Y2=1.805
r163 30 32 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.455 $Y=1.805
+ $X2=1.58 $Y2=1.89
r164 30 31 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=1.455 $Y=1.805
+ $X2=0.885 $Y2=1.805
r165 26 57 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.72 $Y=1.89
+ $X2=0.72 $Y2=1.805
r166 26 28 3.31764 $w=3.28e-07 $l=9.5e-08 $layer=LI1_cond $X=0.72 $Y=1.89
+ $X2=0.72 $Y2=1.985
r167 25 75 4.03528 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=0.355 $Y=1.805
+ $X2=0.24 $Y2=1.805
r168 24 57 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.555 $Y=1.805
+ $X2=0.72 $Y2=1.805
r169 24 25 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=0.555 $Y=1.805
+ $X2=0.355 $Y2=1.805
r170 23 56 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=0.355 $Y=0.925
+ $X2=0.24 $Y2=1.01
r171 22 59 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.53 $Y=0.925
+ $X2=1.615 $Y2=0.925
r172 22 23 76.6578 $w=1.68e-07 $l=1.175e-06 $layer=LI1_cond $X=1.53 $Y=0.925
+ $X2=0.355 $Y2=0.925
r173 7 34 300 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=2 $X=1.47
+ $Y=1.84 $X2=1.62 $Y2=1.985
r174 6 28 300 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=2 $X=0.57
+ $Y=1.84 $X2=0.72 $Y2=1.985
r175 5 70 182 $w=1.7e-07 $l=6.4622e-07 $layer=licon1_NDIFF $count=1 $X=7.435
+ $Y=0.37 $X2=7.575 $Y2=0.95
r176 4 66 182 $w=1.7e-07 $l=6.4622e-07 $layer=licon1_NDIFF $count=1 $X=6.575
+ $Y=0.37 $X2=6.715 $Y2=0.95
r177 3 50 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=4.095
+ $Y=0.37 $X2=4.235 $Y2=0.515
r178 2 61 182 $w=1.7e-07 $l=6.61306e-07 $layer=licon1_NDIFF $count=1 $X=2.335
+ $Y=0.37 $X2=2.475 $Y2=0.965
r179 2 44 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=2.335
+ $Y=0.37 $X2=2.475 $Y2=0.515
r180 1 59 182 $w=1.7e-07 $l=6.21068e-07 $layer=licon1_NDIFF $count=1 $X=1.475
+ $Y=0.37 $X2=1.615 $Y2=0.925
r181 1 38 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=1.475
+ $Y=0.37 $X2=1.615 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_HS__A2111OI_4%A_474_368# 1 2 3 4 15 17 18 21 23 27 29 33
+ 35 36
r64 31 33 17.4613 $w=3.28e-07 $l=5e-07 $layer=LI1_cond $X=5.76 $Y=2.905 $X2=5.76
+ $Y2=2.405
r65 30 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.025 $Y=2.99
+ $X2=4.86 $Y2=2.99
r66 29 31 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=5.595 $Y=2.99
+ $X2=5.76 $Y2=2.905
r67 29 30 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=5.595 $Y=2.99
+ $X2=5.025 $Y2=2.99
r68 25 36 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.86 $Y=2.905
+ $X2=4.86 $Y2=2.99
r69 25 27 17.4613 $w=3.28e-07 $l=5e-07 $layer=LI1_cond $X=4.86 $Y=2.905 $X2=4.86
+ $Y2=2.405
r70 24 35 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.585 $Y=2.99
+ $X2=3.42 $Y2=2.99
r71 23 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.695 $Y=2.99
+ $X2=4.86 $Y2=2.99
r72 23 24 72.4171 $w=1.68e-07 $l=1.11e-06 $layer=LI1_cond $X=4.695 $Y=2.99
+ $X2=3.585 $Y2=2.99
r73 19 35 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.42 $Y=2.905
+ $X2=3.42 $Y2=2.99
r74 19 21 16.9374 $w=3.28e-07 $l=4.85e-07 $layer=LI1_cond $X=3.42 $Y=2.905
+ $X2=3.42 $Y2=2.42
r75 17 35 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.255 $Y=2.99
+ $X2=3.42 $Y2=2.99
r76 17 18 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=3.255 $Y=2.99
+ $X2=2.685 $Y2=2.99
r77 13 18 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=2.56 $Y=2.905
+ $X2=2.685 $Y2=2.99
r78 13 15 20.744 $w=2.48e-07 $l=4.5e-07 $layer=LI1_cond $X=2.56 $Y=2.905
+ $X2=2.56 $Y2=2.455
r79 4 33 300 $w=1.7e-07 $l=6.3559e-07 $layer=licon1_PDIFF $count=2 $X=5.61
+ $Y=1.84 $X2=5.76 $Y2=2.405
r80 3 27 300 $w=1.7e-07 $l=6.3559e-07 $layer=licon1_PDIFF $count=2 $X=4.71
+ $Y=1.84 $X2=4.86 $Y2=2.405
r81 2 21 300 $w=1.7e-07 $l=6.50692e-07 $layer=licon1_PDIFF $count=2 $X=3.27
+ $Y=1.84 $X2=3.42 $Y2=2.42
r82 1 15 300 $w=1.7e-07 $l=6.85912e-07 $layer=licon1_PDIFF $count=2 $X=2.37
+ $Y=1.84 $X2=2.52 $Y2=2.455
.ends

.subckt PM_SKY130_FD_SC_HS__A2111OI_4%A_853_368# 1 2 3 4 5 6 7 22 24 26 30 32 36
+ 38 42 44 48 50 54 56 58 60 65 69 71 73
r94 58 75 3.1514 $w=2.5e-07 $l=1.5e-07 $layer=LI1_cond $X=9.85 $Y=2.12 $X2=9.85
+ $Y2=1.97
r95 58 60 12.9074 $w=2.48e-07 $l=2.8e-07 $layer=LI1_cond $X=9.85 $Y=2.12
+ $X2=9.85 $Y2=2.4
r96 57 73 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.075 $Y=2.035
+ $X2=8.91 $Y2=2.035
r97 56 75 3.99177 $w=1.7e-07 $l=1.5411e-07 $layer=LI1_cond $X=9.725 $Y=2.035
+ $X2=9.85 $Y2=1.97
r98 56 57 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=9.725 $Y=2.035
+ $X2=9.075 $Y2=2.035
r99 52 73 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.91 $Y=2.12 $X2=8.91
+ $Y2=2.035
r100 52 54 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=8.91 $Y=2.12
+ $X2=8.91 $Y2=2.815
r101 51 71 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.095 $Y=2.035
+ $X2=8.01 $Y2=2.035
r102 50 73 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.745 $Y=2.035
+ $X2=8.91 $Y2=2.035
r103 50 51 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=8.745 $Y=2.035
+ $X2=8.095 $Y2=2.035
r104 46 71 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.01 $Y=2.12
+ $X2=8.01 $Y2=2.035
r105 46 48 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=8.01 $Y=2.12
+ $X2=8.01 $Y2=2.43
r106 45 69 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.195 $Y=2.035
+ $X2=7.11 $Y2=2.035
r107 44 71 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.925 $Y=2.035
+ $X2=8.01 $Y2=2.035
r108 44 45 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=7.925 $Y=2.035
+ $X2=7.195 $Y2=2.035
r109 40 69 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.11 $Y=2.12
+ $X2=7.11 $Y2=2.035
r110 40 42 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=7.11 $Y=2.12
+ $X2=7.11 $Y2=2.43
r111 39 67 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.295 $Y=2.035
+ $X2=6.21 $Y2=2.035
r112 38 69 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.025 $Y=2.035
+ $X2=7.11 $Y2=2.035
r113 38 39 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=7.025 $Y=2.035
+ $X2=6.295 $Y2=2.035
r114 34 67 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.21 $Y=2.12
+ $X2=6.21 $Y2=2.035
r115 34 36 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=6.21 $Y=2.12
+ $X2=6.21 $Y2=2.43
r116 33 65 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=5.425 $Y=2.035
+ $X2=5.31 $Y2=2.035
r117 32 67 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.125 $Y=2.035
+ $X2=6.21 $Y2=2.035
r118 32 33 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=6.125 $Y=2.035
+ $X2=5.425 $Y2=2.035
r119 28 65 0.280307 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.31 $Y=2.12
+ $X2=5.31 $Y2=2.035
r120 28 30 22.5478 $w=2.28e-07 $l=4.5e-07 $layer=LI1_cond $X=5.31 $Y=2.12
+ $X2=5.31 $Y2=2.57
r121 27 63 4.57959 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=4.525 $Y=2.035
+ $X2=4.385 $Y2=2.035
r122 26 65 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=5.195 $Y=2.035
+ $X2=5.31 $Y2=2.035
r123 26 27 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.195 $Y=2.035
+ $X2=4.525 $Y2=2.035
r124 22 63 2.78046 $w=2.8e-07 $l=8.5e-08 $layer=LI1_cond $X=4.385 $Y=2.12
+ $X2=4.385 $Y2=2.035
r125 22 24 18.5214 $w=2.78e-07 $l=4.5e-07 $layer=LI1_cond $X=4.385 $Y=2.12
+ $X2=4.385 $Y2=2.57
r126 7 75 600 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=9.66
+ $Y=1.84 $X2=9.81 $Y2=1.985
r127 7 60 300 $w=1.7e-07 $l=6.30555e-07 $layer=licon1_PDIFF $count=2 $X=9.66
+ $Y=1.84 $X2=9.81 $Y2=2.4
r128 6 73 400 $w=1.7e-07 $l=2.59374e-07 $layer=licon1_PDIFF $count=1 $X=8.76
+ $Y=1.84 $X2=8.91 $Y2=2.035
r129 6 54 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=8.76
+ $Y=1.84 $X2=8.91 $Y2=2.815
r130 5 71 600 $w=1.7e-07 $l=2.59374e-07 $layer=licon1_PDIFF $count=1 $X=7.86
+ $Y=1.84 $X2=8.01 $Y2=2.035
r131 5 48 300 $w=1.7e-07 $l=6.60757e-07 $layer=licon1_PDIFF $count=2 $X=7.86
+ $Y=1.84 $X2=8.01 $Y2=2.43
r132 4 69 600 $w=1.7e-07 $l=2.59374e-07 $layer=licon1_PDIFF $count=1 $X=6.96
+ $Y=1.84 $X2=7.11 $Y2=2.035
r133 4 42 300 $w=1.7e-07 $l=6.60757e-07 $layer=licon1_PDIFF $count=2 $X=6.96
+ $Y=1.84 $X2=7.11 $Y2=2.43
r134 3 67 600 $w=1.7e-07 $l=2.59374e-07 $layer=licon1_PDIFF $count=1 $X=6.06
+ $Y=1.84 $X2=6.21 $Y2=2.035
r135 3 36 300 $w=1.7e-07 $l=6.60757e-07 $layer=licon1_PDIFF $count=2 $X=6.06
+ $Y=1.84 $X2=6.21 $Y2=2.43
r136 2 65 600 $w=1.7e-07 $l=2.59374e-07 $layer=licon1_PDIFF $count=1 $X=5.16
+ $Y=1.84 $X2=5.31 $Y2=2.035
r137 2 30 600 $w=1.7e-07 $l=8.01499e-07 $layer=licon1_PDIFF $count=1 $X=5.16
+ $Y=1.84 $X2=5.31 $Y2=2.57
r138 1 63 600 $w=1.7e-07 $l=2.57488e-07 $layer=licon1_PDIFF $count=1 $X=4.265
+ $Y=1.84 $X2=4.41 $Y2=2.035
r139 1 24 600 $w=1.7e-07 $l=7.99218e-07 $layer=licon1_PDIFF $count=1 $X=4.265
+ $Y=1.84 $X2=4.41 $Y2=2.57
.ends

.subckt PM_SKY130_FD_SC_HS__A2111OI_4%VPWR 1 2 3 4 15 17 21 25 29 31 32 33 42 47
+ 54 55 58 61 64
r115 64 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.36 $Y=3.33
+ $X2=9.36 $Y2=3.33
r116 61 62 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=3.33 $X2=8.4
+ $Y2=3.33
r117 58 59 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r118 55 65 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.84 $Y=3.33
+ $X2=9.36 $Y2=3.33
r119 54 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.84 $Y=3.33
+ $X2=9.84 $Y2=3.33
r120 52 64 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=9.525 $Y=3.33
+ $X2=9.4 $Y2=3.33
r121 52 54 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=9.525 $Y=3.33
+ $X2=9.84 $Y2=3.33
r122 51 65 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=3.33
+ $X2=9.36 $Y2=3.33
r123 51 62 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=3.33
+ $X2=8.4 $Y2=3.33
r124 50 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r125 48 61 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.545 $Y=3.33
+ $X2=8.42 $Y2=3.33
r126 48 50 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=8.545 $Y=3.33
+ $X2=8.88 $Y2=3.33
r127 47 64 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=9.275 $Y=3.33
+ $X2=9.4 $Y2=3.33
r128 47 50 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=9.275 $Y=3.33
+ $X2=8.88 $Y2=3.33
r129 46 62 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=3.33
+ $X2=8.4 $Y2=3.33
r130 46 59 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=3.33
+ $X2=7.44 $Y2=3.33
r131 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r132 43 58 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.725 $Y=3.33
+ $X2=7.56 $Y2=3.33
r133 43 45 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=7.725 $Y=3.33
+ $X2=7.92 $Y2=3.33
r134 42 61 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.295 $Y=3.33
+ $X2=8.42 $Y2=3.33
r135 42 45 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=8.295 $Y=3.33
+ $X2=7.92 $Y2=3.33
r136 41 59 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=7.44 $Y2=3.33
r137 40 41 1.32857 $w=1.7e-07 $l=1.19e-06 $layer=mcon $count=7 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r138 36 40 407.102 $w=1.68e-07 $l=6.24e-06 $layer=LI1_cond $X=0.24 $Y=3.33
+ $X2=6.48 $Y2=3.33
r139 36 37 1.32857 $w=1.7e-07 $l=1.19e-06 $layer=mcon $count=7 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r140 33 41 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=6.48 $Y2=3.33
r141 33 37 1.33793 $w=4.9e-07 $l=4.8e-06 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=0.24 $Y2=3.33
r142 31 40 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=6.495 $Y=3.33
+ $X2=6.48 $Y2=3.33
r143 31 32 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.495 $Y=3.33
+ $X2=6.66 $Y2=3.33
r144 27 64 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=9.4 $Y=3.245
+ $X2=9.4 $Y2=3.33
r145 27 29 36.4172 $w=2.48e-07 $l=7.9e-07 $layer=LI1_cond $X=9.4 $Y=3.245
+ $X2=9.4 $Y2=2.455
r146 23 61 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=8.42 $Y=3.245
+ $X2=8.42 $Y2=3.33
r147 23 25 36.4172 $w=2.48e-07 $l=7.9e-07 $layer=LI1_cond $X=8.42 $Y=3.245
+ $X2=8.42 $Y2=2.455
r148 19 58 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.56 $Y=3.245
+ $X2=7.56 $Y2=3.33
r149 19 21 30.3826 $w=3.28e-07 $l=8.7e-07 $layer=LI1_cond $X=7.56 $Y=3.245
+ $X2=7.56 $Y2=2.375
r150 18 32 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.825 $Y=3.33
+ $X2=6.66 $Y2=3.33
r151 17 58 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.395 $Y=3.33
+ $X2=7.56 $Y2=3.33
r152 17 18 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=7.395 $Y=3.33
+ $X2=6.825 $Y2=3.33
r153 13 32 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.66 $Y=3.245
+ $X2=6.66 $Y2=3.33
r154 13 15 30.3826 $w=3.28e-07 $l=8.7e-07 $layer=LI1_cond $X=6.66 $Y=3.245
+ $X2=6.66 $Y2=2.375
r155 4 29 300 $w=1.7e-07 $l=6.85912e-07 $layer=licon1_PDIFF $count=2 $X=9.21
+ $Y=1.84 $X2=9.36 $Y2=2.455
r156 3 25 300 $w=1.7e-07 $l=6.85912e-07 $layer=licon1_PDIFF $count=2 $X=8.31
+ $Y=1.84 $X2=8.46 $Y2=2.455
r157 2 21 300 $w=1.7e-07 $l=6.05372e-07 $layer=licon1_PDIFF $count=2 $X=7.41
+ $Y=1.84 $X2=7.56 $Y2=2.375
r158 1 15 300 $w=1.7e-07 $l=6.05372e-07 $layer=licon1_PDIFF $count=2 $X=6.51
+ $Y=1.84 $X2=6.66 $Y2=2.375
.ends

.subckt PM_SKY130_FD_SC_HS__A2111OI_4%VGND 1 2 3 4 5 6 21 25 27 31 35 39 42 43
+ 44 46 59 67 74 75 78 82 88 90 93 96
r103 96 97 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.36 $Y=0 $X2=9.36
+ $Y2=0
r104 93 94 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r105 90 91 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r106 87 88 11.4973 $w=9.23e-07 $l=9.5e-08 $layer=LI1_cond $X=3.805 $Y=0.377
+ $X2=3.9 $Y2=0.377
r107 85 91 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.56
+ $Y2=0
r108 84 87 2.70378 $w=9.23e-07 $l=2.05e-07 $layer=LI1_cond $X=3.6 $Y=0.377
+ $X2=3.805 $Y2=0.377
r109 84 85 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r110 81 84 9.16649 $w=9.23e-07 $l=6.95e-07 $layer=LI1_cond $X=2.905 $Y=0.377
+ $X2=3.6 $Y2=0.377
r111 81 82 11.4973 $w=9.23e-07 $l=9.5e-08 $layer=LI1_cond $X=2.905 $Y=0.377
+ $X2=2.81 $Y2=0.377
r112 78 79 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r113 75 97 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.84 $Y=0 $X2=9.36
+ $Y2=0
r114 74 75 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.84 $Y=0 $X2=9.84
+ $Y2=0
r115 72 96 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.46 $Y=0 $X2=9.295
+ $Y2=0
r116 72 74 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=9.46 $Y=0 $X2=9.84
+ $Y2=0
r117 71 97 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=0 $X2=9.36
+ $Y2=0
r118 71 94 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=0 $X2=8.4
+ $Y2=0
r119 70 71 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=0 $X2=8.88
+ $Y2=0
r120 68 93 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.6 $Y=0 $X2=8.435
+ $Y2=0
r121 68 70 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=8.6 $Y=0 $X2=8.88
+ $Y2=0
r122 67 96 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.13 $Y=0 $X2=9.295
+ $Y2=0
r123 67 70 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=9.13 $Y=0 $X2=8.88
+ $Y2=0
r124 66 94 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=0 $X2=8.4
+ $Y2=0
r125 65 66 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=7.92 $Y=0
+ $X2=7.92 $Y2=0
r126 62 65 187.893 $w=1.68e-07 $l=2.88e-06 $layer=LI1_cond $X=5.04 $Y=0 $X2=7.92
+ $Y2=0
r127 60 90 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.83 $Y=0 $X2=4.665
+ $Y2=0
r128 60 62 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=4.83 $Y=0 $X2=5.04
+ $Y2=0
r129 59 93 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.27 $Y=0 $X2=8.435
+ $Y2=0
r130 59 65 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=8.27 $Y=0 $X2=7.92
+ $Y2=0
r131 58 85 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.6
+ $Y2=0
r132 57 82 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=2.64 $Y=0 $X2=2.81
+ $Y2=0
r133 57 58 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r134 54 58 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.64
+ $Y2=0
r135 54 79 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r136 53 54 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r137 51 78 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.35 $Y=0 $X2=1.185
+ $Y2=0
r138 51 53 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=1.35 $Y=0 $X2=1.68
+ $Y2=0
r139 49 79 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r140 48 49 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r141 46 78 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.02 $Y=0 $X2=1.185
+ $Y2=0
r142 46 48 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=1.02 $Y=0 $X2=0.72
+ $Y2=0
r143 44 66 0.802756 $w=4.9e-07 $l=2.88e-06 $layer=MET1_cond $X=5.04 $Y=0
+ $X2=7.92 $Y2=0
r144 44 91 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=4.56
+ $Y2=0
r145 44 62 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=5.04 $Y=0
+ $X2=5.04 $Y2=0
r146 42 53 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=1.88 $Y=0 $X2=1.68
+ $Y2=0
r147 42 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.88 $Y=0 $X2=2.045
+ $Y2=0
r148 41 57 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=2.21 $Y=0 $X2=2.64
+ $Y2=0
r149 41 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.21 $Y=0 $X2=2.045
+ $Y2=0
r150 37 96 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.295 $Y=0.085
+ $X2=9.295 $Y2=0
r151 37 39 20.6043 $w=3.28e-07 $l=5.9e-07 $layer=LI1_cond $X=9.295 $Y=0.085
+ $X2=9.295 $Y2=0.675
r152 33 93 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.435 $Y=0.085
+ $X2=8.435 $Y2=0
r153 33 35 20.6043 $w=3.28e-07 $l=5.9e-07 $layer=LI1_cond $X=8.435 $Y=0.085
+ $X2=8.435 $Y2=0.675
r154 29 90 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.665 $Y=0.085
+ $X2=4.665 $Y2=0
r155 29 31 19.382 $w=3.28e-07 $l=5.55e-07 $layer=LI1_cond $X=4.665 $Y=0.085
+ $X2=4.665 $Y2=0.64
r156 27 90 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.5 $Y=0 $X2=4.665
+ $Y2=0
r157 27 88 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=4.5 $Y=0 $X2=3.9
+ $Y2=0
r158 23 43 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.045 $Y=0.085
+ $X2=2.045 $Y2=0
r159 23 25 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=2.045 $Y=0.085
+ $X2=2.045 $Y2=0.55
r160 19 78 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.185 $Y=0.085
+ $X2=1.185 $Y2=0
r161 19 21 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=1.185 $Y=0.085
+ $X2=1.185 $Y2=0.55
r162 6 39 182 $w=1.7e-07 $l=3.68409e-07 $layer=licon1_NDIFF $count=1 $X=9.155
+ $Y=0.37 $X2=9.295 $Y2=0.675
r163 5 35 182 $w=1.7e-07 $l=3.68409e-07 $layer=licon1_NDIFF $count=1 $X=8.295
+ $Y=0.37 $X2=8.435 $Y2=0.675
r164 4 31 182 $w=1.7e-07 $l=3.32716e-07 $layer=licon1_NDIFF $count=1 $X=4.525
+ $Y=0.37 $X2=4.665 $Y2=0.64
r165 3 87 121.333 $w=1.7e-07 $l=1.18271e-06 $layer=licon1_NDIFF $count=1
+ $X=2.765 $Y=0.37 $X2=3.805 $Y2=0.675
r166 3 81 121.333 $w=1.7e-07 $l=3.68409e-07 $layer=licon1_NDIFF $count=1
+ $X=2.765 $Y=0.37 $X2=2.905 $Y2=0.675
r167 2 25 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=1.905
+ $Y=0.37 $X2=2.045 $Y2=0.55
r168 1 21 182 $w=1.7e-07 $l=2.34307e-07 $layer=licon1_NDIFF $count=1 $X=1.06
+ $Y=0.37 $X2=1.185 $Y2=0.55
.ends

.subckt PM_SKY130_FD_SC_HS__A2111OI_4%A_1228_74# 1 2 3 4 5 18 20 24 25 28 30 34
+ 39 42 43 46
c59 20 0 1.6164e-19 $X=8.005 $Y=0.6
r60 41 43 4.37153 $w=3.28e-07 $l=1.05e-07 $layer=LI1_cond $X=7.145 $Y=0.515
+ $X2=7.25 $Y2=0.515
r61 41 42 4.37153 $w=3.28e-07 $l=1.05e-07 $layer=LI1_cond $X=7.145 $Y=0.515
+ $X2=7.04 $Y2=0.515
r62 39 42 30.4245 $w=2.48e-07 $l=6.6e-07 $layer=LI1_cond $X=6.38 $Y=0.475
+ $X2=7.04 $Y2=0.475
r63 37 39 4.02231 $w=3.28e-07 $l=9.5e-08 $layer=LI1_cond $X=6.285 $Y=0.515
+ $X2=6.38 $Y2=0.515
r64 32 34 22.8184 $w=2.48e-07 $l=4.95e-07 $layer=LI1_cond $X=9.765 $Y=1.01
+ $X2=9.765 $Y2=0.515
r65 31 46 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.95 $Y=1.095
+ $X2=8.865 $Y2=1.095
r66 30 32 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=9.64 $Y=1.095
+ $X2=9.765 $Y2=1.01
r67 30 31 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=9.64 $Y=1.095
+ $X2=8.95 $Y2=1.095
r68 26 46 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.865 $Y=1.01
+ $X2=8.865 $Y2=1.095
r69 26 28 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=8.865 $Y=1.01
+ $X2=8.865 $Y2=0.515
r70 24 46 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.78 $Y=1.095
+ $X2=8.865 $Y2=1.095
r71 24 25 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=8.78 $Y=1.095
+ $X2=8.09 $Y2=1.095
r72 21 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.005 $Y=1.01
+ $X2=8.09 $Y2=1.095
r73 21 23 2.93583 $w=1.68e-07 $l=4.5e-08 $layer=LI1_cond $X=8.005 $Y=1.01
+ $X2=8.005 $Y2=0.965
r74 20 45 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.005 $Y=0.6
+ $X2=8.005 $Y2=0.475
r75 20 23 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=8.005 $Y=0.6
+ $X2=8.005 $Y2=0.965
r76 18 45 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=7.92 $Y=0.475
+ $X2=8.005 $Y2=0.475
r77 18 43 30.8855 $w=2.48e-07 $l=6.7e-07 $layer=LI1_cond $X=7.92 $Y=0.475
+ $X2=7.25 $Y2=0.475
r78 5 34 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=9.585
+ $Y=0.37 $X2=9.725 $Y2=0.515
r79 4 28 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=8.725
+ $Y=0.37 $X2=8.865 $Y2=0.515
r80 3 45 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=7.865
+ $Y=0.37 $X2=8.005 $Y2=0.515
r81 3 23 182 $w=1.7e-07 $l=6.61306e-07 $layer=licon1_NDIFF $count=1 $X=7.865
+ $Y=0.37 $X2=8.005 $Y2=0.965
r82 2 41 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=7.005
+ $Y=0.37 $X2=7.145 $Y2=0.515
r83 1 37 182 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=1 $X=6.14
+ $Y=0.37 $X2=6.285 $Y2=0.515
.ends

