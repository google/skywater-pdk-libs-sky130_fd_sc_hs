/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */

`ifndef SKY130_FD_SC_HS__NOR4BB_TB_V
`define SKY130_FD_SC_HS__NOR4BB_TB_V

/**
 * nor4bb: 4-input NOR, first two inputs inverted.
 *
 * Autogenerated test bench.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none

`include "sky130_fd_sc_hs__nor4bb.v"

module top();

    // Inputs are registered
    reg A;
    reg B;
    reg C_N;
    reg D_N;
    reg VPWR;
    reg VGND;

    // Outputs are wires
    wire Y;

    initial
    begin
        // Initial state is x for all inputs.
        A    = 1'bX;
        B    = 1'bX;
        C_N  = 1'bX;
        D_N  = 1'bX;
        VGND = 1'bX;
        VPWR = 1'bX;

        #20   A    = 1'b0;
        #40   B    = 1'b0;
        #60   C_N  = 1'b0;
        #80   D_N  = 1'b0;
        #100  VGND = 1'b0;
        #120  VPWR = 1'b0;
        #140  A    = 1'b1;
        #160  B    = 1'b1;
        #180  C_N  = 1'b1;
        #200  D_N  = 1'b1;
        #220  VGND = 1'b1;
        #240  VPWR = 1'b1;
        #260  A    = 1'b0;
        #280  B    = 1'b0;
        #300  C_N  = 1'b0;
        #320  D_N  = 1'b0;
        #340  VGND = 1'b0;
        #360  VPWR = 1'b0;
        #380  VPWR = 1'b1;
        #400  VGND = 1'b1;
        #420  D_N  = 1'b1;
        #440  C_N  = 1'b1;
        #460  B    = 1'b1;
        #480  A    = 1'b1;
        #500  VPWR = 1'bx;
        #520  VGND = 1'bx;
        #540  D_N  = 1'bx;
        #560  C_N  = 1'bx;
        #580  B    = 1'bx;
        #600  A    = 1'bx;
    end

    sky130_fd_sc_hs__nor4bb dut (.A(A), .B(B), .C_N(C_N), .D_N(D_N), .VPWR(VPWR), .VGND(VGND), .Y(Y));

endmodule

`default_nettype wire
`endif  // SKY130_FD_SC_HS__NOR4BB_TB_V
