* File: sky130_fd_sc_hs__edfxbp_1.pxi.spice
* Created: Thu Aug 27 20:44:28 2020
* 
x_PM_SKY130_FD_SC_HS__EDFXBP_1%D N_D_c_285_n N_D_c_290_n N_D_c_291_n N_D_M1000_g
+ N_D_M1031_g D D N_D_c_287_n N_D_c_288_n N_D_c_293_n
+ PM_SKY130_FD_SC_HS__EDFXBP_1%D
x_PM_SKY130_FD_SC_HS__EDFXBP_1%A_161_446# N_A_161_446#_M1028_s
+ N_A_161_446#_M1032_s N_A_161_446#_c_337_n N_A_161_446#_M1023_g
+ N_A_161_446#_M1001_g N_A_161_446#_c_330_n N_A_161_446#_c_331_n
+ N_A_161_446#_c_332_n N_A_161_446#_c_333_n N_A_161_446#_c_339_n
+ N_A_161_446#_c_340_n N_A_161_446#_c_334_n N_A_161_446#_c_341_n
+ N_A_161_446#_c_342_n N_A_161_446#_c_335_n N_A_161_446#_c_336_n
+ N_A_161_446#_c_376_p PM_SKY130_FD_SC_HS__EDFXBP_1%A_161_446#
x_PM_SKY130_FD_SC_HS__EDFXBP_1%DE N_DE_c_436_n N_DE_M1019_g N_DE_c_437_n
+ N_DE_c_438_n N_DE_c_439_n N_DE_c_440_n N_DE_c_441_n N_DE_M1032_g N_DE_c_442_n
+ N_DE_M1028_g N_DE_c_446_n N_DE_c_447_n N_DE_c_448_n N_DE_M1020_g N_DE_c_443_n
+ N_DE_c_449_n DE PM_SKY130_FD_SC_HS__EDFXBP_1%DE
x_PM_SKY130_FD_SC_HS__EDFXBP_1%A_575_48# N_A_575_48#_M1015_d N_A_575_48#_M1025_d
+ N_A_575_48#_M1002_g N_A_575_48#_c_538_n N_A_575_48#_c_539_n
+ N_A_575_48#_M1007_g N_A_575_48#_c_540_n N_A_575_48#_M1009_g
+ N_A_575_48#_M1010_g N_A_575_48#_c_524_n N_A_575_48#_M1004_g
+ N_A_575_48#_M1022_g N_A_575_48#_c_543_n N_A_575_48#_c_544_n
+ N_A_575_48#_c_526_n N_A_575_48#_c_527_n N_A_575_48#_c_528_n
+ N_A_575_48#_c_529_n N_A_575_48#_c_530_n N_A_575_48#_c_545_n
+ N_A_575_48#_c_531_n N_A_575_48#_c_532_n N_A_575_48#_c_533_n
+ N_A_575_48#_c_534_n N_A_575_48#_c_535_n N_A_575_48#_c_536_n
+ N_A_575_48#_c_550_n N_A_575_48#_c_551_n N_A_575_48#_c_537_n
+ PM_SKY130_FD_SC_HS__EDFXBP_1%A_575_48#
x_PM_SKY130_FD_SC_HS__EDFXBP_1%CLK N_CLK_c_754_n N_CLK_M1029_g N_CLK_c_755_n
+ N_CLK_M1005_g CLK PM_SKY130_FD_SC_HS__EDFXBP_1%CLK
x_PM_SKY130_FD_SC_HS__EDFXBP_1%A_1008_74# N_A_1008_74#_M1030_d
+ N_A_1008_74#_M1003_d N_A_1008_74#_c_813_n N_A_1008_74#_M1011_g
+ N_A_1008_74#_c_787_n N_A_1008_74#_M1013_g N_A_1008_74#_c_788_n
+ N_A_1008_74#_M1008_g N_A_1008_74#_c_789_n N_A_1008_74#_c_814_n
+ N_A_1008_74#_c_815_n N_A_1008_74#_M1012_g N_A_1008_74#_c_790_n
+ N_A_1008_74#_c_791_n N_A_1008_74#_c_792_n N_A_1008_74#_c_816_n
+ N_A_1008_74#_c_793_n N_A_1008_74#_c_794_n N_A_1008_74#_c_795_n
+ N_A_1008_74#_c_796_n N_A_1008_74#_c_889_p N_A_1008_74#_c_797_n
+ N_A_1008_74#_c_798_n N_A_1008_74#_c_799_n N_A_1008_74#_c_800_n
+ N_A_1008_74#_c_801_n N_A_1008_74#_c_802_n N_A_1008_74#_c_803_n
+ N_A_1008_74#_c_804_n N_A_1008_74#_c_820_n N_A_1008_74#_c_821_n
+ N_A_1008_74#_c_805_n N_A_1008_74#_c_806_n N_A_1008_74#_c_807_n
+ N_A_1008_74#_c_808_n N_A_1008_74#_c_809_n N_A_1008_74#_c_810_n
+ N_A_1008_74#_c_811_n N_A_1008_74#_c_812_n
+ PM_SKY130_FD_SC_HS__EDFXBP_1%A_1008_74#
x_PM_SKY130_FD_SC_HS__EDFXBP_1%A_818_74# N_A_818_74#_M1029_d N_A_818_74#_M1005_d
+ N_A_818_74#_M1030_g N_A_818_74#_c_1012_n N_A_818_74#_c_1031_n
+ N_A_818_74#_M1003_g N_A_818_74#_c_1013_n N_A_818_74#_M1033_g
+ N_A_818_74#_c_1015_n N_A_818_74#_c_1034_n N_A_818_74#_c_1035_n
+ N_A_818_74#_M1018_g N_A_818_74#_c_1016_n N_A_818_74#_M1024_g
+ N_A_818_74#_c_1017_n N_A_818_74#_c_1018_n N_A_818_74#_c_1019_n
+ N_A_818_74#_c_1020_n N_A_818_74#_M1027_g N_A_818_74#_c_1021_n
+ N_A_818_74#_c_1022_n N_A_818_74#_c_1023_n N_A_818_74#_c_1039_n
+ N_A_818_74#_c_1024_n N_A_818_74#_c_1041_n N_A_818_74#_c_1129_p
+ N_A_818_74#_c_1203_p N_A_818_74#_c_1042_n N_A_818_74#_c_1043_n
+ N_A_818_74#_c_1025_n N_A_818_74#_c_1026_n N_A_818_74#_c_1027_n
+ N_A_818_74#_c_1046_n N_A_818_74#_c_1047_n N_A_818_74#_c_1123_p
+ N_A_818_74#_c_1028_n N_A_818_74#_c_1029_n
+ PM_SKY130_FD_SC_HS__EDFXBP_1%A_818_74#
x_PM_SKY130_FD_SC_HS__EDFXBP_1%A_1419_71# N_A_1419_71#_M1014_d
+ N_A_1419_71#_M1016_d N_A_1419_71#_M1021_g N_A_1419_71#_c_1232_n
+ N_A_1419_71#_c_1243_n N_A_1419_71#_M1034_g N_A_1419_71#_M1006_g
+ N_A_1419_71#_c_1244_n N_A_1419_71#_c_1245_n N_A_1419_71#_M1026_g
+ N_A_1419_71#_c_1234_n N_A_1419_71#_c_1235_n N_A_1419_71#_c_1236_n
+ N_A_1419_71#_c_1246_n N_A_1419_71#_c_1247_n N_A_1419_71#_c_1237_n
+ N_A_1419_71#_c_1238_n N_A_1419_71#_c_1239_n N_A_1419_71#_c_1240_n
+ N_A_1419_71#_c_1241_n N_A_1419_71#_c_1249_n
+ PM_SKY130_FD_SC_HS__EDFXBP_1%A_1419_71#
x_PM_SKY130_FD_SC_HS__EDFXBP_1%A_1198_97# N_A_1198_97#_M1033_d
+ N_A_1198_97#_M1011_d N_A_1198_97#_c_1368_n N_A_1198_97#_M1014_g
+ N_A_1198_97#_c_1369_n N_A_1198_97#_c_1370_n N_A_1198_97#_M1016_g
+ N_A_1198_97#_c_1371_n N_A_1198_97#_c_1372_n N_A_1198_97#_c_1376_n
+ N_A_1198_97#_c_1373_n N_A_1198_97#_c_1374_n N_A_1198_97#_c_1379_n
+ PM_SKY130_FD_SC_HS__EDFXBP_1%A_1198_97#
x_PM_SKY130_FD_SC_HS__EDFXBP_1%A_1879_74# N_A_1879_74#_M1008_d
+ N_A_1879_74#_M1024_d N_A_1879_74#_M1015_g N_A_1879_74#_c_1480_n
+ N_A_1879_74#_M1025_g N_A_1879_74#_c_1471_n N_A_1879_74#_c_1472_n
+ N_A_1879_74#_c_1473_n N_A_1879_74#_M1017_g N_A_1879_74#_c_1474_n
+ N_A_1879_74#_c_1483_n N_A_1879_74#_M1035_g N_A_1879_74#_c_1475_n
+ N_A_1879_74#_c_1518_n N_A_1879_74#_c_1484_n N_A_1879_74#_c_1485_n
+ N_A_1879_74#_c_1486_n N_A_1879_74#_c_1476_n N_A_1879_74#_c_1477_n
+ N_A_1879_74#_c_1478_n N_A_1879_74#_c_1479_n
+ PM_SKY130_FD_SC_HS__EDFXBP_1%A_1879_74#
x_PM_SKY130_FD_SC_HS__EDFXBP_1%A_27_74# N_A_27_74#_M1031_s N_A_27_74#_M1002_d
+ N_A_27_74#_M1033_s N_A_27_74#_M1000_s N_A_27_74#_M1007_d N_A_27_74#_M1011_s
+ N_A_27_74#_c_1599_n N_A_27_74#_c_1607_n N_A_27_74#_c_1608_n
+ N_A_27_74#_c_1609_n N_A_27_74#_c_1610_n N_A_27_74#_c_1611_n
+ N_A_27_74#_c_1646_n N_A_27_74#_c_1612_n N_A_27_74#_c_1613_n
+ N_A_27_74#_c_1614_n N_A_27_74#_c_1600_n N_A_27_74#_c_1616_n
+ N_A_27_74#_c_1601_n N_A_27_74#_c_1677_n N_A_27_74#_c_1602_n
+ N_A_27_74#_c_1603_n N_A_27_74#_c_1705_n N_A_27_74#_c_1618_n
+ N_A_27_74#_c_1619_n N_A_27_74#_c_1604_n N_A_27_74#_c_1620_n
+ N_A_27_74#_c_1605_n N_A_27_74#_c_1621_n N_A_27_74#_c_1738_p
+ PM_SKY130_FD_SC_HS__EDFXBP_1%A_27_74#
x_PM_SKY130_FD_SC_HS__EDFXBP_1%VPWR N_VPWR_M1023_d N_VPWR_M1032_d N_VPWR_M1005_s
+ N_VPWR_M1003_s N_VPWR_M1034_d N_VPWR_M1026_s N_VPWR_M1009_d N_VPWR_M1035_d
+ N_VPWR_c_1778_n N_VPWR_c_1779_n N_VPWR_c_1780_n N_VPWR_c_1781_n
+ N_VPWR_c_1782_n N_VPWR_c_1783_n N_VPWR_c_1784_n N_VPWR_c_1785_n
+ N_VPWR_c_1786_n N_VPWR_c_1787_n N_VPWR_c_1788_n N_VPWR_c_1789_n VPWR
+ N_VPWR_c_1790_n N_VPWR_c_1791_n N_VPWR_c_1792_n N_VPWR_c_1793_n
+ N_VPWR_c_1794_n N_VPWR_c_1795_n N_VPWR_c_1796_n N_VPWR_c_1777_n
+ N_VPWR_c_1798_n N_VPWR_c_1799_n N_VPWR_c_1800_n N_VPWR_c_1801_n
+ N_VPWR_c_1802_n N_VPWR_c_1803_n PM_SKY130_FD_SC_HS__EDFXBP_1%VPWR
x_PM_SKY130_FD_SC_HS__EDFXBP_1%Q N_Q_M1017_s N_Q_M1035_s N_Q_c_1939_n Q Q Q Q
+ N_Q_c_1940_n PM_SKY130_FD_SC_HS__EDFXBP_1%Q
x_PM_SKY130_FD_SC_HS__EDFXBP_1%Q_N N_Q_N_M1022_d N_Q_N_M1004_d N_Q_N_c_1975_n
+ N_Q_N_c_1976_n N_Q_N_c_1972_n Q_N Q_N Q_N PM_SKY130_FD_SC_HS__EDFXBP_1%Q_N
x_PM_SKY130_FD_SC_HS__EDFXBP_1%VGND N_VGND_M1019_d N_VGND_M1028_d N_VGND_M1029_s
+ N_VGND_M1030_s N_VGND_M1021_d N_VGND_M1006_s N_VGND_M1010_d N_VGND_M1017_d
+ N_VGND_c_1992_n N_VGND_c_1993_n N_VGND_c_1994_n N_VGND_c_1995_n
+ N_VGND_c_1996_n N_VGND_c_1997_n N_VGND_c_1998_n N_VGND_c_1999_n
+ N_VGND_c_2000_n N_VGND_c_2001_n N_VGND_c_2002_n N_VGND_c_2003_n
+ N_VGND_c_2004_n N_VGND_c_2005_n VGND N_VGND_c_2006_n N_VGND_c_2007_n
+ N_VGND_c_2008_n N_VGND_c_2009_n N_VGND_c_2010_n N_VGND_c_2011_n
+ N_VGND_c_2012_n N_VGND_c_2013_n N_VGND_c_2014_n N_VGND_c_2015_n
+ N_VGND_c_2016_n N_VGND_c_2017_n PM_SKY130_FD_SC_HS__EDFXBP_1%VGND
cc_1 VNB N_D_c_285_n 0.041714f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.82
cc_2 VNB N_D_M1031_g 0.0264821f $X=-0.19 $Y=-0.245 $X2=0.65 $Y2=0.58
cc_3 VNB N_D_c_287_n 0.019855f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.145
cc_4 VNB N_D_c_288_n 0.0144514f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.145
cc_5 VNB N_A_161_446#_M1001_g 0.0217822f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_6 VNB N_A_161_446#_c_330_n 0.00292476f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.825
cc_7 VNB N_A_161_446#_c_331_n 0.0209793f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.99
cc_8 VNB N_A_161_446#_c_332_n 0.00930926f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.145
cc_9 VNB N_A_161_446#_c_333_n 0.00574061f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_161_446#_c_334_n 0.00446641f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.825
cc_11 VNB N_A_161_446#_c_335_n 0.00272114f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_161_446#_c_336_n 0.0627118f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_DE_c_436_n 0.0175428f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.15
cc_14 VNB N_DE_c_437_n 0.0279279f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.375
cc_15 VNB N_DE_c_438_n 0.0100448f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.465
cc_16 VNB N_DE_c_439_n 0.0273555f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.75
cc_17 VNB N_DE_c_440_n 0.0224499f $X=-0.19 $Y=-0.245 $X2=0.65 $Y2=0.98
cc_18 VNB N_DE_c_441_n 0.0270689f $X=-0.19 $Y=-0.245 $X2=0.65 $Y2=0.58
cc_19 VNB N_DE_c_442_n 0.0186656f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_20 VNB N_DE_c_443_n 0.00774539f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.99
cc_21 VNB DE 0.00150919f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.295
cc_22 VNB N_A_575_48#_M1002_g 0.0246002f $X=-0.19 $Y=-0.245 $X2=0.65 $Y2=0.58
cc_23 VNB N_A_575_48#_M1010_g 0.045306f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.825
cc_24 VNB N_A_575_48#_c_524_n 0.0344741f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.99
cc_25 VNB N_A_575_48#_M1022_g 0.0284483f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.665
cc_26 VNB N_A_575_48#_c_526_n 0.0200797f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_575_48#_c_527_n 0.00279267f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_575_48#_c_528_n 0.00120373f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_575_48#_c_529_n 0.00168099f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_575_48#_c_530_n 0.0085702f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_575_48#_c_531_n 0.0659711f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_575_48#_c_532_n 0.00254619f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_575_48#_c_533_n 0.00126737f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_575_48#_c_534_n 0.0176138f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_575_48#_c_535_n 0.0016809f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_575_48#_c_536_n 0.0408674f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_575_48#_c_537_n 0.0107368f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_CLK_c_754_n 0.0213924f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.15
cc_39 VNB N_CLK_c_755_n 0.0782816f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.375
cc_40 VNB CLK 0.0118889f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.75
cc_41 VNB N_A_1008_74#_c_787_n 0.0182334f $X=-0.19 $Y=-0.245 $X2=0.65 $Y2=0.58
cc_42 VNB N_A_1008_74#_c_788_n 0.0187258f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_43 VNB N_A_1008_74#_c_789_n 0.0065214f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.145
cc_44 VNB N_A_1008_74#_c_790_n 0.00907777f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_A_1008_74#_c_791_n 0.0170049f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_A_1008_74#_c_792_n 0.00365087f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.665
cc_47 VNB N_A_1008_74#_c_793_n 0.00583653f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_1008_74#_c_794_n 0.0178019f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A_1008_74#_c_795_n 0.00114445f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_A_1008_74#_c_796_n 0.0184433f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_A_1008_74#_c_797_n 0.0111546f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_A_1008_74#_c_798_n 0.00202577f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_A_1008_74#_c_799_n 0.0119359f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_A_1008_74#_c_800_n 0.0036851f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_A_1008_74#_c_801_n 0.00963275f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_A_1008_74#_c_802_n 0.00297237f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_A_1008_74#_c_803_n 0.0163761f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_A_1008_74#_c_804_n 0.00123754f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_A_1008_74#_c_805_n 0.0018569f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_A_1008_74#_c_806_n 0.0389267f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_A_1008_74#_c_807_n 0.00846462f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_A_1008_74#_c_808_n 0.00364081f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_A_1008_74#_c_809_n 0.00938941f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_A_1008_74#_c_810_n 0.035551f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_A_1008_74#_c_811_n 0.00218263f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_A_1008_74#_c_812_n 0.0222493f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_A_818_74#_M1030_g 0.0461962f $X=-0.19 $Y=-0.245 $X2=0.65 $Y2=0.58
cc_68 VNB N_A_818_74#_c_1012_n 0.0107077f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_A_818_74#_c_1013_n 0.00734855f $X=-0.19 $Y=-0.245 $X2=0.585
+ $Y2=1.145
cc_70 VNB N_A_818_74#_M1033_g 0.0560652f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.825
cc_71 VNB N_A_818_74#_c_1015_n 0.024465f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.825
cc_72 VNB N_A_818_74#_c_1016_n 0.0240266f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_A_818_74#_c_1017_n 0.0123623f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_A_818_74#_c_1018_n 0.0279517f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_A_818_74#_c_1019_n 0.00921092f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_A_818_74#_c_1020_n 0.022969f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_A_818_74#_c_1021_n 0.00581916f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_A_818_74#_c_1022_n 7.16371e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VNB N_A_818_74#_c_1023_n 0.00820438f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_A_818_74#_c_1024_n 0.0124455f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_81 VNB N_A_818_74#_c_1025_n 0.00356635f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_82 VNB N_A_818_74#_c_1026_n 7.42552e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_83 VNB N_A_818_74#_c_1027_n 0.00873055f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_84 VNB N_A_818_74#_c_1028_n 0.00166024f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_85 VNB N_A_818_74#_c_1029_n 0.0114709f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_86 VNB N_A_1419_71#_M1021_g 0.0290994f $X=-0.19 $Y=-0.245 $X2=0.65 $Y2=0.58
cc_87 VNB N_A_1419_71#_c_1232_n 0.00200085f $X=-0.19 $Y=-0.245 $X2=0.635
+ $Y2=1.21
cc_88 VNB N_A_1419_71#_M1006_g 0.0492905f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.145
cc_89 VNB N_A_1419_71#_c_1234_n 0.00667676f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_90 VNB N_A_1419_71#_c_1235_n 0.00737941f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_91 VNB N_A_1419_71#_c_1236_n 0.0183664f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_92 VNB N_A_1419_71#_c_1237_n 0.00152844f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_93 VNB N_A_1419_71#_c_1238_n 0.0134958f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_94 VNB N_A_1419_71#_c_1239_n 0.0560647f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_95 VNB N_A_1419_71#_c_1240_n 0.00675239f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_96 VNB N_A_1419_71#_c_1241_n 3.38536e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_97 VNB N_A_1198_97#_c_1368_n 0.0189225f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.75
cc_98 VNB N_A_1198_97#_c_1369_n 0.024814f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_99 VNB N_A_1198_97#_c_1370_n 0.00850451f $X=-0.19 $Y=-0.245 $X2=0.635
+ $Y2=1.21
cc_100 VNB N_A_1198_97#_c_1371_n 0.0216361f $X=-0.19 $Y=-0.245 $X2=0.59
+ $Y2=1.145
cc_101 VNB N_A_1198_97#_c_1372_n 0.0149445f $X=-0.19 $Y=-0.245 $X2=0.59
+ $Y2=1.825
cc_102 VNB N_A_1198_97#_c_1373_n 0.00530369f $X=-0.19 $Y=-0.245 $X2=0.63
+ $Y2=1.295
cc_103 VNB N_A_1198_97#_c_1374_n 2.82323e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_104 VNB N_A_1879_74#_M1015_g 0.0240975f $X=-0.19 $Y=-0.245 $X2=0.65 $Y2=0.58
cc_105 VNB N_A_1879_74#_c_1471_n 0.0609545f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_106 VNB N_A_1879_74#_c_1472_n 0.0696067f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_107 VNB N_A_1879_74#_c_1473_n 0.0182405f $X=-0.19 $Y=-0.245 $X2=0.585
+ $Y2=1.145
cc_108 VNB N_A_1879_74#_c_1474_n 0.00836489f $X=-0.19 $Y=-0.245 $X2=0.585
+ $Y2=1.825
cc_109 VNB N_A_1879_74#_c_1475_n 0.0330367f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_110 VNB N_A_1879_74#_c_1476_n 0.00123731f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_111 VNB N_A_1879_74#_c_1477_n 8.61664e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_112 VNB N_A_1879_74#_c_1478_n 0.0065731f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_113 VNB N_A_1879_74#_c_1479_n 0.00234911f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_114 VNB N_A_27_74#_c_1599_n 0.0427491f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.825
cc_115 VNB N_A_27_74#_c_1600_n 0.0180358f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_116 VNB N_A_27_74#_c_1601_n 0.00312015f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_117 VNB N_A_27_74#_c_1602_n 0.0161129f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_118 VNB N_A_27_74#_c_1603_n 0.0133157f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_119 VNB N_A_27_74#_c_1604_n 0.0141371f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_120 VNB N_A_27_74#_c_1605_n 0.019915f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_121 VNB N_VPWR_c_1777_n 0.601534f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_122 VNB N_Q_c_1939_n 0.00404267f $X=-0.19 $Y=-0.245 $X2=0.65 $Y2=0.58
cc_123 VNB N_Q_c_1940_n 0.0030048f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_124 VNB N_Q_N_c_1972_n 0.0239297f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_125 VNB Q_N 0.0266902f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.145
cc_126 VNB Q_N 0.00940311f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.145
cc_127 VNB N_VGND_c_1992_n 0.014248f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_128 VNB N_VGND_c_1993_n 0.0144254f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_129 VNB N_VGND_c_1994_n 0.00864424f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_130 VNB N_VGND_c_1995_n 0.00998138f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_131 VNB N_VGND_c_1996_n 0.00857507f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_132 VNB N_VGND_c_1997_n 0.00590394f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_133 VNB N_VGND_c_1998_n 0.0176957f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_134 VNB N_VGND_c_1999_n 0.0105004f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_135 VNB N_VGND_c_2000_n 0.0216973f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_136 VNB N_VGND_c_2001_n 0.00616716f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_137 VNB N_VGND_c_2002_n 0.0341929f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_138 VNB N_VGND_c_2003_n 0.00326991f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_139 VNB N_VGND_c_2004_n 0.0196495f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_140 VNB N_VGND_c_2005_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_141 VNB N_VGND_c_2006_n 0.0331655f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_142 VNB N_VGND_c_2007_n 0.0563089f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_143 VNB N_VGND_c_2008_n 0.0296519f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_144 VNB N_VGND_c_2009_n 0.0784082f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_145 VNB N_VGND_c_2010_n 0.0392606f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_146 VNB N_VGND_c_2011_n 0.0193429f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_147 VNB N_VGND_c_2012_n 0.814432f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_148 VNB N_VGND_c_2013_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_149 VNB N_VGND_c_2014_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_150 VNB N_VGND_c_2015_n 0.00461913f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_151 VNB N_VGND_c_2016_n 0.00634377f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_152 VNB N_VGND_c_2017_n 0.00326991f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_153 VPB N_D_c_285_n 0.0114858f $X=-0.19 $Y=1.66 $X2=0.585 $Y2=1.82
cc_154 VPB N_D_c_290_n 0.0240039f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.375
cc_155 VPB N_D_c_291_n 0.0258254f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.465
cc_156 VPB N_D_c_288_n 0.00469484f $X=-0.19 $Y=1.66 $X2=0.59 $Y2=1.145
cc_157 VPB N_D_c_293_n 0.0168466f $X=-0.19 $Y=1.66 $X2=0.59 $Y2=1.825
cc_158 VPB N_A_161_446#_c_337_n 0.0740675f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.75
cc_159 VPB N_A_161_446#_c_331_n 0.0207722f $X=-0.19 $Y=1.66 $X2=0.585 $Y2=1.99
cc_160 VPB N_A_161_446#_c_339_n 0.0112962f $X=-0.19 $Y=1.66 $X2=0.63 $Y2=1.295
cc_161 VPB N_A_161_446#_c_340_n 0.00373221f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_162 VPB N_A_161_446#_c_341_n 0.0040597f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_163 VPB N_A_161_446#_c_342_n 0.00708453f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_164 VPB N_A_161_446#_c_335_n 0.00403255f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_165 VPB N_DE_c_441_n 0.0719849f $X=-0.19 $Y=1.66 $X2=0.65 $Y2=0.58
cc_166 VPB N_DE_c_446_n 0.02786f $X=-0.19 $Y=1.66 $X2=0.585 $Y2=1.145
cc_167 VPB N_DE_c_447_n 0.010137f $X=-0.19 $Y=1.66 $X2=0.585 $Y2=0.98
cc_168 VPB N_DE_c_448_n 0.0151978f $X=-0.19 $Y=1.66 $X2=0.585 $Y2=1.825
cc_169 VPB N_DE_c_449_n 0.0284461f $X=-0.19 $Y=1.66 $X2=0.63 $Y2=1.145
cc_170 VPB DE 9.123e-19 $X=-0.19 $Y=1.66 $X2=0.63 $Y2=1.295
cc_171 VPB N_A_575_48#_c_538_n 0.0229898f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.21
cc_172 VPB N_A_575_48#_c_539_n 0.0225638f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_173 VPB N_A_575_48#_c_540_n 0.0194365f $X=-0.19 $Y=1.66 $X2=0.585 $Y2=1.145
cc_174 VPB N_A_575_48#_M1010_g 0.00317119f $X=-0.19 $Y=1.66 $X2=0.59 $Y2=1.825
cc_175 VPB N_A_575_48#_c_524_n 0.0273367f $X=-0.19 $Y=1.66 $X2=0.585 $Y2=1.99
cc_176 VPB N_A_575_48#_c_543_n 0.00700003f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_177 VPB N_A_575_48#_c_544_n 0.00271237f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_178 VPB N_A_575_48#_c_545_n 0.00640871f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_179 VPB N_A_575_48#_c_531_n 0.0227564f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_180 VPB N_A_575_48#_c_532_n 9.66515e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_181 VPB N_A_575_48#_c_535_n 0.00173239f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_182 VPB N_A_575_48#_c_536_n 0.0149369f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_183 VPB N_A_575_48#_c_550_n 0.0175558f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_184 VPB N_A_575_48#_c_551_n 0.0537012f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_185 VPB N_A_575_48#_c_537_n 0.00109057f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_186 VPB N_CLK_c_755_n 0.0301276f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.375
cc_187 VPB N_A_1008_74#_c_813_n 0.0187952f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.75
cc_188 VPB N_A_1008_74#_c_814_n 0.0149904f $X=-0.19 $Y=1.66 $X2=0.585 $Y2=0.98
cc_189 VPB N_A_1008_74#_c_815_n 0.0225203f $X=-0.19 $Y=1.66 $X2=0.585 $Y2=1.825
cc_190 VPB N_A_1008_74#_c_816_n 0.00534977f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_191 VPB N_A_1008_74#_c_793_n 0.00110243f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_192 VPB N_A_1008_74#_c_802_n 8.50754e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_193 VPB N_A_1008_74#_c_803_n 0.0127272f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_194 VPB N_A_1008_74#_c_820_n 0.00813044f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_195 VPB N_A_1008_74#_c_821_n 0.0637016f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_196 VPB N_A_818_74#_c_1012_n 0.00996914f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_197 VPB N_A_818_74#_c_1031_n 0.0175655f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_198 VPB N_A_818_74#_c_1013_n 0.00712374f $X=-0.19 $Y=1.66 $X2=0.585 $Y2=1.145
cc_199 VPB N_A_818_74#_c_1015_n 0.0634601f $X=-0.19 $Y=1.66 $X2=0.59 $Y2=1.825
cc_200 VPB N_A_818_74#_c_1034_n 0.0140955f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_201 VPB N_A_818_74#_c_1035_n 0.0370204f $X=-0.19 $Y=1.66 $X2=0.63 $Y2=1.295
cc_202 VPB N_A_818_74#_c_1016_n 0.0396814f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_203 VPB N_A_818_74#_c_1021_n 0.00167153f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_204 VPB N_A_818_74#_c_1022_n 0.00551371f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_205 VPB N_A_818_74#_c_1039_n 0.00385875f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_206 VPB N_A_818_74#_c_1024_n 0.00203821f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_207 VPB N_A_818_74#_c_1041_n 0.00306526f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_208 VPB N_A_818_74#_c_1042_n 0.025258f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_209 VPB N_A_818_74#_c_1043_n 0.0211991f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_210 VPB N_A_818_74#_c_1025_n 0.00824485f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_211 VPB N_A_818_74#_c_1026_n 3.03225e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_212 VPB N_A_818_74#_c_1046_n 9.18152e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_213 VPB N_A_818_74#_c_1047_n 0.00609872f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_214 VPB N_A_818_74#_c_1028_n 0.00144674f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_215 VPB N_A_818_74#_c_1029_n 0.0482278f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_216 VPB N_A_1419_71#_c_1232_n 0.0422592f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.21
cc_217 VPB N_A_1419_71#_c_1243_n 0.0243791f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_218 VPB N_A_1419_71#_c_1244_n 0.0622546f $X=-0.19 $Y=1.66 $X2=0.585 $Y2=1.825
cc_219 VPB N_A_1419_71#_c_1245_n 0.0177737f $X=-0.19 $Y=1.66 $X2=0.59 $Y2=1.825
cc_220 VPB N_A_1419_71#_c_1246_n 0.00400808f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_221 VPB N_A_1419_71#_c_1247_n 0.00550153f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_222 VPB N_A_1419_71#_c_1238_n 0.0158398f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_223 VPB N_A_1419_71#_c_1249_n 0.0664579f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_224 VPB N_A_1198_97#_c_1370_n 0.0534383f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.21
cc_225 VPB N_A_1198_97#_c_1376_n 0.00920484f $X=-0.19 $Y=1.66 $X2=0.63 $Y2=1.145
cc_226 VPB N_A_1198_97#_c_1373_n 0.00213164f $X=-0.19 $Y=1.66 $X2=0.63 $Y2=1.295
cc_227 VPB N_A_1198_97#_c_1374_n 0.00427918f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_228 VPB N_A_1198_97#_c_1379_n 0.0152573f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_229 VPB N_A_1879_74#_c_1480_n 0.0172304f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_230 VPB N_A_1879_74#_c_1472_n 0.0146199f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_231 VPB N_A_1879_74#_c_1474_n 8.58573e-19 $X=-0.19 $Y=1.66 $X2=0.585
+ $Y2=1.825
cc_232 VPB N_A_1879_74#_c_1483_n 0.0263925f $X=-0.19 $Y=1.66 $X2=0.59 $Y2=1.825
cc_233 VPB N_A_1879_74#_c_1484_n 2.83835e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_234 VPB N_A_1879_74#_c_1485_n 0.0129297f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_235 VPB N_A_1879_74#_c_1486_n 0.0180664f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_236 VPB N_A_1879_74#_c_1477_n 0.00248469f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_237 VPB N_A_27_74#_c_1599_n 0.0300826f $X=-0.19 $Y=1.66 $X2=0.585 $Y2=1.825
cc_238 VPB N_A_27_74#_c_1607_n 0.0238102f $X=-0.19 $Y=1.66 $X2=0.585 $Y2=1.99
cc_239 VPB N_A_27_74#_c_1608_n 0.0223429f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_240 VPB N_A_27_74#_c_1609_n 0.00993635f $X=-0.19 $Y=1.66 $X2=0.63 $Y2=1.665
cc_241 VPB N_A_27_74#_c_1610_n 0.0107993f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_242 VPB N_A_27_74#_c_1611_n 0.00349119f $X=-0.19 $Y=1.66 $X2=0.63 $Y2=1.825
cc_243 VPB N_A_27_74#_c_1612_n 0.0166766f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_244 VPB N_A_27_74#_c_1613_n 0.00106188f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_245 VPB N_A_27_74#_c_1614_n 0.00954348f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_246 VPB N_A_27_74#_c_1600_n 0.015999f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_247 VPB N_A_27_74#_c_1616_n 0.0275417f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_248 VPB N_A_27_74#_c_1601_n 0.0012069f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_249 VPB N_A_27_74#_c_1618_n 0.00256831f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_250 VPB N_A_27_74#_c_1619_n 0.011152f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_251 VPB N_A_27_74#_c_1620_n 0.0143948f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_252 VPB N_A_27_74#_c_1621_n 0.00501496f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_253 VPB N_VPWR_c_1778_n 0.00600898f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_254 VPB N_VPWR_c_1779_n 0.00647584f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_255 VPB N_VPWR_c_1780_n 0.0102809f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_256 VPB N_VPWR_c_1781_n 0.0223379f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_257 VPB N_VPWR_c_1782_n 0.00744897f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_258 VPB N_VPWR_c_1783_n 0.021152f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_259 VPB N_VPWR_c_1784_n 0.0367693f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_260 VPB N_VPWR_c_1785_n 0.00779972f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_261 VPB N_VPWR_c_1786_n 0.0310451f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_262 VPB N_VPWR_c_1787_n 0.00614127f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_263 VPB N_VPWR_c_1788_n 0.0335097f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_264 VPB N_VPWR_c_1789_n 0.00621339f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_265 VPB N_VPWR_c_1790_n 0.0295786f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_266 VPB N_VPWR_c_1791_n 0.0297419f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_267 VPB N_VPWR_c_1792_n 0.0585373f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_268 VPB N_VPWR_c_1793_n 0.0399942f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_269 VPB N_VPWR_c_1794_n 0.047813f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_270 VPB N_VPWR_c_1795_n 0.03532f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_271 VPB N_VPWR_c_1796_n 0.0188734f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_272 VPB N_VPWR_c_1777_n 0.208332f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_273 VPB N_VPWR_c_1798_n 0.00460249f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_274 VPB N_VPWR_c_1799_n 0.00474673f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_275 VPB N_VPWR_c_1800_n 0.00631318f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_276 VPB N_VPWR_c_1801_n 0.00614127f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_277 VPB N_VPWR_c_1802_n 0.0150734f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_278 VPB N_VPWR_c_1803_n 0.00460249f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_279 VPB Q 0.00642009f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_280 VPB Q 0.0152801f $X=-0.19 $Y=1.66 $X2=0.59 $Y2=1.825
cc_281 VPB N_Q_c_1940_n 0.00392526f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_282 VPB N_Q_N_c_1975_n 0.0089215f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.75
cc_283 VPB N_Q_N_c_1976_n 0.0436171f $X=-0.19 $Y=1.66 $X2=0.65 $Y2=0.58
cc_284 VPB N_Q_N_c_1972_n 0.00779288f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_285 N_D_c_290_n N_A_161_446#_c_337_n 0.0227146f $X=0.505 $Y=2.375 $X2=0 $Y2=0
cc_286 N_D_c_291_n N_A_161_446#_c_337_n 0.0317302f $X=0.505 $Y=2.465 $X2=0 $Y2=0
cc_287 N_D_c_288_n N_A_161_446#_c_337_n 7.04333e-19 $X=0.59 $Y=1.145 $X2=0 $Y2=0
cc_288 N_D_c_293_n N_A_161_446#_c_337_n 0.0135156f $X=0.59 $Y=1.825 $X2=0 $Y2=0
cc_289 N_D_c_285_n N_A_161_446#_c_330_n 0.00156615f $X=0.585 $Y=1.82 $X2=0 $Y2=0
cc_290 N_D_c_288_n N_A_161_446#_c_330_n 0.054575f $X=0.59 $Y=1.145 $X2=0 $Y2=0
cc_291 N_D_c_285_n N_A_161_446#_c_331_n 0.0135156f $X=0.585 $Y=1.82 $X2=0 $Y2=0
cc_292 N_D_c_288_n N_A_161_446#_c_331_n 0.00328897f $X=0.59 $Y=1.145 $X2=0 $Y2=0
cc_293 N_D_c_287_n N_A_161_446#_c_333_n 0.00109278f $X=0.59 $Y=1.145 $X2=0 $Y2=0
cc_294 N_D_c_288_n N_A_161_446#_c_333_n 0.0152737f $X=0.59 $Y=1.145 $X2=0 $Y2=0
cc_295 N_D_c_290_n N_A_161_446#_c_340_n 7.49404e-19 $X=0.505 $Y=2.375 $X2=0
+ $Y2=0
cc_296 N_D_c_288_n N_A_161_446#_c_340_n 0.00337025f $X=0.59 $Y=1.145 $X2=0 $Y2=0
cc_297 N_D_M1031_g N_DE_c_436_n 0.0396236f $X=0.65 $Y=0.58 $X2=-0.19 $Y2=-0.245
cc_298 N_D_c_287_n N_DE_c_438_n 0.00230654f $X=0.59 $Y=1.145 $X2=0 $Y2=0
cc_299 N_D_c_288_n N_DE_c_438_n 9.15464e-19 $X=0.59 $Y=1.145 $X2=0 $Y2=0
cc_300 N_D_M1031_g N_A_27_74#_c_1599_n 0.00626394f $X=0.65 $Y=0.58 $X2=0 $Y2=0
cc_301 N_D_c_287_n N_A_27_74#_c_1599_n 0.0335765f $X=0.59 $Y=1.145 $X2=0 $Y2=0
cc_302 N_D_c_288_n N_A_27_74#_c_1599_n 0.0771094f $X=0.59 $Y=1.145 $X2=0 $Y2=0
cc_303 N_D_c_291_n N_A_27_74#_c_1607_n 0.011553f $X=0.505 $Y=2.465 $X2=0 $Y2=0
cc_304 N_D_c_290_n N_A_27_74#_c_1608_n 0.00467883f $X=0.505 $Y=2.375 $X2=0 $Y2=0
cc_305 N_D_c_291_n N_A_27_74#_c_1608_n 0.00819607f $X=0.505 $Y=2.465 $X2=0 $Y2=0
cc_306 N_D_c_288_n N_A_27_74#_c_1608_n 0.0199372f $X=0.59 $Y=1.145 $X2=0 $Y2=0
cc_307 N_D_c_293_n N_A_27_74#_c_1608_n 9.89815e-19 $X=0.59 $Y=1.825 $X2=0 $Y2=0
cc_308 N_D_M1031_g N_A_27_74#_c_1604_n 0.00616658f $X=0.65 $Y=0.58 $X2=0 $Y2=0
cc_309 N_D_c_287_n N_A_27_74#_c_1604_n 0.00132402f $X=0.59 $Y=1.145 $X2=0 $Y2=0
cc_310 N_D_c_288_n N_A_27_74#_c_1604_n 0.00941984f $X=0.59 $Y=1.145 $X2=0 $Y2=0
cc_311 N_D_c_290_n N_A_27_74#_c_1620_n 0.00289281f $X=0.505 $Y=2.375 $X2=0 $Y2=0
cc_312 N_D_c_291_n N_A_27_74#_c_1620_n 0.00198892f $X=0.505 $Y=2.465 $X2=0 $Y2=0
cc_313 N_D_c_288_n N_A_27_74#_c_1620_n 0.00101811f $X=0.59 $Y=1.145 $X2=0 $Y2=0
cc_314 N_D_c_291_n N_VPWR_c_1778_n 0.0015335f $X=0.505 $Y=2.465 $X2=0 $Y2=0
cc_315 N_D_c_291_n N_VPWR_c_1790_n 0.00445602f $X=0.505 $Y=2.465 $X2=0 $Y2=0
cc_316 N_D_c_291_n N_VPWR_c_1777_n 0.00899186f $X=0.505 $Y=2.465 $X2=0 $Y2=0
cc_317 N_D_M1031_g N_VGND_c_1992_n 0.00214336f $X=0.65 $Y=0.58 $X2=0 $Y2=0
cc_318 N_D_M1031_g N_VGND_c_2006_n 0.004347f $X=0.65 $Y=0.58 $X2=0 $Y2=0
cc_319 N_D_M1031_g N_VGND_c_2012_n 0.00822977f $X=0.65 $Y=0.58 $X2=0 $Y2=0
cc_320 N_A_161_446#_c_334_n N_DE_c_436_n 0.00204929f $X=1.825 $Y=0.645 $X2=-0.19
+ $Y2=-0.245
cc_321 N_A_161_446#_c_332_n N_DE_c_437_n 0.00766827f $X=1.65 $Y=1.195 $X2=0
+ $Y2=0
cc_322 N_A_161_446#_c_331_n N_DE_c_438_n 0.00755967f $X=1.17 $Y=1.615 $X2=0
+ $Y2=0
cc_323 N_A_161_446#_c_333_n N_DE_c_438_n 0.0060493f $X=1.335 $Y=1.195 $X2=0
+ $Y2=0
cc_324 N_A_161_446#_c_330_n N_DE_c_439_n 0.00641523f $X=1.17 $Y=1.615 $X2=0
+ $Y2=0
cc_325 N_A_161_446#_c_332_n N_DE_c_439_n 0.0138982f $X=1.65 $Y=1.195 $X2=0 $Y2=0
cc_326 N_A_161_446#_c_334_n N_DE_c_439_n 0.00444097f $X=1.825 $Y=0.645 $X2=0
+ $Y2=0
cc_327 N_A_161_446#_c_335_n N_DE_c_439_n 5.50673e-19 $X=2.5 $Y=1.145 $X2=0 $Y2=0
cc_328 N_A_161_446#_c_336_n N_DE_c_439_n 0.00405281f $X=2.5 $Y=1.145 $X2=0 $Y2=0
cc_329 N_A_161_446#_c_334_n N_DE_c_440_n 0.0131453f $X=1.825 $Y=0.645 $X2=0
+ $Y2=0
cc_330 N_A_161_446#_c_336_n N_DE_c_440_n 0.00231619f $X=2.5 $Y=1.145 $X2=0 $Y2=0
cc_331 N_A_161_446#_c_337_n N_DE_c_441_n 0.00109586f $X=0.895 $Y=2.465 $X2=0
+ $Y2=0
cc_332 N_A_161_446#_c_330_n N_DE_c_441_n 0.00167413f $X=1.17 $Y=1.615 $X2=0
+ $Y2=0
cc_333 N_A_161_446#_c_331_n N_DE_c_441_n 0.0330072f $X=1.17 $Y=1.615 $X2=0 $Y2=0
cc_334 N_A_161_446#_c_332_n N_DE_c_441_n 0.00335538f $X=1.65 $Y=1.195 $X2=0
+ $Y2=0
cc_335 N_A_161_446#_c_339_n N_DE_c_441_n 0.00618441f $X=1.715 $Y=2.035 $X2=0
+ $Y2=0
cc_336 N_A_161_446#_c_341_n N_DE_c_441_n 0.0088902f $X=1.8 $Y=2.505 $X2=0 $Y2=0
cc_337 N_A_161_446#_c_342_n N_DE_c_441_n 0.0200718f $X=2.335 $Y=2.035 $X2=0
+ $Y2=0
cc_338 N_A_161_446#_c_335_n N_DE_c_441_n 0.00883898f $X=2.5 $Y=1.145 $X2=0 $Y2=0
cc_339 N_A_161_446#_c_336_n N_DE_c_441_n 0.0124395f $X=2.5 $Y=1.145 $X2=0 $Y2=0
cc_340 N_A_161_446#_c_376_p N_DE_c_441_n 0.00789892f $X=1.8 $Y=2.035 $X2=0 $Y2=0
cc_341 N_A_161_446#_M1001_g N_DE_c_442_n 0.0163804f $X=2.56 $Y=0.58 $X2=0 $Y2=0
cc_342 N_A_161_446#_c_334_n N_DE_c_442_n 0.00629753f $X=1.825 $Y=0.645 $X2=0
+ $Y2=0
cc_343 N_A_161_446#_c_342_n N_DE_c_446_n 0.0149963f $X=2.335 $Y=2.035 $X2=0
+ $Y2=0
cc_344 N_A_161_446#_c_335_n N_DE_c_446_n 0.00717101f $X=2.5 $Y=1.145 $X2=0 $Y2=0
cc_345 N_A_161_446#_c_336_n N_DE_c_446_n 0.0140959f $X=2.5 $Y=1.145 $X2=0 $Y2=0
cc_346 N_A_161_446#_c_342_n N_DE_c_447_n 0.00499842f $X=2.335 $Y=2.035 $X2=0
+ $Y2=0
cc_347 N_A_161_446#_c_334_n N_DE_c_443_n 0.00983398f $X=1.825 $Y=0.645 $X2=0
+ $Y2=0
cc_348 N_A_161_446#_c_342_n N_DE_c_449_n 8.8846e-19 $X=2.335 $Y=2.035 $X2=0
+ $Y2=0
cc_349 N_A_161_446#_c_336_n N_DE_c_449_n 0.00104777f $X=2.5 $Y=1.145 $X2=0 $Y2=0
cc_350 N_A_161_446#_c_330_n DE 0.020843f $X=1.17 $Y=1.615 $X2=0 $Y2=0
cc_351 N_A_161_446#_c_331_n DE 0.00200717f $X=1.17 $Y=1.615 $X2=0 $Y2=0
cc_352 N_A_161_446#_c_332_n DE 0.0272396f $X=1.65 $Y=1.195 $X2=0 $Y2=0
cc_353 N_A_161_446#_c_339_n DE 0.0107567f $X=1.715 $Y=2.035 $X2=0 $Y2=0
cc_354 N_A_161_446#_c_342_n DE 0.00139436f $X=2.335 $Y=2.035 $X2=0 $Y2=0
cc_355 N_A_161_446#_c_335_n DE 0.0122102f $X=2.5 $Y=1.145 $X2=0 $Y2=0
cc_356 N_A_161_446#_c_336_n DE 5.17114e-19 $X=2.5 $Y=1.145 $X2=0 $Y2=0
cc_357 N_A_161_446#_c_376_p DE 0.0135702f $X=1.8 $Y=2.035 $X2=0 $Y2=0
cc_358 N_A_161_446#_M1001_g N_A_575_48#_M1002_g 0.0381333f $X=2.56 $Y=0.58 $X2=0
+ $Y2=0
cc_359 N_A_161_446#_c_342_n N_A_575_48#_c_538_n 0.00308805f $X=2.335 $Y=2.035
+ $X2=0 $Y2=0
cc_360 N_A_161_446#_c_335_n N_A_575_48#_c_532_n 0.00135452f $X=2.5 $Y=1.145
+ $X2=0 $Y2=0
cc_361 N_A_161_446#_c_335_n N_A_575_48#_c_534_n 0.00233006f $X=2.5 $Y=1.145
+ $X2=0 $Y2=0
cc_362 N_A_161_446#_c_336_n N_A_575_48#_c_534_n 0.0203846f $X=2.5 $Y=1.145 $X2=0
+ $Y2=0
cc_363 N_A_161_446#_c_342_n N_A_575_48#_c_535_n 0.00287934f $X=2.335 $Y=2.035
+ $X2=0 $Y2=0
cc_364 N_A_161_446#_c_335_n N_A_575_48#_c_535_n 0.0610738f $X=2.5 $Y=1.145 $X2=0
+ $Y2=0
cc_365 N_A_161_446#_c_336_n N_A_575_48#_c_535_n 0.00233006f $X=2.5 $Y=1.145
+ $X2=0 $Y2=0
cc_366 N_A_161_446#_c_335_n N_A_575_48#_c_536_n 0.00571351f $X=2.5 $Y=1.145
+ $X2=0 $Y2=0
cc_367 N_A_161_446#_c_336_n N_A_575_48#_c_536_n 0.0203846f $X=2.5 $Y=1.145 $X2=0
+ $Y2=0
cc_368 N_A_161_446#_c_342_n N_A_575_48#_c_550_n 2.8759e-19 $X=2.335 $Y=2.035
+ $X2=0 $Y2=0
cc_369 N_A_161_446#_c_337_n N_A_27_74#_c_1607_n 0.00177548f $X=0.895 $Y=2.465
+ $X2=0 $Y2=0
cc_370 N_A_161_446#_c_337_n N_A_27_74#_c_1608_n 0.0287627f $X=0.895 $Y=2.465
+ $X2=0 $Y2=0
cc_371 N_A_161_446#_c_339_n N_A_27_74#_c_1608_n 0.017295f $X=1.715 $Y=2.035
+ $X2=0 $Y2=0
cc_372 N_A_161_446#_c_340_n N_A_27_74#_c_1608_n 0.0258112f $X=1.335 $Y=2.035
+ $X2=0 $Y2=0
cc_373 N_A_161_446#_c_341_n N_A_27_74#_c_1608_n 0.0141449f $X=1.8 $Y=2.505 $X2=0
+ $Y2=0
cc_374 N_A_161_446#_c_337_n N_A_27_74#_c_1609_n 0.00412861f $X=0.895 $Y=2.465
+ $X2=0 $Y2=0
cc_375 N_A_161_446#_c_341_n N_A_27_74#_c_1609_n 0.0203028f $X=1.8 $Y=2.505 $X2=0
+ $Y2=0
cc_376 N_A_161_446#_M1032_s N_A_27_74#_c_1610_n 0.00467318f $X=1.655 $Y=2.3
+ $X2=0 $Y2=0
cc_377 N_A_161_446#_c_341_n N_A_27_74#_c_1610_n 0.012787f $X=1.8 $Y=2.505 $X2=0
+ $Y2=0
cc_378 N_A_161_446#_c_337_n N_A_27_74#_c_1611_n 6.5162e-19 $X=0.895 $Y=2.465
+ $X2=0 $Y2=0
cc_379 N_A_161_446#_c_341_n N_A_27_74#_c_1646_n 0.0192722f $X=1.8 $Y=2.505 $X2=0
+ $Y2=0
cc_380 N_A_161_446#_c_342_n N_A_27_74#_c_1612_n 0.0344588f $X=2.335 $Y=2.035
+ $X2=0 $Y2=0
cc_381 N_A_161_446#_c_336_n N_A_27_74#_c_1612_n 2.10848e-19 $X=2.5 $Y=1.145
+ $X2=0 $Y2=0
cc_382 N_A_161_446#_c_341_n N_A_27_74#_c_1613_n 0.0133747f $X=1.8 $Y=2.505 $X2=0
+ $Y2=0
cc_383 N_A_161_446#_c_342_n N_A_27_74#_c_1613_n 0.0139284f $X=2.335 $Y=2.035
+ $X2=0 $Y2=0
cc_384 N_A_161_446#_M1001_g N_A_27_74#_c_1605_n 0.00130006f $X=2.56 $Y=0.58
+ $X2=0 $Y2=0
cc_385 N_A_161_446#_c_337_n N_VPWR_c_1778_n 0.0114317f $X=0.895 $Y=2.465 $X2=0
+ $Y2=0
cc_386 N_A_161_446#_c_337_n N_VPWR_c_1790_n 0.00413917f $X=0.895 $Y=2.465 $X2=0
+ $Y2=0
cc_387 N_A_161_446#_c_337_n N_VPWR_c_1777_n 0.0084921f $X=0.895 $Y=2.465 $X2=0
+ $Y2=0
cc_388 N_A_161_446#_c_331_n N_VGND_c_1992_n 2.96882e-19 $X=1.17 $Y=1.615 $X2=0
+ $Y2=0
cc_389 N_A_161_446#_c_332_n N_VGND_c_1992_n 0.00473841f $X=1.65 $Y=1.195 $X2=0
+ $Y2=0
cc_390 N_A_161_446#_c_333_n N_VGND_c_1992_n 0.0152189f $X=1.335 $Y=1.195 $X2=0
+ $Y2=0
cc_391 N_A_161_446#_c_334_n N_VGND_c_1992_n 0.0223476f $X=1.825 $Y=0.645 $X2=0
+ $Y2=0
cc_392 N_A_161_446#_M1001_g N_VGND_c_1993_n 0.0119836f $X=2.56 $Y=0.58 $X2=0
+ $Y2=0
cc_393 N_A_161_446#_c_334_n N_VGND_c_1993_n 0.0132849f $X=1.825 $Y=0.645 $X2=0
+ $Y2=0
cc_394 N_A_161_446#_c_335_n N_VGND_c_1993_n 0.0144691f $X=2.5 $Y=1.145 $X2=0
+ $Y2=0
cc_395 N_A_161_446#_c_336_n N_VGND_c_1993_n 0.00116651f $X=2.5 $Y=1.145 $X2=0
+ $Y2=0
cc_396 N_A_161_446#_c_334_n N_VGND_c_2000_n 0.00901259f $X=1.825 $Y=0.645 $X2=0
+ $Y2=0
cc_397 N_A_161_446#_M1001_g N_VGND_c_2002_n 0.00413917f $X=2.56 $Y=0.58 $X2=0
+ $Y2=0
cc_398 N_A_161_446#_M1001_g N_VGND_c_2012_n 0.00817239f $X=2.56 $Y=0.58 $X2=0
+ $Y2=0
cc_399 N_A_161_446#_c_334_n N_VGND_c_2012_n 0.011672f $X=1.825 $Y=0.645 $X2=0
+ $Y2=0
cc_400 N_DE_c_446_n N_A_575_48#_c_538_n 0.0071313f $X=2.44 $Y=1.965 $X2=0 $Y2=0
cc_401 N_DE_c_449_n N_A_575_48#_c_538_n 0.0141084f $X=2.515 $Y=2.337 $X2=0 $Y2=0
cc_402 N_DE_c_448_n N_A_575_48#_c_539_n 0.0318153f $X=2.705 $Y=2.445 $X2=0 $Y2=0
cc_403 N_DE_c_446_n N_A_575_48#_c_550_n 0.00425825f $X=2.44 $Y=1.965 $X2=0 $Y2=0
cc_404 N_DE_c_441_n N_A_27_74#_c_1609_n 0.00326422f $X=2.025 $Y=2.225 $X2=0
+ $Y2=0
cc_405 N_DE_c_441_n N_A_27_74#_c_1610_n 0.0146314f $X=2.025 $Y=2.225 $X2=0 $Y2=0
cc_406 N_DE_c_448_n N_A_27_74#_c_1610_n 4.26516e-19 $X=2.705 $Y=2.445 $X2=0
+ $Y2=0
cc_407 N_DE_c_441_n N_A_27_74#_c_1646_n 0.0118088f $X=2.025 $Y=2.225 $X2=0 $Y2=0
cc_408 N_DE_c_448_n N_A_27_74#_c_1646_n 0.00281561f $X=2.705 $Y=2.445 $X2=0
+ $Y2=0
cc_409 N_DE_c_446_n N_A_27_74#_c_1612_n 7.33386e-19 $X=2.44 $Y=1.965 $X2=0 $Y2=0
cc_410 N_DE_c_448_n N_A_27_74#_c_1612_n 0.00653291f $X=2.705 $Y=2.445 $X2=0
+ $Y2=0
cc_411 N_DE_c_449_n N_A_27_74#_c_1612_n 0.0183963f $X=2.515 $Y=2.337 $X2=0 $Y2=0
cc_412 N_DE_c_441_n N_A_27_74#_c_1613_n 0.00591021f $X=2.025 $Y=2.225 $X2=0
+ $Y2=0
cc_413 N_DE_c_448_n N_A_27_74#_c_1614_n 0.00164727f $X=2.705 $Y=2.445 $X2=0
+ $Y2=0
cc_414 N_DE_c_436_n N_A_27_74#_c_1604_n 9.26873e-19 $X=1.04 $Y=0.865 $X2=0 $Y2=0
cc_415 N_DE_c_441_n N_VPWR_c_1779_n 0.00130831f $X=2.025 $Y=2.225 $X2=0 $Y2=0
cc_416 N_DE_c_448_n N_VPWR_c_1779_n 0.00943855f $X=2.705 $Y=2.445 $X2=0 $Y2=0
cc_417 N_DE_c_449_n N_VPWR_c_1779_n 0.00101617f $X=2.515 $Y=2.337 $X2=0 $Y2=0
cc_418 N_DE_c_448_n N_VPWR_c_1786_n 0.00505726f $X=2.705 $Y=2.445 $X2=0 $Y2=0
cc_419 N_DE_c_441_n N_VPWR_c_1791_n 9.78406e-19 $X=2.025 $Y=2.225 $X2=0 $Y2=0
cc_420 N_DE_c_448_n N_VPWR_c_1777_n 0.00489105f $X=2.705 $Y=2.445 $X2=0 $Y2=0
cc_421 N_DE_c_436_n N_VGND_c_1992_n 0.0141921f $X=1.04 $Y=0.865 $X2=0 $Y2=0
cc_422 N_DE_c_437_n N_VGND_c_1992_n 0.00547656f $X=1.575 $Y=0.94 $X2=0 $Y2=0
cc_423 N_DE_c_442_n N_VGND_c_1992_n 0.00616359f $X=2.05 $Y=0.865 $X2=0 $Y2=0
cc_424 N_DE_c_442_n N_VGND_c_1993_n 0.00606571f $X=2.05 $Y=0.865 $X2=0 $Y2=0
cc_425 N_DE_c_442_n N_VGND_c_2000_n 0.00436952f $X=2.05 $Y=0.865 $X2=0 $Y2=0
cc_426 N_DE_c_436_n N_VGND_c_2006_n 0.00383152f $X=1.04 $Y=0.865 $X2=0 $Y2=0
cc_427 N_DE_c_436_n N_VGND_c_2012_n 0.0075725f $X=1.04 $Y=0.865 $X2=0 $Y2=0
cc_428 N_DE_c_437_n N_VGND_c_2012_n 0.00504243f $X=1.575 $Y=0.94 $X2=0 $Y2=0
cc_429 N_DE_c_442_n N_VGND_c_2012_n 0.00829055f $X=2.05 $Y=0.865 $X2=0 $Y2=0
cc_430 N_A_575_48#_c_531_n N_CLK_c_755_n 0.0084639f $X=12.095 $Y=1.665 $X2=0
+ $Y2=0
cc_431 N_A_575_48#_c_536_n N_CLK_c_755_n 0.00571255f $X=3.04 $Y=1.825 $X2=0
+ $Y2=0
cc_432 N_A_575_48#_c_531_n CLK 0.0294885f $X=12.095 $Y=1.665 $X2=0 $Y2=0
cc_433 N_A_575_48#_c_551_n N_A_1008_74#_c_814_n 0.0120634f $X=11.45 $Y=1.932
+ $X2=0 $Y2=0
cc_434 N_A_575_48#_c_540_n N_A_1008_74#_c_815_n 0.022408f $X=11.435 $Y=2.14
+ $X2=0 $Y2=0
cc_435 N_A_575_48#_c_531_n N_A_1008_74#_c_790_n 0.00473892f $X=12.095 $Y=1.665
+ $X2=0 $Y2=0
cc_436 N_A_575_48#_c_531_n N_A_1008_74#_c_816_n 0.0148879f $X=12.095 $Y=1.665
+ $X2=0 $Y2=0
cc_437 N_A_575_48#_c_531_n N_A_1008_74#_c_793_n 0.0227516f $X=12.095 $Y=1.665
+ $X2=0 $Y2=0
cc_438 N_A_575_48#_c_531_n N_A_1008_74#_c_796_n 0.00776037f $X=12.095 $Y=1.665
+ $X2=0 $Y2=0
cc_439 N_A_575_48#_M1010_g N_A_1008_74#_c_801_n 3.28735e-19 $X=11.45 $Y=0.8
+ $X2=0 $Y2=0
cc_440 N_A_575_48#_c_531_n N_A_1008_74#_c_801_n 0.0150995f $X=12.095 $Y=1.665
+ $X2=0 $Y2=0
cc_441 N_A_575_48#_M1010_g N_A_1008_74#_c_802_n 0.00140735f $X=11.45 $Y=0.8
+ $X2=0 $Y2=0
cc_442 N_A_575_48#_c_531_n N_A_1008_74#_c_802_n 0.0168925f $X=12.095 $Y=1.665
+ $X2=0 $Y2=0
cc_443 N_A_575_48#_M1010_g N_A_1008_74#_c_803_n 0.0211981f $X=11.45 $Y=0.8 $X2=0
+ $Y2=0
cc_444 N_A_575_48#_c_531_n N_A_1008_74#_c_803_n 0.00348186f $X=12.095 $Y=1.665
+ $X2=0 $Y2=0
cc_445 N_A_575_48#_c_531_n N_A_1008_74#_c_820_n 0.00865386f $X=12.095 $Y=1.665
+ $X2=0 $Y2=0
cc_446 N_A_575_48#_c_531_n N_A_1008_74#_c_821_n 0.00144307f $X=12.095 $Y=1.665
+ $X2=0 $Y2=0
cc_447 N_A_575_48#_c_531_n N_A_1008_74#_c_805_n 0.00492255f $X=12.095 $Y=1.665
+ $X2=0 $Y2=0
cc_448 N_A_575_48#_c_531_n N_A_1008_74#_c_807_n 0.00711803f $X=12.095 $Y=1.665
+ $X2=0 $Y2=0
cc_449 N_A_575_48#_c_531_n N_A_1008_74#_c_808_n 0.0240931f $X=12.095 $Y=1.665
+ $X2=0 $Y2=0
cc_450 N_A_575_48#_c_531_n N_A_1008_74#_c_810_n 0.00477986f $X=12.095 $Y=1.665
+ $X2=0 $Y2=0
cc_451 N_A_575_48#_c_531_n N_A_818_74#_M1030_g 0.00647453f $X=12.095 $Y=1.665
+ $X2=0 $Y2=0
cc_452 N_A_575_48#_c_531_n N_A_818_74#_c_1012_n 0.00421726f $X=12.095 $Y=1.665
+ $X2=0 $Y2=0
cc_453 N_A_575_48#_c_531_n N_A_818_74#_c_1013_n 0.00498592f $X=12.095 $Y=1.665
+ $X2=0 $Y2=0
cc_454 N_A_575_48#_c_531_n N_A_818_74#_M1033_g 0.00491125f $X=12.095 $Y=1.665
+ $X2=0 $Y2=0
cc_455 N_A_575_48#_c_531_n N_A_818_74#_c_1015_n 0.00839201f $X=12.095 $Y=1.665
+ $X2=0 $Y2=0
cc_456 N_A_575_48#_c_531_n N_A_818_74#_c_1016_n 0.00112103f $X=12.095 $Y=1.665
+ $X2=0 $Y2=0
cc_457 N_A_575_48#_M1010_g N_A_818_74#_c_1020_n 0.0429112f $X=11.45 $Y=0.8 $X2=0
+ $Y2=0
cc_458 N_A_575_48#_c_531_n N_A_818_74#_c_1021_n 0.00375469f $X=12.095 $Y=1.665
+ $X2=0 $Y2=0
cc_459 N_A_575_48#_c_531_n N_A_818_74#_c_1022_n 9.11224e-19 $X=12.095 $Y=1.665
+ $X2=0 $Y2=0
cc_460 N_A_575_48#_c_531_n N_A_818_74#_c_1039_n 0.0157017f $X=12.095 $Y=1.665
+ $X2=0 $Y2=0
cc_461 N_A_575_48#_c_531_n N_A_818_74#_c_1024_n 0.015538f $X=12.095 $Y=1.665
+ $X2=0 $Y2=0
cc_462 N_A_575_48#_c_531_n N_A_818_74#_c_1025_n 0.0522165f $X=12.095 $Y=1.665
+ $X2=0 $Y2=0
cc_463 N_A_575_48#_c_531_n N_A_818_74#_c_1026_n 0.0129744f $X=12.095 $Y=1.665
+ $X2=0 $Y2=0
cc_464 N_A_575_48#_c_531_n N_A_818_74#_c_1027_n 0.00606193f $X=12.095 $Y=1.665
+ $X2=0 $Y2=0
cc_465 N_A_575_48#_c_531_n N_A_818_74#_c_1046_n 0.0124468f $X=12.095 $Y=1.665
+ $X2=0 $Y2=0
cc_466 N_A_575_48#_c_531_n N_A_818_74#_c_1028_n 0.0202139f $X=12.095 $Y=1.665
+ $X2=0 $Y2=0
cc_467 N_A_575_48#_c_531_n N_A_818_74#_c_1029_n 0.00533349f $X=12.095 $Y=1.665
+ $X2=0 $Y2=0
cc_468 N_A_575_48#_c_531_n N_A_1419_71#_c_1232_n 0.00434855f $X=12.095 $Y=1.665
+ $X2=0 $Y2=0
cc_469 N_A_575_48#_c_531_n N_A_1419_71#_c_1244_n 0.0053233f $X=12.095 $Y=1.665
+ $X2=0 $Y2=0
cc_470 N_A_575_48#_c_531_n N_A_1419_71#_c_1234_n 0.0118963f $X=12.095 $Y=1.665
+ $X2=0 $Y2=0
cc_471 N_A_575_48#_c_531_n N_A_1419_71#_c_1236_n 0.0177048f $X=12.095 $Y=1.665
+ $X2=0 $Y2=0
cc_472 N_A_575_48#_c_531_n N_A_1419_71#_c_1246_n 0.0110986f $X=12.095 $Y=1.665
+ $X2=0 $Y2=0
cc_473 N_A_575_48#_c_531_n N_A_1419_71#_c_1237_n 0.0331142f $X=12.095 $Y=1.665
+ $X2=0 $Y2=0
cc_474 N_A_575_48#_c_531_n N_A_1419_71#_c_1238_n 0.00394392f $X=12.095 $Y=1.665
+ $X2=0 $Y2=0
cc_475 N_A_575_48#_c_531_n N_A_1419_71#_c_1239_n 0.00841858f $X=12.095 $Y=1.665
+ $X2=0 $Y2=0
cc_476 N_A_575_48#_c_531_n N_A_1419_71#_c_1240_n 0.00851964f $X=12.095 $Y=1.665
+ $X2=0 $Y2=0
cc_477 N_A_575_48#_c_531_n N_A_1419_71#_c_1241_n 0.00428037f $X=12.095 $Y=1.665
+ $X2=0 $Y2=0
cc_478 N_A_575_48#_c_531_n N_A_1198_97#_c_1369_n 0.00167144f $X=12.095 $Y=1.665
+ $X2=0 $Y2=0
cc_479 N_A_575_48#_c_531_n N_A_1198_97#_c_1370_n 0.00321521f $X=12.095 $Y=1.665
+ $X2=0 $Y2=0
cc_480 N_A_575_48#_c_531_n N_A_1198_97#_c_1373_n 0.0348086f $X=12.095 $Y=1.665
+ $X2=0 $Y2=0
cc_481 N_A_575_48#_c_531_n N_A_1198_97#_c_1374_n 0.0225732f $X=12.095 $Y=1.665
+ $X2=0 $Y2=0
cc_482 N_A_575_48#_c_531_n N_A_1198_97#_c_1379_n 0.0400145f $X=12.095 $Y=1.665
+ $X2=0 $Y2=0
cc_483 N_A_575_48#_M1010_g N_A_1879_74#_M1015_g 0.0108721f $X=11.45 $Y=0.8 $X2=0
+ $Y2=0
cc_484 N_A_575_48#_c_527_n N_A_1879_74#_M1015_g 0.00469864f $X=12.485 $Y=0.34
+ $X2=0 $Y2=0
cc_485 N_A_575_48#_c_537_n N_A_1879_74#_M1015_g 0.0123833f $X=12.32 $Y=0.515
+ $X2=0 $Y2=0
cc_486 N_A_575_48#_c_544_n N_A_1879_74#_c_1480_n 0.0141345f $X=12.615 $Y=2.68
+ $X2=0 $Y2=0
cc_487 N_A_575_48#_c_545_n N_A_1879_74#_c_1480_n 0.0196882f $X=12.615 $Y=1.97
+ $X2=0 $Y2=0
cc_488 N_A_575_48#_c_551_n N_A_1879_74#_c_1480_n 0.0077221f $X=11.45 $Y=1.932
+ $X2=0 $Y2=0
cc_489 N_A_575_48#_c_545_n N_A_1879_74#_c_1471_n 0.00504868f $X=12.615 $Y=1.97
+ $X2=0 $Y2=0
cc_490 N_A_575_48#_c_537_n N_A_1879_74#_c_1471_n 0.00746162f $X=12.32 $Y=0.515
+ $X2=0 $Y2=0
cc_491 N_A_575_48#_M1010_g N_A_1879_74#_c_1472_n 0.0258147f $X=11.45 $Y=0.8
+ $X2=0 $Y2=0
cc_492 N_A_575_48#_c_543_n N_A_1879_74#_c_1472_n 0.00903431f $X=12.155 $Y=1.922
+ $X2=0 $Y2=0
cc_493 N_A_575_48#_c_545_n N_A_1879_74#_c_1472_n 0.00486269f $X=12.615 $Y=1.97
+ $X2=0 $Y2=0
cc_494 N_A_575_48#_c_531_n N_A_1879_74#_c_1472_n 0.00744831f $X=12.095 $Y=1.665
+ $X2=0 $Y2=0
cc_495 N_A_575_48#_c_533_n N_A_1879_74#_c_1472_n 0.0038221f $X=12.24 $Y=1.665
+ $X2=0 $Y2=0
cc_496 N_A_575_48#_c_551_n N_A_1879_74#_c_1472_n 0.00999405f $X=11.45 $Y=1.932
+ $X2=0 $Y2=0
cc_497 N_A_575_48#_c_537_n N_A_1879_74#_c_1472_n 0.0364398f $X=12.32 $Y=0.515
+ $X2=0 $Y2=0
cc_498 N_A_575_48#_M1022_g N_A_1879_74#_c_1473_n 0.00650398f $X=13.905 $Y=0.76
+ $X2=0 $Y2=0
cc_499 N_A_575_48#_c_526_n N_A_1879_74#_c_1473_n 0.0166368f $X=13.265 $Y=0.34
+ $X2=0 $Y2=0
cc_500 N_A_575_48#_c_528_n N_A_1879_74#_c_1473_n 0.00656217f $X=13.35 $Y=1.32
+ $X2=0 $Y2=0
cc_501 N_A_575_48#_c_537_n N_A_1879_74#_c_1473_n 0.00634877f $X=12.32 $Y=0.515
+ $X2=0 $Y2=0
cc_502 N_A_575_48#_c_524_n N_A_1879_74#_c_1474_n 0.00549255f $X=13.85 $Y=1.765
+ $X2=0 $Y2=0
cc_503 N_A_575_48#_c_529_n N_A_1879_74#_c_1474_n 0.0088824f $X=13.435 $Y=1.485
+ $X2=0 $Y2=0
cc_504 N_A_575_48#_c_530_n N_A_1879_74#_c_1474_n 0.00434907f $X=13.865 $Y=1.485
+ $X2=0 $Y2=0
cc_505 N_A_575_48#_c_524_n N_A_1879_74#_c_1483_n 0.00972181f $X=13.85 $Y=1.765
+ $X2=0 $Y2=0
cc_506 N_A_575_48#_c_544_n N_A_1879_74#_c_1483_n 0.00109027f $X=12.615 $Y=2.68
+ $X2=0 $Y2=0
cc_507 N_A_575_48#_c_545_n N_A_1879_74#_c_1483_n 5.62715e-19 $X=12.615 $Y=1.97
+ $X2=0 $Y2=0
cc_508 N_A_575_48#_c_524_n N_A_1879_74#_c_1475_n 0.0214196f $X=13.85 $Y=1.765
+ $X2=0 $Y2=0
cc_509 N_A_575_48#_M1022_g N_A_1879_74#_c_1475_n 0.00432226f $X=13.905 $Y=0.76
+ $X2=0 $Y2=0
cc_510 N_A_575_48#_c_528_n N_A_1879_74#_c_1475_n 0.00922811f $X=13.35 $Y=1.32
+ $X2=0 $Y2=0
cc_511 N_A_575_48#_c_529_n N_A_1879_74#_c_1475_n 0.00593902f $X=13.435 $Y=1.485
+ $X2=0 $Y2=0
cc_512 N_A_575_48#_c_530_n N_A_1879_74#_c_1475_n 0.00498348f $X=13.865 $Y=1.485
+ $X2=0 $Y2=0
cc_513 N_A_575_48#_M1010_g N_A_1879_74#_c_1518_n 0.009371f $X=11.45 $Y=0.8 $X2=0
+ $Y2=0
cc_514 N_A_575_48#_c_531_n N_A_1879_74#_c_1484_n 0.00865863f $X=12.095 $Y=1.665
+ $X2=0 $Y2=0
cc_515 N_A_575_48#_c_540_n N_A_1879_74#_c_1486_n 0.00513045f $X=11.435 $Y=2.14
+ $X2=0 $Y2=0
cc_516 N_A_575_48#_c_543_n N_A_1879_74#_c_1486_n 0.0116309f $X=12.155 $Y=1.922
+ $X2=0 $Y2=0
cc_517 N_A_575_48#_c_531_n N_A_1879_74#_c_1486_n 0.0111042f $X=12.095 $Y=1.665
+ $X2=0 $Y2=0
cc_518 N_A_575_48#_c_551_n N_A_1879_74#_c_1486_n 0.00597696f $X=11.45 $Y=1.932
+ $X2=0 $Y2=0
cc_519 N_A_575_48#_M1010_g N_A_1879_74#_c_1476_n 0.00552175f $X=11.45 $Y=0.8
+ $X2=0 $Y2=0
cc_520 N_A_575_48#_M1010_g N_A_1879_74#_c_1477_n 0.00696667f $X=11.45 $Y=0.8
+ $X2=0 $Y2=0
cc_521 N_A_575_48#_c_543_n N_A_1879_74#_c_1477_n 0.0196011f $X=12.155 $Y=1.922
+ $X2=0 $Y2=0
cc_522 N_A_575_48#_c_531_n N_A_1879_74#_c_1477_n 0.0242989f $X=12.095 $Y=1.665
+ $X2=0 $Y2=0
cc_523 N_A_575_48#_c_551_n N_A_1879_74#_c_1477_n 0.0067904f $X=11.45 $Y=1.932
+ $X2=0 $Y2=0
cc_524 N_A_575_48#_M1010_g N_A_1879_74#_c_1478_n 0.010409f $X=11.45 $Y=0.8 $X2=0
+ $Y2=0
cc_525 N_A_575_48#_c_543_n N_A_1879_74#_c_1478_n 0.0159788f $X=12.155 $Y=1.922
+ $X2=0 $Y2=0
cc_526 N_A_575_48#_c_531_n N_A_1879_74#_c_1478_n 0.0186353f $X=12.095 $Y=1.665
+ $X2=0 $Y2=0
cc_527 N_A_575_48#_c_551_n N_A_1879_74#_c_1478_n 0.00523376f $X=11.45 $Y=1.932
+ $X2=0 $Y2=0
cc_528 N_A_575_48#_c_537_n N_A_1879_74#_c_1478_n 0.0262736f $X=12.32 $Y=0.515
+ $X2=0 $Y2=0
cc_529 N_A_575_48#_M1010_g N_A_1879_74#_c_1479_n 0.00618996f $X=11.45 $Y=0.8
+ $X2=0 $Y2=0
cc_530 N_A_575_48#_c_538_n N_A_27_74#_c_1612_n 0.00419061f $X=3.095 $Y=2.355
+ $X2=0 $Y2=0
cc_531 N_A_575_48#_c_539_n N_A_27_74#_c_1612_n 0.00827774f $X=3.095 $Y=2.445
+ $X2=0 $Y2=0
cc_532 N_A_575_48#_c_532_n N_A_27_74#_c_1612_n 7.91426e-19 $X=3.265 $Y=1.665
+ $X2=0 $Y2=0
cc_533 N_A_575_48#_c_535_n N_A_27_74#_c_1612_n 0.0130849f $X=3.04 $Y=1.145 $X2=0
+ $Y2=0
cc_534 N_A_575_48#_c_550_n N_A_27_74#_c_1612_n 7.98038e-19 $X=3.04 $Y=1.99 $X2=0
+ $Y2=0
cc_535 N_A_575_48#_c_539_n N_A_27_74#_c_1614_n 0.00996615f $X=3.095 $Y=2.445
+ $X2=0 $Y2=0
cc_536 N_A_575_48#_M1002_g N_A_27_74#_c_1600_n 0.00479218f $X=2.95 $Y=0.58 $X2=0
+ $Y2=0
cc_537 N_A_575_48#_c_538_n N_A_27_74#_c_1600_n 0.0102283f $X=3.095 $Y=2.355
+ $X2=0 $Y2=0
cc_538 N_A_575_48#_c_531_n N_A_27_74#_c_1600_n 0.0267718f $X=12.095 $Y=1.665
+ $X2=0 $Y2=0
cc_539 N_A_575_48#_c_532_n N_A_27_74#_c_1600_n 0.00275409f $X=3.265 $Y=1.665
+ $X2=0 $Y2=0
cc_540 N_A_575_48#_c_534_n N_A_27_74#_c_1600_n 0.0168272f $X=3.04 $Y=1.145 $X2=0
+ $Y2=0
cc_541 N_A_575_48#_c_535_n N_A_27_74#_c_1600_n 0.0736675f $X=3.04 $Y=1.145 $X2=0
+ $Y2=0
cc_542 N_A_575_48#_c_531_n N_A_27_74#_c_1616_n 0.0260272f $X=12.095 $Y=1.665
+ $X2=0 $Y2=0
cc_543 N_A_575_48#_c_531_n N_A_27_74#_c_1601_n 0.0192983f $X=12.095 $Y=1.665
+ $X2=0 $Y2=0
cc_544 N_A_575_48#_c_531_n N_A_27_74#_c_1677_n 0.0042797f $X=12.095 $Y=1.665
+ $X2=0 $Y2=0
cc_545 N_A_575_48#_c_531_n N_A_27_74#_c_1602_n 0.0158725f $X=12.095 $Y=1.665
+ $X2=0 $Y2=0
cc_546 N_A_575_48#_M1002_g N_A_27_74#_c_1605_n 0.00984716f $X=2.95 $Y=0.58 $X2=0
+ $Y2=0
cc_547 N_A_575_48#_c_534_n N_A_27_74#_c_1605_n 0.00134541f $X=3.04 $Y=1.145
+ $X2=0 $Y2=0
cc_548 N_A_575_48#_c_535_n N_A_27_74#_c_1605_n 0.0174507f $X=3.04 $Y=1.145 $X2=0
+ $Y2=0
cc_549 N_A_575_48#_c_538_n N_A_27_74#_c_1621_n 0.00223164f $X=3.095 $Y=2.355
+ $X2=0 $Y2=0
cc_550 N_A_575_48#_c_539_n N_A_27_74#_c_1621_n 0.00398191f $X=3.095 $Y=2.445
+ $X2=0 $Y2=0
cc_551 N_A_575_48#_c_531_n N_A_27_74#_c_1621_n 0.00400047f $X=12.095 $Y=1.665
+ $X2=0 $Y2=0
cc_552 N_A_575_48#_c_532_n N_A_27_74#_c_1621_n 0.00266129f $X=3.265 $Y=1.665
+ $X2=0 $Y2=0
cc_553 N_A_575_48#_c_535_n N_A_27_74#_c_1621_n 0.00240844f $X=3.04 $Y=1.145
+ $X2=0 $Y2=0
cc_554 N_A_575_48#_c_543_n N_VPWR_M1009_d 0.00192414f $X=12.155 $Y=1.922 $X2=0
+ $Y2=0
cc_555 N_A_575_48#_c_545_n N_VPWR_M1009_d 0.00123657f $X=12.615 $Y=1.97 $X2=0
+ $Y2=0
cc_556 N_A_575_48#_c_539_n N_VPWR_c_1779_n 0.00146278f $X=3.095 $Y=2.445 $X2=0
+ $Y2=0
cc_557 N_A_575_48#_c_539_n N_VPWR_c_1780_n 0.00323308f $X=3.095 $Y=2.445 $X2=0
+ $Y2=0
cc_558 N_A_575_48#_c_531_n N_VPWR_c_1783_n 0.00246007f $X=12.095 $Y=1.665 $X2=0
+ $Y2=0
cc_559 N_A_575_48#_c_540_n N_VPWR_c_1784_n 0.0125155f $X=11.435 $Y=2.14 $X2=0
+ $Y2=0
cc_560 N_A_575_48#_c_543_n N_VPWR_c_1784_n 0.039418f $X=12.155 $Y=1.922 $X2=0
+ $Y2=0
cc_561 N_A_575_48#_c_544_n N_VPWR_c_1784_n 0.019581f $X=12.615 $Y=2.68 $X2=0
+ $Y2=0
cc_562 N_A_575_48#_c_545_n N_VPWR_c_1784_n 0.0076895f $X=12.615 $Y=1.97 $X2=0
+ $Y2=0
cc_563 N_A_575_48#_c_531_n N_VPWR_c_1784_n 0.0057493f $X=12.095 $Y=1.665 $X2=0
+ $Y2=0
cc_564 N_A_575_48#_c_533_n N_VPWR_c_1784_n 8.11221e-19 $X=12.24 $Y=1.665 $X2=0
+ $Y2=0
cc_565 N_A_575_48#_c_551_n N_VPWR_c_1784_n 0.00450667f $X=11.45 $Y=1.932 $X2=0
+ $Y2=0
cc_566 N_A_575_48#_c_524_n N_VPWR_c_1785_n 0.0211476f $X=13.85 $Y=1.765 $X2=0
+ $Y2=0
cc_567 N_A_575_48#_c_530_n N_VPWR_c_1785_n 0.0215077f $X=13.865 $Y=1.485 $X2=0
+ $Y2=0
cc_568 N_A_575_48#_c_539_n N_VPWR_c_1786_n 0.00548284f $X=3.095 $Y=2.445 $X2=0
+ $Y2=0
cc_569 N_A_575_48#_c_540_n N_VPWR_c_1794_n 0.00341451f $X=11.435 $Y=2.14 $X2=0
+ $Y2=0
cc_570 N_A_575_48#_c_544_n N_VPWR_c_1795_n 0.00710092f $X=12.615 $Y=2.68 $X2=0
+ $Y2=0
cc_571 N_A_575_48#_c_524_n N_VPWR_c_1796_n 0.00413917f $X=13.85 $Y=1.765 $X2=0
+ $Y2=0
cc_572 N_A_575_48#_c_539_n N_VPWR_c_1777_n 0.00539454f $X=3.095 $Y=2.445 $X2=0
+ $Y2=0
cc_573 N_A_575_48#_c_540_n N_VPWR_c_1777_n 0.00408462f $X=11.435 $Y=2.14 $X2=0
+ $Y2=0
cc_574 N_A_575_48#_c_524_n N_VPWR_c_1777_n 0.00821361f $X=13.85 $Y=1.765 $X2=0
+ $Y2=0
cc_575 N_A_575_48#_c_544_n N_VPWR_c_1777_n 0.00836989f $X=12.615 $Y=2.68 $X2=0
+ $Y2=0
cc_576 N_A_575_48#_c_526_n N_Q_M1017_s 0.00276743f $X=13.265 $Y=0.34 $X2=-0.19
+ $Y2=-0.245
cc_577 N_A_575_48#_c_526_n N_Q_c_1939_n 0.017778f $X=13.265 $Y=0.34 $X2=0 $Y2=0
cc_578 N_A_575_48#_c_528_n N_Q_c_1939_n 0.0316832f $X=13.35 $Y=1.32 $X2=0 $Y2=0
cc_579 N_A_575_48#_c_537_n N_Q_c_1939_n 0.022375f $X=12.32 $Y=0.515 $X2=0 $Y2=0
cc_580 N_A_575_48#_c_524_n Q 3.90495e-19 $X=13.85 $Y=1.765 $X2=0 $Y2=0
cc_581 N_A_575_48#_c_529_n Q 0.00673864f $X=13.435 $Y=1.485 $X2=0 $Y2=0
cc_582 N_A_575_48#_c_544_n Q 0.048365f $X=12.615 $Y=2.68 $X2=0 $Y2=0
cc_583 N_A_575_48#_c_529_n N_Q_c_1940_n 0.0263493f $X=13.435 $Y=1.485 $X2=0
+ $Y2=0
cc_584 N_A_575_48#_c_545_n N_Q_c_1940_n 0.0257104f $X=12.615 $Y=1.97 $X2=0 $Y2=0
cc_585 N_A_575_48#_c_533_n N_Q_c_1940_n 0.00128995f $X=12.24 $Y=1.665 $X2=0
+ $Y2=0
cc_586 N_A_575_48#_c_537_n N_Q_c_1940_n 0.025921f $X=12.32 $Y=0.515 $X2=0 $Y2=0
cc_587 N_A_575_48#_c_524_n N_Q_N_c_1975_n 0.00712539f $X=13.85 $Y=1.765 $X2=0
+ $Y2=0
cc_588 N_A_575_48#_c_524_n N_Q_N_c_1972_n 0.0119393f $X=13.85 $Y=1.765 $X2=0
+ $Y2=0
cc_589 N_A_575_48#_M1022_g N_Q_N_c_1972_n 0.00411368f $X=13.905 $Y=0.76 $X2=0
+ $Y2=0
cc_590 N_A_575_48#_c_530_n N_Q_N_c_1972_n 0.0263017f $X=13.865 $Y=1.485 $X2=0
+ $Y2=0
cc_591 N_A_575_48#_M1022_g Q_N 0.00842121f $X=13.905 $Y=0.76 $X2=0 $Y2=0
cc_592 N_A_575_48#_c_524_n Q_N 0.00166529f $X=13.85 $Y=1.765 $X2=0 $Y2=0
cc_593 N_A_575_48#_M1022_g Q_N 0.00287735f $X=13.905 $Y=0.76 $X2=0 $Y2=0
cc_594 N_A_575_48#_c_530_n Q_N 0.00151667f $X=13.865 $Y=1.485 $X2=0 $Y2=0
cc_595 N_A_575_48#_c_526_n N_VGND_M1017_d 4.00445e-19 $X=13.265 $Y=0.34 $X2=0
+ $Y2=0
cc_596 N_A_575_48#_c_528_n N_VGND_M1017_d 0.0104218f $X=13.35 $Y=1.32 $X2=0
+ $Y2=0
cc_597 N_A_575_48#_M1002_g N_VGND_c_1993_n 0.00183544f $X=2.95 $Y=0.58 $X2=0
+ $Y2=0
cc_598 N_A_575_48#_M1002_g N_VGND_c_1994_n 0.00286169f $X=2.95 $Y=0.58 $X2=0
+ $Y2=0
cc_599 N_A_575_48#_M1010_g N_VGND_c_1998_n 0.00773308f $X=11.45 $Y=0.8 $X2=0
+ $Y2=0
cc_600 N_A_575_48#_c_527_n N_VGND_c_1998_n 0.011924f $X=12.485 $Y=0.34 $X2=0
+ $Y2=0
cc_601 N_A_575_48#_c_524_n N_VGND_c_1999_n 0.00174389f $X=13.85 $Y=1.765 $X2=0
+ $Y2=0
cc_602 N_A_575_48#_M1022_g N_VGND_c_1999_n 0.00395306f $X=13.905 $Y=0.76 $X2=0
+ $Y2=0
cc_603 N_A_575_48#_c_526_n N_VGND_c_1999_n 0.0142491f $X=13.265 $Y=0.34 $X2=0
+ $Y2=0
cc_604 N_A_575_48#_c_528_n N_VGND_c_1999_n 0.0526759f $X=13.35 $Y=1.32 $X2=0
+ $Y2=0
cc_605 N_A_575_48#_c_530_n N_VGND_c_1999_n 0.0145561f $X=13.865 $Y=1.485 $X2=0
+ $Y2=0
cc_606 N_A_575_48#_M1002_g N_VGND_c_2002_n 0.00433162f $X=2.95 $Y=0.58 $X2=0
+ $Y2=0
cc_607 N_A_575_48#_M1010_g N_VGND_c_2009_n 0.00387406f $X=11.45 $Y=0.8 $X2=0
+ $Y2=0
cc_608 N_A_575_48#_c_526_n N_VGND_c_2010_n 0.0623747f $X=13.265 $Y=0.34 $X2=0
+ $Y2=0
cc_609 N_A_575_48#_c_527_n N_VGND_c_2010_n 0.0235688f $X=12.485 $Y=0.34 $X2=0
+ $Y2=0
cc_610 N_A_575_48#_M1022_g N_VGND_c_2011_n 0.00537471f $X=13.905 $Y=0.76 $X2=0
+ $Y2=0
cc_611 N_A_575_48#_M1002_g N_VGND_c_2012_n 0.00822327f $X=2.95 $Y=0.58 $X2=0
+ $Y2=0
cc_612 N_A_575_48#_M1010_g N_VGND_c_2012_n 0.00479212f $X=11.45 $Y=0.8 $X2=0
+ $Y2=0
cc_613 N_A_575_48#_M1022_g N_VGND_c_2012_n 0.00539454f $X=13.905 $Y=0.76 $X2=0
+ $Y2=0
cc_614 N_A_575_48#_c_526_n N_VGND_c_2012_n 0.0359274f $X=13.265 $Y=0.34 $X2=0
+ $Y2=0
cc_615 N_A_575_48#_c_527_n N_VGND_c_2012_n 0.0127152f $X=12.485 $Y=0.34 $X2=0
+ $Y2=0
cc_616 N_CLK_c_755_n N_A_818_74#_M1030_g 0.00605661f $X=4.105 $Y=1.765 $X2=0
+ $Y2=0
cc_617 N_CLK_c_754_n N_A_818_74#_c_1023_n 0.00602343f $X=4.015 $Y=1.22 $X2=0
+ $Y2=0
cc_618 N_CLK_c_755_n N_A_818_74#_c_1039_n 0.00946936f $X=4.105 $Y=1.765 $X2=0
+ $Y2=0
cc_619 CLK N_A_818_74#_c_1039_n 0.00802062f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_620 N_CLK_c_754_n N_A_818_74#_c_1024_n 0.00342331f $X=4.015 $Y=1.22 $X2=0
+ $Y2=0
cc_621 N_CLK_c_755_n N_A_818_74#_c_1024_n 0.00721579f $X=4.105 $Y=1.765 $X2=0
+ $Y2=0
cc_622 CLK N_A_818_74#_c_1024_n 0.0295765f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_623 N_CLK_c_754_n N_A_818_74#_c_1027_n 0.00230062f $X=4.015 $Y=1.22 $X2=0
+ $Y2=0
cc_624 N_CLK_c_755_n N_A_818_74#_c_1027_n 0.00173018f $X=4.105 $Y=1.765 $X2=0
+ $Y2=0
cc_625 CLK N_A_818_74#_c_1027_n 0.0224944f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_626 N_CLK_c_755_n N_A_818_74#_c_1029_n 0.00927936f $X=4.105 $Y=1.765 $X2=0
+ $Y2=0
cc_627 N_CLK_c_755_n N_A_27_74#_c_1614_n 0.00424734f $X=4.105 $Y=1.765 $X2=0
+ $Y2=0
cc_628 N_CLK_c_754_n N_A_27_74#_c_1600_n 0.004641f $X=4.015 $Y=1.22 $X2=0 $Y2=0
cc_629 N_CLK_c_755_n N_A_27_74#_c_1600_n 0.017565f $X=4.105 $Y=1.765 $X2=0 $Y2=0
cc_630 CLK N_A_27_74#_c_1600_n 0.0295764f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_631 N_CLK_c_755_n N_A_27_74#_c_1616_n 0.0172284f $X=4.105 $Y=1.765 $X2=0
+ $Y2=0
cc_632 N_CLK_c_755_n N_A_27_74#_c_1621_n 5.90574e-19 $X=4.105 $Y=1.765 $X2=0
+ $Y2=0
cc_633 N_CLK_c_755_n N_VPWR_c_1780_n 0.0217145f $X=4.105 $Y=1.765 $X2=0 $Y2=0
cc_634 N_CLK_c_755_n N_VPWR_c_1788_n 0.00413917f $X=4.105 $Y=1.765 $X2=0 $Y2=0
cc_635 N_CLK_c_755_n N_VPWR_c_1777_n 0.00421563f $X=4.105 $Y=1.765 $X2=0 $Y2=0
cc_636 N_CLK_c_754_n N_VGND_c_1994_n 0.00467989f $X=4.015 $Y=1.22 $X2=0 $Y2=0
cc_637 N_CLK_c_755_n N_VGND_c_1994_n 0.0011901f $X=4.105 $Y=1.765 $X2=0 $Y2=0
cc_638 CLK N_VGND_c_1994_n 0.0143337f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_639 N_CLK_c_754_n N_VGND_c_1995_n 0.00339407f $X=4.015 $Y=1.22 $X2=0 $Y2=0
cc_640 N_CLK_c_754_n N_VGND_c_2004_n 0.00434272f $X=4.015 $Y=1.22 $X2=0 $Y2=0
cc_641 N_CLK_c_754_n N_VGND_c_2012_n 0.00825667f $X=4.015 $Y=1.22 $X2=0 $Y2=0
cc_642 N_A_1008_74#_c_790_n N_A_818_74#_M1030_g 0.00164702f $X=5.18 $Y=0.515
+ $X2=0 $Y2=0
cc_643 N_A_1008_74#_c_792_n N_A_818_74#_M1030_g 0.00266901f $X=5.345 $Y=0.34
+ $X2=0 $Y2=0
cc_644 N_A_1008_74#_c_790_n N_A_818_74#_c_1012_n 0.00217131f $X=5.18 $Y=0.515
+ $X2=0 $Y2=0
cc_645 N_A_1008_74#_c_816_n N_A_818_74#_c_1031_n 0.00397036f $X=5.955 $Y=1.975
+ $X2=0 $Y2=0
cc_646 N_A_1008_74#_c_793_n N_A_818_74#_c_1031_n 9.57923e-19 $X=6.04 $Y=1.81
+ $X2=0 $Y2=0
cc_647 N_A_1008_74#_c_820_n N_A_818_74#_c_1031_n 0.0015561f $X=6.155 $Y=1.975
+ $X2=0 $Y2=0
cc_648 N_A_1008_74#_c_821_n N_A_818_74#_c_1031_n 0.00653061f $X=6.19 $Y=2.215
+ $X2=0 $Y2=0
cc_649 N_A_1008_74#_c_816_n N_A_818_74#_c_1013_n 0.0119307f $X=5.955 $Y=1.975
+ $X2=0 $Y2=0
cc_650 N_A_1008_74#_c_787_n N_A_818_74#_M1033_g 0.013458f $X=6.595 $Y=1.015
+ $X2=0 $Y2=0
cc_651 N_A_1008_74#_c_790_n N_A_818_74#_M1033_g 0.00315974f $X=5.18 $Y=0.515
+ $X2=0 $Y2=0
cc_652 N_A_1008_74#_c_791_n N_A_818_74#_M1033_g 0.00929412f $X=5.955 $Y=0.34
+ $X2=0 $Y2=0
cc_653 N_A_1008_74#_c_793_n N_A_818_74#_M1033_g 0.0315253f $X=6.04 $Y=1.81 $X2=0
+ $Y2=0
cc_654 N_A_1008_74#_c_795_n N_A_818_74#_M1033_g 2.72122e-19 $X=6.76 $Y=0.965
+ $X2=0 $Y2=0
cc_655 N_A_1008_74#_c_804_n N_A_818_74#_M1033_g 0.00206916f $X=6.04 $Y=0.34
+ $X2=0 $Y2=0
cc_656 N_A_1008_74#_c_793_n N_A_818_74#_c_1015_n 0.00923398f $X=6.04 $Y=1.81
+ $X2=0 $Y2=0
cc_657 N_A_1008_74#_c_820_n N_A_818_74#_c_1015_n 0.00574057f $X=6.155 $Y=1.975
+ $X2=0 $Y2=0
cc_658 N_A_1008_74#_c_821_n N_A_818_74#_c_1015_n 0.0214798f $X=6.19 $Y=2.215
+ $X2=0 $Y2=0
cc_659 N_A_1008_74#_c_805_n N_A_818_74#_c_1015_n 3.1263e-19 $X=6.76 $Y=1.05
+ $X2=0 $Y2=0
cc_660 N_A_1008_74#_c_806_n N_A_818_74#_c_1015_n 0.0138685f $X=6.72 $Y=1.18
+ $X2=0 $Y2=0
cc_661 N_A_1008_74#_c_821_n N_A_818_74#_c_1034_n 0.00347128f $X=6.19 $Y=2.215
+ $X2=0 $Y2=0
cc_662 N_A_1008_74#_c_813_n N_A_818_74#_c_1035_n 0.00970175f $X=6.59 $Y=2.465
+ $X2=0 $Y2=0
cc_663 N_A_1008_74#_c_821_n N_A_818_74#_c_1035_n 0.0118636f $X=6.19 $Y=2.215
+ $X2=0 $Y2=0
cc_664 N_A_1008_74#_c_814_n N_A_818_74#_c_1016_n 0.0085831f $X=10.955 $Y=2.05
+ $X2=0 $Y2=0
cc_665 N_A_1008_74#_c_801_n N_A_818_74#_c_1016_n 0.00124684f $X=10.835 $Y=1.205
+ $X2=0 $Y2=0
cc_666 N_A_1008_74#_c_802_n N_A_818_74#_c_1016_n 0.00115671f $X=11 $Y=1.635
+ $X2=0 $Y2=0
cc_667 N_A_1008_74#_c_803_n N_A_818_74#_c_1016_n 0.0212691f $X=11 $Y=1.635 $X2=0
+ $Y2=0
cc_668 N_A_1008_74#_c_801_n N_A_818_74#_c_1017_n 0.00343519f $X=10.835 $Y=1.205
+ $X2=0 $Y2=0
cc_669 N_A_1008_74#_c_802_n N_A_818_74#_c_1017_n 0.00607873f $X=11 $Y=1.635
+ $X2=0 $Y2=0
cc_670 N_A_1008_74#_c_811_n N_A_818_74#_c_1017_n 9.12559e-19 $X=10.085 $Y=1.285
+ $X2=0 $Y2=0
cc_671 N_A_1008_74#_c_801_n N_A_818_74#_c_1018_n 0.0159682f $X=10.835 $Y=1.205
+ $X2=0 $Y2=0
cc_672 N_A_1008_74#_c_803_n N_A_818_74#_c_1018_n 0.0197568f $X=11 $Y=1.635 $X2=0
+ $Y2=0
cc_673 N_A_1008_74#_c_801_n N_A_818_74#_c_1019_n 0.00486996f $X=10.835 $Y=1.205
+ $X2=0 $Y2=0
cc_674 N_A_1008_74#_c_810_n N_A_818_74#_c_1019_n 0.00931461f $X=9.92 $Y=1.285
+ $X2=0 $Y2=0
cc_675 N_A_1008_74#_c_793_n N_A_818_74#_c_1022_n 0.0042578f $X=6.04 $Y=1.81
+ $X2=0 $Y2=0
cc_676 N_A_1008_74#_c_790_n N_A_818_74#_c_1024_n 0.00292736f $X=5.18 $Y=0.515
+ $X2=0 $Y2=0
cc_677 N_A_1008_74#_c_801_n N_A_818_74#_c_1025_n 0.00704471f $X=10.835 $Y=1.205
+ $X2=0 $Y2=0
cc_678 N_A_1008_74#_c_809_n N_A_818_74#_c_1025_n 0.0455289f $X=9.92 $Y=1.285
+ $X2=0 $Y2=0
cc_679 N_A_1008_74#_c_810_n N_A_818_74#_c_1025_n 0.00239497f $X=9.92 $Y=1.285
+ $X2=0 $Y2=0
cc_680 N_A_1008_74#_c_812_n N_A_818_74#_c_1025_n 7.53512e-19 $X=9.755 $Y=1.285
+ $X2=0 $Y2=0
cc_681 N_A_1008_74#_c_789_n N_A_818_74#_c_1026_n 3.83592e-19 $X=9.395 $Y=1.26
+ $X2=0 $Y2=0
cc_682 N_A_1008_74#_c_808_n N_A_818_74#_c_1026_n 0.0122499f $X=9.37 $Y=1.207
+ $X2=0 $Y2=0
cc_683 N_A_1008_74#_c_801_n N_A_818_74#_c_1028_n 0.0226331f $X=10.835 $Y=1.205
+ $X2=0 $Y2=0
cc_684 N_A_1008_74#_c_802_n N_A_818_74#_c_1028_n 0.0191189f $X=11 $Y=1.635 $X2=0
+ $Y2=0
cc_685 N_A_1008_74#_c_803_n N_A_818_74#_c_1028_n 0.00109896f $X=11 $Y=1.635
+ $X2=0 $Y2=0
cc_686 N_A_1008_74#_c_797_n N_A_1419_71#_M1014_d 0.00434104f $X=8.32 $Y=0.34
+ $X2=-0.19 $Y2=-0.245
cc_687 N_A_1008_74#_c_787_n N_A_1419_71#_M1021_g 0.015001f $X=6.595 $Y=1.015
+ $X2=0 $Y2=0
cc_688 N_A_1008_74#_c_794_n N_A_1419_71#_M1021_g 6.76761e-19 $X=6.635 $Y=0.34
+ $X2=0 $Y2=0
cc_689 N_A_1008_74#_c_795_n N_A_1419_71#_M1021_g 0.00700224f $X=6.76 $Y=0.965
+ $X2=0 $Y2=0
cc_690 N_A_1008_74#_c_796_n N_A_1419_71#_M1021_g 0.0155256f $X=7.64 $Y=1.05
+ $X2=0 $Y2=0
cc_691 N_A_1008_74#_c_889_p N_A_1419_71#_M1021_g 0.00342676f $X=7.725 $Y=0.965
+ $X2=0 $Y2=0
cc_692 N_A_1008_74#_c_805_n N_A_1419_71#_M1021_g 0.00148219f $X=6.76 $Y=1.05
+ $X2=0 $Y2=0
cc_693 N_A_1008_74#_c_806_n N_A_1419_71#_M1021_g 0.0216053f $X=6.72 $Y=1.18
+ $X2=0 $Y2=0
cc_694 N_A_1008_74#_c_788_n N_A_1419_71#_M1006_g 0.0671311f $X=9.32 $Y=1.185
+ $X2=0 $Y2=0
cc_695 N_A_1008_74#_c_797_n N_A_1419_71#_M1006_g 7.48878e-19 $X=8.32 $Y=0.34
+ $X2=0 $Y2=0
cc_696 N_A_1008_74#_c_799_n N_A_1419_71#_M1006_g 0.00498056f $X=8.405 $Y=0.965
+ $X2=0 $Y2=0
cc_697 N_A_1008_74#_c_807_n N_A_1419_71#_M1006_g 0.0157296f $X=9.2 $Y=1.207
+ $X2=0 $Y2=0
cc_698 N_A_1008_74#_c_808_n N_A_1419_71#_M1006_g 0.00593839f $X=9.37 $Y=1.207
+ $X2=0 $Y2=0
cc_699 N_A_1008_74#_c_810_n N_A_1419_71#_M1006_g 9.99083e-19 $X=9.92 $Y=1.285
+ $X2=0 $Y2=0
cc_700 N_A_1008_74#_c_789_n N_A_1419_71#_c_1244_n 0.0141167f $X=9.395 $Y=1.26
+ $X2=0 $Y2=0
cc_701 N_A_1008_74#_c_807_n N_A_1419_71#_c_1244_n 0.00297368f $X=9.2 $Y=1.207
+ $X2=0 $Y2=0
cc_702 N_A_1008_74#_c_808_n N_A_1419_71#_c_1244_n 0.00264135f $X=9.37 $Y=1.207
+ $X2=0 $Y2=0
cc_703 N_A_1008_74#_c_809_n N_A_1419_71#_c_1244_n 3.10007e-19 $X=9.92 $Y=1.285
+ $X2=0 $Y2=0
cc_704 N_A_1008_74#_c_810_n N_A_1419_71#_c_1244_n 0.0126239f $X=9.92 $Y=1.285
+ $X2=0 $Y2=0
cc_705 N_A_1008_74#_c_796_n N_A_1419_71#_c_1234_n 0.0135713f $X=7.64 $Y=1.05
+ $X2=0 $Y2=0
cc_706 N_A_1008_74#_c_796_n N_A_1419_71#_c_1235_n 0.0116174f $X=7.64 $Y=1.05
+ $X2=0 $Y2=0
cc_707 N_A_1008_74#_c_797_n N_A_1419_71#_c_1235_n 0.0127109f $X=8.32 $Y=0.34
+ $X2=0 $Y2=0
cc_708 N_A_1008_74#_c_799_n N_A_1419_71#_c_1235_n 0.0273294f $X=8.405 $Y=0.965
+ $X2=0 $Y2=0
cc_709 N_A_1008_74#_c_800_n N_A_1419_71#_c_1235_n 0.0142975f $X=8.49 $Y=1.05
+ $X2=0 $Y2=0
cc_710 N_A_1008_74#_c_800_n N_A_1419_71#_c_1236_n 0.0137179f $X=8.49 $Y=1.05
+ $X2=0 $Y2=0
cc_711 N_A_1008_74#_c_807_n N_A_1419_71#_c_1236_n 0.0408058f $X=9.2 $Y=1.207
+ $X2=0 $Y2=0
cc_712 N_A_1008_74#_c_808_n N_A_1419_71#_c_1236_n 0.0128382f $X=9.37 $Y=1.207
+ $X2=0 $Y2=0
cc_713 N_A_1008_74#_c_807_n N_A_1419_71#_c_1238_n 7.00528e-19 $X=9.2 $Y=1.207
+ $X2=0 $Y2=0
cc_714 N_A_1008_74#_c_796_n N_A_1419_71#_c_1239_n 0.00741769f $X=7.64 $Y=1.05
+ $X2=0 $Y2=0
cc_715 N_A_1008_74#_c_796_n N_A_1419_71#_c_1240_n 0.0307507f $X=7.64 $Y=1.05
+ $X2=0 $Y2=0
cc_716 N_A_1008_74#_c_805_n N_A_1419_71#_c_1240_n 0.00183523f $X=6.76 $Y=1.05
+ $X2=0 $Y2=0
cc_717 N_A_1008_74#_c_793_n N_A_1198_97#_M1033_d 0.0043242f $X=6.04 $Y=1.81
+ $X2=-0.19 $Y2=-0.245
cc_718 N_A_1008_74#_c_796_n N_A_1198_97#_c_1368_n 0.0035241f $X=7.64 $Y=1.05
+ $X2=0 $Y2=0
cc_719 N_A_1008_74#_c_889_p N_A_1198_97#_c_1368_n 0.0138082f $X=7.725 $Y=0.965
+ $X2=0 $Y2=0
cc_720 N_A_1008_74#_c_797_n N_A_1198_97#_c_1368_n 0.0112842f $X=8.32 $Y=0.34
+ $X2=0 $Y2=0
cc_721 N_A_1008_74#_c_798_n N_A_1198_97#_c_1368_n 0.00325013f $X=7.81 $Y=0.34
+ $X2=0 $Y2=0
cc_722 N_A_1008_74#_c_799_n N_A_1198_97#_c_1368_n 0.00344176f $X=8.405 $Y=0.965
+ $X2=0 $Y2=0
cc_723 N_A_1008_74#_c_796_n N_A_1198_97#_c_1371_n 0.00207739f $X=7.64 $Y=1.05
+ $X2=0 $Y2=0
cc_724 N_A_1008_74#_c_797_n N_A_1198_97#_c_1371_n 2.59444e-19 $X=8.32 $Y=0.34
+ $X2=0 $Y2=0
cc_725 N_A_1008_74#_c_800_n N_A_1198_97#_c_1371_n 3.30785e-19 $X=8.49 $Y=1.05
+ $X2=0 $Y2=0
cc_726 N_A_1008_74#_c_787_n N_A_1198_97#_c_1372_n 0.00490388f $X=6.595 $Y=1.015
+ $X2=0 $Y2=0
cc_727 N_A_1008_74#_c_793_n N_A_1198_97#_c_1372_n 0.0684079f $X=6.04 $Y=1.81
+ $X2=0 $Y2=0
cc_728 N_A_1008_74#_c_794_n N_A_1198_97#_c_1372_n 0.012971f $X=6.635 $Y=0.34
+ $X2=0 $Y2=0
cc_729 N_A_1008_74#_c_795_n N_A_1198_97#_c_1372_n 0.0434146f $X=6.76 $Y=0.965
+ $X2=0 $Y2=0
cc_730 N_A_1008_74#_c_813_n N_A_1198_97#_c_1376_n 0.0241319f $X=6.59 $Y=2.465
+ $X2=0 $Y2=0
cc_731 N_A_1008_74#_c_820_n N_A_1198_97#_c_1376_n 0.0313425f $X=6.155 $Y=1.975
+ $X2=0 $Y2=0
cc_732 N_A_1008_74#_c_821_n N_A_1198_97#_c_1376_n 0.011425f $X=6.19 $Y=2.215
+ $X2=0 $Y2=0
cc_733 N_A_1008_74#_c_793_n N_A_1198_97#_c_1373_n 0.016642f $X=6.04 $Y=1.81
+ $X2=0 $Y2=0
cc_734 N_A_1008_74#_c_820_n N_A_1198_97#_c_1373_n 0.0071888f $X=6.155 $Y=1.975
+ $X2=0 $Y2=0
cc_735 N_A_1008_74#_c_821_n N_A_1198_97#_c_1373_n 0.00212672f $X=6.19 $Y=2.215
+ $X2=0 $Y2=0
cc_736 N_A_1008_74#_c_805_n N_A_1198_97#_c_1373_n 0.00693964f $X=6.76 $Y=1.05
+ $X2=0 $Y2=0
cc_737 N_A_1008_74#_c_806_n N_A_1198_97#_c_1373_n 0.00345208f $X=6.72 $Y=1.18
+ $X2=0 $Y2=0
cc_738 N_A_1008_74#_c_796_n N_A_1198_97#_c_1379_n 0.00403611f $X=7.64 $Y=1.05
+ $X2=0 $Y2=0
cc_739 N_A_1008_74#_c_805_n N_A_1198_97#_c_1379_n 0.0035157f $X=6.76 $Y=1.05
+ $X2=0 $Y2=0
cc_740 N_A_1008_74#_c_806_n N_A_1198_97#_c_1379_n 5.63474e-19 $X=6.72 $Y=1.18
+ $X2=0 $Y2=0
cc_741 N_A_1008_74#_c_788_n N_A_1879_74#_c_1518_n 0.0116277f $X=9.32 $Y=1.185
+ $X2=0 $Y2=0
cc_742 N_A_1008_74#_c_801_n N_A_1879_74#_c_1518_n 0.0195638f $X=10.835 $Y=1.205
+ $X2=0 $Y2=0
cc_743 N_A_1008_74#_c_809_n N_A_1879_74#_c_1518_n 0.10001f $X=9.92 $Y=1.285
+ $X2=0 $Y2=0
cc_744 N_A_1008_74#_c_810_n N_A_1879_74#_c_1518_n 0.00751815f $X=9.92 $Y=1.285
+ $X2=0 $Y2=0
cc_745 N_A_1008_74#_c_812_n N_A_1879_74#_c_1518_n 0.00135557f $X=9.755 $Y=1.285
+ $X2=0 $Y2=0
cc_746 N_A_1008_74#_c_815_n N_A_1879_74#_c_1485_n 0.0164887f $X=10.955 $Y=2.14
+ $X2=0 $Y2=0
cc_747 N_A_1008_74#_c_814_n N_A_1879_74#_c_1486_n 0.00537389f $X=10.955 $Y=2.05
+ $X2=0 $Y2=0
cc_748 N_A_1008_74#_c_815_n N_A_1879_74#_c_1486_n 0.011442f $X=10.955 $Y=2.14
+ $X2=0 $Y2=0
cc_749 N_A_1008_74#_c_802_n N_A_1879_74#_c_1486_n 0.0177996f $X=11 $Y=1.635
+ $X2=0 $Y2=0
cc_750 N_A_1008_74#_c_803_n N_A_1879_74#_c_1486_n 0.00286383f $X=11 $Y=1.635
+ $X2=0 $Y2=0
cc_751 N_A_1008_74#_c_801_n N_A_1879_74#_c_1476_n 0.00275916f $X=10.835 $Y=1.205
+ $X2=0 $Y2=0
cc_752 N_A_1008_74#_c_814_n N_A_1879_74#_c_1477_n 0.00365186f $X=10.955 $Y=2.05
+ $X2=0 $Y2=0
cc_753 N_A_1008_74#_c_802_n N_A_1879_74#_c_1477_n 0.022413f $X=11 $Y=1.635 $X2=0
+ $Y2=0
cc_754 N_A_1008_74#_c_803_n N_A_1879_74#_c_1477_n 0.00169441f $X=11 $Y=1.635
+ $X2=0 $Y2=0
cc_755 N_A_1008_74#_c_801_n N_A_1879_74#_c_1479_n 0.0122123f $X=10.835 $Y=1.205
+ $X2=0 $Y2=0
cc_756 N_A_1008_74#_c_802_n N_A_1879_74#_c_1479_n 0.0169626f $X=11 $Y=1.635
+ $X2=0 $Y2=0
cc_757 N_A_1008_74#_c_816_n N_A_27_74#_c_1601_n 0.0143193f $X=5.955 $Y=1.975
+ $X2=0 $Y2=0
cc_758 N_A_1008_74#_c_793_n N_A_27_74#_c_1601_n 0.00755755f $X=6.04 $Y=1.81
+ $X2=0 $Y2=0
cc_759 N_A_1008_74#_M1003_d N_A_27_74#_c_1677_n 0.00611851f $X=5.57 $Y=1.83
+ $X2=0 $Y2=0
cc_760 N_A_1008_74#_c_816_n N_A_27_74#_c_1677_n 0.013259f $X=5.955 $Y=1.975
+ $X2=0 $Y2=0
cc_761 N_A_1008_74#_c_820_n N_A_27_74#_c_1677_n 0.00592943f $X=6.155 $Y=1.975
+ $X2=0 $Y2=0
cc_762 N_A_1008_74#_c_821_n N_A_27_74#_c_1677_n 9.74821e-19 $X=6.19 $Y=2.215
+ $X2=0 $Y2=0
cc_763 N_A_1008_74#_c_790_n N_A_27_74#_c_1602_n 0.0104179f $X=5.18 $Y=0.515
+ $X2=0 $Y2=0
cc_764 N_A_1008_74#_c_816_n N_A_27_74#_c_1602_n 0.00607166f $X=5.955 $Y=1.975
+ $X2=0 $Y2=0
cc_765 N_A_1008_74#_c_793_n N_A_27_74#_c_1602_n 0.0133477f $X=6.04 $Y=1.81 $X2=0
+ $Y2=0
cc_766 N_A_1008_74#_c_790_n N_A_27_74#_c_1603_n 0.0395004f $X=5.18 $Y=0.515
+ $X2=0 $Y2=0
cc_767 N_A_1008_74#_c_791_n N_A_27_74#_c_1603_n 0.0192805f $X=5.955 $Y=0.34
+ $X2=0 $Y2=0
cc_768 N_A_1008_74#_c_793_n N_A_27_74#_c_1603_n 0.0396105f $X=6.04 $Y=1.81 $X2=0
+ $Y2=0
cc_769 N_A_1008_74#_M1003_d N_A_27_74#_c_1705_n 0.0176753f $X=5.57 $Y=1.83 $X2=0
+ $Y2=0
cc_770 N_A_1008_74#_M1003_d N_A_27_74#_c_1618_n 4.91511e-19 $X=5.57 $Y=1.83
+ $X2=0 $Y2=0
cc_771 N_A_1008_74#_M1003_d N_A_27_74#_c_1619_n 0.00368649f $X=5.57 $Y=1.83
+ $X2=0 $Y2=0
cc_772 N_A_1008_74#_c_813_n N_A_27_74#_c_1619_n 0.0056934f $X=6.59 $Y=2.465
+ $X2=0 $Y2=0
cc_773 N_A_1008_74#_c_820_n N_A_27_74#_c_1619_n 0.013596f $X=6.155 $Y=1.975
+ $X2=0 $Y2=0
cc_774 N_A_1008_74#_c_821_n N_A_27_74#_c_1619_n 0.00817649f $X=6.19 $Y=2.215
+ $X2=0 $Y2=0
cc_775 N_A_1008_74#_c_815_n N_VPWR_c_1784_n 0.00204117f $X=10.955 $Y=2.14 $X2=0
+ $Y2=0
cc_776 N_A_1008_74#_c_813_n N_VPWR_c_1792_n 0.00352402f $X=6.59 $Y=2.465 $X2=0
+ $Y2=0
cc_777 N_A_1008_74#_c_815_n N_VPWR_c_1794_n 0.00380268f $X=10.955 $Y=2.14 $X2=0
+ $Y2=0
cc_778 N_A_1008_74#_c_813_n N_VPWR_c_1777_n 0.00525012f $X=6.59 $Y=2.465 $X2=0
+ $Y2=0
cc_779 N_A_1008_74#_c_815_n N_VPWR_c_1777_n 0.0045051f $X=10.955 $Y=2.14 $X2=0
+ $Y2=0
cc_780 N_A_1008_74#_c_821_n N_VPWR_c_1777_n 3.14866e-19 $X=6.19 $Y=2.215 $X2=0
+ $Y2=0
cc_781 N_A_1008_74#_c_796_n N_VGND_M1021_d 0.00452021f $X=7.64 $Y=1.05 $X2=0
+ $Y2=0
cc_782 N_A_1008_74#_c_889_p N_VGND_M1021_d 0.00573796f $X=7.725 $Y=0.965 $X2=0
+ $Y2=0
cc_783 N_A_1008_74#_c_798_n N_VGND_M1021_d 5.22721e-19 $X=7.81 $Y=0.34 $X2=0
+ $Y2=0
cc_784 N_A_1008_74#_c_807_n N_VGND_M1006_s 0.00504668f $X=9.2 $Y=1.207 $X2=0
+ $Y2=0
cc_785 N_A_1008_74#_c_792_n N_VGND_c_1995_n 0.0112234f $X=5.345 $Y=0.34 $X2=0
+ $Y2=0
cc_786 N_A_1008_74#_c_787_n N_VGND_c_1996_n 3.67983e-19 $X=6.595 $Y=1.015 $X2=0
+ $Y2=0
cc_787 N_A_1008_74#_c_794_n N_VGND_c_1996_n 0.00891265f $X=6.635 $Y=0.34 $X2=0
+ $Y2=0
cc_788 N_A_1008_74#_c_795_n N_VGND_c_1996_n 0.0164377f $X=6.76 $Y=0.965 $X2=0
+ $Y2=0
cc_789 N_A_1008_74#_c_796_n N_VGND_c_1996_n 0.0177503f $X=7.64 $Y=1.05 $X2=0
+ $Y2=0
cc_790 N_A_1008_74#_c_889_p N_VGND_c_1996_n 0.0277232f $X=7.725 $Y=0.965 $X2=0
+ $Y2=0
cc_791 N_A_1008_74#_c_798_n N_VGND_c_1996_n 0.0146475f $X=7.81 $Y=0.34 $X2=0
+ $Y2=0
cc_792 N_A_1008_74#_c_788_n N_VGND_c_1997_n 0.00237914f $X=9.32 $Y=1.185 $X2=0
+ $Y2=0
cc_793 N_A_1008_74#_c_797_n N_VGND_c_1997_n 0.0146661f $X=8.32 $Y=0.34 $X2=0
+ $Y2=0
cc_794 N_A_1008_74#_c_799_n N_VGND_c_1997_n 0.0262253f $X=8.405 $Y=0.965 $X2=0
+ $Y2=0
cc_795 N_A_1008_74#_c_807_n N_VGND_c_1997_n 0.0138644f $X=9.2 $Y=1.207 $X2=0
+ $Y2=0
cc_796 N_A_1008_74#_c_787_n N_VGND_c_2007_n 7.53287e-19 $X=6.595 $Y=1.015 $X2=0
+ $Y2=0
cc_797 N_A_1008_74#_c_791_n N_VGND_c_2007_n 0.0392369f $X=5.955 $Y=0.34 $X2=0
+ $Y2=0
cc_798 N_A_1008_74#_c_792_n N_VGND_c_2007_n 0.0179217f $X=5.345 $Y=0.34 $X2=0
+ $Y2=0
cc_799 N_A_1008_74#_c_794_n N_VGND_c_2007_n 0.0507167f $X=6.635 $Y=0.34 $X2=0
+ $Y2=0
cc_800 N_A_1008_74#_c_804_n N_VGND_c_2007_n 0.0121867f $X=6.04 $Y=0.34 $X2=0
+ $Y2=0
cc_801 N_A_1008_74#_c_797_n N_VGND_c_2008_n 0.0446499f $X=8.32 $Y=0.34 $X2=0
+ $Y2=0
cc_802 N_A_1008_74#_c_798_n N_VGND_c_2008_n 0.0120637f $X=7.81 $Y=0.34 $X2=0
+ $Y2=0
cc_803 N_A_1008_74#_c_788_n N_VGND_c_2009_n 0.00461464f $X=9.32 $Y=1.185 $X2=0
+ $Y2=0
cc_804 N_A_1008_74#_c_788_n N_VGND_c_2012_n 0.00913717f $X=9.32 $Y=1.185 $X2=0
+ $Y2=0
cc_805 N_A_1008_74#_c_791_n N_VGND_c_2012_n 0.0229266f $X=5.955 $Y=0.34 $X2=0
+ $Y2=0
cc_806 N_A_1008_74#_c_792_n N_VGND_c_2012_n 0.00971942f $X=5.345 $Y=0.34 $X2=0
+ $Y2=0
cc_807 N_A_1008_74#_c_794_n N_VGND_c_2012_n 0.0288862f $X=6.635 $Y=0.34 $X2=0
+ $Y2=0
cc_808 N_A_1008_74#_c_797_n N_VGND_c_2012_n 0.0252533f $X=8.32 $Y=0.34 $X2=0
+ $Y2=0
cc_809 N_A_1008_74#_c_798_n N_VGND_c_2012_n 0.00644906f $X=7.81 $Y=0.34 $X2=0
+ $Y2=0
cc_810 N_A_1008_74#_c_804_n N_VGND_c_2012_n 0.00660921f $X=6.04 $Y=0.34 $X2=0
+ $Y2=0
cc_811 N_A_1008_74#_c_795_n A_1334_97# 0.00555912f $X=6.76 $Y=0.965 $X2=-0.19
+ $Y2=-0.245
cc_812 N_A_1008_74#_c_807_n A_1807_74# 0.00366293f $X=9.2 $Y=1.207 $X2=-0.19
+ $Y2=-0.245
cc_813 N_A_818_74#_c_1042_n N_A_1419_71#_M1016_d 0.00638803f $X=9.235 $Y=2.84
+ $X2=0 $Y2=0
cc_814 N_A_818_74#_c_1123_p N_A_1419_71#_M1016_d 0.00896756f $X=8.28 $Y=2.63
+ $X2=0 $Y2=0
cc_815 N_A_818_74#_c_1015_n N_A_1419_71#_c_1232_n 0.0171753f $X=6.595 $Y=1.68
+ $X2=0 $Y2=0
cc_816 N_A_818_74#_c_1047_n N_A_1419_71#_c_1232_n 0.00757834f $X=7.235 $Y=2.23
+ $X2=0 $Y2=0
cc_817 N_A_818_74#_c_1034_n N_A_1419_71#_c_1243_n 0.0142752f $X=7.055 $Y=2.215
+ $X2=0 $Y2=0
cc_818 N_A_818_74#_c_1035_n N_A_1419_71#_c_1243_n 0.0220573f $X=7.04 $Y=2.465
+ $X2=0 $Y2=0
cc_819 N_A_818_74#_c_1041_n N_A_1419_71#_c_1243_n 0.0036165f $X=7.235 $Y=2.545
+ $X2=0 $Y2=0
cc_820 N_A_818_74#_c_1129_p N_A_1419_71#_c_1243_n 0.0146186f $X=8.195 $Y=2.63
+ $X2=0 $Y2=0
cc_821 N_A_818_74#_c_1123_p N_A_1419_71#_c_1243_n 8.85409e-19 $X=8.28 $Y=2.63
+ $X2=0 $Y2=0
cc_822 N_A_818_74#_c_1016_n N_A_1419_71#_c_1244_n 0.00942133f $X=10.385 $Y=1.885
+ $X2=0 $Y2=0
cc_823 N_A_818_74#_c_1043_n N_A_1419_71#_c_1244_n 0.0109739f $X=9.32 $Y=2.755
+ $X2=0 $Y2=0
cc_824 N_A_818_74#_c_1025_n N_A_1419_71#_c_1244_n 0.0250829f $X=10.295 $Y=1.705
+ $X2=0 $Y2=0
cc_825 N_A_818_74#_c_1026_n N_A_1419_71#_c_1244_n 0.00336657f $X=9.405 $Y=1.705
+ $X2=0 $Y2=0
cc_826 N_A_818_74#_c_1016_n N_A_1419_71#_c_1245_n 0.0524942f $X=10.385 $Y=1.885
+ $X2=0 $Y2=0
cc_827 N_A_818_74#_c_1043_n N_A_1419_71#_c_1245_n 0.0018203f $X=9.32 $Y=2.755
+ $X2=0 $Y2=0
cc_828 N_A_818_74#_c_1042_n N_A_1419_71#_c_1246_n 0.0143404f $X=9.235 $Y=2.84
+ $X2=0 $Y2=0
cc_829 N_A_818_74#_c_1123_p N_A_1419_71#_c_1246_n 0.00603276f $X=8.28 $Y=2.63
+ $X2=0 $Y2=0
cc_830 N_A_818_74#_c_1042_n N_A_1419_71#_c_1247_n 0.0253999f $X=9.235 $Y=2.84
+ $X2=0 $Y2=0
cc_831 N_A_818_74#_c_1043_n N_A_1419_71#_c_1247_n 0.0311064f $X=9.32 $Y=2.755
+ $X2=0 $Y2=0
cc_832 N_A_818_74#_c_1123_p N_A_1419_71#_c_1247_n 0.00175868f $X=8.28 $Y=2.63
+ $X2=0 $Y2=0
cc_833 N_A_818_74#_c_1043_n N_A_1419_71#_c_1237_n 0.021419f $X=9.32 $Y=2.755
+ $X2=0 $Y2=0
cc_834 N_A_818_74#_c_1026_n N_A_1419_71#_c_1237_n 0.010381f $X=9.405 $Y=1.705
+ $X2=0 $Y2=0
cc_835 N_A_818_74#_c_1026_n N_A_1419_71#_c_1238_n 0.00188287f $X=9.405 $Y=1.705
+ $X2=0 $Y2=0
cc_836 N_A_818_74#_c_1015_n N_A_1419_71#_c_1239_n 0.00374419f $X=6.595 $Y=1.68
+ $X2=0 $Y2=0
cc_837 N_A_818_74#_c_1042_n N_A_1419_71#_c_1249_n 0.00250279f $X=9.235 $Y=2.84
+ $X2=0 $Y2=0
cc_838 N_A_818_74#_c_1043_n N_A_1419_71#_c_1249_n 0.0154498f $X=9.32 $Y=2.755
+ $X2=0 $Y2=0
cc_839 N_A_818_74#_c_1129_p N_A_1198_97#_c_1370_n 0.0124298f $X=8.195 $Y=2.63
+ $X2=0 $Y2=0
cc_840 N_A_818_74#_c_1042_n N_A_1198_97#_c_1370_n 0.00102155f $X=9.235 $Y=2.84
+ $X2=0 $Y2=0
cc_841 N_A_818_74#_c_1123_p N_A_1198_97#_c_1370_n 0.0133205f $X=8.28 $Y=2.63
+ $X2=0 $Y2=0
cc_842 N_A_818_74#_M1033_g N_A_1198_97#_c_1372_n 0.00292584f $X=5.915 $Y=0.695
+ $X2=0 $Y2=0
cc_843 N_A_818_74#_c_1015_n N_A_1198_97#_c_1376_n 0.0117545f $X=6.595 $Y=1.68
+ $X2=0 $Y2=0
cc_844 N_A_818_74#_c_1034_n N_A_1198_97#_c_1376_n 0.00307881f $X=7.055 $Y=2.215
+ $X2=0 $Y2=0
cc_845 N_A_818_74#_c_1035_n N_A_1198_97#_c_1376_n 0.0100095f $X=7.04 $Y=2.465
+ $X2=0 $Y2=0
cc_846 N_A_818_74#_c_1041_n N_A_1198_97#_c_1376_n 0.00627244f $X=7.235 $Y=2.545
+ $X2=0 $Y2=0
cc_847 N_A_818_74#_c_1047_n N_A_1198_97#_c_1376_n 0.0276179f $X=7.235 $Y=2.23
+ $X2=0 $Y2=0
cc_848 N_A_818_74#_M1033_g N_A_1198_97#_c_1373_n 4.8526e-19 $X=5.915 $Y=0.695
+ $X2=0 $Y2=0
cc_849 N_A_818_74#_c_1015_n N_A_1198_97#_c_1373_n 0.0228797f $X=6.595 $Y=1.68
+ $X2=0 $Y2=0
cc_850 N_A_818_74#_c_1129_p N_A_1198_97#_c_1374_n 0.00628566f $X=8.195 $Y=2.63
+ $X2=0 $Y2=0
cc_851 N_A_818_74#_c_1123_p N_A_1198_97#_c_1374_n 9.20527e-19 $X=8.28 $Y=2.63
+ $X2=0 $Y2=0
cc_852 N_A_818_74#_c_1015_n N_A_1198_97#_c_1379_n 0.0197908f $X=6.595 $Y=1.68
+ $X2=0 $Y2=0
cc_853 N_A_818_74#_c_1129_p N_A_1198_97#_c_1379_n 0.0148484f $X=8.195 $Y=2.63
+ $X2=0 $Y2=0
cc_854 N_A_818_74#_c_1047_n N_A_1198_97#_c_1379_n 0.0293015f $X=7.235 $Y=2.23
+ $X2=0 $Y2=0
cc_855 N_A_818_74#_c_1019_n N_A_1879_74#_c_1518_n 0.0109116f $X=10.625 $Y=1.185
+ $X2=0 $Y2=0
cc_856 N_A_818_74#_c_1020_n N_A_1879_74#_c_1518_n 0.0126814f $X=11.06 $Y=1.11
+ $X2=0 $Y2=0
cc_857 N_A_818_74#_c_1016_n N_A_1879_74#_c_1484_n 0.00409881f $X=10.385 $Y=1.885
+ $X2=0 $Y2=0
cc_858 N_A_818_74#_c_1028_n N_A_1879_74#_c_1484_n 0.00999652f $X=10.46 $Y=1.625
+ $X2=0 $Y2=0
cc_859 N_A_818_74#_c_1016_n N_A_1879_74#_c_1485_n 0.014436f $X=10.385 $Y=1.885
+ $X2=0 $Y2=0
cc_860 N_A_818_74#_c_1020_n N_A_1879_74#_c_1476_n 0.00379106f $X=11.06 $Y=1.11
+ $X2=0 $Y2=0
cc_861 N_A_818_74#_c_1017_n N_A_1879_74#_c_1479_n 3.31074e-19 $X=10.55 $Y=1.46
+ $X2=0 $Y2=0
cc_862 N_A_818_74#_c_1018_n N_A_1879_74#_c_1479_n 7.91946e-19 $X=10.985 $Y=1.185
+ $X2=0 $Y2=0
cc_863 N_A_818_74#_c_1039_n N_A_27_74#_c_1600_n 0.00971937f $X=4.555 $Y=1.975
+ $X2=0 $Y2=0
cc_864 N_A_818_74#_M1005_d N_A_27_74#_c_1616_n 0.00838378f $X=4.18 $Y=1.84 $X2=0
+ $Y2=0
cc_865 N_A_818_74#_c_1012_n N_A_27_74#_c_1616_n 0.00193622f $X=5.42 $Y=1.68
+ $X2=0 $Y2=0
cc_866 N_A_818_74#_c_1039_n N_A_27_74#_c_1616_n 0.0551459f $X=4.555 $Y=1.975
+ $X2=0 $Y2=0
cc_867 N_A_818_74#_c_1029_n N_A_27_74#_c_1616_n 0.0114083f $X=4.837 $Y=1.68
+ $X2=0 $Y2=0
cc_868 N_A_818_74#_M1030_g N_A_27_74#_c_1601_n 0.002953f $X=4.965 $Y=0.74 $X2=0
+ $Y2=0
cc_869 N_A_818_74#_c_1012_n N_A_27_74#_c_1601_n 0.0137254f $X=5.42 $Y=1.68 $X2=0
+ $Y2=0
cc_870 N_A_818_74#_c_1031_n N_A_27_74#_c_1601_n 0.00603813f $X=5.495 $Y=1.755
+ $X2=0 $Y2=0
cc_871 N_A_818_74#_M1033_g N_A_27_74#_c_1601_n 0.00213848f $X=5.915 $Y=0.695
+ $X2=0 $Y2=0
cc_872 N_A_818_74#_c_1024_n N_A_27_74#_c_1601_n 0.00915757f $X=4.64 $Y=1.81
+ $X2=0 $Y2=0
cc_873 N_A_818_74#_c_1046_n N_A_27_74#_c_1601_n 0.0191537f $X=4.8 $Y=1.975 $X2=0
+ $Y2=0
cc_874 N_A_818_74#_c_1029_n N_A_27_74#_c_1601_n 0.0034344f $X=4.837 $Y=1.68
+ $X2=0 $Y2=0
cc_875 N_A_818_74#_c_1031_n N_A_27_74#_c_1677_n 0.0156812f $X=5.495 $Y=1.755
+ $X2=0 $Y2=0
cc_876 N_A_818_74#_M1030_g N_A_27_74#_c_1602_n 0.00405031f $X=4.965 $Y=0.74
+ $X2=0 $Y2=0
cc_877 N_A_818_74#_c_1012_n N_A_27_74#_c_1602_n 0.0109179f $X=5.42 $Y=1.68 $X2=0
+ $Y2=0
cc_878 N_A_818_74#_M1033_g N_A_27_74#_c_1602_n 0.0038364f $X=5.915 $Y=0.695
+ $X2=0 $Y2=0
cc_879 N_A_818_74#_c_1024_n N_A_27_74#_c_1602_n 0.00665823f $X=4.64 $Y=1.81
+ $X2=0 $Y2=0
cc_880 N_A_818_74#_M1030_g N_A_27_74#_c_1603_n 0.00511417f $X=4.965 $Y=0.74
+ $X2=0 $Y2=0
cc_881 N_A_818_74#_M1033_g N_A_27_74#_c_1603_n 0.00876272f $X=5.915 $Y=0.695
+ $X2=0 $Y2=0
cc_882 N_A_818_74#_c_1031_n N_A_27_74#_c_1618_n 0.00377169f $X=5.495 $Y=1.755
+ $X2=0 $Y2=0
cc_883 N_A_818_74#_c_1129_p N_VPWR_M1034_d 0.0117246f $X=8.195 $Y=2.63 $X2=0
+ $Y2=0
cc_884 N_A_818_74#_c_1031_n N_VPWR_c_1781_n 0.00804469f $X=5.495 $Y=1.755 $X2=0
+ $Y2=0
cc_885 N_A_818_74#_c_1129_p N_VPWR_c_1782_n 0.024844f $X=8.195 $Y=2.63 $X2=0
+ $Y2=0
cc_886 N_A_818_74#_c_1123_p N_VPWR_c_1782_n 0.00295969f $X=8.28 $Y=2.63 $X2=0
+ $Y2=0
cc_887 N_A_818_74#_c_1016_n N_VPWR_c_1783_n 0.00353387f $X=10.385 $Y=1.885 $X2=0
+ $Y2=0
cc_888 N_A_818_74#_c_1042_n N_VPWR_c_1783_n 0.0150383f $X=9.235 $Y=2.84 $X2=0
+ $Y2=0
cc_889 N_A_818_74#_c_1043_n N_VPWR_c_1783_n 0.0629935f $X=9.32 $Y=2.755 $X2=0
+ $Y2=0
cc_890 N_A_818_74#_c_1025_n N_VPWR_c_1783_n 0.021234f $X=10.295 $Y=1.705 $X2=0
+ $Y2=0
cc_891 N_A_818_74#_c_1031_n N_VPWR_c_1792_n 0.00512473f $X=5.495 $Y=1.755 $X2=0
+ $Y2=0
cc_892 N_A_818_74#_c_1035_n N_VPWR_c_1792_n 0.00444469f $X=7.04 $Y=2.465 $X2=0
+ $Y2=0
cc_893 N_A_818_74#_c_1129_p N_VPWR_c_1792_n 0.00575245f $X=8.195 $Y=2.63 $X2=0
+ $Y2=0
cc_894 N_A_818_74#_c_1203_p N_VPWR_c_1792_n 0.00305489f $X=7.32 $Y=2.63 $X2=0
+ $Y2=0
cc_895 N_A_818_74#_c_1129_p N_VPWR_c_1793_n 0.00252675f $X=8.195 $Y=2.63 $X2=0
+ $Y2=0
cc_896 N_A_818_74#_c_1042_n N_VPWR_c_1793_n 0.0348172f $X=9.235 $Y=2.84 $X2=0
+ $Y2=0
cc_897 N_A_818_74#_c_1123_p N_VPWR_c_1793_n 0.00478198f $X=8.28 $Y=2.63 $X2=0
+ $Y2=0
cc_898 N_A_818_74#_c_1016_n N_VPWR_c_1794_n 0.00445602f $X=10.385 $Y=1.885 $X2=0
+ $Y2=0
cc_899 N_A_818_74#_c_1031_n N_VPWR_c_1777_n 0.00492022f $X=5.495 $Y=1.755 $X2=0
+ $Y2=0
cc_900 N_A_818_74#_c_1035_n N_VPWR_c_1777_n 0.00892093f $X=7.04 $Y=2.465 $X2=0
+ $Y2=0
cc_901 N_A_818_74#_c_1016_n N_VPWR_c_1777_n 0.00862959f $X=10.385 $Y=1.885 $X2=0
+ $Y2=0
cc_902 N_A_818_74#_c_1129_p N_VPWR_c_1777_n 0.0161685f $X=8.195 $Y=2.63 $X2=0
+ $Y2=0
cc_903 N_A_818_74#_c_1203_p N_VPWR_c_1777_n 0.00506135f $X=7.32 $Y=2.63 $X2=0
+ $Y2=0
cc_904 N_A_818_74#_c_1042_n N_VPWR_c_1777_n 0.0356528f $X=9.235 $Y=2.84 $X2=0
+ $Y2=0
cc_905 N_A_818_74#_c_1123_p N_VPWR_c_1777_n 0.00563039f $X=8.28 $Y=2.63 $X2=0
+ $Y2=0
cc_906 N_A_818_74#_c_1129_p A_1423_508# 0.00363958f $X=8.195 $Y=2.63 $X2=-0.19
+ $Y2=-0.245
cc_907 N_A_818_74#_c_1203_p A_1423_508# 0.00361866f $X=7.32 $Y=2.63 $X2=-0.19
+ $Y2=-0.245
cc_908 N_A_818_74#_c_1024_n N_VGND_M1030_s 0.00199309f $X=4.64 $Y=1.81 $X2=0
+ $Y2=0
cc_909 N_A_818_74#_c_1027_n N_VGND_M1030_s 0.00426582f $X=4.64 $Y=0.925 $X2=0
+ $Y2=0
cc_910 N_A_818_74#_c_1023_n N_VGND_c_1994_n 0.0182488f $X=4.23 $Y=0.515 $X2=0
+ $Y2=0
cc_911 N_A_818_74#_M1030_g N_VGND_c_1995_n 0.00936698f $X=4.965 $Y=0.74 $X2=0
+ $Y2=0
cc_912 N_A_818_74#_c_1023_n N_VGND_c_1995_n 0.0246408f $X=4.23 $Y=0.515 $X2=0
+ $Y2=0
cc_913 N_A_818_74#_c_1027_n N_VGND_c_1995_n 0.0111795f $X=4.64 $Y=0.925 $X2=0
+ $Y2=0
cc_914 N_A_818_74#_c_1023_n N_VGND_c_2004_n 0.0142249f $X=4.23 $Y=0.515 $X2=0
+ $Y2=0
cc_915 N_A_818_74#_M1030_g N_VGND_c_2007_n 0.00383152f $X=4.965 $Y=0.74 $X2=0
+ $Y2=0
cc_916 N_A_818_74#_M1033_g N_VGND_c_2007_n 7.53287e-19 $X=5.915 $Y=0.695 $X2=0
+ $Y2=0
cc_917 N_A_818_74#_c_1020_n N_VGND_c_2009_n 0.00333934f $X=11.06 $Y=1.11 $X2=0
+ $Y2=0
cc_918 N_A_818_74#_M1030_g N_VGND_c_2012_n 0.00762539f $X=4.965 $Y=0.74 $X2=0
+ $Y2=0
cc_919 N_A_818_74#_c_1020_n N_VGND_c_2012_n 0.00479212f $X=11.06 $Y=1.11 $X2=0
+ $Y2=0
cc_920 N_A_818_74#_c_1023_n N_VGND_c_2012_n 0.011867f $X=4.23 $Y=0.515 $X2=0
+ $Y2=0
cc_921 N_A_818_74#_c_1027_n N_VGND_c_2012_n 0.00711058f $X=4.64 $Y=0.925 $X2=0
+ $Y2=0
cc_922 N_A_1419_71#_M1021_g N_A_1198_97#_c_1368_n 0.0128473f $X=7.17 $Y=0.695
+ $X2=0 $Y2=0
cc_923 N_A_1419_71#_c_1235_n N_A_1198_97#_c_1368_n 0.00210086f $X=8.065 $Y=0.81
+ $X2=0 $Y2=0
cc_924 N_A_1419_71#_c_1234_n N_A_1198_97#_c_1369_n 0.00588549f $X=7.98 $Y=1.39
+ $X2=0 $Y2=0
cc_925 N_A_1419_71#_c_1235_n N_A_1198_97#_c_1369_n 0.00279446f $X=8.065 $Y=0.81
+ $X2=0 $Y2=0
cc_926 N_A_1419_71#_c_1237_n N_A_1198_97#_c_1369_n 0.00259234f $X=8.865 $Y=1.74
+ $X2=0 $Y2=0
cc_927 N_A_1419_71#_c_1238_n N_A_1198_97#_c_1369_n 9.68537e-19 $X=8.865 $Y=1.74
+ $X2=0 $Y2=0
cc_928 N_A_1419_71#_c_1239_n N_A_1198_97#_c_1369_n 0.017706f $X=7.37 $Y=1.435
+ $X2=0 $Y2=0
cc_929 N_A_1419_71#_c_1240_n N_A_1198_97#_c_1369_n 4.74622e-19 $X=7.535 $Y=1.437
+ $X2=0 $Y2=0
cc_930 N_A_1419_71#_c_1241_n N_A_1198_97#_c_1369_n 0.00706594f $X=8.065 $Y=1.39
+ $X2=0 $Y2=0
cc_931 N_A_1419_71#_c_1232_n N_A_1198_97#_c_1370_n 0.0266926f $X=7.55 $Y=2.375
+ $X2=0 $Y2=0
cc_932 N_A_1419_71#_c_1243_n N_A_1198_97#_c_1370_n 0.0140299f $X=7.55 $Y=2.465
+ $X2=0 $Y2=0
cc_933 N_A_1419_71#_c_1236_n N_A_1198_97#_c_1370_n 0.00209193f $X=8.7 $Y=1.39
+ $X2=0 $Y2=0
cc_934 N_A_1419_71#_c_1246_n N_A_1198_97#_c_1370_n 0.00581956f $X=8.7 $Y=2.25
+ $X2=0 $Y2=0
cc_935 N_A_1419_71#_c_1247_n N_A_1198_97#_c_1370_n 6.47508e-19 $X=8.865 $Y=2.125
+ $X2=0 $Y2=0
cc_936 N_A_1419_71#_c_1237_n N_A_1198_97#_c_1370_n 0.00155708f $X=8.865 $Y=1.74
+ $X2=0 $Y2=0
cc_937 N_A_1419_71#_c_1238_n N_A_1198_97#_c_1370_n 0.0113869f $X=8.865 $Y=1.74
+ $X2=0 $Y2=0
cc_938 N_A_1419_71#_c_1241_n N_A_1198_97#_c_1370_n 0.001391f $X=8.065 $Y=1.39
+ $X2=0 $Y2=0
cc_939 N_A_1419_71#_c_1249_n N_A_1198_97#_c_1370_n 0.00857715f $X=8.865 $Y=2.42
+ $X2=0 $Y2=0
cc_940 N_A_1419_71#_c_1234_n N_A_1198_97#_c_1371_n 0.00655034f $X=7.98 $Y=1.39
+ $X2=0 $Y2=0
cc_941 N_A_1419_71#_c_1235_n N_A_1198_97#_c_1371_n 0.0101181f $X=8.065 $Y=0.81
+ $X2=0 $Y2=0
cc_942 N_A_1419_71#_c_1239_n N_A_1198_97#_c_1371_n 6.75815e-19 $X=7.37 $Y=1.435
+ $X2=0 $Y2=0
cc_943 N_A_1419_71#_c_1239_n N_A_1198_97#_c_1372_n 4.83812e-19 $X=7.37 $Y=1.435
+ $X2=0 $Y2=0
cc_944 N_A_1419_71#_c_1243_n N_A_1198_97#_c_1376_n 0.00134027f $X=7.55 $Y=2.465
+ $X2=0 $Y2=0
cc_945 N_A_1419_71#_c_1239_n N_A_1198_97#_c_1373_n 0.0014698f $X=7.37 $Y=1.435
+ $X2=0 $Y2=0
cc_946 N_A_1419_71#_c_1240_n N_A_1198_97#_c_1373_n 0.00200168f $X=7.535 $Y=1.437
+ $X2=0 $Y2=0
cc_947 N_A_1419_71#_c_1232_n N_A_1198_97#_c_1374_n 0.00118446f $X=7.55 $Y=2.375
+ $X2=0 $Y2=0
cc_948 N_A_1419_71#_c_1234_n N_A_1198_97#_c_1374_n 0.00294848f $X=7.98 $Y=1.39
+ $X2=0 $Y2=0
cc_949 N_A_1419_71#_c_1236_n N_A_1198_97#_c_1374_n 0.00684268f $X=8.7 $Y=1.39
+ $X2=0 $Y2=0
cc_950 N_A_1419_71#_c_1246_n N_A_1198_97#_c_1374_n 0.00156617f $X=8.7 $Y=2.25
+ $X2=0 $Y2=0
cc_951 N_A_1419_71#_c_1237_n N_A_1198_97#_c_1374_n 0.00969696f $X=8.865 $Y=1.74
+ $X2=0 $Y2=0
cc_952 N_A_1419_71#_c_1238_n N_A_1198_97#_c_1374_n 0.00135816f $X=8.865 $Y=1.74
+ $X2=0 $Y2=0
cc_953 N_A_1419_71#_c_1241_n N_A_1198_97#_c_1374_n 0.0114927f $X=8.065 $Y=1.39
+ $X2=0 $Y2=0
cc_954 N_A_1419_71#_c_1232_n N_A_1198_97#_c_1379_n 0.0152333f $X=7.55 $Y=2.375
+ $X2=0 $Y2=0
cc_955 N_A_1419_71#_c_1234_n N_A_1198_97#_c_1379_n 0.0134128f $X=7.98 $Y=1.39
+ $X2=0 $Y2=0
cc_956 N_A_1419_71#_c_1239_n N_A_1198_97#_c_1379_n 0.00580021f $X=7.37 $Y=1.435
+ $X2=0 $Y2=0
cc_957 N_A_1419_71#_c_1240_n N_A_1198_97#_c_1379_n 0.0186728f $X=7.535 $Y=1.437
+ $X2=0 $Y2=0
cc_958 N_A_1419_71#_c_1245_n N_A_1879_74#_c_1484_n 4.88662e-19 $X=9.965 $Y=1.885
+ $X2=0 $Y2=0
cc_959 N_A_1419_71#_c_1245_n N_A_1879_74#_c_1485_n 0.00237971f $X=9.965 $Y=1.885
+ $X2=0 $Y2=0
cc_960 N_A_1419_71#_c_1243_n N_VPWR_c_1782_n 0.00588667f $X=7.55 $Y=2.465 $X2=0
+ $Y2=0
cc_961 N_A_1419_71#_c_1244_n N_VPWR_c_1783_n 0.00503097f $X=9.89 $Y=1.81 $X2=0
+ $Y2=0
cc_962 N_A_1419_71#_c_1245_n N_VPWR_c_1783_n 0.0222536f $X=9.965 $Y=1.885 $X2=0
+ $Y2=0
cc_963 N_A_1419_71#_c_1243_n N_VPWR_c_1792_n 0.00324023f $X=7.55 $Y=2.465 $X2=0
+ $Y2=0
cc_964 N_A_1419_71#_c_1245_n N_VPWR_c_1794_n 0.00413917f $X=9.965 $Y=1.885 $X2=0
+ $Y2=0
cc_965 N_A_1419_71#_c_1243_n N_VPWR_c_1777_n 0.0041065f $X=7.55 $Y=2.465 $X2=0
+ $Y2=0
cc_966 N_A_1419_71#_c_1245_n N_VPWR_c_1777_n 0.00817532f $X=9.965 $Y=1.885 $X2=0
+ $Y2=0
cc_967 N_A_1419_71#_M1021_g N_VGND_c_1996_n 0.00887076f $X=7.17 $Y=0.695 $X2=0
+ $Y2=0
cc_968 N_A_1419_71#_M1006_g N_VGND_c_1997_n 0.0130682f $X=8.96 $Y=0.74 $X2=0
+ $Y2=0
cc_969 N_A_1419_71#_M1021_g N_VGND_c_2007_n 0.00413255f $X=7.17 $Y=0.695 $X2=0
+ $Y2=0
cc_970 N_A_1419_71#_M1006_g N_VGND_c_2009_n 0.00383152f $X=8.96 $Y=0.74 $X2=0
+ $Y2=0
cc_971 N_A_1419_71#_M1021_g N_VGND_c_2012_n 0.00428305f $X=7.17 $Y=0.695 $X2=0
+ $Y2=0
cc_972 N_A_1419_71#_M1006_g N_VGND_c_2012_n 0.0075694f $X=8.96 $Y=0.74 $X2=0
+ $Y2=0
cc_973 N_A_1198_97#_c_1376_n N_A_27_74#_c_1619_n 0.00642296f $X=6.635 $Y=2.55
+ $X2=0 $Y2=0
cc_974 N_A_1198_97#_c_1370_n N_VPWR_c_1782_n 0.00511117f $X=8.17 $Y=2.045 $X2=0
+ $Y2=0
cc_975 N_A_1198_97#_c_1376_n N_VPWR_c_1792_n 0.0161533f $X=6.635 $Y=2.55 $X2=0
+ $Y2=0
cc_976 N_A_1198_97#_c_1370_n N_VPWR_c_1793_n 0.00316704f $X=8.17 $Y=2.045 $X2=0
+ $Y2=0
cc_977 N_A_1198_97#_c_1370_n N_VPWR_c_1777_n 0.00399574f $X=8.17 $Y=2.045 $X2=0
+ $Y2=0
cc_978 N_A_1198_97#_c_1376_n N_VPWR_c_1777_n 0.0144706f $X=6.635 $Y=2.55 $X2=0
+ $Y2=0
cc_979 N_A_1198_97#_c_1368_n N_VGND_c_1996_n 0.00222522f $X=7.85 $Y=1.085 $X2=0
+ $Y2=0
cc_980 N_A_1198_97#_c_1368_n N_VGND_c_2008_n 0.00278237f $X=7.85 $Y=1.085 $X2=0
+ $Y2=0
cc_981 N_A_1198_97#_c_1368_n N_VGND_c_2012_n 0.00363424f $X=7.85 $Y=1.085 $X2=0
+ $Y2=0
cc_982 N_A_1879_74#_c_1484_n N_VPWR_c_1783_n 0.00524238f $X=10.61 $Y=2.155 $X2=0
+ $Y2=0
cc_983 N_A_1879_74#_c_1485_n N_VPWR_c_1783_n 0.0239768f $X=10.61 $Y=2.815 $X2=0
+ $Y2=0
cc_984 N_A_1879_74#_c_1480_n N_VPWR_c_1784_n 0.0137799f $X=12.39 $Y=1.75 $X2=0
+ $Y2=0
cc_985 N_A_1879_74#_c_1472_n N_VPWR_c_1784_n 5.26364e-19 $X=12.48 $Y=1.36 $X2=0
+ $Y2=0
cc_986 N_A_1879_74#_c_1483_n N_VPWR_c_1785_n 0.00718907f $X=13.4 $Y=1.765 $X2=0
+ $Y2=0
cc_987 N_A_1879_74#_c_1485_n N_VPWR_c_1794_n 0.0145938f $X=10.61 $Y=2.815 $X2=0
+ $Y2=0
cc_988 N_A_1879_74#_c_1480_n N_VPWR_c_1795_n 0.00472847f $X=12.39 $Y=1.75 $X2=0
+ $Y2=0
cc_989 N_A_1879_74#_c_1483_n N_VPWR_c_1795_n 0.00445602f $X=13.4 $Y=1.765 $X2=0
+ $Y2=0
cc_990 N_A_1879_74#_c_1480_n N_VPWR_c_1777_n 0.00503886f $X=12.39 $Y=1.75 $X2=0
+ $Y2=0
cc_991 N_A_1879_74#_c_1483_n N_VPWR_c_1777_n 0.00862475f $X=13.4 $Y=1.765 $X2=0
+ $Y2=0
cc_992 N_A_1879_74#_c_1485_n N_VPWR_c_1777_n 0.0120466f $X=10.61 $Y=2.815 $X2=0
+ $Y2=0
cc_993 N_A_1879_74#_c_1471_n N_Q_c_1939_n 0.00625823f $X=13.07 $Y=1.36 $X2=0
+ $Y2=0
cc_994 N_A_1879_74#_c_1473_n N_Q_c_1939_n 0.00440101f $X=13.145 $Y=1.205 $X2=0
+ $Y2=0
cc_995 N_A_1879_74#_c_1483_n Q 0.003159f $X=13.4 $Y=1.765 $X2=0 $Y2=0
cc_996 N_A_1879_74#_c_1475_n Q 0.00523601f $X=13.4 $Y=1.36 $X2=0 $Y2=0
cc_997 N_A_1879_74#_c_1480_n Q 0.00193457f $X=12.39 $Y=1.75 $X2=0 $Y2=0
cc_998 N_A_1879_74#_c_1483_n Q 0.0112875f $X=13.4 $Y=1.765 $X2=0 $Y2=0
cc_999 N_A_1879_74#_c_1480_n N_Q_c_1940_n 0.002508f $X=12.39 $Y=1.75 $X2=0 $Y2=0
cc_1000 N_A_1879_74#_c_1471_n N_Q_c_1940_n 0.018157f $X=13.07 $Y=1.36 $X2=0
+ $Y2=0
cc_1001 N_A_1879_74#_c_1472_n N_Q_c_1940_n 0.00153496f $X=12.48 $Y=1.36 $X2=0
+ $Y2=0
cc_1002 N_A_1879_74#_c_1473_n N_Q_c_1940_n 0.00561072f $X=13.145 $Y=1.205 $X2=0
+ $Y2=0
cc_1003 N_A_1879_74#_c_1474_n N_Q_c_1940_n 0.00465733f $X=13.4 $Y=1.675 $X2=0
+ $Y2=0
cc_1004 N_A_1879_74#_c_1483_n N_Q_c_1940_n 0.0017333f $X=13.4 $Y=1.765 $X2=0
+ $Y2=0
cc_1005 N_A_1879_74#_c_1475_n N_Q_c_1940_n 0.00544113f $X=13.4 $Y=1.36 $X2=0
+ $Y2=0
cc_1006 N_A_1879_74#_c_1518_n N_VGND_c_1997_n 0.00427951f $X=11.275 $Y=0.785
+ $X2=0 $Y2=0
cc_1007 N_A_1879_74#_M1015_g N_VGND_c_1998_n 0.00864682f $X=12.105 $Y=0.69 $X2=0
+ $Y2=0
cc_1008 N_A_1879_74#_c_1472_n N_VGND_c_1998_n 0.0057671f $X=12.48 $Y=1.36 $X2=0
+ $Y2=0
cc_1009 N_A_1879_74#_c_1518_n N_VGND_c_1998_n 0.0230855f $X=11.275 $Y=0.785
+ $X2=0 $Y2=0
cc_1010 N_A_1879_74#_c_1476_n N_VGND_c_1998_n 0.0021734f $X=11.36 $Y=1.155 $X2=0
+ $Y2=0
cc_1011 N_A_1879_74#_c_1478_n N_VGND_c_1998_n 0.0262585f $X=11.9 $Y=1.32 $X2=0
+ $Y2=0
cc_1012 N_A_1879_74#_c_1473_n N_VGND_c_1999_n 0.00145725f $X=13.145 $Y=1.205
+ $X2=0 $Y2=0
cc_1013 N_A_1879_74#_c_1518_n N_VGND_c_2009_n 0.0343006f $X=11.275 $Y=0.785
+ $X2=0 $Y2=0
cc_1014 N_A_1879_74#_M1015_g N_VGND_c_2010_n 0.00430908f $X=12.105 $Y=0.69 $X2=0
+ $Y2=0
cc_1015 N_A_1879_74#_c_1473_n N_VGND_c_2010_n 9.59479e-19 $X=13.145 $Y=1.205
+ $X2=0 $Y2=0
cc_1016 N_A_1879_74#_M1015_g N_VGND_c_2012_n 0.00825456f $X=12.105 $Y=0.69 $X2=0
+ $Y2=0
cc_1017 N_A_1879_74#_c_1518_n N_VGND_c_2012_n 0.0564515f $X=11.275 $Y=0.785
+ $X2=0 $Y2=0
cc_1018 N_A_1879_74#_c_1518_n A_2227_118# 0.0055961f $X=11.275 $Y=0.785
+ $X2=-0.19 $Y2=-0.245
cc_1019 N_A_1879_74#_c_1476_n A_2227_118# 6.71699e-19 $X=11.36 $Y=1.155
+ $X2=-0.19 $Y2=-0.245
cc_1020 N_A_27_74#_c_1610_n N_VPWR_M1032_d 3.33888e-19 $X=2.055 $Y=2.99 $X2=0
+ $Y2=0
cc_1021 N_A_27_74#_c_1646_n N_VPWR_M1032_d 0.00490162f $X=2.14 $Y=2.905 $X2=0
+ $Y2=0
cc_1022 N_A_27_74#_c_1612_n N_VPWR_M1032_d 0.00530362f $X=3.155 $Y=2.375 $X2=0
+ $Y2=0
cc_1023 N_A_27_74#_c_1616_n N_VPWR_M1005_s 0.00827001f $X=5.215 $Y=2.395 $X2=0
+ $Y2=0
cc_1024 N_A_27_74#_c_1616_n N_VPWR_M1003_s 0.00255417f $X=5.215 $Y=2.395 $X2=0
+ $Y2=0
cc_1025 N_A_27_74#_c_1601_n N_VPWR_M1003_s 0.0112943f $X=5.3 $Y=2.31 $X2=0 $Y2=0
cc_1026 N_A_27_74#_c_1738_p N_VPWR_M1003_s 0.00184106f $X=5.3 $Y=2.395 $X2=0
+ $Y2=0
cc_1027 N_A_27_74#_c_1607_n N_VPWR_c_1778_n 0.0105554f $X=0.28 $Y=2.75 $X2=0
+ $Y2=0
cc_1028 N_A_27_74#_c_1608_n N_VPWR_c_1778_n 0.017759f $X=1.375 $Y=2.375 $X2=0
+ $Y2=0
cc_1029 N_A_27_74#_c_1609_n N_VPWR_c_1778_n 0.0208967f $X=1.46 $Y=2.905 $X2=0
+ $Y2=0
cc_1030 N_A_27_74#_c_1611_n N_VPWR_c_1778_n 0.0146662f $X=1.545 $Y=2.99 $X2=0
+ $Y2=0
cc_1031 N_A_27_74#_c_1610_n N_VPWR_c_1779_n 0.0146323f $X=2.055 $Y=2.99 $X2=0
+ $Y2=0
cc_1032 N_A_27_74#_c_1646_n N_VPWR_c_1779_n 0.0205316f $X=2.14 $Y=2.905 $X2=0
+ $Y2=0
cc_1033 N_A_27_74#_c_1612_n N_VPWR_c_1779_n 0.0178153f $X=3.155 $Y=2.375 $X2=0
+ $Y2=0
cc_1034 N_A_27_74#_c_1614_n N_VPWR_c_1779_n 0.0100153f $X=3.32 $Y=2.73 $X2=0
+ $Y2=0
cc_1035 N_A_27_74#_c_1614_n N_VPWR_c_1780_n 0.0261435f $X=3.32 $Y=2.73 $X2=0
+ $Y2=0
cc_1036 N_A_27_74#_c_1616_n N_VPWR_c_1780_n 0.0215279f $X=5.215 $Y=2.395 $X2=0
+ $Y2=0
cc_1037 N_A_27_74#_c_1616_n N_VPWR_c_1781_n 0.00870407f $X=5.215 $Y=2.395 $X2=0
+ $Y2=0
cc_1038 N_A_27_74#_c_1677_n N_VPWR_c_1781_n 0.00100191f $X=5.605 $Y=2.395 $X2=0
+ $Y2=0
cc_1039 N_A_27_74#_c_1618_n N_VPWR_c_1781_n 0.0114906f $X=5.775 $Y=2.975 $X2=0
+ $Y2=0
cc_1040 N_A_27_74#_c_1738_p N_VPWR_c_1781_n 0.0129915f $X=5.3 $Y=2.395 $X2=0
+ $Y2=0
cc_1041 N_A_27_74#_c_1614_n N_VPWR_c_1786_n 0.0159746f $X=3.32 $Y=2.73 $X2=0
+ $Y2=0
cc_1042 N_A_27_74#_c_1607_n N_VPWR_c_1790_n 0.0159414f $X=0.28 $Y=2.75 $X2=0
+ $Y2=0
cc_1043 N_A_27_74#_c_1610_n N_VPWR_c_1791_n 0.0449818f $X=2.055 $Y=2.99 $X2=0
+ $Y2=0
cc_1044 N_A_27_74#_c_1611_n N_VPWR_c_1791_n 0.0121867f $X=1.545 $Y=2.99 $X2=0
+ $Y2=0
cc_1045 N_A_27_74#_c_1618_n N_VPWR_c_1792_n 0.0111306f $X=5.775 $Y=2.975 $X2=0
+ $Y2=0
cc_1046 N_A_27_74#_c_1619_n N_VPWR_c_1792_n 0.0391423f $X=6.28 $Y=2.975 $X2=0
+ $Y2=0
cc_1047 N_A_27_74#_M1011_s N_VPWR_c_1777_n 0.00257265f $X=6.135 $Y=2.54 $X2=0
+ $Y2=0
cc_1048 N_A_27_74#_c_1607_n N_VPWR_c_1777_n 0.0131581f $X=0.28 $Y=2.75 $X2=0
+ $Y2=0
cc_1049 N_A_27_74#_c_1610_n N_VPWR_c_1777_n 0.025776f $X=2.055 $Y=2.99 $X2=0
+ $Y2=0
cc_1050 N_A_27_74#_c_1611_n N_VPWR_c_1777_n 0.00660921f $X=1.545 $Y=2.99 $X2=0
+ $Y2=0
cc_1051 N_A_27_74#_c_1614_n N_VPWR_c_1777_n 0.0141401f $X=3.32 $Y=2.73 $X2=0
+ $Y2=0
cc_1052 N_A_27_74#_c_1616_n N_VPWR_c_1777_n 0.0426251f $X=5.215 $Y=2.395 $X2=0
+ $Y2=0
cc_1053 N_A_27_74#_c_1677_n N_VPWR_c_1777_n 0.00553357f $X=5.605 $Y=2.395 $X2=0
+ $Y2=0
cc_1054 N_A_27_74#_c_1618_n N_VPWR_c_1777_n 0.00656177f $X=5.775 $Y=2.975 $X2=0
+ $Y2=0
cc_1055 N_A_27_74#_c_1619_n N_VPWR_c_1777_n 0.0249596f $X=6.28 $Y=2.975 $X2=0
+ $Y2=0
cc_1056 N_A_27_74#_c_1738_p N_VPWR_c_1777_n 6.0606e-19 $X=5.3 $Y=2.395 $X2=0
+ $Y2=0
cc_1057 N_A_27_74#_c_1604_n N_VGND_c_1992_n 0.0107796f $X=0.435 $Y=0.585 $X2=0
+ $Y2=0
cc_1058 N_A_27_74#_c_1605_n N_VGND_c_1993_n 0.0148546f $X=3.46 $Y=0.58 $X2=0
+ $Y2=0
cc_1059 N_A_27_74#_c_1600_n N_VGND_c_1994_n 0.014793f $X=3.46 $Y=2.29 $X2=0
+ $Y2=0
cc_1060 N_A_27_74#_c_1605_n N_VGND_c_1994_n 0.0373981f $X=3.46 $Y=0.58 $X2=0
+ $Y2=0
cc_1061 N_A_27_74#_c_1605_n N_VGND_c_2002_n 0.0234711f $X=3.46 $Y=0.58 $X2=0
+ $Y2=0
cc_1062 N_A_27_74#_c_1604_n N_VGND_c_2006_n 0.0156682f $X=0.435 $Y=0.585 $X2=0
+ $Y2=0
cc_1063 N_A_27_74#_c_1604_n N_VGND_c_2012_n 0.0175747f $X=0.435 $Y=0.585 $X2=0
+ $Y2=0
cc_1064 N_A_27_74#_c_1605_n N_VGND_c_2012_n 0.0197338f $X=3.46 $Y=0.58 $X2=0
+ $Y2=0
cc_1065 N_VPWR_c_1785_n Q 0.0791681f $X=13.625 $Y=1.985 $X2=0 $Y2=0
cc_1066 N_VPWR_c_1784_n Q 0.004725f $X=12.115 $Y=2.49 $X2=0 $Y2=0
cc_1067 N_VPWR_c_1795_n Q 0.0183866f $X=13.54 $Y=3.33 $X2=0 $Y2=0
cc_1068 N_VPWR_c_1777_n Q 0.0151859f $X=14.16 $Y=3.33 $X2=0 $Y2=0
cc_1069 N_VPWR_c_1785_n N_Q_N_c_1975_n 0.0777954f $X=13.625 $Y=1.985 $X2=0 $Y2=0
cc_1070 N_VPWR_c_1796_n N_Q_N_c_1976_n 0.0144126f $X=14.16 $Y=3.33 $X2=0 $Y2=0
cc_1071 N_VPWR_c_1777_n N_Q_N_c_1976_n 0.0119295f $X=14.16 $Y=3.33 $X2=0 $Y2=0
cc_1072 Q_N N_VGND_c_1999_n 0.0296679f $X=14.075 $Y=0.47 $X2=0 $Y2=0
cc_1073 Q_N N_VGND_c_2011_n 0.0147163f $X=14.075 $Y=0.47 $X2=0 $Y2=0
cc_1074 Q_N N_VGND_c_2012_n 0.0130412f $X=14.075 $Y=0.47 $X2=0 $Y2=0
