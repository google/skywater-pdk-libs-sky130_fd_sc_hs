* File: sky130_fd_sc_hs__sedfxtp_1.pxi.spice
* Created: Tue Sep  1 20:24:33 2020
* 
x_PM_SKY130_FD_SC_HS__SEDFXTP_1%D N_D_c_329_n N_D_c_334_n N_D_c_335_n
+ N_D_M1037_g N_D_M1017_g N_D_c_331_n D D N_D_c_332_n N_D_c_333_n
+ PM_SKY130_FD_SC_HS__SEDFXTP_1%D
x_PM_SKY130_FD_SC_HS__SEDFXTP_1%A_159_404# N_A_159_404#_M1010_s
+ N_A_159_404#_M1036_s N_A_159_404#_c_381_n N_A_159_404#_M1023_g
+ N_A_159_404#_M1012_g N_A_159_404#_c_382_n N_A_159_404#_c_374_n
+ N_A_159_404#_c_375_n N_A_159_404#_c_376_n N_A_159_404#_c_377_n
+ N_A_159_404#_c_384_n N_A_159_404#_c_385_n N_A_159_404#_c_378_n
+ N_A_159_404#_c_386_n N_A_159_404#_c_387_n N_A_159_404#_c_379_n
+ N_A_159_404#_c_389_n N_A_159_404#_c_380_n
+ PM_SKY130_FD_SC_HS__SEDFXTP_1%A_159_404#
x_PM_SKY130_FD_SC_HS__SEDFXTP_1%DE N_DE_M1004_g N_DE_c_490_n N_DE_c_491_n
+ N_DE_c_492_n N_DE_c_498_n N_DE_M1036_g N_DE_c_493_n N_DE_M1010_g N_DE_c_499_n
+ N_DE_c_500_n N_DE_c_501_n N_DE_M1013_g N_DE_c_494_n DE N_DE_c_495_n
+ N_DE_c_502_n N_DE_c_496_n PM_SKY130_FD_SC_HS__SEDFXTP_1%DE
x_PM_SKY130_FD_SC_HS__SEDFXTP_1%A_547_301# N_A_547_301#_M1019_d
+ N_A_547_301#_M1005_d N_A_547_301#_M1038_g N_A_547_301#_c_592_n
+ N_A_547_301#_c_593_n N_A_547_301#_M1000_g N_A_547_301#_c_580_n
+ N_A_547_301#_M1035_g N_A_547_301#_c_581_n N_A_547_301#_c_582_n
+ N_A_547_301#_c_594_n N_A_547_301#_M1021_g N_A_547_301#_c_583_n
+ N_A_547_301#_c_596_n N_A_547_301#_c_597_n N_A_547_301#_c_598_n
+ N_A_547_301#_c_584_n N_A_547_301#_c_599_n N_A_547_301#_c_585_n
+ N_A_547_301#_c_586_n N_A_547_301#_c_587_n N_A_547_301#_c_588_n
+ N_A_547_301#_c_589_n N_A_547_301#_c_590_n N_A_547_301#_c_591_n
+ PM_SKY130_FD_SC_HS__SEDFXTP_1%A_547_301#
x_PM_SKY130_FD_SC_HS__SEDFXTP_1%A_639_85# N_A_639_85#_M1041_s
+ N_A_639_85#_M1027_s N_A_639_85#_c_817_n N_A_639_85#_M1025_g
+ N_A_639_85#_c_818_n N_A_639_85#_c_819_n N_A_639_85#_c_828_n
+ N_A_639_85#_M1002_g N_A_639_85#_c_820_n N_A_639_85#_c_829_n
+ N_A_639_85#_c_821_n N_A_639_85#_c_822_n N_A_639_85#_c_823_n
+ N_A_639_85#_c_824_n N_A_639_85#_c_832_n N_A_639_85#_c_833_n
+ N_A_639_85#_c_825_n N_A_639_85#_c_826_n N_A_639_85#_c_827_n
+ N_A_639_85#_c_835_n N_A_639_85#_c_836_n
+ PM_SKY130_FD_SC_HS__SEDFXTP_1%A_639_85#
x_PM_SKY130_FD_SC_HS__SEDFXTP_1%SCD N_SCD_M1031_g N_SCD_c_934_n N_SCD_c_935_n
+ N_SCD_M1016_g SCD N_SCD_c_933_n PM_SKY130_FD_SC_HS__SEDFXTP_1%SCD
x_PM_SKY130_FD_SC_HS__SEDFXTP_1%SCE N_SCE_c_984_n N_SCE_M1008_g N_SCE_c_985_n
+ N_SCE_c_986_n N_SCE_c_977_n N_SCE_c_988_n N_SCE_M1027_g N_SCE_M1041_g
+ N_SCE_c_979_n N_SCE_c_980_n N_SCE_M1028_g SCE N_SCE_c_983_n
+ PM_SKY130_FD_SC_HS__SEDFXTP_1%SCE
x_PM_SKY130_FD_SC_HS__SEDFXTP_1%CLK N_CLK_c_1063_n N_CLK_M1018_g N_CLK_c_1064_n
+ N_CLK_M1020_g CLK PM_SKY130_FD_SC_HS__SEDFXTP_1%CLK
x_PM_SKY130_FD_SC_HS__SEDFXTP_1%A_1492_74# N_A_1492_74#_M1007_d
+ N_A_1492_74#_M1030_d N_A_1492_74#_c_1120_n N_A_1492_74#_M1015_g
+ N_A_1492_74#_c_1096_n N_A_1492_74#_M1032_g N_A_1492_74#_M1024_g
+ N_A_1492_74#_c_1098_n N_A_1492_74#_c_1122_n N_A_1492_74#_M1040_g
+ N_A_1492_74#_c_1099_n N_A_1492_74#_c_1100_n N_A_1492_74#_c_1101_n
+ N_A_1492_74#_c_1123_n N_A_1492_74#_c_1102_n N_A_1492_74#_c_1103_n
+ N_A_1492_74#_c_1104_n N_A_1492_74#_c_1105_n N_A_1492_74#_c_1106_n
+ N_A_1492_74#_c_1107_n N_A_1492_74#_c_1202_p N_A_1492_74#_c_1108_n
+ N_A_1492_74#_c_1109_n N_A_1492_74#_c_1110_n N_A_1492_74#_c_1111_n
+ N_A_1492_74#_c_1112_n N_A_1492_74#_c_1113_n N_A_1492_74#_c_1114_n
+ N_A_1492_74#_c_1115_n N_A_1492_74#_c_1116_n N_A_1492_74#_c_1117_n
+ N_A_1492_74#_c_1127_n N_A_1492_74#_c_1239_p N_A_1492_74#_c_1118_n
+ N_A_1492_74#_c_1119_n PM_SKY130_FD_SC_HS__SEDFXTP_1%A_1492_74#
x_PM_SKY130_FD_SC_HS__SEDFXTP_1%A_1295_74# N_A_1295_74#_M1018_d
+ N_A_1295_74#_M1020_d N_A_1295_74#_M1007_g N_A_1295_74#_c_1330_n
+ N_A_1295_74#_c_1344_n N_A_1295_74#_M1030_g N_A_1295_74#_c_1331_n
+ N_A_1295_74#_M1026_g N_A_1295_74#_c_1333_n N_A_1295_74#_c_1347_n
+ N_A_1295_74#_c_1348_n N_A_1295_74#_M1014_g N_A_1295_74#_c_1334_n
+ N_A_1295_74#_M1001_g N_A_1295_74#_M1034_g N_A_1295_74#_c_1336_n
+ N_A_1295_74#_c_1337_n N_A_1295_74#_c_1338_n N_A_1295_74#_c_1339_n
+ N_A_1295_74#_c_1340_n N_A_1295_74#_c_1354_n N_A_1295_74#_c_1355_n
+ N_A_1295_74#_c_1356_n N_A_1295_74#_c_1357_n N_A_1295_74#_c_1358_n
+ N_A_1295_74#_c_1359_n N_A_1295_74#_c_1360_n N_A_1295_74#_c_1341_n
+ N_A_1295_74#_c_1361_n N_A_1295_74#_c_1342_n
+ PM_SKY130_FD_SC_HS__SEDFXTP_1%A_1295_74#
x_PM_SKY130_FD_SC_HS__SEDFXTP_1%A_1910_71# N_A_1910_71#_M1033_d
+ N_A_1910_71#_M1039_d N_A_1910_71#_M1029_g N_A_1910_71#_c_1530_n
+ N_A_1910_71#_c_1543_n N_A_1910_71#_M1003_g N_A_1910_71#_c_1531_n
+ N_A_1910_71#_c_1545_n N_A_1910_71#_M1009_g N_A_1910_71#_c_1532_n
+ N_A_1910_71#_M1022_g N_A_1910_71#_c_1533_n N_A_1910_71#_c_1534_n
+ N_A_1910_71#_c_1535_n N_A_1910_71#_c_1536_n N_A_1910_71#_c_1537_n
+ N_A_1910_71#_c_1538_n N_A_1910_71#_c_1539_n N_A_1910_71#_c_1547_n
+ N_A_1910_71#_c_1540_n N_A_1910_71#_c_1541_n
+ PM_SKY130_FD_SC_HS__SEDFXTP_1%A_1910_71#
x_PM_SKY130_FD_SC_HS__SEDFXTP_1%A_1688_97# N_A_1688_97#_M1026_d
+ N_A_1688_97#_M1015_d N_A_1688_97#_c_1642_n N_A_1688_97#_M1039_g
+ N_A_1688_97#_M1033_g N_A_1688_97#_c_1644_n N_A_1688_97#_c_1648_n
+ N_A_1688_97#_c_1649_n N_A_1688_97#_c_1650_n N_A_1688_97#_c_1651_n
+ N_A_1688_97#_c_1645_n N_A_1688_97#_c_1646_n
+ PM_SKY130_FD_SC_HS__SEDFXTP_1%A_1688_97#
x_PM_SKY130_FD_SC_HS__SEDFXTP_1%A_2385_74# N_A_2385_74#_M1024_d
+ N_A_2385_74#_M1001_d N_A_2385_74#_M1019_g N_A_2385_74#_c_1741_n
+ N_A_2385_74#_c_1752_n N_A_2385_74#_M1005_g N_A_2385_74#_c_1742_n
+ N_A_2385_74#_c_1743_n N_A_2385_74#_c_1744_n N_A_2385_74#_M1006_g
+ N_A_2385_74#_c_1753_n N_A_2385_74#_M1011_g N_A_2385_74#_c_1745_n
+ N_A_2385_74#_c_1825_n N_A_2385_74#_c_1746_n N_A_2385_74#_c_1747_n
+ N_A_2385_74#_c_1755_n N_A_2385_74#_c_1756_n N_A_2385_74#_c_1757_n
+ N_A_2385_74#_c_1748_n N_A_2385_74#_c_1759_n N_A_2385_74#_c_1749_n
+ N_A_2385_74#_c_1761_n N_A_2385_74#_c_1750_n
+ PM_SKY130_FD_SC_HS__SEDFXTP_1%A_2385_74#
x_PM_SKY130_FD_SC_HS__SEDFXTP_1%A_27_74# N_A_27_74#_M1017_s N_A_27_74#_M1038_d
+ N_A_27_74#_M1037_s N_A_27_74#_M1000_d N_A_27_74#_c_1884_n N_A_27_74#_c_1890_n
+ N_A_27_74#_c_1891_n N_A_27_74#_c_1892_n N_A_27_74#_c_1893_n
+ N_A_27_74#_c_1894_n N_A_27_74#_c_1925_n N_A_27_74#_c_1895_n
+ N_A_27_74#_c_1896_n N_A_27_74#_c_1885_n N_A_27_74#_c_1897_n
+ N_A_27_74#_c_1886_n N_A_27_74#_c_1887_n N_A_27_74#_c_1899_n
+ N_A_27_74#_c_1888_n N_A_27_74#_c_1900_n PM_SKY130_FD_SC_HS__SEDFXTP_1%A_27_74#
x_PM_SKY130_FD_SC_HS__SEDFXTP_1%VPWR N_VPWR_M1023_d N_VPWR_M1036_d
+ N_VPWR_M1027_d N_VPWR_M1020_s N_VPWR_M1030_s N_VPWR_M1003_d N_VPWR_M1009_s
+ N_VPWR_M1021_d N_VPWR_M1011_d N_VPWR_c_2008_n N_VPWR_c_2009_n N_VPWR_c_2010_n
+ N_VPWR_c_2011_n N_VPWR_c_2012_n N_VPWR_c_2013_n N_VPWR_c_2014_n
+ N_VPWR_c_2015_n N_VPWR_c_2016_n N_VPWR_c_2017_n N_VPWR_c_2018_n
+ N_VPWR_c_2019_n N_VPWR_c_2020_n N_VPWR_c_2021_n N_VPWR_c_2022_n
+ N_VPWR_c_2023_n N_VPWR_c_2024_n N_VPWR_c_2025_n N_VPWR_c_2026_n
+ N_VPWR_c_2027_n VPWR N_VPWR_c_2028_n N_VPWR_c_2029_n N_VPWR_c_2030_n
+ N_VPWR_c_2031_n N_VPWR_c_2032_n N_VPWR_c_2033_n N_VPWR_c_2034_n
+ N_VPWR_c_2007_n PM_SKY130_FD_SC_HS__SEDFXTP_1%VPWR
x_PM_SKY130_FD_SC_HS__SEDFXTP_1%A_669_111# N_A_669_111#_M1025_d
+ N_A_669_111#_M1028_d N_A_669_111#_M1026_s N_A_669_111#_M1008_d
+ N_A_669_111#_M1002_d N_A_669_111#_M1015_s N_A_669_111#_c_2178_n
+ N_A_669_111#_c_2249_n N_A_669_111#_c_2179_n N_A_669_111#_c_2191_n
+ N_A_669_111#_c_2209_n N_A_669_111#_c_2180_n N_A_669_111#_c_2169_n
+ N_A_669_111#_c_2170_n N_A_669_111#_c_2171_n N_A_669_111#_c_2172_n
+ N_A_669_111#_c_2182_n N_A_669_111#_c_2183_n N_A_669_111#_c_2173_n
+ N_A_669_111#_c_2174_n N_A_669_111#_c_2199_n N_A_669_111#_c_2175_n
+ N_A_669_111#_c_2282_n N_A_669_111#_c_2184_n N_A_669_111#_c_2185_n
+ N_A_669_111#_c_2176_n N_A_669_111#_c_2177_n N_A_669_111#_c_2187_n
+ N_A_669_111#_c_2188_n N_A_669_111#_c_2189_n N_A_669_111#_c_2351_n
+ PM_SKY130_FD_SC_HS__SEDFXTP_1%A_669_111#
x_PM_SKY130_FD_SC_HS__SEDFXTP_1%Q N_Q_M1006_s N_Q_M1011_s Q Q Q Q Q Q Q
+ PM_SKY130_FD_SC_HS__SEDFXTP_1%Q
x_PM_SKY130_FD_SC_HS__SEDFXTP_1%VGND N_VGND_M1004_d N_VGND_M1010_d
+ N_VGND_M1041_d N_VGND_M1018_s N_VGND_M1007_s N_VGND_M1029_d N_VGND_M1022_s
+ N_VGND_M1035_d N_VGND_M1006_d N_VGND_c_2387_n N_VGND_c_2388_n N_VGND_c_2389_n
+ N_VGND_c_2390_n N_VGND_c_2391_n N_VGND_c_2392_n N_VGND_c_2393_n
+ N_VGND_c_2394_n N_VGND_c_2395_n N_VGND_c_2396_n N_VGND_c_2397_n
+ N_VGND_c_2398_n N_VGND_c_2399_n N_VGND_c_2400_n N_VGND_c_2401_n VGND
+ N_VGND_c_2402_n N_VGND_c_2403_n N_VGND_c_2404_n N_VGND_c_2405_n
+ N_VGND_c_2406_n N_VGND_c_2407_n N_VGND_c_2408_n N_VGND_c_2409_n
+ N_VGND_c_2410_n N_VGND_c_2411_n N_VGND_c_2412_n N_VGND_c_2413_n
+ PM_SKY130_FD_SC_HS__SEDFXTP_1%VGND
cc_1 VNB N_D_c_329_n 0.0261273f $X=-0.19 $Y=-0.245 $X2=0.575 $Y2=1.61
cc_2 VNB N_D_M1017_g 0.0339978f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=0.58
cc_3 VNB N_D_c_331_n 0.00355983f $X=-0.19 $Y=-0.245 $X2=0.575 $Y2=1.78
cc_4 VNB N_D_c_332_n 0.0188363f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=1.275
cc_5 VNB N_D_c_333_n 0.00936403f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=1.275
cc_6 VNB N_A_159_404#_M1012_g 0.0413951f $X=-0.19 $Y=-0.245 $X2=0.575 $Y2=1.78
cc_7 VNB N_A_159_404#_c_374_n 0.00358262f $X=-0.19 $Y=-0.245 $X2=0.575 $Y2=1.11
cc_8 VNB N_A_159_404#_c_375_n 0.0190364f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=1.275
cc_9 VNB N_A_159_404#_c_376_n 0.0112302f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_159_404#_c_377_n 0.00187438f $X=-0.19 $Y=-0.245 $X2=0.615
+ $Y2=1.295
cc_11 VNB N_A_159_404#_c_378_n 0.00794325f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_159_404#_c_379_n 0.00469829f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_159_404#_c_380_n 0.0196188f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_DE_M1004_g 0.0290737f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.78
cc_15 VNB N_DE_c_490_n 0.0277406f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.245
cc_16 VNB N_DE_c_491_n 0.00761418f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.64
cc_17 VNB N_DE_c_492_n 3.94837e-19 $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=0.58
cc_18 VNB N_DE_c_493_n 0.0158343f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_19 VNB N_DE_c_494_n 0.0340384f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=1.295
cc_20 VNB N_DE_c_495_n 0.0244846f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_DE_c_496_n 0.0164531f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_547_301#_M1038_g 0.0398126f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=0.58
cc_23 VNB N_A_547_301#_c_580_n 0.0170882f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_547_301#_c_581_n 0.0378978f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=1.275
cc_25 VNB N_A_547_301#_c_582_n 0.00715985f $X=-0.19 $Y=-0.245 $X2=0.575 $Y2=1.11
cc_26 VNB N_A_547_301#_c_583_n 0.034466f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=1.665
cc_27 VNB N_A_547_301#_c_584_n 0.00952178f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_547_301#_c_585_n 0.0787936f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_547_301#_c_586_n 0.00111649f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_547_301#_c_587_n 3.13795e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_547_301#_c_588_n 3.48754e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_547_301#_c_589_n 0.00740414f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_547_301#_c_590_n 0.0212294f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_547_301#_c_591_n 0.007854f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_639_85#_c_817_n 0.0159586f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.64
cc_36 VNB N_A_639_85#_c_818_n 0.0316995f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=0.58
cc_37 VNB N_A_639_85#_c_819_n 0.00865069f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_639_85#_c_820_n 0.00772331f $X=-0.19 $Y=-0.245 $X2=0.575 $Y2=1.275
cc_39 VNB N_A_639_85#_c_821_n 0.00576423f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=1.275
cc_40 VNB N_A_639_85#_c_822_n 0.074433f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_639_85#_c_823_n 0.00606184f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_639_85#_c_824_n 0.0328354f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_639_85#_c_825_n 0.00307366f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_639_85#_c_826_n 0.02808f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_A_639_85#_c_827_n 0.00639732f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_SCD_M1031_g 0.0287203f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.78
cc_47 VNB SCD 0.0174228f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=0.58
cc_48 VNB N_SCD_c_933_n 0.0207883f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_49 VNB N_SCE_c_977_n 0.00811558f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.64
cc_50 VNB N_SCE_M1041_g 0.0308745f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_SCE_c_979_n 0.0565784f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_SCE_c_980_n 0.012806f $X=-0.19 $Y=-0.245 $X2=0.575 $Y2=1.275
cc_53 VNB N_SCE_M1028_g 0.0390656f $X=-0.19 $Y=-0.245 $X2=0.575 $Y2=1.11
cc_54 VNB SCE 0.00391934f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_SCE_c_983_n 0.0326445f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=1.665
cc_56 VNB N_CLK_c_1063_n 0.0207827f $X=-0.19 $Y=-0.245 $X2=0.575 $Y2=1.28
cc_57 VNB N_CLK_c_1064_n 0.0433052f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.155
cc_58 VNB CLK 0.00360057f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.64
cc_59 VNB N_A_1492_74#_c_1096_n 0.0183029f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=0.58
cc_60 VNB N_A_1492_74#_M1024_g 0.0349335f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_A_1492_74#_c_1098_n 0.00527446f $X=-0.19 $Y=-0.245 $X2=0.58
+ $Y2=1.275
cc_62 VNB N_A_1492_74#_c_1099_n 0.00932933f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_A_1492_74#_c_1100_n 0.0184356f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_A_1492_74#_c_1101_n 0.00362036f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_A_1492_74#_c_1102_n 0.00587229f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_A_1492_74#_c_1103_n 0.01738f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_A_1492_74#_c_1104_n 5.57375e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_A_1492_74#_c_1105_n 0.00159984f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_A_1492_74#_c_1106_n 0.0392354f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_A_1492_74#_c_1107_n 0.00807263f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_A_1492_74#_c_1108_n 0.00904398f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_A_1492_74#_c_1109_n 0.00203f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_A_1492_74#_c_1110_n 0.00961154f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_A_1492_74#_c_1111_n 0.00471223f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_A_1492_74#_c_1112_n 0.00314294f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_A_1492_74#_c_1113_n 0.0028814f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_A_1492_74#_c_1114_n 0.00305718f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_A_1492_74#_c_1115_n 0.0165047f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VNB N_A_1492_74#_c_1116_n 0.0116007f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_A_1492_74#_c_1117_n 0.00123754f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_81 VNB N_A_1492_74#_c_1118_n 0.00398359f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_82 VNB N_A_1492_74#_c_1119_n 0.030036f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_83 VNB N_A_1295_74#_M1007_g 0.0496814f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=0.58
cc_84 VNB N_A_1295_74#_c_1330_n 0.00990377f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_85 VNB N_A_1295_74#_c_1331_n 0.00787256f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_86 VNB N_A_1295_74#_M1026_g 0.0561689f $X=-0.19 $Y=-0.245 $X2=0.575 $Y2=1.11
cc_87 VNB N_A_1295_74#_c_1333_n 0.026052f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_88 VNB N_A_1295_74#_c_1334_n 0.0179088f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_89 VNB N_A_1295_74#_M1034_g 0.0484177f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_90 VNB N_A_1295_74#_c_1336_n 0.00962966f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_91 VNB N_A_1295_74#_c_1337_n 0.00499721f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_92 VNB N_A_1295_74#_c_1338_n 7.16371e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_93 VNB N_A_1295_74#_c_1339_n 0.00817988f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_94 VNB N_A_1295_74#_c_1340_n 0.0147857f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_95 VNB N_A_1295_74#_c_1341_n 0.00882492f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_96 VNB N_A_1295_74#_c_1342_n 0.00402307f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_97 VNB N_A_1910_71#_M1029_g 0.0275892f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=0.58
cc_98 VNB N_A_1910_71#_c_1530_n 0.0127731f $X=-0.19 $Y=-0.245 $X2=0.575 $Y2=1.78
cc_99 VNB N_A_1910_71#_c_1531_n 0.00843181f $X=-0.19 $Y=-0.245 $X2=0.58
+ $Y2=1.275
cc_100 VNB N_A_1910_71#_c_1532_n 0.0197313f $X=-0.19 $Y=-0.245 $X2=0.615
+ $Y2=1.295
cc_101 VNB N_A_1910_71#_c_1533_n 0.00940458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_102 VNB N_A_1910_71#_c_1534_n 0.0054522f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_103 VNB N_A_1910_71#_c_1535_n 0.00231007f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_104 VNB N_A_1910_71#_c_1536_n 0.00461404f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_105 VNB N_A_1910_71#_c_1537_n 0.00180512f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_106 VNB N_A_1910_71#_c_1538_n 0.0576016f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_107 VNB N_A_1910_71#_c_1539_n 0.00107588f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_108 VNB N_A_1910_71#_c_1540_n 0.0354176f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_109 VNB N_A_1910_71#_c_1541_n 0.0286377f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_110 VNB N_A_1688_97#_c_1642_n 0.0163425f $X=-0.19 $Y=-0.245 $X2=0.495
+ $Y2=2.64
cc_111 VNB N_A_1688_97#_M1033_g 0.0419527f $X=-0.19 $Y=-0.245 $X2=0.575 $Y2=1.78
cc_112 VNB N_A_1688_97#_c_1644_n 0.0160612f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_113 VNB N_A_1688_97#_c_1645_n 0.00173865f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_114 VNB N_A_1688_97#_c_1646_n 0.00375455f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_115 VNB N_A_2385_74#_M1019_g 0.0321574f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=0.58
cc_116 VNB N_A_2385_74#_c_1741_n 0.00281699f $X=-0.19 $Y=-0.245 $X2=0.575
+ $Y2=1.78
cc_117 VNB N_A_2385_74#_c_1742_n 0.0865631f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_118 VNB N_A_2385_74#_c_1743_n 0.0449607f $X=-0.19 $Y=-0.245 $X2=0.575
+ $Y2=1.275
cc_119 VNB N_A_2385_74#_c_1744_n 0.0260131f $X=-0.19 $Y=-0.245 $X2=0.58
+ $Y2=1.275
cc_120 VNB N_A_2385_74#_c_1745_n 0.034067f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_121 VNB N_A_2385_74#_c_1746_n 0.00286498f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_122 VNB N_A_2385_74#_c_1747_n 0.0035576f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_123 VNB N_A_2385_74#_c_1748_n 0.00756009f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_124 VNB N_A_2385_74#_c_1749_n 0.00394269f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_125 VNB N_A_2385_74#_c_1750_n 0.00399884f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_126 VNB N_A_27_74#_c_1884_n 0.0412306f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_127 VNB N_A_27_74#_c_1885_n 0.00379155f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_128 VNB N_A_27_74#_c_1886_n 0.0065331f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_129 VNB N_A_27_74#_c_1887_n 0.0216354f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_130 VNB N_A_27_74#_c_1888_n 0.00390083f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_131 VNB N_VPWR_c_2007_n 0.641339f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_132 VNB N_A_669_111#_c_2169_n 0.00908825f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_133 VNB N_A_669_111#_c_2170_n 0.0135895f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_134 VNB N_A_669_111#_c_2171_n 0.00322709f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_135 VNB N_A_669_111#_c_2172_n 0.0114953f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_136 VNB N_A_669_111#_c_2173_n 0.00737783f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_137 VNB N_A_669_111#_c_2174_n 0.00417594f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_138 VNB N_A_669_111#_c_2175_n 0.0175669f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_139 VNB N_A_669_111#_c_2176_n 0.00888231f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_140 VNB N_A_669_111#_c_2177_n 0.00806826f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_141 VNB Q 0.0104501f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.64
cc_142 VNB N_VGND_c_2387_n 0.013355f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_143 VNB N_VGND_c_2388_n 0.0180526f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_144 VNB N_VGND_c_2389_n 0.00683062f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_145 VNB N_VGND_c_2390_n 0.0158101f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_146 VNB N_VGND_c_2391_n 0.0103972f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_147 VNB N_VGND_c_2392_n 0.0105613f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_148 VNB N_VGND_c_2393_n 0.00590394f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_149 VNB N_VGND_c_2394_n 0.010678f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_150 VNB N_VGND_c_2395_n 0.0505973f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_151 VNB N_VGND_c_2396_n 0.0655119f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_152 VNB N_VGND_c_2397_n 0.00332923f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_153 VNB N_VGND_c_2398_n 0.029639f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_154 VNB N_VGND_c_2399_n 0.00500104f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_155 VNB N_VGND_c_2400_n 0.020445f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_156 VNB N_VGND_c_2401_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_157 VNB N_VGND_c_2402_n 0.0333036f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_158 VNB N_VGND_c_2403_n 0.0195928f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_159 VNB N_VGND_c_2404_n 0.0602803f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_160 VNB N_VGND_c_2405_n 0.0296519f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_161 VNB N_VGND_c_2406_n 0.0339585f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_162 VNB N_VGND_c_2407_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_163 VNB N_VGND_c_2408_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_164 VNB N_VGND_c_2409_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_165 VNB N_VGND_c_2410_n 0.00461913f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_166 VNB N_VGND_c_2411_n 0.0403351f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_167 VNB N_VGND_c_2412_n 0.0313022f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_168 VNB N_VGND_c_2413_n 0.835548f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_169 VPB N_D_c_334_n 0.023206f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=2.155
cc_170 VPB N_D_c_335_n 0.0251378f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=2.245
cc_171 VPB N_D_c_331_n 0.01311f $X=-0.19 $Y=1.66 $X2=0.575 $Y2=1.78
cc_172 VPB N_D_c_333_n 0.00398042f $X=-0.19 $Y=1.66 $X2=0.58 $Y2=1.275
cc_173 VPB N_A_159_404#_c_381_n 0.0181955f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=2.64
cc_174 VPB N_A_159_404#_c_382_n 0.0368589f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_175 VPB N_A_159_404#_c_375_n 0.0274972f $X=-0.19 $Y=1.66 $X2=0.615 $Y2=1.275
cc_176 VPB N_A_159_404#_c_384_n 0.0147373f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_177 VPB N_A_159_404#_c_385_n 0.00263747f $X=-0.19 $Y=1.66 $X2=0.615 $Y2=1.665
cc_178 VPB N_A_159_404#_c_386_n 0.00254697f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_179 VPB N_A_159_404#_c_387_n 0.00845557f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_180 VPB N_A_159_404#_c_379_n 0.00260289f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_181 VPB N_A_159_404#_c_389_n 0.00145276f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_182 VPB N_A_159_404#_c_380_n 0.0218988f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_183 VPB N_DE_c_492_n 0.0236903f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=0.58
cc_184 VPB N_DE_c_498_n 0.0183363f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_185 VPB N_DE_c_499_n 0.0342754f $X=-0.19 $Y=1.66 $X2=0.575 $Y2=1.275
cc_186 VPB N_DE_c_500_n 0.0263402f $X=-0.19 $Y=1.66 $X2=0.58 $Y2=1.275
cc_187 VPB N_DE_c_501_n 0.0161255f $X=-0.19 $Y=1.66 $X2=0.58 $Y2=1.275
cc_188 VPB N_DE_c_502_n 0.00316831f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_189 VPB N_A_547_301#_c_592_n 0.0222841f $X=-0.19 $Y=1.66 $X2=0.575 $Y2=1.78
cc_190 VPB N_A_547_301#_c_593_n 0.0212328f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.21
cc_191 VPB N_A_547_301#_c_594_n 0.0564056f $X=-0.19 $Y=1.66 $X2=0.615 $Y2=1.275
cc_192 VPB N_A_547_301#_c_583_n 0.0215025f $X=-0.19 $Y=1.66 $X2=0.615 $Y2=1.665
cc_193 VPB N_A_547_301#_c_596_n 0.00747546f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_194 VPB N_A_547_301#_c_597_n 0.00813529f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_195 VPB N_A_547_301#_c_598_n 0.0072007f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_196 VPB N_A_547_301#_c_599_n 0.00382486f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_197 VPB N_A_547_301#_c_585_n 0.0492038f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_198 VPB N_A_547_301#_c_586_n 3.27019e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_199 VPB N_A_547_301#_c_587_n 0.00230607f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_200 VPB N_A_547_301#_c_589_n 0.00235438f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_201 VPB N_A_547_301#_c_590_n 0.0222105f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_202 VPB N_A_639_85#_c_828_n 0.0162092f $X=-0.19 $Y=1.66 $X2=0.575 $Y2=1.78
cc_203 VPB N_A_639_85#_c_829_n 0.0232862f $X=-0.19 $Y=1.66 $X2=0.58 $Y2=1.275
cc_204 VPB N_A_639_85#_c_823_n 0.0028825f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_205 VPB N_A_639_85#_c_824_n 0.0325706f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_206 VPB N_A_639_85#_c_832_n 0.00466068f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_207 VPB N_A_639_85#_c_833_n 0.0218649f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_208 VPB N_A_639_85#_c_826_n 0.0200498f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_209 VPB N_A_639_85#_c_835_n 0.00579469f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_210 VPB N_A_639_85#_c_836_n 0.00833187f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_211 VPB N_SCD_c_934_n 0.0204059f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=2.64
cc_212 VPB N_SCD_c_935_n 0.0215923f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=2.64
cc_213 VPB SCD 0.00271418f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=0.58
cc_214 VPB N_SCD_c_933_n 0.00959317f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.21
cc_215 VPB N_SCE_c_984_n 0.0185503f $X=-0.19 $Y=1.66 $X2=0.575 $Y2=1.28
cc_216 VPB N_SCE_c_985_n 0.0805259f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=2.155
cc_217 VPB N_SCE_c_986_n 0.0132883f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=2.245
cc_218 VPB N_SCE_c_977_n 0.0278252f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=2.64
cc_219 VPB N_SCE_c_988_n 0.00745008f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.11
cc_220 VPB N_SCE_M1027_g 0.00949617f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_221 VPB N_CLK_c_1064_n 0.0282333f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=2.155
cc_222 VPB N_A_1492_74#_c_1120_n 0.0202275f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=2.64
cc_223 VPB N_A_1492_74#_c_1098_n 0.0373999f $X=-0.19 $Y=1.66 $X2=0.58 $Y2=1.275
cc_224 VPB N_A_1492_74#_c_1122_n 0.0219866f $X=-0.19 $Y=1.66 $X2=0.58 $Y2=1.275
cc_225 VPB N_A_1492_74#_c_1123_n 0.0116938f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_226 VPB N_A_1492_74#_c_1102_n 0.00103576f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_227 VPB N_A_1492_74#_c_1114_n 0.00647556f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_228 VPB N_A_1492_74#_c_1115_n 0.01808f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_229 VPB N_A_1492_74#_c_1127_n 0.0562983f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_230 VPB N_A_1295_74#_c_1330_n 0.0118008f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_231 VPB N_A_1295_74#_c_1344_n 0.0210946f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.21
cc_232 VPB N_A_1295_74#_c_1331_n 0.00858255f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_233 VPB N_A_1295_74#_c_1333_n 0.0236102f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_234 VPB N_A_1295_74#_c_1347_n 0.00967628f $X=-0.19 $Y=1.66 $X2=0.615
+ $Y2=1.665
cc_235 VPB N_A_1295_74#_c_1348_n 0.0592091f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_236 VPB N_A_1295_74#_c_1334_n 0.0412617f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_237 VPB N_A_1295_74#_c_1336_n 0.00811031f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_238 VPB N_A_1295_74#_c_1337_n 0.00167153f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_239 VPB N_A_1295_74#_c_1338_n 0.00489057f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_240 VPB N_A_1295_74#_c_1340_n 0.00390172f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_241 VPB N_A_1295_74#_c_1354_n 0.00377732f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_242 VPB N_A_1295_74#_c_1355_n 0.0374691f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_243 VPB N_A_1295_74#_c_1356_n 0.00553717f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_244 VPB N_A_1295_74#_c_1357_n 0.00264345f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_245 VPB N_A_1295_74#_c_1358_n 0.0141068f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_246 VPB N_A_1295_74#_c_1359_n 0.00103733f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_247 VPB N_A_1295_74#_c_1360_n 0.00271783f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_248 VPB N_A_1295_74#_c_1361_n 0.00410269f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_249 VPB N_A_1295_74#_c_1342_n 0.00120704f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_250 VPB N_A_1910_71#_c_1530_n 0.0406498f $X=-0.19 $Y=1.66 $X2=0.575 $Y2=1.78
cc_251 VPB N_A_1910_71#_c_1543_n 0.0218546f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.21
cc_252 VPB N_A_1910_71#_c_1531_n 0.00843705f $X=-0.19 $Y=1.66 $X2=0.58 $Y2=1.275
cc_253 VPB N_A_1910_71#_c_1545_n 0.0301608f $X=-0.19 $Y=1.66 $X2=0.575 $Y2=1.11
cc_254 VPB N_A_1910_71#_c_1535_n 0.00811658f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_255 VPB N_A_1910_71#_c_1547_n 0.00827933f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_256 VPB N_A_1688_97#_c_1642_n 0.0409392f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=2.64
cc_257 VPB N_A_1688_97#_c_1648_n 0.00288391f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_258 VPB N_A_1688_97#_c_1649_n 0.00147601f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_259 VPB N_A_1688_97#_c_1650_n 0.00837991f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_260 VPB N_A_1688_97#_c_1651_n 0.00281594f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_261 VPB N_A_1688_97#_c_1645_n 8.10289e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_262 VPB N_A_1688_97#_c_1646_n 0.00971417f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_263 VPB N_A_2385_74#_c_1741_n 0.0327476f $X=-0.19 $Y=1.66 $X2=0.575 $Y2=1.78
cc_264 VPB N_A_2385_74#_c_1752_n 0.0276311f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.21
cc_265 VPB N_A_2385_74#_c_1753_n 0.0218963f $X=-0.19 $Y=1.66 $X2=0.615 $Y2=1.275
cc_266 VPB N_A_2385_74#_c_1745_n 0.0112814f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_267 VPB N_A_2385_74#_c_1755_n 0.00508324f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_268 VPB N_A_2385_74#_c_1756_n 0.00304367f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_269 VPB N_A_2385_74#_c_1757_n 0.0102729f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_270 VPB N_A_2385_74#_c_1748_n 9.47506e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_271 VPB N_A_2385_74#_c_1759_n 0.00879642f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_272 VPB N_A_2385_74#_c_1749_n 0.00118718f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_273 VPB N_A_2385_74#_c_1761_n 2.36926e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_274 VPB N_A_27_74#_c_1884_n 0.0308767f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_275 VPB N_A_27_74#_c_1890_n 0.0233575f $X=-0.19 $Y=1.66 $X2=0.575 $Y2=1.275
cc_276 VPB N_A_27_74#_c_1891_n 0.0136238f $X=-0.19 $Y=1.66 $X2=0.58 $Y2=1.275
cc_277 VPB N_A_27_74#_c_1892_n 0.00998336f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_278 VPB N_A_27_74#_c_1893_n 0.00955076f $X=-0.19 $Y=1.66 $X2=0.615 $Y2=1.295
cc_279 VPB N_A_27_74#_c_1894_n 0.00349119f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_280 VPB N_A_27_74#_c_1895_n 0.00557118f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_281 VPB N_A_27_74#_c_1896_n 8.44548e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_282 VPB N_A_27_74#_c_1897_n 0.00216571f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_283 VPB N_A_27_74#_c_1886_n 0.0123983f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_284 VPB N_A_27_74#_c_1899_n 0.0136359f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_285 VPB N_A_27_74#_c_1900_n 0.00125429f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_286 VPB N_VPWR_c_2008_n 0.00600898f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_287 VPB N_VPWR_c_2009_n 0.00554607f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_288 VPB N_VPWR_c_2010_n 0.00745483f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_289 VPB N_VPWR_c_2011_n 0.0137442f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_290 VPB N_VPWR_c_2012_n 0.0216876f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_291 VPB N_VPWR_c_2013_n 0.0115296f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_292 VPB N_VPWR_c_2014_n 0.0140087f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_293 VPB N_VPWR_c_2015_n 0.0112438f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_294 VPB N_VPWR_c_2016_n 0.0103331f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_295 VPB N_VPWR_c_2017_n 0.0649859f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_296 VPB N_VPWR_c_2018_n 0.0293385f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_297 VPB N_VPWR_c_2019_n 0.00460249f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_298 VPB N_VPWR_c_2020_n 0.0296515f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_299 VPB N_VPWR_c_2021_n 0.00463855f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_300 VPB N_VPWR_c_2022_n 0.0323948f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_301 VPB N_VPWR_c_2023_n 0.00614127f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_302 VPB N_VPWR_c_2024_n 0.0552187f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_303 VPB N_VPWR_c_2025_n 0.00614151f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_304 VPB N_VPWR_c_2026_n 0.02253f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_305 VPB N_VPWR_c_2027_n 0.00614151f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_306 VPB N_VPWR_c_2028_n 0.0581188f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_307 VPB N_VPWR_c_2029_n 0.0301986f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_308 VPB N_VPWR_c_2030_n 0.0630629f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_309 VPB N_VPWR_c_2031_n 0.0335565f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_310 VPB N_VPWR_c_2032_n 0.0047828f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_311 VPB N_VPWR_c_2033_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_312 VPB N_VPWR_c_2034_n 0.00872592f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_313 VPB N_VPWR_c_2007_n 0.201629f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_314 VPB N_A_669_111#_c_2178_n 0.0021597f $X=-0.19 $Y=1.66 $X2=0.615 $Y2=1.275
cc_315 VPB N_A_669_111#_c_2179_n 0.00773134f $X=-0.19 $Y=1.66 $X2=0.615
+ $Y2=1.665
cc_316 VPB N_A_669_111#_c_2180_n 0.00104828f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_317 VPB N_A_669_111#_c_2172_n 0.0146872f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_318 VPB N_A_669_111#_c_2182_n 0.0211884f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_319 VPB N_A_669_111#_c_2183_n 0.0013145f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_320 VPB N_A_669_111#_c_2184_n 0.00168782f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_321 VPB N_A_669_111#_c_2185_n 0.0113166f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_322 VPB N_A_669_111#_c_2177_n 0.00997524f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_323 VPB N_A_669_111#_c_2187_n 0.00851243f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_324 VPB N_A_669_111#_c_2188_n 0.00520801f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_325 VPB N_A_669_111#_c_2189_n 0.0104462f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_326 VPB Q 0.0143136f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=2.64
cc_327 N_D_c_335_n N_A_159_404#_c_381_n 0.0437624f $X=0.495 $Y=2.245 $X2=0 $Y2=0
cc_328 N_D_c_334_n N_A_159_404#_c_382_n 0.0148107f $X=0.495 $Y=2.155 $X2=0 $Y2=0
cc_329 N_D_c_333_n N_A_159_404#_c_382_n 2.17226e-19 $X=0.58 $Y=1.275 $X2=0 $Y2=0
cc_330 N_D_c_329_n N_A_159_404#_c_374_n 3.80673e-19 $X=0.575 $Y=1.61 $X2=0 $Y2=0
cc_331 N_D_c_334_n N_A_159_404#_c_374_n 9.9879e-19 $X=0.495 $Y=2.155 $X2=0 $Y2=0
cc_332 N_D_c_332_n N_A_159_404#_c_374_n 0.0015654f $X=0.58 $Y=1.275 $X2=0 $Y2=0
cc_333 N_D_c_333_n N_A_159_404#_c_374_n 0.0513741f $X=0.58 $Y=1.275 $X2=0 $Y2=0
cc_334 N_D_c_329_n N_A_159_404#_c_375_n 0.0188968f $X=0.575 $Y=1.61 $X2=0 $Y2=0
cc_335 N_D_c_334_n N_A_159_404#_c_375_n 0.00771914f $X=0.495 $Y=2.155 $X2=0
+ $Y2=0
cc_336 N_D_c_333_n N_A_159_404#_c_375_n 0.00203546f $X=0.58 $Y=1.275 $X2=0 $Y2=0
cc_337 N_D_M1017_g N_A_159_404#_c_377_n 7.90161e-19 $X=0.64 $Y=0.58 $X2=0 $Y2=0
cc_338 N_D_c_333_n N_A_159_404#_c_377_n 0.00339256f $X=0.58 $Y=1.275 $X2=0 $Y2=0
cc_339 N_D_c_334_n N_A_159_404#_c_385_n 8.60369e-19 $X=0.495 $Y=2.155 $X2=0
+ $Y2=0
cc_340 N_D_M1017_g N_DE_M1004_g 0.0460069f $X=0.64 $Y=0.58 $X2=0 $Y2=0
cc_341 N_D_c_332_n N_DE_c_491_n 0.00594772f $X=0.58 $Y=1.275 $X2=0 $Y2=0
cc_342 N_D_c_333_n N_DE_c_491_n 5.91251e-19 $X=0.58 $Y=1.275 $X2=0 $Y2=0
cc_343 N_D_c_335_n N_A_27_74#_c_1884_n 0.00151458f $X=0.495 $Y=2.245 $X2=0 $Y2=0
cc_344 N_D_M1017_g N_A_27_74#_c_1884_n 0.00883069f $X=0.64 $Y=0.58 $X2=0 $Y2=0
cc_345 N_D_c_332_n N_A_27_74#_c_1884_n 0.0320048f $X=0.58 $Y=1.275 $X2=0 $Y2=0
cc_346 N_D_c_333_n N_A_27_74#_c_1884_n 0.0508256f $X=0.58 $Y=1.275 $X2=0 $Y2=0
cc_347 N_D_c_335_n N_A_27_74#_c_1890_n 0.00909651f $X=0.495 $Y=2.245 $X2=0 $Y2=0
cc_348 N_D_c_335_n N_A_27_74#_c_1891_n 0.013421f $X=0.495 $Y=2.245 $X2=0 $Y2=0
cc_349 N_D_c_331_n N_A_27_74#_c_1891_n 8.5751e-19 $X=0.575 $Y=1.78 $X2=0 $Y2=0
cc_350 N_D_c_333_n N_A_27_74#_c_1891_n 0.0125489f $X=0.58 $Y=1.275 $X2=0 $Y2=0
cc_351 N_D_M1017_g N_A_27_74#_c_1887_n 0.013685f $X=0.64 $Y=0.58 $X2=0 $Y2=0
cc_352 N_D_c_332_n N_A_27_74#_c_1887_n 0.00173628f $X=0.58 $Y=1.275 $X2=0 $Y2=0
cc_353 N_D_c_333_n N_A_27_74#_c_1887_n 0.00887419f $X=0.58 $Y=1.275 $X2=0 $Y2=0
cc_354 N_D_c_335_n N_A_27_74#_c_1899_n 0.00217861f $X=0.495 $Y=2.245 $X2=0 $Y2=0
cc_355 N_D_c_333_n N_A_27_74#_c_1899_n 3.08769e-19 $X=0.58 $Y=1.275 $X2=0 $Y2=0
cc_356 N_D_c_335_n N_VPWR_c_2008_n 0.0015335f $X=0.495 $Y=2.245 $X2=0 $Y2=0
cc_357 N_D_c_335_n N_VPWR_c_2018_n 0.00445602f $X=0.495 $Y=2.245 $X2=0 $Y2=0
cc_358 N_D_c_335_n N_VPWR_c_2007_n 0.00861324f $X=0.495 $Y=2.245 $X2=0 $Y2=0
cc_359 N_D_M1017_g N_VGND_c_2387_n 0.00214336f $X=0.64 $Y=0.58 $X2=0 $Y2=0
cc_360 N_D_M1017_g N_VGND_c_2402_n 0.00435951f $X=0.64 $Y=0.58 $X2=0 $Y2=0
cc_361 N_D_M1017_g N_VGND_c_2413_n 0.0082474f $X=0.64 $Y=0.58 $X2=0 $Y2=0
cc_362 N_A_159_404#_c_377_n N_DE_M1004_g 0.00936862f $X=1.305 $Y=1.065 $X2=0
+ $Y2=0
cc_363 N_A_159_404#_c_378_n N_DE_M1004_g 0.00467324f $X=1.805 $Y=0.765 $X2=0
+ $Y2=0
cc_364 N_A_159_404#_c_374_n N_DE_c_490_n 0.00529154f $X=1.14 $Y=1.605 $X2=0
+ $Y2=0
cc_365 N_A_159_404#_c_376_n N_DE_c_490_n 0.0128862f $X=1.64 $Y=1.065 $X2=0 $Y2=0
cc_366 N_A_159_404#_c_377_n N_DE_c_490_n 0.0035816f $X=1.305 $Y=1.065 $X2=0
+ $Y2=0
cc_367 N_A_159_404#_c_374_n N_DE_c_491_n 0.00217967f $X=1.14 $Y=1.605 $X2=0
+ $Y2=0
cc_368 N_A_159_404#_c_375_n N_DE_c_491_n 0.0182467f $X=1.14 $Y=1.605 $X2=0 $Y2=0
cc_369 N_A_159_404#_c_377_n N_DE_c_491_n 0.00230966f $X=1.305 $Y=1.065 $X2=0
+ $Y2=0
cc_370 N_A_159_404#_c_374_n N_DE_c_492_n 0.00113501f $X=1.14 $Y=1.605 $X2=0
+ $Y2=0
cc_371 N_A_159_404#_c_375_n N_DE_c_492_n 0.0076847f $X=1.14 $Y=1.605 $X2=0 $Y2=0
cc_372 N_A_159_404#_c_384_n N_DE_c_492_n 0.00300051f $X=1.705 $Y=2.035 $X2=0
+ $Y2=0
cc_373 N_A_159_404#_c_379_n N_DE_c_492_n 0.00403373f $X=2.22 $Y=1.685 $X2=0
+ $Y2=0
cc_374 N_A_159_404#_c_389_n N_DE_c_492_n 0.0062364f $X=1.79 $Y=2.035 $X2=0 $Y2=0
cc_375 N_A_159_404#_c_380_n N_DE_c_492_n 0.0110636f $X=2.45 $Y=1.685 $X2=0 $Y2=0
cc_376 N_A_159_404#_c_386_n N_DE_c_498_n 0.00415054f $X=1.79 $Y=2.515 $X2=0
+ $Y2=0
cc_377 N_A_159_404#_M1012_g N_DE_c_493_n 0.0189277f $X=2.45 $Y=0.765 $X2=0 $Y2=0
cc_378 N_A_159_404#_c_376_n N_DE_c_493_n 0.00267945f $X=1.64 $Y=1.065 $X2=0
+ $Y2=0
cc_379 N_A_159_404#_c_378_n N_DE_c_493_n 0.00112392f $X=1.805 $Y=0.765 $X2=0
+ $Y2=0
cc_380 N_A_159_404#_c_387_n N_DE_c_499_n 0.00748816f $X=2.055 $Y=2.035 $X2=0
+ $Y2=0
cc_381 N_A_159_404#_c_382_n N_DE_c_500_n 0.0110122f $X=0.885 $Y=2.132 $X2=0
+ $Y2=0
cc_382 N_A_159_404#_c_384_n N_DE_c_500_n 0.00205074f $X=1.705 $Y=2.035 $X2=0
+ $Y2=0
cc_383 N_A_159_404#_c_386_n N_DE_c_500_n 0.0143357f $X=1.79 $Y=2.515 $X2=0 $Y2=0
cc_384 N_A_159_404#_c_387_n N_DE_c_500_n 0.0116886f $X=2.055 $Y=2.035 $X2=0
+ $Y2=0
cc_385 N_A_159_404#_c_389_n N_DE_c_500_n 0.00129501f $X=1.79 $Y=2.035 $X2=0
+ $Y2=0
cc_386 N_A_159_404#_c_380_n N_DE_c_500_n 0.0265887f $X=2.45 $Y=1.685 $X2=0 $Y2=0
cc_387 N_A_159_404#_c_376_n N_DE_c_494_n 0.0163184f $X=1.64 $Y=1.065 $X2=0 $Y2=0
cc_388 N_A_159_404#_c_379_n N_DE_c_494_n 2.29827e-19 $X=2.22 $Y=1.685 $X2=0
+ $Y2=0
cc_389 N_A_159_404#_c_380_n N_DE_c_494_n 0.00159577f $X=2.45 $Y=1.685 $X2=0
+ $Y2=0
cc_390 N_A_159_404#_M1012_g N_DE_c_495_n 0.00853426f $X=2.45 $Y=0.765 $X2=0
+ $Y2=0
cc_391 N_A_159_404#_c_374_n N_DE_c_495_n 0.00802476f $X=1.14 $Y=1.605 $X2=0
+ $Y2=0
cc_392 N_A_159_404#_c_375_n N_DE_c_495_n 0.0127671f $X=1.14 $Y=1.605 $X2=0 $Y2=0
cc_393 N_A_159_404#_M1012_g N_DE_c_502_n 0.00104309f $X=2.45 $Y=0.765 $X2=0
+ $Y2=0
cc_394 N_A_159_404#_c_374_n N_DE_c_502_n 0.0301697f $X=1.14 $Y=1.605 $X2=0 $Y2=0
cc_395 N_A_159_404#_c_375_n N_DE_c_502_n 0.00170436f $X=1.14 $Y=1.605 $X2=0
+ $Y2=0
cc_396 N_A_159_404#_c_376_n N_DE_c_502_n 0.024732f $X=1.64 $Y=1.065 $X2=0 $Y2=0
cc_397 N_A_159_404#_c_384_n N_DE_c_502_n 0.0151027f $X=1.705 $Y=2.035 $X2=0
+ $Y2=0
cc_398 N_A_159_404#_c_379_n N_DE_c_502_n 0.0170229f $X=2.22 $Y=1.685 $X2=0 $Y2=0
cc_399 N_A_159_404#_c_389_n N_DE_c_502_n 0.0116821f $X=1.79 $Y=2.035 $X2=0 $Y2=0
cc_400 N_A_159_404#_c_380_n N_DE_c_502_n 0.00131025f $X=2.45 $Y=1.685 $X2=0
+ $Y2=0
cc_401 N_A_159_404#_c_384_n N_DE_c_496_n 7.50963e-19 $X=1.705 $Y=2.035 $X2=0
+ $Y2=0
cc_402 N_A_159_404#_c_379_n N_DE_c_496_n 4.52778e-19 $X=2.22 $Y=1.685 $X2=0
+ $Y2=0
cc_403 N_A_159_404#_c_380_n N_DE_c_496_n 0.00813987f $X=2.45 $Y=1.685 $X2=0
+ $Y2=0
cc_404 N_A_159_404#_M1012_g N_A_547_301#_M1038_g 0.0562452f $X=2.45 $Y=0.765
+ $X2=0 $Y2=0
cc_405 N_A_159_404#_c_387_n N_A_547_301#_c_592_n 0.0038026f $X=2.055 $Y=2.035
+ $X2=0 $Y2=0
cc_406 N_A_159_404#_c_379_n N_A_547_301#_c_592_n 0.00244729f $X=2.22 $Y=1.685
+ $X2=0 $Y2=0
cc_407 N_A_159_404#_c_380_n N_A_547_301#_c_592_n 4.41976e-19 $X=2.45 $Y=1.685
+ $X2=0 $Y2=0
cc_408 N_A_159_404#_c_379_n N_A_547_301#_c_586_n 0.00678737f $X=2.22 $Y=1.685
+ $X2=0 $Y2=0
cc_409 N_A_159_404#_c_380_n N_A_547_301#_c_586_n 0.00472168f $X=2.45 $Y=1.685
+ $X2=0 $Y2=0
cc_410 N_A_159_404#_M1012_g N_A_547_301#_c_589_n 0.00255748f $X=2.45 $Y=0.765
+ $X2=0 $Y2=0
cc_411 N_A_159_404#_c_379_n N_A_547_301#_c_589_n 0.0222225f $X=2.22 $Y=1.685
+ $X2=0 $Y2=0
cc_412 N_A_159_404#_M1012_g N_A_547_301#_c_590_n 0.0219933f $X=2.45 $Y=0.765
+ $X2=0 $Y2=0
cc_413 N_A_159_404#_c_379_n N_A_547_301#_c_590_n 2.27104e-19 $X=2.22 $Y=1.685
+ $X2=0 $Y2=0
cc_414 N_A_159_404#_c_381_n N_A_27_74#_c_1890_n 0.00180228f $X=0.885 $Y=2.245
+ $X2=0 $Y2=0
cc_415 N_A_159_404#_c_381_n N_A_27_74#_c_1891_n 0.0199182f $X=0.885 $Y=2.245
+ $X2=0 $Y2=0
cc_416 N_A_159_404#_c_382_n N_A_27_74#_c_1891_n 0.00652688f $X=0.885 $Y=2.132
+ $X2=0 $Y2=0
cc_417 N_A_159_404#_c_384_n N_A_27_74#_c_1891_n 0.018801f $X=1.705 $Y=2.035
+ $X2=0 $Y2=0
cc_418 N_A_159_404#_c_385_n N_A_27_74#_c_1891_n 0.0271868f $X=1.305 $Y=2.035
+ $X2=0 $Y2=0
cc_419 N_A_159_404#_c_386_n N_A_27_74#_c_1891_n 0.0141649f $X=1.79 $Y=2.515
+ $X2=0 $Y2=0
cc_420 N_A_159_404#_c_381_n N_A_27_74#_c_1892_n 0.00426176f $X=0.885 $Y=2.245
+ $X2=0 $Y2=0
cc_421 N_A_159_404#_c_386_n N_A_27_74#_c_1892_n 0.0203028f $X=1.79 $Y=2.515
+ $X2=0 $Y2=0
cc_422 N_A_159_404#_M1036_s N_A_27_74#_c_1893_n 0.00361559f $X=1.645 $Y=2.315
+ $X2=0 $Y2=0
cc_423 N_A_159_404#_c_386_n N_A_27_74#_c_1893_n 0.012787f $X=1.79 $Y=2.515 $X2=0
+ $Y2=0
cc_424 N_A_159_404#_c_381_n N_A_27_74#_c_1894_n 6.5162e-19 $X=0.885 $Y=2.245
+ $X2=0 $Y2=0
cc_425 N_A_159_404#_c_386_n N_A_27_74#_c_1925_n 0.0192722f $X=1.79 $Y=2.515
+ $X2=0 $Y2=0
cc_426 N_A_159_404#_c_387_n N_A_27_74#_c_1895_n 0.0134118f $X=2.055 $Y=2.035
+ $X2=0 $Y2=0
cc_427 N_A_159_404#_c_386_n N_A_27_74#_c_1896_n 0.0133944f $X=1.79 $Y=2.515
+ $X2=0 $Y2=0
cc_428 N_A_159_404#_c_387_n N_A_27_74#_c_1896_n 0.0146675f $X=2.055 $Y=2.035
+ $X2=0 $Y2=0
cc_429 N_A_159_404#_c_380_n N_A_27_74#_c_1896_n 2.29212e-19 $X=2.45 $Y=1.685
+ $X2=0 $Y2=0
cc_430 N_A_159_404#_M1012_g N_A_27_74#_c_1885_n 0.00214472f $X=2.45 $Y=0.765
+ $X2=0 $Y2=0
cc_431 N_A_159_404#_M1012_g N_A_27_74#_c_1888_n 8.29074e-19 $X=2.45 $Y=0.765
+ $X2=0 $Y2=0
cc_432 N_A_159_404#_c_381_n N_VPWR_c_2008_n 0.0104537f $X=0.885 $Y=2.245 $X2=0
+ $Y2=0
cc_433 N_A_159_404#_c_381_n N_VPWR_c_2018_n 0.00413917f $X=0.885 $Y=2.245 $X2=0
+ $Y2=0
cc_434 N_A_159_404#_c_381_n N_VPWR_c_2007_n 0.00817239f $X=0.885 $Y=2.245 $X2=0
+ $Y2=0
cc_435 N_A_159_404#_c_376_n N_VGND_c_2387_n 0.00874483f $X=1.64 $Y=1.065 $X2=0
+ $Y2=0
cc_436 N_A_159_404#_c_377_n N_VGND_c_2387_n 0.0207698f $X=1.305 $Y=1.065 $X2=0
+ $Y2=0
cc_437 N_A_159_404#_c_378_n N_VGND_c_2387_n 0.0181585f $X=1.805 $Y=0.765 $X2=0
+ $Y2=0
cc_438 N_A_159_404#_M1012_g N_VGND_c_2388_n 0.0132084f $X=2.45 $Y=0.765 $X2=0
+ $Y2=0
cc_439 N_A_159_404#_c_376_n N_VGND_c_2388_n 0.00121149f $X=1.64 $Y=1.065 $X2=0
+ $Y2=0
cc_440 N_A_159_404#_c_378_n N_VGND_c_2388_n 0.0167923f $X=1.805 $Y=0.765 $X2=0
+ $Y2=0
cc_441 N_A_159_404#_c_379_n N_VGND_c_2388_n 0.0116552f $X=2.22 $Y=1.685 $X2=0
+ $Y2=0
cc_442 N_A_159_404#_c_380_n N_VGND_c_2388_n 0.0018691f $X=2.45 $Y=1.685 $X2=0
+ $Y2=0
cc_443 N_A_159_404#_M1012_g N_VGND_c_2396_n 0.00377474f $X=2.45 $Y=0.765 $X2=0
+ $Y2=0
cc_444 N_A_159_404#_c_378_n N_VGND_c_2403_n 0.00619316f $X=1.805 $Y=0.765 $X2=0
+ $Y2=0
cc_445 N_A_159_404#_M1012_g N_VGND_c_2413_n 0.00410937f $X=2.45 $Y=0.765 $X2=0
+ $Y2=0
cc_446 N_A_159_404#_c_378_n N_VGND_c_2413_n 0.00802722f $X=1.805 $Y=0.765 $X2=0
+ $Y2=0
cc_447 N_DE_c_499_n N_A_547_301#_c_592_n 0.010561f $X=2.62 $Y=2.165 $X2=0 $Y2=0
cc_448 N_DE_c_501_n N_A_547_301#_c_593_n 0.0437219f $X=2.695 $Y=2.24 $X2=0 $Y2=0
cc_449 N_DE_c_499_n N_A_547_301#_c_586_n 9.30616e-19 $X=2.62 $Y=2.165 $X2=0
+ $Y2=0
cc_450 N_DE_c_499_n N_A_547_301#_c_589_n 0.00510927f $X=2.62 $Y=2.165 $X2=0
+ $Y2=0
cc_451 N_DE_c_499_n N_A_547_301#_c_590_n 0.0026439f $X=2.62 $Y=2.165 $X2=0 $Y2=0
cc_452 N_DE_c_498_n N_A_27_74#_c_1892_n 0.00326422f $X=2.015 $Y=2.24 $X2=0 $Y2=0
cc_453 N_DE_c_498_n N_A_27_74#_c_1893_n 0.0134964f $X=2.015 $Y=2.24 $X2=0 $Y2=0
cc_454 N_DE_c_500_n N_A_27_74#_c_1893_n 0.00222708f $X=2.09 $Y=2.165 $X2=0 $Y2=0
cc_455 N_DE_c_501_n N_A_27_74#_c_1893_n 4.28313e-19 $X=2.695 $Y=2.24 $X2=0 $Y2=0
cc_456 N_DE_c_498_n N_A_27_74#_c_1925_n 0.0118088f $X=2.015 $Y=2.24 $X2=0 $Y2=0
cc_457 N_DE_c_501_n N_A_27_74#_c_1925_n 0.00283455f $X=2.695 $Y=2.24 $X2=0 $Y2=0
cc_458 N_DE_c_499_n N_A_27_74#_c_1895_n 0.00979321f $X=2.62 $Y=2.165 $X2=0 $Y2=0
cc_459 N_DE_c_501_n N_A_27_74#_c_1895_n 0.0156958f $X=2.695 $Y=2.24 $X2=0 $Y2=0
cc_460 N_DE_c_498_n N_A_27_74#_c_1896_n 0.0058392f $X=2.015 $Y=2.24 $X2=0 $Y2=0
cc_461 N_DE_c_499_n N_A_27_74#_c_1896_n 8.10671e-19 $X=2.62 $Y=2.165 $X2=0 $Y2=0
cc_462 N_DE_c_501_n N_A_27_74#_c_1897_n 0.00179485f $X=2.695 $Y=2.24 $X2=0 $Y2=0
cc_463 N_DE_M1004_g N_A_27_74#_c_1887_n 9.27003e-19 $X=1.03 $Y=0.58 $X2=0 $Y2=0
cc_464 N_DE_c_498_n N_VPWR_c_2009_n 0.00153478f $X=2.015 $Y=2.24 $X2=0 $Y2=0
cc_465 N_DE_c_501_n N_VPWR_c_2009_n 0.00967911f $X=2.695 $Y=2.24 $X2=0 $Y2=0
cc_466 N_DE_c_498_n N_VPWR_c_2020_n 0.00275664f $X=2.015 $Y=2.24 $X2=0 $Y2=0
cc_467 N_DE_c_501_n N_VPWR_c_2028_n 0.00410286f $X=2.695 $Y=2.24 $X2=0 $Y2=0
cc_468 N_DE_c_498_n N_VPWR_c_2007_n 0.00544287f $X=2.015 $Y=2.24 $X2=0 $Y2=0
cc_469 N_DE_c_501_n N_VPWR_c_2007_n 0.00493487f $X=2.695 $Y=2.24 $X2=0 $Y2=0
cc_470 N_DE_M1004_g N_VGND_c_2387_n 0.0141988f $X=1.03 $Y=0.58 $X2=0 $Y2=0
cc_471 N_DE_c_490_n N_VGND_c_2387_n 0.00144101f $X=1.515 $Y=1.125 $X2=0 $Y2=0
cc_472 N_DE_c_493_n N_VGND_c_2387_n 0.00223024f $X=2.02 $Y=1.05 $X2=0 $Y2=0
cc_473 N_DE_c_493_n N_VGND_c_2388_n 0.0105305f $X=2.02 $Y=1.05 $X2=0 $Y2=0
cc_474 N_DE_M1004_g N_VGND_c_2402_n 0.00383152f $X=1.03 $Y=0.58 $X2=0 $Y2=0
cc_475 N_DE_c_493_n N_VGND_c_2403_n 0.00377474f $X=2.02 $Y=1.05 $X2=0 $Y2=0
cc_476 N_DE_M1004_g N_VGND_c_2413_n 0.0075725f $X=1.03 $Y=0.58 $X2=0 $Y2=0
cc_477 N_DE_c_493_n N_VGND_c_2413_n 0.00410937f $X=2.02 $Y=1.05 $X2=0 $Y2=0
cc_478 N_A_547_301#_M1038_g N_A_639_85#_c_817_n 0.0180128f $X=2.84 $Y=0.765
+ $X2=0 $Y2=0
cc_479 N_A_547_301#_c_585_n N_A_639_85#_c_818_n 0.00570953f $X=14.015 $Y=1.665
+ $X2=0 $Y2=0
cc_480 N_A_547_301#_c_585_n N_A_639_85#_c_823_n 0.0247491f $X=14.015 $Y=1.665
+ $X2=0 $Y2=0
cc_481 N_A_547_301#_c_585_n N_A_639_85#_c_824_n 0.00715008f $X=14.015 $Y=1.665
+ $X2=0 $Y2=0
cc_482 N_A_547_301#_c_590_n N_A_639_85#_c_824_n 0.00548413f $X=3.085 $Y=1.67
+ $X2=0 $Y2=0
cc_483 N_A_547_301#_c_585_n N_A_639_85#_c_833_n 0.0386859f $X=14.015 $Y=1.665
+ $X2=0 $Y2=0
cc_484 N_A_547_301#_c_585_n N_A_639_85#_c_825_n 0.0184731f $X=14.015 $Y=1.665
+ $X2=0 $Y2=0
cc_485 N_A_547_301#_c_585_n N_A_639_85#_c_826_n 0.00228959f $X=14.015 $Y=1.665
+ $X2=0 $Y2=0
cc_486 N_A_547_301#_c_585_n N_A_639_85#_c_827_n 0.008134f $X=14.015 $Y=1.665
+ $X2=0 $Y2=0
cc_487 N_A_547_301#_c_585_n N_A_639_85#_c_836_n 7.90379e-19 $X=14.015 $Y=1.665
+ $X2=0 $Y2=0
cc_488 N_A_547_301#_c_585_n SCD 0.0305151f $X=14.015 $Y=1.665 $X2=0 $Y2=0
cc_489 N_A_547_301#_c_585_n N_SCD_c_933_n 6.94548e-19 $X=14.015 $Y=1.665 $X2=0
+ $Y2=0
cc_490 N_A_547_301#_c_593_n N_SCE_c_984_n 0.0074134f $X=3.085 $Y=2.24 $X2=-0.19
+ $Y2=-0.245
cc_491 N_A_547_301#_c_585_n N_SCE_c_984_n 0.00250527f $X=14.015 $Y=1.665
+ $X2=-0.19 $Y2=-0.245
cc_492 N_A_547_301#_c_593_n N_SCE_c_986_n 0.00288121f $X=3.085 $Y=2.24 $X2=0
+ $Y2=0
cc_493 N_A_547_301#_c_585_n N_SCE_c_977_n 0.00600851f $X=14.015 $Y=1.665 $X2=0
+ $Y2=0
cc_494 N_A_547_301#_c_585_n N_SCE_M1028_g 0.0030065f $X=14.015 $Y=1.665 $X2=0
+ $Y2=0
cc_495 N_A_547_301#_c_585_n SCE 0.00971008f $X=14.015 $Y=1.665 $X2=0 $Y2=0
cc_496 N_A_547_301#_c_585_n N_CLK_c_1064_n 0.00780772f $X=14.015 $Y=1.665 $X2=0
+ $Y2=0
cc_497 N_A_547_301#_c_585_n CLK 0.0153239f $X=14.015 $Y=1.665 $X2=0 $Y2=0
cc_498 N_A_547_301#_c_594_n N_A_1492_74#_c_1098_n 0.0199822f $X=13.185 $Y=2.465
+ $X2=0 $Y2=0
cc_499 N_A_547_301#_c_583_n N_A_1492_74#_c_1098_n 0.0167078f $X=13.29 $Y=2.05
+ $X2=0 $Y2=0
cc_500 N_A_547_301#_c_596_n N_A_1492_74#_c_1098_n 9.79303e-19 $X=13.955 $Y=2.227
+ $X2=0 $Y2=0
cc_501 N_A_547_301#_c_585_n N_A_1492_74#_c_1098_n 0.00460492f $X=14.015 $Y=1.665
+ $X2=0 $Y2=0
cc_502 N_A_547_301#_c_594_n N_A_1492_74#_c_1122_n 0.0324071f $X=13.185 $Y=2.465
+ $X2=0 $Y2=0
cc_503 N_A_547_301#_c_585_n N_A_1492_74#_c_1099_n 0.00510576f $X=14.015 $Y=1.665
+ $X2=0 $Y2=0
cc_504 N_A_547_301#_c_585_n N_A_1492_74#_c_1123_n 0.0187939f $X=14.015 $Y=1.665
+ $X2=0 $Y2=0
cc_505 N_A_547_301#_c_585_n N_A_1492_74#_c_1102_n 0.0196832f $X=14.015 $Y=1.665
+ $X2=0 $Y2=0
cc_506 N_A_547_301#_c_585_n N_A_1492_74#_c_1105_n 0.00629785f $X=14.015 $Y=1.665
+ $X2=0 $Y2=0
cc_507 N_A_547_301#_c_585_n N_A_1492_74#_c_1106_n 0.00151815f $X=14.015 $Y=1.665
+ $X2=0 $Y2=0
cc_508 N_A_547_301#_c_585_n N_A_1492_74#_c_1107_n 0.00522051f $X=14.015 $Y=1.665
+ $X2=0 $Y2=0
cc_509 N_A_547_301#_c_585_n N_A_1492_74#_c_1111_n 0.0054723f $X=14.015 $Y=1.665
+ $X2=0 $Y2=0
cc_510 N_A_547_301#_c_585_n N_A_1492_74#_c_1114_n 0.0387589f $X=14.015 $Y=1.665
+ $X2=0 $Y2=0
cc_511 N_A_547_301#_c_585_n N_A_1492_74#_c_1115_n 0.00372651f $X=14.015 $Y=1.665
+ $X2=0 $Y2=0
cc_512 N_A_547_301#_c_585_n N_A_1492_74#_c_1116_n 0.0140456f $X=14.015 $Y=1.665
+ $X2=0 $Y2=0
cc_513 N_A_547_301#_c_585_n N_A_1492_74#_c_1127_n 4.33735e-19 $X=14.015 $Y=1.665
+ $X2=0 $Y2=0
cc_514 N_A_547_301#_c_582_n N_A_1492_74#_c_1118_n 0.00221599f $X=12.825 $Y=0.94
+ $X2=0 $Y2=0
cc_515 N_A_547_301#_c_583_n N_A_1492_74#_c_1118_n 0.00115933f $X=13.29 $Y=2.05
+ $X2=0 $Y2=0
cc_516 N_A_547_301#_c_585_n N_A_1492_74#_c_1118_n 0.00907344f $X=14.015 $Y=1.665
+ $X2=0 $Y2=0
cc_517 N_A_547_301#_c_582_n N_A_1492_74#_c_1119_n 0.0204399f $X=12.825 $Y=0.94
+ $X2=0 $Y2=0
cc_518 N_A_547_301#_c_583_n N_A_1492_74#_c_1119_n 0.020543f $X=13.29 $Y=2.05
+ $X2=0 $Y2=0
cc_519 N_A_547_301#_c_585_n N_A_1295_74#_M1007_g 0.00681622f $X=14.015 $Y=1.665
+ $X2=0 $Y2=0
cc_520 N_A_547_301#_c_585_n N_A_1295_74#_c_1330_n 0.00343737f $X=14.015 $Y=1.665
+ $X2=0 $Y2=0
cc_521 N_A_547_301#_c_585_n N_A_1295_74#_c_1331_n 0.00234493f $X=14.015 $Y=1.665
+ $X2=0 $Y2=0
cc_522 N_A_547_301#_c_585_n N_A_1295_74#_M1026_g 0.00507242f $X=14.015 $Y=1.665
+ $X2=0 $Y2=0
cc_523 N_A_547_301#_c_585_n N_A_1295_74#_c_1333_n 0.00396108f $X=14.015 $Y=1.665
+ $X2=0 $Y2=0
cc_524 N_A_547_301#_c_585_n N_A_1295_74#_c_1334_n 0.00810975f $X=14.015 $Y=1.665
+ $X2=0 $Y2=0
cc_525 N_A_547_301#_c_580_n N_A_1295_74#_M1034_g 0.0416832f $X=12.75 $Y=0.865
+ $X2=0 $Y2=0
cc_526 N_A_547_301#_c_585_n N_A_1295_74#_c_1336_n 0.00855361f $X=14.015 $Y=1.665
+ $X2=0 $Y2=0
cc_527 N_A_547_301#_c_585_n N_A_1295_74#_c_1337_n 0.00210802f $X=14.015 $Y=1.665
+ $X2=0 $Y2=0
cc_528 N_A_547_301#_c_585_n N_A_1295_74#_c_1338_n 8.23884e-19 $X=14.015 $Y=1.665
+ $X2=0 $Y2=0
cc_529 N_A_547_301#_c_585_n N_A_1295_74#_c_1340_n 0.0149279f $X=14.015 $Y=1.665
+ $X2=0 $Y2=0
cc_530 N_A_547_301#_c_585_n N_A_1295_74#_c_1354_n 0.0179094f $X=14.015 $Y=1.665
+ $X2=0 $Y2=0
cc_531 N_A_547_301#_c_585_n N_A_1295_74#_c_1356_n 0.00326617f $X=14.015 $Y=1.665
+ $X2=0 $Y2=0
cc_532 N_A_547_301#_c_585_n N_A_1295_74#_c_1360_n 0.00447604f $X=14.015 $Y=1.665
+ $X2=0 $Y2=0
cc_533 N_A_547_301#_c_585_n N_A_1295_74#_c_1341_n 0.00590512f $X=14.015 $Y=1.665
+ $X2=0 $Y2=0
cc_534 N_A_547_301#_c_585_n N_A_1295_74#_c_1361_n 0.0140274f $X=14.015 $Y=1.665
+ $X2=0 $Y2=0
cc_535 N_A_547_301#_c_585_n N_A_1295_74#_c_1342_n 0.0202419f $X=14.015 $Y=1.665
+ $X2=0 $Y2=0
cc_536 N_A_547_301#_c_585_n N_A_1910_71#_c_1530_n 0.00192843f $X=14.015 $Y=1.665
+ $X2=0 $Y2=0
cc_537 N_A_547_301#_c_585_n N_A_1910_71#_c_1531_n 0.0126659f $X=14.015 $Y=1.665
+ $X2=0 $Y2=0
cc_538 N_A_547_301#_c_585_n N_A_1910_71#_c_1533_n 0.00936086f $X=14.015 $Y=1.665
+ $X2=0 $Y2=0
cc_539 N_A_547_301#_c_585_n N_A_1910_71#_c_1535_n 0.0169862f $X=14.015 $Y=1.665
+ $X2=0 $Y2=0
cc_540 N_A_547_301#_c_585_n N_A_1910_71#_c_1536_n 0.00392515f $X=14.015 $Y=1.665
+ $X2=0 $Y2=0
cc_541 N_A_547_301#_c_585_n N_A_1910_71#_c_1537_n 0.0282283f $X=14.015 $Y=1.665
+ $X2=0 $Y2=0
cc_542 N_A_547_301#_c_585_n N_A_1910_71#_c_1538_n 0.010664f $X=14.015 $Y=1.665
+ $X2=0 $Y2=0
cc_543 N_A_547_301#_c_585_n N_A_1910_71#_c_1539_n 0.0078177f $X=14.015 $Y=1.665
+ $X2=0 $Y2=0
cc_544 N_A_547_301#_c_585_n N_A_1910_71#_c_1547_n 0.00624077f $X=14.015 $Y=1.665
+ $X2=0 $Y2=0
cc_545 N_A_547_301#_c_585_n N_A_1910_71#_c_1540_n 0.00470461f $X=14.015 $Y=1.665
+ $X2=0 $Y2=0
cc_546 N_A_547_301#_c_585_n N_A_1910_71#_c_1541_n 0.00425165f $X=14.015 $Y=1.665
+ $X2=0 $Y2=0
cc_547 N_A_547_301#_c_585_n N_A_1688_97#_c_1642_n 0.00243608f $X=14.015 $Y=1.665
+ $X2=0 $Y2=0
cc_548 N_A_547_301#_c_585_n N_A_1688_97#_c_1644_n 0.0103123f $X=14.015 $Y=1.665
+ $X2=0 $Y2=0
cc_549 N_A_547_301#_c_585_n N_A_1688_97#_c_1649_n 0.013499f $X=14.015 $Y=1.665
+ $X2=0 $Y2=0
cc_550 N_A_547_301#_c_585_n N_A_1688_97#_c_1645_n 0.0226429f $X=14.015 $Y=1.665
+ $X2=0 $Y2=0
cc_551 N_A_547_301#_c_585_n N_A_1688_97#_c_1646_n 0.0543747f $X=14.015 $Y=1.665
+ $X2=0 $Y2=0
cc_552 N_A_547_301#_c_581_n N_A_2385_74#_M1019_g 0.00587027f $X=13.215 $Y=0.94
+ $X2=0 $Y2=0
cc_553 N_A_547_301#_c_584_n N_A_2385_74#_M1019_g 0.0132432f $X=14.09 $Y=0.58
+ $X2=0 $Y2=0
cc_554 N_A_547_301#_c_591_n N_A_2385_74#_M1019_g 0.00822691f $X=14.165 $Y=1.55
+ $X2=0 $Y2=0
cc_555 N_A_547_301#_c_594_n N_A_2385_74#_c_1741_n 0.00539777f $X=13.185 $Y=2.465
+ $X2=0 $Y2=0
cc_556 N_A_547_301#_c_596_n N_A_2385_74#_c_1741_n 0.00529843f $X=13.955 $Y=2.227
+ $X2=0 $Y2=0
cc_557 N_A_547_301#_c_599_n N_A_2385_74#_c_1741_n 0.00247226f $X=14.12 $Y=2.227
+ $X2=0 $Y2=0
cc_558 N_A_547_301#_c_585_n N_A_2385_74#_c_1741_n 0.00471849f $X=14.015 $Y=1.665
+ $X2=0 $Y2=0
cc_559 N_A_547_301#_c_587_n N_A_2385_74#_c_1741_n 0.0011953f $X=14.16 $Y=1.665
+ $X2=0 $Y2=0
cc_560 N_A_547_301#_c_588_n N_A_2385_74#_c_1741_n 0.013343f $X=14.16 $Y=1.665
+ $X2=0 $Y2=0
cc_561 N_A_547_301#_c_594_n N_A_2385_74#_c_1752_n 0.0148188f $X=13.185 $Y=2.465
+ $X2=0 $Y2=0
cc_562 N_A_547_301#_c_596_n N_A_2385_74#_c_1752_n 0.0130594f $X=13.955 $Y=2.227
+ $X2=0 $Y2=0
cc_563 N_A_547_301#_c_597_n N_A_2385_74#_c_1752_n 0.00957711f $X=14.12 $Y=2.465
+ $X2=0 $Y2=0
cc_564 N_A_547_301#_c_599_n N_A_2385_74#_c_1752_n 0.00411219f $X=14.12 $Y=2.227
+ $X2=0 $Y2=0
cc_565 N_A_547_301#_c_599_n N_A_2385_74#_c_1742_n 0.00162285f $X=14.12 $Y=2.227
+ $X2=0 $Y2=0
cc_566 N_A_547_301#_c_585_n N_A_2385_74#_c_1742_n 0.00131041f $X=14.015 $Y=1.665
+ $X2=0 $Y2=0
cc_567 N_A_547_301#_c_587_n N_A_2385_74#_c_1742_n 0.00624135f $X=14.16 $Y=1.665
+ $X2=0 $Y2=0
cc_568 N_A_547_301#_c_588_n N_A_2385_74#_c_1742_n 0.0102169f $X=14.16 $Y=1.665
+ $X2=0 $Y2=0
cc_569 N_A_547_301#_c_591_n N_A_2385_74#_c_1742_n 0.0186482f $X=14.165 $Y=1.55
+ $X2=0 $Y2=0
cc_570 N_A_547_301#_c_583_n N_A_2385_74#_c_1743_n 0.0324311f $X=13.29 $Y=2.05
+ $X2=0 $Y2=0
cc_571 N_A_547_301#_c_596_n N_A_2385_74#_c_1743_n 7.11771e-19 $X=13.955 $Y=2.227
+ $X2=0 $Y2=0
cc_572 N_A_547_301#_c_584_n N_A_2385_74#_c_1743_n 0.00553752f $X=14.09 $Y=0.58
+ $X2=0 $Y2=0
cc_573 N_A_547_301#_c_585_n N_A_2385_74#_c_1743_n 0.0031725f $X=14.015 $Y=1.665
+ $X2=0 $Y2=0
cc_574 N_A_547_301#_c_591_n N_A_2385_74#_c_1743_n 0.0041084f $X=14.165 $Y=1.55
+ $X2=0 $Y2=0
cc_575 N_A_547_301#_c_584_n N_A_2385_74#_c_1744_n 0.00172591f $X=14.09 $Y=0.58
+ $X2=0 $Y2=0
cc_576 N_A_547_301#_c_597_n N_A_2385_74#_c_1753_n 0.00101948f $X=14.12 $Y=2.465
+ $X2=0 $Y2=0
cc_577 N_A_547_301#_c_598_n N_A_2385_74#_c_1753_n 6.01012e-19 $X=14.165 $Y=2.075
+ $X2=0 $Y2=0
cc_578 N_A_547_301#_c_599_n N_A_2385_74#_c_1753_n 6.1382e-19 $X=14.12 $Y=2.227
+ $X2=0 $Y2=0
cc_579 N_A_547_301#_c_588_n N_A_2385_74#_c_1745_n 4.68247e-19 $X=14.16 $Y=1.665
+ $X2=0 $Y2=0
cc_580 N_A_547_301#_c_580_n N_A_2385_74#_c_1747_n 0.00739677f $X=12.75 $Y=0.865
+ $X2=0 $Y2=0
cc_581 N_A_547_301#_c_581_n N_A_2385_74#_c_1747_n 0.0207909f $X=13.215 $Y=0.94
+ $X2=0 $Y2=0
cc_582 N_A_547_301#_c_582_n N_A_2385_74#_c_1747_n 0.00277863f $X=12.825 $Y=0.94
+ $X2=0 $Y2=0
cc_583 N_A_547_301#_c_584_n N_A_2385_74#_c_1747_n 0.00130753f $X=14.09 $Y=0.58
+ $X2=0 $Y2=0
cc_584 N_A_547_301#_c_594_n N_A_2385_74#_c_1755_n 2.58731e-19 $X=13.185 $Y=2.465
+ $X2=0 $Y2=0
cc_585 N_A_547_301#_c_583_n N_A_2385_74#_c_1755_n 7.7774e-19 $X=13.29 $Y=2.05
+ $X2=0 $Y2=0
cc_586 N_A_547_301#_c_596_n N_A_2385_74#_c_1755_n 0.00470681f $X=13.955 $Y=2.227
+ $X2=0 $Y2=0
cc_587 N_A_547_301#_c_585_n N_A_2385_74#_c_1755_n 0.0134505f $X=14.015 $Y=1.665
+ $X2=0 $Y2=0
cc_588 N_A_547_301#_c_594_n N_A_2385_74#_c_1756_n 0.00299156f $X=13.185 $Y=2.465
+ $X2=0 $Y2=0
cc_589 N_A_547_301#_c_596_n N_A_2385_74#_c_1756_n 0.0128f $X=13.955 $Y=2.227
+ $X2=0 $Y2=0
cc_590 N_A_547_301#_c_594_n N_A_2385_74#_c_1757_n 0.00281727f $X=13.185 $Y=2.465
+ $X2=0 $Y2=0
cc_591 N_A_547_301#_c_596_n N_A_2385_74#_c_1757_n 0.0076835f $X=13.955 $Y=2.227
+ $X2=0 $Y2=0
cc_592 N_A_547_301#_c_585_n N_A_2385_74#_c_1757_n 0.0151547f $X=14.015 $Y=1.665
+ $X2=0 $Y2=0
cc_593 N_A_547_301#_c_581_n N_A_2385_74#_c_1748_n 0.00628125f $X=13.215 $Y=0.94
+ $X2=0 $Y2=0
cc_594 N_A_547_301#_c_583_n N_A_2385_74#_c_1748_n 0.0185585f $X=13.29 $Y=2.05
+ $X2=0 $Y2=0
cc_595 N_A_547_301#_c_585_n N_A_2385_74#_c_1748_n 0.0173314f $X=14.015 $Y=1.665
+ $X2=0 $Y2=0
cc_596 N_A_547_301#_c_594_n N_A_2385_74#_c_1759_n 6.92651e-19 $X=13.185 $Y=2.465
+ $X2=0 $Y2=0
cc_597 N_A_547_301#_c_583_n N_A_2385_74#_c_1759_n 0.00338995f $X=13.29 $Y=2.05
+ $X2=0 $Y2=0
cc_598 N_A_547_301#_c_596_n N_A_2385_74#_c_1759_n 0.0336224f $X=13.955 $Y=2.227
+ $X2=0 $Y2=0
cc_599 N_A_547_301#_c_598_n N_A_2385_74#_c_1759_n 0.0101588f $X=14.165 $Y=2.075
+ $X2=0 $Y2=0
cc_600 N_A_547_301#_c_585_n N_A_2385_74#_c_1759_n 0.016712f $X=14.015 $Y=1.665
+ $X2=0 $Y2=0
cc_601 N_A_547_301#_c_587_n N_A_2385_74#_c_1759_n 0.00131723f $X=14.16 $Y=1.665
+ $X2=0 $Y2=0
cc_602 N_A_547_301#_c_583_n N_A_2385_74#_c_1749_n 0.00227385f $X=13.29 $Y=2.05
+ $X2=0 $Y2=0
cc_603 N_A_547_301#_c_585_n N_A_2385_74#_c_1749_n 0.0106844f $X=14.015 $Y=1.665
+ $X2=0 $Y2=0
cc_604 N_A_547_301#_c_587_n N_A_2385_74#_c_1749_n 0.00108878f $X=14.16 $Y=1.665
+ $X2=0 $Y2=0
cc_605 N_A_547_301#_c_588_n N_A_2385_74#_c_1749_n 0.00819793f $X=14.16 $Y=1.665
+ $X2=0 $Y2=0
cc_606 N_A_547_301#_c_591_n N_A_2385_74#_c_1749_n 0.00737285f $X=14.165 $Y=1.55
+ $X2=0 $Y2=0
cc_607 N_A_547_301#_c_594_n N_A_2385_74#_c_1761_n 0.00111922f $X=13.185 $Y=2.465
+ $X2=0 $Y2=0
cc_608 N_A_547_301#_c_583_n N_A_2385_74#_c_1761_n 0.00636734f $X=13.29 $Y=2.05
+ $X2=0 $Y2=0
cc_609 N_A_547_301#_c_596_n N_A_2385_74#_c_1761_n 0.0128325f $X=13.955 $Y=2.227
+ $X2=0 $Y2=0
cc_610 N_A_547_301#_c_585_n N_A_2385_74#_c_1761_n 0.00230187f $X=14.015 $Y=1.665
+ $X2=0 $Y2=0
cc_611 N_A_547_301#_c_583_n N_A_2385_74#_c_1750_n 0.00108101f $X=13.29 $Y=2.05
+ $X2=0 $Y2=0
cc_612 N_A_547_301#_c_584_n N_A_2385_74#_c_1750_n 0.0010601f $X=14.09 $Y=0.58
+ $X2=0 $Y2=0
cc_613 N_A_547_301#_c_585_n N_A_2385_74#_c_1750_n 0.00627479f $X=14.015 $Y=1.665
+ $X2=0 $Y2=0
cc_614 N_A_547_301#_c_591_n N_A_2385_74#_c_1750_n 0.0242399f $X=14.165 $Y=1.55
+ $X2=0 $Y2=0
cc_615 N_A_547_301#_c_593_n N_A_27_74#_c_1895_n 0.0131657f $X=3.085 $Y=2.24
+ $X2=0 $Y2=0
cc_616 N_A_547_301#_c_585_n N_A_27_74#_c_1895_n 0.00373727f $X=14.015 $Y=1.665
+ $X2=0 $Y2=0
cc_617 N_A_547_301#_c_586_n N_A_27_74#_c_1895_n 0.00324212f $X=2.785 $Y=1.665
+ $X2=0 $Y2=0
cc_618 N_A_547_301#_c_589_n N_A_27_74#_c_1895_n 0.0148801f $X=2.9 $Y=1.67 $X2=0
+ $Y2=0
cc_619 N_A_547_301#_c_590_n N_A_27_74#_c_1895_n 0.00432537f $X=3.085 $Y=1.67
+ $X2=0 $Y2=0
cc_620 N_A_547_301#_M1038_g N_A_27_74#_c_1885_n 0.0139482f $X=2.84 $Y=0.765
+ $X2=0 $Y2=0
cc_621 N_A_547_301#_c_593_n N_A_27_74#_c_1897_n 0.00870642f $X=3.085 $Y=2.24
+ $X2=0 $Y2=0
cc_622 N_A_547_301#_M1038_g N_A_27_74#_c_1886_n 0.00499775f $X=2.84 $Y=0.765
+ $X2=0 $Y2=0
cc_623 N_A_547_301#_c_593_n N_A_27_74#_c_1886_n 0.00116727f $X=3.085 $Y=2.24
+ $X2=0 $Y2=0
cc_624 N_A_547_301#_c_585_n N_A_27_74#_c_1886_n 0.0165869f $X=14.015 $Y=1.665
+ $X2=0 $Y2=0
cc_625 N_A_547_301#_c_586_n N_A_27_74#_c_1886_n 3.76633e-19 $X=2.785 $Y=1.665
+ $X2=0 $Y2=0
cc_626 N_A_547_301#_c_589_n N_A_27_74#_c_1886_n 0.0239479f $X=2.9 $Y=1.67 $X2=0
+ $Y2=0
cc_627 N_A_547_301#_c_590_n N_A_27_74#_c_1886_n 0.0181596f $X=3.085 $Y=1.67
+ $X2=0 $Y2=0
cc_628 N_A_547_301#_M1038_g N_A_27_74#_c_1888_n 0.00693595f $X=2.84 $Y=0.765
+ $X2=0 $Y2=0
cc_629 N_A_547_301#_c_585_n N_A_27_74#_c_1888_n 0.00829724f $X=14.015 $Y=1.665
+ $X2=0 $Y2=0
cc_630 N_A_547_301#_c_589_n N_A_27_74#_c_1888_n 0.011369f $X=2.9 $Y=1.67 $X2=0
+ $Y2=0
cc_631 N_A_547_301#_c_590_n N_A_27_74#_c_1888_n 0.00835602f $X=3.085 $Y=1.67
+ $X2=0 $Y2=0
cc_632 N_A_547_301#_c_593_n N_A_27_74#_c_1900_n 0.00166465f $X=3.085 $Y=2.24
+ $X2=0 $Y2=0
cc_633 N_A_547_301#_c_585_n N_A_27_74#_c_1900_n 0.00276825f $X=14.015 $Y=1.665
+ $X2=0 $Y2=0
cc_634 N_A_547_301#_c_596_n N_VPWR_M1021_d 0.00294158f $X=13.955 $Y=2.227 $X2=0
+ $Y2=0
cc_635 N_A_547_301#_c_593_n N_VPWR_c_2009_n 0.00150486f $X=3.085 $Y=2.24 $X2=0
+ $Y2=0
cc_636 N_A_547_301#_c_594_n N_VPWR_c_2015_n 0.0103114f $X=13.185 $Y=2.465 $X2=0
+ $Y2=0
cc_637 N_A_547_301#_c_596_n N_VPWR_c_2015_n 0.0260798f $X=13.955 $Y=2.227 $X2=0
+ $Y2=0
cc_638 N_A_547_301#_c_597_n N_VPWR_c_2015_n 0.0132122f $X=14.12 $Y=2.465 $X2=0
+ $Y2=0
cc_639 N_A_547_301#_c_593_n N_VPWR_c_2028_n 0.0044174f $X=3.085 $Y=2.24 $X2=0
+ $Y2=0
cc_640 N_A_547_301#_c_594_n N_VPWR_c_2030_n 0.00461464f $X=13.185 $Y=2.465 $X2=0
+ $Y2=0
cc_641 N_A_547_301#_c_597_n N_VPWR_c_2031_n 0.0145938f $X=14.12 $Y=2.465 $X2=0
+ $Y2=0
cc_642 N_A_547_301#_c_593_n N_VPWR_c_2007_n 0.00544287f $X=3.085 $Y=2.24 $X2=0
+ $Y2=0
cc_643 N_A_547_301#_c_594_n N_VPWR_c_2007_n 0.0098334f $X=13.185 $Y=2.465 $X2=0
+ $Y2=0
cc_644 N_A_547_301#_c_597_n N_VPWR_c_2007_n 0.0120466f $X=14.12 $Y=2.465 $X2=0
+ $Y2=0
cc_645 N_A_547_301#_c_585_n N_A_669_111#_c_2178_n 0.00392161f $X=14.015 $Y=1.665
+ $X2=0 $Y2=0
cc_646 N_A_547_301#_c_593_n N_A_669_111#_c_2191_n 5.18926e-19 $X=3.085 $Y=2.24
+ $X2=0 $Y2=0
cc_647 N_A_547_301#_c_585_n N_A_669_111#_c_2170_n 0.00659142f $X=14.015 $Y=1.665
+ $X2=0 $Y2=0
cc_648 N_A_547_301#_c_585_n N_A_669_111#_c_2171_n 0.00245341f $X=14.015 $Y=1.665
+ $X2=0 $Y2=0
cc_649 N_A_547_301#_c_585_n N_A_669_111#_c_2172_n 0.0190561f $X=14.015 $Y=1.665
+ $X2=0 $Y2=0
cc_650 N_A_547_301#_c_585_n N_A_669_111#_c_2182_n 0.0198621f $X=14.015 $Y=1.665
+ $X2=0 $Y2=0
cc_651 N_A_547_301#_c_585_n N_A_669_111#_c_2183_n 0.0143314f $X=14.015 $Y=1.665
+ $X2=0 $Y2=0
cc_652 N_A_547_301#_c_585_n N_A_669_111#_c_2173_n 0.0287955f $X=14.015 $Y=1.665
+ $X2=0 $Y2=0
cc_653 N_A_547_301#_c_585_n N_A_669_111#_c_2174_n 0.00573242f $X=14.015 $Y=1.665
+ $X2=0 $Y2=0
cc_654 N_A_547_301#_c_585_n N_A_669_111#_c_2199_n 0.00419251f $X=14.015 $Y=1.665
+ $X2=0 $Y2=0
cc_655 N_A_547_301#_c_585_n N_A_669_111#_c_2176_n 0.0057569f $X=14.015 $Y=1.665
+ $X2=0 $Y2=0
cc_656 N_A_547_301#_M1038_g N_A_669_111#_c_2177_n 6.24576e-19 $X=2.84 $Y=0.765
+ $X2=0 $Y2=0
cc_657 N_A_547_301#_c_585_n N_A_669_111#_c_2177_n 0.0179445f $X=14.015 $Y=1.665
+ $X2=0 $Y2=0
cc_658 N_A_547_301#_c_585_n N_A_669_111#_c_2188_n 0.00120995f $X=14.015 $Y=1.665
+ $X2=0 $Y2=0
cc_659 N_A_547_301#_c_585_n N_A_669_111#_c_2189_n 0.00614572f $X=14.015 $Y=1.665
+ $X2=0 $Y2=0
cc_660 N_A_547_301#_c_597_n Q 0.0462676f $X=14.12 $Y=2.465 $X2=0 $Y2=0
cc_661 N_A_547_301#_c_584_n Q 0.123443f $X=14.09 $Y=0.58 $X2=0 $Y2=0
cc_662 N_A_547_301#_c_599_n Q 0.0249916f $X=14.12 $Y=2.227 $X2=0 $Y2=0
cc_663 N_A_547_301#_c_587_n Q 0.0070972f $X=14.16 $Y=1.665 $X2=0 $Y2=0
cc_664 N_A_547_301#_M1038_g N_VGND_c_2388_n 0.0018473f $X=2.84 $Y=0.765 $X2=0
+ $Y2=0
cc_665 N_A_547_301#_c_585_n N_VGND_c_2389_n 0.00632657f $X=14.015 $Y=1.665 $X2=0
+ $Y2=0
cc_666 N_A_547_301#_M1038_g N_VGND_c_2396_n 0.00436277f $X=2.84 $Y=0.765 $X2=0
+ $Y2=0
cc_667 N_A_547_301#_c_584_n N_VGND_c_2406_n 0.0156722f $X=14.09 $Y=0.58 $X2=0
+ $Y2=0
cc_668 N_A_547_301#_c_580_n N_VGND_c_2411_n 0.00383152f $X=12.75 $Y=0.865 $X2=0
+ $Y2=0
cc_669 N_A_547_301#_c_580_n N_VGND_c_2412_n 0.0105517f $X=12.75 $Y=0.865 $X2=0
+ $Y2=0
cc_670 N_A_547_301#_c_581_n N_VGND_c_2412_n 0.0039717f $X=13.215 $Y=0.94 $X2=0
+ $Y2=0
cc_671 N_A_547_301#_c_584_n N_VGND_c_2412_n 0.0103991f $X=14.09 $Y=0.58 $X2=0
+ $Y2=0
cc_672 N_A_547_301#_M1038_g N_VGND_c_2413_n 0.00489211f $X=2.84 $Y=0.765 $X2=0
+ $Y2=0
cc_673 N_A_547_301#_c_580_n N_VGND_c_2413_n 0.00367447f $X=12.75 $Y=0.865 $X2=0
+ $Y2=0
cc_674 N_A_547_301#_c_584_n N_VGND_c_2413_n 0.0130167f $X=14.09 $Y=0.58 $X2=0
+ $Y2=0
cc_675 N_A_639_85#_c_829_n N_SCD_c_934_n 0.0256258f $X=5.655 $Y=1.92 $X2=0 $Y2=0
cc_676 N_A_639_85#_c_833_n N_SCD_c_934_n 0.01197f $X=5.49 $Y=2 $X2=0 $Y2=0
cc_677 N_A_639_85#_c_828_n N_SCD_c_935_n 0.0439755f $X=5.58 $Y=2.2 $X2=0 $Y2=0
cc_678 N_A_639_85#_c_833_n SCD 0.0249062f $X=5.49 $Y=2 $X2=0 $Y2=0
cc_679 N_A_639_85#_c_825_n SCD 0.0193362f $X=5.655 $Y=1.58 $X2=0 $Y2=0
cc_680 N_A_639_85#_c_826_n SCD 0.00113478f $X=5.655 $Y=1.58 $X2=0 $Y2=0
cc_681 N_A_639_85#_c_833_n N_SCD_c_933_n 0.00104612f $X=5.49 $Y=2 $X2=0 $Y2=0
cc_682 N_A_639_85#_c_825_n N_SCD_c_933_n 0.00227755f $X=5.655 $Y=1.58 $X2=0
+ $Y2=0
cc_683 N_A_639_85#_c_826_n N_SCD_c_933_n 0.0256258f $X=5.655 $Y=1.58 $X2=0 $Y2=0
cc_684 N_A_639_85#_c_832_n N_SCE_c_984_n 3.50071e-19 $X=4.1 $Y=2.255 $X2=-0.19
+ $Y2=-0.245
cc_685 N_A_639_85#_c_836_n N_SCE_c_984_n 0.00100796f $X=4.285 $Y=2.495 $X2=-0.19
+ $Y2=-0.245
cc_686 N_A_639_85#_c_836_n N_SCE_c_985_n 0.00201936f $X=4.285 $Y=2.495 $X2=0
+ $Y2=0
cc_687 N_A_639_85#_c_823_n N_SCE_c_977_n 0.00765996f $X=3.995 $Y=1.78 $X2=0
+ $Y2=0
cc_688 N_A_639_85#_c_824_n N_SCE_c_977_n 0.0210125f $X=3.995 $Y=1.78 $X2=0 $Y2=0
cc_689 N_A_639_85#_c_832_n N_SCE_c_977_n 0.00371596f $X=4.1 $Y=2.255 $X2=0 $Y2=0
cc_690 N_A_639_85#_c_833_n N_SCE_c_977_n 0.0188979f $X=5.49 $Y=2 $X2=0 $Y2=0
cc_691 N_A_639_85#_c_832_n N_SCE_M1027_g 0.00171259f $X=4.1 $Y=2.255 $X2=0 $Y2=0
cc_692 N_A_639_85#_c_836_n N_SCE_M1027_g 0.00320341f $X=4.285 $Y=2.495 $X2=0
+ $Y2=0
cc_693 N_A_639_85#_c_821_n N_SCE_M1041_g 0.00283026f $X=3.995 $Y=0.42 $X2=0
+ $Y2=0
cc_694 N_A_639_85#_c_822_n N_SCE_M1041_g 0.0203141f $X=3.995 $Y=0.42 $X2=0 $Y2=0
cc_695 N_A_639_85#_c_823_n N_SCE_M1041_g 0.00321528f $X=3.995 $Y=1.78 $X2=0
+ $Y2=0
cc_696 N_A_639_85#_c_827_n N_SCE_M1041_g 0.00549407f $X=4.41 $Y=0.805 $X2=0
+ $Y2=0
cc_697 N_A_639_85#_c_820_n SCE 4.01743e-19 $X=3.995 $Y=1.125 $X2=0 $Y2=0
cc_698 N_A_639_85#_c_823_n SCE 0.0216259f $X=3.995 $Y=1.78 $X2=0 $Y2=0
cc_699 N_A_639_85#_c_833_n SCE 0.00603941f $X=5.49 $Y=2 $X2=0 $Y2=0
cc_700 N_A_639_85#_c_827_n SCE 0.0111158f $X=4.41 $Y=0.805 $X2=0 $Y2=0
cc_701 N_A_639_85#_c_820_n N_SCE_c_983_n 0.0175073f $X=3.995 $Y=1.125 $X2=0
+ $Y2=0
cc_702 N_A_639_85#_c_823_n N_SCE_c_983_n 0.00197408f $X=3.995 $Y=1.78 $X2=0
+ $Y2=0
cc_703 N_A_639_85#_c_833_n N_SCE_c_983_n 8.54293e-19 $X=5.49 $Y=2 $X2=0 $Y2=0
cc_704 N_A_639_85#_c_827_n N_SCE_c_983_n 9.58107e-19 $X=4.41 $Y=0.805 $X2=0
+ $Y2=0
cc_705 N_A_639_85#_c_826_n N_CLK_c_1064_n 0.00897042f $X=5.655 $Y=1.58 $X2=0
+ $Y2=0
cc_706 N_A_639_85#_c_817_n N_A_27_74#_c_1885_n 0.00736452f $X=3.27 $Y=1.05 $X2=0
+ $Y2=0
cc_707 N_A_639_85#_c_819_n N_A_27_74#_c_1885_n 0.0040964f $X=3.345 $Y=1.125
+ $X2=0 $Y2=0
cc_708 N_A_639_85#_c_819_n N_A_27_74#_c_1886_n 9.15581e-19 $X=3.345 $Y=1.125
+ $X2=0 $Y2=0
cc_709 N_A_639_85#_c_818_n N_A_27_74#_c_1888_n 0.00362743f $X=3.83 $Y=1.125
+ $X2=0 $Y2=0
cc_710 N_A_639_85#_c_819_n N_A_27_74#_c_1888_n 0.00908768f $X=3.345 $Y=1.125
+ $X2=0 $Y2=0
cc_711 N_A_639_85#_c_828_n N_VPWR_c_2010_n 0.00149083f $X=5.58 $Y=2.2 $X2=0
+ $Y2=0
cc_712 N_A_639_85#_c_828_n N_VPWR_c_2011_n 0.00328352f $X=5.58 $Y=2.2 $X2=0
+ $Y2=0
cc_713 N_A_639_85#_c_828_n N_VPWR_c_2029_n 0.00530811f $X=5.58 $Y=2.2 $X2=0
+ $Y2=0
cc_714 N_A_639_85#_c_828_n N_VPWR_c_2007_n 0.005315f $X=5.58 $Y=2.2 $X2=0 $Y2=0
cc_715 N_A_639_85#_c_824_n N_A_669_111#_c_2178_n 5.59349e-19 $X=3.995 $Y=1.78
+ $X2=0 $Y2=0
cc_716 N_A_639_85#_c_836_n N_A_669_111#_c_2178_n 0.0358182f $X=4.285 $Y=2.495
+ $X2=0 $Y2=0
cc_717 N_A_639_85#_M1027_s N_A_669_111#_c_2179_n 0.00259631f $X=4.155 $Y=2.275
+ $X2=0 $Y2=0
cc_718 N_A_639_85#_c_836_n N_A_669_111#_c_2179_n 0.0265612f $X=4.285 $Y=2.495
+ $X2=0 $Y2=0
cc_719 N_A_639_85#_c_836_n N_A_669_111#_c_2209_n 0.0230808f $X=4.285 $Y=2.495
+ $X2=0 $Y2=0
cc_720 N_A_639_85#_c_833_n N_A_669_111#_c_2180_n 0.0134263f $X=5.49 $Y=2 $X2=0
+ $Y2=0
cc_721 N_A_639_85#_c_836_n N_A_669_111#_c_2180_n 0.0140999f $X=4.285 $Y=2.495
+ $X2=0 $Y2=0
cc_722 N_A_639_85#_c_825_n N_A_669_111#_c_2170_n 0.00177664f $X=5.655 $Y=1.58
+ $X2=0 $Y2=0
cc_723 N_A_639_85#_c_833_n N_A_669_111#_c_2171_n 3.08031e-19 $X=5.49 $Y=2 $X2=0
+ $Y2=0
cc_724 N_A_639_85#_c_825_n N_A_669_111#_c_2171_n 0.0253172f $X=5.655 $Y=1.58
+ $X2=0 $Y2=0
cc_725 N_A_639_85#_c_826_n N_A_669_111#_c_2171_n 0.0023541f $X=5.655 $Y=1.58
+ $X2=0 $Y2=0
cc_726 N_A_639_85#_c_828_n N_A_669_111#_c_2172_n 0.00156538f $X=5.58 $Y=2.2
+ $X2=0 $Y2=0
cc_727 N_A_639_85#_c_829_n N_A_669_111#_c_2172_n 0.00342548f $X=5.655 $Y=1.92
+ $X2=0 $Y2=0
cc_728 N_A_639_85#_c_833_n N_A_669_111#_c_2172_n 0.0135436f $X=5.49 $Y=2 $X2=0
+ $Y2=0
cc_729 N_A_639_85#_c_825_n N_A_669_111#_c_2172_n 0.0365245f $X=5.655 $Y=1.58
+ $X2=0 $Y2=0
cc_730 N_A_639_85#_c_826_n N_A_669_111#_c_2172_n 0.00527835f $X=5.655 $Y=1.58
+ $X2=0 $Y2=0
cc_731 N_A_639_85#_c_817_n N_A_669_111#_c_2176_n 0.00326664f $X=3.27 $Y=1.05
+ $X2=0 $Y2=0
cc_732 N_A_639_85#_c_818_n N_A_669_111#_c_2176_n 0.00571191f $X=3.83 $Y=1.125
+ $X2=0 $Y2=0
cc_733 N_A_639_85#_c_821_n N_A_669_111#_c_2176_n 0.00549356f $X=3.995 $Y=0.42
+ $X2=0 $Y2=0
cc_734 N_A_639_85#_c_822_n N_A_669_111#_c_2176_n 0.00535604f $X=3.995 $Y=0.42
+ $X2=0 $Y2=0
cc_735 N_A_639_85#_c_827_n N_A_669_111#_c_2176_n 0.0337923f $X=4.41 $Y=0.805
+ $X2=0 $Y2=0
cc_736 N_A_639_85#_c_817_n N_A_669_111#_c_2177_n 4.66894e-19 $X=3.27 $Y=1.05
+ $X2=0 $Y2=0
cc_737 N_A_639_85#_c_818_n N_A_669_111#_c_2177_n 0.0149432f $X=3.83 $Y=1.125
+ $X2=0 $Y2=0
cc_738 N_A_639_85#_c_823_n N_A_669_111#_c_2177_n 0.065605f $X=3.995 $Y=1.78
+ $X2=0 $Y2=0
cc_739 N_A_639_85#_c_824_n N_A_669_111#_c_2177_n 0.0123304f $X=3.995 $Y=1.78
+ $X2=0 $Y2=0
cc_740 N_A_639_85#_c_832_n N_A_669_111#_c_2177_n 0.00902514f $X=4.1 $Y=2.255
+ $X2=0 $Y2=0
cc_741 N_A_639_85#_c_835_n N_A_669_111#_c_2177_n 0.0142217f $X=4.045 $Y=2 $X2=0
+ $Y2=0
cc_742 N_A_639_85#_c_836_n N_A_669_111#_c_2177_n 0.00217874f $X=4.285 $Y=2.495
+ $X2=0 $Y2=0
cc_743 N_A_639_85#_c_828_n N_A_669_111#_c_2187_n 0.00772809f $X=5.58 $Y=2.2
+ $X2=0 $Y2=0
cc_744 N_A_639_85#_c_828_n N_A_669_111#_c_2188_n 0.011357f $X=5.58 $Y=2.2 $X2=0
+ $Y2=0
cc_745 N_A_639_85#_c_829_n N_A_669_111#_c_2188_n 4.52395e-19 $X=5.655 $Y=1.92
+ $X2=0 $Y2=0
cc_746 N_A_639_85#_c_833_n N_A_669_111#_c_2188_n 0.0808616f $X=5.49 $Y=2 $X2=0
+ $Y2=0
cc_747 N_A_639_85#_c_828_n N_A_669_111#_c_2189_n 0.00227738f $X=5.58 $Y=2.2
+ $X2=0 $Y2=0
cc_748 N_A_639_85#_c_829_n N_A_669_111#_c_2189_n 0.00152938f $X=5.655 $Y=1.92
+ $X2=0 $Y2=0
cc_749 N_A_639_85#_c_821_n N_VGND_c_2389_n 0.0120611f $X=3.995 $Y=0.42 $X2=0
+ $Y2=0
cc_750 N_A_639_85#_c_827_n N_VGND_c_2389_n 0.0168669f $X=4.41 $Y=0.805 $X2=0
+ $Y2=0
cc_751 N_A_639_85#_c_817_n N_VGND_c_2396_n 0.00436277f $X=3.27 $Y=1.05 $X2=0
+ $Y2=0
cc_752 N_A_639_85#_c_821_n N_VGND_c_2396_n 0.0181555f $X=3.995 $Y=0.42 $X2=0
+ $Y2=0
cc_753 N_A_639_85#_c_822_n N_VGND_c_2396_n 0.00451316f $X=3.995 $Y=0.42 $X2=0
+ $Y2=0
cc_754 N_A_639_85#_c_827_n N_VGND_c_2396_n 0.00805954f $X=4.41 $Y=0.805 $X2=0
+ $Y2=0
cc_755 N_A_639_85#_c_817_n N_VGND_c_2413_n 0.00489211f $X=3.27 $Y=1.05 $X2=0
+ $Y2=0
cc_756 N_A_639_85#_c_821_n N_VGND_c_2413_n 0.0104822f $X=3.995 $Y=0.42 $X2=0
+ $Y2=0
cc_757 N_A_639_85#_c_822_n N_VGND_c_2413_n 0.00274137f $X=3.995 $Y=0.42 $X2=0
+ $Y2=0
cc_758 N_A_639_85#_c_827_n N_VGND_c_2413_n 0.0117476f $X=4.41 $Y=0.805 $X2=0
+ $Y2=0
cc_759 N_SCD_c_935_n N_SCE_c_985_n 0.00100522f $X=5.19 $Y=2.2 $X2=0 $Y2=0
cc_760 N_SCD_c_934_n N_SCE_c_977_n 0.00601231f $X=5.19 $Y=2.11 $X2=0 $Y2=0
cc_761 SCD N_SCE_c_977_n 0.00385693f $X=4.955 $Y=1.21 $X2=0 $Y2=0
cc_762 N_SCD_c_933_n N_SCE_c_977_n 0.00810881f $X=5.115 $Y=1.58 $X2=0 $Y2=0
cc_763 N_SCD_c_935_n N_SCE_c_988_n 0.00601231f $X=5.19 $Y=2.2 $X2=0 $Y2=0
cc_764 N_SCD_c_935_n N_SCE_M1027_g 0.0111767f $X=5.19 $Y=2.2 $X2=0 $Y2=0
cc_765 N_SCD_M1031_g N_SCE_M1041_g 0.0142089f $X=5.055 $Y=0.835 $X2=0 $Y2=0
cc_766 N_SCD_M1031_g N_SCE_c_979_n 0.00894529f $X=5.055 $Y=0.835 $X2=0 $Y2=0
cc_767 N_SCD_M1031_g N_SCE_M1028_g 0.0397809f $X=5.055 $Y=0.835 $X2=0 $Y2=0
cc_768 N_SCD_M1031_g SCE 2.73422e-19 $X=5.055 $Y=0.835 $X2=0 $Y2=0
cc_769 SCD SCE 0.023703f $X=4.955 $Y=1.21 $X2=0 $Y2=0
cc_770 N_SCD_M1031_g N_SCE_c_983_n 0.0117224f $X=5.055 $Y=0.835 $X2=0 $Y2=0
cc_771 SCD N_SCE_c_983_n 0.00202477f $X=4.955 $Y=1.21 $X2=0 $Y2=0
cc_772 N_SCD_c_933_n N_SCE_c_983_n 0.00561978f $X=5.115 $Y=1.58 $X2=0 $Y2=0
cc_773 N_SCD_c_935_n N_VPWR_c_2010_n 0.00959399f $X=5.19 $Y=2.2 $X2=0 $Y2=0
cc_774 N_SCD_c_935_n N_VPWR_c_2029_n 0.00489294f $X=5.19 $Y=2.2 $X2=0 $Y2=0
cc_775 N_SCD_c_935_n N_VPWR_c_2007_n 0.00481893f $X=5.19 $Y=2.2 $X2=0 $Y2=0
cc_776 N_SCD_c_935_n N_A_669_111#_c_2179_n 3.76568e-19 $X=5.19 $Y=2.2 $X2=0
+ $Y2=0
cc_777 N_SCD_c_935_n N_A_669_111#_c_2209_n 0.00283455f $X=5.19 $Y=2.2 $X2=0
+ $Y2=0
cc_778 N_SCD_M1031_g N_A_669_111#_c_2169_n 0.00142522f $X=5.055 $Y=0.835 $X2=0
+ $Y2=0
cc_779 N_SCD_M1031_g N_A_669_111#_c_2171_n 0.00103169f $X=5.055 $Y=0.835 $X2=0
+ $Y2=0
cc_780 SCD N_A_669_111#_c_2171_n 0.00545313f $X=4.955 $Y=1.21 $X2=0 $Y2=0
cc_781 N_SCD_c_935_n N_A_669_111#_c_2187_n 0.00141291f $X=5.19 $Y=2.2 $X2=0
+ $Y2=0
cc_782 N_SCD_c_935_n N_A_669_111#_c_2188_n 0.0160628f $X=5.19 $Y=2.2 $X2=0 $Y2=0
cc_783 N_SCD_c_935_n N_A_669_111#_c_2189_n 3.56261e-19 $X=5.19 $Y=2.2 $X2=0
+ $Y2=0
cc_784 N_SCD_M1031_g N_VGND_c_2389_n 0.0101548f $X=5.055 $Y=0.835 $X2=0 $Y2=0
cc_785 SCD N_VGND_c_2389_n 0.00441285f $X=4.955 $Y=1.21 $X2=0 $Y2=0
cc_786 N_SCD_M1031_g N_VGND_c_2413_n 7.97988e-19 $X=5.055 $Y=0.835 $X2=0 $Y2=0
cc_787 N_SCE_c_984_n N_A_27_74#_c_1897_n 0.00161473f $X=3.535 $Y=3.03 $X2=0
+ $Y2=0
cc_788 N_SCE_c_984_n N_A_27_74#_c_1886_n 7.32247e-19 $X=3.535 $Y=3.03 $X2=0
+ $Y2=0
cc_789 N_SCE_c_984_n N_A_27_74#_c_1900_n 7.52181e-19 $X=3.535 $Y=3.03 $X2=0
+ $Y2=0
cc_790 N_SCE_c_985_n N_VPWR_c_2010_n 0.00310923f $X=4.42 $Y=3.105 $X2=0 $Y2=0
cc_791 N_SCE_M1027_g N_VPWR_c_2010_n 0.00117443f $X=4.51 $Y=2.595 $X2=0 $Y2=0
cc_792 N_SCE_c_986_n N_VPWR_c_2028_n 0.0240584f $X=3.61 $Y=3.105 $X2=0 $Y2=0
cc_793 N_SCE_c_985_n N_VPWR_c_2007_n 0.0252128f $X=4.42 $Y=3.105 $X2=0 $Y2=0
cc_794 N_SCE_c_986_n N_VPWR_c_2007_n 0.0100661f $X=3.61 $Y=3.105 $X2=0 $Y2=0
cc_795 N_SCE_c_984_n N_A_669_111#_c_2178_n 0.00196983f $X=3.535 $Y=3.03 $X2=0
+ $Y2=0
cc_796 N_SCE_M1027_g N_A_669_111#_c_2178_n 0.00450557f $X=4.51 $Y=2.595 $X2=0
+ $Y2=0
cc_797 N_SCE_c_984_n N_A_669_111#_c_2249_n 0.00538071f $X=3.535 $Y=3.03 $X2=0
+ $Y2=0
cc_798 N_SCE_c_985_n N_A_669_111#_c_2179_n 0.0217336f $X=4.42 $Y=3.105 $X2=0
+ $Y2=0
cc_799 N_SCE_M1027_g N_A_669_111#_c_2179_n 0.00872278f $X=4.51 $Y=2.595 $X2=0
+ $Y2=0
cc_800 N_SCE_c_984_n N_A_669_111#_c_2191_n 0.00373701f $X=3.535 $Y=3.03 $X2=0
+ $Y2=0
cc_801 N_SCE_c_985_n N_A_669_111#_c_2191_n 0.00837949f $X=4.42 $Y=3.105 $X2=0
+ $Y2=0
cc_802 N_SCE_c_986_n N_A_669_111#_c_2191_n 0.0013142f $X=3.61 $Y=3.105 $X2=0
+ $Y2=0
cc_803 N_SCE_M1027_g N_A_669_111#_c_2209_n 0.0162802f $X=4.51 $Y=2.595 $X2=0
+ $Y2=0
cc_804 N_SCE_c_988_n N_A_669_111#_c_2180_n 4.69291e-19 $X=4.51 $Y=2.2 $X2=0
+ $Y2=0
cc_805 N_SCE_M1027_g N_A_669_111#_c_2180_n 0.00578626f $X=4.51 $Y=2.595 $X2=0
+ $Y2=0
cc_806 N_SCE_M1028_g N_A_669_111#_c_2169_n 0.0096824f $X=5.415 $Y=0.835 $X2=0
+ $Y2=0
cc_807 N_SCE_M1028_g N_A_669_111#_c_2171_n 0.00463814f $X=5.415 $Y=0.835 $X2=0
+ $Y2=0
cc_808 N_SCE_c_984_n N_A_669_111#_c_2177_n 0.00415211f $X=3.535 $Y=3.03 $X2=0
+ $Y2=0
cc_809 N_SCE_c_977_n N_A_669_111#_c_2177_n 5.38351e-19 $X=4.51 $Y=2.11 $X2=0
+ $Y2=0
cc_810 N_SCE_M1041_g N_VGND_c_2389_n 0.00563898f $X=4.625 $Y=0.835 $X2=0 $Y2=0
cc_811 N_SCE_c_979_n N_VGND_c_2389_n 0.0197475f $X=5.34 $Y=0.18 $X2=0 $Y2=0
cc_812 N_SCE_M1028_g N_VGND_c_2389_n 0.00666558f $X=5.415 $Y=0.835 $X2=0 $Y2=0
cc_813 N_SCE_c_979_n N_VGND_c_2390_n 0.0112176f $X=5.34 $Y=0.18 $X2=0 $Y2=0
cc_814 N_SCE_M1028_g N_VGND_c_2390_n 5.64384e-19 $X=5.415 $Y=0.835 $X2=0 $Y2=0
cc_815 N_SCE_c_980_n N_VGND_c_2396_n 0.00768659f $X=4.7 $Y=0.18 $X2=0 $Y2=0
cc_816 N_SCE_c_979_n N_VGND_c_2398_n 0.0177114f $X=5.34 $Y=0.18 $X2=0 $Y2=0
cc_817 N_SCE_c_979_n N_VGND_c_2413_n 0.0299336f $X=5.34 $Y=0.18 $X2=0 $Y2=0
cc_818 N_SCE_c_980_n N_VGND_c_2413_n 0.0106458f $X=4.7 $Y=0.18 $X2=0 $Y2=0
cc_819 N_CLK_c_1064_n N_A_1295_74#_M1007_g 0.00432739f $X=6.55 $Y=1.705 $X2=0
+ $Y2=0
cc_820 N_CLK_c_1064_n N_A_1295_74#_c_1336_n 0.00943695f $X=6.55 $Y=1.705 $X2=0
+ $Y2=0
cc_821 N_CLK_c_1063_n N_A_1295_74#_c_1339_n 0.00601567f $X=6.4 $Y=1.22 $X2=0
+ $Y2=0
cc_822 N_CLK_c_1063_n N_A_1295_74#_c_1340_n 0.00268707f $X=6.4 $Y=1.22 $X2=0
+ $Y2=0
cc_823 N_CLK_c_1064_n N_A_1295_74#_c_1340_n 0.00558976f $X=6.55 $Y=1.705 $X2=0
+ $Y2=0
cc_824 CLK N_A_1295_74#_c_1340_n 0.027973f $X=6.395 $Y=1.21 $X2=0 $Y2=0
cc_825 N_CLK_c_1063_n N_A_1295_74#_c_1341_n 0.00344395f $X=6.4 $Y=1.22 $X2=0
+ $Y2=0
cc_826 N_CLK_c_1064_n N_A_1295_74#_c_1341_n 0.00103195f $X=6.55 $Y=1.705 $X2=0
+ $Y2=0
cc_827 CLK N_A_1295_74#_c_1341_n 0.0139664f $X=6.395 $Y=1.21 $X2=0 $Y2=0
cc_828 N_CLK_c_1064_n N_A_1295_74#_c_1361_n 0.00796702f $X=6.55 $Y=1.705 $X2=0
+ $Y2=0
cc_829 CLK N_A_1295_74#_c_1361_n 0.00235215f $X=6.395 $Y=1.21 $X2=0 $Y2=0
cc_830 N_CLK_c_1064_n N_VPWR_c_2011_n 0.0184328f $X=6.55 $Y=1.705 $X2=0 $Y2=0
cc_831 N_CLK_c_1064_n N_VPWR_c_2022_n 0.00479724f $X=6.55 $Y=1.705 $X2=0 $Y2=0
cc_832 N_CLK_c_1064_n N_VPWR_c_2007_n 0.00477621f $X=6.55 $Y=1.705 $X2=0 $Y2=0
cc_833 N_CLK_c_1063_n N_A_669_111#_c_2169_n 0.00384469f $X=6.4 $Y=1.22 $X2=0
+ $Y2=0
cc_834 N_CLK_c_1063_n N_A_669_111#_c_2170_n 0.00420168f $X=6.4 $Y=1.22 $X2=0
+ $Y2=0
cc_835 CLK N_A_669_111#_c_2170_n 0.00545388f $X=6.395 $Y=1.21 $X2=0 $Y2=0
cc_836 N_CLK_c_1064_n N_A_669_111#_c_2172_n 0.0141174f $X=6.55 $Y=1.705 $X2=0
+ $Y2=0
cc_837 CLK N_A_669_111#_c_2172_n 0.022885f $X=6.395 $Y=1.21 $X2=0 $Y2=0
cc_838 N_CLK_c_1064_n N_A_669_111#_c_2182_n 0.017191f $X=6.55 $Y=1.705 $X2=0
+ $Y2=0
cc_839 N_CLK_c_1064_n N_A_669_111#_c_2187_n 0.00369503f $X=6.55 $Y=1.705 $X2=0
+ $Y2=0
cc_840 N_CLK_c_1064_n N_A_669_111#_c_2189_n 0.00260589f $X=6.55 $Y=1.705 $X2=0
+ $Y2=0
cc_841 N_CLK_c_1063_n N_VGND_c_2390_n 0.00776346f $X=6.4 $Y=1.22 $X2=0 $Y2=0
cc_842 N_CLK_c_1063_n N_VGND_c_2391_n 0.00334136f $X=6.4 $Y=1.22 $X2=0 $Y2=0
cc_843 N_CLK_c_1063_n N_VGND_c_2400_n 0.00434272f $X=6.4 $Y=1.22 $X2=0 $Y2=0
cc_844 N_CLK_c_1063_n N_VGND_c_2413_n 0.00825443f $X=6.4 $Y=1.22 $X2=0 $Y2=0
cc_845 N_A_1492_74#_c_1099_n N_A_1295_74#_M1007_g 0.00168241f $X=7.6 $Y=0.515
+ $X2=0 $Y2=0
cc_846 N_A_1492_74#_c_1101_n N_A_1295_74#_M1007_g 0.00266901f $X=7.765 $Y=0.34
+ $X2=0 $Y2=0
cc_847 N_A_1492_74#_c_1099_n N_A_1295_74#_c_1330_n 0.00257504f $X=7.6 $Y=0.515
+ $X2=0 $Y2=0
cc_848 N_A_1492_74#_c_1123_n N_A_1295_74#_c_1344_n 0.00533913f $X=8.405 $Y=1.99
+ $X2=0 $Y2=0
cc_849 N_A_1492_74#_c_1102_n N_A_1295_74#_c_1344_n 9.21756e-19 $X=8.49 $Y=1.82
+ $X2=0 $Y2=0
cc_850 N_A_1492_74#_c_1127_n N_A_1295_74#_c_1344_n 0.00571652f $X=8.575 $Y=2.17
+ $X2=0 $Y2=0
cc_851 N_A_1492_74#_c_1123_n N_A_1295_74#_c_1331_n 0.0126221f $X=8.405 $Y=1.99
+ $X2=0 $Y2=0
cc_852 N_A_1492_74#_c_1096_n N_A_1295_74#_M1026_g 0.0134631f $X=9.045 $Y=1.015
+ $X2=0 $Y2=0
cc_853 N_A_1492_74#_c_1099_n N_A_1295_74#_M1026_g 0.00317282f $X=7.6 $Y=0.515
+ $X2=0 $Y2=0
cc_854 N_A_1492_74#_c_1100_n N_A_1295_74#_M1026_g 0.00929412f $X=8.405 $Y=0.34
+ $X2=0 $Y2=0
cc_855 N_A_1492_74#_c_1102_n N_A_1295_74#_M1026_g 0.0306171f $X=8.49 $Y=1.82
+ $X2=0 $Y2=0
cc_856 N_A_1492_74#_c_1117_n N_A_1295_74#_M1026_g 0.00206916f $X=8.49 $Y=0.34
+ $X2=0 $Y2=0
cc_857 N_A_1492_74#_c_1123_n N_A_1295_74#_c_1333_n 0.00197072f $X=8.405 $Y=1.99
+ $X2=0 $Y2=0
cc_858 N_A_1492_74#_c_1102_n N_A_1295_74#_c_1333_n 0.0077472f $X=8.49 $Y=1.82
+ $X2=0 $Y2=0
cc_859 N_A_1492_74#_c_1105_n N_A_1295_74#_c_1333_n 7.2465e-19 $X=9.175 $Y=1.18
+ $X2=0 $Y2=0
cc_860 N_A_1492_74#_c_1106_n N_A_1295_74#_c_1333_n 0.0181826f $X=9.175 $Y=1.18
+ $X2=0 $Y2=0
cc_861 N_A_1492_74#_c_1127_n N_A_1295_74#_c_1333_n 0.00583382f $X=8.575 $Y=2.17
+ $X2=0 $Y2=0
cc_862 N_A_1492_74#_c_1120_n N_A_1295_74#_c_1348_n 0.0134813f $X=8.875 $Y=2.465
+ $X2=0 $Y2=0
cc_863 N_A_1492_74#_c_1106_n N_A_1295_74#_c_1348_n 2.22258e-19 $X=9.175 $Y=1.18
+ $X2=0 $Y2=0
cc_864 N_A_1492_74#_c_1127_n N_A_1295_74#_c_1348_n 0.0161286f $X=8.575 $Y=2.17
+ $X2=0 $Y2=0
cc_865 N_A_1492_74#_M1024_g N_A_1295_74#_c_1334_n 0.0212555f $X=11.85 $Y=0.69
+ $X2=0 $Y2=0
cc_866 N_A_1492_74#_c_1098_n N_A_1295_74#_c_1334_n 0.0139323f $X=12.765 $Y=2.375
+ $X2=0 $Y2=0
cc_867 N_A_1492_74#_c_1122_n N_A_1295_74#_c_1334_n 0.0119156f $X=12.765 $Y=2.465
+ $X2=0 $Y2=0
cc_868 N_A_1492_74#_c_1114_n N_A_1295_74#_c_1334_n 5.46133e-19 $X=11.76 $Y=1.635
+ $X2=0 $Y2=0
cc_869 N_A_1492_74#_c_1115_n N_A_1295_74#_c_1334_n 0.00269787f $X=11.76 $Y=1.635
+ $X2=0 $Y2=0
cc_870 N_A_1492_74#_c_1116_n N_A_1295_74#_c_1334_n 0.00470669f $X=12.675
+ $Y=1.195 $X2=0 $Y2=0
cc_871 N_A_1492_74#_c_1118_n N_A_1295_74#_c_1334_n 3.16884e-19 $X=12.84 $Y=1.195
+ $X2=0 $Y2=0
cc_872 N_A_1492_74#_c_1119_n N_A_1295_74#_c_1334_n 0.021347f $X=12.84 $Y=1.39
+ $X2=0 $Y2=0
cc_873 N_A_1492_74#_M1024_g N_A_1295_74#_M1034_g 0.0277654f $X=11.85 $Y=0.69
+ $X2=0 $Y2=0
cc_874 N_A_1492_74#_c_1114_n N_A_1295_74#_M1034_g 7.5412e-19 $X=11.76 $Y=1.635
+ $X2=0 $Y2=0
cc_875 N_A_1492_74#_c_1116_n N_A_1295_74#_M1034_g 0.0115589f $X=12.675 $Y=1.195
+ $X2=0 $Y2=0
cc_876 N_A_1492_74#_c_1118_n N_A_1295_74#_M1034_g 0.00143858f $X=12.84 $Y=1.195
+ $X2=0 $Y2=0
cc_877 N_A_1492_74#_c_1119_n N_A_1295_74#_M1034_g 0.0110933f $X=12.84 $Y=1.39
+ $X2=0 $Y2=0
cc_878 N_A_1492_74#_c_1102_n N_A_1295_74#_c_1338_n 0.00354171f $X=8.49 $Y=1.82
+ $X2=0 $Y2=0
cc_879 N_A_1492_74#_c_1127_n N_A_1295_74#_c_1338_n 0.0180723f $X=8.575 $Y=2.17
+ $X2=0 $Y2=0
cc_880 N_A_1492_74#_c_1099_n N_A_1295_74#_c_1340_n 0.00243738f $X=7.6 $Y=0.515
+ $X2=0 $Y2=0
cc_881 N_A_1492_74#_c_1114_n N_A_1295_74#_c_1358_n 0.00891578f $X=11.76 $Y=1.635
+ $X2=0 $Y2=0
cc_882 N_A_1492_74#_c_1115_n N_A_1295_74#_c_1358_n 0.00311532f $X=11.76 $Y=1.635
+ $X2=0 $Y2=0
cc_883 N_A_1492_74#_c_1098_n N_A_1295_74#_c_1360_n 5.35617e-19 $X=12.765
+ $Y=2.375 $X2=0 $Y2=0
cc_884 N_A_1492_74#_c_1114_n N_A_1295_74#_c_1360_n 0.00484942f $X=11.76 $Y=1.635
+ $X2=0 $Y2=0
cc_885 N_A_1492_74#_c_1115_n N_A_1295_74#_c_1360_n 3.94242e-19 $X=11.76 $Y=1.635
+ $X2=0 $Y2=0
cc_886 N_A_1492_74#_M1024_g N_A_1295_74#_c_1342_n 0.00163405f $X=11.85 $Y=0.69
+ $X2=0 $Y2=0
cc_887 N_A_1492_74#_c_1114_n N_A_1295_74#_c_1342_n 0.0212328f $X=11.76 $Y=1.635
+ $X2=0 $Y2=0
cc_888 N_A_1492_74#_c_1116_n N_A_1295_74#_c_1342_n 0.0301176f $X=12.675 $Y=1.195
+ $X2=0 $Y2=0
cc_889 N_A_1492_74#_c_1118_n N_A_1295_74#_c_1342_n 0.00676121f $X=12.84 $Y=1.195
+ $X2=0 $Y2=0
cc_890 N_A_1492_74#_c_1119_n N_A_1295_74#_c_1342_n 0.00218464f $X=12.84 $Y=1.39
+ $X2=0 $Y2=0
cc_891 N_A_1492_74#_c_1108_n N_A_1910_71#_M1033_d 0.0039106f $X=10.85 $Y=0.34
+ $X2=-0.19 $Y2=-0.245
cc_892 N_A_1492_74#_c_1096_n N_A_1910_71#_M1029_g 0.0152991f $X=9.045 $Y=1.015
+ $X2=0 $Y2=0
cc_893 N_A_1492_74#_c_1103_n N_A_1910_71#_M1029_g 7.05141e-19 $X=9.085 $Y=0.34
+ $X2=0 $Y2=0
cc_894 N_A_1492_74#_c_1104_n N_A_1910_71#_M1029_g 0.00533215f $X=9.17 $Y=0.85
+ $X2=0 $Y2=0
cc_895 N_A_1492_74#_c_1105_n N_A_1910_71#_M1029_g 0.00170347f $X=9.175 $Y=1.18
+ $X2=0 $Y2=0
cc_896 N_A_1492_74#_c_1106_n N_A_1910_71#_M1029_g 0.0210364f $X=9.175 $Y=1.18
+ $X2=0 $Y2=0
cc_897 N_A_1492_74#_c_1107_n N_A_1910_71#_M1029_g 0.0138944f $X=10.17 $Y=0.935
+ $X2=0 $Y2=0
cc_898 N_A_1492_74#_c_1202_p N_A_1910_71#_M1029_g 0.00310164f $X=10.255 $Y=0.85
+ $X2=0 $Y2=0
cc_899 N_A_1492_74#_M1024_g N_A_1910_71#_c_1532_n 0.0606927f $X=11.85 $Y=0.69
+ $X2=0 $Y2=0
cc_900 N_A_1492_74#_c_1108_n N_A_1910_71#_c_1532_n 6.63977e-19 $X=10.85 $Y=0.34
+ $X2=0 $Y2=0
cc_901 N_A_1492_74#_c_1110_n N_A_1910_71#_c_1532_n 0.00423957f $X=10.935
+ $Y=0.855 $X2=0 $Y2=0
cc_902 N_A_1492_74#_c_1111_n N_A_1910_71#_c_1532_n 0.0123071f $X=11.56 $Y=0.94
+ $X2=0 $Y2=0
cc_903 N_A_1492_74#_c_1113_n N_A_1910_71#_c_1532_n 0.00500819f $X=11.71 $Y=1.28
+ $X2=0 $Y2=0
cc_904 N_A_1492_74#_c_1107_n N_A_1910_71#_c_1533_n 0.0329621f $X=10.17 $Y=0.935
+ $X2=0 $Y2=0
cc_905 N_A_1492_74#_c_1107_n N_A_1910_71#_c_1534_n 0.00750114f $X=10.17 $Y=0.935
+ $X2=0 $Y2=0
cc_906 N_A_1492_74#_c_1108_n N_A_1910_71#_c_1534_n 0.0127109f $X=10.85 $Y=0.34
+ $X2=0 $Y2=0
cc_907 N_A_1492_74#_c_1110_n N_A_1910_71#_c_1534_n 0.0191933f $X=10.935 $Y=0.855
+ $X2=0 $Y2=0
cc_908 N_A_1492_74#_c_1112_n N_A_1910_71#_c_1534_n 0.0141515f $X=11.02 $Y=0.94
+ $X2=0 $Y2=0
cc_909 N_A_1492_74#_M1024_g N_A_1910_71#_c_1537_n 2.40007e-19 $X=11.85 $Y=0.69
+ $X2=0 $Y2=0
cc_910 N_A_1492_74#_c_1111_n N_A_1910_71#_c_1537_n 0.0266054f $X=11.56 $Y=0.94
+ $X2=0 $Y2=0
cc_911 N_A_1492_74#_c_1112_n N_A_1910_71#_c_1537_n 0.0139074f $X=11.02 $Y=0.94
+ $X2=0 $Y2=0
cc_912 N_A_1492_74#_c_1113_n N_A_1910_71#_c_1537_n 0.00703577f $X=11.71 $Y=1.28
+ $X2=0 $Y2=0
cc_913 N_A_1492_74#_c_1114_n N_A_1910_71#_c_1537_n 0.0198463f $X=11.76 $Y=1.635
+ $X2=0 $Y2=0
cc_914 N_A_1492_74#_c_1108_n N_A_1910_71#_c_1538_n 0.00306165f $X=10.85 $Y=0.34
+ $X2=0 $Y2=0
cc_915 N_A_1492_74#_c_1111_n N_A_1910_71#_c_1538_n 0.0111491f $X=11.56 $Y=0.94
+ $X2=0 $Y2=0
cc_916 N_A_1492_74#_c_1112_n N_A_1910_71#_c_1538_n 0.00459457f $X=11.02 $Y=0.94
+ $X2=0 $Y2=0
cc_917 N_A_1492_74#_c_1105_n N_A_1910_71#_c_1539_n 0.00963411f $X=9.175 $Y=1.18
+ $X2=0 $Y2=0
cc_918 N_A_1492_74#_c_1106_n N_A_1910_71#_c_1539_n 5.34652e-19 $X=9.175 $Y=1.18
+ $X2=0 $Y2=0
cc_919 N_A_1492_74#_c_1107_n N_A_1910_71#_c_1539_n 0.0232123f $X=10.17 $Y=0.935
+ $X2=0 $Y2=0
cc_920 N_A_1492_74#_c_1107_n N_A_1910_71#_c_1540_n 0.00529227f $X=10.17 $Y=0.935
+ $X2=0 $Y2=0
cc_921 N_A_1492_74#_M1024_g N_A_1910_71#_c_1541_n 0.00606257f $X=11.85 $Y=0.69
+ $X2=0 $Y2=0
cc_922 N_A_1492_74#_c_1113_n N_A_1910_71#_c_1541_n 0.00706327f $X=11.71 $Y=1.28
+ $X2=0 $Y2=0
cc_923 N_A_1492_74#_c_1114_n N_A_1910_71#_c_1541_n 0.00623901f $X=11.76 $Y=1.635
+ $X2=0 $Y2=0
cc_924 N_A_1492_74#_c_1115_n N_A_1910_71#_c_1541_n 0.0210318f $X=11.76 $Y=1.635
+ $X2=0 $Y2=0
cc_925 N_A_1492_74#_c_1102_n N_A_1688_97#_M1026_d 0.0043242f $X=8.49 $Y=1.82
+ $X2=-0.19 $Y2=-0.245
cc_926 N_A_1492_74#_c_1107_n N_A_1688_97#_M1033_g 0.0057601f $X=10.17 $Y=0.935
+ $X2=0 $Y2=0
cc_927 N_A_1492_74#_c_1202_p N_A_1688_97#_M1033_g 0.0115776f $X=10.255 $Y=0.85
+ $X2=0 $Y2=0
cc_928 N_A_1492_74#_c_1108_n N_A_1688_97#_M1033_g 0.0112842f $X=10.85 $Y=0.34
+ $X2=0 $Y2=0
cc_929 N_A_1492_74#_c_1109_n N_A_1688_97#_M1033_g 0.00331918f $X=10.34 $Y=0.34
+ $X2=0 $Y2=0
cc_930 N_A_1492_74#_c_1110_n N_A_1688_97#_M1033_g 0.00328401f $X=10.935 $Y=0.855
+ $X2=0 $Y2=0
cc_931 N_A_1492_74#_c_1096_n N_A_1688_97#_c_1644_n 0.0049112f $X=9.045 $Y=1.015
+ $X2=0 $Y2=0
cc_932 N_A_1492_74#_c_1102_n N_A_1688_97#_c_1644_n 0.076172f $X=8.49 $Y=1.82
+ $X2=0 $Y2=0
cc_933 N_A_1492_74#_c_1103_n N_A_1688_97#_c_1644_n 0.012971f $X=9.085 $Y=0.34
+ $X2=0 $Y2=0
cc_934 N_A_1492_74#_c_1105_n N_A_1688_97#_c_1644_n 0.0239141f $X=9.175 $Y=1.18
+ $X2=0 $Y2=0
cc_935 N_A_1492_74#_c_1239_p N_A_1688_97#_c_1644_n 0.0114261f $X=9.212 $Y=0.935
+ $X2=0 $Y2=0
cc_936 N_A_1492_74#_c_1120_n N_A_1688_97#_c_1648_n 0.00231881f $X=8.875 $Y=2.465
+ $X2=0 $Y2=0
cc_937 N_A_1492_74#_c_1102_n N_A_1688_97#_c_1649_n 0.0119523f $X=8.49 $Y=1.82
+ $X2=0 $Y2=0
cc_938 N_A_1492_74#_c_1106_n N_A_1688_97#_c_1649_n 4.32369e-19 $X=9.175 $Y=1.18
+ $X2=0 $Y2=0
cc_939 N_A_1492_74#_c_1127_n N_A_1688_97#_c_1649_n 0.00205522f $X=8.575 $Y=2.17
+ $X2=0 $Y2=0
cc_940 N_A_1492_74#_c_1123_n N_A_1688_97#_c_1650_n 0.0366921f $X=8.405 $Y=1.99
+ $X2=0 $Y2=0
cc_941 N_A_1492_74#_c_1102_n N_A_1688_97#_c_1650_n 0.00162478f $X=8.49 $Y=1.82
+ $X2=0 $Y2=0
cc_942 N_A_1492_74#_c_1127_n N_A_1688_97#_c_1650_n 0.0101106f $X=8.575 $Y=2.17
+ $X2=0 $Y2=0
cc_943 N_A_1492_74#_c_1120_n N_A_1688_97#_c_1651_n 0.00682301f $X=8.875 $Y=2.465
+ $X2=0 $Y2=0
cc_944 N_A_1492_74#_c_1127_n N_A_1688_97#_c_1651_n 0.00347676f $X=8.575 $Y=2.17
+ $X2=0 $Y2=0
cc_945 N_A_1492_74#_c_1105_n N_A_1688_97#_c_1646_n 0.00969703f $X=9.175 $Y=1.18
+ $X2=0 $Y2=0
cc_946 N_A_1492_74#_c_1106_n N_A_1688_97#_c_1646_n 0.00142351f $X=9.175 $Y=1.18
+ $X2=0 $Y2=0
cc_947 N_A_1492_74#_c_1107_n N_A_1688_97#_c_1646_n 0.00388953f $X=10.17 $Y=0.935
+ $X2=0 $Y2=0
cc_948 N_A_1492_74#_M1024_g N_A_2385_74#_c_1825_n 0.00277139f $X=11.85 $Y=0.69
+ $X2=0 $Y2=0
cc_949 N_A_1492_74#_c_1116_n N_A_2385_74#_c_1825_n 0.0243071f $X=12.675 $Y=1.195
+ $X2=0 $Y2=0
cc_950 N_A_1492_74#_M1024_g N_A_2385_74#_c_1746_n 0.00725553f $X=11.85 $Y=0.69
+ $X2=0 $Y2=0
cc_951 N_A_1492_74#_c_1116_n N_A_2385_74#_c_1747_n 0.0323431f $X=12.675 $Y=1.195
+ $X2=0 $Y2=0
cc_952 N_A_1492_74#_c_1118_n N_A_2385_74#_c_1747_n 0.0254828f $X=12.84 $Y=1.195
+ $X2=0 $Y2=0
cc_953 N_A_1492_74#_c_1119_n N_A_2385_74#_c_1747_n 2.90561e-19 $X=12.84 $Y=1.39
+ $X2=0 $Y2=0
cc_954 N_A_1492_74#_c_1098_n N_A_2385_74#_c_1755_n 0.0133233f $X=12.765 $Y=2.375
+ $X2=0 $Y2=0
cc_955 N_A_1492_74#_c_1116_n N_A_2385_74#_c_1755_n 0.0030736f $X=12.675 $Y=1.195
+ $X2=0 $Y2=0
cc_956 N_A_1492_74#_c_1118_n N_A_2385_74#_c_1755_n 0.00774105f $X=12.84 $Y=1.195
+ $X2=0 $Y2=0
cc_957 N_A_1492_74#_c_1098_n N_A_2385_74#_c_1756_n 0.00697239f $X=12.765
+ $Y=2.375 $X2=0 $Y2=0
cc_958 N_A_1492_74#_c_1122_n N_A_2385_74#_c_1756_n 0.0239509f $X=12.765 $Y=2.465
+ $X2=0 $Y2=0
cc_959 N_A_1492_74#_c_1098_n N_A_2385_74#_c_1757_n 0.00595698f $X=12.765
+ $Y=2.375 $X2=0 $Y2=0
cc_960 N_A_1492_74#_c_1118_n N_A_2385_74#_c_1757_n 0.0109926f $X=12.84 $Y=1.195
+ $X2=0 $Y2=0
cc_961 N_A_1492_74#_c_1119_n N_A_2385_74#_c_1757_n 0.00103738f $X=12.84 $Y=1.39
+ $X2=0 $Y2=0
cc_962 N_A_1492_74#_c_1098_n N_A_2385_74#_c_1748_n 0.00249889f $X=12.765
+ $Y=2.375 $X2=0 $Y2=0
cc_963 N_A_1492_74#_c_1118_n N_A_2385_74#_c_1748_n 0.0339179f $X=12.84 $Y=1.195
+ $X2=0 $Y2=0
cc_964 N_A_1492_74#_c_1119_n N_A_2385_74#_c_1748_n 0.00174016f $X=12.84 $Y=1.39
+ $X2=0 $Y2=0
cc_965 N_A_1492_74#_c_1120_n N_VPWR_c_2024_n 0.00444483f $X=8.875 $Y=2.465 $X2=0
+ $Y2=0
cc_966 N_A_1492_74#_c_1122_n N_VPWR_c_2030_n 0.00332301f $X=12.765 $Y=2.465
+ $X2=0 $Y2=0
cc_967 N_A_1492_74#_c_1120_n N_VPWR_c_2007_n 0.00508527f $X=8.875 $Y=2.465 $X2=0
+ $Y2=0
cc_968 N_A_1492_74#_c_1122_n N_VPWR_c_2007_n 0.0052991f $X=12.765 $Y=2.465 $X2=0
+ $Y2=0
cc_969 N_A_1492_74#_c_1123_n N_A_669_111#_c_2183_n 0.0148492f $X=8.405 $Y=1.99
+ $X2=0 $Y2=0
cc_970 N_A_1492_74#_c_1102_n N_A_669_111#_c_2183_n 0.00321631f $X=8.49 $Y=1.82
+ $X2=0 $Y2=0
cc_971 N_A_1492_74#_c_1123_n N_A_669_111#_c_2173_n 0.018064f $X=8.405 $Y=1.99
+ $X2=0 $Y2=0
cc_972 N_A_1492_74#_c_1102_n N_A_669_111#_c_2173_n 0.0128904f $X=8.49 $Y=1.82
+ $X2=0 $Y2=0
cc_973 N_A_1492_74#_c_1099_n N_A_669_111#_c_2174_n 0.00697011f $X=7.6 $Y=0.515
+ $X2=0 $Y2=0
cc_974 N_A_1492_74#_M1030_d N_A_669_111#_c_2199_n 0.00488381f $X=7.975 $Y=1.84
+ $X2=0 $Y2=0
cc_975 N_A_1492_74#_c_1120_n N_A_669_111#_c_2199_n 5.2088e-19 $X=8.875 $Y=2.465
+ $X2=0 $Y2=0
cc_976 N_A_1492_74#_c_1123_n N_A_669_111#_c_2199_n 0.0136228f $X=8.405 $Y=1.99
+ $X2=0 $Y2=0
cc_977 N_A_1492_74#_c_1127_n N_A_669_111#_c_2199_n 0.00209126f $X=8.575 $Y=2.17
+ $X2=0 $Y2=0
cc_978 N_A_1492_74#_c_1099_n N_A_669_111#_c_2175_n 0.035665f $X=7.6 $Y=0.515
+ $X2=0 $Y2=0
cc_979 N_A_1492_74#_c_1100_n N_A_669_111#_c_2175_n 0.019204f $X=8.405 $Y=0.34
+ $X2=0 $Y2=0
cc_980 N_A_1492_74#_c_1102_n N_A_669_111#_c_2175_n 0.0528515f $X=8.49 $Y=1.82
+ $X2=0 $Y2=0
cc_981 N_A_1492_74#_M1030_d N_A_669_111#_c_2282_n 0.00458284f $X=7.975 $Y=1.84
+ $X2=0 $Y2=0
cc_982 N_A_1492_74#_c_1120_n N_A_669_111#_c_2282_n 0.0033043f $X=8.875 $Y=2.465
+ $X2=0 $Y2=0
cc_983 N_A_1492_74#_M1030_d N_A_669_111#_c_2184_n 0.00188412f $X=7.975 $Y=1.84
+ $X2=0 $Y2=0
cc_984 N_A_1492_74#_M1030_d N_A_669_111#_c_2185_n 0.00222941f $X=7.975 $Y=1.84
+ $X2=0 $Y2=0
cc_985 N_A_1492_74#_c_1120_n N_A_669_111#_c_2185_n 0.0035741f $X=8.875 $Y=2.465
+ $X2=0 $Y2=0
cc_986 N_A_1492_74#_c_1123_n N_A_669_111#_c_2185_n 0.0186228f $X=8.405 $Y=1.99
+ $X2=0 $Y2=0
cc_987 N_A_1492_74#_c_1127_n N_A_669_111#_c_2185_n 0.00452329f $X=8.575 $Y=2.17
+ $X2=0 $Y2=0
cc_988 N_A_1492_74#_c_1107_n N_VGND_M1029_d 0.00712543f $X=10.17 $Y=0.935 $X2=0
+ $Y2=0
cc_989 N_A_1492_74#_c_1202_p N_VGND_M1029_d 0.00491722f $X=10.255 $Y=0.85 $X2=0
+ $Y2=0
cc_990 N_A_1492_74#_c_1109_n N_VGND_M1029_d 5.36892e-19 $X=10.34 $Y=0.34 $X2=0
+ $Y2=0
cc_991 N_A_1492_74#_c_1111_n N_VGND_M1022_s 0.00389007f $X=11.56 $Y=0.94 $X2=0
+ $Y2=0
cc_992 N_A_1492_74#_c_1101_n N_VGND_c_2391_n 0.0112234f $X=7.765 $Y=0.34 $X2=0
+ $Y2=0
cc_993 N_A_1492_74#_c_1103_n N_VGND_c_2392_n 0.00700152f $X=9.085 $Y=0.34 $X2=0
+ $Y2=0
cc_994 N_A_1492_74#_c_1104_n N_VGND_c_2392_n 0.00537476f $X=9.17 $Y=0.85 $X2=0
+ $Y2=0
cc_995 N_A_1492_74#_c_1107_n N_VGND_c_2392_n 0.0192736f $X=10.17 $Y=0.935 $X2=0
+ $Y2=0
cc_996 N_A_1492_74#_c_1202_p N_VGND_c_2392_n 0.0190358f $X=10.255 $Y=0.85 $X2=0
+ $Y2=0
cc_997 N_A_1492_74#_c_1109_n N_VGND_c_2392_n 0.0145685f $X=10.34 $Y=0.34 $X2=0
+ $Y2=0
cc_998 N_A_1492_74#_M1024_g N_VGND_c_2393_n 0.00148407f $X=11.85 $Y=0.69 $X2=0
+ $Y2=0
cc_999 N_A_1492_74#_c_1108_n N_VGND_c_2393_n 0.0146661f $X=10.85 $Y=0.34 $X2=0
+ $Y2=0
cc_1000 N_A_1492_74#_c_1110_n N_VGND_c_2393_n 0.0197547f $X=10.935 $Y=0.855
+ $X2=0 $Y2=0
cc_1001 N_A_1492_74#_c_1111_n N_VGND_c_2393_n 0.0150542f $X=11.56 $Y=0.94 $X2=0
+ $Y2=0
cc_1002 N_A_1492_74#_c_1096_n N_VGND_c_2404_n 7.53287e-19 $X=9.045 $Y=1.015
+ $X2=0 $Y2=0
cc_1003 N_A_1492_74#_c_1100_n N_VGND_c_2404_n 0.0411694f $X=8.405 $Y=0.34 $X2=0
+ $Y2=0
cc_1004 N_A_1492_74#_c_1101_n N_VGND_c_2404_n 0.0179217f $X=7.765 $Y=0.34 $X2=0
+ $Y2=0
cc_1005 N_A_1492_74#_c_1103_n N_VGND_c_2404_n 0.0449818f $X=9.085 $Y=0.34 $X2=0
+ $Y2=0
cc_1006 N_A_1492_74#_c_1117_n N_VGND_c_2404_n 0.0121867f $X=8.49 $Y=0.34 $X2=0
+ $Y2=0
cc_1007 N_A_1492_74#_c_1108_n N_VGND_c_2405_n 0.0446499f $X=10.85 $Y=0.34 $X2=0
+ $Y2=0
cc_1008 N_A_1492_74#_c_1109_n N_VGND_c_2405_n 0.0120637f $X=10.34 $Y=0.34 $X2=0
+ $Y2=0
cc_1009 N_A_1492_74#_M1024_g N_VGND_c_2411_n 0.00434272f $X=11.85 $Y=0.69 $X2=0
+ $Y2=0
cc_1010 N_A_1492_74#_M1024_g N_VGND_c_2413_n 0.00821463f $X=11.85 $Y=0.69 $X2=0
+ $Y2=0
cc_1011 N_A_1492_74#_c_1100_n N_VGND_c_2413_n 0.0240545f $X=8.405 $Y=0.34 $X2=0
+ $Y2=0
cc_1012 N_A_1492_74#_c_1101_n N_VGND_c_2413_n 0.00971942f $X=7.765 $Y=0.34 $X2=0
+ $Y2=0
cc_1013 N_A_1492_74#_c_1103_n N_VGND_c_2413_n 0.025776f $X=9.085 $Y=0.34 $X2=0
+ $Y2=0
cc_1014 N_A_1492_74#_c_1107_n N_VGND_c_2413_n 0.0201846f $X=10.17 $Y=0.935 $X2=0
+ $Y2=0
cc_1015 N_A_1492_74#_c_1108_n N_VGND_c_2413_n 0.0252533f $X=10.85 $Y=0.34 $X2=0
+ $Y2=0
cc_1016 N_A_1492_74#_c_1109_n N_VGND_c_2413_n 0.00644906f $X=10.34 $Y=0.34 $X2=0
+ $Y2=0
cc_1017 N_A_1492_74#_c_1111_n N_VGND_c_2413_n 0.00983886f $X=11.56 $Y=0.94 $X2=0
+ $Y2=0
cc_1018 N_A_1492_74#_c_1113_n N_VGND_c_2413_n 0.00657755f $X=11.71 $Y=1.28 $X2=0
+ $Y2=0
cc_1019 N_A_1492_74#_c_1117_n N_VGND_c_2413_n 0.00660921f $X=8.49 $Y=0.34 $X2=0
+ $Y2=0
cc_1020 N_A_1492_74#_c_1239_p N_VGND_c_2413_n 0.00322096f $X=9.212 $Y=0.935
+ $X2=0 $Y2=0
cc_1021 N_A_1492_74#_c_1104_n A_1824_97# 0.00486153f $X=9.17 $Y=0.85 $X2=-0.19
+ $Y2=-0.245
cc_1022 N_A_1492_74#_c_1107_n A_1824_97# 0.00308187f $X=10.17 $Y=0.935 $X2=-0.19
+ $Y2=-0.245
cc_1023 N_A_1492_74#_c_1239_p A_1824_97# 0.00193682f $X=9.212 $Y=0.935 $X2=-0.19
+ $Y2=-0.245
cc_1024 N_A_1492_74#_c_1113_n A_2313_74# 0.00230895f $X=11.71 $Y=1.28 $X2=-0.19
+ $Y2=-0.245
cc_1025 N_A_1295_74#_c_1358_n N_A_1910_71#_M1039_d 0.00731573f $X=12.03 $Y=2.475
+ $X2=0 $Y2=0
cc_1026 N_A_1295_74#_c_1333_n N_A_1910_71#_c_1530_n 0.0102336f $X=9.175 $Y=1.69
+ $X2=0 $Y2=0
cc_1027 N_A_1295_74#_c_1348_n N_A_1910_71#_c_1530_n 0.0291411f $X=9.375 $Y=2.465
+ $X2=0 $Y2=0
cc_1028 N_A_1295_74#_c_1356_n N_A_1910_71#_c_1530_n 0.0073441f $X=9.485 $Y=2.09
+ $X2=0 $Y2=0
cc_1029 N_A_1295_74#_c_1357_n N_A_1910_71#_c_1530_n 0.00392779f $X=9.57 $Y=2.39
+ $X2=0 $Y2=0
cc_1030 N_A_1295_74#_c_1348_n N_A_1910_71#_c_1543_n 0.026729f $X=9.375 $Y=2.465
+ $X2=0 $Y2=0
cc_1031 N_A_1295_74#_c_1358_n N_A_1910_71#_c_1543_n 0.014972f $X=12.03 $Y=2.475
+ $X2=0 $Y2=0
cc_1032 N_A_1295_74#_c_1358_n N_A_1910_71#_c_1545_n 0.0202137f $X=12.03 $Y=2.475
+ $X2=0 $Y2=0
cc_1033 N_A_1295_74#_c_1360_n N_A_1910_71#_c_1545_n 0.0122277f $X=12.115 $Y=2.39
+ $X2=0 $Y2=0
cc_1034 N_A_1295_74#_c_1358_n N_A_1910_71#_c_1547_n 0.027361f $X=12.03 $Y=2.475
+ $X2=0 $Y2=0
cc_1035 N_A_1295_74#_c_1358_n N_A_1688_97#_c_1642_n 0.0173821f $X=12.03 $Y=2.475
+ $X2=0 $Y2=0
cc_1036 N_A_1295_74#_M1026_g N_A_1688_97#_c_1644_n 0.00342569f $X=8.365 $Y=0.695
+ $X2=0 $Y2=0
cc_1037 N_A_1295_74#_c_1333_n N_A_1688_97#_c_1644_n 0.00411041f $X=9.175 $Y=1.69
+ $X2=0 $Y2=0
cc_1038 N_A_1295_74#_c_1348_n N_A_1688_97#_c_1648_n 0.00778975f $X=9.375
+ $Y=2.465 $X2=0 $Y2=0
cc_1039 N_A_1295_74#_c_1333_n N_A_1688_97#_c_1649_n 0.00995496f $X=9.175 $Y=1.69
+ $X2=0 $Y2=0
cc_1040 N_A_1295_74#_c_1347_n N_A_1688_97#_c_1650_n 0.0059401f $X=9.25 $Y=1.925
+ $X2=0 $Y2=0
cc_1041 N_A_1295_74#_c_1348_n N_A_1688_97#_c_1650_n 0.00240421f $X=9.375
+ $Y=2.465 $X2=0 $Y2=0
cc_1042 N_A_1295_74#_c_1356_n N_A_1688_97#_c_1650_n 0.0200573f $X=9.485 $Y=2.09
+ $X2=0 $Y2=0
cc_1043 N_A_1295_74#_c_1357_n N_A_1688_97#_c_1650_n 0.00602344f $X=9.57 $Y=2.39
+ $X2=0 $Y2=0
cc_1044 N_A_1295_74#_c_1333_n N_A_1688_97#_c_1651_n 4.82451e-19 $X=9.175 $Y=1.69
+ $X2=0 $Y2=0
cc_1045 N_A_1295_74#_c_1348_n N_A_1688_97#_c_1651_n 0.00772562f $X=9.375
+ $Y=2.465 $X2=0 $Y2=0
cc_1046 N_A_1295_74#_c_1356_n N_A_1688_97#_c_1651_n 0.0112687f $X=9.485 $Y=2.09
+ $X2=0 $Y2=0
cc_1047 N_A_1295_74#_c_1359_n N_A_1688_97#_c_1651_n 0.0136934f $X=9.655 $Y=2.475
+ $X2=0 $Y2=0
cc_1048 N_A_1295_74#_c_1358_n N_A_1688_97#_c_1645_n 0.00566213f $X=12.03
+ $Y=2.475 $X2=0 $Y2=0
cc_1049 N_A_1295_74#_c_1333_n N_A_1688_97#_c_1646_n 0.00959259f $X=9.175 $Y=1.69
+ $X2=0 $Y2=0
cc_1050 N_A_1295_74#_c_1347_n N_A_1688_97#_c_1646_n 0.00322616f $X=9.25 $Y=1.925
+ $X2=0 $Y2=0
cc_1051 N_A_1295_74#_c_1348_n N_A_1688_97#_c_1646_n 0.0045192f $X=9.375 $Y=2.465
+ $X2=0 $Y2=0
cc_1052 N_A_1295_74#_c_1356_n N_A_1688_97#_c_1646_n 0.0332493f $X=9.485 $Y=2.09
+ $X2=0 $Y2=0
cc_1053 N_A_1295_74#_c_1358_n N_A_1688_97#_c_1646_n 0.0134405f $X=12.03 $Y=2.475
+ $X2=0 $Y2=0
cc_1054 N_A_1295_74#_M1034_g N_A_2385_74#_c_1746_n 0.00236994f $X=12.36 $Y=0.58
+ $X2=0 $Y2=0
cc_1055 N_A_1295_74#_M1034_g N_A_2385_74#_c_1747_n 0.0117469f $X=12.36 $Y=0.58
+ $X2=0 $Y2=0
cc_1056 N_A_1295_74#_c_1334_n N_A_2385_74#_c_1755_n 0.00505146f $X=12.23
+ $Y=1.885 $X2=0 $Y2=0
cc_1057 N_A_1295_74#_c_1360_n N_A_2385_74#_c_1755_n 0.0245872f $X=12.115 $Y=2.39
+ $X2=0 $Y2=0
cc_1058 N_A_1295_74#_c_1342_n N_A_2385_74#_c_1755_n 0.00549953f $X=12.3 $Y=1.59
+ $X2=0 $Y2=0
cc_1059 N_A_1295_74#_c_1334_n N_A_2385_74#_c_1756_n 0.0115967f $X=12.23 $Y=1.885
+ $X2=0 $Y2=0
cc_1060 N_A_1295_74#_c_1358_n N_A_2385_74#_c_1756_n 0.0142964f $X=12.03 $Y=2.475
+ $X2=0 $Y2=0
cc_1061 N_A_1295_74#_c_1360_n N_A_2385_74#_c_1756_n 0.0175574f $X=12.115 $Y=2.39
+ $X2=0 $Y2=0
cc_1062 N_A_1295_74#_c_1358_n N_VPWR_M1003_d 0.00663158f $X=12.03 $Y=2.475 $X2=0
+ $Y2=0
cc_1063 N_A_1295_74#_c_1358_n N_VPWR_M1009_s 0.011473f $X=12.03 $Y=2.475 $X2=0
+ $Y2=0
cc_1064 N_A_1295_74#_c_1344_n N_VPWR_c_2012_n 0.0107626f $X=7.9 $Y=1.765 $X2=0
+ $Y2=0
cc_1065 N_A_1295_74#_c_1348_n N_VPWR_c_2013_n 0.00126791f $X=9.375 $Y=2.465
+ $X2=0 $Y2=0
cc_1066 N_A_1295_74#_c_1358_n N_VPWR_c_2013_n 0.0212411f $X=12.03 $Y=2.475 $X2=0
+ $Y2=0
cc_1067 N_A_1295_74#_c_1358_n N_VPWR_c_2014_n 0.021438f $X=12.03 $Y=2.475 $X2=0
+ $Y2=0
cc_1068 N_A_1295_74#_c_1344_n N_VPWR_c_2024_n 0.00413917f $X=7.9 $Y=1.765 $X2=0
+ $Y2=0
cc_1069 N_A_1295_74#_c_1348_n N_VPWR_c_2024_n 0.00445602f $X=9.375 $Y=2.465
+ $X2=0 $Y2=0
cc_1070 N_A_1295_74#_c_1334_n N_VPWR_c_2030_n 0.00461464f $X=12.23 $Y=1.885
+ $X2=0 $Y2=0
cc_1071 N_A_1295_74#_c_1344_n N_VPWR_c_2007_n 0.00417047f $X=7.9 $Y=1.765 $X2=0
+ $Y2=0
cc_1072 N_A_1295_74#_c_1348_n N_VPWR_c_2007_n 0.0089489f $X=9.375 $Y=2.465 $X2=0
+ $Y2=0
cc_1073 N_A_1295_74#_c_1334_n N_VPWR_c_2007_n 0.00776565f $X=12.23 $Y=1.885
+ $X2=0 $Y2=0
cc_1074 N_A_1295_74#_c_1358_n N_VPWR_c_2007_n 0.0697413f $X=12.03 $Y=2.475 $X2=0
+ $Y2=0
cc_1075 N_A_1295_74#_c_1359_n N_VPWR_c_2007_n 0.00704359f $X=9.655 $Y=2.475
+ $X2=0 $Y2=0
cc_1076 N_A_1295_74#_c_1341_n N_A_669_111#_c_2169_n 0.0030604f $X=6.915 $Y=0.925
+ $X2=0 $Y2=0
cc_1077 N_A_1295_74#_c_1340_n N_A_669_111#_c_2170_n 0.00329338f $X=6.915 $Y=1.76
+ $X2=0 $Y2=0
cc_1078 N_A_1295_74#_c_1340_n N_A_669_111#_c_2172_n 0.00400982f $X=6.915 $Y=1.76
+ $X2=0 $Y2=0
cc_1079 N_A_1295_74#_c_1361_n N_A_669_111#_c_2172_n 0.0151305f $X=7 $Y=1.96
+ $X2=0 $Y2=0
cc_1080 N_A_1295_74#_M1020_d N_A_669_111#_c_2182_n 0.00751145f $X=6.625 $Y=1.78
+ $X2=0 $Y2=0
cc_1081 N_A_1295_74#_c_1330_n N_A_669_111#_c_2182_n 0.00350193f $X=7.825 $Y=1.69
+ $X2=0 $Y2=0
cc_1082 N_A_1295_74#_c_1355_n N_A_669_111#_c_2182_n 0.00832711f $X=7.225
+ $Y=1.995 $X2=0 $Y2=0
cc_1083 N_A_1295_74#_c_1361_n N_A_669_111#_c_2182_n 0.0541919f $X=7 $Y=1.96
+ $X2=0 $Y2=0
cc_1084 N_A_1295_74#_c_1330_n N_A_669_111#_c_2183_n 0.0092843f $X=7.825 $Y=1.69
+ $X2=0 $Y2=0
cc_1085 N_A_1295_74#_c_1344_n N_A_669_111#_c_2183_n 0.00638726f $X=7.9 $Y=1.765
+ $X2=0 $Y2=0
cc_1086 N_A_1295_74#_c_1340_n N_A_669_111#_c_2183_n 0.00177709f $X=6.915 $Y=1.76
+ $X2=0 $Y2=0
cc_1087 N_A_1295_74#_c_1354_n N_A_669_111#_c_2183_n 0.0204093f $X=7.225 $Y=1.995
+ $X2=0 $Y2=0
cc_1088 N_A_1295_74#_c_1355_n N_A_669_111#_c_2183_n 0.00195483f $X=7.225
+ $Y=1.995 $X2=0 $Y2=0
cc_1089 N_A_1295_74#_c_1361_n N_A_669_111#_c_2183_n 0.00220948f $X=7 $Y=1.96
+ $X2=0 $Y2=0
cc_1090 N_A_1295_74#_c_1330_n N_A_669_111#_c_2173_n 0.00146076f $X=7.825 $Y=1.69
+ $X2=0 $Y2=0
cc_1091 N_A_1295_74#_c_1331_n N_A_669_111#_c_2173_n 0.00790604f $X=8.29 $Y=1.69
+ $X2=0 $Y2=0
cc_1092 N_A_1295_74#_M1026_g N_A_669_111#_c_2173_n 0.00300237f $X=8.365 $Y=0.695
+ $X2=0 $Y2=0
cc_1093 N_A_1295_74#_c_1337_n N_A_669_111#_c_2173_n 0.00639244f $X=7.9 $Y=1.69
+ $X2=0 $Y2=0
cc_1094 N_A_1295_74#_M1007_g N_A_669_111#_c_2174_n 0.00341137f $X=7.385 $Y=0.74
+ $X2=0 $Y2=0
cc_1095 N_A_1295_74#_c_1330_n N_A_669_111#_c_2174_n 0.00413549f $X=7.825 $Y=1.69
+ $X2=0 $Y2=0
cc_1096 N_A_1295_74#_c_1340_n N_A_669_111#_c_2174_n 0.00465635f $X=6.915 $Y=1.76
+ $X2=0 $Y2=0
cc_1097 N_A_1295_74#_c_1344_n N_A_669_111#_c_2199_n 0.0162046f $X=7.9 $Y=1.765
+ $X2=0 $Y2=0
cc_1098 N_A_1295_74#_M1007_g N_A_669_111#_c_2175_n 0.00949229f $X=7.385 $Y=0.74
+ $X2=0 $Y2=0
cc_1099 N_A_1295_74#_M1026_g N_A_669_111#_c_2175_n 0.0127542f $X=8.365 $Y=0.695
+ $X2=0 $Y2=0
cc_1100 N_A_1295_74#_c_1344_n N_A_669_111#_c_2184_n 0.00497744f $X=7.9 $Y=1.765
+ $X2=0 $Y2=0
cc_1101 N_A_1295_74#_c_1358_n A_1890_508# 3.21084e-19 $X=12.03 $Y=2.475
+ $X2=-0.19 $Y2=-0.245
cc_1102 N_A_1295_74#_c_1359_n A_1890_508# 0.00328363f $X=9.655 $Y=2.475
+ $X2=-0.19 $Y2=-0.245
cc_1103 N_A_1295_74#_c_1358_n A_2274_392# 0.0321447f $X=12.03 $Y=2.475 $X2=-0.19
+ $Y2=-0.245
cc_1104 N_A_1295_74#_c_1360_n A_2274_392# 0.00754191f $X=12.115 $Y=2.39
+ $X2=-0.19 $Y2=-0.245
cc_1105 N_A_1295_74#_c_1339_n N_VGND_c_2390_n 0.0191484f $X=6.615 $Y=0.515 $X2=0
+ $Y2=0
cc_1106 N_A_1295_74#_M1007_g N_VGND_c_2391_n 0.00936698f $X=7.385 $Y=0.74 $X2=0
+ $Y2=0
cc_1107 N_A_1295_74#_c_1339_n N_VGND_c_2391_n 0.0219045f $X=6.615 $Y=0.515 $X2=0
+ $Y2=0
cc_1108 N_A_1295_74#_c_1339_n N_VGND_c_2400_n 0.0142249f $X=6.615 $Y=0.515 $X2=0
+ $Y2=0
cc_1109 N_A_1295_74#_M1007_g N_VGND_c_2404_n 0.00383152f $X=7.385 $Y=0.74 $X2=0
+ $Y2=0
cc_1110 N_A_1295_74#_M1026_g N_VGND_c_2404_n 7.53287e-19 $X=8.365 $Y=0.695 $X2=0
+ $Y2=0
cc_1111 N_A_1295_74#_M1034_g N_VGND_c_2411_n 0.00461464f $X=12.36 $Y=0.58 $X2=0
+ $Y2=0
cc_1112 N_A_1295_74#_M1034_g N_VGND_c_2412_n 0.00128745f $X=12.36 $Y=0.58 $X2=0
+ $Y2=0
cc_1113 N_A_1295_74#_M1007_g N_VGND_c_2413_n 0.00762539f $X=7.385 $Y=0.74 $X2=0
+ $Y2=0
cc_1114 N_A_1295_74#_M1034_g N_VGND_c_2413_n 0.00447595f $X=12.36 $Y=0.58 $X2=0
+ $Y2=0
cc_1115 N_A_1295_74#_c_1339_n N_VGND_c_2413_n 0.011867f $X=6.615 $Y=0.515 $X2=0
+ $Y2=0
cc_1116 N_A_1295_74#_c_1341_n N_VGND_c_2413_n 0.00766711f $X=6.915 $Y=0.925
+ $X2=0 $Y2=0
cc_1117 N_A_1910_71#_c_1530_n N_A_1688_97#_c_1642_n 0.0412719f $X=9.805 $Y=2.375
+ $X2=0 $Y2=0
cc_1118 N_A_1910_71#_c_1543_n N_A_1688_97#_c_1642_n 0.0101394f $X=9.805 $Y=2.465
+ $X2=0 $Y2=0
cc_1119 N_A_1910_71#_c_1533_n N_A_1688_97#_c_1642_n 0.00444722f $X=10.51 $Y=1.28
+ $X2=0 $Y2=0
cc_1120 N_A_1910_71#_c_1535_n N_A_1688_97#_c_1642_n 0.00805767f $X=10.72 $Y=1.97
+ $X2=0 $Y2=0
cc_1121 N_A_1910_71#_c_1536_n N_A_1688_97#_c_1642_n 6.95256e-19 $X=10.805
+ $Y=1.36 $X2=0 $Y2=0
cc_1122 N_A_1910_71#_c_1538_n N_A_1688_97#_c_1642_n 0.00125393f $X=11.22 $Y=1.36
+ $X2=0 $Y2=0
cc_1123 N_A_1910_71#_c_1547_n N_A_1688_97#_c_1642_n 0.00735278f $X=10.72
+ $Y=2.095 $X2=0 $Y2=0
cc_1124 N_A_1910_71#_M1029_g N_A_1688_97#_M1033_g 0.0117986f $X=9.625 $Y=0.695
+ $X2=0 $Y2=0
cc_1125 N_A_1910_71#_c_1533_n N_A_1688_97#_M1033_g 0.0143882f $X=10.51 $Y=1.28
+ $X2=0 $Y2=0
cc_1126 N_A_1910_71#_c_1534_n N_A_1688_97#_M1033_g 0.00617454f $X=10.595 $Y=0.81
+ $X2=0 $Y2=0
cc_1127 N_A_1910_71#_c_1536_n N_A_1688_97#_M1033_g 0.00364236f $X=10.805 $Y=1.36
+ $X2=0 $Y2=0
cc_1128 N_A_1910_71#_c_1538_n N_A_1688_97#_M1033_g 0.0182885f $X=11.22 $Y=1.36
+ $X2=0 $Y2=0
cc_1129 N_A_1910_71#_c_1539_n N_A_1688_97#_M1033_g 4.79872e-19 $X=9.895 $Y=1.32
+ $X2=0 $Y2=0
cc_1130 N_A_1910_71#_c_1540_n N_A_1688_97#_M1033_g 0.00990298f $X=9.805 $Y=1.32
+ $X2=0 $Y2=0
cc_1131 N_A_1910_71#_M1029_g N_A_1688_97#_c_1644_n 0.00248627f $X=9.625 $Y=0.695
+ $X2=0 $Y2=0
cc_1132 N_A_1910_71#_c_1539_n N_A_1688_97#_c_1644_n 0.0028446f $X=9.895 $Y=1.32
+ $X2=0 $Y2=0
cc_1133 N_A_1910_71#_c_1543_n N_A_1688_97#_c_1651_n 0.00165875f $X=9.805
+ $Y=2.465 $X2=0 $Y2=0
cc_1134 N_A_1910_71#_c_1530_n N_A_1688_97#_c_1645_n 6.52417e-19 $X=9.805
+ $Y=2.375 $X2=0 $Y2=0
cc_1135 N_A_1910_71#_c_1533_n N_A_1688_97#_c_1645_n 0.021831f $X=10.51 $Y=1.28
+ $X2=0 $Y2=0
cc_1136 N_A_1910_71#_c_1535_n N_A_1688_97#_c_1645_n 0.0187591f $X=10.72 $Y=1.97
+ $X2=0 $Y2=0
cc_1137 N_A_1910_71#_c_1547_n N_A_1688_97#_c_1645_n 0.00536709f $X=10.72
+ $Y=2.095 $X2=0 $Y2=0
cc_1138 N_A_1910_71#_c_1530_n N_A_1688_97#_c_1646_n 0.0133695f $X=9.805 $Y=2.375
+ $X2=0 $Y2=0
cc_1139 N_A_1910_71#_c_1533_n N_A_1688_97#_c_1646_n 0.0104157f $X=10.51 $Y=1.28
+ $X2=0 $Y2=0
cc_1140 N_A_1910_71#_c_1539_n N_A_1688_97#_c_1646_n 0.0207029f $X=9.895 $Y=1.32
+ $X2=0 $Y2=0
cc_1141 N_A_1910_71#_c_1540_n N_A_1688_97#_c_1646_n 0.00444912f $X=9.805 $Y=1.32
+ $X2=0 $Y2=0
cc_1142 N_A_1910_71#_c_1532_n N_A_2385_74#_c_1825_n 4.8666e-19 $X=11.49 $Y=1.11
+ $X2=0 $Y2=0
cc_1143 N_A_1910_71#_c_1532_n N_A_2385_74#_c_1746_n 0.001335f $X=11.49 $Y=1.11
+ $X2=0 $Y2=0
cc_1144 N_A_1910_71#_c_1543_n N_VPWR_c_2013_n 0.00932856f $X=9.805 $Y=2.465
+ $X2=0 $Y2=0
cc_1145 N_A_1910_71#_c_1545_n N_VPWR_c_2014_n 0.0183124f $X=11.295 $Y=1.885
+ $X2=0 $Y2=0
cc_1146 N_A_1910_71#_c_1543_n N_VPWR_c_2024_n 0.00413917f $X=9.805 $Y=2.465
+ $X2=0 $Y2=0
cc_1147 N_A_1910_71#_c_1545_n N_VPWR_c_2030_n 0.00413917f $X=11.295 $Y=1.885
+ $X2=0 $Y2=0
cc_1148 N_A_1910_71#_c_1543_n N_VPWR_c_2007_n 0.00398542f $X=9.805 $Y=2.465
+ $X2=0 $Y2=0
cc_1149 N_A_1910_71#_c_1545_n N_VPWR_c_2007_n 0.00403443f $X=11.295 $Y=1.885
+ $X2=0 $Y2=0
cc_1150 N_A_1910_71#_M1029_g N_VGND_c_2392_n 0.00360445f $X=9.625 $Y=0.695 $X2=0
+ $Y2=0
cc_1151 N_A_1910_71#_c_1532_n N_VGND_c_2393_n 0.0104726f $X=11.49 $Y=1.11 $X2=0
+ $Y2=0
cc_1152 N_A_1910_71#_M1029_g N_VGND_c_2404_n 0.00497279f $X=9.625 $Y=0.695 $X2=0
+ $Y2=0
cc_1153 N_A_1910_71#_c_1532_n N_VGND_c_2411_n 0.00383152f $X=11.49 $Y=1.11 $X2=0
+ $Y2=0
cc_1154 N_A_1910_71#_M1029_g N_VGND_c_2413_n 0.00509887f $X=9.625 $Y=0.695 $X2=0
+ $Y2=0
cc_1155 N_A_1910_71#_c_1532_n N_VGND_c_2413_n 0.00386494f $X=11.49 $Y=1.11 $X2=0
+ $Y2=0
cc_1156 N_A_1688_97#_c_1642_n N_VPWR_c_2013_n 0.00418529f $X=10.325 $Y=1.915
+ $X2=0 $Y2=0
cc_1157 N_A_1688_97#_c_1648_n N_VPWR_c_2013_n 0.00715172f $X=9.15 $Y=2.75 $X2=0
+ $Y2=0
cc_1158 N_A_1688_97#_c_1642_n N_VPWR_c_2014_n 0.00600586f $X=10.325 $Y=1.915
+ $X2=0 $Y2=0
cc_1159 N_A_1688_97#_c_1648_n N_VPWR_c_2024_n 0.014453f $X=9.15 $Y=2.75 $X2=0
+ $Y2=0
cc_1160 N_A_1688_97#_c_1642_n N_VPWR_c_2026_n 0.00487664f $X=10.325 $Y=1.915
+ $X2=0 $Y2=0
cc_1161 N_A_1688_97#_c_1642_n N_VPWR_c_2007_n 0.00505379f $X=10.325 $Y=1.915
+ $X2=0 $Y2=0
cc_1162 N_A_1688_97#_c_1648_n N_VPWR_c_2007_n 0.011992f $X=9.15 $Y=2.75 $X2=0
+ $Y2=0
cc_1163 N_A_1688_97#_c_1651_n N_VPWR_c_2007_n 0.00536095f $X=9.075 $Y=2.56 $X2=0
+ $Y2=0
cc_1164 N_A_1688_97#_c_1650_n N_A_669_111#_c_2199_n 0.0046794f $X=9.075 $Y=2.39
+ $X2=0 $Y2=0
cc_1165 N_A_1688_97#_c_1651_n N_A_669_111#_c_2282_n 0.00155083f $X=9.075 $Y=2.56
+ $X2=0 $Y2=0
cc_1166 N_A_1688_97#_c_1648_n N_A_669_111#_c_2185_n 0.0111988f $X=9.15 $Y=2.75
+ $X2=0 $Y2=0
cc_1167 N_A_1688_97#_M1033_g N_VGND_c_2392_n 0.00193096f $X=10.38 $Y=0.69 $X2=0
+ $Y2=0
cc_1168 N_A_1688_97#_M1033_g N_VGND_c_2405_n 0.00278237f $X=10.38 $Y=0.69 $X2=0
+ $Y2=0
cc_1169 N_A_1688_97#_M1033_g N_VGND_c_2413_n 0.00363424f $X=10.38 $Y=0.69 $X2=0
+ $Y2=0
cc_1170 N_A_2385_74#_c_1752_n N_VPWR_c_2015_n 0.00623607f $X=13.895 $Y=2.245
+ $X2=0 $Y2=0
cc_1171 N_A_2385_74#_c_1756_n N_VPWR_c_2015_n 0.0111431f $X=12.455 $Y=2.815
+ $X2=0 $Y2=0
cc_1172 N_A_2385_74#_c_1753_n N_VPWR_c_2017_n 0.00990979f $X=14.865 $Y=1.765
+ $X2=0 $Y2=0
cc_1173 N_A_2385_74#_c_1756_n N_VPWR_c_2030_n 0.0189801f $X=12.455 $Y=2.815
+ $X2=0 $Y2=0
cc_1174 N_A_2385_74#_c_1752_n N_VPWR_c_2031_n 0.00445602f $X=13.895 $Y=2.245
+ $X2=0 $Y2=0
cc_1175 N_A_2385_74#_c_1753_n N_VPWR_c_2031_n 0.00434272f $X=14.865 $Y=1.765
+ $X2=0 $Y2=0
cc_1176 N_A_2385_74#_c_1752_n N_VPWR_c_2007_n 0.00863669f $X=13.895 $Y=2.245
+ $X2=0 $Y2=0
cc_1177 N_A_2385_74#_c_1753_n N_VPWR_c_2007_n 0.00829165f $X=14.865 $Y=1.765
+ $X2=0 $Y2=0
cc_1178 N_A_2385_74#_c_1756_n N_VPWR_c_2007_n 0.0154423f $X=12.455 $Y=2.815
+ $X2=0 $Y2=0
cc_1179 N_A_2385_74#_M1019_g Q 8.40247e-19 $X=13.875 $Y=0.58 $X2=0 $Y2=0
cc_1180 N_A_2385_74#_c_1741_n Q 6.6515e-19 $X=13.895 $Y=2.155 $X2=0 $Y2=0
cc_1181 N_A_2385_74#_c_1752_n Q 0.00134701f $X=13.895 $Y=2.245 $X2=0 $Y2=0
cc_1182 N_A_2385_74#_c_1742_n Q 0.0314646f $X=14.775 $Y=1.425 $X2=0 $Y2=0
cc_1183 N_A_2385_74#_c_1744_n Q 0.0170778f $X=14.865 $Y=1.23 $X2=0 $Y2=0
cc_1184 N_A_2385_74#_c_1753_n Q 0.0184448f $X=14.865 $Y=1.765 $X2=0 $Y2=0
cc_1185 N_A_2385_74#_c_1745_n Q 0.0278379f $X=14.865 $Y=1.497 $X2=0 $Y2=0
cc_1186 N_A_2385_74#_c_1747_n N_VGND_M1035_d 0.00523342f $X=13.175 $Y=0.855
+ $X2=0 $Y2=0
cc_1187 N_A_2385_74#_c_1746_n N_VGND_c_2393_n 0.0109748f $X=12.065 $Y=0.515
+ $X2=0 $Y2=0
cc_1188 N_A_2385_74#_c_1744_n N_VGND_c_2395_n 0.00647412f $X=14.865 $Y=1.23
+ $X2=0 $Y2=0
cc_1189 N_A_2385_74#_M1019_g N_VGND_c_2406_n 0.00434272f $X=13.875 $Y=0.58 $X2=0
+ $Y2=0
cc_1190 N_A_2385_74#_c_1744_n N_VGND_c_2406_n 0.00434272f $X=14.865 $Y=1.23
+ $X2=0 $Y2=0
cc_1191 N_A_2385_74#_c_1746_n N_VGND_c_2411_n 0.014415f $X=12.065 $Y=0.515 $X2=0
+ $Y2=0
cc_1192 N_A_2385_74#_M1019_g N_VGND_c_2412_n 0.010036f $X=13.875 $Y=0.58 $X2=0
+ $Y2=0
cc_1193 N_A_2385_74#_c_1743_n N_VGND_c_2412_n 8.9533e-19 $X=13.985 $Y=1.425
+ $X2=0 $Y2=0
cc_1194 N_A_2385_74#_c_1746_n N_VGND_c_2412_n 0.00419512f $X=12.065 $Y=0.515
+ $X2=0 $Y2=0
cc_1195 N_A_2385_74#_c_1747_n N_VGND_c_2412_n 0.0395975f $X=13.175 $Y=0.855
+ $X2=0 $Y2=0
cc_1196 N_A_2385_74#_c_1750_n N_VGND_c_2412_n 0.00542593f $X=13.78 $Y=1.215
+ $X2=0 $Y2=0
cc_1197 N_A_2385_74#_M1019_g N_VGND_c_2413_n 0.00830035f $X=13.875 $Y=0.58 $X2=0
+ $Y2=0
cc_1198 N_A_2385_74#_c_1744_n N_VGND_c_2413_n 0.00828941f $X=14.865 $Y=1.23
+ $X2=0 $Y2=0
cc_1199 N_A_2385_74#_c_1746_n N_VGND_c_2413_n 0.0119404f $X=12.065 $Y=0.515
+ $X2=0 $Y2=0
cc_1200 N_A_2385_74#_c_1747_n N_VGND_c_2413_n 0.0209571f $X=13.175 $Y=0.855
+ $X2=0 $Y2=0
cc_1201 N_A_2385_74#_c_1747_n A_2487_74# 0.0023798f $X=13.175 $Y=0.855 $X2=-0.19
+ $Y2=-0.245
cc_1202 N_A_27_74#_c_1891_n A_114_464# 0.0048076f $X=1.365 $Y=2.375 $X2=-0.19
+ $Y2=-0.245
cc_1203 N_A_27_74#_c_1891_n N_VPWR_M1023_d 0.00509381f $X=1.365 $Y=2.375
+ $X2=-0.19 $Y2=-0.245
cc_1204 N_A_27_74#_c_1893_n N_VPWR_M1036_d 4.76982e-19 $X=2.045 $Y=2.99 $X2=0
+ $Y2=0
cc_1205 N_A_27_74#_c_1925_n N_VPWR_M1036_d 0.00490162f $X=2.13 $Y=2.905 $X2=0
+ $Y2=0
cc_1206 N_A_27_74#_c_1895_n N_VPWR_M1036_d 0.00972296f $X=3.145 $Y=2.375 $X2=0
+ $Y2=0
cc_1207 N_A_27_74#_c_1890_n N_VPWR_c_2008_n 0.0105321f $X=0.27 $Y=2.465 $X2=0
+ $Y2=0
cc_1208 N_A_27_74#_c_1891_n N_VPWR_c_2008_n 0.0154248f $X=1.365 $Y=2.375 $X2=0
+ $Y2=0
cc_1209 N_A_27_74#_c_1892_n N_VPWR_c_2008_n 0.0208967f $X=1.45 $Y=2.905 $X2=0
+ $Y2=0
cc_1210 N_A_27_74#_c_1894_n N_VPWR_c_2008_n 0.0146662f $X=1.535 $Y=2.99 $X2=0
+ $Y2=0
cc_1211 N_A_27_74#_c_1893_n N_VPWR_c_2009_n 0.0145842f $X=2.045 $Y=2.99 $X2=0
+ $Y2=0
cc_1212 N_A_27_74#_c_1925_n N_VPWR_c_2009_n 0.0205316f $X=2.13 $Y=2.905 $X2=0
+ $Y2=0
cc_1213 N_A_27_74#_c_1895_n N_VPWR_c_2009_n 0.0154248f $X=3.145 $Y=2.375 $X2=0
+ $Y2=0
cc_1214 N_A_27_74#_c_1897_n N_VPWR_c_2009_n 0.0101141f $X=3.31 $Y=2.46 $X2=0
+ $Y2=0
cc_1215 N_A_27_74#_c_1890_n N_VPWR_c_2018_n 0.0154947f $X=0.27 $Y=2.465 $X2=0
+ $Y2=0
cc_1216 N_A_27_74#_c_1893_n N_VPWR_c_2020_n 0.0445209f $X=2.045 $Y=2.99 $X2=0
+ $Y2=0
cc_1217 N_A_27_74#_c_1894_n N_VPWR_c_2020_n 0.0121867f $X=1.535 $Y=2.99 $X2=0
+ $Y2=0
cc_1218 N_A_27_74#_c_1897_n N_VPWR_c_2028_n 0.0108086f $X=3.31 $Y=2.46 $X2=0
+ $Y2=0
cc_1219 N_A_27_74#_c_1890_n N_VPWR_c_2007_n 0.0127886f $X=0.27 $Y=2.465 $X2=0
+ $Y2=0
cc_1220 N_A_27_74#_c_1893_n N_VPWR_c_2007_n 0.0250929f $X=2.045 $Y=2.99 $X2=0
+ $Y2=0
cc_1221 N_A_27_74#_c_1894_n N_VPWR_c_2007_n 0.00660921f $X=1.535 $Y=2.99 $X2=0
+ $Y2=0
cc_1222 N_A_27_74#_c_1897_n N_VPWR_c_2007_n 0.00906495f $X=3.31 $Y=2.46 $X2=0
+ $Y2=0
cc_1223 N_A_27_74#_c_1895_n A_554_463# 0.0048076f $X=3.145 $Y=2.375 $X2=-0.19
+ $Y2=-0.245
cc_1224 N_A_27_74#_c_1897_n N_A_669_111#_c_2249_n 0.033328f $X=3.31 $Y=2.46
+ $X2=0 $Y2=0
cc_1225 N_A_27_74#_c_1897_n N_A_669_111#_c_2191_n 0.00568204f $X=3.31 $Y=2.46
+ $X2=0 $Y2=0
cc_1226 N_A_27_74#_c_1885_n N_A_669_111#_c_2176_n 0.018852f $X=3.055 $Y=0.765
+ $X2=0 $Y2=0
cc_1227 N_A_27_74#_c_1885_n N_A_669_111#_c_2177_n 0.0070485f $X=3.055 $Y=0.765
+ $X2=0 $Y2=0
cc_1228 N_A_27_74#_c_1886_n N_A_669_111#_c_2177_n 0.0708093f $X=3.31 $Y=2.29
+ $X2=0 $Y2=0
cc_1229 N_A_27_74#_c_1888_n N_A_669_111#_c_2177_n 0.0135705f $X=3.31 $Y=1.25
+ $X2=0 $Y2=0
cc_1230 N_A_27_74#_c_1900_n N_A_669_111#_c_2177_n 0.0138383f $X=3.27 $Y=2.375
+ $X2=0 $Y2=0
cc_1231 N_A_27_74#_c_1887_n N_VGND_c_2387_n 0.010763f $X=0.35 $Y=0.645 $X2=0
+ $Y2=0
cc_1232 N_A_27_74#_c_1885_n N_VGND_c_2388_n 0.0145731f $X=3.055 $Y=0.765 $X2=0
+ $Y2=0
cc_1233 N_A_27_74#_c_1885_n N_VGND_c_2396_n 0.00814422f $X=3.055 $Y=0.765 $X2=0
+ $Y2=0
cc_1234 N_A_27_74#_c_1887_n N_VGND_c_2402_n 0.0128299f $X=0.35 $Y=0.645 $X2=0
+ $Y2=0
cc_1235 N_A_27_74#_c_1885_n N_VGND_c_2413_n 0.0106161f $X=3.055 $Y=0.765 $X2=0
+ $Y2=0
cc_1236 N_A_27_74#_c_1887_n N_VGND_c_2413_n 0.0165133f $X=0.35 $Y=0.645 $X2=0
+ $Y2=0
cc_1237 N_VPWR_c_2010_n N_A_669_111#_c_2179_n 0.0147124f $X=4.965 $Y=2.765 $X2=0
+ $Y2=0
cc_1238 N_VPWR_c_2028_n N_A_669_111#_c_2179_n 0.0546448f $X=4.88 $Y=3.33 $X2=0
+ $Y2=0
cc_1239 N_VPWR_c_2007_n N_A_669_111#_c_2179_n 0.0292625f $X=15.12 $Y=3.33 $X2=0
+ $Y2=0
cc_1240 N_VPWR_c_2028_n N_A_669_111#_c_2191_n 0.0190556f $X=4.88 $Y=3.33 $X2=0
+ $Y2=0
cc_1241 N_VPWR_c_2007_n N_A_669_111#_c_2191_n 0.00957028f $X=15.12 $Y=3.33 $X2=0
+ $Y2=0
cc_1242 N_VPWR_M1027_d N_A_669_111#_c_2209_n 0.00522241f $X=4.585 $Y=2.275 $X2=0
+ $Y2=0
cc_1243 N_VPWR_c_2010_n N_A_669_111#_c_2209_n 0.0231493f $X=4.965 $Y=2.765 $X2=0
+ $Y2=0
cc_1244 N_VPWR_M1020_s N_A_669_111#_c_2182_n 0.00755048f $X=6.2 $Y=1.78 $X2=0
+ $Y2=0
cc_1245 N_VPWR_M1030_s N_A_669_111#_c_2182_n 0.00194795f $X=7.55 $Y=1.84 $X2=0
+ $Y2=0
cc_1246 N_VPWR_c_2011_n N_A_669_111#_c_2182_n 0.0215517f $X=6.325 $Y=2.755 $X2=0
+ $Y2=0
cc_1247 N_VPWR_c_2012_n N_A_669_111#_c_2182_n 0.00874994f $X=7.675 $Y=2.785
+ $X2=0 $Y2=0
cc_1248 N_VPWR_c_2007_n N_A_669_111#_c_2182_n 0.0365828f $X=15.12 $Y=3.33 $X2=0
+ $Y2=0
cc_1249 N_VPWR_M1030_s N_A_669_111#_c_2183_n 0.0114686f $X=7.55 $Y=1.84 $X2=0
+ $Y2=0
cc_1250 N_VPWR_c_2012_n N_A_669_111#_c_2199_n 0.00100013f $X=7.675 $Y=2.785
+ $X2=0 $Y2=0
cc_1251 N_VPWR_c_2007_n N_A_669_111#_c_2199_n 0.00512221f $X=15.12 $Y=3.33 $X2=0
+ $Y2=0
cc_1252 N_VPWR_c_2012_n N_A_669_111#_c_2184_n 0.0103109f $X=7.675 $Y=2.785 $X2=0
+ $Y2=0
cc_1253 N_VPWR_c_2024_n N_A_669_111#_c_2184_n 0.00756061f $X=9.865 $Y=3.33 $X2=0
+ $Y2=0
cc_1254 N_VPWR_c_2007_n N_A_669_111#_c_2184_n 0.00626901f $X=15.12 $Y=3.33 $X2=0
+ $Y2=0
cc_1255 N_VPWR_c_2024_n N_A_669_111#_c_2185_n 0.0262326f $X=9.865 $Y=3.33 $X2=0
+ $Y2=0
cc_1256 N_VPWR_c_2007_n N_A_669_111#_c_2185_n 0.0226252f $X=15.12 $Y=3.33 $X2=0
+ $Y2=0
cc_1257 N_VPWR_c_2010_n N_A_669_111#_c_2187_n 0.0102312f $X=4.965 $Y=2.765 $X2=0
+ $Y2=0
cc_1258 N_VPWR_c_2011_n N_A_669_111#_c_2187_n 0.0221648f $X=6.325 $Y=2.755 $X2=0
+ $Y2=0
cc_1259 N_VPWR_c_2029_n N_A_669_111#_c_2187_n 0.0126964f $X=6.16 $Y=3.33 $X2=0
+ $Y2=0
cc_1260 N_VPWR_c_2007_n N_A_669_111#_c_2187_n 0.0122875f $X=15.12 $Y=3.33 $X2=0
+ $Y2=0
cc_1261 N_VPWR_M1027_d N_A_669_111#_c_2188_n 0.00977001f $X=4.585 $Y=2.275 $X2=0
+ $Y2=0
cc_1262 N_VPWR_c_2010_n N_A_669_111#_c_2188_n 0.0154248f $X=4.965 $Y=2.765 $X2=0
+ $Y2=0
cc_1263 N_VPWR_c_2007_n N_A_669_111#_c_2189_n 0.00619814f $X=15.12 $Y=3.33 $X2=0
+ $Y2=0
cc_1264 N_VPWR_M1030_s N_A_669_111#_c_2351_n 0.00183865f $X=7.55 $Y=1.84 $X2=0
+ $Y2=0
cc_1265 N_VPWR_c_2012_n N_A_669_111#_c_2351_n 0.012967f $X=7.675 $Y=2.785 $X2=0
+ $Y2=0
cc_1266 N_VPWR_c_2007_n N_A_669_111#_c_2351_n 6.24256e-19 $X=15.12 $Y=3.33 $X2=0
+ $Y2=0
cc_1267 N_VPWR_c_2017_n Q 0.0811475f $X=15.09 $Y=1.985 $X2=0 $Y2=0
cc_1268 N_VPWR_c_2031_n Q 0.0150101f $X=15.005 $Y=3.33 $X2=0 $Y2=0
cc_1269 N_VPWR_c_2007_n Q 0.0123677f $X=15.12 $Y=3.33 $X2=0 $Y2=0
cc_1270 N_A_669_111#_c_2188_n A_1053_455# 0.0048076f $X=5.64 $Y=2.377 $X2=-0.19
+ $Y2=-0.245
cc_1271 N_A_669_111#_c_2170_n N_VGND_M1018_s 0.00208524f $X=5.99 $Y=1.16 $X2=0
+ $Y2=0
cc_1272 N_A_669_111#_c_2169_n N_VGND_c_2389_n 0.013268f $X=5.63 $Y=0.835 $X2=0
+ $Y2=0
cc_1273 N_A_669_111#_c_2169_n N_VGND_c_2390_n 0.0201715f $X=5.63 $Y=0.835 $X2=0
+ $Y2=0
cc_1274 N_A_669_111#_c_2170_n N_VGND_c_2390_n 0.0125997f $X=5.99 $Y=1.16 $X2=0
+ $Y2=0
cc_1275 N_A_669_111#_c_2176_n N_VGND_c_2396_n 0.00856317f $X=3.555 $Y=0.765
+ $X2=0 $Y2=0
cc_1276 N_A_669_111#_c_2169_n N_VGND_c_2398_n 0.00698925f $X=5.63 $Y=0.835 $X2=0
+ $Y2=0
cc_1277 N_A_669_111#_c_2169_n N_VGND_c_2413_n 0.0100239f $X=5.63 $Y=0.835 $X2=0
+ $Y2=0
cc_1278 N_A_669_111#_c_2176_n N_VGND_c_2413_n 0.0111006f $X=3.555 $Y=0.765 $X2=0
+ $Y2=0
cc_1279 Q N_VGND_c_2395_n 0.0295402f $X=14.555 $Y=0.47 $X2=0 $Y2=0
cc_1280 Q N_VGND_c_2406_n 0.0150101f $X=14.555 $Y=0.47 $X2=0 $Y2=0
cc_1281 Q N_VGND_c_2413_n 0.0123677f $X=14.555 $Y=0.47 $X2=0 $Y2=0
