* File: sky130_fd_sc_hs__o311ai_2.pex.spice
* Created: Thu Aug 27 21:02:12 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HS__O311AI_2%A1 3 5 7 8 10 13 15 16 24
c42 8 0 3.17312e-19 $X=0.97 $Y=1.765
r43 24 25 1.91777 $w=3.77e-07 $l=1.5e-08 $layer=POLY_cond $X=0.97 $Y=1.557
+ $X2=0.985 $Y2=1.557
r44 22 24 49.2228 $w=3.77e-07 $l=3.85e-07 $layer=POLY_cond $X=0.585 $Y=1.557
+ $X2=0.97 $Y2=1.557
r45 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.585
+ $Y=1.515 $X2=0.585 $Y2=1.515
r46 20 22 9.58886 $w=3.77e-07 $l=7.5e-08 $layer=POLY_cond $X=0.51 $Y=1.557
+ $X2=0.585 $Y2=1.557
r47 19 20 1.91777 $w=3.77e-07 $l=1.5e-08 $layer=POLY_cond $X=0.495 $Y=1.557
+ $X2=0.51 $Y2=1.557
r48 16 23 3.61813 $w=4.28e-07 $l=1.35e-07 $layer=LI1_cond $X=0.72 $Y=1.565
+ $X2=0.585 $Y2=1.565
r49 15 23 9.24634 $w=4.28e-07 $l=3.45e-07 $layer=LI1_cond $X=0.24 $Y=1.565
+ $X2=0.585 $Y2=1.565
r50 11 25 24.4204 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.985 $Y=1.35
+ $X2=0.985 $Y2=1.557
r51 11 13 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=0.985 $Y=1.35
+ $X2=0.985 $Y2=0.74
r52 8 24 24.4204 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=0.97 $Y=1.765
+ $X2=0.97 $Y2=1.557
r53 8 10 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.97 $Y=1.765
+ $X2=0.97 $Y2=2.4
r54 5 20 24.4204 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=0.51 $Y=1.765
+ $X2=0.51 $Y2=1.557
r55 5 7 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.51 $Y=1.765
+ $X2=0.51 $Y2=2.4
r56 1 19 24.4204 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.495 $Y=1.35
+ $X2=0.495 $Y2=1.557
r57 1 3 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=0.495 $Y=1.35
+ $X2=0.495 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HS__O311AI_2%A2 1 3 6 10 12 14 15 16 17 26
c54 17 0 1.96049e-19 $X=2.16 $Y=1.665
c55 12 0 6.66869e-20 $X=1.98 $Y=1.765
r56 26 27 8.58356 $w=3.65e-07 $l=6.5e-08 $layer=POLY_cond $X=1.915 $Y=1.557
+ $X2=1.98 $Y2=1.557
r57 24 26 1.32055 $w=3.65e-07 $l=1e-08 $layer=POLY_cond $X=1.905 $Y=1.557
+ $X2=1.915 $Y2=1.557
r58 24 25 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.905
+ $Y=1.515 $X2=1.905 $Y2=1.515
r59 22 24 56.7836 $w=3.65e-07 $l=4.3e-07 $layer=POLY_cond $X=1.475 $Y=1.557
+ $X2=1.905 $Y2=1.557
r60 21 22 1.98082 $w=3.65e-07 $l=1.5e-08 $layer=POLY_cond $X=1.46 $Y=1.557
+ $X2=1.475 $Y2=1.557
r61 17 25 6.83426 $w=4.28e-07 $l=2.55e-07 $layer=LI1_cond $X=2.16 $Y=1.565
+ $X2=1.905 $Y2=1.565
r62 16 25 6.03022 $w=4.28e-07 $l=2.25e-07 $layer=LI1_cond $X=1.68 $Y=1.565
+ $X2=1.905 $Y2=1.565
r63 15 16 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=1.2 $Y=1.565
+ $X2=1.68 $Y2=1.565
r64 12 27 23.6381 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=1.98 $Y=1.765
+ $X2=1.98 $Y2=1.557
r65 12 14 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.98 $Y=1.765
+ $X2=1.98 $Y2=2.4
r66 8 26 23.6381 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.915 $Y=1.35
+ $X2=1.915 $Y2=1.557
r67 8 10 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.915 $Y=1.35
+ $X2=1.915 $Y2=0.74
r68 4 22 23.6381 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.475 $Y=1.35
+ $X2=1.475 $Y2=1.557
r69 4 6 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.475 $Y=1.35
+ $X2=1.475 $Y2=0.74
r70 1 21 23.6381 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=1.46 $Y=1.765
+ $X2=1.46 $Y2=1.557
r71 1 3 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.46 $Y=1.765
+ $X2=1.46 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_HS__O311AI_2%A3 3 7 9 11 12 13 14 16 17 18
c62 18 0 1.50622e-19 $X=3.12 $Y=1.665
c63 12 0 1.72564e-20 $X=3.35 $Y=1.65
c64 9 0 6.12971e-20 $X=2.99 $Y=1.765
r65 23 25 22.1691 $w=3.37e-07 $l=1.55e-07 $layer=POLY_cond $X=2.69 $Y=1.557
+ $X2=2.845 $Y2=1.557
r66 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.69
+ $Y=1.515 $X2=2.69 $Y2=1.515
r67 21 23 43.6231 $w=3.37e-07 $l=3.05e-07 $layer=POLY_cond $X=2.385 $Y=1.557
+ $X2=2.69 $Y2=1.557
r68 18 24 11.5244 $w=4.28e-07 $l=4.3e-07 $layer=LI1_cond $X=3.12 $Y=1.565
+ $X2=2.69 $Y2=1.565
r69 17 24 1.34005 $w=4.28e-07 $l=5e-08 $layer=LI1_cond $X=2.64 $Y=1.565 $X2=2.69
+ $Y2=1.565
r70 14 16 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.44 $Y=1.765
+ $X2=3.44 $Y2=2.4
r71 12 14 26.9307 $w=1.5e-07 $l=1.53542e-07 $layer=POLY_cond $X=3.35 $Y=1.65
+ $X2=3.44 $Y2=1.765
r72 12 13 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=3.35 $Y=1.65
+ $X2=3.08 $Y2=1.65
r73 9 13 27.9259 $w=3.37e-07 $l=1.53542e-07 $layer=POLY_cond $X=2.99 $Y=1.765
+ $X2=3.08 $Y2=1.65
r74 9 25 20.7389 $w=3.37e-07 $l=2.70969e-07 $layer=POLY_cond $X=2.99 $Y=1.765
+ $X2=2.845 $Y2=1.557
r75 9 11 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.99 $Y=1.765
+ $X2=2.99 $Y2=2.4
r76 5 25 21.7231 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.845 $Y=1.35
+ $X2=2.845 $Y2=1.557
r77 5 7 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.845 $Y=1.35
+ $X2=2.845 $Y2=0.74
r78 1 21 21.7231 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.385 $Y=1.35
+ $X2=2.385 $Y2=1.557
r79 1 3 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.385 $Y=1.35
+ $X2=2.385 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HS__O311AI_2%B1 1 3 4 5 6 8 9 11 12 14 16 19 21 22 26
c70 22 0 1.09862e-20 $X=4.08 $Y=1.665
c71 19 0 1.4261e-19 $X=3.935 $Y=1.53
r72 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.935
+ $Y=1.515 $X2=3.935 $Y2=1.515
r73 22 27 3.88615 $w=4.28e-07 $l=1.45e-07 $layer=LI1_cond $X=4.08 $Y=1.565
+ $X2=3.935 $Y2=1.565
r74 21 27 8.97834 $w=4.28e-07 $l=3.35e-07 $layer=LI1_cond $X=3.6 $Y=1.565
+ $X2=3.935 $Y2=1.565
r75 19 26 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=3.935 $Y=1.53
+ $X2=3.935 $Y2=1.515
r76 19 20 99.5969 $w=1.96e-07 $l=4.05e-07 $layer=POLY_cond $X=3.935 $Y=1.647
+ $X2=4.34 $Y2=1.647
r77 17 19 11.0663 $w=1.96e-07 $l=4.5e-08 $layer=POLY_cond $X=3.89 $Y=1.647
+ $X2=3.935 $Y2=1.647
r78 15 26 31.475 $w=3.3e-07 $l=1.8e-07 $layer=POLY_cond $X=3.935 $Y=1.335
+ $X2=3.935 $Y2=1.515
r79 15 16 13.5877 $w=2.4e-07 $l=7.5e-08 $layer=POLY_cond $X=3.935 $Y=1.335
+ $X2=3.935 $Y2=1.26
r80 12 20 9.11062 $w=1.5e-07 $l=1.18e-07 $layer=POLY_cond $X=4.34 $Y=1.765
+ $X2=4.34 $Y2=1.647
r81 12 14 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=4.34 $Y=1.765
+ $X2=4.34 $Y2=2.4
r82 9 17 9.11062 $w=1.5e-07 $l=1.18e-07 $layer=POLY_cond $X=3.89 $Y=1.765
+ $X2=3.89 $Y2=1.647
r83 9 11 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.89 $Y=1.765
+ $X2=3.89 $Y2=2.4
r84 6 16 13.5877 $w=2.4e-07 $l=1.21861e-07 $layer=POLY_cond $X=3.845 $Y=1.185
+ $X2=3.935 $Y2=1.26
r85 6 8 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=3.845 $Y=1.185
+ $X2=3.845 $Y2=0.74
r86 4 16 12.1617 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.77 $Y=1.26
+ $X2=3.935 $Y2=1.26
r87 4 5 215.362 $w=1.5e-07 $l=4.2e-07 $layer=POLY_cond $X=3.77 $Y=1.26 $X2=3.35
+ $Y2=1.26
r88 1 5 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.275 $Y=1.185
+ $X2=3.35 $Y2=1.26
r89 1 3 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=3.275 $Y=1.185
+ $X2=3.275 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HS__O311AI_2%C1 1 3 6 8 10 13 15 16 22
c50 16 0 5.86747e-20 $X=5.52 $Y=1.665
r51 24 25 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.43
+ $Y=1.465 $X2=5.43 $Y2=1.465
r52 22 24 20.7109 $w=3.84e-07 $l=1.65e-07 $layer=POLY_cond $X=5.265 $Y=1.532
+ $X2=5.43 $Y2=1.532
r53 21 22 3.13802 $w=3.84e-07 $l=2.5e-08 $layer=POLY_cond $X=5.24 $Y=1.532
+ $X2=5.265 $Y2=1.532
r54 20 21 50.8359 $w=3.84e-07 $l=4.05e-07 $layer=POLY_cond $X=4.835 $Y=1.532
+ $X2=5.24 $Y2=1.532
r55 19 20 5.64844 $w=3.84e-07 $l=4.5e-08 $layer=POLY_cond $X=4.79 $Y=1.532
+ $X2=4.835 $Y2=1.532
r56 16 25 2.24265 $w=4.78e-07 $l=9e-08 $layer=LI1_cond $X=5.52 $Y=1.54 $X2=5.43
+ $Y2=1.54
r57 15 25 9.71814 $w=4.78e-07 $l=3.9e-07 $layer=LI1_cond $X=5.04 $Y=1.54
+ $X2=5.43 $Y2=1.54
r58 11 22 24.8669 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=5.265 $Y=1.3
+ $X2=5.265 $Y2=1.532
r59 11 13 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=5.265 $Y=1.3
+ $X2=5.265 $Y2=0.74
r60 8 21 24.8669 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=5.24 $Y=1.765
+ $X2=5.24 $Y2=1.532
r61 8 10 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=5.24 $Y=1.765
+ $X2=5.24 $Y2=2.4
r62 4 20 24.8669 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=4.835 $Y=1.3
+ $X2=4.835 $Y2=1.532
r63 4 6 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=4.835 $Y=1.3 $X2=4.835
+ $Y2=0.74
r64 1 19 24.8669 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=4.79 $Y=1.765
+ $X2=4.79 $Y2=1.532
r65 1 3 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=4.79 $Y=1.765
+ $X2=4.79 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_HS__O311AI_2%A_28_368# 1 2 3 10 12 14 18 20 27 29
c39 18 0 1.71574e-19 $X=1.235 $Y=2.815
r40 21 27 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.4 $Y=2.035
+ $X2=1.235 $Y2=2.035
r41 20 29 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.12 $Y=2.035
+ $X2=2.245 $Y2=2.035
r42 20 21 46.9733 $w=1.68e-07 $l=7.2e-07 $layer=LI1_cond $X=2.12 $Y=2.035
+ $X2=1.4 $Y2=2.035
r43 16 27 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.235 $Y=2.12
+ $X2=1.235 $Y2=2.035
r44 16 18 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=1.235 $Y=2.12
+ $X2=1.235 $Y2=2.815
r45 15 25 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.45 $Y=2.035
+ $X2=0.285 $Y2=2.035
r46 14 27 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.07 $Y=2.035
+ $X2=1.235 $Y2=2.035
r47 14 15 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=1.07 $Y=2.035
+ $X2=0.45 $Y2=2.035
r48 10 25 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.285 $Y=2.12
+ $X2=0.285 $Y2=2.035
r49 10 12 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=0.285 $Y=2.12
+ $X2=0.285 $Y2=2.815
r50 3 29 300 $w=1.7e-07 $l=3.4187e-07 $layer=licon1_PDIFF $count=2 $X=2.055
+ $Y=1.84 $X2=2.205 $Y2=2.115
r51 2 27 400 $w=1.7e-07 $l=3.57596e-07 $layer=licon1_PDIFF $count=1 $X=1.045
+ $Y=1.84 $X2=1.235 $Y2=2.115
r52 2 18 400 $w=1.7e-07 $l=1.06577e-06 $layer=licon1_PDIFF $count=1 $X=1.045
+ $Y=1.84 $X2=1.235 $Y2=2.815
r53 1 25 400 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_PDIFF $count=1 $X=0.14
+ $Y=1.84 $X2=0.285 $Y2=2.115
r54 1 12 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=0.14
+ $Y=1.84 $X2=0.285 $Y2=2.815
.ends

.subckt PM_SKY130_FD_SC_HS__O311AI_2%VPWR 1 2 3 14 18 22 25 26 27 29 42 43 46 49
r68 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r69 46 47 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r70 42 43 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r71 40 43 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=5.52 $Y2=3.33
r72 40 50 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=4.08 $Y2=3.33
r73 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r74 37 49 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.28 $Y=3.33
+ $X2=4.115 $Y2=3.33
r75 37 39 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=4.28 $Y=3.33
+ $X2=4.56 $Y2=3.33
r76 36 50 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.08 $Y2=3.33
r77 35 36 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r78 33 47 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r79 32 35 156.578 $w=1.68e-07 $l=2.4e-06 $layer=LI1_cond $X=1.2 $Y=3.33 $X2=3.6
+ $Y2=3.33
r80 32 33 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r81 30 46 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.9 $Y=3.33
+ $X2=0.775 $Y2=3.33
r82 30 32 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=0.9 $Y=3.33 $X2=1.2
+ $Y2=3.33
r83 29 49 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.95 $Y=3.33
+ $X2=4.115 $Y2=3.33
r84 29 35 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=3.95 $Y=3.33 $X2=3.6
+ $Y2=3.33
r85 27 36 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=2.88 $Y=3.33
+ $X2=3.6 $Y2=3.33
r86 27 33 0.468274 $w=4.9e-07 $l=1.68e-06 $layer=MET1_cond $X=2.88 $Y=3.33
+ $X2=1.2 $Y2=3.33
r87 25 39 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=4.85 $Y=3.33
+ $X2=4.56 $Y2=3.33
r88 25 26 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.85 $Y=3.33
+ $X2=4.975 $Y2=3.33
r89 24 42 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=5.1 $Y=3.33 $X2=5.52
+ $Y2=3.33
r90 24 26 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.1 $Y=3.33
+ $X2=4.975 $Y2=3.33
r91 20 26 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.975 $Y=3.245
+ $X2=4.975 $Y2=3.33
r92 20 22 36.4172 $w=2.48e-07 $l=7.9e-07 $layer=LI1_cond $X=4.975 $Y=3.245
+ $X2=4.975 $Y2=2.455
r93 16 49 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.115 $Y=3.245
+ $X2=4.115 $Y2=3.33
r94 16 18 27.5888 $w=3.28e-07 $l=7.9e-07 $layer=LI1_cond $X=4.115 $Y=3.245
+ $X2=4.115 $Y2=2.455
r95 12 46 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.775 $Y=3.245
+ $X2=0.775 $Y2=3.33
r96 12 14 36.4172 $w=2.48e-07 $l=7.9e-07 $layer=LI1_cond $X=0.775 $Y=3.245
+ $X2=0.775 $Y2=2.455
r97 3 22 300 $w=1.7e-07 $l=6.85912e-07 $layer=licon1_PDIFF $count=2 $X=4.865
+ $Y=1.84 $X2=5.015 $Y2=2.455
r98 2 18 300 $w=1.7e-07 $l=6.85912e-07 $layer=licon1_PDIFF $count=2 $X=3.965
+ $Y=1.84 $X2=4.115 $Y2=2.455
r99 1 14 300 $w=1.7e-07 $l=6.85912e-07 $layer=licon1_PDIFF $count=2 $X=0.585
+ $Y=1.84 $X2=0.735 $Y2=2.455
.ends

.subckt PM_SKY130_FD_SC_HS__O311AI_2%A_307_368# 1 2 9 11 12 15
r26 13 15 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=3.215 $Y=2.905
+ $X2=3.215 $Y2=2.455
r27 11 13 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.13 $Y=2.99
+ $X2=3.215 $Y2=2.905
r28 11 12 78.9412 $w=1.68e-07 $l=1.21e-06 $layer=LI1_cond $X=3.13 $Y=2.99
+ $X2=1.92 $Y2=2.99
r29 7 12 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.755 $Y=2.905
+ $X2=1.92 $Y2=2.99
r30 7 9 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=1.755 $Y=2.905
+ $X2=1.755 $Y2=2.455
r31 2 15 300 $w=1.7e-07 $l=6.85912e-07 $layer=licon1_PDIFF $count=2 $X=3.065
+ $Y=1.84 $X2=3.215 $Y2=2.455
r32 1 9 300 $w=1.7e-07 $l=7.16607e-07 $layer=licon1_PDIFF $count=2 $X=1.535
+ $Y=1.84 $X2=1.755 $Y2=2.455
.ends

.subckt PM_SKY130_FD_SC_HS__O311AI_2%Y 1 2 3 4 5 6 21 25 27 31 33 35 37 39 43 46
+ 48 51 54 55 56 66
r92 61 66 1.32248 $w=3.03e-07 $l=3.5e-08 $layer=LI1_cond $X=4.552 $Y=0.96
+ $X2=4.552 $Y2=0.925
r93 55 56 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=4.565 $Y=1.295
+ $X2=4.565 $Y2=1.665
r94 55 67 5.76222 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=4.565 $Y=1.295
+ $X2=4.565 $Y2=1.13
r95 54 61 2.99104 $w=3.17e-07 $l=9.12688e-08 $layer=LI1_cond $X=4.565 $Y=1.045
+ $X2=4.552 $Y2=0.96
r96 54 67 2.99104 $w=3.17e-07 $l=8.5e-08 $layer=LI1_cond $X=4.565 $Y=1.045
+ $X2=4.565 $Y2=1.13
r97 54 66 2.45603 $w=3.03e-07 $l=6.5e-08 $layer=LI1_cond $X=4.552 $Y=0.86
+ $X2=4.552 $Y2=0.925
r98 49 56 9.95292 $w=3.28e-07 $l=2.85e-07 $layer=LI1_cond $X=4.565 $Y=1.95
+ $X2=4.565 $Y2=1.665
r99 49 51 1.96316 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.565 $Y=1.95
+ $X2=4.565 $Y2=2.035
r100 41 43 20.5135 $w=2.48e-07 $l=4.45e-07 $layer=LI1_cond $X=5.52 $Y=0.96
+ $X2=5.52 $Y2=0.515
r101 37 53 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.465 $Y=2.12
+ $X2=5.465 $Y2=2.035
r102 37 39 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=5.465 $Y=2.12
+ $X2=5.465 $Y2=2.815
r103 36 51 4.30018 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.73 $Y=2.035
+ $X2=4.565 $Y2=2.035
r104 35 53 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.3 $Y=2.035
+ $X2=5.465 $Y2=2.035
r105 35 36 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=5.3 $Y=2.035
+ $X2=4.73 $Y2=2.035
r106 34 54 3.66292 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.73 $Y=1.045
+ $X2=4.565 $Y2=1.045
r107 33 41 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=5.395 $Y=1.045
+ $X2=5.52 $Y2=0.96
r108 33 34 43.385 $w=1.68e-07 $l=6.65e-07 $layer=LI1_cond $X=5.395 $Y=1.045
+ $X2=4.73 $Y2=1.045
r109 29 51 1.96316 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.565 $Y=2.12
+ $X2=4.565 $Y2=2.035
r110 29 31 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=4.565 $Y=2.12
+ $X2=4.565 $Y2=2.4
r111 28 48 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.75 $Y=2.035
+ $X2=3.625 $Y2=2.035
r112 27 51 4.30018 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.4 $Y=2.035
+ $X2=4.565 $Y2=2.035
r113 27 28 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=4.4 $Y=2.035
+ $X2=3.75 $Y2=2.035
r114 23 48 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.625 $Y=2.12
+ $X2=3.625 $Y2=2.035
r115 23 25 32.0379 $w=2.48e-07 $l=6.95e-07 $layer=LI1_cond $X=3.625 $Y=2.12
+ $X2=3.625 $Y2=2.815
r116 22 46 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.93 $Y=2.035
+ $X2=2.765 $Y2=2.035
r117 21 48 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.5 $Y=2.035
+ $X2=3.625 $Y2=2.035
r118 21 22 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=3.5 $Y=2.035
+ $X2=2.93 $Y2=2.035
r119 6 53 400 $w=1.7e-07 $l=3.4187e-07 $layer=licon1_PDIFF $count=1 $X=5.315
+ $Y=1.84 $X2=5.465 $Y2=2.115
r120 6 39 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=5.315
+ $Y=1.84 $X2=5.465 $Y2=2.815
r121 5 51 600 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=4.415
+ $Y=1.84 $X2=4.565 $Y2=1.985
r122 5 31 300 $w=1.7e-07 $l=6.30555e-07 $layer=licon1_PDIFF $count=2 $X=4.415
+ $Y=1.84 $X2=4.565 $Y2=2.4
r123 4 48 400 $w=1.7e-07 $l=3.4187e-07 $layer=licon1_PDIFF $count=1 $X=3.515
+ $Y=1.84 $X2=3.665 $Y2=2.115
r124 4 25 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=3.515
+ $Y=1.84 $X2=3.665 $Y2=2.815
r125 3 46 300 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_PDIFF $count=2 $X=2.62
+ $Y=1.84 $X2=2.765 $Y2=2.115
r126 2 43 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=5.34
+ $Y=0.37 $X2=5.48 $Y2=0.515
r127 1 54 182 $w=1.7e-07 $l=5.57808e-07 $layer=licon1_NDIFF $count=1 $X=4.475
+ $Y=0.37 $X2=4.62 $Y2=0.86
.ends

.subckt PM_SKY130_FD_SC_HS__O311AI_2%A_27_74# 1 2 3 4 5 18 20 21 24 26 30 32 36
+ 38 42 44 45 46
c81 46 0 1.72564e-20 $X=3.1 $Y=1.095
r82 40 42 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=4.06 $Y=1.01
+ $X2=4.06 $Y2=0.86
r83 39 46 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.225 $Y=1.095
+ $X2=3.1 $Y2=1.095
r84 38 40 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.895 $Y=1.095
+ $X2=4.06 $Y2=1.01
r85 38 39 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.895 $Y=1.095
+ $X2=3.225 $Y2=1.095
r86 34 46 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.1 $Y=1.01
+ $X2=3.1 $Y2=1.095
r87 34 36 22.8184 $w=2.48e-07 $l=4.95e-07 $layer=LI1_cond $X=3.1 $Y=1.01 $X2=3.1
+ $Y2=0.515
r88 33 45 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.295 $Y=1.095
+ $X2=2.17 $Y2=1.095
r89 32 46 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.975 $Y=1.095
+ $X2=3.1 $Y2=1.095
r90 32 33 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=2.975 $Y=1.095
+ $X2=2.295 $Y2=1.095
r91 28 45 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.17 $Y=1.01
+ $X2=2.17 $Y2=1.095
r92 28 30 22.8184 $w=2.48e-07 $l=4.95e-07 $layer=LI1_cond $X=2.17 $Y=1.01
+ $X2=2.17 $Y2=0.515
r93 27 44 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.365 $Y=1.095
+ $X2=1.24 $Y2=1.095
r94 26 45 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.045 $Y=1.095
+ $X2=2.17 $Y2=1.095
r95 26 27 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=2.045 $Y=1.095
+ $X2=1.365 $Y2=1.095
r96 22 44 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.24 $Y=1.01
+ $X2=1.24 $Y2=1.095
r97 22 24 22.8184 $w=2.48e-07 $l=4.95e-07 $layer=LI1_cond $X=1.24 $Y=1.01
+ $X2=1.24 $Y2=0.515
r98 20 44 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.115 $Y=1.095
+ $X2=1.24 $Y2=1.095
r99 20 21 48.9305 $w=1.68e-07 $l=7.5e-07 $layer=LI1_cond $X=1.115 $Y=1.095
+ $X2=0.365 $Y2=1.095
r100 16 21 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.24 $Y=1.01
+ $X2=0.365 $Y2=1.095
r101 16 18 22.8184 $w=2.48e-07 $l=4.95e-07 $layer=LI1_cond $X=0.24 $Y=1.01
+ $X2=0.24 $Y2=0.515
r102 5 42 182 $w=1.7e-07 $l=5.55608e-07 $layer=licon1_NDIFF $count=1 $X=3.92
+ $Y=0.37 $X2=4.06 $Y2=0.86
r103 4 36 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.92
+ $Y=0.37 $X2=3.06 $Y2=0.515
r104 3 30 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.99
+ $Y=0.37 $X2=2.13 $Y2=0.515
r105 2 24 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.06
+ $Y=0.37 $X2=1.2 $Y2=0.515
r106 1 18 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__O311AI_2%VGND 1 2 3 12 16 20 22 24 29 34 44 45 48 51
+ 54
r67 54 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r68 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r69 48 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r70 44 45 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r71 42 45 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=3.12 $Y=0 $X2=5.52
+ $Y2=0
r72 41 44 156.578 $w=1.68e-07 $l=2.4e-06 $layer=LI1_cond $X=3.12 $Y=0 $X2=5.52
+ $Y2=0
r73 41 42 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r74 39 54 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.795 $Y=0 $X2=2.63
+ $Y2=0
r75 39 41 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=2.795 $Y=0 $X2=3.12
+ $Y2=0
r76 38 55 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r77 38 52 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.68
+ $Y2=0
r78 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r79 35 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.865 $Y=0 $X2=1.7
+ $Y2=0
r80 35 37 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=1.865 $Y=0 $X2=2.16
+ $Y2=0
r81 34 54 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.465 $Y=0 $X2=2.63
+ $Y2=0
r82 34 37 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=2.465 $Y=0 $X2=2.16
+ $Y2=0
r83 33 52 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=1.68
+ $Y2=0
r84 33 49 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r85 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r86 30 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.875 $Y=0 $X2=0.71
+ $Y2=0
r87 30 32 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.875 $Y=0 $X2=1.2
+ $Y2=0
r88 29 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.535 $Y=0 $X2=1.7
+ $Y2=0
r89 29 32 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=1.535 $Y=0 $X2=1.2
+ $Y2=0
r90 27 49 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r91 26 27 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r92 24 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.545 $Y=0 $X2=0.71
+ $Y2=0
r93 24 26 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.545 $Y=0 $X2=0.24
+ $Y2=0
r94 22 42 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.88 $Y=0 $X2=3.12
+ $Y2=0
r95 22 55 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.88 $Y=0 $X2=2.64
+ $Y2=0
r96 18 54 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.63 $Y=0.085
+ $X2=2.63 $Y2=0
r97 18 20 17.8105 $w=3.28e-07 $l=5.1e-07 $layer=LI1_cond $X=2.63 $Y=0.085
+ $X2=2.63 $Y2=0.595
r98 14 51 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.7 $Y=0.085 $X2=1.7
+ $Y2=0
r99 14 16 17.8105 $w=3.28e-07 $l=5.1e-07 $layer=LI1_cond $X=1.7 $Y=0.085 $X2=1.7
+ $Y2=0.595
r100 10 48 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.71 $Y=0.085
+ $X2=0.71 $Y2=0
r101 10 12 17.8105 $w=3.28e-07 $l=5.1e-07 $layer=LI1_cond $X=0.71 $Y=0.085
+ $X2=0.71 $Y2=0.595
r102 3 20 182 $w=1.7e-07 $l=2.98119e-07 $layer=licon1_NDIFF $count=1 $X=2.46
+ $Y=0.37 $X2=2.63 $Y2=0.595
r103 2 16 182 $w=1.7e-07 $l=2.90474e-07 $layer=licon1_NDIFF $count=1 $X=1.55
+ $Y=0.37 $X2=1.7 $Y2=0.595
r104 1 12 182 $w=1.7e-07 $l=2.86575e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.37 $X2=0.71 $Y2=0.595
.ends

.subckt PM_SKY130_FD_SC_HS__O311AI_2%A_670_74# 1 2 9 11 12 15
r25 13 15 5.06376 $w=3.28e-07 $l=1.45e-07 $layer=LI1_cond $X=5.05 $Y=0.425
+ $X2=5.05 $Y2=0.57
r26 11 13 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.885 $Y=0.34
+ $X2=5.05 $Y2=0.425
r27 11 12 75.6791 $w=1.68e-07 $l=1.16e-06 $layer=LI1_cond $X=4.885 $Y=0.34
+ $X2=3.725 $Y2=0.34
r28 7 12 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.56 $Y=0.425
+ $X2=3.725 $Y2=0.34
r29 7 9 5.93683 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=3.56 $Y=0.425 $X2=3.56
+ $Y2=0.595
r30 2 15 182 $w=1.7e-07 $l=2.60768e-07 $layer=licon1_NDIFF $count=1 $X=4.91
+ $Y=0.37 $X2=5.05 $Y2=0.57
r31 1 9 182 $w=1.7e-07 $l=3.1285e-07 $layer=licon1_NDIFF $count=1 $X=3.35
+ $Y=0.37 $X2=3.56 $Y2=0.595
.ends

