* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hs__o41ai_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
M1000 a_157_74# A1 VGND VNB nlowvt w=740000u l=150000u
+  ad=7.104e+11p pd=6.36e+06u as=6.327e+11p ps=4.67e+06u
M1001 a_157_74# A3 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1002 a_260_368# A4 Y VPB pshort w=1.12e+06u l=150000u
+  ad=3.808e+11p pd=2.92e+06u as=3.92e+11p ps=2.94e+06u
M1003 Y B1 VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=9.072e+11p ps=6.1e+06u
M1004 a_358_368# A3 a_260_368# VPB pshort w=1.12e+06u l=150000u
+  ad=4.704e+11p pd=3.08e+06u as=0p ps=0u
M1005 VPWR A1 a_472_368# VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=4.704e+11p ps=3.08e+06u
M1006 a_472_368# A2 a_358_368# VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VGND A2 a_157_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VGND A4 a_157_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_157_74# B1 Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
.ends
