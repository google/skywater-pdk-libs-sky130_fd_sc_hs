# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_hs__fahcon_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__fahcon_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  11.52000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425000 1.350000 0.805000 1.780000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.969000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.445000 1.180000 5.060000 1.550000 ;
    END
  END B
  PIN CI
    ANTENNAGATEAREA  0.525000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.675000 1.180000 8.005000 1.550000 ;
    END
  END CI
  PIN COUT_N
    ANTENNADIFFAREA  0.782600 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.790000 2.085000 6.175000 2.255000 ;
        RECT 5.790000 2.255000 6.120000 2.965000 ;
        RECT 6.005000 1.210000 6.650000 1.380000 ;
        RECT 6.005000 1.380000 6.175000 2.085000 ;
        RECT 6.320000 0.350000 6.650000 1.210000 ;
    END
  END COUT_N
  PIN SUM
    ANTENNADIFFAREA  0.541300 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 11.075000 1.820000 11.435000 2.980000 ;
        RECT 11.155000 0.350000 11.435000 1.130000 ;
        RECT 11.265000 1.130000 11.435000 1.820000 ;
    END
  END SUM
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 11.520000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 11.520000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 11.520000 0.085000 ;
      RECT  0.000000  3.245000 11.520000 3.415000 ;
      RECT  0.085000  0.480000  0.365000 0.980000 ;
      RECT  0.085000  0.980000  1.245000 1.150000 ;
      RECT  0.085000  1.150000  1.180000 1.180000 ;
      RECT  0.085000  1.180000  0.255000 1.950000 ;
      RECT  0.085000  1.950000  0.485000 2.980000 ;
      RECT  0.545000  0.085000  0.715000 0.480000 ;
      RECT  0.545000  0.480000  0.905000 0.810000 ;
      RECT  0.655000  1.950000  0.985000 3.245000 ;
      RECT  0.975000  1.180000  1.180000 1.680000 ;
      RECT  1.075000  0.255000  2.615000 0.425000 ;
      RECT  1.075000  0.425000  1.245000 0.980000 ;
      RECT  1.190000  1.850000  1.520000 2.905000 ;
      RECT  1.190000  2.905000  3.810000 3.075000 ;
      RECT  1.350000  1.320000  1.745000 1.490000 ;
      RECT  1.350000  1.490000  1.520000 1.850000 ;
      RECT  1.415000  0.595000  1.745000 1.320000 ;
      RECT  1.690000  1.660000  2.095000 1.830000 ;
      RECT  1.690000  1.830000  1.860000 2.565000 ;
      RECT  1.690000  2.565000  3.260000 2.735000 ;
      RECT  1.925000  0.595000  2.275000 1.325000 ;
      RECT  1.925000  1.325000  2.095000 1.660000 ;
      RECT  2.030000  2.000000  2.200000 2.225000 ;
      RECT  2.030000  2.225000  3.275000 2.395000 ;
      RECT  2.400000  1.805000  2.775000 2.055000 ;
      RECT  2.445000  0.425000  2.615000 0.725000 ;
      RECT  2.445000  0.725000  2.775000 1.805000 ;
      RECT  2.785000  0.255000  4.735000 0.425000 ;
      RECT  2.785000  0.425000  3.115000 0.555000 ;
      RECT  2.945000  0.725000  3.275000 2.225000 ;
      RECT  3.460000  0.645000  3.810000 2.905000 ;
      RECT  4.040000  0.425000  4.735000 1.010000 ;
      RECT  4.040000  1.010000  4.210000 1.805000 ;
      RECT  4.040000  1.805000  4.375000 2.965000 ;
      RECT  4.545000  1.805000  4.875000 3.245000 ;
      RECT  4.905000  0.085000  5.155000 0.965000 ;
      RECT  5.100000  1.975000  5.430000 2.965000 ;
      RECT  5.230000  1.135000  5.495000 1.305000 ;
      RECT  5.230000  1.305000  5.400000 1.975000 ;
      RECT  5.325000  0.390000  6.150000 0.640000 ;
      RECT  5.325000  0.640000  5.495000 1.135000 ;
      RECT  5.570000  1.475000  5.835000 1.805000 ;
      RECT  5.665000  0.810000  6.115000 1.040000 ;
      RECT  5.665000  1.040000  5.835000 1.475000 ;
      RECT  6.345000  1.550000  6.610000 1.880000 ;
      RECT  6.345000  2.085000  7.475000 2.970000 ;
      RECT  6.820000  0.810000  7.075000 1.130000 ;
      RECT  6.820000  1.130000  7.135000 1.800000 ;
      RECT  7.245000  0.350000  7.575000 0.960000 ;
      RECT  7.305000  0.960000  7.475000 2.085000 ;
      RECT  7.645000  1.940000  7.815000 3.245000 ;
      RECT  7.745000  0.085000  7.995000 1.010000 ;
      RECT  8.015000  1.820000  8.345000 2.320000 ;
      RECT  8.015000  2.320000 10.030000 2.490000 ;
      RECT  8.015000  2.490000  8.345000 2.980000 ;
      RECT  8.175000  0.350000  8.515000 1.130000 ;
      RECT  8.175000  1.130000  8.345000 1.820000 ;
      RECT  8.515000  1.300000  8.765000 1.550000 ;
      RECT  8.515000  1.550000  8.965000 1.780000 ;
      RECT  8.575000  2.660000  8.905000 2.870000 ;
      RECT  8.575000  2.870000 10.455000 3.040000 ;
      RECT  8.775000  0.255000 10.325000 0.425000 ;
      RECT  8.775000  0.425000  9.105000 1.130000 ;
      RECT  8.935000  1.130000  9.105000 1.210000 ;
      RECT  8.935000  1.210000  9.305000 1.380000 ;
      RECT  9.135000  1.380000  9.305000 1.820000 ;
      RECT  9.135000  1.820000  9.360000 2.150000 ;
      RECT  9.275000  0.810000  9.645000 1.040000 ;
      RECT  9.475000  1.040000  9.645000 1.260000 ;
      RECT  9.475000  1.260000  9.690000 1.590000 ;
      RECT  9.560000  1.820000 10.030000 2.320000 ;
      RECT  9.560000  2.490000 10.030000 2.700000 ;
      RECT  9.815000  0.595000  9.985000 0.920000 ;
      RECT  9.815000  0.920000 10.625000 1.090000 ;
      RECT  9.860000  1.260000 10.285000 1.590000 ;
      RECT  9.860000  1.590000 10.030000 1.820000 ;
      RECT 10.155000  0.425000 10.325000 0.580000 ;
      RECT 10.155000  0.580000 10.980000 0.750000 ;
      RECT 10.200000  1.760000 10.625000 1.930000 ;
      RECT 10.200000  1.930000 10.455000 2.870000 ;
      RECT 10.455000  1.090000 10.625000 1.760000 ;
      RECT 10.495000  0.085000 10.895000 0.410000 ;
      RECT 10.650000  2.100000 10.900000 3.245000 ;
      RECT 10.810000  0.750000 10.980000 1.300000 ;
      RECT 10.810000  1.300000 11.095000 1.630000 ;
    LAYER mcon ;
      RECT  0.155000 -0.085000  0.325000 0.085000 ;
      RECT  0.155000  3.245000  0.325000 3.415000 ;
      RECT  0.635000 -0.085000  0.805000 0.085000 ;
      RECT  0.635000  3.245000  0.805000 3.415000 ;
      RECT  1.115000 -0.085000  1.285000 0.085000 ;
      RECT  1.115000  3.245000  1.285000 3.415000 ;
      RECT  1.595000 -0.085000  1.765000 0.085000 ;
      RECT  1.595000  3.245000  1.765000 3.415000 ;
      RECT  2.075000 -0.085000  2.245000 0.085000 ;
      RECT  2.075000  0.840000  2.245000 1.010000 ;
      RECT  2.075000  3.245000  2.245000 3.415000 ;
      RECT  2.555000 -0.085000  2.725000 0.085000 ;
      RECT  2.555000  3.245000  2.725000 3.415000 ;
      RECT  3.035000 -0.085000  3.205000 0.085000 ;
      RECT  3.035000  1.580000  3.205000 1.750000 ;
      RECT  3.035000  3.245000  3.205000 3.415000 ;
      RECT  3.515000 -0.085000  3.685000 0.085000 ;
      RECT  3.515000  3.245000  3.685000 3.415000 ;
      RECT  3.995000 -0.085000  4.165000 0.085000 ;
      RECT  3.995000  3.245000  4.165000 3.415000 ;
      RECT  4.475000 -0.085000  4.645000 0.085000 ;
      RECT  4.475000  3.245000  4.645000 3.415000 ;
      RECT  4.955000 -0.085000  5.125000 0.085000 ;
      RECT  4.955000  3.245000  5.125000 3.415000 ;
      RECT  5.435000 -0.085000  5.605000 0.085000 ;
      RECT  5.435000  3.245000  5.605000 3.415000 ;
      RECT  5.915000 -0.085000  6.085000 0.085000 ;
      RECT  5.915000  0.840000  6.085000 1.010000 ;
      RECT  5.915000  3.245000  6.085000 3.415000 ;
      RECT  6.395000 -0.085000  6.565000 0.085000 ;
      RECT  6.395000  1.580000  6.565000 1.750000 ;
      RECT  6.395000  3.245000  6.565000 3.415000 ;
      RECT  6.875000 -0.085000  7.045000 0.085000 ;
      RECT  6.875000  0.840000  7.045000 1.010000 ;
      RECT  6.875000  3.245000  7.045000 3.415000 ;
      RECT  7.355000 -0.085000  7.525000 0.085000 ;
      RECT  7.355000  3.245000  7.525000 3.415000 ;
      RECT  7.835000 -0.085000  8.005000 0.085000 ;
      RECT  7.835000  3.245000  8.005000 3.415000 ;
      RECT  8.315000 -0.085000  8.485000 0.085000 ;
      RECT  8.315000  3.245000  8.485000 3.415000 ;
      RECT  8.795000 -0.085000  8.965000 0.085000 ;
      RECT  8.795000  1.580000  8.965000 1.750000 ;
      RECT  8.795000  3.245000  8.965000 3.415000 ;
      RECT  9.275000 -0.085000  9.445000 0.085000 ;
      RECT  9.275000  0.840000  9.445000 1.010000 ;
      RECT  9.275000  3.245000  9.445000 3.415000 ;
      RECT  9.755000 -0.085000  9.925000 0.085000 ;
      RECT  9.755000  3.245000  9.925000 3.415000 ;
      RECT 10.235000 -0.085000 10.405000 0.085000 ;
      RECT 10.235000  3.245000 10.405000 3.415000 ;
      RECT 10.715000 -0.085000 10.885000 0.085000 ;
      RECT 10.715000  3.245000 10.885000 3.415000 ;
      RECT 11.195000 -0.085000 11.365000 0.085000 ;
      RECT 11.195000  3.245000 11.365000 3.415000 ;
    LAYER met1 ;
      RECT 2.015000 0.810000 2.305000 0.855000 ;
      RECT 2.015000 0.855000 9.505000 0.995000 ;
      RECT 2.015000 0.995000 2.305000 1.040000 ;
      RECT 2.975000 1.550000 3.265000 1.595000 ;
      RECT 2.975000 1.595000 9.025000 1.735000 ;
      RECT 2.975000 1.735000 3.265000 1.780000 ;
      RECT 5.855000 0.810000 6.145000 0.855000 ;
      RECT 5.855000 0.995000 6.145000 1.040000 ;
      RECT 6.335000 1.550000 6.625000 1.595000 ;
      RECT 6.335000 1.735000 6.625000 1.780000 ;
      RECT 6.815000 0.810000 7.105000 0.855000 ;
      RECT 6.815000 0.995000 7.105000 1.040000 ;
      RECT 8.735000 1.550000 9.025000 1.595000 ;
      RECT 8.735000 1.735000 9.025000 1.780000 ;
      RECT 9.215000 0.810000 9.505000 0.855000 ;
      RECT 9.215000 0.995000 9.505000 1.040000 ;
  END
END sky130_fd_sc_hs__fahcon_1
END LIBRARY
