* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hs__and3b_2 A_N B C VGND VNB VPB VPWR X
M1000 VGND C a_454_74# VNB nlowvt w=740000u l=150000u
+  ad=6.8395e+11p pd=6.06e+06u as=3.108e+11p ps=2.32e+06u
M1001 VPWR a_284_368# X VPB pshort w=1.12e+06u l=150000u
+  ad=1.432e+12p pd=1.098e+07u as=3.528e+11p ps=2.87e+06u
M1002 X a_284_368# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.072e+11p pd=2.04e+06u as=0p ps=0u
M1003 a_284_368# B VPWR VPB pshort w=1e+06u l=150000u
+  ad=5.95e+11p pd=5.19e+06u as=0p ps=0u
M1004 VPWR C a_284_368# VPB pshort w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VPWR a_27_88# a_284_368# VPB pshort w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_454_74# B a_376_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=1.776e+11p ps=1.96e+06u
M1007 a_376_74# a_27_88# a_284_368# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1008 VPWR A_N a_27_88# VPB pshort w=840000u l=150000u
+  ad=0p pd=0u as=2.478e+11p ps=2.27e+06u
M1009 X a_284_368# VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VGND A_N a_27_88# VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=1.5675e+11p ps=1.67e+06u
M1011 VGND a_284_368# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
