* NGSPICE file created from sky130_fd_sc_hs__o311ai_4.ext - technology: sky130A

.subckt sky130_fd_sc_hs__o311ai_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
M1000 VGND A1 a_459_74# VNB nlowvt w=740000u l=150000u
+  ad=2.19225e+12p pd=1.657e+07u as=1.7316e+12p ps=1.652e+07u
M1001 a_459_74# A1 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1002 a_459_74# B1 a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=1.02765e+12p ps=1.022e+07u
M1003 VGND A2 a_459_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 Y C1 a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=4.181e+11p pd=4.09e+06u as=0p ps=0u
M1005 a_459_74# A2 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VGND A1 a_459_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 Y B1 VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=1.8536e+12p pd=1.227e+07u as=3.6176e+12p ps=1.99e+07u
M1008 VPWR C1 Y VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VPWR B1 Y VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_1350_368# A2 a_841_368# VPB pshort w=1.12e+06u l=150000u
+  ad=1.4e+12p pd=1.146e+07u as=1.8592e+12p ps=1.452e+07u
M1011 a_841_368# A3 Y VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_841_368# A2 a_1350_368# VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_841_368# A2 a_1350_368# VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_1350_368# A1 VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VGND A3 a_459_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_1350_368# A2 a_841_368# VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_459_74# A3 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_459_74# A1 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_27_74# B1 a_459_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_27_74# B1 a_459_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_459_74# A2 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 Y A3 a_841_368# VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_27_74# C1 Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 VPWR A1 a_1350_368# VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 a_27_74# C1 Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 Y C1 VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 a_841_368# A3 Y VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1028 Y A3 a_841_368# VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1029 VGND A3 a_459_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1030 VGND A2 a_459_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1031 a_1350_368# A1 VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1032 a_459_74# B1 a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1033 VPWR A1 a_1350_368# VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1034 Y C1 a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1035 a_459_74# A3 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

