# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_hs__o2111a_1
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_hs__o2111a_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.840000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.261000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.405000 1.300000 3.735000 1.780000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.261000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.715000 1.415000 3.235000 1.780000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.237000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.045000 1.415000 2.505000 1.780000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.237000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.545000 0.440000 1.875000 1.900000 ;
    END
  END C1
  PIN D1
    ANTENNAGATEAREA  0.237000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.005000 1.550000 1.335000 1.880000 ;
    END
  END D1
  PIN X
    ANTENNADIFFAREA  0.533900 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.095000 0.350000 0.355000 1.040000 ;
        RECT 0.095000 1.040000 0.265000 1.820000 ;
        RECT 0.095000 1.820000 0.445000 2.980000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 3.840000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 3.840000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.840000 0.085000 ;
      RECT 0.000000  3.245000 3.840000 3.415000 ;
      RECT 0.435000  1.210000 1.330000 1.380000 ;
      RECT 0.435000  1.380000 0.785000 1.550000 ;
      RECT 0.535000  0.085000 0.865000 1.040000 ;
      RECT 0.615000  1.550000 0.785000 2.070000 ;
      RECT 0.615000  2.070000 2.865000 2.240000 ;
      RECT 0.615000  2.410000 0.945000 3.245000 ;
      RECT 1.080000  0.350000 1.330000 1.210000 ;
      RECT 1.195000  2.240000 2.865000 2.245000 ;
      RECT 1.195000  2.245000 1.525000 2.925000 ;
      RECT 1.740000  2.455000 2.290000 3.245000 ;
      RECT 2.380000  0.350000 2.710000 0.960000 ;
      RECT 2.380000  0.960000 3.710000 1.130000 ;
      RECT 2.535000  2.045000 2.865000 2.070000 ;
      RECT 2.535000  2.245000 2.865000 2.925000 ;
      RECT 2.880000  0.085000 3.210000 0.790000 ;
      RECT 3.380000  0.350000 3.710000 0.960000 ;
      RECT 3.405000  1.950000 3.735000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
  END
END sky130_fd_sc_hs__o2111a_1
END LIBRARY
