* File: sky130_fd_sc_hs__and2b_2.pxi.spice
* Created: Thu Aug 27 20:32:00 2020
* 
x_PM_SKY130_FD_SC_HS__AND2B_2%A_N N_A_N_M1008_g N_A_N_c_59_n N_A_N_M1004_g A_N
+ N_A_N_c_60_n PM_SKY130_FD_SC_HS__AND2B_2%A_N
x_PM_SKY130_FD_SC_HS__AND2B_2%A_198_48# N_A_198_48#_M1001_d N_A_198_48#_M1006_d
+ N_A_198_48#_M1002_g N_A_198_48#_c_93_n N_A_198_48#_M1003_g N_A_198_48#_M1009_g
+ N_A_198_48#_c_94_n N_A_198_48#_M1005_g N_A_198_48#_c_87_n N_A_198_48#_c_88_n
+ N_A_198_48#_c_149_p N_A_198_48#_c_130_p N_A_198_48#_c_96_n N_A_198_48#_c_89_n
+ N_A_198_48#_c_90_n N_A_198_48#_c_91_n N_A_198_48#_c_92_n
+ PM_SKY130_FD_SC_HS__AND2B_2%A_198_48#
x_PM_SKY130_FD_SC_HS__AND2B_2%B N_B_c_183_n N_B_c_188_n N_B_M1006_g N_B_M1000_g
+ B N_B_c_184_n N_B_c_185_n N_B_c_186_n PM_SKY130_FD_SC_HS__AND2B_2%B
x_PM_SKY130_FD_SC_HS__AND2B_2%A_27_74# N_A_27_74#_M1008_s N_A_27_74#_M1004_s
+ N_A_27_74#_M1001_g N_A_27_74#_c_224_n N_A_27_74#_M1007_g N_A_27_74#_c_225_n
+ N_A_27_74#_c_226_n N_A_27_74#_c_227_n N_A_27_74#_c_228_n N_A_27_74#_c_256_n
+ N_A_27_74#_c_233_n N_A_27_74#_c_229_n N_A_27_74#_c_230_n
+ PM_SKY130_FD_SC_HS__AND2B_2%A_27_74#
x_PM_SKY130_FD_SC_HS__AND2B_2%VPWR N_VPWR_M1004_d N_VPWR_M1005_s N_VPWR_M1007_d
+ N_VPWR_c_308_n N_VPWR_c_309_n N_VPWR_c_310_n N_VPWR_c_311_n VPWR
+ N_VPWR_c_312_n N_VPWR_c_313_n N_VPWR_c_314_n N_VPWR_c_307_n
+ PM_SKY130_FD_SC_HS__AND2B_2%VPWR
x_PM_SKY130_FD_SC_HS__AND2B_2%X N_X_M1002_s N_X_M1003_d N_X_c_349_n N_X_c_350_n
+ X N_X_c_352_n N_X_c_351_n PM_SKY130_FD_SC_HS__AND2B_2%X
x_PM_SKY130_FD_SC_HS__AND2B_2%VGND N_VGND_M1008_d N_VGND_M1009_d N_VGND_c_385_n
+ VGND N_VGND_c_386_n N_VGND_c_387_n N_VGND_c_388_n N_VGND_c_389_n
+ N_VGND_c_390_n N_VGND_c_391_n PM_SKY130_FD_SC_HS__AND2B_2%VGND
cc_1 VNB N_A_N_M1008_g 0.0471947f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.645
cc_2 VNB N_A_N_c_59_n 0.0350404f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.765
cc_3 VNB N_A_N_c_60_n 0.0146504f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.515
cc_4 VNB N_A_198_48#_M1002_g 0.0222235f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_5 VNB N_A_198_48#_M1009_g 0.0229301f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_6 VNB N_A_198_48#_c_87_n 5.83691e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_7 VNB N_A_198_48#_c_88_n 0.016583f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_A_198_48#_c_89_n 0.0212534f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A_198_48#_c_90_n 0.00813058f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_198_48#_c_91_n 0.00335621f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_198_48#_c_92_n 0.0666858f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_B_c_183_n 0.00715513f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.645
cc_13 VNB N_B_c_184_n 0.0308569f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.515
cc_14 VNB N_B_c_185_n 0.0105112f $X=-0.19 $Y=-0.245 $X2=0.337 $Y2=1.515
cc_15 VNB N_B_c_186_n 0.0195323f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_27_74#_M1001_g 0.0298947f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_27_74#_c_224_n 0.0353906f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.515
cc_18 VNB N_A_27_74#_c_225_n 0.0280542f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_27_74#_c_226_n 0.00803206f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_27_74#_c_227_n 0.0102182f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_27_74#_c_228_n 0.0092086f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_27_74#_c_229_n 0.00141274f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_27_74#_c_230_n 0.0155316f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_VPWR_c_307_n 0.143779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_X_c_349_n 0.00240191f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_X_c_350_n 0.00417716f $X=-0.19 $Y=-0.245 $X2=0.337 $Y2=1.515
cc_27 VNB N_X_c_351_n 0.00120427f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_385_n 0.00900547f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_386_n 0.0191515f $X=-0.19 $Y=-0.245 $X2=0.337 $Y2=1.665
cc_30 VNB N_VGND_c_387_n 0.0299712f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_388_n 0.205711f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_389_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_390_n 0.0186948f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_391_n 0.0254342f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VPB N_A_N_c_59_n 0.0363148f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.765
cc_36 VPB N_A_N_c_60_n 0.00743971f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.515
cc_37 VPB N_A_198_48#_c_93_n 0.0163182f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.515
cc_38 VPB N_A_198_48#_c_94_n 0.0172945f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_39 VPB N_A_198_48#_c_87_n 0.00382312f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_40 VPB N_A_198_48#_c_96_n 0.0169966f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_41 VPB N_A_198_48#_c_92_n 0.0144806f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_42 VPB N_B_c_183_n 0.00435005f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.645
cc_43 VPB N_B_c_188_n 0.0239451f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.645
cc_44 VPB N_A_27_74#_c_224_n 0.0265849f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.515
cc_45 VPB N_A_27_74#_c_228_n 0.00342431f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_46 VPB N_A_27_74#_c_233_n 0.0351409f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_47 VPB N_A_27_74#_c_229_n 0.0103864f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_48 VPB N_VPWR_c_308_n 0.0195702f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_49 VPB N_VPWR_c_309_n 0.0206527f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_50 VPB N_VPWR_c_310_n 0.0121909f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_51 VPB N_VPWR_c_311_n 0.0233261f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_52 VPB N_VPWR_c_312_n 0.0208116f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_53 VPB N_VPWR_c_313_n 0.0276654f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_54 VPB N_VPWR_c_314_n 0.021352f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_55 VPB N_VPWR_c_307_n 0.065822f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_56 VPB N_X_c_352_n 0.00207956f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_57 VPB N_X_c_351_n 9.04994e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_58 N_A_N_M1008_g N_A_198_48#_M1002_g 0.0229244f $X=0.495 $Y=0.645 $X2=0 $Y2=0
cc_59 N_A_N_c_59_n N_A_198_48#_c_93_n 0.0206387f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_60 N_A_N_c_59_n N_A_198_48#_c_92_n 0.00907721f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_61 N_A_N_M1008_g N_A_27_74#_c_225_n 0.0141875f $X=0.495 $Y=0.645 $X2=0 $Y2=0
cc_62 N_A_N_M1008_g N_A_27_74#_c_226_n 0.0120599f $X=0.495 $Y=0.645 $X2=0 $Y2=0
cc_63 N_A_N_c_59_n N_A_27_74#_c_226_n 9.9484e-19 $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_64 N_A_N_c_60_n N_A_27_74#_c_226_n 0.00759305f $X=0.385 $Y=1.515 $X2=0 $Y2=0
cc_65 N_A_N_M1008_g N_A_27_74#_c_227_n 0.00419608f $X=0.495 $Y=0.645 $X2=0 $Y2=0
cc_66 N_A_N_c_59_n N_A_27_74#_c_227_n 0.00158281f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_67 N_A_N_c_60_n N_A_27_74#_c_227_n 0.02782f $X=0.385 $Y=1.515 $X2=0 $Y2=0
cc_68 N_A_N_M1008_g N_A_27_74#_c_228_n 0.00382916f $X=0.495 $Y=0.645 $X2=0 $Y2=0
cc_69 N_A_N_c_59_n N_A_27_74#_c_228_n 0.0076877f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_70 N_A_N_c_60_n N_A_27_74#_c_228_n 0.0329132f $X=0.385 $Y=1.515 $X2=0 $Y2=0
cc_71 N_A_N_c_59_n N_A_27_74#_c_233_n 0.0285771f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_72 N_A_N_c_60_n N_A_27_74#_c_233_n 0.0339846f $X=0.385 $Y=1.515 $X2=0 $Y2=0
cc_73 N_A_N_c_59_n N_VPWR_c_308_n 0.00357566f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_74 N_A_N_c_59_n N_VPWR_c_313_n 0.00393265f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_75 N_A_N_c_59_n N_VPWR_c_307_n 0.00462577f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_76 N_A_N_M1008_g N_X_c_349_n 6.3158e-19 $X=0.495 $Y=0.645 $X2=0 $Y2=0
cc_77 N_A_N_M1008_g N_VGND_c_385_n 0.00622602f $X=0.495 $Y=0.645 $X2=0 $Y2=0
cc_78 N_A_N_M1008_g N_VGND_c_386_n 0.00434272f $X=0.495 $Y=0.645 $X2=0 $Y2=0
cc_79 N_A_N_M1008_g N_VGND_c_388_n 0.0082497f $X=0.495 $Y=0.645 $X2=0 $Y2=0
cc_80 N_A_198_48#_c_90_n N_B_c_183_n 0.00233439f $X=1.62 $Y=1.465 $X2=0 $Y2=0
cc_81 N_A_198_48#_c_92_n N_B_c_183_n 0.00285107f $X=1.575 $Y=1.532 $X2=0 $Y2=0
cc_82 N_A_198_48#_c_94_n N_B_c_188_n 0.0164553f $X=1.575 $Y=1.765 $X2=0 $Y2=0
cc_83 N_A_198_48#_c_87_n N_B_c_188_n 0.00323752f $X=1.77 $Y=1.87 $X2=0 $Y2=0
cc_84 N_A_198_48#_c_96_n N_B_c_188_n 0.0157449f $X=2.63 $Y=2.05 $X2=0 $Y2=0
cc_85 N_A_198_48#_M1009_g N_B_c_184_n 8.98792e-19 $X=1.495 $Y=0.74 $X2=0 $Y2=0
cc_86 N_A_198_48#_c_88_n N_B_c_184_n 0.00101648f $X=2.89 $Y=0.925 $X2=0 $Y2=0
cc_87 N_A_198_48#_c_96_n N_B_c_184_n 0.00317892f $X=2.63 $Y=2.05 $X2=0 $Y2=0
cc_88 N_A_198_48#_c_91_n N_B_c_184_n 9.40265e-19 $X=1.655 $Y=1.3 $X2=0 $Y2=0
cc_89 N_A_198_48#_c_92_n N_B_c_184_n 0.00674836f $X=1.575 $Y=1.532 $X2=0 $Y2=0
cc_90 N_A_198_48#_c_88_n N_B_c_185_n 0.0347049f $X=2.89 $Y=0.925 $X2=0 $Y2=0
cc_91 N_A_198_48#_c_96_n N_B_c_185_n 0.0236465f $X=2.63 $Y=2.05 $X2=0 $Y2=0
cc_92 N_A_198_48#_c_91_n N_B_c_185_n 0.0290845f $X=1.655 $Y=1.3 $X2=0 $Y2=0
cc_93 N_A_198_48#_c_92_n N_B_c_185_n 8.78648e-19 $X=1.575 $Y=1.532 $X2=0 $Y2=0
cc_94 N_A_198_48#_c_88_n N_B_c_186_n 0.0140192f $X=2.89 $Y=0.925 $X2=0 $Y2=0
cc_95 N_A_198_48#_c_89_n N_B_c_186_n 0.00189613f $X=3.055 $Y=0.515 $X2=0 $Y2=0
cc_96 N_A_198_48#_c_91_n N_B_c_186_n 0.00418196f $X=1.655 $Y=1.3 $X2=0 $Y2=0
cc_97 N_A_198_48#_c_88_n N_A_27_74#_M1001_g 0.0120679f $X=2.89 $Y=0.925 $X2=0
+ $Y2=0
cc_98 N_A_198_48#_c_89_n N_A_27_74#_M1001_g 0.010211f $X=3.055 $Y=0.515 $X2=0
+ $Y2=0
cc_99 N_A_198_48#_c_88_n N_A_27_74#_c_224_n 0.00428484f $X=2.89 $Y=0.925 $X2=0
+ $Y2=0
cc_100 N_A_198_48#_c_96_n N_A_27_74#_c_224_n 0.00392882f $X=2.63 $Y=2.05 $X2=0
+ $Y2=0
cc_101 N_A_198_48#_M1002_g N_A_27_74#_c_225_n 6.28869e-19 $X=1.065 $Y=0.74 $X2=0
+ $Y2=0
cc_102 N_A_198_48#_M1002_g N_A_27_74#_c_226_n 0.00169872f $X=1.065 $Y=0.74 $X2=0
+ $Y2=0
cc_103 N_A_198_48#_M1002_g N_A_27_74#_c_228_n 0.00265413f $X=1.065 $Y=0.74 $X2=0
+ $Y2=0
cc_104 N_A_198_48#_c_93_n N_A_27_74#_c_228_n 0.00146566f $X=1.125 $Y=1.765 $X2=0
+ $Y2=0
cc_105 N_A_198_48#_c_92_n N_A_27_74#_c_228_n 0.00300277f $X=1.575 $Y=1.532 $X2=0
+ $Y2=0
cc_106 N_A_198_48#_M1006_d N_A_27_74#_c_256_n 0.00572155f $X=2.48 $Y=1.89 $X2=0
+ $Y2=0
cc_107 N_A_198_48#_c_93_n N_A_27_74#_c_256_n 0.0139601f $X=1.125 $Y=1.765 $X2=0
+ $Y2=0
cc_108 N_A_198_48#_c_94_n N_A_27_74#_c_256_n 0.017468f $X=1.575 $Y=1.765 $X2=0
+ $Y2=0
cc_109 N_A_198_48#_c_130_p N_A_27_74#_c_256_n 0.0119962f $X=1.855 $Y=2.01 $X2=0
+ $Y2=0
cc_110 N_A_198_48#_c_96_n N_A_27_74#_c_256_n 0.0570887f $X=2.63 $Y=2.05 $X2=0
+ $Y2=0
cc_111 N_A_198_48#_c_92_n N_A_27_74#_c_256_n 5.21741e-19 $X=1.575 $Y=1.532 $X2=0
+ $Y2=0
cc_112 N_A_198_48#_c_93_n N_A_27_74#_c_233_n 0.00758832f $X=1.125 $Y=1.765 $X2=0
+ $Y2=0
cc_113 N_A_198_48#_c_96_n N_A_27_74#_c_229_n 0.0123906f $X=2.63 $Y=2.05 $X2=0
+ $Y2=0
cc_114 N_A_198_48#_c_88_n N_A_27_74#_c_230_n 0.0265166f $X=2.89 $Y=0.925 $X2=0
+ $Y2=0
cc_115 N_A_198_48#_c_96_n N_A_27_74#_c_230_n 0.00174944f $X=2.63 $Y=2.05 $X2=0
+ $Y2=0
cc_116 N_A_198_48#_c_87_n N_VPWR_M1005_s 6.72919e-19 $X=1.77 $Y=1.87 $X2=0 $Y2=0
cc_117 N_A_198_48#_c_130_p N_VPWR_M1005_s 0.00386318f $X=1.855 $Y=2.01 $X2=0
+ $Y2=0
cc_118 N_A_198_48#_c_96_n N_VPWR_M1005_s 0.0111803f $X=2.63 $Y=2.05 $X2=0 $Y2=0
cc_119 N_A_198_48#_c_93_n N_VPWR_c_308_n 0.0104237f $X=1.125 $Y=1.765 $X2=0
+ $Y2=0
cc_120 N_A_198_48#_c_93_n N_VPWR_c_309_n 0.00461464f $X=1.125 $Y=1.765 $X2=0
+ $Y2=0
cc_121 N_A_198_48#_c_94_n N_VPWR_c_309_n 0.00415318f $X=1.575 $Y=1.765 $X2=0
+ $Y2=0
cc_122 N_A_198_48#_c_93_n N_VPWR_c_314_n 0.00130667f $X=1.125 $Y=1.765 $X2=0
+ $Y2=0
cc_123 N_A_198_48#_c_94_n N_VPWR_c_314_n 0.0173938f $X=1.575 $Y=1.765 $X2=0
+ $Y2=0
cc_124 N_A_198_48#_c_93_n N_VPWR_c_307_n 0.00469135f $X=1.125 $Y=1.765 $X2=0
+ $Y2=0
cc_125 N_A_198_48#_c_94_n N_VPWR_c_307_n 0.00414505f $X=1.575 $Y=1.765 $X2=0
+ $Y2=0
cc_126 N_A_198_48#_M1002_g N_X_c_349_n 0.0087663f $X=1.065 $Y=0.74 $X2=0 $Y2=0
cc_127 N_A_198_48#_M1009_g N_X_c_349_n 0.0158227f $X=1.495 $Y=0.74 $X2=0 $Y2=0
cc_128 N_A_198_48#_c_149_p N_X_c_349_n 0.0107372f $X=1.855 $Y=0.925 $X2=0 $Y2=0
cc_129 N_A_198_48#_M1002_g N_X_c_350_n 0.00252883f $X=1.065 $Y=0.74 $X2=0 $Y2=0
cc_130 N_A_198_48#_M1009_g N_X_c_350_n 0.00345782f $X=1.495 $Y=0.74 $X2=0 $Y2=0
cc_131 N_A_198_48#_c_91_n N_X_c_350_n 0.00679675f $X=1.655 $Y=1.3 $X2=0 $Y2=0
cc_132 N_A_198_48#_c_92_n N_X_c_350_n 0.00199986f $X=1.575 $Y=1.532 $X2=0 $Y2=0
cc_133 N_A_198_48#_c_93_n N_X_c_352_n 0.00880762f $X=1.125 $Y=1.765 $X2=0 $Y2=0
cc_134 N_A_198_48#_c_94_n N_X_c_352_n 0.00391362f $X=1.575 $Y=1.765 $X2=0 $Y2=0
cc_135 N_A_198_48#_c_87_n N_X_c_352_n 0.00266849f $X=1.77 $Y=1.87 $X2=0 $Y2=0
cc_136 N_A_198_48#_c_90_n N_X_c_352_n 0.00420181f $X=1.62 $Y=1.465 $X2=0 $Y2=0
cc_137 N_A_198_48#_c_92_n N_X_c_352_n 0.00793677f $X=1.575 $Y=1.532 $X2=0 $Y2=0
cc_138 N_A_198_48#_M1002_g N_X_c_351_n 0.00341038f $X=1.065 $Y=0.74 $X2=0 $Y2=0
cc_139 N_A_198_48#_c_93_n N_X_c_351_n 0.00142571f $X=1.125 $Y=1.765 $X2=0 $Y2=0
cc_140 N_A_198_48#_M1009_g N_X_c_351_n 0.00102916f $X=1.495 $Y=0.74 $X2=0 $Y2=0
cc_141 N_A_198_48#_c_87_n N_X_c_351_n 0.00578887f $X=1.77 $Y=1.87 $X2=0 $Y2=0
cc_142 N_A_198_48#_c_90_n N_X_c_351_n 0.0239361f $X=1.62 $Y=1.465 $X2=0 $Y2=0
cc_143 N_A_198_48#_c_91_n N_X_c_351_n 0.00495842f $X=1.655 $Y=1.3 $X2=0 $Y2=0
cc_144 N_A_198_48#_c_92_n N_X_c_351_n 0.0199288f $X=1.575 $Y=1.532 $X2=0 $Y2=0
cc_145 N_A_198_48#_c_88_n N_VGND_M1009_d 0.0186433f $X=2.89 $Y=0.925 $X2=0 $Y2=0
cc_146 N_A_198_48#_c_149_p N_VGND_M1009_d 0.00543344f $X=1.855 $Y=0.925 $X2=0
+ $Y2=0
cc_147 N_A_198_48#_c_91_n N_VGND_M1009_d 0.00340602f $X=1.655 $Y=1.3 $X2=0 $Y2=0
cc_148 N_A_198_48#_M1002_g N_VGND_c_385_n 0.00484286f $X=1.065 $Y=0.74 $X2=0
+ $Y2=0
cc_149 N_A_198_48#_c_89_n N_VGND_c_387_n 0.0145639f $X=3.055 $Y=0.515 $X2=0
+ $Y2=0
cc_150 N_A_198_48#_M1002_g N_VGND_c_388_n 0.00821312f $X=1.065 $Y=0.74 $X2=0
+ $Y2=0
cc_151 N_A_198_48#_M1009_g N_VGND_c_388_n 0.00825037f $X=1.495 $Y=0.74 $X2=0
+ $Y2=0
cc_152 N_A_198_48#_c_88_n N_VGND_c_388_n 0.0171606f $X=2.89 $Y=0.925 $X2=0 $Y2=0
cc_153 N_A_198_48#_c_149_p N_VGND_c_388_n 7.40526e-19 $X=1.855 $Y=0.925 $X2=0
+ $Y2=0
cc_154 N_A_198_48#_c_89_n N_VGND_c_388_n 0.0119984f $X=3.055 $Y=0.515 $X2=0
+ $Y2=0
cc_155 N_A_198_48#_M1002_g N_VGND_c_390_n 0.00434272f $X=1.065 $Y=0.74 $X2=0
+ $Y2=0
cc_156 N_A_198_48#_M1009_g N_VGND_c_390_n 0.00434272f $X=1.495 $Y=0.74 $X2=0
+ $Y2=0
cc_157 N_A_198_48#_M1009_g N_VGND_c_391_n 0.00838515f $X=1.495 $Y=0.74 $X2=0
+ $Y2=0
cc_158 N_A_198_48#_c_88_n N_VGND_c_391_n 0.0288531f $X=2.89 $Y=0.925 $X2=0 $Y2=0
cc_159 N_A_198_48#_c_149_p N_VGND_c_391_n 0.0111249f $X=1.855 $Y=0.925 $X2=0
+ $Y2=0
cc_160 N_A_198_48#_c_89_n N_VGND_c_391_n 0.00836615f $X=3.055 $Y=0.515 $X2=0
+ $Y2=0
cc_161 N_A_198_48#_c_88_n A_505_74# 0.00734082f $X=2.89 $Y=0.925 $X2=-0.19
+ $Y2=-0.245
cc_162 N_B_c_185_n N_A_27_74#_M1001_g 7.68955e-19 $X=2.36 $Y=1.385 $X2=0 $Y2=0
cc_163 N_B_c_186_n N_A_27_74#_M1001_g 0.0346115f $X=2.36 $Y=1.22 $X2=0 $Y2=0
cc_164 N_B_c_183_n N_A_27_74#_c_224_n 0.0126436f $X=2.405 $Y=1.725 $X2=0 $Y2=0
cc_165 N_B_c_188_n N_A_27_74#_c_224_n 0.0352665f $X=2.405 $Y=1.815 $X2=0 $Y2=0
cc_166 N_B_c_184_n N_A_27_74#_c_224_n 0.0346115f $X=2.36 $Y=1.385 $X2=0 $Y2=0
cc_167 N_B_c_185_n N_A_27_74#_c_224_n 3.1618e-19 $X=2.36 $Y=1.385 $X2=0 $Y2=0
cc_168 N_B_c_188_n N_A_27_74#_c_256_n 0.0133581f $X=2.405 $Y=1.815 $X2=0 $Y2=0
cc_169 N_B_c_183_n N_A_27_74#_c_230_n 5.05504e-19 $X=2.405 $Y=1.725 $X2=0 $Y2=0
cc_170 N_B_c_184_n N_A_27_74#_c_230_n 3.17209e-19 $X=2.36 $Y=1.385 $X2=0 $Y2=0
cc_171 N_B_c_185_n N_A_27_74#_c_230_n 0.0147792f $X=2.36 $Y=1.385 $X2=0 $Y2=0
cc_172 N_B_c_188_n N_VPWR_c_311_n 0.00109671f $X=2.405 $Y=1.815 $X2=0 $Y2=0
cc_173 N_B_c_188_n N_VPWR_c_312_n 0.00527445f $X=2.405 $Y=1.815 $X2=0 $Y2=0
cc_174 N_B_c_188_n N_VPWR_c_314_n 0.00712556f $X=2.405 $Y=1.815 $X2=0 $Y2=0
cc_175 N_B_c_188_n N_VPWR_c_307_n 0.00523671f $X=2.405 $Y=1.815 $X2=0 $Y2=0
cc_176 N_B_c_186_n N_VGND_c_387_n 0.00383152f $X=2.36 $Y=1.22 $X2=0 $Y2=0
cc_177 N_B_c_186_n N_VGND_c_388_n 0.00382027f $X=2.36 $Y=1.22 $X2=0 $Y2=0
cc_178 N_B_c_186_n N_VGND_c_391_n 0.0103112f $X=2.36 $Y=1.22 $X2=0 $Y2=0
cc_179 N_A_27_74#_c_228_n N_VPWR_M1004_d 0.00297742f $X=0.805 $Y=1.95 $X2=-0.19
+ $Y2=-0.245
cc_180 N_A_27_74#_c_256_n N_VPWR_M1004_d 0.00509611f $X=2.965 $Y=2.405 $X2=-0.19
+ $Y2=-0.245
cc_181 N_A_27_74#_c_233_n N_VPWR_M1004_d 0.0141925f $X=0.89 $Y=2.405 $X2=-0.19
+ $Y2=-0.245
cc_182 N_A_27_74#_c_256_n N_VPWR_M1005_s 0.0150071f $X=2.965 $Y=2.405 $X2=0
+ $Y2=0
cc_183 N_A_27_74#_c_256_n N_VPWR_M1007_d 0.00950867f $X=2.965 $Y=2.405 $X2=0
+ $Y2=0
cc_184 N_A_27_74#_c_229_n N_VPWR_M1007_d 0.0186475f $X=3.05 $Y=2.32 $X2=0 $Y2=0
cc_185 N_A_27_74#_c_256_n N_VPWR_c_308_n 0.00704757f $X=2.965 $Y=2.405 $X2=0
+ $Y2=0
cc_186 N_A_27_74#_c_233_n N_VPWR_c_308_n 0.023618f $X=0.89 $Y=2.405 $X2=0 $Y2=0
cc_187 N_A_27_74#_c_224_n N_VPWR_c_311_n 0.00988711f $X=2.855 $Y=1.815 $X2=0
+ $Y2=0
cc_188 N_A_27_74#_c_256_n N_VPWR_c_311_n 0.0139805f $X=2.965 $Y=2.405 $X2=0
+ $Y2=0
cc_189 N_A_27_74#_c_224_n N_VPWR_c_312_n 0.00473462f $X=2.855 $Y=1.815 $X2=0
+ $Y2=0
cc_190 N_A_27_74#_c_233_n N_VPWR_c_313_n 0.00671799f $X=0.89 $Y=2.405 $X2=0
+ $Y2=0
cc_191 N_A_27_74#_c_256_n N_VPWR_c_314_n 0.0449691f $X=2.965 $Y=2.405 $X2=0
+ $Y2=0
cc_192 N_A_27_74#_c_224_n N_VPWR_c_307_n 0.00474795f $X=2.855 $Y=1.815 $X2=0
+ $Y2=0
cc_193 N_A_27_74#_c_256_n N_VPWR_c_307_n 0.0454349f $X=2.965 $Y=2.405 $X2=0
+ $Y2=0
cc_194 N_A_27_74#_c_233_n N_VPWR_c_307_n 0.0183179f $X=0.89 $Y=2.405 $X2=0 $Y2=0
cc_195 N_A_27_74#_c_256_n N_X_M1003_d 0.00558496f $X=2.965 $Y=2.405 $X2=0 $Y2=0
cc_196 N_A_27_74#_c_225_n N_X_c_349_n 0.00402818f $X=0.28 $Y=0.645 $X2=0 $Y2=0
cc_197 N_A_27_74#_c_226_n N_X_c_350_n 0.011582f $X=0.72 $Y=1.095 $X2=0 $Y2=0
cc_198 N_A_27_74#_c_228_n N_X_c_352_n 0.00880966f $X=0.805 $Y=1.95 $X2=0 $Y2=0
cc_199 N_A_27_74#_c_256_n N_X_c_352_n 0.0238935f $X=2.965 $Y=2.405 $X2=0 $Y2=0
cc_200 N_A_27_74#_c_233_n N_X_c_352_n 0.0151329f $X=0.89 $Y=2.405 $X2=0 $Y2=0
cc_201 N_A_27_74#_c_228_n N_X_c_351_n 0.0373262f $X=0.805 $Y=1.95 $X2=0 $Y2=0
cc_202 N_A_27_74#_c_226_n N_VGND_M1008_d 0.00338852f $X=0.72 $Y=1.095 $X2=-0.19
+ $Y2=-0.245
cc_203 N_A_27_74#_c_225_n N_VGND_c_385_n 0.0191765f $X=0.28 $Y=0.645 $X2=0 $Y2=0
cc_204 N_A_27_74#_c_226_n N_VGND_c_385_n 0.0234311f $X=0.72 $Y=1.095 $X2=0 $Y2=0
cc_205 N_A_27_74#_c_225_n N_VGND_c_386_n 0.0145639f $X=0.28 $Y=0.645 $X2=0 $Y2=0
cc_206 N_A_27_74#_M1001_g N_VGND_c_387_n 0.00434272f $X=2.84 $Y=0.74 $X2=0 $Y2=0
cc_207 N_A_27_74#_M1001_g N_VGND_c_388_n 0.00449497f $X=2.84 $Y=0.74 $X2=0 $Y2=0
cc_208 N_A_27_74#_c_225_n N_VGND_c_388_n 0.0119984f $X=0.28 $Y=0.645 $X2=0 $Y2=0
cc_209 N_A_27_74#_M1001_g N_VGND_c_391_n 0.00126064f $X=2.84 $Y=0.74 $X2=0 $Y2=0
cc_210 N_X_c_349_n N_VGND_c_385_n 0.0191765f $X=1.28 $Y=0.515 $X2=0 $Y2=0
cc_211 N_X_c_349_n N_VGND_c_388_n 0.0118826f $X=1.28 $Y=0.515 $X2=0 $Y2=0
cc_212 N_X_c_349_n N_VGND_c_390_n 0.0144922f $X=1.28 $Y=0.515 $X2=0 $Y2=0
cc_213 N_X_c_349_n N_VGND_c_391_n 0.0102732f $X=1.28 $Y=0.515 $X2=0 $Y2=0
