* File: sky130_fd_sc_hs__a41oi_4.pxi.spice
* Created: Tue Sep  1 19:54:28 2020
* 
x_PM_SKY130_FD_SC_HS__A41OI_4%B1 N_B1_M1016_g N_B1_c_154_n N_B1_M1014_g
+ N_B1_M1035_g N_B1_c_155_n N_B1_M1018_g N_B1_c_156_n N_B1_M1019_g N_B1_c_151_n
+ N_B1_c_152_n N_B1_c_159_n N_B1_M1023_g B1 B1 B1 N_B1_c_153_n
+ PM_SKY130_FD_SC_HS__A41OI_4%B1
x_PM_SKY130_FD_SC_HS__A41OI_4%A1 N_A1_c_227_n N_A1_M1027_g N_A1_c_228_n
+ N_A1_c_229_n N_A1_c_235_n N_A1_M1012_g N_A1_c_230_n N_A1_M1029_g N_A1_c_236_n
+ N_A1_M1020_g N_A1_c_231_n N_A1_M1032_g N_A1_c_237_n N_A1_M1025_g N_A1_c_232_n
+ N_A1_M1037_g N_A1_c_238_n N_A1_M1026_g A1 A1 N_A1_c_233_n N_A1_c_234_n
+ PM_SKY130_FD_SC_HS__A41OI_4%A1
x_PM_SKY130_FD_SC_HS__A41OI_4%A2 N_A2_c_335_n N_A2_M1006_g N_A2_c_342_n
+ N_A2_M1000_g N_A2_c_336_n N_A2_M1007_g N_A2_c_343_n N_A2_M1001_g N_A2_c_337_n
+ N_A2_M1030_g N_A2_c_344_n N_A2_M1015_g N_A2_c_338_n N_A2_M1033_g N_A2_c_345_n
+ N_A2_M1031_g N_A2_c_339_n A2 A2 N_A2_c_340_n N_A2_c_341_n N_A2_c_348_n
+ PM_SKY130_FD_SC_HS__A41OI_4%A2
x_PM_SKY130_FD_SC_HS__A41OI_4%A3 N_A3_c_432_n N_A3_M1002_g N_A3_M1010_g
+ N_A3_c_433_n N_A3_M1004_g N_A3_M1024_g N_A3_c_434_n N_A3_M1008_g N_A3_M1028_g
+ N_A3_c_435_n N_A3_M1009_g N_A3_M1036_g A3 A3 A3 A3 A3 N_A3_c_431_n
+ PM_SKY130_FD_SC_HS__A41OI_4%A3
x_PM_SKY130_FD_SC_HS__A41OI_4%A4 N_A4_c_519_n N_A4_M1005_g N_A4_M1003_g
+ N_A4_c_520_n N_A4_M1011_g N_A4_M1017_g N_A4_M1022_g N_A4_c_521_n N_A4_M1013_g
+ N_A4_c_522_n N_A4_M1021_g N_A4_M1034_g A4 A4 A4 A4 N_A4_c_518_n
+ PM_SKY130_FD_SC_HS__A41OI_4%A4
x_PM_SKY130_FD_SC_HS__A41OI_4%A_27_368# N_A_27_368#_M1014_s N_A_27_368#_M1018_s
+ N_A_27_368#_M1023_s N_A_27_368#_M1020_d N_A_27_368#_M1026_d
+ N_A_27_368#_M1001_s N_A_27_368#_M1031_s N_A_27_368#_M1004_d
+ N_A_27_368#_M1009_d N_A_27_368#_M1011_s N_A_27_368#_M1021_s
+ N_A_27_368#_c_591_n N_A_27_368#_c_592_n N_A_27_368#_c_593_n
+ N_A_27_368#_c_612_n N_A_27_368#_c_594_n N_A_27_368#_c_616_n
+ N_A_27_368#_c_617_n N_A_27_368#_c_624_n N_A_27_368#_c_626_n
+ N_A_27_368#_c_629_n N_A_27_368#_c_630_n N_A_27_368#_c_595_n
+ N_A_27_368#_c_645_n N_A_27_368#_c_596_n N_A_27_368#_c_654_n
+ N_A_27_368#_c_597_n N_A_27_368#_c_670_n N_A_27_368#_c_598_n
+ N_A_27_368#_c_678_n N_A_27_368#_c_599_n N_A_27_368#_c_694_n
+ N_A_27_368#_c_600_n N_A_27_368#_c_702_n N_A_27_368#_c_601_n
+ N_A_27_368#_c_602_n N_A_27_368#_c_603_n N_A_27_368#_c_604_n
+ N_A_27_368#_c_638_n N_A_27_368#_c_605_n N_A_27_368#_c_667_n
+ N_A_27_368#_c_686_n N_A_27_368#_c_690_n N_A_27_368#_c_710_n
+ PM_SKY130_FD_SC_HS__A41OI_4%A_27_368#
x_PM_SKY130_FD_SC_HS__A41OI_4%Y N_Y_M1016_s N_Y_M1027_d N_Y_M1032_d N_Y_M1014_d
+ N_Y_M1019_d N_Y_c_788_n N_Y_c_789_n N_Y_c_790_n N_Y_c_806_n N_Y_c_791_n
+ N_Y_c_792_n N_Y_c_837_n N_Y_c_838_n N_Y_c_814_n N_Y_c_818_n N_Y_c_795_n
+ N_Y_c_846_n Y N_Y_c_793_n Y PM_SKY130_FD_SC_HS__A41OI_4%Y
x_PM_SKY130_FD_SC_HS__A41OI_4%VPWR N_VPWR_M1012_s N_VPWR_M1025_s N_VPWR_M1000_d
+ N_VPWR_M1015_d N_VPWR_M1002_s N_VPWR_M1008_s N_VPWR_M1005_d N_VPWR_M1013_d
+ N_VPWR_c_899_n N_VPWR_c_900_n N_VPWR_c_901_n N_VPWR_c_902_n N_VPWR_c_903_n
+ N_VPWR_c_904_n N_VPWR_c_905_n N_VPWR_c_906_n N_VPWR_c_907_n N_VPWR_c_908_n
+ N_VPWR_c_909_n N_VPWR_c_910_n N_VPWR_c_911_n N_VPWR_c_912_n N_VPWR_c_913_n
+ VPWR N_VPWR_c_914_n N_VPWR_c_915_n N_VPWR_c_916_n N_VPWR_c_898_n
+ N_VPWR_c_918_n N_VPWR_c_919_n N_VPWR_c_920_n N_VPWR_c_921_n N_VPWR_c_922_n
+ N_VPWR_c_923_n N_VPWR_c_924_n PM_SKY130_FD_SC_HS__A41OI_4%VPWR
x_PM_SKY130_FD_SC_HS__A41OI_4%VGND N_VGND_M1016_d N_VGND_M1035_d N_VGND_M1003_s
+ N_VGND_M1022_s N_VGND_c_1042_n N_VGND_c_1043_n N_VGND_c_1044_n N_VGND_c_1045_n
+ N_VGND_c_1046_n VGND N_VGND_c_1047_n N_VGND_c_1048_n N_VGND_c_1049_n
+ N_VGND_c_1050_n N_VGND_c_1051_n N_VGND_c_1052_n N_VGND_c_1053_n
+ N_VGND_c_1054_n PM_SKY130_FD_SC_HS__A41OI_4%VGND
x_PM_SKY130_FD_SC_HS__A41OI_4%A_325_74# N_A_325_74#_M1027_s N_A_325_74#_M1029_s
+ N_A_325_74#_M1037_s N_A_325_74#_M1007_s N_A_325_74#_M1033_s
+ N_A_325_74#_c_1141_n N_A_325_74#_c_1142_n N_A_325_74#_c_1143_n
+ N_A_325_74#_c_1144_n N_A_325_74#_c_1145_n N_A_325_74#_c_1146_n
+ N_A_325_74#_c_1147_n N_A_325_74#_c_1148_n
+ PM_SKY130_FD_SC_HS__A41OI_4%A_325_74#
x_PM_SKY130_FD_SC_HS__A41OI_4%A_852_74# N_A_852_74#_M1006_d N_A_852_74#_M1030_d
+ N_A_852_74#_M1010_s N_A_852_74#_M1028_s N_A_852_74#_c_1204_n
+ N_A_852_74#_c_1205_n PM_SKY130_FD_SC_HS__A41OI_4%A_852_74#
x_PM_SKY130_FD_SC_HS__A41OI_4%A_1235_74# N_A_1235_74#_M1010_d
+ N_A_1235_74#_M1024_d N_A_1235_74#_M1036_d N_A_1235_74#_M1017_d
+ N_A_1235_74#_M1034_d N_A_1235_74#_c_1235_n N_A_1235_74#_c_1236_n
+ N_A_1235_74#_c_1237_n N_A_1235_74#_c_1238_n N_A_1235_74#_c_1239_n
+ N_A_1235_74#_c_1240_n N_A_1235_74#_c_1241_n N_A_1235_74#_c_1242_n
+ N_A_1235_74#_c_1243_n PM_SKY130_FD_SC_HS__A41OI_4%A_1235_74#
cc_1 VNB N_B1_M1016_g 0.0315575f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_2 VNB N_B1_M1035_g 0.0315591f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=0.74
cc_3 VNB N_B1_c_151_n 0.0153571f $X=-0.19 $Y=-0.245 $X2=1.865 $Y2=1.64
cc_4 VNB N_B1_c_152_n 0.0714135f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=1.64
cc_5 VNB N_B1_c_153_n 0.0184974f $X=-0.19 $Y=-0.245 $X2=1.265 $Y2=1.515
cc_6 VNB N_A1_c_227_n 0.01857f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.35
cc_7 VNB N_A1_c_228_n 0.0132358f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_A1_c_229_n 0.00839791f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=1.765
cc_9 VNB N_A1_c_230_n 0.0179822f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=0.74
cc_10 VNB N_A1_c_231_n 0.0176901f $X=-0.19 $Y=-0.245 $X2=1.505 $Y2=1.765
cc_11 VNB N_A1_c_232_n 0.0157849f $X=-0.19 $Y=-0.245 $X2=1.955 $Y2=2.4
cc_12 VNB N_A1_c_233_n 0.00231182f $X=-0.19 $Y=-0.245 $X2=1.505 $Y2=1.557
cc_13 VNB N_A1_c_234_n 0.112291f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A2_c_335_n 0.0166764f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.35
cc_15 VNB N_A2_c_336_n 0.0158586f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=2.4
cc_16 VNB N_A2_c_337_n 0.015257f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=2.4
cc_17 VNB N_A2_c_338_n 0.0199171f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=1.64
cc_18 VNB N_A2_c_339_n 0.00252762f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A2_c_340_n 0.141226f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.565
cc_20 VNB N_A2_c_341_n 0.00352257f $X=-0.19 $Y=-0.245 $X2=1.2 $Y2=1.565
cc_21 VNB N_A3_M1010_g 0.0320084f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=2.4
cc_22 VNB N_A3_M1024_g 0.0234256f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=2.4
cc_23 VNB N_A3_M1028_g 0.0234234f $X=-0.19 $Y=-0.245 $X2=1.955 $Y2=1.765
cc_24 VNB N_A3_M1036_g 0.0240886f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB A3 0.00908404f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.515
cc_26 VNB N_A3_c_431_n 0.0804939f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A4_M1003_g 0.0230056f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=2.4
cc_28 VNB N_A4_M1017_g 0.0224899f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=2.4
cc_29 VNB N_A4_M1022_g 0.0230771f $X=-0.19 $Y=-0.245 $X2=1.505 $Y2=2.4
cc_30 VNB N_A4_M1034_g 0.0331137f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB A4 0.0166485f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.515
cc_32 VNB N_A4_c_518_n 0.074139f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_Y_c_788_n 0.00280455f $X=-0.19 $Y=-0.245 $X2=1.865 $Y2=1.64
cc_34 VNB N_Y_c_789_n 0.0168364f $X=-0.19 $Y=-0.245 $X2=1.955 $Y2=2.4
cc_35 VNB N_Y_c_790_n 0.00231148f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_36 VNB N_Y_c_791_n 0.0105726f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.557
cc_37 VNB N_Y_c_792_n 0.00412271f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.515
cc_38 VNB N_Y_c_793_n 8.52578e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_VPWR_c_898_n 0.422413f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_1042_n 0.010678f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=2.4
cc_41 VNB N_VGND_c_1043_n 0.043326f $X=-0.19 $Y=-0.245 $X2=1.505 $Y2=1.765
cc_42 VNB N_VGND_c_1044_n 0.0107076f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=1.64
cc_43 VNB N_VGND_c_1045_n 0.00323505f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_44 VNB N_VGND_c_1046_n 0.00574819f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_VGND_c_1047_n 0.018855f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.557
cc_46 VNB N_VGND_c_1048_n 0.163203f $X=-0.19 $Y=-0.245 $X2=1.265 $Y2=1.557
cc_47 VNB N_VGND_c_1049_n 0.0151736f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.565
cc_48 VNB N_VGND_c_1050_n 0.0188218f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_VGND_c_1051_n 0.533259f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_VGND_c_1052_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_VGND_c_1053_n 0.00604233f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_VGND_c_1054_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_A_325_74#_c_1141_n 0.00384069f $X=-0.19 $Y=-0.245 $X2=1.865 $Y2=1.64
cc_54 VNB N_A_325_74#_c_1142_n 0.00280532f $X=-0.19 $Y=-0.245 $X2=1.955
+ $Y2=1.765
cc_55 VNB N_A_325_74#_c_1143_n 0.00417961f $X=-0.19 $Y=-0.245 $X2=1.955 $Y2=2.4
cc_56 VNB N_A_325_74#_c_1144_n 0.00437333f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_57 VNB N_A_325_74#_c_1145_n 0.0026202f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_A_325_74#_c_1146_n 0.0133561f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=1.557
cc_59 VNB N_A_325_74#_c_1147_n 0.00496413f $X=-0.19 $Y=-0.245 $X2=1.265
+ $Y2=1.557
cc_60 VNB N_A_325_74#_c_1148_n 0.00609172f $X=-0.19 $Y=-0.245 $X2=1.265
+ $Y2=1.515
cc_61 VNB N_A_852_74#_c_1204_n 0.00251362f $X=-0.19 $Y=-0.245 $X2=1.955 $Y2=2.4
cc_62 VNB N_A_852_74#_c_1205_n 0.0283516f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_63 VNB N_A_1235_74#_c_1235_n 0.00754101f $X=-0.19 $Y=-0.245 $X2=1.505 $Y2=2.4
cc_64 VNB N_A_1235_74#_c_1236_n 0.0016059f $X=-0.19 $Y=-0.245 $X2=1.955
+ $Y2=1.765
cc_65 VNB N_A_1235_74#_c_1237_n 0.00323033f $X=-0.19 $Y=-0.245 $X2=0.635
+ $Y2=1.58
cc_66 VNB N_A_1235_74#_c_1238_n 0.00517531f $X=-0.19 $Y=-0.245 $X2=1.115
+ $Y2=1.58
cc_67 VNB N_A_1235_74#_c_1239_n 0.00178908f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_A_1235_74#_c_1240_n 0.0134691f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=1.557
cc_69 VNB N_A_1235_74#_c_1241_n 0.0266181f $X=-0.19 $Y=-0.245 $X2=0.995
+ $Y2=1.557
cc_70 VNB N_A_1235_74#_c_1242_n 0.00523512f $X=-0.19 $Y=-0.245 $X2=1.505
+ $Y2=1.557
cc_71 VNB N_A_1235_74#_c_1243_n 0.00127131f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VPB N_B1_c_154_n 0.0189957f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=1.765
cc_73 VPB N_B1_c_155_n 0.0153942f $X=-0.19 $Y=1.66 $X2=1.005 $Y2=1.765
cc_74 VPB N_B1_c_156_n 0.015061f $X=-0.19 $Y=1.66 $X2=1.505 $Y2=1.765
cc_75 VPB N_B1_c_151_n 0.0124581f $X=-0.19 $Y=1.66 $X2=1.865 $Y2=1.64
cc_76 VPB N_B1_c_152_n 0.0371843f $X=-0.19 $Y=1.66 $X2=1.595 $Y2=1.64
cc_77 VPB N_B1_c_159_n 0.0141058f $X=-0.19 $Y=1.66 $X2=1.955 $Y2=1.765
cc_78 VPB N_B1_c_153_n 0.0155975f $X=-0.19 $Y=1.66 $X2=1.265 $Y2=1.515
cc_79 VPB N_A1_c_235_n 0.0159363f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=2.4
cc_80 VPB N_A1_c_236_n 0.0162339f $X=-0.19 $Y=1.66 $X2=1.005 $Y2=1.765
cc_81 VPB N_A1_c_237_n 0.0156973f $X=-0.19 $Y=1.66 $X2=1.865 $Y2=1.64
cc_82 VPB N_A1_c_238_n 0.0162235f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_83 VPB N_A1_c_233_n 0.00759863f $X=-0.19 $Y=1.66 $X2=1.505 $Y2=1.557
cc_84 VPB N_A1_c_234_n 0.0535961f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_85 VPB N_A2_c_342_n 0.016235f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_86 VPB N_A2_c_343_n 0.0159674f $X=-0.19 $Y=1.66 $X2=0.995 $Y2=0.74
cc_87 VPB N_A2_c_344_n 0.0159004f $X=-0.19 $Y=1.66 $X2=1.505 $Y2=2.4
cc_88 VPB N_A2_c_345_n 0.0162194f $X=-0.19 $Y=1.66 $X2=1.955 $Y2=2.4
cc_89 VPB N_A2_c_340_n 0.0250732f $X=-0.19 $Y=1.66 $X2=0.72 $Y2=1.565
cc_90 VPB N_A2_c_341_n 0.00288228f $X=-0.19 $Y=1.66 $X2=1.2 $Y2=1.565
cc_91 VPB N_A2_c_348_n 0.0034614f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_92 VPB N_A3_c_432_n 0.0161662f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.35
cc_93 VPB N_A3_c_433_n 0.0158901f $X=-0.19 $Y=1.66 $X2=0.995 $Y2=1.35
cc_94 VPB N_A3_c_434_n 0.0158909f $X=-0.19 $Y=1.66 $X2=1.505 $Y2=1.765
cc_95 VPB N_A3_c_435_n 0.0165284f $X=-0.19 $Y=1.66 $X2=1.955 $Y2=2.4
cc_96 VPB A3 0.0151653f $X=-0.19 $Y=1.66 $X2=0.585 $Y2=1.515
cc_97 VPB N_A3_c_431_n 0.0522122f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_98 VPB N_A4_c_519_n 0.0157384f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.35
cc_99 VPB N_A4_c_520_n 0.0155127f $X=-0.19 $Y=1.66 $X2=0.995 $Y2=1.35
cc_100 VPB N_A4_c_521_n 0.0155127f $X=-0.19 $Y=1.66 $X2=1.595 $Y2=1.64
cc_101 VPB N_A4_c_522_n 0.0208611f $X=-0.19 $Y=1.66 $X2=1.955 $Y2=2.4
cc_102 VPB A4 0.0166366f $X=-0.19 $Y=1.66 $X2=0.585 $Y2=1.515
cc_103 VPB N_A4_c_518_n 0.047895f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_104 VPB N_A_27_368#_c_591_n 0.0366851f $X=-0.19 $Y=1.66 $X2=1.265 $Y2=1.557
cc_105 VPB N_A_27_368#_c_592_n 0.00269852f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=1.565
cc_106 VPB N_A_27_368#_c_593_n 0.00988933f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_107 VPB N_A_27_368#_c_594_n 0.00431993f $X=-0.19 $Y=1.66 $X2=1.2 $Y2=1.565
cc_108 VPB N_A_27_368#_c_595_n 0.00257348f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_109 VPB N_A_27_368#_c_596_n 0.00257348f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_110 VPB N_A_27_368#_c_597_n 0.00257348f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_111 VPB N_A_27_368#_c_598_n 0.00257348f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_112 VPB N_A_27_368#_c_599_n 0.00289722f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_113 VPB N_A_27_368#_c_600_n 0.00257348f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_114 VPB N_A_27_368#_c_601_n 0.00739392f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_115 VPB N_A_27_368#_c_602_n 0.0353617f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_116 VPB N_A_27_368#_c_603_n 0.0022931f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_117 VPB N_A_27_368#_c_604_n 0.00257417f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_118 VPB N_A_27_368#_c_605_n 0.00183525f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_119 VPB N_Y_c_791_n 0.00254319f $X=-0.19 $Y=1.66 $X2=0.585 $Y2=1.557
cc_120 VPB N_Y_c_795_n 0.00214877f $X=-0.19 $Y=1.66 $X2=1.2 $Y2=1.565
cc_121 VPB Y 8.23063e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_122 VPB N_VPWR_c_899_n 0.00928771f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_123 VPB N_VPWR_c_900_n 0.0196495f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.557
cc_124 VPB N_VPWR_c_901_n 0.00890006f $X=-0.19 $Y=1.66 $X2=0.585 $Y2=1.515
cc_125 VPB N_VPWR_c_902_n 0.0198086f $X=-0.19 $Y=1.66 $X2=1.005 $Y2=1.557
cc_126 VPB N_VPWR_c_903_n 0.00892434f $X=-0.19 $Y=1.66 $X2=1.505 $Y2=1.557
cc_127 VPB N_VPWR_c_904_n 0.0199677f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_128 VPB N_VPWR_c_905_n 0.00886117f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_129 VPB N_VPWR_c_906_n 0.0196495f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_130 VPB N_VPWR_c_907_n 0.00886117f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_131 VPB N_VPWR_c_908_n 0.0196495f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_132 VPB N_VPWR_c_909_n 0.0082016f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_133 VPB N_VPWR_c_910_n 0.00516621f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_134 VPB N_VPWR_c_911_n 0.00799266f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_135 VPB N_VPWR_c_912_n 0.0206041f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_136 VPB N_VPWR_c_913_n 0.00324402f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_137 VPB N_VPWR_c_914_n 0.0604982f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_138 VPB N_VPWR_c_915_n 0.0185368f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_139 VPB N_VPWR_c_916_n 0.0202453f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_140 VPB N_VPWR_c_898_n 0.109292f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_141 VPB N_VPWR_c_918_n 0.00631788f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_142 VPB N_VPWR_c_919_n 0.0047828f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_143 VPB N_VPWR_c_920_n 0.0047828f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_144 VPB N_VPWR_c_921_n 0.0047828f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_145 VPB N_VPWR_c_922_n 0.0047828f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_146 VPB N_VPWR_c_923_n 0.0047828f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_147 VPB N_VPWR_c_924_n 0.00460249f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_148 N_B1_c_151_n N_A1_c_229_n 0.00882381f $X=1.865 $Y=1.64 $X2=0 $Y2=0
cc_149 N_B1_c_159_n N_A1_c_235_n 0.0240212f $X=1.955 $Y=1.765 $X2=0 $Y2=0
cc_150 N_B1_c_151_n N_A1_c_233_n 2.71309e-19 $X=1.865 $Y=1.64 $X2=0 $Y2=0
cc_151 N_B1_c_151_n N_A1_c_234_n 0.010913f $X=1.865 $Y=1.64 $X2=0 $Y2=0
cc_152 N_B1_c_152_n N_A1_c_234_n 0.00226331f $X=1.595 $Y=1.64 $X2=0 $Y2=0
cc_153 N_B1_c_154_n N_A_27_368#_c_591_n 0.0106095f $X=0.51 $Y=1.765 $X2=0 $Y2=0
cc_154 N_B1_c_155_n N_A_27_368#_c_591_n 6.04056e-19 $X=1.005 $Y=1.765 $X2=0
+ $Y2=0
cc_155 N_B1_c_153_n N_A_27_368#_c_591_n 0.025553f $X=1.265 $Y=1.515 $X2=0 $Y2=0
cc_156 N_B1_c_154_n N_A_27_368#_c_592_n 0.0114142f $X=0.51 $Y=1.765 $X2=0 $Y2=0
cc_157 N_B1_c_155_n N_A_27_368#_c_592_n 0.0141012f $X=1.005 $Y=1.765 $X2=0 $Y2=0
cc_158 N_B1_c_154_n N_A_27_368#_c_593_n 0.00253309f $X=0.51 $Y=1.765 $X2=0 $Y2=0
cc_159 N_B1_c_156_n N_A_27_368#_c_612_n 0.00791006f $X=1.505 $Y=1.765 $X2=0
+ $Y2=0
cc_160 N_B1_c_159_n N_A_27_368#_c_612_n 5.7112e-19 $X=1.955 $Y=1.765 $X2=0 $Y2=0
cc_161 N_B1_c_156_n N_A_27_368#_c_594_n 0.0108414f $X=1.505 $Y=1.765 $X2=0 $Y2=0
cc_162 N_B1_c_159_n N_A_27_368#_c_594_n 0.0125587f $X=1.955 $Y=1.765 $X2=0 $Y2=0
cc_163 N_B1_c_159_n N_A_27_368#_c_616_n 0.00193585f $X=1.955 $Y=1.765 $X2=0
+ $Y2=0
cc_164 N_B1_c_156_n N_A_27_368#_c_617_n 5.19141e-19 $X=1.505 $Y=1.765 $X2=0
+ $Y2=0
cc_165 N_B1_c_159_n N_A_27_368#_c_617_n 0.00636367f $X=1.955 $Y=1.765 $X2=0
+ $Y2=0
cc_166 N_B1_c_156_n N_A_27_368#_c_603_n 0.00193739f $X=1.505 $Y=1.765 $X2=0
+ $Y2=0
cc_167 N_B1_M1016_g N_Y_c_788_n 0.00838277f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_168 N_B1_M1035_g N_Y_c_788_n 0.00350341f $X=0.995 $Y=0.74 $X2=0 $Y2=0
cc_169 N_B1_M1035_g N_Y_c_789_n 0.0167736f $X=0.995 $Y=0.74 $X2=0 $Y2=0
cc_170 N_B1_c_151_n N_Y_c_789_n 0.00445057f $X=1.865 $Y=1.64 $X2=0 $Y2=0
cc_171 N_B1_c_152_n N_Y_c_789_n 0.0150996f $X=1.595 $Y=1.64 $X2=0 $Y2=0
cc_172 N_B1_c_153_n N_Y_c_789_n 0.041974f $X=1.265 $Y=1.515 $X2=0 $Y2=0
cc_173 N_B1_M1016_g N_Y_c_790_n 0.00502286f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_174 N_B1_c_152_n N_Y_c_790_n 0.00404034f $X=1.595 $Y=1.64 $X2=0 $Y2=0
cc_175 N_B1_c_153_n N_Y_c_790_n 0.0282341f $X=1.265 $Y=1.515 $X2=0 $Y2=0
cc_176 N_B1_c_156_n N_Y_c_806_n 0.00556293f $X=1.505 $Y=1.765 $X2=0 $Y2=0
cc_177 N_B1_c_159_n N_Y_c_806_n 0.0055605f $X=1.955 $Y=1.765 $X2=0 $Y2=0
cc_178 N_B1_c_156_n N_Y_c_791_n 9.82568e-19 $X=1.505 $Y=1.765 $X2=0 $Y2=0
cc_179 N_B1_c_151_n N_Y_c_791_n 0.0128215f $X=1.865 $Y=1.64 $X2=0 $Y2=0
cc_180 N_B1_c_152_n N_Y_c_791_n 0.003371f $X=1.595 $Y=1.64 $X2=0 $Y2=0
cc_181 N_B1_c_159_n N_Y_c_791_n 0.00184424f $X=1.955 $Y=1.765 $X2=0 $Y2=0
cc_182 N_B1_c_153_n N_Y_c_791_n 0.0186052f $X=1.265 $Y=1.515 $X2=0 $Y2=0
cc_183 N_B1_c_151_n N_Y_c_792_n 3.13305e-19 $X=1.865 $Y=1.64 $X2=0 $Y2=0
cc_184 N_B1_c_155_n N_Y_c_814_n 0.00975321f $X=1.005 $Y=1.765 $X2=0 $Y2=0
cc_185 N_B1_c_156_n N_Y_c_814_n 7.14259e-19 $X=1.505 $Y=1.765 $X2=0 $Y2=0
cc_186 N_B1_c_152_n N_Y_c_814_n 0.00180944f $X=1.595 $Y=1.64 $X2=0 $Y2=0
cc_187 N_B1_c_153_n N_Y_c_814_n 0.0252535f $X=1.265 $Y=1.515 $X2=0 $Y2=0
cc_188 N_B1_c_155_n N_Y_c_818_n 0.0122806f $X=1.005 $Y=1.765 $X2=0 $Y2=0
cc_189 N_B1_c_156_n N_Y_c_818_n 0.0172462f $X=1.505 $Y=1.765 $X2=0 $Y2=0
cc_190 N_B1_c_151_n N_Y_c_818_n 8.8529e-19 $X=1.865 $Y=1.64 $X2=0 $Y2=0
cc_191 N_B1_c_152_n N_Y_c_818_n 0.00173082f $X=1.595 $Y=1.64 $X2=0 $Y2=0
cc_192 N_B1_c_153_n N_Y_c_818_n 0.0335538f $X=1.265 $Y=1.515 $X2=0 $Y2=0
cc_193 N_B1_c_156_n N_Y_c_795_n 0.0032427f $X=1.505 $Y=1.765 $X2=0 $Y2=0
cc_194 N_B1_c_151_n N_Y_c_795_n 0.00519069f $X=1.865 $Y=1.64 $X2=0 $Y2=0
cc_195 N_B1_c_159_n N_Y_c_795_n 0.0141959f $X=1.955 $Y=1.765 $X2=0 $Y2=0
cc_196 N_B1_c_154_n N_VPWR_c_914_n 0.00278262f $X=0.51 $Y=1.765 $X2=0 $Y2=0
cc_197 N_B1_c_155_n N_VPWR_c_914_n 0.00278271f $X=1.005 $Y=1.765 $X2=0 $Y2=0
cc_198 N_B1_c_156_n N_VPWR_c_914_n 0.00278257f $X=1.505 $Y=1.765 $X2=0 $Y2=0
cc_199 N_B1_c_159_n N_VPWR_c_914_n 0.00278257f $X=1.955 $Y=1.765 $X2=0 $Y2=0
cc_200 N_B1_c_154_n N_VPWR_c_898_n 0.0035775f $X=0.51 $Y=1.765 $X2=0 $Y2=0
cc_201 N_B1_c_155_n N_VPWR_c_898_n 0.00354701f $X=1.005 $Y=1.765 $X2=0 $Y2=0
cc_202 N_B1_c_156_n N_VPWR_c_898_n 0.00354283f $X=1.505 $Y=1.765 $X2=0 $Y2=0
cc_203 N_B1_c_159_n N_VPWR_c_898_n 0.00353905f $X=1.955 $Y=1.765 $X2=0 $Y2=0
cc_204 N_B1_M1016_g N_VGND_c_1043_n 0.00647381f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_205 N_B1_c_153_n N_VGND_c_1043_n 0.0179756f $X=1.265 $Y=1.515 $X2=0 $Y2=0
cc_206 N_B1_M1016_g N_VGND_c_1044_n 6.83978e-19 $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_207 N_B1_M1035_g N_VGND_c_1044_n 0.012834f $X=0.995 $Y=0.74 $X2=0 $Y2=0
cc_208 N_B1_M1016_g N_VGND_c_1047_n 0.00434272f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_209 N_B1_M1035_g N_VGND_c_1047_n 0.00383152f $X=0.995 $Y=0.74 $X2=0 $Y2=0
cc_210 N_B1_M1016_g N_VGND_c_1051_n 0.008246f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_211 N_B1_M1035_g N_VGND_c_1051_n 0.00758198f $X=0.995 $Y=0.74 $X2=0 $Y2=0
cc_212 N_B1_M1035_g N_A_325_74#_c_1141_n 8.38994e-19 $X=0.995 $Y=0.74 $X2=0
+ $Y2=0
cc_213 N_B1_M1035_g N_A_325_74#_c_1143_n 7.24903e-19 $X=0.995 $Y=0.74 $X2=0
+ $Y2=0
cc_214 N_A1_c_232_n N_A2_c_335_n 0.0123861f $X=3.685 $Y=1.205 $X2=-0.19
+ $Y2=-0.245
cc_215 N_A1_c_238_n N_A2_c_342_n 0.00873349f $X=3.91 $Y=1.765 $X2=0 $Y2=0
cc_216 N_A1_c_234_n N_A2_c_340_n 0.0250019f $X=3.685 $Y=1.485 $X2=0 $Y2=0
cc_217 N_A1_c_238_n N_A2_c_341_n 6.6009e-19 $X=3.91 $Y=1.765 $X2=0 $Y2=0
cc_218 N_A1_c_234_n N_A2_c_341_n 0.00968288f $X=3.685 $Y=1.485 $X2=0 $Y2=0
cc_219 N_A1_c_235_n N_A_27_368#_c_594_n 0.00313312f $X=2.405 $Y=1.765 $X2=0
+ $Y2=0
cc_220 N_A1_c_235_n N_A_27_368#_c_616_n 4.27055e-19 $X=2.405 $Y=1.765 $X2=0
+ $Y2=0
cc_221 N_A1_c_235_n N_A_27_368#_c_617_n 0.00656166f $X=2.405 $Y=1.765 $X2=0
+ $Y2=0
cc_222 N_A1_c_236_n N_A_27_368#_c_617_n 5.78806e-19 $X=2.955 $Y=1.765 $X2=0
+ $Y2=0
cc_223 N_A1_c_235_n N_A_27_368#_c_624_n 0.0123082f $X=2.405 $Y=1.765 $X2=0 $Y2=0
cc_224 N_A1_c_236_n N_A_27_368#_c_624_n 0.0123082f $X=2.955 $Y=1.765 $X2=0 $Y2=0
cc_225 N_A1_c_237_n N_A_27_368#_c_626_n 0.0120804f $X=3.405 $Y=1.765 $X2=0 $Y2=0
cc_226 N_A1_c_238_n N_A_27_368#_c_626_n 0.0158396f $X=3.91 $Y=1.765 $X2=0 $Y2=0
cc_227 N_A1_c_234_n N_A_27_368#_c_626_n 0.00282462f $X=3.685 $Y=1.485 $X2=0
+ $Y2=0
cc_228 N_A1_c_238_n N_A_27_368#_c_629_n 0.00216792f $X=3.91 $Y=1.765 $X2=0 $Y2=0
cc_229 N_A1_c_237_n N_A_27_368#_c_630_n 7.83052e-19 $X=3.405 $Y=1.765 $X2=0
+ $Y2=0
cc_230 N_A1_c_238_n N_A_27_368#_c_630_n 0.0032558f $X=3.91 $Y=1.765 $X2=0 $Y2=0
cc_231 N_A1_c_237_n N_A_27_368#_c_595_n 5.28386e-19 $X=3.405 $Y=1.765 $X2=0
+ $Y2=0
cc_232 N_A1_c_238_n N_A_27_368#_c_595_n 0.00690874f $X=3.91 $Y=1.765 $X2=0 $Y2=0
cc_233 N_A1_c_235_n N_A_27_368#_c_604_n 5.94284e-19 $X=2.405 $Y=1.765 $X2=0
+ $Y2=0
cc_234 N_A1_c_236_n N_A_27_368#_c_604_n 0.00809959f $X=2.955 $Y=1.765 $X2=0
+ $Y2=0
cc_235 N_A1_c_237_n N_A_27_368#_c_604_n 0.00817155f $X=3.405 $Y=1.765 $X2=0
+ $Y2=0
cc_236 N_A1_c_238_n N_A_27_368#_c_604_n 6.08656e-19 $X=3.91 $Y=1.765 $X2=0 $Y2=0
cc_237 N_A1_c_238_n N_A_27_368#_c_638_n 2.24111e-19 $X=3.91 $Y=1.765 $X2=0 $Y2=0
cc_238 N_A1_c_227_n N_Y_c_791_n 0.00133985f $X=1.985 $Y=1.205 $X2=0 $Y2=0
cc_239 N_A1_c_228_n N_Y_c_791_n 0.00843072f $X=2.285 $Y=1.28 $X2=0 $Y2=0
cc_240 N_A1_c_229_n N_Y_c_791_n 0.00605915f $X=2.06 $Y=1.28 $X2=0 $Y2=0
cc_241 N_A1_c_235_n N_Y_c_791_n 9.32379e-19 $X=2.405 $Y=1.765 $X2=0 $Y2=0
cc_242 N_A1_c_230_n N_Y_c_791_n 5.00179e-19 $X=2.485 $Y=1.205 $X2=0 $Y2=0
cc_243 N_A1_c_233_n N_Y_c_791_n 0.0341986f $X=3.13 $Y=1.515 $X2=0 $Y2=0
cc_244 N_A1_c_234_n N_Y_c_791_n 0.00160355f $X=3.685 $Y=1.485 $X2=0 $Y2=0
cc_245 N_A1_c_227_n N_Y_c_792_n 0.0129676f $X=1.985 $Y=1.205 $X2=0 $Y2=0
cc_246 N_A1_c_228_n N_Y_c_792_n 0.00642903f $X=2.285 $Y=1.28 $X2=0 $Y2=0
cc_247 N_A1_c_230_n N_Y_c_792_n 0.00641298f $X=2.485 $Y=1.205 $X2=0 $Y2=0
cc_248 N_A1_c_233_n N_Y_c_792_n 0.0114135f $X=3.13 $Y=1.515 $X2=0 $Y2=0
cc_249 N_A1_c_230_n N_Y_c_837_n 0.0054833f $X=2.485 $Y=1.205 $X2=0 $Y2=0
cc_250 N_A1_c_228_n N_Y_c_838_n 0.00401797f $X=2.285 $Y=1.28 $X2=0 $Y2=0
cc_251 N_A1_c_235_n N_Y_c_838_n 0.011193f $X=2.405 $Y=1.765 $X2=0 $Y2=0
cc_252 N_A1_c_236_n N_Y_c_838_n 0.011193f $X=2.955 $Y=1.765 $X2=0 $Y2=0
cc_253 N_A1_c_237_n N_Y_c_838_n 0.0143026f $X=3.405 $Y=1.765 $X2=0 $Y2=0
cc_254 N_A1_c_238_n N_Y_c_838_n 0.0015992f $X=3.91 $Y=1.765 $X2=0 $Y2=0
cc_255 N_A1_c_233_n N_Y_c_838_n 0.0697975f $X=3.13 $Y=1.515 $X2=0 $Y2=0
cc_256 N_A1_c_234_n N_Y_c_838_n 0.0036203f $X=3.685 $Y=1.485 $X2=0 $Y2=0
cc_257 N_A1_c_235_n N_Y_c_795_n 0.00306874f $X=2.405 $Y=1.765 $X2=0 $Y2=0
cc_258 N_A1_c_231_n N_Y_c_846_n 0.00605027f $X=3.255 $Y=1.205 $X2=0 $Y2=0
cc_259 N_A1_c_232_n N_Y_c_846_n 0.0047069f $X=3.685 $Y=1.205 $X2=0 $Y2=0
cc_260 N_A1_c_234_n N_Y_c_846_n 0.00196781f $X=3.685 $Y=1.485 $X2=0 $Y2=0
cc_261 N_A1_c_236_n Y 8.21497e-19 $X=2.955 $Y=1.765 $X2=0 $Y2=0
cc_262 N_A1_c_237_n Y 0.00506969f $X=3.405 $Y=1.765 $X2=0 $Y2=0
cc_263 N_A1_c_238_n Y 0.00428868f $X=3.91 $Y=1.765 $X2=0 $Y2=0
cc_264 N_A1_c_234_n Y 0.0195821f $X=3.685 $Y=1.485 $X2=0 $Y2=0
cc_265 N_A1_c_231_n N_Y_c_793_n 0.00263107f $X=3.255 $Y=1.205 $X2=0 $Y2=0
cc_266 N_A1_c_232_n N_Y_c_793_n 0.00413936f $X=3.685 $Y=1.205 $X2=0 $Y2=0
cc_267 N_A1_c_233_n N_Y_c_793_n 0.0331256f $X=3.13 $Y=1.515 $X2=0 $Y2=0
cc_268 N_A1_c_234_n N_Y_c_793_n 0.0204398f $X=3.685 $Y=1.485 $X2=0 $Y2=0
cc_269 N_A1_c_235_n N_VPWR_c_899_n 0.00344554f $X=2.405 $Y=1.765 $X2=0 $Y2=0
cc_270 N_A1_c_236_n N_VPWR_c_899_n 0.0053505f $X=2.955 $Y=1.765 $X2=0 $Y2=0
cc_271 N_A1_c_236_n N_VPWR_c_900_n 0.00445602f $X=2.955 $Y=1.765 $X2=0 $Y2=0
cc_272 N_A1_c_237_n N_VPWR_c_900_n 0.00445602f $X=3.405 $Y=1.765 $X2=0 $Y2=0
cc_273 N_A1_c_237_n N_VPWR_c_901_n 0.00417862f $X=3.405 $Y=1.765 $X2=0 $Y2=0
cc_274 N_A1_c_238_n N_VPWR_c_901_n 0.00489307f $X=3.91 $Y=1.765 $X2=0 $Y2=0
cc_275 N_A1_c_238_n N_VPWR_c_902_n 0.00445602f $X=3.91 $Y=1.765 $X2=0 $Y2=0
cc_276 N_A1_c_235_n N_VPWR_c_914_n 0.0044313f $X=2.405 $Y=1.765 $X2=0 $Y2=0
cc_277 N_A1_c_235_n N_VPWR_c_898_n 0.00853652f $X=2.405 $Y=1.765 $X2=0 $Y2=0
cc_278 N_A1_c_236_n N_VPWR_c_898_n 0.00857797f $X=2.955 $Y=1.765 $X2=0 $Y2=0
cc_279 N_A1_c_237_n N_VPWR_c_898_n 0.00858094f $X=3.405 $Y=1.765 $X2=0 $Y2=0
cc_280 N_A1_c_238_n N_VPWR_c_898_n 0.00857618f $X=3.91 $Y=1.765 $X2=0 $Y2=0
cc_281 N_A1_c_227_n N_VGND_c_1044_n 0.00179989f $X=1.985 $Y=1.205 $X2=0 $Y2=0
cc_282 N_A1_c_227_n N_VGND_c_1048_n 0.00278247f $X=1.985 $Y=1.205 $X2=0 $Y2=0
cc_283 N_A1_c_230_n N_VGND_c_1048_n 0.00278271f $X=2.485 $Y=1.205 $X2=0 $Y2=0
cc_284 N_A1_c_231_n N_VGND_c_1048_n 0.00278271f $X=3.255 $Y=1.205 $X2=0 $Y2=0
cc_285 N_A1_c_232_n N_VGND_c_1048_n 0.00278271f $X=3.685 $Y=1.205 $X2=0 $Y2=0
cc_286 N_A1_c_227_n N_VGND_c_1051_n 0.00359084f $X=1.985 $Y=1.205 $X2=0 $Y2=0
cc_287 N_A1_c_230_n N_VGND_c_1051_n 0.00356595f $X=2.485 $Y=1.205 $X2=0 $Y2=0
cc_288 N_A1_c_231_n N_VGND_c_1051_n 0.00355937f $X=3.255 $Y=1.205 $X2=0 $Y2=0
cc_289 N_A1_c_232_n N_VGND_c_1051_n 0.0035414f $X=3.685 $Y=1.205 $X2=0 $Y2=0
cc_290 N_A1_c_227_n N_A_325_74#_c_1141_n 0.00690005f $X=1.985 $Y=1.205 $X2=0
+ $Y2=0
cc_291 N_A1_c_230_n N_A_325_74#_c_1141_n 4.62714e-19 $X=2.485 $Y=1.205 $X2=0
+ $Y2=0
cc_292 N_A1_c_227_n N_A_325_74#_c_1142_n 0.00831967f $X=1.985 $Y=1.205 $X2=0
+ $Y2=0
cc_293 N_A1_c_230_n N_A_325_74#_c_1142_n 0.0136015f $X=2.485 $Y=1.205 $X2=0
+ $Y2=0
cc_294 N_A1_c_227_n N_A_325_74#_c_1143_n 0.00395315f $X=1.985 $Y=1.205 $X2=0
+ $Y2=0
cc_295 N_A1_c_230_n N_A_325_74#_c_1144_n 7.29988e-19 $X=2.485 $Y=1.205 $X2=0
+ $Y2=0
cc_296 N_A1_c_231_n N_A_325_74#_c_1144_n 7.86496e-19 $X=3.255 $Y=1.205 $X2=0
+ $Y2=0
cc_297 N_A1_c_233_n N_A_325_74#_c_1144_n 0.0373748f $X=3.13 $Y=1.515 $X2=0 $Y2=0
cc_298 N_A1_c_234_n N_A_325_74#_c_1144_n 0.0133776f $X=3.685 $Y=1.485 $X2=0
+ $Y2=0
cc_299 N_A1_c_231_n N_A_325_74#_c_1145_n 0.0132525f $X=3.255 $Y=1.205 $X2=0
+ $Y2=0
cc_300 N_A1_c_232_n N_A_325_74#_c_1145_n 0.0133672f $X=3.685 $Y=1.205 $X2=0
+ $Y2=0
cc_301 N_A1_c_232_n N_A_325_74#_c_1148_n 0.00272146f $X=3.685 $Y=1.205 $X2=0
+ $Y2=0
cc_302 N_A1_c_234_n N_A_325_74#_c_1148_n 0.0056439f $X=3.685 $Y=1.485 $X2=0
+ $Y2=0
cc_303 N_A2_c_345_n N_A3_c_432_n 0.00855924f $X=5.82 $Y=1.765 $X2=-0.19
+ $Y2=-0.245
cc_304 N_A2_c_345_n A3 5.49243e-19 $X=5.82 $Y=1.765 $X2=0 $Y2=0
cc_305 N_A2_c_339_n A3 0.018331f $X=5.455 $Y=1.485 $X2=0 $Y2=0
cc_306 N_A2_c_340_n A3 0.010488f $X=5.545 $Y=1.485 $X2=0 $Y2=0
cc_307 N_A2_c_339_n N_A3_c_431_n 2.09661e-19 $X=5.455 $Y=1.485 $X2=0 $Y2=0
cc_308 N_A2_c_340_n N_A3_c_431_n 0.0150065f $X=5.545 $Y=1.485 $X2=0 $Y2=0
cc_309 N_A2_c_342_n N_A_27_368#_c_629_n 4.27055e-19 $X=4.36 $Y=1.765 $X2=0 $Y2=0
cc_310 N_A2_c_340_n N_A_27_368#_c_629_n 4.71954e-19 $X=5.545 $Y=1.485 $X2=0
+ $Y2=0
cc_311 N_A2_c_341_n N_A_27_368#_c_629_n 0.0239058f $X=4.445 $Y=1.55 $X2=0 $Y2=0
cc_312 N_A2_c_342_n N_A_27_368#_c_630_n 0.00327744f $X=4.36 $Y=1.765 $X2=0 $Y2=0
cc_313 N_A2_c_343_n N_A_27_368#_c_630_n 5.16365e-19 $X=4.87 $Y=1.765 $X2=0 $Y2=0
cc_314 N_A2_c_342_n N_A_27_368#_c_595_n 0.0056972f $X=4.36 $Y=1.765 $X2=0 $Y2=0
cc_315 N_A2_c_342_n N_A_27_368#_c_645_n 0.012331f $X=4.36 $Y=1.765 $X2=0 $Y2=0
cc_316 N_A2_c_343_n N_A_27_368#_c_645_n 0.0129915f $X=4.87 $Y=1.765 $X2=0 $Y2=0
cc_317 N_A2_c_339_n N_A_27_368#_c_645_n 0.0104417f $X=5.455 $Y=1.485 $X2=0 $Y2=0
cc_318 N_A2_c_340_n N_A_27_368#_c_645_n 0.0034529f $X=5.545 $Y=1.485 $X2=0 $Y2=0
cc_319 N_A2_c_341_n N_A_27_368#_c_645_n 0.0269797f $X=4.445 $Y=1.55 $X2=0 $Y2=0
cc_320 N_A2_c_342_n N_A_27_368#_c_596_n 6.10709e-19 $X=4.36 $Y=1.765 $X2=0 $Y2=0
cc_321 N_A2_c_343_n N_A_27_368#_c_596_n 0.0109394f $X=4.87 $Y=1.765 $X2=0 $Y2=0
cc_322 N_A2_c_344_n N_A_27_368#_c_596_n 0.0112197f $X=5.32 $Y=1.765 $X2=0 $Y2=0
cc_323 N_A2_c_345_n N_A_27_368#_c_596_n 6.99794e-19 $X=5.82 $Y=1.765 $X2=0 $Y2=0
cc_324 N_A2_c_344_n N_A_27_368#_c_654_n 0.0129411f $X=5.32 $Y=1.765 $X2=0 $Y2=0
cc_325 N_A2_c_345_n N_A_27_368#_c_654_n 0.0159921f $X=5.82 $Y=1.765 $X2=0 $Y2=0
cc_326 N_A2_c_339_n N_A_27_368#_c_654_n 0.0154783f $X=5.455 $Y=1.485 $X2=0 $Y2=0
cc_327 N_A2_c_340_n N_A_27_368#_c_654_n 0.00754244f $X=5.545 $Y=1.485 $X2=0
+ $Y2=0
cc_328 N_A2_c_344_n N_A_27_368#_c_597_n 6.04643e-19 $X=5.32 $Y=1.765 $X2=0 $Y2=0
cc_329 N_A2_c_345_n N_A_27_368#_c_597_n 0.0100488f $X=5.82 $Y=1.765 $X2=0 $Y2=0
cc_330 N_A2_c_342_n N_A_27_368#_c_638_n 0.00175111f $X=4.36 $Y=1.765 $X2=0 $Y2=0
cc_331 N_A2_c_342_n N_A_27_368#_c_605_n 6.0194e-19 $X=4.36 $Y=1.765 $X2=0 $Y2=0
cc_332 N_A2_c_343_n N_A_27_368#_c_605_n 0.00312796f $X=4.87 $Y=1.765 $X2=0 $Y2=0
cc_333 N_A2_c_344_n N_A_27_368#_c_605_n 0.00310836f $X=5.32 $Y=1.765 $X2=0 $Y2=0
cc_334 N_A2_c_345_n N_A_27_368#_c_605_n 6.04745e-19 $X=5.82 $Y=1.765 $X2=0 $Y2=0
cc_335 N_A2_c_339_n N_A_27_368#_c_605_n 0.0276944f $X=5.455 $Y=1.485 $X2=0 $Y2=0
cc_336 N_A2_c_340_n N_A_27_368#_c_605_n 0.0082857f $X=5.545 $Y=1.485 $X2=0 $Y2=0
cc_337 N_A2_c_345_n N_A_27_368#_c_667_n 5.96565e-19 $X=5.82 $Y=1.765 $X2=0 $Y2=0
cc_338 N_A2_c_341_n Y 0.0134646f $X=4.445 $Y=1.55 $X2=0 $Y2=0
cc_339 N_A2_c_335_n N_Y_c_793_n 0.00102246f $X=4.185 $Y=1.205 $X2=0 $Y2=0
cc_340 N_A2_c_341_n N_Y_c_793_n 0.0112767f $X=4.445 $Y=1.55 $X2=0 $Y2=0
cc_341 N_A2_c_342_n N_VPWR_c_902_n 0.00445602f $X=4.36 $Y=1.765 $X2=0 $Y2=0
cc_342 N_A2_c_342_n N_VPWR_c_903_n 0.00535595f $X=4.36 $Y=1.765 $X2=0 $Y2=0
cc_343 N_A2_c_343_n N_VPWR_c_903_n 0.00669982f $X=4.87 $Y=1.765 $X2=0 $Y2=0
cc_344 N_A2_c_343_n N_VPWR_c_904_n 0.00445602f $X=4.87 $Y=1.765 $X2=0 $Y2=0
cc_345 N_A2_c_344_n N_VPWR_c_904_n 0.00445602f $X=5.32 $Y=1.765 $X2=0 $Y2=0
cc_346 N_A2_c_344_n N_VPWR_c_905_n 0.00534288f $X=5.32 $Y=1.765 $X2=0 $Y2=0
cc_347 N_A2_c_345_n N_VPWR_c_905_n 0.00671059f $X=5.82 $Y=1.765 $X2=0 $Y2=0
cc_348 N_A2_c_345_n N_VPWR_c_906_n 0.00445602f $X=5.82 $Y=1.765 $X2=0 $Y2=0
cc_349 N_A2_c_342_n N_VPWR_c_898_n 0.00858221f $X=4.36 $Y=1.765 $X2=0 $Y2=0
cc_350 N_A2_c_343_n N_VPWR_c_898_n 0.00857689f $X=4.87 $Y=1.765 $X2=0 $Y2=0
cc_351 N_A2_c_344_n N_VPWR_c_898_n 0.0085805f $X=5.32 $Y=1.765 $X2=0 $Y2=0
cc_352 N_A2_c_345_n N_VPWR_c_898_n 0.00857462f $X=5.82 $Y=1.765 $X2=0 $Y2=0
cc_353 N_A2_c_335_n N_VGND_c_1048_n 0.00278247f $X=4.185 $Y=1.205 $X2=0 $Y2=0
cc_354 N_A2_c_336_n N_VGND_c_1048_n 0.00278271f $X=4.685 $Y=1.205 $X2=0 $Y2=0
cc_355 N_A2_c_337_n N_VGND_c_1048_n 0.00278271f $X=5.115 $Y=1.205 $X2=0 $Y2=0
cc_356 N_A2_c_338_n N_VGND_c_1048_n 0.00278271f $X=5.545 $Y=1.205 $X2=0 $Y2=0
cc_357 N_A2_c_335_n N_VGND_c_1051_n 0.00354796f $X=4.185 $Y=1.205 $X2=0 $Y2=0
cc_358 N_A2_c_336_n N_VGND_c_1051_n 0.00354087f $X=4.685 $Y=1.205 $X2=0 $Y2=0
cc_359 N_A2_c_337_n N_VGND_c_1051_n 0.00353428f $X=5.115 $Y=1.205 $X2=0 $Y2=0
cc_360 N_A2_c_338_n N_VGND_c_1051_n 0.00358427f $X=5.545 $Y=1.205 $X2=0 $Y2=0
cc_361 N_A2_c_335_n N_A_325_74#_c_1146_n 0.016033f $X=4.185 $Y=1.205 $X2=0 $Y2=0
cc_362 N_A2_c_336_n N_A_325_74#_c_1146_n 0.0144954f $X=4.685 $Y=1.205 $X2=0
+ $Y2=0
cc_363 N_A2_c_337_n N_A_325_74#_c_1146_n 0.0136457f $X=5.115 $Y=1.205 $X2=0
+ $Y2=0
cc_364 N_A2_c_338_n N_A_325_74#_c_1146_n 0.014579f $X=5.545 $Y=1.205 $X2=0 $Y2=0
cc_365 N_A2_c_335_n N_A_325_74#_c_1148_n 0.0106f $X=4.185 $Y=1.205 $X2=0 $Y2=0
cc_366 N_A2_c_336_n N_A_325_74#_c_1148_n 8.0943e-19 $X=4.685 $Y=1.205 $X2=0
+ $Y2=0
cc_367 N_A2_c_341_n N_A_325_74#_c_1148_n 0.0139392f $X=4.445 $Y=1.55 $X2=0 $Y2=0
cc_368 N_A2_c_335_n N_A_852_74#_c_1205_n 0.00183659f $X=4.185 $Y=1.205 $X2=0
+ $Y2=0
cc_369 N_A2_c_336_n N_A_852_74#_c_1205_n 0.013333f $X=4.685 $Y=1.205 $X2=0 $Y2=0
cc_370 N_A2_c_337_n N_A_852_74#_c_1205_n 0.0133316f $X=5.115 $Y=1.205 $X2=0
+ $Y2=0
cc_371 N_A2_c_338_n N_A_852_74#_c_1205_n 0.017437f $X=5.545 $Y=1.205 $X2=0 $Y2=0
cc_372 N_A2_c_340_n N_A_852_74#_c_1205_n 0.0199303f $X=5.545 $Y=1.485 $X2=0
+ $Y2=0
cc_373 N_A2_c_341_n N_A_852_74#_c_1205_n 0.0946862f $X=4.445 $Y=1.55 $X2=0 $Y2=0
cc_374 N_A2_c_338_n N_A_1235_74#_c_1242_n 5.88287e-19 $X=5.545 $Y=1.205 $X2=0
+ $Y2=0
cc_375 N_A3_c_435_n N_A4_c_519_n 0.0227028f $X=7.72 $Y=1.765 $X2=-0.19
+ $Y2=-0.245
cc_376 N_A3_M1036_g N_A4_M1003_g 0.019323f $X=7.825 $Y=0.74 $X2=0 $Y2=0
cc_377 A3 A4 0.0284999f $X=7.835 $Y=1.58 $X2=0 $Y2=0
cc_378 N_A3_c_431_n A4 3.28267e-19 $X=7.72 $Y=1.557 $X2=0 $Y2=0
cc_379 A3 N_A4_c_518_n 0.00399933f $X=7.835 $Y=1.58 $X2=0 $Y2=0
cc_380 N_A3_c_431_n N_A4_c_518_n 0.0222322f $X=7.72 $Y=1.557 $X2=0 $Y2=0
cc_381 N_A3_c_432_n N_A_27_368#_c_597_n 0.0105763f $X=6.27 $Y=1.765 $X2=0 $Y2=0
cc_382 N_A3_c_433_n N_A_27_368#_c_597_n 6.99794e-19 $X=6.77 $Y=1.765 $X2=0 $Y2=0
cc_383 N_A3_c_432_n N_A_27_368#_c_670_n 0.0122806f $X=6.27 $Y=1.765 $X2=0 $Y2=0
cc_384 N_A3_c_433_n N_A_27_368#_c_670_n 0.0122806f $X=6.77 $Y=1.765 $X2=0 $Y2=0
cc_385 A3 N_A_27_368#_c_670_n 0.04337f $X=7.835 $Y=1.58 $X2=0 $Y2=0
cc_386 N_A3_c_431_n N_A_27_368#_c_670_n 0.00157772f $X=7.72 $Y=1.557 $X2=0 $Y2=0
cc_387 N_A3_c_432_n N_A_27_368#_c_598_n 6.04643e-19 $X=6.27 $Y=1.765 $X2=0 $Y2=0
cc_388 N_A3_c_433_n N_A_27_368#_c_598_n 0.0100939f $X=6.77 $Y=1.765 $X2=0 $Y2=0
cc_389 N_A3_c_434_n N_A_27_368#_c_598_n 0.010582f $X=7.22 $Y=1.765 $X2=0 $Y2=0
cc_390 N_A3_c_435_n N_A_27_368#_c_598_n 6.99794e-19 $X=7.72 $Y=1.765 $X2=0 $Y2=0
cc_391 N_A3_c_434_n N_A_27_368#_c_678_n 0.0122806f $X=7.22 $Y=1.765 $X2=0 $Y2=0
cc_392 N_A3_c_435_n N_A_27_368#_c_678_n 0.0122806f $X=7.72 $Y=1.765 $X2=0 $Y2=0
cc_393 A3 N_A_27_368#_c_678_n 0.04337f $X=7.835 $Y=1.58 $X2=0 $Y2=0
cc_394 N_A3_c_431_n N_A_27_368#_c_678_n 0.0015756f $X=7.72 $Y=1.557 $X2=0 $Y2=0
cc_395 N_A3_c_434_n N_A_27_368#_c_599_n 6.04643e-19 $X=7.22 $Y=1.765 $X2=0 $Y2=0
cc_396 N_A3_c_435_n N_A_27_368#_c_599_n 0.0100845f $X=7.72 $Y=1.765 $X2=0 $Y2=0
cc_397 N_A3_c_432_n N_A_27_368#_c_667_n 4.27055e-19 $X=6.27 $Y=1.765 $X2=0 $Y2=0
cc_398 A3 N_A_27_368#_c_667_n 0.023353f $X=7.835 $Y=1.58 $X2=0 $Y2=0
cc_399 N_A3_c_433_n N_A_27_368#_c_686_n 4.27055e-19 $X=6.77 $Y=1.765 $X2=0 $Y2=0
cc_400 N_A3_c_434_n N_A_27_368#_c_686_n 4.27055e-19 $X=7.22 $Y=1.765 $X2=0 $Y2=0
cc_401 A3 N_A_27_368#_c_686_n 0.0237598f $X=7.835 $Y=1.58 $X2=0 $Y2=0
cc_402 N_A3_c_431_n N_A_27_368#_c_686_n 0.00143454f $X=7.72 $Y=1.557 $X2=0 $Y2=0
cc_403 N_A3_c_435_n N_A_27_368#_c_690_n 4.27055e-19 $X=7.72 $Y=1.765 $X2=0 $Y2=0
cc_404 A3 N_A_27_368#_c_690_n 0.0198357f $X=7.835 $Y=1.58 $X2=0 $Y2=0
cc_405 N_A3_c_431_n N_A_27_368#_c_690_n 4.43066e-19 $X=7.72 $Y=1.557 $X2=0 $Y2=0
cc_406 N_A3_c_432_n N_VPWR_c_906_n 0.00445602f $X=6.27 $Y=1.765 $X2=0 $Y2=0
cc_407 N_A3_c_432_n N_VPWR_c_907_n 0.00534288f $X=6.27 $Y=1.765 $X2=0 $Y2=0
cc_408 N_A3_c_433_n N_VPWR_c_907_n 0.00671059f $X=6.77 $Y=1.765 $X2=0 $Y2=0
cc_409 N_A3_c_433_n N_VPWR_c_908_n 0.00445602f $X=6.77 $Y=1.765 $X2=0 $Y2=0
cc_410 N_A3_c_434_n N_VPWR_c_908_n 0.00445602f $X=7.22 $Y=1.765 $X2=0 $Y2=0
cc_411 N_A3_c_434_n N_VPWR_c_909_n 0.00534288f $X=7.22 $Y=1.765 $X2=0 $Y2=0
cc_412 N_A3_c_435_n N_VPWR_c_909_n 0.00540678f $X=7.72 $Y=1.765 $X2=0 $Y2=0
cc_413 N_A3_c_435_n N_VPWR_c_910_n 5.09142e-19 $X=7.72 $Y=1.765 $X2=0 $Y2=0
cc_414 N_A3_c_435_n N_VPWR_c_915_n 0.00445602f $X=7.72 $Y=1.765 $X2=0 $Y2=0
cc_415 N_A3_c_432_n N_VPWR_c_898_n 0.00858134f $X=6.27 $Y=1.765 $X2=0 $Y2=0
cc_416 N_A3_c_433_n N_VPWR_c_898_n 0.00857378f $X=6.77 $Y=1.765 $X2=0 $Y2=0
cc_417 N_A3_c_434_n N_VPWR_c_898_n 0.0085805f $X=7.22 $Y=1.765 $X2=0 $Y2=0
cc_418 N_A3_c_435_n N_VPWR_c_898_n 0.00857893f $X=7.72 $Y=1.765 $X2=0 $Y2=0
cc_419 N_A3_M1036_g N_VGND_c_1045_n 6.35276e-19 $X=7.825 $Y=0.74 $X2=0 $Y2=0
cc_420 N_A3_M1010_g N_VGND_c_1048_n 0.00291649f $X=6.535 $Y=0.74 $X2=0 $Y2=0
cc_421 N_A3_M1024_g N_VGND_c_1048_n 0.00291649f $X=6.965 $Y=0.74 $X2=0 $Y2=0
cc_422 N_A3_M1028_g N_VGND_c_1048_n 0.00291649f $X=7.395 $Y=0.74 $X2=0 $Y2=0
cc_423 N_A3_M1036_g N_VGND_c_1048_n 0.00291649f $X=7.825 $Y=0.74 $X2=0 $Y2=0
cc_424 N_A3_M1010_g N_VGND_c_1051_n 0.0036412f $X=6.535 $Y=0.74 $X2=0 $Y2=0
cc_425 N_A3_M1024_g N_VGND_c_1051_n 0.00359121f $X=6.965 $Y=0.74 $X2=0 $Y2=0
cc_426 N_A3_M1028_g N_VGND_c_1051_n 0.00359121f $X=7.395 $Y=0.74 $X2=0 $Y2=0
cc_427 N_A3_M1036_g N_VGND_c_1051_n 0.00359219f $X=7.825 $Y=0.74 $X2=0 $Y2=0
cc_428 N_A3_M1010_g N_A_325_74#_c_1146_n 0.00326143f $X=6.535 $Y=0.74 $X2=0
+ $Y2=0
cc_429 N_A3_M1028_g N_A_852_74#_c_1204_n 0.00207464f $X=7.395 $Y=0.74 $X2=0
+ $Y2=0
cc_430 N_A3_M1036_g N_A_852_74#_c_1204_n 0.00466497f $X=7.825 $Y=0.74 $X2=0
+ $Y2=0
cc_431 N_A3_c_431_n N_A_852_74#_c_1204_n 0.0022876f $X=7.72 $Y=1.557 $X2=0 $Y2=0
cc_432 N_A3_M1010_g N_A_852_74#_c_1205_n 0.0177225f $X=6.535 $Y=0.74 $X2=0 $Y2=0
cc_433 N_A3_M1024_g N_A_852_74#_c_1205_n 0.0136379f $X=6.965 $Y=0.74 $X2=0 $Y2=0
cc_434 N_A3_M1028_g N_A_852_74#_c_1205_n 0.0118331f $X=7.395 $Y=0.74 $X2=0 $Y2=0
cc_435 A3 N_A_852_74#_c_1205_n 0.125425f $X=7.835 $Y=1.58 $X2=0 $Y2=0
cc_436 N_A3_c_431_n N_A_852_74#_c_1205_n 0.0119159f $X=7.72 $Y=1.557 $X2=0 $Y2=0
cc_437 N_A3_M1010_g N_A_1235_74#_c_1235_n 0.00891446f $X=6.535 $Y=0.74 $X2=0
+ $Y2=0
cc_438 N_A3_M1024_g N_A_1235_74#_c_1235_n 0.0103412f $X=6.965 $Y=0.74 $X2=0
+ $Y2=0
cc_439 N_A3_M1028_g N_A_1235_74#_c_1235_n 0.0102518f $X=7.395 $Y=0.74 $X2=0
+ $Y2=0
cc_440 N_A3_M1036_g N_A_1235_74#_c_1235_n 0.014175f $X=7.825 $Y=0.74 $X2=0 $Y2=0
cc_441 N_A3_M1036_g N_A_1235_74#_c_1238_n 0.0017668f $X=7.825 $Y=0.74 $X2=0
+ $Y2=0
cc_442 A3 N_A_1235_74#_c_1238_n 0.00721346f $X=7.835 $Y=1.58 $X2=0 $Y2=0
cc_443 N_A3_M1010_g N_A_1235_74#_c_1242_n 0.0018597f $X=6.535 $Y=0.74 $X2=0
+ $Y2=0
cc_444 N_A4_c_519_n N_A_27_368#_c_599_n 0.00464047f $X=8.22 $Y=1.765 $X2=0 $Y2=0
cc_445 N_A4_c_519_n N_A_27_368#_c_694_n 0.0192576f $X=8.22 $Y=1.765 $X2=0 $Y2=0
cc_446 N_A4_c_520_n N_A_27_368#_c_694_n 0.0120074f $X=8.67 $Y=1.765 $X2=0 $Y2=0
cc_447 A4 N_A_27_368#_c_694_n 0.0303009f $X=9.755 $Y=1.58 $X2=0 $Y2=0
cc_448 N_A4_c_518_n N_A_27_368#_c_694_n 0.00130859f $X=9.57 $Y=1.557 $X2=0 $Y2=0
cc_449 N_A4_c_519_n N_A_27_368#_c_600_n 6.63853e-19 $X=8.22 $Y=1.765 $X2=0 $Y2=0
cc_450 N_A4_c_520_n N_A_27_368#_c_600_n 0.0104721f $X=8.67 $Y=1.765 $X2=0 $Y2=0
cc_451 N_A4_c_521_n N_A_27_368#_c_600_n 0.0103431f $X=9.12 $Y=1.765 $X2=0 $Y2=0
cc_452 N_A4_c_522_n N_A_27_368#_c_600_n 6.45594e-19 $X=9.57 $Y=1.765 $X2=0 $Y2=0
cc_453 N_A4_c_521_n N_A_27_368#_c_702_n 0.0120074f $X=9.12 $Y=1.765 $X2=0 $Y2=0
cc_454 N_A4_c_522_n N_A_27_368#_c_702_n 0.0120074f $X=9.57 $Y=1.765 $X2=0 $Y2=0
cc_455 A4 N_A_27_368#_c_702_n 0.0393875f $X=9.755 $Y=1.58 $X2=0 $Y2=0
cc_456 N_A4_c_518_n N_A_27_368#_c_702_n 0.00131142f $X=9.57 $Y=1.557 $X2=0 $Y2=0
cc_457 N_A4_c_522_n N_A_27_368#_c_601_n 4.27055e-19 $X=9.57 $Y=1.765 $X2=0 $Y2=0
cc_458 A4 N_A_27_368#_c_601_n 0.0260502f $X=9.755 $Y=1.58 $X2=0 $Y2=0
cc_459 N_A4_c_521_n N_A_27_368#_c_602_n 6.45594e-19 $X=9.12 $Y=1.765 $X2=0 $Y2=0
cc_460 N_A4_c_522_n N_A_27_368#_c_602_n 0.0104891f $X=9.57 $Y=1.765 $X2=0 $Y2=0
cc_461 N_A4_c_520_n N_A_27_368#_c_710_n 4.27055e-19 $X=8.67 $Y=1.765 $X2=0 $Y2=0
cc_462 N_A4_c_521_n N_A_27_368#_c_710_n 4.27055e-19 $X=9.12 $Y=1.765 $X2=0 $Y2=0
cc_463 A4 N_A_27_368#_c_710_n 0.0237598f $X=9.755 $Y=1.58 $X2=0 $Y2=0
cc_464 N_A4_c_518_n N_A_27_368#_c_710_n 0.00144162f $X=9.57 $Y=1.557 $X2=0 $Y2=0
cc_465 N_A4_c_519_n N_VPWR_c_910_n 0.0103564f $X=8.22 $Y=1.765 $X2=0 $Y2=0
cc_466 N_A4_c_520_n N_VPWR_c_910_n 0.00526215f $X=8.67 $Y=1.765 $X2=0 $Y2=0
cc_467 N_A4_c_521_n N_VPWR_c_911_n 0.00486623f $X=9.12 $Y=1.765 $X2=0 $Y2=0
cc_468 N_A4_c_522_n N_VPWR_c_911_n 0.00486623f $X=9.57 $Y=1.765 $X2=0 $Y2=0
cc_469 N_A4_c_520_n N_VPWR_c_912_n 0.00445602f $X=8.67 $Y=1.765 $X2=0 $Y2=0
cc_470 N_A4_c_521_n N_VPWR_c_912_n 0.00445602f $X=9.12 $Y=1.765 $X2=0 $Y2=0
cc_471 N_A4_c_519_n N_VPWR_c_915_n 0.00413917f $X=8.22 $Y=1.765 $X2=0 $Y2=0
cc_472 N_A4_c_522_n N_VPWR_c_916_n 0.00445602f $X=9.57 $Y=1.765 $X2=0 $Y2=0
cc_473 N_A4_c_519_n N_VPWR_c_898_n 0.00818241f $X=8.22 $Y=1.765 $X2=0 $Y2=0
cc_474 N_A4_c_520_n N_VPWR_c_898_n 0.00857589f $X=8.67 $Y=1.765 $X2=0 $Y2=0
cc_475 N_A4_c_521_n N_VPWR_c_898_n 0.00857589f $X=9.12 $Y=1.765 $X2=0 $Y2=0
cc_476 N_A4_c_522_n N_VPWR_c_898_n 0.008611f $X=9.57 $Y=1.765 $X2=0 $Y2=0
cc_477 N_A4_M1003_g N_VGND_c_1045_n 0.010782f $X=8.255 $Y=0.74 $X2=0 $Y2=0
cc_478 N_A4_M1017_g N_VGND_c_1045_n 0.0106755f $X=8.685 $Y=0.74 $X2=0 $Y2=0
cc_479 N_A4_M1022_g N_VGND_c_1045_n 4.71636e-19 $X=9.115 $Y=0.74 $X2=0 $Y2=0
cc_480 N_A4_M1017_g N_VGND_c_1046_n 4.71636e-19 $X=8.685 $Y=0.74 $X2=0 $Y2=0
cc_481 N_A4_M1022_g N_VGND_c_1046_n 0.0105384f $X=9.115 $Y=0.74 $X2=0 $Y2=0
cc_482 N_A4_M1034_g N_VGND_c_1046_n 0.00392488f $X=9.585 $Y=0.74 $X2=0 $Y2=0
cc_483 N_A4_M1003_g N_VGND_c_1048_n 0.00383152f $X=8.255 $Y=0.74 $X2=0 $Y2=0
cc_484 N_A4_M1017_g N_VGND_c_1049_n 0.00383152f $X=8.685 $Y=0.74 $X2=0 $Y2=0
cc_485 N_A4_M1022_g N_VGND_c_1049_n 0.00383152f $X=9.115 $Y=0.74 $X2=0 $Y2=0
cc_486 N_A4_M1034_g N_VGND_c_1050_n 0.00461464f $X=9.585 $Y=0.74 $X2=0 $Y2=0
cc_487 N_A4_M1003_g N_VGND_c_1051_n 0.00757637f $X=8.255 $Y=0.74 $X2=0 $Y2=0
cc_488 N_A4_M1017_g N_VGND_c_1051_n 0.0075754f $X=8.685 $Y=0.74 $X2=0 $Y2=0
cc_489 N_A4_M1022_g N_VGND_c_1051_n 0.0075754f $X=9.115 $Y=0.74 $X2=0 $Y2=0
cc_490 N_A4_M1034_g N_VGND_c_1051_n 0.00911481f $X=9.585 $Y=0.74 $X2=0 $Y2=0
cc_491 N_A4_M1003_g N_A_1235_74#_c_1237_n 0.0161035f $X=8.255 $Y=0.74 $X2=0
+ $Y2=0
cc_492 N_A4_M1017_g N_A_1235_74#_c_1237_n 0.0130453f $X=8.685 $Y=0.74 $X2=0
+ $Y2=0
cc_493 A4 N_A_1235_74#_c_1237_n 0.0398909f $X=9.755 $Y=1.58 $X2=0 $Y2=0
cc_494 N_A4_c_518_n N_A_1235_74#_c_1237_n 0.00427455f $X=9.57 $Y=1.557 $X2=0
+ $Y2=0
cc_495 N_A4_M1017_g N_A_1235_74#_c_1239_n 3.92313e-19 $X=8.685 $Y=0.74 $X2=0
+ $Y2=0
cc_496 N_A4_M1022_g N_A_1235_74#_c_1239_n 3.92313e-19 $X=9.115 $Y=0.74 $X2=0
+ $Y2=0
cc_497 N_A4_M1022_g N_A_1235_74#_c_1240_n 0.0133256f $X=9.115 $Y=0.74 $X2=0
+ $Y2=0
cc_498 N_A4_M1034_g N_A_1235_74#_c_1240_n 0.0146212f $X=9.585 $Y=0.74 $X2=0
+ $Y2=0
cc_499 A4 N_A_1235_74#_c_1240_n 0.0766773f $X=9.755 $Y=1.58 $X2=0 $Y2=0
cc_500 N_A4_c_518_n N_A_1235_74#_c_1240_n 0.00313888f $X=9.57 $Y=1.557 $X2=0
+ $Y2=0
cc_501 N_A4_M1034_g N_A_1235_74#_c_1241_n 0.00160529f $X=9.585 $Y=0.74 $X2=0
+ $Y2=0
cc_502 A4 N_A_1235_74#_c_1243_n 0.0146029f $X=9.755 $Y=1.58 $X2=0 $Y2=0
cc_503 N_A4_c_518_n N_A_1235_74#_c_1243_n 0.00232957f $X=9.57 $Y=1.557 $X2=0
+ $Y2=0
cc_504 N_A_27_368#_c_592_n N_Y_M1014_d 0.00245557f $X=1.115 $Y=2.99 $X2=0 $Y2=0
cc_505 N_A_27_368#_c_594_n N_Y_M1019_d 0.00243452f $X=2.015 $Y=2.99 $X2=0 $Y2=0
cc_506 N_A_27_368#_c_612_n N_Y_c_806_n 0.0289859f $X=1.28 $Y=2.405 $X2=0 $Y2=0
cc_507 N_A_27_368#_c_594_n N_Y_c_806_n 0.0126885f $X=2.015 $Y=2.99 $X2=0 $Y2=0
cc_508 N_A_27_368#_c_616_n N_Y_c_806_n 0.0117758f $X=2.18 $Y=2.46 $X2=0 $Y2=0
cc_509 N_A_27_368#_c_617_n N_Y_c_806_n 0.0178797f $X=2.18 $Y=2.905 $X2=0 $Y2=0
cc_510 N_A_27_368#_M1023_s N_Y_c_838_n 0.00456372f $X=2.03 $Y=1.84 $X2=0 $Y2=0
cc_511 N_A_27_368#_M1020_d N_Y_c_838_n 0.00355329f $X=3.03 $Y=1.84 $X2=0 $Y2=0
cc_512 N_A_27_368#_c_624_n N_Y_c_838_n 0.039006f $X=3.015 $Y=2.375 $X2=0 $Y2=0
cc_513 N_A_27_368#_c_626_n N_Y_c_838_n 0.0235117f $X=3.97 $Y=2.375 $X2=0 $Y2=0
cc_514 N_A_27_368#_c_629_n N_Y_c_838_n 0.0108534f $X=4.135 $Y=2.12 $X2=0 $Y2=0
cc_515 N_A_27_368#_c_604_n N_Y_c_838_n 0.0173542f $X=3.18 $Y=2.375 $X2=0 $Y2=0
cc_516 N_A_27_368#_c_592_n N_Y_c_814_n 0.0185424f $X=1.115 $Y=2.99 $X2=0 $Y2=0
cc_517 N_A_27_368#_M1018_s N_Y_c_818_n 0.00453144f $X=1.08 $Y=1.84 $X2=0 $Y2=0
cc_518 N_A_27_368#_c_612_n N_Y_c_818_n 0.0202249f $X=1.28 $Y=2.405 $X2=0 $Y2=0
cc_519 N_A_27_368#_M1023_s N_Y_c_795_n 0.00169183f $X=2.03 $Y=1.84 $X2=0 $Y2=0
cc_520 N_A_27_368#_c_616_n N_Y_c_795_n 0.017402f $X=2.18 $Y=2.46 $X2=0 $Y2=0
cc_521 N_A_27_368#_c_624_n N_VPWR_M1012_s 0.00615777f $X=3.015 $Y=2.375
+ $X2=-0.19 $Y2=1.66
cc_522 N_A_27_368#_c_626_n N_VPWR_M1025_s 0.00551389f $X=3.97 $Y=2.375 $X2=0
+ $Y2=0
cc_523 N_A_27_368#_c_645_n N_VPWR_M1000_d 0.00517295f $X=4.93 $Y=2.035 $X2=0
+ $Y2=0
cc_524 N_A_27_368#_c_654_n N_VPWR_M1015_d 0.00549892f $X=5.88 $Y=2.035 $X2=0
+ $Y2=0
cc_525 N_A_27_368#_c_670_n N_VPWR_M1002_s 0.00480741f $X=6.83 $Y=2.035 $X2=0
+ $Y2=0
cc_526 N_A_27_368#_c_678_n N_VPWR_M1008_s 0.00480741f $X=7.78 $Y=2.035 $X2=0
+ $Y2=0
cc_527 N_A_27_368#_c_694_n N_VPWR_M1005_d 0.00384138f $X=8.73 $Y=2.035 $X2=0
+ $Y2=0
cc_528 N_A_27_368#_c_702_n N_VPWR_M1013_d 0.00408911f $X=9.63 $Y=2.035 $X2=0
+ $Y2=0
cc_529 N_A_27_368#_c_594_n N_VPWR_c_899_n 0.0119239f $X=2.015 $Y=2.99 $X2=0
+ $Y2=0
cc_530 N_A_27_368#_c_624_n N_VPWR_c_899_n 0.0232685f $X=3.015 $Y=2.375 $X2=0
+ $Y2=0
cc_531 N_A_27_368#_c_604_n N_VPWR_c_899_n 0.0139233f $X=3.18 $Y=2.375 $X2=0
+ $Y2=0
cc_532 N_A_27_368#_c_604_n N_VPWR_c_900_n 0.0145674f $X=3.18 $Y=2.375 $X2=0
+ $Y2=0
cc_533 N_A_27_368#_c_626_n N_VPWR_c_901_n 0.0188752f $X=3.97 $Y=2.375 $X2=0
+ $Y2=0
cc_534 N_A_27_368#_c_595_n N_VPWR_c_901_n 0.0135735f $X=4.135 $Y=2.815 $X2=0
+ $Y2=0
cc_535 N_A_27_368#_c_604_n N_VPWR_c_901_n 0.0234974f $X=3.18 $Y=2.375 $X2=0
+ $Y2=0
cc_536 N_A_27_368#_c_595_n N_VPWR_c_902_n 0.014552f $X=4.135 $Y=2.815 $X2=0
+ $Y2=0
cc_537 N_A_27_368#_c_595_n N_VPWR_c_903_n 0.0348632f $X=4.135 $Y=2.815 $X2=0
+ $Y2=0
cc_538 N_A_27_368#_c_645_n N_VPWR_c_903_n 0.019282f $X=4.93 $Y=2.035 $X2=0 $Y2=0
cc_539 N_A_27_368#_c_596_n N_VPWR_c_903_n 0.0254585f $X=5.095 $Y=2.815 $X2=0
+ $Y2=0
cc_540 N_A_27_368#_c_638_n N_VPWR_c_903_n 0.0121024f $X=4.135 $Y=2.375 $X2=0
+ $Y2=0
cc_541 N_A_27_368#_c_596_n N_VPWR_c_904_n 0.014552f $X=5.095 $Y=2.815 $X2=0
+ $Y2=0
cc_542 N_A_27_368#_c_596_n N_VPWR_c_905_n 0.0462948f $X=5.095 $Y=2.815 $X2=0
+ $Y2=0
cc_543 N_A_27_368#_c_654_n N_VPWR_c_905_n 0.0184684f $X=5.88 $Y=2.035 $X2=0
+ $Y2=0
cc_544 N_A_27_368#_c_597_n N_VPWR_c_905_n 0.0266484f $X=6.045 $Y=2.815 $X2=0
+ $Y2=0
cc_545 N_A_27_368#_c_597_n N_VPWR_c_906_n 0.014552f $X=6.045 $Y=2.815 $X2=0
+ $Y2=0
cc_546 N_A_27_368#_c_597_n N_VPWR_c_907_n 0.0462948f $X=6.045 $Y=2.815 $X2=0
+ $Y2=0
cc_547 N_A_27_368#_c_670_n N_VPWR_c_907_n 0.0184684f $X=6.83 $Y=2.035 $X2=0
+ $Y2=0
cc_548 N_A_27_368#_c_598_n N_VPWR_c_907_n 0.0266484f $X=6.995 $Y=2.815 $X2=0
+ $Y2=0
cc_549 N_A_27_368#_c_598_n N_VPWR_c_908_n 0.014552f $X=6.995 $Y=2.815 $X2=0
+ $Y2=0
cc_550 N_A_27_368#_c_598_n N_VPWR_c_909_n 0.0462948f $X=6.995 $Y=2.815 $X2=0
+ $Y2=0
cc_551 N_A_27_368#_c_678_n N_VPWR_c_909_n 0.0184684f $X=7.78 $Y=2.035 $X2=0
+ $Y2=0
cc_552 N_A_27_368#_c_599_n N_VPWR_c_909_n 0.0266484f $X=7.945 $Y=2.425 $X2=0
+ $Y2=0
cc_553 N_A_27_368#_c_599_n N_VPWR_c_910_n 0.0256025f $X=7.945 $Y=2.425 $X2=0
+ $Y2=0
cc_554 N_A_27_368#_c_694_n N_VPWR_c_910_n 0.0154248f $X=8.73 $Y=2.035 $X2=0
+ $Y2=0
cc_555 N_A_27_368#_c_600_n N_VPWR_c_910_n 0.0462948f $X=8.895 $Y=2.815 $X2=0
+ $Y2=0
cc_556 N_A_27_368#_c_600_n N_VPWR_c_911_n 0.0449718f $X=8.895 $Y=2.815 $X2=0
+ $Y2=0
cc_557 N_A_27_368#_c_702_n N_VPWR_c_911_n 0.0136682f $X=9.63 $Y=2.035 $X2=0
+ $Y2=0
cc_558 N_A_27_368#_c_602_n N_VPWR_c_911_n 0.0449718f $X=9.795 $Y=2.815 $X2=0
+ $Y2=0
cc_559 N_A_27_368#_c_600_n N_VPWR_c_912_n 0.014552f $X=8.895 $Y=2.815 $X2=0
+ $Y2=0
cc_560 N_A_27_368#_c_592_n N_VPWR_c_914_n 0.0422607f $X=1.115 $Y=2.99 $X2=0
+ $Y2=0
cc_561 N_A_27_368#_c_593_n N_VPWR_c_914_n 0.0236215f $X=0.445 $Y=2.99 $X2=0
+ $Y2=0
cc_562 N_A_27_368#_c_594_n N_VPWR_c_914_n 0.0594312f $X=2.015 $Y=2.99 $X2=0
+ $Y2=0
cc_563 N_A_27_368#_c_603_n N_VPWR_c_914_n 0.0236039f $X=1.28 $Y=2.99 $X2=0 $Y2=0
cc_564 N_A_27_368#_c_599_n N_VPWR_c_915_n 0.0145938f $X=7.945 $Y=2.425 $X2=0
+ $Y2=0
cc_565 N_A_27_368#_c_602_n N_VPWR_c_916_n 0.0145938f $X=9.795 $Y=2.815 $X2=0
+ $Y2=0
cc_566 N_A_27_368#_c_592_n N_VPWR_c_898_n 0.0238634f $X=1.115 $Y=2.99 $X2=0
+ $Y2=0
cc_567 N_A_27_368#_c_593_n N_VPWR_c_898_n 0.0127839f $X=0.445 $Y=2.99 $X2=0
+ $Y2=0
cc_568 N_A_27_368#_c_594_n N_VPWR_c_898_n 0.0328875f $X=2.015 $Y=2.99 $X2=0
+ $Y2=0
cc_569 N_A_27_368#_c_595_n N_VPWR_c_898_n 0.0119791f $X=4.135 $Y=2.815 $X2=0
+ $Y2=0
cc_570 N_A_27_368#_c_596_n N_VPWR_c_898_n 0.0119791f $X=5.095 $Y=2.815 $X2=0
+ $Y2=0
cc_571 N_A_27_368#_c_597_n N_VPWR_c_898_n 0.0119791f $X=6.045 $Y=2.815 $X2=0
+ $Y2=0
cc_572 N_A_27_368#_c_598_n N_VPWR_c_898_n 0.0119791f $X=6.995 $Y=2.815 $X2=0
+ $Y2=0
cc_573 N_A_27_368#_c_599_n N_VPWR_c_898_n 0.0120466f $X=7.945 $Y=2.425 $X2=0
+ $Y2=0
cc_574 N_A_27_368#_c_600_n N_VPWR_c_898_n 0.0119791f $X=8.895 $Y=2.815 $X2=0
+ $Y2=0
cc_575 N_A_27_368#_c_602_n N_VPWR_c_898_n 0.0120466f $X=9.795 $Y=2.815 $X2=0
+ $Y2=0
cc_576 N_A_27_368#_c_603_n N_VPWR_c_898_n 0.012761f $X=1.28 $Y=2.99 $X2=0 $Y2=0
cc_577 N_A_27_368#_c_604_n N_VPWR_c_898_n 0.0119851f $X=3.18 $Y=2.375 $X2=0
+ $Y2=0
cc_578 N_Y_c_838_n N_VPWR_M1012_s 0.00584303f $X=3.465 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_579 N_Y_c_838_n N_VPWR_M1025_s 0.00416285f $X=3.465 $Y=2.035 $X2=0 $Y2=0
cc_580 Y N_VPWR_M1025_s 0.00134133f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_581 N_Y_c_789_n N_VGND_M1035_d 0.00299905f $X=1.815 $Y=1.095 $X2=0 $Y2=0
cc_582 N_Y_c_788_n N_VGND_c_1043_n 0.0243474f $X=0.71 $Y=0.515 $X2=0 $Y2=0
cc_583 N_Y_c_790_n N_VGND_c_1043_n 0.00555794f $X=0.875 $Y=1.095 $X2=0 $Y2=0
cc_584 N_Y_c_788_n N_VGND_c_1044_n 0.0191765f $X=0.71 $Y=0.515 $X2=0 $Y2=0
cc_585 N_Y_c_789_n N_VGND_c_1044_n 0.0219406f $X=1.815 $Y=1.095 $X2=0 $Y2=0
cc_586 N_Y_c_788_n N_VGND_c_1047_n 0.0145639f $X=0.71 $Y=0.515 $X2=0 $Y2=0
cc_587 N_Y_c_788_n N_VGND_c_1051_n 0.0119984f $X=0.71 $Y=0.515 $X2=0 $Y2=0
cc_588 N_Y_c_789_n N_A_325_74#_M1027_s 0.00258447f $X=1.815 $Y=1.095 $X2=-0.19
+ $Y2=-0.245
cc_589 N_Y_c_792_n N_A_325_74#_M1027_s 4.03947e-19 $X=2.27 $Y=1.01 $X2=-0.19
+ $Y2=-0.245
cc_590 N_Y_c_789_n N_A_325_74#_c_1141_n 0.0216365f $X=1.815 $Y=1.095 $X2=0 $Y2=0
cc_591 N_Y_M1027_d N_A_325_74#_c_1142_n 0.00250873f $X=2.06 $Y=0.37 $X2=0 $Y2=0
cc_592 N_Y_c_792_n N_A_325_74#_c_1142_n 0.00306797f $X=2.27 $Y=1.01 $X2=0 $Y2=0
cc_593 N_Y_c_837_n N_A_325_74#_c_1142_n 0.018913f $X=2.27 $Y=0.76 $X2=0 $Y2=0
cc_594 N_Y_c_792_n N_A_325_74#_c_1144_n 0.00586549f $X=2.27 $Y=1.01 $X2=0 $Y2=0
cc_595 N_Y_c_793_n N_A_325_74#_c_1144_n 0.00343886f $X=3.59 $Y=1.55 $X2=0 $Y2=0
cc_596 N_Y_M1032_d N_A_325_74#_c_1145_n 0.00176461f $X=3.33 $Y=0.37 $X2=0 $Y2=0
cc_597 N_Y_c_846_n N_A_325_74#_c_1145_n 0.0156869f $X=3.47 $Y=0.785 $X2=0 $Y2=0
cc_598 N_Y_c_846_n N_A_325_74#_c_1148_n 0.0194208f $X=3.47 $Y=0.785 $X2=0 $Y2=0
cc_599 N_VGND_c_1044_n N_A_325_74#_c_1141_n 0.027945f $X=1.21 $Y=0.675 $X2=0
+ $Y2=0
cc_600 N_VGND_c_1048_n N_A_325_74#_c_1142_n 0.0423044f $X=8.305 $Y=0 $X2=0 $Y2=0
cc_601 N_VGND_c_1051_n N_A_325_74#_c_1142_n 0.0239316f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_602 N_VGND_c_1044_n N_A_325_74#_c_1143_n 0.0121616f $X=1.21 $Y=0.675 $X2=0
+ $Y2=0
cc_603 N_VGND_c_1048_n N_A_325_74#_c_1143_n 0.0233048f $X=8.305 $Y=0 $X2=0 $Y2=0
cc_604 N_VGND_c_1051_n N_A_325_74#_c_1143_n 0.0126653f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_605 N_VGND_c_1048_n N_A_325_74#_c_1145_n 0.0422287f $X=8.305 $Y=0 $X2=0 $Y2=0
cc_606 N_VGND_c_1051_n N_A_325_74#_c_1145_n 0.0238173f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_607 N_VGND_c_1048_n N_A_325_74#_c_1146_n 0.119831f $X=8.305 $Y=0 $X2=0 $Y2=0
cc_608 N_VGND_c_1051_n N_A_325_74#_c_1146_n 0.0658365f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_609 N_VGND_c_1048_n N_A_325_74#_c_1147_n 0.037994f $X=8.305 $Y=0 $X2=0 $Y2=0
cc_610 N_VGND_c_1051_n N_A_325_74#_c_1147_n 0.0206052f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_611 N_VGND_c_1048_n N_A_325_74#_c_1148_n 0.0235688f $X=8.305 $Y=0 $X2=0 $Y2=0
cc_612 N_VGND_c_1051_n N_A_325_74#_c_1148_n 0.0127152f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_613 N_VGND_c_1051_n N_A_852_74#_c_1205_n 0.0137814f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_614 N_VGND_c_1045_n N_A_1235_74#_c_1236_n 0.00985092f $X=8.47 $Y=0.675 $X2=0
+ $Y2=0
cc_615 N_VGND_c_1048_n N_A_1235_74#_c_1236_n 0.00758556f $X=8.305 $Y=0 $X2=0
+ $Y2=0
cc_616 N_VGND_c_1051_n N_A_1235_74#_c_1236_n 0.00627867f $X=9.84 $Y=0 $X2=0
+ $Y2=0
cc_617 N_VGND_M1003_s N_A_1235_74#_c_1237_n 0.00176461f $X=8.33 $Y=0.37 $X2=0
+ $Y2=0
cc_618 N_VGND_c_1045_n N_A_1235_74#_c_1237_n 0.0170777f $X=8.47 $Y=0.675 $X2=0
+ $Y2=0
cc_619 N_VGND_c_1045_n N_A_1235_74#_c_1239_n 0.0182488f $X=8.47 $Y=0.675 $X2=0
+ $Y2=0
cc_620 N_VGND_c_1046_n N_A_1235_74#_c_1239_n 0.0182488f $X=9.33 $Y=0.675 $X2=0
+ $Y2=0
cc_621 N_VGND_c_1049_n N_A_1235_74#_c_1239_n 0.00749631f $X=9.165 $Y=0 $X2=0
+ $Y2=0
cc_622 N_VGND_c_1051_n N_A_1235_74#_c_1239_n 0.0062048f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_623 N_VGND_M1022_s N_A_1235_74#_c_1240_n 0.00218982f $X=9.19 $Y=0.37 $X2=0
+ $Y2=0
cc_624 N_VGND_c_1046_n N_A_1235_74#_c_1240_n 0.0185459f $X=9.33 $Y=0.675 $X2=0
+ $Y2=0
cc_625 N_VGND_c_1046_n N_A_1235_74#_c_1241_n 0.00129215f $X=9.33 $Y=0.675 $X2=0
+ $Y2=0
cc_626 N_VGND_c_1050_n N_A_1235_74#_c_1241_n 0.011066f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_627 N_VGND_c_1051_n N_A_1235_74#_c_1241_n 0.00915947f $X=9.84 $Y=0 $X2=0
+ $Y2=0
cc_628 N_VGND_c_1048_n N_A_1235_74#_c_1242_n 0.0730035f $X=8.305 $Y=0 $X2=0
+ $Y2=0
cc_629 N_VGND_c_1051_n N_A_1235_74#_c_1242_n 0.0614975f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_630 N_A_325_74#_c_1146_n N_A_852_74#_M1006_d 0.00240933f $X=5.76 $Y=0.515
+ $X2=-0.19 $Y2=-0.245
cc_631 N_A_325_74#_c_1146_n N_A_852_74#_M1030_d 0.00171374f $X=5.76 $Y=0.515
+ $X2=0 $Y2=0
cc_632 N_A_325_74#_M1007_s N_A_852_74#_c_1205_n 0.0017749f $X=4.76 $Y=0.37 $X2=0
+ $Y2=0
cc_633 N_A_325_74#_M1033_s N_A_852_74#_c_1205_n 0.00429177f $X=5.62 $Y=0.37
+ $X2=0 $Y2=0
cc_634 N_A_325_74#_c_1146_n N_A_852_74#_c_1205_n 0.0970525f $X=5.76 $Y=0.515
+ $X2=0 $Y2=0
cc_635 N_A_325_74#_c_1148_n N_A_852_74#_c_1205_n 0.0135819f $X=3.97 $Y=0.515
+ $X2=0 $Y2=0
cc_636 N_A_325_74#_c_1146_n N_A_1235_74#_c_1242_n 0.0202095f $X=5.76 $Y=0.515
+ $X2=0 $Y2=0
cc_637 N_A_852_74#_c_1205_n N_A_1235_74#_M1010_d 0.00429177f $X=7.445 $Y=0.95
+ $X2=-0.19 $Y2=-0.245
cc_638 N_A_852_74#_c_1205_n N_A_1235_74#_M1024_d 0.00185845f $X=7.445 $Y=0.95
+ $X2=0 $Y2=0
cc_639 N_A_852_74#_M1010_s N_A_1235_74#_c_1235_n 0.00187648f $X=6.61 $Y=0.37
+ $X2=0 $Y2=0
cc_640 N_A_852_74#_M1028_s N_A_1235_74#_c_1235_n 0.00179007f $X=7.47 $Y=0.37
+ $X2=0 $Y2=0
cc_641 N_A_852_74#_c_1204_n N_A_1235_74#_c_1235_n 0.016201f $X=7.61 $Y=0.95
+ $X2=0 $Y2=0
cc_642 N_A_852_74#_c_1205_n N_A_1235_74#_c_1235_n 0.0487326f $X=7.445 $Y=0.95
+ $X2=0 $Y2=0
cc_643 N_A_852_74#_c_1204_n N_A_1235_74#_c_1238_n 0.00561736f $X=7.61 $Y=0.95
+ $X2=0 $Y2=0
cc_644 N_A_852_74#_c_1205_n N_A_1235_74#_c_1242_n 0.0208608f $X=7.445 $Y=0.95
+ $X2=0 $Y2=0
