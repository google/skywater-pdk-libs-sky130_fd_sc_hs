* File: sky130_fd_sc_hs__a211o_1.pxi.spice
* Created: Thu Aug 27 20:23:14 2020
* 
x_PM_SKY130_FD_SC_HS__A211O_1%A_81_264# N_A_81_264#_M1009_d N_A_81_264#_M1006_d
+ N_A_81_264#_M1007_d N_A_81_264#_c_71_n N_A_81_264#_M1000_g N_A_81_264#_M1004_g
+ N_A_81_264#_c_65_n N_A_81_264#_c_66_n N_A_81_264#_c_112_p N_A_81_264#_c_67_n
+ N_A_81_264#_c_88_p N_A_81_264#_c_68_n N_A_81_264#_c_69_n N_A_81_264#_c_70_n
+ N_A_81_264#_c_80_p PM_SKY130_FD_SC_HS__A211O_1%A_81_264#
x_PM_SKY130_FD_SC_HS__A211O_1%A2 N_A2_c_144_n N_A2_M1002_g N_A2_M1008_g A2
+ PM_SKY130_FD_SC_HS__A211O_1%A2
x_PM_SKY130_FD_SC_HS__A211O_1%A1 N_A1_c_176_n N_A1_M1001_g N_A1_M1009_g A1 A1
+ PM_SKY130_FD_SC_HS__A211O_1%A1
x_PM_SKY130_FD_SC_HS__A211O_1%B1 N_B1_M1005_g N_B1_c_216_n N_B1_c_217_n
+ N_B1_c_222_n N_B1_M1003_g N_B1_c_218_n N_B1_c_219_n B1 N_B1_c_220_n
+ PM_SKY130_FD_SC_HS__A211O_1%B1
x_PM_SKY130_FD_SC_HS__A211O_1%C1 N_C1_c_262_n N_C1_c_269_n N_C1_M1007_g
+ N_C1_M1006_g N_C1_c_264_n N_C1_c_265_n C1 N_C1_c_266_n N_C1_c_267_n
+ PM_SKY130_FD_SC_HS__A211O_1%C1
x_PM_SKY130_FD_SC_HS__A211O_1%X N_X_M1004_s N_X_M1000_s N_X_c_300_n X X X X
+ N_X_c_301_n PM_SKY130_FD_SC_HS__A211O_1%X
x_PM_SKY130_FD_SC_HS__A211O_1%VPWR N_VPWR_M1000_d N_VPWR_M1002_d N_VPWR_c_322_n
+ N_VPWR_c_323_n N_VPWR_c_324_n N_VPWR_c_325_n VPWR N_VPWR_c_326_n
+ N_VPWR_c_327_n N_VPWR_c_321_n N_VPWR_c_329_n PM_SKY130_FD_SC_HS__A211O_1%VPWR
x_PM_SKY130_FD_SC_HS__A211O_1%A_279_392# N_A_279_392#_M1002_s
+ N_A_279_392#_M1001_d N_A_279_392#_c_360_n N_A_279_392#_c_361_n
+ N_A_279_392#_c_362_n N_A_279_392#_c_363_n N_A_279_392#_c_364_n
+ PM_SKY130_FD_SC_HS__A211O_1%A_279_392#
x_PM_SKY130_FD_SC_HS__A211O_1%VGND N_VGND_M1004_d N_VGND_M1005_d N_VGND_c_396_n
+ N_VGND_c_397_n N_VGND_c_398_n N_VGND_c_411_n VGND N_VGND_c_399_n
+ N_VGND_c_400_n N_VGND_c_401_n N_VGND_c_402_n N_VGND_c_403_n
+ PM_SKY130_FD_SC_HS__A211O_1%VGND
cc_1 VNB N_A_81_264#_M1004_g 0.0324185f $X=-0.19 $Y=-0.245 $X2=1.205 $Y2=0.74
cc_2 VNB N_A_81_264#_c_65_n 0.0204685f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.485
cc_3 VNB N_A_81_264#_c_66_n 0.0718582f $X=-0.19 $Y=-0.245 $X2=1.13 $Y2=1.485
cc_4 VNB N_A_81_264#_c_67_n 7.10275e-19 $X=-0.19 $Y=-0.245 $X2=2.28 $Y2=1.195
cc_5 VNB N_A_81_264#_c_68_n 0.00884873f $X=-0.19 $Y=-0.245 $X2=3.332 $Y2=1.28
cc_6 VNB N_A_81_264#_c_69_n 0.0161422f $X=-0.19 $Y=-0.245 $X2=3.29 $Y2=2.105
cc_7 VNB N_A_81_264#_c_70_n 0.00827298f $X=-0.19 $Y=-0.245 $X2=1.33 $Y2=1.195
cc_8 VNB N_A2_c_144_n 0.019391f $X=-0.19 $Y=-0.245 $X2=2.305 $Y2=0.68
cc_9 VNB N_A2_M1008_g 0.0194469f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB A2 8.71858e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A1_c_176_n 0.0159842f $X=-0.19 $Y=-0.245 $X2=2.305 $Y2=0.68
cc_12 VNB N_A1_M1009_g 0.0178919f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB A1 0.00334688f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_B1_M1005_g 0.0103467f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_B1_c_216_n 0.00535021f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_B1_c_217_n 0.00795002f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_B1_c_218_n 0.00691726f $X=-0.19 $Y=-0.245 $X2=1.205 $Y2=1.32
cc_18 VNB N_B1_c_219_n 0.0402549f $X=-0.19 $Y=-0.245 $X2=1.205 $Y2=0.74
cc_19 VNB N_B1_c_220_n 0.00873306f $X=-0.19 $Y=-0.245 $X2=2.28 $Y2=1.195
cc_20 VNB N_C1_c_262_n 0.00730236f $X=-0.19 $Y=-0.245 $X2=3.235 $Y2=0.68
cc_21 VNB N_C1_M1006_g 0.0109671f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_C1_c_264_n 0.0159635f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.4
cc_23 VNB N_C1_c_265_n 0.0129564f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.4
cc_24 VNB N_C1_c_266_n 0.0649024f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_C1_c_267_n 0.0130621f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.485
cc_26 VNB N_X_c_300_n 0.0728325f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_X_c_301_n 0.0287783f $X=-0.19 $Y=-0.245 $X2=3.29 $Y2=2.105
cc_28 VNB N_VPWR_c_321_n 0.163682f $X=-0.19 $Y=-0.245 $X2=1.33 $Y2=1.525
cc_29 VNB N_VGND_c_396_n 0.0106392f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_397_n 0.03389f $X=-0.19 $Y=-0.245 $X2=1.205 $Y2=1.32
cc_31 VNB N_VGND_c_398_n 0.00716336f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_399_n 0.0350575f $X=-0.19 $Y=-0.245 $X2=2.28 $Y2=1.195
cc_33 VNB N_VGND_c_400_n 0.018627f $X=-0.19 $Y=-0.245 $X2=1.33 $Y2=1.195
cc_34 VNB N_VGND_c_401_n 0.236325f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_402_n 0.00846609f $X=-0.19 $Y=-0.245 $X2=2.445 $Y2=1.02
cc_36 VNB N_VGND_c_403_n 0.00311272f $X=-0.19 $Y=-0.245 $X2=2.445 $Y2=1.18
cc_37 VPB N_A_81_264#_c_71_n 0.0227063f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.765
cc_38 VPB N_A_81_264#_c_65_n 0.0105479f $X=-0.19 $Y=1.66 $X2=0.585 $Y2=1.485
cc_39 VPB N_A_81_264#_c_69_n 0.0608363f $X=-0.19 $Y=1.66 $X2=3.29 $Y2=2.105
cc_40 VPB N_A2_c_144_n 0.0475003f $X=-0.19 $Y=1.66 $X2=2.305 $Y2=0.68
cc_41 VPB A2 6.38721e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_42 VPB N_A1_c_176_n 0.0333648f $X=-0.19 $Y=1.66 $X2=2.305 $Y2=0.68
cc_43 VPB A1 0.00274431f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_44 VPB N_B1_c_217_n 0.00623388f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_45 VPB N_B1_c_222_n 0.0218019f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_46 VPB N_C1_c_262_n 0.0085689f $X=-0.19 $Y=1.66 $X2=3.235 $Y2=0.68
cc_47 VPB N_C1_c_269_n 0.0266571f $X=-0.19 $Y=1.66 $X2=3.14 $Y2=1.96
cc_48 VPB X 0.0132919f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=2.4
cc_49 VPB X 0.0420202f $X=-0.19 $Y=1.66 $X2=1.115 $Y2=1.485
cc_50 VPB N_X_c_301_n 0.00772285f $X=-0.19 $Y=1.66 $X2=3.29 $Y2=2.105
cc_51 VPB N_VPWR_c_322_n 0.034239f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_52 VPB N_VPWR_c_323_n 0.00835244f $X=-0.19 $Y=1.66 $X2=1.205 $Y2=0.74
cc_53 VPB N_VPWR_c_324_n 0.0291961f $X=-0.19 $Y=1.66 $X2=1.13 $Y2=1.485
cc_54 VPB N_VPWR_c_325_n 0.00382106f $X=-0.19 $Y=1.66 $X2=1.245 $Y2=1.525
cc_55 VPB N_VPWR_c_326_n 0.0196317f $X=-0.19 $Y=1.66 $X2=1.115 $Y2=1.485
cc_56 VPB N_VPWR_c_327_n 0.0522023f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_57 VPB N_VPWR_c_321_n 0.0996142f $X=-0.19 $Y=1.66 $X2=1.33 $Y2=1.525
cc_58 VPB N_VPWR_c_329_n 0.0047828f $X=-0.19 $Y=1.66 $X2=2.445 $Y2=1.02
cc_59 VPB N_A_279_392#_c_360_n 0.0063052f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_60 VPB N_A_279_392#_c_361_n 0.0162509f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_61 VPB N_A_279_392#_c_362_n 0.0042359f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=2.4
cc_62 VPB N_A_279_392#_c_363_n 0.00251823f $X=-0.19 $Y=1.66 $X2=1.205 $Y2=1.32
cc_63 VPB N_A_279_392#_c_364_n 0.00257348f $X=-0.19 $Y=1.66 $X2=1.205 $Y2=0.74
cc_64 N_A_81_264#_c_66_n N_A2_c_144_n 0.011377f $X=1.13 $Y=1.485 $X2=-0.19
+ $Y2=-0.245
cc_65 N_A_81_264#_c_67_n N_A2_c_144_n 0.00275112f $X=2.28 $Y=1.195 $X2=-0.19
+ $Y2=-0.245
cc_66 N_A_81_264#_c_70_n N_A2_c_144_n 0.00128716f $X=1.33 $Y=1.195 $X2=-0.19
+ $Y2=-0.245
cc_67 N_A_81_264#_M1004_g N_A2_M1008_g 0.0184608f $X=1.205 $Y=0.74 $X2=0 $Y2=0
cc_68 N_A_81_264#_c_67_n N_A2_M1008_g 0.0143446f $X=2.28 $Y=1.195 $X2=0 $Y2=0
cc_69 N_A_81_264#_c_70_n N_A2_M1008_g 0.00348718f $X=1.33 $Y=1.195 $X2=0 $Y2=0
cc_70 N_A_81_264#_c_80_p N_A2_M1008_g 0.00119896f $X=2.445 $Y=1.02 $X2=0 $Y2=0
cc_71 N_A_81_264#_c_67_n A2 0.0158156f $X=2.28 $Y=1.195 $X2=0 $Y2=0
cc_72 N_A_81_264#_c_70_n A2 0.0147172f $X=1.33 $Y=1.195 $X2=0 $Y2=0
cc_73 N_A_81_264#_c_67_n N_A1_c_176_n 0.00238064f $X=2.28 $Y=1.195 $X2=-0.19
+ $Y2=-0.245
cc_74 N_A_81_264#_c_80_p N_A1_c_176_n 0.00146597f $X=2.445 $Y=1.02 $X2=-0.19
+ $Y2=-0.245
cc_75 N_A_81_264#_c_67_n N_A1_M1009_g 0.00929703f $X=2.28 $Y=1.195 $X2=0 $Y2=0
cc_76 N_A_81_264#_c_80_p N_A1_M1009_g 0.00740969f $X=2.445 $Y=1.02 $X2=0 $Y2=0
cc_77 N_A_81_264#_c_67_n A1 0.0149787f $X=2.28 $Y=1.195 $X2=0 $Y2=0
cc_78 N_A_81_264#_c_88_p A1 0.00978427f $X=3.125 $Y=1.18 $X2=0 $Y2=0
cc_79 N_A_81_264#_c_69_n A1 0.0142203f $X=3.29 $Y=2.105 $X2=0 $Y2=0
cc_80 N_A_81_264#_c_80_p A1 0.0221054f $X=2.445 $Y=1.02 $X2=0 $Y2=0
cc_81 N_A_81_264#_c_88_p N_B1_M1005_g 0.0105499f $X=3.125 $Y=1.18 $X2=0 $Y2=0
cc_82 N_A_81_264#_c_69_n N_B1_M1005_g 6.23577e-19 $X=3.29 $Y=2.105 $X2=0 $Y2=0
cc_83 N_A_81_264#_c_80_p N_B1_M1005_g 0.00657043f $X=2.445 $Y=1.02 $X2=0 $Y2=0
cc_84 N_A_81_264#_c_69_n N_B1_c_216_n 0.00160032f $X=3.29 $Y=2.105 $X2=0 $Y2=0
cc_85 N_A_81_264#_c_69_n N_B1_c_222_n 0.00318869f $X=3.29 $Y=2.105 $X2=0 $Y2=0
cc_86 N_A_81_264#_c_88_p N_B1_c_218_n 0.00435412f $X=3.125 $Y=1.18 $X2=0 $Y2=0
cc_87 N_A_81_264#_c_80_p N_B1_c_218_n 0.0147688f $X=2.445 $Y=1.02 $X2=0 $Y2=0
cc_88 N_A_81_264#_c_88_p N_B1_c_219_n 7.3851e-19 $X=3.125 $Y=1.18 $X2=0 $Y2=0
cc_89 N_A_81_264#_c_67_n N_B1_c_220_n 0.0074564f $X=2.28 $Y=1.195 $X2=0 $Y2=0
cc_90 N_A_81_264#_c_69_n N_C1_c_262_n 0.00916022f $X=3.29 $Y=2.105 $X2=0 $Y2=0
cc_91 N_A_81_264#_c_69_n N_C1_c_269_n 0.0239338f $X=3.29 $Y=2.105 $X2=0 $Y2=0
cc_92 N_A_81_264#_c_88_p N_C1_M1006_g 0.00577939f $X=3.125 $Y=1.18 $X2=0 $Y2=0
cc_93 N_A_81_264#_c_68_n N_C1_M1006_g 0.00432932f $X=3.332 $Y=1.28 $X2=0 $Y2=0
cc_94 N_A_81_264#_c_69_n N_C1_M1006_g 0.00442215f $X=3.29 $Y=2.105 $X2=0 $Y2=0
cc_95 N_A_81_264#_c_80_p N_C1_M1006_g 6.44932e-19 $X=2.445 $Y=1.02 $X2=0 $Y2=0
cc_96 N_A_81_264#_c_88_p N_C1_c_264_n 0.00380231f $X=3.125 $Y=1.18 $X2=0 $Y2=0
cc_97 N_A_81_264#_c_69_n N_C1_c_264_n 0.00866992f $X=3.29 $Y=2.105 $X2=0 $Y2=0
cc_98 N_A_81_264#_c_68_n N_C1_c_266_n 0.00462642f $X=3.332 $Y=1.28 $X2=0 $Y2=0
cc_99 N_A_81_264#_c_68_n N_C1_c_267_n 0.00731659f $X=3.332 $Y=1.28 $X2=0 $Y2=0
cc_100 N_A_81_264#_M1004_g N_X_c_300_n 0.00216353f $X=1.205 $Y=0.74 $X2=0 $Y2=0
cc_101 N_A_81_264#_c_65_n N_X_c_300_n 0.0172391f $X=0.585 $Y=1.485 $X2=0 $Y2=0
cc_102 N_A_81_264#_c_112_p N_X_c_300_n 0.0381409f $X=1.245 $Y=1.525 $X2=0 $Y2=0
cc_103 N_A_81_264#_c_70_n N_X_c_300_n 0.00156681f $X=1.33 $Y=1.195 $X2=0 $Y2=0
cc_104 N_A_81_264#_c_71_n X 0.00264835f $X=0.495 $Y=1.765 $X2=0 $Y2=0
cc_105 N_A_81_264#_c_65_n X 7.80018e-19 $X=0.585 $Y=1.485 $X2=0 $Y2=0
cc_106 N_A_81_264#_c_112_p X 7.04289e-19 $X=1.245 $Y=1.525 $X2=0 $Y2=0
cc_107 N_A_81_264#_c_71_n X 0.0121388f $X=0.495 $Y=1.765 $X2=0 $Y2=0
cc_108 N_A_81_264#_c_65_n N_X_c_301_n 0.0142734f $X=0.585 $Y=1.485 $X2=0 $Y2=0
cc_109 N_A_81_264#_c_112_p N_X_c_301_n 0.0198186f $X=1.245 $Y=1.525 $X2=0 $Y2=0
cc_110 N_A_81_264#_c_71_n N_VPWR_c_322_n 0.0100916f $X=0.495 $Y=1.765 $X2=0
+ $Y2=0
cc_111 N_A_81_264#_c_66_n N_VPWR_c_322_n 0.00577732f $X=1.13 $Y=1.485 $X2=0
+ $Y2=0
cc_112 N_A_81_264#_c_112_p N_VPWR_c_322_n 0.0205252f $X=1.245 $Y=1.525 $X2=0
+ $Y2=0
cc_113 N_A_81_264#_c_71_n N_VPWR_c_326_n 0.00445602f $X=0.495 $Y=1.765 $X2=0
+ $Y2=0
cc_114 N_A_81_264#_c_69_n N_VPWR_c_327_n 0.0183866f $X=3.29 $Y=2.105 $X2=0 $Y2=0
cc_115 N_A_81_264#_c_71_n N_VPWR_c_321_n 0.00865852f $X=0.495 $Y=1.765 $X2=0
+ $Y2=0
cc_116 N_A_81_264#_c_69_n N_VPWR_c_321_n 0.0151859f $X=3.29 $Y=2.105 $X2=0 $Y2=0
cc_117 N_A_81_264#_c_67_n N_A_279_392#_c_360_n 0.00525329f $X=2.28 $Y=1.195
+ $X2=0 $Y2=0
cc_118 N_A_81_264#_c_70_n N_A_279_392#_c_360_n 0.00365135f $X=1.33 $Y=1.195
+ $X2=0 $Y2=0
cc_119 N_A_81_264#_c_67_n N_A_279_392#_c_362_n 0.0050898f $X=2.28 $Y=1.195 $X2=0
+ $Y2=0
cc_120 N_A_81_264#_c_69_n N_A_279_392#_c_363_n 0.00560794f $X=3.29 $Y=2.105
+ $X2=0 $Y2=0
cc_121 N_A_81_264#_c_69_n N_A_279_392#_c_364_n 0.0267619f $X=3.29 $Y=2.105 $X2=0
+ $Y2=0
cc_122 N_A_81_264#_c_67_n N_VGND_M1004_d 0.00549f $X=2.28 $Y=1.195 $X2=-0.19
+ $Y2=-0.245
cc_123 N_A_81_264#_c_70_n N_VGND_M1004_d 0.00147249f $X=1.33 $Y=1.195 $X2=-0.19
+ $Y2=-0.245
cc_124 N_A_81_264#_c_88_p N_VGND_M1005_d 0.0101595f $X=3.125 $Y=1.18 $X2=0 $Y2=0
cc_125 N_A_81_264#_M1004_g N_VGND_c_396_n 0.0185781f $X=1.205 $Y=0.74 $X2=0
+ $Y2=0
cc_126 N_A_81_264#_c_67_n N_VGND_c_396_n 0.0187286f $X=2.28 $Y=1.195 $X2=0 $Y2=0
cc_127 N_A_81_264#_c_70_n N_VGND_c_396_n 0.0113056f $X=1.33 $Y=1.195 $X2=0 $Y2=0
cc_128 N_A_81_264#_c_80_p N_VGND_c_396_n 0.00281502f $X=2.445 $Y=1.02 $X2=0
+ $Y2=0
cc_129 N_A_81_264#_c_88_p N_VGND_c_411_n 0.0200298f $X=3.125 $Y=1.18 $X2=0 $Y2=0
cc_130 N_A_81_264#_c_68_n N_VGND_c_411_n 0.00682172f $X=3.332 $Y=1.28 $X2=0
+ $Y2=0
cc_131 N_A_81_264#_M1004_g N_VGND_c_399_n 0.00383152f $X=1.205 $Y=0.74 $X2=0
+ $Y2=0
cc_132 N_A_81_264#_M1004_g N_VGND_c_401_n 0.00762539f $X=1.205 $Y=0.74 $X2=0
+ $Y2=0
cc_133 N_A_81_264#_c_67_n A_366_136# 0.0107009f $X=2.28 $Y=1.195 $X2=-0.19
+ $Y2=-0.245
cc_134 N_A2_c_144_n N_A1_c_176_n 0.0432681f $X=1.745 $Y=1.885 $X2=-0.19
+ $Y2=-0.245
cc_135 A2 N_A1_c_176_n 4.15752e-19 $X=1.595 $Y=1.58 $X2=-0.19 $Y2=-0.245
cc_136 N_A2_M1008_g N_A1_M1009_g 0.0345428f $X=1.755 $Y=1 $X2=0 $Y2=0
cc_137 N_A2_c_144_n A1 0.0011401f $X=1.745 $Y=1.885 $X2=0 $Y2=0
cc_138 A2 A1 0.0217322f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_139 N_A2_M1008_g N_B1_c_220_n 9.20121e-19 $X=1.755 $Y=1 $X2=0 $Y2=0
cc_140 N_A2_c_144_n N_VPWR_c_323_n 0.00507786f $X=1.745 $Y=1.885 $X2=0 $Y2=0
cc_141 N_A2_c_144_n N_VPWR_c_324_n 0.00445602f $X=1.745 $Y=1.885 $X2=0 $Y2=0
cc_142 N_A2_c_144_n N_VPWR_c_321_n 0.00862738f $X=1.745 $Y=1.885 $X2=0 $Y2=0
cc_143 N_A2_c_144_n N_A_279_392#_c_360_n 0.00403451f $X=1.745 $Y=1.885 $X2=0
+ $Y2=0
cc_144 A2 N_A_279_392#_c_360_n 0.00832201f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_145 N_A2_c_144_n N_A_279_392#_c_361_n 0.0106338f $X=1.745 $Y=1.885 $X2=0
+ $Y2=0
cc_146 N_A2_c_144_n N_A_279_392#_c_362_n 0.0125514f $X=1.745 $Y=1.885 $X2=0
+ $Y2=0
cc_147 A2 N_A_279_392#_c_362_n 0.0107144f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_148 N_A2_c_144_n N_A_279_392#_c_364_n 6.36743e-19 $X=1.745 $Y=1.885 $X2=0
+ $Y2=0
cc_149 N_A2_M1008_g N_VGND_c_396_n 0.00973412f $X=1.755 $Y=1 $X2=0 $Y2=0
cc_150 N_A2_M1008_g N_VGND_c_397_n 0.00322089f $X=1.755 $Y=1 $X2=0 $Y2=0
cc_151 N_A2_M1008_g N_VGND_c_401_n 0.00381775f $X=1.755 $Y=1 $X2=0 $Y2=0
cc_152 N_A1_M1009_g N_B1_M1005_g 0.0234991f $X=2.23 $Y=1 $X2=0 $Y2=0
cc_153 N_A1_c_176_n N_B1_c_216_n 0.0213265f $X=2.225 $Y=1.885 $X2=0 $Y2=0
cc_154 A1 N_B1_c_216_n 0.00337715f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_155 N_A1_c_176_n N_B1_c_217_n 0.00563966f $X=2.225 $Y=1.885 $X2=0 $Y2=0
cc_156 A1 N_B1_c_217_n 0.0168748f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_157 N_A1_c_176_n N_B1_c_222_n 0.00907122f $X=2.225 $Y=1.885 $X2=0 $Y2=0
cc_158 N_A1_M1009_g N_B1_c_218_n 0.00125823f $X=2.23 $Y=1 $X2=0 $Y2=0
cc_159 N_A1_M1009_g N_B1_c_219_n 0.00110296f $X=2.23 $Y=1 $X2=0 $Y2=0
cc_160 N_A1_M1009_g N_B1_c_220_n 0.00886977f $X=2.23 $Y=1 $X2=0 $Y2=0
cc_161 A1 N_C1_c_264_n 0.0011425f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_162 N_A1_c_176_n N_VPWR_c_323_n 0.00507786f $X=2.225 $Y=1.885 $X2=0 $Y2=0
cc_163 N_A1_c_176_n N_VPWR_c_327_n 0.00445602f $X=2.225 $Y=1.885 $X2=0 $Y2=0
cc_164 N_A1_c_176_n N_VPWR_c_321_n 0.0085802f $X=2.225 $Y=1.885 $X2=0 $Y2=0
cc_165 N_A1_c_176_n N_A_279_392#_c_361_n 6.36743e-19 $X=2.225 $Y=1.885 $X2=0
+ $Y2=0
cc_166 N_A1_c_176_n N_A_279_392#_c_362_n 0.0144848f $X=2.225 $Y=1.885 $X2=0
+ $Y2=0
cc_167 A1 N_A_279_392#_c_362_n 0.0174981f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_168 N_A1_c_176_n N_A_279_392#_c_363_n 0.00238554f $X=2.225 $Y=1.885 $X2=0
+ $Y2=0
cc_169 A1 N_A_279_392#_c_363_n 0.0285613f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_170 N_A1_c_176_n N_A_279_392#_c_364_n 0.0104821f $X=2.225 $Y=1.885 $X2=0
+ $Y2=0
cc_171 N_A1_M1009_g N_VGND_c_396_n 0.00122805f $X=2.23 $Y=1 $X2=0 $Y2=0
cc_172 N_A1_M1009_g N_VGND_c_397_n 4.93445e-19 $X=2.23 $Y=1 $X2=0 $Y2=0
cc_173 N_B1_c_217_n N_C1_c_262_n 0.00972148f $X=2.675 $Y=1.795 $X2=0 $Y2=0
cc_174 N_B1_c_222_n N_C1_c_269_n 0.0696973f $X=2.675 $Y=1.885 $X2=0 $Y2=0
cc_175 N_B1_M1005_g N_C1_M1006_g 0.0216012f $X=2.66 $Y=1 $X2=0 $Y2=0
cc_176 N_B1_c_216_n N_C1_c_264_n 0.00972148f $X=2.675 $Y=1.485 $X2=0 $Y2=0
cc_177 N_B1_c_218_n N_C1_c_265_n 3.55191e-19 $X=2.71 $Y=0.405 $X2=0 $Y2=0
cc_178 N_B1_c_219_n N_C1_c_265_n 0.0214776f $X=2.71 $Y=0.405 $X2=0 $Y2=0
cc_179 N_B1_c_222_n N_VPWR_c_327_n 0.00445602f $X=2.675 $Y=1.885 $X2=0 $Y2=0
cc_180 N_B1_c_222_n N_VPWR_c_321_n 0.00857948f $X=2.675 $Y=1.885 $X2=0 $Y2=0
cc_181 N_B1_c_222_n N_A_279_392#_c_363_n 0.00354727f $X=2.675 $Y=1.885 $X2=0
+ $Y2=0
cc_182 N_B1_c_222_n N_A_279_392#_c_364_n 0.0143199f $X=2.675 $Y=1.885 $X2=0
+ $Y2=0
cc_183 N_B1_c_220_n N_VGND_c_396_n 0.0221185f $X=2.275 $Y=0.462 $X2=0 $Y2=0
cc_184 N_B1_c_219_n N_VGND_c_397_n 0.00584621f $X=2.71 $Y=0.405 $X2=0 $Y2=0
cc_185 N_B1_c_220_n N_VGND_c_397_n 0.055077f $X=2.275 $Y=0.462 $X2=0 $Y2=0
cc_186 N_B1_M1005_g N_VGND_c_398_n 0.00215652f $X=2.66 $Y=1 $X2=0 $Y2=0
cc_187 N_B1_c_218_n N_VGND_c_398_n 0.0250136f $X=2.71 $Y=0.405 $X2=0 $Y2=0
cc_188 N_B1_c_219_n N_VGND_c_398_n 0.00121901f $X=2.71 $Y=0.405 $X2=0 $Y2=0
cc_189 N_B1_c_218_n N_VGND_c_411_n 0.00633625f $X=2.71 $Y=0.405 $X2=0 $Y2=0
cc_190 N_B1_c_219_n N_VGND_c_411_n 0.00210363f $X=2.71 $Y=0.405 $X2=0 $Y2=0
cc_191 N_B1_c_219_n N_VGND_c_401_n 0.00754635f $X=2.71 $Y=0.405 $X2=0 $Y2=0
cc_192 N_B1_c_220_n N_VGND_c_401_n 0.0301837f $X=2.275 $Y=0.462 $X2=0 $Y2=0
cc_193 N_C1_c_269_n N_VPWR_c_327_n 0.00445602f $X=3.065 $Y=1.885 $X2=0 $Y2=0
cc_194 N_C1_c_269_n N_VPWR_c_321_n 0.00861971f $X=3.065 $Y=1.885 $X2=0 $Y2=0
cc_195 N_C1_c_269_n N_A_279_392#_c_363_n 4.73984e-19 $X=3.065 $Y=1.885 $X2=0
+ $Y2=0
cc_196 N_C1_c_269_n N_A_279_392#_c_364_n 0.00240695f $X=3.065 $Y=1.885 $X2=0
+ $Y2=0
cc_197 N_C1_M1006_g N_VGND_c_398_n 0.00617796f $X=3.16 $Y=1 $X2=0 $Y2=0
cc_198 N_C1_c_265_n N_VGND_c_398_n 0.0123056f $X=3.235 $Y=0.405 $X2=0 $Y2=0
cc_199 N_C1_c_267_n N_VGND_c_398_n 0.0300116f $X=3.55 $Y=0.405 $X2=0 $Y2=0
cc_200 N_C1_M1006_g N_VGND_c_411_n 0.0110866f $X=3.16 $Y=1 $X2=0 $Y2=0
cc_201 N_C1_c_265_n N_VGND_c_400_n 0.0106085f $X=3.235 $Y=0.405 $X2=0 $Y2=0
cc_202 N_C1_c_267_n N_VGND_c_400_n 0.0215843f $X=3.55 $Y=0.405 $X2=0 $Y2=0
cc_203 N_C1_c_265_n N_VGND_c_401_n 0.00124593f $X=3.235 $Y=0.405 $X2=0 $Y2=0
cc_204 N_C1_c_266_n N_VGND_c_401_n 0.0154555f $X=3.55 $Y=0.405 $X2=0 $Y2=0
cc_205 N_C1_c_267_n N_VGND_c_401_n 0.0110944f $X=3.55 $Y=0.405 $X2=0 $Y2=0
cc_206 X N_VPWR_c_322_n 0.0781509f $X=0.155 $Y=1.95 $X2=0 $Y2=0
cc_207 X N_VPWR_c_326_n 0.0154862f $X=0.24 $Y=2.035 $X2=0 $Y2=0
cc_208 X N_VPWR_c_321_n 0.0127853f $X=0.24 $Y=2.035 $X2=0 $Y2=0
cc_209 N_X_c_300_n N_VGND_c_396_n 0.0233861f $X=0.17 $Y=0.737 $X2=0 $Y2=0
cc_210 N_X_c_300_n N_VGND_c_399_n 0.0359798f $X=0.17 $Y=0.737 $X2=0 $Y2=0
cc_211 N_X_c_300_n N_VGND_c_401_n 0.0351661f $X=0.17 $Y=0.737 $X2=0 $Y2=0
cc_212 N_VPWR_c_322_n N_A_279_392#_c_360_n 0.00728152f $X=0.72 $Y=1.985 $X2=0
+ $Y2=0
cc_213 N_VPWR_c_322_n N_A_279_392#_c_361_n 0.0347066f $X=0.72 $Y=1.985 $X2=0
+ $Y2=0
cc_214 N_VPWR_c_323_n N_A_279_392#_c_361_n 0.0455206f $X=1.985 $Y=2.455 $X2=0
+ $Y2=0
cc_215 N_VPWR_c_324_n N_A_279_392#_c_361_n 0.0145938f $X=1.885 $Y=3.33 $X2=0
+ $Y2=0
cc_216 N_VPWR_c_321_n N_A_279_392#_c_361_n 0.0120466f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_217 N_VPWR_M1002_d N_A_279_392#_c_362_n 0.00279158f $X=1.82 $Y=1.96 $X2=0
+ $Y2=0
cc_218 N_VPWR_c_323_n N_A_279_392#_c_362_n 0.016109f $X=1.985 $Y=2.455 $X2=0
+ $Y2=0
cc_219 N_VPWR_c_323_n N_A_279_392#_c_364_n 0.0455206f $X=1.985 $Y=2.455 $X2=0
+ $Y2=0
cc_220 N_VPWR_c_327_n N_A_279_392#_c_364_n 0.014552f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_221 N_VPWR_c_321_n N_A_279_392#_c_364_n 0.0119791f $X=3.6 $Y=3.33 $X2=0 $Y2=0
