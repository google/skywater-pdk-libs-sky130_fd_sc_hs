* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hs__einvp_2 A TE VGND VNB VPB VPWR Z
M1000 VGND TE a_263_323# VNB nlowvt w=420000u l=150000u
+  ad=3.332e+11p pd=3.48e+06u as=1.197e+11p ps=1.41e+06u
M1001 a_36_74# A Z VNB nlowvt w=740000u l=150000u
+  ad=6.29e+11p pd=6.14e+06u as=2.072e+11p ps=2.04e+06u
M1002 VGND TE a_36_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1003 a_27_368# A Z VPB pshort w=1.12e+06u l=150000u
+  ad=9.912e+11p pd=8.49e+06u as=3.36e+11p ps=2.84e+06u
M1004 VPWR TE a_263_323# VPB pshort w=640000u l=150000u
+  ad=5.248e+11p pd=4.71e+06u as=1.856e+11p ps=1.86e+06u
M1005 Z A a_27_368# VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VPWR a_263_323# a_27_368# VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_27_368# a_263_323# VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_36_74# TE VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 Z A a_36_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
