* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hs__mux2_1 A0 A1 S VGND VNB VPB VPWR X
X0 a_27_112# S VPWR VPB sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X1 a_304_74# A1 a_524_368# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=150000u
X2 a_443_74# a_27_112# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X3 a_226_74# A1 a_304_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X4 VPWR S a_223_368# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=150000u
X5 VGND S a_226_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X6 a_524_368# a_27_112# VPWR VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=150000u
X7 a_27_112# S VGND VNB sky130_fd_pr__nfet_01v8_lvt w=550000u l=150000u
X8 VGND a_304_74# X VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X9 a_223_368# A0 a_304_74# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=150000u
X10 a_304_74# A0 a_443_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X11 VPWR a_304_74# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
.ends
