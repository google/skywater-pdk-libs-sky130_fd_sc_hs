* NGSPICE file created from sky130_fd_sc_hs__dfxbp_2.ext - technology: sky130A

.subckt sky130_fd_sc_hs__dfxbp_2 CLK D VGND VNB VPB VPWR Q Q_N
M1000 a_1000_424# a_27_74# a_753_284# VPB pshort w=840000u l=150000u
+  ad=4.851e+11p pd=3.46e+06u as=2.52e+11p ps=2.28e+06u
M1001 Q a_1290_102# VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=3.36e+11p pd=2.84e+06u as=2.84038e+12p ps=2.25e+07u
M1002 a_1248_128# a_27_74# a_1000_424# VNB nlowvt w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=3.9205e+11p ps=3.36e+06u
M1003 Q a_1290_102# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.072e+11p pd=2.04e+06u as=2.11565e+12p ps=1.739e+07u
M1004 VGND a_753_284# a_717_102# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1005 VPWR a_753_284# a_702_445# VPB pshort w=420000u l=150000u
+  ad=0p pd=0u as=1.134e+11p ps=1.38e+06u
M1006 Q_N a_1835_368# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.072e+11p pd=2.04e+06u as=0p ps=0u
M1007 a_753_284# a_558_445# VGND VNB nlowvt w=550000u l=150000u
+  ad=3.87e+11p pd=2.98e+06u as=0p ps=0u
M1008 VGND a_1835_368# Q_N VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VPWR a_1290_102# Q VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VGND a_1290_102# a_1248_128# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_206_368# a_27_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=3.252e+11p pd=2.59e+06u as=0p ps=0u
M1012 a_1000_424# a_206_368# a_753_284# VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VGND a_1290_102# Q VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_717_102# a_206_368# a_558_445# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.66075e+11p ps=1.73e+06u
M1015 a_1290_102# a_1000_424# VPWR VPB pshort w=840000u l=150000u
+  ad=2.52e+11p pd=2.28e+06u as=0p ps=0u
M1016 a_206_368# a_27_74# VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=3.304e+11p pd=2.83e+06u as=0p ps=0u
M1017 VPWR CLK a_27_74# VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=3.304e+11p ps=2.83e+06u
M1018 Q_N a_1835_368# VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=3.36e+11p pd=2.84e+06u as=0p ps=0u
M1019 VPWR a_1290_102# a_1835_368# VPB pshort w=1e+06u l=150000u
+  ad=0p pd=0u as=2.95e+11p ps=2.59e+06u
M1020 VPWR a_1000_424# a_1290_102# VPB pshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 VGND a_1000_424# a_1290_102# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1022 a_451_503# D VPWR VPB pshort w=420000u l=150000u
+  ad=2.1245e+11p pd=2.19e+06u as=0p ps=0u
M1023 VPWR a_1835_368# Q_N VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 a_451_503# D VGND VNB nlowvt w=420000u l=150000u
+  ad=1.176e+11p pd=1.4e+06u as=0p ps=0u
M1025 VGND CLK a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1026 a_558_445# a_27_74# a_451_503# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 VGND a_1290_102# a_1835_368# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=1.824e+11p ps=1.85e+06u
M1028 a_558_445# a_206_368# a_451_503# VPB pshort w=420000u l=150000u
+  ad=2.394e+11p pd=1.98e+06u as=0p ps=0u
M1029 a_702_445# a_27_74# a_558_445# VPB pshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1030 a_1208_479# a_206_368# a_1000_424# VPB pshort w=420000u l=150000u
+  ad=1.785e+11p pd=1.69e+06u as=0p ps=0u
M1031 a_753_284# a_558_445# VPWR VPB pshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1032 VPWR a_1290_102# a_1208_479# VPB pshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

