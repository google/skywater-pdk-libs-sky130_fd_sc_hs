* File: sky130_fd_sc_hs__o221ai_1.pex.spice
* Created: Tue Sep  1 20:15:45 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HS__O221AI_1%C1 3 5 7 8 12 13
c27 5 0 9.64256e-20 $X=0.635 $Y=1.765
r28 13 14 20.8272 $w=3.24e-07 $l=1.4e-07 $layer=POLY_cond $X=0.495 $Y=1.532
+ $X2=0.635 $Y2=1.532
r29 11 13 33.4722 $w=3.24e-07 $l=2.25e-07 $layer=POLY_cond $X=0.27 $Y=1.532
+ $X2=0.495 $Y2=1.532
r30 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.27
+ $Y=1.465 $X2=0.27 $Y2=1.465
r31 8 12 6.9845 $w=3.28e-07 $l=2e-07 $layer=LI1_cond $X=0.27 $Y=1.665 $X2=0.27
+ $Y2=1.465
r32 5 14 20.7868 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=0.635 $Y=1.765
+ $X2=0.635 $Y2=1.532
r33 5 7 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.635 $Y=1.765
+ $X2=0.635 $Y2=2.4
r34 1 13 20.7868 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=0.495 $Y=1.3
+ $X2=0.495 $Y2=1.532
r35 1 3 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=0.495 $Y=1.3 $X2=0.495
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HS__O221AI_1%B1 3 5 8 10 13 14
c34 14 0 9.64256e-20 $X=1.47 $Y=1.515
c35 3 0 5.62133e-20 $X=1.545 $Y=1.765
r36 13 14 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.47
+ $Y=1.515 $X2=1.47 $Y2=1.515
r37 10 14 2.67779 $w=6.68e-07 $l=1.5e-07 $layer=LI1_cond $X=1.3 $Y=1.665 $X2=1.3
+ $Y2=1.515
r38 6 13 37.0704 $w=1.5e-07 $l=2.11941e-07 $layer=POLY_cond $X=1.555 $Y=1.35
+ $X2=1.545 $Y2=1.557
r39 6 8 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.555 $Y=1.35
+ $X2=1.555 $Y2=0.74
r40 3 13 37.0704 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=1.545 $Y=1.765
+ $X2=1.545 $Y2=1.557
r41 3 5 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.545 $Y=1.765
+ $X2=1.545 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_HS__O221AI_1%B2 1 3 6 8 12
c36 12 0 5.62133e-20 $X=2.04 $Y=1.515
c37 6 0 6.24822e-20 $X=2.055 $Y=0.74
r38 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.04
+ $Y=1.515 $X2=2.04 $Y2=1.515
r39 8 12 4.32166 $w=3.98e-07 $l=1.5e-07 $layer=LI1_cond $X=2.075 $Y=1.665
+ $X2=2.075 $Y2=1.515
r40 4 11 38.5562 $w=2.99e-07 $l=1.72337e-07 $layer=POLY_cond $X=2.055 $Y=1.35
+ $X2=2.04 $Y2=1.515
r41 4 6 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.055 $Y=1.35
+ $X2=2.055 $Y2=0.74
r42 1 11 52.2586 $w=2.99e-07 $l=2.85044e-07 $layer=POLY_cond $X=1.965 $Y=1.765
+ $X2=2.04 $Y2=1.515
r43 1 3 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.965 $Y=1.765
+ $X2=1.965 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_HS__O221AI_1%A2 1 3 6 8 9 10 11 19 33
c43 6 0 1.42066e-19 $X=2.555 $Y=0.74
r44 33 34 1.2285 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=2.61 $Y=1.665
+ $X2=2.61 $Y2=1.68
r45 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.61
+ $Y=1.515 $X2=2.61 $Y2=1.515
r46 10 11 17.0562 $w=2.48e-07 $l=3.7e-07 $layer=LI1_cond $X=2.65 $Y=2.405
+ $X2=2.65 $Y2=2.775
r47 9 10 17.0562 $w=2.48e-07 $l=3.7e-07 $layer=LI1_cond $X=2.65 $Y=2.035
+ $X2=2.65 $Y2=2.405
r48 8 33 1.22229 $w=3.28e-07 $l=3.5e-08 $layer=LI1_cond $X=2.61 $Y=1.63 $X2=2.61
+ $Y2=1.665
r49 8 19 4.01609 $w=3.28e-07 $l=1.15e-07 $layer=LI1_cond $X=2.61 $Y=1.63
+ $X2=2.61 $Y2=1.515
r50 8 9 14.7513 $w=2.48e-07 $l=3.2e-07 $layer=LI1_cond $X=2.65 $Y=1.715 $X2=2.65
+ $Y2=2.035
r51 8 34 1.61342 $w=2.48e-07 $l=3.5e-08 $layer=LI1_cond $X=2.65 $Y=1.715
+ $X2=2.65 $Y2=1.68
r52 4 18 38.5562 $w=2.99e-07 $l=1.90526e-07 $layer=POLY_cond $X=2.555 $Y=1.35
+ $X2=2.61 $Y2=1.515
r53 4 6 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.555 $Y=1.35
+ $X2=2.555 $Y2=0.74
r54 1 18 52.2586 $w=2.99e-07 $l=2.85044e-07 $layer=POLY_cond $X=2.535 $Y=1.765
+ $X2=2.61 $Y2=1.515
r55 1 3 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.535 $Y=1.765
+ $X2=2.535 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_HS__O221AI_1%A1 1 3 6 8 9 13
r28 15 16 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.52
+ $Y=1.465 $X2=3.52 $Y2=1.465
r29 13 15 23.0464 $w=3.66e-07 $l=1.75e-07 $layer=POLY_cond $X=3.345 $Y=1.532
+ $X2=3.52 $Y2=1.532
r30 12 13 31.6066 $w=3.66e-07 $l=2.4e-07 $layer=POLY_cond $X=3.105 $Y=1.532
+ $X2=3.345 $Y2=1.532
r31 9 16 1.99346 $w=4.78e-07 $l=8e-08 $layer=LI1_cond $X=3.6 $Y=1.54 $X2=3.52
+ $Y2=1.54
r32 8 16 9.96732 $w=4.78e-07 $l=4e-07 $layer=LI1_cond $X=3.12 $Y=1.54 $X2=3.52
+ $Y2=1.54
r33 4 13 23.7042 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=3.345 $Y=1.3
+ $X2=3.345 $Y2=1.532
r34 4 6 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=3.345 $Y=1.3 $X2=3.345
+ $Y2=0.74
r35 1 12 23.7042 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=3.105 $Y=1.765
+ $X2=3.105 $Y2=1.532
r36 1 3 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.105 $Y=1.765
+ $X2=3.105 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_HS__O221AI_1%Y 1 2 3 12 15 16 17 18 20 28 29 40 44
c51 17 0 9.51097e-20 $X=0.775 $Y=2.035
r52 33 44 26.7487 $w=1.68e-07 $l=4.1e-07 $layer=LI1_cond $X=0.28 $Y=1.045
+ $X2=0.69 $Y2=1.045
r53 33 40 1.22229 $w=3.28e-07 $l=3.5e-08 $layer=LI1_cond $X=0.28 $Y=0.96
+ $X2=0.28 $Y2=0.925
r54 29 33 2.60963 $w=1.68e-07 $l=4e-08 $layer=LI1_cond $X=0.24 $Y=1.045 $X2=0.28
+ $Y2=1.045
r55 29 40 0.873063 $w=3.28e-07 $l=2.5e-08 $layer=LI1_cond $X=0.28 $Y=0.9
+ $X2=0.28 $Y2=0.925
r56 28 29 13.4452 $w=3.28e-07 $l=3.85e-07 $layer=LI1_cond $X=0.28 $Y=0.515
+ $X2=0.28 $Y2=0.9
r57 23 25 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=0.41 $Y=2.035
+ $X2=0.69 $Y2=2.035
r58 18 27 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.19 $Y=2.12 $X2=2.19
+ $Y2=2.035
r59 18 20 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=2.19 $Y=2.12
+ $X2=2.19 $Y2=2.815
r60 17 25 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=0.775 $Y=2.035
+ $X2=0.69 $Y2=2.035
r61 16 27 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.025 $Y=2.035
+ $X2=2.19 $Y2=2.035
r62 16 17 81.5508 $w=1.68e-07 $l=1.25e-06 $layer=LI1_cond $X=2.025 $Y=2.035
+ $X2=0.775 $Y2=2.035
r63 15 25 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.69 $Y=1.95
+ $X2=0.69 $Y2=2.035
r64 14 44 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.69 $Y=1.13
+ $X2=0.69 $Y2=1.045
r65 14 15 53.4973 $w=1.68e-07 $l=8.2e-07 $layer=LI1_cond $X=0.69 $Y=1.13
+ $X2=0.69 $Y2=1.95
r66 12 23 32.0379 $w=2.48e-07 $l=6.95e-07 $layer=LI1_cond $X=0.45 $Y=2.815
+ $X2=0.45 $Y2=2.12
r67 3 27 400 $w=1.7e-07 $l=3.4187e-07 $layer=licon1_PDIFF $count=1 $X=2.04
+ $Y=1.84 $X2=2.19 $Y2=2.115
r68 3 20 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=2.04
+ $Y=1.84 $X2=2.19 $Y2=2.815
r69 2 23 400 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_PDIFF $count=1 $X=0.265
+ $Y=1.84 $X2=0.41 $Y2=2.115
r70 2 12 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=0.265
+ $Y=1.84 $X2=0.41 $Y2=2.815
r71 1 28 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__O221AI_1%VPWR 1 2 9 13 18 19 20 22 35 36 39
c38 1 0 9.51097e-20 $X=0.71 $Y=1.84
r39 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r40 35 36 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r41 33 36 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=3.6 $Y2=3.33
r42 32 33 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r43 30 40 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r44 29 32 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.68 $Y=3.33
+ $X2=3.12 $Y2=3.33
r45 29 30 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r46 27 39 14.7712 $w=1.7e-07 $l=4.08e-07 $layer=LI1_cond $X=1.56 $Y=3.33
+ $X2=1.152 $Y2=3.33
r47 27 29 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=1.56 $Y=3.33
+ $X2=1.68 $Y2=3.33
r48 25 40 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r49 24 25 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r50 22 39 14.7712 $w=1.7e-07 $l=4.07e-07 $layer=LI1_cond $X=0.745 $Y=3.33
+ $X2=1.152 $Y2=3.33
r51 22 24 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=0.745 $Y=3.33
+ $X2=0.72 $Y2=3.33
r52 20 33 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=3.12 $Y2=3.33
r53 20 30 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=1.68 $Y2=3.33
r54 18 32 2.93583 $w=1.68e-07 $l=4.5e-08 $layer=LI1_cond $X=3.165 $Y=3.33
+ $X2=3.12 $Y2=3.33
r55 18 19 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.165 $Y=3.33
+ $X2=3.33 $Y2=3.33
r56 17 35 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=3.495 $Y=3.33
+ $X2=3.6 $Y2=3.33
r57 17 19 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.495 $Y=3.33
+ $X2=3.33 $Y2=3.33
r58 13 16 24.4458 $w=3.28e-07 $l=7e-07 $layer=LI1_cond $X=3.33 $Y=2.115 $X2=3.33
+ $Y2=2.815
r59 11 19 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.33 $Y=3.245
+ $X2=3.33 $Y2=3.33
r60 11 16 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=3.33 $Y=3.245
+ $X2=3.33 $Y2=2.815
r61 7 39 3.16747 $w=8.15e-07 $l=8.5e-08 $layer=LI1_cond $X=1.152 $Y=3.245
+ $X2=1.152 $Y2=3.33
r62 7 9 12.768 $w=8.13e-07 $l=8.7e-07 $layer=LI1_cond $X=1.152 $Y=3.245
+ $X2=1.152 $Y2=2.375
r63 2 16 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=3.18
+ $Y=1.84 $X2=3.33 $Y2=2.815
r64 2 13 400 $w=1.7e-07 $l=3.4187e-07 $layer=licon1_PDIFF $count=1 $X=3.18
+ $Y=1.84 $X2=3.33 $Y2=2.115
r65 1 9 150 $w=1.7e-07 $l=8.35733e-07 $layer=licon1_PDIFF $count=4 $X=0.71
+ $Y=1.84 $X2=1.32 $Y2=2.375
.ends

.subckt PM_SKY130_FD_SC_HS__O221AI_1%A_114_74# 1 2 7 9 14
c23 14 0 1.42066e-19 $X=1.84 $Y=0.435
c24 7 0 6.24822e-20 $X=1.675 $Y=0.435
r25 14 17 6.80989 $w=3.28e-07 $l=1.95e-07 $layer=LI1_cond $X=1.84 $Y=0.435
+ $X2=1.84 $Y2=0.63
r26 9 12 5.93683 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=0.78 $Y=0.435
+ $X2=0.78 $Y2=0.605
r27 8 9 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.945 $Y=0.435
+ $X2=0.78 $Y2=0.435
r28 7 14 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.675 $Y=0.435
+ $X2=1.84 $Y2=0.435
r29 7 8 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=1.675 $Y=0.435
+ $X2=0.945 $Y2=0.435
r30 2 17 182 $w=1.7e-07 $l=3.49571e-07 $layer=licon1_NDIFF $count=1 $X=1.63
+ $Y=0.37 $X2=1.84 $Y2=0.63
r31 1 12 182 $w=1.7e-07 $l=2.96859e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.37 $X2=0.71 $Y2=0.605
.ends

.subckt PM_SKY130_FD_SC_HS__O221AI_1%A_239_74# 1 2 3 10 14 16 20 23 27
r46 23 25 4.53993 $w=3.28e-07 $l=1.3e-07 $layer=LI1_cond $X=1.34 $Y=0.965
+ $X2=1.34 $Y2=1.095
r47 18 20 15.5405 $w=3.28e-07 $l=4.45e-07 $layer=LI1_cond $X=3.56 $Y=0.96
+ $X2=3.56 $Y2=0.515
r48 17 27 8.61065 $w=1.7e-07 $l=1.77059e-07 $layer=LI1_cond $X=2.505 $Y=1.045
+ $X2=2.34 $Y2=1.07
r49 16 18 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.395 $Y=1.045
+ $X2=3.56 $Y2=0.96
r50 16 17 58.0642 $w=1.68e-07 $l=8.9e-07 $layer=LI1_cond $X=3.395 $Y=1.045
+ $X2=2.505 $Y2=1.045
r51 12 27 0.89609 $w=3.3e-07 $l=1.1e-07 $layer=LI1_cond $X=2.34 $Y=0.96 $X2=2.34
+ $Y2=1.07
r52 12 14 15.5405 $w=3.28e-07 $l=4.45e-07 $layer=LI1_cond $X=2.34 $Y=0.96
+ $X2=2.34 $Y2=0.515
r53 11 25 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.505 $Y=1.095
+ $X2=1.34 $Y2=1.095
r54 10 27 8.61065 $w=1.7e-07 $l=1.77059e-07 $layer=LI1_cond $X=2.175 $Y=1.095
+ $X2=2.34 $Y2=1.07
r55 10 11 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.175 $Y=1.095
+ $X2=1.505 $Y2=1.095
r56 3 20 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.42
+ $Y=0.37 $X2=3.56 $Y2=0.515
r57 2 14 91 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=2 $X=2.13
+ $Y=0.37 $X2=2.34 $Y2=0.515
r58 1 23 182 $w=1.7e-07 $l=6.63551e-07 $layer=licon1_NDIFF $count=1 $X=1.195
+ $Y=0.37 $X2=1.34 $Y2=0.965
.ends

.subckt PM_SKY130_FD_SC_HS__O221AI_1%VGND 1 6 8 10 20 21 24
r33 24 25 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r34 21 25 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=3.12
+ $Y2=0
r35 20 21 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r36 18 24 11.9488 $w=1.7e-07 $l=2.75e-07 $layer=LI1_cond $X=3.225 $Y=0 $X2=2.95
+ $Y2=0
r37 18 20 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=3.225 $Y=0 $X2=3.6
+ $Y2=0
r38 17 25 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r39 16 17 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r40 12 16 156.578 $w=1.68e-07 $l=2.4e-06 $layer=LI1_cond $X=0.24 $Y=0 $X2=2.64
+ $Y2=0
r41 12 13 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r42 10 24 11.9488 $w=1.7e-07 $l=2.75e-07 $layer=LI1_cond $X=2.675 $Y=0 $X2=2.95
+ $Y2=0
r43 10 16 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=2.675 $Y=0 $X2=2.64
+ $Y2=0
r44 8 17 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=2.64
+ $Y2=0
r45 8 13 0.468274 $w=4.9e-07 $l=1.68e-06 $layer=MET1_cond $X=1.92 $Y=0 $X2=0.24
+ $Y2=0
r46 4 24 2.31338 $w=5.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.95 $Y=0.085 $X2=2.95
+ $Y2=0
r47 4 6 11.7433 $w=5.48e-07 $l=5.4e-07 $layer=LI1_cond $X=2.95 $Y=0.085 $X2=2.95
+ $Y2=0.625
r48 1 6 91 $w=1.7e-07 $l=6.1441e-07 $layer=licon1_NDIFF $count=2 $X=2.63 $Y=0.37
+ $X2=3.13 $Y2=0.625
.ends

