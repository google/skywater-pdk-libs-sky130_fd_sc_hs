* File: sky130_fd_sc_hs__a211oi_4.pxi.spice
* Created: Thu Aug 27 20:23:54 2020
* 
x_PM_SKY130_FD_SC_HS__A211OI_4%A2 N_A2_c_116_n N_A2_M1002_g N_A2_M1004_g
+ N_A2_c_117_n N_A2_M1006_g N_A2_M1005_g N_A2_c_118_n N_A2_M1023_g N_A2_M1013_g
+ N_A2_c_119_n N_A2_M1026_g N_A2_M1015_g A2 A2 A2 A2 A2 N_A2_c_115_n
+ PM_SKY130_FD_SC_HS__A211OI_4%A2
x_PM_SKY130_FD_SC_HS__A211OI_4%A1 N_A1_M1000_g N_A1_c_196_n N_A1_M1008_g
+ N_A1_M1010_g N_A1_c_197_n N_A1_M1011_g N_A1_M1021_g N_A1_c_198_n N_A1_M1014_g
+ N_A1_M1025_g N_A1_c_199_n N_A1_M1016_g A1 A1 A1 N_A1_c_200_n N_A1_c_195_n
+ PM_SKY130_FD_SC_HS__A211OI_4%A1
x_PM_SKY130_FD_SC_HS__A211OI_4%B1 N_B1_c_269_n N_B1_M1017_g N_B1_c_270_n
+ N_B1_M1022_g N_B1_c_271_n N_B1_M1024_g N_B1_M1001_g N_B1_M1020_g N_B1_c_272_n
+ N_B1_M1027_g B1 B1 B1 B1 N_B1_c_268_n PM_SKY130_FD_SC_HS__A211OI_4%B1
x_PM_SKY130_FD_SC_HS__A211OI_4%C1 N_C1_M1018_g N_C1_c_346_n N_C1_M1003_g
+ N_C1_M1019_g N_C1_c_347_n N_C1_M1007_g N_C1_c_348_n N_C1_M1009_g N_C1_c_349_n
+ N_C1_M1012_g C1 C1 C1 N_C1_c_345_n PM_SKY130_FD_SC_HS__A211OI_4%C1
x_PM_SKY130_FD_SC_HS__A211OI_4%A_77_368# N_A_77_368#_M1002_s N_A_77_368#_M1006_s
+ N_A_77_368#_M1026_s N_A_77_368#_M1011_s N_A_77_368#_M1016_s
+ N_A_77_368#_M1017_d N_A_77_368#_M1024_d N_A_77_368#_c_406_n
+ N_A_77_368#_c_407_n N_A_77_368#_c_418_n N_A_77_368#_c_408_n
+ N_A_77_368#_c_425_n N_A_77_368#_c_409_n N_A_77_368#_c_435_n
+ N_A_77_368#_c_410_n N_A_77_368#_c_441_n N_A_77_368#_c_411_n
+ N_A_77_368#_c_412_n N_A_77_368#_c_452_n N_A_77_368#_c_454_n
+ N_A_77_368#_c_458_n N_A_77_368#_c_461_n N_A_77_368#_c_430_n
+ N_A_77_368#_c_433_n N_A_77_368#_c_446_n N_A_77_368#_c_413_n
+ N_A_77_368#_c_464_n PM_SKY130_FD_SC_HS__A211OI_4%A_77_368#
x_PM_SKY130_FD_SC_HS__A211OI_4%VPWR N_VPWR_M1002_d N_VPWR_M1023_d N_VPWR_M1008_d
+ N_VPWR_M1014_d N_VPWR_c_506_n N_VPWR_c_507_n N_VPWR_c_508_n N_VPWR_c_509_n
+ N_VPWR_c_510_n N_VPWR_c_511_n N_VPWR_c_512_n N_VPWR_c_513_n N_VPWR_c_514_n
+ VPWR N_VPWR_c_515_n N_VPWR_c_516_n N_VPWR_c_505_n N_VPWR_c_518_n
+ N_VPWR_c_519_n PM_SKY130_FD_SC_HS__A211OI_4%VPWR
x_PM_SKY130_FD_SC_HS__A211OI_4%A_901_368# N_A_901_368#_M1017_s
+ N_A_901_368#_M1022_s N_A_901_368#_M1027_s N_A_901_368#_M1007_s
+ N_A_901_368#_M1012_s N_A_901_368#_c_608_n N_A_901_368#_c_609_n
+ N_A_901_368#_c_610_n N_A_901_368#_c_624_n N_A_901_368#_c_611_n
+ N_A_901_368#_c_632_n N_A_901_368#_c_612_n N_A_901_368#_c_637_n
+ N_A_901_368#_c_613_n N_A_901_368#_c_614_n N_A_901_368#_c_615_n
+ N_A_901_368#_c_616_n N_A_901_368#_c_617_n
+ PM_SKY130_FD_SC_HS__A211OI_4%A_901_368#
x_PM_SKY130_FD_SC_HS__A211OI_4%Y N_Y_M1000_s N_Y_M1021_s N_Y_M1001_d N_Y_M1020_d
+ N_Y_M1019_s N_Y_M1003_d N_Y_M1009_d N_Y_c_688_n N_Y_c_689_n N_Y_c_690_n
+ N_Y_c_691_n N_Y_c_692_n N_Y_c_693_n N_Y_c_694_n N_Y_c_695_n N_Y_c_696_n
+ N_Y_c_697_n N_Y_c_730_n Y Y Y Y Y Y Y Y PM_SKY130_FD_SC_HS__A211OI_4%Y
x_PM_SKY130_FD_SC_HS__A211OI_4%A_92_74# N_A_92_74#_M1004_s N_A_92_74#_M1005_s
+ N_A_92_74#_M1015_s N_A_92_74#_M1010_d N_A_92_74#_M1025_d N_A_92_74#_c_765_n
+ N_A_92_74#_c_766_n N_A_92_74#_c_767_n N_A_92_74#_c_768_n N_A_92_74#_c_769_n
+ N_A_92_74#_c_770_n N_A_92_74#_c_771_n N_A_92_74#_c_772_n
+ PM_SKY130_FD_SC_HS__A211OI_4%A_92_74#
x_PM_SKY130_FD_SC_HS__A211OI_4%VGND N_VGND_M1004_d N_VGND_M1013_d N_VGND_M1001_s
+ N_VGND_M1018_d N_VGND_c_816_n N_VGND_c_817_n N_VGND_c_818_n N_VGND_c_819_n
+ N_VGND_c_820_n N_VGND_c_821_n N_VGND_c_822_n N_VGND_c_823_n VGND
+ N_VGND_c_824_n N_VGND_c_825_n N_VGND_c_826_n N_VGND_c_827_n N_VGND_c_828_n
+ N_VGND_c_829_n PM_SKY130_FD_SC_HS__A211OI_4%VGND
cc_1 VNB N_A2_M1004_g 0.0318708f $X=-0.19 $Y=-0.245 $X2=0.8 $Y2=0.74
cc_2 VNB N_A2_M1005_g 0.0224899f $X=-0.19 $Y=-0.245 $X2=1.23 $Y2=0.74
cc_3 VNB N_A2_M1013_g 0.0224899f $X=-0.19 $Y=-0.245 $X2=1.66 $Y2=0.74
cc_4 VNB N_A2_M1015_g 0.0230056f $X=-0.19 $Y=-0.245 $X2=2.09 $Y2=0.74
cc_5 VNB A2 0.0329433f $X=-0.19 $Y=-0.245 $X2=2.075 $Y2=1.58
cc_6 VNB N_A2_c_115_n 0.0727053f $X=-0.19 $Y=-0.245 $X2=2.085 $Y2=1.557
cc_7 VNB N_A1_M1000_g 0.0240886f $X=-0.19 $Y=-0.245 $X2=0.735 $Y2=2.4
cc_8 VNB N_A1_M1010_g 0.0234234f $X=-0.19 $Y=-0.245 $X2=1.185 $Y2=2.4
cc_9 VNB N_A1_M1021_g 0.0234256f $X=-0.19 $Y=-0.245 $X2=1.635 $Y2=2.4
cc_10 VNB N_A1_M1025_g 0.0328863f $X=-0.19 $Y=-0.245 $X2=2.085 $Y2=2.4
cc_11 VNB N_A1_c_195_n 0.0762638f $X=-0.19 $Y=-0.245 $X2=1.66 $Y2=1.557
cc_12 VNB N_B1_M1001_g 0.0289588f $X=-0.19 $Y=-0.245 $X2=1.23 $Y2=0.74
cc_13 VNB N_B1_M1020_g 0.0208323f $X=-0.19 $Y=-0.245 $X2=1.635 $Y2=2.4
cc_14 VNB B1 0.00922652f $X=-0.19 $Y=-0.245 $X2=2.085 $Y2=2.4
cc_15 VNB N_B1_c_268_n 0.124313f $X=-0.19 $Y=-0.245 $X2=0.735 $Y2=1.557
cc_16 VNB N_C1_M1018_g 0.0214f $X=-0.19 $Y=-0.245 $X2=0.735 $Y2=2.4
cc_17 VNB N_C1_M1019_g 0.0270575f $X=-0.19 $Y=-0.245 $X2=1.185 $Y2=2.4
cc_18 VNB C1 0.00375419f $X=-0.19 $Y=-0.245 $X2=2.085 $Y2=2.4
cc_19 VNB N_C1_c_345_n 0.0976733f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_VPWR_c_505_n 0.362705f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.565
cc_21 VNB N_Y_c_688_n 0.00622517f $X=-0.19 $Y=-0.245 $X2=2.085 $Y2=1.765
cc_22 VNB N_Y_c_689_n 0.0721116f $X=-0.19 $Y=-0.245 $X2=2.09 $Y2=0.74
cc_23 VNB N_Y_c_690_n 0.0252102f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_24 VNB N_Y_c_691_n 0.00369528f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=1.58
cc_25 VNB N_Y_c_692_n 0.00178908f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_Y_c_693_n 0.00306324f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_Y_c_694_n 0.109424f $X=-0.19 $Y=-0.245 $X2=0.81 $Y2=1.515
cc_28 VNB N_Y_c_695_n 0.00130318f $X=-0.19 $Y=-0.245 $X2=1.83 $Y2=1.557
cc_29 VNB N_Y_c_696_n 0.00180772f $X=-0.19 $Y=-0.245 $X2=1.83 $Y2=1.515
cc_30 VNB N_Y_c_697_n 0.00354475f $X=-0.19 $Y=-0.245 $X2=1.83 $Y2=1.515
cc_31 VNB N_A_92_74#_c_765_n 0.0270834f $X=-0.19 $Y=-0.245 $X2=1.66 $Y2=1.35
cc_32 VNB N_A_92_74#_c_766_n 0.00307486f $X=-0.19 $Y=-0.245 $X2=1.66 $Y2=0.74
cc_33 VNB N_A_92_74#_c_767_n 0.00963497f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_92_74#_c_768_n 0.00178908f $X=-0.19 $Y=-0.245 $X2=2.085 $Y2=2.4
cc_35 VNB N_A_92_74#_c_769_n 0.00917346f $X=-0.19 $Y=-0.245 $X2=2.09 $Y2=0.74
cc_36 VNB N_A_92_74#_c_770_n 0.0016059f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_92_74#_c_771_n 0.0213494f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_92_74#_c_772_n 0.00127131f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_816_n 0.00323505f $X=-0.19 $Y=-0.245 $X2=1.635 $Y2=1.765
cc_40 VNB N_VGND_c_817_n 0.00323505f $X=-0.19 $Y=-0.245 $X2=1.66 $Y2=0.74
cc_41 VNB N_VGND_c_818_n 0.00323505f $X=-0.19 $Y=-0.245 $X2=2.085 $Y2=2.4
cc_42 VNB N_VGND_c_819_n 0.00323505f $X=-0.19 $Y=-0.245 $X2=2.09 $Y2=0.74
cc_43 VNB N_VGND_c_820_n 0.0270966f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_44 VNB N_VGND_c_821_n 0.00604233f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.58
cc_45 VNB N_VGND_c_822_n 0.0151736f $X=-0.19 $Y=-0.245 $X2=2.075 $Y2=1.58
cc_46 VNB N_VGND_c_823_n 0.00604233f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_VGND_c_824_n 0.10229f $X=-0.19 $Y=-0.245 $X2=1.185 $Y2=1.557
cc_48 VNB N_VGND_c_825_n 0.0151736f $X=-0.19 $Y=-0.245 $X2=2.085 $Y2=1.557
cc_49 VNB N_VGND_c_826_n 0.0437444f $X=-0.19 $Y=-0.245 $X2=0.81 $Y2=1.565
cc_50 VNB N_VGND_c_827_n 0.517711f $X=-0.19 $Y=-0.245 $X2=1.2 $Y2=1.565
cc_51 VNB N_VGND_c_828_n 0.00604233f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_VGND_c_829_n 0.00604233f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VPB N_A2_c_116_n 0.0208611f $X=-0.19 $Y=1.66 $X2=0.735 $Y2=1.765
cc_54 VPB N_A2_c_117_n 0.0155096f $X=-0.19 $Y=1.66 $X2=1.185 $Y2=1.765
cc_55 VPB N_A2_c_118_n 0.015f $X=-0.19 $Y=1.66 $X2=1.635 $Y2=1.765
cc_56 VPB N_A2_c_119_n 0.015303f $X=-0.19 $Y=1.66 $X2=2.085 $Y2=1.765
cc_57 VPB A2 0.028021f $X=-0.19 $Y=1.66 $X2=2.075 $Y2=1.58
cc_58 VPB N_A2_c_115_n 0.047221f $X=-0.19 $Y=1.66 $X2=2.085 $Y2=1.557
cc_59 VPB N_A1_c_196_n 0.0153741f $X=-0.19 $Y=1.66 $X2=0.8 $Y2=0.74
cc_60 VPB N_A1_c_197_n 0.0149968f $X=-0.19 $Y=1.66 $X2=1.23 $Y2=0.74
cc_61 VPB N_A1_c_198_n 0.014996f $X=-0.19 $Y=1.66 $X2=1.66 $Y2=0.74
cc_62 VPB N_A1_c_199_n 0.0178321f $X=-0.19 $Y=1.66 $X2=2.09 $Y2=0.74
cc_63 VPB N_A1_c_200_n 0.00839819f $X=-0.19 $Y=1.66 $X2=1.635 $Y2=1.557
cc_64 VPB N_A1_c_195_n 0.0477846f $X=-0.19 $Y=1.66 $X2=1.66 $Y2=1.557
cc_65 VPB N_B1_c_269_n 0.018273f $X=-0.19 $Y=1.66 $X2=0.735 $Y2=1.765
cc_66 VPB N_B1_c_270_n 0.0146598f $X=-0.19 $Y=1.66 $X2=0.8 $Y2=1.35
cc_67 VPB N_B1_c_271_n 0.0146598f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_68 VPB N_B1_c_272_n 0.0149106f $X=-0.19 $Y=1.66 $X2=1.66 $Y2=1.35
cc_69 VPB B1 0.0134962f $X=-0.19 $Y=1.66 $X2=2.085 $Y2=2.4
cc_70 VPB N_B1_c_268_n 0.0248224f $X=-0.19 $Y=1.66 $X2=0.735 $Y2=1.557
cc_71 VPB N_C1_c_346_n 0.0147854f $X=-0.19 $Y=1.66 $X2=0.8 $Y2=0.74
cc_72 VPB N_C1_c_347_n 0.0146577f $X=-0.19 $Y=1.66 $X2=1.23 $Y2=0.74
cc_73 VPB N_C1_c_348_n 0.0146889f $X=-0.19 $Y=1.66 $X2=1.635 $Y2=1.765
cc_74 VPB N_C1_c_349_n 0.0172095f $X=-0.19 $Y=1.66 $X2=1.66 $Y2=1.35
cc_75 VPB C1 0.0102962f $X=-0.19 $Y=1.66 $X2=2.085 $Y2=2.4
cc_76 VPB N_C1_c_345_n 0.0479083f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_77 VPB N_A_77_368#_c_406_n 0.0075508f $X=-0.19 $Y=1.66 $X2=2.085 $Y2=1.765
cc_78 VPB N_A_77_368#_c_407_n 0.0360166f $X=-0.19 $Y=1.66 $X2=2.085 $Y2=2.4
cc_79 VPB N_A_77_368#_c_408_n 0.00216998f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_80 VPB N_A_77_368#_c_409_n 0.00180921f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_81 VPB N_A_77_368#_c_410_n 0.00180921f $X=-0.19 $Y=1.66 $X2=0.81 $Y2=1.515
cc_82 VPB N_A_77_368#_c_411_n 0.0110935f $X=-0.19 $Y=1.66 $X2=1.83 $Y2=1.557
cc_83 VPB N_A_77_368#_c_412_n 0.0146646f $X=-0.19 $Y=1.66 $X2=1.83 $Y2=1.515
cc_84 VPB N_A_77_368#_c_413_n 0.0126446f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_85 VPB N_VPWR_c_506_n 0.00734662f $X=-0.19 $Y=1.66 $X2=1.635 $Y2=1.765
cc_86 VPB N_VPWR_c_507_n 0.00271781f $X=-0.19 $Y=1.66 $X2=1.66 $Y2=0.74
cc_87 VPB N_VPWR_c_508_n 0.0164465f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_88 VPB N_VPWR_c_509_n 0.00261791f $X=-0.19 $Y=1.66 $X2=2.09 $Y2=1.35
cc_89 VPB N_VPWR_c_510_n 0.00329129f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_90 VPB N_VPWR_c_511_n 0.0274252f $X=-0.19 $Y=1.66 $X2=1.595 $Y2=1.58
cc_91 VPB N_VPWR_c_512_n 0.00324402f $X=-0.19 $Y=1.66 $X2=2.075 $Y2=1.58
cc_92 VPB N_VPWR_c_513_n 0.0185253f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_93 VPB N_VPWR_c_514_n 0.00601644f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_94 VPB N_VPWR_c_515_n 0.0164465f $X=-0.19 $Y=1.66 $X2=1.23 $Y2=1.557
cc_95 VPB N_VPWR_c_516_n 0.115166f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_96 VPB N_VPWR_c_505_n 0.118472f $X=-0.19 $Y=1.66 $X2=0.72 $Y2=1.565
cc_97 VPB N_VPWR_c_518_n 0.00601644f $X=-0.19 $Y=1.66 $X2=1.2 $Y2=1.565
cc_98 VPB N_VPWR_c_519_n 0.00601644f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_99 VPB N_A_901_368#_c_608_n 0.00587218f $X=-0.19 $Y=1.66 $X2=1.66 $Y2=1.35
cc_100 VPB N_A_901_368#_c_609_n 0.00213603f $X=-0.19 $Y=1.66 $X2=1.66 $Y2=0.74
cc_101 VPB N_A_901_368#_c_610_n 0.00468476f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_102 VPB N_A_901_368#_c_611_n 0.00237811f $X=-0.19 $Y=1.66 $X2=2.09 $Y2=0.74
cc_103 VPB N_A_901_368#_c_612_n 0.00213603f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_104 VPB N_A_901_368#_c_613_n 0.0120084f $X=-0.19 $Y=1.66 $X2=0.8 $Y2=1.557
cc_105 VPB N_A_901_368#_c_614_n 0.030715f $X=-0.19 $Y=1.66 $X2=1.185 $Y2=1.557
cc_106 VPB N_A_901_368#_c_615_n 0.0021839f $X=-0.19 $Y=1.66 $X2=1.635 $Y2=1.557
cc_107 VPB N_A_901_368#_c_616_n 0.00192911f $X=-0.19 $Y=1.66 $X2=1.66 $Y2=1.557
cc_108 VPB N_A_901_368#_c_617_n 0.0021839f $X=-0.19 $Y=1.66 $X2=1.83 $Y2=1.557
cc_109 VPB N_Y_c_694_n 0.0206069f $X=-0.19 $Y=1.66 $X2=0.81 $Y2=1.515
cc_110 N_A2_M1015_g N_A1_M1000_g 0.019323f $X=2.09 $Y=0.74 $X2=0 $Y2=0
cc_111 N_A2_c_119_n N_A1_c_196_n 0.00882725f $X=2.085 $Y=1.765 $X2=0 $Y2=0
cc_112 A2 N_A1_c_200_n 0.0303408f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_113 N_A2_c_115_n N_A1_c_200_n 4.0511e-19 $X=2.085 $Y=1.557 $X2=0 $Y2=0
cc_114 A2 N_A1_c_195_n 0.00346994f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_115 N_A2_c_115_n N_A1_c_195_n 0.0195417f $X=2.085 $Y=1.557 $X2=0 $Y2=0
cc_116 N_A2_c_116_n N_A_77_368#_c_406_n 4.27055e-19 $X=0.735 $Y=1.765 $X2=0
+ $Y2=0
cc_117 A2 N_A_77_368#_c_406_n 0.0265364f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_118 N_A2_c_116_n N_A_77_368#_c_407_n 0.0108977f $X=0.735 $Y=1.765 $X2=0 $Y2=0
cc_119 N_A2_c_117_n N_A_77_368#_c_407_n 6.45594e-19 $X=1.185 $Y=1.765 $X2=0
+ $Y2=0
cc_120 N_A2_c_116_n N_A_77_368#_c_418_n 0.0120074f $X=0.735 $Y=1.765 $X2=0 $Y2=0
cc_121 N_A2_c_117_n N_A_77_368#_c_418_n 0.0120074f $X=1.185 $Y=1.765 $X2=0 $Y2=0
cc_122 A2 N_A_77_368#_c_418_n 0.0393875f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_123 N_A2_c_115_n N_A_77_368#_c_418_n 0.00130859f $X=2.085 $Y=1.557 $X2=0
+ $Y2=0
cc_124 N_A2_c_116_n N_A_77_368#_c_408_n 6.47982e-19 $X=0.735 $Y=1.765 $X2=0
+ $Y2=0
cc_125 N_A2_c_117_n N_A_77_368#_c_408_n 0.0104832f $X=1.185 $Y=1.765 $X2=0 $Y2=0
cc_126 N_A2_c_118_n N_A_77_368#_c_408_n 0.00614488f $X=1.635 $Y=1.765 $X2=0
+ $Y2=0
cc_127 N_A2_c_118_n N_A_77_368#_c_425_n 0.0126853f $X=1.635 $Y=1.765 $X2=0 $Y2=0
cc_128 N_A2_c_119_n N_A_77_368#_c_425_n 0.0126853f $X=2.085 $Y=1.765 $X2=0 $Y2=0
cc_129 A2 N_A_77_368#_c_425_n 0.0477183f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_130 N_A2_c_115_n N_A_77_368#_c_425_n 0.00150005f $X=2.085 $Y=1.557 $X2=0
+ $Y2=0
cc_131 N_A2_c_119_n N_A_77_368#_c_409_n 0.00563739f $X=2.085 $Y=1.765 $X2=0
+ $Y2=0
cc_132 N_A2_c_117_n N_A_77_368#_c_430_n 4.27055e-19 $X=1.185 $Y=1.765 $X2=0
+ $Y2=0
cc_133 A2 N_A_77_368#_c_430_n 0.0193936f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_134 N_A2_c_115_n N_A_77_368#_c_430_n 0.00124229f $X=2.085 $Y=1.557 $X2=0
+ $Y2=0
cc_135 A2 N_A_77_368#_c_433_n 0.00441988f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_136 N_A2_c_116_n N_VPWR_c_506_n 0.00486623f $X=0.735 $Y=1.765 $X2=0 $Y2=0
cc_137 N_A2_c_117_n N_VPWR_c_506_n 0.00366706f $X=1.185 $Y=1.765 $X2=0 $Y2=0
cc_138 N_A2_c_117_n N_VPWR_c_507_n 5.55114e-19 $X=1.185 $Y=1.765 $X2=0 $Y2=0
cc_139 N_A2_c_118_n N_VPWR_c_507_n 0.0113491f $X=1.635 $Y=1.765 $X2=0 $Y2=0
cc_140 N_A2_c_119_n N_VPWR_c_507_n 0.0112179f $X=2.085 $Y=1.765 $X2=0 $Y2=0
cc_141 N_A2_c_119_n N_VPWR_c_508_n 0.00413917f $X=2.085 $Y=1.765 $X2=0 $Y2=0
cc_142 N_A2_c_119_n N_VPWR_c_509_n 5.35985e-19 $X=2.085 $Y=1.765 $X2=0 $Y2=0
cc_143 N_A2_c_116_n N_VPWR_c_511_n 0.00445602f $X=0.735 $Y=1.765 $X2=0 $Y2=0
cc_144 N_A2_c_117_n N_VPWR_c_513_n 0.00445602f $X=1.185 $Y=1.765 $X2=0 $Y2=0
cc_145 N_A2_c_118_n N_VPWR_c_513_n 0.00413917f $X=1.635 $Y=1.765 $X2=0 $Y2=0
cc_146 N_A2_c_116_n N_VPWR_c_505_n 0.00861635f $X=0.735 $Y=1.765 $X2=0 $Y2=0
cc_147 N_A2_c_117_n N_VPWR_c_505_n 0.00857589f $X=1.185 $Y=1.765 $X2=0 $Y2=0
cc_148 N_A2_c_118_n N_VPWR_c_505_n 0.00817726f $X=1.635 $Y=1.765 $X2=0 $Y2=0
cc_149 N_A2_c_119_n N_VPWR_c_505_n 0.0081781f $X=2.085 $Y=1.765 $X2=0 $Y2=0
cc_150 N_A2_M1004_g N_A_92_74#_c_765_n 0.00159319f $X=0.8 $Y=0.74 $X2=0 $Y2=0
cc_151 N_A2_M1004_g N_A_92_74#_c_766_n 0.0136535f $X=0.8 $Y=0.74 $X2=0 $Y2=0
cc_152 N_A2_M1005_g N_A_92_74#_c_766_n 0.0130918f $X=1.23 $Y=0.74 $X2=0 $Y2=0
cc_153 A2 N_A_92_74#_c_766_n 0.0517333f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_154 N_A2_c_115_n N_A_92_74#_c_766_n 0.00368969f $X=2.085 $Y=1.557 $X2=0 $Y2=0
cc_155 A2 N_A_92_74#_c_767_n 0.0224351f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_156 N_A2_c_115_n N_A_92_74#_c_767_n 6.38135e-19 $X=2.085 $Y=1.557 $X2=0 $Y2=0
cc_157 N_A2_M1005_g N_A_92_74#_c_768_n 3.92313e-19 $X=1.23 $Y=0.74 $X2=0 $Y2=0
cc_158 N_A2_M1013_g N_A_92_74#_c_768_n 3.92313e-19 $X=1.66 $Y=0.74 $X2=0 $Y2=0
cc_159 N_A2_M1013_g N_A_92_74#_c_769_n 0.0130453f $X=1.66 $Y=0.74 $X2=0 $Y2=0
cc_160 N_A2_M1015_g N_A_92_74#_c_769_n 0.0128967f $X=2.09 $Y=0.74 $X2=0 $Y2=0
cc_161 A2 N_A_92_74#_c_769_n 0.0568851f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_162 N_A2_c_115_n N_A_92_74#_c_769_n 0.00247712f $X=2.085 $Y=1.557 $X2=0 $Y2=0
cc_163 A2 N_A_92_74#_c_772_n 0.0146029f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_164 N_A2_c_115_n N_A_92_74#_c_772_n 0.00232957f $X=2.085 $Y=1.557 $X2=0 $Y2=0
cc_165 N_A2_M1004_g N_VGND_c_816_n 0.0137191f $X=0.8 $Y=0.74 $X2=0 $Y2=0
cc_166 N_A2_M1005_g N_VGND_c_816_n 0.0106755f $X=1.23 $Y=0.74 $X2=0 $Y2=0
cc_167 N_A2_M1013_g N_VGND_c_816_n 4.71636e-19 $X=1.66 $Y=0.74 $X2=0 $Y2=0
cc_168 N_A2_M1005_g N_VGND_c_817_n 4.71636e-19 $X=1.23 $Y=0.74 $X2=0 $Y2=0
cc_169 N_A2_M1013_g N_VGND_c_817_n 0.0106755f $X=1.66 $Y=0.74 $X2=0 $Y2=0
cc_170 N_A2_M1015_g N_VGND_c_817_n 0.0107817f $X=2.09 $Y=0.74 $X2=0 $Y2=0
cc_171 N_A2_M1004_g N_VGND_c_820_n 0.00383152f $X=0.8 $Y=0.74 $X2=0 $Y2=0
cc_172 N_A2_M1005_g N_VGND_c_822_n 0.00383152f $X=1.23 $Y=0.74 $X2=0 $Y2=0
cc_173 N_A2_M1013_g N_VGND_c_822_n 0.00383152f $X=1.66 $Y=0.74 $X2=0 $Y2=0
cc_174 N_A2_M1015_g N_VGND_c_824_n 0.00383152f $X=2.09 $Y=0.74 $X2=0 $Y2=0
cc_175 N_A2_M1004_g N_VGND_c_827_n 0.00762539f $X=0.8 $Y=0.74 $X2=0 $Y2=0
cc_176 N_A2_M1005_g N_VGND_c_827_n 0.0075754f $X=1.23 $Y=0.74 $X2=0 $Y2=0
cc_177 N_A2_M1013_g N_VGND_c_827_n 0.0075754f $X=1.66 $Y=0.74 $X2=0 $Y2=0
cc_178 N_A2_M1015_g N_VGND_c_827_n 0.00757637f $X=2.09 $Y=0.74 $X2=0 $Y2=0
cc_179 N_A1_M1025_g B1 0.00133012f $X=3.81 $Y=0.74 $X2=0 $Y2=0
cc_180 N_A1_c_199_n B1 2.30672e-19 $X=3.885 $Y=1.765 $X2=0 $Y2=0
cc_181 N_A1_c_200_n B1 0.0148046f $X=3.69 $Y=1.515 $X2=0 $Y2=0
cc_182 N_A1_c_195_n B1 0.00913805f $X=3.81 $Y=1.557 $X2=0 $Y2=0
cc_183 N_A1_c_196_n N_A_77_368#_c_409_n 0.00563739f $X=2.535 $Y=1.765 $X2=0
+ $Y2=0
cc_184 N_A1_c_196_n N_A_77_368#_c_435_n 0.0140291f $X=2.535 $Y=1.765 $X2=0 $Y2=0
cc_185 N_A1_c_197_n N_A_77_368#_c_435_n 0.0126853f $X=2.985 $Y=1.765 $X2=0 $Y2=0
cc_186 N_A1_c_200_n N_A_77_368#_c_435_n 0.0413979f $X=3.69 $Y=1.515 $X2=0 $Y2=0
cc_187 N_A1_c_195_n N_A_77_368#_c_435_n 0.00150076f $X=3.81 $Y=1.557 $X2=0 $Y2=0
cc_188 N_A1_c_197_n N_A_77_368#_c_410_n 0.00563739f $X=2.985 $Y=1.765 $X2=0
+ $Y2=0
cc_189 N_A1_c_198_n N_A_77_368#_c_410_n 0.00563739f $X=3.435 $Y=1.765 $X2=0
+ $Y2=0
cc_190 N_A1_c_198_n N_A_77_368#_c_441_n 0.0126853f $X=3.435 $Y=1.765 $X2=0 $Y2=0
cc_191 N_A1_c_199_n N_A_77_368#_c_441_n 0.015731f $X=3.885 $Y=1.765 $X2=0 $Y2=0
cc_192 N_A1_c_200_n N_A_77_368#_c_441_n 0.0370201f $X=3.69 $Y=1.515 $X2=0 $Y2=0
cc_193 N_A1_c_195_n N_A_77_368#_c_441_n 0.00150005f $X=3.81 $Y=1.557 $X2=0 $Y2=0
cc_194 N_A1_c_199_n N_A_77_368#_c_411_n 0.00729586f $X=3.885 $Y=1.765 $X2=0
+ $Y2=0
cc_195 N_A1_c_200_n N_A_77_368#_c_446_n 0.0150275f $X=3.69 $Y=1.515 $X2=0 $Y2=0
cc_196 N_A1_c_195_n N_A_77_368#_c_446_n 0.00104225f $X=3.81 $Y=1.557 $X2=0 $Y2=0
cc_197 N_A1_c_199_n N_A_77_368#_c_413_n 0.00314968f $X=3.885 $Y=1.765 $X2=0
+ $Y2=0
cc_198 N_A1_c_196_n N_VPWR_c_507_n 5.35985e-19 $X=2.535 $Y=1.765 $X2=0 $Y2=0
cc_199 N_A1_c_196_n N_VPWR_c_508_n 0.00413917f $X=2.535 $Y=1.765 $X2=0 $Y2=0
cc_200 N_A1_c_196_n N_VPWR_c_509_n 0.0112179f $X=2.535 $Y=1.765 $X2=0 $Y2=0
cc_201 N_A1_c_197_n N_VPWR_c_509_n 0.0112179f $X=2.985 $Y=1.765 $X2=0 $Y2=0
cc_202 N_A1_c_198_n N_VPWR_c_509_n 5.35985e-19 $X=3.435 $Y=1.765 $X2=0 $Y2=0
cc_203 N_A1_c_197_n N_VPWR_c_510_n 5.35985e-19 $X=2.985 $Y=1.765 $X2=0 $Y2=0
cc_204 N_A1_c_198_n N_VPWR_c_510_n 0.0112179f $X=3.435 $Y=1.765 $X2=0 $Y2=0
cc_205 N_A1_c_199_n N_VPWR_c_510_n 0.0122511f $X=3.885 $Y=1.765 $X2=0 $Y2=0
cc_206 N_A1_c_197_n N_VPWR_c_515_n 0.00413917f $X=2.985 $Y=1.765 $X2=0 $Y2=0
cc_207 N_A1_c_198_n N_VPWR_c_515_n 0.00413917f $X=3.435 $Y=1.765 $X2=0 $Y2=0
cc_208 N_A1_c_199_n N_VPWR_c_516_n 0.00413917f $X=3.885 $Y=1.765 $X2=0 $Y2=0
cc_209 N_A1_c_196_n N_VPWR_c_505_n 0.0081781f $X=2.535 $Y=1.765 $X2=0 $Y2=0
cc_210 N_A1_c_197_n N_VPWR_c_505_n 0.00817726f $X=2.985 $Y=1.765 $X2=0 $Y2=0
cc_211 N_A1_c_198_n N_VPWR_c_505_n 0.00817726f $X=3.435 $Y=1.765 $X2=0 $Y2=0
cc_212 N_A1_c_199_n N_VPWR_c_505_n 0.00822528f $X=3.885 $Y=1.765 $X2=0 $Y2=0
cc_213 N_A1_c_199_n N_A_901_368#_c_610_n 0.00177935f $X=3.885 $Y=1.765 $X2=0
+ $Y2=0
cc_214 N_A1_M1000_g N_Y_c_688_n 0.00450806f $X=2.52 $Y=0.74 $X2=0 $Y2=0
cc_215 N_A1_M1010_g N_Y_c_688_n 0.0136469f $X=2.95 $Y=0.74 $X2=0 $Y2=0
cc_216 N_A1_M1021_g N_Y_c_688_n 0.0136469f $X=3.38 $Y=0.74 $X2=0 $Y2=0
cc_217 N_A1_c_200_n N_Y_c_688_n 0.0835653f $X=3.69 $Y=1.515 $X2=0 $Y2=0
cc_218 N_A1_c_195_n N_Y_c_688_n 0.00663681f $X=3.81 $Y=1.557 $X2=0 $Y2=0
cc_219 N_A1_M1025_g N_Y_c_689_n 0.0113071f $X=3.81 $Y=0.74 $X2=0 $Y2=0
cc_220 N_A1_c_195_n N_Y_c_689_n 0.00349933f $X=3.81 $Y=1.557 $X2=0 $Y2=0
cc_221 N_A1_M1025_g N_Y_c_695_n 0.00953159f $X=3.81 $Y=0.74 $X2=0 $Y2=0
cc_222 N_A1_M1000_g N_A_92_74#_c_769_n 0.0017668f $X=2.52 $Y=0.74 $X2=0 $Y2=0
cc_223 N_A1_M1000_g N_A_92_74#_c_771_n 0.0146042f $X=2.52 $Y=0.74 $X2=0 $Y2=0
cc_224 N_A1_M1010_g N_A_92_74#_c_771_n 0.0105399f $X=2.95 $Y=0.74 $X2=0 $Y2=0
cc_225 N_A1_M1021_g N_A_92_74#_c_771_n 0.0106128f $X=3.38 $Y=0.74 $X2=0 $Y2=0
cc_226 N_A1_M1025_g N_A_92_74#_c_771_n 0.0115786f $X=3.81 $Y=0.74 $X2=0 $Y2=0
cc_227 N_A1_M1000_g N_VGND_c_817_n 6.39729e-19 $X=2.52 $Y=0.74 $X2=0 $Y2=0
cc_228 N_A1_M1000_g N_VGND_c_824_n 0.00291649f $X=2.52 $Y=0.74 $X2=0 $Y2=0
cc_229 N_A1_M1010_g N_VGND_c_824_n 0.00291649f $X=2.95 $Y=0.74 $X2=0 $Y2=0
cc_230 N_A1_M1021_g N_VGND_c_824_n 0.00291649f $X=3.38 $Y=0.74 $X2=0 $Y2=0
cc_231 N_A1_M1025_g N_VGND_c_824_n 0.00291649f $X=3.81 $Y=0.74 $X2=0 $Y2=0
cc_232 N_A1_M1000_g N_VGND_c_827_n 0.00359219f $X=2.52 $Y=0.74 $X2=0 $Y2=0
cc_233 N_A1_M1010_g N_VGND_c_827_n 0.00359121f $X=2.95 $Y=0.74 $X2=0 $Y2=0
cc_234 N_A1_M1021_g N_VGND_c_827_n 0.00359121f $X=3.38 $Y=0.74 $X2=0 $Y2=0
cc_235 N_A1_M1025_g N_VGND_c_827_n 0.0036412f $X=3.81 $Y=0.74 $X2=0 $Y2=0
cc_236 N_B1_M1020_g N_C1_M1018_g 0.0173064f $X=6.19 $Y=0.74 $X2=0 $Y2=0
cc_237 B1 N_C1_M1018_g 2.47186e-19 $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_238 N_B1_c_272_n N_C1_c_346_n 0.0126585f $X=6.205 $Y=1.765 $X2=0 $Y2=0
cc_239 B1 C1 0.0285942f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_240 N_B1_c_268_n C1 0.00420777f $X=6.19 $Y=1.532 $X2=0 $Y2=0
cc_241 B1 N_C1_c_345_n 3.05886e-19 $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_242 N_B1_c_268_n N_C1_c_345_n 0.0226518f $X=6.19 $Y=1.532 $X2=0 $Y2=0
cc_243 N_B1_c_269_n N_A_77_368#_c_411_n 0.00431037f $X=4.855 $Y=1.765 $X2=0
+ $Y2=0
cc_244 N_B1_c_269_n N_A_77_368#_c_412_n 0.0146058f $X=4.855 $Y=1.765 $X2=0 $Y2=0
cc_245 B1 N_A_77_368#_c_412_n 0.0390644f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_246 N_B1_c_269_n N_A_77_368#_c_452_n 0.00532448f $X=4.855 $Y=1.765 $X2=0
+ $Y2=0
cc_247 N_B1_c_270_n N_A_77_368#_c_452_n 0.00532448f $X=5.305 $Y=1.765 $X2=0
+ $Y2=0
cc_248 N_B1_c_270_n N_A_77_368#_c_454_n 0.0126853f $X=5.305 $Y=1.765 $X2=0 $Y2=0
cc_249 N_B1_c_271_n N_A_77_368#_c_454_n 0.0126853f $X=5.755 $Y=1.765 $X2=0 $Y2=0
cc_250 B1 N_A_77_368#_c_454_n 0.0482292f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_251 N_B1_c_268_n N_A_77_368#_c_454_n 0.00152513f $X=6.19 $Y=1.532 $X2=0 $Y2=0
cc_252 N_B1_c_272_n N_A_77_368#_c_458_n 0.00234136f $X=6.205 $Y=1.765 $X2=0
+ $Y2=0
cc_253 B1 N_A_77_368#_c_458_n 0.0177227f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_254 N_B1_c_268_n N_A_77_368#_c_458_n 0.00111367f $X=6.19 $Y=1.532 $X2=0 $Y2=0
cc_255 N_B1_c_271_n N_A_77_368#_c_461_n 0.00576017f $X=5.755 $Y=1.765 $X2=0
+ $Y2=0
cc_256 N_B1_c_272_n N_A_77_368#_c_461_n 0.00741046f $X=6.205 $Y=1.765 $X2=0
+ $Y2=0
cc_257 N_B1_c_269_n N_A_77_368#_c_413_n 0.00328692f $X=4.855 $Y=1.765 $X2=0
+ $Y2=0
cc_258 B1 N_A_77_368#_c_464_n 0.0151514f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_259 N_B1_c_268_n N_A_77_368#_c_464_n 9.40498e-19 $X=6.19 $Y=1.532 $X2=0 $Y2=0
cc_260 N_B1_c_269_n N_VPWR_c_516_n 0.00278257f $X=4.855 $Y=1.765 $X2=0 $Y2=0
cc_261 N_B1_c_270_n N_VPWR_c_516_n 0.00278257f $X=5.305 $Y=1.765 $X2=0 $Y2=0
cc_262 N_B1_c_271_n N_VPWR_c_516_n 0.00278257f $X=5.755 $Y=1.765 $X2=0 $Y2=0
cc_263 N_B1_c_272_n N_VPWR_c_516_n 0.00278271f $X=6.205 $Y=1.765 $X2=0 $Y2=0
cc_264 N_B1_c_269_n N_VPWR_c_505_n 0.00358623f $X=4.855 $Y=1.765 $X2=0 $Y2=0
cc_265 N_B1_c_270_n N_VPWR_c_505_n 0.00353822f $X=5.305 $Y=1.765 $X2=0 $Y2=0
cc_266 N_B1_c_271_n N_VPWR_c_505_n 0.00353822f $X=5.755 $Y=1.765 $X2=0 $Y2=0
cc_267 N_B1_c_272_n N_VPWR_c_505_n 0.00353907f $X=6.205 $Y=1.765 $X2=0 $Y2=0
cc_268 N_B1_c_269_n N_A_901_368#_c_608_n 0.008278f $X=4.855 $Y=1.765 $X2=0 $Y2=0
cc_269 N_B1_c_270_n N_A_901_368#_c_608_n 5.7112e-19 $X=5.305 $Y=1.765 $X2=0
+ $Y2=0
cc_270 N_B1_c_269_n N_A_901_368#_c_609_n 0.0108414f $X=4.855 $Y=1.765 $X2=0
+ $Y2=0
cc_271 N_B1_c_270_n N_A_901_368#_c_609_n 0.0108414f $X=5.305 $Y=1.765 $X2=0
+ $Y2=0
cc_272 N_B1_c_269_n N_A_901_368#_c_610_n 0.00262934f $X=4.855 $Y=1.765 $X2=0
+ $Y2=0
cc_273 N_B1_c_269_n N_A_901_368#_c_624_n 5.7112e-19 $X=4.855 $Y=1.765 $X2=0
+ $Y2=0
cc_274 N_B1_c_270_n N_A_901_368#_c_624_n 0.00830261f $X=5.305 $Y=1.765 $X2=0
+ $Y2=0
cc_275 N_B1_c_271_n N_A_901_368#_c_624_n 0.00843162f $X=5.755 $Y=1.765 $X2=0
+ $Y2=0
cc_276 N_B1_c_272_n N_A_901_368#_c_624_n 6.18425e-19 $X=6.205 $Y=1.765 $X2=0
+ $Y2=0
cc_277 N_B1_c_271_n N_A_901_368#_c_611_n 0.0108414f $X=5.755 $Y=1.765 $X2=0
+ $Y2=0
cc_278 N_B1_c_272_n N_A_901_368#_c_611_n 0.0128006f $X=6.205 $Y=1.765 $X2=0
+ $Y2=0
cc_279 N_B1_c_270_n N_A_901_368#_c_615_n 0.00175197f $X=5.305 $Y=1.765 $X2=0
+ $Y2=0
cc_280 N_B1_c_271_n N_A_901_368#_c_615_n 0.00175197f $X=5.755 $Y=1.765 $X2=0
+ $Y2=0
cc_281 B1 N_Y_c_689_n 0.0736923f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_282 N_B1_c_268_n N_Y_c_689_n 0.0150425f $X=6.19 $Y=1.532 $X2=0 $Y2=0
cc_283 N_B1_M1001_g N_Y_c_690_n 0.00159319f $X=5.76 $Y=0.74 $X2=0 $Y2=0
cc_284 N_B1_M1001_g N_Y_c_691_n 0.012695f $X=5.76 $Y=0.74 $X2=0 $Y2=0
cc_285 N_B1_M1020_g N_Y_c_691_n 0.0170429f $X=6.19 $Y=0.74 $X2=0 $Y2=0
cc_286 B1 N_Y_c_691_n 0.036928f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_287 N_B1_c_268_n N_Y_c_691_n 0.00469911f $X=6.19 $Y=1.532 $X2=0 $Y2=0
cc_288 N_B1_M1020_g N_Y_c_692_n 3.92313e-19 $X=6.19 $Y=0.74 $X2=0 $Y2=0
cc_289 B1 N_Y_c_696_n 0.0216392f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_290 N_B1_c_268_n N_Y_c_696_n 0.00584863f $X=6.19 $Y=1.532 $X2=0 $Y2=0
cc_291 N_B1_M1020_g N_Y_c_697_n 0.00158218f $X=6.19 $Y=0.74 $X2=0 $Y2=0
cc_292 N_B1_M1001_g N_VGND_c_818_n 0.0125716f $X=5.76 $Y=0.74 $X2=0 $Y2=0
cc_293 N_B1_M1020_g N_VGND_c_818_n 0.00955691f $X=6.19 $Y=0.74 $X2=0 $Y2=0
cc_294 N_B1_M1020_g N_VGND_c_819_n 4.71636e-19 $X=6.19 $Y=0.74 $X2=0 $Y2=0
cc_295 N_B1_M1001_g N_VGND_c_824_n 0.00383152f $X=5.76 $Y=0.74 $X2=0 $Y2=0
cc_296 N_B1_M1020_g N_VGND_c_825_n 0.00383152f $X=6.19 $Y=0.74 $X2=0 $Y2=0
cc_297 N_B1_M1001_g N_VGND_c_827_n 0.00762539f $X=5.76 $Y=0.74 $X2=0 $Y2=0
cc_298 N_B1_M1020_g N_VGND_c_827_n 0.00757637f $X=6.19 $Y=0.74 $X2=0 $Y2=0
cc_299 N_C1_c_346_n N_VPWR_c_516_n 0.00278257f $X=6.655 $Y=1.765 $X2=0 $Y2=0
cc_300 N_C1_c_347_n N_VPWR_c_516_n 0.00278257f $X=7.105 $Y=1.765 $X2=0 $Y2=0
cc_301 N_C1_c_348_n N_VPWR_c_516_n 0.00278257f $X=7.555 $Y=1.765 $X2=0 $Y2=0
cc_302 N_C1_c_349_n N_VPWR_c_516_n 0.00278257f $X=8.005 $Y=1.765 $X2=0 $Y2=0
cc_303 N_C1_c_346_n N_VPWR_c_505_n 0.00353905f $X=6.655 $Y=1.765 $X2=0 $Y2=0
cc_304 N_C1_c_347_n N_VPWR_c_505_n 0.00353822f $X=7.105 $Y=1.765 $X2=0 $Y2=0
cc_305 N_C1_c_348_n N_VPWR_c_505_n 0.00353822f $X=7.555 $Y=1.765 $X2=0 $Y2=0
cc_306 N_C1_c_349_n N_VPWR_c_505_n 0.00357674f $X=8.005 $Y=1.765 $X2=0 $Y2=0
cc_307 N_C1_c_346_n N_A_901_368#_c_632_n 0.0110935f $X=6.655 $Y=1.765 $X2=0
+ $Y2=0
cc_308 N_C1_c_347_n N_A_901_368#_c_632_n 6.24416e-19 $X=7.105 $Y=1.765 $X2=0
+ $Y2=0
cc_309 C1 N_A_901_368#_c_632_n 0.0175444f $X=7.355 $Y=1.58 $X2=0 $Y2=0
cc_310 N_C1_c_346_n N_A_901_368#_c_612_n 0.0108414f $X=6.655 $Y=1.765 $X2=0
+ $Y2=0
cc_311 N_C1_c_347_n N_A_901_368#_c_612_n 0.0108414f $X=7.105 $Y=1.765 $X2=0
+ $Y2=0
cc_312 N_C1_c_346_n N_A_901_368#_c_637_n 5.7112e-19 $X=6.655 $Y=1.765 $X2=0
+ $Y2=0
cc_313 N_C1_c_347_n N_A_901_368#_c_637_n 0.00766499f $X=7.105 $Y=1.765 $X2=0
+ $Y2=0
cc_314 N_C1_c_348_n N_A_901_368#_c_637_n 0.00766499f $X=7.555 $Y=1.765 $X2=0
+ $Y2=0
cc_315 N_C1_c_349_n N_A_901_368#_c_637_n 5.7112e-19 $X=8.005 $Y=1.765 $X2=0
+ $Y2=0
cc_316 N_C1_c_348_n N_A_901_368#_c_613_n 0.0108414f $X=7.555 $Y=1.765 $X2=0
+ $Y2=0
cc_317 N_C1_c_349_n N_A_901_368#_c_613_n 0.0134708f $X=8.005 $Y=1.765 $X2=0
+ $Y2=0
cc_318 N_C1_c_348_n N_A_901_368#_c_614_n 5.96501e-19 $X=7.555 $Y=1.765 $X2=0
+ $Y2=0
cc_319 N_C1_c_349_n N_A_901_368#_c_614_n 0.011822f $X=8.005 $Y=1.765 $X2=0 $Y2=0
cc_320 N_C1_c_346_n N_A_901_368#_c_616_n 0.00171731f $X=6.655 $Y=1.765 $X2=0
+ $Y2=0
cc_321 N_C1_c_347_n N_A_901_368#_c_617_n 0.00175197f $X=7.105 $Y=1.765 $X2=0
+ $Y2=0
cc_322 N_C1_c_348_n N_A_901_368#_c_617_n 0.00175197f $X=7.555 $Y=1.765 $X2=0
+ $Y2=0
cc_323 N_C1_M1018_g N_Y_c_692_n 3.92313e-19 $X=6.62 $Y=0.74 $X2=0 $Y2=0
cc_324 N_C1_M1018_g N_Y_c_693_n 0.0129459f $X=6.62 $Y=0.74 $X2=0 $Y2=0
cc_325 N_C1_M1019_g N_Y_c_693_n 0.0139042f $X=7.05 $Y=0.74 $X2=0 $Y2=0
cc_326 C1 N_Y_c_693_n 0.0519673f $X=7.355 $Y=1.58 $X2=0 $Y2=0
cc_327 N_C1_c_345_n N_Y_c_693_n 0.00386327f $X=7.555 $Y=1.542 $X2=0 $Y2=0
cc_328 N_C1_M1019_g N_Y_c_694_n 0.00528327f $X=7.05 $Y=0.74 $X2=0 $Y2=0
cc_329 N_C1_c_347_n N_Y_c_694_n 0.0126342f $X=7.105 $Y=1.765 $X2=0 $Y2=0
cc_330 N_C1_c_348_n N_Y_c_694_n 0.0251045f $X=7.555 $Y=1.765 $X2=0 $Y2=0
cc_331 N_C1_c_349_n N_Y_c_694_n 0.0152401f $X=8.005 $Y=1.765 $X2=0 $Y2=0
cc_332 C1 N_Y_c_694_n 0.10805f $X=7.355 $Y=1.58 $X2=0 $Y2=0
cc_333 N_C1_c_345_n N_Y_c_694_n 0.0671294f $X=7.555 $Y=1.542 $X2=0 $Y2=0
cc_334 C1 N_Y_c_697_n 0.011271f $X=7.355 $Y=1.58 $X2=0 $Y2=0
cc_335 N_C1_c_346_n N_Y_c_730_n 0.00222151f $X=6.655 $Y=1.765 $X2=0 $Y2=0
cc_336 N_C1_c_347_n N_Y_c_730_n 0.00497407f $X=7.105 $Y=1.765 $X2=0 $Y2=0
cc_337 C1 N_Y_c_730_n 0.0150275f $X=7.355 $Y=1.58 $X2=0 $Y2=0
cc_338 N_C1_c_345_n N_Y_c_730_n 0.00104154f $X=7.555 $Y=1.542 $X2=0 $Y2=0
cc_339 N_C1_M1018_g N_VGND_c_818_n 4.56715e-19 $X=6.62 $Y=0.74 $X2=0 $Y2=0
cc_340 N_C1_M1018_g N_VGND_c_819_n 0.0106755f $X=6.62 $Y=0.74 $X2=0 $Y2=0
cc_341 N_C1_M1019_g N_VGND_c_819_n 0.0137064f $X=7.05 $Y=0.74 $X2=0 $Y2=0
cc_342 N_C1_M1018_g N_VGND_c_825_n 0.00383152f $X=6.62 $Y=0.74 $X2=0 $Y2=0
cc_343 N_C1_M1019_g N_VGND_c_826_n 0.00383152f $X=7.05 $Y=0.74 $X2=0 $Y2=0
cc_344 N_C1_M1018_g N_VGND_c_827_n 0.00757637f $X=6.62 $Y=0.74 $X2=0 $Y2=0
cc_345 N_C1_M1019_g N_VGND_c_827_n 0.00762539f $X=7.05 $Y=0.74 $X2=0 $Y2=0
cc_346 N_A_77_368#_c_418_n N_VPWR_M1002_d 0.00408911f $X=1.245 $Y=2.035
+ $X2=-0.19 $Y2=1.66
cc_347 N_A_77_368#_c_425_n N_VPWR_M1023_d 0.00359365f $X=2.225 $Y=2.035 $X2=0
+ $Y2=0
cc_348 N_A_77_368#_c_435_n N_VPWR_M1008_d 0.00359365f $X=3.125 $Y=2.035 $X2=0
+ $Y2=0
cc_349 N_A_77_368#_c_441_n N_VPWR_M1014_d 0.00359365f $X=4.025 $Y=2.035 $X2=0
+ $Y2=0
cc_350 N_A_77_368#_c_407_n N_VPWR_c_506_n 0.0449718f $X=0.51 $Y=2.815 $X2=0
+ $Y2=0
cc_351 N_A_77_368#_c_418_n N_VPWR_c_506_n 0.0136682f $X=1.245 $Y=2.035 $X2=0
+ $Y2=0
cc_352 N_A_77_368#_c_408_n N_VPWR_c_506_n 0.0440249f $X=1.41 $Y=2.445 $X2=0
+ $Y2=0
cc_353 N_A_77_368#_c_408_n N_VPWR_c_507_n 0.0462948f $X=1.41 $Y=2.445 $X2=0
+ $Y2=0
cc_354 N_A_77_368#_c_425_n N_VPWR_c_507_n 0.0171813f $X=2.225 $Y=2.035 $X2=0
+ $Y2=0
cc_355 N_A_77_368#_c_409_n N_VPWR_c_507_n 0.0449718f $X=2.31 $Y=2.445 $X2=0
+ $Y2=0
cc_356 N_A_77_368#_c_409_n N_VPWR_c_508_n 0.00749631f $X=2.31 $Y=2.445 $X2=0
+ $Y2=0
cc_357 N_A_77_368#_c_409_n N_VPWR_c_509_n 0.0449718f $X=2.31 $Y=2.445 $X2=0
+ $Y2=0
cc_358 N_A_77_368#_c_435_n N_VPWR_c_509_n 0.0171813f $X=3.125 $Y=2.035 $X2=0
+ $Y2=0
cc_359 N_A_77_368#_c_410_n N_VPWR_c_509_n 0.0449718f $X=3.21 $Y=2.445 $X2=0
+ $Y2=0
cc_360 N_A_77_368#_c_410_n N_VPWR_c_510_n 0.0449718f $X=3.21 $Y=2.445 $X2=0
+ $Y2=0
cc_361 N_A_77_368#_c_441_n N_VPWR_c_510_n 0.0171813f $X=4.025 $Y=2.035 $X2=0
+ $Y2=0
cc_362 N_A_77_368#_c_411_n N_VPWR_c_510_n 0.0462948f $X=4.11 $Y=2.4 $X2=0 $Y2=0
cc_363 N_A_77_368#_c_407_n N_VPWR_c_511_n 0.0145938f $X=0.51 $Y=2.815 $X2=0
+ $Y2=0
cc_364 N_A_77_368#_c_408_n N_VPWR_c_513_n 0.0110241f $X=1.41 $Y=2.445 $X2=0
+ $Y2=0
cc_365 N_A_77_368#_c_410_n N_VPWR_c_515_n 0.00749631f $X=3.21 $Y=2.445 $X2=0
+ $Y2=0
cc_366 N_A_77_368#_c_411_n N_VPWR_c_516_n 0.011066f $X=4.11 $Y=2.4 $X2=0 $Y2=0
cc_367 N_A_77_368#_c_407_n N_VPWR_c_505_n 0.0120466f $X=0.51 $Y=2.815 $X2=0
+ $Y2=0
cc_368 N_A_77_368#_c_408_n N_VPWR_c_505_n 0.00909194f $X=1.41 $Y=2.445 $X2=0
+ $Y2=0
cc_369 N_A_77_368#_c_409_n N_VPWR_c_505_n 0.0062048f $X=2.31 $Y=2.445 $X2=0
+ $Y2=0
cc_370 N_A_77_368#_c_410_n N_VPWR_c_505_n 0.0062048f $X=3.21 $Y=2.445 $X2=0
+ $Y2=0
cc_371 N_A_77_368#_c_411_n N_VPWR_c_505_n 0.00915947f $X=4.11 $Y=2.4 $X2=0 $Y2=0
cc_372 N_A_77_368#_c_412_n N_A_901_368#_M1017_s 0.0055238f $X=4.995 $Y=2.035
+ $X2=-0.19 $Y2=1.66
cc_373 N_A_77_368#_c_454_n N_A_901_368#_M1022_s 0.00362653f $X=5.895 $Y=2.035
+ $X2=0 $Y2=0
cc_374 N_A_77_368#_c_411_n N_A_901_368#_c_608_n 0.0463434f $X=4.11 $Y=2.4 $X2=0
+ $Y2=0
cc_375 N_A_77_368#_c_412_n N_A_901_368#_c_608_n 0.0220544f $X=4.995 $Y=2.035
+ $X2=0 $Y2=0
cc_376 N_A_77_368#_c_452_n N_A_901_368#_c_608_n 0.0289859f $X=5.08 $Y=2.57 $X2=0
+ $Y2=0
cc_377 N_A_77_368#_M1017_d N_A_901_368#_c_609_n 0.00247267f $X=4.93 $Y=1.84
+ $X2=0 $Y2=0
cc_378 N_A_77_368#_c_452_n N_A_901_368#_c_609_n 0.012787f $X=5.08 $Y=2.57 $X2=0
+ $Y2=0
cc_379 N_A_77_368#_c_411_n N_A_901_368#_c_610_n 0.00601305f $X=4.11 $Y=2.4 $X2=0
+ $Y2=0
cc_380 N_A_77_368#_c_452_n N_A_901_368#_c_624_n 0.0289859f $X=5.08 $Y=2.57 $X2=0
+ $Y2=0
cc_381 N_A_77_368#_c_454_n N_A_901_368#_c_624_n 0.0171814f $X=5.895 $Y=2.035
+ $X2=0 $Y2=0
cc_382 N_A_77_368#_c_461_n N_A_901_368#_c_624_n 0.0298377f $X=5.98 $Y=2.57 $X2=0
+ $Y2=0
cc_383 N_A_77_368#_M1024_d N_A_901_368#_c_611_n 0.00222494f $X=5.83 $Y=1.84
+ $X2=0 $Y2=0
cc_384 N_A_77_368#_c_461_n N_A_901_368#_c_611_n 0.0144323f $X=5.98 $Y=2.57 $X2=0
+ $Y2=0
cc_385 N_VPWR_c_516_n N_A_901_368#_c_609_n 0.03588f $X=8.4 $Y=3.33 $X2=0 $Y2=0
cc_386 N_VPWR_c_505_n N_A_901_368#_c_609_n 0.0201952f $X=8.4 $Y=3.33 $X2=0 $Y2=0
cc_387 N_VPWR_c_510_n N_A_901_368#_c_610_n 0.00293437f $X=3.66 $Y=2.41 $X2=0
+ $Y2=0
cc_388 N_VPWR_c_516_n N_A_901_368#_c_610_n 0.0236039f $X=8.4 $Y=3.33 $X2=0 $Y2=0
cc_389 N_VPWR_c_505_n N_A_901_368#_c_610_n 0.012761f $X=8.4 $Y=3.33 $X2=0 $Y2=0
cc_390 N_VPWR_c_516_n N_A_901_368#_c_611_n 0.0390543f $X=8.4 $Y=3.33 $X2=0 $Y2=0
cc_391 N_VPWR_c_505_n N_A_901_368#_c_611_n 0.0220062f $X=8.4 $Y=3.33 $X2=0 $Y2=0
cc_392 N_VPWR_c_516_n N_A_901_368#_c_612_n 0.03588f $X=8.4 $Y=3.33 $X2=0 $Y2=0
cc_393 N_VPWR_c_505_n N_A_901_368#_c_612_n 0.0201952f $X=8.4 $Y=3.33 $X2=0 $Y2=0
cc_394 N_VPWR_c_516_n N_A_901_368#_c_613_n 0.0594839f $X=8.4 $Y=3.33 $X2=0 $Y2=0
cc_395 N_VPWR_c_505_n N_A_901_368#_c_613_n 0.0329562f $X=8.4 $Y=3.33 $X2=0 $Y2=0
cc_396 N_VPWR_c_516_n N_A_901_368#_c_615_n 0.0235512f $X=8.4 $Y=3.33 $X2=0 $Y2=0
cc_397 N_VPWR_c_505_n N_A_901_368#_c_615_n 0.0126924f $X=8.4 $Y=3.33 $X2=0 $Y2=0
cc_398 N_VPWR_c_516_n N_A_901_368#_c_616_n 0.0200196f $X=8.4 $Y=3.33 $X2=0 $Y2=0
cc_399 N_VPWR_c_505_n N_A_901_368#_c_616_n 0.0108171f $X=8.4 $Y=3.33 $X2=0 $Y2=0
cc_400 N_VPWR_c_516_n N_A_901_368#_c_617_n 0.0235512f $X=8.4 $Y=3.33 $X2=0 $Y2=0
cc_401 N_VPWR_c_505_n N_A_901_368#_c_617_n 0.0126924f $X=8.4 $Y=3.33 $X2=0 $Y2=0
cc_402 N_A_901_368#_c_612_n N_Y_M1003_d 0.00247267f $X=7.165 $Y=2.99 $X2=0 $Y2=0
cc_403 N_A_901_368#_c_613_n N_Y_M1009_d 0.00222494f $X=8.065 $Y=2.99 $X2=0 $Y2=0
cc_404 N_A_901_368#_M1007_s N_Y_c_694_n 0.00359365f $X=7.18 $Y=1.84 $X2=0 $Y2=0
cc_405 N_A_901_368#_M1012_s N_Y_c_694_n 0.00290367f $X=8.08 $Y=1.84 $X2=0 $Y2=0
cc_406 N_A_901_368#_c_637_n N_Y_c_694_n 0.0465206f $X=7.33 $Y=2.455 $X2=0 $Y2=0
cc_407 N_A_901_368#_c_613_n N_Y_c_694_n 0.013472f $X=8.065 $Y=2.99 $X2=0 $Y2=0
cc_408 N_A_901_368#_c_614_n N_Y_c_694_n 0.0244523f $X=8.23 $Y=2.285 $X2=0 $Y2=0
cc_409 N_A_901_368#_c_632_n N_Y_c_730_n 0.0517654f $X=6.43 $Y=2.115 $X2=0 $Y2=0
cc_410 N_A_901_368#_c_612_n N_Y_c_730_n 0.012787f $X=7.165 $Y=2.99 $X2=0 $Y2=0
cc_411 N_A_901_368#_c_637_n N_Y_c_730_n 0.0289859f $X=7.33 $Y=2.455 $X2=0 $Y2=0
cc_412 N_Y_c_688_n N_A_92_74#_M1010_d 0.00177483f $X=3.588 $Y=0.957 $X2=0 $Y2=0
cc_413 N_Y_c_689_n N_A_92_74#_M1025_d 0.00425265f $X=5.38 $Y=1.045 $X2=0 $Y2=0
cc_414 N_Y_c_688_n N_A_92_74#_c_769_n 0.00561736f $X=3.588 $Y=0.957 $X2=0 $Y2=0
cc_415 N_Y_M1000_s N_A_92_74#_c_771_n 0.00179328f $X=2.595 $Y=0.37 $X2=0 $Y2=0
cc_416 N_Y_M1021_s N_A_92_74#_c_771_n 0.00179328f $X=3.455 $Y=0.37 $X2=0 $Y2=0
cc_417 N_Y_c_688_n N_A_92_74#_c_771_n 0.0630655f $X=3.588 $Y=0.957 $X2=0 $Y2=0
cc_418 N_Y_c_689_n N_A_92_74#_c_771_n 0.0160707f $X=5.38 $Y=1.045 $X2=0 $Y2=0
cc_419 N_Y_c_691_n N_VGND_M1001_s 0.00176461f $X=6.32 $Y=1.045 $X2=0 $Y2=0
cc_420 N_Y_c_693_n N_VGND_M1018_d 0.00176461f $X=7.18 $Y=1.095 $X2=0 $Y2=0
cc_421 N_Y_c_690_n N_VGND_c_818_n 0.0164982f $X=5.545 $Y=0.515 $X2=0 $Y2=0
cc_422 N_Y_c_691_n N_VGND_c_818_n 0.0170777f $X=6.32 $Y=1.045 $X2=0 $Y2=0
cc_423 N_Y_c_692_n N_VGND_c_818_n 0.0164567f $X=6.405 $Y=0.515 $X2=0 $Y2=0
cc_424 N_Y_c_692_n N_VGND_c_819_n 0.0182488f $X=6.405 $Y=0.515 $X2=0 $Y2=0
cc_425 N_Y_c_693_n N_VGND_c_819_n 0.0170777f $X=7.18 $Y=1.095 $X2=0 $Y2=0
cc_426 N_Y_c_694_n N_VGND_c_819_n 0.0184913f $X=7.695 $Y=2.035 $X2=0 $Y2=0
cc_427 N_Y_c_690_n N_VGND_c_824_n 0.011066f $X=5.545 $Y=0.515 $X2=0 $Y2=0
cc_428 N_Y_c_692_n N_VGND_c_825_n 0.00749631f $X=6.405 $Y=0.515 $X2=0 $Y2=0
cc_429 N_Y_c_694_n N_VGND_c_826_n 0.0595689f $X=7.695 $Y=2.035 $X2=0 $Y2=0
cc_430 N_Y_c_690_n N_VGND_c_827_n 0.00915947f $X=5.545 $Y=0.515 $X2=0 $Y2=0
cc_431 N_Y_c_692_n N_VGND_c_827_n 0.0062048f $X=6.405 $Y=0.515 $X2=0 $Y2=0
cc_432 N_Y_c_694_n N_VGND_c_827_n 0.049306f $X=7.695 $Y=2.035 $X2=0 $Y2=0
cc_433 N_A_92_74#_c_766_n N_VGND_M1004_d 0.00176461f $X=1.36 $Y=1.095 $X2=-0.19
+ $Y2=-0.245
cc_434 N_A_92_74#_c_769_n N_VGND_M1013_d 0.00176461f $X=2.22 $Y=1.095 $X2=0
+ $Y2=0
cc_435 N_A_92_74#_c_765_n N_VGND_c_816_n 0.0182902f $X=0.585 $Y=0.515 $X2=0
+ $Y2=0
cc_436 N_A_92_74#_c_766_n N_VGND_c_816_n 0.0170777f $X=1.36 $Y=1.095 $X2=0 $Y2=0
cc_437 N_A_92_74#_c_768_n N_VGND_c_816_n 0.0182488f $X=1.445 $Y=0.515 $X2=0
+ $Y2=0
cc_438 N_A_92_74#_c_768_n N_VGND_c_817_n 0.0182488f $X=1.445 $Y=0.515 $X2=0
+ $Y2=0
cc_439 N_A_92_74#_c_769_n N_VGND_c_817_n 0.0170777f $X=2.22 $Y=1.095 $X2=0 $Y2=0
cc_440 N_A_92_74#_c_770_n N_VGND_c_817_n 0.0103909f $X=2.305 $Y=0.615 $X2=0
+ $Y2=0
cc_441 N_A_92_74#_c_765_n N_VGND_c_820_n 0.011066f $X=0.585 $Y=0.515 $X2=0 $Y2=0
cc_442 N_A_92_74#_c_768_n N_VGND_c_822_n 0.00749631f $X=1.445 $Y=0.515 $X2=0
+ $Y2=0
cc_443 N_A_92_74#_c_770_n N_VGND_c_824_n 0.00758556f $X=2.305 $Y=0.615 $X2=0
+ $Y2=0
cc_444 N_A_92_74#_c_771_n N_VGND_c_824_n 0.0732318f $X=4.025 $Y=0.515 $X2=0
+ $Y2=0
cc_445 N_A_92_74#_c_765_n N_VGND_c_827_n 0.00915947f $X=0.585 $Y=0.515 $X2=0
+ $Y2=0
cc_446 N_A_92_74#_c_768_n N_VGND_c_827_n 0.0062048f $X=1.445 $Y=0.515 $X2=0
+ $Y2=0
cc_447 N_A_92_74#_c_770_n N_VGND_c_827_n 0.00627867f $X=2.305 $Y=0.615 $X2=0
+ $Y2=0
cc_448 N_A_92_74#_c_771_n N_VGND_c_827_n 0.0615843f $X=4.025 $Y=0.515 $X2=0
+ $Y2=0
