* File: sky130_fd_sc_hs__o22ai_4.pxi.spice
* Created: Thu Aug 27 21:00:43 2020
* 
x_PM_SKY130_FD_SC_HS__O22AI_4%A1 N_A1_M1000_g N_A1_c_125_n N_A1_M1005_g
+ N_A1_c_126_n N_A1_M1006_g N_A1_M1011_g N_A1_M1025_g N_A1_c_127_n N_A1_M1007_g
+ N_A1_c_120_n N_A1_M1017_g N_A1_M1029_g N_A1_c_122_n N_A1_c_130_n N_A1_c_123_n
+ A1 A1 N_A1_c_124_n N_A1_c_133_n N_A1_c_134_n PM_SKY130_FD_SC_HS__O22AI_4%A1
x_PM_SKY130_FD_SC_HS__O22AI_4%A2 N_A2_c_249_n N_A2_M1008_g N_A2_c_243_n
+ N_A2_M1002_g N_A2_c_244_n N_A2_M1004_g N_A2_c_250_n N_A2_M1009_g N_A2_c_245_n
+ N_A2_M1020_g N_A2_c_251_n N_A2_M1010_g N_A2_c_252_n N_A2_M1014_g N_A2_c_246_n
+ N_A2_M1031_g A2 A2 A2 N_A2_c_248_n PM_SKY130_FD_SC_HS__O22AI_4%A2
x_PM_SKY130_FD_SC_HS__O22AI_4%B1 N_B1_M1003_g N_B1_c_341_n N_B1_M1001_g
+ N_B1_c_342_n N_B1_M1012_g N_B1_M1016_g N_B1_c_343_n N_B1_M1015_g N_B1_M1023_g
+ N_B1_c_334_n N_B1_M1024_g N_B1_c_335_n N_B1_M1028_g N_B1_c_336_n N_B1_c_337_n
+ N_B1_c_338_n B1 N_B1_c_339_n N_B1_c_340_n PM_SKY130_FD_SC_HS__O22AI_4%B1
x_PM_SKY130_FD_SC_HS__O22AI_4%B2 N_B2_M1013_g N_B2_c_457_n N_B2_M1018_g
+ N_B2_M1019_g N_B2_c_458_n N_B2_M1022_g N_B2_M1021_g N_B2_c_459_n N_B2_M1027_g
+ N_B2_c_460_n N_B2_M1030_g N_B2_M1026_g B2 B2 N_B2_c_461_n N_B2_c_456_n
+ N_B2_c_463_n N_B2_c_483_n PM_SKY130_FD_SC_HS__O22AI_4%B2
x_PM_SKY130_FD_SC_HS__O22AI_4%VPWR N_VPWR_M1005_d N_VPWR_M1006_d N_VPWR_M1017_d
+ N_VPWR_M1012_d N_VPWR_M1024_d N_VPWR_c_540_n N_VPWR_c_541_n N_VPWR_c_542_n
+ N_VPWR_c_543_n N_VPWR_c_544_n N_VPWR_c_545_n N_VPWR_c_546_n VPWR
+ N_VPWR_c_547_n N_VPWR_c_548_n N_VPWR_c_549_n N_VPWR_c_550_n N_VPWR_c_551_n
+ N_VPWR_c_552_n N_VPWR_c_553_n N_VPWR_c_539_n PM_SKY130_FD_SC_HS__O22AI_4%VPWR
x_PM_SKY130_FD_SC_HS__O22AI_4%A_117_368# N_A_117_368#_M1005_s
+ N_A_117_368#_M1007_s N_A_117_368#_M1009_d N_A_117_368#_M1014_d
+ N_A_117_368#_c_636_n N_A_117_368#_c_645_n N_A_117_368#_c_649_n
+ N_A_117_368#_c_652_n N_A_117_368#_c_637_n N_A_117_368#_c_638_n
+ N_A_117_368#_c_639_n PM_SKY130_FD_SC_HS__O22AI_4%A_117_368#
x_PM_SKY130_FD_SC_HS__O22AI_4%Y N_Y_M1003_s N_Y_M1023_s N_Y_M1019_s N_Y_M1026_s
+ N_Y_M1008_s N_Y_M1010_s N_Y_M1018_s N_Y_M1027_s N_Y_c_695_n N_Y_c_700_n
+ N_Y_c_715_n N_Y_c_701_n N_Y_c_746_n N_Y_c_691_n N_Y_c_687_n N_Y_c_688_n
+ N_Y_c_703_n N_Y_c_729_n N_Y_c_731_n N_Y_c_760_n N_Y_c_735_n N_Y_c_767_n
+ N_Y_c_736_n Y Y N_Y_c_689_n Y N_Y_c_690_n PM_SKY130_FD_SC_HS__O22AI_4%Y
x_PM_SKY130_FD_SC_HS__O22AI_4%A_877_368# N_A_877_368#_M1001_s
+ N_A_877_368#_M1015_s N_A_877_368#_M1022_d N_A_877_368#_M1030_d
+ N_A_877_368#_c_835_n N_A_877_368#_c_869_n N_A_877_368#_c_843_n
+ N_A_877_368#_c_829_n N_A_877_368#_c_830_n N_A_877_368#_c_874_n
+ N_A_877_368#_c_831_n N_A_877_368#_c_839_n N_A_877_368#_c_832_n
+ N_A_877_368#_c_833_n PM_SKY130_FD_SC_HS__O22AI_4%A_877_368#
x_PM_SKY130_FD_SC_HS__O22AI_4%A_27_74# N_A_27_74#_M1000_d N_A_27_74#_M1011_d
+ N_A_27_74#_M1002_d N_A_27_74#_M1020_d N_A_27_74#_M1029_d N_A_27_74#_M1016_d
+ N_A_27_74#_M1013_d N_A_27_74#_M1021_d N_A_27_74#_M1028_d N_A_27_74#_c_883_n
+ N_A_27_74#_c_884_n N_A_27_74#_c_885_n N_A_27_74#_c_886_n N_A_27_74#_c_907_n
+ N_A_27_74#_c_887_n N_A_27_74#_c_923_n N_A_27_74#_c_888_n N_A_27_74#_c_889_n
+ N_A_27_74#_c_890_n N_A_27_74#_c_913_n N_A_27_74#_c_891_n N_A_27_74#_c_892_n
+ N_A_27_74#_c_932_n N_A_27_74#_c_935_n N_A_27_74#_c_893_n N_A_27_74#_c_894_n
+ N_A_27_74#_c_895_n N_A_27_74#_c_896_n N_A_27_74#_c_897_n
+ PM_SKY130_FD_SC_HS__O22AI_4%A_27_74#
x_PM_SKY130_FD_SC_HS__O22AI_4%VGND N_VGND_M1000_s N_VGND_M1025_s N_VGND_M1004_s
+ N_VGND_M1031_s N_VGND_c_1009_n N_VGND_c_1010_n N_VGND_c_1011_n N_VGND_c_1012_n
+ VGND N_VGND_c_1013_n N_VGND_c_1014_n N_VGND_c_1015_n N_VGND_c_1016_n
+ N_VGND_c_1017_n N_VGND_c_1018_n N_VGND_c_1019_n N_VGND_c_1020_n
+ N_VGND_c_1021_n N_VGND_c_1022_n PM_SKY130_FD_SC_HS__O22AI_4%VGND
cc_1 VNB N_A1_M1000_g 0.0318055f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_2 VNB N_A1_M1011_g 0.0221345f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=0.74
cc_3 VNB N_A1_M1025_g 0.023347f $X=-0.19 $Y=-0.245 $X2=1.425 $Y2=0.74
cc_4 VNB N_A1_c_120_n 0.0233052f $X=-0.19 $Y=-0.245 $X2=3.76 $Y2=1.765
cc_5 VNB N_A1_M1029_g 0.0256089f $X=-0.19 $Y=-0.245 $X2=3.855 $Y2=0.74
cc_6 VNB N_A1_c_122_n 5.80078e-19 $X=-0.19 $Y=-0.245 $X2=1.38 $Y2=1.485
cc_7 VNB N_A1_c_123_n 0.00755711f $X=-0.19 $Y=-0.245 $X2=3.805 $Y2=1.515
cc_8 VNB N_A1_c_124_n 0.0908218f $X=-0.19 $Y=-0.245 $X2=1.425 $Y2=1.542
cc_9 VNB N_A2_c_243_n 0.0171512f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A2_c_244_n 0.0173859f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=2.4
cc_11 VNB N_A2_c_245_n 0.0172061f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=0.74
cc_12 VNB N_A2_c_246_n 0.0187428f $X=-0.19 $Y=-0.245 $X2=3.76 $Y2=1.765
cc_13 VNB A2 0.00911391f $X=-0.19 $Y=-0.245 $X2=3.855 $Y2=0.74
cc_14 VNB N_A2_c_248_n 0.112625f $X=-0.19 $Y=-0.245 $X2=3.805 $Y2=1.515
cc_15 VNB N_B1_M1003_g 0.0213686f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_16 VNB N_B1_M1016_g 0.0209615f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=0.74
cc_17 VNB N_B1_M1023_g 0.0206172f $X=-0.19 $Y=-0.245 $X2=1.46 $Y2=2.4
cc_18 VNB N_B1_c_334_n 0.0414793f $X=-0.19 $Y=-0.245 $X2=3.76 $Y2=1.765
cc_19 VNB N_B1_c_335_n 0.0197466f $X=-0.19 $Y=-0.245 $X2=3.855 $Y2=1.35
cc_20 VNB N_B1_c_336_n 0.00305806f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_B1_c_337_n 0.0164724f $X=-0.19 $Y=-0.245 $X2=3.64 $Y2=1.805
cc_22 VNB N_B1_c_338_n 0.00320503f $X=-0.19 $Y=-0.245 $X2=1.465 $Y2=1.485
cc_23 VNB N_B1_c_339_n 0.07386f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.542
cc_24 VNB N_B1_c_340_n 0.00417394f $X=-0.19 $Y=-0.245 $X2=0.96 $Y2=1.542
cc_25 VNB N_B2_M1013_g 0.0212007f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_26 VNB N_B2_M1019_g 0.0225267f $X=-0.19 $Y=-0.245 $X2=0.96 $Y2=2.4
cc_27 VNB N_B2_M1021_g 0.0235253f $X=-0.19 $Y=-0.245 $X2=1.425 $Y2=0.74
cc_28 VNB N_B2_M1026_g 0.02313f $X=-0.19 $Y=-0.245 $X2=3.855 $Y2=0.74
cc_29 VNB N_B2_c_456_n 0.0725265f $X=-0.19 $Y=-0.245 $X2=2.555 $Y2=1.95
cc_30 VNB N_VPWR_c_539_n 0.342803f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_Y_c_687_n 0.00775967f $X=-0.19 $Y=-0.245 $X2=3.805 $Y2=1.805
cc_32 VNB N_Y_c_688_n 0.0327392f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_Y_c_689_n 0.00340136f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_Y_c_690_n 0.00141707f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_27_74#_c_883_n 0.0265694f $X=-0.19 $Y=-0.245 $X2=0.705 $Y2=1.485
cc_36 VNB N_A_27_74#_c_884_n 0.00324652f $X=-0.19 $Y=-0.245 $X2=0.705 $Y2=1.485
cc_37 VNB N_A_27_74#_c_885_n 0.0138252f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_27_74#_c_886_n 0.00206666f $X=-0.19 $Y=-0.245 $X2=3.64 $Y2=1.805
cc_39 VNB N_A_27_74#_c_887_n 0.00206561f $X=-0.19 $Y=-0.245 $X2=1.465 $Y2=1.805
cc_40 VNB N_A_27_74#_c_888_n 0.00253097f $X=-0.19 $Y=-0.245 $X2=2.555 $Y2=1.95
cc_41 VNB N_A_27_74#_c_889_n 0.0104547f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_27_74#_c_890_n 0.00211111f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.542
cc_43 VNB N_A_27_74#_c_891_n 0.00757463f $X=-0.19 $Y=-0.245 $X2=0.705 $Y2=1.542
cc_44 VNB N_A_27_74#_c_892_n 0.00184947f $X=-0.19 $Y=-0.245 $X2=3.12 $Y2=1.935
cc_45 VNB N_A_27_74#_c_893_n 9.8643e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_A_27_74#_c_894_n 0.00281291f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_27_74#_c_895_n 0.00219607f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_27_74#_c_896_n 0.0155228f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A_27_74#_c_897_n 0.00288497f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_VGND_c_1009_n 0.00578139f $X=-0.19 $Y=-0.245 $X2=1.425 $Y2=1.32
cc_51 VNB N_VGND_c_1010_n 0.00494723f $X=-0.19 $Y=-0.245 $X2=1.46 $Y2=1.765
cc_52 VNB N_VGND_c_1011_n 0.00494723f $X=-0.19 $Y=-0.245 $X2=3.76 $Y2=2.4
cc_53 VNB N_VGND_c_1012_n 0.00851143f $X=-0.19 $Y=-0.245 $X2=3.855 $Y2=0.74
cc_54 VNB N_VGND_c_1013_n 0.0191515f $X=-0.19 $Y=-0.245 $X2=0.705 $Y2=1.485
cc_55 VNB N_VGND_c_1014_n 0.0169342f $X=-0.19 $Y=-0.245 $X2=3.64 $Y2=1.805
cc_56 VNB N_VGND_c_1015_n 0.0169342f $X=-0.19 $Y=-0.245 $X2=1.385 $Y2=1.485
cc_57 VNB N_VGND_c_1016_n 0.016883f $X=-0.19 $Y=-0.245 $X2=3.805 $Y2=1.515
cc_58 VNB N_VGND_c_1017_n 0.10275f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=1.542
cc_59 VNB N_VGND_c_1018_n 0.42396f $X=-0.19 $Y=-0.245 $X2=1.385 $Y2=1.542
cc_60 VNB N_VGND_c_1019_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=3.805 $Y2=1.515
cc_61 VNB N_VGND_c_1020_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_VGND_c_1021_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=3.235 $Y2=1.935
cc_63 VNB N_VGND_c_1022_n 0.00634377f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VPB N_A1_c_125_n 0.0176575f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=1.765
cc_65 VPB N_A1_c_126_n 0.0153793f $X=-0.19 $Y=1.66 $X2=0.96 $Y2=1.765
cc_66 VPB N_A1_c_127_n 0.0155121f $X=-0.19 $Y=1.66 $X2=1.46 $Y2=1.765
cc_67 VPB N_A1_c_120_n 0.0275121f $X=-0.19 $Y=1.66 $X2=3.76 $Y2=1.765
cc_68 VPB N_A1_c_122_n 9.45824e-19 $X=-0.19 $Y=1.66 $X2=1.38 $Y2=1.485
cc_69 VPB N_A1_c_130_n 0.0082105f $X=-0.19 $Y=1.66 $X2=3.64 $Y2=1.805
cc_70 VPB N_A1_c_123_n 0.0028448f $X=-0.19 $Y=1.66 $X2=3.805 $Y2=1.515
cc_71 VPB N_A1_c_124_n 0.0230649f $X=-0.19 $Y=1.66 $X2=1.425 $Y2=1.542
cc_72 VPB N_A1_c_133_n 0.0121284f $X=-0.19 $Y=1.66 $X2=2.525 $Y2=1.935
cc_73 VPB N_A1_c_134_n 0.00422601f $X=-0.19 $Y=1.66 $X2=3.235 $Y2=1.935
cc_74 VPB N_A2_c_249_n 0.0154584f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.32
cc_75 VPB N_A2_c_250_n 0.0152892f $X=-0.19 $Y=1.66 $X2=0.96 $Y2=2.4
cc_76 VPB N_A2_c_251_n 0.0149042f $X=-0.19 $Y=1.66 $X2=1.425 $Y2=0.74
cc_77 VPB N_A2_c_252_n 0.015079f $X=-0.19 $Y=1.66 $X2=1.46 $Y2=1.765
cc_78 VPB N_A2_c_248_n 0.0248721f $X=-0.19 $Y=1.66 $X2=3.805 $Y2=1.515
cc_79 VPB N_B1_c_341_n 0.0166048f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=1.765
cc_80 VPB N_B1_c_342_n 0.0156204f $X=-0.19 $Y=1.66 $X2=0.96 $Y2=1.765
cc_81 VPB N_B1_c_343_n 0.0157536f $X=-0.19 $Y=1.66 $X2=1.425 $Y2=1.32
cc_82 VPB N_B1_c_334_n 0.0240018f $X=-0.19 $Y=1.66 $X2=3.76 $Y2=1.765
cc_83 VPB N_B1_c_339_n 0.019837f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.542
cc_84 VPB N_B2_c_457_n 0.0152881f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=1.765
cc_85 VPB N_B2_c_458_n 0.0147686f $X=-0.19 $Y=1.66 $X2=0.995 $Y2=0.74
cc_86 VPB N_B2_c_459_n 0.0147442f $X=-0.19 $Y=1.66 $X2=1.46 $Y2=1.765
cc_87 VPB N_B2_c_460_n 0.0151692f $X=-0.19 $Y=1.66 $X2=3.76 $Y2=1.765
cc_88 VPB N_B2_c_461_n 0.00286486f $X=-0.19 $Y=1.66 $X2=3.805 $Y2=1.805
cc_89 VPB N_B2_c_456_n 0.0483549f $X=-0.19 $Y=1.66 $X2=2.555 $Y2=1.95
cc_90 VPB N_B2_c_463_n 0.00295096f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_91 VPB N_VPWR_c_540_n 0.0108116f $X=-0.19 $Y=1.66 $X2=1.425 $Y2=0.74
cc_92 VPB N_VPWR_c_541_n 0.0580724f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_93 VPB N_VPWR_c_542_n 0.00593699f $X=-0.19 $Y=1.66 $X2=3.76 $Y2=2.4
cc_94 VPB N_VPWR_c_543_n 0.00969839f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_95 VPB N_VPWR_c_544_n 0.00571271f $X=-0.19 $Y=1.66 $X2=0.705 $Y2=1.485
cc_96 VPB N_VPWR_c_545_n 0.0136226f $X=-0.19 $Y=1.66 $X2=2.525 $Y2=1.805
cc_97 VPB N_VPWR_c_546_n 0.0384779f $X=-0.19 $Y=1.66 $X2=3.64 $Y2=1.805
cc_98 VPB N_VPWR_c_547_n 0.0182909f $X=-0.19 $Y=1.66 $X2=1.385 $Y2=1.485
cc_99 VPB N_VPWR_c_548_n 0.0631261f $X=-0.19 $Y=1.66 $X2=3.805 $Y2=1.515
cc_100 VPB N_VPWR_c_549_n 0.0196495f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=1.542
cc_101 VPB N_VPWR_c_550_n 0.0588051f $X=-0.19 $Y=1.66 $X2=1.425 $Y2=1.542
cc_102 VPB N_VPWR_c_551_n 0.00614127f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_103 VPB N_VPWR_c_552_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_104 VPB N_VPWR_c_553_n 0.00460249f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_105 VPB N_VPWR_c_539_n 0.0871957f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_106 VPB N_A_117_368#_c_636_n 0.00243101f $X=-0.19 $Y=1.66 $X2=1.425 $Y2=1.32
cc_107 VPB N_A_117_368#_c_637_n 0.00257348f $X=-0.19 $Y=1.66 $X2=1.46 $Y2=2.4
cc_108 VPB N_A_117_368#_c_638_n 0.0105922f $X=-0.19 $Y=1.66 $X2=3.855 $Y2=1.35
cc_109 VPB N_A_117_368#_c_639_n 0.00183343f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_110 VPB N_Y_c_691_n 0.0105186f $X=-0.19 $Y=1.66 $X2=3.805 $Y2=1.515
cc_111 VPB N_Y_c_688_n 0.0132318f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_112 VPB N_A_877_368#_c_829_n 0.0030474f $X=-0.19 $Y=1.66 $X2=1.46 $Y2=1.765
cc_113 VPB N_A_877_368#_c_830_n 0.00302802f $X=-0.19 $Y=1.66 $X2=1.46 $Y2=2.4
cc_114 VPB N_A_877_368#_c_831_n 0.0051269f $X=-0.19 $Y=1.66 $X2=3.855 $Y2=1.35
cc_115 VPB N_A_877_368#_c_832_n 0.00257348f $X=-0.19 $Y=1.66 $X2=0.705 $Y2=1.485
cc_116 VPB N_A_877_368#_c_833_n 0.00123754f $X=-0.19 $Y=1.66 $X2=1.55 $Y2=1.805
cc_117 N_A1_c_127_n N_A2_c_249_n 0.0256164f $X=1.46 $Y=1.765 $X2=-0.19
+ $Y2=-0.245
cc_118 N_A1_c_133_n N_A2_c_249_n 0.0109765f $X=2.525 $Y=1.935 $X2=-0.19
+ $Y2=-0.245
cc_119 N_A1_M1025_g N_A2_c_243_n 0.0293754f $X=1.425 $Y=0.74 $X2=0 $Y2=0
cc_120 N_A1_c_133_n N_A2_c_250_n 0.00831895f $X=2.525 $Y=1.935 $X2=0 $Y2=0
cc_121 N_A1_c_134_n N_A2_c_251_n 0.0165263f $X=3.235 $Y=1.935 $X2=0 $Y2=0
cc_122 N_A1_c_120_n N_A2_c_252_n 0.0398433f $X=3.76 $Y=1.765 $X2=0 $Y2=0
cc_123 N_A1_c_130_n N_A2_c_252_n 0.00664095f $X=3.64 $Y=1.805 $X2=0 $Y2=0
cc_124 N_A1_c_134_n N_A2_c_252_n 0.00955036f $X=3.235 $Y=1.935 $X2=0 $Y2=0
cc_125 N_A1_M1029_g N_A2_c_246_n 0.0274388f $X=3.855 $Y=0.74 $X2=0 $Y2=0
cc_126 N_A1_M1025_g A2 7.61463e-19 $X=1.425 $Y=0.74 $X2=0 $Y2=0
cc_127 N_A1_M1029_g A2 5.59403e-19 $X=3.855 $Y=0.74 $X2=0 $Y2=0
cc_128 N_A1_c_122_n A2 0.0101061f $X=1.38 $Y=1.485 $X2=0 $Y2=0
cc_129 N_A1_c_123_n A2 0.00788709f $X=3.805 $Y=1.515 $X2=0 $Y2=0
cc_130 N_A1_c_124_n A2 9.98877e-19 $X=1.425 $Y=1.542 $X2=0 $Y2=0
cc_131 N_A1_c_133_n A2 0.10443f $X=2.525 $Y=1.935 $X2=0 $Y2=0
cc_132 N_A1_c_120_n N_A2_c_248_n 0.021845f $X=3.76 $Y=1.765 $X2=0 $Y2=0
cc_133 N_A1_c_122_n N_A2_c_248_n 0.00222133f $X=1.38 $Y=1.485 $X2=0 $Y2=0
cc_134 N_A1_c_130_n N_A2_c_248_n 0.00868406f $X=3.64 $Y=1.805 $X2=0 $Y2=0
cc_135 N_A1_c_123_n N_A2_c_248_n 0.00255637f $X=3.805 $Y=1.515 $X2=0 $Y2=0
cc_136 N_A1_c_124_n N_A2_c_248_n 0.0210999f $X=1.425 $Y=1.542 $X2=0 $Y2=0
cc_137 N_A1_c_133_n N_A2_c_248_n 0.0147227f $X=2.525 $Y=1.935 $X2=0 $Y2=0
cc_138 N_A1_c_134_n N_A2_c_248_n 0.0102026f $X=3.235 $Y=1.935 $X2=0 $Y2=0
cc_139 N_A1_M1029_g N_B1_M1003_g 0.0199157f $X=3.855 $Y=0.74 $X2=0 $Y2=0
cc_140 N_A1_c_120_n N_B1_c_341_n 0.0313624f $X=3.76 $Y=1.765 $X2=0 $Y2=0
cc_141 N_A1_c_123_n N_B1_c_341_n 4.93923e-19 $X=3.805 $Y=1.515 $X2=0 $Y2=0
cc_142 N_A1_c_120_n N_B1_c_336_n 3.18267e-19 $X=3.76 $Y=1.765 $X2=0 $Y2=0
cc_143 N_A1_M1029_g N_B1_c_336_n 2.59363e-19 $X=3.855 $Y=0.74 $X2=0 $Y2=0
cc_144 N_A1_c_123_n N_B1_c_336_n 0.0134326f $X=3.805 $Y=1.515 $X2=0 $Y2=0
cc_145 N_A1_c_120_n N_B1_c_339_n 0.0204385f $X=3.76 $Y=1.765 $X2=0 $Y2=0
cc_146 N_A1_c_123_n N_B1_c_339_n 0.00206488f $X=3.805 $Y=1.515 $X2=0 $Y2=0
cc_147 N_A1_c_125_n N_VPWR_c_541_n 0.008783f $X=0.51 $Y=1.765 $X2=0 $Y2=0
cc_148 N_A1_c_125_n N_VPWR_c_542_n 5.0805e-19 $X=0.51 $Y=1.765 $X2=0 $Y2=0
cc_149 N_A1_c_126_n N_VPWR_c_542_n 0.00957326f $X=0.96 $Y=1.765 $X2=0 $Y2=0
cc_150 N_A1_c_127_n N_VPWR_c_542_n 0.00628391f $X=1.46 $Y=1.765 $X2=0 $Y2=0
cc_151 N_A1_c_120_n N_VPWR_c_543_n 0.00519161f $X=3.76 $Y=1.765 $X2=0 $Y2=0
cc_152 N_A1_c_125_n N_VPWR_c_547_n 0.00445602f $X=0.51 $Y=1.765 $X2=0 $Y2=0
cc_153 N_A1_c_126_n N_VPWR_c_547_n 0.00413917f $X=0.96 $Y=1.765 $X2=0 $Y2=0
cc_154 N_A1_c_127_n N_VPWR_c_548_n 0.00444469f $X=1.46 $Y=1.765 $X2=0 $Y2=0
cc_155 N_A1_c_120_n N_VPWR_c_548_n 0.00444483f $X=3.76 $Y=1.765 $X2=0 $Y2=0
cc_156 N_A1_c_125_n N_VPWR_c_539_n 0.008611f $X=0.51 $Y=1.765 $X2=0 $Y2=0
cc_157 N_A1_c_126_n N_VPWR_c_539_n 0.00817726f $X=0.96 $Y=1.765 $X2=0 $Y2=0
cc_158 N_A1_c_127_n N_VPWR_c_539_n 0.00853793f $X=1.46 $Y=1.765 $X2=0 $Y2=0
cc_159 N_A1_c_120_n N_VPWR_c_539_n 0.00453994f $X=3.76 $Y=1.765 $X2=0 $Y2=0
cc_160 N_A1_c_133_n N_A_117_368#_M1007_s 0.00197722f $X=2.525 $Y=1.935 $X2=0
+ $Y2=0
cc_161 N_A1_c_134_n N_A_117_368#_M1009_d 0.00229049f $X=3.235 $Y=1.935 $X2=0
+ $Y2=0
cc_162 N_A1_c_130_n N_A_117_368#_M1014_d 0.0031003f $X=3.64 $Y=1.805 $X2=0 $Y2=0
cc_163 N_A1_c_125_n N_A_117_368#_c_636_n 0.00863998f $X=0.51 $Y=1.765 $X2=0
+ $Y2=0
cc_164 N_A1_c_126_n N_A_117_368#_c_636_n 2.71519e-19 $X=0.96 $Y=1.765 $X2=0
+ $Y2=0
cc_165 N_A1_c_126_n N_A_117_368#_c_645_n 0.0140516f $X=0.96 $Y=1.765 $X2=0 $Y2=0
cc_166 N_A1_c_127_n N_A_117_368#_c_645_n 0.0122751f $X=1.46 $Y=1.765 $X2=0 $Y2=0
cc_167 N_A1_c_122_n N_A_117_368#_c_645_n 0.0256838f $X=1.38 $Y=1.485 $X2=0 $Y2=0
cc_168 N_A1_c_124_n N_A_117_368#_c_645_n 0.00642683f $X=1.425 $Y=1.542 $X2=0
+ $Y2=0
cc_169 N_A1_c_127_n N_A_117_368#_c_649_n 4.2644e-19 $X=1.46 $Y=1.765 $X2=0 $Y2=0
cc_170 N_A1_c_122_n N_A_117_368#_c_649_n 0.00121062f $X=1.38 $Y=1.485 $X2=0
+ $Y2=0
cc_171 N_A1_c_133_n N_A_117_368#_c_649_n 0.0162332f $X=2.525 $Y=1.935 $X2=0
+ $Y2=0
cc_172 N_A1_c_126_n N_A_117_368#_c_652_n 2.69714e-19 $X=0.96 $Y=1.765 $X2=0
+ $Y2=0
cc_173 N_A1_c_127_n N_A_117_368#_c_652_n 0.00821933f $X=1.46 $Y=1.765 $X2=0
+ $Y2=0
cc_174 N_A1_c_127_n N_A_117_368#_c_637_n 0.00344897f $X=1.46 $Y=1.765 $X2=0
+ $Y2=0
cc_175 N_A1_c_120_n N_A_117_368#_c_638_n 0.0036373f $X=3.76 $Y=1.765 $X2=0 $Y2=0
cc_176 N_A1_c_125_n N_A_117_368#_c_639_n 0.00516862f $X=0.51 $Y=1.765 $X2=0
+ $Y2=0
cc_177 N_A1_c_126_n N_A_117_368#_c_639_n 0.00639387f $X=0.96 $Y=1.765 $X2=0
+ $Y2=0
cc_178 N_A1_c_127_n N_A_117_368#_c_639_n 9.43425e-19 $X=1.46 $Y=1.765 $X2=0
+ $Y2=0
cc_179 N_A1_c_122_n N_A_117_368#_c_639_n 0.0288487f $X=1.38 $Y=1.485 $X2=0 $Y2=0
cc_180 N_A1_c_124_n N_A_117_368#_c_639_n 0.0076085f $X=1.425 $Y=1.542 $X2=0
+ $Y2=0
cc_181 N_A1_c_133_n N_Y_M1008_s 0.00250873f $X=2.525 $Y=1.935 $X2=0 $Y2=0
cc_182 N_A1_c_134_n N_Y_M1010_s 0.00229049f $X=3.235 $Y=1.935 $X2=0 $Y2=0
cc_183 N_A1_c_120_n N_Y_c_695_n 0.0139858f $X=3.76 $Y=1.765 $X2=0 $Y2=0
cc_184 N_A1_c_130_n N_Y_c_695_n 0.011587f $X=3.64 $Y=1.805 $X2=0 $Y2=0
cc_185 N_A1_c_123_n N_Y_c_695_n 0.00772626f $X=3.805 $Y=1.515 $X2=0 $Y2=0
cc_186 N_A1_c_133_n N_Y_c_695_n 0.00432188f $X=2.525 $Y=1.935 $X2=0 $Y2=0
cc_187 N_A1_c_134_n N_Y_c_695_n 0.0399401f $X=3.235 $Y=1.935 $X2=0 $Y2=0
cc_188 N_A1_c_120_n N_Y_c_700_n 0.00674458f $X=3.76 $Y=1.765 $X2=0 $Y2=0
cc_189 N_A1_c_120_n N_Y_c_701_n 0.00417391f $X=3.76 $Y=1.765 $X2=0 $Y2=0
cc_190 N_A1_c_123_n N_Y_c_701_n 0.00349616f $X=3.805 $Y=1.515 $X2=0 $Y2=0
cc_191 N_A1_c_133_n N_Y_c_703_n 0.0195313f $X=2.525 $Y=1.935 $X2=0 $Y2=0
cc_192 N_A1_c_120_n N_A_877_368#_c_832_n 9.30091e-19 $X=3.76 $Y=1.765 $X2=0
+ $Y2=0
cc_193 N_A1_M1000_g N_A_27_74#_c_883_n 0.00980115f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_194 N_A1_M1011_g N_A_27_74#_c_883_n 9.32548e-19 $X=0.995 $Y=0.74 $X2=0 $Y2=0
cc_195 N_A1_M1000_g N_A_27_74#_c_884_n 0.0143535f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_196 N_A1_M1011_g N_A_27_74#_c_884_n 0.01285f $X=0.995 $Y=0.74 $X2=0 $Y2=0
cc_197 N_A1_c_122_n N_A_27_74#_c_884_n 0.0432965f $X=1.38 $Y=1.485 $X2=0 $Y2=0
cc_198 N_A1_c_124_n N_A_27_74#_c_884_n 0.00381149f $X=1.425 $Y=1.542 $X2=0 $Y2=0
cc_199 N_A1_M1000_g N_A_27_74#_c_885_n 0.00243964f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_200 N_A1_M1011_g N_A_27_74#_c_886_n 3.97481e-19 $X=0.995 $Y=0.74 $X2=0 $Y2=0
cc_201 N_A1_M1025_g N_A_27_74#_c_886_n 0.00739853f $X=1.425 $Y=0.74 $X2=0 $Y2=0
cc_202 N_A1_M1025_g N_A_27_74#_c_907_n 0.0104473f $X=1.425 $Y=0.74 $X2=0 $Y2=0
cc_203 N_A1_c_122_n N_A_27_74#_c_907_n 0.0069724f $X=1.38 $Y=1.485 $X2=0 $Y2=0
cc_204 N_A1_c_120_n N_A_27_74#_c_889_n 9.8174e-19 $X=3.76 $Y=1.765 $X2=0 $Y2=0
cc_205 N_A1_M1029_g N_A_27_74#_c_889_n 0.0131779f $X=3.855 $Y=0.74 $X2=0 $Y2=0
cc_206 N_A1_c_123_n N_A_27_74#_c_889_n 0.0146621f $X=3.805 $Y=1.515 $X2=0 $Y2=0
cc_207 N_A1_M1029_g N_A_27_74#_c_890_n 0.00485335f $X=3.855 $Y=0.74 $X2=0 $Y2=0
cc_208 N_A1_M1029_g N_A_27_74#_c_913_n 0.00504463f $X=3.855 $Y=0.74 $X2=0 $Y2=0
cc_209 N_A1_M1025_g N_A_27_74#_c_892_n 0.00416046f $X=1.425 $Y=0.74 $X2=0 $Y2=0
cc_210 N_A1_c_122_n N_A_27_74#_c_892_n 0.0208089f $X=1.38 $Y=1.485 $X2=0 $Y2=0
cc_211 N_A1_c_124_n N_A_27_74#_c_892_n 0.00232957f $X=1.425 $Y=1.542 $X2=0 $Y2=0
cc_212 N_A1_M1000_g N_VGND_c_1009_n 0.00555396f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_213 N_A1_M1011_g N_VGND_c_1009_n 0.0098353f $X=0.995 $Y=0.74 $X2=0 $Y2=0
cc_214 N_A1_M1025_g N_VGND_c_1009_n 5.08869e-19 $X=1.425 $Y=0.74 $X2=0 $Y2=0
cc_215 N_A1_M1025_g N_VGND_c_1010_n 0.00335277f $X=1.425 $Y=0.74 $X2=0 $Y2=0
cc_216 N_A1_M1029_g N_VGND_c_1012_n 0.00309798f $X=3.855 $Y=0.74 $X2=0 $Y2=0
cc_217 N_A1_M1000_g N_VGND_c_1013_n 0.00434272f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_218 N_A1_M1011_g N_VGND_c_1014_n 0.00383152f $X=0.995 $Y=0.74 $X2=0 $Y2=0
cc_219 N_A1_M1025_g N_VGND_c_1014_n 0.00434272f $X=1.425 $Y=0.74 $X2=0 $Y2=0
cc_220 N_A1_M1029_g N_VGND_c_1017_n 0.00430908f $X=3.855 $Y=0.74 $X2=0 $Y2=0
cc_221 N_A1_M1000_g N_VGND_c_1018_n 0.00824376f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_222 N_A1_M1011_g N_VGND_c_1018_n 0.0075754f $X=0.995 $Y=0.74 $X2=0 $Y2=0
cc_223 N_A1_M1025_g N_VGND_c_1018_n 0.00445549f $X=1.425 $Y=0.74 $X2=0 $Y2=0
cc_224 N_A1_M1029_g N_VGND_c_1018_n 0.00445992f $X=3.855 $Y=0.74 $X2=0 $Y2=0
cc_225 N_A2_c_249_n N_VPWR_c_548_n 0.00291635f $X=1.91 $Y=1.765 $X2=0 $Y2=0
cc_226 N_A2_c_250_n N_VPWR_c_548_n 0.00291649f $X=2.41 $Y=1.765 $X2=0 $Y2=0
cc_227 N_A2_c_251_n N_VPWR_c_548_n 0.00291649f $X=2.86 $Y=1.765 $X2=0 $Y2=0
cc_228 N_A2_c_252_n N_VPWR_c_548_n 0.00291649f $X=3.31 $Y=1.765 $X2=0 $Y2=0
cc_229 N_A2_c_249_n N_VPWR_c_539_n 0.0036005f $X=1.91 $Y=1.765 $X2=0 $Y2=0
cc_230 N_A2_c_250_n N_VPWR_c_539_n 0.00359029f $X=2.41 $Y=1.765 $X2=0 $Y2=0
cc_231 N_A2_c_251_n N_VPWR_c_539_n 0.00359515f $X=2.86 $Y=1.765 $X2=0 $Y2=0
cc_232 N_A2_c_252_n N_VPWR_c_539_n 0.00359599f $X=3.31 $Y=1.765 $X2=0 $Y2=0
cc_233 N_A2_c_249_n N_A_117_368#_c_649_n 0.00183099f $X=1.91 $Y=1.765 $X2=0
+ $Y2=0
cc_234 N_A2_c_249_n N_A_117_368#_c_652_n 0.0080872f $X=1.91 $Y=1.765 $X2=0 $Y2=0
cc_235 N_A2_c_250_n N_A_117_368#_c_652_n 8.55793e-19 $X=2.41 $Y=1.765 $X2=0
+ $Y2=0
cc_236 N_A2_c_249_n N_A_117_368#_c_637_n 8.06278e-19 $X=1.91 $Y=1.765 $X2=0
+ $Y2=0
cc_237 N_A2_c_249_n N_A_117_368#_c_638_n 0.0162584f $X=1.91 $Y=1.765 $X2=0 $Y2=0
cc_238 N_A2_c_250_n N_A_117_368#_c_638_n 0.0128011f $X=2.41 $Y=1.765 $X2=0 $Y2=0
cc_239 N_A2_c_251_n N_A_117_368#_c_638_n 0.0122986f $X=2.86 $Y=1.765 $X2=0 $Y2=0
cc_240 N_A2_c_252_n N_A_117_368#_c_638_n 0.0122931f $X=3.31 $Y=1.765 $X2=0 $Y2=0
cc_241 N_A2_c_250_n N_Y_c_695_n 0.00968513f $X=2.41 $Y=1.765 $X2=0 $Y2=0
cc_242 N_A2_c_251_n N_Y_c_695_n 0.00855704f $X=2.86 $Y=1.765 $X2=0 $Y2=0
cc_243 N_A2_c_252_n N_Y_c_695_n 0.00986206f $X=3.31 $Y=1.765 $X2=0 $Y2=0
cc_244 N_A2_c_250_n N_Y_c_703_n 0.00551791f $X=2.41 $Y=1.765 $X2=0 $Y2=0
cc_245 N_A2_c_251_n N_Y_c_703_n 9.55407e-19 $X=2.86 $Y=1.765 $X2=0 $Y2=0
cc_246 N_A2_c_243_n N_A_27_74#_c_886_n 7.18081e-19 $X=1.925 $Y=1.22 $X2=0 $Y2=0
cc_247 N_A2_c_243_n N_A_27_74#_c_907_n 0.0110188f $X=1.925 $Y=1.22 $X2=0 $Y2=0
cc_248 A2 N_A_27_74#_c_907_n 0.0105847f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_249 N_A2_c_243_n N_A_27_74#_c_887_n 2.29136e-19 $X=1.925 $Y=1.22 $X2=0 $Y2=0
cc_250 N_A2_c_244_n N_A_27_74#_c_887_n 0.00703259f $X=2.355 $Y=1.22 $X2=0 $Y2=0
cc_251 N_A2_c_245_n N_A_27_74#_c_887_n 7.13338e-19 $X=2.855 $Y=1.22 $X2=0 $Y2=0
cc_252 N_A2_c_244_n N_A_27_74#_c_923_n 0.00892313f $X=2.355 $Y=1.22 $X2=0 $Y2=0
cc_253 N_A2_c_245_n N_A_27_74#_c_923_n 0.0100105f $X=2.855 $Y=1.22 $X2=0 $Y2=0
cc_254 A2 N_A_27_74#_c_923_n 0.0454799f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_255 N_A2_c_248_n N_A_27_74#_c_923_n 0.00106692f $X=3.31 $Y=1.492 $X2=0 $Y2=0
cc_256 N_A2_c_245_n N_A_27_74#_c_888_n 2.49954e-19 $X=2.855 $Y=1.22 $X2=0 $Y2=0
cc_257 N_A2_c_246_n N_A_27_74#_c_888_n 2.68395e-19 $X=3.325 $Y=1.22 $X2=0 $Y2=0
cc_258 N_A2_c_246_n N_A_27_74#_c_889_n 0.0154305f $X=3.325 $Y=1.22 $X2=0 $Y2=0
cc_259 N_A2_c_246_n N_A_27_74#_c_913_n 3.72705e-19 $X=3.325 $Y=1.22 $X2=0 $Y2=0
cc_260 N_A2_c_243_n N_A_27_74#_c_892_n 7.4692e-19 $X=1.925 $Y=1.22 $X2=0 $Y2=0
cc_261 N_A2_c_244_n N_A_27_74#_c_932_n 7.17169e-19 $X=2.355 $Y=1.22 $X2=0 $Y2=0
cc_262 A2 N_A_27_74#_c_932_n 0.0189543f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_263 N_A2_c_248_n N_A_27_74#_c_932_n 7.06072e-19 $X=3.31 $Y=1.492 $X2=0 $Y2=0
cc_264 A2 N_A_27_74#_c_935_n 0.0198393f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_265 N_A2_c_248_n N_A_27_74#_c_935_n 9.84341e-19 $X=3.31 $Y=1.492 $X2=0 $Y2=0
cc_266 N_A2_c_243_n N_VGND_c_1010_n 0.00771106f $X=1.925 $Y=1.22 $X2=0 $Y2=0
cc_267 N_A2_c_244_n N_VGND_c_1010_n 4.39845e-19 $X=2.355 $Y=1.22 $X2=0 $Y2=0
cc_268 N_A2_c_244_n N_VGND_c_1011_n 0.00335277f $X=2.355 $Y=1.22 $X2=0 $Y2=0
cc_269 N_A2_c_245_n N_VGND_c_1011_n 0.00775702f $X=2.855 $Y=1.22 $X2=0 $Y2=0
cc_270 N_A2_c_246_n N_VGND_c_1011_n 4.2363e-19 $X=3.325 $Y=1.22 $X2=0 $Y2=0
cc_271 N_A2_c_246_n N_VGND_c_1012_n 0.00199261f $X=3.325 $Y=1.22 $X2=0 $Y2=0
cc_272 N_A2_c_243_n N_VGND_c_1015_n 0.00383152f $X=1.925 $Y=1.22 $X2=0 $Y2=0
cc_273 N_A2_c_244_n N_VGND_c_1015_n 0.00434272f $X=2.355 $Y=1.22 $X2=0 $Y2=0
cc_274 N_A2_c_245_n N_VGND_c_1016_n 0.00383152f $X=2.855 $Y=1.22 $X2=0 $Y2=0
cc_275 N_A2_c_246_n N_VGND_c_1016_n 0.00461464f $X=3.325 $Y=1.22 $X2=0 $Y2=0
cc_276 N_A2_c_243_n N_VGND_c_1018_n 0.00383967f $X=1.925 $Y=1.22 $X2=0 $Y2=0
cc_277 N_A2_c_244_n N_VGND_c_1018_n 0.00445496f $X=2.355 $Y=1.22 $X2=0 $Y2=0
cc_278 N_A2_c_245_n N_VGND_c_1018_n 0.00384354f $X=2.855 $Y=1.22 $X2=0 $Y2=0
cc_279 N_A2_c_246_n N_VGND_c_1018_n 0.00463822f $X=3.325 $Y=1.22 $X2=0 $Y2=0
cc_280 N_B1_M1023_g N_B2_M1013_g 0.0236891f $X=5.225 $Y=0.74 $X2=0 $Y2=0
cc_281 N_B1_c_336_n N_B2_M1013_g 3.11251e-19 $X=5.405 $Y=1.465 $X2=0 $Y2=0
cc_282 N_B1_c_337_n N_B2_M1013_g 0.00788083f $X=7.4 $Y=1.175 $X2=0 $Y2=0
cc_283 N_B1_c_340_n N_B2_M1013_g 0.00599736f $X=5.52 $Y=1.175 $X2=0 $Y2=0
cc_284 N_B1_c_343_n N_B2_c_457_n 0.0299545f $X=5.21 $Y=1.765 $X2=0 $Y2=0
cc_285 N_B1_c_337_n N_B2_M1019_g 0.0108858f $X=7.4 $Y=1.175 $X2=0 $Y2=0
cc_286 N_B1_c_340_n N_B2_M1019_g 5.5004e-19 $X=5.52 $Y=1.175 $X2=0 $Y2=0
cc_287 N_B1_c_337_n N_B2_M1021_g 0.0112791f $X=7.4 $Y=1.175 $X2=0 $Y2=0
cc_288 N_B1_c_334_n N_B2_c_460_n 0.0235108f $X=7.56 $Y=1.765 $X2=0 $Y2=0
cc_289 N_B1_c_334_n N_B2_M1026_g 0.0187736f $X=7.56 $Y=1.765 $X2=0 $Y2=0
cc_290 N_B1_c_335_n N_B2_M1026_g 0.0270173f $X=7.585 $Y=1.22 $X2=0 $Y2=0
cc_291 N_B1_c_337_n N_B2_M1026_g 0.0108221f $X=7.4 $Y=1.175 $X2=0 $Y2=0
cc_292 N_B1_c_338_n N_B2_M1026_g 0.00185513f $X=7.565 $Y=1.175 $X2=0 $Y2=0
cc_293 N_B1_c_334_n N_B2_c_461_n 0.00207557f $X=7.56 $Y=1.765 $X2=0 $Y2=0
cc_294 N_B1_c_338_n N_B2_c_461_n 0.0070832f $X=7.565 $Y=1.175 $X2=0 $Y2=0
cc_295 N_B1_c_334_n N_B2_c_456_n 0.00955853f $X=7.56 $Y=1.765 $X2=0 $Y2=0
cc_296 N_B1_c_337_n N_B2_c_456_n 0.0108448f $X=7.4 $Y=1.175 $X2=0 $Y2=0
cc_297 N_B1_c_339_n N_B2_c_456_n 0.0276235f $X=5.21 $Y=1.532 $X2=0 $Y2=0
cc_298 N_B1_c_340_n N_B2_c_456_n 0.0105603f $X=5.52 $Y=1.175 $X2=0 $Y2=0
cc_299 N_B1_c_337_n N_B2_c_483_n 0.0991186f $X=7.4 $Y=1.175 $X2=0 $Y2=0
cc_300 N_B1_c_339_n N_B2_c_483_n 2.04599e-19 $X=5.21 $Y=1.532 $X2=0 $Y2=0
cc_301 N_B1_c_340_n N_B2_c_483_n 0.0154812f $X=5.52 $Y=1.175 $X2=0 $Y2=0
cc_302 N_B1_c_341_n N_VPWR_c_543_n 0.00517191f $X=4.31 $Y=1.765 $X2=0 $Y2=0
cc_303 N_B1_c_342_n N_VPWR_c_544_n 0.00460996f $X=4.76 $Y=1.765 $X2=0 $Y2=0
cc_304 N_B1_c_343_n N_VPWR_c_544_n 0.0076142f $X=5.21 $Y=1.765 $X2=0 $Y2=0
cc_305 N_B1_c_334_n N_VPWR_c_546_n 0.0163641f $X=7.56 $Y=1.765 $X2=0 $Y2=0
cc_306 N_B1_c_341_n N_VPWR_c_549_n 0.00445602f $X=4.31 $Y=1.765 $X2=0 $Y2=0
cc_307 N_B1_c_342_n N_VPWR_c_549_n 0.00445602f $X=4.76 $Y=1.765 $X2=0 $Y2=0
cc_308 N_B1_c_343_n N_VPWR_c_550_n 0.00413917f $X=5.21 $Y=1.765 $X2=0 $Y2=0
cc_309 N_B1_c_334_n N_VPWR_c_550_n 0.0044313f $X=7.56 $Y=1.765 $X2=0 $Y2=0
cc_310 N_B1_c_341_n N_VPWR_c_539_n 0.00857825f $X=4.31 $Y=1.765 $X2=0 $Y2=0
cc_311 N_B1_c_342_n N_VPWR_c_539_n 0.00857589f $X=4.76 $Y=1.765 $X2=0 $Y2=0
cc_312 N_B1_c_343_n N_VPWR_c_539_n 0.00818241f $X=5.21 $Y=1.765 $X2=0 $Y2=0
cc_313 N_B1_c_334_n N_VPWR_c_539_n 0.00856889f $X=7.56 $Y=1.765 $X2=0 $Y2=0
cc_314 N_B1_c_340_n N_Y_M1023_s 0.00148168f $X=5.52 $Y=1.175 $X2=0 $Y2=0
cc_315 N_B1_c_337_n N_Y_M1019_s 0.00251484f $X=7.4 $Y=1.175 $X2=0 $Y2=0
cc_316 N_B1_c_337_n N_Y_M1026_s 0.00199526f $X=7.4 $Y=1.175 $X2=0 $Y2=0
cc_317 N_B1_c_338_n N_Y_M1026_s 6.17026e-19 $X=7.565 $Y=1.175 $X2=0 $Y2=0
cc_318 N_B1_c_341_n N_Y_c_695_n 0.0016959f $X=4.31 $Y=1.765 $X2=0 $Y2=0
cc_319 N_B1_c_341_n N_Y_c_700_n 0.00525286f $X=4.31 $Y=1.765 $X2=0 $Y2=0
cc_320 N_B1_c_341_n N_Y_c_715_n 0.0166356f $X=4.31 $Y=1.765 $X2=0 $Y2=0
cc_321 N_B1_c_342_n N_Y_c_715_n 0.0109799f $X=4.76 $Y=1.765 $X2=0 $Y2=0
cc_322 N_B1_c_343_n N_Y_c_715_n 0.0112441f $X=5.21 $Y=1.765 $X2=0 $Y2=0
cc_323 N_B1_c_336_n N_Y_c_715_n 0.0584372f $X=5.405 $Y=1.465 $X2=0 $Y2=0
cc_324 N_B1_c_337_n N_Y_c_715_n 0.00341175f $X=7.4 $Y=1.175 $X2=0 $Y2=0
cc_325 N_B1_c_339_n N_Y_c_715_n 0.0122957f $X=5.21 $Y=1.532 $X2=0 $Y2=0
cc_326 N_B1_c_340_n N_Y_c_715_n 0.0135056f $X=5.52 $Y=1.175 $X2=0 $Y2=0
cc_327 N_B1_c_334_n N_Y_c_691_n 0.0184267f $X=7.56 $Y=1.765 $X2=0 $Y2=0
cc_328 N_B1_c_338_n N_Y_c_691_n 0.0103133f $X=7.565 $Y=1.175 $X2=0 $Y2=0
cc_329 N_B1_c_334_n N_Y_c_687_n 2.54483e-19 $X=7.56 $Y=1.765 $X2=0 $Y2=0
cc_330 N_B1_c_335_n N_Y_c_687_n 0.00967079f $X=7.585 $Y=1.22 $X2=0 $Y2=0
cc_331 N_B1_c_334_n N_Y_c_688_n 0.0199854f $X=7.56 $Y=1.765 $X2=0 $Y2=0
cc_332 N_B1_c_335_n N_Y_c_688_n 0.00614976f $X=7.585 $Y=1.22 $X2=0 $Y2=0
cc_333 N_B1_c_338_n N_Y_c_688_n 0.0350504f $X=7.565 $Y=1.175 $X2=0 $Y2=0
cc_334 N_B1_c_343_n N_Y_c_729_n 0.0010098f $X=5.21 $Y=1.765 $X2=0 $Y2=0
cc_335 N_B1_c_337_n N_Y_c_729_n 7.66151e-19 $X=7.4 $Y=1.175 $X2=0 $Y2=0
cc_336 N_B1_M1023_g N_Y_c_731_n 0.00725011f $X=5.225 $Y=0.74 $X2=0 $Y2=0
cc_337 N_B1_c_336_n N_Y_c_731_n 0.00885985f $X=5.405 $Y=1.465 $X2=0 $Y2=0
cc_338 N_B1_c_337_n N_Y_c_731_n 0.09861f $X=7.4 $Y=1.175 $X2=0 $Y2=0
cc_339 N_B1_c_340_n N_Y_c_731_n 0.0133434f $X=5.52 $Y=1.175 $X2=0 $Y2=0
cc_340 N_B1_c_334_n N_Y_c_735_n 7.09751e-19 $X=7.56 $Y=1.765 $X2=0 $Y2=0
cc_341 N_B1_c_334_n N_Y_c_736_n 4.70019e-19 $X=7.56 $Y=1.765 $X2=0 $Y2=0
cc_342 N_B1_c_335_n N_Y_c_736_n 0.00788319f $X=7.585 $Y=1.22 $X2=0 $Y2=0
cc_343 N_B1_c_338_n N_Y_c_736_n 0.0163546f $X=7.565 $Y=1.175 $X2=0 $Y2=0
cc_344 N_B1_M1003_g N_Y_c_689_n 0.00203855f $X=4.295 $Y=0.74 $X2=0 $Y2=0
cc_345 N_B1_M1016_g N_Y_c_689_n 0.0143968f $X=4.785 $Y=0.74 $X2=0 $Y2=0
cc_346 N_B1_c_336_n N_Y_c_689_n 0.0593442f $X=5.405 $Y=1.465 $X2=0 $Y2=0
cc_347 N_B1_c_339_n N_Y_c_689_n 0.00617128f $X=5.21 $Y=1.532 $X2=0 $Y2=0
cc_348 N_B1_M1023_g N_Y_c_690_n 0.008409f $X=5.225 $Y=0.74 $X2=0 $Y2=0
cc_349 N_B1_c_340_n N_Y_c_690_n 0.00235206f $X=5.52 $Y=1.175 $X2=0 $Y2=0
cc_350 N_B1_c_342_n N_A_877_368#_c_835_n 0.0120074f $X=4.76 $Y=1.765 $X2=0 $Y2=0
cc_351 N_B1_c_343_n N_A_877_368#_c_835_n 0.0147239f $X=5.21 $Y=1.765 $X2=0 $Y2=0
cc_352 N_B1_c_343_n N_A_877_368#_c_830_n 0.0013657f $X=5.21 $Y=1.765 $X2=0 $Y2=0
cc_353 N_B1_c_334_n N_A_877_368#_c_831_n 0.00333933f $X=7.56 $Y=1.765 $X2=0
+ $Y2=0
cc_354 N_B1_c_334_n N_A_877_368#_c_839_n 0.00630596f $X=7.56 $Y=1.765 $X2=0
+ $Y2=0
cc_355 N_B1_c_341_n N_A_877_368#_c_832_n 0.011029f $X=4.31 $Y=1.765 $X2=0 $Y2=0
cc_356 N_B1_c_342_n N_A_877_368#_c_832_n 0.00935636f $X=4.76 $Y=1.765 $X2=0
+ $Y2=0
cc_357 N_B1_c_343_n N_A_877_368#_c_832_n 6.74271e-19 $X=5.21 $Y=1.765 $X2=0
+ $Y2=0
cc_358 N_B1_c_337_n N_A_27_74#_M1013_d 0.00176891f $X=7.4 $Y=1.175 $X2=0 $Y2=0
cc_359 N_B1_c_337_n N_A_27_74#_M1021_d 0.00251484f $X=7.4 $Y=1.175 $X2=0 $Y2=0
cc_360 N_B1_c_338_n N_A_27_74#_M1028_d 3.49062e-19 $X=7.565 $Y=1.175 $X2=0 $Y2=0
cc_361 N_B1_M1003_g N_A_27_74#_c_889_n 0.00373455f $X=4.295 $Y=0.74 $X2=0 $Y2=0
cc_362 N_B1_M1003_g N_A_27_74#_c_890_n 0.00188298f $X=4.295 $Y=0.74 $X2=0 $Y2=0
cc_363 N_B1_M1003_g N_A_27_74#_c_913_n 0.00469212f $X=4.295 $Y=0.74 $X2=0 $Y2=0
cc_364 N_B1_M1016_g N_A_27_74#_c_913_n 7.81702e-19 $X=4.785 $Y=0.74 $X2=0 $Y2=0
cc_365 N_B1_M1003_g N_A_27_74#_c_891_n 0.0156461f $X=4.295 $Y=0.74 $X2=0 $Y2=0
cc_366 N_B1_M1016_g N_A_27_74#_c_891_n 0.0132936f $X=4.785 $Y=0.74 $X2=0 $Y2=0
cc_367 N_B1_M1023_g N_A_27_74#_c_891_n 0.0125475f $X=5.225 $Y=0.74 $X2=0 $Y2=0
cc_368 N_B1_c_335_n N_A_27_74#_c_895_n 3.47155e-19 $X=7.585 $Y=1.22 $X2=0 $Y2=0
cc_369 N_B1_c_335_n N_A_27_74#_c_897_n 0.0118166f $X=7.585 $Y=1.22 $X2=0 $Y2=0
cc_370 N_B1_M1003_g N_VGND_c_1017_n 0.00278257f $X=4.295 $Y=0.74 $X2=0 $Y2=0
cc_371 N_B1_M1016_g N_VGND_c_1017_n 0.00278271f $X=4.785 $Y=0.74 $X2=0 $Y2=0
cc_372 N_B1_M1023_g N_VGND_c_1017_n 0.00278271f $X=5.225 $Y=0.74 $X2=0 $Y2=0
cc_373 N_B1_c_335_n N_VGND_c_1017_n 0.00278271f $X=7.585 $Y=1.22 $X2=0 $Y2=0
cc_374 N_B1_M1003_g N_VGND_c_1018_n 0.00354187f $X=4.295 $Y=0.74 $X2=0 $Y2=0
cc_375 N_B1_M1016_g N_VGND_c_1018_n 0.00354097f $X=4.785 $Y=0.74 $X2=0 $Y2=0
cc_376 N_B1_M1023_g N_VGND_c_1018_n 0.00353625f $X=5.225 $Y=0.74 $X2=0 $Y2=0
cc_377 N_B1_c_335_n N_VGND_c_1018_n 0.00358041f $X=7.585 $Y=1.22 $X2=0 $Y2=0
cc_378 N_B2_c_457_n N_VPWR_c_550_n 0.00278271f $X=5.71 $Y=1.765 $X2=0 $Y2=0
cc_379 N_B2_c_458_n N_VPWR_c_550_n 0.00278271f $X=6.16 $Y=1.765 $X2=0 $Y2=0
cc_380 N_B2_c_459_n N_VPWR_c_550_n 0.00278271f $X=6.61 $Y=1.765 $X2=0 $Y2=0
cc_381 N_B2_c_460_n N_VPWR_c_550_n 0.00278271f $X=7.07 $Y=1.765 $X2=0 $Y2=0
cc_382 N_B2_c_457_n N_VPWR_c_539_n 0.00354337f $X=5.71 $Y=1.765 $X2=0 $Y2=0
cc_383 N_B2_c_458_n N_VPWR_c_539_n 0.00353823f $X=6.16 $Y=1.765 $X2=0 $Y2=0
cc_384 N_B2_c_459_n N_VPWR_c_539_n 0.00353919f $X=6.61 $Y=1.765 $X2=0 $Y2=0
cc_385 N_B2_c_460_n N_VPWR_c_539_n 0.00350714f $X=7.07 $Y=1.765 $X2=0 $Y2=0
cc_386 N_B2_c_457_n N_Y_c_715_n 0.014011f $X=5.71 $Y=1.765 $X2=0 $Y2=0
cc_387 N_B2_c_458_n N_Y_c_746_n 0.012525f $X=6.16 $Y=1.765 $X2=0 $Y2=0
cc_388 N_B2_c_459_n N_Y_c_746_n 0.0120074f $X=6.61 $Y=1.765 $X2=0 $Y2=0
cc_389 N_B2_c_456_n N_Y_c_746_n 0.00305342f $X=7.07 $Y=1.557 $X2=0 $Y2=0
cc_390 N_B2_c_463_n N_Y_c_746_n 0.0208976f $X=6.715 $Y=1.605 $X2=0 $Y2=0
cc_391 N_B2_c_483_n N_Y_c_746_n 0.0115835f $X=6.365 $Y=1.605 $X2=0 $Y2=0
cc_392 N_B2_c_460_n N_Y_c_691_n 0.0129073f $X=7.07 $Y=1.765 $X2=0 $Y2=0
cc_393 N_B2_c_461_n N_Y_c_691_n 0.0107902f $X=6.99 $Y=1.515 $X2=0 $Y2=0
cc_394 N_B2_c_457_n N_Y_c_729_n 0.0117736f $X=5.71 $Y=1.765 $X2=0 $Y2=0
cc_395 N_B2_c_458_n N_Y_c_729_n 0.0121294f $X=6.16 $Y=1.765 $X2=0 $Y2=0
cc_396 N_B2_c_459_n N_Y_c_729_n 0.00104171f $X=6.61 $Y=1.765 $X2=0 $Y2=0
cc_397 N_B2_c_456_n N_Y_c_729_n 0.00670438f $X=7.07 $Y=1.557 $X2=0 $Y2=0
cc_398 N_B2_c_483_n N_Y_c_729_n 0.0195958f $X=6.365 $Y=1.605 $X2=0 $Y2=0
cc_399 N_B2_M1013_g N_Y_c_731_n 0.00841587f $X=5.655 $Y=0.74 $X2=0 $Y2=0
cc_400 N_B2_M1019_g N_Y_c_731_n 0.0118672f $X=6.085 $Y=0.74 $X2=0 $Y2=0
cc_401 N_B2_M1021_g N_Y_c_760_n 0.00427826f $X=6.585 $Y=0.74 $X2=0 $Y2=0
cc_402 N_B2_M1026_g N_Y_c_760_n 2.63525e-19 $X=7.085 $Y=0.74 $X2=0 $Y2=0
cc_403 N_B2_c_458_n N_Y_c_735_n 5.7112e-19 $X=6.16 $Y=1.765 $X2=0 $Y2=0
cc_404 N_B2_c_459_n N_Y_c_735_n 0.00894037f $X=6.61 $Y=1.765 $X2=0 $Y2=0
cc_405 N_B2_c_460_n N_Y_c_735_n 0.00776489f $X=7.07 $Y=1.765 $X2=0 $Y2=0
cc_406 N_B2_c_456_n N_Y_c_735_n 0.00152565f $X=7.07 $Y=1.557 $X2=0 $Y2=0
cc_407 N_B2_c_463_n N_Y_c_735_n 0.0233502f $X=6.715 $Y=1.605 $X2=0 $Y2=0
cc_408 N_B2_M1021_g N_Y_c_767_n 0.00757292f $X=6.585 $Y=0.74 $X2=0 $Y2=0
cc_409 N_B2_M1026_g N_Y_c_767_n 0.0121078f $X=7.085 $Y=0.74 $X2=0 $Y2=0
cc_410 N_B2_M1013_g N_Y_c_690_n 5.9325e-19 $X=5.655 $Y=0.74 $X2=0 $Y2=0
cc_411 N_B2_c_457_n N_A_877_368#_c_843_n 0.0052306f $X=5.71 $Y=1.765 $X2=0 $Y2=0
cc_412 N_B2_c_457_n N_A_877_368#_c_829_n 0.0127803f $X=5.71 $Y=1.765 $X2=0 $Y2=0
cc_413 N_B2_c_458_n N_A_877_368#_c_829_n 0.0128349f $X=6.16 $Y=1.765 $X2=0 $Y2=0
cc_414 N_B2_c_459_n N_A_877_368#_c_831_n 0.0128926f $X=6.61 $Y=1.765 $X2=0 $Y2=0
cc_415 N_B2_c_460_n N_A_877_368#_c_831_n 0.0132531f $X=7.07 $Y=1.765 $X2=0 $Y2=0
cc_416 N_B2_M1013_g N_A_27_74#_c_891_n 0.0124925f $X=5.655 $Y=0.74 $X2=0 $Y2=0
cc_417 N_B2_M1019_g N_A_27_74#_c_893_n 0.00528709f $X=6.085 $Y=0.74 $X2=0 $Y2=0
cc_418 N_B2_M1021_g N_A_27_74#_c_893_n 3.43302e-19 $X=6.585 $Y=0.74 $X2=0 $Y2=0
cc_419 N_B2_M1019_g N_A_27_74#_c_894_n 0.00644043f $X=6.085 $Y=0.74 $X2=0 $Y2=0
cc_420 N_B2_M1021_g N_A_27_74#_c_894_n 0.0110646f $X=6.585 $Y=0.74 $X2=0 $Y2=0
cc_421 N_B2_M1026_g N_A_27_74#_c_895_n 0.00557328f $X=7.085 $Y=0.74 $X2=0 $Y2=0
cc_422 N_B2_M1026_g N_A_27_74#_c_897_n 0.00642625f $X=7.085 $Y=0.74 $X2=0 $Y2=0
cc_423 N_B2_M1013_g N_VGND_c_1017_n 0.00278271f $X=5.655 $Y=0.74 $X2=0 $Y2=0
cc_424 N_B2_M1019_g N_VGND_c_1017_n 0.00278271f $X=6.085 $Y=0.74 $X2=0 $Y2=0
cc_425 N_B2_M1021_g N_VGND_c_1017_n 0.00278271f $X=6.585 $Y=0.74 $X2=0 $Y2=0
cc_426 N_B2_M1026_g N_VGND_c_1017_n 0.00278271f $X=7.085 $Y=0.74 $X2=0 $Y2=0
cc_427 N_B2_M1013_g N_VGND_c_1018_n 0.00353526f $X=5.655 $Y=0.74 $X2=0 $Y2=0
cc_428 N_B2_M1019_g N_VGND_c_1018_n 0.00354087f $X=6.085 $Y=0.74 $X2=0 $Y2=0
cc_429 N_B2_M1021_g N_VGND_c_1018_n 0.00354745f $X=6.585 $Y=0.74 $X2=0 $Y2=0
cc_430 N_B2_M1026_g N_VGND_c_1018_n 0.00354798f $X=7.085 $Y=0.74 $X2=0 $Y2=0
cc_431 N_VPWR_c_542_n N_A_117_368#_c_636_n 0.022534f $X=1.185 $Y=2.485 $X2=0
+ $Y2=0
cc_432 N_VPWR_c_547_n N_A_117_368#_c_636_n 0.0123628f $X=1.02 $Y=3.33 $X2=0
+ $Y2=0
cc_433 N_VPWR_c_539_n N_A_117_368#_c_636_n 0.0101999f $X=7.92 $Y=3.33 $X2=0
+ $Y2=0
cc_434 N_VPWR_M1006_d N_A_117_368#_c_645_n 0.00567466f $X=1.035 $Y=1.84 $X2=0
+ $Y2=0
cc_435 N_VPWR_c_542_n N_A_117_368#_c_645_n 0.0202249f $X=1.185 $Y=2.485 $X2=0
+ $Y2=0
cc_436 N_VPWR_c_542_n N_A_117_368#_c_637_n 0.0142735f $X=1.185 $Y=2.485 $X2=0
+ $Y2=0
cc_437 N_VPWR_c_548_n N_A_117_368#_c_637_n 0.0146352f $X=3.87 $Y=3.33 $X2=0
+ $Y2=0
cc_438 N_VPWR_c_539_n N_A_117_368#_c_637_n 0.0120433f $X=7.92 $Y=3.33 $X2=0
+ $Y2=0
cc_439 N_VPWR_c_543_n N_A_117_368#_c_638_n 0.0141475f $X=4.035 $Y=2.78 $X2=0
+ $Y2=0
cc_440 N_VPWR_c_548_n N_A_117_368#_c_638_n 0.0762741f $X=3.87 $Y=3.33 $X2=0
+ $Y2=0
cc_441 N_VPWR_c_539_n N_A_117_368#_c_638_n 0.0637471f $X=7.92 $Y=3.33 $X2=0
+ $Y2=0
cc_442 N_VPWR_c_541_n N_A_117_368#_c_639_n 0.0771921f $X=0.285 $Y=1.985 $X2=0
+ $Y2=0
cc_443 N_VPWR_M1017_d N_Y_c_695_n 0.00737459f $X=3.835 $Y=1.84 $X2=0 $Y2=0
cc_444 N_VPWR_c_543_n N_Y_c_695_n 0.0218609f $X=4.035 $Y=2.78 $X2=0 $Y2=0
cc_445 N_VPWR_c_539_n N_Y_c_695_n 0.00766693f $X=7.92 $Y=3.33 $X2=0 $Y2=0
cc_446 N_VPWR_M1017_d N_Y_c_700_n 0.00792585f $X=3.835 $Y=1.84 $X2=0 $Y2=0
cc_447 N_VPWR_M1017_d N_Y_c_715_n 0.00158596f $X=3.835 $Y=1.84 $X2=0 $Y2=0
cc_448 N_VPWR_M1012_d N_Y_c_715_n 0.00373566f $X=4.835 $Y=1.84 $X2=0 $Y2=0
cc_449 N_VPWR_c_543_n N_Y_c_715_n 8.26031e-19 $X=4.035 $Y=2.78 $X2=0 $Y2=0
cc_450 N_VPWR_M1017_d N_Y_c_701_n 0.0102791f $X=3.835 $Y=1.84 $X2=0 $Y2=0
cc_451 N_VPWR_M1024_d N_Y_c_691_n 0.0115832f $X=7.635 $Y=1.84 $X2=0 $Y2=0
cc_452 N_VPWR_c_546_n N_Y_c_691_n 0.0258342f $X=7.835 $Y=2.455 $X2=0 $Y2=0
cc_453 N_VPWR_M1024_d N_Y_c_688_n 0.00183644f $X=7.635 $Y=1.84 $X2=0 $Y2=0
cc_454 N_VPWR_M1012_d N_A_877_368#_c_835_n 0.00401812f $X=4.835 $Y=1.84 $X2=0
+ $Y2=0
cc_455 N_VPWR_c_544_n N_A_877_368#_c_835_n 0.0154669f $X=4.985 $Y=2.755 $X2=0
+ $Y2=0
cc_456 N_VPWR_c_550_n N_A_877_368#_c_829_n 0.0460938f $X=7.67 $Y=3.33 $X2=0
+ $Y2=0
cc_457 N_VPWR_c_539_n N_A_877_368#_c_829_n 0.0260732f $X=7.92 $Y=3.33 $X2=0
+ $Y2=0
cc_458 N_VPWR_c_544_n N_A_877_368#_c_830_n 0.0114567f $X=4.985 $Y=2.755 $X2=0
+ $Y2=0
cc_459 N_VPWR_c_550_n N_A_877_368#_c_830_n 0.0179217f $X=7.67 $Y=3.33 $X2=0
+ $Y2=0
cc_460 N_VPWR_c_539_n N_A_877_368#_c_830_n 0.00971942f $X=7.92 $Y=3.33 $X2=0
+ $Y2=0
cc_461 N_VPWR_c_546_n N_A_877_368#_c_831_n 0.0119239f $X=7.835 $Y=2.455 $X2=0
+ $Y2=0
cc_462 N_VPWR_c_550_n N_A_877_368#_c_831_n 0.0677651f $X=7.67 $Y=3.33 $X2=0
+ $Y2=0
cc_463 N_VPWR_c_539_n N_A_877_368#_c_831_n 0.0377062f $X=7.92 $Y=3.33 $X2=0
+ $Y2=0
cc_464 N_VPWR_c_543_n N_A_877_368#_c_832_n 0.0127976f $X=4.035 $Y=2.78 $X2=0
+ $Y2=0
cc_465 N_VPWR_c_544_n N_A_877_368#_c_832_n 0.0302025f $X=4.985 $Y=2.755 $X2=0
+ $Y2=0
cc_466 N_VPWR_c_549_n N_A_877_368#_c_832_n 0.014552f $X=4.9 $Y=3.33 $X2=0 $Y2=0
cc_467 N_VPWR_c_539_n N_A_877_368#_c_832_n 0.0119791f $X=7.92 $Y=3.33 $X2=0
+ $Y2=0
cc_468 N_VPWR_c_550_n N_A_877_368#_c_833_n 0.0121867f $X=7.67 $Y=3.33 $X2=0
+ $Y2=0
cc_469 N_VPWR_c_539_n N_A_877_368#_c_833_n 0.00660921f $X=7.92 $Y=3.33 $X2=0
+ $Y2=0
cc_470 N_VPWR_c_541_n N_A_27_74#_c_885_n 0.00886035f $X=0.285 $Y=1.985 $X2=0
+ $Y2=0
cc_471 N_A_117_368#_c_638_n N_Y_M1008_s 0.00255805f $X=3.535 $Y=2.78 $X2=0 $Y2=0
cc_472 N_A_117_368#_c_638_n N_Y_M1010_s 0.00202102f $X=3.535 $Y=2.78 $X2=0 $Y2=0
cc_473 N_A_117_368#_M1009_d N_Y_c_695_n 0.00393711f $X=2.485 $Y=1.84 $X2=0 $Y2=0
cc_474 N_A_117_368#_M1014_d N_Y_c_695_n 0.00505538f $X=3.385 $Y=1.84 $X2=0 $Y2=0
cc_475 N_A_117_368#_c_638_n N_Y_c_695_n 0.072617f $X=3.535 $Y=2.78 $X2=0 $Y2=0
cc_476 N_A_117_368#_c_638_n N_Y_c_703_n 0.0199219f $X=3.535 $Y=2.78 $X2=0 $Y2=0
cc_477 N_Y_c_715_n N_A_877_368#_M1001_s 0.00373084f $X=5.77 $Y=1.935 $X2=-0.19
+ $Y2=-0.245
cc_478 N_Y_c_715_n N_A_877_368#_M1015_s 0.00552655f $X=5.77 $Y=1.935 $X2=0 $Y2=0
cc_479 N_Y_c_746_n N_A_877_368#_M1022_d 0.00422016f $X=6.67 $Y=2.035 $X2=0 $Y2=0
cc_480 N_Y_c_691_n N_A_877_368#_M1030_d 0.0103516f $X=7.9 $Y=2.035 $X2=0 $Y2=0
cc_481 N_Y_c_715_n N_A_877_368#_c_835_n 0.0327933f $X=5.77 $Y=1.935 $X2=0 $Y2=0
cc_482 N_Y_c_715_n N_A_877_368#_c_869_n 0.0185498f $X=5.77 $Y=1.935 $X2=0 $Y2=0
cc_483 N_Y_c_729_n N_A_877_368#_c_869_n 0.0123817f $X=5.935 $Y=2.015 $X2=0 $Y2=0
cc_484 N_Y_c_729_n N_A_877_368#_c_843_n 0.0251101f $X=5.935 $Y=2.015 $X2=0 $Y2=0
cc_485 N_Y_M1018_s N_A_877_368#_c_829_n 0.00197722f $X=5.785 $Y=1.84 $X2=0 $Y2=0
cc_486 N_Y_c_729_n N_A_877_368#_c_829_n 0.0160777f $X=5.935 $Y=2.015 $X2=0 $Y2=0
cc_487 N_Y_c_746_n N_A_877_368#_c_874_n 0.0136682f $X=6.67 $Y=2.035 $X2=0 $Y2=0
cc_488 N_Y_c_729_n N_A_877_368#_c_874_n 0.0289859f $X=5.935 $Y=2.015 $X2=0 $Y2=0
cc_489 N_Y_c_735_n N_A_877_368#_c_874_n 0.0289859f $X=6.835 $Y=2.115 $X2=0 $Y2=0
cc_490 N_Y_M1027_s N_A_877_368#_c_831_n 0.00208352f $X=6.685 $Y=1.84 $X2=0 $Y2=0
cc_491 N_Y_c_735_n N_A_877_368#_c_831_n 0.0161263f $X=6.835 $Y=2.115 $X2=0 $Y2=0
cc_492 N_Y_c_691_n N_A_877_368#_c_839_n 0.0194114f $X=7.9 $Y=2.035 $X2=0 $Y2=0
cc_493 N_Y_c_695_n N_A_877_368#_c_832_n 0.0116309f $X=3.98 $Y=2.405 $X2=0 $Y2=0
cc_494 N_Y_c_700_n N_A_877_368#_c_832_n 0.00833538f $X=4.065 $Y=2.32 $X2=0 $Y2=0
cc_495 N_Y_c_715_n N_A_877_368#_c_832_n 0.0173337f $X=5.77 $Y=1.935 $X2=0 $Y2=0
cc_496 N_Y_c_689_n N_A_27_74#_M1016_d 5.0211e-19 $X=4.965 $Y=0.94 $X2=0 $Y2=0
cc_497 N_Y_c_690_n N_A_27_74#_M1016_d 0.00136745f $X=5.155 $Y=0.94 $X2=0 $Y2=0
cc_498 N_Y_c_731_n N_A_27_74#_M1013_d 0.00335829f $X=6.205 $Y=0.757 $X2=0 $Y2=0
cc_499 N_Y_c_767_n N_A_27_74#_M1021_d 0.00473528f $X=7.205 $Y=0.757 $X2=0 $Y2=0
cc_500 N_Y_c_687_n N_A_27_74#_M1028_d 0.0115696f $X=7.9 $Y=0.835 $X2=0 $Y2=0
cc_501 N_Y_c_688_n N_A_27_74#_M1028_d 0.00349433f $X=7.985 $Y=1.95 $X2=0 $Y2=0
cc_502 N_Y_c_689_n N_A_27_74#_c_889_n 0.01255f $X=4.965 $Y=0.94 $X2=0 $Y2=0
cc_503 N_Y_M1003_s N_A_27_74#_c_891_n 0.00245681f $X=4.37 $Y=0.37 $X2=0 $Y2=0
cc_504 N_Y_M1023_s N_A_27_74#_c_891_n 0.00180456f $X=5.3 $Y=0.37 $X2=0 $Y2=0
cc_505 N_Y_c_689_n N_A_27_74#_c_891_n 0.0444771f $X=4.965 $Y=0.94 $X2=0 $Y2=0
cc_506 N_Y_c_690_n N_A_27_74#_c_893_n 0.0444771f $X=5.155 $Y=0.94 $X2=0 $Y2=0
cc_507 N_Y_M1019_s N_A_27_74#_c_894_n 0.00251484f $X=6.16 $Y=0.37 $X2=0 $Y2=0
cc_508 N_Y_c_731_n N_A_27_74#_c_894_n 0.00265349f $X=6.205 $Y=0.757 $X2=0 $Y2=0
cc_509 N_Y_c_760_n N_A_27_74#_c_894_n 0.0185397f $X=6.535 $Y=0.757 $X2=0 $Y2=0
cc_510 N_Y_c_767_n N_A_27_74#_c_894_n 0.00247659f $X=7.205 $Y=0.757 $X2=0 $Y2=0
cc_511 N_Y_c_767_n N_A_27_74#_c_895_n 0.0191051f $X=7.205 $Y=0.757 $X2=0 $Y2=0
cc_512 N_Y_c_687_n N_A_27_74#_c_896_n 0.0254247f $X=7.9 $Y=0.835 $X2=0 $Y2=0
cc_513 N_Y_M1026_s N_A_27_74#_c_897_n 0.00250419f $X=7.16 $Y=0.37 $X2=0 $Y2=0
cc_514 N_Y_c_687_n N_A_27_74#_c_897_n 0.00440728f $X=7.9 $Y=0.835 $X2=0 $Y2=0
cc_515 N_Y_c_767_n N_A_27_74#_c_897_n 0.00247659f $X=7.205 $Y=0.757 $X2=0 $Y2=0
cc_516 N_Y_c_736_n N_A_27_74#_c_897_n 0.0185397f $X=7.535 $Y=0.757 $X2=0 $Y2=0
cc_517 N_Y_c_687_n N_VGND_c_1017_n 4.05485e-19 $X=7.9 $Y=0.835 $X2=0 $Y2=0
cc_518 N_Y_c_687_n N_VGND_c_1018_n 0.00100481f $X=7.9 $Y=0.835 $X2=0 $Y2=0
cc_519 N_A_27_74#_c_884_n N_VGND_M1000_s 0.00250873f $X=1.125 $Y=1.065 $X2=-0.19
+ $Y2=-0.245
cc_520 N_A_27_74#_c_907_n N_VGND_M1025_s 0.0114794f $X=2.055 $Y=0.925 $X2=0
+ $Y2=0
cc_521 N_A_27_74#_c_923_n N_VGND_M1004_s 0.00462121f $X=2.985 $Y=0.925 $X2=0
+ $Y2=0
cc_522 N_A_27_74#_c_889_n N_VGND_M1031_s 0.0109491f $X=3.905 $Y=0.925 $X2=0
+ $Y2=0
cc_523 N_A_27_74#_c_883_n N_VGND_c_1009_n 0.0180508f $X=0.28 $Y=0.515 $X2=0
+ $Y2=0
cc_524 N_A_27_74#_c_884_n N_VGND_c_1009_n 0.0209867f $X=1.125 $Y=1.065 $X2=0
+ $Y2=0
cc_525 N_A_27_74#_c_886_n N_VGND_c_1009_n 0.017215f $X=1.21 $Y=0.515 $X2=0 $Y2=0
cc_526 N_A_27_74#_c_886_n N_VGND_c_1010_n 0.0122975f $X=1.21 $Y=0.515 $X2=0
+ $Y2=0
cc_527 N_A_27_74#_c_907_n N_VGND_c_1010_n 0.0205261f $X=2.055 $Y=0.925 $X2=0
+ $Y2=0
cc_528 N_A_27_74#_c_887_n N_VGND_c_1010_n 0.0121972f $X=2.14 $Y=0.515 $X2=0
+ $Y2=0
cc_529 N_A_27_74#_c_887_n N_VGND_c_1011_n 0.0122975f $X=2.14 $Y=0.515 $X2=0
+ $Y2=0
cc_530 N_A_27_74#_c_923_n N_VGND_c_1011_n 0.0205261f $X=2.985 $Y=0.925 $X2=0
+ $Y2=0
cc_531 N_A_27_74#_c_888_n N_VGND_c_1011_n 0.0121972f $X=3.07 $Y=0.515 $X2=0
+ $Y2=0
cc_532 N_A_27_74#_c_888_n N_VGND_c_1012_n 0.00154841f $X=3.07 $Y=0.515 $X2=0
+ $Y2=0
cc_533 N_A_27_74#_c_889_n N_VGND_c_1012_n 0.0211672f $X=3.905 $Y=0.925 $X2=0
+ $Y2=0
cc_534 N_A_27_74#_c_890_n N_VGND_c_1012_n 0.0184532f $X=4.07 $Y=0.58 $X2=0 $Y2=0
cc_535 N_A_27_74#_c_883_n N_VGND_c_1013_n 0.0145639f $X=0.28 $Y=0.515 $X2=0
+ $Y2=0
cc_536 N_A_27_74#_c_886_n N_VGND_c_1014_n 0.0109942f $X=1.21 $Y=0.515 $X2=0
+ $Y2=0
cc_537 N_A_27_74#_c_887_n N_VGND_c_1015_n 0.0109704f $X=2.14 $Y=0.515 $X2=0
+ $Y2=0
cc_538 N_A_27_74#_c_888_n N_VGND_c_1016_n 0.0110419f $X=3.07 $Y=0.515 $X2=0
+ $Y2=0
cc_539 N_A_27_74#_c_890_n N_VGND_c_1017_n 0.023516f $X=4.07 $Y=0.58 $X2=0 $Y2=0
cc_540 N_A_27_74#_c_891_n N_VGND_c_1017_n 0.250323f $X=5.873 $Y=0.417 $X2=0
+ $Y2=0
cc_541 N_A_27_74#_c_883_n N_VGND_c_1018_n 0.0119984f $X=0.28 $Y=0.515 $X2=0
+ $Y2=0
cc_542 N_A_27_74#_c_886_n N_VGND_c_1018_n 0.00904371f $X=1.21 $Y=0.515 $X2=0
+ $Y2=0
cc_543 N_A_27_74#_c_907_n N_VGND_c_1018_n 0.0113663f $X=2.055 $Y=0.925 $X2=0
+ $Y2=0
cc_544 N_A_27_74#_c_887_n N_VGND_c_1018_n 0.00903439f $X=2.14 $Y=0.515 $X2=0
+ $Y2=0
cc_545 N_A_27_74#_c_923_n N_VGND_c_1018_n 0.0113542f $X=2.985 $Y=0.925 $X2=0
+ $Y2=0
cc_546 N_A_27_74#_c_888_n N_VGND_c_1018_n 0.00915013f $X=3.07 $Y=0.515 $X2=0
+ $Y2=0
cc_547 N_A_27_74#_c_889_n N_VGND_c_1018_n 0.010844f $X=3.905 $Y=0.925 $X2=0
+ $Y2=0
cc_548 N_A_27_74#_c_890_n N_VGND_c_1018_n 0.0126466f $X=4.07 $Y=0.58 $X2=0 $Y2=0
cc_549 N_A_27_74#_c_891_n N_VGND_c_1018_n 0.139412f $X=5.873 $Y=0.417 $X2=0
+ $Y2=0
