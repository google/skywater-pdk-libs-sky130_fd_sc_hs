* NGSPICE file created from sky130_fd_sc_hs__sdfrbp_2.ext - technology: sky130A

.subckt sky130_fd_sc_hs__sdfrbp_2 CLK D RESET_B SCD SCE VGND VNB VPB VPWR Q Q_N
M1000 a_1223_118# a_1025_74# a_388_79# VPB pshort w=420000u l=150000u
+  ad=2.436e+11p pd=2.84e+06u as=6.808e+11p ps=5.72e+06u
M1001 a_1401_118# a_1370_289# a_1323_118# VNB nlowvt w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=1.008e+11p ps=1.32e+06u
M1002 a_2000_74# a_852_74# a_1790_74# VNB nlowvt w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=4.33e+11p ps=3.08e+06u
M1003 a_1370_289# a_1223_118# VGND VNB nlowvt w=640000u l=150000u
+  ad=1.792e+11p pd=1.84e+06u as=2.1894e+12p ps=1.849e+07u
M1004 VGND CLK a_852_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1005 VPWR SCD a_538_464# VPB pshort w=640000u l=150000u
+  ad=3.4579e+12p pd=2.698e+07u as=1.728e+11p ps=1.82e+06u
M1006 a_1025_74# a_852_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1007 a_307_464# SCE VPWR VPB pshort w=640000u l=150000u
+  ad=1.728e+11p pd=1.82e+06u as=0p ps=0u
M1008 a_1325_457# a_852_74# a_1223_118# VPB pshort w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=0p ps=0u
M1009 a_1955_471# a_1025_74# a_1790_74# VPB pshort w=420000u l=150000u
+  ad=1.134e+11p pd=1.38e+06u as=4.029e+11p ps=3.28e+06u
M1010 a_2604_392# a_1790_74# VGND VNB nlowvt w=640000u l=150000u
+  ad=1.696e+11p pd=1.81e+06u as=0p ps=0u
M1011 a_1370_289# a_1223_118# VPWR VPB pshort w=1e+06u l=150000u
+  ad=3e+11p pd=2.6e+06u as=0p ps=0u
M1012 VGND RESET_B a_1401_118# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_1223_118# RESET_B VPWR VPB pshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_310_79# a_27_79# a_223_79# VNB nlowvt w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=2.835e+11p ps=3.03e+06u
M1015 a_223_79# SCD a_547_79# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1016 a_1790_74# a_852_74# a_1370_289# VPB pshort w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 Q_N a_1790_74# VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=3.36e+11p pd=2.84e+06u as=0p ps=0u
M1018 a_2006_373# a_1790_74# a_2158_74# VNB nlowvt w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=8.82e+10p ps=1.26e+06u
M1019 a_1223_118# a_852_74# a_388_79# VNB nlowvt w=420000u l=150000u
+  ad=1.47e+11p pd=1.54e+06u as=3.906e+11p ps=3.54e+06u
M1020 a_1323_118# a_1025_74# a_1223_118# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 VPWR a_1790_74# Q_N VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 VPWR CLK a_852_74# VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=3.304e+11p ps=2.83e+06u
M1023 VPWR SCE a_27_79# VPB pshort w=640000u l=150000u
+  ad=0p pd=0u as=1.888e+11p ps=1.87e+06u
M1024 a_1790_74# a_1025_74# a_1370_289# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 Q a_2604_392# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.072e+11p pd=2.04e+06u as=0p ps=0u
M1026 a_538_464# a_27_79# a_388_79# VPB pshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 a_2158_74# RESET_B VGND VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1028 Q_N a_1790_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.072e+11p pd=2.04e+06u as=0p ps=0u
M1029 a_388_79# D a_310_79# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1030 Q a_2604_392# VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=3.36e+11p pd=2.84e+06u as=0p ps=0u
M1031 VPWR a_2604_392# Q VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1032 a_1025_74# a_852_74# VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=3.08e+11p pd=2.79e+06u as=0p ps=0u
M1033 VGND SCE a_27_79# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.197e+11p ps=1.41e+06u
M1034 a_547_79# SCE a_388_79# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1035 a_388_79# D a_307_464# VPB pshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1036 a_2006_373# RESET_B VPWR VPB pshort w=420000u l=150000u
+  ad=1.26e+11p pd=1.44e+06u as=0p ps=0u
M1037 VPWR a_1370_289# a_1325_457# VPB pshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1038 VPWR a_2006_373# a_1955_471# VPB pshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1039 VGND a_1790_74# Q_N VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1040 VGND a_2604_392# Q VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1041 VPWR a_1790_74# a_2006_373# VPB pshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1042 a_2604_392# a_1790_74# VPWR VPB pshort w=1e+06u l=150000u
+  ad=2.75e+11p pd=2.55e+06u as=0p ps=0u
M1043 VGND RESET_B a_223_79# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1044 a_388_79# RESET_B VPWR VPB pshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1045 VGND a_2006_373# a_2000_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

