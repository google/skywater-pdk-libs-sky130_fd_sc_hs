* File: sky130_fd_sc_hs__a2111oi_2.pxi.spice
* Created: Tue Sep  1 19:48:12 2020
* 
x_PM_SKY130_FD_SC_HS__A2111OI_2%D1 N_D1_c_92_n N_D1_M1008_g N_D1_M1007_g
+ N_D1_c_93_n N_D1_M1009_g D1 D1 N_D1_c_91_n PM_SKY130_FD_SC_HS__A2111OI_2%D1
x_PM_SKY130_FD_SC_HS__A2111OI_2%C1 N_C1_M1001_g N_C1_c_131_n N_C1_M1011_g
+ N_C1_c_132_n N_C1_M1014_g C1 C1 C1 N_C1_c_130_n
+ PM_SKY130_FD_SC_HS__A2111OI_2%C1
x_PM_SKY130_FD_SC_HS__A2111OI_2%B1 N_B1_c_171_n N_B1_M1010_g N_B1_c_172_n
+ N_B1_c_173_n N_B1_c_176_n N_B1_M1015_g N_B1_c_177_n N_B1_M1016_g B1 B1
+ N_B1_c_175_n PM_SKY130_FD_SC_HS__A2111OI_2%B1
x_PM_SKY130_FD_SC_HS__A2111OI_2%A1 N_A1_c_224_n N_A1_M1000_g N_A1_M1003_g
+ N_A1_c_225_n N_A1_M1002_g N_A1_M1013_g A1 A1 N_A1_c_223_n
+ PM_SKY130_FD_SC_HS__A2111OI_2%A1
x_PM_SKY130_FD_SC_HS__A2111OI_2%A2 N_A2_M1005_g N_A2_c_279_n N_A2_M1004_g
+ N_A2_M1012_g N_A2_c_280_n N_A2_M1006_g A2 N_A2_c_277_n N_A2_c_278_n
+ PM_SKY130_FD_SC_HS__A2111OI_2%A2
x_PM_SKY130_FD_SC_HS__A2111OI_2%A_69_368# N_A_69_368#_M1008_s
+ N_A_69_368#_M1009_s N_A_69_368#_M1014_s N_A_69_368#_c_313_n
+ N_A_69_368#_c_314_n N_A_69_368#_c_315_n N_A_69_368#_c_321_n
+ N_A_69_368#_c_316_n N_A_69_368#_c_317_n N_A_69_368#_c_318_n
+ PM_SKY130_FD_SC_HS__A2111OI_2%A_69_368#
x_PM_SKY130_FD_SC_HS__A2111OI_2%Y N_Y_M1007_d N_Y_M1010_d N_Y_M1003_s
+ N_Y_M1008_d N_Y_c_349_n N_Y_c_350_n N_Y_c_364_n N_Y_c_359_n N_Y_c_351_n
+ N_Y_c_352_n N_Y_c_353_n N_Y_c_354_n N_Y_c_367_n N_Y_c_355_n N_Y_c_356_n
+ N_Y_c_357_n Y Y PM_SKY130_FD_SC_HS__A2111OI_2%Y
x_PM_SKY130_FD_SC_HS__A2111OI_2%A_334_368# N_A_334_368#_M1011_d
+ N_A_334_368#_M1015_d N_A_334_368#_c_422_n N_A_334_368#_c_426_n
+ N_A_334_368#_c_423_n PM_SKY130_FD_SC_HS__A2111OI_2%A_334_368#
x_PM_SKY130_FD_SC_HS__A2111OI_2%A_533_368# N_A_533_368#_M1015_s
+ N_A_533_368#_M1016_s N_A_533_368#_M1002_s N_A_533_368#_M1006_s
+ N_A_533_368#_c_449_n N_A_533_368#_c_450_n N_A_533_368#_c_451_n
+ N_A_533_368#_c_458_n N_A_533_368#_c_460_n N_A_533_368#_c_466_n
+ N_A_533_368#_c_452_n N_A_533_368#_c_475_n N_A_533_368#_c_453_n
+ N_A_533_368#_c_454_n N_A_533_368#_c_472_n
+ PM_SKY130_FD_SC_HS__A2111OI_2%A_533_368#
x_PM_SKY130_FD_SC_HS__A2111OI_2%VPWR N_VPWR_M1000_d N_VPWR_M1004_d
+ N_VPWR_c_508_n N_VPWR_c_509_n VPWR N_VPWR_c_510_n N_VPWR_c_511_n
+ N_VPWR_c_512_n N_VPWR_c_507_n N_VPWR_c_514_n N_VPWR_c_515_n
+ PM_SKY130_FD_SC_HS__A2111OI_2%VPWR
x_PM_SKY130_FD_SC_HS__A2111OI_2%VGND N_VGND_M1007_s N_VGND_M1001_d
+ N_VGND_M1005_s N_VGND_c_566_n N_VGND_c_567_n N_VGND_c_568_n N_VGND_c_569_n
+ VGND N_VGND_c_570_n N_VGND_c_571_n N_VGND_c_572_n N_VGND_c_573_n
+ N_VGND_c_574_n N_VGND_c_575_n PM_SKY130_FD_SC_HS__A2111OI_2%VGND
x_PM_SKY130_FD_SC_HS__A2111OI_2%A_722_74# N_A_722_74#_M1003_d
+ N_A_722_74#_M1013_d N_A_722_74#_M1012_d N_A_722_74#_c_619_n
+ N_A_722_74#_c_620_n N_A_722_74#_c_621_n N_A_722_74#_c_622_n
+ N_A_722_74#_c_623_n PM_SKY130_FD_SC_HS__A2111OI_2%A_722_74#
cc_1 VNB N_D1_M1007_g 0.0296222f $X=-0.19 $Y=-0.245 $X2=1.04 $Y2=0.74
cc_2 VNB D1 0.00551793f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.58
cc_3 VNB N_D1_c_91_n 0.0482427f $X=-0.19 $Y=-0.245 $X2=1.13 $Y2=1.515
cc_4 VNB N_C1_M1001_g 0.0273389f $X=-0.19 $Y=-0.245 $X2=0.695 $Y2=2.4
cc_5 VNB C1 0.0165977f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_6 VNB N_C1_c_130_n 0.0370211f $X=-0.19 $Y=-0.245 $X2=1.145 $Y2=1.557
cc_7 VNB N_B1_c_171_n 0.0201467f $X=-0.19 $Y=-0.245 $X2=0.695 $Y2=1.765
cc_8 VNB N_B1_c_172_n 0.0446588f $X=-0.19 $Y=-0.245 $X2=1.04 $Y2=1.35
cc_9 VNB N_B1_c_173_n 0.00913645f $X=-0.19 $Y=-0.245 $X2=1.04 $Y2=0.74
cc_10 VNB B1 0.0124371f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_B1_c_175_n 0.0681176f $X=-0.19 $Y=-0.245 $X2=1.13 $Y2=1.515
cc_12 VNB N_A1_M1003_g 0.0295402f $X=-0.19 $Y=-0.245 $X2=1.04 $Y2=0.74
cc_13 VNB N_A1_M1013_g 0.024081f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB A1 0.00589944f $X=-0.19 $Y=-0.245 $X2=1.04 $Y2=1.557
cc_15 VNB N_A1_c_223_n 0.0346751f $X=-0.19 $Y=-0.245 $X2=1.13 $Y2=1.565
cc_16 VNB N_A2_M1005_g 0.023157f $X=-0.19 $Y=-0.245 $X2=0.695 $Y2=2.4
cc_17 VNB N_A2_M1012_g 0.0320221f $X=-0.19 $Y=-0.245 $X2=1.145 $Y2=2.4
cc_18 VNB N_A2_c_277_n 0.00102489f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.565
cc_19 VNB N_A2_c_278_n 0.0472696f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_Y_c_349_n 0.0238079f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_Y_c_350_n 0.0177372f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_Y_c_351_n 0.00327056f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.565
cc_23 VNB N_Y_c_352_n 0.00305444f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_Y_c_353_n 0.0188906f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_Y_c_354_n 0.0355113f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_Y_c_355_n 0.00821167f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_Y_c_356_n 0.0108587f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_Y_c_357_n 0.00250929f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB Y 0.025793f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_VPWR_c_507_n 0.243291f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_566_n 0.0274256f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_567_n 0.0184856f $X=-0.19 $Y=-0.245 $X2=1.04 $Y2=1.557
cc_33 VNB N_VGND_c_568_n 0.00917051f $X=-0.19 $Y=-0.245 $X2=1.145 $Y2=1.557
cc_34 VNB N_VGND_c_569_n 0.00396562f $X=-0.19 $Y=-0.245 $X2=1.13 $Y2=1.565
cc_35 VNB N_VGND_c_570_n 0.0795701f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_571_n 0.0178682f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_572_n 0.348653f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_573_n 0.0293037f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_574_n 0.00653982f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_575_n 0.00622543f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_722_74#_c_619_n 0.016287f $X=-0.19 $Y=-0.245 $X2=1.145 $Y2=2.4
cc_42 VNB N_A_722_74#_c_620_n 0.0016059f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_722_74#_c_621_n 0.0172894f $X=-0.19 $Y=-0.245 $X2=1.13 $Y2=1.515
cc_44 VNB N_A_722_74#_c_622_n 0.00250711f $X=-0.19 $Y=-0.245 $X2=1.13 $Y2=1.515
cc_45 VNB N_A_722_74#_c_623_n 0.0270834f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VPB N_D1_c_92_n 0.017242f $X=-0.19 $Y=1.66 $X2=0.695 $Y2=1.765
cc_47 VPB N_D1_c_93_n 0.0147911f $X=-0.19 $Y=1.66 $X2=1.145 $Y2=1.765
cc_48 VPB D1 0.00779977f $X=-0.19 $Y=1.66 $X2=1.115 $Y2=1.58
cc_49 VPB N_D1_c_91_n 0.0223493f $X=-0.19 $Y=1.66 $X2=1.13 $Y2=1.515
cc_50 VPB N_C1_c_131_n 0.0147911f $X=-0.19 $Y=1.66 $X2=1.04 $Y2=0.74
cc_51 VPB N_C1_c_132_n 0.0186669f $X=-0.19 $Y=1.66 $X2=1.145 $Y2=1.765
cc_52 VPB C1 0.0133825f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_53 VPB N_C1_c_130_n 0.0206438f $X=-0.19 $Y=1.66 $X2=1.145 $Y2=1.557
cc_54 VPB N_B1_c_176_n 0.0185418f $X=-0.19 $Y=1.66 $X2=1.04 $Y2=0.74
cc_55 VPB N_B1_c_177_n 0.0149057f $X=-0.19 $Y=1.66 $X2=1.145 $Y2=2.4
cc_56 VPB N_B1_c_175_n 0.0139017f $X=-0.19 $Y=1.66 $X2=1.13 $Y2=1.515
cc_57 VPB N_A1_c_224_n 0.0153195f $X=-0.19 $Y=1.66 $X2=0.695 $Y2=1.765
cc_58 VPB N_A1_c_225_n 0.0157847f $X=-0.19 $Y=1.66 $X2=1.145 $Y2=1.765
cc_59 VPB A1 0.00584804f $X=-0.19 $Y=1.66 $X2=1.04 $Y2=1.557
cc_60 VPB N_A1_c_223_n 0.0194941f $X=-0.19 $Y=1.66 $X2=1.13 $Y2=1.565
cc_61 VPB N_A2_c_279_n 0.0153712f $X=-0.19 $Y=1.66 $X2=1.04 $Y2=0.74
cc_62 VPB N_A2_c_280_n 0.0198958f $X=-0.19 $Y=1.66 $X2=1.115 $Y2=1.58
cc_63 VPB N_A2_c_277_n 0.00283943f $X=-0.19 $Y=1.66 $X2=0.72 $Y2=1.565
cc_64 VPB N_A2_c_278_n 0.0230699f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_65 VPB N_A_69_368#_c_313_n 0.0233684f $X=-0.19 $Y=1.66 $X2=1.115 $Y2=1.58
cc_66 VPB N_A_69_368#_c_314_n 0.0030474f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_67 VPB N_A_69_368#_c_315_n 0.00939918f $X=-0.19 $Y=1.66 $X2=0.695 $Y2=1.557
cc_68 VPB N_A_69_368#_c_316_n 0.0067982f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_69 VPB N_A_69_368#_c_317_n 0.00584978f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_70 VPB N_A_69_368#_c_318_n 0.00123754f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_71 VPB N_Y_c_359_n 0.0160034f $X=-0.19 $Y=1.66 $X2=1.04 $Y2=1.557
cc_72 VPB Y 0.0142074f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_73 VPB N_A_334_368#_c_422_n 0.0110263f $X=-0.19 $Y=1.66 $X2=1.145 $Y2=2.4
cc_74 VPB N_A_334_368#_c_423_n 0.00246895f $X=-0.19 $Y=1.66 $X2=1.04 $Y2=1.557
cc_75 VPB N_A_533_368#_c_449_n 0.00585892f $X=-0.19 $Y=1.66 $X2=0.695 $Y2=1.557
cc_76 VPB N_A_533_368#_c_450_n 0.00456202f $X=-0.19 $Y=1.66 $X2=1.13 $Y2=1.557
cc_77 VPB N_A_533_368#_c_451_n 0.00396918f $X=-0.19 $Y=1.66 $X2=1.13 $Y2=1.515
cc_78 VPB N_A_533_368#_c_452_n 0.00216998f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_79 VPB N_A_533_368#_c_453_n 0.0171433f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_80 VPB N_A_533_368#_c_454_n 0.0345863f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_81 VPB N_VPWR_c_508_n 0.00705934f $X=-0.19 $Y=1.66 $X2=1.145 $Y2=2.4
cc_82 VPB N_VPWR_c_509_n 0.00339119f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_83 VPB N_VPWR_c_510_n 0.0986568f $X=-0.19 $Y=1.66 $X2=1.13 $Y2=1.557
cc_84 VPB N_VPWR_c_511_n 0.0185125f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_85 VPB N_VPWR_c_512_n 0.0177091f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_86 VPB N_VPWR_c_507_n 0.0932175f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_87 VPB N_VPWR_c_514_n 0.00324402f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_88 VPB N_VPWR_c_515_n 0.00601644f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_89 N_D1_M1007_g N_C1_M1001_g 0.0207626f $X=1.04 $Y=0.74 $X2=0 $Y2=0
cc_90 N_D1_c_93_n N_C1_c_131_n 0.0127228f $X=1.145 $Y=1.765 $X2=0 $Y2=0
cc_91 D1 C1 0.0352545f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_92 N_D1_c_91_n C1 4.84655e-19 $X=1.13 $Y=1.515 $X2=0 $Y2=0
cc_93 D1 N_C1_c_130_n 0.00163028f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_94 N_D1_c_91_n N_C1_c_130_n 0.0255576f $X=1.13 $Y=1.515 $X2=0 $Y2=0
cc_95 N_D1_c_92_n N_A_69_368#_c_314_n 0.0137046f $X=0.695 $Y=1.765 $X2=0 $Y2=0
cc_96 N_D1_c_93_n N_A_69_368#_c_314_n 0.0128006f $X=1.145 $Y=1.765 $X2=0 $Y2=0
cc_97 D1 N_A_69_368#_c_321_n 0.00256352f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_98 N_D1_M1007_g N_Y_c_349_n 0.0169004f $X=1.04 $Y=0.74 $X2=0 $Y2=0
cc_99 D1 N_Y_c_349_n 0.0419733f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_100 N_D1_c_91_n N_Y_c_349_n 0.00987898f $X=1.13 $Y=1.515 $X2=0 $Y2=0
cc_101 N_D1_c_92_n N_Y_c_364_n 0.0136569f $X=0.695 $Y=1.765 $X2=0 $Y2=0
cc_102 D1 N_Y_c_364_n 0.0104662f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_103 N_D1_M1007_g N_Y_c_351_n 0.00383226f $X=1.04 $Y=0.74 $X2=0 $Y2=0
cc_104 N_D1_c_92_n N_Y_c_367_n 0.0134092f $X=0.695 $Y=1.765 $X2=0 $Y2=0
cc_105 N_D1_c_93_n N_Y_c_367_n 0.00918116f $X=1.145 $Y=1.765 $X2=0 $Y2=0
cc_106 D1 N_Y_c_367_n 0.0237598f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_107 N_D1_c_91_n N_Y_c_367_n 0.00144727f $X=1.13 $Y=1.515 $X2=0 $Y2=0
cc_108 D1 N_Y_c_355_n 0.0133987f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_109 N_D1_c_91_n N_Y_c_355_n 0.00339787f $X=1.13 $Y=1.515 $X2=0 $Y2=0
cc_110 N_D1_c_92_n Y 0.00555197f $X=0.695 $Y=1.765 $X2=0 $Y2=0
cc_111 N_D1_M1007_g Y 0.00380025f $X=1.04 $Y=0.74 $X2=0 $Y2=0
cc_112 D1 Y 0.0263051f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_113 N_D1_c_91_n Y 0.00275245f $X=1.13 $Y=1.515 $X2=0 $Y2=0
cc_114 N_D1_c_92_n N_VPWR_c_510_n 0.00278271f $X=0.695 $Y=1.765 $X2=0 $Y2=0
cc_115 N_D1_c_93_n N_VPWR_c_510_n 0.00278271f $X=1.145 $Y=1.765 $X2=0 $Y2=0
cc_116 N_D1_c_92_n N_VPWR_c_507_n 0.00357798f $X=0.695 $Y=1.765 $X2=0 $Y2=0
cc_117 N_D1_c_93_n N_VPWR_c_507_n 0.00353907f $X=1.145 $Y=1.765 $X2=0 $Y2=0
cc_118 N_D1_M1007_g N_VGND_c_566_n 0.0129243f $X=1.04 $Y=0.74 $X2=0 $Y2=0
cc_119 N_D1_M1007_g N_VGND_c_567_n 0.00383152f $X=1.04 $Y=0.74 $X2=0 $Y2=0
cc_120 N_D1_M1007_g N_VGND_c_572_n 0.00758569f $X=1.04 $Y=0.74 $X2=0 $Y2=0
cc_121 N_C1_M1001_g N_B1_c_171_n 0.0247539f $X=1.58 $Y=0.74 $X2=-0.19 $Y2=-0.245
cc_122 C1 N_B1_c_173_n 0.0170771f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_123 N_C1_c_130_n N_B1_c_173_n 0.00495638f $X=1.67 $Y=1.515 $X2=0 $Y2=0
cc_124 C1 N_B1_c_176_n 5.49627e-19 $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_125 C1 B1 0.0132423f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_126 C1 N_B1_c_175_n 0.0145426f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_127 N_C1_c_131_n N_A_69_368#_c_316_n 0.0127563f $X=1.595 $Y=1.765 $X2=0 $Y2=0
cc_128 N_C1_c_132_n N_A_69_368#_c_316_n 0.0137046f $X=2.045 $Y=1.765 $X2=0 $Y2=0
cc_129 N_C1_M1001_g N_Y_c_351_n 5.52855e-19 $X=1.58 $Y=0.74 $X2=0 $Y2=0
cc_130 N_C1_M1001_g N_Y_c_352_n 0.0145564f $X=1.58 $Y=0.74 $X2=0 $Y2=0
cc_131 C1 N_Y_c_352_n 0.0514073f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_132 N_C1_c_130_n N_Y_c_352_n 0.00514858f $X=1.67 $Y=1.515 $X2=0 $Y2=0
cc_133 N_C1_M1001_g N_Y_c_353_n 8.24518e-19 $X=1.58 $Y=0.74 $X2=0 $Y2=0
cc_134 C1 N_Y_c_354_n 0.0120661f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_135 C1 N_Y_c_356_n 0.0294457f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_136 N_C1_c_132_n N_A_334_368#_c_422_n 0.0138963f $X=2.045 $Y=1.765 $X2=0
+ $Y2=0
cc_137 C1 N_A_334_368#_c_422_n 0.0586847f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_138 N_C1_c_131_n N_A_334_368#_c_426_n 0.00918116f $X=1.595 $Y=1.765 $X2=0
+ $Y2=0
cc_139 N_C1_c_132_n N_A_334_368#_c_426_n 0.0134092f $X=2.045 $Y=1.765 $X2=0
+ $Y2=0
cc_140 C1 N_A_334_368#_c_426_n 0.0237597f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_141 N_C1_c_130_n N_A_334_368#_c_426_n 0.00162844f $X=1.67 $Y=1.515 $X2=0
+ $Y2=0
cc_142 N_C1_c_132_n N_A_533_368#_c_451_n 5.67935e-19 $X=2.045 $Y=1.765 $X2=0
+ $Y2=0
cc_143 N_C1_c_131_n N_VPWR_c_510_n 0.00278271f $X=1.595 $Y=1.765 $X2=0 $Y2=0
cc_144 N_C1_c_132_n N_VPWR_c_510_n 0.00278271f $X=2.045 $Y=1.765 $X2=0 $Y2=0
cc_145 N_C1_c_131_n N_VPWR_c_507_n 0.00353907f $X=1.595 $Y=1.765 $X2=0 $Y2=0
cc_146 N_C1_c_132_n N_VPWR_c_507_n 0.00358624f $X=2.045 $Y=1.765 $X2=0 $Y2=0
cc_147 N_C1_M1001_g N_VGND_c_566_n 4.50149e-19 $X=1.58 $Y=0.74 $X2=0 $Y2=0
cc_148 N_C1_M1001_g N_VGND_c_567_n 0.00461464f $X=1.58 $Y=0.74 $X2=0 $Y2=0
cc_149 N_C1_M1001_g N_VGND_c_568_n 0.00279591f $X=1.58 $Y=0.74 $X2=0 $Y2=0
cc_150 N_C1_M1001_g N_VGND_c_572_n 0.0090927f $X=1.58 $Y=0.74 $X2=0 $Y2=0
cc_151 N_B1_c_177_n N_A1_c_224_n 0.00960549f $X=3.465 $Y=1.765 $X2=-0.19
+ $Y2=-0.245
cc_152 B1 N_A1_M1003_g 0.00481817f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_153 N_B1_c_175_n N_A1_M1003_g 0.00561135f $X=3.39 $Y=1.385 $X2=0 $Y2=0
cc_154 B1 A1 0.0132858f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_155 N_B1_c_175_n A1 0.001199f $X=3.39 $Y=1.385 $X2=0 $Y2=0
cc_156 B1 N_A1_c_223_n 0.00199478f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_157 N_B1_c_175_n N_A1_c_223_n 0.0206493f $X=3.39 $Y=1.385 $X2=0 $Y2=0
cc_158 N_B1_c_176_n N_A_69_368#_c_316_n 5.67935e-19 $X=3.015 $Y=1.765 $X2=0
+ $Y2=0
cc_159 N_B1_c_171_n N_Y_c_352_n 0.0116603f $X=2.12 $Y=1.185 $X2=0 $Y2=0
cc_160 N_B1_c_171_n N_Y_c_353_n 0.00612384f $X=2.12 $Y=1.185 $X2=0 $Y2=0
cc_161 N_B1_c_172_n N_Y_c_354_n 0.0141305f $X=2.925 $Y=1.26 $X2=0 $Y2=0
cc_162 B1 N_Y_c_354_n 0.0503328f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_163 N_B1_c_175_n N_Y_c_354_n 0.00370328f $X=3.39 $Y=1.385 $X2=0 $Y2=0
cc_164 N_B1_c_171_n N_Y_c_356_n 0.00662344f $X=2.12 $Y=1.185 $X2=0 $Y2=0
cc_165 N_B1_c_172_n N_Y_c_356_n 0.00744713f $X=2.925 $Y=1.26 $X2=0 $Y2=0
cc_166 N_B1_c_172_n N_A_334_368#_c_422_n 0.00376848f $X=2.925 $Y=1.26 $X2=0
+ $Y2=0
cc_167 N_B1_c_176_n N_A_334_368#_c_422_n 0.0164789f $X=3.015 $Y=1.765 $X2=0
+ $Y2=0
cc_168 B1 N_A_334_368#_c_422_n 0.00251507f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_169 N_B1_c_176_n N_A_334_368#_c_423_n 0.0195587f $X=3.015 $Y=1.765 $X2=0
+ $Y2=0
cc_170 N_B1_c_177_n N_A_334_368#_c_423_n 0.00657118f $X=3.465 $Y=1.765 $X2=0
+ $Y2=0
cc_171 B1 N_A_334_368#_c_423_n 0.0149843f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_172 N_B1_c_175_n N_A_334_368#_c_423_n 0.00250027f $X=3.39 $Y=1.385 $X2=0
+ $Y2=0
cc_173 N_B1_c_176_n N_A_533_368#_c_450_n 0.0137046f $X=3.015 $Y=1.765 $X2=0
+ $Y2=0
cc_174 N_B1_c_177_n N_A_533_368#_c_450_n 0.0125587f $X=3.465 $Y=1.765 $X2=0
+ $Y2=0
cc_175 N_B1_c_177_n N_A_533_368#_c_458_n 0.00205467f $X=3.465 $Y=1.765 $X2=0
+ $Y2=0
cc_176 B1 N_A_533_368#_c_458_n 0.00744503f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_177 N_B1_c_176_n N_A_533_368#_c_460_n 7.1895e-19 $X=3.015 $Y=1.765 $X2=0
+ $Y2=0
cc_178 N_B1_c_177_n N_A_533_368#_c_460_n 0.00956952f $X=3.465 $Y=1.765 $X2=0
+ $Y2=0
cc_179 N_B1_c_176_n N_VPWR_c_510_n 0.00278271f $X=3.015 $Y=1.765 $X2=0 $Y2=0
cc_180 N_B1_c_177_n N_VPWR_c_510_n 0.00278257f $X=3.465 $Y=1.765 $X2=0 $Y2=0
cc_181 N_B1_c_176_n N_VPWR_c_507_n 0.00358624f $X=3.015 $Y=1.765 $X2=0 $Y2=0
cc_182 N_B1_c_177_n N_VPWR_c_507_n 0.00353905f $X=3.465 $Y=1.765 $X2=0 $Y2=0
cc_183 N_B1_c_171_n N_VGND_c_568_n 0.00602646f $X=2.12 $Y=1.185 $X2=0 $Y2=0
cc_184 N_B1_c_171_n N_VGND_c_570_n 0.00434272f $X=2.12 $Y=1.185 $X2=0 $Y2=0
cc_185 N_B1_c_171_n N_VGND_c_572_n 0.00826088f $X=2.12 $Y=1.185 $X2=0 $Y2=0
cc_186 N_A1_M1013_g N_A2_M1005_g 0.019323f $X=4.38 $Y=0.74 $X2=0 $Y2=0
cc_187 N_A1_c_225_n N_A2_c_279_n 0.00908392f $X=4.365 $Y=1.765 $X2=0 $Y2=0
cc_188 A1 N_A2_c_277_n 0.0353991f $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_189 N_A1_c_223_n N_A2_c_277_n 3.04398e-19 $X=4.365 $Y=1.557 $X2=0 $Y2=0
cc_190 A1 N_A2_c_278_n 0.0038932f $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_191 N_A1_c_223_n N_A2_c_278_n 0.0190382f $X=4.365 $Y=1.557 $X2=0 $Y2=0
cc_192 N_A1_M1003_g N_Y_c_354_n 0.0149884f $X=3.95 $Y=0.74 $X2=0 $Y2=0
cc_193 A1 N_Y_c_354_n 0.00137046f $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_194 N_A1_M1003_g N_Y_c_357_n 0.00878264f $X=3.95 $Y=0.74 $X2=0 $Y2=0
cc_195 N_A1_M1013_g N_Y_c_357_n 0.00464929f $X=4.38 $Y=0.74 $X2=0 $Y2=0
cc_196 A1 N_Y_c_357_n 0.0218587f $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_197 N_A1_c_223_n N_Y_c_357_n 0.00221794f $X=4.365 $Y=1.557 $X2=0 $Y2=0
cc_198 N_A1_c_224_n N_A_533_368#_c_450_n 0.0032261f $X=3.915 $Y=1.765 $X2=0
+ $Y2=0
cc_199 N_A1_c_224_n N_A_533_368#_c_458_n 9.1767e-19 $X=3.915 $Y=1.765 $X2=0
+ $Y2=0
cc_200 N_A1_c_224_n N_A_533_368#_c_460_n 0.00944051f $X=3.915 $Y=1.765 $X2=0
+ $Y2=0
cc_201 N_A1_c_225_n N_A_533_368#_c_460_n 6.22492e-19 $X=4.365 $Y=1.765 $X2=0
+ $Y2=0
cc_202 N_A1_c_224_n N_A_533_368#_c_466_n 0.0153029f $X=3.915 $Y=1.765 $X2=0
+ $Y2=0
cc_203 N_A1_c_225_n N_A_533_368#_c_466_n 0.0120074f $X=4.365 $Y=1.765 $X2=0
+ $Y2=0
cc_204 A1 N_A_533_368#_c_466_n 0.0313954f $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_205 N_A1_c_223_n N_A_533_368#_c_466_n 0.00130859f $X=4.365 $Y=1.557 $X2=0
+ $Y2=0
cc_206 N_A1_c_224_n N_A_533_368#_c_452_n 6.47982e-19 $X=3.915 $Y=1.765 $X2=0
+ $Y2=0
cc_207 N_A1_c_225_n N_A_533_368#_c_452_n 0.0104832f $X=4.365 $Y=1.765 $X2=0
+ $Y2=0
cc_208 N_A1_c_225_n N_A_533_368#_c_472_n 4.27055e-19 $X=4.365 $Y=1.765 $X2=0
+ $Y2=0
cc_209 A1 N_A_533_368#_c_472_n 0.0193938f $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_210 N_A1_c_224_n N_VPWR_c_508_n 0.00331651f $X=3.915 $Y=1.765 $X2=0 $Y2=0
cc_211 N_A1_c_225_n N_VPWR_c_508_n 0.00366706f $X=4.365 $Y=1.765 $X2=0 $Y2=0
cc_212 N_A1_c_225_n N_VPWR_c_509_n 5.55114e-19 $X=4.365 $Y=1.765 $X2=0 $Y2=0
cc_213 N_A1_c_224_n N_VPWR_c_510_n 0.0044313f $X=3.915 $Y=1.765 $X2=0 $Y2=0
cc_214 N_A1_c_225_n N_VPWR_c_511_n 0.00445602f $X=4.365 $Y=1.765 $X2=0 $Y2=0
cc_215 N_A1_c_224_n N_VPWR_c_507_n 0.00853445f $X=3.915 $Y=1.765 $X2=0 $Y2=0
cc_216 N_A1_c_225_n N_VPWR_c_507_n 0.00857673f $X=4.365 $Y=1.765 $X2=0 $Y2=0
cc_217 N_A1_M1013_g N_VGND_c_569_n 6.35092e-19 $X=4.38 $Y=0.74 $X2=0 $Y2=0
cc_218 N_A1_M1003_g N_VGND_c_570_n 0.00291649f $X=3.95 $Y=0.74 $X2=0 $Y2=0
cc_219 N_A1_M1013_g N_VGND_c_570_n 0.00291649f $X=4.38 $Y=0.74 $X2=0 $Y2=0
cc_220 N_A1_M1003_g N_VGND_c_572_n 0.00363173f $X=3.95 $Y=0.74 $X2=0 $Y2=0
cc_221 N_A1_M1013_g N_VGND_c_572_n 0.00359219f $X=4.38 $Y=0.74 $X2=0 $Y2=0
cc_222 N_A1_M1003_g N_A_722_74#_c_619_n 0.010283f $X=3.95 $Y=0.74 $X2=0 $Y2=0
cc_223 N_A1_M1013_g N_A_722_74#_c_619_n 0.0142063f $X=4.38 $Y=0.74 $X2=0 $Y2=0
cc_224 N_A1_M1013_g N_A_722_74#_c_622_n 0.00174382f $X=4.38 $Y=0.74 $X2=0 $Y2=0
cc_225 A1 N_A_722_74#_c_622_n 0.0148778f $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_226 N_A2_c_279_n N_A_533_368#_c_452_n 0.00614488f $X=4.815 $Y=1.765 $X2=0
+ $Y2=0
cc_227 N_A2_c_279_n N_A_533_368#_c_475_n 0.0160432f $X=4.815 $Y=1.765 $X2=0
+ $Y2=0
cc_228 N_A2_c_280_n N_A_533_368#_c_475_n 0.0171961f $X=5.265 $Y=1.765 $X2=0
+ $Y2=0
cc_229 N_A2_c_277_n N_A_533_368#_c_475_n 0.0222295f $X=5.015 $Y=1.515 $X2=0
+ $Y2=0
cc_230 N_A2_c_278_n N_A_533_368#_c_475_n 0.00130746f $X=5.25 $Y=1.557 $X2=0
+ $Y2=0
cc_231 N_A2_c_280_n N_A_533_368#_c_453_n 0.00314968f $X=5.265 $Y=1.765 $X2=0
+ $Y2=0
cc_232 N_A2_c_280_n N_A_533_368#_c_454_n 0.00729586f $X=5.265 $Y=1.765 $X2=0
+ $Y2=0
cc_233 N_A2_c_279_n N_VPWR_c_509_n 0.0114128f $X=4.815 $Y=1.765 $X2=0 $Y2=0
cc_234 N_A2_c_280_n N_VPWR_c_509_n 0.0143569f $X=5.265 $Y=1.765 $X2=0 $Y2=0
cc_235 N_A2_c_279_n N_VPWR_c_511_n 0.00413917f $X=4.815 $Y=1.765 $X2=0 $Y2=0
cc_236 N_A2_c_280_n N_VPWR_c_512_n 0.00413917f $X=5.265 $Y=1.765 $X2=0 $Y2=0
cc_237 N_A2_c_279_n N_VPWR_c_507_n 0.0081781f $X=4.815 $Y=1.765 $X2=0 $Y2=0
cc_238 N_A2_c_280_n N_VPWR_c_507_n 0.00821187f $X=5.265 $Y=1.765 $X2=0 $Y2=0
cc_239 N_A2_M1005_g N_VGND_c_569_n 0.0108748f $X=4.81 $Y=0.74 $X2=0 $Y2=0
cc_240 N_A2_M1012_g N_VGND_c_569_n 0.0137776f $X=5.25 $Y=0.74 $X2=0 $Y2=0
cc_241 N_A2_M1005_g N_VGND_c_570_n 0.00383152f $X=4.81 $Y=0.74 $X2=0 $Y2=0
cc_242 N_A2_M1012_g N_VGND_c_571_n 0.00383152f $X=5.25 $Y=0.74 $X2=0 $Y2=0
cc_243 N_A2_M1005_g N_VGND_c_572_n 0.00757637f $X=4.81 $Y=0.74 $X2=0 $Y2=0
cc_244 N_A2_M1012_g N_VGND_c_572_n 0.00761248f $X=5.25 $Y=0.74 $X2=0 $Y2=0
cc_245 N_A2_M1005_g N_A_722_74#_c_621_n 0.0164896f $X=4.81 $Y=0.74 $X2=0 $Y2=0
cc_246 N_A2_M1012_g N_A_722_74#_c_621_n 0.0180492f $X=5.25 $Y=0.74 $X2=0 $Y2=0
cc_247 N_A2_c_277_n N_A_722_74#_c_621_n 0.0251424f $X=5.015 $Y=1.515 $X2=0 $Y2=0
cc_248 N_A2_c_278_n N_A_722_74#_c_621_n 0.00216008f $X=5.25 $Y=1.557 $X2=0 $Y2=0
cc_249 N_A2_M1012_g N_A_722_74#_c_623_n 0.00159319f $X=5.25 $Y=0.74 $X2=0 $Y2=0
cc_250 N_A_69_368#_c_314_n N_Y_M1008_d 0.00197722f $X=1.285 $Y=2.99 $X2=0 $Y2=0
cc_251 N_A_69_368#_M1008_s N_Y_c_364_n 0.0111275f $X=0.345 $Y=1.84 $X2=0 $Y2=0
cc_252 N_A_69_368#_c_313_n N_Y_c_364_n 0.0161539f $X=0.47 $Y=2.455 $X2=0 $Y2=0
cc_253 N_A_69_368#_c_313_n N_Y_c_359_n 0.00451074f $X=0.47 $Y=2.455 $X2=0 $Y2=0
cc_254 N_A_69_368#_c_313_n N_Y_c_367_n 0.0298377f $X=0.47 $Y=2.455 $X2=0 $Y2=0
cc_255 N_A_69_368#_c_314_n N_Y_c_367_n 0.0160777f $X=1.285 $Y=2.99 $X2=0 $Y2=0
cc_256 N_A_69_368#_c_321_n N_Y_c_367_n 0.051802f $X=1.37 $Y=2.115 $X2=0 $Y2=0
cc_257 N_A_69_368#_M1008_s Y 0.00146477f $X=0.345 $Y=1.84 $X2=0 $Y2=0
cc_258 N_A_69_368#_c_316_n N_A_334_368#_M1011_d 0.00197722f $X=2.185 $Y=2.99
+ $X2=-0.19 $Y2=1.66
cc_259 N_A_69_368#_M1014_s N_A_334_368#_c_422_n 0.00558057f $X=2.12 $Y=1.84
+ $X2=0 $Y2=0
cc_260 N_A_69_368#_c_317_n N_A_334_368#_c_422_n 0.0202979f $X=2.27 $Y=2.455
+ $X2=0 $Y2=0
cc_261 N_A_69_368#_c_321_n N_A_334_368#_c_426_n 0.051802f $X=1.37 $Y=2.115 $X2=0
+ $Y2=0
cc_262 N_A_69_368#_c_316_n N_A_334_368#_c_426_n 0.0160777f $X=2.185 $Y=2.99
+ $X2=0 $Y2=0
cc_263 N_A_69_368#_c_317_n N_A_334_368#_c_426_n 0.0298377f $X=2.27 $Y=2.455
+ $X2=0 $Y2=0
cc_264 N_A_69_368#_c_317_n N_A_533_368#_c_449_n 0.0457258f $X=2.27 $Y=2.455
+ $X2=0 $Y2=0
cc_265 N_A_69_368#_c_316_n N_A_533_368#_c_451_n 0.0147157f $X=2.185 $Y=2.99
+ $X2=0 $Y2=0
cc_266 N_A_69_368#_c_314_n N_VPWR_c_510_n 0.0460938f $X=1.285 $Y=2.99 $X2=0
+ $Y2=0
cc_267 N_A_69_368#_c_315_n N_VPWR_c_510_n 0.0179217f $X=0.555 $Y=2.99 $X2=0
+ $Y2=0
cc_268 N_A_69_368#_c_316_n N_VPWR_c_510_n 0.0640155f $X=2.185 $Y=2.99 $X2=0
+ $Y2=0
cc_269 N_A_69_368#_c_318_n N_VPWR_c_510_n 0.0121867f $X=1.37 $Y=2.99 $X2=0 $Y2=0
cc_270 N_A_69_368#_c_314_n N_VPWR_c_507_n 0.0260732f $X=1.285 $Y=2.99 $X2=0
+ $Y2=0
cc_271 N_A_69_368#_c_315_n N_VPWR_c_507_n 0.00971942f $X=0.555 $Y=2.99 $X2=0
+ $Y2=0
cc_272 N_A_69_368#_c_316_n N_VPWR_c_507_n 0.0357926f $X=2.185 $Y=2.99 $X2=0
+ $Y2=0
cc_273 N_A_69_368#_c_318_n N_VPWR_c_507_n 0.00660921f $X=1.37 $Y=2.99 $X2=0
+ $Y2=0
cc_274 N_Y_c_349_n N_VGND_M1007_s 0.00299905f $X=1.16 $Y=1.095 $X2=-0.19
+ $Y2=-0.245
cc_275 N_Y_c_352_n N_VGND_M1001_d 0.00309832f $X=2.17 $Y=1.095 $X2=0 $Y2=0
cc_276 N_Y_c_349_n N_VGND_c_566_n 0.0219406f $X=1.16 $Y=1.095 $X2=0 $Y2=0
cc_277 N_Y_c_351_n N_VGND_c_566_n 0.0191765f $X=1.325 $Y=0.515 $X2=0 $Y2=0
cc_278 N_Y_c_351_n N_VGND_c_567_n 0.0146357f $X=1.325 $Y=0.515 $X2=0 $Y2=0
cc_279 N_Y_c_351_n N_VGND_c_568_n 0.00158453f $X=1.325 $Y=0.515 $X2=0 $Y2=0
cc_280 N_Y_c_352_n N_VGND_c_568_n 0.022455f $X=2.17 $Y=1.095 $X2=0 $Y2=0
cc_281 N_Y_c_353_n N_VGND_c_568_n 0.0191425f $X=2.335 $Y=0.515 $X2=0 $Y2=0
cc_282 N_Y_c_353_n N_VGND_c_570_n 0.0145639f $X=2.335 $Y=0.515 $X2=0 $Y2=0
cc_283 N_Y_c_351_n N_VGND_c_572_n 0.0121141f $X=1.325 $Y=0.515 $X2=0 $Y2=0
cc_284 N_Y_c_353_n N_VGND_c_572_n 0.0119984f $X=2.335 $Y=0.515 $X2=0 $Y2=0
cc_285 N_Y_c_354_n N_VGND_c_572_n 0.0406621f $X=4 $Y=0.872 $X2=0 $Y2=0
cc_286 N_Y_c_354_n N_A_722_74#_M1003_d 0.00838011f $X=4 $Y=0.872 $X2=-0.19
+ $Y2=-0.245
cc_287 N_Y_M1003_s N_A_722_74#_c_619_n 0.00178571f $X=4.025 $Y=0.37 $X2=0 $Y2=0
cc_288 N_Y_c_354_n N_A_722_74#_c_619_n 0.0268535f $X=4 $Y=0.872 $X2=0 $Y2=0
cc_289 N_Y_c_357_n N_A_722_74#_c_619_n 0.0161432f $X=4.165 $Y=0.872 $X2=0 $Y2=0
cc_290 N_Y_c_357_n N_A_722_74#_c_622_n 0.00517071f $X=4.165 $Y=0.872 $X2=0 $Y2=0
cc_291 N_A_334_368#_c_422_n N_A_533_368#_M1015_s 0.00625313f $X=3.075 $Y=2.035
+ $X2=-0.19 $Y2=1.66
cc_292 N_A_334_368#_c_422_n N_A_533_368#_c_449_n 0.0210301f $X=3.075 $Y=2.035
+ $X2=0 $Y2=0
cc_293 N_A_334_368#_M1015_d N_A_533_368#_c_450_n 0.00218679f $X=3.09 $Y=1.84
+ $X2=0 $Y2=0
cc_294 N_A_334_368#_c_423_n N_A_533_368#_c_450_n 0.0144323f $X=3.24 $Y=1.985
+ $X2=0 $Y2=0
cc_295 N_A_334_368#_c_423_n N_A_533_368#_c_458_n 0.013092f $X=3.24 $Y=1.985
+ $X2=0 $Y2=0
cc_296 N_A_334_368#_c_423_n N_A_533_368#_c_460_n 0.0411694f $X=3.24 $Y=1.985
+ $X2=0 $Y2=0
cc_297 N_A_533_368#_c_466_n N_VPWR_M1000_d 0.00408911f $X=4.425 $Y=2.035
+ $X2=-0.19 $Y2=1.66
cc_298 N_A_533_368#_c_475_n N_VPWR_M1004_d 0.00359006f $X=5.405 $Y=2.035 $X2=0
+ $Y2=0
cc_299 N_A_533_368#_c_450_n N_VPWR_c_508_n 0.0119328f $X=3.525 $Y=2.99 $X2=0
+ $Y2=0
cc_300 N_A_533_368#_c_460_n N_VPWR_c_508_n 0.0400262f $X=3.69 $Y=2.815 $X2=0
+ $Y2=0
cc_301 N_A_533_368#_c_466_n N_VPWR_c_508_n 0.0136682f $X=4.425 $Y=2.035 $X2=0
+ $Y2=0
cc_302 N_A_533_368#_c_452_n N_VPWR_c_508_n 0.0440249f $X=4.59 $Y=2.445 $X2=0
+ $Y2=0
cc_303 N_A_533_368#_c_452_n N_VPWR_c_509_n 0.0462948f $X=4.59 $Y=2.445 $X2=0
+ $Y2=0
cc_304 N_A_533_368#_c_475_n N_VPWR_c_509_n 0.0171813f $X=5.405 $Y=2.035 $X2=0
+ $Y2=0
cc_305 N_A_533_368#_c_454_n N_VPWR_c_509_n 0.0462948f $X=5.49 $Y=2.4 $X2=0 $Y2=0
cc_306 N_A_533_368#_c_450_n N_VPWR_c_510_n 0.0626055f $X=3.525 $Y=2.99 $X2=0
+ $Y2=0
cc_307 N_A_533_368#_c_451_n N_VPWR_c_510_n 0.0200723f $X=2.905 $Y=2.99 $X2=0
+ $Y2=0
cc_308 N_A_533_368#_c_452_n N_VPWR_c_511_n 0.0110241f $X=4.59 $Y=2.445 $X2=0
+ $Y2=0
cc_309 N_A_533_368#_c_454_n N_VPWR_c_512_n 0.011066f $X=5.49 $Y=2.4 $X2=0 $Y2=0
cc_310 N_A_533_368#_c_450_n N_VPWR_c_507_n 0.0346986f $X=3.525 $Y=2.99 $X2=0
+ $Y2=0
cc_311 N_A_533_368#_c_451_n N_VPWR_c_507_n 0.0108858f $X=2.905 $Y=2.99 $X2=0
+ $Y2=0
cc_312 N_A_533_368#_c_452_n N_VPWR_c_507_n 0.00909194f $X=4.59 $Y=2.445 $X2=0
+ $Y2=0
cc_313 N_A_533_368#_c_454_n N_VPWR_c_507_n 0.00915947f $X=5.49 $Y=2.4 $X2=0
+ $Y2=0
cc_314 N_A_533_368#_c_453_n N_A_722_74#_c_621_n 0.00831718f $X=5.53 $Y=2.12
+ $X2=0 $Y2=0
cc_315 N_VGND_c_570_n N_A_722_74#_c_619_n 0.038121f $X=4.86 $Y=0 $X2=0 $Y2=0
cc_316 N_VGND_c_572_n N_A_722_74#_c_619_n 0.0321651f $X=5.52 $Y=0 $X2=0 $Y2=0
cc_317 N_VGND_c_569_n N_A_722_74#_c_620_n 0.00989215f $X=5.03 $Y=0.675 $X2=0
+ $Y2=0
cc_318 N_VGND_c_570_n N_A_722_74#_c_620_n 0.00758556f $X=4.86 $Y=0 $X2=0 $Y2=0
cc_319 N_VGND_c_572_n N_A_722_74#_c_620_n 0.00627867f $X=5.52 $Y=0 $X2=0 $Y2=0
cc_320 N_VGND_M1005_s N_A_722_74#_c_621_n 0.00187091f $X=4.885 $Y=0.37 $X2=0
+ $Y2=0
cc_321 N_VGND_c_569_n N_A_722_74#_c_621_n 0.0178913f $X=5.03 $Y=0.675 $X2=0
+ $Y2=0
cc_322 N_VGND_c_569_n N_A_722_74#_c_623_n 0.0183707f $X=5.03 $Y=0.675 $X2=0
+ $Y2=0
cc_323 N_VGND_c_571_n N_A_722_74#_c_623_n 0.011066f $X=5.52 $Y=0 $X2=0 $Y2=0
cc_324 N_VGND_c_572_n N_A_722_74#_c_623_n 0.00915947f $X=5.52 $Y=0 $X2=0 $Y2=0
