* File: sky130_fd_sc_hs__fa_4.spice
* Created: Tue Sep  1 20:05:32 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hs__fa_4.pex.spice"
.subckt sky130_fd_sc_hs__fa_4  VNB VPB B CIN A VPWR SUM COUT VGND
* 
* VGND	VGND
* COUT	COUT
* SUM	SUM
* VPWR	VPWR
* A	A
* CIN	CIN
* B	B
* VPB	VPB
* VNB	VNB
MM1029 N_VGND_M1029_d N_A_M1029_g N_A_27_74#_M1029_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.39435 AS=0.2109 PD=1.87 PS=2.05 NRD=77.496 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75010.1 A=0.111 P=1.78 MULT=1
MM1025 N_A_27_74#_M1025_d N_B_M1025_g N_VGND_M1029_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.39435 PD=1.02 PS=1.87 NRD=0 NRS=77.496 M=1 R=4.93333 SA=75001.3
+ SB=75009 A=0.111 P=1.78 MULT=1
MM1004 N_A_418_74#_M1004_d N_CIN_M1004_g N_A_27_74#_M1025_d VNB NLOWVT L=0.15
+ W=0.74 AD=0.1554 AS=0.1036 PD=1.16 PS=1.02 NRD=11.34 NRS=0 M=1 R=4.93333
+ SA=75001.7 SB=75008.5 A=0.111 P=1.78 MULT=1
MM1019 A_532_74# N_B_M1019_g N_A_418_74#_M1004_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.1443 AS=0.1554 PD=1.13 PS=1.16 NRD=22.692 NRS=11.34 M=1 R=4.93333
+ SA=75002.3 SB=75008 A=0.111 P=1.78 MULT=1
MM1030 N_VGND_M1030_d N_A_M1030_g A_532_74# VNB NLOWVT L=0.15 W=0.74 AD=0.1184
+ AS=0.1443 PD=1.06 PS=1.13 NRD=0 NRS=22.692 M=1 R=4.93333 SA=75002.8 SB=75007.4
+ A=0.111 P=1.78 MULT=1
MM1026 N_A_734_74#_M1026_d N_CIN_M1026_g N_VGND_M1030_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1184 PD=1.02 PS=1.06 NRD=0 NRS=6.48 M=1 R=4.93333 SA=75003.3
+ SB=75007 A=0.111 P=1.78 MULT=1
MM1027 N_VGND_M1027_d N_B_M1027_g N_A_734_74#_M1026_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.19035 AS=0.1036 PD=1.37 PS=1.02 NRD=32.784 NRS=0 M=1 R=4.93333 SA=75003.7
+ SB=75006.5 A=0.111 P=1.78 MULT=1
MM1012 N_A_734_74#_M1012_d N_A_M1012_g N_VGND_M1027_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.19035 PD=1.02 PS=1.37 NRD=0 NRS=32.784 M=1 R=4.93333 SA=75004.3
+ SB=75005.9 A=0.111 P=1.78 MULT=1
MM1013 N_A_1024_74#_M1013_d N_A_418_74#_M1013_g N_A_734_74#_M1012_d VNB NLOWVT
+ L=0.15 W=0.74 AD=0.1961 AS=0.1036 PD=1.27 PS=1.02 NRD=40.536 NRS=0 M=1
+ R=4.93333 SA=75004.8 SB=75005.5 A=0.111 P=1.78 MULT=1
MM1022 A_1160_74# N_CIN_M1022_g N_A_1024_74#_M1013_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.0888 AS=0.1961 PD=0.98 PS=1.27 NRD=10.536 NRS=0 M=1 R=4.93333 SA=75005.4
+ SB=75004.8 A=0.111 P=1.78 MULT=1
MM1039 A_1238_74# N_B_M1039_g A_1160_74# VNB NLOWVT L=0.15 W=0.74 AD=0.1332
+ AS=0.0888 PD=1.1 PS=0.98 NRD=20.268 NRS=10.536 M=1 R=4.93333 SA=75005.8
+ SB=75004.4 A=0.111 P=1.78 MULT=1
MM1005 N_VGND_M1005_d N_A_M1005_g A_1238_74# VNB NLOWVT L=0.15 W=0.74 AD=0.19385
+ AS=0.1332 PD=1.41 PS=1.1 NRD=13.776 NRS=20.268 M=1 R=4.93333 SA=75006.3
+ SB=75003.9 A=0.111 P=1.78 MULT=1
MM1016 N_VGND_M1005_d N_A_1024_74#_M1016_g N_SUM_M1016_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.19385 AS=0.1036 PD=1.41 PS=1.02 NRD=33.552 NRS=0 M=1 R=4.93333
+ SA=75006.6 SB=75003.5 A=0.111 P=1.78 MULT=1
MM1017 N_VGND_M1017_d N_A_1024_74#_M1017_g N_SUM_M1016_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.19615 AS=0.1036 PD=1.41 PS=1.02 NRD=34.056 NRS=0 M=1 R=4.93333
+ SA=75007 SB=75003.1 A=0.111 P=1.78 MULT=1
MM1032 N_VGND_M1017_d N_A_1024_74#_M1032_g N_SUM_M1032_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.19615 AS=0.1036 PD=1.41 PS=1.02 NRD=34.056 NRS=0 M=1 R=4.93333
+ SA=75007.6 SB=75002.5 A=0.111 P=1.78 MULT=1
MM1035 N_VGND_M1035_d N_A_1024_74#_M1035_g N_SUM_M1032_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.19615 AS=0.1036 PD=1.41 PS=1.02 NRD=34.056 NRS=0 M=1 R=4.93333
+ SA=75008 SB=75002.1 A=0.111 P=1.78 MULT=1
MM1010 N_COUT_M1010_d N_A_418_74#_M1010_g N_VGND_M1035_d VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.19615 PD=1.02 PS=1.41 NRD=0 NRS=34.056 M=1 R=4.93333
+ SA=75008.6 SB=75001.5 A=0.111 P=1.78 MULT=1
MM1011 N_COUT_M1010_d N_A_418_74#_M1011_g N_VGND_M1011_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75009
+ SB=75001.1 A=0.111 P=1.78 MULT=1
MM1018 N_COUT_M1018_d N_A_418_74#_M1018_g N_VGND_M1011_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75009.5 SB=75000.6 A=0.111 P=1.78 MULT=1
MM1033 N_COUT_M1018_d N_A_418_74#_M1033_g N_VGND_M1033_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.2109 PD=1.02 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75009.9 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1009 N_VPWR_M1009_d N_A_M1009_g N_A_27_392#_M1009_s VPB PSHORT L=0.15 W=1
+ AD=0.253375 AS=0.295 PD=1.725 PS=2.59 NRD=1.9503 NRS=1.9503 M=1 R=6.66667
+ SA=75000.2 SB=75007.9 A=0.15 P=2.3 MULT=1
MM1023 N_A_27_392#_M1023_d N_B_M1023_g N_VPWR_M1009_d VPB PSHORT L=0.15 W=1
+ AD=0.490662 AS=0.253375 PD=2.05 PS=1.725 NRD=85.8132 NRS=15.2478 M=1 R=6.66667
+ SA=75000.7 SB=75009.1 A=0.15 P=2.3 MULT=1
MM1036 N_A_418_74#_M1036_d N_CIN_M1036_g N_A_27_392#_M1023_d VPB PSHORT L=0.15
+ W=1 AD=0.15 AS=0.490662 PD=1.3 PS=2.05 NRD=0 NRS=85.8132 M=1 R=6.66667
+ SA=75001.7 SB=75008.1 A=0.15 P=2.3 MULT=1
MM1002 A_535_347# N_B_M1002_g N_A_418_74#_M1036_d VPB PSHORT L=0.15 W=1 AD=0.18
+ AS=0.15 PD=1.36 PS=1.3 NRD=24.6053 NRS=1.9503 M=1 R=6.66667 SA=75002.2
+ SB=75007.6 A=0.15 P=2.3 MULT=1
MM1015 N_VPWR_M1015_d N_A_M1015_g A_535_347# VPB PSHORT L=0.15 W=1 AD=0.175
+ AS=0.18 PD=1.35 PS=1.36 NRD=1.9503 NRS=24.6053 M=1 R=6.66667 SA=75002.7
+ SB=75007.1 A=0.15 P=2.3 MULT=1
MM1014 N_A_737_347#_M1014_d N_CIN_M1014_g N_VPWR_M1015_d VPB PSHORT L=0.15 W=1
+ AD=0.15 AS=0.175 PD=1.3 PS=1.35 NRD=1.9503 NRS=11.8003 M=1 R=6.66667
+ SA=75003.2 SB=75006.6 A=0.15 P=2.3 MULT=1
MM1021 N_VPWR_M1021_d N_B_M1021_g N_A_737_347#_M1014_d VPB PSHORT L=0.15 W=1
+ AD=0.21 AS=0.15 PD=1.42 PS=1.3 NRD=18.715 NRS=1.9503 M=1 R=6.66667 SA=75003.6
+ SB=75006.2 A=0.15 P=2.3 MULT=1
MM1028 N_A_737_347#_M1028_d N_A_M1028_g N_VPWR_M1021_d VPB PSHORT L=0.15 W=1
+ AD=0.175 AS=0.21 PD=1.35 PS=1.42 NRD=11.8003 NRS=8.8453 M=1 R=6.66667
+ SA=75004.2 SB=75005.6 A=0.15 P=2.3 MULT=1
MM1000 N_A_1024_74#_M1000_d N_A_418_74#_M1000_g N_A_737_347#_M1028_d VPB PSHORT
+ L=0.15 W=1 AD=0.175 AS=0.175 PD=1.35 PS=1.35 NRD=11.8003 NRS=1.9503 M=1
+ R=6.66667 SA=75004.7 SB=75005.1 A=0.15 P=2.3 MULT=1
MM1037 A_1141_347# N_CIN_M1037_g N_A_1024_74#_M1000_d VPB PSHORT L=0.15 W=1
+ AD=0.16 AS=0.175 PD=1.32 PS=1.35 NRD=20.6653 NRS=1.9503 M=1 R=6.66667
+ SA=75005.2 SB=75004.6 A=0.15 P=2.3 MULT=1
MM1006 A_1235_347# N_B_M1006_g A_1141_347# VPB PSHORT L=0.15 W=1 AD=0.20235
+ AS=0.16 PD=1.495 PS=1.32 NRD=29.0181 NRS=20.6653 M=1 R=6.66667 SA=75005.7
+ SB=75004.1 A=0.15 P=2.3 MULT=1
MM1024 N_VPWR_M1024_d N_A_M1024_g A_1235_347# VPB PSHORT L=0.15 W=1 AD=0.203019
+ AS=0.20235 PD=1.42925 PS=1.495 NRD=21.1578 NRS=29.0181 M=1 R=6.66667
+ SA=75005.6 SB=75004.1 A=0.15 P=2.3 MULT=1
MM1003 N_VPWR_M1024_d N_A_1024_74#_M1003_g N_SUM_M1003_s VPB PSHORT L=0.15
+ W=1.12 AD=0.227381 AS=0.168 PD=1.60075 PS=1.42 NRD=1.7533 NRS=1.7533 M=1
+ R=7.46667 SA=75005.5 SB=75003.5 A=0.168 P=2.54 MULT=1
MM1031 N_VPWR_M1031_d N_A_1024_74#_M1031_g N_SUM_M1003_s VPB PSHORT L=0.15
+ W=1.12 AD=0.196 AS=0.168 PD=1.47 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75006 SB=75003.1 A=0.168 P=2.54 MULT=1
MM1034 N_VPWR_M1031_d N_A_1024_74#_M1034_g N_SUM_M1034_s VPB PSHORT L=0.15
+ W=1.12 AD=0.196 AS=0.168 PD=1.47 PS=1.42 NRD=10.5395 NRS=1.7533 M=1 R=7.46667
+ SA=75006.5 SB=75002.6 A=0.168 P=2.54 MULT=1
MM1038 N_VPWR_M1038_d N_A_1024_74#_M1038_g N_SUM_M1034_s VPB PSHORT L=0.15
+ W=1.12 AD=0.196 AS=0.168 PD=1.47 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75006.9 SB=75002.1 A=0.168 P=2.54 MULT=1
MM1001 N_COUT_M1001_d N_A_418_74#_M1001_g N_VPWR_M1038_d VPB PSHORT L=0.15
+ W=1.12 AD=0.168 AS=0.196 PD=1.42 PS=1.47 NRD=1.7533 NRS=10.5395 M=1 R=7.46667
+ SA=75007.4 SB=75001.6 A=0.168 P=2.54 MULT=1
MM1007 N_COUT_M1001_d N_A_418_74#_M1007_g N_VPWR_M1007_s VPB PSHORT L=0.15
+ W=1.12 AD=0.168 AS=0.196 PD=1.42 PS=1.47 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75007.9 SB=75001.2 A=0.168 P=2.54 MULT=1
MM1008 N_COUT_M1008_d N_A_418_74#_M1008_g N_VPWR_M1007_s VPB PSHORT L=0.15
+ W=1.12 AD=0.168 AS=0.196 PD=1.42 PS=1.47 NRD=1.7533 NRS=10.5395 M=1 R=7.46667
+ SA=75008.4 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1020 N_COUT_M1008_d N_A_418_74#_M1020_g N_VPWR_M1020_s VPB PSHORT L=0.15
+ W=1.12 AD=0.168 AS=0.3304 PD=1.42 PS=2.83 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75008.8 SB=75000.2 A=0.168 P=2.54 MULT=1
DX40_noxref VNB VPB NWDIODE A=21.8696 P=26.77
c_94 VNB 0 9.5881e-20 $X=0 $Y=0
c_192 VPB 0 3.55722e-19 $X=0 $Y=3.085
c_1426 A_535_347# 0 1.17721e-19 $X=2.675 $Y=1.735
*
.include "sky130_fd_sc_hs__fa_4.pxi.spice"
*
.ends
*
*
