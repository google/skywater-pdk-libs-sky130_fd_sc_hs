* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hs__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
X0 X a_83_264# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X1 a_398_392# A2 a_83_264# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=150000u
X2 a_257_136# A1 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X3 a_662_136# C1 a_83_264# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X4 VPWR A1 a_398_392# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=150000u
X5 a_257_136# B1 a_662_136# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X6 a_83_264# B1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=150000u
X7 VGND A2 a_257_136# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X8 VPWR C1 a_83_264# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=150000u
X9 X a_83_264# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
.ends
