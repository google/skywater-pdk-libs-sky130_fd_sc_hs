* File: sky130_fd_sc_hs__fa_1.pex.spice
* Created: Tue Sep  1 20:05:20 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HS__FA_1%A_69_260# 1 2 9 11 13 15 16 17 18 20 24 27 30
+ 35 40
c100 24 0 7.81052e-20 $X=2.245 $Y=2.59
r101 40 42 4.36531 $w=3.28e-07 $l=1.25e-07 $layer=LI1_cond $X=2.245 $Y=1.91
+ $X2=2.245 $Y2=2.035
r102 35 37 4.01609 $w=3.28e-07 $l=1.15e-07 $layer=LI1_cond $X=2.105 $Y=0.55
+ $X2=2.105 $Y2=0.665
r103 30 32 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=1.14 $Y=1.795
+ $X2=1.14 $Y2=2.035
r104 27 29 17.3534 $w=2.32e-07 $l=3.3e-07 $layer=LI1_cond $X=0.565 $Y=1.465
+ $X2=0.565 $Y2=1.795
r105 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.51
+ $Y=1.465 $X2=0.51 $Y2=1.465
r106 22 42 2.96841 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=2.245 $Y=2.12
+ $X2=2.245 $Y2=2.035
r107 22 24 16.4136 $w=3.28e-07 $l=4.7e-07 $layer=LI1_cond $X=2.245 $Y=2.12
+ $X2=2.245 $Y2=2.59
r108 21 32 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.225 $Y=2.035
+ $X2=1.14 $Y2=2.035
r109 20 42 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.08 $Y=2.035
+ $X2=2.245 $Y2=2.035
r110 20 21 55.7807 $w=1.68e-07 $l=8.55e-07 $layer=LI1_cond $X=2.08 $Y=2.035
+ $X2=1.225 $Y2=2.035
r111 19 29 2.55969 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=0.705 $Y=1.795
+ $X2=0.565 $Y2=1.795
r112 18 30 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.055 $Y=1.795
+ $X2=1.14 $Y2=1.795
r113 18 19 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=1.055 $Y=1.795
+ $X2=0.705 $Y2=1.795
r114 16 37 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.94 $Y=0.665
+ $X2=2.105 $Y2=0.665
r115 16 17 80.5722 $w=1.68e-07 $l=1.235e-06 $layer=LI1_cond $X=1.94 $Y=0.665
+ $X2=0.705 $Y2=0.665
r116 15 27 9.57122 $w=2.32e-07 $l=1.90526e-07 $layer=LI1_cond $X=0.62 $Y=1.3
+ $X2=0.565 $Y2=1.465
r117 14 17 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.62 $Y=0.75
+ $X2=0.705 $Y2=0.665
r118 14 15 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=0.62 $Y=0.75
+ $X2=0.62 $Y2=1.3
r119 11 28 61.4066 $w=2.86e-07 $l=3.07409e-07 $layer=POLY_cond $X=0.495 $Y=1.765
+ $X2=0.51 $Y2=1.465
r120 11 13 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.495 $Y=1.765
+ $X2=0.495 $Y2=2.4
r121 7 28 38.6549 $w=2.86e-07 $l=1.72337e-07 $layer=POLY_cond $X=0.495 $Y=1.3
+ $X2=0.51 $Y2=1.465
r122 7 9 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=0.495 $Y=1.3
+ $X2=0.495 $Y2=0.74
r123 2 40 400 $w=1.7e-07 $l=2.38485e-07 $layer=licon1_PDIFF $count=1 $X=2.095
+ $Y=1.735 $X2=2.245 $Y2=1.91
r124 2 24 400 $w=1.7e-07 $l=9.26971e-07 $layer=licon1_PDIFF $count=1 $X=2.095
+ $Y=1.735 $X2=2.245 $Y2=2.59
r125 1 35 182 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_NDIFF $count=1 $X=1.965
+ $Y=0.375 $X2=2.105 $Y2=0.55
.ends

.subckt PM_SKY130_FD_SC_HS__FA_1%A 1 3 6 8 10 11 13 14 16 17 19 20 22 23 25 27
+ 28 32 35 37 40 41 45 47 51 54
c215 47 0 1.97438e-19 $X=4.545 $Y=1.012
c216 40 0 2.98399e-20 $X=5.895 $Y=1.32
c217 28 0 8.44456e-20 $X=3.3 $Y=1.005
c218 20 0 1.00637e-19 $X=6.055 $Y=1.66
r219 54 59 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.545
+ $Y=1.29 $X2=4.545 $Y2=1.29
r220 52 61 35.4412 $w=3.06e-07 $l=2.25e-07 $layer=POLY_cond $X=6.045 $Y=1.41
+ $X2=6.045 $Y2=1.185
r221 51 52 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.045
+ $Y=1.41 $X2=6.045 $Y2=1.41
r222 46 54 6.46067 $w=3.28e-07 $l=1.85e-07 $layer=LI1_cond $X=4.545 $Y=1.105
+ $X2=4.545 $Y2=1.29
r223 46 47 0.89609 $w=3.3e-07 $l=9.3e-08 $layer=LI1_cond $X=4.545 $Y=1.105
+ $X2=4.545 $Y2=1.012
r224 43 44 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.05
+ $Y=1.385 $X2=1.05 $Y2=1.385
r225 41 43 18.3968 $w=2.52e-07 $l=3.8e-07 $layer=LI1_cond $X=1.05 $Y=1.005
+ $X2=1.05 $Y2=1.385
r226 40 51 6.77908 $w=2.53e-07 $l=1.5e-07 $layer=LI1_cond $X=5.895 $Y=1.447
+ $X2=6.045 $Y2=1.447
r227 39 40 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=5.895 $Y=1.105
+ $X2=5.895 $Y2=1.32
r228 38 47 8.61065 $w=1.7e-07 $l=1.68953e-07 $layer=LI1_cond $X=4.71 $Y=1.02
+ $X2=4.545 $Y2=1.012
r229 37 39 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.81 $Y=1.02
+ $X2=5.895 $Y2=1.105
r230 37 38 71.7647 $w=1.68e-07 $l=1.1e-06 $layer=LI1_cond $X=5.81 $Y=1.02
+ $X2=4.71 $Y2=1.02
r231 36 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.63 $Y=1.005
+ $X2=3.465 $Y2=1.005
r232 35 47 8.61065 $w=1.7e-07 $l=1.68464e-07 $layer=LI1_cond $X=4.38 $Y=1.005
+ $X2=4.545 $Y2=1.012
r233 35 36 48.9305 $w=1.68e-07 $l=7.5e-07 $layer=LI1_cond $X=4.38 $Y=1.005
+ $X2=3.63 $Y2=1.005
r234 32 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.465
+ $Y=1.29 $X2=3.465 $Y2=1.29
r235 30 45 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.465 $Y=1.09
+ $X2=3.465 $Y2=1.005
r236 30 32 6.9845 $w=3.28e-07 $l=2e-07 $layer=LI1_cond $X=3.465 $Y=1.09
+ $X2=3.465 $Y2=1.29
r237 29 41 3.04159 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.215 $Y=1.005
+ $X2=1.05 $Y2=1.005
r238 28 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.3 $Y=1.005
+ $X2=3.465 $Y2=1.005
r239 28 29 136.027 $w=1.68e-07 $l=2.085e-06 $layer=LI1_cond $X=3.3 $Y=1.005
+ $X2=1.215 $Y2=1.005
r240 25 27 133.353 $w=1.5e-07 $l=4.15e-07 $layer=POLY_cond $X=6.485 $Y=1.11
+ $X2=6.485 $Y2=0.695
r241 24 61 19.4347 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.21 $Y=1.185
+ $X2=6.045 $Y2=1.185
r242 23 25 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=6.41 $Y=1.185
+ $X2=6.485 $Y2=1.11
r243 23 24 102.553 $w=1.5e-07 $l=2e-07 $layer=POLY_cond $X=6.41 $Y=1.185
+ $X2=6.21 $Y2=1.185
r244 20 52 51.9239 $w=3.06e-07 $l=2.54951e-07 $layer=POLY_cond $X=6.055 $Y=1.66
+ $X2=6.045 $Y2=1.41
r245 20 22 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=6.055 $Y=1.66
+ $X2=6.055 $Y2=2.235
r246 17 59 38.8629 $w=2.72e-07 $l=1.92678e-07 $layer=POLY_cond $X=4.605 $Y=1.125
+ $X2=4.545 $Y2=1.29
r247 17 19 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=4.605 $Y=1.125
+ $X2=4.605 $Y2=0.695
r248 14 59 75.1901 $w=2.72e-07 $l=3.89487e-07 $layer=POLY_cond $X=4.505 $Y=1.66
+ $X2=4.545 $Y2=1.29
r249 14 16 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=4.505 $Y=1.66
+ $X2=4.505 $Y2=2.235
r250 11 33 75.1901 $w=2.72e-07 $l=4.05771e-07 $layer=POLY_cond $X=3.54 $Y=1.66
+ $X2=3.465 $Y2=1.29
r251 11 13 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=3.54 $Y=1.66
+ $X2=3.54 $Y2=2.235
r252 8 33 38.8629 $w=2.72e-07 $l=1.94808e-07 $layer=POLY_cond $X=3.53 $Y=1.125
+ $X2=3.465 $Y2=1.29
r253 8 10 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=3.53 $Y=1.125
+ $X2=3.53 $Y2=0.695
r254 4 44 38.9026 $w=2.7e-07 $l=1.92678e-07 $layer=POLY_cond $X=1.11 $Y=1.22
+ $X2=1.05 $Y2=1.385
r255 4 6 269.202 $w=1.5e-07 $l=5.25e-07 $layer=POLY_cond $X=1.11 $Y=1.22
+ $X2=1.11 $Y2=0.695
r256 1 44 77.2841 $w=2.7e-07 $l=3.995e-07 $layer=POLY_cond $X=1.01 $Y=1.765
+ $X2=1.05 $Y2=1.385
r257 1 3 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=1.01 $Y=1.765
+ $X2=1.01 $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_HS__FA_1%CIN 3 5 7 10 12 14 17 19 21 22 24 27 28 29 30
+ 33 36 39 46
c170 36 0 9.44466e-20 $X=5.04 $Y=1.665
c171 28 0 1.02197e-19 $X=1.825 $Y=1.665
c172 22 0 2.98399e-20 $X=5.155 $Y=1.425
c173 3 0 8.59909e-20 $X=1.89 $Y=0.695
r174 46 51 8.27811 $w=3.53e-07 $l=2.55e-07 $layer=LI1_cond $X=4.017 $Y=1.41
+ $X2=4.017 $Y2=1.665
r175 45 46 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.005
+ $Y=1.41 $X2=4.005 $Y2=1.41
r176 42 43 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.95
+ $Y=1.41 $X2=1.95 $Y2=1.41
r177 39 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=1.665
+ $X2=4.08 $Y2=1.665
r178 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=1.665
+ $X2=5.04 $Y2=1.665
r179 33 43 8.235 $w=4e-07 $l=2.7e-07 $layer=LI1_cond $X=1.68 $Y=1.52 $X2=1.95
+ $Y2=1.52
r180 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=1.665
+ $X2=1.68 $Y2=1.665
r181 30 39 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.225 $Y=1.665
+ $X2=4.08 $Y2=1.665
r182 29 36 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.895 $Y=1.665
+ $X2=5.04 $Y2=1.665
r183 29 30 0.829206 $w=1.4e-07 $l=6.7e-07 $layer=MET1_cond $X=4.895 $Y=1.665
+ $X2=4.225 $Y2=1.665
r184 28 32 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.825 $Y=1.665
+ $X2=1.68 $Y2=1.665
r185 27 39 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.935 $Y=1.665
+ $X2=4.08 $Y2=1.665
r186 27 28 2.61138 $w=1.4e-07 $l=2.11e-06 $layer=MET1_cond $X=3.935 $Y=1.665
+ $X2=1.825 $Y2=1.665
r187 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.475
+ $Y=1.41 $X2=5.475 $Y2=1.41
r188 22 37 12.0255 $w=2.28e-07 $l=2.4e-07 $layer=LI1_cond $X=5.04 $Y=1.425
+ $X2=5.04 $Y2=1.665
r189 22 24 12.2927 $w=2.98e-07 $l=3.2e-07 $layer=LI1_cond $X=5.155 $Y=1.425
+ $X2=5.475 $Y2=1.425
r190 19 25 52.2586 $w=2.99e-07 $l=2.57391e-07 $layer=POLY_cond $X=5.46 $Y=1.66
+ $X2=5.475 $Y2=1.41
r191 19 21 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=5.46 $Y=1.66
+ $X2=5.46 $Y2=2.235
r192 15 25 38.5562 $w=2.99e-07 $l=1.88348e-07 $layer=POLY_cond $X=5.425 $Y=1.245
+ $X2=5.475 $Y2=1.41
r193 15 17 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=5.425 $Y=1.245
+ $X2=5.425 $Y2=0.695
r194 12 45 52.2586 $w=2.99e-07 $l=2.69258e-07 $layer=POLY_cond $X=4.045 $Y=1.66
+ $X2=4.005 $Y2=1.41
r195 12 14 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=4.045 $Y=1.66
+ $X2=4.045 $Y2=2.235
r196 8 45 38.5562 $w=2.99e-07 $l=1.86145e-07 $layer=POLY_cond $X=3.96 $Y=1.245
+ $X2=4.005 $Y2=1.41
r197 8 10 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=3.96 $Y=1.245
+ $X2=3.96 $Y2=0.695
r198 5 42 52.2586 $w=2.99e-07 $l=2.82843e-07 $layer=POLY_cond $X=2.02 $Y=1.66
+ $X2=1.95 $Y2=1.41
r199 5 7 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=2.02 $Y=1.66
+ $X2=2.02 $Y2=2.235
r200 1 42 38.5562 $w=2.99e-07 $l=1.92678e-07 $layer=POLY_cond $X=1.89 $Y=1.245
+ $X2=1.95 $Y2=1.41
r201 1 3 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=1.89 $Y=1.245
+ $X2=1.89 $Y2=0.695
.ends

.subckt PM_SKY130_FD_SC_HS__FA_1%A_465_249# 1 2 9 11 13 14 16 19 21 22 23 26 27
+ 28 31 33 36 38 39 40 43 47 51
c183 47 0 1.02197e-19 $X=2.49 $Y=1.41
c184 38 0 1.47446e-19 $X=6.465 $Y=1.745
r185 58 60 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=6.235 $Y=1.065
+ $X2=6.465 $Y2=1.065
r186 51 53 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=5.21 $Y=0.6 $X2=5.21
+ $Y2=0.68
r187 47 48 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.49
+ $Y=1.41 $X2=2.49 $Y2=1.41
r188 43 44 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.875
+ $Y=1.385 $X2=7.875 $Y2=1.385
r189 41 43 8.20679 $w=3.28e-07 $l=2.35e-07 $layer=LI1_cond $X=7.875 $Y=1.15
+ $X2=7.875 $Y2=1.385
r190 40 60 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=6.55 $Y=1.065
+ $X2=6.465 $Y2=1.065
r191 39 41 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=7.71 $Y=1.065
+ $X2=7.875 $Y2=1.15
r192 39 40 75.6791 $w=1.68e-07 $l=1.16e-06 $layer=LI1_cond $X=7.71 $Y=1.065
+ $X2=6.55 $Y2=1.065
r193 37 60 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.465 $Y=1.15
+ $X2=6.465 $Y2=1.065
r194 37 38 38.8182 $w=1.68e-07 $l=5.95e-07 $layer=LI1_cond $X=6.465 $Y=1.15
+ $X2=6.465 $Y2=1.745
r195 36 58 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.235 $Y=0.98
+ $X2=6.235 $Y2=1.065
r196 35 36 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=6.235 $Y=0.765
+ $X2=6.235 $Y2=0.98
r197 33 38 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.38 $Y=1.83
+ $X2=6.465 $Y2=1.745
r198 33 34 57.738 $w=1.68e-07 $l=8.85e-07 $layer=LI1_cond $X=6.38 $Y=1.83
+ $X2=5.495 $Y2=1.83
r199 32 53 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.375 $Y=0.68
+ $X2=5.21 $Y2=0.68
r200 31 35 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.15 $Y=0.68
+ $X2=6.235 $Y2=0.765
r201 31 32 50.5615 $w=1.68e-07 $l=7.75e-07 $layer=LI1_cond $X=6.15 $Y=0.68
+ $X2=5.375 $Y2=0.68
r202 27 34 8.77544 $w=2.85e-07 $l=3.87161e-07 $layer=LI1_cond $X=5.197 $Y=2.035
+ $X2=5.495 $Y2=1.83
r203 27 28 122 $w=1.68e-07 $l=1.87e-06 $layer=LI1_cond $X=5.07 $Y=2.035 $X2=3.2
+ $Y2=2.035
r204 26 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.115 $Y=1.95
+ $X2=3.2 $Y2=2.035
r205 25 26 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=3.115 $Y=1.795
+ $X2=3.115 $Y2=1.95
r206 24 47 11.4375 $w=3.2e-07 $l=3.92301e-07 $layer=LI1_cond $X=2.75 $Y=1.71
+ $X2=2.537 $Y2=1.41
r207 23 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.03 $Y=1.71
+ $X2=3.115 $Y2=1.795
r208 23 24 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=3.03 $Y=1.71
+ $X2=2.75 $Y2=1.71
r209 21 44 31.475 $w=3.3e-07 $l=1.8e-07 $layer=POLY_cond $X=8.055 $Y=1.385
+ $X2=7.875 $Y2=1.385
r210 21 22 66.2869 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=8.145 $Y=1.385
+ $X2=8.145 $Y2=1.22
r211 19 22 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=8.16 $Y=0.74
+ $X2=8.16 $Y2=1.22
r212 14 21 149.859 $w=1.8e-07 $l=3.8e-07 $layer=POLY_cond $X=8.145 $Y=1.765
+ $X2=8.145 $Y2=1.385
r213 14 16 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=8.145 $Y=1.765
+ $X2=8.145 $Y2=2.4
r214 11 48 52.2586 $w=2.99e-07 $l=2.59808e-07 $layer=POLY_cond $X=2.47 $Y=1.66
+ $X2=2.49 $Y2=1.41
r215 11 13 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=2.47 $Y=1.66
+ $X2=2.47 $Y2=2.235
r216 7 48 38.5562 $w=2.99e-07 $l=1.92678e-07 $layer=POLY_cond $X=2.43 $Y=1.245
+ $X2=2.49 $Y2=1.41
r217 7 9 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=2.43 $Y=1.245
+ $X2=2.43 $Y2=0.695
r218 2 27 300 $w=1.7e-07 $l=3.67423e-07 $layer=licon1_PDIFF $count=2 $X=5.085
+ $Y=1.735 $X2=5.235 $Y2=2.035
r219 1 51 182 $w=1.7e-07 $l=2.86575e-07 $layer=licon1_NDIFF $count=1 $X=5.07
+ $Y=0.375 $X2=5.21 $Y2=0.6
.ends

.subckt PM_SKY130_FD_SC_HS__FA_1%B 3 5 8 9 10 13 14 15 16 17 18 21 22 26 27 28
+ 29 30 31 34 35 40 43 46 47 48 49 50 52 55 58
c175 58 0 1.00637e-19 $X=7.305 $Y=1.485
c176 40 0 3.65707e-20 $X=6.89 $Y=2.31
c177 28 0 9.44466e-20 $X=5.01 $Y=1.57
c178 21 0 2.62363e-19 $X=2.955 $Y=2.235
c179 5 0 8.44456e-20 $X=1.515 $Y=1.87
r180 57 58 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=7.305
+ $Y=1.485 $X2=7.305 $Y2=1.485
r181 55 57 13.0085 $w=3.52e-07 $l=9.5e-08 $layer=POLY_cond $X=7.21 $Y=1.527
+ $X2=7.305 $Y2=1.527
r182 54 55 43.8182 $w=3.52e-07 $l=3.2e-07 $layer=POLY_cond $X=6.89 $Y=1.527
+ $X2=7.21 $Y2=1.527
r183 52 58 3.21335 $w=6.68e-07 $l=1.8e-07 $layer=LI1_cond $X=7.135 $Y=1.665
+ $X2=7.135 $Y2=1.485
r184 41 55 22.7654 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=7.21 $Y=1.32
+ $X2=7.21 $Y2=1.527
r185 41 43 320.479 $w=1.5e-07 $l=6.25e-07 $layer=POLY_cond $X=7.21 $Y=1.32
+ $X2=7.21 $Y2=0.695
r186 38 50 105.158 $w=1.8e-07 $l=2.65e-07 $layer=POLY_cond $X=6.89 $Y=2.885
+ $X2=6.89 $Y2=3.15
r187 38 40 294.84 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=6.89 $Y=2.885
+ $X2=6.89 $Y2=2.31
r188 37 54 22.7654 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=6.89 $Y=1.735
+ $X2=6.89 $Y2=1.527
r189 37 40 294.84 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=6.89 $Y=1.735
+ $X2=6.89 $Y2=2.31
r190 36 49 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=5.1 $Y=3.15 $X2=5.01
+ $Y2=3.15
r191 35 50 7.1379 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=6.8 $Y=3.15 $X2=6.89
+ $Y2=3.15
r192 35 36 871.702 $w=1.5e-07 $l=1.7e-06 $layer=POLY_cond $X=6.8 $Y=3.15 $X2=5.1
+ $Y2=3.15
r193 32 34 294.84 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=5.01 $Y=2.81
+ $X2=5.01 $Y2=2.235
r194 31 34 294.84 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=5.01 $Y=1.66
+ $X2=5.01 $Y2=2.235
r195 30 49 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=5.01 $Y=3.075
+ $X2=5.01 $Y2=3.15
r196 29 32 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=5.01 $Y=2.9 $X2=5.01
+ $Y2=2.81
r197 29 30 68.0242 $w=1.8e-07 $l=1.75e-07 $layer=POLY_cond $X=5.01 $Y=2.9
+ $X2=5.01 $Y2=3.075
r198 28 31 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=5.01 $Y=1.57 $X2=5.01
+ $Y2=1.66
r199 27 48 37.1337 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=5.01 $Y=1.18 $X2=5.01
+ $Y2=1.09
r200 27 28 151.597 $w=1.8e-07 $l=3.9e-07 $layer=POLY_cond $X=5.01 $Y=1.18
+ $X2=5.01 $Y2=1.57
r201 26 48 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=4.995 $Y=0.695
+ $X2=4.995 $Y2=1.09
r202 23 47 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=3.045 $Y=3.15
+ $X2=2.955 $Y2=3.15
r203 22 49 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=4.92 $Y=3.15 $X2=5.01
+ $Y2=3.15
r204 22 23 961.436 $w=1.5e-07 $l=1.875e-06 $layer=POLY_cond $X=4.92 $Y=3.15
+ $X2=3.045 $Y2=3.15
r205 19 21 294.84 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=2.955 $Y=2.81
+ $X2=2.955 $Y2=2.235
r206 18 21 294.84 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=2.955 $Y=1.66
+ $X2=2.955 $Y2=2.235
r207 17 47 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=2.955 $Y=3.075
+ $X2=2.955 $Y2=3.15
r208 16 19 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=2.955 $Y=2.9
+ $X2=2.955 $Y2=2.81
r209 16 17 68.0242 $w=1.8e-07 $l=1.75e-07 $layer=POLY_cond $X=2.955 $Y=2.9
+ $X2=2.955 $Y2=3.075
r210 15 18 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=2.955 $Y=1.57
+ $X2=2.955 $Y2=1.66
r211 14 46 37.1337 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=2.955 $Y=1.18
+ $X2=2.955 $Y2=1.09
r212 14 15 151.597 $w=1.8e-07 $l=3.9e-07 $layer=POLY_cond $X=2.955 $Y=1.18
+ $X2=2.955 $Y2=1.57
r213 13 46 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=2.94 $Y=0.695
+ $X2=2.94 $Y2=1.09
r214 9 47 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=2.865 $Y=3.15
+ $X2=2.955 $Y2=3.15
r215 9 10 646.085 $w=1.5e-07 $l=1.26e-06 $layer=POLY_cond $X=2.865 $Y=3.15
+ $X2=1.605 $Y2=3.15
r216 6 10 26.9307 $w=1.5e-07 $l=1.69115e-07 $layer=POLY_cond $X=1.515 $Y=3.02
+ $X2=1.605 $Y2=3.15
r217 6 8 294.84 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=1.515 $Y=3.02
+ $X2=1.515 $Y2=2.445
r218 5 45 60.25 $w=1.8e-07 $l=1.55e-07 $layer=POLY_cond $X=1.515 $Y=1.87
+ $X2=1.515 $Y2=1.715
r219 5 8 294.84 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=1.515 $Y=1.87
+ $X2=1.515 $Y2=2.445
r220 3 45 523.021 $w=1.5e-07 $l=1.02e-06 $layer=POLY_cond $X=1.5 $Y=0.695
+ $X2=1.5 $Y2=1.715
.ends

.subckt PM_SKY130_FD_SC_HS__FA_1%SUM 1 2 9 11 15 16 17 28
r20 21 28 2.67531 $w=2.78e-07 $l=6.5e-08 $layer=LI1_cond $X=0.225 $Y=0.99
+ $X2=0.225 $Y2=0.925
r21 17 30 7.11633 $w=2.78e-07 $l=1.3e-07 $layer=LI1_cond $X=0.225 $Y=1 $X2=0.225
+ $Y2=1.13
r22 17 21 0.411587 $w=2.78e-07 $l=1e-08 $layer=LI1_cond $X=0.225 $Y=1 $X2=0.225
+ $Y2=0.99
r23 17 28 0.411587 $w=2.78e-07 $l=1e-08 $layer=LI1_cond $X=0.225 $Y=0.915
+ $X2=0.225 $Y2=0.925
r24 16 17 16.4635 $w=2.78e-07 $l=4e-07 $layer=LI1_cond $X=0.225 $Y=0.515
+ $X2=0.225 $Y2=0.915
r25 15 30 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=0.17 $Y=1.82 $X2=0.17
+ $Y2=1.13
r26 11 13 35.427 $w=2.68e-07 $l=8.3e-07 $layer=LI1_cond $X=0.22 $Y=1.985
+ $X2=0.22 $Y2=2.815
r27 9 15 7.33542 $w=2.68e-07 $l=1.35e-07 $layer=LI1_cond $X=0.22 $Y=1.955
+ $X2=0.22 $Y2=1.82
r28 9 11 1.28049 $w=2.68e-07 $l=3e-08 $layer=LI1_cond $X=0.22 $Y=1.955 $X2=0.22
+ $Y2=1.985
r29 2 13 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.27 $Y2=2.815
r30 2 11 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.27 $Y2=1.985
r31 1 16 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__FA_1%VPWR 1 2 3 4 5 18 24 28 32 36 41 42 43 45 50 59
+ 66 73 74 77 80 83 86
c108 4 0 1.10875e-19 $X=6.13 $Y=1.735
r109 86 87 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r110 83 84 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r111 80 81 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r112 77 78 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r113 74 87 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=3.33
+ $X2=7.92 $Y2=3.33
r114 73 74 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=3.33 $X2=8.4
+ $Y2=3.33
r115 71 86 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.085 $Y=3.33
+ $X2=7.92 $Y2=3.33
r116 71 73 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=8.085 $Y=3.33
+ $X2=8.4 $Y2=3.33
r117 70 87 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=7.92 $Y2=3.33
r118 70 84 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=6.48 $Y2=3.33
r119 69 70 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r120 67 83 13.7128 $w=1.7e-07 $l=3.53e-07 $layer=LI1_cond $X=6.825 $Y=3.33
+ $X2=6.472 $Y2=3.33
r121 67 69 40.123 $w=1.68e-07 $l=6.15e-07 $layer=LI1_cond $X=6.825 $Y=3.33
+ $X2=7.44 $Y2=3.33
r122 66 86 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.755 $Y=3.33
+ $X2=7.92 $Y2=3.33
r123 66 69 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=7.755 $Y=3.33
+ $X2=7.44 $Y2=3.33
r124 65 84 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=3.33 $X2=6.48
+ $Y2=3.33
r125 64 65 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r126 62 65 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=6 $Y2=3.33
r127 61 64 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=4.56 $Y=3.33 $X2=6
+ $Y2=3.33
r128 61 62 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r129 59 83 13.7128 $w=1.7e-07 $l=3.52e-07 $layer=LI1_cond $X=6.12 $Y=3.33
+ $X2=6.472 $Y2=3.33
r130 59 64 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=6.12 $Y=3.33 $X2=6
+ $Y2=3.33
r131 58 81 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=3.12 $Y2=3.33
r132 57 58 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r133 55 80 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.41 $Y=3.33
+ $X2=3.245 $Y2=3.33
r134 55 57 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.41 $Y=3.33
+ $X2=4.08 $Y2=3.33
r135 54 81 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=3.12 $Y2=3.33
r136 54 78 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r137 53 54 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r138 51 77 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.885 $Y=3.33
+ $X2=0.72 $Y2=3.33
r139 51 53 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=0.885 $Y=3.33
+ $X2=1.2 $Y2=3.33
r140 50 80 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.08 $Y=3.33
+ $X2=3.245 $Y2=3.33
r141 50 53 122.652 $w=1.68e-07 $l=1.88e-06 $layer=LI1_cond $X=3.08 $Y=3.33
+ $X2=1.2 $Y2=3.33
r142 48 78 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r143 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r144 45 77 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.555 $Y=3.33
+ $X2=0.72 $Y2=3.33
r145 45 47 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=0.555 $Y=3.33
+ $X2=0.24 $Y2=3.33
r146 43 62 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=4.32 $Y=3.33
+ $X2=4.56 $Y2=3.33
r147 43 58 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=4.32 $Y=3.33
+ $X2=4.08 $Y2=3.33
r148 41 57 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=4.105 $Y=3.33
+ $X2=4.08 $Y2=3.33
r149 41 42 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.105 $Y=3.33
+ $X2=4.27 $Y2=3.33
r150 40 61 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=4.435 $Y=3.33
+ $X2=4.56 $Y2=3.33
r151 40 42 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.435 $Y=3.33
+ $X2=4.27 $Y2=3.33
r152 36 39 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=7.92 $Y=1.985
+ $X2=7.92 $Y2=2.815
r153 34 86 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.92 $Y=3.245
+ $X2=7.92 $Y2=3.33
r154 34 39 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=7.92 $Y=3.245
+ $X2=7.92 $Y2=2.815
r155 30 83 2.87722 $w=7.05e-07 $l=8.5e-08 $layer=LI1_cond $X=6.472 $Y=3.245
+ $X2=6.472 $Y2=3.33
r156 30 32 10.9428 $w=7.03e-07 $l=6.45e-07 $layer=LI1_cond $X=6.472 $Y=3.245
+ $X2=6.472 $Y2=2.6
r157 26 42 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.27 $Y=3.245
+ $X2=4.27 $Y2=3.33
r158 26 28 27.0649 $w=3.28e-07 $l=7.75e-07 $layer=LI1_cond $X=4.27 $Y=3.245
+ $X2=4.27 $Y2=2.47
r159 22 80 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.245 $Y=3.245
+ $X2=3.245 $Y2=3.33
r160 22 24 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=3.245 $Y=3.245
+ $X2=3.245 $Y2=2.795
r161 18 21 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=0.72 $Y=2.135
+ $X2=0.72 $Y2=2.815
r162 16 77 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.72 $Y=3.245
+ $X2=0.72 $Y2=3.33
r163 16 21 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=0.72 $Y=3.245
+ $X2=0.72 $Y2=2.815
r164 5 39 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=7.775
+ $Y=1.84 $X2=7.92 $Y2=2.815
r165 5 36 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=7.775
+ $Y=1.84 $X2=7.92 $Y2=1.985
r166 4 32 300 $w=1.7e-07 $l=1.09849e-06 $layer=licon1_PDIFF $count=2 $X=6.13
+ $Y=1.735 $X2=6.66 $Y2=2.6
r167 3 28 600 $w=1.7e-07 $l=8.0652e-07 $layer=licon1_PDIFF $count=1 $X=4.12
+ $Y=1.735 $X2=4.27 $Y2=2.47
r168 2 24 600 $w=1.7e-07 $l=1.16254e-06 $layer=licon1_PDIFF $count=1 $X=3.03
+ $Y=1.735 $X2=3.245 $Y2=2.795
r169 1 21 600 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=0.57
+ $Y=1.84 $X2=0.72 $Y2=2.815
r170 1 18 300 $w=1.7e-07 $l=3.62319e-07 $layer=licon1_PDIFF $count=2 $X=0.57
+ $Y=1.84 $X2=0.72 $Y2=2.135
.ends

.subckt PM_SKY130_FD_SC_HS__FA_1%A_509_347# 1 2 9 13 15 17 18
c39 13 0 1.84258e-19 $X=2.695 $Y=2.59
r40 18 21 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=3.765 $Y=2.375
+ $X2=3.765 $Y2=2.455
r41 16 17 2.76166 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.86 $Y=2.375
+ $X2=2.735 $Y2=2.375
r42 15 18 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.6 $Y=2.375
+ $X2=3.765 $Y2=2.375
r43 15 16 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=3.6 $Y=2.375
+ $X2=2.86 $Y2=2.375
r44 11 17 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.735 $Y=2.46
+ $X2=2.735 $Y2=2.375
r45 11 13 5.9927 $w=2.48e-07 $l=1.3e-07 $layer=LI1_cond $X=2.735 $Y=2.46
+ $X2=2.735 $Y2=2.59
r46 7 17 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.735 $Y=2.29
+ $X2=2.735 $Y2=2.375
r47 7 9 7.37564 $w=2.48e-07 $l=1.6e-07 $layer=LI1_cond $X=2.735 $Y=2.29
+ $X2=2.735 $Y2=2.13
r48 2 21 600 $w=1.7e-07 $l=7.91454e-07 $layer=licon1_PDIFF $count=1 $X=3.615
+ $Y=1.735 $X2=3.765 $Y2=2.455
r49 1 13 600 $w=1.7e-07 $l=9.26971e-07 $layer=licon1_PDIFF $count=1 $X=2.545
+ $Y=1.735 $X2=2.695 $Y2=2.59
r50 1 9 600 $w=1.7e-07 $l=4.63977e-07 $layer=licon1_PDIFF $count=1 $X=2.545
+ $Y=1.735 $X2=2.695 $Y2=2.13
.ends

.subckt PM_SKY130_FD_SC_HS__FA_1%A_1107_347# 1 2 7 9 11 13 15
r28 13 20 3.10428 $w=3.2e-07 $l=1.5548e-07 $layer=LI1_cond $X=7.16 $Y=2.255
+ $X2=7.155 $Y2=2.102
r29 13 15 14.7657 $w=3.18e-07 $l=4.1e-07 $layer=LI1_cond $X=7.16 $Y=2.255
+ $X2=7.16 $Y2=2.665
r30 12 18 4.64039 $w=1.7e-07 $l=1.43e-07 $layer=LI1_cond $X=5.95 $Y=2.17
+ $X2=5.807 $Y2=2.17
r31 11 20 4.57783 $w=1.7e-07 $l=1.96074e-07 $layer=LI1_cond $X=6.99 $Y=2.17
+ $X2=7.155 $Y2=2.102
r32 11 12 67.8503 $w=1.68e-07 $l=1.04e-06 $layer=LI1_cond $X=6.99 $Y=2.17
+ $X2=5.95 $Y2=2.17
r33 7 18 2.75828 $w=2.85e-07 $l=8.5e-08 $layer=LI1_cond $X=5.807 $Y=2.255
+ $X2=5.807 $Y2=2.17
r34 7 9 13.5463 $w=2.83e-07 $l=3.35e-07 $layer=LI1_cond $X=5.807 $Y=2.255
+ $X2=5.807 $Y2=2.59
r35 2 20 600 $w=1.7e-07 $l=3.88555e-07 $layer=licon1_PDIFF $count=1 $X=6.965
+ $Y=1.81 $X2=7.155 $Y2=2.115
r36 2 15 600 $w=1.7e-07 $l=9.45238e-07 $layer=licon1_PDIFF $count=1 $X=6.965
+ $Y=1.81 $X2=7.155 $Y2=2.665
r37 1 18 600 $w=1.7e-07 $l=5.63516e-07 $layer=licon1_PDIFF $count=1 $X=5.535
+ $Y=1.735 $X2=5.83 $Y2=2.17
r38 1 9 600 $w=1.7e-07 $l=9.9159e-07 $layer=licon1_PDIFF $count=1 $X=5.535
+ $Y=1.735 $X2=5.83 $Y2=2.59
.ends

.subckt PM_SKY130_FD_SC_HS__FA_1%COUT 1 2 7 8 9 10 11 12 13 29
r18 22 29 1.3969 $w=3.28e-07 $l=4e-08 $layer=LI1_cond $X=8.375 $Y=0.965
+ $X2=8.375 $Y2=0.925
r19 12 13 16.7217 $w=2.53e-07 $l=3.7e-07 $layer=LI1_cond $X=8.412 $Y=2.405
+ $X2=8.412 $Y2=2.775
r20 11 12 18.9814 $w=2.53e-07 $l=4.2e-07 $layer=LI1_cond $X=8.412 $Y=1.985
+ $X2=8.412 $Y2=2.405
r21 10 11 14.462 $w=2.53e-07 $l=3.2e-07 $layer=LI1_cond $X=8.412 $Y=1.665
+ $X2=8.412 $Y2=1.985
r22 9 10 16.7217 $w=2.53e-07 $l=3.7e-07 $layer=LI1_cond $X=8.412 $Y=1.295
+ $X2=8.412 $Y2=1.665
r23 9 45 7.45698 $w=2.53e-07 $l=1.65e-07 $layer=LI1_cond $X=8.412 $Y=1.295
+ $X2=8.412 $Y2=1.13
r24 8 45 5.6192 $w=3.28e-07 $l=1.43e-07 $layer=LI1_cond $X=8.375 $Y=0.987
+ $X2=8.375 $Y2=1.13
r25 8 22 0.768295 $w=3.28e-07 $l=2.2e-08 $layer=LI1_cond $X=8.375 $Y=0.987
+ $X2=8.375 $Y2=0.965
r26 8 29 0.803218 $w=3.28e-07 $l=2.3e-08 $layer=LI1_cond $X=8.375 $Y=0.902
+ $X2=8.375 $Y2=0.925
r27 7 8 13.515 $w=3.28e-07 $l=3.87e-07 $layer=LI1_cond $X=8.375 $Y=0.515
+ $X2=8.375 $Y2=0.902
r28 2 13 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=8.22
+ $Y=1.84 $X2=8.37 $Y2=2.815
r29 2 11 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=8.22
+ $Y=1.84 $X2=8.37 $Y2=1.985
r30 1 7 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=8.235
+ $Y=0.37 $X2=8.375 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__FA_1%VGND 1 2 3 4 5 16 20 24 28 30 32 37 42 50 57 58
+ 69 75 78 81
r108 81 82 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=0 $X2=7.92
+ $Y2=0
r109 78 79 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=0 $X2=6.96
+ $Y2=0
r110 75 76 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r111 70 76 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=4.08
+ $Y2=0
r112 69 72 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=3.235 $Y=0
+ $X2=3.235 $Y2=0.325
r113 69 70 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.12 $Y=0
+ $X2=3.12 $Y2=0
r114 58 82 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=0 $X2=7.92
+ $Y2=0
r115 57 58 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r116 55 81 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.03 $Y=0 $X2=7.905
+ $Y2=0
r117 55 57 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=8.03 $Y=0 $X2=8.4
+ $Y2=0
r118 54 82 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=0 $X2=7.92
+ $Y2=0
r119 54 79 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=0 $X2=6.96
+ $Y2=0
r120 53 54 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=0 $X2=7.44
+ $Y2=0
r121 51 78 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.08 $Y=0 $X2=6.955
+ $Y2=0
r122 51 53 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=7.08 $Y=0 $X2=7.44
+ $Y2=0
r123 50 81 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.78 $Y=0 $X2=7.905
+ $Y2=0
r124 50 53 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=7.78 $Y=0 $X2=7.44
+ $Y2=0
r125 49 79 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=0 $X2=6.96
+ $Y2=0
r126 48 49 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6.48 $Y=0
+ $X2=6.48 $Y2=0
r127 46 49 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=4.56 $Y=0
+ $X2=6.48 $Y2=0
r128 45 48 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=4.56 $Y=0 $X2=6.48
+ $Y2=0
r129 45 46 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.56 $Y=0
+ $X2=4.56 $Y2=0
r130 43 75 10.9443 $w=1.7e-07 $l=2.38e-07 $layer=LI1_cond $X=4.555 $Y=0
+ $X2=4.317 $Y2=0
r131 43 45 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=4.555 $Y=0 $X2=4.56
+ $Y2=0
r132 42 78 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.83 $Y=0 $X2=6.955
+ $Y2=0
r133 42 48 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=6.83 $Y=0 $X2=6.48
+ $Y2=0
r134 41 70 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=1.2 $Y=0 $X2=3.12
+ $Y2=0
r135 41 63 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r136 40 41 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r137 38 40 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=0.98 $Y=0 $X2=1.2
+ $Y2=0
r138 37 69 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.07 $Y=0 $X2=3.235
+ $Y2=0
r139 37 40 122 $w=1.68e-07 $l=1.87e-06 $layer=LI1_cond $X=3.07 $Y=0 $X2=1.2
+ $Y2=0
r140 35 63 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r141 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r142 32 65 10.5505 $w=3.53e-07 $l=3.25e-07 $layer=LI1_cond $X=0.802 $Y=0
+ $X2=0.802 $Y2=0.325
r143 32 38 5.0588 $w=1.7e-07 $l=1.78e-07 $layer=LI1_cond $X=0.802 $Y=0 $X2=0.98
+ $Y2=0
r144 32 63 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r145 32 34 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=0.625 $Y=0
+ $X2=0.24 $Y2=0
r146 30 46 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=4.32 $Y=0
+ $X2=4.56 $Y2=0
r147 30 76 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=4.32 $Y=0
+ $X2=4.08 $Y2=0
r148 26 81 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=7.905 $Y=0.085
+ $X2=7.905 $Y2=0
r149 26 28 23.9708 $w=2.48e-07 $l=5.2e-07 $layer=LI1_cond $X=7.905 $Y=0.085
+ $X2=7.905 $Y2=0.605
r150 22 78 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.955 $Y=0.085
+ $X2=6.955 $Y2=0
r151 22 24 10.1415 $w=2.48e-07 $l=2.2e-07 $layer=LI1_cond $X=6.955 $Y=0.085
+ $X2=6.955 $Y2=0.305
r152 18 75 1.94084 $w=4.75e-07 $l=8.5e-08 $layer=LI1_cond $X=4.317 $Y=0.085
+ $X2=4.317 $Y2=0
r153 18 20 11.5831 $w=4.73e-07 $l=4.6e-07 $layer=LI1_cond $X=4.317 $Y=0.085
+ $X2=4.317 $Y2=0.545
r154 17 69 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.4 $Y=0 $X2=3.235
+ $Y2=0
r155 16 75 10.9443 $w=1.7e-07 $l=2.37e-07 $layer=LI1_cond $X=4.08 $Y=0 $X2=4.317
+ $Y2=0
r156 16 17 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=4.08 $Y=0 $X2=3.4
+ $Y2=0
r157 5 28 182 $w=1.7e-07 $l=2.90861e-07 $layer=licon1_NDIFF $count=1 $X=7.82
+ $Y=0.37 $X2=7.945 $Y2=0.605
r158 4 24 182 $w=1.7e-07 $l=3.88426e-07 $layer=licon1_NDIFF $count=1 $X=6.56
+ $Y=0.375 $X2=6.915 $Y2=0.305
r159 3 20 182 $w=1.7e-07 $l=3.54965e-07 $layer=licon1_NDIFF $count=1 $X=4.035
+ $Y=0.375 $X2=4.315 $Y2=0.545
r160 2 72 182 $w=1.7e-07 $l=2.43721e-07 $layer=licon1_NDIFF $count=1 $X=3.015
+ $Y=0.375 $X2=3.235 $Y2=0.325
r161 1 65 182 $w=1.7e-07 $l=2.51496e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.37 $X2=0.8 $Y2=0.325
.ends

.subckt PM_SKY130_FD_SC_HS__FA_1%A_501_75# 1 2 7 12 14
c26 12 0 8.59909e-20 $X=2.89 $Y=0.585
r27 14 16 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=3.745 $Y=0.585
+ $X2=3.745 $Y2=0.665
r28 10 12 9.85908 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=2.685 $Y=0.585
+ $X2=2.89 $Y2=0.585
r29 7 16 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.58 $Y=0.665
+ $X2=3.745 $Y2=0.665
r30 7 12 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=3.58 $Y=0.665 $X2=2.89
+ $Y2=0.665
r31 2 14 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=3.605
+ $Y=0.375 $X2=3.745 $Y2=0.585
r32 1 10 182 $w=1.7e-07 $l=2.86182e-07 $layer=licon1_NDIFF $count=1 $X=2.505
+ $Y=0.375 $X2=2.685 $Y2=0.585
.ends

.subckt PM_SKY130_FD_SC_HS__FA_1%A_1100_75# 1 2 7 12 13 14 16
r41 16 18 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=7.425 $Y=0.645
+ $X2=7.425 $Y2=0.725
r42 13 18 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.26 $Y=0.725
+ $X2=7.425 $Y2=0.725
r43 13 14 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=7.26 $Y=0.725 $X2=6.66
+ $Y2=0.725
r44 12 14 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.575 $Y=0.64
+ $X2=6.66 $Y2=0.725
r45 11 12 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=6.575 $Y=0.425
+ $X2=6.575 $Y2=0.64
r46 7 11 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.49 $Y=0.34
+ $X2=6.575 $Y2=0.425
r47 7 9 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=6.49 $Y=0.34 $X2=6.19
+ $Y2=0.34
r48 2 16 182 $w=1.7e-07 $l=3.32716e-07 $layer=licon1_NDIFF $count=1 $X=7.285
+ $Y=0.375 $X2=7.425 $Y2=0.645
r49 1 9 91 $w=1.7e-07 $l=7.07284e-07 $layer=licon1_NDIFF $count=2 $X=5.5
+ $Y=0.375 $X2=6.19 $Y2=0.34
.ends

