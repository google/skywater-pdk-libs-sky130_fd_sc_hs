# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_sc_hs__buf_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__buf_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  2.400000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.825000 1.350000 2.275000 1.780000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  0.543200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.945000 0.350000 1.275000 1.180000 ;
        RECT 0.945000 1.180000 1.315000 2.150000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 2.400000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.000000 0.000000 2.400000 0.245000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.660000 2.590000 3.520000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 2.400000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.400000 0.085000 ;
      RECT 0.000000  3.245000 2.400000 3.415000 ;
      RECT 0.105000  1.300000 0.775000 1.630000 ;
      RECT 0.115000  1.820000 0.420000 2.735000 ;
      RECT 0.115000  2.735000 0.825000 3.245000 ;
      RECT 0.515000  0.085000 0.765000 1.130000 ;
      RECT 0.605000  1.630000 0.775000 2.320000 ;
      RECT 0.605000  2.320000 2.285000 2.490000 ;
      RECT 1.395000  2.660000 1.725000 3.245000 ;
      RECT 1.445000  0.085000 1.775000 0.840000 ;
      RECT 1.485000  1.010000 2.285000 1.180000 ;
      RECT 1.485000  1.180000 1.655000 2.320000 ;
      RECT 1.930000  1.950000 2.285000 2.320000 ;
      RECT 1.930000  2.490000 2.285000 2.880000 ;
      RECT 1.955000  0.450000 2.285000 1.010000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
  END
END sky130_fd_sc_hs__buf_2
END LIBRARY
