* File: sky130_fd_sc_hs__o22a_4.spice
* Created: Tue Sep  1 20:16:16 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hs__o22a_4.pex.spice"
.subckt sky130_fd_sc_hs__o22a_4  VNB VPB A2 A1 B2 B1 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* B1	B1
* B2	B2
* A1	A1
* A2	A2
* VPB	VPB
* VNB	VNB
MM1020 N_A_27_136#_M1020_d N_A1_M1020_g N_VGND_M1020_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.1824 AS=0.112 PD=1.85 PS=0.99 NRD=0 NRS=13.116 M=1 R=4.26667 SA=75000.2
+ SB=75003.6 A=0.096 P=1.58 MULT=1
MM1018 N_A_27_136#_M1018_d N_A2_M1018_g N_VGND_M1020_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.0896 AS=0.112 PD=0.92 PS=0.99 NRD=0 NRS=0 M=1 R=4.26667 SA=75000.7
+ SB=75003.1 A=0.096 P=1.58 MULT=1
MM1019 N_A_27_136#_M1018_d N_A2_M1019_g N_VGND_M1019_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.0896 AS=0.1248 PD=0.92 PS=1.03 NRD=0 NRS=13.116 M=1 R=4.26667 SA=75001.1
+ SB=75002.6 A=0.096 P=1.58 MULT=1
MM1021 N_A_27_136#_M1021_d N_A1_M1021_g N_VGND_M1019_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.12 AS=0.1248 PD=1.015 PS=1.03 NRD=5.616 NRS=7.488 M=1 R=4.26667
+ SA=75001.7 SB=75002.1 A=0.096 P=1.58 MULT=1
MM1001 N_A_27_136#_M1021_d N_B1_M1001_g N_A_206_392#_M1001_s VNB NLOWVT L=0.15
+ W=0.64 AD=0.12 AS=0.0912 PD=1.015 PS=0.925 NRD=12.18 NRS=0.936 M=1 R=4.26667
+ SA=75002.2 SB=75001.6 A=0.096 P=1.58 MULT=1
MM1013 N_A_206_392#_M1001_s N_B2_M1013_g N_A_27_136#_M1013_s VNB NLOWVT L=0.15
+ W=0.64 AD=0.0912 AS=0.1136 PD=0.925 PS=0.995 NRD=0 NRS=6.552 M=1 R=4.26667
+ SA=75002.6 SB=75001.1 A=0.096 P=1.58 MULT=1
MM1017 N_A_206_392#_M1017_d N_B2_M1017_g N_A_27_136#_M1013_s VNB NLOWVT L=0.15
+ W=0.64 AD=0.0896 AS=0.1136 PD=0.92 PS=0.995 NRD=0 NRS=7.488 M=1 R=4.26667
+ SA=75003.1 SB=75000.6 A=0.096 P=1.58 MULT=1
MM1023 N_A_27_136#_M1023_d N_B1_M1023_g N_A_206_392#_M1017_d VNB NLOWVT L=0.15
+ W=0.64 AD=0.1824 AS=0.0896 PD=1.85 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75003.6 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1004 N_VGND_M1004_d N_A_206_392#_M1004_g N_X_M1004_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.2991 AS=0.1036 PD=2.41 PS=1.02 NRD=13.776 NRS=0 M=1 R=4.93333 SA=75000.3
+ SB=75001.5 A=0.111 P=1.78 MULT=1
MM1007 N_VGND_M1007_d N_A_206_392#_M1007_g N_X_M1004_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.7
+ SB=75001.1 A=0.111 P=1.78 MULT=1
MM1016 N_VGND_M1007_d N_A_206_392#_M1016_g N_X_M1016_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.1
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1022 N_VGND_M1022_d N_A_206_392#_M1022_g N_X_M1016_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.2146 AS=0.1036 PD=2.06 PS=1.02 NRD=0.804 NRS=0 M=1 R=4.93333 SA=75001.6
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1008 N_VPWR_M1008_d N_A1_M1008_g N_A_116_392#_M1008_s VPB PSHORT L=0.15 W=1
+ AD=0.295 AS=0.15 PD=2.59 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=6.66667 SA=75000.2
+ SB=75005.9 A=0.15 P=2.3 MULT=1
MM1010 N_A_206_392#_M1010_d N_A2_M1010_g N_A_116_392#_M1008_s VPB PSHORT L=0.15
+ W=1 AD=0.175 AS=0.15 PD=1.35 PS=1.3 NRD=11.8003 NRS=1.9503 M=1 R=6.66667
+ SA=75000.7 SB=75005.5 A=0.15 P=2.3 MULT=1
MM1011 N_A_206_392#_M1010_d N_A2_M1011_g N_A_116_392#_M1011_s VPB PSHORT L=0.15
+ W=1 AD=0.175 AS=0.175 PD=1.35 PS=1.35 NRD=1.9503 NRS=11.8003 M=1 R=6.66667
+ SA=75001.2 SB=75005 A=0.15 P=2.3 MULT=1
MM1009 N_VPWR_M1009_d N_A1_M1009_g N_A_116_392#_M1011_s VPB PSHORT L=0.15 W=1
+ AD=0.2 AS=0.175 PD=1.4 PS=1.35 NRD=11.8003 NRS=1.9503 M=1 R=6.66667 SA=75001.7
+ SB=75004.5 A=0.15 P=2.3 MULT=1
MM1002 N_A_516_392#_M1002_d N_B1_M1002_g N_VPWR_M1009_d VPB PSHORT L=0.15 W=1
+ AD=0.15 AS=0.2 PD=1.3 PS=1.4 NRD=1.9503 NRS=11.8003 M=1 R=6.66667 SA=75002.2
+ SB=75003.9 A=0.15 P=2.3 MULT=1
MM1005 N_A_206_392#_M1005_d N_B2_M1005_g N_A_516_392#_M1002_d VPB PSHORT L=0.15
+ W=1 AD=0.175 AS=0.15 PD=1.35 PS=1.3 NRD=11.8003 NRS=1.9503 M=1 R=6.66667
+ SA=75002.7 SB=75003.5 A=0.15 P=2.3 MULT=1
MM1006 N_A_206_392#_M1005_d N_B2_M1006_g N_A_516_392#_M1006_s VPB PSHORT L=0.15
+ W=1 AD=0.175 AS=0.175 PD=1.35 PS=1.35 NRD=1.9503 NRS=11.8003 M=1 R=6.66667
+ SA=75003.2 SB=75003 A=0.15 P=2.3 MULT=1
MM1003 N_A_516_392#_M1006_s N_B1_M1003_g N_VPWR_M1003_s VPB PSHORT L=0.15 W=1
+ AD=0.175 AS=0.206226 PD=1.35 PS=1.43396 NRD=1.9503 NRS=19.0302 M=1 R=6.66667
+ SA=75003.7 SB=75002.5 A=0.15 P=2.3 MULT=1
MM1000 N_VPWR_M1003_s N_A_206_392#_M1000_g N_X_M1000_s VPB PSHORT L=0.15 W=1.12
+ AD=0.230974 AS=0.1876 PD=1.60604 PS=1.455 NRD=4.3931 NRS=7.8997 M=1 R=7.46667
+ SA=75003.8 SB=75001.9 A=0.168 P=2.54 MULT=1
MM1012 N_VPWR_M1012_d N_A_206_392#_M1012_g N_X_M1000_s VPB PSHORT L=0.15 W=1.12
+ AD=0.322 AS=0.1876 PD=1.695 PS=1.455 NRD=28.1316 NRS=1.7533 M=1 R=7.46667
+ SA=75004.3 SB=75001.4 A=0.168 P=2.54 MULT=1
MM1014 N_VPWR_M1012_d N_A_206_392#_M1014_g N_X_M1014_s VPB PSHORT L=0.15 W=1.12
+ AD=0.322 AS=0.168 PD=1.695 PS=1.42 NRD=23.7385 NRS=1.7533 M=1 R=7.46667
+ SA=75005 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1015 N_VPWR_M1015_d N_A_206_392#_M1015_g N_X_M1014_s VPB PSHORT L=0.15 W=1.12
+ AD=0.3864 AS=0.168 PD=2.93 PS=1.42 NRD=10.5395 NRS=1.7533 M=1 R=7.46667
+ SA=75005.5 SB=75000.3 A=0.168 P=2.54 MULT=1
DX24_noxref VNB VPB NWDIODE A=13.206 P=17.92
c_114 VPB 0 1.20589e-19 $X=0 $Y=3.085
*
.include "sky130_fd_sc_hs__o22a_4.pxi.spice"
*
.ends
*
*
