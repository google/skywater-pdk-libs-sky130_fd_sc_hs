* File: sky130_fd_sc_hs__a32oi_4.spice
* Created: Thu Aug 27 20:30:33 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hs__a32oi_4.pex.spice"
.subckt sky130_fd_sc_hs__a32oi_4  VNB VPB B2 B1 A1 A2 A3 Y VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* Y	Y
* A3	A3
* A2	A2
* A1	A1
* B1	B1
* B2	B2
* VPB	VPB
* VNB	VNB
MM1004 N_A_27_74#_M1004_d N_B2_M1004_g N_VGND_M1004_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.1295 PD=2.05 PS=1.09 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75000.2
+ SB=75003.4 A=0.111 P=1.78 MULT=1
MM1006 N_A_27_74#_M1006_d N_B2_M1006_g N_VGND_M1004_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1295 PD=1.02 PS=1.09 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.7
+ SB=75002.9 A=0.111 P=1.78 MULT=1
MM1025 N_A_27_74#_M1006_d N_B2_M1025_g N_VGND_M1025_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.12765 PD=1.02 PS=1.085 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.1
+ SB=75002.5 A=0.111 P=1.78 MULT=1
MM1034 N_A_27_74#_M1034_d N_B2_M1034_g N_VGND_M1025_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.12765 PD=1.02 PS=1.085 NRD=0 NRS=10.536 M=1 R=4.93333
+ SA=75001.6 SB=75002 A=0.111 P=1.78 MULT=1
MM1009 N_A_27_74#_M1034_d N_B1_M1009_g N_Y_M1009_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75002.1
+ SB=75001.6 A=0.111 P=1.78 MULT=1
MM1018 N_A_27_74#_M1018_d N_B1_M1018_g N_Y_M1009_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1295 AS=0.1036 PD=1.09 PS=1.02 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75002.5
+ SB=75001.1 A=0.111 P=1.78 MULT=1
MM1031 N_A_27_74#_M1018_d N_B1_M1031_g N_Y_M1031_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1295 AS=0.1036 PD=1.09 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75003
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1037 N_A_27_74#_M1037_d N_B1_M1037_g N_Y_M1031_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.1036 PD=2.05 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75003.4
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1002 N_A_868_74#_M1002_d N_A1_M1002_g N_Y_M1002_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.1295 PD=2.05 PS=1.09 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75000.2
+ SB=75003.3 A=0.111 P=1.78 MULT=1
MM1019 N_A_868_74#_M1019_d N_A1_M1019_g N_Y_M1002_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1295 PD=1.02 PS=1.09 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.7
+ SB=75002.8 A=0.111 P=1.78 MULT=1
MM1032 N_A_868_74#_M1019_d N_A1_M1032_g N_Y_M1032_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.1
+ SB=75002.4 A=0.111 P=1.78 MULT=1
MM1035 N_A_868_74#_M1035_d N_A1_M1035_g N_Y_M1032_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.6
+ SB=75001.9 A=0.111 P=1.78 MULT=1
MM1000 N_A_868_74#_M1035_d N_A2_M1000_g N_A_1313_74#_M1000_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75002
+ SB=75001.5 A=0.111 P=1.78 MULT=1
MM1003 N_A_868_74#_M1003_d N_A2_M1003_g N_A_1313_74#_M1000_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.10545 AS=0.1036 PD=1.025 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75002.4 SB=75001.1 A=0.111 P=1.78 MULT=1
MM1012 N_A_868_74#_M1003_d N_A2_M1012_g N_A_1313_74#_M1012_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.10545 AS=0.1036 PD=1.025 PS=1.02 NRD=0.804 NRS=0 M=1 R=4.93333
+ SA=75002.9 SB=75000.6 A=0.111 P=1.78 MULT=1
MM1013 N_A_868_74#_M1013_d N_A2_M1013_g N_A_1313_74#_M1012_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.2109 AS=0.1036 PD=2.05 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75003.3 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1001 N_VGND_M1001_d N_A3_M1001_g N_A_1313_74#_M1001_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.1036 PD=2.05 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75001.5 A=0.111 P=1.78 MULT=1
MM1014 N_VGND_M1014_d N_A3_M1014_g N_A_1313_74#_M1001_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.6
+ SB=75001.1 A=0.111 P=1.78 MULT=1
MM1036 N_VGND_M1014_d N_A3_M1036_g N_A_1313_74#_M1036_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.1
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1038 N_VGND_M1038_d N_A3_M1038_g N_A_1313_74#_M1036_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.1036 PD=2.05 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.5
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1005 N_Y_M1005_d N_B2_M1005_g N_A_27_368#_M1005_s VPB PSHORT L=0.15 W=1.12
+ AD=0.1932 AS=0.336 PD=1.465 PS=2.84 NRD=9.6727 NRS=2.6201 M=1 R=7.46667
+ SA=75000.2 SB=75009.8 A=0.168 P=2.54 MULT=1
MM1010 N_Y_M1005_d N_B2_M1010_g N_A_27_368#_M1010_s VPB PSHORT L=0.15 W=1.12
+ AD=0.1932 AS=0.168 PD=1.465 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.7 SB=75009.3 A=0.168 P=2.54 MULT=1
MM1015 N_Y_M1015_d N_B2_M1015_g N_A_27_368#_M1010_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.2 SB=75008.8 A=0.168 P=2.54 MULT=1
MM1021 N_Y_M1015_d N_B2_M1021_g N_A_27_368#_M1021_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.196 PD=1.42 PS=1.47 NRD=1.7533 NRS=10.5395 M=1 R=7.46667
+ SA=75001.6 SB=75008.4 A=0.168 P=2.54 MULT=1
MM1011 N_A_27_368#_M1021_s N_B1_M1011_g N_Y_M1011_s VPB PSHORT L=0.15 W=1.12
+ AD=0.196 AS=0.196 PD=1.47 PS=1.47 NRD=1.7533 NRS=10.5395 M=1 R=7.46667
+ SA=75002.1 SB=75007.9 A=0.168 P=2.54 MULT=1
MM1016 N_A_27_368#_M1016_d N_B1_M1016_g N_Y_M1011_s VPB PSHORT L=0.15 W=1.12
+ AD=0.196 AS=0.196 PD=1.47 PS=1.47 NRD=10.5395 NRS=1.7533 M=1 R=7.46667
+ SA=75002.6 SB=75007.4 A=0.168 P=2.54 MULT=1
MM1017 N_A_27_368#_M1016_d N_B1_M1017_g N_Y_M1017_s VPB PSHORT L=0.15 W=1.12
+ AD=0.196 AS=0.196 PD=1.47 PS=1.47 NRD=1.7533 NRS=10.5395 M=1 R=7.46667
+ SA=75003.1 SB=75006.9 A=0.168 P=2.54 MULT=1
MM1020 N_A_27_368#_M1020_d N_B1_M1020_g N_Y_M1017_s VPB PSHORT L=0.15 W=1.12
+ AD=0.2744 AS=0.196 PD=1.61 PS=1.47 NRD=10.5395 NRS=1.7533 M=1 R=7.46667
+ SA=75003.6 SB=75006.4 A=0.168 P=2.54 MULT=1
MM1022 N_A_27_368#_M1020_d N_A1_M1022_g N_VPWR_M1022_s VPB PSHORT L=0.15 W=1.12
+ AD=0.2744 AS=0.196 PD=1.61 PS=1.47 NRD=26.3783 NRS=1.7533 M=1 R=7.46667
+ SA=75004.3 SB=75005.7 A=0.168 P=2.54 MULT=1
MM1023 N_A_27_368#_M1023_d N_A1_M1023_g N_VPWR_M1022_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.196 PD=1.42 PS=1.47 NRD=1.7533 NRS=10.5395 M=1 R=7.46667
+ SA=75004.8 SB=75005.2 A=0.168 P=2.54 MULT=1
MM1029 N_A_27_368#_M1023_d N_A1_M1029_g N_VPWR_M1029_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.224 PD=1.42 PS=1.52 NRD=1.7533 NRS=10.5395 M=1 R=7.46667
+ SA=75005.2 SB=75004.8 A=0.168 P=2.54 MULT=1
MM1039 N_A_27_368#_M1039_d N_A1_M1039_g N_VPWR_M1029_s VPB PSHORT L=0.15 W=1.12
+ AD=0.1736 AS=0.224 PD=1.43 PS=1.52 NRD=1.7533 NRS=10.5395 M=1 R=7.46667
+ SA=75005.8 SB=75004.2 A=0.168 P=2.54 MULT=1
MM1007 N_VPWR_M1007_d N_A2_M1007_g N_A_27_368#_M1039_d VPB PSHORT L=0.15 W=1.12
+ AD=0.2184 AS=0.1736 PD=1.51 PS=1.43 NRD=8.7862 NRS=3.5066 M=1 R=7.46667
+ SA=75006.2 SB=75003.8 A=0.168 P=2.54 MULT=1
MM1026 N_VPWR_M1007_d N_A2_M1026_g N_A_27_368#_M1026_s VPB PSHORT L=0.15 W=1.12
+ AD=0.2184 AS=0.168 PD=1.51 PS=1.42 NRD=10.5395 NRS=1.7533 M=1 R=7.46667
+ SA=75006.8 SB=75003.2 A=0.168 P=2.54 MULT=1
MM1030 N_VPWR_M1030_d N_A2_M1030_g N_A_27_368#_M1026_s VPB PSHORT L=0.15 W=1.12
+ AD=0.196 AS=0.168 PD=1.47 PS=1.42 NRD=10.5395 NRS=1.7533 M=1 R=7.46667
+ SA=75007.2 SB=75002.8 A=0.168 P=2.54 MULT=1
MM1033 N_VPWR_M1030_d N_A2_M1033_g N_A_27_368#_M1033_s VPB PSHORT L=0.15 W=1.12
+ AD=0.196 AS=0.196 PD=1.47 PS=1.47 NRD=1.7533 NRS=10.5395 M=1 R=7.46667
+ SA=75007.7 SB=75002.3 A=0.168 P=2.54 MULT=1
MM1008 N_A_27_368#_M1033_s N_A3_M1008_g N_VPWR_M1008_s VPB PSHORT L=0.15 W=1.12
+ AD=0.196 AS=0.196 PD=1.47 PS=1.47 NRD=1.7533 NRS=10.5395 M=1 R=7.46667
+ SA=75008.2 SB=75001.8 A=0.168 P=2.54 MULT=1
MM1024 N_A_27_368#_M1024_d N_A3_M1024_g N_VPWR_M1008_s VPB PSHORT L=0.15 W=1.12
+ AD=0.196 AS=0.196 PD=1.47 PS=1.47 NRD=10.5395 NRS=1.7533 M=1 R=7.46667
+ SA=75008.7 SB=75001.3 A=0.168 P=2.54 MULT=1
MM1027 N_A_27_368#_M1024_d N_A3_M1027_g N_VPWR_M1027_s VPB PSHORT L=0.15 W=1.12
+ AD=0.196 AS=0.2268 PD=1.47 PS=1.525 NRD=1.7533 NRS=10.5395 M=1 R=7.46667
+ SA=75009.2 SB=75000.8 A=0.168 P=2.54 MULT=1
MM1028 N_A_27_368#_M1028_d N_A3_M1028_g N_VPWR_M1027_s VPB PSHORT L=0.15 W=1.12
+ AD=0.3304 AS=0.2268 PD=2.83 PS=1.525 NRD=1.7533 NRS=11.426 M=1 R=7.46667
+ SA=75009.8 SB=75000.2 A=0.168 P=2.54 MULT=1
DX40_noxref VNB VPB NWDIODE A=20.3484 P=25.6
*
.include "sky130_fd_sc_hs__a32oi_4.pxi.spice"
*
.ends
*
*
