* File: sky130_fd_sc_hs__or2_1.spice
* Created: Tue Sep  1 20:19:48 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hs__or2_1.pex.spice"
.subckt sky130_fd_sc_hs__or2_1  VNB VPB B A VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A	A
* B	B
* VPB	VPB
* VNB	VNB
MM1005 N_A_63_368#_M1005_d N_B_M1005_g N_VGND_M1005_s VNB NLOWVT L=0.15 W=0.55
+ AD=0.130625 AS=0.2695 PD=1.025 PS=2.08 NRD=34.908 NRS=0 M=1 R=3.66667
+ SA=75000.4 SB=75001.4 A=0.0825 P=1.4 MULT=1
MM1004 N_VGND_M1004_d N_A_M1004_g N_A_63_368#_M1005_d VNB NLOWVT L=0.15 W=0.55
+ AD=0.129591 AS=0.130625 PD=0.997674 PS=1.025 NRD=17.448 NRS=7.632 M=1
+ R=3.66667 SA=75001 SB=75000.8 A=0.0825 P=1.4 MULT=1
MM1002 N_X_M1002_d N_A_63_368#_M1002_g N_VGND_M1004_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.174359 PD=2.05 PS=1.34233 NRD=0 NRS=11.34 M=1 R=4.93333
+ SA=75001.3 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1000 A_152_368# N_B_M1000_g N_A_63_368#_M1000_s VPB PSHORT L=0.15 W=0.84
+ AD=0.1134 AS=0.2478 PD=1.11 PS=2.27 NRD=18.7544 NRS=2.3443 M=1 R=5.6
+ SA=75000.2 SB=75001.4 A=0.126 P=1.98 MULT=1
MM1003 N_VPWR_M1003_d N_A_M1003_g A_152_368# VPB PSHORT L=0.15 W=0.84 AD=0.2868
+ AS=0.1134 PD=1.50857 PS=1.11 NRD=67.1573 NRS=18.7544 M=1 R=5.6 SA=75000.6
+ SB=75001 A=0.126 P=1.98 MULT=1
MM1001 N_X_M1001_d N_A_63_368#_M1001_g N_VPWR_M1003_d VPB PSHORT L=0.15 W=1.12
+ AD=0.3304 AS=0.3824 PD=2.83 PS=2.01143 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.2 SB=75000.2 A=0.168 P=2.54 MULT=1
DX6_noxref VNB VPB NWDIODE A=5.1708 P=9.28
*
.include "sky130_fd_sc_hs__or2_1.pxi.spice"
*
.ends
*
*
