* File: sky130_fd_sc_hs__and4bb_2.spice
* Created: Thu Aug 27 20:33:57 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hs__and4bb_2.pex.spice"
.subckt sky130_fd_sc_hs__and4bb_2  VNB VPB A_N C D B_N VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* B_N	B_N
* D	D
* C	C
* A_N	A_N
* VPB	VPB
* VNB	VNB
MM1015 N_VGND_M1015_d N_A_N_M1015_g N_A_27_74#_M1015_s VNB NLOWVT L=0.15 W=0.55
+ AD=0.15675 AS=0.15675 PD=1.67 PS=1.67 NRD=0 NRS=0 M=1 R=3.66667 SA=75000.2
+ SB=75000.2 A=0.0825 P=1.4 MULT=1
MM1006 A_312_82# N_A_27_74#_M1006_g N_A_225_82#_M1006_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.0888 AS=0.2109 PD=0.98 PS=2.05 NRD=10.536 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75003.4 A=0.111 P=1.78 MULT=1
MM1003 A_390_82# N_A_354_252#_M1003_g A_312_82# VNB NLOWVT L=0.15 W=0.74
+ AD=0.1443 AS=0.0888 PD=1.13 PS=0.98 NRD=22.692 NRS=10.536 M=1 R=4.93333
+ SA=75000.6 SB=75003 A=0.111 P=1.78 MULT=1
MM1013 A_498_82# N_C_M1013_g A_390_82# VNB NLOWVT L=0.15 W=0.74 AD=0.1332
+ AS=0.1443 PD=1.1 PS=1.13 NRD=20.268 NRS=22.692 M=1 R=4.93333 SA=75001.1
+ SB=75002.4 A=0.111 P=1.78 MULT=1
MM1014 N_VGND_M1014_d N_D_M1014_g A_498_82# VNB NLOWVT L=0.15 W=0.74 AD=0.2553
+ AS=0.1332 PD=1.43 PS=1.1 NRD=0 NRS=20.268 M=1 R=4.93333 SA=75001.6 SB=75001.9
+ A=0.111 P=1.78 MULT=1
MM1004 N_X_M1004_d N_A_225_82#_M1004_g N_VGND_M1014_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.2553 PD=1.02 PS=1.43 NRD=0 NRS=66.48 M=1 R=4.93333 SA=75002.5
+ SB=75001.1 A=0.111 P=1.78 MULT=1
MM1012 N_X_M1004_d N_A_225_82#_M1012_g N_VGND_M1012_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.216866 PD=1.02 PS=1.61767 NRD=0 NRS=38.604 M=1 R=4.93333
+ SA=75002.9 SB=75000.7 A=0.111 P=1.78 MULT=1
MM1010 N_A_354_252#_M1010_d N_B_N_M1010_g N_VGND_M1012_s VNB NLOWVT L=0.15
+ W=0.55 AD=0.15675 AS=0.161184 PD=1.67 PS=1.20233 NRD=0 NRS=51.936 M=1
+ R=3.66667 SA=75003.5 SB=75000.2 A=0.0825 P=1.4 MULT=1
MM1005 N_VPWR_M1005_d N_A_N_M1005_g N_A_27_74#_M1005_s VPB PSHORT L=0.15 W=0.84
+ AD=0.182609 AS=0.2478 PD=1.29652 PS=2.27 NRD=31.0669 NRS=2.3443 M=1 R=5.6
+ SA=75000.2 SB=75004.3 A=0.126 P=1.98 MULT=1
MM1001 N_A_225_82#_M1001_d N_A_27_74#_M1001_g N_VPWR_M1005_d VPB PSHORT L=0.15
+ W=1 AD=0.285 AS=0.217391 PD=1.57 PS=1.54348 NRD=41.3503 NRS=1.9503 M=1
+ R=6.66667 SA=75000.7 SB=75003.7 A=0.15 P=2.3 MULT=1
MM1000 N_VPWR_M1000_d N_A_354_252#_M1000_g N_A_225_82#_M1001_d VPB PSHORT L=0.15
+ W=1 AD=0.255 AS=0.285 PD=1.51 PS=1.57 NRD=24.6053 NRS=15.7403 M=1 R=6.66667
+ SA=75001.4 SB=75003 A=0.15 P=2.3 MULT=1
MM1008 N_A_225_82#_M1008_d N_C_M1008_g N_VPWR_M1000_d VPB PSHORT L=0.15 W=1
+ AD=0.15 AS=0.255 PD=1.3 PS=1.51 NRD=1.9503 NRS=20.685 M=1 R=6.66667 SA=75002.1
+ SB=75002.3 A=0.15 P=2.3 MULT=1
MM1009 N_VPWR_M1009_d N_D_M1009_g N_A_225_82#_M1008_d VPB PSHORT L=0.15 W=1
+ AD=0.309811 AS=0.15 PD=1.64623 PS=1.3 NRD=29.55 NRS=1.9503 M=1 R=6.66667
+ SA=75002.5 SB=75001.8 A=0.15 P=2.3 MULT=1
MM1002 N_X_M1002_d N_A_225_82#_M1002_g N_VPWR_M1009_d VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.346989 PD=1.42 PS=1.84377 NRD=1.7533 NRS=34.2977 M=1 R=7.46667
+ SA=75003 SB=75001.1 A=0.168 P=2.54 MULT=1
MM1007 N_X_M1002_d N_A_225_82#_M1007_g N_VPWR_M1007_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.232 PD=1.42 PS=1.72 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75003.4 SB=75000.6 A=0.168 P=2.54 MULT=1
MM1011 N_A_354_252#_M1011_d N_B_N_M1011_g N_VPWR_M1007_s VPB PSHORT L=0.15
+ W=0.84 AD=0.2604 AS=0.174 PD=2.3 PS=1.29 NRD=3.5066 NRS=22.261 M=1 R=5.6
+ SA=75003.9 SB=75000.2 A=0.126 P=1.98 MULT=1
DX16_noxref VNB VPB NWDIODE A=10.5276 P=15.04
c_47 VNB 0 1.18904e-19 $X=0 $Y=0
c_95 VPB 0 1.46091e-19 $X=0 $Y=3.085
*
.include "sky130_fd_sc_hs__and4bb_2.pxi.spice"
*
.ends
*
*
