* File: sky130_fd_sc_hs__or3_1.pex.spice
* Created: Tue Sep  1 20:20:25 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HS__OR3_1%C 3 5 7 8 12
r26 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.405
+ $Y=1.515 $X2=0.405 $Y2=1.515
r27 8 12 4.42216 $w=4.28e-07 $l=1.65e-07 $layer=LI1_cond $X=0.24 $Y=1.565
+ $X2=0.405 $Y2=1.565
r28 5 11 52.4131 $w=2.96e-07 $l=2.93684e-07 $layer=POLY_cond $X=0.505 $Y=1.765
+ $X2=0.41 $Y2=1.515
r29 5 7 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=0.505 $Y=1.765
+ $X2=0.505 $Y2=2.34
r30 1 11 38.5718 $w=2.96e-07 $l=2.03101e-07 $layer=POLY_cond $X=0.495 $Y=1.35
+ $X2=0.41 $Y2=1.515
r31 1 3 361.5 $w=1.5e-07 $l=7.05e-07 $layer=POLY_cond $X=0.495 $Y=1.35 $X2=0.495
+ $Y2=0.645
.ends

.subckt PM_SKY130_FD_SC_HS__OR3_1%B 1 3 6 8
c30 8 0 1.14577e-19 $X=1.2 $Y=1.665
r31 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1 $Y=1.515
+ $X2=1 $Y2=1.515
r32 8 12 5.3602 $w=4.28e-07 $l=2e-07 $layer=LI1_cond $X=1.2 $Y=1.565 $X2=1
+ $Y2=1.565
r33 4 11 38.5562 $w=2.99e-07 $l=1.67481e-07 $layer=POLY_cond $X=0.995 $Y=1.35
+ $X2=1 $Y2=1.515
r34 4 6 361.5 $w=1.5e-07 $l=7.05e-07 $layer=POLY_cond $X=0.995 $Y=1.35 $X2=0.995
+ $Y2=0.645
r35 1 11 52.2586 $w=2.99e-07 $l=2.85044e-07 $layer=POLY_cond $X=0.925 $Y=1.765
+ $X2=1 $Y2=1.515
r36 1 3 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=0.925 $Y=1.765
+ $X2=0.925 $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_HS__OR3_1%A 1 3 6 8 12 13
c35 6 0 7.84672e-20 $X=1.81 $Y=0.645
c36 1 0 1.14577e-19 $X=1.495 $Y=1.765
r37 12 14 21.3629 $w=3.61e-07 $l=1.6e-07 $layer=POLY_cond $X=1.65 $Y=1.557
+ $X2=1.81 $Y2=1.557
r38 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.65
+ $Y=1.515 $X2=1.65 $Y2=1.515
r39 10 12 20.6953 $w=3.61e-07 $l=1.55e-07 $layer=POLY_cond $X=1.495 $Y=1.557
+ $X2=1.65 $Y2=1.557
r40 8 13 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=1.65 $Y=1.665
+ $X2=1.65 $Y2=1.515
r41 4 14 23.3725 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.81 $Y=1.35
+ $X2=1.81 $Y2=1.557
r42 4 6 361.5 $w=1.5e-07 $l=7.05e-07 $layer=POLY_cond $X=1.81 $Y=1.35 $X2=1.81
+ $Y2=0.645
r43 1 10 23.3725 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=1.495 $Y=1.765
+ $X2=1.495 $Y2=1.557
r44 1 3 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=1.495 $Y=1.765
+ $X2=1.495 $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_HS__OR3_1%A_27_74# 1 2 3 10 12 15 19 24 25 27 29 30 32
+ 35 36
r83 39 40 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.29
+ $Y=1.465 $X2=2.29 $Y2=1.465
r84 34 36 10.9648 $w=7.23e-07 $l=1.65e-07 $layer=LI1_cond $X=1.595 $Y=0.817
+ $X2=1.76 $Y2=0.817
r85 34 35 17.3164 $w=7.23e-07 $l=5.5e-07 $layer=LI1_cond $X=1.595 $Y=0.817
+ $X2=1.045 $Y2=0.817
r86 29 39 9.1003 $w=2.73e-07 $l=2.07918e-07 $layer=LI1_cond $X=2.175 $Y=1.63
+ $X2=2.272 $Y2=1.465
r87 29 30 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=2.175 $Y=1.63
+ $X2=2.175 $Y2=1.95
r88 27 39 16.5348 $w=2.73e-07 $l=4.51929e-07 $layer=LI1_cond $X=2.09 $Y=1.095
+ $X2=2.272 $Y2=1.465
r89 27 36 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=2.09 $Y=1.095
+ $X2=1.76 $Y2=1.095
r90 26 32 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.445 $Y=2.035
+ $X2=0.28 $Y2=2.035
r91 25 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.09 $Y=2.035
+ $X2=2.175 $Y2=1.95
r92 25 26 107.321 $w=1.68e-07 $l=1.645e-06 $layer=LI1_cond $X=2.09 $Y=2.035
+ $X2=0.445 $Y2=2.035
r93 24 35 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=0.365 $Y=1.095
+ $X2=1.045 $Y2=1.095
r94 17 24 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.24 $Y=1.01
+ $X2=0.365 $Y2=1.095
r95 17 19 16.8257 $w=2.48e-07 $l=3.65e-07 $layer=LI1_cond $X=0.24 $Y=1.01
+ $X2=0.24 $Y2=0.645
r96 13 40 38.5916 $w=2.93e-07 $l=2.03101e-07 $layer=POLY_cond $X=2.38 $Y=1.3
+ $X2=2.295 $Y2=1.465
r97 13 15 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=2.38 $Y=1.3 $X2=2.38
+ $Y2=0.74
r98 10 40 60.7998 $w=2.93e-07 $l=3.37639e-07 $layer=POLY_cond $X=2.375 $Y=1.765
+ $X2=2.295 $Y2=1.465
r99 10 12 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.375 $Y=1.765
+ $X2=2.375 $Y2=2.4
r100 3 32 300 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.115
r101 2 34 91 $w=1.7e-07 $l=6.37868e-07 $layer=licon1_NDIFF $count=2 $X=1.07
+ $Y=0.37 $X2=1.595 $Y2=0.62
r102 1 19 182 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.645
.ends

.subckt PM_SKY130_FD_SC_HS__OR3_1%VPWR 1 6 8 10 20 21 24
r26 24 25 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r27 21 25 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=2.16 $Y2=3.33
r28 20 21 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r29 18 24 14.259 $w=1.7e-07 $l=3.8e-07 $layer=LI1_cond $X=2.315 $Y=3.33
+ $X2=1.935 $Y2=3.33
r30 18 20 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=2.315 $Y=3.33
+ $X2=2.64 $Y2=3.33
r31 16 17 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r32 13 17 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=1.2 $Y2=3.33
r33 12 16 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.24 $Y=3.33 $X2=1.2
+ $Y2=3.33
r34 12 13 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r35 10 24 14.259 $w=1.7e-07 $l=3.8e-07 $layer=LI1_cond $X=1.555 $Y=3.33
+ $X2=1.935 $Y2=3.33
r36 10 16 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=1.555 $Y=3.33
+ $X2=1.2 $Y2=3.33
r37 8 25 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.44 $Y=3.33
+ $X2=2.16 $Y2=3.33
r38 8 17 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.44 $Y=3.33
+ $X2=1.2 $Y2=3.33
r39 4 24 3.03114 $w=7.6e-07 $l=8.5e-08 $layer=LI1_cond $X=1.935 $Y=3.245
+ $X2=1.935 $Y2=3.33
r40 4 6 13.6919 $w=7.58e-07 $l=8.7e-07 $layer=LI1_cond $X=1.935 $Y=3.245
+ $X2=1.935 $Y2=2.375
r41 1 6 150 $w=1.7e-07 $l=8.04177e-07 $layer=licon1_PDIFF $count=4 $X=1.57
+ $Y=1.84 $X2=2.15 $Y2=2.375
.ends

.subckt PM_SKY130_FD_SC_HS__OR3_1%X 1 2 7 9 15 16 17 28
c24 17 0 7.84672e-20 $X=2.555 $Y=0.84
r25 21 28 0.726197 $w=3.63e-07 $l=2.3e-08 $layer=LI1_cond $X=2.612 $Y=0.948
+ $X2=2.612 $Y2=0.925
r26 17 30 8.08227 $w=3.63e-07 $l=1.51e-07 $layer=LI1_cond $X=2.612 $Y=0.979
+ $X2=2.612 $Y2=1.13
r27 17 21 0.978787 $w=3.63e-07 $l=3.1e-08 $layer=LI1_cond $X=2.612 $Y=0.979
+ $X2=2.612 $Y2=0.948
r28 17 28 0.978787 $w=3.63e-07 $l=3.1e-08 $layer=LI1_cond $X=2.612 $Y=0.894
+ $X2=2.612 $Y2=0.925
r29 16 17 11.9665 $w=3.63e-07 $l=3.79e-07 $layer=LI1_cond $X=2.612 $Y=0.515
+ $X2=2.612 $Y2=0.894
r30 15 30 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=2.71 $Y=1.82 $X2=2.71
+ $Y2=1.13
r31 9 11 34.1617 $w=2.78e-07 $l=8.3e-07 $layer=LI1_cond $X=2.655 $Y=1.985
+ $X2=2.655 $Y2=2.815
r32 7 15 7.52792 $w=2.78e-07 $l=1.4e-07 $layer=LI1_cond $X=2.655 $Y=1.96
+ $X2=2.655 $Y2=1.82
r33 7 9 1.02897 $w=2.78e-07 $l=2.5e-08 $layer=LI1_cond $X=2.655 $Y=1.96
+ $X2=2.655 $Y2=1.985
r34 2 11 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=2.45
+ $Y=1.84 $X2=2.6 $Y2=2.815
r35 2 9 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=2.45
+ $Y=1.84 $X2=2.6 $Y2=1.985
r36 1 16 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.455
+ $Y=0.37 $X2=2.595 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__OR3_1%VGND 1 2 9 13 15 17 22 29 30 33 36
r34 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r35 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r36 30 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=2.16
+ $Y2=0
r37 29 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r38 27 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.26 $Y=0 $X2=2.095
+ $Y2=0
r39 27 29 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=2.26 $Y=0 $X2=2.64
+ $Y2=0
r40 26 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r41 25 26 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r42 23 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.875 $Y=0 $X2=0.71
+ $Y2=0
r43 23 25 52.5187 $w=1.68e-07 $l=8.05e-07 $layer=LI1_cond $X=0.875 $Y=0 $X2=1.68
+ $Y2=0
r44 22 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.93 $Y=0 $X2=2.095
+ $Y2=0
r45 22 25 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=1.93 $Y=0 $X2=1.68
+ $Y2=0
r46 20 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r47 19 20 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r48 17 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.545 $Y=0 $X2=0.71
+ $Y2=0
r49 17 19 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.545 $Y=0 $X2=0.24
+ $Y2=0
r50 15 26 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.44 $Y=0 $X2=1.68
+ $Y2=0
r51 15 34 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.44 $Y=0 $X2=0.72
+ $Y2=0
r52 11 36 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.095 $Y=0.085
+ $X2=2.095 $Y2=0
r53 11 13 19.5566 $w=3.28e-07 $l=5.6e-07 $layer=LI1_cond $X=2.095 $Y=0.085
+ $X2=2.095 $Y2=0.645
r54 7 33 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.71 $Y=0.085 $X2=0.71
+ $Y2=0
r55 7 9 19.5566 $w=3.28e-07 $l=5.6e-07 $layer=LI1_cond $X=0.71 $Y=0.085 $X2=0.71
+ $Y2=0.645
r56 2 13 182 $w=1.7e-07 $l=3.65205e-07 $layer=licon1_NDIFF $count=1 $X=1.885
+ $Y=0.37 $X2=2.095 $Y2=0.645
r57 1 9 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.37 $X2=0.71 $Y2=0.645
.ends

