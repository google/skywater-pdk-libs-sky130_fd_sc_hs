* NGSPICE file created from sky130_fd_sc_hs__nor3b_4.ext - technology: sky130A

.subckt sky130_fd_sc_hs__nor3b_4 A B C_N VGND VNB VPB VPWR Y
M1000 VGND a_468_264# Y VNB nlowvt w=740000u l=150000u
+  ad=2.0498e+12p pd=1.59e+07u as=1.3135e+12p ps=1.243e+07u
M1001 Y a_468_264# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1002 Y A VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1003 VGND B Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_468_264# C_N VPWR VPB pshort w=840000u l=150000u
+  ad=2.52e+11p pd=2.28e+06u as=1.3762e+12p ps=1.105e+07u
M1005 VPWR C_N a_468_264# VPB pshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_468_264# C_N VGND VNB nlowvt w=740000u l=150000u
+  ad=6.771e+11p pd=3.31e+06u as=0p ps=0u
M1007 a_126_368# A VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=1.428e+12p pd=1.151e+07u as=0p ps=0u
M1008 VGND B Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 Y a_468_264# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_27_368# B a_126_368# VPB pshort w=1.12e+06u l=150000u
+  ad=1.7248e+12p pd=1.428e+07u as=0p ps=0u
M1011 VGND A Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_126_368# B a_27_368# VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VGND a_468_264# Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_126_368# B a_27_368# VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 Y A VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_27_368# B a_126_368# VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 VPWR A a_126_368# VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 Y a_468_264# a_27_368# VPB pshort w=1.12e+06u l=150000u
+  ad=6.72e+11p pd=5.68e+06u as=0p ps=0u
M1019 a_126_368# A VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_27_368# a_468_264# Y VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 VPWR A a_126_368# VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 VGND A Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 Y a_468_264# a_27_368# VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 Y B VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 a_27_368# a_468_264# Y VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 Y B VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

