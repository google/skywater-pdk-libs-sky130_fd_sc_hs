* File: sky130_fd_sc_hs__or4b_4.spice
* Created: Thu Aug 27 21:07:20 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hs__or4b_4.pex.spice"
.subckt sky130_fd_sc_hs__or4b_4  VNB VPB B A C D_N VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* D_N	D_N
* C	C
* A	A
* B	B
* VPB	VPB
* VNB	VNB
MM1020 N_VGND_M1020_d N_B_M1020_g N_A_27_74#_M1020_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1554 AS=0.2109 PD=1.16 PS=2.05 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75002.6 A=0.111 P=1.78 MULT=1
MM1021 N_A_27_74#_M1021_d N_A_M1021_g N_VGND_M1020_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.40885 AS=0.1554 PD=1.845 PS=1.16 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75000.8
+ SB=75002 A=0.111 P=1.78 MULT=1
MM1018 N_VGND_M1018_d N_C_M1018_g N_A_27_74#_M1021_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.1554 AS=0.40885 PD=1.16 PS=1.845 NRD=1.62 NRS=11.34 M=1 R=4.93333
+ SA=75002 SB=75000.8 A=0.111 P=1.78 MULT=1
MM1019 N_A_27_74#_M1019_d N_A_563_48#_M1019_g N_VGND_M1018_d VNB NLOWVT L=0.15
+ W=0.74 AD=0.2109 AS=0.1554 PD=2.05 PS=1.16 NRD=0 NRS=21.072 M=1 R=4.93333
+ SA=75002.6 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1016 N_VGND_M1016_d N_D_N_M1016_g N_A_563_48#_M1016_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.125217 AS=0.32135 PD=1.0342 PS=2.98 NRD=15.936 NRS=15.936 M=1 R=4.26667
+ SA=75000.3 SB=75002.2 A=0.096 P=1.58 MULT=1
MM1001 N_VGND_M1016_d N_A_27_74#_M1001_g N_X_M1001_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.144783 AS=0.14985 PD=1.1958 PS=1.145 NRD=2.424 NRS=8.916 M=1 R=4.93333
+ SA=75000.8 SB=75001.7 A=0.111 P=1.78 MULT=1
MM1013 N_VGND_M1013_d N_A_27_74#_M1013_g N_X_M1001_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1295 AS=0.14985 PD=1.09 PS=1.145 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75001.3
+ SB=75001.1 A=0.111 P=1.78 MULT=1
MM1014 N_VGND_M1013_d N_A_27_74#_M1014_g N_X_M1014_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1295 AS=0.1036 PD=1.09 PS=1.02 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75001.8
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1017 N_VGND_M1017_d N_A_27_74#_M1017_g N_X_M1014_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.1036 PD=2.05 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75002.2
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1006 N_A_116_392#_M1006_d N_B_M1006_g N_A_27_392#_M1006_s VPB PSHORT L=0.15
+ W=1 AD=0.15 AS=0.295 PD=1.3 PS=2.59 NRD=1.9503 NRS=1.9503 M=1 R=6.66667
+ SA=75000.2 SB=75003.5 A=0.15 P=2.3 MULT=1
MM1007 N_VPWR_M1007_d N_A_M1007_g N_A_116_392#_M1006_d VPB PSHORT L=0.15 W=1
+ AD=0.15 AS=0.15 PD=1.3 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=6.66667 SA=75000.7
+ SB=75003.1 A=0.15 P=2.3 MULT=1
MM1010 N_VPWR_M1007_d N_A_M1010_g N_A_116_392#_M1010_s VPB PSHORT L=0.15 W=1
+ AD=0.15 AS=0.175 PD=1.3 PS=1.35 NRD=1.9503 NRS=11.8003 M=1 R=6.66667
+ SA=75001.1 SB=75002.6 A=0.15 P=2.3 MULT=1
MM1011 N_A_116_392#_M1010_s N_B_M1011_g N_A_27_392#_M1011_s VPB PSHORT L=0.15
+ W=1 AD=0.175 AS=0.175 PD=1.35 PS=1.35 NRD=1.9503 NRS=11.8003 M=1 R=6.66667
+ SA=75001.6 SB=75002.1 A=0.15 P=2.3 MULT=1
MM1009 N_A_496_392#_M1009_d N_C_M1009_g N_A_27_392#_M1011_s VPB PSHORT L=0.15
+ W=1 AD=0.175 AS=0.175 PD=1.35 PS=1.35 NRD=11.8003 NRS=1.9503 M=1 R=6.66667
+ SA=75002.1 SB=75001.6 A=0.15 P=2.3 MULT=1
MM1008 N_A_27_74#_M1008_d N_A_563_48#_M1008_g N_A_496_392#_M1009_d VPB PSHORT
+ L=0.15 W=1 AD=0.15 AS=0.175 PD=1.3 PS=1.35 NRD=1.9503 NRS=1.9503 M=1 R=6.66667
+ SA=75002.6 SB=75001.1 A=0.15 P=2.3 MULT=1
MM1012 N_A_27_74#_M1008_d N_A_563_48#_M1012_g N_A_496_392#_M1012_s VPB PSHORT
+ L=0.15 W=1 AD=0.15 AS=0.15 PD=1.3 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=6.66667
+ SA=75003.1 SB=75000.7 A=0.15 P=2.3 MULT=1
MM1015 N_A_496_392#_M1012_s N_C_M1015_g N_A_27_392#_M1015_s VPB PSHORT L=0.15
+ W=1 AD=0.15 AS=0.295 PD=1.3 PS=2.59 NRD=1.9503 NRS=1.9503 M=1 R=6.66667
+ SA=75003.5 SB=75000.2 A=0.15 P=2.3 MULT=1
MM1004 N_VPWR_M1004_d N_D_N_M1004_g N_A_563_48#_M1004_s VPB PSHORT L=0.15 W=1
+ AD=0.198302 AS=0.295 PD=1.41981 PS=2.59 NRD=19.0302 NRS=1.9503 M=1 R=6.66667
+ SA=75000.2 SB=75002.1 A=0.15 P=2.3 MULT=1
MM1000 N_X_M1000_d N_A_27_74#_M1000_g N_VPWR_M1004_d VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.222098 PD=1.42 PS=1.59019 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.7 SB=75001.6 A=0.168 P=2.54 MULT=1
MM1002 N_X_M1000_d N_A_27_74#_M1002_g N_VPWR_M1002_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.1 SB=75001.1 A=0.168 P=2.54 MULT=1
MM1003 N_X_M1003_d N_A_27_74#_M1003_g N_VPWR_M1002_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.6 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1005 N_X_M1003_d N_A_27_74#_M1005_g N_VPWR_M1005_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.3248 PD=1.42 PS=2.82 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75002 SB=75000.2 A=0.168 P=2.54 MULT=1
DX22_noxref VNB VPB NWDIODE A=14.0988 P=18.88
c_72 VNB 0 1.8329e-19 $X=0 $Y=0
c_129 VPB 0 3.16766e-20 $X=0 $Y=3.085
*
.include "sky130_fd_sc_hs__or4b_4.pxi.spice"
*
.ends
*
*
