* File: sky130_fd_sc_hs__nor4b_1.pxi.spice
* Created: Tue Sep  1 20:12:21 2020
* 
x_PM_SKY130_FD_SC_HS__NOR4B_1%D_N N_D_N_c_58_n N_D_N_c_63_n N_D_N_M1002_g
+ N_D_N_M1008_g D_N N_D_N_c_61_n PM_SKY130_FD_SC_HS__NOR4B_1%D_N
x_PM_SKY130_FD_SC_HS__NOR4B_1%A N_A_c_98_n N_A_M1004_g N_A_M1009_g A N_A_c_100_n
+ PM_SKY130_FD_SC_HS__NOR4B_1%A
x_PM_SKY130_FD_SC_HS__NOR4B_1%B N_B_c_132_n N_B_M1007_g N_B_M1006_g B
+ N_B_c_134_n PM_SKY130_FD_SC_HS__NOR4B_1%B
x_PM_SKY130_FD_SC_HS__NOR4B_1%C N_C_c_163_n N_C_M1000_g N_C_M1001_g C
+ N_C_c_165_n PM_SKY130_FD_SC_HS__NOR4B_1%C
x_PM_SKY130_FD_SC_HS__NOR4B_1%A_57_368# N_A_57_368#_M1008_s N_A_57_368#_M1002_s
+ N_A_57_368#_M1005_g N_A_57_368#_c_196_n N_A_57_368#_M1003_g
+ N_A_57_368#_c_206_n N_A_57_368#_c_201_n N_A_57_368#_c_197_n
+ N_A_57_368#_c_202_n N_A_57_368#_c_198_n N_A_57_368#_c_204_n
+ N_A_57_368#_c_199_n PM_SKY130_FD_SC_HS__NOR4B_1%A_57_368#
x_PM_SKY130_FD_SC_HS__NOR4B_1%VPWR N_VPWR_M1002_d N_VPWR_c_266_n N_VPWR_c_267_n
+ N_VPWR_c_268_n VPWR N_VPWR_c_269_n N_VPWR_c_265_n
+ PM_SKY130_FD_SC_HS__NOR4B_1%VPWR
x_PM_SKY130_FD_SC_HS__NOR4B_1%Y N_Y_M1009_d N_Y_M1001_d N_Y_M1003_d N_Y_c_295_n
+ N_Y_c_296_n N_Y_c_297_n N_Y_c_298_n N_Y_c_299_n N_Y_c_300_n Y Y Y N_Y_c_301_n
+ PM_SKY130_FD_SC_HS__NOR4B_1%Y
x_PM_SKY130_FD_SC_HS__NOR4B_1%VGND N_VGND_M1008_d N_VGND_M1006_d N_VGND_M1005_d
+ N_VGND_c_354_n N_VGND_c_355_n N_VGND_c_356_n N_VGND_c_357_n N_VGND_c_358_n
+ N_VGND_c_359_n N_VGND_c_360_n N_VGND_c_361_n VGND N_VGND_c_362_n
+ N_VGND_c_363_n PM_SKY130_FD_SC_HS__NOR4B_1%VGND
cc_1 VNB N_D_N_c_58_n 0.0134167f $X=-0.19 $Y=-0.245 $X2=0.655 $Y2=1.675
cc_2 VNB N_D_N_M1008_g 0.0280622f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=0.645
cc_3 VNB D_N 0.00776204f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_4 VNB N_D_N_c_61_n 0.035461f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.275
cc_5 VNB N_A_c_98_n 0.0265542f $X=-0.19 $Y=-0.245 $X2=0.655 $Y2=1.44
cc_6 VNB N_A_M1009_g 0.0259031f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=1.11
cc_7 VNB N_A_c_100_n 0.00355186f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.275
cc_8 VNB N_B_c_132_n 0.026233f $X=-0.19 $Y=-0.245 $X2=0.655 $Y2=1.44
cc_9 VNB N_B_M1006_g 0.0258898f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=1.11
cc_10 VNB N_B_c_134_n 0.00165719f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.275
cc_11 VNB N_C_c_163_n 0.0242458f $X=-0.19 $Y=-0.245 $X2=0.655 $Y2=1.44
cc_12 VNB N_C_M1001_g 0.0258908f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=1.11
cc_13 VNB N_C_c_165_n 0.00381276f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.275
cc_14 VNB N_A_57_368#_M1005_g 0.0264924f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_57_368#_c_196_n 0.0272591f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_57_368#_c_197_n 0.0401545f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_57_368#_c_198_n 0.0356004f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_57_368#_c_199_n 0.00512013f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_VPWR_c_265_n 0.143779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_Y_c_295_n 0.00240191f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.275
cc_21 VNB N_Y_c_296_n 0.00823886f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.275
cc_22 VNB N_Y_c_297_n 0.0090164f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.11
cc_23 VNB N_Y_c_298_n 0.00240191f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_Y_c_299_n 0.0181248f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_Y_c_300_n 0.00775352f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_Y_c_301_n 0.0230123f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_VGND_c_354_n 0.0134539f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.275
cc_28 VNB N_VGND_c_355_n 0.00907103f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.44
cc_29 VNB N_VGND_c_356_n 0.0158851f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_357_n 0.0313058f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_358_n 0.0232674f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_359_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_360_n 0.0186948f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_361_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_362_n 0.019013f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_363_n 0.211126f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VPB N_D_N_c_58_n 8.57692e-19 $X=-0.19 $Y=1.66 $X2=0.655 $Y2=1.675
cc_38 VPB N_D_N_c_63_n 0.0271117f $X=-0.19 $Y=1.66 $X2=0.655 $Y2=1.765
cc_39 VPB N_A_c_98_n 0.0284143f $X=-0.19 $Y=1.66 $X2=0.655 $Y2=1.44
cc_40 VPB N_A_c_100_n 0.00286025f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=1.275
cc_41 VPB N_B_c_132_n 0.0268225f $X=-0.19 $Y=1.66 $X2=0.655 $Y2=1.44
cc_42 VPB N_B_c_134_n 0.00296273f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=1.275
cc_43 VPB N_C_c_163_n 0.0282492f $X=-0.19 $Y=1.66 $X2=0.655 $Y2=1.44
cc_44 VPB N_C_c_165_n 0.00328097f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=1.275
cc_45 VPB N_A_57_368#_c_196_n 0.0341574f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_46 VPB N_A_57_368#_c_201_n 0.00142313f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_47 VPB N_A_57_368#_c_202_n 0.0219494f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_48 VPB N_A_57_368#_c_198_n 0.00813831f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_49 VPB N_A_57_368#_c_204_n 0.0328014f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_50 VPB N_A_57_368#_c_199_n 4.03371e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_51 VPB N_VPWR_c_266_n 0.0171181f $X=-0.19 $Y=1.66 $X2=0.67 $Y2=1.11
cc_52 VPB N_VPWR_c_267_n 0.0265205f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_53 VPB N_VPWR_c_268_n 0.00614127f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.21
cc_54 VPB N_VPWR_c_269_n 0.0689598f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_55 VPB N_VPWR_c_265_n 0.10567f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_56 VPB Y 0.0487223f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_57 VPB N_Y_c_301_n 0.00903339f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_58 N_D_N_c_58_n N_A_c_98_n 0.0135175f $X=0.655 $Y=1.675 $X2=-0.19 $Y2=-0.245
cc_59 N_D_N_c_63_n N_A_c_98_n 0.0220221f $X=0.655 $Y=1.765 $X2=-0.19 $Y2=-0.245
cc_60 D_N N_A_c_98_n 5.07587e-19 $X=0.635 $Y=1.21 $X2=-0.19 $Y2=-0.245
cc_61 N_D_N_c_61_n N_A_c_98_n 0.00563717f $X=0.61 $Y=1.275 $X2=-0.19 $Y2=-0.245
cc_62 N_D_N_M1008_g N_A_M1009_g 0.0184418f $X=0.67 $Y=0.645 $X2=0 $Y2=0
cc_63 D_N N_A_M1009_g 0.00400388f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_64 N_D_N_c_61_n N_A_M1009_g 0.00644195f $X=0.61 $Y=1.275 $X2=0 $Y2=0
cc_65 N_D_N_c_58_n N_A_c_100_n 0.00157569f $X=0.655 $Y=1.675 $X2=0 $Y2=0
cc_66 N_D_N_c_63_n N_A_c_100_n 0.00227246f $X=0.655 $Y=1.765 $X2=0 $Y2=0
cc_67 D_N N_A_c_100_n 0.00714274f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_68 N_D_N_c_63_n N_A_57_368#_c_206_n 0.0146705f $X=0.655 $Y=1.765 $X2=0 $Y2=0
cc_69 D_N N_A_57_368#_c_206_n 0.00584907f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_70 N_D_N_M1008_g N_A_57_368#_c_197_n 0.0111596f $X=0.67 $Y=0.645 $X2=0 $Y2=0
cc_71 D_N N_A_57_368#_c_197_n 0.0144068f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_72 N_D_N_c_61_n N_A_57_368#_c_197_n 0.0035824f $X=0.61 $Y=1.275 $X2=0 $Y2=0
cc_73 N_D_N_c_63_n N_A_57_368#_c_202_n 0.00467115f $X=0.655 $Y=1.765 $X2=0 $Y2=0
cc_74 D_N N_A_57_368#_c_202_n 0.00684172f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_75 N_D_N_c_61_n N_A_57_368#_c_202_n 0.00245637f $X=0.61 $Y=1.275 $X2=0 $Y2=0
cc_76 N_D_N_c_58_n N_A_57_368#_c_198_n 0.00996102f $X=0.655 $Y=1.675 $X2=0 $Y2=0
cc_77 N_D_N_c_63_n N_A_57_368#_c_198_n 0.00160056f $X=0.655 $Y=1.765 $X2=0 $Y2=0
cc_78 N_D_N_M1008_g N_A_57_368#_c_198_n 0.0049454f $X=0.67 $Y=0.645 $X2=0 $Y2=0
cc_79 D_N N_A_57_368#_c_198_n 0.0249903f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_80 N_D_N_c_61_n N_A_57_368#_c_198_n 0.00231223f $X=0.61 $Y=1.275 $X2=0 $Y2=0
cc_81 N_D_N_c_63_n N_A_57_368#_c_204_n 0.0123352f $X=0.655 $Y=1.765 $X2=0 $Y2=0
cc_82 N_D_N_c_63_n N_VPWR_c_266_n 0.0068216f $X=0.655 $Y=1.765 $X2=0 $Y2=0
cc_83 N_D_N_c_63_n N_VPWR_c_267_n 0.00393873f $X=0.655 $Y=1.765 $X2=0 $Y2=0
cc_84 N_D_N_c_63_n N_VPWR_c_265_n 0.00462577f $X=0.655 $Y=1.765 $X2=0 $Y2=0
cc_85 N_D_N_M1008_g N_Y_c_295_n 4.34666e-19 $X=0.67 $Y=0.645 $X2=0 $Y2=0
cc_86 N_D_N_M1008_g N_Y_c_297_n 4.50506e-19 $X=0.67 $Y=0.645 $X2=0 $Y2=0
cc_87 D_N N_Y_c_297_n 0.00269803f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_88 N_D_N_M1008_g N_VGND_c_354_n 0.00693523f $X=0.67 $Y=0.645 $X2=0 $Y2=0
cc_89 D_N N_VGND_c_354_n 0.00212308f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_90 N_D_N_M1008_g N_VGND_c_358_n 0.00433162f $X=0.67 $Y=0.645 $X2=0 $Y2=0
cc_91 N_D_N_M1008_g N_VGND_c_363_n 0.00821785f $X=0.67 $Y=0.645 $X2=0 $Y2=0
cc_92 N_A_c_98_n N_B_c_132_n 0.0889312f $X=1.225 $Y=1.765 $X2=-0.19 $Y2=-0.245
cc_93 N_A_c_100_n N_B_c_132_n 0.00130194f $X=1.15 $Y=1.515 $X2=-0.19 $Y2=-0.245
cc_94 N_A_M1009_g N_B_M1006_g 0.019972f $X=1.24 $Y=0.74 $X2=0 $Y2=0
cc_95 N_A_c_98_n N_B_c_134_n 0.00168387f $X=1.225 $Y=1.765 $X2=0 $Y2=0
cc_96 N_A_c_100_n N_B_c_134_n 0.0277335f $X=1.15 $Y=1.515 $X2=0 $Y2=0
cc_97 N_A_c_98_n N_A_57_368#_c_206_n 0.0159168f $X=1.225 $Y=1.765 $X2=0 $Y2=0
cc_98 N_A_c_100_n N_A_57_368#_c_206_n 0.0226548f $X=1.15 $Y=1.515 $X2=0 $Y2=0
cc_99 N_A_c_98_n N_A_57_368#_c_202_n 0.00135095f $X=1.225 $Y=1.765 $X2=0 $Y2=0
cc_100 N_A_c_98_n N_VPWR_c_266_n 0.0170305f $X=1.225 $Y=1.765 $X2=0 $Y2=0
cc_101 N_A_c_98_n N_VPWR_c_269_n 0.00413917f $X=1.225 $Y=1.765 $X2=0 $Y2=0
cc_102 N_A_c_98_n N_VPWR_c_265_n 0.00817532f $X=1.225 $Y=1.765 $X2=0 $Y2=0
cc_103 N_A_M1009_g N_Y_c_295_n 0.00863911f $X=1.24 $Y=0.74 $X2=0 $Y2=0
cc_104 N_A_M1009_g N_Y_c_297_n 0.00453747f $X=1.24 $Y=0.74 $X2=0 $Y2=0
cc_105 N_A_c_100_n N_Y_c_297_n 0.00196319f $X=1.15 $Y=1.515 $X2=0 $Y2=0
cc_106 N_A_c_98_n N_VGND_c_354_n 8.85031e-19 $X=1.225 $Y=1.765 $X2=0 $Y2=0
cc_107 N_A_M1009_g N_VGND_c_354_n 0.00545144f $X=1.24 $Y=0.74 $X2=0 $Y2=0
cc_108 N_A_c_100_n N_VGND_c_354_n 0.00542787f $X=1.15 $Y=1.515 $X2=0 $Y2=0
cc_109 N_A_M1009_g N_VGND_c_360_n 0.00434272f $X=1.24 $Y=0.74 $X2=0 $Y2=0
cc_110 N_A_M1009_g N_VGND_c_363_n 0.0082141f $X=1.24 $Y=0.74 $X2=0 $Y2=0
cc_111 N_B_c_132_n N_C_c_163_n 0.0758679f $X=1.645 $Y=1.765 $X2=-0.19 $Y2=-0.245
cc_112 N_B_c_134_n N_C_c_163_n 7.55505e-19 $X=1.69 $Y=1.515 $X2=-0.19 $Y2=-0.245
cc_113 N_B_M1006_g N_C_M1001_g 0.0252177f $X=1.67 $Y=0.74 $X2=0 $Y2=0
cc_114 N_B_c_132_n N_C_c_165_n 0.00217395f $X=1.645 $Y=1.765 $X2=0 $Y2=0
cc_115 N_B_c_134_n N_C_c_165_n 0.0318722f $X=1.69 $Y=1.515 $X2=0 $Y2=0
cc_116 N_B_c_132_n N_A_57_368#_c_206_n 0.0159139f $X=1.645 $Y=1.765 $X2=0 $Y2=0
cc_117 N_B_c_134_n N_A_57_368#_c_206_n 0.0215605f $X=1.69 $Y=1.515 $X2=0 $Y2=0
cc_118 N_B_c_132_n N_VPWR_c_266_n 0.00385876f $X=1.645 $Y=1.765 $X2=0 $Y2=0
cc_119 N_B_c_132_n N_VPWR_c_269_n 0.00461464f $X=1.645 $Y=1.765 $X2=0 $Y2=0
cc_120 N_B_c_132_n N_VPWR_c_265_n 0.00910115f $X=1.645 $Y=1.765 $X2=0 $Y2=0
cc_121 N_B_M1006_g N_Y_c_295_n 0.00969128f $X=1.67 $Y=0.74 $X2=0 $Y2=0
cc_122 N_B_c_132_n N_Y_c_296_n 7.68393e-19 $X=1.645 $Y=1.765 $X2=0 $Y2=0
cc_123 N_B_M1006_g N_Y_c_296_n 0.0118338f $X=1.67 $Y=0.74 $X2=0 $Y2=0
cc_124 N_B_c_134_n N_Y_c_296_n 0.0175347f $X=1.69 $Y=1.515 $X2=0 $Y2=0
cc_125 N_B_c_132_n N_Y_c_297_n 5.43336e-19 $X=1.645 $Y=1.765 $X2=0 $Y2=0
cc_126 N_B_M1006_g N_Y_c_297_n 0.0015571f $X=1.67 $Y=0.74 $X2=0 $Y2=0
cc_127 N_B_c_134_n N_Y_c_297_n 0.00799991f $X=1.69 $Y=1.515 $X2=0 $Y2=0
cc_128 N_B_M1006_g N_Y_c_298_n 8.70047e-19 $X=1.67 $Y=0.74 $X2=0 $Y2=0
cc_129 N_B_M1006_g N_VGND_c_355_n 0.00491516f $X=1.67 $Y=0.74 $X2=0 $Y2=0
cc_130 N_B_M1006_g N_VGND_c_360_n 0.00434272f $X=1.67 $Y=0.74 $X2=0 $Y2=0
cc_131 N_B_M1006_g N_VGND_c_363_n 0.00821482f $X=1.67 $Y=0.74 $X2=0 $Y2=0
cc_132 N_C_M1001_g N_A_57_368#_M1005_g 0.0199815f $X=2.25 $Y=0.74 $X2=0 $Y2=0
cc_133 N_C_c_163_n N_A_57_368#_c_196_n 0.0623738f $X=2.155 $Y=1.765 $X2=0 $Y2=0
cc_134 N_C_c_165_n N_A_57_368#_c_196_n 7.0116e-19 $X=2.23 $Y=1.515 $X2=0 $Y2=0
cc_135 N_C_c_163_n N_A_57_368#_c_206_n 0.0168272f $X=2.155 $Y=1.765 $X2=0 $Y2=0
cc_136 N_C_c_165_n N_A_57_368#_c_206_n 0.0235257f $X=2.23 $Y=1.515 $X2=0 $Y2=0
cc_137 N_C_c_163_n N_A_57_368#_c_201_n 0.0032952f $X=2.155 $Y=1.765 $X2=0 $Y2=0
cc_138 N_C_c_165_n N_A_57_368#_c_201_n 0.00796423f $X=2.23 $Y=1.515 $X2=0 $Y2=0
cc_139 N_C_c_163_n N_A_57_368#_c_199_n 0.00187066f $X=2.155 $Y=1.765 $X2=0 $Y2=0
cc_140 N_C_c_165_n N_A_57_368#_c_199_n 0.0264357f $X=2.23 $Y=1.515 $X2=0 $Y2=0
cc_141 N_C_c_163_n N_VPWR_c_269_n 0.00461464f $X=2.155 $Y=1.765 $X2=0 $Y2=0
cc_142 N_C_c_163_n N_VPWR_c_265_n 0.00911364f $X=2.155 $Y=1.765 $X2=0 $Y2=0
cc_143 N_C_M1001_g N_Y_c_295_n 8.64794e-19 $X=2.25 $Y=0.74 $X2=0 $Y2=0
cc_144 N_C_c_163_n N_Y_c_296_n 7.6608e-19 $X=2.155 $Y=1.765 $X2=0 $Y2=0
cc_145 N_C_M1001_g N_Y_c_296_n 0.0118338f $X=2.25 $Y=0.74 $X2=0 $Y2=0
cc_146 N_C_c_165_n N_Y_c_296_n 0.0191575f $X=2.23 $Y=1.515 $X2=0 $Y2=0
cc_147 N_C_M1001_g N_Y_c_298_n 0.00980887f $X=2.25 $Y=0.74 $X2=0 $Y2=0
cc_148 N_C_c_163_n N_Y_c_300_n 5.46117e-19 $X=2.155 $Y=1.765 $X2=0 $Y2=0
cc_149 N_C_M1001_g N_Y_c_300_n 0.0015571f $X=2.25 $Y=0.74 $X2=0 $Y2=0
cc_150 N_C_c_165_n N_Y_c_300_n 0.00799991f $X=2.23 $Y=1.515 $X2=0 $Y2=0
cc_151 N_C_M1001_g N_VGND_c_355_n 0.0061968f $X=2.25 $Y=0.74 $X2=0 $Y2=0
cc_152 N_C_M1001_g N_VGND_c_362_n 0.00434272f $X=2.25 $Y=0.74 $X2=0 $Y2=0
cc_153 N_C_M1001_g N_VGND_c_363_n 0.00821706f $X=2.25 $Y=0.74 $X2=0 $Y2=0
cc_154 N_A_57_368#_c_206_n N_VPWR_M1002_d 0.0131231f $X=2.565 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_155 N_A_57_368#_c_206_n N_VPWR_c_266_n 0.0219335f $X=2.565 $Y=2.035 $X2=0
+ $Y2=0
cc_156 N_A_57_368#_c_204_n N_VPWR_c_266_n 0.025186f $X=0.35 $Y=2.035 $X2=0 $Y2=0
cc_157 N_A_57_368#_c_204_n N_VPWR_c_267_n 0.00995358f $X=0.35 $Y=2.035 $X2=0
+ $Y2=0
cc_158 N_A_57_368#_c_196_n N_VPWR_c_269_n 0.00461464f $X=2.725 $Y=1.765 $X2=0
+ $Y2=0
cc_159 N_A_57_368#_c_196_n N_VPWR_c_265_n 0.0091462f $X=2.725 $Y=1.765 $X2=0
+ $Y2=0
cc_160 N_A_57_368#_c_204_n N_VPWR_c_265_n 0.0148468f $X=0.35 $Y=2.035 $X2=0
+ $Y2=0
cc_161 N_A_57_368#_c_206_n A_260_368# 0.0119045f $X=2.565 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_162 N_A_57_368#_c_206_n A_344_368# 0.0165022f $X=2.565 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_163 N_A_57_368#_c_206_n A_446_368# 0.0196974f $X=2.565 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_164 N_A_57_368#_c_201_n A_446_368# 0.00144634f $X=2.65 $Y=1.95 $X2=-0.19
+ $Y2=-0.245
cc_165 N_A_57_368#_M1005_g N_Y_c_298_n 0.01371f $X=2.68 $Y=0.74 $X2=0 $Y2=0
cc_166 N_A_57_368#_M1005_g N_Y_c_299_n 0.0129008f $X=2.68 $Y=0.74 $X2=0 $Y2=0
cc_167 N_A_57_368#_c_196_n N_Y_c_299_n 0.00422928f $X=2.725 $Y=1.765 $X2=0 $Y2=0
cc_168 N_A_57_368#_c_199_n N_Y_c_299_n 0.0224209f $X=2.77 $Y=1.515 $X2=0 $Y2=0
cc_169 N_A_57_368#_M1005_g N_Y_c_300_n 0.00155819f $X=2.68 $Y=0.74 $X2=0 $Y2=0
cc_170 N_A_57_368#_c_199_n N_Y_c_300_n 0.00553408f $X=2.77 $Y=1.515 $X2=0 $Y2=0
cc_171 N_A_57_368#_c_196_n Y 0.0411062f $X=2.725 $Y=1.765 $X2=0 $Y2=0
cc_172 N_A_57_368#_c_206_n Y 0.0140855f $X=2.565 $Y=2.035 $X2=0 $Y2=0
cc_173 N_A_57_368#_c_201_n Y 0.00743442f $X=2.65 $Y=1.95 $X2=0 $Y2=0
cc_174 N_A_57_368#_c_199_n Y 0.00239484f $X=2.77 $Y=1.515 $X2=0 $Y2=0
cc_175 N_A_57_368#_M1005_g N_Y_c_301_n 0.00477786f $X=2.68 $Y=0.74 $X2=0 $Y2=0
cc_176 N_A_57_368#_c_196_n N_Y_c_301_n 0.00544381f $X=2.725 $Y=1.765 $X2=0 $Y2=0
cc_177 N_A_57_368#_c_201_n N_Y_c_301_n 0.00676462f $X=2.65 $Y=1.95 $X2=0 $Y2=0
cc_178 N_A_57_368#_c_199_n N_Y_c_301_n 0.0249903f $X=2.77 $Y=1.515 $X2=0 $Y2=0
cc_179 N_A_57_368#_c_197_n N_VGND_c_354_n 0.0252474f $X=0.455 $Y=0.645 $X2=0
+ $Y2=0
cc_180 N_A_57_368#_M1005_g N_VGND_c_357_n 0.0141934f $X=2.68 $Y=0.74 $X2=0 $Y2=0
cc_181 N_A_57_368#_c_197_n N_VGND_c_358_n 0.0225742f $X=0.455 $Y=0.645 $X2=0
+ $Y2=0
cc_182 N_A_57_368#_M1005_g N_VGND_c_362_n 0.00434272f $X=2.68 $Y=0.74 $X2=0
+ $Y2=0
cc_183 N_A_57_368#_M1005_g N_VGND_c_363_n 0.00824301f $X=2.68 $Y=0.74 $X2=0
+ $Y2=0
cc_184 N_A_57_368#_c_197_n N_VGND_c_363_n 0.0187953f $X=0.455 $Y=0.645 $X2=0
+ $Y2=0
cc_185 N_VPWR_c_269_n Y 0.0164205f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_186 N_VPWR_c_265_n Y 0.0135915f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_187 N_Y_c_296_n N_VGND_M1006_d 0.00374272f $X=2.3 $Y=1.095 $X2=0 $Y2=0
cc_188 N_Y_c_299_n N_VGND_M1005_d 0.00411309f $X=3.105 $Y=1.095 $X2=0 $Y2=0
cc_189 N_Y_c_295_n N_VGND_c_354_n 0.0229287f $X=1.455 $Y=0.515 $X2=0 $Y2=0
cc_190 N_Y_c_295_n N_VGND_c_355_n 0.0191765f $X=1.455 $Y=0.515 $X2=0 $Y2=0
cc_191 N_Y_c_296_n N_VGND_c_355_n 0.0257093f $X=2.3 $Y=1.095 $X2=0 $Y2=0
cc_192 N_Y_c_298_n N_VGND_c_355_n 0.0183215f $X=2.465 $Y=0.515 $X2=0 $Y2=0
cc_193 N_Y_c_298_n N_VGND_c_357_n 0.0191765f $X=2.465 $Y=0.515 $X2=0 $Y2=0
cc_194 N_Y_c_299_n N_VGND_c_357_n 0.0260326f $X=3.105 $Y=1.095 $X2=0 $Y2=0
cc_195 N_Y_c_295_n N_VGND_c_360_n 0.0144922f $X=1.455 $Y=0.515 $X2=0 $Y2=0
cc_196 N_Y_c_298_n N_VGND_c_362_n 0.0144922f $X=2.465 $Y=0.515 $X2=0 $Y2=0
cc_197 N_Y_c_295_n N_VGND_c_363_n 0.0118826f $X=1.455 $Y=0.515 $X2=0 $Y2=0
cc_198 N_Y_c_298_n N_VGND_c_363_n 0.0118826f $X=2.465 $Y=0.515 $X2=0 $Y2=0
