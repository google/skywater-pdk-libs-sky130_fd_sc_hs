* File: sky130_fd_sc_hs__o21ba_1.pxi.spice
* Created: Tue Sep  1 20:14:49 2020
* 
x_PM_SKY130_FD_SC_HS__O21BA_1%A1 N_A1_c_73_n N_A1_M1008_g N_A1_c_78_n
+ N_A1_M1002_g A1 A1 N_A1_c_75_n N_A1_c_76_n PM_SKY130_FD_SC_HS__O21BA_1%A1
x_PM_SKY130_FD_SC_HS__O21BA_1%A2 N_A2_c_106_n N_A2_M1007_g N_A2_M1009_g
+ N_A2_c_102_n N_A2_c_103_n A2 A2 N_A2_c_105_n PM_SKY130_FD_SC_HS__O21BA_1%A2
x_PM_SKY130_FD_SC_HS__O21BA_1%A_281_244# N_A_281_244#_M1005_s
+ N_A_281_244#_M1001_s N_A_281_244#_c_141_n N_A_281_244#_c_151_n
+ N_A_281_244#_M1006_g N_A_281_244#_M1003_g N_A_281_244#_c_143_n
+ N_A_281_244#_c_144_n N_A_281_244#_c_145_n N_A_281_244#_c_146_n
+ N_A_281_244#_c_153_n N_A_281_244#_c_154_n N_A_281_244#_c_147_n
+ N_A_281_244#_c_148_n N_A_281_244#_c_149_n
+ PM_SKY130_FD_SC_HS__O21BA_1%A_281_244#
x_PM_SKY130_FD_SC_HS__O21BA_1%B1_N N_B1_N_c_202_n N_B1_N_M1001_g N_B1_N_c_203_n
+ N_B1_N_M1005_g B1_N PM_SKY130_FD_SC_HS__O21BA_1%B1_N
x_PM_SKY130_FD_SC_HS__O21BA_1%A_200_392# N_A_200_392#_M1003_d
+ N_A_200_392#_M1007_d N_A_200_392#_c_233_n N_A_200_392#_M1004_g
+ N_A_200_392#_M1000_g N_A_200_392#_c_235_n N_A_200_392#_c_236_n
+ N_A_200_392#_c_242_n N_A_200_392#_c_237_n N_A_200_392#_c_244_n
+ N_A_200_392#_c_248_n N_A_200_392#_c_238_n N_A_200_392#_c_239_n
+ PM_SKY130_FD_SC_HS__O21BA_1%A_200_392#
x_PM_SKY130_FD_SC_HS__O21BA_1%VPWR N_VPWR_M1002_s N_VPWR_M1006_d N_VPWR_M1001_d
+ N_VPWR_c_314_n N_VPWR_c_315_n N_VPWR_c_316_n N_VPWR_c_317_n VPWR
+ N_VPWR_c_318_n N_VPWR_c_319_n N_VPWR_c_320_n N_VPWR_c_313_n N_VPWR_c_322_n
+ N_VPWR_c_323_n PM_SKY130_FD_SC_HS__O21BA_1%VPWR
x_PM_SKY130_FD_SC_HS__O21BA_1%X N_X_M1000_d N_X_M1004_d N_X_c_358_n N_X_c_359_n
+ X X X X N_X_c_360_n PM_SKY130_FD_SC_HS__O21BA_1%X
x_PM_SKY130_FD_SC_HS__O21BA_1%A_27_74# N_A_27_74#_M1008_s N_A_27_74#_M1009_d
+ N_A_27_74#_c_384_n N_A_27_74#_c_388_n N_A_27_74#_c_385_n N_A_27_74#_c_386_n
+ PM_SKY130_FD_SC_HS__O21BA_1%A_27_74#
x_PM_SKY130_FD_SC_HS__O21BA_1%VGND N_VGND_M1008_d N_VGND_M1005_d N_VGND_c_411_n
+ N_VGND_c_412_n VGND N_VGND_c_413_n N_VGND_c_414_n N_VGND_c_415_n
+ N_VGND_c_416_n N_VGND_c_417_n N_VGND_c_418_n PM_SKY130_FD_SC_HS__O21BA_1%VGND
cc_1 VNB N_A1_c_73_n 0.0298684f $X=-0.19 $Y=-0.245 $X2=0.395 $Y2=1.625
cc_2 VNB A1 0.0231282f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_3 VNB N_A1_c_75_n 0.020516f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.295
cc_4 VNB N_A1_c_76_n 0.0261918f $X=-0.19 $Y=-0.245 $X2=0.395 $Y2=1.13
cc_5 VNB N_A2_c_102_n 0.019683f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.46
cc_6 VNB N_A2_c_103_n 0.0237722f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_7 VNB A2 0.00689173f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_8 VNB N_A2_c_105_n 0.0160326f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.295
cc_9 VNB N_A_281_244#_c_141_n 0.00864087f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.46
cc_10 VNB N_A_281_244#_M1003_g 0.0268815f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.295
cc_11 VNB N_A_281_244#_c_143_n 0.01163f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_281_244#_c_144_n 0.00211765f $X=-0.19 $Y=-0.245 $X2=0.337
+ $Y2=1.665
cc_13 VNB N_A_281_244#_c_145_n 0.00647567f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_281_244#_c_146_n 0.0367177f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_281_244#_c_147_n 0.00327435f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_281_244#_c_148_n 0.00421238f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_281_244#_c_149_n 0.0388575f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_B1_N_c_202_n 0.039745f $X=-0.19 $Y=-0.245 $X2=0.395 $Y2=1.305
cc_19 VNB N_B1_N_c_203_n 0.0229476f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.69
cc_20 VNB B1_N 0.00365732f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.46
cc_21 VNB N_A_200_392#_c_233_n 0.0355852f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.46
cc_22 VNB N_A_200_392#_M1000_g 0.0299727f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_200_392#_c_235_n 0.0176071f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_200_392#_c_236_n 0.00623122f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_200_392#_c_237_n 2.56499e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_200_392#_c_238_n 0.00393771f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_200_392#_c_239_n 0.00302585f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_VPWR_c_313_n 0.163682f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_X_c_358_n 0.0267037f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_30 VNB N_X_c_359_n 0.01394f $X=-0.19 $Y=-0.245 $X2=0.395 $Y2=1.295
cc_31 VNB N_X_c_360_n 0.024976f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_27_74#_c_384_n 0.0193497f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_33 VNB N_A_27_74#_c_385_n 0.00752814f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_27_74#_c_386_n 0.00252555f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.295
cc_35 VNB N_VGND_c_411_n 0.00970653f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_36 VNB N_VGND_c_412_n 0.0172154f $X=-0.19 $Y=-0.245 $X2=0.395 $Y2=1.295
cc_37 VNB N_VGND_c_413_n 0.0191515f $X=-0.19 $Y=-0.245 $X2=0.337 $Y2=1.295
cc_38 VNB N_VGND_c_414_n 0.0543292f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_415_n 0.0190372f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_416_n 0.24119f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_417_n 0.00632279f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_418_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VPB N_A1_c_73_n 0.025423f $X=-0.19 $Y=1.66 $X2=0.395 $Y2=1.625
cc_44 VPB N_A1_c_78_n 0.019221f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.885
cc_45 VPB A1 0.00808948f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.21
cc_46 VPB N_A2_c_106_n 0.0169988f $X=-0.19 $Y=1.66 $X2=0.395 $Y2=1.305
cc_47 VPB N_A2_c_103_n 0.020226f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.21
cc_48 VPB A2 0.00506394f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_49 VPB N_A_281_244#_c_141_n 0.00778925f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.46
cc_50 VPB N_A_281_244#_c_151_n 0.0248446f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.21
cc_51 VPB N_A_281_244#_c_144_n 0.00414995f $X=-0.19 $Y=1.66 $X2=0.337 $Y2=1.665
cc_52 VPB N_A_281_244#_c_153_n 0.00946383f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_53 VPB N_A_281_244#_c_154_n 0.00913392f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_54 VPB N_B1_N_c_202_n 0.0289087f $X=-0.19 $Y=1.66 $X2=0.395 $Y2=1.305
cc_55 VPB N_A_200_392#_c_233_n 0.0294154f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.46
cc_56 VPB N_A_200_392#_c_236_n 0.00611446f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_57 VPB N_A_200_392#_c_242_n 0.0169246f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_58 VPB N_A_200_392#_c_237_n 0.00320286f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_59 VPB N_A_200_392#_c_244_n 0.00332091f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_60 VPB N_VPWR_c_314_n 0.0120106f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_61 VPB N_VPWR_c_315_n 0.0481714f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_62 VPB N_VPWR_c_316_n 0.021665f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_63 VPB N_VPWR_c_317_n 0.0203522f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_64 VPB N_VPWR_c_318_n 0.0323805f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_65 VPB N_VPWR_c_319_n 0.0320766f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_66 VPB N_VPWR_c_320_n 0.0189171f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_67 VPB N_VPWR_c_313_n 0.0785599f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_68 VPB N_VPWR_c_322_n 0.00614127f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_69 VPB N_VPWR_c_323_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_70 VPB X 0.0138434f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.295
cc_71 VPB X 0.041687f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_72 VPB N_X_c_360_n 0.0075617f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_73 N_A1_c_78_n N_A2_c_106_n 0.0531395f $X=0.505 $Y=1.885 $X2=-0.19 $Y2=-0.245
cc_74 N_A1_c_76_n N_A2_c_102_n 0.0218539f $X=0.395 $Y=1.13 $X2=0 $Y2=0
cc_75 N_A1_c_73_n N_A2_c_103_n 0.0202485f $X=0.395 $Y=1.625 $X2=0 $Y2=0
cc_76 A1 A2 0.0348017f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_77 N_A1_c_75_n A2 0.00260358f $X=0.385 $Y=1.295 $X2=0 $Y2=0
cc_78 A1 N_A2_c_105_n 0.00246986f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_79 N_A1_c_75_n N_A2_c_105_n 0.0154493f $X=0.385 $Y=1.295 $X2=0 $Y2=0
cc_80 N_A1_c_73_n N_VPWR_c_315_n 0.00139936f $X=0.395 $Y=1.625 $X2=0 $Y2=0
cc_81 N_A1_c_78_n N_VPWR_c_315_n 0.0231372f $X=0.505 $Y=1.885 $X2=0 $Y2=0
cc_82 A1 N_VPWR_c_315_n 0.0255544f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_83 N_A1_c_78_n N_VPWR_c_318_n 0.00413917f $X=0.505 $Y=1.885 $X2=0 $Y2=0
cc_84 N_A1_c_78_n N_VPWR_c_313_n 0.00817532f $X=0.505 $Y=1.885 $X2=0 $Y2=0
cc_85 N_A1_c_76_n N_A_27_74#_c_384_n 0.00684796f $X=0.395 $Y=1.13 $X2=0 $Y2=0
cc_86 A1 N_A_27_74#_c_388_n 0.00787831f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_87 N_A1_c_76_n N_A_27_74#_c_388_n 0.00967287f $X=0.395 $Y=1.13 $X2=0 $Y2=0
cc_88 A1 N_A_27_74#_c_385_n 0.0254243f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_89 N_A1_c_75_n N_A_27_74#_c_385_n 0.00137692f $X=0.385 $Y=1.295 $X2=0 $Y2=0
cc_90 N_A1_c_76_n N_A_27_74#_c_385_n 7.15033e-19 $X=0.395 $Y=1.13 $X2=0 $Y2=0
cc_91 N_A1_c_76_n N_A_27_74#_c_386_n 5.85113e-19 $X=0.395 $Y=1.13 $X2=0 $Y2=0
cc_92 N_A1_c_76_n N_VGND_c_411_n 0.00488987f $X=0.395 $Y=1.13 $X2=0 $Y2=0
cc_93 N_A1_c_76_n N_VGND_c_413_n 0.00434272f $X=0.395 $Y=1.13 $X2=0 $Y2=0
cc_94 N_A1_c_76_n N_VGND_c_416_n 0.00439339f $X=0.395 $Y=1.13 $X2=0 $Y2=0
cc_95 N_A2_c_103_n N_A_281_244#_c_141_n 0.0151949f $X=1 $Y=1.635 $X2=0 $Y2=0
cc_96 N_A2_c_106_n N_A_281_244#_c_151_n 0.0268274f $X=0.925 $Y=1.885 $X2=0 $Y2=0
cc_97 N_A2_c_103_n N_A_281_244#_c_151_n 0.00289334f $X=1 $Y=1.635 $X2=0 $Y2=0
cc_98 N_A2_c_102_n N_A_281_244#_M1003_g 0.0109162f $X=1 $Y=1.13 $X2=0 $Y2=0
cc_99 A2 N_A_281_244#_M1003_g 7.79834e-19 $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_100 N_A2_c_105_n N_A_281_244#_M1003_g 0.00380119f $X=1 $Y=1.295 $X2=0 $Y2=0
cc_101 A2 N_A_281_244#_c_143_n 0.00560366f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_102 N_A2_c_105_n N_A_281_244#_c_143_n 0.0151949f $X=1 $Y=1.295 $X2=0 $Y2=0
cc_103 A2 N_A_200_392#_c_236_n 0.0357245f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_104 N_A2_c_105_n N_A_200_392#_c_236_n 2.2434e-19 $X=1 $Y=1.295 $X2=0 $Y2=0
cc_105 N_A2_c_106_n N_A_200_392#_c_244_n 0.00309874f $X=0.925 $Y=1.885 $X2=0
+ $Y2=0
cc_106 N_A2_c_103_n N_A_200_392#_c_248_n 8.29952e-19 $X=1 $Y=1.635 $X2=0 $Y2=0
cc_107 A2 N_A_200_392#_c_248_n 0.0226372f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_108 N_A2_c_106_n N_VPWR_c_315_n 0.0035452f $X=0.925 $Y=1.885 $X2=0 $Y2=0
cc_109 N_A2_c_106_n N_VPWR_c_316_n 5.64735e-19 $X=0.925 $Y=1.885 $X2=0 $Y2=0
cc_110 N_A2_c_106_n N_VPWR_c_318_n 0.00461464f $X=0.925 $Y=1.885 $X2=0 $Y2=0
cc_111 N_A2_c_106_n N_VPWR_c_313_n 0.00910574f $X=0.925 $Y=1.885 $X2=0 $Y2=0
cc_112 N_A2_c_102_n N_A_27_74#_c_384_n 5.85113e-19 $X=1 $Y=1.13 $X2=0 $Y2=0
cc_113 N_A2_c_102_n N_A_27_74#_c_388_n 0.00974567f $X=1 $Y=1.13 $X2=0 $Y2=0
cc_114 A2 N_A_27_74#_c_388_n 0.0347531f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_115 N_A2_c_105_n N_A_27_74#_c_388_n 9.46749e-19 $X=1 $Y=1.295 $X2=0 $Y2=0
cc_116 N_A2_c_102_n N_A_27_74#_c_386_n 0.00669591f $X=1 $Y=1.13 $X2=0 $Y2=0
cc_117 N_A2_c_102_n N_VGND_c_411_n 0.00488987f $X=1 $Y=1.13 $X2=0 $Y2=0
cc_118 N_A2_c_102_n N_VGND_c_414_n 0.00434272f $X=1 $Y=1.13 $X2=0 $Y2=0
cc_119 N_A2_c_102_n N_VGND_c_416_n 0.00435917f $X=1 $Y=1.13 $X2=0 $Y2=0
cc_120 N_A_281_244#_c_144_n N_B1_N_c_202_n 0.00829829f $X=2.14 $Y=1.82 $X2=-0.19
+ $Y2=-0.245
cc_121 N_A_281_244#_c_145_n N_B1_N_c_202_n 0.00114872f $X=2.14 $Y=1.385
+ $X2=-0.19 $Y2=-0.245
cc_122 N_A_281_244#_c_146_n N_B1_N_c_202_n 0.0212168f $X=2.14 $Y=1.385 $X2=-0.19
+ $Y2=-0.245
cc_123 N_A_281_244#_c_154_n N_B1_N_c_202_n 0.00701349f $X=2.52 $Y=1.985
+ $X2=-0.19 $Y2=-0.245
cc_124 N_A_281_244#_c_148_n N_B1_N_c_202_n 0.00105159f $X=2.555 $Y=0.845
+ $X2=-0.19 $Y2=-0.245
cc_125 N_A_281_244#_c_147_n N_B1_N_c_203_n 0.00438837f $X=2.14 $Y=1.22 $X2=0
+ $Y2=0
cc_126 N_A_281_244#_c_148_n N_B1_N_c_203_n 0.00422447f $X=2.555 $Y=0.845 $X2=0
+ $Y2=0
cc_127 N_A_281_244#_c_146_n B1_N 0.00131019f $X=2.14 $Y=1.385 $X2=0 $Y2=0
cc_128 N_A_281_244#_c_154_n B1_N 0.0098063f $X=2.52 $Y=1.985 $X2=0 $Y2=0
cc_129 N_A_281_244#_c_147_n B1_N 0.0235839f $X=2.14 $Y=1.22 $X2=0 $Y2=0
cc_130 N_A_281_244#_c_148_n B1_N 0.0143996f $X=2.555 $Y=0.845 $X2=0 $Y2=0
cc_131 N_A_281_244#_M1003_g N_A_200_392#_c_235_n 0.00745905f $X=1.51 $Y=0.69
+ $X2=0 $Y2=0
cc_132 N_A_281_244#_c_148_n N_A_200_392#_c_235_n 0.0264642f $X=2.555 $Y=0.845
+ $X2=0 $Y2=0
cc_133 N_A_281_244#_c_141_n N_A_200_392#_c_236_n 0.0102224f $X=1.495 $Y=1.795
+ $X2=0 $Y2=0
cc_134 N_A_281_244#_c_151_n N_A_200_392#_c_236_n 0.00309755f $X=1.495 $Y=1.885
+ $X2=0 $Y2=0
cc_135 N_A_281_244#_c_145_n N_A_200_392#_c_236_n 0.0414317f $X=2.14 $Y=1.385
+ $X2=0 $Y2=0
cc_136 N_A_281_244#_c_146_n N_A_200_392#_c_236_n 2.99159e-19 $X=2.14 $Y=1.385
+ $X2=0 $Y2=0
cc_137 N_A_281_244#_c_153_n N_A_200_392#_c_236_n 0.0117447f $X=2.305 $Y=1.985
+ $X2=0 $Y2=0
cc_138 N_A_281_244#_c_147_n N_A_200_392#_c_236_n 0.00863714f $X=2.14 $Y=1.22
+ $X2=0 $Y2=0
cc_139 N_A_281_244#_c_149_n N_A_200_392#_c_236_n 0.0203485f $X=1.975 $Y=1.385
+ $X2=0 $Y2=0
cc_140 N_A_281_244#_M1001_s N_A_200_392#_c_242_n 0.011395f $X=2.305 $Y=1.84
+ $X2=0 $Y2=0
cc_141 N_A_281_244#_c_153_n N_A_200_392#_c_242_n 0.0277408f $X=2.305 $Y=1.985
+ $X2=0 $Y2=0
cc_142 N_A_281_244#_c_154_n N_A_200_392#_c_242_n 0.0249136f $X=2.52 $Y=1.985
+ $X2=0 $Y2=0
cc_143 N_A_281_244#_c_154_n N_A_200_392#_c_237_n 0.014348f $X=2.52 $Y=1.985
+ $X2=0 $Y2=0
cc_144 N_A_281_244#_c_151_n N_A_200_392#_c_244_n 0.003101f $X=1.495 $Y=1.885
+ $X2=0 $Y2=0
cc_145 N_A_281_244#_c_151_n N_A_200_392#_c_248_n 0.0365676f $X=1.495 $Y=1.885
+ $X2=0 $Y2=0
cc_146 N_A_281_244#_c_153_n N_A_200_392#_c_248_n 0.0152282f $X=2.305 $Y=1.985
+ $X2=0 $Y2=0
cc_147 N_A_281_244#_c_149_n N_A_200_392#_c_248_n 4.14132e-19 $X=1.975 $Y=1.385
+ $X2=0 $Y2=0
cc_148 N_A_281_244#_c_147_n N_A_200_392#_c_238_n 0.00146638f $X=2.14 $Y=1.22
+ $X2=0 $Y2=0
cc_149 N_A_281_244#_c_149_n N_A_200_392#_c_238_n 0.00677504f $X=1.975 $Y=1.385
+ $X2=0 $Y2=0
cc_150 N_A_281_244#_c_151_n N_VPWR_c_316_n 0.00835607f $X=1.495 $Y=1.885 $X2=0
+ $Y2=0
cc_151 N_A_281_244#_c_151_n N_VPWR_c_318_n 0.00413917f $X=1.495 $Y=1.885 $X2=0
+ $Y2=0
cc_152 N_A_281_244#_c_151_n N_VPWR_c_313_n 0.0041556f $X=1.495 $Y=1.885 $X2=0
+ $Y2=0
cc_153 N_A_281_244#_M1003_g N_A_27_74#_c_388_n 0.00205241f $X=1.51 $Y=0.69 $X2=0
+ $Y2=0
cc_154 N_A_281_244#_M1003_g N_A_27_74#_c_386_n 0.00454372f $X=1.51 $Y=0.69 $X2=0
+ $Y2=0
cc_155 N_A_281_244#_M1003_g N_VGND_c_414_n 0.00451267f $X=1.51 $Y=0.69 $X2=0
+ $Y2=0
cc_156 N_A_281_244#_c_148_n N_VGND_c_414_n 0.00927306f $X=2.555 $Y=0.845 $X2=0
+ $Y2=0
cc_157 N_A_281_244#_M1003_g N_VGND_c_416_n 0.00881535f $X=1.51 $Y=0.69 $X2=0
+ $Y2=0
cc_158 N_A_281_244#_c_148_n N_VGND_c_416_n 0.0165534f $X=2.555 $Y=0.845 $X2=0
+ $Y2=0
cc_159 N_B1_N_c_202_n N_A_200_392#_c_233_n 0.0412109f $X=2.75 $Y=1.765 $X2=0
+ $Y2=0
cc_160 B1_N N_A_200_392#_c_233_n 2.75885e-19 $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_161 N_B1_N_c_203_n N_A_200_392#_M1000_g 0.0181853f $X=2.77 $Y=1.22 $X2=0
+ $Y2=0
cc_162 B1_N N_A_200_392#_M1000_g 7.87159e-19 $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_163 N_B1_N_c_202_n N_A_200_392#_c_242_n 0.0183847f $X=2.75 $Y=1.765 $X2=0
+ $Y2=0
cc_164 N_B1_N_c_202_n N_A_200_392#_c_237_n 0.00977421f $X=2.75 $Y=1.765 $X2=0
+ $Y2=0
cc_165 N_B1_N_c_202_n N_A_200_392#_c_239_n 0.00363632f $X=2.75 $Y=1.765 $X2=0
+ $Y2=0
cc_166 B1_N N_A_200_392#_c_239_n 0.0156452f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_167 N_B1_N_c_202_n N_VPWR_c_317_n 0.00427039f $X=2.75 $Y=1.765 $X2=0 $Y2=0
cc_168 N_B1_N_c_202_n N_VPWR_c_319_n 0.00402388f $X=2.75 $Y=1.765 $X2=0 $Y2=0
cc_169 N_B1_N_c_202_n N_VPWR_c_313_n 0.00462577f $X=2.75 $Y=1.765 $X2=0 $Y2=0
cc_170 N_B1_N_c_203_n N_X_c_358_n 6.61818e-19 $X=2.77 $Y=1.22 $X2=0 $Y2=0
cc_171 N_B1_N_c_202_n X 8.93994e-19 $X=2.75 $Y=1.765 $X2=0 $Y2=0
cc_172 N_B1_N_c_203_n N_VGND_c_412_n 0.00650911f $X=2.77 $Y=1.22 $X2=0 $Y2=0
cc_173 N_B1_N_c_203_n N_VGND_c_414_n 0.00434489f $X=2.77 $Y=1.22 $X2=0 $Y2=0
cc_174 N_B1_N_c_203_n N_VGND_c_416_n 0.00487769f $X=2.77 $Y=1.22 $X2=0 $Y2=0
cc_175 N_A_200_392#_c_236_n N_VPWR_M1006_d 5.94494e-19 $X=1.7 $Y=1.97 $X2=0
+ $Y2=0
cc_176 N_A_200_392#_c_242_n N_VPWR_M1006_d 0.0045773f $X=3.055 $Y=2.405 $X2=0
+ $Y2=0
cc_177 N_A_200_392#_c_248_n N_VPWR_M1006_d 0.0128722f $X=1.785 $Y=2.23 $X2=0
+ $Y2=0
cc_178 N_A_200_392#_c_242_n N_VPWR_M1001_d 0.0119539f $X=3.055 $Y=2.405 $X2=0
+ $Y2=0
cc_179 N_A_200_392#_c_237_n N_VPWR_M1001_d 0.00958635f $X=3.14 $Y=2.32 $X2=0
+ $Y2=0
cc_180 N_A_200_392#_c_244_n N_VPWR_c_315_n 0.00669492f $X=1.22 $Y=2.135 $X2=0
+ $Y2=0
cc_181 N_A_200_392#_c_244_n N_VPWR_c_316_n 0.0127976f $X=1.22 $Y=2.135 $X2=0
+ $Y2=0
cc_182 N_A_200_392#_c_248_n N_VPWR_c_316_n 0.0225152f $X=1.785 $Y=2.23 $X2=0
+ $Y2=0
cc_183 N_A_200_392#_c_233_n N_VPWR_c_317_n 0.00904313f $X=3.335 $Y=1.765 $X2=0
+ $Y2=0
cc_184 N_A_200_392#_c_242_n N_VPWR_c_317_n 0.0255974f $X=3.055 $Y=2.405 $X2=0
+ $Y2=0
cc_185 N_A_200_392#_c_244_n N_VPWR_c_318_n 0.0142934f $X=1.22 $Y=2.135 $X2=0
+ $Y2=0
cc_186 N_A_200_392#_c_233_n N_VPWR_c_320_n 0.00445602f $X=3.335 $Y=1.765 $X2=0
+ $Y2=0
cc_187 N_A_200_392#_c_233_n N_VPWR_c_313_n 0.00865213f $X=3.335 $Y=1.765 $X2=0
+ $Y2=0
cc_188 N_A_200_392#_c_242_n N_VPWR_c_313_n 0.0355705f $X=3.055 $Y=2.405 $X2=0
+ $Y2=0
cc_189 N_A_200_392#_c_244_n N_VPWR_c_313_n 0.0119825f $X=1.22 $Y=2.135 $X2=0
+ $Y2=0
cc_190 N_A_200_392#_c_248_n N_VPWR_c_313_n 0.00670731f $X=1.785 $Y=2.23 $X2=0
+ $Y2=0
cc_191 N_A_200_392#_M1000_g N_X_c_358_n 0.00806387f $X=3.34 $Y=0.74 $X2=0 $Y2=0
cc_192 N_A_200_392#_c_233_n N_X_c_359_n 4.48913e-19 $X=3.335 $Y=1.765 $X2=0
+ $Y2=0
cc_193 N_A_200_392#_M1000_g N_X_c_359_n 0.00386394f $X=3.34 $Y=0.74 $X2=0 $Y2=0
cc_194 N_A_200_392#_c_239_n N_X_c_359_n 0.00175157f $X=3.25 $Y=1.485 $X2=0 $Y2=0
cc_195 N_A_200_392#_c_233_n X 0.00301202f $X=3.335 $Y=1.765 $X2=0 $Y2=0
cc_196 N_A_200_392#_c_237_n X 0.0196895f $X=3.14 $Y=2.32 $X2=0 $Y2=0
cc_197 N_A_200_392#_c_239_n X 0.00153915f $X=3.25 $Y=1.485 $X2=0 $Y2=0
cc_198 N_A_200_392#_c_233_n X 0.0128211f $X=3.335 $Y=1.765 $X2=0 $Y2=0
cc_199 N_A_200_392#_c_233_n N_X_c_360_n 0.0101986f $X=3.335 $Y=1.765 $X2=0 $Y2=0
cc_200 N_A_200_392#_M1000_g N_X_c_360_n 0.00477624f $X=3.34 $Y=0.74 $X2=0 $Y2=0
cc_201 N_A_200_392#_c_237_n N_X_c_360_n 0.00535848f $X=3.14 $Y=2.32 $X2=0 $Y2=0
cc_202 N_A_200_392#_c_239_n N_X_c_360_n 0.0249376f $X=3.25 $Y=1.485 $X2=0 $Y2=0
cc_203 N_A_200_392#_c_235_n N_A_27_74#_c_386_n 0.0172628f $X=1.78 $Y=0.515 $X2=0
+ $Y2=0
cc_204 N_A_200_392#_c_233_n N_VGND_c_412_n 0.00283306f $X=3.335 $Y=1.765 $X2=0
+ $Y2=0
cc_205 N_A_200_392#_M1000_g N_VGND_c_412_n 0.00703428f $X=3.34 $Y=0.74 $X2=0
+ $Y2=0
cc_206 N_A_200_392#_c_239_n N_VGND_c_412_n 0.00834888f $X=3.25 $Y=1.485 $X2=0
+ $Y2=0
cc_207 N_A_200_392#_c_235_n N_VGND_c_414_n 0.0146357f $X=1.78 $Y=0.515 $X2=0
+ $Y2=0
cc_208 N_A_200_392#_M1000_g N_VGND_c_415_n 0.00434272f $X=3.34 $Y=0.74 $X2=0
+ $Y2=0
cc_209 N_A_200_392#_M1000_g N_VGND_c_416_n 0.00828734f $X=3.34 $Y=0.74 $X2=0
+ $Y2=0
cc_210 N_A_200_392#_c_235_n N_VGND_c_416_n 0.0121141f $X=1.78 $Y=0.515 $X2=0
+ $Y2=0
cc_211 N_VPWR_c_317_n X 0.0129586f $X=3.06 $Y=2.78 $X2=0 $Y2=0
cc_212 N_VPWR_c_320_n X 0.0159324f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_213 N_VPWR_c_313_n X 0.0131546f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_214 N_X_c_358_n N_VGND_c_412_n 0.0259022f $X=3.555 $Y=0.515 $X2=0 $Y2=0
cc_215 N_X_c_358_n N_VGND_c_415_n 0.0161257f $X=3.555 $Y=0.515 $X2=0 $Y2=0
cc_216 N_X_c_358_n N_VGND_c_416_n 0.013291f $X=3.555 $Y=0.515 $X2=0 $Y2=0
cc_217 N_A_27_74#_c_388_n N_VGND_M1008_d 0.0125077f $X=1.115 $Y=0.875 $X2=-0.19
+ $Y2=-0.245
cc_218 N_A_27_74#_c_384_n N_VGND_c_411_n 0.0109215f $X=0.28 $Y=0.515 $X2=0 $Y2=0
cc_219 N_A_27_74#_c_388_n N_VGND_c_411_n 0.0243105f $X=1.115 $Y=0.875 $X2=0
+ $Y2=0
cc_220 N_A_27_74#_c_386_n N_VGND_c_411_n 0.0109215f $X=1.28 $Y=0.515 $X2=0 $Y2=0
cc_221 N_A_27_74#_c_384_n N_VGND_c_413_n 0.0144497f $X=0.28 $Y=0.515 $X2=0 $Y2=0
cc_222 N_A_27_74#_c_386_n N_VGND_c_414_n 0.0144232f $X=1.28 $Y=0.515 $X2=0 $Y2=0
cc_223 N_A_27_74#_c_384_n N_VGND_c_416_n 0.0119539f $X=0.28 $Y=0.515 $X2=0 $Y2=0
cc_224 N_A_27_74#_c_388_n N_VGND_c_416_n 0.0116461f $X=1.115 $Y=0.875 $X2=0
+ $Y2=0
cc_225 N_A_27_74#_c_386_n N_VGND_c_416_n 0.0119105f $X=1.28 $Y=0.515 $X2=0 $Y2=0
