* File: sky130_fd_sc_hs__a32o_1.spice
* Created: Tue Sep  1 19:53:24 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hs__a32o_1.pex.spice"
.subckt sky130_fd_sc_hs__a32o_1  VNB VPB A3 A2 A1 B1 B2 X VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* X	X
* B2	B2
* B1	B1
* A1	A1
* A2	A2
* A3	A3
* VPB	VPB
* VNB	VNB
MM1010 N_VGND_M1010_d N_A_84_48#_M1010_g N_X_M1010_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.224145 AS=0.2109 PD=1.41029 PS=2.05 NRD=22.692 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75002.7 A=0.111 P=1.78 MULT=1
MM1006 A_259_94# N_A3_M1006_g N_VGND_M1010_d VNB NLOWVT L=0.15 W=0.64 AD=0.0768
+ AS=0.193855 PD=0.88 PS=1.21971 NRD=12.18 NRS=29.988 M=1 R=4.26667 SA=75000.9
+ SB=75002.3 A=0.096 P=1.58 MULT=1
MM1007 A_337_94# N_A2_M1007_g A_259_94# VNB NLOWVT L=0.15 W=0.64 AD=0.1248
+ AS=0.0768 PD=1.03 PS=0.88 NRD=26.244 NRS=12.18 M=1 R=4.26667 SA=75001.3
+ SB=75001.9 A=0.096 P=1.58 MULT=1
MM1011 N_A_84_48#_M1011_d N_A1_M1011_g A_337_94# VNB NLOWVT L=0.15 W=0.64
+ AD=0.2016 AS=0.1248 PD=1.27 PS=1.03 NRD=0 NRS=26.244 M=1 R=4.26667 SA=75001.9
+ SB=75001.4 A=0.096 P=1.58 MULT=1
MM1001 A_601_94# N_B1_M1001_g N_A_84_48#_M1011_d VNB NLOWVT L=0.15 W=0.64
+ AD=0.0768 AS=0.2016 PD=0.88 PS=1.27 NRD=12.18 NRS=0 M=1 R=4.26667 SA=75002.6
+ SB=75000.6 A=0.096 P=1.58 MULT=1
MM1009 N_VGND_M1009_d N_B2_M1009_g A_601_94# VNB NLOWVT L=0.15 W=0.64 AD=0.1824
+ AS=0.0768 PD=1.85 PS=0.88 NRD=0 NRS=12.18 M=1 R=4.26667 SA=75003 SB=75000.2
+ A=0.096 P=1.58 MULT=1
MM1000 N_VPWR_M1000_d N_A_84_48#_M1000_g N_X_M1000_s VPB PSHORT L=0.15 W=1.12
+ AD=0.275457 AS=0.3304 PD=1.69057 PS=2.83 NRD=15.8191 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75002.7 A=0.168 P=2.54 MULT=1
MM1002 N_A_244_368#_M1002_d N_A3_M1002_g N_VPWR_M1000_d VPB PSHORT L=0.15 W=1
+ AD=0.15 AS=0.245943 PD=1.3 PS=1.50943 NRD=1.9503 NRS=22.1625 M=1 R=6.66667
+ SA=75000.8 SB=75002.4 A=0.15 P=2.3 MULT=1
MM1004 N_VPWR_M1004_d N_A2_M1004_g N_A_244_368#_M1002_d VPB PSHORT L=0.15 W=1
+ AD=0.295 AS=0.15 PD=1.59 PS=1.3 NRD=30.535 NRS=1.9503 M=1 R=6.66667 SA=75001.3
+ SB=75002 A=0.15 P=2.3 MULT=1
MM1005 N_A_244_368#_M1005_d N_A1_M1005_g N_VPWR_M1004_d VPB PSHORT L=0.15 W=1
+ AD=0.15 AS=0.295 PD=1.3 PS=1.59 NRD=1.9503 NRS=30.535 M=1 R=6.66667 SA=75002
+ SB=75001.2 A=0.15 P=2.3 MULT=1
MM1008 N_A_84_48#_M1008_d N_B1_M1008_g N_A_244_368#_M1005_d VPB PSHORT L=0.15
+ W=1 AD=0.2 AS=0.15 PD=1.4 PS=1.3 NRD=11.8003 NRS=1.9503 M=1 R=6.66667
+ SA=75002.5 SB=75000.8 A=0.15 P=2.3 MULT=1
MM1003 N_A_244_368#_M1003_d N_B2_M1003_g N_A_84_48#_M1008_d VPB PSHORT L=0.15
+ W=1 AD=0.295 AS=0.2 PD=2.59 PS=1.4 NRD=1.9503 NRS=11.8003 M=1 R=6.66667
+ SA=75003 SB=75000.2 A=0.15 P=2.3 MULT=1
DX12_noxref VNB VPB NWDIODE A=7.8492 P=12.16
*
.include "sky130_fd_sc_hs__a32o_1.pxi.spice"
*
.ends
*
*
