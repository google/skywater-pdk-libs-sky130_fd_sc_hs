# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_hs__sedfxtp_4
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_hs__sedfxtp_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  16.80000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425000 0.980000 0.825000 1.990000 ;
    END
  END D
  PIN DE
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.535000 1.320000 1.865000 1.780000 ;
    END
  END DE
  PIN Q
    ANTENNADIFFAREA  1.097500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 15.065000 1.820000 16.675000 2.150000 ;
        RECT 15.065000 2.150000 15.285000 2.980000 ;
        RECT 15.075000 0.560000 15.325000 1.090000 ;
        RECT 15.075000 1.090000 16.675000 1.340000 ;
        RECT 15.165000 1.340000 16.675000 1.820000 ;
        RECT 15.970000 2.150000 16.185000 2.980000 ;
        RECT 15.995000 0.575000 16.200000 1.090000 ;
    END
  END Q
  PIN SCD
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.955000 1.180000 5.370000 1.745000 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.445000 1.180000 4.785000 1.510000 ;
    END
  END SCE
  PIN CLK
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 6.455000 1.180000 7.075000 1.550000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT  0.000000 -0.085000 16.800000 0.085000 ;
        RECT  1.040000  0.085000  1.370000 0.810000 ;
        RECT  2.030000  0.085000  2.360000 1.005000 ;
        RECT  4.765000  0.085000  5.095000 1.010000 ;
        RECT  6.110000  0.085000  6.360000 0.905000 ;
        RECT  7.095000  0.085000  7.425000 0.670000 ;
        RECT  9.840000  0.085000 10.090000 0.690000 ;
        RECT 11.280000  0.085000 11.530000 0.690000 ;
        RECT 12.855000  0.085000 13.835000 0.680000 ;
        RECT 14.565000  0.085000 14.895000 1.340000 ;
        RECT 15.495000  0.085000 15.825000 0.920000 ;
        RECT 16.370000  0.085000 16.700000 0.920000 ;
      LAYER mcon ;
        RECT  0.155000 -0.085000  0.325000 0.085000 ;
        RECT  0.635000 -0.085000  0.805000 0.085000 ;
        RECT  1.115000 -0.085000  1.285000 0.085000 ;
        RECT  1.595000 -0.085000  1.765000 0.085000 ;
        RECT  2.075000 -0.085000  2.245000 0.085000 ;
        RECT  2.555000 -0.085000  2.725000 0.085000 ;
        RECT  3.035000 -0.085000  3.205000 0.085000 ;
        RECT  3.515000 -0.085000  3.685000 0.085000 ;
        RECT  3.995000 -0.085000  4.165000 0.085000 ;
        RECT  4.475000 -0.085000  4.645000 0.085000 ;
        RECT  4.955000 -0.085000  5.125000 0.085000 ;
        RECT  5.435000 -0.085000  5.605000 0.085000 ;
        RECT  5.915000 -0.085000  6.085000 0.085000 ;
        RECT  6.395000 -0.085000  6.565000 0.085000 ;
        RECT  6.875000 -0.085000  7.045000 0.085000 ;
        RECT  7.355000 -0.085000  7.525000 0.085000 ;
        RECT  7.835000 -0.085000  8.005000 0.085000 ;
        RECT  8.315000 -0.085000  8.485000 0.085000 ;
        RECT  8.795000 -0.085000  8.965000 0.085000 ;
        RECT  9.275000 -0.085000  9.445000 0.085000 ;
        RECT  9.755000 -0.085000  9.925000 0.085000 ;
        RECT 10.235000 -0.085000 10.405000 0.085000 ;
        RECT 10.715000 -0.085000 10.885000 0.085000 ;
        RECT 11.195000 -0.085000 11.365000 0.085000 ;
        RECT 11.675000 -0.085000 11.845000 0.085000 ;
        RECT 12.155000 -0.085000 12.325000 0.085000 ;
        RECT 12.635000 -0.085000 12.805000 0.085000 ;
        RECT 13.115000 -0.085000 13.285000 0.085000 ;
        RECT 13.595000 -0.085000 13.765000 0.085000 ;
        RECT 14.075000 -0.085000 14.245000 0.085000 ;
        RECT 14.555000 -0.085000 14.725000 0.085000 ;
        RECT 15.035000 -0.085000 15.205000 0.085000 ;
        RECT 15.515000 -0.085000 15.685000 0.085000 ;
        RECT 15.995000 -0.085000 16.165000 0.085000 ;
        RECT 16.475000 -0.085000 16.645000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.245000 16.800000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT  0.000000 3.245000 16.800000 3.415000 ;
        RECT  1.035000 2.630000  1.285000 3.245000 ;
        RECT  2.475000 2.630000  2.725000 3.245000 ;
        RECT  4.970000 2.595000  5.220000 3.245000 ;
        RECT  6.260000 2.675000  6.590000 3.245000 ;
        RECT  7.610000 2.675000  7.940000 3.245000 ;
        RECT  9.960000 2.730000 10.290000 3.245000 ;
        RECT 10.995000 2.730000 11.325000 3.245000 ;
        RECT 13.335000 2.650000 13.875000 3.245000 ;
        RECT 14.565000 1.950000 14.895000 3.245000 ;
        RECT 15.465000 2.320000 15.795000 3.245000 ;
        RECT 16.365000 2.320000 16.695000 3.245000 ;
      LAYER mcon ;
        RECT  0.155000 3.245000  0.325000 3.415000 ;
        RECT  0.635000 3.245000  0.805000 3.415000 ;
        RECT  1.115000 3.245000  1.285000 3.415000 ;
        RECT  1.595000 3.245000  1.765000 3.415000 ;
        RECT  2.075000 3.245000  2.245000 3.415000 ;
        RECT  2.555000 3.245000  2.725000 3.415000 ;
        RECT  3.035000 3.245000  3.205000 3.415000 ;
        RECT  3.515000 3.245000  3.685000 3.415000 ;
        RECT  3.995000 3.245000  4.165000 3.415000 ;
        RECT  4.475000 3.245000  4.645000 3.415000 ;
        RECT  4.955000 3.245000  5.125000 3.415000 ;
        RECT  5.435000 3.245000  5.605000 3.415000 ;
        RECT  5.915000 3.245000  6.085000 3.415000 ;
        RECT  6.395000 3.245000  6.565000 3.415000 ;
        RECT  6.875000 3.245000  7.045000 3.415000 ;
        RECT  7.355000 3.245000  7.525000 3.415000 ;
        RECT  7.835000 3.245000  8.005000 3.415000 ;
        RECT  8.315000 3.245000  8.485000 3.415000 ;
        RECT  8.795000 3.245000  8.965000 3.415000 ;
        RECT  9.275000 3.245000  9.445000 3.415000 ;
        RECT  9.755000 3.245000  9.925000 3.415000 ;
        RECT 10.235000 3.245000 10.405000 3.415000 ;
        RECT 10.715000 3.245000 10.885000 3.415000 ;
        RECT 11.195000 3.245000 11.365000 3.415000 ;
        RECT 11.675000 3.245000 11.845000 3.415000 ;
        RECT 12.155000 3.245000 12.325000 3.415000 ;
        RECT 12.635000 3.245000 12.805000 3.415000 ;
        RECT 13.115000 3.245000 13.285000 3.415000 ;
        RECT 13.595000 3.245000 13.765000 3.415000 ;
        RECT 14.075000 3.245000 14.245000 3.415000 ;
        RECT 14.555000 3.245000 14.725000 3.415000 ;
        RECT 15.035000 3.245000 15.205000 3.415000 ;
        RECT 15.515000 3.245000 15.685000 3.415000 ;
        RECT 15.995000 3.245000 16.165000 3.415000 ;
        RECT 16.475000 3.245000 16.645000 3.415000 ;
      LAYER met1 ;
        RECT 0.000000 3.085000 16.800000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.085000 0.340000  0.550000 0.810000 ;
      RECT  0.085000 0.810000  0.255000 2.290000 ;
      RECT  0.085000 2.290000  1.625000 2.460000 ;
      RECT  0.085000 2.460000  0.495000 2.980000 ;
      RECT  0.995000 0.980000  1.850000 1.150000 ;
      RECT  0.995000 1.150000  1.325000 1.950000 ;
      RECT  0.995000 1.950000  2.365000 2.120000 ;
      RECT  1.455000 2.460000  1.625000 2.905000 ;
      RECT  1.455000 2.905000  2.305000 3.075000 ;
      RECT  1.600000 0.545000  1.850000 0.980000 ;
      RECT  1.795000 2.120000  1.965000 2.735000 ;
      RECT  2.115000 1.520000  2.365000 1.950000 ;
      RECT  2.135000 2.290000  3.485000 2.460000 ;
      RECT  2.135000 2.460000  2.305000 2.905000 ;
      RECT  2.535000 1.520000  3.055000 1.850000 ;
      RECT  2.850000 0.545000  3.180000 1.175000 ;
      RECT  2.850000 1.175000  3.485000 1.345000 ;
      RECT  3.235000 2.460000  3.485000 2.975000 ;
      RECT  3.315000 1.345000  3.485000 2.290000 ;
      RECT  3.350000 0.675000  3.825000 1.005000 ;
      RECT  3.655000 1.005000  3.825000 2.295000 ;
      RECT  3.655000 2.295000  3.935000 2.905000 ;
      RECT  3.655000 2.905000  4.800000 3.075000 ;
      RECT  3.995000 0.255000  4.275000 0.605000 ;
      RECT  3.995000 0.605000  4.585000 1.010000 ;
      RECT  3.995000 1.010000  4.275000 1.915000 ;
      RECT  3.995000 1.915000  5.860000 2.085000 ;
      RECT  4.105000 2.085000  4.275000 2.255000 ;
      RECT  4.105000 2.255000  4.460000 2.735000 ;
      RECT  4.630000 2.255000  6.200000 2.335000 ;
      RECT  4.630000 2.335000  8.325000 2.425000 ;
      RECT  4.630000 2.425000  4.800000 2.905000 ;
      RECT  5.555000 0.605000  5.885000 1.075000 ;
      RECT  5.555000 1.075000  6.200000 1.245000 ;
      RECT  5.580000 1.415000  5.860000 1.915000 ;
      RECT  5.730000 2.425000  8.325000 2.505000 ;
      RECT  5.730000 2.505000  6.060000 2.935000 ;
      RECT  6.030000 1.245000  6.200000 2.255000 ;
      RECT  6.540000 0.350000  6.870000 0.840000 ;
      RECT  6.540000 0.840000  7.415000 1.010000 ;
      RECT  6.710000 1.785000  7.490000 2.165000 ;
      RECT  7.245000 1.010000  7.415000 1.785000 ;
      RECT  7.605000 0.255000  9.505000 0.425000 ;
      RECT  7.605000 0.425000  7.855000 1.130000 ;
      RECT  7.720000 1.480000  8.325000 1.650000 ;
      RECT  7.720000 1.650000  7.890000 2.335000 ;
      RECT  8.060000 1.820000  8.665000 1.995000 ;
      RECT  8.060000 1.995000  8.830000 2.165000 ;
      RECT  8.075000 0.595000  8.325000 1.480000 ;
      RECT  8.155000 2.505000  8.830000 2.980000 ;
      RECT  8.495000 0.425000  8.665000 1.820000 ;
      RECT  8.495000 2.165000  8.830000 2.335000 ;
      RECT  8.835000 0.595000  9.005000 1.630000 ;
      RECT  8.835000 1.630000 10.585000 1.800000 ;
      RECT  9.000000 1.800000  9.170000 2.520000 ;
      RECT  9.000000 2.520000  9.360000 2.980000 ;
      RECT  9.175000 0.425000  9.505000 0.860000 ;
      RECT  9.175000 0.860000 10.430000 1.030000 ;
      RECT  9.175000 1.030000  9.505000 1.255000 ;
      RECT  9.340000 2.000000  9.700000 2.330000 ;
      RECT  9.530000 2.330000  9.700000 2.390000 ;
      RECT  9.530000 2.390000 12.295000 2.560000 ;
      RECT  9.715000 1.200000 11.475000 1.370000 ;
      RECT  9.715000 1.370000 10.045000 1.405000 ;
      RECT 10.255000 1.540000 10.585000 1.630000 ;
      RECT 10.260000 0.255000 11.110000 0.425000 ;
      RECT 10.260000 0.425000 10.430000 0.860000 ;
      RECT 10.475000 1.970000 10.925000 2.220000 ;
      RECT 10.600000 0.595000 10.770000 1.200000 ;
      RECT 10.755000 1.370000 11.475000 1.530000 ;
      RECT 10.755000 1.530000 10.925000 1.970000 ;
      RECT 10.940000 0.425000 11.110000 0.860000 ;
      RECT 10.940000 0.860000 11.855000 1.030000 ;
      RECT 11.685000 1.030000 11.855000 1.190000 ;
      RECT 11.685000 1.190000 13.095000 1.360000 ;
      RECT 11.685000 1.360000 11.955000 1.800000 ;
      RECT 12.035000 0.350000 12.365000 0.850000 ;
      RECT 12.035000 0.850000 13.435000 0.990000 ;
      RECT 12.035000 0.990000 14.055000 1.020000 ;
      RECT 12.125000 1.530000 12.555000 1.755000 ;
      RECT 12.125000 1.755000 12.295000 2.390000 ;
      RECT 12.465000 1.925000 12.895000 2.980000 ;
      RECT 12.725000 1.755000 14.055000 1.925000 ;
      RECT 12.765000 1.360000 13.095000 1.585000 ;
      RECT 13.155000 2.095000 13.485000 2.180000 ;
      RECT 13.155000 2.180000 14.395000 2.350000 ;
      RECT 13.265000 1.020000 14.055000 1.755000 ;
      RECT 13.725000 0.980000 14.055000 0.990000 ;
      RECT 13.725000 1.925000 14.055000 1.990000 ;
      RECT 14.005000 0.350000 14.395000 0.810000 ;
      RECT 14.045000 2.350000 14.395000 2.980000 ;
      RECT 14.225000 0.810000 14.395000 1.550000 ;
      RECT 14.225000 1.550000 14.755000 1.780000 ;
      RECT 14.225000 1.780000 14.395000 2.180000 ;
    LAYER mcon ;
      RECT  2.555000 1.580000  2.725000 1.750000 ;
      RECT 14.555000 1.580000 14.725000 1.750000 ;
    LAYER met1 ;
      RECT  2.495000 1.550000  2.785000 1.595000 ;
      RECT  2.495000 1.595000 14.785000 1.735000 ;
      RECT  2.495000 1.735000  2.785000 1.780000 ;
      RECT 14.495000 1.550000 14.785000 1.595000 ;
      RECT 14.495000 1.735000 14.785000 1.780000 ;
  END
END sky130_fd_sc_hs__sedfxtp_4
