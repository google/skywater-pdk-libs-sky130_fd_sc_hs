# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_hs__sdfxbp_1
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_hs__sdfxbp_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  12.48000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.085000 1.455000 1.630000 1.785000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.518900 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 10.500000 0.350000 10.915000 1.130000 ;
        RECT 10.650000 1.820000 10.915000 2.980000 ;
        RECT 10.745000 1.130000 10.915000 1.820000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.530100 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 12.035000 0.350000 12.375000 1.050000 ;
        RECT 12.045000 1.820000 12.375000 2.980000 ;
        RECT 12.155000 1.050000 12.375000 1.820000 ;
    END
  END Q_N
  PIN SCD
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.380000 1.550000 2.725000 2.150000 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425000 0.955000 2.050000 1.285000 ;
        RECT 1.565000 0.810000 2.050000 0.955000 ;
    END
  END SCE
  PIN CLK
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 3.235000 1.180000 3.685000 1.550000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT  0.000000 -0.085000 12.480000 0.085000 ;
        RECT  0.635000  0.085000  0.965000 0.730000 ;
        RECT  2.615000  0.085000  2.865000 0.810000 ;
        RECT  3.595000  0.085000  3.935000 0.670000 ;
        RECT  6.430000  0.085000  6.680000 0.520000 ;
        RECT  8.740000  0.085000  9.410000 0.810000 ;
        RECT 10.150000  0.085000 10.320000 1.130000 ;
        RECT 11.490000  0.085000 11.865000 1.020000 ;
      LAYER mcon ;
        RECT  0.155000 -0.085000  0.325000 0.085000 ;
        RECT  0.635000 -0.085000  0.805000 0.085000 ;
        RECT  1.115000 -0.085000  1.285000 0.085000 ;
        RECT  1.595000 -0.085000  1.765000 0.085000 ;
        RECT  2.075000 -0.085000  2.245000 0.085000 ;
        RECT  2.555000 -0.085000  2.725000 0.085000 ;
        RECT  3.035000 -0.085000  3.205000 0.085000 ;
        RECT  3.515000 -0.085000  3.685000 0.085000 ;
        RECT  3.995000 -0.085000  4.165000 0.085000 ;
        RECT  4.475000 -0.085000  4.645000 0.085000 ;
        RECT  4.955000 -0.085000  5.125000 0.085000 ;
        RECT  5.435000 -0.085000  5.605000 0.085000 ;
        RECT  5.915000 -0.085000  6.085000 0.085000 ;
        RECT  6.395000 -0.085000  6.565000 0.085000 ;
        RECT  6.875000 -0.085000  7.045000 0.085000 ;
        RECT  7.355000 -0.085000  7.525000 0.085000 ;
        RECT  7.835000 -0.085000  8.005000 0.085000 ;
        RECT  8.315000 -0.085000  8.485000 0.085000 ;
        RECT  8.795000 -0.085000  8.965000 0.085000 ;
        RECT  9.275000 -0.085000  9.445000 0.085000 ;
        RECT  9.755000 -0.085000  9.925000 0.085000 ;
        RECT 10.235000 -0.085000 10.405000 0.085000 ;
        RECT 10.715000 -0.085000 10.885000 0.085000 ;
        RECT 11.195000 -0.085000 11.365000 0.085000 ;
        RECT 11.675000 -0.085000 11.845000 0.085000 ;
        RECT 12.155000 -0.085000 12.325000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.245000 12.480000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT  0.000000 3.245000 12.480000 3.415000 ;
        RECT  0.700000 2.300000  1.030000 3.245000 ;
        RECT  2.560000 2.730000  3.150000 3.245000 ;
        RECT  3.830000 2.730000  4.335000 3.245000 ;
        RECT  6.450000 2.860000  6.780000 3.245000 ;
        RECT  8.860000 2.650000  9.430000 3.245000 ;
        RECT 10.120000 1.820000 10.450000 3.245000 ;
        RECT 11.540000 1.995000 11.870000 3.245000 ;
      LAYER mcon ;
        RECT  0.155000 3.245000  0.325000 3.415000 ;
        RECT  0.635000 3.245000  0.805000 3.415000 ;
        RECT  1.115000 3.245000  1.285000 3.415000 ;
        RECT  1.595000 3.245000  1.765000 3.415000 ;
        RECT  2.075000 3.245000  2.245000 3.415000 ;
        RECT  2.555000 3.245000  2.725000 3.415000 ;
        RECT  3.035000 3.245000  3.205000 3.415000 ;
        RECT  3.515000 3.245000  3.685000 3.415000 ;
        RECT  3.995000 3.245000  4.165000 3.415000 ;
        RECT  4.475000 3.245000  4.645000 3.415000 ;
        RECT  4.955000 3.245000  5.125000 3.415000 ;
        RECT  5.435000 3.245000  5.605000 3.415000 ;
        RECT  5.915000 3.245000  6.085000 3.415000 ;
        RECT  6.395000 3.245000  6.565000 3.415000 ;
        RECT  6.875000 3.245000  7.045000 3.415000 ;
        RECT  7.355000 3.245000  7.525000 3.415000 ;
        RECT  7.835000 3.245000  8.005000 3.415000 ;
        RECT  8.315000 3.245000  8.485000 3.415000 ;
        RECT  8.795000 3.245000  8.965000 3.415000 ;
        RECT  9.275000 3.245000  9.445000 3.415000 ;
        RECT  9.755000 3.245000  9.925000 3.415000 ;
        RECT 10.235000 3.245000 10.405000 3.415000 ;
        RECT 10.715000 3.245000 10.885000 3.415000 ;
        RECT 11.195000 3.245000 11.365000 3.415000 ;
        RECT 11.675000 3.245000 11.845000 3.415000 ;
        RECT 12.155000 3.245000 12.325000 3.415000 ;
      LAYER met1 ;
        RECT 0.000000 3.085000 12.480000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.085000 0.350000  0.465000 0.785000 ;
      RECT  0.085000 0.785000  0.255000 1.525000 ;
      RECT  0.085000 1.525000  0.915000 1.855000 ;
      RECT  0.085000 1.855000  0.530000 2.980000 ;
      RECT  0.745000 1.855000  0.915000 1.955000 ;
      RECT  0.745000 1.955000  2.170000 2.125000 ;
      RECT  1.455000 0.390000  2.390000 0.640000 ;
      RECT  1.570000 2.300000  1.900000 2.390000 ;
      RECT  1.570000 2.390000  4.675000 2.460000 ;
      RECT  1.570000 2.460000  5.235000 2.560000 ;
      RECT  1.570000 2.560000  1.900000 2.980000 ;
      RECT  1.840000 1.795000  2.170000 1.955000 ;
      RECT  2.220000 0.640000  2.390000 1.180000 ;
      RECT  2.220000 1.180000  3.065000 1.350000 ;
      RECT  2.895000 1.350000  3.065000 2.390000 ;
      RECT  3.035000 0.350000  3.365000 0.840000 ;
      RECT  3.035000 0.840000  4.025000 1.010000 ;
      RECT  3.270000 1.820000  4.025000 1.990000 ;
      RECT  3.270000 1.990000  3.600000 2.220000 ;
      RECT  3.855000 1.010000  4.025000 1.820000 ;
      RECT  4.195000 0.255000  6.035000 0.425000 ;
      RECT  4.195000 0.425000  4.445000 1.130000 ;
      RECT  4.195000 1.480000  4.900000 1.650000 ;
      RECT  4.195000 1.650000  4.365000 2.390000 ;
      RECT  4.505000 2.560000  5.235000 2.630000 ;
      RECT  4.535000 1.820000  5.240000 2.220000 ;
      RECT  4.650000 0.595000  4.900000 1.480000 ;
      RECT  4.910000 2.220000  5.240000 2.280000 ;
      RECT  4.985000 2.630000  5.235000 2.920000 ;
      RECT  5.070000 0.425000  5.240000 1.820000 ;
      RECT  5.410000 0.595000  5.580000 1.530000 ;
      RECT  5.410000 1.530000  7.020000 1.700000 ;
      RECT  5.410000 1.700000  5.580000 2.460000 ;
      RECT  5.410000 2.460000  5.765000 2.920000 ;
      RECT  5.750000 0.425000  6.035000 0.690000 ;
      RECT  5.750000 0.690000  7.020000 0.860000 ;
      RECT  5.750000 0.860000  6.035000 1.360000 ;
      RECT  5.750000 1.870000  6.105000 2.200000 ;
      RECT  5.935000 2.200000  6.105000 2.520000 ;
      RECT  5.935000 2.520000  7.735000 2.690000 ;
      RECT  6.245000 1.030000  7.360000 1.360000 ;
      RECT  6.690000 1.700000  7.020000 1.930000 ;
      RECT  6.850000 0.255000  7.860000 0.425000 ;
      RECT  6.850000 0.425000  7.020000 0.690000 ;
      RECT  6.985000 2.100000  7.395000 2.350000 ;
      RECT  7.190000 0.595000  7.520000 0.920000 ;
      RECT  7.190000 0.920000  7.360000 1.030000 ;
      RECT  7.190000 1.360000  7.360000 2.100000 ;
      RECT  7.530000 1.090000  7.860000 1.250000 ;
      RECT  7.530000 1.250000  8.220000 1.355000 ;
      RECT  7.530000 1.355000  8.680000 1.420000 ;
      RECT  7.565000 1.630000  7.880000 1.960000 ;
      RECT  7.565000 1.960000  7.735000 2.520000 ;
      RECT  7.690000 0.425000  7.860000 1.090000 ;
      RECT  7.905000 2.130000  8.235000 2.980000 ;
      RECT  8.030000 0.350000  8.560000 0.810000 ;
      RECT  8.050000 1.420000  8.680000 1.610000 ;
      RECT  8.065000 1.780000  9.020000 1.950000 ;
      RECT  8.065000 1.950000  8.235000 2.130000 ;
      RECT  8.390000 0.810000  8.560000 0.980000 ;
      RECT  8.390000 0.980000  9.020000 1.100000 ;
      RECT  8.390000 1.100000  9.610000 1.150000 ;
      RECT  8.710000 2.120000  9.950000 2.350000 ;
      RECT  8.850000 1.150000  9.610000 1.270000 ;
      RECT  8.850000 1.270000  9.020000 1.780000 ;
      RECT  9.280000 1.270000  9.610000 1.770000 ;
      RECT  9.590000 0.350000  9.950000 0.930000 ;
      RECT  9.600000 1.940000  9.950000 2.120000 ;
      RECT  9.600000 2.350000  9.950000 2.980000 ;
      RECT  9.780000 0.930000  9.950000 1.320000 ;
      RECT  9.780000 1.320000 10.575000 1.650000 ;
      RECT  9.780000 1.650000  9.950000 1.940000 ;
      RECT 11.090000 0.540000 11.310000 1.220000 ;
      RECT 11.090000 1.220000 11.985000 1.550000 ;
      RECT 11.090000 1.550000 11.340000 2.875000 ;
  END
END sky130_fd_sc_hs__sdfxbp_1
