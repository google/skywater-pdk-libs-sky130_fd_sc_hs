* File: sky130_fd_sc_hs__and2b_2.spice
* Created: Tue Sep  1 19:54:57 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hs__and2b_2.pex.spice"
.subckt sky130_fd_sc_hs__and2b_2  VNB VPB A_N B VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* B	B
* A_N	A_N
* VPB	VPB
* VNB	VNB
MM1008 N_VGND_M1008_d N_A_N_M1008_g N_A_27_74#_M1008_s VNB NLOWVT L=0.15 W=0.55
+ AD=0.11874 AS=0.15675 PD=0.989147 PS=1.67 NRD=15.264 NRS=0 M=1 R=3.66667
+ SA=75000.2 SB=75002.6 A=0.0825 P=1.4 MULT=1
MM1002 N_VGND_M1008_d N_A_198_48#_M1002_g N_X_M1002_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.15976 AS=0.1036 PD=1.33085 PS=1.02 NRD=11.34 NRS=0 M=1 R=4.93333
+ SA=75000.6 SB=75002 A=0.111 P=1.78 MULT=1
MM1009 N_VGND_M1009_d N_A_198_48#_M1009_g N_X_M1002_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.29785 AS=0.1036 PD=1.545 PS=1.02 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75001.1
+ SB=75001.6 A=0.111 P=1.78 MULT=1
MM1000 A_505_74# N_B_M1000_g N_VGND_M1009_d VNB NLOWVT L=0.15 W=0.74 AD=0.0888
+ AS=0.29785 PD=0.98 PS=1.545 NRD=10.536 NRS=0 M=1 R=4.93333 SA=75002 SB=75000.6
+ A=0.111 P=1.78 MULT=1
MM1001 N_A_198_48#_M1001_d N_A_27_74#_M1001_g A_505_74# VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.0888 PD=2.05 PS=0.98 NRD=0 NRS=10.536 M=1 R=4.93333 SA=75002.4
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1004 N_VPWR_M1004_d N_A_N_M1004_g N_A_27_74#_M1004_s VPB PSHORT L=0.15 W=0.84
+ AD=0.216043 AS=0.2478 PD=1.37143 PS=2.27 NRD=47.4179 NRS=2.3443 M=1 R=5.6
+ SA=75000.2 SB=75002.5 A=0.126 P=1.98 MULT=1
MM1003 N_X_M1003_d N_A_198_48#_M1003_g N_VPWR_M1004_d VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.288057 PD=1.42 PS=1.82857 NRD=1.7533 NRS=16.7056 M=1 R=7.46667
+ SA=75000.7 SB=75001.8 A=0.168 P=2.54 MULT=1
MM1005 N_X_M1003_d N_A_198_48#_M1005_g N_VPWR_M1005_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.388064 PD=1.42 PS=1.90189 NRD=1.7533 NRS=27.2451 M=1 R=7.46667
+ SA=75001.2 SB=75001.4 A=0.168 P=2.54 MULT=1
MM1006 N_A_198_48#_M1006_d N_B_M1006_g N_VPWR_M1005_s VPB PSHORT L=0.15 W=1
+ AD=0.15 AS=0.346486 PD=1.3 PS=1.69811 NRD=1.9503 NRS=48.2453 M=1 R=6.66667
+ SA=75002 SB=75000.7 A=0.15 P=2.3 MULT=1
MM1007 N_VPWR_M1007_d N_A_27_74#_M1007_g N_A_198_48#_M1006_d VPB PSHORT L=0.15
+ W=1 AD=0.295 AS=0.15 PD=2.59 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=6.66667
+ SA=75002.5 SB=75000.2 A=0.15 P=2.3 MULT=1
DX10_noxref VNB VPB NWDIODE A=6.9564 P=11.2
*
.include "sky130_fd_sc_hs__and2b_2.pxi.spice"
*
.ends
*
*
