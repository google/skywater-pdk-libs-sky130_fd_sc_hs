* File: sky130_fd_sc_hs__buf_2.pxi.spice
* Created: Thu Aug 27 20:34:26 2020
* 
x_PM_SKY130_FD_SC_HS__BUF_2%A_21_260# N_A_21_260#_M1001_d N_A_21_260#_M1005_d
+ N_A_21_260#_c_53_n N_A_21_260#_M1002_g N_A_21_260#_M1000_g N_A_21_260#_M1004_g
+ N_A_21_260#_c_54_n N_A_21_260#_M1003_g N_A_21_260#_c_44_n N_A_21_260#_c_45_n
+ N_A_21_260#_c_46_n N_A_21_260#_c_47_n N_A_21_260#_c_79_p N_A_21_260#_c_78_p
+ N_A_21_260#_c_48_n N_A_21_260#_c_49_n N_A_21_260#_c_50_n N_A_21_260#_c_65_p
+ N_A_21_260#_c_58_n N_A_21_260#_c_59_n N_A_21_260#_c_51_n N_A_21_260#_c_52_n
+ N_A_21_260#_c_82_p N_A_21_260#_c_60_n PM_SKY130_FD_SC_HS__BUF_2%A_21_260#
x_PM_SKY130_FD_SC_HS__BUF_2%A N_A_c_137_n N_A_M1005_g N_A_M1001_g A
+ PM_SKY130_FD_SC_HS__BUF_2%A
x_PM_SKY130_FD_SC_HS__BUF_2%VPWR N_VPWR_M1002_s N_VPWR_M1003_s N_VPWR_c_166_n
+ N_VPWR_c_167_n N_VPWR_c_168_n N_VPWR_c_169_n VPWR N_VPWR_c_170_n
+ N_VPWR_c_171_n N_VPWR_c_165_n PM_SKY130_FD_SC_HS__BUF_2%VPWR
x_PM_SKY130_FD_SC_HS__BUF_2%X N_X_M1000_s N_X_M1002_d N_X_c_207_n X X X X
+ PM_SKY130_FD_SC_HS__BUF_2%X
x_PM_SKY130_FD_SC_HS__BUF_2%VGND N_VGND_M1000_d N_VGND_M1004_d N_VGND_c_226_n
+ N_VGND_c_227_n N_VGND_c_228_n N_VGND_c_229_n VGND N_VGND_c_230_n
+ N_VGND_c_231_n N_VGND_c_232_n N_VGND_c_233_n PM_SKY130_FD_SC_HS__BUF_2%VGND
cc_1 VNB N_A_21_260#_M1000_g 0.0260206f $X=-0.19 $Y=-0.245 $X2=0.895 $Y2=0.74
cc_2 VNB N_A_21_260#_M1004_g 0.0221622f $X=-0.19 $Y=-0.245 $X2=1.325 $Y2=0.74
cc_3 VNB N_A_21_260#_c_44_n 0.0854223f $X=-0.19 $Y=-0.245 $X2=0.795 $Y2=1.465
cc_4 VNB N_A_21_260#_c_45_n 0.045662f $X=-0.19 $Y=-0.245 $X2=1.325 $Y2=1.532
cc_5 VNB N_A_21_260#_c_46_n 0.00193814f $X=-0.19 $Y=-0.245 $X2=0.69 $Y2=1.63
cc_6 VNB N_A_21_260#_c_47_n 0.0011634f $X=-0.19 $Y=-0.245 $X2=0.69 $Y2=2.32
cc_7 VNB N_A_21_260#_c_48_n 0.00890624f $X=-0.19 $Y=-0.245 $X2=1.57 $Y2=2.32
cc_8 VNB N_A_21_260#_c_49_n 0.01461f $X=-0.19 $Y=-0.245 $X2=1.955 $Y2=1.095
cc_9 VNB N_A_21_260#_c_50_n 8.47669e-19 $X=-0.19 $Y=-0.245 $X2=1.655 $Y2=1.095
cc_10 VNB N_A_21_260#_c_51_n 0.0243828f $X=-0.19 $Y=-0.245 $X2=2.12 $Y2=0.615
cc_11 VNB N_A_21_260#_c_52_n 0.0133345f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.465
cc_12 VNB N_A_c_137_n 0.0335823f $X=-0.19 $Y=-0.245 $X2=1.98 $Y2=0.47
cc_13 VNB N_A_M1001_g 0.0339921f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB A 0.0130859f $X=-0.19 $Y=-0.245 $X2=0.885 $Y2=2.4
cc_15 VNB N_VPWR_c_165_n 0.103974f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_X_c_207_n 0.00240191f $X=-0.19 $Y=-0.245 $X2=0.885 $Y2=2.4
cc_17 VNB N_VGND_c_226_n 0.0419262f $X=-0.19 $Y=-0.245 $X2=0.885 $Y2=2.4
cc_18 VNB N_VGND_c_227_n 0.0134303f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_VGND_c_228_n 0.0185316f $X=-0.19 $Y=-0.245 $X2=1.325 $Y2=0.74
cc_20 VNB N_VGND_c_229_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_VGND_c_230_n 0.019013f $X=-0.19 $Y=-0.245 $X2=1.325 $Y2=1.532
cc_22 VNB N_VGND_c_231_n 0.0199267f $X=-0.19 $Y=-0.245 $X2=1.485 $Y2=2.405
cc_23 VNB N_VGND_c_232_n 0.179377f $X=-0.19 $Y=-0.245 $X2=0.775 $Y2=2.405
cc_24 VNB N_VGND_c_233_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=1.955 $Y2=1.095
cc_25 VPB N_A_21_260#_c_53_n 0.0169052f $X=-0.19 $Y=1.66 $X2=0.885 $Y2=1.765
cc_26 VPB N_A_21_260#_c_54_n 0.0168495f $X=-0.19 $Y=1.66 $X2=1.335 $Y2=1.765
cc_27 VPB N_A_21_260#_c_45_n 0.0130549f $X=-0.19 $Y=1.66 $X2=1.325 $Y2=1.532
cc_28 VPB N_A_21_260#_c_47_n 0.00689501f $X=-0.19 $Y=1.66 $X2=0.69 $Y2=2.32
cc_29 VPB N_A_21_260#_c_48_n 0.00332521f $X=-0.19 $Y=1.66 $X2=1.57 $Y2=2.32
cc_30 VPB N_A_21_260#_c_58_n 0.0145954f $X=-0.19 $Y=1.66 $X2=2.105 $Y2=2.035
cc_31 VPB N_A_21_260#_c_59_n 0.0185418f $X=-0.19 $Y=1.66 $X2=2.105 $Y2=2.715
cc_32 VPB N_A_21_260#_c_60_n 0.00704942f $X=-0.19 $Y=1.66 $X2=2.107 $Y2=2.405
cc_33 VPB N_A_c_137_n 0.0347897f $X=-0.19 $Y=1.66 $X2=1.98 $Y2=0.47
cc_34 VPB A 0.00768344f $X=-0.19 $Y=1.66 $X2=0.885 $Y2=2.4
cc_35 VPB N_VPWR_c_166_n 0.0366721f $X=-0.19 $Y=1.66 $X2=0.885 $Y2=2.4
cc_36 VPB N_VPWR_c_167_n 0.0102715f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_37 VPB N_VPWR_c_168_n 0.017758f $X=-0.19 $Y=1.66 $X2=1.325 $Y2=0.74
cc_38 VPB N_VPWR_c_169_n 0.00614127f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_39 VPB N_VPWR_c_170_n 0.0426589f $X=-0.19 $Y=1.66 $X2=1.335 $Y2=2.4
cc_40 VPB N_VPWR_c_171_n 0.0213573f $X=-0.19 $Y=1.66 $X2=1.335 $Y2=1.532
cc_41 VPB N_VPWR_c_165_n 0.0551542f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_42 N_A_21_260#_c_54_n N_A_c_137_n 0.0253316f $X=1.335 $Y=1.765 $X2=-0.19
+ $Y2=-0.245
cc_43 N_A_21_260#_c_45_n N_A_c_137_n 0.01166f $X=1.325 $Y=1.532 $X2=-0.19
+ $Y2=-0.245
cc_44 N_A_21_260#_c_48_n N_A_c_137_n 0.0102819f $X=1.57 $Y=2.32 $X2=-0.19
+ $Y2=-0.245
cc_45 N_A_21_260#_c_49_n N_A_c_137_n 0.00603351f $X=1.955 $Y=1.095 $X2=-0.19
+ $Y2=-0.245
cc_46 N_A_21_260#_c_65_p N_A_c_137_n 0.0116695f $X=1.93 $Y=2.405 $X2=-0.19
+ $Y2=-0.245
cc_47 N_A_21_260#_c_58_n N_A_c_137_n 0.00573434f $X=2.105 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_48 N_A_21_260#_c_59_n N_A_c_137_n 0.00651964f $X=2.105 $Y=2.715 $X2=-0.19
+ $Y2=-0.245
cc_49 N_A_21_260#_c_60_n N_A_c_137_n 2.24111e-19 $X=2.107 $Y=2.405 $X2=-0.19
+ $Y2=-0.245
cc_50 N_A_21_260#_M1004_g N_A_M1001_g 0.0202585f $X=1.325 $Y=0.74 $X2=0 $Y2=0
cc_51 N_A_21_260#_c_48_n N_A_M1001_g 0.00372624f $X=1.57 $Y=2.32 $X2=0 $Y2=0
cc_52 N_A_21_260#_c_49_n N_A_M1001_g 0.0134941f $X=1.955 $Y=1.095 $X2=0 $Y2=0
cc_53 N_A_21_260#_c_51_n N_A_M1001_g 0.00826634f $X=2.12 $Y=0.615 $X2=0 $Y2=0
cc_54 N_A_21_260#_c_48_n A 0.0330647f $X=1.57 $Y=2.32 $X2=0 $Y2=0
cc_55 N_A_21_260#_c_49_n A 0.0373558f $X=1.955 $Y=1.095 $X2=0 $Y2=0
cc_56 N_A_21_260#_c_65_p A 0.00295695f $X=1.93 $Y=2.405 $X2=0 $Y2=0
cc_57 N_A_21_260#_c_58_n A 0.0277278f $X=2.105 $Y=2.035 $X2=0 $Y2=0
cc_58 N_A_21_260#_c_47_n N_VPWR_M1002_s 0.0079747f $X=0.69 $Y=2.32 $X2=-0.19
+ $Y2=-0.245
cc_59 N_A_21_260#_c_78_p N_VPWR_M1002_s 0.00407439f $X=0.775 $Y=2.405 $X2=-0.19
+ $Y2=-0.245
cc_60 N_A_21_260#_c_79_p N_VPWR_M1003_s 8.26908e-19 $X=1.485 $Y=2.405 $X2=0
+ $Y2=0
cc_61 N_A_21_260#_c_48_n N_VPWR_M1003_s 0.0116593f $X=1.57 $Y=2.32 $X2=0 $Y2=0
cc_62 N_A_21_260#_c_65_p N_VPWR_M1003_s 0.00412328f $X=1.93 $Y=2.405 $X2=0 $Y2=0
cc_63 N_A_21_260#_c_82_p N_VPWR_M1003_s 0.00206912f $X=1.57 $Y=2.405 $X2=0 $Y2=0
cc_64 N_A_21_260#_c_53_n N_VPWR_c_166_n 0.00734501f $X=0.885 $Y=1.765 $X2=0
+ $Y2=0
cc_65 N_A_21_260#_c_44_n N_VPWR_c_166_n 0.00698803f $X=0.795 $Y=1.465 $X2=0
+ $Y2=0
cc_66 N_A_21_260#_c_47_n N_VPWR_c_166_n 0.0356886f $X=0.69 $Y=2.32 $X2=0 $Y2=0
cc_67 N_A_21_260#_c_78_p N_VPWR_c_166_n 0.0135162f $X=0.775 $Y=2.405 $X2=0 $Y2=0
cc_68 N_A_21_260#_c_52_n N_VPWR_c_166_n 0.0235035f $X=0.61 $Y=1.465 $X2=0 $Y2=0
cc_69 N_A_21_260#_c_53_n N_VPWR_c_167_n 0.00140553f $X=0.885 $Y=1.765 $X2=0
+ $Y2=0
cc_70 N_A_21_260#_c_54_n N_VPWR_c_167_n 0.0105708f $X=1.335 $Y=1.765 $X2=0 $Y2=0
cc_71 N_A_21_260#_c_79_p N_VPWR_c_167_n 0.00239871f $X=1.485 $Y=2.405 $X2=0
+ $Y2=0
cc_72 N_A_21_260#_c_65_p N_VPWR_c_167_n 0.00545605f $X=1.93 $Y=2.405 $X2=0 $Y2=0
cc_73 N_A_21_260#_c_59_n N_VPWR_c_167_n 0.0149288f $X=2.105 $Y=2.715 $X2=0 $Y2=0
cc_74 N_A_21_260#_c_82_p N_VPWR_c_167_n 0.0148723f $X=1.57 $Y=2.405 $X2=0 $Y2=0
cc_75 N_A_21_260#_c_53_n N_VPWR_c_168_n 0.00413917f $X=0.885 $Y=1.765 $X2=0
+ $Y2=0
cc_76 N_A_21_260#_c_54_n N_VPWR_c_168_n 0.00413917f $X=1.335 $Y=1.765 $X2=0
+ $Y2=0
cc_77 N_A_21_260#_c_53_n N_VPWR_c_170_n 0.00984811f $X=0.885 $Y=1.765 $X2=0
+ $Y2=0
cc_78 N_A_21_260#_c_54_n N_VPWR_c_170_n 0.00104702f $X=1.335 $Y=1.765 $X2=0
+ $Y2=0
cc_79 N_A_21_260#_c_79_p N_VPWR_c_170_n 7.73906e-19 $X=1.485 $Y=2.405 $X2=0
+ $Y2=0
cc_80 N_A_21_260#_c_78_p N_VPWR_c_170_n 0.00951352f $X=0.775 $Y=2.405 $X2=0
+ $Y2=0
cc_81 N_A_21_260#_c_59_n N_VPWR_c_171_n 0.0111689f $X=2.105 $Y=2.715 $X2=0 $Y2=0
cc_82 N_A_21_260#_c_53_n N_VPWR_c_165_n 0.00412855f $X=0.885 $Y=1.765 $X2=0
+ $Y2=0
cc_83 N_A_21_260#_c_54_n N_VPWR_c_165_n 0.00414505f $X=1.335 $Y=1.765 $X2=0
+ $Y2=0
cc_84 N_A_21_260#_c_79_p N_VPWR_c_165_n 0.01825f $X=1.485 $Y=2.405 $X2=0 $Y2=0
cc_85 N_A_21_260#_c_78_p N_VPWR_c_165_n 7.42064e-19 $X=0.775 $Y=2.405 $X2=0
+ $Y2=0
cc_86 N_A_21_260#_c_65_p N_VPWR_c_165_n 0.00687032f $X=1.93 $Y=2.405 $X2=0 $Y2=0
cc_87 N_A_21_260#_c_59_n N_VPWR_c_165_n 0.0122112f $X=2.105 $Y=2.715 $X2=0 $Y2=0
cc_88 N_A_21_260#_c_82_p N_VPWR_c_165_n 6.15054e-19 $X=1.57 $Y=2.405 $X2=0 $Y2=0
cc_89 N_A_21_260#_c_79_p N_X_M1002_d 0.00558496f $X=1.485 $Y=2.405 $X2=0 $Y2=0
cc_90 N_A_21_260#_M1000_g N_X_c_207_n 0.0126407f $X=0.895 $Y=0.74 $X2=0 $Y2=0
cc_91 N_A_21_260#_M1004_g N_X_c_207_n 0.012447f $X=1.325 $Y=0.74 $X2=0 $Y2=0
cc_92 N_A_21_260#_c_50_n N_X_c_207_n 0.012021f $X=1.655 $Y=1.095 $X2=0 $Y2=0
cc_93 N_A_21_260#_c_53_n X 0.00494541f $X=0.885 $Y=1.765 $X2=0 $Y2=0
cc_94 N_A_21_260#_M1000_g X 0.00665606f $X=0.895 $Y=0.74 $X2=0 $Y2=0
cc_95 N_A_21_260#_M1004_g X 0.00500622f $X=1.325 $Y=0.74 $X2=0 $Y2=0
cc_96 N_A_21_260#_c_54_n X 0.00642091f $X=1.335 $Y=1.765 $X2=0 $Y2=0
cc_97 N_A_21_260#_c_45_n X 0.0343295f $X=1.325 $Y=1.532 $X2=0 $Y2=0
cc_98 N_A_21_260#_c_46_n X 0.0264924f $X=0.69 $Y=1.63 $X2=0 $Y2=0
cc_99 N_A_21_260#_c_47_n X 0.0276437f $X=0.69 $Y=2.32 $X2=0 $Y2=0
cc_100 N_A_21_260#_c_79_p X 0.0202284f $X=1.485 $Y=2.405 $X2=0 $Y2=0
cc_101 N_A_21_260#_c_48_n X 0.0729774f $X=1.57 $Y=2.32 $X2=0 $Y2=0
cc_102 N_A_21_260#_c_49_n N_VGND_M1004_d 0.00124373f $X=1.955 $Y=1.095 $X2=0
+ $Y2=0
cc_103 N_A_21_260#_c_50_n N_VGND_M1004_d 0.00366903f $X=1.655 $Y=1.095 $X2=0
+ $Y2=0
cc_104 N_A_21_260#_M1000_g N_VGND_c_226_n 0.00647412f $X=0.895 $Y=0.74 $X2=0
+ $Y2=0
cc_105 N_A_21_260#_c_44_n N_VGND_c_226_n 0.00333176f $X=0.795 $Y=1.465 $X2=0
+ $Y2=0
cc_106 N_A_21_260#_c_46_n N_VGND_c_226_n 0.0141756f $X=0.69 $Y=1.63 $X2=0 $Y2=0
cc_107 N_A_21_260#_c_52_n N_VGND_c_226_n 0.00746796f $X=0.61 $Y=1.465 $X2=0
+ $Y2=0
cc_108 N_A_21_260#_M1004_g N_VGND_c_227_n 0.00760577f $X=1.325 $Y=0.74 $X2=0
+ $Y2=0
cc_109 N_A_21_260#_c_49_n N_VGND_c_227_n 0.00956383f $X=1.955 $Y=1.095 $X2=0
+ $Y2=0
cc_110 N_A_21_260#_c_50_n N_VGND_c_227_n 0.0153275f $X=1.655 $Y=1.095 $X2=0
+ $Y2=0
cc_111 N_A_21_260#_c_51_n N_VGND_c_227_n 0.0147373f $X=2.12 $Y=0.615 $X2=0 $Y2=0
cc_112 N_A_21_260#_M1000_g N_VGND_c_230_n 0.00434272f $X=0.895 $Y=0.74 $X2=0
+ $Y2=0
cc_113 N_A_21_260#_M1004_g N_VGND_c_230_n 0.00434272f $X=1.325 $Y=0.74 $X2=0
+ $Y2=0
cc_114 N_A_21_260#_c_51_n N_VGND_c_231_n 0.0103491f $X=2.12 $Y=0.615 $X2=0 $Y2=0
cc_115 N_A_21_260#_M1000_g N_VGND_c_232_n 0.00825283f $X=0.895 $Y=0.74 $X2=0
+ $Y2=0
cc_116 N_A_21_260#_M1004_g N_VGND_c_232_n 0.00825059f $X=1.325 $Y=0.74 $X2=0
+ $Y2=0
cc_117 N_A_21_260#_c_51_n N_VGND_c_232_n 0.0113354f $X=2.12 $Y=0.615 $X2=0 $Y2=0
cc_118 N_A_c_137_n N_VPWR_c_167_n 0.00451031f $X=1.87 $Y=1.765 $X2=0 $Y2=0
cc_119 N_A_c_137_n N_VPWR_c_171_n 0.00481822f $X=1.87 $Y=1.765 $X2=0 $Y2=0
cc_120 N_A_c_137_n N_VPWR_c_165_n 0.00508379f $X=1.87 $Y=1.765 $X2=0 $Y2=0
cc_121 N_A_M1001_g N_X_c_207_n 9.86633e-19 $X=1.905 $Y=0.79 $X2=0 $Y2=0
cc_122 N_A_M1001_g N_VGND_c_227_n 0.00561794f $X=1.905 $Y=0.79 $X2=0 $Y2=0
cc_123 N_A_M1001_g N_VGND_c_231_n 0.00485498f $X=1.905 $Y=0.79 $X2=0 $Y2=0
cc_124 N_A_M1001_g N_VGND_c_232_n 0.00514438f $X=1.905 $Y=0.79 $X2=0 $Y2=0
cc_125 N_X_c_207_n N_VGND_c_226_n 0.0294122f $X=1.11 $Y=0.515 $X2=0 $Y2=0
cc_126 N_X_c_207_n N_VGND_c_227_n 0.0191765f $X=1.11 $Y=0.515 $X2=0 $Y2=0
cc_127 N_X_c_207_n N_VGND_c_230_n 0.0144922f $X=1.11 $Y=0.515 $X2=0 $Y2=0
cc_128 N_X_c_207_n N_VGND_c_232_n 0.0118826f $X=1.11 $Y=0.515 $X2=0 $Y2=0
