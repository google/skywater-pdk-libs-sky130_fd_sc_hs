# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_hs__dlxtn_1
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_hs__dlxtn_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  6.720000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.208500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105000 1.180000 0.435000 1.565000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.545000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.270000 0.350000 6.605000 2.980000 ;
    END
  END Q
  PIN GATE_N
    ANTENNAGATEAREA  0.237000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.945000 1.500000 1.315000 1.830000 ;
    END
  END GATE_N
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 6.720000 0.085000 ;
        RECT 0.625000  0.085000 0.955000 0.490000 ;
        RECT 2.815000  0.085000 3.145000 1.055000 ;
        RECT 4.850000  0.085000 5.100000 1.135000 ;
        RECT 5.840000  0.085000 6.090000 1.130000 ;
      LAYER mcon ;
        RECT 0.155000 -0.085000 0.325000 0.085000 ;
        RECT 0.635000 -0.085000 0.805000 0.085000 ;
        RECT 1.115000 -0.085000 1.285000 0.085000 ;
        RECT 1.595000 -0.085000 1.765000 0.085000 ;
        RECT 2.075000 -0.085000 2.245000 0.085000 ;
        RECT 2.555000 -0.085000 2.725000 0.085000 ;
        RECT 3.035000 -0.085000 3.205000 0.085000 ;
        RECT 3.515000 -0.085000 3.685000 0.085000 ;
        RECT 3.995000 -0.085000 4.165000 0.085000 ;
        RECT 4.475000 -0.085000 4.645000 0.085000 ;
        RECT 4.955000 -0.085000 5.125000 0.085000 ;
        RECT 5.435000 -0.085000 5.605000 0.085000 ;
        RECT 5.915000 -0.085000 6.085000 0.085000 ;
        RECT 6.395000 -0.085000 6.565000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.245000 6.720000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 3.245000 6.720000 3.415000 ;
        RECT 0.620000 2.075000 0.950000 3.245000 ;
        RECT 2.360000 2.780000 2.705000 3.245000 ;
        RECT 4.470000 2.525000 5.065000 3.245000 ;
        RECT 5.825000 1.820000 6.075000 3.245000 ;
      LAYER mcon ;
        RECT 0.155000 3.245000 0.325000 3.415000 ;
        RECT 0.635000 3.245000 0.805000 3.415000 ;
        RECT 1.115000 3.245000 1.285000 3.415000 ;
        RECT 1.595000 3.245000 1.765000 3.415000 ;
        RECT 2.075000 3.245000 2.245000 3.415000 ;
        RECT 2.555000 3.245000 2.725000 3.415000 ;
        RECT 3.035000 3.245000 3.205000 3.415000 ;
        RECT 3.515000 3.245000 3.685000 3.415000 ;
        RECT 3.995000 3.245000 4.165000 3.415000 ;
        RECT 4.475000 3.245000 4.645000 3.415000 ;
        RECT 4.955000 3.245000 5.125000 3.415000 ;
        RECT 5.435000 3.245000 5.605000 3.415000 ;
        RECT 5.915000 3.245000 6.085000 3.415000 ;
        RECT 6.395000 3.245000 6.565000 3.415000 ;
      LAYER met1 ;
        RECT 0.000000 3.085000 6.720000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.115000 0.555000 0.445000 0.660000 ;
      RECT 0.115000 0.660000 1.315000 0.830000 ;
      RECT 0.115000 0.830000 0.775000 1.010000 ;
      RECT 0.120000 1.735000 0.775000 1.905000 ;
      RECT 0.120000 1.905000 0.450000 2.955000 ;
      RECT 0.605000 1.010000 0.775000 1.735000 ;
      RECT 1.135000 1.000000 1.885000 1.330000 ;
      RECT 1.145000 0.255000 2.645000 0.425000 ;
      RECT 1.145000 0.425000 1.315000 0.660000 ;
      RECT 1.155000 2.075000 1.655000 2.440000 ;
      RECT 1.155000 2.440000 3.045000 2.610000 ;
      RECT 1.155000 2.610000 1.655000 2.955000 ;
      RECT 1.485000 0.760000 1.885000 1.000000 ;
      RECT 1.485000 1.330000 1.885000 1.770000 ;
      RECT 1.485000 1.770000 1.655000 2.075000 ;
      RECT 1.825000 1.940000 2.225000 2.270000 ;
      RECT 2.055000 0.595000 2.305000 1.725000 ;
      RECT 2.055000 1.725000 3.500000 1.895000 ;
      RECT 2.055000 1.895000 2.225000 1.940000 ;
      RECT 2.475000 0.425000 2.645000 1.225000 ;
      RECT 2.475000 1.225000 2.970000 1.555000 ;
      RECT 2.875000 2.610000 3.045000 2.905000 ;
      RECT 2.875000 2.905000 4.180000 3.075000 ;
      RECT 3.180000 1.470000 3.500000 1.725000 ;
      RECT 3.315000 0.255000 4.355000 0.585000 ;
      RECT 3.315000 0.585000 3.485000 1.470000 ;
      RECT 3.330000 2.065000 3.840000 2.735000 ;
      RECT 3.655000 0.805000 4.680000 1.055000 ;
      RECT 3.670000 1.055000 3.840000 2.065000 ;
      RECT 4.010000 1.455000 4.340000 1.785000 ;
      RECT 4.010000 1.785000 4.180000 2.905000 ;
      RECT 4.350000 2.025000 5.655000 2.355000 ;
      RECT 4.510000 1.055000 4.680000 1.305000 ;
      RECT 4.510000 1.305000 5.315000 1.635000 ;
      RECT 5.265000 1.940000 5.655000 2.025000 ;
      RECT 5.265000 2.355000 5.655000 2.980000 ;
      RECT 5.280000 0.455000 5.655000 1.135000 ;
      RECT 5.485000 1.135000 5.655000 1.300000 ;
      RECT 5.485000 1.300000 5.885000 1.630000 ;
      RECT 5.485000 1.630000 5.655000 1.940000 ;
  END
END sky130_fd_sc_hs__dlxtn_1
