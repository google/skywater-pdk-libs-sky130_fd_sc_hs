# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_hs__fa_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  9.120000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAPARTIALMETALSIDEAREA  4.683000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.095000 1.550000 0.385000 1.595000 ;
        RECT 0.095000 1.595000 6.625000 1.735000 ;
        RECT 0.095000 1.735000 0.385000 1.780000 ;
        RECT 2.495000 1.550000 2.785000 1.595000 ;
        RECT 2.495000 1.735000 2.785000 1.780000 ;
        RECT 3.935000 1.550000 4.225000 1.595000 ;
        RECT 3.935000 1.735000 4.225000 1.780000 ;
        RECT 6.335000 1.550000 6.625000 1.595000 ;
        RECT 6.335000 1.735000 6.625000 1.780000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  1.044000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605000 1.920000 0.835000 2.150000 ;
        RECT 0.665000 1.245000 1.165000 1.575000 ;
        RECT 0.665000 1.575000 0.835000 1.920000 ;
    END
  END B
  PIN CIN
    ANTENNAGATEAREA  0.783000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.715000 1.260000 2.225000 1.575000 ;
        RECT 2.055000 1.575000 2.225000 1.950000 ;
        RECT 2.055000 1.950000 4.535000 2.105000 ;
        RECT 2.055000 2.105000 4.195000 2.120000 ;
        RECT 3.215000 1.260000 3.545000 1.575000 ;
        RECT 3.375000 1.575000 3.545000 1.935000 ;
        RECT 3.375000 1.935000 4.535000 1.950000 ;
        RECT 3.375000 2.120000 4.195000 2.150000 ;
        RECT 4.365000 1.745000 5.635000 1.915000 ;
        RECT 4.365000 1.915000 4.535000 1.935000 ;
        RECT 5.305000 1.260000 5.635000 1.745000 ;
    END
  END CIN
  PIN COUT
    ANTENNADIFFAREA  0.649600 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.985000 1.820000 7.555000 2.150000 ;
        RECT 7.105000 0.915000 7.555000 1.085000 ;
        RECT 7.385000 1.085000 7.555000 1.820000 ;
    END
  END COUT
  PIN SUM
    ANTENNADIFFAREA  0.543200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.220000 1.820000 8.575000 2.980000 ;
        RECT 8.245000 0.375000 8.575000 1.150000 ;
        RECT 8.405000 1.150000 8.575000 1.820000 ;
    END
  END SUM
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 9.120000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 9.120000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 9.120000 0.085000 ;
      RECT 0.000000  3.245000 9.120000 3.415000 ;
      RECT 0.095000  1.950000 0.425000 2.320000 ;
      RECT 0.095000  2.320000 1.545000 2.490000 ;
      RECT 0.095000  2.490000 0.445000 2.910000 ;
      RECT 0.105000  1.300000 0.435000 1.780000 ;
      RECT 0.115000  0.375000 0.445000 0.905000 ;
      RECT 0.115000  0.905000 1.205000 1.075000 ;
      RECT 0.115000  1.075000 0.445000 1.130000 ;
      RECT 0.615000  0.085000 0.865000 0.735000 ;
      RECT 0.615000  2.660000 1.010000 3.245000 ;
      RECT 1.035000  0.420000 1.810000 0.750000 ;
      RECT 1.035000  0.750000 1.205000 0.905000 ;
      RECT 1.215000  2.085000 1.545000 2.320000 ;
      RECT 1.215000  2.490000 1.545000 2.755000 ;
      RECT 1.375000  0.920000 6.935000 1.090000 ;
      RECT 1.375000  1.090000 1.545000 1.745000 ;
      RECT 1.375000  1.745000 1.885000 1.915000 ;
      RECT 1.715000  1.915000 1.885000 2.290000 ;
      RECT 1.715000  2.290000 2.185000 2.620000 ;
      RECT 1.980000  0.375000 2.310000 0.920000 ;
      RECT 2.525000  1.260000 3.005000 1.575000 ;
      RECT 2.525000  1.575000 2.755000 1.780000 ;
      RECT 2.800000  0.085000 3.310000 0.705000 ;
      RECT 2.825000  2.290000 3.155000 3.245000 ;
      RECT 3.405000  2.320000 4.825000 2.490000 ;
      RECT 3.405000  2.490000 3.735000 2.755000 ;
      RECT 3.480000  0.375000 3.810000 0.580000 ;
      RECT 3.480000  0.580000 4.970000 0.750000 ;
      RECT 3.905000  2.660000 4.290000 3.245000 ;
      RECT 3.965000  1.260000 4.525000 1.575000 ;
      RECT 3.965000  1.575000 4.195000 1.765000 ;
      RECT 3.990000  0.085000 4.320000 0.410000 ;
      RECT 4.495000  2.275000 4.825000 2.320000 ;
      RECT 4.495000  2.490000 4.825000 2.755000 ;
      RECT 4.500000  0.420000 4.970000 0.580000 ;
      RECT 4.765000  1.090000 5.095000 1.575000 ;
      RECT 5.005000  2.085000 5.335000 2.320000 ;
      RECT 5.005000  2.320000 8.050000 2.490000 ;
      RECT 5.005000  2.490000 5.335000 2.755000 ;
      RECT 5.140000  0.375000 5.470000 0.575000 ;
      RECT 5.140000  0.575000 8.050000 0.745000 ;
      RECT 5.140000  0.745000 5.470000 0.750000 ;
      RECT 6.265000  1.350000 6.595000 1.780000 ;
      RECT 6.470000  0.085000 6.925000 0.405000 ;
      RECT 6.535000  2.660000 6.865000 3.245000 ;
      RECT 6.765000  1.090000 6.935000 1.255000 ;
      RECT 6.765000  1.255000 7.165000 1.585000 ;
      RECT 7.530000  2.730000 8.050000 3.245000 ;
      RECT 7.615000  0.085000 8.065000 0.405000 ;
      RECT 7.880000  0.745000 8.050000 1.320000 ;
      RECT 7.880000  1.320000 8.235000 1.650000 ;
      RECT 7.880000  1.650000 8.050000 2.320000 ;
      RECT 8.750000  1.820000 9.000000 3.245000 ;
      RECT 8.755000  0.085000 9.005000 1.155000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  1.580000 0.325000 1.750000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  1.580000 2.725000 1.750000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  1.580000 4.165000 1.750000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  1.580000 6.565000 1.750000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
      RECT 7.835000 -0.085000 8.005000 0.085000 ;
      RECT 7.835000  3.245000 8.005000 3.415000 ;
      RECT 8.315000 -0.085000 8.485000 0.085000 ;
      RECT 8.315000  3.245000 8.485000 3.415000 ;
      RECT 8.795000 -0.085000 8.965000 0.085000 ;
      RECT 8.795000  3.245000 8.965000 3.415000 ;
  END
END sky130_fd_sc_hs__fa_2
