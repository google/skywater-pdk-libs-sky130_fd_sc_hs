* File: sky130_fd_sc_hs__a2111oi_4.pxi.spice
* Created: Thu Aug 27 20:23:07 2020
* 
x_PM_SKY130_FD_SC_HS__A2111OI_4%D1 N_D1_c_140_n N_D1_M1000_g N_D1_c_141_n
+ N_D1_M1001_g N_D1_c_142_n N_D1_M1002_g N_D1_c_136_n N_D1_M1017_g N_D1_c_137_n
+ N_D1_M1028_g N_D1_c_143_n N_D1_M1003_g D1 D1 D1 N_D1_c_138_n N_D1_c_139_n
+ PM_SKY130_FD_SC_HS__A2111OI_4%D1
x_PM_SKY130_FD_SC_HS__A2111OI_4%C1 N_C1_M1015_g N_C1_c_210_n N_C1_M1007_g
+ N_C1_M1025_g N_C1_c_211_n N_C1_M1009_g N_C1_c_212_n N_C1_M1012_g N_C1_c_213_n
+ N_C1_M1014_g C1 C1 N_C1_c_208_n N_C1_c_209_n PM_SKY130_FD_SC_HS__A2111OI_4%C1
x_PM_SKY130_FD_SC_HS__A2111OI_4%B1 N_B1_M1011_g N_B1_M1022_g N_B1_c_288_n
+ N_B1_M1004_g N_B1_c_289_n N_B1_M1010_g N_B1_c_290_n N_B1_M1013_g N_B1_c_291_n
+ N_B1_M1030_g B1 B1 B1 N_B1_c_286_n N_B1_c_287_n
+ PM_SKY130_FD_SC_HS__A2111OI_4%B1
x_PM_SKY130_FD_SC_HS__A2111OI_4%A1 N_A1_c_362_n N_A1_M1016_g N_A1_M1006_g
+ N_A1_c_363_n N_A1_M1019_g N_A1_M1008_g N_A1_c_364_n N_A1_M1020_g N_A1_M1029_g
+ N_A1_c_365_n N_A1_M1021_g N_A1_M1032_g A1 A1 A1 N_A1_c_361_n
+ PM_SKY130_FD_SC_HS__A2111OI_4%A1
x_PM_SKY130_FD_SC_HS__A2111OI_4%A2 N_A2_M1005_g N_A2_c_446_n N_A2_M1023_g
+ N_A2_M1018_g N_A2_c_447_n N_A2_M1026_g N_A2_M1024_g N_A2_c_448_n N_A2_M1031_g
+ N_A2_M1027_g N_A2_c_449_n N_A2_M1033_g A2 A2 A2 N_A2_c_450_n N_A2_c_445_n
+ PM_SKY130_FD_SC_HS__A2111OI_4%A2
x_PM_SKY130_FD_SC_HS__A2111OI_4%A_29_368# N_A_29_368#_M1000_s
+ N_A_29_368#_M1001_s N_A_29_368#_M1003_s N_A_29_368#_M1009_s
+ N_A_29_368#_M1014_s N_A_29_368#_c_517_n N_A_29_368#_c_518_n
+ N_A_29_368#_c_519_n N_A_29_368#_c_526_n N_A_29_368#_c_520_n
+ N_A_29_368#_c_530_n N_A_29_368#_c_531_n N_A_29_368#_c_537_n
+ N_A_29_368#_c_572_p N_A_29_368#_c_541_n N_A_29_368#_c_521_n
+ N_A_29_368#_c_545_n N_A_29_368#_c_522_n
+ PM_SKY130_FD_SC_HS__A2111OI_4%A_29_368#
x_PM_SKY130_FD_SC_HS__A2111OI_4%Y N_Y_M1017_d N_Y_M1015_d N_Y_M1011_d
+ N_Y_M1006_s N_Y_M1029_s N_Y_M1000_d N_Y_M1002_d N_Y_c_587_n N_Y_c_588_n
+ N_Y_c_600_n N_Y_c_610_n N_Y_c_601_n N_Y_c_618_n N_Y_c_589_n N_Y_c_623_n
+ N_Y_c_590_n N_Y_c_591_n N_Y_c_592_n N_Y_c_593_n N_Y_c_602_n N_Y_c_629_n
+ N_Y_c_594_n N_Y_c_595_n N_Y_c_596_n N_Y_c_597_n N_Y_c_598_n Y Y N_Y_c_604_n Y
+ PM_SKY130_FD_SC_HS__A2111OI_4%Y
x_PM_SKY130_FD_SC_HS__A2111OI_4%A_474_368# N_A_474_368#_M1007_d
+ N_A_474_368#_M1012_d N_A_474_368#_M1004_s N_A_474_368#_M1013_s
+ N_A_474_368#_c_726_n N_A_474_368#_c_720_n N_A_474_368#_c_721_n
+ N_A_474_368#_c_732_n N_A_474_368#_c_722_n N_A_474_368#_c_739_n
+ N_A_474_368#_c_723_n N_A_474_368#_c_745_n N_A_474_368#_c_724_n
+ N_A_474_368#_c_725_n PM_SKY130_FD_SC_HS__A2111OI_4%A_474_368#
x_PM_SKY130_FD_SC_HS__A2111OI_4%A_853_368# N_A_853_368#_M1004_d
+ N_A_853_368#_M1010_d N_A_853_368#_M1030_d N_A_853_368#_M1019_s
+ N_A_853_368#_M1021_s N_A_853_368#_M1026_s N_A_853_368#_M1033_s
+ N_A_853_368#_c_784_n N_A_853_368#_c_785_n N_A_853_368#_c_794_n
+ N_A_853_368#_c_846_n N_A_853_368#_c_798_n N_A_853_368#_c_786_n
+ N_A_853_368#_c_806_n N_A_853_368#_c_787_n N_A_853_368#_c_812_n
+ N_A_853_368#_c_788_n N_A_853_368#_c_821_n N_A_853_368#_c_789_n
+ N_A_853_368#_c_829_n N_A_853_368#_c_790_n N_A_853_368#_c_791_n
+ N_A_853_368#_c_803_n N_A_853_368#_c_817_n N_A_853_368#_c_819_n
+ N_A_853_368#_c_835_n PM_SKY130_FD_SC_HS__A2111OI_4%A_853_368#
x_PM_SKY130_FD_SC_HS__A2111OI_4%VPWR N_VPWR_M1016_d N_VPWR_M1020_d
+ N_VPWR_M1023_d N_VPWR_M1031_d N_VPWR_c_879_n N_VPWR_c_880_n N_VPWR_c_881_n
+ N_VPWR_c_882_n N_VPWR_c_883_n N_VPWR_c_884_n N_VPWR_c_885_n VPWR
+ N_VPWR_c_886_n N_VPWR_c_887_n N_VPWR_c_888_n N_VPWR_c_878_n N_VPWR_c_890_n
+ N_VPWR_c_891_n N_VPWR_c_892_n PM_SKY130_FD_SC_HS__A2111OI_4%VPWR
x_PM_SKY130_FD_SC_HS__A2111OI_4%VGND N_VGND_M1017_s N_VGND_M1028_s
+ N_VGND_M1025_s N_VGND_M1022_s N_VGND_M1005_s N_VGND_M1024_s N_VGND_c_993_n
+ N_VGND_c_994_n N_VGND_c_995_n N_VGND_c_996_n N_VGND_c_997_n N_VGND_c_998_n
+ N_VGND_c_999_n N_VGND_c_1000_n VGND N_VGND_c_1001_n N_VGND_c_1002_n
+ N_VGND_c_1003_n N_VGND_c_1004_n N_VGND_c_1005_n N_VGND_c_1006_n
+ N_VGND_c_1007_n N_VGND_c_1008_n N_VGND_c_1009_n N_VGND_c_1010_n
+ N_VGND_c_1011_n PM_SKY130_FD_SC_HS__A2111OI_4%VGND
x_PM_SKY130_FD_SC_HS__A2111OI_4%A_1228_74# N_A_1228_74#_M1006_d
+ N_A_1228_74#_M1008_d N_A_1228_74#_M1032_d N_A_1228_74#_M1018_d
+ N_A_1228_74#_M1027_d N_A_1228_74#_c_1096_n N_A_1228_74#_c_1097_n
+ N_A_1228_74#_c_1098_n N_A_1228_74#_c_1099_n N_A_1228_74#_c_1100_n
+ N_A_1228_74#_c_1101_n N_A_1228_74#_c_1102_n N_A_1228_74#_c_1103_n
+ N_A_1228_74#_c_1104_n N_A_1228_74#_c_1105_n N_A_1228_74#_c_1106_n
+ PM_SKY130_FD_SC_HS__A2111OI_4%A_1228_74#
cc_1 VNB N_D1_c_136_n 0.0208421f $X=-0.19 $Y=-0.245 $X2=1.4 $Y2=1.22
cc_2 VNB N_D1_c_137_n 0.0162859f $X=-0.19 $Y=-0.245 $X2=1.83 $Y2=1.22
cc_3 VNB N_D1_c_138_n 0.0126583f $X=-0.19 $Y=-0.245 $X2=1.74 $Y2=1.385
cc_4 VNB N_D1_c_139_n 0.127057f $X=-0.19 $Y=-0.245 $X2=1.83 $Y2=1.492
cc_5 VNB N_C1_M1015_g 0.0218891f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.4
cc_6 VNB N_C1_M1025_g 0.0273339f $X=-0.19 $Y=-0.245 $X2=1.4 $Y2=1.22
cc_7 VNB N_C1_c_208_n 0.0948507f $X=-0.19 $Y=-0.245 $X2=1.74 $Y2=1.492
cc_8 VNB N_C1_c_209_n 0.00205555f $X=-0.19 $Y=-0.245 $X2=1.74 $Y2=1.385
cc_9 VNB N_B1_M1011_g 0.0288572f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.4
cc_10 VNB N_B1_M1022_g 0.0305521f $X=-0.19 $Y=-0.245 $X2=1.395 $Y2=1.765
cc_11 VNB N_B1_c_286_n 0.123711f $X=-0.19 $Y=-0.245 $X2=1.74 $Y2=1.385
cc_12 VNB N_B1_c_287_n 0.00264168f $X=-0.19 $Y=-0.245 $X2=1.83 $Y2=1.492
cc_13 VNB N_A1_M1006_g 0.0326041f $X=-0.19 $Y=-0.245 $X2=0.945 $Y2=2.4
cc_14 VNB N_A1_M1008_g 0.0232165f $X=-0.19 $Y=-0.245 $X2=1.83 $Y2=1.22
cc_15 VNB N_A1_M1029_g 0.0233981f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.21
cc_16 VNB N_A1_M1032_g 0.0240711f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.385
cc_17 VNB A1 0.00465397f $X=-0.19 $Y=-0.245 $X2=1.4 $Y2=1.492
cc_18 VNB N_A1_c_361_n 0.0703327f $X=-0.19 $Y=-0.245 $X2=1.74 $Y2=1.365
cc_19 VNB N_A2_M1005_g 0.0230056f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.4
cc_20 VNB N_A2_M1018_g 0.0224899f $X=-0.19 $Y=-0.245 $X2=1.4 $Y2=1.22
cc_21 VNB N_A2_M1024_g 0.0224899f $X=-0.19 $Y=-0.245 $X2=1.845 $Y2=2.4
cc_22 VNB N_A2_M1027_g 0.0318708f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A2_c_445_n 0.0830291f $X=-0.19 $Y=-0.245 $X2=1.74 $Y2=1.365
cc_24 VNB N_Y_c_587_n 0.0224339f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_Y_c_588_n 0.0130653f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_Y_c_589_n 0.00210053f $X=-0.19 $Y=-0.245 $X2=1.845 $Y2=1.492
cc_27 VNB N_Y_c_590_n 0.00206666f $X=-0.19 $Y=-0.245 $X2=1.4 $Y2=1.365
cc_28 VNB N_Y_c_591_n 0.0118592f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_Y_c_592_n 0.00206666f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_Y_c_593_n 0.00249052f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_Y_c_594_n 0.00242779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_Y_c_595_n 0.00507892f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_Y_c_596_n 0.0762531f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_Y_c_597_n 0.00228886f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_Y_c_598_n 0.00250929f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB Y 0.0375295f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_VPWR_c_878_n 0.422413f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_993_n 0.0211662f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=1.21
cc_39 VNB N_VGND_c_994_n 0.00259973f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.492
cc_40 VNB N_VGND_c_995_n 0.0169342f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.385
cc_41 VNB N_VGND_c_996_n 0.0264859f $X=-0.19 $Y=-0.245 $X2=1.4 $Y2=1.492
cc_42 VNB N_VGND_c_997_n 0.00323505f $X=-0.19 $Y=-0.245 $X2=1.74 $Y2=1.385
cc_43 VNB N_VGND_c_998_n 0.00323505f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.365
cc_44 VNB N_VGND_c_999_n 0.0151212f $X=-0.19 $Y=-0.245 $X2=1.2 $Y2=1.365
cc_45 VNB N_VGND_c_1000_n 0.00604233f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_VGND_c_1001_n 0.0346017f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_VGND_c_1002_n 0.0938841f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_VGND_c_1003_n 0.0151736f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_VGND_c_1004_n 0.0197776f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_VGND_c_1005_n 0.573484f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_VGND_c_1006_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_VGND_c_1007_n 0.0169342f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_VGND_c_1008_n 0.037009f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_VGND_c_1009_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_VGND_c_1010_n 0.00604233f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_VGND_c_1011_n 0.00604233f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_A_1228_74#_c_1096_n 0.00310413f $X=-0.19 $Y=-0.245 $X2=1.845 $Y2=2.4
cc_58 VNB N_A_1228_74#_c_1097_n 0.0016059f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.21
cc_59 VNB N_A_1228_74#_c_1098_n 0.00460553f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_A_1228_74#_c_1099_n 0.00406794f $X=-0.19 $Y=-0.245 $X2=0.495
+ $Y2=1.492
cc_61 VNB N_A_1228_74#_c_1100_n 0.00178908f $X=-0.19 $Y=-0.245 $X2=0.72
+ $Y2=1.385
cc_62 VNB N_A_1228_74#_c_1101_n 0.0158169f $X=-0.19 $Y=-0.245 $X2=1.395
+ $Y2=1.492
cc_63 VNB N_A_1228_74#_c_1102_n 0.0266107f $X=-0.19 $Y=-0.245 $X2=1.74 $Y2=1.492
cc_64 VNB N_A_1228_74#_c_1103_n 0.0157537f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.365
cc_65 VNB N_A_1228_74#_c_1104_n 0.00301978f $X=-0.19 $Y=-0.245 $X2=1.2 $Y2=1.365
cc_66 VNB N_A_1228_74#_c_1105_n 0.0017805f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_A_1228_74#_c_1106_n 0.00127131f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VPB N_D1_c_140_n 0.0172279f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.765
cc_69 VPB N_D1_c_141_n 0.0141098f $X=-0.19 $Y=1.66 $X2=0.945 $Y2=1.765
cc_70 VPB N_D1_c_142_n 0.0141098f $X=-0.19 $Y=1.66 $X2=1.395 $Y2=1.765
cc_71 VPB N_D1_c_143_n 0.0148859f $X=-0.19 $Y=1.66 $X2=1.845 $Y2=1.765
cc_72 VPB N_D1_c_139_n 0.0261813f $X=-0.19 $Y=1.66 $X2=1.83 $Y2=1.492
cc_73 VPB N_C1_c_210_n 0.0153205f $X=-0.19 $Y=1.66 $X2=0.945 $Y2=2.4
cc_74 VPB N_C1_c_211_n 0.0146598f $X=-0.19 $Y=1.66 $X2=1.4 $Y2=0.74
cc_75 VPB N_C1_c_212_n 0.0146584f $X=-0.19 $Y=1.66 $X2=1.83 $Y2=0.74
cc_76 VPB N_C1_c_213_n 0.0183217f $X=-0.19 $Y=1.66 $X2=1.845 $Y2=2.4
cc_77 VPB N_C1_c_208_n 0.0475172f $X=-0.19 $Y=1.66 $X2=1.74 $Y2=1.492
cc_78 VPB N_C1_c_209_n 0.00883118f $X=-0.19 $Y=1.66 $X2=1.74 $Y2=1.385
cc_79 VPB N_B1_c_288_n 0.0182952f $X=-0.19 $Y=1.66 $X2=1.395 $Y2=2.4
cc_80 VPB N_B1_c_289_n 0.0146598f $X=-0.19 $Y=1.66 $X2=1.4 $Y2=0.74
cc_81 VPB N_B1_c_290_n 0.0146598f $X=-0.19 $Y=1.66 $X2=1.83 $Y2=0.74
cc_82 VPB N_B1_c_291_n 0.0154562f $X=-0.19 $Y=1.66 $X2=1.845 $Y2=2.4
cc_83 VPB N_B1_c_286_n 0.0660292f $X=-0.19 $Y=1.66 $X2=1.74 $Y2=1.385
cc_84 VPB N_B1_c_287_n 0.0137732f $X=-0.19 $Y=1.66 $X2=1.83 $Y2=1.492
cc_85 VPB N_A1_c_362_n 0.0153762f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.765
cc_86 VPB N_A1_c_363_n 0.0149968f $X=-0.19 $Y=1.66 $X2=1.395 $Y2=2.4
cc_87 VPB N_A1_c_364_n 0.0149968f $X=-0.19 $Y=1.66 $X2=1.83 $Y2=0.74
cc_88 VPB N_A1_c_365_n 0.015303f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_89 VPB A1 0.0107427f $X=-0.19 $Y=1.66 $X2=1.4 $Y2=1.492
cc_90 VPB N_A1_c_361_n 0.0461433f $X=-0.19 $Y=1.66 $X2=1.74 $Y2=1.365
cc_91 VPB N_A2_c_446_n 0.0153734f $X=-0.19 $Y=1.66 $X2=0.945 $Y2=2.4
cc_92 VPB N_A2_c_447_n 0.0155127f $X=-0.19 $Y=1.66 $X2=1.4 $Y2=0.74
cc_93 VPB N_A2_c_448_n 0.0155119f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.21
cc_94 VPB N_A2_c_449_n 0.0198646f $X=-0.19 $Y=1.66 $X2=0.72 $Y2=1.492
cc_95 VPB N_A2_c_450_n 0.0083958f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_96 VPB N_A2_c_445_n 0.0499225f $X=-0.19 $Y=1.66 $X2=1.74 $Y2=1.365
cc_97 VPB N_A_29_368#_c_517_n 0.0325715f $X=-0.19 $Y=1.66 $X2=1.845 $Y2=2.4
cc_98 VPB N_A_29_368#_c_518_n 0.0030474f $X=-0.19 $Y=1.66 $X2=1.115 $Y2=1.21
cc_99 VPB N_A_29_368#_c_519_n 0.0093919f $X=-0.19 $Y=1.66 $X2=1.595 $Y2=1.21
cc_100 VPB N_A_29_368#_c_520_n 0.00477562f $X=-0.19 $Y=1.66 $X2=0.72 $Y2=1.492
cc_101 VPB N_A_29_368#_c_521_n 0.00123754f $X=-0.19 $Y=1.66 $X2=1.2 $Y2=1.365
cc_102 VPB N_A_29_368#_c_522_n 0.0143923f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_103 VPB N_Y_c_600_n 0.00168332f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_104 VPB N_Y_c_601_n 0.00531797f $X=-0.19 $Y=1.66 $X2=1.395 $Y2=1.492
cc_105 VPB N_Y_c_602_n 0.00224287f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_106 VPB Y 0.00287511f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_107 VPB N_Y_c_604_n 0.00758256f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_108 VPB N_A_474_368#_c_720_n 0.00213603f $X=-0.19 $Y=1.66 $X2=1.845 $Y2=2.4
cc_109 VPB N_A_474_368#_c_721_n 0.00266046f $X=-0.19 $Y=1.66 $X2=1.845 $Y2=2.4
cc_110 VPB N_A_474_368#_c_722_n 0.0163588f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_111 VPB N_A_474_368#_c_723_n 0.00431993f $X=-0.19 $Y=1.66 $X2=0.945 $Y2=1.492
cc_112 VPB N_A_474_368#_c_724_n 0.0021839f $X=-0.19 $Y=1.66 $X2=1.74 $Y2=1.385
cc_113 VPB N_A_474_368#_c_725_n 0.0021839f $X=-0.19 $Y=1.66 $X2=1.74 $Y2=1.385
cc_114 VPB N_A_853_368#_c_784_n 0.00171922f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_115 VPB N_A_853_368#_c_785_n 0.00539749f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_116 VPB N_A_853_368#_c_786_n 0.00180901f $X=-0.19 $Y=1.66 $X2=1.74 $Y2=1.385
cc_117 VPB N_A_853_368#_c_787_n 0.00180921f $X=-0.19 $Y=1.66 $X2=1.2 $Y2=1.365
cc_118 VPB N_A_853_368#_c_788_n 0.00180921f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_119 VPB N_A_853_368#_c_789_n 0.00257348f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_120 VPB N_A_853_368#_c_790_n 0.0185714f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_121 VPB N_A_853_368#_c_791_n 0.0345863f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_122 VPB N_VPWR_c_879_n 0.00329129f $X=-0.19 $Y=1.66 $X2=1.83 $Y2=0.74
cc_123 VPB N_VPWR_c_880_n 0.0164465f $X=-0.19 $Y=1.66 $X2=1.845 $Y2=2.4
cc_124 VPB N_VPWR_c_881_n 0.00261791f $X=-0.19 $Y=1.66 $X2=1.595 $Y2=1.21
cc_125 VPB N_VPWR_c_882_n 0.00504372f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.492
cc_126 VPB N_VPWR_c_883_n 0.00571271f $X=-0.19 $Y=1.66 $X2=0.945 $Y2=1.492
cc_127 VPB N_VPWR_c_884_n 0.152862f $X=-0.19 $Y=1.66 $X2=1.4 $Y2=1.492
cc_128 VPB N_VPWR_c_885_n 0.00601644f $X=-0.19 $Y=1.66 $X2=1.4 $Y2=1.385
cc_129 VPB N_VPWR_c_886_n 0.0164465f $X=-0.19 $Y=1.66 $X2=1.2 $Y2=1.365
cc_130 VPB N_VPWR_c_887_n 0.0206041f $X=-0.19 $Y=1.66 $X2=1.74 $Y2=1.365
cc_131 VPB N_VPWR_c_888_n 0.0177091f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_132 VPB N_VPWR_c_878_n 0.109443f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_133 VPB N_VPWR_c_890_n 0.00601644f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_134 VPB N_VPWR_c_891_n 0.00460249f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_135 VPB N_VPWR_c_892_n 0.00460249f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_136 N_D1_c_137_n N_C1_M1015_g 0.0174718f $X=1.83 $Y=1.22 $X2=0 $Y2=0
cc_137 N_D1_c_138_n N_C1_M1015_g 0.00131191f $X=1.74 $Y=1.385 $X2=0 $Y2=0
cc_138 N_D1_c_143_n N_C1_c_210_n 0.010221f $X=1.845 $Y=1.765 $X2=0 $Y2=0
cc_139 N_D1_c_138_n N_C1_c_208_n 3.91262e-19 $X=1.74 $Y=1.385 $X2=0 $Y2=0
cc_140 N_D1_c_139_n N_C1_c_208_n 0.0335167f $X=1.83 $Y=1.492 $X2=0 $Y2=0
cc_141 N_D1_c_138_n N_C1_c_209_n 0.00980746f $X=1.74 $Y=1.385 $X2=0 $Y2=0
cc_142 N_D1_c_139_n N_C1_c_209_n 0.00194335f $X=1.83 $Y=1.492 $X2=0 $Y2=0
cc_143 N_D1_c_140_n N_A_29_368#_c_517_n 0.00970707f $X=0.495 $Y=1.765 $X2=0
+ $Y2=0
cc_144 N_D1_c_140_n N_A_29_368#_c_518_n 0.0137046f $X=0.495 $Y=1.765 $X2=0 $Y2=0
cc_145 N_D1_c_141_n N_A_29_368#_c_518_n 0.0128349f $X=0.945 $Y=1.765 $X2=0 $Y2=0
cc_146 N_D1_c_141_n N_A_29_368#_c_526_n 0.0062909f $X=0.945 $Y=1.765 $X2=0 $Y2=0
cc_147 N_D1_c_142_n N_A_29_368#_c_526_n 0.00443541f $X=1.395 $Y=1.765 $X2=0
+ $Y2=0
cc_148 N_D1_c_142_n N_A_29_368#_c_520_n 0.0128349f $X=1.395 $Y=1.765 $X2=0 $Y2=0
cc_149 N_D1_c_143_n N_A_29_368#_c_520_n 0.0125587f $X=1.845 $Y=1.765 $X2=0 $Y2=0
cc_150 N_D1_c_143_n N_A_29_368#_c_530_n 0.00242156f $X=1.845 $Y=1.765 $X2=0
+ $Y2=0
cc_151 N_D1_c_142_n N_A_29_368#_c_531_n 7.24405e-19 $X=1.395 $Y=1.765 $X2=0
+ $Y2=0
cc_152 N_D1_c_143_n N_A_29_368#_c_531_n 0.00989155f $X=1.845 $Y=1.765 $X2=0
+ $Y2=0
cc_153 N_D1_c_136_n N_Y_c_587_n 0.0116578f $X=1.4 $Y=1.22 $X2=0 $Y2=0
cc_154 N_D1_c_138_n N_Y_c_587_n 0.0722866f $X=1.74 $Y=1.385 $X2=0 $Y2=0
cc_155 N_D1_c_139_n N_Y_c_587_n 0.0106419f $X=1.83 $Y=1.492 $X2=0 $Y2=0
cc_156 N_D1_c_140_n N_Y_c_600_n 0.00994474f $X=0.495 $Y=1.765 $X2=0 $Y2=0
cc_157 N_D1_c_139_n N_Y_c_600_n 0.00796487f $X=1.83 $Y=1.492 $X2=0 $Y2=0
cc_158 N_D1_c_140_n N_Y_c_610_n 0.0171108f $X=0.495 $Y=1.765 $X2=0 $Y2=0
cc_159 N_D1_c_141_n N_Y_c_610_n 0.0124829f $X=0.945 $Y=1.765 $X2=0 $Y2=0
cc_160 N_D1_c_142_n N_Y_c_610_n 6.41034e-19 $X=1.395 $Y=1.765 $X2=0 $Y2=0
cc_161 N_D1_c_141_n N_Y_c_601_n 0.00899835f $X=0.945 $Y=1.765 $X2=0 $Y2=0
cc_162 N_D1_c_142_n N_Y_c_601_n 0.00991644f $X=1.395 $Y=1.765 $X2=0 $Y2=0
cc_163 N_D1_c_143_n N_Y_c_601_n 0.00347702f $X=1.845 $Y=1.765 $X2=0 $Y2=0
cc_164 N_D1_c_138_n N_Y_c_601_n 0.0631462f $X=1.74 $Y=1.385 $X2=0 $Y2=0
cc_165 N_D1_c_139_n N_Y_c_601_n 0.0129335f $X=1.83 $Y=1.492 $X2=0 $Y2=0
cc_166 N_D1_c_141_n N_Y_c_618_n 6.4339e-19 $X=0.945 $Y=1.765 $X2=0 $Y2=0
cc_167 N_D1_c_142_n N_Y_c_618_n 0.011908f $X=1.395 $Y=1.765 $X2=0 $Y2=0
cc_168 N_D1_c_143_n N_Y_c_618_n 0.00481138f $X=1.845 $Y=1.765 $X2=0 $Y2=0
cc_169 N_D1_c_136_n N_Y_c_589_n 4.50863e-19 $X=1.4 $Y=1.22 $X2=0 $Y2=0
cc_170 N_D1_c_137_n N_Y_c_589_n 4.50863e-19 $X=1.83 $Y=1.22 $X2=0 $Y2=0
cc_171 N_D1_c_137_n N_Y_c_623_n 0.00957073f $X=1.83 $Y=1.22 $X2=0 $Y2=0
cc_172 N_D1_c_138_n N_Y_c_623_n 0.0131073f $X=1.74 $Y=1.385 $X2=0 $Y2=0
cc_173 N_D1_c_140_n N_Y_c_602_n 0.00109449f $X=0.495 $Y=1.765 $X2=0 $Y2=0
cc_174 N_D1_c_141_n N_Y_c_602_n 0.00109449f $X=0.945 $Y=1.765 $X2=0 $Y2=0
cc_175 N_D1_c_138_n N_Y_c_602_n 0.0277828f $X=1.74 $Y=1.385 $X2=0 $Y2=0
cc_176 N_D1_c_139_n N_Y_c_602_n 0.00501057f $X=1.83 $Y=1.492 $X2=0 $Y2=0
cc_177 N_D1_c_138_n N_Y_c_629_n 0.0146818f $X=1.74 $Y=1.385 $X2=0 $Y2=0
cc_178 N_D1_c_139_n N_Y_c_629_n 7.07126e-19 $X=1.83 $Y=1.492 $X2=0 $Y2=0
cc_179 N_D1_c_138_n Y 0.0267576f $X=1.74 $Y=1.385 $X2=0 $Y2=0
cc_180 N_D1_c_139_n Y 0.0172496f $X=1.83 $Y=1.492 $X2=0 $Y2=0
cc_181 N_D1_c_140_n N_VPWR_c_884_n 0.00278271f $X=0.495 $Y=1.765 $X2=0 $Y2=0
cc_182 N_D1_c_141_n N_VPWR_c_884_n 0.00278271f $X=0.945 $Y=1.765 $X2=0 $Y2=0
cc_183 N_D1_c_142_n N_VPWR_c_884_n 0.00278271f $X=1.395 $Y=1.765 $X2=0 $Y2=0
cc_184 N_D1_c_143_n N_VPWR_c_884_n 0.00278257f $X=1.845 $Y=1.765 $X2=0 $Y2=0
cc_185 N_D1_c_140_n N_VPWR_c_878_n 0.00357283f $X=0.495 $Y=1.765 $X2=0 $Y2=0
cc_186 N_D1_c_141_n N_VPWR_c_878_n 0.00353823f $X=0.945 $Y=1.765 $X2=0 $Y2=0
cc_187 N_D1_c_142_n N_VPWR_c_878_n 0.00353823f $X=1.395 $Y=1.765 $X2=0 $Y2=0
cc_188 N_D1_c_143_n N_VPWR_c_878_n 0.00353905f $X=1.845 $Y=1.765 $X2=0 $Y2=0
cc_189 N_D1_c_136_n N_VGND_c_993_n 0.00850375f $X=1.4 $Y=1.22 $X2=0 $Y2=0
cc_190 N_D1_c_137_n N_VGND_c_993_n 3.67997e-19 $X=1.83 $Y=1.22 $X2=0 $Y2=0
cc_191 N_D1_c_136_n N_VGND_c_994_n 3.67997e-19 $X=1.4 $Y=1.22 $X2=0 $Y2=0
cc_192 N_D1_c_137_n N_VGND_c_994_n 0.0074045f $X=1.83 $Y=1.22 $X2=0 $Y2=0
cc_193 N_D1_c_136_n N_VGND_c_999_n 0.00383152f $X=1.4 $Y=1.22 $X2=0 $Y2=0
cc_194 N_D1_c_137_n N_VGND_c_999_n 0.00383152f $X=1.83 $Y=1.22 $X2=0 $Y2=0
cc_195 N_D1_c_136_n N_VGND_c_1005_n 0.00383967f $X=1.4 $Y=1.22 $X2=0 $Y2=0
cc_196 N_D1_c_137_n N_VGND_c_1005_n 0.00383967f $X=1.83 $Y=1.22 $X2=0 $Y2=0
cc_197 N_C1_c_208_n N_B1_M1011_g 0.01353f $X=3.42 $Y=1.515 $X2=0 $Y2=0
cc_198 N_C1_c_208_n N_B1_c_286_n 0.00780189f $X=3.42 $Y=1.515 $X2=0 $Y2=0
cc_199 N_C1_c_209_n N_B1_c_286_n 0.00157841f $X=3.42 $Y=1.515 $X2=0 $Y2=0
cc_200 N_C1_c_213_n N_B1_c_287_n 3.73855e-19 $X=3.645 $Y=1.765 $X2=0 $Y2=0
cc_201 N_C1_c_208_n N_B1_c_287_n 0.00402291f $X=3.42 $Y=1.515 $X2=0 $Y2=0
cc_202 N_C1_c_210_n N_A_29_368#_c_520_n 0.00322215f $X=2.295 $Y=1.765 $X2=0
+ $Y2=0
cc_203 N_C1_c_210_n N_A_29_368#_c_530_n 4.96706e-19 $X=2.295 $Y=1.765 $X2=0
+ $Y2=0
cc_204 N_C1_c_210_n N_A_29_368#_c_531_n 0.00981849f $X=2.295 $Y=1.765 $X2=0
+ $Y2=0
cc_205 N_C1_c_211_n N_A_29_368#_c_531_n 4.45174e-19 $X=2.745 $Y=1.765 $X2=0
+ $Y2=0
cc_206 N_C1_c_210_n N_A_29_368#_c_537_n 0.0120074f $X=2.295 $Y=1.765 $X2=0 $Y2=0
cc_207 N_C1_c_211_n N_A_29_368#_c_537_n 0.0126853f $X=2.745 $Y=1.765 $X2=0 $Y2=0
cc_208 N_C1_c_208_n N_A_29_368#_c_537_n 0.0013078f $X=3.42 $Y=1.515 $X2=0 $Y2=0
cc_209 N_C1_c_209_n N_A_29_368#_c_537_n 0.0419986f $X=3.42 $Y=1.515 $X2=0 $Y2=0
cc_210 N_C1_c_212_n N_A_29_368#_c_541_n 0.0126853f $X=3.195 $Y=1.765 $X2=0 $Y2=0
cc_211 N_C1_c_213_n N_A_29_368#_c_541_n 0.0154604f $X=3.645 $Y=1.765 $X2=0 $Y2=0
cc_212 N_C1_c_208_n N_A_29_368#_c_541_n 0.00215835f $X=3.42 $Y=1.515 $X2=0 $Y2=0
cc_213 N_C1_c_209_n N_A_29_368#_c_541_n 0.0294734f $X=3.42 $Y=1.515 $X2=0 $Y2=0
cc_214 N_C1_c_208_n N_A_29_368#_c_545_n 0.00130557f $X=3.42 $Y=1.515 $X2=0 $Y2=0
cc_215 N_C1_c_209_n N_A_29_368#_c_545_n 0.0183565f $X=3.42 $Y=1.515 $X2=0 $Y2=0
cc_216 N_C1_c_212_n N_A_29_368#_c_522_n 6.18219e-19 $X=3.195 $Y=1.765 $X2=0
+ $Y2=0
cc_217 N_C1_c_213_n N_A_29_368#_c_522_n 0.00430911f $X=3.645 $Y=1.765 $X2=0
+ $Y2=0
cc_218 N_C1_c_208_n N_A_29_368#_c_522_n 5.14738e-19 $X=3.42 $Y=1.515 $X2=0 $Y2=0
cc_219 N_C1_c_209_n N_Y_c_601_n 0.00219629f $X=3.42 $Y=1.515 $X2=0 $Y2=0
cc_220 N_C1_M1015_g N_Y_c_623_n 0.0112633f $X=2.26 $Y=0.74 $X2=0 $Y2=0
cc_221 N_C1_c_209_n N_Y_c_623_n 0.00539983f $X=3.42 $Y=1.515 $X2=0 $Y2=0
cc_222 N_C1_M1015_g N_Y_c_590_n 3.97481e-19 $X=2.26 $Y=0.74 $X2=0 $Y2=0
cc_223 N_C1_M1025_g N_Y_c_590_n 0.00615586f $X=2.69 $Y=0.74 $X2=0 $Y2=0
cc_224 N_C1_M1025_g N_Y_c_591_n 0.0142398f $X=2.69 $Y=0.74 $X2=0 $Y2=0
cc_225 N_C1_c_208_n N_Y_c_591_n 0.0276022f $X=3.42 $Y=1.515 $X2=0 $Y2=0
cc_226 N_C1_c_209_n N_Y_c_591_n 0.0662651f $X=3.42 $Y=1.515 $X2=0 $Y2=0
cc_227 N_C1_M1015_g N_Y_c_594_n 0.00177693f $X=2.26 $Y=0.74 $X2=0 $Y2=0
cc_228 N_C1_M1025_g N_Y_c_594_n 0.00906122f $X=2.69 $Y=0.74 $X2=0 $Y2=0
cc_229 N_C1_c_208_n N_Y_c_594_n 0.00245733f $X=3.42 $Y=1.515 $X2=0 $Y2=0
cc_230 N_C1_c_209_n N_Y_c_594_n 0.0211949f $X=3.42 $Y=1.515 $X2=0 $Y2=0
cc_231 N_C1_c_211_n N_A_474_368#_c_726_n 0.00735508f $X=2.745 $Y=1.765 $X2=0
+ $Y2=0
cc_232 N_C1_c_212_n N_A_474_368#_c_726_n 5.53825e-19 $X=3.195 $Y=1.765 $X2=0
+ $Y2=0
cc_233 N_C1_c_211_n N_A_474_368#_c_720_n 0.0108414f $X=2.745 $Y=1.765 $X2=0
+ $Y2=0
cc_234 N_C1_c_212_n N_A_474_368#_c_720_n 0.0107904f $X=3.195 $Y=1.765 $X2=0
+ $Y2=0
cc_235 N_C1_c_210_n N_A_474_368#_c_721_n 0.00124692f $X=2.295 $Y=1.765 $X2=0
+ $Y2=0
cc_236 N_C1_c_211_n N_A_474_368#_c_721_n 0.0014181f $X=2.745 $Y=1.765 $X2=0
+ $Y2=0
cc_237 N_C1_c_211_n N_A_474_368#_c_732_n 5.52094e-19 $X=2.745 $Y=1.765 $X2=0
+ $Y2=0
cc_238 N_C1_c_212_n N_A_474_368#_c_732_n 0.00767389f $X=3.195 $Y=1.765 $X2=0
+ $Y2=0
cc_239 N_C1_c_213_n N_A_474_368#_c_732_n 0.0121282f $X=3.645 $Y=1.765 $X2=0
+ $Y2=0
cc_240 N_C1_c_213_n N_A_474_368#_c_722_n 0.012762f $X=3.645 $Y=1.765 $X2=0 $Y2=0
cc_241 N_C1_c_212_n N_A_474_368#_c_724_n 0.00175197f $X=3.195 $Y=1.765 $X2=0
+ $Y2=0
cc_242 N_C1_c_213_n N_A_474_368#_c_724_n 0.00175197f $X=3.645 $Y=1.765 $X2=0
+ $Y2=0
cc_243 N_C1_c_210_n N_VPWR_c_884_n 0.0044313f $X=2.295 $Y=1.765 $X2=0 $Y2=0
cc_244 N_C1_c_211_n N_VPWR_c_884_n 0.00278257f $X=2.745 $Y=1.765 $X2=0 $Y2=0
cc_245 N_C1_c_212_n N_VPWR_c_884_n 0.00278257f $X=3.195 $Y=1.765 $X2=0 $Y2=0
cc_246 N_C1_c_213_n N_VPWR_c_884_n 0.00278257f $X=3.645 $Y=1.765 $X2=0 $Y2=0
cc_247 N_C1_c_210_n N_VPWR_c_878_n 0.00854206f $X=2.295 $Y=1.765 $X2=0 $Y2=0
cc_248 N_C1_c_211_n N_VPWR_c_878_n 0.00353822f $X=2.745 $Y=1.765 $X2=0 $Y2=0
cc_249 N_C1_c_212_n N_VPWR_c_878_n 0.00353822f $X=3.195 $Y=1.765 $X2=0 $Y2=0
cc_250 N_C1_c_213_n N_VPWR_c_878_n 0.00358623f $X=3.645 $Y=1.765 $X2=0 $Y2=0
cc_251 N_C1_M1015_g N_VGND_c_994_n 0.00766594f $X=2.26 $Y=0.74 $X2=0 $Y2=0
cc_252 N_C1_M1025_g N_VGND_c_994_n 4.39708e-19 $X=2.69 $Y=0.74 $X2=0 $Y2=0
cc_253 N_C1_M1015_g N_VGND_c_1005_n 0.00383967f $X=2.26 $Y=0.74 $X2=0 $Y2=0
cc_254 N_C1_M1025_g N_VGND_c_1005_n 0.00825037f $X=2.69 $Y=0.74 $X2=0 $Y2=0
cc_255 N_C1_M1015_g N_VGND_c_1007_n 0.00383152f $X=2.26 $Y=0.74 $X2=0 $Y2=0
cc_256 N_C1_M1025_g N_VGND_c_1007_n 0.00434272f $X=2.69 $Y=0.74 $X2=0 $Y2=0
cc_257 N_C1_M1025_g N_VGND_c_1008_n 0.00597094f $X=2.69 $Y=0.74 $X2=0 $Y2=0
cc_258 N_B1_c_291_n N_A1_c_362_n 0.00841319f $X=5.985 $Y=1.765 $X2=-0.19
+ $Y2=-0.245
cc_259 N_B1_c_286_n A1 4.47344e-19 $X=5.91 $Y=1.515 $X2=0 $Y2=0
cc_260 N_B1_c_287_n A1 0.019126f $X=5.91 $Y=1.515 $X2=0 $Y2=0
cc_261 N_B1_c_286_n N_A1_c_361_n 0.0199753f $X=5.91 $Y=1.515 $X2=0 $Y2=0
cc_262 N_B1_c_287_n N_A1_c_361_n 0.00184572f $X=5.91 $Y=1.515 $X2=0 $Y2=0
cc_263 N_B1_c_288_n N_A_29_368#_c_522_n 0.002051f $X=4.635 $Y=1.765 $X2=0 $Y2=0
cc_264 N_B1_c_286_n N_A_29_368#_c_522_n 0.00251593f $X=5.91 $Y=1.515 $X2=0 $Y2=0
cc_265 N_B1_M1011_g N_Y_c_591_n 0.0149534f $X=4.02 $Y=0.74 $X2=0 $Y2=0
cc_266 N_B1_M1011_g N_Y_c_592_n 0.0118293f $X=4.02 $Y=0.74 $X2=0 $Y2=0
cc_267 N_B1_M1022_g N_Y_c_592_n 3.97481e-19 $X=4.45 $Y=0.74 $X2=0 $Y2=0
cc_268 N_B1_M1011_g N_Y_c_595_n 0.0040828f $X=4.02 $Y=0.74 $X2=0 $Y2=0
cc_269 N_B1_c_286_n N_Y_c_595_n 0.00423267f $X=5.91 $Y=1.515 $X2=0 $Y2=0
cc_270 N_B1_c_287_n N_Y_c_595_n 0.00386581f $X=5.91 $Y=1.515 $X2=0 $Y2=0
cc_271 N_B1_M1022_g N_Y_c_596_n 0.0166073f $X=4.45 $Y=0.74 $X2=0 $Y2=0
cc_272 N_B1_c_286_n N_Y_c_596_n 0.0373961f $X=5.91 $Y=1.515 $X2=0 $Y2=0
cc_273 N_B1_c_287_n N_Y_c_596_n 0.135914f $X=5.91 $Y=1.515 $X2=0 $Y2=0
cc_274 N_B1_c_288_n N_A_474_368#_c_722_n 0.012762f $X=4.635 $Y=1.765 $X2=0 $Y2=0
cc_275 N_B1_c_288_n N_A_474_368#_c_739_n 0.0123195f $X=4.635 $Y=1.765 $X2=0
+ $Y2=0
cc_276 N_B1_c_289_n N_A_474_368#_c_739_n 0.00786518f $X=5.085 $Y=1.765 $X2=0
+ $Y2=0
cc_277 N_B1_c_290_n N_A_474_368#_c_739_n 5.52094e-19 $X=5.535 $Y=1.765 $X2=0
+ $Y2=0
cc_278 N_B1_c_289_n N_A_474_368#_c_723_n 0.0108414f $X=5.085 $Y=1.765 $X2=0
+ $Y2=0
cc_279 N_B1_c_290_n N_A_474_368#_c_723_n 0.0125934f $X=5.535 $Y=1.765 $X2=0
+ $Y2=0
cc_280 N_B1_c_291_n N_A_474_368#_c_723_n 0.00396164f $X=5.985 $Y=1.765 $X2=0
+ $Y2=0
cc_281 N_B1_c_289_n N_A_474_368#_c_745_n 5.52094e-19 $X=5.085 $Y=1.765 $X2=0
+ $Y2=0
cc_282 N_B1_c_290_n N_A_474_368#_c_745_n 0.00786518f $X=5.535 $Y=1.765 $X2=0
+ $Y2=0
cc_283 N_B1_c_291_n N_A_474_368#_c_745_n 0.00692938f $X=5.985 $Y=1.765 $X2=0
+ $Y2=0
cc_284 N_B1_c_288_n N_A_474_368#_c_725_n 0.00175197f $X=4.635 $Y=1.765 $X2=0
+ $Y2=0
cc_285 N_B1_c_289_n N_A_474_368#_c_725_n 0.00175197f $X=5.085 $Y=1.765 $X2=0
+ $Y2=0
cc_286 N_B1_c_286_n N_A_853_368#_c_784_n 0.00266667f $X=5.91 $Y=1.515 $X2=0
+ $Y2=0
cc_287 N_B1_c_287_n N_A_853_368#_c_784_n 0.0211118f $X=5.91 $Y=1.515 $X2=0 $Y2=0
cc_288 N_B1_c_288_n N_A_853_368#_c_794_n 0.0126853f $X=4.635 $Y=1.765 $X2=0
+ $Y2=0
cc_289 N_B1_c_289_n N_A_853_368#_c_794_n 0.0126853f $X=5.085 $Y=1.765 $X2=0
+ $Y2=0
cc_290 N_B1_c_286_n N_A_853_368#_c_794_n 0.00132059f $X=5.91 $Y=1.515 $X2=0
+ $Y2=0
cc_291 N_B1_c_287_n N_A_853_368#_c_794_n 0.0446098f $X=5.91 $Y=1.515 $X2=0 $Y2=0
cc_292 N_B1_c_290_n N_A_853_368#_c_798_n 0.0126853f $X=5.535 $Y=1.765 $X2=0
+ $Y2=0
cc_293 N_B1_c_291_n N_A_853_368#_c_798_n 0.0126853f $X=5.985 $Y=1.765 $X2=0
+ $Y2=0
cc_294 N_B1_c_286_n N_A_853_368#_c_798_n 0.00132059f $X=5.91 $Y=1.515 $X2=0
+ $Y2=0
cc_295 N_B1_c_287_n N_A_853_368#_c_798_n 0.0437431f $X=5.91 $Y=1.515 $X2=0 $Y2=0
cc_296 N_B1_c_291_n N_A_853_368#_c_786_n 0.00557061f $X=5.985 $Y=1.765 $X2=0
+ $Y2=0
cc_297 N_B1_c_286_n N_A_853_368#_c_803_n 0.0013074f $X=5.91 $Y=1.515 $X2=0 $Y2=0
cc_298 N_B1_c_287_n N_A_853_368#_c_803_n 0.0183565f $X=5.91 $Y=1.515 $X2=0 $Y2=0
cc_299 N_B1_c_291_n N_VPWR_c_879_n 5.74542e-19 $X=5.985 $Y=1.765 $X2=0 $Y2=0
cc_300 N_B1_c_288_n N_VPWR_c_884_n 0.00278257f $X=4.635 $Y=1.765 $X2=0 $Y2=0
cc_301 N_B1_c_289_n N_VPWR_c_884_n 0.00278257f $X=5.085 $Y=1.765 $X2=0 $Y2=0
cc_302 N_B1_c_290_n N_VPWR_c_884_n 0.00278257f $X=5.535 $Y=1.765 $X2=0 $Y2=0
cc_303 N_B1_c_291_n N_VPWR_c_884_n 0.0044313f $X=5.985 $Y=1.765 $X2=0 $Y2=0
cc_304 N_B1_c_288_n N_VPWR_c_878_n 0.00358623f $X=4.635 $Y=1.765 $X2=0 $Y2=0
cc_305 N_B1_c_289_n N_VPWR_c_878_n 0.00353822f $X=5.085 $Y=1.765 $X2=0 $Y2=0
cc_306 N_B1_c_290_n N_VPWR_c_878_n 0.00353822f $X=5.535 $Y=1.765 $X2=0 $Y2=0
cc_307 N_B1_c_291_n N_VPWR_c_878_n 0.00854206f $X=5.985 $Y=1.765 $X2=0 $Y2=0
cc_308 N_B1_M1011_g N_VGND_c_995_n 0.00434272f $X=4.02 $Y=0.74 $X2=0 $Y2=0
cc_309 N_B1_M1022_g N_VGND_c_995_n 0.00383152f $X=4.45 $Y=0.74 $X2=0 $Y2=0
cc_310 N_B1_M1011_g N_VGND_c_996_n 5.07239e-19 $X=4.02 $Y=0.74 $X2=0 $Y2=0
cc_311 N_B1_M1022_g N_VGND_c_996_n 0.0117017f $X=4.45 $Y=0.74 $X2=0 $Y2=0
cc_312 N_B1_M1011_g N_VGND_c_1005_n 0.00825037f $X=4.02 $Y=0.74 $X2=0 $Y2=0
cc_313 N_B1_M1022_g N_VGND_c_1005_n 0.0075754f $X=4.45 $Y=0.74 $X2=0 $Y2=0
cc_314 N_B1_M1011_g N_VGND_c_1008_n 0.00597094f $X=4.02 $Y=0.74 $X2=0 $Y2=0
cc_315 N_A1_M1032_g N_A2_M1005_g 0.019323f $X=7.79 $Y=0.74 $X2=0 $Y2=0
cc_316 N_A1_c_365_n N_A2_c_446_n 0.00834682f $X=7.785 $Y=1.765 $X2=0 $Y2=0
cc_317 A1 N_A2_c_450_n 0.0381127f $X=7.835 $Y=1.58 $X2=0 $Y2=0
cc_318 N_A1_c_361_n N_A2_c_450_n 3.59125e-19 $X=7.785 $Y=1.557 $X2=0 $Y2=0
cc_319 A1 N_A2_c_445_n 0.00345732f $X=7.835 $Y=1.58 $X2=0 $Y2=0
cc_320 N_A1_c_361_n N_A2_c_445_n 0.019348f $X=7.785 $Y=1.557 $X2=0 $Y2=0
cc_321 N_A1_M1008_g N_Y_c_593_n 0.00939349f $X=6.93 $Y=0.74 $X2=0 $Y2=0
cc_322 N_A1_M1029_g N_Y_c_593_n 0.0106855f $X=7.36 $Y=0.74 $X2=0 $Y2=0
cc_323 A1 N_Y_c_593_n 0.0330906f $X=7.835 $Y=1.58 $X2=0 $Y2=0
cc_324 N_A1_c_361_n N_Y_c_593_n 0.00218272f $X=7.785 $Y=1.557 $X2=0 $Y2=0
cc_325 N_A1_M1006_g N_Y_c_596_n 0.0123964f $X=6.5 $Y=0.74 $X2=0 $Y2=0
cc_326 A1 N_Y_c_596_n 0.0342389f $X=7.835 $Y=1.58 $X2=0 $Y2=0
cc_327 N_A1_c_361_n N_Y_c_596_n 0.00333888f $X=7.785 $Y=1.557 $X2=0 $Y2=0
cc_328 N_A1_M1006_g N_Y_c_597_n 0.0110564f $X=6.5 $Y=0.74 $X2=0 $Y2=0
cc_329 N_A1_M1008_g N_Y_c_597_n 0.00548858f $X=6.93 $Y=0.74 $X2=0 $Y2=0
cc_330 N_A1_M1029_g N_Y_c_597_n 6.61345e-19 $X=7.36 $Y=0.74 $X2=0 $Y2=0
cc_331 N_A1_c_361_n N_Y_c_597_n 0.00229127f $X=7.785 $Y=1.557 $X2=0 $Y2=0
cc_332 N_A1_M1008_g N_Y_c_598_n 5.30577e-19 $X=6.93 $Y=0.74 $X2=0 $Y2=0
cc_333 N_A1_M1029_g N_Y_c_598_n 0.0045607f $X=7.36 $Y=0.74 $X2=0 $Y2=0
cc_334 N_A1_M1032_g N_Y_c_598_n 0.00463734f $X=7.79 $Y=0.74 $X2=0 $Y2=0
cc_335 A1 N_Y_c_598_n 0.0218587f $X=7.835 $Y=1.58 $X2=0 $Y2=0
cc_336 N_A1_c_361_n N_Y_c_598_n 0.00221794f $X=7.785 $Y=1.557 $X2=0 $Y2=0
cc_337 N_A1_c_362_n N_A_474_368#_c_723_n 3.01915e-19 $X=6.435 $Y=1.765 $X2=0
+ $Y2=0
cc_338 N_A1_c_362_n N_A_853_368#_c_786_n 0.00557168f $X=6.435 $Y=1.765 $X2=0
+ $Y2=0
cc_339 N_A1_c_362_n N_A_853_368#_c_806_n 0.0152905f $X=6.435 $Y=1.765 $X2=0
+ $Y2=0
cc_340 N_A1_c_363_n N_A_853_368#_c_806_n 0.0126853f $X=6.885 $Y=1.765 $X2=0
+ $Y2=0
cc_341 A1 N_A_853_368#_c_806_n 0.0381145f $X=7.835 $Y=1.58 $X2=0 $Y2=0
cc_342 N_A1_c_361_n N_A_853_368#_c_806_n 0.00150005f $X=7.785 $Y=1.557 $X2=0
+ $Y2=0
cc_343 N_A1_c_363_n N_A_853_368#_c_787_n 0.00557168f $X=6.885 $Y=1.765 $X2=0
+ $Y2=0
cc_344 N_A1_c_364_n N_A_853_368#_c_787_n 0.00557168f $X=7.335 $Y=1.765 $X2=0
+ $Y2=0
cc_345 N_A1_c_364_n N_A_853_368#_c_812_n 0.0126853f $X=7.335 $Y=1.765 $X2=0
+ $Y2=0
cc_346 N_A1_c_365_n N_A_853_368#_c_812_n 0.0126853f $X=7.785 $Y=1.765 $X2=0
+ $Y2=0
cc_347 A1 N_A_853_368#_c_812_n 0.0477183f $X=7.835 $Y=1.58 $X2=0 $Y2=0
cc_348 N_A1_c_361_n N_A_853_368#_c_812_n 0.00150005f $X=7.785 $Y=1.557 $X2=0
+ $Y2=0
cc_349 N_A1_c_365_n N_A_853_368#_c_788_n 0.00557168f $X=7.785 $Y=1.765 $X2=0
+ $Y2=0
cc_350 A1 N_A_853_368#_c_817_n 0.0150275f $X=7.835 $Y=1.58 $X2=0 $Y2=0
cc_351 N_A1_c_361_n N_A_853_368#_c_817_n 0.00104296f $X=7.785 $Y=1.557 $X2=0
+ $Y2=0
cc_352 A1 N_A_853_368#_c_819_n 0.00972373f $X=7.835 $Y=1.58 $X2=0 $Y2=0
cc_353 N_A1_c_362_n N_VPWR_c_879_n 0.0117047f $X=6.435 $Y=1.765 $X2=0 $Y2=0
cc_354 N_A1_c_363_n N_VPWR_c_879_n 0.0116643f $X=6.885 $Y=1.765 $X2=0 $Y2=0
cc_355 N_A1_c_364_n N_VPWR_c_879_n 5.35985e-19 $X=7.335 $Y=1.765 $X2=0 $Y2=0
cc_356 N_A1_c_363_n N_VPWR_c_880_n 0.00413917f $X=6.885 $Y=1.765 $X2=0 $Y2=0
cc_357 N_A1_c_364_n N_VPWR_c_880_n 0.00413917f $X=7.335 $Y=1.765 $X2=0 $Y2=0
cc_358 N_A1_c_363_n N_VPWR_c_881_n 5.35985e-19 $X=6.885 $Y=1.765 $X2=0 $Y2=0
cc_359 N_A1_c_364_n N_VPWR_c_881_n 0.0116643f $X=7.335 $Y=1.765 $X2=0 $Y2=0
cc_360 N_A1_c_365_n N_VPWR_c_881_n 0.0116643f $X=7.785 $Y=1.765 $X2=0 $Y2=0
cc_361 N_A1_c_365_n N_VPWR_c_882_n 5.37805e-19 $X=7.785 $Y=1.765 $X2=0 $Y2=0
cc_362 N_A1_c_362_n N_VPWR_c_884_n 0.00413917f $X=6.435 $Y=1.765 $X2=0 $Y2=0
cc_363 N_A1_c_365_n N_VPWR_c_886_n 0.00413917f $X=7.785 $Y=1.765 $X2=0 $Y2=0
cc_364 N_A1_c_362_n N_VPWR_c_878_n 0.0081781f $X=6.435 $Y=1.765 $X2=0 $Y2=0
cc_365 N_A1_c_363_n N_VPWR_c_878_n 0.00817726f $X=6.885 $Y=1.765 $X2=0 $Y2=0
cc_366 N_A1_c_364_n N_VPWR_c_878_n 0.00817726f $X=7.335 $Y=1.765 $X2=0 $Y2=0
cc_367 N_A1_c_365_n N_VPWR_c_878_n 0.0081781f $X=7.785 $Y=1.765 $X2=0 $Y2=0
cc_368 N_A1_M1032_g N_VGND_c_997_n 6.35276e-19 $X=7.79 $Y=0.74 $X2=0 $Y2=0
cc_369 N_A1_M1006_g N_VGND_c_1002_n 0.00291649f $X=6.5 $Y=0.74 $X2=0 $Y2=0
cc_370 N_A1_M1008_g N_VGND_c_1002_n 0.00291649f $X=6.93 $Y=0.74 $X2=0 $Y2=0
cc_371 N_A1_M1029_g N_VGND_c_1002_n 0.00291649f $X=7.36 $Y=0.74 $X2=0 $Y2=0
cc_372 N_A1_M1032_g N_VGND_c_1002_n 0.00291649f $X=7.79 $Y=0.74 $X2=0 $Y2=0
cc_373 N_A1_M1006_g N_VGND_c_1005_n 0.0036412f $X=6.5 $Y=0.74 $X2=0 $Y2=0
cc_374 N_A1_M1008_g N_VGND_c_1005_n 0.00359121f $X=6.93 $Y=0.74 $X2=0 $Y2=0
cc_375 N_A1_M1029_g N_VGND_c_1005_n 0.00359121f $X=7.36 $Y=0.74 $X2=0 $Y2=0
cc_376 N_A1_M1032_g N_VGND_c_1005_n 0.00359219f $X=7.79 $Y=0.74 $X2=0 $Y2=0
cc_377 N_A1_M1029_g N_A_1228_74#_c_1096_n 0.010822f $X=7.36 $Y=0.74 $X2=0 $Y2=0
cc_378 N_A1_M1032_g N_A_1228_74#_c_1096_n 0.0142063f $X=7.79 $Y=0.74 $X2=0 $Y2=0
cc_379 N_A1_M1032_g N_A_1228_74#_c_1099_n 0.00174382f $X=7.79 $Y=0.74 $X2=0
+ $Y2=0
cc_380 A1 N_A_1228_74#_c_1099_n 0.0103694f $X=7.835 $Y=1.58 $X2=0 $Y2=0
cc_381 N_A1_M1006_g N_A_1228_74#_c_1104_n 0.0113038f $X=6.5 $Y=0.74 $X2=0 $Y2=0
cc_382 N_A1_M1008_g N_A_1228_74#_c_1104_n 0.0109057f $X=6.93 $Y=0.74 $X2=0 $Y2=0
cc_383 N_A2_c_446_n N_A_853_368#_c_788_n 0.00371619f $X=8.235 $Y=1.765 $X2=0
+ $Y2=0
cc_384 N_A2_c_446_n N_A_853_368#_c_821_n 0.0140291f $X=8.235 $Y=1.765 $X2=0
+ $Y2=0
cc_385 N_A2_c_447_n N_A_853_368#_c_821_n 0.0120074f $X=8.685 $Y=1.765 $X2=0
+ $Y2=0
cc_386 N_A2_c_450_n N_A_853_368#_c_821_n 0.0372325f $X=9.39 $Y=1.515 $X2=0 $Y2=0
cc_387 N_A2_c_445_n N_A_853_368#_c_821_n 0.00130859f $X=9.51 $Y=1.557 $X2=0
+ $Y2=0
cc_388 N_A2_c_446_n N_A_853_368#_c_789_n 6.69308e-19 $X=8.235 $Y=1.765 $X2=0
+ $Y2=0
cc_389 N_A2_c_447_n N_A_853_368#_c_789_n 0.010609f $X=8.685 $Y=1.765 $X2=0 $Y2=0
cc_390 N_A2_c_448_n N_A_853_368#_c_789_n 0.010609f $X=9.135 $Y=1.765 $X2=0 $Y2=0
cc_391 N_A2_c_449_n N_A_853_368#_c_789_n 6.69308e-19 $X=9.585 $Y=1.765 $X2=0
+ $Y2=0
cc_392 N_A2_c_448_n N_A_853_368#_c_829_n 0.0120074f $X=9.135 $Y=1.765 $X2=0
+ $Y2=0
cc_393 N_A2_c_449_n N_A_853_368#_c_829_n 0.015731f $X=9.585 $Y=1.765 $X2=0 $Y2=0
cc_394 N_A2_c_450_n N_A_853_368#_c_829_n 0.0328547f $X=9.39 $Y=1.515 $X2=0 $Y2=0
cc_395 N_A2_c_445_n N_A_853_368#_c_829_n 0.00130859f $X=9.51 $Y=1.557 $X2=0
+ $Y2=0
cc_396 N_A2_c_449_n N_A_853_368#_c_790_n 0.00314968f $X=9.585 $Y=1.765 $X2=0
+ $Y2=0
cc_397 N_A2_c_449_n N_A_853_368#_c_791_n 0.00526798f $X=9.585 $Y=1.765 $X2=0
+ $Y2=0
cc_398 N_A2_c_447_n N_A_853_368#_c_835_n 4.27055e-19 $X=8.685 $Y=1.765 $X2=0
+ $Y2=0
cc_399 N_A2_c_448_n N_A_853_368#_c_835_n 4.27055e-19 $X=9.135 $Y=1.765 $X2=0
+ $Y2=0
cc_400 N_A2_c_450_n N_A_853_368#_c_835_n 0.0237598f $X=9.39 $Y=1.515 $X2=0 $Y2=0
cc_401 N_A2_c_445_n N_A_853_368#_c_835_n 0.00144162f $X=9.51 $Y=1.557 $X2=0
+ $Y2=0
cc_402 N_A2_c_446_n N_VPWR_c_881_n 5.35985e-19 $X=8.235 $Y=1.765 $X2=0 $Y2=0
cc_403 N_A2_c_446_n N_VPWR_c_882_n 0.0106464f $X=8.235 $Y=1.765 $X2=0 $Y2=0
cc_404 N_A2_c_447_n N_VPWR_c_882_n 0.00526215f $X=8.685 $Y=1.765 $X2=0 $Y2=0
cc_405 N_A2_c_448_n N_VPWR_c_883_n 0.00526215f $X=9.135 $Y=1.765 $X2=0 $Y2=0
cc_406 N_A2_c_449_n N_VPWR_c_883_n 0.0135832f $X=9.585 $Y=1.765 $X2=0 $Y2=0
cc_407 N_A2_c_446_n N_VPWR_c_886_n 0.00413917f $X=8.235 $Y=1.765 $X2=0 $Y2=0
cc_408 N_A2_c_447_n N_VPWR_c_887_n 0.00445602f $X=8.685 $Y=1.765 $X2=0 $Y2=0
cc_409 N_A2_c_448_n N_VPWR_c_887_n 0.00445602f $X=9.135 $Y=1.765 $X2=0 $Y2=0
cc_410 N_A2_c_449_n N_VPWR_c_888_n 0.00413917f $X=9.585 $Y=1.765 $X2=0 $Y2=0
cc_411 N_A2_c_446_n N_VPWR_c_878_n 0.0081781f $X=8.235 $Y=1.765 $X2=0 $Y2=0
cc_412 N_A2_c_447_n N_VPWR_c_878_n 0.00857589f $X=8.685 $Y=1.765 $X2=0 $Y2=0
cc_413 N_A2_c_448_n N_VPWR_c_878_n 0.00857589f $X=9.135 $Y=1.765 $X2=0 $Y2=0
cc_414 N_A2_c_449_n N_VPWR_c_878_n 0.00821187f $X=9.585 $Y=1.765 $X2=0 $Y2=0
cc_415 N_A2_M1005_g N_VGND_c_997_n 0.010782f $X=8.22 $Y=0.74 $X2=0 $Y2=0
cc_416 N_A2_M1018_g N_VGND_c_997_n 0.0106755f $X=8.65 $Y=0.74 $X2=0 $Y2=0
cc_417 N_A2_M1024_g N_VGND_c_997_n 4.71636e-19 $X=9.08 $Y=0.74 $X2=0 $Y2=0
cc_418 N_A2_M1018_g N_VGND_c_998_n 4.71636e-19 $X=8.65 $Y=0.74 $X2=0 $Y2=0
cc_419 N_A2_M1024_g N_VGND_c_998_n 0.0106755f $X=9.08 $Y=0.74 $X2=0 $Y2=0
cc_420 N_A2_M1027_g N_VGND_c_998_n 0.0137191f $X=9.51 $Y=0.74 $X2=0 $Y2=0
cc_421 N_A2_M1005_g N_VGND_c_1002_n 0.00383152f $X=8.22 $Y=0.74 $X2=0 $Y2=0
cc_422 N_A2_M1018_g N_VGND_c_1003_n 0.00383152f $X=8.65 $Y=0.74 $X2=0 $Y2=0
cc_423 N_A2_M1024_g N_VGND_c_1003_n 0.00383152f $X=9.08 $Y=0.74 $X2=0 $Y2=0
cc_424 N_A2_M1027_g N_VGND_c_1004_n 0.00383152f $X=9.51 $Y=0.74 $X2=0 $Y2=0
cc_425 N_A2_M1005_g N_VGND_c_1005_n 0.00757637f $X=8.22 $Y=0.74 $X2=0 $Y2=0
cc_426 N_A2_M1018_g N_VGND_c_1005_n 0.0075754f $X=8.65 $Y=0.74 $X2=0 $Y2=0
cc_427 N_A2_M1024_g N_VGND_c_1005_n 0.0075754f $X=9.08 $Y=0.74 $X2=0 $Y2=0
cc_428 N_A2_M1027_g N_VGND_c_1005_n 0.00761428f $X=9.51 $Y=0.74 $X2=0 $Y2=0
cc_429 N_A2_M1005_g N_A_1228_74#_c_1098_n 0.0147012f $X=8.22 $Y=0.74 $X2=0 $Y2=0
cc_430 N_A2_M1018_g N_A_1228_74#_c_1098_n 0.0130453f $X=8.65 $Y=0.74 $X2=0 $Y2=0
cc_431 N_A2_c_450_n N_A_1228_74#_c_1098_n 0.0431743f $X=9.39 $Y=1.515 $X2=0
+ $Y2=0
cc_432 N_A2_c_445_n N_A_1228_74#_c_1098_n 0.00224206f $X=9.51 $Y=1.557 $X2=0
+ $Y2=0
cc_433 N_A2_M1018_g N_A_1228_74#_c_1100_n 3.92313e-19 $X=8.65 $Y=0.74 $X2=0
+ $Y2=0
cc_434 N_A2_M1024_g N_A_1228_74#_c_1100_n 3.92313e-19 $X=9.08 $Y=0.74 $X2=0
+ $Y2=0
cc_435 N_A2_M1024_g N_A_1228_74#_c_1101_n 0.0130918f $X=9.08 $Y=0.74 $X2=0 $Y2=0
cc_436 N_A2_M1027_g N_A_1228_74#_c_1101_n 0.0145697f $X=9.51 $Y=0.74 $X2=0 $Y2=0
cc_437 N_A2_c_450_n N_A_1228_74#_c_1101_n 0.0453632f $X=9.39 $Y=1.515 $X2=0
+ $Y2=0
cc_438 N_A2_c_445_n N_A_1228_74#_c_1101_n 0.00615819f $X=9.51 $Y=1.557 $X2=0
+ $Y2=0
cc_439 N_A2_M1027_g N_A_1228_74#_c_1102_n 0.00159319f $X=9.51 $Y=0.74 $X2=0
+ $Y2=0
cc_440 N_A2_c_450_n N_A_1228_74#_c_1106_n 0.0146029f $X=9.39 $Y=1.515 $X2=0
+ $Y2=0
cc_441 N_A2_c_445_n N_A_1228_74#_c_1106_n 0.00232957f $X=9.51 $Y=1.557 $X2=0
+ $Y2=0
cc_442 N_A_29_368#_c_518_n N_Y_M1000_d 0.00197722f $X=1.085 $Y=2.99 $X2=0 $Y2=0
cc_443 N_A_29_368#_c_520_n N_Y_M1002_d 0.00218679f $X=1.905 $Y=2.99 $X2=0 $Y2=0
cc_444 N_A_29_368#_M1000_s N_Y_c_600_n 2.67089e-19 $X=0.145 $Y=1.84 $X2=0 $Y2=0
cc_445 N_A_29_368#_c_517_n N_Y_c_610_n 0.0452595f $X=0.27 $Y=2.225 $X2=0 $Y2=0
cc_446 N_A_29_368#_c_518_n N_Y_c_610_n 0.0160777f $X=1.085 $Y=2.99 $X2=0 $Y2=0
cc_447 N_A_29_368#_c_526_n N_Y_c_610_n 0.0439674f $X=1.17 $Y=2.225 $X2=0 $Y2=0
cc_448 N_A_29_368#_M1001_s N_Y_c_601_n 0.00247267f $X=1.02 $Y=1.84 $X2=0 $Y2=0
cc_449 N_A_29_368#_c_526_n N_Y_c_601_n 0.0136682f $X=1.17 $Y=2.225 $X2=0 $Y2=0
cc_450 N_A_29_368#_c_526_n N_Y_c_618_n 0.0430411f $X=1.17 $Y=2.225 $X2=0 $Y2=0
cc_451 N_A_29_368#_c_520_n N_Y_c_618_n 0.0144323f $X=1.905 $Y=2.99 $X2=0 $Y2=0
cc_452 N_A_29_368#_c_530_n N_Y_c_618_n 0.0121024f $X=2.07 $Y=2.12 $X2=0 $Y2=0
cc_453 N_A_29_368#_c_531_n N_Y_c_618_n 0.0412035f $X=2.07 $Y=2.815 $X2=0 $Y2=0
cc_454 N_A_29_368#_c_522_n N_Y_c_591_n 0.010505f $X=3.87 $Y=2.05 $X2=0 $Y2=0
cc_455 N_A_29_368#_M1000_s N_Y_c_604_n 0.00253425f $X=0.145 $Y=1.84 $X2=0 $Y2=0
cc_456 N_A_29_368#_c_517_n N_Y_c_604_n 0.0206709f $X=0.27 $Y=2.225 $X2=0 $Y2=0
cc_457 N_A_29_368#_c_537_n N_A_474_368#_M1007_d 0.00384138f $X=2.855 $Y=2.035
+ $X2=-0.19 $Y2=1.66
cc_458 N_A_29_368#_c_541_n N_A_474_368#_M1012_d 0.00354874f $X=3.705 $Y=2.035
+ $X2=0 $Y2=0
cc_459 N_A_29_368#_c_531_n N_A_474_368#_c_726_n 0.0411694f $X=2.07 $Y=2.815
+ $X2=0 $Y2=0
cc_460 N_A_29_368#_c_537_n N_A_474_368#_c_726_n 0.0154248f $X=2.855 $Y=2.035
+ $X2=0 $Y2=0
cc_461 N_A_29_368#_M1009_s N_A_474_368#_c_720_n 0.00197722f $X=2.82 $Y=1.84
+ $X2=0 $Y2=0
cc_462 N_A_29_368#_c_572_p N_A_474_368#_c_720_n 0.014157f $X=2.97 $Y=2.57 $X2=0
+ $Y2=0
cc_463 N_A_29_368#_c_520_n N_A_474_368#_c_721_n 0.0132987f $X=1.905 $Y=2.99
+ $X2=0 $Y2=0
cc_464 N_A_29_368#_c_541_n N_A_474_368#_c_732_n 0.0171813f $X=3.705 $Y=2.035
+ $X2=0 $Y2=0
cc_465 N_A_29_368#_M1014_s N_A_474_368#_c_722_n 0.00260133f $X=3.72 $Y=1.84
+ $X2=0 $Y2=0
cc_466 N_A_29_368#_c_522_n N_A_474_368#_c_722_n 0.0196739f $X=3.87 $Y=2.05 $X2=0
+ $Y2=0
cc_467 N_A_29_368#_c_522_n N_A_853_368#_c_784_n 0.0137127f $X=3.87 $Y=2.05 $X2=0
+ $Y2=0
cc_468 N_A_29_368#_c_522_n N_A_853_368#_c_785_n 0.0430074f $X=3.87 $Y=2.05 $X2=0
+ $Y2=0
cc_469 N_A_29_368#_c_518_n N_VPWR_c_884_n 0.0460938f $X=1.085 $Y=2.99 $X2=0
+ $Y2=0
cc_470 N_A_29_368#_c_519_n N_VPWR_c_884_n 0.0178855f $X=0.355 $Y=2.99 $X2=0
+ $Y2=0
cc_471 N_A_29_368#_c_520_n N_VPWR_c_884_n 0.0645381f $X=1.905 $Y=2.99 $X2=0
+ $Y2=0
cc_472 N_A_29_368#_c_521_n N_VPWR_c_884_n 0.0121867f $X=1.17 $Y=2.99 $X2=0 $Y2=0
cc_473 N_A_29_368#_c_518_n N_VPWR_c_878_n 0.0260732f $X=1.085 $Y=2.99 $X2=0
+ $Y2=0
cc_474 N_A_29_368#_c_519_n N_VPWR_c_878_n 0.00971414f $X=0.355 $Y=2.99 $X2=0
+ $Y2=0
cc_475 N_A_29_368#_c_520_n N_VPWR_c_878_n 0.0358265f $X=1.905 $Y=2.99 $X2=0
+ $Y2=0
cc_476 N_A_29_368#_c_521_n N_VPWR_c_878_n 0.00660921f $X=1.17 $Y=2.99 $X2=0
+ $Y2=0
cc_477 N_Y_c_587_n N_VGND_M1017_s 0.00473729f $X=1.53 $Y=0.925 $X2=-0.19
+ $Y2=-0.245
cc_478 N_Y_c_623_n N_VGND_M1028_s 0.00807452f $X=2.39 $Y=0.925 $X2=0 $Y2=0
cc_479 N_Y_c_591_n N_VGND_M1025_s 0.0158527f $X=4.07 $Y=1.095 $X2=0 $Y2=0
cc_480 N_Y_c_596_n N_VGND_M1022_s 0.00285432f $X=6.55 $Y=0.975 $X2=0 $Y2=0
cc_481 N_Y_c_587_n N_VGND_c_993_n 0.0215198f $X=1.53 $Y=0.925 $X2=0 $Y2=0
cc_482 N_Y_c_589_n N_VGND_c_993_n 0.0135953f $X=1.615 $Y=0.495 $X2=0 $Y2=0
cc_483 N_Y_c_589_n N_VGND_c_994_n 0.0135953f $X=1.615 $Y=0.495 $X2=0 $Y2=0
cc_484 N_Y_c_623_n N_VGND_c_994_n 0.0167019f $X=2.39 $Y=0.925 $X2=0 $Y2=0
cc_485 N_Y_c_590_n N_VGND_c_994_n 0.0121972f $X=2.475 $Y=0.515 $X2=0 $Y2=0
cc_486 N_Y_c_592_n N_VGND_c_995_n 0.0109942f $X=4.235 $Y=0.515 $X2=0 $Y2=0
cc_487 N_Y_c_592_n N_VGND_c_996_n 0.0170358f $X=4.235 $Y=0.515 $X2=0 $Y2=0
cc_488 N_Y_c_596_n N_VGND_c_996_n 0.022285f $X=6.55 $Y=0.975 $X2=0 $Y2=0
cc_489 N_Y_c_589_n N_VGND_c_999_n 0.00814895f $X=1.615 $Y=0.495 $X2=0 $Y2=0
cc_490 N_Y_c_587_n N_VGND_c_1005_n 0.0293519f $X=1.53 $Y=0.925 $X2=0 $Y2=0
cc_491 N_Y_c_588_n N_VGND_c_1005_n 0.00906892f $X=0.355 $Y=0.925 $X2=0 $Y2=0
cc_492 N_Y_c_589_n N_VGND_c_1005_n 0.00627841f $X=1.615 $Y=0.495 $X2=0 $Y2=0
cc_493 N_Y_c_623_n N_VGND_c_1005_n 0.0116543f $X=2.39 $Y=0.925 $X2=0 $Y2=0
cc_494 N_Y_c_590_n N_VGND_c_1005_n 0.00904371f $X=2.475 $Y=0.515 $X2=0 $Y2=0
cc_495 N_Y_c_592_n N_VGND_c_1005_n 0.00904371f $X=4.235 $Y=0.515 $X2=0 $Y2=0
cc_496 N_Y_c_590_n N_VGND_c_1007_n 0.0109942f $X=2.475 $Y=0.515 $X2=0 $Y2=0
cc_497 N_Y_c_590_n N_VGND_c_1008_n 0.0185534f $X=2.475 $Y=0.515 $X2=0 $Y2=0
cc_498 N_Y_c_591_n N_VGND_c_1008_n 0.0863478f $X=4.07 $Y=1.095 $X2=0 $Y2=0
cc_499 N_Y_c_592_n N_VGND_c_1008_n 0.0185534f $X=4.235 $Y=0.515 $X2=0 $Y2=0
cc_500 N_Y_c_596_n N_A_1228_74#_M1006_d 0.00392596f $X=6.55 $Y=0.975 $X2=-0.19
+ $Y2=-0.245
cc_501 N_Y_c_593_n N_A_1228_74#_M1008_d 0.00205565f $X=7.41 $Y=1.022 $X2=0 $Y2=0
cc_502 N_Y_M1029_s N_A_1228_74#_c_1096_n 0.00178571f $X=7.435 $Y=0.37 $X2=0
+ $Y2=0
cc_503 N_Y_c_593_n N_A_1228_74#_c_1096_n 0.00540301f $X=7.41 $Y=1.022 $X2=0
+ $Y2=0
cc_504 N_Y_c_598_n N_A_1228_74#_c_1096_n 0.0161432f $X=7.575 $Y=0.95 $X2=0 $Y2=0
cc_505 N_Y_c_598_n N_A_1228_74#_c_1099_n 0.00517071f $X=7.575 $Y=0.95 $X2=0
+ $Y2=0
cc_506 N_Y_c_596_n N_A_1228_74#_c_1103_n 0.0128721f $X=6.55 $Y=0.975 $X2=0 $Y2=0
cc_507 N_Y_M1006_s N_A_1228_74#_c_1104_n 0.00179007f $X=6.575 $Y=0.37 $X2=0
+ $Y2=0
cc_508 N_Y_c_593_n N_A_1228_74#_c_1104_n 0.00538156f $X=7.41 $Y=1.022 $X2=0
+ $Y2=0
cc_509 N_Y_c_596_n N_A_1228_74#_c_1104_n 0.00465091f $X=6.55 $Y=0.975 $X2=0
+ $Y2=0
cc_510 N_Y_c_597_n N_A_1228_74#_c_1104_n 0.0163588f $X=6.88 $Y=0.975 $X2=0 $Y2=0
cc_511 N_Y_c_593_n N_A_1228_74#_c_1105_n 0.0101598f $X=7.41 $Y=1.022 $X2=0 $Y2=0
cc_512 N_A_474_368#_c_722_n N_A_853_368#_M1004_d 0.00287371f $X=4.695 $Y=2.99
+ $X2=-0.19 $Y2=1.66
cc_513 N_A_474_368#_c_723_n N_A_853_368#_M1010_d 0.00197722f $X=5.595 $Y=2.99
+ $X2=0 $Y2=0
cc_514 N_A_474_368#_c_722_n N_A_853_368#_c_785_n 0.019616f $X=4.695 $Y=2.99
+ $X2=0 $Y2=0
cc_515 N_A_474_368#_M1004_s N_A_853_368#_c_794_n 0.00359365f $X=4.71 $Y=1.84
+ $X2=0 $Y2=0
cc_516 N_A_474_368#_c_739_n N_A_853_368#_c_794_n 0.0171813f $X=4.86 $Y=2.405
+ $X2=0 $Y2=0
cc_517 N_A_474_368#_c_723_n N_A_853_368#_c_846_n 0.014157f $X=5.595 $Y=2.99
+ $X2=0 $Y2=0
cc_518 N_A_474_368#_M1013_s N_A_853_368#_c_798_n 0.00359365f $X=5.61 $Y=1.84
+ $X2=0 $Y2=0
cc_519 N_A_474_368#_c_745_n N_A_853_368#_c_798_n 0.0171813f $X=5.76 $Y=2.405
+ $X2=0 $Y2=0
cc_520 N_A_474_368#_c_723_n N_A_853_368#_c_786_n 0.00522251f $X=5.595 $Y=2.99
+ $X2=0 $Y2=0
cc_521 N_A_474_368#_c_745_n N_A_853_368#_c_786_n 0.0400262f $X=5.76 $Y=2.405
+ $X2=0 $Y2=0
cc_522 N_A_474_368#_c_723_n N_VPWR_c_879_n 0.00279034f $X=5.595 $Y=2.99 $X2=0
+ $Y2=0
cc_523 N_A_474_368#_c_720_n N_VPWR_c_884_n 0.03588f $X=3.255 $Y=2.99 $X2=0 $Y2=0
cc_524 N_A_474_368#_c_721_n N_VPWR_c_884_n 0.017869f $X=2.685 $Y=2.99 $X2=0
+ $Y2=0
cc_525 N_A_474_368#_c_722_n N_VPWR_c_884_n 0.0706659f $X=4.695 $Y=2.99 $X2=0
+ $Y2=0
cc_526 N_A_474_368#_c_723_n N_VPWR_c_884_n 0.0594312f $X=5.595 $Y=2.99 $X2=0
+ $Y2=0
cc_527 N_A_474_368#_c_724_n N_VPWR_c_884_n 0.0235512f $X=3.42 $Y=2.99 $X2=0
+ $Y2=0
cc_528 N_A_474_368#_c_725_n N_VPWR_c_884_n 0.0235512f $X=4.86 $Y=2.99 $X2=0
+ $Y2=0
cc_529 N_A_474_368#_c_720_n N_VPWR_c_878_n 0.0201952f $X=3.255 $Y=2.99 $X2=0
+ $Y2=0
cc_530 N_A_474_368#_c_721_n N_VPWR_c_878_n 0.00965079f $X=2.685 $Y=2.99 $X2=0
+ $Y2=0
cc_531 N_A_474_368#_c_722_n N_VPWR_c_878_n 0.040498f $X=4.695 $Y=2.99 $X2=0
+ $Y2=0
cc_532 N_A_474_368#_c_723_n N_VPWR_c_878_n 0.0328875f $X=5.595 $Y=2.99 $X2=0
+ $Y2=0
cc_533 N_A_474_368#_c_724_n N_VPWR_c_878_n 0.0126924f $X=3.42 $Y=2.99 $X2=0
+ $Y2=0
cc_534 N_A_474_368#_c_725_n N_VPWR_c_878_n 0.0126924f $X=4.86 $Y=2.99 $X2=0
+ $Y2=0
cc_535 N_A_853_368#_c_806_n N_VPWR_M1016_d 0.00359365f $X=7.025 $Y=2.035
+ $X2=-0.19 $Y2=1.66
cc_536 N_A_853_368#_c_812_n N_VPWR_M1020_d 0.00359365f $X=7.925 $Y=2.035 $X2=0
+ $Y2=0
cc_537 N_A_853_368#_c_821_n N_VPWR_M1023_d 0.00384138f $X=8.745 $Y=2.035 $X2=0
+ $Y2=0
cc_538 N_A_853_368#_c_829_n N_VPWR_M1031_d 0.00384138f $X=9.725 $Y=2.035 $X2=0
+ $Y2=0
cc_539 N_A_853_368#_c_786_n N_VPWR_c_879_n 0.0449718f $X=6.21 $Y=2.43 $X2=0
+ $Y2=0
cc_540 N_A_853_368#_c_806_n N_VPWR_c_879_n 0.0171813f $X=7.025 $Y=2.035 $X2=0
+ $Y2=0
cc_541 N_A_853_368#_c_787_n N_VPWR_c_879_n 0.0449718f $X=7.11 $Y=2.43 $X2=0
+ $Y2=0
cc_542 N_A_853_368#_c_787_n N_VPWR_c_880_n 0.00749631f $X=7.11 $Y=2.43 $X2=0
+ $Y2=0
cc_543 N_A_853_368#_c_787_n N_VPWR_c_881_n 0.0449718f $X=7.11 $Y=2.43 $X2=0
+ $Y2=0
cc_544 N_A_853_368#_c_812_n N_VPWR_c_881_n 0.0171813f $X=7.925 $Y=2.035 $X2=0
+ $Y2=0
cc_545 N_A_853_368#_c_788_n N_VPWR_c_881_n 0.0449718f $X=8.01 $Y=2.43 $X2=0
+ $Y2=0
cc_546 N_A_853_368#_c_788_n N_VPWR_c_882_n 0.0440249f $X=8.01 $Y=2.43 $X2=0
+ $Y2=0
cc_547 N_A_853_368#_c_821_n N_VPWR_c_882_n 0.0154248f $X=8.745 $Y=2.035 $X2=0
+ $Y2=0
cc_548 N_A_853_368#_c_789_n N_VPWR_c_882_n 0.0462948f $X=8.91 $Y=2.815 $X2=0
+ $Y2=0
cc_549 N_A_853_368#_c_789_n N_VPWR_c_883_n 0.0462948f $X=8.91 $Y=2.815 $X2=0
+ $Y2=0
cc_550 N_A_853_368#_c_829_n N_VPWR_c_883_n 0.0154248f $X=9.725 $Y=2.035 $X2=0
+ $Y2=0
cc_551 N_A_853_368#_c_791_n N_VPWR_c_883_n 0.0453479f $X=9.81 $Y=2.4 $X2=0 $Y2=0
cc_552 N_A_853_368#_c_786_n N_VPWR_c_884_n 0.00749631f $X=6.21 $Y=2.43 $X2=0
+ $Y2=0
cc_553 N_A_853_368#_c_788_n N_VPWR_c_886_n 0.00749631f $X=8.01 $Y=2.43 $X2=0
+ $Y2=0
cc_554 N_A_853_368#_c_789_n N_VPWR_c_887_n 0.014552f $X=8.91 $Y=2.815 $X2=0
+ $Y2=0
cc_555 N_A_853_368#_c_791_n N_VPWR_c_888_n 0.011066f $X=9.81 $Y=2.4 $X2=0 $Y2=0
cc_556 N_A_853_368#_c_786_n N_VPWR_c_878_n 0.0062048f $X=6.21 $Y=2.43 $X2=0
+ $Y2=0
cc_557 N_A_853_368#_c_787_n N_VPWR_c_878_n 0.0062048f $X=7.11 $Y=2.43 $X2=0
+ $Y2=0
cc_558 N_A_853_368#_c_788_n N_VPWR_c_878_n 0.0062048f $X=8.01 $Y=2.43 $X2=0
+ $Y2=0
cc_559 N_A_853_368#_c_789_n N_VPWR_c_878_n 0.0119791f $X=8.91 $Y=2.815 $X2=0
+ $Y2=0
cc_560 N_A_853_368#_c_791_n N_VPWR_c_878_n 0.00915947f $X=9.81 $Y=2.4 $X2=0
+ $Y2=0
cc_561 N_A_853_368#_c_790_n N_A_1228_74#_c_1101_n 0.00609927f $X=9.85 $Y=2.12
+ $X2=0 $Y2=0
cc_562 N_VGND_c_997_n N_A_1228_74#_c_1097_n 0.00985092f $X=8.435 $Y=0.675 $X2=0
+ $Y2=0
cc_563 N_VGND_c_1002_n N_A_1228_74#_c_1097_n 0.00758556f $X=8.27 $Y=0 $X2=0
+ $Y2=0
cc_564 N_VGND_c_1005_n N_A_1228_74#_c_1097_n 0.00627867f $X=9.84 $Y=0 $X2=0
+ $Y2=0
cc_565 N_VGND_M1005_s N_A_1228_74#_c_1098_n 0.00176461f $X=8.295 $Y=0.37 $X2=0
+ $Y2=0
cc_566 N_VGND_c_997_n N_A_1228_74#_c_1098_n 0.0170777f $X=8.435 $Y=0.675 $X2=0
+ $Y2=0
cc_567 N_VGND_c_997_n N_A_1228_74#_c_1100_n 0.0182488f $X=8.435 $Y=0.675 $X2=0
+ $Y2=0
cc_568 N_VGND_c_998_n N_A_1228_74#_c_1100_n 0.0182488f $X=9.295 $Y=0.675 $X2=0
+ $Y2=0
cc_569 N_VGND_c_1003_n N_A_1228_74#_c_1100_n 0.00749631f $X=9.13 $Y=0 $X2=0
+ $Y2=0
cc_570 N_VGND_c_1005_n N_A_1228_74#_c_1100_n 0.0062048f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_571 N_VGND_M1024_s N_A_1228_74#_c_1101_n 0.00176461f $X=9.155 $Y=0.37 $X2=0
+ $Y2=0
cc_572 N_VGND_c_998_n N_A_1228_74#_c_1101_n 0.0170777f $X=9.295 $Y=0.675 $X2=0
+ $Y2=0
cc_573 N_VGND_c_998_n N_A_1228_74#_c_1102_n 0.0182902f $X=9.295 $Y=0.675 $X2=0
+ $Y2=0
cc_574 N_VGND_c_1004_n N_A_1228_74#_c_1102_n 0.011066f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_575 N_VGND_c_1005_n N_A_1228_74#_c_1102_n 0.00915947f $X=9.84 $Y=0 $X2=0
+ $Y2=0
cc_576 N_VGND_c_1002_n N_A_1228_74#_c_1103_n 0.0732673f $X=8.27 $Y=0 $X2=0 $Y2=0
cc_577 N_VGND_c_1005_n N_A_1228_74#_c_1103_n 0.0615998f $X=9.84 $Y=0 $X2=0 $Y2=0
