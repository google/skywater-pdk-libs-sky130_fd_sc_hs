* File: sky130_fd_sc_hs__o32ai_2.pex.spice
* Created: Tue Sep  1 20:18:58 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HS__O32AI_2%B2 3 5 7 10 12 14 15 16 17 26
c46 17 0 1.22193e-19 $X=1.2 $Y=1.665
c47 12 0 1.88367e-19 $X=0.955 $Y=1.765
r48 26 27 3.8871 $w=3.72e-07 $l=3e-08 $layer=POLY_cond $X=0.925 $Y=1.557
+ $X2=0.955 $Y2=1.557
r49 24 26 11.6613 $w=3.72e-07 $l=9e-08 $layer=POLY_cond $X=0.835 $Y=1.557
+ $X2=0.925 $Y2=1.557
r50 24 25 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.835
+ $Y=1.515 $X2=0.835 $Y2=1.515
r51 22 24 42.7581 $w=3.72e-07 $l=3.3e-07 $layer=POLY_cond $X=0.505 $Y=1.557
+ $X2=0.835 $Y2=1.557
r52 21 22 1.2957 $w=3.72e-07 $l=1e-08 $layer=POLY_cond $X=0.495 $Y=1.557
+ $X2=0.505 $Y2=1.557
r53 17 25 9.78236 $w=4.28e-07 $l=3.65e-07 $layer=LI1_cond $X=1.2 $Y=1.565
+ $X2=0.835 $Y2=1.565
r54 16 25 3.08211 $w=4.28e-07 $l=1.15e-07 $layer=LI1_cond $X=0.72 $Y=1.565
+ $X2=0.835 $Y2=1.565
r55 15 16 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=0.24 $Y=1.565
+ $X2=0.72 $Y2=1.565
r56 12 27 24.0971 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=0.955 $Y=1.765
+ $X2=0.955 $Y2=1.557
r57 12 14 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.955 $Y=1.765
+ $X2=0.955 $Y2=2.4
r58 8 26 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.925 $Y=1.35
+ $X2=0.925 $Y2=1.557
r59 8 10 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=0.925 $Y=1.35
+ $X2=0.925 $Y2=0.74
r60 5 22 24.0971 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=0.505 $Y=1.765
+ $X2=0.505 $Y2=1.557
r61 5 7 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.505 $Y=1.765
+ $X2=0.505 $Y2=2.4
r62 1 21 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.495 $Y=1.35
+ $X2=0.495 $Y2=1.557
r63 1 3 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=0.495 $Y=1.35
+ $X2=0.495 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HS__O32AI_2%B1 1 3 6 8 10 13 15 21 22
c55 1 0 1.22193e-19 $X=1.405 $Y=1.765
r56 22 23 9.37222 $w=3.6e-07 $l=7e-08 $layer=POLY_cond $X=1.855 $Y=1.557
+ $X2=1.925 $Y2=1.557
r57 20 22 27.4472 $w=3.6e-07 $l=2.05e-07 $layer=POLY_cond $X=1.65 $Y=1.557
+ $X2=1.855 $Y2=1.557
r58 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.65
+ $Y=1.515 $X2=1.65 $Y2=1.515
r59 18 20 30.125 $w=3.6e-07 $l=2.25e-07 $layer=POLY_cond $X=1.425 $Y=1.557
+ $X2=1.65 $Y2=1.557
r60 17 18 2.67778 $w=3.6e-07 $l=2e-08 $layer=POLY_cond $X=1.405 $Y=1.557
+ $X2=1.425 $Y2=1.557
r61 15 21 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=1.65 $Y=1.665
+ $X2=1.65 $Y2=1.515
r62 11 23 23.3057 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.925 $Y=1.35
+ $X2=1.925 $Y2=1.557
r63 11 13 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.925 $Y=1.35
+ $X2=1.925 $Y2=0.74
r64 8 22 23.3057 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=1.855 $Y=1.765
+ $X2=1.855 $Y2=1.557
r65 8 10 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.855 $Y=1.765
+ $X2=1.855 $Y2=2.4
r66 4 18 23.3057 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.425 $Y=1.35
+ $X2=1.425 $Y2=1.557
r67 4 6 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.425 $Y=1.35
+ $X2=1.425 $Y2=0.74
r68 1 17 23.3057 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=1.405 $Y=1.765
+ $X2=1.405 $Y2=1.557
r69 1 3 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.405 $Y=1.765
+ $X2=1.405 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_HS__O32AI_2%A3 3 5 7 10 12 14 15 16 24
c60 12 0 1.57212e-19 $X=3.315 $Y=1.765
c61 5 0 1.68844e-19 $X=2.865 $Y=1.765
r62 24 25 8.35838 $w=3.46e-07 $l=6e-08 $layer=POLY_cond $X=3.255 $Y=1.557
+ $X2=3.315 $Y2=1.557
r63 23 24 54.3295 $w=3.46e-07 $l=3.9e-07 $layer=POLY_cond $X=2.865 $Y=1.557
+ $X2=3.255 $Y2=1.557
r64 21 23 48.7572 $w=3.46e-07 $l=3.5e-07 $layer=POLY_cond $X=2.515 $Y=1.557
+ $X2=2.865 $Y2=1.557
r65 21 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.515
+ $Y=1.515 $X2=2.515 $Y2=1.515
r66 19 21 12.5376 $w=3.46e-07 $l=9e-08 $layer=POLY_cond $X=2.425 $Y=1.557
+ $X2=2.515 $Y2=1.557
r67 16 22 3.35013 $w=4.28e-07 $l=1.25e-07 $layer=LI1_cond $X=2.64 $Y=1.565
+ $X2=2.515 $Y2=1.565
r68 15 22 9.51435 $w=4.28e-07 $l=3.55e-07 $layer=LI1_cond $X=2.16 $Y=1.565
+ $X2=2.515 $Y2=1.565
r69 12 25 22.3532 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=3.315 $Y=1.765
+ $X2=3.315 $Y2=1.557
r70 12 14 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.315 $Y=1.765
+ $X2=3.315 $Y2=2.4
r71 8 24 22.3532 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.255 $Y=1.35
+ $X2=3.255 $Y2=1.557
r72 8 10 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=3.255 $Y=1.35
+ $X2=3.255 $Y2=0.74
r73 5 23 22.3532 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=2.865 $Y=1.765
+ $X2=2.865 $Y2=1.557
r74 5 7 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.865 $Y=1.765
+ $X2=2.865 $Y2=2.4
r75 1 19 22.3532 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.425 $Y=1.35
+ $X2=2.425 $Y2=1.557
r76 1 3 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.425 $Y=1.35
+ $X2=2.425 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HS__O32AI_2%A2 3 5 7 8 10 13 15 16 24
c51 24 0 1.91457e-19 $X=4.215 $Y=1.557
c52 16 0 1.57212e-19 $X=4.08 $Y=1.665
r53 24 25 1.9127 $w=3.78e-07 $l=1.5e-08 $layer=POLY_cond $X=4.215 $Y=1.557
+ $X2=4.23 $Y2=1.557
r54 22 24 47.8175 $w=3.78e-07 $l=3.75e-07 $layer=POLY_cond $X=3.84 $Y=1.557
+ $X2=4.215 $Y2=1.557
r55 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.84
+ $Y=1.515 $X2=3.84 $Y2=1.515
r56 20 22 9.56349 $w=3.78e-07 $l=7.5e-08 $layer=POLY_cond $X=3.765 $Y=1.557
+ $X2=3.84 $Y2=1.557
r57 19 20 1.9127 $w=3.78e-07 $l=1.5e-08 $layer=POLY_cond $X=3.75 $Y=1.557
+ $X2=3.765 $Y2=1.557
r58 16 23 6.43224 $w=4.28e-07 $l=2.4e-07 $layer=LI1_cond $X=4.08 $Y=1.565
+ $X2=3.84 $Y2=1.565
r59 15 23 6.43224 $w=4.28e-07 $l=2.4e-07 $layer=LI1_cond $X=3.6 $Y=1.565
+ $X2=3.84 $Y2=1.565
r60 11 25 24.4846 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.23 $Y=1.35
+ $X2=4.23 $Y2=1.557
r61 11 13 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=4.23 $Y=1.35
+ $X2=4.23 $Y2=0.74
r62 8 24 24.4846 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=4.215 $Y=1.765
+ $X2=4.215 $Y2=1.557
r63 8 10 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=4.215 $Y=1.765
+ $X2=4.215 $Y2=2.4
r64 5 20 24.4846 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=3.765 $Y=1.765
+ $X2=3.765 $Y2=1.557
r65 5 7 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.765 $Y=1.765
+ $X2=3.765 $Y2=2.4
r66 1 19 24.4846 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.75 $Y=1.35
+ $X2=3.75 $Y2=1.557
r67 1 3 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=3.75 $Y=1.35 $X2=3.75
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HS__O32AI_2%A1 3 5 7 8 10 13 15 16 17 18 19 24 32
r48 32 33 1.9127 $w=3.78e-07 $l=1.5e-08 $layer=POLY_cond $X=5.73 $Y=1.557
+ $X2=5.745 $Y2=1.557
r49 30 32 35.0661 $w=3.78e-07 $l=2.75e-07 $layer=POLY_cond $X=5.455 $Y=1.557
+ $X2=5.73 $Y2=1.557
r50 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.455
+ $Y=1.515 $X2=5.455 $Y2=1.515
r51 28 30 22.9524 $w=3.78e-07 $l=1.8e-07 $layer=POLY_cond $X=5.275 $Y=1.557
+ $X2=5.455 $Y2=1.557
r52 27 31 9.11234 $w=4.28e-07 $l=3.4e-07 $layer=LI1_cond $X=5.115 $Y=1.565
+ $X2=5.455 $Y2=1.565
r53 26 27 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.115
+ $Y=1.515 $X2=5.115 $Y2=1.515
r54 24 28 12.3802 $w=3.78e-07 $l=1.08995e-07 $layer=POLY_cond $X=5.185 $Y=1.515
+ $X2=5.275 $Y2=1.557
r55 24 26 12.2403 $w=3.3e-07 $l=7e-08 $layer=POLY_cond $X=5.185 $Y=1.515
+ $X2=5.115 $Y2=1.515
r56 18 19 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=5.52 $Y=1.565 $X2=6
+ $Y2=1.565
r57 18 31 1.74206 $w=4.28e-07 $l=6.5e-08 $layer=LI1_cond $X=5.52 $Y=1.565
+ $X2=5.455 $Y2=1.565
r58 17 27 2.01008 $w=4.28e-07 $l=7.5e-08 $layer=LI1_cond $X=5.04 $Y=1.565
+ $X2=5.115 $Y2=1.565
r59 16 17 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=4.56 $Y=1.565
+ $X2=5.04 $Y2=1.565
r60 15 26 62.0758 $w=3.3e-07 $l=3.55e-07 $layer=POLY_cond $X=4.76 $Y=1.515
+ $X2=5.115 $Y2=1.515
r61 11 33 24.4846 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=5.745 $Y=1.35
+ $X2=5.745 $Y2=1.557
r62 11 13 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=5.745 $Y=1.35
+ $X2=5.745 $Y2=0.74
r63 8 32 24.4846 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=5.73 $Y=1.765
+ $X2=5.73 $Y2=1.557
r64 8 10 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=5.73 $Y=1.765
+ $X2=5.73 $Y2=2.4
r65 5 28 24.4846 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=5.275 $Y=1.765
+ $X2=5.275 $Y2=1.557
r66 5 7 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=5.275 $Y=1.765
+ $X2=5.275 $Y2=2.4
r67 1 15 32.1775 $w=3.3e-07 $l=1.98997e-07 $layer=POLY_cond $X=4.685 $Y=1.35
+ $X2=4.76 $Y2=1.515
r68 1 3 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=4.685 $Y=1.35
+ $X2=4.685 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HS__O32AI_2%A_27_368# 1 2 3 12 16 17 18 19 20 27
c36 27 0 1.68844e-19 $X=2.08 $Y=2.455
r37 21 25 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.265 $Y=2.375
+ $X2=1.18 $Y2=2.375
r38 20 27 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.915 $Y=2.375
+ $X2=2.08 $Y2=2.375
r39 20 21 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=1.915 $Y=2.375
+ $X2=1.265 $Y2=2.375
r40 18 25 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.18 $Y=2.46 $X2=1.18
+ $Y2=2.375
r41 18 19 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=1.18 $Y=2.46
+ $X2=1.18 $Y2=2.905
r42 16 19 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.095 $Y=2.99
+ $X2=1.18 $Y2=2.905
r43 16 17 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=1.095 $Y=2.99
+ $X2=0.365 $Y2=2.99
r44 12 15 32.2684 $w=2.48e-07 $l=7e-07 $layer=LI1_cond $X=0.24 $Y=2.115 $X2=0.24
+ $Y2=2.815
r45 10 17 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.24 $Y=2.905
+ $X2=0.365 $Y2=2.99
r46 10 15 4.14879 $w=2.48e-07 $l=9e-08 $layer=LI1_cond $X=0.24 $Y=2.905 $X2=0.24
+ $Y2=2.815
r47 3 27 300 $w=1.7e-07 $l=6.85912e-07 $layer=licon1_PDIFF $count=2 $X=1.93
+ $Y=1.84 $X2=2.08 $Y2=2.455
r48 2 25 300 $w=1.7e-07 $l=6.85912e-07 $layer=licon1_PDIFF $count=2 $X=1.03
+ $Y=1.84 $X2=1.18 $Y2=2.455
r49 1 15 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.815
r50 1 12 400 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.115
.ends

.subckt PM_SKY130_FD_SC_HS__O32AI_2%Y 1 2 3 4 15 19 20 21 25 27 32 33 34 35 45
+ 46
r91 45 46 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=3.09 $Y=1.985
+ $X2=3.09 $Y2=1.82
r92 34 45 1.74613 $w=3.28e-07 $l=5e-08 $layer=LI1_cond $X=3.09 $Y=2.035 $X2=3.09
+ $Y2=1.985
r93 34 35 8.20134 $w=4.98e-07 $l=2.85e-07 $layer=LI1_cond $X=3.09 $Y=2.12
+ $X2=3.09 $Y2=2.405
r94 29 46 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=3.01 $Y=1.18 $X2=3.01
+ $Y2=1.82
r95 28 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.875 $Y=1.095
+ $X2=1.71 $Y2=1.095
r96 27 29 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.925 $Y=1.095
+ $X2=3.01 $Y2=1.18
r97 27 28 68.5027 $w=1.68e-07 $l=1.05e-06 $layer=LI1_cond $X=2.925 $Y=1.095
+ $X2=1.875 $Y2=1.095
r98 23 33 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.71 $Y=1.01 $X2=1.71
+ $Y2=1.095
r99 23 25 8.20679 $w=3.28e-07 $l=2.35e-07 $layer=LI1_cond $X=1.71 $Y=1.01
+ $X2=1.71 $Y2=0.775
r100 22 32 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.895 $Y=2.035
+ $X2=0.73 $Y2=2.035
r101 21 34 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.925 $Y=2.035
+ $X2=3.09 $Y2=2.035
r102 21 22 132.439 $w=1.68e-07 $l=2.03e-06 $layer=LI1_cond $X=2.925 $Y=2.035
+ $X2=0.895 $Y2=2.035
r103 19 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.545 $Y=1.095
+ $X2=1.71 $Y2=1.095
r104 19 20 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.545 $Y=1.095
+ $X2=0.875 $Y2=1.095
r105 13 20 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.71 $Y=1.01
+ $X2=0.875 $Y2=1.095
r106 13 15 8.20679 $w=3.28e-07 $l=2.35e-07 $layer=LI1_cond $X=0.71 $Y=1.01
+ $X2=0.71 $Y2=0.775
r107 4 45 300 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=2 $X=2.94
+ $Y=1.84 $X2=3.09 $Y2=1.985
r108 3 32 300 $w=1.7e-07 $l=3.4187e-07 $layer=licon1_PDIFF $count=2 $X=0.58
+ $Y=1.84 $X2=0.73 $Y2=2.115
r109 2 25 182 $w=1.7e-07 $l=4.99074e-07 $layer=licon1_NDIFF $count=1 $X=1.5
+ $Y=0.37 $X2=1.71 $Y2=0.775
r110 1 15 182 $w=1.7e-07 $l=4.69814e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.37 $X2=0.71 $Y2=0.775
.ends

.subckt PM_SKY130_FD_SC_HS__O32AI_2%VPWR 1 2 3 12 16 18 20 24 26 34 39 45 48 52
c66 12 0 1.88367e-19 $X=1.63 $Y=2.805
r67 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r68 48 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r69 45 46 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r70 43 52 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=3.33 $X2=6
+ $Y2=3.33
r71 43 49 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=5.04 $Y2=3.33
r72 42 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r73 40 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.165 $Y=3.33 $X2=5
+ $Y2=3.33
r74 40 42 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=5.165 $Y=3.33
+ $X2=5.52 $Y2=3.33
r75 39 51 4.0045 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=5.87 $Y=3.33
+ $X2=6.055 $Y2=3.33
r76 39 42 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=5.87 $Y=3.33
+ $X2=5.52 $Y2=3.33
r77 38 49 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=5.04 $Y2=3.33
r78 37 38 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r79 35 45 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.715 $Y=3.33
+ $X2=1.59 $Y2=3.33
r80 35 37 185.61 $w=1.68e-07 $l=2.845e-06 $layer=LI1_cond $X=1.715 $Y=3.33
+ $X2=4.56 $Y2=3.33
r81 34 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.835 $Y=3.33 $X2=5
+ $Y2=3.33
r82 34 37 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=4.835 $Y=3.33
+ $X2=4.56 $Y2=3.33
r83 33 46 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=1.68 $Y2=3.33
r84 32 33 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r85 29 33 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=1.2 $Y2=3.33
r86 28 32 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.24 $Y=3.33 $X2=1.2
+ $Y2=3.33
r87 28 29 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r88 26 45 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.465 $Y=3.33
+ $X2=1.59 $Y2=3.33
r89 26 32 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=1.465 $Y=3.33
+ $X2=1.2 $Y2=3.33
r90 24 38 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=4.56 $Y2=3.33
r91 24 46 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=1.68 $Y2=3.33
r92 20 23 32.2684 $w=2.48e-07 $l=7e-07 $layer=LI1_cond $X=5.995 $Y=2.115
+ $X2=5.995 $Y2=2.815
r93 18 51 3.13866 $w=2.5e-07 $l=1.11018e-07 $layer=LI1_cond $X=5.995 $Y=3.245
+ $X2=6.055 $Y2=3.33
r94 18 23 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=5.995 $Y=3.245
+ $X2=5.995 $Y2=2.815
r95 14 48 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5 $Y=3.245 $X2=5
+ $Y2=3.33
r96 14 16 27.5888 $w=3.28e-07 $l=7.9e-07 $layer=LI1_cond $X=5 $Y=3.245 $X2=5
+ $Y2=2.455
r97 10 45 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.59 $Y=3.245
+ $X2=1.59 $Y2=3.33
r98 10 12 20.283 $w=2.48e-07 $l=4.4e-07 $layer=LI1_cond $X=1.59 $Y=3.245
+ $X2=1.59 $Y2=2.805
r99 3 23 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=5.805
+ $Y=1.84 $X2=5.955 $Y2=2.815
r100 3 20 400 $w=1.7e-07 $l=3.4187e-07 $layer=licon1_PDIFF $count=1 $X=5.805
+ $Y=1.84 $X2=5.955 $Y2=2.115
r101 2 16 300 $w=1.7e-07 $l=6.83667e-07 $layer=licon1_PDIFF $count=2 $X=4.855
+ $Y=1.84 $X2=5 $Y2=2.455
r102 1 12 600 $w=1.7e-07 $l=1.03729e-06 $layer=licon1_PDIFF $count=1 $X=1.48
+ $Y=1.84 $X2=1.63 $Y2=2.805
.ends

.subckt PM_SKY130_FD_SC_HS__O32AI_2%A_499_368# 1 2 3 12 14 15 18 22 26 28
r38 24 26 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=4.44 $Y=2.905
+ $X2=4.44 $Y2=2.455
r39 23 28 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.625 $Y=2.99
+ $X2=3.54 $Y2=2.99
r40 22 24 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.275 $Y=2.99
+ $X2=4.44 $Y2=2.905
r41 22 23 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=4.275 $Y=2.99
+ $X2=3.625 $Y2=2.99
r42 18 21 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=3.54 $Y=2.115 $X2=3.54
+ $Y2=2.815
r43 16 28 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.54 $Y=2.905
+ $X2=3.54 $Y2=2.99
r44 16 21 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=3.54 $Y=2.905 $X2=3.54
+ $Y2=2.815
r45 14 28 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.455 $Y=2.99
+ $X2=3.54 $Y2=2.99
r46 14 15 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=3.455 $Y=2.99
+ $X2=2.725 $Y2=2.99
r47 10 15 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=2.6 $Y=2.905
+ $X2=2.725 $Y2=2.99
r48 10 12 20.744 $w=2.48e-07 $l=4.5e-07 $layer=LI1_cond $X=2.6 $Y=2.905 $X2=2.6
+ $Y2=2.455
r49 3 26 300 $w=1.7e-07 $l=6.85912e-07 $layer=licon1_PDIFF $count=2 $X=4.29
+ $Y=1.84 $X2=4.44 $Y2=2.455
r50 2 21 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=3.39
+ $Y=1.84 $X2=3.54 $Y2=2.815
r51 2 18 400 $w=1.7e-07 $l=3.4187e-07 $layer=licon1_PDIFF $count=1 $X=3.39
+ $Y=1.84 $X2=3.54 $Y2=2.115
r52 1 12 300 $w=1.7e-07 $l=6.83667e-07 $layer=licon1_PDIFF $count=2 $X=2.495
+ $Y=1.84 $X2=2.64 $Y2=2.455
.ends

.subckt PM_SKY130_FD_SC_HS__O32AI_2%A_768_368# 1 2 9 11 13 16
c30 9 0 1.91457e-19 $X=5.335 $Y=2.035
r31 11 18 2.63384 $w=3.35e-07 $l=8.5e-08 $layer=LI1_cond $X=5.502 $Y=2.12
+ $X2=5.502 $Y2=2.035
r32 11 13 23.9089 $w=3.33e-07 $l=6.95e-07 $layer=LI1_cond $X=5.502 $Y=2.12
+ $X2=5.502 $Y2=2.815
r33 10 16 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.075 $Y=2.035
+ $X2=3.95 $Y2=2.035
r34 9 18 5.17472 $w=1.7e-07 $l=1.67e-07 $layer=LI1_cond $X=5.335 $Y=2.035
+ $X2=5.502 $Y2=2.035
r35 9 10 82.2032 $w=1.68e-07 $l=1.26e-06 $layer=LI1_cond $X=5.335 $Y=2.035
+ $X2=4.075 $Y2=2.035
r36 2 18 400 $w=1.7e-07 $l=2.59374e-07 $layer=licon1_PDIFF $count=1 $X=5.35
+ $Y=1.84 $X2=5.5 $Y2=2.035
r37 2 13 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=5.35
+ $Y=1.84 $X2=5.5 $Y2=2.815
r38 1 16 300 $w=1.7e-07 $l=3.4187e-07 $layer=licon1_PDIFF $count=2 $X=3.84
+ $Y=1.84 $X2=3.99 $Y2=2.115
.ends

.subckt PM_SKY130_FD_SC_HS__O32AI_2%A_27_74# 1 2 3 4 5 6 21 23 24 27 29 34 35 36
+ 38 39 40 43 45 49 51 53 56
r91 53 55 8.3814 $w=3.28e-07 $l=2.4e-07 $layer=LI1_cond $X=3.47 $Y=0.515
+ $X2=3.47 $Y2=0.755
r92 47 49 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=5.96 $Y=1.01
+ $X2=5.96 $Y2=0.515
r93 46 56 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.635 $Y=1.095
+ $X2=4.47 $Y2=1.095
r94 45 47 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=5.795 $Y=1.095
+ $X2=5.96 $Y2=1.01
r95 45 46 75.6791 $w=1.68e-07 $l=1.16e-06 $layer=LI1_cond $X=5.795 $Y=1.095
+ $X2=4.635 $Y2=1.095
r96 41 56 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.47 $Y=1.01 $X2=4.47
+ $Y2=1.095
r97 41 43 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=4.47 $Y=1.01
+ $X2=4.47 $Y2=0.515
r98 39 56 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.305 $Y=1.095
+ $X2=4.47 $Y2=1.095
r99 39 40 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.305 $Y=1.095
+ $X2=3.635 $Y2=1.095
r100 38 40 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.47 $Y=1.01
+ $X2=3.635 $Y2=1.095
r101 37 55 2.96841 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=3.47 $Y=0.84
+ $X2=3.47 $Y2=0.755
r102 37 38 5.93683 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=3.47 $Y=0.84
+ $X2=3.47 $Y2=1.01
r103 35 55 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.305 $Y=0.755
+ $X2=3.47 $Y2=0.755
r104 35 36 60.6738 $w=1.68e-07 $l=9.3e-07 $layer=LI1_cond $X=3.305 $Y=0.755
+ $X2=2.375 $Y2=0.755
r105 32 36 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.21 $Y=0.67
+ $X2=2.375 $Y2=0.755
r106 32 34 2.61919 $w=3.28e-07 $l=7.5e-08 $layer=LI1_cond $X=2.21 $Y=0.67
+ $X2=2.21 $Y2=0.595
r107 31 34 5.93683 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=2.21 $Y=0.425
+ $X2=2.21 $Y2=0.595
r108 30 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.375 $Y=0.34
+ $X2=1.21 $Y2=0.34
r109 29 31 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.045 $Y=0.34
+ $X2=2.21 $Y2=0.425
r110 29 30 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.045 $Y=0.34
+ $X2=1.375 $Y2=0.34
r111 25 51 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.21 $Y=0.425
+ $X2=1.21 $Y2=0.34
r112 25 27 8.20679 $w=3.28e-07 $l=2.35e-07 $layer=LI1_cond $X=1.21 $Y=0.425
+ $X2=1.21 $Y2=0.66
r113 23 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.045 $Y=0.34
+ $X2=1.21 $Y2=0.34
r114 23 24 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.045 $Y=0.34
+ $X2=0.365 $Y2=0.34
r115 19 24 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.24 $Y=0.425
+ $X2=0.365 $Y2=0.34
r116 19 21 4.14879 $w=2.48e-07 $l=9e-08 $layer=LI1_cond $X=0.24 $Y=0.425
+ $X2=0.24 $Y2=0.515
r117 6 49 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=5.82
+ $Y=0.37 $X2=5.96 $Y2=0.515
r118 5 43 91 $w=1.7e-07 $l=2.26164e-07 $layer=licon1_NDIFF $count=2 $X=4.305
+ $Y=0.37 $X2=4.47 $Y2=0.515
r119 4 53 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.33
+ $Y=0.37 $X2=3.47 $Y2=0.515
r120 3 34 182 $w=1.7e-07 $l=3.1285e-07 $layer=licon1_NDIFF $count=1 $X=2 $Y=0.37
+ $X2=2.21 $Y2=0.595
r121 2 27 182 $w=1.7e-07 $l=3.80789e-07 $layer=licon1_NDIFF $count=1 $X=1
+ $Y=0.37 $X2=1.21 $Y2=0.66
r122 1 21 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__O32AI_2%VGND 1 2 3 12 15 16 17 37 38 43 46 50 56
r66 55 56 11.2541 $w=8.88e-07 $l=9.5e-08 $layer=LI1_cond $X=5.53 $Y=0.36
+ $X2=5.625 $Y2=0.36
r67 52 55 0.137079 $w=8.88e-07 $l=1e-08 $layer=LI1_cond $X=5.52 $Y=0.36 $X2=5.53
+ $Y2=0.36
r68 52 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r69 49 53 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=5.52
+ $Y2=0
r70 48 52 6.57978 $w=8.88e-07 $l=4.8e-07 $layer=LI1_cond $X=5.04 $Y=0.36
+ $X2=5.52 $Y2=0.36
r71 48 50 13.1732 $w=8.88e-07 $l=2.35e-07 $layer=LI1_cond $X=5.04 $Y=0.36
+ $X2=4.805 $Y2=0.36
r72 48 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r73 45 46 12.5119 $w=5.83e-07 $l=2.85e-07 $layer=LI1_cond $X=2.84 $Y=0.207
+ $X2=3.125 $Y2=0.207
r74 41 45 4.08916 $w=5.83e-07 $l=2e-07 $layer=LI1_cond $X=2.64 $Y=0.207 $X2=2.84
+ $Y2=0.207
r75 41 43 8.42273 $w=5.83e-07 $l=8.5e-08 $layer=LI1_cond $X=2.64 $Y=0.207
+ $X2=2.555 $Y2=0.207
r76 41 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r77 38 53 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=0 $X2=5.52
+ $Y2=0
r78 37 56 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=6 $Y=0 $X2=5.625
+ $Y2=0
r79 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=0 $X2=6 $Y2=0
r80 34 49 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=5.04
+ $Y2=0
r81 33 50 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=4.56 $Y=0 $X2=4.805
+ $Y2=0
r82 33 34 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r83 30 34 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.56
+ $Y2=0
r84 29 46 30.9893 $w=1.68e-07 $l=4.75e-07 $layer=LI1_cond $X=3.6 $Y=0 $X2=3.125
+ $Y2=0
r85 29 30 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r86 26 42 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r87 25 43 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=2.16 $Y=0 $X2=2.555
+ $Y2=0
r88 25 26 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r89 22 26 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=0.24 $Y=0 $X2=2.16
+ $Y2=0
r90 21 25 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=0.24 $Y=0 $X2=2.16
+ $Y2=0
r91 21 22 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r92 17 30 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=3.6
+ $Y2=0
r93 17 42 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=2.64
+ $Y2=0
r94 15 29 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=3.805 $Y=0 $X2=3.6
+ $Y2=0
r95 15 16 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.805 $Y=0 $X2=3.97
+ $Y2=0
r96 14 33 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=4.135 $Y=0 $X2=4.56
+ $Y2=0
r97 14 16 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.135 $Y=0 $X2=3.97
+ $Y2=0
r98 10 16 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.97 $Y=0.085
+ $X2=3.97 $Y2=0
r99 10 12 19.2074 $w=3.28e-07 $l=5.5e-07 $layer=LI1_cond $X=3.97 $Y=0.085
+ $X2=3.97 $Y2=0.635
r100 3 55 91 $w=1.7e-07 $l=8.94874e-07 $layer=licon1_NDIFF $count=2 $X=4.76
+ $Y=0.37 $X2=5.53 $Y2=0.64
r101 2 12 182 $w=1.7e-07 $l=3.29621e-07 $layer=licon1_NDIFF $count=1 $X=3.825
+ $Y=0.37 $X2=3.97 $Y2=0.635
r102 1 45 182 $w=1.7e-07 $l=3.57071e-07 $layer=licon1_NDIFF $count=1 $X=2.5
+ $Y=0.37 $X2=2.84 $Y2=0.335
.ends

