* File: sky130_fd_sc_hs__dlclkp_4.pxi.spice
* Created: Tue Sep  1 20:01:33 2020
* 
x_PM_SKY130_FD_SC_HS__DLCLKP_4%A_84_48# N_A_84_48#_M1018_d N_A_84_48#_M1009_d
+ N_A_84_48#_c_147_n N_A_84_48#_M1021_g N_A_84_48#_c_148_n N_A_84_48#_M1011_g
+ N_A_84_48#_c_149_n N_A_84_48#_c_150_n N_A_84_48#_c_159_p N_A_84_48#_c_213_p
+ N_A_84_48#_c_151_n N_A_84_48#_c_183_p N_A_84_48#_c_201_p N_A_84_48#_c_170_p
+ N_A_84_48#_c_218_p N_A_84_48#_c_155_n N_A_84_48#_c_152_n
+ PM_SKY130_FD_SC_HS__DLCLKP_4%A_84_48#
x_PM_SKY130_FD_SC_HS__DLCLKP_4%GATE N_GATE_c_233_n N_GATE_M1002_g N_GATE_M1017_g
+ GATE PM_SKY130_FD_SC_HS__DLCLKP_4%GATE
x_PM_SKY130_FD_SC_HS__DLCLKP_4%A_334_54# N_A_334_54#_M1019_s N_A_334_54#_M1016_s
+ N_A_334_54#_c_265_n N_A_334_54#_M1018_g N_A_334_54#_c_274_n
+ N_A_334_54#_M1003_g N_A_334_54#_c_266_n N_A_334_54#_M1004_g
+ N_A_334_54#_M1025_g N_A_334_54#_c_268_n N_A_334_54#_c_269_n
+ N_A_334_54#_c_277_n N_A_334_54#_c_293_n N_A_334_54#_c_270_n
+ N_A_334_54#_c_338_p N_A_334_54#_c_279_n N_A_334_54#_c_342_p
+ N_A_334_54#_c_271_n N_A_334_54#_c_272_n N_A_334_54#_c_280_n
+ N_A_334_54#_c_273_n PM_SKY130_FD_SC_HS__DLCLKP_4%A_334_54#
x_PM_SKY130_FD_SC_HS__DLCLKP_4%A_334_338# N_A_334_338#_M1025_d
+ N_A_334_338#_M1004_d N_A_334_338#_c_394_n N_A_334_338#_M1009_g
+ N_A_334_338#_c_387_n N_A_334_338#_c_396_n N_A_334_338#_M1012_g
+ N_A_334_338#_c_389_n N_A_334_338#_c_390_n N_A_334_338#_c_391_n
+ N_A_334_338#_c_399_n N_A_334_338#_c_392_n N_A_334_338#_c_393_n
+ PM_SKY130_FD_SC_HS__DLCLKP_4%A_334_338#
x_PM_SKY130_FD_SC_HS__DLCLKP_4%A_27_74# N_A_27_74#_M1021_s N_A_27_74#_M1011_s
+ N_A_27_74#_c_465_n N_A_27_74#_c_466_n N_A_27_74#_c_480_n N_A_27_74#_M1010_g
+ N_A_27_74#_M1000_g N_A_27_74#_M1023_g N_A_27_74#_c_469_n N_A_27_74#_M1007_g
+ N_A_27_74#_c_470_n N_A_27_74#_c_482_n N_A_27_74#_c_489_n N_A_27_74#_c_493_n
+ N_A_27_74#_c_471_n N_A_27_74#_c_472_n N_A_27_74#_c_473_n N_A_27_74#_c_474_n
+ N_A_27_74#_c_475_n N_A_27_74#_c_534_n N_A_27_74#_c_476_n N_A_27_74#_c_483_n
+ N_A_27_74#_c_477_n N_A_27_74#_c_478_n PM_SKY130_FD_SC_HS__DLCLKP_4%A_27_74#
x_PM_SKY130_FD_SC_HS__DLCLKP_4%CLK N_CLK_c_608_n N_CLK_c_609_n N_CLK_M1016_g
+ N_CLK_M1019_g N_CLK_c_610_n N_CLK_M1014_g N_CLK_M1005_g CLK N_CLK_c_606_n
+ N_CLK_c_607_n PM_SKY130_FD_SC_HS__DLCLKP_4%CLK
x_PM_SKY130_FD_SC_HS__DLCLKP_4%A_1044_368# N_A_1044_368#_M1023_d
+ N_A_1044_368#_M1014_d N_A_1044_368#_c_651_n N_A_1044_368#_c_664_n
+ N_A_1044_368#_M1001_g N_A_1044_368#_M1006_g N_A_1044_368#_c_665_n
+ N_A_1044_368#_M1020_g N_A_1044_368#_M1008_g N_A_1044_368#_c_654_n
+ N_A_1044_368#_c_655_n N_A_1044_368#_c_668_n N_A_1044_368#_M1022_g
+ N_A_1044_368#_M1013_g N_A_1044_368#_c_669_n N_A_1044_368#_M1024_g
+ N_A_1044_368#_M1015_g N_A_1044_368#_c_658_n N_A_1044_368#_c_671_n
+ N_A_1044_368#_c_672_n N_A_1044_368#_c_673_n N_A_1044_368#_c_659_n
+ N_A_1044_368#_c_660_n N_A_1044_368#_c_661_n N_A_1044_368#_c_662_n
+ PM_SKY130_FD_SC_HS__DLCLKP_4%A_1044_368#
x_PM_SKY130_FD_SC_HS__DLCLKP_4%VPWR N_VPWR_M1011_d N_VPWR_M1010_d N_VPWR_M1016_d
+ N_VPWR_M1007_d N_VPWR_M1020_d N_VPWR_M1024_d N_VPWR_c_772_n N_VPWR_c_773_n
+ N_VPWR_c_774_n N_VPWR_c_775_n N_VPWR_c_776_n N_VPWR_c_777_n N_VPWR_c_778_n
+ N_VPWR_c_779_n N_VPWR_c_780_n N_VPWR_c_781_n N_VPWR_c_782_n VPWR
+ N_VPWR_c_783_n N_VPWR_c_784_n N_VPWR_c_785_n N_VPWR_c_786_n N_VPWR_c_787_n
+ N_VPWR_c_788_n N_VPWR_c_789_n N_VPWR_c_771_n PM_SKY130_FD_SC_HS__DLCLKP_4%VPWR
x_PM_SKY130_FD_SC_HS__DLCLKP_4%GCLK N_GCLK_M1006_d N_GCLK_M1013_d N_GCLK_M1001_s
+ N_GCLK_M1022_s N_GCLK_c_884_n N_GCLK_c_877_n N_GCLK_c_885_n N_GCLK_c_903_n
+ N_GCLK_c_878_n N_GCLK_c_879_n N_GCLK_c_886_n N_GCLK_c_880_n N_GCLK_c_881_n
+ N_GCLK_c_882_n GCLK GCLK PM_SKY130_FD_SC_HS__DLCLKP_4%GCLK
x_PM_SKY130_FD_SC_HS__DLCLKP_4%VGND N_VGND_M1021_d N_VGND_M1000_d N_VGND_M1019_d
+ N_VGND_M1006_s N_VGND_M1008_s N_VGND_M1015_s N_VGND_c_948_n N_VGND_c_949_n
+ N_VGND_c_950_n N_VGND_c_951_n N_VGND_c_952_n N_VGND_c_953_n VGND
+ N_VGND_c_954_n N_VGND_c_955_n N_VGND_c_956_n N_VGND_c_957_n N_VGND_c_958_n
+ N_VGND_c_959_n N_VGND_c_960_n N_VGND_c_961_n N_VGND_c_962_n N_VGND_c_963_n
+ N_VGND_c_964_n PM_SKY130_FD_SC_HS__DLCLKP_4%VGND
cc_1 VNB N_A_84_48#_c_147_n 0.0230635f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.22
cc_2 VNB N_A_84_48#_c_148_n 0.0514445f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=1.765
cc_3 VNB N_A_84_48#_c_149_n 0.00150907f $X=-0.19 $Y=-0.245 $X2=0.795 $Y2=1.97
cc_4 VNB N_A_84_48#_c_150_n 0.01229f $X=-0.19 $Y=-0.245 $X2=1.435 $Y2=1.275
cc_5 VNB N_A_84_48#_c_151_n 0.00256251f $X=-0.19 $Y=-0.245 $X2=1.52 $Y2=1.19
cc_6 VNB N_A_84_48#_c_152_n 0.00621205f $X=-0.19 $Y=-0.245 $X2=0.707 $Y2=1.275
cc_7 VNB N_GATE_c_233_n 0.0194459f $X=-0.19 $Y=-0.245 $X2=1.82 $Y2=0.4
cc_8 VNB N_GATE_M1017_g 0.0348671f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB GATE 0.00265138f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_10 VNB N_A_334_54#_c_265_n 0.0179936f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.22
cc_11 VNB N_A_334_54#_c_266_n 0.0330076f $X=-0.19 $Y=-0.245 $X2=0.795 $Y2=1.55
cc_12 VNB N_A_334_54#_M1025_g 0.0241088f $X=-0.19 $Y=-0.245 $X2=1.52 $Y2=0.98
cc_13 VNB N_A_334_54#_c_268_n 0.00525847f $X=-0.19 $Y=-0.245 $X2=1.52 $Y2=2.52
cc_14 VNB N_A_334_54#_c_269_n 0.0373992f $X=-0.19 $Y=-0.245 $X2=1.605 $Y2=0.815
cc_15 VNB N_A_334_54#_c_270_n 0.00268632f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_334_54#_c_271_n 0.00716059f $X=-0.19 $Y=-0.245 $X2=0.695 $Y2=1.385
cc_17 VNB N_A_334_54#_c_272_n 0.0618249f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.385
cc_18 VNB N_A_334_54#_c_273_n 0.00537146f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_334_338#_c_387_n 0.00433237f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=1.765
cc_20 VNB N_A_334_338#_M1012_g 0.0377623f $X=-0.19 $Y=-0.245 $X2=0.795 $Y2=1.97
cc_21 VNB N_A_334_338#_c_389_n 0.00766943f $X=-0.19 $Y=-0.245 $X2=1.52 $Y2=0.98
cc_22 VNB N_A_334_338#_c_390_n 0.00409063f $X=-0.19 $Y=-0.245 $X2=1.52 $Y2=1.19
cc_23 VNB N_A_334_338#_c_391_n 0.0223667f $X=-0.19 $Y=-0.245 $X2=2.06 $Y2=0.815
cc_24 VNB N_A_334_338#_c_392_n 0.0113424f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_334_338#_c_393_n 0.00929218f $X=-0.19 $Y=-0.245 $X2=0.695
+ $Y2=1.385
cc_26 VNB N_A_27_74#_c_465_n 0.00576023f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.22
cc_27 VNB N_A_27_74#_c_466_n 0.0106067f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_28 VNB N_A_27_74#_M1000_g 0.0266169f $X=-0.19 $Y=-0.245 $X2=1.435 $Y2=1.275
cc_29 VNB N_A_27_74#_M1023_g 0.023672f $X=-0.19 $Y=-0.245 $X2=0.88 $Y2=2.055
cc_30 VNB N_A_27_74#_c_469_n 0.0300223f $X=-0.19 $Y=-0.245 $X2=1.52 $Y2=1.19
cc_31 VNB N_A_27_74#_c_470_n 0.0207357f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_27_74#_c_471_n 0.0309217f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_27_74#_c_472_n 0.00233902f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_27_74#_c_473_n 0.00122215f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_27_74#_c_474_n 0.00767704f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_27_74#_c_475_n 0.0354209f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_27_74#_c_476_n 0.00704942f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_27_74#_c_477_n 0.031259f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_27_74#_c_478_n 0.0460418f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_CLK_M1019_g 0.0293985f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_41 VNB N_CLK_M1005_g 0.0222599f $X=-0.19 $Y=-0.245 $X2=1.435 $Y2=1.275
cc_42 VNB N_CLK_c_606_n 0.00487367f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_CLK_c_607_n 0.0518691f $X=-0.19 $Y=-0.245 $X2=1.605 $Y2=2.685
cc_44 VNB N_A_1044_368#_c_651_n 0.0171186f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.22
cc_45 VNB N_A_1044_368#_M1006_g 0.0265413f $X=-0.19 $Y=-0.245 $X2=0.795 $Y2=1.97
cc_46 VNB N_A_1044_368#_M1008_g 0.025436f $X=-0.19 $Y=-0.245 $X2=1.52 $Y2=2.14
cc_47 VNB N_A_1044_368#_c_654_n 0.0121954f $X=-0.19 $Y=-0.245 $X2=1.605
+ $Y2=0.815
cc_48 VNB N_A_1044_368#_c_655_n 0.0200533f $X=-0.19 $Y=-0.245 $X2=2.06 $Y2=0.815
cc_49 VNB N_A_1044_368#_M1013_g 0.0254487f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_A_1044_368#_M1015_g 0.036104f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.385
cc_51 VNB N_A_1044_368#_c_658_n 0.0317783f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_A_1044_368#_c_659_n 0.0281117f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_A_1044_368#_c_660_n 0.00409086f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_A_1044_368#_c_661_n 0.0599216f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_A_1044_368#_c_662_n 0.01192f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_VPWR_c_771_n 0.362705f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_GCLK_c_877_n 0.00240191f $X=-0.19 $Y=-0.245 $X2=1.52 $Y2=2.14
cc_58 VNB N_GCLK_c_878_n 0.00766134f $X=-0.19 $Y=-0.245 $X2=2.06 $Y2=0.815
cc_59 VNB N_GCLK_c_879_n 0.00158543f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_GCLK_c_880_n 0.00316097f $X=-0.19 $Y=-0.245 $X2=0.695 $Y2=1.385
cc_61 VNB N_GCLK_c_881_n 3.53034e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_GCLK_c_882_n 0.00194448f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB GCLK 0.00915128f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_VGND_c_948_n 0.00727256f $X=-0.19 $Y=-0.245 $X2=1.52 $Y2=2.14
cc_65 VNB N_VGND_c_949_n 0.00972604f $X=-0.19 $Y=-0.245 $X2=2.06 $Y2=0.815
cc_66 VNB N_VGND_c_950_n 0.00396467f $X=-0.19 $Y=-0.245 $X2=2.15 $Y2=2.685
cc_67 VNB N_VGND_c_951_n 0.00807502f $X=-0.19 $Y=-0.245 $X2=0.707 $Y2=1.385
cc_68 VNB N_VGND_c_952_n 0.0120272f $X=-0.19 $Y=-0.245 $X2=0.695 $Y2=1.385
cc_69 VNB N_VGND_c_953_n 0.0353267f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.385
cc_70 VNB N_VGND_c_954_n 0.01755f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_VGND_c_955_n 0.0565077f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_VGND_c_956_n 0.0277574f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_VGND_c_957_n 0.0549955f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_VGND_c_958_n 0.0190448f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_VGND_c_959_n 0.0172524f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_VGND_c_960_n 0.0070281f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_VGND_c_961_n 0.00573719f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_VGND_c_962_n 0.00604233f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VNB N_VGND_c_963_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_VGND_c_964_n 0.467177f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_81 VPB N_A_84_48#_c_148_n 0.0291156f $X=-0.19 $Y=1.66 $X2=0.6 $Y2=1.765
cc_82 VPB N_A_84_48#_c_149_n 0.00329408f $X=-0.19 $Y=1.66 $X2=0.795 $Y2=1.97
cc_83 VPB N_A_84_48#_c_155_n 0.00267723f $X=-0.19 $Y=1.66 $X2=2.15 $Y2=2.685
cc_84 VPB N_GATE_c_233_n 0.0371834f $X=-0.19 $Y=1.66 $X2=1.82 $Y2=0.4
cc_85 VPB GATE 0.00239649f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.74
cc_86 VPB N_A_334_54#_c_274_n 0.0559551f $X=-0.19 $Y=1.66 $X2=0.6 $Y2=1.765
cc_87 VPB N_A_334_54#_c_266_n 0.0372031f $X=-0.19 $Y=1.66 $X2=0.795 $Y2=1.55
cc_88 VPB N_A_334_54#_c_268_n 0.00486805f $X=-0.19 $Y=1.66 $X2=1.52 $Y2=2.52
cc_89 VPB N_A_334_54#_c_277_n 0.0246311f $X=-0.19 $Y=1.66 $X2=2.06 $Y2=0.815
cc_90 VPB N_A_334_54#_c_270_n 0.00271009f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_91 VPB N_A_334_54#_c_279_n 0.0195272f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_92 VPB N_A_334_54#_c_280_n 0.0138077f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_93 VPB N_A_334_338#_c_394_n 0.0181106f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.22
cc_94 VPB N_A_334_338#_c_387_n 0.0278659f $X=-0.19 $Y=1.66 $X2=0.6 $Y2=1.765
cc_95 VPB N_A_334_338#_c_396_n 0.0120128f $X=-0.19 $Y=1.66 $X2=0.6 $Y2=2.4
cc_96 VPB N_A_334_338#_c_389_n 0.00547328f $X=-0.19 $Y=1.66 $X2=1.52 $Y2=0.98
cc_97 VPB N_A_334_338#_c_391_n 0.0127529f $X=-0.19 $Y=1.66 $X2=2.06 $Y2=0.815
cc_98 VPB N_A_334_338#_c_399_n 0.00203646f $X=-0.19 $Y=1.66 $X2=2.15 $Y2=2.685
cc_99 VPB N_A_27_74#_c_466_n 0.0423815f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.74
cc_100 VPB N_A_27_74#_c_480_n 0.0240069f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.74
cc_101 VPB N_A_27_74#_c_469_n 0.0242725f $X=-0.19 $Y=1.66 $X2=1.52 $Y2=1.19
cc_102 VPB N_A_27_74#_c_482_n 0.0439898f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_103 VPB N_A_27_74#_c_483_n 0.0126367f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_104 VPB N_A_27_74#_c_477_n 0.00828958f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_105 VPB N_CLK_c_608_n 0.0177893f $X=-0.19 $Y=1.66 $X2=1.835 $Y2=1.96
cc_106 VPB N_CLK_c_609_n 0.0268357f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_107 VPB N_CLK_c_610_n 0.0169757f $X=-0.19 $Y=1.66 $X2=0.6 $Y2=1.765
cc_108 VPB N_CLK_c_606_n 0.00636285f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_109 VPB N_CLK_c_607_n 0.0194408f $X=-0.19 $Y=1.66 $X2=1.605 $Y2=2.685
cc_110 VPB N_A_1044_368#_c_651_n 0.00997041f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.22
cc_111 VPB N_A_1044_368#_c_664_n 0.0163821f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.74
cc_112 VPB N_A_1044_368#_c_665_n 0.016027f $X=-0.19 $Y=1.66 $X2=0.88 $Y2=1.275
cc_113 VPB N_A_1044_368#_c_654_n 0.0093007f $X=-0.19 $Y=1.66 $X2=1.605 $Y2=0.815
cc_114 VPB N_A_1044_368#_c_655_n 0.0209962f $X=-0.19 $Y=1.66 $X2=2.06 $Y2=0.815
cc_115 VPB N_A_1044_368#_c_668_n 0.0155432f $X=-0.19 $Y=1.66 $X2=2.06 $Y2=0.815
cc_116 VPB N_A_1044_368#_c_669_n 0.0187811f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_117 VPB N_A_1044_368#_c_658_n 0.0209591f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_118 VPB N_A_1044_368#_c_671_n 0.00323293f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_119 VPB N_A_1044_368#_c_672_n 0.00290214f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_120 VPB N_A_1044_368#_c_673_n 0.00661549f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_121 VPB N_A_1044_368#_c_660_n 0.00308751f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_122 VPB N_A_1044_368#_c_662_n 0.0103718f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_123 VPB N_VPWR_c_772_n 0.0104956f $X=-0.19 $Y=1.66 $X2=1.52 $Y2=2.14
cc_124 VPB N_VPWR_c_773_n 0.00776002f $X=-0.19 $Y=1.66 $X2=2.06 $Y2=0.815
cc_125 VPB N_VPWR_c_774_n 0.0096853f $X=-0.19 $Y=1.66 $X2=2.15 $Y2=2.685
cc_126 VPB N_VPWR_c_775_n 0.0141371f $X=-0.19 $Y=1.66 $X2=0.707 $Y2=1.385
cc_127 VPB N_VPWR_c_776_n 0.00755968f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.385
cc_128 VPB N_VPWR_c_777_n 0.0120106f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_129 VPB N_VPWR_c_778_n 0.0483332f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_130 VPB N_VPWR_c_779_n 0.0238191f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_131 VPB N_VPWR_c_780_n 0.00718714f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_132 VPB N_VPWR_c_781_n 0.0354159f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_133 VPB N_VPWR_c_782_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_134 VPB N_VPWR_c_783_n 0.0556468f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_135 VPB N_VPWR_c_784_n 0.0186948f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_136 VPB N_VPWR_c_785_n 0.018682f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_137 VPB N_VPWR_c_786_n 0.0185253f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_138 VPB N_VPWR_c_787_n 0.00631473f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_139 VPB N_VPWR_c_788_n 0.0169969f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_140 VPB N_VPWR_c_789_n 0.0047828f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_141 VPB N_VPWR_c_771_n 0.110407f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_142 VPB N_GCLK_c_884_n 0.00351007f $X=-0.19 $Y=1.66 $X2=1.435 $Y2=1.275
cc_143 VPB N_GCLK_c_885_n 0.00423197f $X=-0.19 $Y=1.66 $X2=1.605 $Y2=0.815
cc_144 VPB N_GCLK_c_886_n 0.00273338f $X=-0.19 $Y=1.66 $X2=2.15 $Y2=2.685
cc_145 VPB GCLK 8.14549e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_146 VPB GCLK 0.0097106f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_147 N_A_84_48#_c_148_n N_GATE_c_233_n 0.0273784f $X=0.6 $Y=1.765 $X2=-0.19
+ $Y2=-0.245
cc_148 N_A_84_48#_c_149_n N_GATE_c_233_n 0.00309285f $X=0.795 $Y=1.97 $X2=-0.19
+ $Y2=-0.245
cc_149 N_A_84_48#_c_150_n N_GATE_c_233_n 0.00441226f $X=1.435 $Y=1.275 $X2=-0.19
+ $Y2=-0.245
cc_150 N_A_84_48#_c_159_p N_GATE_c_233_n 0.0188213f $X=1.435 $Y=2.055 $X2=-0.19
+ $Y2=-0.245
cc_151 N_A_84_48#_c_152_n N_GATE_c_233_n 0.00229665f $X=0.707 $Y=1.275 $X2=-0.19
+ $Y2=-0.245
cc_152 N_A_84_48#_c_147_n N_GATE_M1017_g 0.00900631f $X=0.495 $Y=1.22 $X2=0
+ $Y2=0
cc_153 N_A_84_48#_c_148_n N_GATE_M1017_g 0.00628804f $X=0.6 $Y=1.765 $X2=0 $Y2=0
cc_154 N_A_84_48#_c_150_n N_GATE_M1017_g 0.0148109f $X=1.435 $Y=1.275 $X2=0
+ $Y2=0
cc_155 N_A_84_48#_c_151_n N_GATE_M1017_g 0.00393105f $X=1.52 $Y=1.19 $X2=0 $Y2=0
cc_156 N_A_84_48#_c_152_n N_GATE_M1017_g 0.00224326f $X=0.707 $Y=1.275 $X2=0
+ $Y2=0
cc_157 N_A_84_48#_c_150_n GATE 0.0250347f $X=1.435 $Y=1.275 $X2=0 $Y2=0
cc_158 N_A_84_48#_c_159_p GATE 0.0221636f $X=1.435 $Y=2.055 $X2=0 $Y2=0
cc_159 N_A_84_48#_c_152_n GATE 0.0188052f $X=0.707 $Y=1.275 $X2=0 $Y2=0
cc_160 N_A_84_48#_c_151_n N_A_334_54#_c_265_n 0.00417838f $X=1.52 $Y=1.19 $X2=0
+ $Y2=0
cc_161 N_A_84_48#_c_170_p N_A_334_54#_c_265_n 0.0208157f $X=2.06 $Y=0.815 $X2=0
+ $Y2=0
cc_162 N_A_84_48#_c_155_n N_A_334_54#_c_274_n 0.0171226f $X=2.15 $Y=2.685 $X2=0
+ $Y2=0
cc_163 N_A_84_48#_M1009_d N_A_334_54#_c_268_n 0.00367686f $X=1.835 $Y=1.96 $X2=0
+ $Y2=0
cc_164 N_A_84_48#_c_150_n N_A_334_54#_c_268_n 0.0142091f $X=1.435 $Y=1.275 $X2=0
+ $Y2=0
cc_165 N_A_84_48#_c_159_p N_A_334_54#_c_268_n 0.00651027f $X=1.435 $Y=2.055
+ $X2=0 $Y2=0
cc_166 N_A_84_48#_c_151_n N_A_334_54#_c_268_n 0.00293885f $X=1.52 $Y=1.19 $X2=0
+ $Y2=0
cc_167 N_A_84_48#_c_170_p N_A_334_54#_c_268_n 0.021323f $X=2.06 $Y=0.815 $X2=0
+ $Y2=0
cc_168 N_A_84_48#_c_150_n N_A_334_54#_c_269_n 0.00140598f $X=1.435 $Y=1.275
+ $X2=0 $Y2=0
cc_169 N_A_84_48#_c_170_p N_A_334_54#_c_269_n 0.00166298f $X=2.06 $Y=0.815 $X2=0
+ $Y2=0
cc_170 N_A_84_48#_M1009_d N_A_334_54#_c_277_n 0.00136409f $X=1.835 $Y=1.96 $X2=0
+ $Y2=0
cc_171 N_A_84_48#_c_155_n N_A_334_54#_c_277_n 0.0337813f $X=2.15 $Y=2.685 $X2=0
+ $Y2=0
cc_172 N_A_84_48#_M1009_d N_A_334_54#_c_293_n 0.00272588f $X=1.835 $Y=1.96 $X2=0
+ $Y2=0
cc_173 N_A_84_48#_c_159_p N_A_334_54#_c_293_n 0.00786628f $X=1.435 $Y=2.055
+ $X2=0 $Y2=0
cc_174 N_A_84_48#_c_183_p N_A_334_54#_c_293_n 0.0164691f $X=1.52 $Y=2.52 $X2=0
+ $Y2=0
cc_175 N_A_84_48#_c_155_n N_A_334_54#_c_293_n 0.0194358f $X=2.15 $Y=2.685 $X2=0
+ $Y2=0
cc_176 N_A_84_48#_c_159_p N_A_334_338#_c_394_n 0.00128014f $X=1.435 $Y=2.055
+ $X2=0 $Y2=0
cc_177 N_A_84_48#_c_183_p N_A_334_338#_c_394_n 0.00525093f $X=1.52 $Y=2.52 $X2=0
+ $Y2=0
cc_178 N_A_84_48#_c_155_n N_A_334_338#_c_394_n 0.0216785f $X=2.15 $Y=2.685 $X2=0
+ $Y2=0
cc_179 N_A_84_48#_c_155_n N_A_334_338#_c_387_n 8.04691e-19 $X=2.15 $Y=2.685
+ $X2=0 $Y2=0
cc_180 N_A_84_48#_c_170_p N_A_334_338#_M1012_g 0.0121963f $X=2.06 $Y=0.815 $X2=0
+ $Y2=0
cc_181 N_A_84_48#_c_170_p N_A_334_338#_c_390_n 9.67748e-19 $X=2.06 $Y=0.815
+ $X2=0 $Y2=0
cc_182 N_A_84_48#_c_155_n N_A_27_74#_c_480_n 0.00156179f $X=2.15 $Y=2.685 $X2=0
+ $Y2=0
cc_183 N_A_84_48#_c_170_p N_A_27_74#_M1000_g 3.05797e-19 $X=2.06 $Y=0.815 $X2=0
+ $Y2=0
cc_184 N_A_84_48#_c_147_n N_A_27_74#_c_470_n 0.00159473f $X=0.495 $Y=1.22 $X2=0
+ $Y2=0
cc_185 N_A_84_48#_c_148_n N_A_27_74#_c_482_n 0.0181236f $X=0.6 $Y=1.765 $X2=0
+ $Y2=0
cc_186 N_A_84_48#_c_147_n N_A_27_74#_c_489_n 0.0144795f $X=0.495 $Y=1.22 $X2=0
+ $Y2=0
cc_187 N_A_84_48#_c_148_n N_A_27_74#_c_489_n 0.00175055f $X=0.6 $Y=1.765 $X2=0
+ $Y2=0
cc_188 N_A_84_48#_c_150_n N_A_27_74#_c_489_n 0.0280388f $X=1.435 $Y=1.275 $X2=0
+ $Y2=0
cc_189 N_A_84_48#_c_152_n N_A_27_74#_c_489_n 0.0254697f $X=0.707 $Y=1.275 $X2=0
+ $Y2=0
cc_190 N_A_84_48#_c_147_n N_A_27_74#_c_493_n 0.00257528f $X=0.495 $Y=1.22 $X2=0
+ $Y2=0
cc_191 N_A_84_48#_M1018_d N_A_27_74#_c_471_n 0.00241797f $X=1.82 $Y=0.4 $X2=0
+ $Y2=0
cc_192 N_A_84_48#_c_201_p N_A_27_74#_c_471_n 0.00707909f $X=1.605 $Y=0.815 $X2=0
+ $Y2=0
cc_193 N_A_84_48#_c_170_p N_A_27_74#_c_471_n 0.0325781f $X=2.06 $Y=0.815 $X2=0
+ $Y2=0
cc_194 N_A_84_48#_c_147_n N_A_27_74#_c_472_n 3.78932e-19 $X=0.495 $Y=1.22 $X2=0
+ $Y2=0
cc_195 N_A_84_48#_c_170_p N_A_27_74#_c_474_n 0.012421f $X=2.06 $Y=0.815 $X2=0
+ $Y2=0
cc_196 N_A_84_48#_c_148_n N_A_27_74#_c_483_n 0.0079847f $X=0.6 $Y=1.765 $X2=0
+ $Y2=0
cc_197 N_A_84_48#_c_149_n N_A_27_74#_c_483_n 0.00656532f $X=0.795 $Y=1.97 $X2=0
+ $Y2=0
cc_198 N_A_84_48#_c_147_n N_A_27_74#_c_477_n 0.0129583f $X=0.495 $Y=1.22 $X2=0
+ $Y2=0
cc_199 N_A_84_48#_c_148_n N_A_27_74#_c_477_n 0.00608413f $X=0.6 $Y=1.765 $X2=0
+ $Y2=0
cc_200 N_A_84_48#_c_149_n N_A_27_74#_c_477_n 0.012745f $X=0.795 $Y=1.97 $X2=0
+ $Y2=0
cc_201 N_A_84_48#_c_152_n N_A_27_74#_c_477_n 0.027924f $X=0.707 $Y=1.275 $X2=0
+ $Y2=0
cc_202 N_A_84_48#_c_149_n N_VPWR_M1011_d 0.00283262f $X=0.795 $Y=1.97 $X2=-0.19
+ $Y2=-0.245
cc_203 N_A_84_48#_c_159_p N_VPWR_M1011_d 0.0115688f $X=1.435 $Y=2.055 $X2=-0.19
+ $Y2=-0.245
cc_204 N_A_84_48#_c_213_p N_VPWR_M1011_d 0.00485774f $X=0.88 $Y=2.055 $X2=-0.19
+ $Y2=-0.245
cc_205 N_A_84_48#_c_148_n N_VPWR_c_772_n 0.0106564f $X=0.6 $Y=1.765 $X2=0 $Y2=0
cc_206 N_A_84_48#_c_159_p N_VPWR_c_772_n 0.0226626f $X=1.435 $Y=2.055 $X2=0
+ $Y2=0
cc_207 N_A_84_48#_c_213_p N_VPWR_c_772_n 0.00843013f $X=0.88 $Y=2.055 $X2=0
+ $Y2=0
cc_208 N_A_84_48#_c_148_n N_VPWR_c_779_n 0.00445602f $X=0.6 $Y=1.765 $X2=0 $Y2=0
cc_209 N_A_84_48#_c_218_p N_VPWR_c_783_n 0.00429642f $X=1.605 $Y=2.685 $X2=0
+ $Y2=0
cc_210 N_A_84_48#_c_155_n N_VPWR_c_783_n 0.0212578f $X=2.15 $Y=2.685 $X2=0 $Y2=0
cc_211 N_A_84_48#_c_148_n N_VPWR_c_771_n 0.00864234f $X=0.6 $Y=1.765 $X2=0 $Y2=0
cc_212 N_A_84_48#_c_218_p N_VPWR_c_771_n 0.00576021f $X=1.605 $Y=2.685 $X2=0
+ $Y2=0
cc_213 N_A_84_48#_c_155_n N_VPWR_c_771_n 0.0281637f $X=2.15 $Y=2.685 $X2=0 $Y2=0
cc_214 N_A_84_48#_c_159_p A_283_392# 0.00394468f $X=1.435 $Y=2.055 $X2=-0.19
+ $Y2=-0.245
cc_215 N_A_84_48#_c_183_p A_283_392# 0.0040492f $X=1.52 $Y=2.52 $X2=-0.19
+ $Y2=-0.245
cc_216 N_A_84_48#_c_218_p A_283_392# 0.00257104f $X=1.605 $Y=2.685 $X2=-0.19
+ $Y2=-0.245
cc_217 N_A_84_48#_c_155_n A_283_392# 0.00122781f $X=2.15 $Y=2.685 $X2=-0.19
+ $Y2=-0.245
cc_218 N_A_84_48#_c_147_n N_VGND_c_948_n 0.0112574f $X=0.495 $Y=1.22 $X2=0 $Y2=0
cc_219 N_A_84_48#_c_147_n N_VGND_c_954_n 0.00398535f $X=0.495 $Y=1.22 $X2=0
+ $Y2=0
cc_220 N_A_84_48#_c_147_n N_VGND_c_964_n 0.00404969f $X=0.495 $Y=1.22 $X2=0
+ $Y2=0
cc_221 N_A_84_48#_c_151_n A_286_80# 6.49906e-19 $X=1.52 $Y=1.19 $X2=-0.19
+ $Y2=-0.245
cc_222 N_A_84_48#_c_201_p A_286_80# 0.00147622f $X=1.605 $Y=0.815 $X2=-0.19
+ $Y2=-0.245
cc_223 N_A_84_48#_c_170_p A_286_80# 3.7187e-19 $X=2.06 $Y=0.815 $X2=-0.19
+ $Y2=-0.245
cc_224 N_GATE_M1017_g N_A_334_54#_c_265_n 0.0308885f $X=1.355 $Y=0.72 $X2=0
+ $Y2=0
cc_225 N_GATE_c_233_n N_A_334_54#_c_268_n 0.00379041f $X=1.34 $Y=1.885 $X2=0
+ $Y2=0
cc_226 N_GATE_M1017_g N_A_334_54#_c_268_n 7.74843e-19 $X=1.355 $Y=0.72 $X2=0
+ $Y2=0
cc_227 GATE N_A_334_54#_c_268_n 0.0120209f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_228 N_GATE_c_233_n N_A_334_54#_c_269_n 0.0308885f $X=1.34 $Y=1.885 $X2=0
+ $Y2=0
cc_229 N_GATE_c_233_n N_A_334_338#_c_394_n 0.0505819f $X=1.34 $Y=1.885 $X2=0
+ $Y2=0
cc_230 N_GATE_c_233_n N_A_334_338#_c_396_n 0.0111662f $X=1.34 $Y=1.885 $X2=0
+ $Y2=0
cc_231 GATE N_A_334_338#_c_396_n 4.93257e-19 $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_232 N_GATE_M1017_g N_A_27_74#_c_471_n 0.0147887f $X=1.355 $Y=0.72 $X2=0 $Y2=0
cc_233 N_GATE_c_233_n N_VPWR_c_772_n 0.0133474f $X=1.34 $Y=1.885 $X2=0 $Y2=0
cc_234 N_GATE_c_233_n N_VPWR_c_783_n 0.00461464f $X=1.34 $Y=1.885 $X2=0 $Y2=0
cc_235 N_GATE_c_233_n N_VPWR_c_771_n 0.00911633f $X=1.34 $Y=1.885 $X2=0 $Y2=0
cc_236 N_GATE_M1017_g N_VGND_c_948_n 9.39772e-19 $X=1.355 $Y=0.72 $X2=0 $Y2=0
cc_237 N_GATE_M1017_g N_VGND_c_955_n 9.29978e-19 $X=1.355 $Y=0.72 $X2=0 $Y2=0
cc_238 N_A_334_54#_c_279_n N_A_334_338#_M1004_d 0.00771987f $X=4.205 $Y=2.605
+ $X2=0 $Y2=0
cc_239 N_A_334_54#_c_274_n N_A_334_338#_c_394_n 0.0205629f $X=2.545 $Y=2.465
+ $X2=0 $Y2=0
cc_240 N_A_334_54#_c_268_n N_A_334_338#_c_394_n 0.00579991f $X=1.9 $Y=1.315
+ $X2=0 $Y2=0
cc_241 N_A_334_54#_c_293_n N_A_334_338#_c_394_n 0.00970937f $X=2.065 $Y=2.2
+ $X2=0 $Y2=0
cc_242 N_A_334_54#_c_268_n N_A_334_338#_c_387_n 0.0132375f $X=1.9 $Y=1.315 $X2=0
+ $Y2=0
cc_243 N_A_334_54#_c_277_n N_A_334_338#_c_387_n 0.00839201f $X=3.305 $Y=2.2
+ $X2=0 $Y2=0
cc_244 N_A_334_54#_c_268_n N_A_334_338#_c_396_n 0.00570704f $X=1.9 $Y=1.315
+ $X2=0 $Y2=0
cc_245 N_A_334_54#_c_269_n N_A_334_338#_c_396_n 0.0274437f $X=1.9 $Y=1.315 $X2=0
+ $Y2=0
cc_246 N_A_334_54#_c_265_n N_A_334_338#_M1012_g 0.016863f $X=1.745 $Y=1.15 $X2=0
+ $Y2=0
cc_247 N_A_334_54#_c_268_n N_A_334_338#_M1012_g 0.00174539f $X=1.9 $Y=1.315
+ $X2=0 $Y2=0
cc_248 N_A_334_54#_c_269_n N_A_334_338#_M1012_g 0.0178648f $X=1.9 $Y=1.315 $X2=0
+ $Y2=0
cc_249 N_A_334_54#_c_266_n N_A_334_338#_c_389_n 0.00372691f $X=3.585 $Y=2.045
+ $X2=0 $Y2=0
cc_250 N_A_334_54#_M1025_g N_A_334_338#_c_389_n 0.0100418f $X=3.695 $Y=0.995
+ $X2=0 $Y2=0
cc_251 N_A_334_54#_c_270_n N_A_334_338#_c_389_n 0.0286552f $X=3.39 $Y=2.35 $X2=0
+ $Y2=0
cc_252 N_A_334_54#_c_280_n N_A_334_338#_c_389_n 0.00615352f $X=4.37 $Y=2.255
+ $X2=0 $Y2=0
cc_253 N_A_334_54#_c_274_n N_A_334_338#_c_390_n 0.00116631f $X=2.545 $Y=2.465
+ $X2=0 $Y2=0
cc_254 N_A_334_54#_c_268_n N_A_334_338#_c_390_n 0.0259472f $X=1.9 $Y=1.315 $X2=0
+ $Y2=0
cc_255 N_A_334_54#_c_269_n N_A_334_338#_c_390_n 4.56399e-19 $X=1.9 $Y=1.315
+ $X2=0 $Y2=0
cc_256 N_A_334_54#_c_277_n N_A_334_338#_c_390_n 0.018746f $X=3.305 $Y=2.2 $X2=0
+ $Y2=0
cc_257 N_A_334_54#_c_270_n N_A_334_338#_c_390_n 0.0029232f $X=3.39 $Y=2.35 $X2=0
+ $Y2=0
cc_258 N_A_334_54#_c_274_n N_A_334_338#_c_391_n 0.0215139f $X=2.545 $Y=2.465
+ $X2=0 $Y2=0
cc_259 N_A_334_54#_c_268_n N_A_334_338#_c_391_n 0.0045632f $X=1.9 $Y=1.315 $X2=0
+ $Y2=0
cc_260 N_A_334_54#_c_277_n N_A_334_338#_c_391_n 0.00128281f $X=3.305 $Y=2.2
+ $X2=0 $Y2=0
cc_261 N_A_334_54#_c_266_n N_A_334_338#_c_399_n 0.00448808f $X=3.585 $Y=2.045
+ $X2=0 $Y2=0
cc_262 N_A_334_54#_c_270_n N_A_334_338#_c_399_n 5.72571e-19 $X=3.39 $Y=2.35
+ $X2=0 $Y2=0
cc_263 N_A_334_54#_c_279_n N_A_334_338#_c_399_n 0.0212439f $X=4.205 $Y=2.605
+ $X2=0 $Y2=0
cc_264 N_A_334_54#_c_280_n N_A_334_338#_c_399_n 0.0121633f $X=4.37 $Y=2.255
+ $X2=0 $Y2=0
cc_265 N_A_334_54#_c_266_n N_A_334_338#_c_392_n 0.00766568f $X=3.585 $Y=2.045
+ $X2=0 $Y2=0
cc_266 N_A_334_54#_M1025_g N_A_334_338#_c_392_n 0.0138443f $X=3.695 $Y=0.995
+ $X2=0 $Y2=0
cc_267 N_A_334_54#_c_277_n N_A_334_338#_c_392_n 0.0228749f $X=3.305 $Y=2.2 $X2=0
+ $Y2=0
cc_268 N_A_334_54#_c_270_n N_A_334_338#_c_392_n 0.0268965f $X=3.39 $Y=2.35 $X2=0
+ $Y2=0
cc_269 N_A_334_54#_M1025_g N_A_334_338#_c_393_n 0.002462f $X=3.695 $Y=0.995
+ $X2=0 $Y2=0
cc_270 N_A_334_54#_c_274_n N_A_27_74#_c_466_n 0.0231363f $X=2.545 $Y=2.465 $X2=0
+ $Y2=0
cc_271 N_A_334_54#_c_266_n N_A_27_74#_c_466_n 0.0249148f $X=3.585 $Y=2.045 $X2=0
+ $Y2=0
cc_272 N_A_334_54#_c_277_n N_A_27_74#_c_466_n 0.0256803f $X=3.305 $Y=2.2 $X2=0
+ $Y2=0
cc_273 N_A_334_54#_c_270_n N_A_27_74#_c_466_n 0.0062763f $X=3.39 $Y=2.35 $X2=0
+ $Y2=0
cc_274 N_A_334_54#_c_338_p N_A_27_74#_c_466_n 0.00233459f $X=3.39 $Y=2.52 $X2=0
+ $Y2=0
cc_275 N_A_334_54#_c_274_n N_A_27_74#_c_480_n 0.0295229f $X=2.545 $Y=2.465 $X2=0
+ $Y2=0
cc_276 N_A_334_54#_c_266_n N_A_27_74#_c_480_n 0.0133467f $X=3.585 $Y=2.045 $X2=0
+ $Y2=0
cc_277 N_A_334_54#_c_338_p N_A_27_74#_c_480_n 0.0010822f $X=3.39 $Y=2.52 $X2=0
+ $Y2=0
cc_278 N_A_334_54#_c_342_p N_A_27_74#_c_480_n 0.00446046f $X=3.475 $Y=2.605
+ $X2=0 $Y2=0
cc_279 N_A_334_54#_M1025_g N_A_27_74#_M1000_g 0.0171519f $X=3.695 $Y=0.995 $X2=0
+ $Y2=0
cc_280 N_A_334_54#_c_265_n N_A_27_74#_c_471_n 0.0119481f $X=1.745 $Y=1.15 $X2=0
+ $Y2=0
cc_281 N_A_334_54#_M1025_g N_A_27_74#_c_474_n 0.00318939f $X=3.695 $Y=0.995
+ $X2=0 $Y2=0
cc_282 N_A_334_54#_M1019_s N_A_27_74#_c_475_n 0.00239646f $X=4.3 $Y=0.37 $X2=0
+ $Y2=0
cc_283 N_A_334_54#_M1025_g N_A_27_74#_c_475_n 0.0175247f $X=3.695 $Y=0.995 $X2=0
+ $Y2=0
cc_284 N_A_334_54#_c_271_n N_A_27_74#_c_475_n 0.0151779f $X=4.28 $Y=0.385 $X2=0
+ $Y2=0
cc_285 N_A_334_54#_c_272_n N_A_27_74#_c_475_n 0.00634638f $X=3.98 $Y=0.35 $X2=0
+ $Y2=0
cc_286 N_A_334_54#_c_273_n N_A_27_74#_c_475_n 0.0258904f $X=4.445 $Y=0.685 $X2=0
+ $Y2=0
cc_287 N_A_334_54#_c_272_n N_A_27_74#_c_478_n 0.00690617f $X=3.98 $Y=0.35 $X2=0
+ $Y2=0
cc_288 N_A_334_54#_c_279_n N_CLK_c_609_n 0.00743413f $X=4.205 $Y=2.605 $X2=0
+ $Y2=0
cc_289 N_A_334_54#_c_280_n N_CLK_c_609_n 0.00706416f $X=4.37 $Y=2.255 $X2=0
+ $Y2=0
cc_290 N_A_334_54#_c_271_n N_CLK_M1019_g 0.0023f $X=4.28 $Y=0.385 $X2=0 $Y2=0
cc_291 N_A_334_54#_c_272_n N_CLK_M1019_g 0.00464769f $X=3.98 $Y=0.35 $X2=0 $Y2=0
cc_292 N_A_334_54#_c_280_n N_CLK_c_606_n 0.0077433f $X=4.37 $Y=2.255 $X2=0 $Y2=0
cc_293 N_A_334_54#_M1025_g N_CLK_c_607_n 0.00408582f $X=3.695 $Y=0.995 $X2=0
+ $Y2=0
cc_294 N_A_334_54#_c_280_n N_CLK_c_607_n 6.37339e-19 $X=4.37 $Y=2.255 $X2=0
+ $Y2=0
cc_295 N_A_334_54#_c_277_n N_VPWR_M1010_d 0.00177961f $X=3.305 $Y=2.2 $X2=0
+ $Y2=0
cc_296 N_A_334_54#_c_270_n N_VPWR_M1010_d 0.00165901f $X=3.39 $Y=2.35 $X2=0
+ $Y2=0
cc_297 N_A_334_54#_c_338_p N_VPWR_M1010_d 0.00230127f $X=3.39 $Y=2.52 $X2=0
+ $Y2=0
cc_298 N_A_334_54#_c_342_p N_VPWR_M1010_d 0.00440567f $X=3.475 $Y=2.605 $X2=0
+ $Y2=0
cc_299 N_A_334_54#_c_266_n N_VPWR_c_773_n 0.00660808f $X=3.585 $Y=2.045 $X2=0
+ $Y2=0
cc_300 N_A_334_54#_c_277_n N_VPWR_c_773_n 0.00734096f $X=3.305 $Y=2.2 $X2=0
+ $Y2=0
cc_301 N_A_334_54#_c_342_p N_VPWR_c_773_n 0.0113006f $X=3.475 $Y=2.605 $X2=0
+ $Y2=0
cc_302 N_A_334_54#_c_279_n N_VPWR_c_774_n 0.0310448f $X=4.205 $Y=2.605 $X2=0
+ $Y2=0
cc_303 N_A_334_54#_c_280_n N_VPWR_c_774_n 0.0288995f $X=4.37 $Y=2.255 $X2=0
+ $Y2=0
cc_304 N_A_334_54#_c_266_n N_VPWR_c_781_n 0.00326738f $X=3.585 $Y=2.045 $X2=0
+ $Y2=0
cc_305 N_A_334_54#_c_279_n N_VPWR_c_781_n 0.0260353f $X=4.205 $Y=2.605 $X2=0
+ $Y2=0
cc_306 N_A_334_54#_c_342_p N_VPWR_c_781_n 4.5124e-19 $X=3.475 $Y=2.605 $X2=0
+ $Y2=0
cc_307 N_A_334_54#_c_274_n N_VPWR_c_783_n 0.00446156f $X=2.545 $Y=2.465 $X2=0
+ $Y2=0
cc_308 N_A_334_54#_c_274_n N_VPWR_c_771_n 0.00893546f $X=2.545 $Y=2.465 $X2=0
+ $Y2=0
cc_309 N_A_334_54#_c_266_n N_VPWR_c_771_n 0.00420856f $X=3.585 $Y=2.045 $X2=0
+ $Y2=0
cc_310 N_A_334_54#_c_279_n N_VPWR_c_771_n 0.0321175f $X=4.205 $Y=2.605 $X2=0
+ $Y2=0
cc_311 N_A_334_54#_c_342_p N_VPWR_c_771_n 0.00178054f $X=3.475 $Y=2.605 $X2=0
+ $Y2=0
cc_312 N_A_334_54#_M1025_g N_VGND_c_949_n 0.00921355f $X=3.695 $Y=0.995 $X2=0
+ $Y2=0
cc_313 N_A_334_54#_c_271_n N_VGND_c_949_n 0.0205948f $X=4.28 $Y=0.385 $X2=0
+ $Y2=0
cc_314 N_A_334_54#_c_272_n N_VGND_c_949_n 0.0115834f $X=3.98 $Y=0.35 $X2=0 $Y2=0
cc_315 N_A_334_54#_c_273_n N_VGND_c_949_n 0.00972897f $X=4.445 $Y=0.685 $X2=0
+ $Y2=0
cc_316 N_A_334_54#_c_271_n N_VGND_c_950_n 0.0151168f $X=4.28 $Y=0.385 $X2=0
+ $Y2=0
cc_317 N_A_334_54#_c_272_n N_VGND_c_950_n 9.77729e-19 $X=3.98 $Y=0.35 $X2=0
+ $Y2=0
cc_318 N_A_334_54#_c_265_n N_VGND_c_955_n 9.29978e-19 $X=1.745 $Y=1.15 $X2=0
+ $Y2=0
cc_319 N_A_334_54#_c_271_n N_VGND_c_956_n 0.0532296f $X=4.28 $Y=0.385 $X2=0
+ $Y2=0
cc_320 N_A_334_54#_c_272_n N_VGND_c_956_n 0.0118937f $X=3.98 $Y=0.35 $X2=0 $Y2=0
cc_321 N_A_334_54#_c_271_n N_VGND_c_964_n 0.0289216f $X=4.28 $Y=0.385 $X2=0
+ $Y2=0
cc_322 N_A_334_54#_c_272_n N_VGND_c_964_n 0.0190295f $X=3.98 $Y=0.35 $X2=0 $Y2=0
cc_323 N_A_334_338#_M1012_g N_A_27_74#_c_465_n 8.86417e-19 $X=2.38 $Y=0.83 $X2=0
+ $Y2=0
cc_324 N_A_334_338#_c_390_n N_A_27_74#_c_465_n 0.00163581f $X=2.47 $Y=1.445
+ $X2=0 $Y2=0
cc_325 N_A_334_338#_c_391_n N_A_27_74#_c_465_n 0.0209296f $X=2.47 $Y=1.64 $X2=0
+ $Y2=0
cc_326 N_A_334_338#_c_392_n N_A_27_74#_c_465_n 0.00918689f $X=3.825 $Y=1.485
+ $X2=0 $Y2=0
cc_327 N_A_334_338#_M1012_g N_A_27_74#_M1000_g 0.0213372f $X=2.38 $Y=0.83 $X2=0
+ $Y2=0
cc_328 N_A_334_338#_c_392_n N_A_27_74#_M1000_g 0.00564586f $X=3.825 $Y=1.485
+ $X2=0 $Y2=0
cc_329 N_A_334_338#_M1012_g N_A_27_74#_c_471_n 0.00658236f $X=2.38 $Y=0.83 $X2=0
+ $Y2=0
cc_330 N_A_334_338#_M1012_g N_A_27_74#_c_474_n 0.00591925f $X=2.38 $Y=0.83 $X2=0
+ $Y2=0
cc_331 N_A_334_338#_M1025_d N_A_27_74#_c_475_n 0.0056672f $X=3.77 $Y=0.625 $X2=0
+ $Y2=0
cc_332 N_A_334_338#_c_392_n N_A_27_74#_c_475_n 0.0652325f $X=3.825 $Y=1.485
+ $X2=0 $Y2=0
cc_333 N_A_334_338#_M1012_g N_A_27_74#_c_534_n 0.00396757f $X=2.38 $Y=0.83 $X2=0
+ $Y2=0
cc_334 N_A_334_338#_c_392_n N_A_27_74#_c_534_n 0.0167062f $X=3.825 $Y=1.485
+ $X2=0 $Y2=0
cc_335 N_A_334_338#_M1012_g N_A_27_74#_c_478_n 0.00202272f $X=2.38 $Y=0.83 $X2=0
+ $Y2=0
cc_336 N_A_334_338#_c_389_n N_CLK_c_608_n 0.00673379f $X=3.91 $Y=2.18 $X2=0
+ $Y2=0
cc_337 N_A_334_338#_c_389_n N_CLK_c_609_n 0.00145717f $X=3.91 $Y=2.18 $X2=0
+ $Y2=0
cc_338 N_A_334_338#_c_389_n N_CLK_c_606_n 0.00747805f $X=3.91 $Y=2.18 $X2=0
+ $Y2=0
cc_339 N_A_334_338#_c_393_n N_CLK_c_606_n 0.0164788f $X=3.99 $Y=1.445 $X2=0
+ $Y2=0
cc_340 N_A_334_338#_c_389_n N_CLK_c_607_n 2.7829e-19 $X=3.91 $Y=2.18 $X2=0 $Y2=0
cc_341 N_A_334_338#_c_393_n N_CLK_c_607_n 0.00121403f $X=3.99 $Y=1.445 $X2=0
+ $Y2=0
cc_342 N_A_334_338#_c_394_n N_VPWR_c_783_n 0.00308386f $X=1.76 $Y=1.885 $X2=0
+ $Y2=0
cc_343 N_A_334_338#_c_394_n N_VPWR_c_771_n 0.00381773f $X=1.76 $Y=1.885 $X2=0
+ $Y2=0
cc_344 N_A_334_338#_c_392_n N_VGND_M1000_d 0.00483981f $X=3.825 $Y=1.485 $X2=0
+ $Y2=0
cc_345 N_A_334_338#_c_390_n A_491_124# 0.00338728f $X=2.47 $Y=1.445 $X2=-0.19
+ $Y2=-0.245
cc_346 N_A_334_338#_c_392_n A_491_124# 0.00720817f $X=3.825 $Y=1.485 $X2=-0.19
+ $Y2=-0.245
cc_347 N_A_27_74#_c_475_n N_CLK_M1019_g 0.0163338f $X=5.26 $Y=1.105 $X2=0 $Y2=0
cc_348 N_A_27_74#_c_469_n N_CLK_c_610_n 0.00879087f $X=5.63 $Y=1.765 $X2=0 $Y2=0
cc_349 N_A_27_74#_M1023_g N_CLK_M1005_g 0.0350457f $X=5.55 $Y=0.74 $X2=0 $Y2=0
cc_350 N_A_27_74#_c_475_n N_CLK_M1005_g 0.0253438f $X=5.26 $Y=1.105 $X2=0 $Y2=0
cc_351 N_A_27_74#_c_469_n N_CLK_c_606_n 8.58876e-19 $X=5.63 $Y=1.765 $X2=0 $Y2=0
cc_352 N_A_27_74#_c_475_n N_CLK_c_606_n 0.0723728f $X=5.26 $Y=1.105 $X2=0 $Y2=0
cc_353 N_A_27_74#_c_469_n N_CLK_c_607_n 0.0411752f $X=5.63 $Y=1.765 $X2=0 $Y2=0
cc_354 N_A_27_74#_c_475_n N_CLK_c_607_n 0.00864636f $X=5.26 $Y=1.105 $X2=0 $Y2=0
cc_355 N_A_27_74#_c_469_n N_A_1044_368#_c_671_n 0.00165784f $X=5.63 $Y=1.765
+ $X2=0 $Y2=0
cc_356 N_A_27_74#_c_475_n N_A_1044_368#_c_671_n 0.0262851f $X=5.26 $Y=1.105
+ $X2=0 $Y2=0
cc_357 N_A_27_74#_c_469_n N_A_1044_368#_c_672_n 0.0163193f $X=5.63 $Y=1.765
+ $X2=0 $Y2=0
cc_358 N_A_27_74#_c_469_n N_A_1044_368#_c_673_n 0.0149402f $X=5.63 $Y=1.765
+ $X2=0 $Y2=0
cc_359 N_A_27_74#_c_475_n N_A_1044_368#_c_673_n 0.0157721f $X=5.26 $Y=1.105
+ $X2=0 $Y2=0
cc_360 N_A_27_74#_M1023_g N_A_1044_368#_c_659_n 0.0148811f $X=5.55 $Y=0.74 $X2=0
+ $Y2=0
cc_361 N_A_27_74#_c_469_n N_A_1044_368#_c_659_n 0.00141647f $X=5.63 $Y=1.765
+ $X2=0 $Y2=0
cc_362 N_A_27_74#_c_475_n N_A_1044_368#_c_659_n 0.0228054f $X=5.26 $Y=1.105
+ $X2=0 $Y2=0
cc_363 N_A_27_74#_M1023_g N_A_1044_368#_c_660_n 0.00143549f $X=5.55 $Y=0.74
+ $X2=0 $Y2=0
cc_364 N_A_27_74#_c_469_n N_A_1044_368#_c_660_n 0.00702988f $X=5.63 $Y=1.765
+ $X2=0 $Y2=0
cc_365 N_A_27_74#_c_475_n N_A_1044_368#_c_660_n 0.0337495f $X=5.26 $Y=1.105
+ $X2=0 $Y2=0
cc_366 N_A_27_74#_M1023_g N_A_1044_368#_c_661_n 0.0121306f $X=5.55 $Y=0.74 $X2=0
+ $Y2=0
cc_367 N_A_27_74#_c_469_n N_A_1044_368#_c_661_n 0.0208223f $X=5.63 $Y=1.765
+ $X2=0 $Y2=0
cc_368 N_A_27_74#_c_475_n N_A_1044_368#_c_661_n 3.72912e-19 $X=5.26 $Y=1.105
+ $X2=0 $Y2=0
cc_369 N_A_27_74#_c_469_n N_A_1044_368#_c_662_n 0.00192399f $X=5.63 $Y=1.765
+ $X2=0 $Y2=0
cc_370 N_A_27_74#_c_482_n N_VPWR_c_772_n 0.0404609f $X=0.375 $Y=2.815 $X2=0
+ $Y2=0
cc_371 N_A_27_74#_c_480_n N_VPWR_c_773_n 0.00660808f $X=2.965 $Y=2.465 $X2=0
+ $Y2=0
cc_372 N_A_27_74#_c_469_n N_VPWR_c_775_n 0.0196637f $X=5.63 $Y=1.765 $X2=0 $Y2=0
cc_373 N_A_27_74#_c_482_n N_VPWR_c_779_n 0.0188328f $X=0.375 $Y=2.815 $X2=0
+ $Y2=0
cc_374 N_A_27_74#_c_480_n N_VPWR_c_783_n 0.00461464f $X=2.965 $Y=2.465 $X2=0
+ $Y2=0
cc_375 N_A_27_74#_c_469_n N_VPWR_c_784_n 0.00445602f $X=5.63 $Y=1.765 $X2=0
+ $Y2=0
cc_376 N_A_27_74#_c_480_n N_VPWR_c_771_n 0.00985926f $X=2.965 $Y=2.465 $X2=0
+ $Y2=0
cc_377 N_A_27_74#_c_469_n N_VPWR_c_771_n 0.00862108f $X=5.63 $Y=1.765 $X2=0
+ $Y2=0
cc_378 N_A_27_74#_c_482_n N_VPWR_c_771_n 0.0155553f $X=0.375 $Y=2.815 $X2=0
+ $Y2=0
cc_379 N_A_27_74#_c_489_n N_VGND_M1021_d 0.0166022f $X=1.095 $Y=0.935 $X2=-0.19
+ $Y2=-0.245
cc_380 N_A_27_74#_c_493_n N_VGND_M1021_d 0.00684638f $X=1.18 $Y=0.85 $X2=-0.19
+ $Y2=-0.245
cc_381 N_A_27_74#_c_472_n N_VGND_M1021_d 2.48347e-19 $X=1.265 $Y=0.34 $X2=-0.19
+ $Y2=-0.245
cc_382 N_A_27_74#_c_474_n N_VGND_M1000_d 0.00120802f $X=2.98 $Y=1.02 $X2=0 $Y2=0
cc_383 N_A_27_74#_c_475_n N_VGND_M1000_d 0.015135f $X=5.26 $Y=1.105 $X2=0 $Y2=0
cc_384 N_A_27_74#_c_534_n N_VGND_M1000_d 3.54991e-19 $X=3.145 $Y=1.105 $X2=0
+ $Y2=0
cc_385 N_A_27_74#_c_475_n N_VGND_M1019_d 0.00176461f $X=5.26 $Y=1.105 $X2=0
+ $Y2=0
cc_386 N_A_27_74#_c_470_n N_VGND_c_948_n 0.0125137f $X=0.28 $Y=0.515 $X2=0 $Y2=0
cc_387 N_A_27_74#_c_489_n N_VGND_c_948_n 0.0250287f $X=1.095 $Y=0.935 $X2=0
+ $Y2=0
cc_388 N_A_27_74#_c_493_n N_VGND_c_948_n 0.0196481f $X=1.18 $Y=0.85 $X2=0 $Y2=0
cc_389 N_A_27_74#_c_472_n N_VGND_c_948_n 0.0150932f $X=1.265 $Y=0.34 $X2=0 $Y2=0
cc_390 N_A_27_74#_M1000_g N_VGND_c_949_n 0.00104285f $X=2.98 $Y=1.155 $X2=0
+ $Y2=0
cc_391 N_A_27_74#_c_473_n N_VGND_c_949_n 0.0142656f $X=2.98 $Y=0.425 $X2=0 $Y2=0
cc_392 N_A_27_74#_c_474_n N_VGND_c_949_n 0.0348535f $X=2.98 $Y=1.02 $X2=0 $Y2=0
cc_393 N_A_27_74#_c_475_n N_VGND_c_949_n 0.0219153f $X=5.26 $Y=1.105 $X2=0 $Y2=0
cc_394 N_A_27_74#_c_478_n N_VGND_c_949_n 0.00260146f $X=2.98 $Y=0.38 $X2=0 $Y2=0
cc_395 N_A_27_74#_M1023_g N_VGND_c_950_n 0.00197566f $X=5.55 $Y=0.74 $X2=0 $Y2=0
cc_396 N_A_27_74#_c_475_n N_VGND_c_950_n 0.0170777f $X=5.26 $Y=1.105 $X2=0 $Y2=0
cc_397 N_A_27_74#_c_470_n N_VGND_c_954_n 0.011066f $X=0.28 $Y=0.515 $X2=0 $Y2=0
cc_398 N_A_27_74#_c_471_n N_VGND_c_955_n 0.0997901f $X=2.815 $Y=0.34 $X2=0 $Y2=0
cc_399 N_A_27_74#_c_472_n N_VGND_c_955_n 0.0121867f $X=1.265 $Y=0.34 $X2=0 $Y2=0
cc_400 N_A_27_74#_c_473_n N_VGND_c_955_n 0.0224969f $X=2.98 $Y=0.425 $X2=0 $Y2=0
cc_401 N_A_27_74#_c_478_n N_VGND_c_955_n 0.00612073f $X=2.98 $Y=0.38 $X2=0 $Y2=0
cc_402 N_A_27_74#_M1023_g N_VGND_c_957_n 0.00748462f $X=5.55 $Y=0.74 $X2=0 $Y2=0
cc_403 N_A_27_74#_M1023_g N_VGND_c_964_n 0.0082231f $X=5.55 $Y=0.74 $X2=0 $Y2=0
cc_404 N_A_27_74#_c_470_n N_VGND_c_964_n 0.00915947f $X=0.28 $Y=0.515 $X2=0
+ $Y2=0
cc_405 N_A_27_74#_c_489_n N_VGND_c_964_n 0.0124076f $X=1.095 $Y=0.935 $X2=0
+ $Y2=0
cc_406 N_A_27_74#_c_471_n N_VGND_c_964_n 0.0582686f $X=2.815 $Y=0.34 $X2=0 $Y2=0
cc_407 N_A_27_74#_c_472_n N_VGND_c_964_n 0.00660921f $X=1.265 $Y=0.34 $X2=0
+ $Y2=0
cc_408 N_A_27_74#_c_473_n N_VGND_c_964_n 0.0113197f $X=2.98 $Y=0.425 $X2=0 $Y2=0
cc_409 N_A_27_74#_c_478_n N_VGND_c_964_n 0.00853275f $X=2.98 $Y=0.38 $X2=0 $Y2=0
cc_410 N_A_27_74#_c_471_n A_286_80# 0.00150293f $X=2.815 $Y=0.34 $X2=-0.19
+ $Y2=-0.245
cc_411 N_A_27_74#_c_474_n A_491_124# 0.00107962f $X=2.98 $Y=1.02 $X2=-0.19
+ $Y2=-0.245
cc_412 N_A_27_74#_c_534_n A_491_124# 0.00308074f $X=3.145 $Y=1.105 $X2=-0.19
+ $Y2=-0.245
cc_413 N_A_27_74#_c_475_n A_1047_74# 0.0056254f $X=5.26 $Y=1.105 $X2=-0.19
+ $Y2=-0.245
cc_414 N_CLK_c_610_n N_A_1044_368#_c_671_n 6.47605e-19 $X=5.145 $Y=1.765 $X2=0
+ $Y2=0
cc_415 N_CLK_c_610_n N_A_1044_368#_c_672_n 4.36461e-19 $X=5.145 $Y=1.765 $X2=0
+ $Y2=0
cc_416 N_CLK_M1005_g N_A_1044_368#_c_659_n 0.00233225f $X=5.16 $Y=0.74 $X2=0
+ $Y2=0
cc_417 N_CLK_c_609_n N_VPWR_c_774_n 0.0112334f $X=4.595 $Y=2.035 $X2=0 $Y2=0
cc_418 N_CLK_c_610_n N_VPWR_c_774_n 0.00335681f $X=5.145 $Y=1.765 $X2=0 $Y2=0
cc_419 N_CLK_c_606_n N_VPWR_c_774_n 0.0172311f $X=4.905 $Y=1.515 $X2=0 $Y2=0
cc_420 N_CLK_c_607_n N_VPWR_c_774_n 0.00175302f $X=5.145 $Y=1.557 $X2=0 $Y2=0
cc_421 N_CLK_c_609_n N_VPWR_c_781_n 0.00554343f $X=4.595 $Y=2.035 $X2=0 $Y2=0
cc_422 N_CLK_c_610_n N_VPWR_c_784_n 0.00460063f $X=5.145 $Y=1.765 $X2=0 $Y2=0
cc_423 N_CLK_c_609_n N_VPWR_c_771_n 0.00542671f $X=4.595 $Y=2.035 $X2=0 $Y2=0
cc_424 N_CLK_c_610_n N_VPWR_c_771_n 0.00912686f $X=5.145 $Y=1.765 $X2=0 $Y2=0
cc_425 N_CLK_M1019_g N_VGND_c_950_n 0.0104121f $X=4.73 $Y=0.74 $X2=0 $Y2=0
cc_426 N_CLK_M1005_g N_VGND_c_950_n 0.0140817f $X=5.16 $Y=0.74 $X2=0 $Y2=0
cc_427 N_CLK_M1019_g N_VGND_c_956_n 0.00383152f $X=4.73 $Y=0.74 $X2=0 $Y2=0
cc_428 N_CLK_M1005_g N_VGND_c_957_n 0.00383152f $X=5.16 $Y=0.74 $X2=0 $Y2=0
cc_429 N_CLK_M1019_g N_VGND_c_964_n 0.00759393f $X=4.73 $Y=0.74 $X2=0 $Y2=0
cc_430 N_CLK_M1005_g N_VGND_c_964_n 0.0075725f $X=5.16 $Y=0.74 $X2=0 $Y2=0
cc_431 N_A_1044_368#_c_673_n N_VPWR_M1007_d 0.0118246f $X=5.975 $Y=1.905 $X2=0
+ $Y2=0
cc_432 N_A_1044_368#_c_672_n N_VPWR_c_774_n 0.0307037f $X=5.405 $Y=2.815 $X2=0
+ $Y2=0
cc_433 N_A_1044_368#_c_664_n N_VPWR_c_775_n 0.0196637f $X=6.735 $Y=1.765 $X2=0
+ $Y2=0
cc_434 N_A_1044_368#_c_672_n N_VPWR_c_775_n 0.0316504f $X=5.405 $Y=2.815 $X2=0
+ $Y2=0
cc_435 N_A_1044_368#_c_673_n N_VPWR_c_775_n 0.0511035f $X=5.975 $Y=1.905 $X2=0
+ $Y2=0
cc_436 N_A_1044_368#_c_662_n N_VPWR_c_775_n 0.00992125f $X=6.185 $Y=1.4 $X2=0
+ $Y2=0
cc_437 N_A_1044_368#_c_665_n N_VPWR_c_776_n 0.00187195f $X=7.2 $Y=1.765 $X2=0
+ $Y2=0
cc_438 N_A_1044_368#_c_654_n N_VPWR_c_776_n 0.00165934f $X=7.595 $Y=1.54 $X2=0
+ $Y2=0
cc_439 N_A_1044_368#_c_668_n N_VPWR_c_776_n 0.00538946f $X=7.685 $Y=1.765 $X2=0
+ $Y2=0
cc_440 N_A_1044_368#_c_668_n N_VPWR_c_778_n 6.80807e-19 $X=7.685 $Y=1.765 $X2=0
+ $Y2=0
cc_441 N_A_1044_368#_c_669_n N_VPWR_c_778_n 0.015599f $X=8.135 $Y=1.765 $X2=0
+ $Y2=0
cc_442 N_A_1044_368#_c_672_n N_VPWR_c_784_n 0.0145938f $X=5.405 $Y=2.815 $X2=0
+ $Y2=0
cc_443 N_A_1044_368#_c_664_n N_VPWR_c_785_n 0.00445602f $X=6.735 $Y=1.765 $X2=0
+ $Y2=0
cc_444 N_A_1044_368#_c_665_n N_VPWR_c_785_n 0.00461464f $X=7.2 $Y=1.765 $X2=0
+ $Y2=0
cc_445 N_A_1044_368#_c_668_n N_VPWR_c_786_n 0.00445602f $X=7.685 $Y=1.765 $X2=0
+ $Y2=0
cc_446 N_A_1044_368#_c_669_n N_VPWR_c_786_n 0.00413917f $X=8.135 $Y=1.765 $X2=0
+ $Y2=0
cc_447 N_A_1044_368#_c_664_n N_VPWR_c_771_n 0.00861862f $X=6.735 $Y=1.765 $X2=0
+ $Y2=0
cc_448 N_A_1044_368#_c_665_n N_VPWR_c_771_n 0.00908413f $X=7.2 $Y=1.765 $X2=0
+ $Y2=0
cc_449 N_A_1044_368#_c_668_n N_VPWR_c_771_n 0.00857917f $X=7.685 $Y=1.765 $X2=0
+ $Y2=0
cc_450 N_A_1044_368#_c_669_n N_VPWR_c_771_n 0.00817726f $X=8.135 $Y=1.765 $X2=0
+ $Y2=0
cc_451 N_A_1044_368#_c_672_n N_VPWR_c_771_n 0.0120466f $X=5.405 $Y=2.815 $X2=0
+ $Y2=0
cc_452 N_A_1044_368#_c_664_n N_GCLK_c_884_n 0.0209486f $X=6.735 $Y=1.765 $X2=0
+ $Y2=0
cc_453 N_A_1044_368#_c_665_n N_GCLK_c_884_n 0.00161111f $X=7.2 $Y=1.765 $X2=0
+ $Y2=0
cc_454 N_A_1044_368#_c_655_n N_GCLK_c_884_n 0.00346335f $X=7.29 $Y=1.54 $X2=0
+ $Y2=0
cc_455 N_A_1044_368#_c_673_n N_GCLK_c_884_n 0.00670806f $X=5.975 $Y=1.905 $X2=0
+ $Y2=0
cc_456 N_A_1044_368#_c_660_n N_GCLK_c_884_n 0.00384271f $X=6.185 $Y=1.515 $X2=0
+ $Y2=0
cc_457 N_A_1044_368#_M1006_g N_GCLK_c_877_n 0.0205429f $X=6.785 $Y=0.74 $X2=0
+ $Y2=0
cc_458 N_A_1044_368#_M1008_g N_GCLK_c_877_n 0.0126177f $X=7.215 $Y=0.74 $X2=0
+ $Y2=0
cc_459 N_A_1044_368#_M1013_g N_GCLK_c_877_n 6.13796e-19 $X=7.715 $Y=0.74 $X2=0
+ $Y2=0
cc_460 N_A_1044_368#_c_659_n N_GCLK_c_877_n 0.015596f $X=6.162 $Y=1.13 $X2=0
+ $Y2=0
cc_461 N_A_1044_368#_c_660_n N_GCLK_c_877_n 0.00255045f $X=6.185 $Y=1.515 $X2=0
+ $Y2=0
cc_462 N_A_1044_368#_c_661_n N_GCLK_c_877_n 7.55566e-19 $X=6.185 $Y=0.835 $X2=0
+ $Y2=0
cc_463 N_A_1044_368#_c_654_n N_GCLK_c_885_n 0.0112701f $X=7.595 $Y=1.54 $X2=0
+ $Y2=0
cc_464 N_A_1044_368#_c_655_n N_GCLK_c_885_n 0.0121787f $X=7.29 $Y=1.54 $X2=0
+ $Y2=0
cc_465 N_A_1044_368#_c_658_n N_GCLK_c_885_n 0.0111023f $X=8.135 $Y=1.582 $X2=0
+ $Y2=0
cc_466 N_A_1044_368#_c_655_n N_GCLK_c_903_n 0.0213393f $X=7.29 $Y=1.54 $X2=0
+ $Y2=0
cc_467 N_A_1044_368#_c_660_n N_GCLK_c_903_n 0.00643488f $X=6.185 $Y=1.515 $X2=0
+ $Y2=0
cc_468 N_A_1044_368#_M1008_g N_GCLK_c_878_n 0.0113403f $X=7.215 $Y=0.74 $X2=0
+ $Y2=0
cc_469 N_A_1044_368#_c_654_n N_GCLK_c_878_n 0.0044116f $X=7.595 $Y=1.54 $X2=0
+ $Y2=0
cc_470 N_A_1044_368#_M1013_g N_GCLK_c_878_n 0.0113115f $X=7.715 $Y=0.74 $X2=0
+ $Y2=0
cc_471 N_A_1044_368#_M1006_g N_GCLK_c_879_n 0.00524345f $X=6.785 $Y=0.74 $X2=0
+ $Y2=0
cc_472 N_A_1044_368#_M1008_g N_GCLK_c_879_n 0.00272521f $X=7.215 $Y=0.74 $X2=0
+ $Y2=0
cc_473 N_A_1044_368#_c_655_n N_GCLK_c_879_n 0.00271192f $X=7.29 $Y=1.54 $X2=0
+ $Y2=0
cc_474 N_A_1044_368#_c_660_n N_GCLK_c_879_n 0.00581761f $X=6.185 $Y=1.515 $X2=0
+ $Y2=0
cc_475 N_A_1044_368#_c_661_n N_GCLK_c_879_n 5.80746e-19 $X=6.185 $Y=0.835 $X2=0
+ $Y2=0
cc_476 N_A_1044_368#_c_665_n N_GCLK_c_886_n 5.69921e-19 $X=7.2 $Y=1.765 $X2=0
+ $Y2=0
cc_477 N_A_1044_368#_c_668_n N_GCLK_c_886_n 0.0145294f $X=7.685 $Y=1.765 $X2=0
+ $Y2=0
cc_478 N_A_1044_368#_c_669_n N_GCLK_c_886_n 0.00771123f $X=8.135 $Y=1.765 $X2=0
+ $Y2=0
cc_479 N_A_1044_368#_M1008_g N_GCLK_c_880_n 6.95109e-19 $X=7.215 $Y=0.74 $X2=0
+ $Y2=0
cc_480 N_A_1044_368#_M1013_g N_GCLK_c_880_n 0.0122683f $X=7.715 $Y=0.74 $X2=0
+ $Y2=0
cc_481 N_A_1044_368#_M1015_g N_GCLK_c_880_n 0.00292368f $X=8.145 $Y=0.74 $X2=0
+ $Y2=0
cc_482 N_A_1044_368#_M1013_g N_GCLK_c_881_n 4.96773e-19 $X=7.715 $Y=0.74 $X2=0
+ $Y2=0
cc_483 N_A_1044_368#_M1015_g N_GCLK_c_881_n 4.72088e-19 $X=8.145 $Y=0.74 $X2=0
+ $Y2=0
cc_484 N_A_1044_368#_c_658_n N_GCLK_c_881_n 0.0180848f $X=8.135 $Y=1.582 $X2=0
+ $Y2=0
cc_485 N_A_1044_368#_M1013_g N_GCLK_c_882_n 0.00223615f $X=7.715 $Y=0.74 $X2=0
+ $Y2=0
cc_486 N_A_1044_368#_M1015_g N_GCLK_c_882_n 0.0053794f $X=8.145 $Y=0.74 $X2=0
+ $Y2=0
cc_487 N_A_1044_368#_c_668_n GCLK 4.18229e-19 $X=7.685 $Y=1.765 $X2=0 $Y2=0
cc_488 N_A_1044_368#_c_658_n GCLK 0.0121871f $X=8.135 $Y=1.582 $X2=0 $Y2=0
cc_489 N_A_1044_368#_c_669_n GCLK 0.00703386f $X=8.135 $Y=1.765 $X2=0 $Y2=0
cc_490 N_A_1044_368#_c_658_n GCLK 0.019053f $X=8.135 $Y=1.582 $X2=0 $Y2=0
cc_491 N_A_1044_368#_c_659_n N_VGND_c_950_n 0.0163082f $X=6.162 $Y=1.13 $X2=0
+ $Y2=0
cc_492 N_A_1044_368#_M1008_g N_VGND_c_951_n 0.00659576f $X=7.215 $Y=0.74 $X2=0
+ $Y2=0
cc_493 N_A_1044_368#_M1013_g N_VGND_c_951_n 0.00170206f $X=7.715 $Y=0.74 $X2=0
+ $Y2=0
cc_494 N_A_1044_368#_M1013_g N_VGND_c_953_n 5.78878e-19 $X=7.715 $Y=0.74 $X2=0
+ $Y2=0
cc_495 N_A_1044_368#_M1015_g N_VGND_c_953_n 0.0128863f $X=8.145 $Y=0.74 $X2=0
+ $Y2=0
cc_496 N_A_1044_368#_M1006_g N_VGND_c_957_n 0.00777188f $X=6.785 $Y=0.74 $X2=0
+ $Y2=0
cc_497 N_A_1044_368#_c_659_n N_VGND_c_957_n 0.0480661f $X=6.162 $Y=1.13 $X2=0
+ $Y2=0
cc_498 N_A_1044_368#_c_661_n N_VGND_c_957_n 0.00197975f $X=6.185 $Y=0.835 $X2=0
+ $Y2=0
cc_499 N_A_1044_368#_M1006_g N_VGND_c_958_n 0.00434272f $X=6.785 $Y=0.74 $X2=0
+ $Y2=0
cc_500 N_A_1044_368#_M1008_g N_VGND_c_958_n 0.00434272f $X=7.215 $Y=0.74 $X2=0
+ $Y2=0
cc_501 N_A_1044_368#_M1013_g N_VGND_c_959_n 0.00434272f $X=7.715 $Y=0.74 $X2=0
+ $Y2=0
cc_502 N_A_1044_368#_M1015_g N_VGND_c_959_n 0.00383152f $X=8.145 $Y=0.74 $X2=0
+ $Y2=0
cc_503 N_A_1044_368#_M1006_g N_VGND_c_964_n 0.00825283f $X=6.785 $Y=0.74 $X2=0
+ $Y2=0
cc_504 N_A_1044_368#_M1008_g N_VGND_c_964_n 0.00820718f $X=7.215 $Y=0.74 $X2=0
+ $Y2=0
cc_505 N_A_1044_368#_M1013_g N_VGND_c_964_n 0.00820942f $X=7.715 $Y=0.74 $X2=0
+ $Y2=0
cc_506 N_A_1044_368#_M1015_g N_VGND_c_964_n 0.0075754f $X=8.145 $Y=0.74 $X2=0
+ $Y2=0
cc_507 N_A_1044_368#_c_659_n N_VGND_c_964_n 0.0198939f $X=6.162 $Y=1.13 $X2=0
+ $Y2=0
cc_508 N_VPWR_c_775_n N_GCLK_c_884_n 0.0316504f $X=6.46 $Y=2.26 $X2=0 $Y2=0
cc_509 N_VPWR_c_776_n N_GCLK_c_884_n 0.0439845f $X=7.46 $Y=2.055 $X2=0 $Y2=0
cc_510 N_VPWR_c_785_n N_GCLK_c_884_n 0.0145938f $X=7.295 $Y=3.33 $X2=0 $Y2=0
cc_511 N_VPWR_c_771_n N_GCLK_c_884_n 0.0120466f $X=8.4 $Y=3.33 $X2=0 $Y2=0
cc_512 N_VPWR_c_776_n N_GCLK_c_885_n 0.018891f $X=7.46 $Y=2.055 $X2=0 $Y2=0
cc_513 N_VPWR_c_776_n N_GCLK_c_886_n 0.0716194f $X=7.46 $Y=2.055 $X2=0 $Y2=0
cc_514 N_VPWR_c_778_n N_GCLK_c_886_n 0.0690922f $X=8.36 $Y=2.035 $X2=0 $Y2=0
cc_515 N_VPWR_c_786_n N_GCLK_c_886_n 0.0110241f $X=8.195 $Y=3.33 $X2=0 $Y2=0
cc_516 N_VPWR_c_771_n N_GCLK_c_886_n 0.00909194f $X=8.4 $Y=3.33 $X2=0 $Y2=0
cc_517 N_VPWR_c_778_n GCLK 0.0242686f $X=8.36 $Y=2.035 $X2=0 $Y2=0
cc_518 N_GCLK_c_877_n N_VGND_c_951_n 0.0266484f $X=7 $Y=0.515 $X2=0 $Y2=0
cc_519 N_GCLK_c_878_n N_VGND_c_951_n 0.0199684f $X=7.765 $Y=1.295 $X2=0 $Y2=0
cc_520 N_GCLK_c_880_n N_VGND_c_951_n 0.0244284f $X=7.93 $Y=0.515 $X2=0 $Y2=0
cc_521 N_GCLK_c_880_n N_VGND_c_953_n 0.0254585f $X=7.93 $Y=0.515 $X2=0 $Y2=0
cc_522 GCLK N_VGND_c_953_n 0.0109035f $X=8.315 $Y=1.58 $X2=0 $Y2=0
cc_523 N_GCLK_c_877_n N_VGND_c_957_n 0.00618339f $X=7 $Y=0.515 $X2=0 $Y2=0
cc_524 N_GCLK_c_877_n N_VGND_c_958_n 0.0144922f $X=7 $Y=0.515 $X2=0 $Y2=0
cc_525 N_GCLK_c_880_n N_VGND_c_959_n 0.0109942f $X=7.93 $Y=0.515 $X2=0 $Y2=0
cc_526 N_GCLK_c_877_n N_VGND_c_964_n 0.0118826f $X=7 $Y=0.515 $X2=0 $Y2=0
cc_527 N_GCLK_c_880_n N_VGND_c_964_n 0.00904371f $X=7.93 $Y=0.515 $X2=0 $Y2=0
