* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hs__dfxbp_1 CLK D VGND VNB VPB VPWR Q Q_N
M1000 a_701_463# a_543_447# VPWR VPB pshort w=840000u l=150000u
+  ad=5.082e+11p pd=2.89e+06u as=1.90825e+12p ps=1.568e+07u
M1001 Q a_1191_120# VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=3.192e+11p pd=2.81e+06u as=0p ps=0u
M1002 a_543_447# a_27_74# a_420_503# VNB nlowvt w=420000u l=150000u
+  ad=1.51375e+11p pd=1.66e+06u as=1.176e+11p ps=1.4e+06u
M1003 a_543_447# a_205_368# a_420_503# VPB pshort w=420000u l=150000u
+  ad=2.15075e+11p pd=2.22e+06u as=2.9275e+11p ps=2.67e+06u
M1004 VGND a_701_463# a_713_102# VNB nlowvt w=420000u l=150000u
+  ad=1.73478e+12p pd=1.365e+07u as=8.82e+10p ps=1.26e+06u
M1005 Q a_1191_120# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1006 Q_N a_1644_94# VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=3.248e+11p pd=2.82e+06u as=0p ps=0u
M1007 a_701_463# a_543_447# VGND VNB nlowvt w=550000u l=150000u
+  ad=2.365e+11p pd=2.26e+06u as=0p ps=0u
M1008 a_420_503# D VGND VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VPWR a_1005_120# a_1191_120# VPB pshort w=1e+06u l=150000u
+  ad=0p pd=0u as=2.9e+11p ps=2.58e+06u
M1010 a_420_503# D VPWR VPB pshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_1005_120# a_27_74# a_701_463# VPB pshort w=840000u l=150000u
+  ad=2.817e+11p pd=2.45e+06u as=0p ps=0u
M1012 a_1005_120# a_205_368# a_701_463# VNB nlowvt w=550000u l=150000u
+  ad=2.593e+11p pd=2.18e+06u as=0p ps=0u
M1013 a_713_102# a_205_368# a_543_447# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 VPWR a_1191_120# a_1158_482# VPB pshort w=420000u l=150000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1015 VGND a_1191_120# a_1143_146# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1016 VPWR a_1191_120# a_1644_94# VPB pshort w=840000u l=150000u
+  ad=0p pd=0u as=2.394e+11p ps=2.25e+06u
M1017 a_205_368# a_27_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=3.252e+11p pd=2.59e+06u as=0p ps=0u
M1018 VGND a_1005_120# a_1191_120# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=1.824e+11p ps=1.85e+06u
M1019 a_1143_146# a_27_74# a_1005_120# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_650_508# a_27_74# a_543_447# VPB pshort w=420000u l=150000u
+  ad=1.134e+11p pd=1.38e+06u as=0p ps=0u
M1021 VPWR CLK a_27_74# VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=3.248e+11p ps=2.82e+06u
M1022 a_205_368# a_27_74# VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=3.192e+11p pd=2.81e+06u as=0p ps=0u
M1023 a_1158_482# a_205_368# a_1005_120# VPB pshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 VGND CLK a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1025 Q_N a_1644_94# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1026 VPWR a_701_463# a_650_508# VPB pshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 VGND a_1191_120# a_1644_94# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=1.824e+11p ps=1.85e+06u
.ends
