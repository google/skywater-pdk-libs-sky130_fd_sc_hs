* File: sky130_fd_sc_hs__sdfstp_4.pex.spice
* Created: Thu Aug 27 21:09:43 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HS__SDFSTP_4%SCE 3 5 7 8 10 13 15 16 18 23 27 31
r78 23 27 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.69
+ $Y=1.645 $X2=0.69 $Y2=1.645
r79 19 31 22.732 $w=3.3e-07 $l=1.3e-07 $layer=POLY_cond $X=1.88 $Y=1.415
+ $X2=2.01 $Y2=1.415
r80 18 21 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=1.88 $Y=1.415 $X2=1.88
+ $Y2=1.495
r81 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.88
+ $Y=1.415 $X2=1.88 $Y2=1.415
r82 16 23 9.23067 $w=1.7e-07 $l=1.72337e-07 $layer=LI1_cond $X=0.855 $Y=1.495
+ $X2=0.72 $Y2=1.58
r83 15 21 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.715 $Y=1.495
+ $X2=1.88 $Y2=1.495
r84 15 16 56.107 $w=1.68e-07 $l=8.6e-07 $layer=LI1_cond $X=1.715 $Y=1.495
+ $X2=0.855 $Y2=1.495
r85 11 31 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.01 $Y=1.25
+ $X2=2.01 $Y2=1.415
r86 11 13 343.553 $w=1.5e-07 $l=6.7e-07 $layer=POLY_cond $X=2.01 $Y=1.25
+ $X2=2.01 $Y2=0.58
r87 8 27 102.927 $w=2.88e-07 $l=7.03562e-07 $layer=POLY_cond $X=0.945 $Y=2.245
+ $X2=0.72 $Y2=1.645
r88 8 10 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=0.945 $Y=2.245
+ $X2=0.945 $Y2=2.64
r89 5 27 102.927 $w=2.88e-07 $l=7.03562e-07 $layer=POLY_cond $X=0.495 $Y=2.245
+ $X2=0.72 $Y2=1.645
r90 5 7 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=0.495 $Y=2.245
+ $X2=0.495 $Y2=2.64
r91 1 27 43.9382 $w=5.76e-07 $l=2.96226e-07 $layer=POLY_cond $X=0.495 $Y=1.48
+ $X2=0.72 $Y2=1.645
r92 1 3 461.489 $w=1.5e-07 $l=9e-07 $layer=POLY_cond $X=0.495 $Y=1.48 $X2=0.495
+ $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_HS__SDFSTP_4%A_27_74# 1 2 9 10 12 15 18 21 25 26 30 33
+ 35 37
c74 30 0 7.33056e-20 $X=1.95 $Y=1.995
c75 21 0 1.69735e-19 $X=1.785 $Y=2.405
r76 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.95
+ $Y=1.995 $X2=1.95 $Y2=1.995
r77 28 30 14.4055 $w=2.58e-07 $l=3.25e-07 $layer=LI1_cond $X=1.915 $Y=2.32
+ $X2=1.915 $Y2=1.995
r78 26 37 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.975 $Y=1.075
+ $X2=0.975 $Y2=0.91
r79 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.975
+ $Y=1.075 $X2=0.975 $Y2=1.075
r80 23 33 0.94211 $w=3.3e-07 $l=1.7e-07 $layer=LI1_cond $X=0.445 $Y=1.075
+ $X2=0.275 $Y2=1.075
r81 23 25 18.5089 $w=3.28e-07 $l=5.3e-07 $layer=LI1_cond $X=0.445 $Y=1.075
+ $X2=0.975 $Y2=1.075
r82 22 35 2.76166 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.355 $Y=2.405
+ $X2=0.23 $Y2=2.405
r83 21 28 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=1.785 $Y=2.405
+ $X2=1.915 $Y2=2.32
r84 21 22 93.2941 $w=1.68e-07 $l=1.43e-06 $layer=LI1_cond $X=1.785 $Y=2.405
+ $X2=0.355 $Y2=2.405
r85 18 35 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.23 $Y=2.32 $X2=0.23
+ $Y2=2.405
r86 17 33 5.66538 $w=2.95e-07 $l=1.86145e-07 $layer=LI1_cond $X=0.23 $Y=1.24
+ $X2=0.275 $Y2=1.075
r87 17 18 49.7855 $w=2.48e-07 $l=1.08e-06 $layer=LI1_cond $X=0.23 $Y=1.24
+ $X2=0.23 $Y2=2.32
r88 13 33 5.66538 $w=2.95e-07 $l=1.65e-07 $layer=LI1_cond $X=0.275 $Y=0.91
+ $X2=0.275 $Y2=1.075
r89 13 15 11.1855 $w=3.38e-07 $l=3.3e-07 $layer=LI1_cond $X=0.275 $Y=0.91
+ $X2=0.275 $Y2=0.58
r90 10 31 52.2586 $w=2.99e-07 $l=2.7157e-07 $layer=POLY_cond $X=1.995 $Y=2.245
+ $X2=1.95 $Y2=1.995
r91 10 12 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=1.995 $Y=2.245
+ $X2=1.995 $Y2=2.64
r92 9 37 106.04 $w=1.5e-07 $l=3.3e-07 $layer=POLY_cond $X=1.035 $Y=0.58
+ $X2=1.035 $Y2=0.91
r93 2 35 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=2.32 $X2=0.27 $Y2=2.465
r94 1 15 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_HS__SDFSTP_4%D 1 3 6 8 12
c36 1 0 4.43302e-20 $X=1.365 $Y=2.245
r37 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.41
+ $Y=1.985 $X2=1.41 $Y2=1.985
r38 8 12 7.33373 $w=3.28e-07 $l=2.1e-07 $layer=LI1_cond $X=1.2 $Y=1.985 $X2=1.41
+ $Y2=1.985
r39 4 11 38.5718 $w=2.96e-07 $l=1.72337e-07 $layer=POLY_cond $X=1.425 $Y=1.82
+ $X2=1.41 $Y2=1.985
r40 4 6 635.83 $w=1.5e-07 $l=1.24e-06 $layer=POLY_cond $X=1.425 $Y=1.82
+ $X2=1.425 $Y2=0.58
r41 1 11 54.0414 $w=2.96e-07 $l=2.81603e-07 $layer=POLY_cond $X=1.365 $Y=2.245
+ $X2=1.41 $Y2=1.985
r42 1 3 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=1.365 $Y=2.245
+ $X2=1.365 $Y2=2.64
.ends

.subckt PM_SKY130_FD_SC_HS__SDFSTP_4%SCD 3 6 7 9 10 11 12 17
c42 10 0 6.61961e-20 $X=2.64 $Y=1.295
c43 7 0 2.43041e-19 $X=2.415 $Y=2.245
r44 21 22 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=2.695
+ $Y=1.945 $X2=2.695 $Y2=1.945
r45 17 19 47.5561 $w=5.35e-07 $l=1.65e-07 $layer=POLY_cond $X=2.592 $Y=1.265
+ $X2=2.592 $Y2=1.1
r46 12 22 3.70428 $w=2.78e-07 $l=9e-08 $layer=LI1_cond $X=2.695 $Y=2.035
+ $X2=2.695 $Y2=1.945
r47 11 22 11.5244 $w=2.78e-07 $l=2.8e-07 $layer=LI1_cond $X=2.695 $Y=1.665
+ $X2=2.695 $Y2=1.945
r48 10 11 16.4635 $w=2.78e-07 $l=4e-07 $layer=LI1_cond $X=2.695 $Y=1.265
+ $X2=2.695 $Y2=1.665
r49 10 17 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=2.695
+ $Y=1.265 $X2=2.695 $Y2=1.265
r50 7 21 55.5708 $w=4.15e-07 $l=3.78286e-07 $layer=POLY_cond $X=2.415 $Y=2.245
+ $X2=2.592 $Y2=1.945
r51 7 9 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=2.415 $Y=2.245
+ $X2=2.415 $Y2=2.64
r52 6 21 11.7419 $w=5.35e-07 $l=1.02e-07 $layer=POLY_cond $X=2.592 $Y=1.843
+ $X2=2.592 $Y2=1.945
r53 5 17 10.2006 $w=5.35e-07 $l=1.02e-07 $layer=POLY_cond $X=2.592 $Y=1.367
+ $X2=2.592 $Y2=1.265
r54 5 6 47.6026 $w=5.35e-07 $l=4.76e-07 $layer=POLY_cond $X=2.592 $Y=1.367
+ $X2=2.592 $Y2=1.843
r55 3 19 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=2.4 $Y=0.58 $X2=2.4
+ $Y2=1.1
.ends

.subckt PM_SKY130_FD_SC_HS__SDFSTP_4%CLK 1 3 4 6 7
c34 4 0 6.61961e-20 $X=3.51 $Y=1.765
r35 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.49
+ $Y=1.385 $X2=3.49 $Y2=1.385
r36 7 11 3.42618 $w=3.68e-07 $l=1.1e-07 $layer=LI1_cond $X=3.6 $Y=1.365 $X2=3.49
+ $Y2=1.365
r37 4 10 77.2841 $w=2.7e-07 $l=3.89872e-07 $layer=POLY_cond $X=3.51 $Y=1.765
+ $X2=3.49 $Y2=1.385
r38 4 6 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.51 $Y=1.765
+ $X2=3.51 $Y2=2.4
r39 1 10 38.9026 $w=2.7e-07 $l=1.88348e-07 $layer=POLY_cond $X=3.44 $Y=1.22
+ $X2=3.49 $Y2=1.385
r40 1 3 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=3.44 $Y=1.22 $X2=3.44
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HS__SDFSTP_4%A_803_74# 1 2 8 9 11 12 16 20 21 22 24 25
+ 27 29 31 32 34 36 37 40 42 43 44 48 54 56 57 60 61 62 64 65 66 67 69 72 76 77
+ 79 80 83 84 89 90 95 99 106 108
c298 99 0 3.98141e-20 $X=10.6 $Y=1.97
c299 79 0 2.67659e-20 $X=5.665 $Y=1.94
c300 66 0 1.23112e-19 $X=7.545 $Y=2.035
c301 32 0 9.10184e-20 $X=10.44 $Y=2.465
c302 31 0 1.98549e-19 $X=10.44 $Y=2.375
c303 21 0 1.22616e-19 $X=9.375 $Y=1.16
r304 105 106 33.0969 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=5.09 $Y=1.565
+ $X2=5.18 $Y2=1.565
r305 99 110 27.9778 $w=3.3e-07 $l=1.6e-07 $layer=POLY_cond $X=10.6 $Y=1.97
+ $X2=10.44 $Y2=1.97
r306 98 99 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.6
+ $Y=1.97 $X2=10.6 $Y2=1.97
r307 95 98 4.36531 $w=3.28e-07 $l=1.25e-07 $layer=LI1_cond $X=10.6 $Y=1.845
+ $X2=10.6 $Y2=1.97
r308 92 93 0.69845 $w=3.28e-07 $l=2e-08 $layer=LI1_cond $X=9.21 $Y=1.845
+ $X2=9.21 $Y2=1.865
r309 90 108 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=9.21 $Y=1.615
+ $X2=9.21 $Y2=1.45
r310 89 92 8.03218 $w=3.28e-07 $l=2.3e-07 $layer=LI1_cond $X=9.21 $Y=1.615
+ $X2=9.21 $Y2=1.845
r311 89 90 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.21
+ $Y=1.615 $X2=9.21 $Y2=1.615
r312 84 86 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=7.81 $Y=1.865
+ $X2=7.81 $Y2=2.035
r313 79 82 8.51388 $w=2.88e-07 $l=1.65e-07 $layer=LI1_cond $X=5.685 $Y=1.94
+ $X2=5.685 $Y2=2.105
r314 79 80 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.665
+ $Y=1.94 $X2=5.665 $Y2=1.94
r315 76 77 8.76268 $w=2.78e-07 $l=1.7e-07 $layer=LI1_cond $X=4.945 $Y=1.095
+ $X2=4.945 $Y2=1.265
r316 72 74 6.9845 $w=3.28e-07 $l=2e-07 $layer=LI1_cond $X=4.235 $Y=2.78
+ $X2=4.235 $Y2=2.98
r317 70 92 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.375 $Y=1.845
+ $X2=9.21 $Y2=1.845
r318 69 95 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.435 $Y=1.845
+ $X2=10.6 $Y2=1.845
r319 69 70 69.1551 $w=1.68e-07 $l=1.06e-06 $layer=LI1_cond $X=10.435 $Y=1.845
+ $X2=9.375 $Y2=1.845
r320 68 84 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.895 $Y=1.865
+ $X2=7.81 $Y2=1.865
r321 67 93 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.045 $Y=1.865
+ $X2=9.21 $Y2=1.865
r322 67 68 75.0267 $w=1.68e-07 $l=1.15e-06 $layer=LI1_cond $X=9.045 $Y=1.865
+ $X2=7.895 $Y2=1.865
r323 65 86 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.725 $Y=2.035
+ $X2=7.81 $Y2=2.035
r324 65 66 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=7.725 $Y=2.035
+ $X2=7.545 $Y2=2.035
r325 63 66 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.46 $Y=2.12
+ $X2=7.545 $Y2=2.035
r326 63 64 50.5615 $w=1.68e-07 $l=7.75e-07 $layer=LI1_cond $X=7.46 $Y=2.12
+ $X2=7.46 $Y2=2.895
r327 61 64 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.375 $Y=2.98
+ $X2=7.46 $Y2=2.895
r328 61 62 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=7.375 $Y=2.98
+ $X2=6.865 $Y2=2.98
r329 60 62 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.78 $Y=2.895
+ $X2=6.865 $Y2=2.98
r330 59 60 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=6.78 $Y=2.46
+ $X2=6.78 $Y2=2.895
r331 58 83 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.83 $Y=2.375
+ $X2=5.745 $Y2=2.375
r332 57 59 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.695 $Y=2.375
+ $X2=6.78 $Y2=2.46
r333 57 58 56.4332 $w=1.68e-07 $l=8.65e-07 $layer=LI1_cond $X=6.695 $Y=2.375
+ $X2=5.83 $Y2=2.375
r334 55 83 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.745 $Y=2.46
+ $X2=5.745 $Y2=2.375
r335 55 56 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=5.745 $Y=2.46
+ $X2=5.745 $Y2=2.895
r336 54 83 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.745 $Y=2.29
+ $X2=5.745 $Y2=2.375
r337 54 82 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=5.745 $Y=2.29
+ $X2=5.745 $Y2=2.105
r338 51 76 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.055 $Y=0.425
+ $X2=5.055 $Y2=1.095
r339 49 105 33.2236 $w=3.3e-07 $l=1.9e-07 $layer=POLY_cond $X=4.9 $Y=1.565
+ $X2=5.09 $Y2=1.565
r340 48 77 12.3476 $w=2.78e-07 $l=3e-07 $layer=LI1_cond $X=4.89 $Y=1.565
+ $X2=4.89 $Y2=1.265
r341 48 49 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.9
+ $Y=1.565 $X2=4.9 $Y2=1.565
r342 45 74 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.4 $Y=2.98
+ $X2=4.235 $Y2=2.98
r343 44 56 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.66 $Y=2.98
+ $X2=5.745 $Y2=2.895
r344 44 45 82.2032 $w=1.68e-07 $l=1.26e-06 $layer=LI1_cond $X=5.66 $Y=2.98
+ $X2=4.4 $Y2=2.98
r345 42 51 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.97 $Y=0.34
+ $X2=5.055 $Y2=0.425
r346 42 43 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=4.97 $Y=0.34
+ $X2=4.24 $Y2=0.34
r347 38 43 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.155 $Y=0.425
+ $X2=4.24 $Y2=0.34
r348 38 40 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=4.155 $Y=0.425
+ $X2=4.155 $Y2=0.515
r349 35 80 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=5.665 $Y=1.73
+ $X2=5.665 $Y2=1.94
r350 35 36 13.5877 $w=2.4e-07 $l=7.5e-08 $layer=POLY_cond $X=5.665 $Y=1.73
+ $X2=5.665 $Y2=1.655
r351 32 34 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=10.44 $Y=2.465
+ $X2=10.44 $Y2=2.75
r352 31 32 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=10.44 $Y=2.375
+ $X2=10.44 $Y2=2.465
r353 30 110 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=10.44 $Y=2.135
+ $X2=10.44 $Y2=1.97
r354 30 31 93.2903 $w=1.8e-07 $l=2.4e-07 $layer=POLY_cond $X=10.44 $Y=2.135
+ $X2=10.44 $Y2=2.375
r355 27 29 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=10.16 $Y=1.085
+ $X2=10.16 $Y2=0.69
r356 26 37 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=9.805 $Y=1.16
+ $X2=9.73 $Y2=1.16
r357 25 27 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=10.085 $Y=1.16
+ $X2=10.16 $Y2=1.085
r358 25 26 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=10.085 $Y=1.16
+ $X2=9.805 $Y2=1.16
r359 22 37 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=9.73 $Y=1.085
+ $X2=9.73 $Y2=1.16
r360 22 24 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=9.73 $Y=1.085
+ $X2=9.73 $Y2=0.69
r361 20 37 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=9.655 $Y=1.16
+ $X2=9.73 $Y2=1.16
r362 20 21 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=9.655 $Y=1.16
+ $X2=9.375 $Y2=1.16
r363 18 21 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=9.3 $Y=1.235
+ $X2=9.375 $Y2=1.16
r364 18 108 110.245 $w=1.5e-07 $l=2.15e-07 $layer=POLY_cond $X=9.3 $Y=1.235
+ $X2=9.3 $Y2=1.45
r365 14 36 13.5877 $w=2.4e-07 $l=8.66025e-08 $layer=POLY_cond $X=5.69 $Y=1.58
+ $X2=5.665 $Y2=1.655
r366 14 16 494.819 $w=1.5e-07 $l=9.65e-07 $layer=POLY_cond $X=5.69 $Y=1.58
+ $X2=5.69 $Y2=0.615
r367 12 36 12.1617 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.5 $Y=1.655
+ $X2=5.665 $Y2=1.655
r368 12 106 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=5.5 $Y=1.655
+ $X2=5.18 $Y2=1.655
r369 9 11 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=5.09 $Y=2.21 $X2=5.09
+ $Y2=2.495
r370 8 9 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=5.09 $Y=2.12 $X2=5.09
+ $Y2=2.21
r371 7 105 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=5.09 $Y=1.73
+ $X2=5.09 $Y2=1.565
r372 7 8 151.597 $w=1.8e-07 $l=3.9e-07 $layer=POLY_cond $X=5.09 $Y=1.73 $X2=5.09
+ $Y2=2.12
r373 2 72 600 $w=1.7e-07 $l=1.03518e-06 $layer=licon1_PDIFF $count=1 $X=4.035
+ $Y=1.84 $X2=4.235 $Y2=2.78
r374 1 40 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=4.015
+ $Y=0.37 $X2=4.155 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__SDFSTP_4%A_1201_55# 1 2 9 10 12 14 15 17 21 25 27 31
+ 34 40
c86 14 0 2.67659e-20 $X=6.26 $Y=1.78
r87 34 37 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=6.205 $Y=1.945
+ $X2=6.205 $Y2=2.035
r88 34 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.205
+ $Y=1.945 $X2=6.205 $Y2=1.945
r89 31 41 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.17 $Y=1.1
+ $X2=6.17 $Y2=1.265
r90 31 40 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.17 $Y=1.1
+ $X2=6.17 $Y2=0.935
r91 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.17
+ $Y=1.1 $X2=6.17 $Y2=1.1
r92 27 30 8.55602 $w=3.28e-07 $l=2.45e-07 $layer=LI1_cond $X=6.17 $Y=0.855
+ $X2=6.17 $Y2=1.1
r93 23 25 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=7.12 $Y=2.12
+ $X2=7.12 $Y2=2.495
r94 19 21 6.63528 $w=3.28e-07 $l=1.9e-07 $layer=LI1_cond $X=6.935 $Y=0.77
+ $X2=6.935 $Y2=0.58
r95 18 37 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.37 $Y=2.035
+ $X2=6.205 $Y2=2.035
r96 17 23 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.035 $Y=2.035
+ $X2=7.12 $Y2=2.12
r97 17 18 43.385 $w=1.68e-07 $l=6.65e-07 $layer=LI1_cond $X=7.035 $Y=2.035
+ $X2=6.37 $Y2=2.035
r98 16 27 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.335 $Y=0.855
+ $X2=6.17 $Y2=0.855
r99 15 19 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=6.77 $Y=0.855
+ $X2=6.935 $Y2=0.77
r100 15 16 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=6.77 $Y=0.855
+ $X2=6.335 $Y2=0.855
r101 14 35 38.578 $w=2.95e-07 $l=1.90526e-07 $layer=POLY_cond $X=6.26 $Y=1.78
+ $X2=6.205 $Y2=1.945
r102 14 41 264.074 $w=1.5e-07 $l=5.15e-07 $layer=POLY_cond $X=6.26 $Y=1.78
+ $X2=6.26 $Y2=1.265
r103 10 35 54.9169 $w=2.95e-07 $l=3.00167e-07 $layer=POLY_cond $X=6.13 $Y=2.21
+ $X2=6.205 $Y2=1.945
r104 10 12 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=6.13 $Y=2.21
+ $X2=6.13 $Y2=2.495
r105 9 40 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=6.08 $Y=0.615
+ $X2=6.08 $Y2=0.935
r106 2 25 600 $w=1.7e-07 $l=2.86182e-07 $layer=licon1_PDIFF $count=1 $X=6.94
+ $Y=2.285 $X2=7.12 $Y2=2.495
r107 1 21 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=6.79
+ $Y=0.37 $X2=6.935 $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_HS__SDFSTP_4%A_1017_81# 1 2 8 9 11 12 14 16 17 19 20 22
+ 24 25 27 28 30 34 35 38 40 44 46 48 50 51 52 56 59 69
c174 25 0 7.58781e-20 $X=8.475 $Y=1.79
c175 8 0 1.23112e-19 $X=6.865 $Y=2.12
r176 68 69 27.3299 $w=2.91e-07 $l=1.65e-07 $layer=POLY_cond $X=8.31 $Y=1.267
+ $X2=8.475 $Y2=1.267
r177 63 68 34.7835 $w=2.91e-07 $l=2.1e-07 $layer=POLY_cond $X=8.1 $Y=1.267
+ $X2=8.31 $Y2=1.267
r178 63 66 12.4227 $w=2.91e-07 $l=7.5e-08 $layer=POLY_cond $X=8.1 $Y=1.267
+ $X2=8.025 $Y2=1.267
r179 62 63 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.1
+ $Y=1.285 $X2=8.1 $Y2=1.285
r180 59 62 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=8.1 $Y=1.195 $X2=8.1
+ $Y2=1.285
r181 55 57 8.55602 $w=3.28e-07 $l=2.45e-07 $layer=LI1_cond $X=6.79 $Y=1.275
+ $X2=6.79 $Y2=1.52
r182 55 56 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.79
+ $Y=1.275 $X2=6.79 $Y2=1.275
r183 52 55 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=6.79 $Y=1.195 $X2=6.79
+ $Y2=1.275
r184 49 52 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.955 $Y=1.195
+ $X2=6.79 $Y2=1.195
r185 48 59 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.935 $Y=1.195
+ $X2=8.1 $Y2=1.195
r186 48 49 63.9358 $w=1.68e-07 $l=9.8e-07 $layer=LI1_cond $X=7.935 $Y=1.195
+ $X2=6.955 $Y2=1.195
r187 47 50 2.76166 $w=1.7e-07 $l=2.2e-07 $layer=LI1_cond $X=5.64 $Y=1.52
+ $X2=5.42 $Y2=1.52
r188 46 57 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.625 $Y=1.52
+ $X2=6.79 $Y2=1.52
r189 46 47 64.262 $w=1.68e-07 $l=9.85e-07 $layer=LI1_cond $X=6.625 $Y=1.52
+ $X2=5.64 $Y2=1.52
r190 42 50 3.70735 $w=2.5e-07 $l=1.09087e-07 $layer=LI1_cond $X=5.475 $Y=1.435
+ $X2=5.42 $Y2=1.52
r191 42 44 28.6365 $w=3.28e-07 $l=8.2e-07 $layer=LI1_cond $X=5.475 $Y=1.435
+ $X2=5.475 $Y2=0.615
r192 38 51 7.52792 $w=2.78e-07 $l=1.4e-07 $layer=LI1_cond $X=5.34 $Y=2.415
+ $X2=5.34 $Y2=2.275
r193 38 40 3.49849 $w=2.78e-07 $l=8.5e-08 $layer=LI1_cond $X=5.34 $Y=2.415
+ $X2=5.34 $Y2=2.5
r194 36 50 3.70735 $w=2.5e-07 $l=1.72337e-07 $layer=LI1_cond $X=5.285 $Y=1.605
+ $X2=5.42 $Y2=1.52
r195 36 51 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.285 $Y=1.605
+ $X2=5.285 $Y2=2.275
r196 34 56 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=6.79 $Y=1.615
+ $X2=6.79 $Y2=1.275
r197 34 35 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.79 $Y=1.615
+ $X2=6.79 $Y2=1.78
r198 28 69 43.8935 $w=2.91e-07 $l=3.44173e-07 $layer=POLY_cond $X=8.74 $Y=1.085
+ $X2=8.475 $Y2=1.267
r199 28 30 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=8.74 $Y=1.085
+ $X2=8.74 $Y2=0.69
r200 25 27 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=8.475 $Y=1.79
+ $X2=8.475 $Y2=2.285
r201 24 25 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=8.475 $Y=1.7
+ $X2=8.475 $Y2=1.79
r202 23 69 14.0159 $w=1.8e-07 $l=1.83e-07 $layer=POLY_cond $X=8.475 $Y=1.45
+ $X2=8.475 $Y2=1.267
r203 23 24 97.1774 $w=1.8e-07 $l=2.5e-07 $layer=POLY_cond $X=8.475 $Y=1.45
+ $X2=8.475 $Y2=1.7
r204 20 68 18.2534 $w=1.5e-07 $l=1.82e-07 $layer=POLY_cond $X=8.31 $Y=1.085
+ $X2=8.31 $Y2=1.267
r205 20 22 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=8.31 $Y=1.085
+ $X2=8.31 $Y2=0.69
r206 17 19 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=8.025 $Y=1.79
+ $X2=8.025 $Y2=2.285
r207 16 17 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=8.025 $Y=1.7
+ $X2=8.025 $Y2=1.79
r208 15 66 14.0159 $w=1.8e-07 $l=1.83e-07 $layer=POLY_cond $X=8.025 $Y=1.45
+ $X2=8.025 $Y2=1.267
r209 15 16 97.1774 $w=1.8e-07 $l=2.5e-07 $layer=POLY_cond $X=8.025 $Y=1.45
+ $X2=8.025 $Y2=1.7
r210 12 56 79.2329 $w=2.19e-07 $l=5.61872e-07 $layer=POLY_cond $X=7.15 $Y=0.865
+ $X2=6.79 $Y2=1.275
r211 12 14 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=7.15 $Y=0.865
+ $X2=7.15 $Y2=0.58
r212 9 11 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=6.865 $Y=2.21
+ $X2=6.865 $Y2=2.495
r213 8 9 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=6.865 $Y=2.12 $X2=6.865
+ $Y2=2.21
r214 8 35 132.161 $w=1.8e-07 $l=3.4e-07 $layer=POLY_cond $X=6.865 $Y=2.12
+ $X2=6.865 $Y2=1.78
r215 2 40 600 $w=1.7e-07 $l=2.80134e-07 $layer=licon1_PDIFF $count=1 $X=5.165
+ $Y=2.285 $X2=5.315 $Y2=2.5
r216 1 44 182 $w=1.7e-07 $l=4.83735e-07 $layer=licon1_NDIFF $count=1 $X=5.085
+ $Y=0.405 $X2=5.475 $Y2=0.615
.ends

.subckt PM_SKY130_FD_SC_HS__SDFSTP_4%SET_B 2 3 5 8 11 13 14 16 19 21 22 23 28 34
+ 35 38 39
c143 28 0 1.12416e-19 $X=11.76 $Y=1.665
c144 22 0 6.13349e-20 $X=11.615 $Y=1.665
c145 11 0 7.95967e-20 $X=11.612 $Y=1.953
c146 3 0 1.49656e-19 $X=7.345 $Y=2.21
r147 38 40 45.1558 $w=3.75e-07 $l=1.65e-07 $layer=POLY_cond $X=11.612 $Y=1.635
+ $X2=11.612 $Y2=1.47
r148 38 39 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=11.635
+ $Y=1.635 $X2=11.635 $Y2=1.635
r149 33 35 31.475 $w=3.3e-07 $l=1.8e-07 $layer=POLY_cond $X=7.36 $Y=1.615
+ $X2=7.54 $Y2=1.615
r150 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.36
+ $Y=1.615 $X2=7.36 $Y2=1.615
r151 30 33 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=7.345 $Y=1.615
+ $X2=7.36 $Y2=1.615
r152 28 39 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.76 $Y=1.665
+ $X2=11.76 $Y2=1.665
r153 25 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=1.665
+ $X2=7.44 $Y2=1.665
r154 23 25 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=7.585 $Y=1.665
+ $X2=7.44 $Y2=1.665
r155 22 28 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=11.615 $Y=1.665
+ $X2=11.76 $Y2=1.665
r156 22 23 4.98761 $w=1.4e-07 $l=4.03e-06 $layer=MET1_cond $X=11.615 $Y=1.665
+ $X2=7.585 $Y2=1.665
r157 19 40 456.362 $w=1.5e-07 $l=8.9e-07 $layer=POLY_cond $X=11.6 $Y=0.58
+ $X2=11.6 $Y2=1.47
r158 14 16 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=11.515 $Y=2.465
+ $X2=11.515 $Y2=2.75
r159 13 14 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=11.515 $Y=2.375
+ $X2=11.515 $Y2=2.465
r160 13 21 91.3468 $w=1.8e-07 $l=2.35e-07 $layer=POLY_cond $X=11.515 $Y=2.375
+ $X2=11.515 $Y2=2.14
r161 11 21 42.8297 $w=3.75e-07 $l=1.87e-07 $layer=POLY_cond $X=11.612 $Y=1.953
+ $X2=11.612 $Y2=2.14
r162 10 38 3.26277 $w=3.75e-07 $l=2.2e-08 $layer=POLY_cond $X=11.612 $Y=1.657
+ $X2=11.612 $Y2=1.635
r163 10 11 43.8991 $w=3.75e-07 $l=2.96e-07 $layer=POLY_cond $X=11.612 $Y=1.657
+ $X2=11.612 $Y2=1.953
r164 6 35 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.54 $Y=1.45
+ $X2=7.54 $Y2=1.615
r165 6 8 446.106 $w=1.5e-07 $l=8.7e-07 $layer=POLY_cond $X=7.54 $Y=1.45 $X2=7.54
+ $Y2=0.58
r166 3 5 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=7.345 $Y=2.21
+ $X2=7.345 $Y2=2.495
r167 2 3 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=7.345 $Y=2.12 $X2=7.345
+ $Y2=2.21
r168 1 30 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=7.345 $Y=1.78
+ $X2=7.345 $Y2=1.615
r169 1 2 132.161 $w=1.8e-07 $l=3.4e-07 $layer=POLY_cond $X=7.345 $Y=1.78
+ $X2=7.345 $Y2=2.12
.ends

.subckt PM_SKY130_FD_SC_HS__SDFSTP_4%A_616_74# 1 2 9 11 13 15 16 17 19 20 21 22
+ 23 26 28 30 31 33 35 36 39 40 43 44 45 48 52 54 56 59 62 63 64 69 72
c200 19 0 1.33164e-19 $X=4.53 $Y=3.075
c201 11 0 1.2825e-19 $X=3.96 $Y=1.765
r202 73 74 2.73088 $w=3.53e-07 $l=2e-08 $layer=POLY_cond $X=3.94 $Y=1.557
+ $X2=3.96 $Y2=1.557
r203 70 74 12.289 $w=3.53e-07 $l=9e-08 $layer=POLY_cond $X=4.05 $Y=1.557
+ $X2=3.96 $Y2=1.557
r204 69 70 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.05
+ $Y=1.515 $X2=4.05 $Y2=1.515
r205 67 69 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=4.05 $Y=1.82
+ $X2=4.05 $Y2=1.515
r206 64 66 5.07075 $w=2.48e-07 $l=1.1e-07 $layer=LI1_cond $X=3.175 $Y=1.945
+ $X2=3.285 $Y2=1.945
r207 63 67 6.98653 $w=2.5e-07 $l=2.18746e-07 $layer=LI1_cond $X=3.885 $Y=1.945
+ $X2=4.05 $Y2=1.82
r208 63 66 27.6586 $w=2.48e-07 $l=6e-07 $layer=LI1_cond $X=3.885 $Y=1.945
+ $X2=3.285 $Y2=1.945
r209 62 64 7.14316 $w=2.5e-07 $l=1.62019e-07 $layer=LI1_cond $X=3.09 $Y=1.82
+ $X2=3.175 $Y2=1.945
r210 62 72 52.8449 $w=1.68e-07 $l=8.1e-07 $layer=LI1_cond $X=3.09 $Y=1.82
+ $X2=3.09 $Y2=1.01
r211 57 72 9.39714 $w=3.83e-07 $l=1.92e-07 $layer=LI1_cond $X=3.197 $Y=0.818
+ $X2=3.197 $Y2=1.01
r212 57 59 9.06988 $w=3.83e-07 $l=3.03e-07 $layer=LI1_cond $X=3.197 $Y=0.818
+ $X2=3.197 $Y2=0.515
r213 50 52 41.0213 $w=1.5e-07 $l=8e-08 $layer=POLY_cond $X=4.45 $Y=2.045
+ $X2=4.53 $Y2=2.045
r214 46 48 443.543 $w=1.5e-07 $l=8.65e-07 $layer=POLY_cond $X=10.67 $Y=1.445
+ $X2=10.67 $Y2=0.58
r215 44 46 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=10.595 $Y=1.52
+ $X2=10.67 $Y2=1.445
r216 44 45 292.277 $w=1.5e-07 $l=5.7e-07 $layer=POLY_cond $X=10.595 $Y=1.52
+ $X2=10.025 $Y2=1.52
r217 41 43 253.819 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=9.935 $Y=3.035
+ $X2=9.935 $Y2=2.54
r218 40 43 253.819 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=9.935 $Y=2.045
+ $X2=9.935 $Y2=2.54
r219 39 40 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=9.935 $Y=1.955
+ $X2=9.935 $Y2=2.045
r220 38 45 22.7899 $w=1.97e-07 $l=2.05122e-07 $layer=POLY_cond $X=9.935 $Y=1.685
+ $X2=10.025 $Y2=1.52
r221 38 39 104.952 $w=1.8e-07 $l=2.7e-07 $layer=POLY_cond $X=9.935 $Y=1.685
+ $X2=9.935 $Y2=1.955
r222 37 56 20.4101 $w=1.5e-07 $l=9.94987e-08 $layer=POLY_cond $X=9.575 $Y=3.15
+ $X2=9.485 $Y2=3.13
r223 36 41 26.9307 $w=1.5e-07 $l=1.53542e-07 $layer=POLY_cond $X=9.845 $Y=3.15
+ $X2=9.935 $Y2=3.035
r224 36 37 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=9.845 $Y=3.15
+ $X2=9.575 $Y2=3.15
r225 33 56 5.30422 $w=1.5e-07 $l=9.5e-08 $layer=POLY_cond $X=9.485 $Y=3.035
+ $X2=9.485 $Y2=3.13
r226 33 35 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=9.485 $Y=3.035
+ $X2=9.485 $Y2=2.54
r227 32 54 7.1379 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=5.715 $Y=3.15
+ $X2=5.625 $Y2=3.15
r228 31 56 20.4101 $w=1.5e-07 $l=9.94987e-08 $layer=POLY_cond $X=9.395 $Y=3.15
+ $X2=9.485 $Y2=3.13
r229 31 32 1886.98 $w=1.5e-07 $l=3.68e-06 $layer=POLY_cond $X=9.395 $Y=3.15
+ $X2=5.715 $Y2=3.15
r230 28 54 72.1175 $w=1.8e-07 $l=1.8e-07 $layer=POLY_cond $X=5.625 $Y=2.97
+ $X2=5.625 $Y2=3.15
r231 28 30 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=5.625 $Y=2.97
+ $X2=5.625 $Y2=2.685
r232 24 26 217.926 $w=1.5e-07 $l=4.25e-07 $layer=POLY_cond $X=5.01 $Y=1.04
+ $X2=5.01 $Y2=0.615
r233 22 54 7.1379 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=5.535 $Y=3.15
+ $X2=5.625 $Y2=3.15
r234 22 23 476.872 $w=1.5e-07 $l=9.3e-07 $layer=POLY_cond $X=5.535 $Y=3.15
+ $X2=4.605 $Y2=3.15
r235 20 24 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.935 $Y=1.115
+ $X2=5.01 $Y2=1.04
r236 20 21 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=4.935 $Y=1.115
+ $X2=4.525 $Y2=1.115
r237 19 23 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.53 $Y=3.075
+ $X2=4.605 $Y2=3.15
r238 18 52 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.53 $Y=2.12
+ $X2=4.53 $Y2=2.045
r239 18 19 489.691 $w=1.5e-07 $l=9.55e-07 $layer=POLY_cond $X=4.53 $Y=2.12
+ $X2=4.53 $Y2=3.075
r240 17 50 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.45 $Y=1.97
+ $X2=4.45 $Y2=2.045
r241 16 70 54.6176 $w=3.53e-07 $l=4e-07 $layer=POLY_cond $X=4.45 $Y=1.557
+ $X2=4.05 $Y2=1.557
r242 16 17 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=4.45 $Y=1.68
+ $X2=4.45 $Y2=1.97
r243 15 16 22.8335 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.45 $Y=1.35
+ $X2=4.45 $Y2=1.557
r244 14 21 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.45 $Y=1.19
+ $X2=4.525 $Y2=1.115
r245 14 15 82.0426 $w=1.5e-07 $l=1.6e-07 $layer=POLY_cond $X=4.45 $Y=1.19
+ $X2=4.45 $Y2=1.35
r246 11 74 22.8335 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=3.96 $Y=1.765
+ $X2=3.96 $Y2=1.557
r247 11 13 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.96 $Y=1.765
+ $X2=3.96 $Y2=2.4
r248 7 73 22.8335 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.94 $Y=1.35
+ $X2=3.94 $Y2=1.557
r249 7 9 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=3.94 $Y=1.35 $X2=3.94
+ $Y2=0.74
r250 2 66 600 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=3.14
+ $Y=1.84 $X2=3.285 $Y2=1.985
r251 1 59 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=3.08
+ $Y=0.37 $X2=3.225 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__SDFSTP_4%A_2191_180# 1 2 8 11 12 14 15 19 22 24 25
+ 29 34 36 39 42
c106 34 0 1.11167e-19 $X=12.465 $Y=2.815
c107 29 0 1.71901e-19 $X=11.12 $Y=1.065
c108 24 0 4.1327e-20 $X=12.625 $Y=2.18
r109 37 39 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=12.465 $Y=2.265
+ $X2=12.625 $Y2=2.265
r110 32 34 5.76222 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=12.3 $Y=2.815
+ $X2=12.465 $Y2=2.815
r111 29 43 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=11.12 $Y=1.065
+ $X2=11.12 $Y2=1.23
r112 29 42 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=11.12 $Y=1.065
+ $X2=11.12 $Y2=0.9
r113 28 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=11.12
+ $Y=1.065 $X2=11.12 $Y2=1.065
r114 25 28 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=11.12 $Y=0.985
+ $X2=11.12 $Y2=1.065
r115 24 39 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=12.625 $Y=2.18
+ $X2=12.625 $Y2=2.265
r116 23 36 3.351 $w=2.8e-07 $l=1.46458e-07 $layer=LI1_cond $X=12.625 $Y=1.07
+ $X2=12.515 $Y2=0.985
r117 23 24 72.4171 $w=1.68e-07 $l=1.11e-06 $layer=LI1_cond $X=12.625 $Y=1.07
+ $X2=12.625 $Y2=2.18
r118 22 34 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12.465 $Y=2.65
+ $X2=12.465 $Y2=2.815
r119 21 37 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=12.465 $Y=2.35
+ $X2=12.465 $Y2=2.265
r120 21 22 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=12.465 $Y=2.35
+ $X2=12.465 $Y2=2.65
r121 17 36 3.351 $w=2.8e-07 $l=8.5e-08 $layer=LI1_cond $X=12.515 $Y=0.9
+ $X2=12.515 $Y2=0.985
r122 17 19 9.45594 $w=3.88e-07 $l=3.2e-07 $layer=LI1_cond $X=12.515 $Y=0.9
+ $X2=12.515 $Y2=0.58
r123 16 25 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.285 $Y=0.985
+ $X2=11.12 $Y2=0.985
r124 15 36 3.18746 $w=1.7e-07 $l=1.95e-07 $layer=LI1_cond $X=12.32 $Y=0.985
+ $X2=12.515 $Y2=0.985
r125 15 16 67.5241 $w=1.68e-07 $l=1.035e-06 $layer=LI1_cond $X=12.32 $Y=0.985
+ $X2=11.285 $Y2=0.985
r126 12 14 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=11.065 $Y=2.465
+ $X2=11.065 $Y2=2.75
r127 11 42 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=11.06 $Y=0.58
+ $X2=11.06 $Y2=0.9
r128 8 12 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=11.065 $Y=2.375
+ $X2=11.065 $Y2=2.465
r129 8 43 445.073 $w=1.8e-07 $l=1.145e-06 $layer=POLY_cond $X=11.065 $Y=2.375
+ $X2=11.065 $Y2=1.23
r130 2 32 600 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_PDIFF $count=1 $X=12.155
+ $Y=2.54 $X2=12.3 $Y2=2.815
r131 1 19 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=12.345
+ $Y=0.37 $X2=12.485 $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_HS__SDFSTP_4%A_1823_524# 1 2 3 4 5 18 21 22 24 25 27 29
+ 32 34 36 38 42 44 46 47 51 55 56 57 58 59 61 62 66 70 71 74 76 80 82 84
c216 58 0 2.62796e-19 $X=10.935 $Y=1.485
c217 38 0 4.1327e-20 $X=13.26 $Y=1.967
c218 27 0 1.11167e-19 $X=13.03 $Y=2.045
r219 87 88 34.5038 $w=5.75e-07 $l=7.5e-08 $layer=POLY_cond $X=12.327 $Y=1.965
+ $X2=12.327 $Y2=2.04
r220 76 78 7.28509 $w=2.78e-07 $l=1.77e-07 $layer=LI1_cond $X=9.235 $Y=2.79
+ $X2=9.235 $Y2=2.967
r221 74 82 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=12.125 $Y=2.31
+ $X2=12.125 $Y2=2.395
r222 74 84 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=12.125 $Y=2.31
+ $X2=12.125 $Y2=2.01
r223 71 87 42.8024 $w=5.75e-07 $l=4.6e-07 $layer=POLY_cond $X=12.327 $Y=1.505
+ $X2=12.327 $Y2=1.965
r224 71 86 48.7424 $w=5.75e-07 $l=1.65e-07 $layer=POLY_cond $X=12.327 $Y=1.505
+ $X2=12.327 $Y2=1.34
r225 70 71 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=12.205
+ $Y=1.505 $X2=12.205 $Y2=1.505
r226 68 84 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=12.205 $Y=1.845
+ $X2=12.205 $Y2=2.01
r227 68 70 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=12.205 $Y=1.845
+ $X2=12.205 $Y2=1.505
r228 64 82 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=11.74 $Y=2.395
+ $X2=12.125 $Y2=2.395
r229 64 66 9.42908 $w=3.28e-07 $l=2.7e-07 $layer=LI1_cond $X=11.74 $Y=2.48
+ $X2=11.74 $Y2=2.75
r230 63 80 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=11.105 $Y=2.395
+ $X2=11.02 $Y2=2.395
r231 62 64 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=11.575 $Y=2.395
+ $X2=11.74 $Y2=2.395
r232 62 63 30.6631 $w=1.68e-07 $l=4.7e-07 $layer=LI1_cond $X=11.575 $Y=2.395
+ $X2=11.105 $Y2=2.395
r233 61 80 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=11.02 $Y=2.31
+ $X2=11.02 $Y2=2.395
r234 60 61 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=11.02 $Y=1.57
+ $X2=11.02 $Y2=2.31
r235 58 60 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=10.935 $Y=1.485
+ $X2=11.02 $Y2=1.57
r236 58 59 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=10.935 $Y=1.485
+ $X2=10.54 $Y2=1.485
r237 56 80 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.935 $Y=2.395
+ $X2=11.02 $Y2=2.395
r238 56 57 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=10.935 $Y=2.395
+ $X2=10.375 $Y2=2.395
r239 53 59 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=10.375 $Y=1.4
+ $X2=10.54 $Y2=1.485
r240 53 55 30.9064 $w=3.28e-07 $l=8.85e-07 $layer=LI1_cond $X=10.375 $Y=1.4
+ $X2=10.375 $Y2=0.515
r241 52 55 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=10.375 $Y=0.425
+ $X2=10.375 $Y2=0.515
r242 49 51 4.01609 $w=3.28e-07 $l=1.15e-07 $layer=LI1_cond $X=10.21 $Y=2.86
+ $X2=10.21 $Y2=2.745
r243 48 57 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=10.21 $Y=2.48
+ $X2=10.375 $Y2=2.395
r244 48 51 9.25447 $w=3.28e-07 $l=2.65e-07 $layer=LI1_cond $X=10.21 $Y=2.48
+ $X2=10.21 $Y2=2.745
r245 46 52 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=10.21 $Y=0.34
+ $X2=10.375 $Y2=0.425
r246 46 47 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=10.21 $Y=0.34
+ $X2=9.68 $Y2=0.34
r247 45 78 2.30834 $w=2.15e-07 $l=1.4e-07 $layer=LI1_cond $X=9.375 $Y=2.967
+ $X2=9.235 $Y2=2.967
r248 44 49 7.21882 $w=2.15e-07 $l=2.11849e-07 $layer=LI1_cond $X=10.045 $Y=2.967
+ $X2=10.21 $Y2=2.86
r249 44 45 35.9133 $w=2.13e-07 $l=6.7e-07 $layer=LI1_cond $X=10.045 $Y=2.967
+ $X2=9.375 $Y2=2.967
r250 40 47 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=9.515 $Y=0.425
+ $X2=9.68 $Y2=0.34
r251 40 42 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=9.515 $Y=0.425
+ $X2=9.515 $Y2=0.515
r252 38 39 69.7632 $w=1.52e-07 $l=2.2e-07 $layer=POLY_cond $X=13.26 $Y=1.967
+ $X2=13.48 $Y2=1.967
r253 37 38 72.9342 $w=1.52e-07 $l=2.3e-07 $layer=POLY_cond $X=13.03 $Y=1.967
+ $X2=13.26 $Y2=1.967
r254 34 39 3.14937 $w=1.5e-07 $l=7.8e-08 $layer=POLY_cond $X=13.48 $Y=2.045
+ $X2=13.48 $Y2=1.967
r255 34 36 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=13.48 $Y=2.045
+ $X2=13.48 $Y2=2.54
r256 30 38 3.14937 $w=1.5e-07 $l=7.7e-08 $layer=POLY_cond $X=13.26 $Y=1.89
+ $X2=13.26 $Y2=1.967
r257 30 32 589.681 $w=1.5e-07 $l=1.15e-06 $layer=POLY_cond $X=13.26 $Y=1.89
+ $X2=13.26 $Y2=0.74
r258 27 37 3.14937 $w=1.5e-07 $l=7.8e-08 $layer=POLY_cond $X=13.03 $Y=2.045
+ $X2=13.03 $Y2=1.967
r259 27 29 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=13.03 $Y=2.045
+ $X2=13.03 $Y2=2.54
r260 26 87 34.9747 $w=1.5e-07 $l=2.88e-07 $layer=POLY_cond $X=12.615 $Y=1.965
+ $X2=12.327 $Y2=1.965
r261 25 37 28.5395 $w=1.52e-07 $l=9.09945e-08 $layer=POLY_cond $X=12.94 $Y=1.965
+ $X2=13.03 $Y2=1.967
r262 25 26 166.649 $w=1.5e-07 $l=3.25e-07 $layer=POLY_cond $X=12.94 $Y=1.965
+ $X2=12.615 $Y2=1.965
r263 22 24 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=12.525 $Y=2.465
+ $X2=12.525 $Y2=2.75
r264 21 22 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=12.525 $Y=2.375
+ $X2=12.525 $Y2=2.465
r265 21 88 130.218 $w=1.8e-07 $l=3.35e-07 $layer=POLY_cond $X=12.525 $Y=2.375
+ $X2=12.525 $Y2=2.04
r266 18 86 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=12.27 $Y=0.58
+ $X2=12.27 $Y2=1.34
r267 5 66 600 $w=1.7e-07 $l=2.74955e-07 $layer=licon1_PDIFF $count=1 $X=11.59
+ $Y=2.54 $X2=11.74 $Y2=2.75
r268 4 51 600 $w=1.7e-07 $l=7.1807e-07 $layer=licon1_PDIFF $count=1 $X=10.01
+ $Y=2.12 $X2=10.21 $Y2=2.745
r269 3 76 600 $w=1.7e-07 $l=2.31409e-07 $layer=licon1_PDIFF $count=1 $X=9.115
+ $Y=2.62 $X2=9.26 $Y2=2.79
r270 2 55 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=10.235
+ $Y=0.37 $X2=10.375 $Y2=0.515
r271 1 42 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=9.37
+ $Y=0.37 $X2=9.515 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__SDFSTP_4%A_2580_74# 1 2 9 11 13 16 18 20 23 25 27 28
+ 29 32 35 36 38 39 42 46 53 56
c121 39 0 1.69241e-19 $X=15.312 $Y=1.395
c122 32 0 2.40437e-20 $X=15.275 $Y=0.74
c123 23 0 2.92295e-20 $X=14.845 $Y=0.74
r124 63 64 5.10053 $w=3.78e-07 $l=4e-08 $layer=POLY_cond $X=14.845 $Y=1.542
+ $X2=14.885 $Y2=1.542
r125 60 61 11.4762 $w=3.78e-07 $l=9e-08 $layer=POLY_cond $X=14.345 $Y=1.542
+ $X2=14.435 $Y2=1.542
r126 59 60 45.9048 $w=3.78e-07 $l=3.6e-07 $layer=POLY_cond $X=13.985 $Y=1.542
+ $X2=14.345 $Y2=1.542
r127 54 63 40.1667 $w=3.78e-07 $l=3.15e-07 $layer=POLY_cond $X=14.53 $Y=1.542
+ $X2=14.845 $Y2=1.542
r128 54 61 12.1138 $w=3.78e-07 $l=9.5e-08 $layer=POLY_cond $X=14.53 $Y=1.542
+ $X2=14.435 $Y2=1.542
r129 53 54 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=14.53
+ $Y=1.485 $X2=14.53 $Y2=1.485
r130 51 59 17.2143 $w=3.78e-07 $l=1.35e-07 $layer=POLY_cond $X=13.85 $Y=1.542
+ $X2=13.985 $Y2=1.542
r131 51 57 11.4762 $w=3.78e-07 $l=9e-08 $layer=POLY_cond $X=13.85 $Y=1.542
+ $X2=13.76 $Y2=1.542
r132 50 53 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=13.85 $Y=1.485
+ $X2=14.53 $Y2=1.485
r133 50 51 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=13.85
+ $Y=1.485 $X2=13.85 $Y2=1.485
r134 48 56 0.364692 $w=3.3e-07 $l=5.3619e-07 $layer=LI1_cond $X=13.34 $Y=1.485
+ $X2=12.88 $Y2=1.32
r135 48 50 17.8105 $w=3.28e-07 $l=5.1e-07 $layer=LI1_cond $X=13.34 $Y=1.485
+ $X2=13.85 $Y2=1.485
r136 44 56 6.46576 $w=2.5e-07 $l=5.14174e-07 $layer=LI1_cond $X=13.255 $Y=1.65
+ $X2=12.88 $Y2=1.32
r137 44 46 40.123 $w=1.68e-07 $l=6.15e-07 $layer=LI1_cond $X=13.255 $Y=1.65
+ $X2=13.255 $Y2=2.265
r138 40 56 6.46576 $w=2.5e-07 $l=1.65e-07 $layer=LI1_cond $X=13.045 $Y=1.32
+ $X2=12.88 $Y2=1.32
r139 40 42 28.1126 $w=3.28e-07 $l=8.05e-07 $layer=LI1_cond $X=13.045 $Y=1.32
+ $X2=13.045 $Y2=0.515
r140 36 38 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=15.335 $Y=1.765
+ $X2=15.335 $Y2=2.4
r141 35 36 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=15.335 $Y=1.675
+ $X2=15.335 $Y2=1.765
r142 34 39 18.8402 $w=1.65e-07 $l=8.57321e-08 $layer=POLY_cond $X=15.335 $Y=1.47
+ $X2=15.312 $Y2=1.395
r143 34 35 79.6855 $w=1.8e-07 $l=2.05e-07 $layer=POLY_cond $X=15.335 $Y=1.47
+ $X2=15.335 $Y2=1.675
r144 30 39 18.8402 $w=1.65e-07 $l=9.16515e-08 $layer=POLY_cond $X=15.275 $Y=1.32
+ $X2=15.312 $Y2=1.395
r145 30 32 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=15.275 $Y=1.32
+ $X2=15.275 $Y2=0.74
r146 29 64 29.6209 $w=3.78e-07 $l=1.86652e-07 $layer=POLY_cond $X=14.975
+ $Y=1.395 $X2=14.885 $Y2=1.542
r147 28 39 6.66866 $w=1.5e-07 $l=1.12e-07 $layer=POLY_cond $X=15.2 $Y=1.395
+ $X2=15.312 $Y2=1.395
r148 28 29 115.372 $w=1.5e-07 $l=2.25e-07 $layer=POLY_cond $X=15.2 $Y=1.395
+ $X2=14.975 $Y2=1.395
r149 25 64 24.4846 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=14.885 $Y=1.765
+ $X2=14.885 $Y2=1.542
r150 25 27 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=14.885 $Y=1.765
+ $X2=14.885 $Y2=2.4
r151 21 63 24.4846 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=14.845 $Y=1.32
+ $X2=14.845 $Y2=1.542
r152 21 23 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=14.845 $Y=1.32
+ $X2=14.845 $Y2=0.74
r153 18 61 24.4846 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=14.435 $Y=1.765
+ $X2=14.435 $Y2=1.542
r154 18 20 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=14.435 $Y=1.765
+ $X2=14.435 $Y2=2.4
r155 14 60 24.4846 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=14.345 $Y=1.32
+ $X2=14.345 $Y2=1.542
r156 14 16 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=14.345 $Y=1.32
+ $X2=14.345 $Y2=0.74
r157 11 59 24.4846 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=13.985 $Y=1.765
+ $X2=13.985 $Y2=1.542
r158 11 13 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=13.985 $Y=1.765
+ $X2=13.985 $Y2=2.4
r159 7 57 24.4846 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=13.76 $Y=1.32
+ $X2=13.76 $Y2=1.542
r160 7 9 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=13.76 $Y=1.32
+ $X2=13.76 $Y2=0.74
r161 2 46 300 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=2 $X=13.105
+ $Y=2.12 $X2=13.255 $Y2=2.265
r162 1 42 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=12.9
+ $Y=0.37 $X2=13.045 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__SDFSTP_4%VPWR 1 2 3 4 5 6 7 8 9 10 11 36 40 42 46 50
+ 54 58 62 66 70 74 76 78 83 84 86 87 88 90 95 100 115 122 127 132 137 143 146
+ 149 152 155 158 161 164 168
c213 46 0 1.33164e-19 $X=3.735 $Y=2.78
r214 167 168 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=15.6 $Y=3.33
+ $X2=15.6 $Y2=3.33
r215 164 165 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=14.64 $Y=3.33
+ $X2=14.64 $Y2=3.33
r216 161 162 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.68 $Y=3.33
+ $X2=13.68 $Y2=3.33
r217 158 159 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=12.72 $Y=3.33
+ $X2=12.72 $Y2=3.33
r218 155 156 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.28 $Y=3.33
+ $X2=11.28 $Y2=3.33
r219 152 153 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r220 149 150 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r221 147 150 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.6 $Y2=3.33
r222 146 147 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r223 143 144 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r224 141 168 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=15.12 $Y=3.33
+ $X2=15.6 $Y2=3.33
r225 141 165 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=15.12 $Y=3.33
+ $X2=14.64 $Y2=3.33
r226 140 141 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=15.12 $Y=3.33
+ $X2=15.12 $Y2=3.33
r227 138 164 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=14.825 $Y=3.33
+ $X2=14.66 $Y2=3.33
r228 138 140 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=14.825 $Y=3.33
+ $X2=15.12 $Y2=3.33
r229 137 167 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=15.395 $Y=3.33
+ $X2=15.617 $Y2=3.33
r230 137 140 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=15.395 $Y=3.33
+ $X2=15.12 $Y2=3.33
r231 136 165 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=14.16 $Y=3.33
+ $X2=14.64 $Y2=3.33
r232 136 162 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=14.16 $Y=3.33
+ $X2=13.68 $Y2=3.33
r233 135 136 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=14.16 $Y=3.33
+ $X2=14.16 $Y2=3.33
r234 133 161 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=13.87 $Y=3.33
+ $X2=13.705 $Y2=3.33
r235 133 135 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=13.87 $Y=3.33
+ $X2=14.16 $Y2=3.33
r236 132 164 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=14.495 $Y=3.33
+ $X2=14.66 $Y2=3.33
r237 132 135 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=14.495 $Y=3.33
+ $X2=14.16 $Y2=3.33
r238 131 162 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=13.2 $Y=3.33
+ $X2=13.68 $Y2=3.33
r239 131 159 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=13.2 $Y=3.33
+ $X2=12.72 $Y2=3.33
r240 130 131 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.2 $Y=3.33
+ $X2=13.2 $Y2=3.33
r241 128 158 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=12.97 $Y=3.33
+ $X2=12.845 $Y2=3.33
r242 128 130 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=12.97 $Y=3.33
+ $X2=13.2 $Y2=3.33
r243 127 161 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=13.54 $Y=3.33
+ $X2=13.705 $Y2=3.33
r244 127 130 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=13.54 $Y=3.33
+ $X2=13.2 $Y2=3.33
r245 126 159 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=11.76 $Y=3.33
+ $X2=12.72 $Y2=3.33
r246 126 156 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.76 $Y=3.33
+ $X2=11.28 $Y2=3.33
r247 125 126 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=11.76 $Y=3.33
+ $X2=11.76 $Y2=3.33
r248 123 155 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=11.375 $Y=3.33
+ $X2=11.25 $Y2=3.33
r249 123 125 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=11.375 $Y=3.33
+ $X2=11.76 $Y2=3.33
r250 122 158 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=12.72 $Y=3.33
+ $X2=12.845 $Y2=3.33
r251 122 125 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=12.72 $Y=3.33
+ $X2=11.76 $Y2=3.33
r252 121 156 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.8 $Y=3.33
+ $X2=11.28 $Y2=3.33
r253 120 121 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=10.8 $Y=3.33
+ $X2=10.8 $Y2=3.33
r254 118 121 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=8.88 $Y=3.33
+ $X2=10.8 $Y2=3.33
r255 117 120 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=8.88 $Y=3.33
+ $X2=10.8 $Y2=3.33
r256 117 118 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r257 115 155 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=11.125 $Y=3.33
+ $X2=11.25 $Y2=3.33
r258 115 120 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=11.125 $Y=3.33
+ $X2=10.8 $Y2=3.33
r259 114 118 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=3.33
+ $X2=8.88 $Y2=3.33
r260 113 114 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.4 $Y=3.33
+ $X2=8.4 $Y2=3.33
r261 111 153 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=6.48 $Y2=3.33
r262 110 111 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r263 108 152 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.525 $Y=3.33
+ $X2=6.4 $Y2=3.33
r264 108 110 59.6952 $w=1.68e-07 $l=9.15e-07 $layer=LI1_cond $X=6.525 $Y=3.33
+ $X2=7.44 $Y2=3.33
r265 107 153 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=3.33
+ $X2=6.48 $Y2=3.33
r266 106 107 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r267 104 107 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=6 $Y2=3.33
r268 104 150 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=3.6 $Y2=3.33
r269 103 106 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=4.08 $Y=3.33
+ $X2=6 $Y2=3.33
r270 103 104 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r271 101 149 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.9 $Y=3.33
+ $X2=3.735 $Y2=3.33
r272 101 103 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=3.9 $Y=3.33
+ $X2=4.08 $Y2=3.33
r273 100 152 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.275 $Y=3.33
+ $X2=6.4 $Y2=3.33
r274 100 106 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=6.275 $Y=3.33
+ $X2=6 $Y2=3.33
r275 99 147 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.64 $Y2=3.33
r276 99 144 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r277 98 99 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r278 96 143 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.885 $Y=3.33
+ $X2=0.72 $Y2=3.33
r279 96 98 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=0.885 $Y=3.33
+ $X2=1.2 $Y2=3.33
r280 95 146 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.56 $Y=3.33
+ $X2=2.725 $Y2=3.33
r281 95 98 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=2.56 $Y=3.33
+ $X2=1.2 $Y2=3.33
r282 93 144 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r283 92 93 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r284 90 143 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.555 $Y=3.33
+ $X2=0.72 $Y2=3.33
r285 90 92 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=0.555 $Y=3.33
+ $X2=0.24 $Y2=3.33
r286 88 114 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=3.33
+ $X2=8.4 $Y2=3.33
r287 88 111 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=3.33
+ $X2=7.44 $Y2=3.33
r288 86 113 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=8.535 $Y=3.33
+ $X2=8.4 $Y2=3.33
r289 86 87 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.535 $Y=3.33
+ $X2=8.7 $Y2=3.33
r290 85 117 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=8.865 $Y=3.33
+ $X2=8.88 $Y2=3.33
r291 85 87 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.865 $Y=3.33
+ $X2=8.7 $Y2=3.33
r292 83 110 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=7.715 $Y=3.33
+ $X2=7.44 $Y2=3.33
r293 83 84 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.715 $Y=3.33
+ $X2=7.8 $Y2=3.33
r294 82 113 33.5989 $w=1.68e-07 $l=5.15e-07 $layer=LI1_cond $X=7.885 $Y=3.33
+ $X2=8.4 $Y2=3.33
r295 82 84 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.885 $Y=3.33
+ $X2=7.8 $Y2=3.33
r296 78 81 24.4458 $w=3.28e-07 $l=7e-07 $layer=LI1_cond $X=15.56 $Y=2.115
+ $X2=15.56 $Y2=2.815
r297 76 167 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=15.56 $Y=3.245
+ $X2=15.617 $Y2=3.33
r298 76 81 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=15.56 $Y=3.245
+ $X2=15.56 $Y2=2.815
r299 72 164 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=14.66 $Y=3.245
+ $X2=14.66 $Y2=3.33
r300 72 74 29.3349 $w=3.28e-07 $l=8.4e-07 $layer=LI1_cond $X=14.66 $Y=3.245
+ $X2=14.66 $Y2=2.405
r301 68 161 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=13.705 $Y=3.245
+ $X2=13.705 $Y2=3.33
r302 68 70 34.2241 $w=3.28e-07 $l=9.8e-07 $layer=LI1_cond $X=13.705 $Y=3.245
+ $X2=13.705 $Y2=2.265
r303 64 158 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=12.845 $Y=3.245
+ $X2=12.845 $Y2=3.33
r304 64 66 22.8184 $w=2.48e-07 $l=4.95e-07 $layer=LI1_cond $X=12.845 $Y=3.245
+ $X2=12.845 $Y2=2.75
r305 60 155 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=11.25 $Y=3.245
+ $X2=11.25 $Y2=3.33
r306 60 62 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=11.25 $Y=3.245
+ $X2=11.25 $Y2=2.815
r307 56 87 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.7 $Y=3.245 $X2=8.7
+ $Y2=3.33
r308 56 58 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=8.7 $Y=3.245
+ $X2=8.7 $Y2=2.55
r309 52 84 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.8 $Y=3.245 $X2=7.8
+ $Y2=3.33
r310 52 54 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=7.8 $Y=3.245
+ $X2=7.8 $Y2=2.505
r311 48 152 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.4 $Y=3.245
+ $X2=6.4 $Y2=3.33
r312 48 50 20.744 $w=2.48e-07 $l=4.5e-07 $layer=LI1_cond $X=6.4 $Y=3.245 $X2=6.4
+ $Y2=2.795
r313 44 149 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.735 $Y=3.245
+ $X2=3.735 $Y2=3.33
r314 44 46 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=3.735 $Y=3.245
+ $X2=3.735 $Y2=2.78
r315 43 146 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.89 $Y=3.33
+ $X2=2.725 $Y2=3.33
r316 42 149 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.57 $Y=3.33
+ $X2=3.735 $Y2=3.33
r317 42 43 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=3.57 $Y=3.33
+ $X2=2.89 $Y2=3.33
r318 38 146 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.725 $Y=3.245
+ $X2=2.725 $Y2=3.33
r319 38 40 8.73063 $w=3.28e-07 $l=2.5e-07 $layer=LI1_cond $X=2.725 $Y=3.245
+ $X2=2.725 $Y2=2.995
r320 34 143 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.72 $Y=3.245
+ $X2=0.72 $Y2=3.33
r321 34 36 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=0.72 $Y=3.245
+ $X2=0.72 $Y2=2.78
r322 11 81 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=15.41
+ $Y=1.84 $X2=15.56 $Y2=2.815
r323 11 78 400 $w=1.7e-07 $l=3.4187e-07 $layer=licon1_PDIFF $count=1 $X=15.41
+ $Y=1.84 $X2=15.56 $Y2=2.115
r324 10 74 300 $w=1.7e-07 $l=6.3559e-07 $layer=licon1_PDIFF $count=2 $X=14.51
+ $Y=1.84 $X2=14.66 $Y2=2.405
r325 9 70 300 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=2 $X=13.555
+ $Y=2.12 $X2=13.705 $Y2=2.265
r326 8 66 600 $w=1.7e-07 $l=2.95212e-07 $layer=licon1_PDIFF $count=1 $X=12.6
+ $Y=2.54 $X2=12.805 $Y2=2.75
r327 7 62 600 $w=1.7e-07 $l=3.4187e-07 $layer=licon1_PDIFF $count=1 $X=11.14
+ $Y=2.54 $X2=11.29 $Y2=2.815
r328 6 58 600 $w=1.7e-07 $l=7.5629e-07 $layer=licon1_PDIFF $count=1 $X=8.55
+ $Y=1.865 $X2=8.7 $Y2=2.55
r329 5 54 600 $w=1.7e-07 $l=4.77493e-07 $layer=licon1_PDIFF $count=1 $X=7.42
+ $Y=2.285 $X2=7.8 $Y2=2.505
r330 4 50 600 $w=1.7e-07 $l=6.16401e-07 $layer=licon1_PDIFF $count=1 $X=6.205
+ $Y=2.285 $X2=6.44 $Y2=2.795
r331 3 46 600 $w=1.7e-07 $l=1.01223e-06 $layer=licon1_PDIFF $count=1 $X=3.585
+ $Y=1.84 $X2=3.735 $Y2=2.78
r332 2 40 600 $w=1.7e-07 $l=7.83741e-07 $layer=licon1_PDIFF $count=1 $X=2.49
+ $Y=2.32 $X2=2.725 $Y2=2.995
r333 1 36 600 $w=1.7e-07 $l=5.29717e-07 $layer=licon1_PDIFF $count=1 $X=0.57
+ $Y=2.32 $X2=0.72 $Y2=2.78
.ends

.subckt PM_SKY130_FD_SC_HS__SDFSTP_4%A_288_464# 1 2 3 4 13 18 19 20 22 23 25 28
+ 32 34 37 44 46
c123 28 0 1.2825e-19 $X=4.495 $Y=1.9
c124 22 0 4.43302e-20 $X=2.3 $Y=2.49
r125 46 48 4.07466 $w=5.09e-07 $l=1.7e-07 $layer=LI1_cond $X=4.72 $Y=2.325
+ $X2=4.72 $Y2=2.495
r126 41 44 7.68295 $w=3.28e-07 $l=2.2e-07 $layer=LI1_cond $X=4.495 $Y=0.76
+ $X2=4.715 $Y2=0.76
r127 37 39 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=3.09 $Y=2.325
+ $X2=3.09 $Y2=2.575
r128 30 32 5.5876 $w=3.28e-07 $l=1.6e-07 $layer=LI1_cond $X=1.715 $Y=0.575
+ $X2=1.875 $Y2=0.575
r129 28 46 15.9959 $w=5.09e-07 $l=5.25595e-07 $layer=LI1_cond $X=4.495 $Y=1.9
+ $X2=4.72 $Y2=2.325
r130 27 41 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.495 $Y=0.925
+ $X2=4.495 $Y2=0.76
r131 27 28 63.6096 $w=1.68e-07 $l=9.75e-07 $layer=LI1_cond $X=4.495 $Y=0.925
+ $X2=4.495 $Y2=1.9
r132 26 37 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.175 $Y=2.325
+ $X2=3.09 $Y2=2.325
r133 25 46 7.26882 $w=1.7e-07 $l=3.1e-07 $layer=LI1_cond $X=4.41 $Y=2.325
+ $X2=4.72 $Y2=2.325
r134 25 26 80.5722 $w=1.68e-07 $l=1.235e-06 $layer=LI1_cond $X=4.41 $Y=2.325
+ $X2=3.175 $Y2=2.325
r135 24 34 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.385 $Y=2.575
+ $X2=2.3 $Y2=2.575
r136 23 39 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.005 $Y=2.575
+ $X2=3.09 $Y2=2.575
r137 23 24 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=3.005 $Y=2.575
+ $X2=2.385 $Y2=2.575
r138 22 34 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=2.3 $Y=2.49 $X2=2.3
+ $Y2=2.575
r139 21 22 91.9893 $w=1.68e-07 $l=1.41e-06 $layer=LI1_cond $X=2.3 $Y=1.08
+ $X2=2.3 $Y2=2.49
r140 19 21 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.215 $Y=0.995
+ $X2=2.3 $Y2=1.08
r141 19 20 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=2.215 $Y=0.995
+ $X2=1.96 $Y2=0.995
r142 18 20 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.875 $Y=0.91
+ $X2=1.96 $Y2=0.995
r143 17 32 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.875 $Y=0.74
+ $X2=1.875 $Y2=0.575
r144 17 18 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=1.875 $Y=0.74
+ $X2=1.875 $Y2=0.91
r145 13 34 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=2.3 $Y=2.785
+ $X2=2.3 $Y2=2.575
r146 13 15 24.6623 $w=2.48e-07 $l=5.35e-07 $layer=LI1_cond $X=2.215 $Y=2.785
+ $X2=1.68 $Y2=2.785
r147 4 48 600 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_PDIFF $count=1 $X=4.72
+ $Y=2.285 $X2=4.865 $Y2=2.495
r148 3 15 600 $w=1.7e-07 $l=5.31625e-07 $layer=licon1_PDIFF $count=1 $X=1.44
+ $Y=2.32 $X2=1.68 $Y2=2.745
r149 2 44 182 $w=1.7e-07 $l=4.21307e-07 $layer=licon1_NDIFF $count=1 $X=4.57
+ $Y=0.405 $X2=4.715 $Y2=0.76
r150 1 30 182 $w=1.7e-07 $l=3.005e-07 $layer=licon1_NDIFF $count=1 $X=1.5
+ $Y=0.37 $X2=1.715 $Y2=0.575
.ends

.subckt PM_SKY130_FD_SC_HS__SDFSTP_4%A_1620_373# 1 2 7 9 11 18
c33 18 0 2.89568e-19 $X=9.71 $Y=2.265
c34 9 0 7.58781e-20 $X=8.25 $Y=2.55
c35 7 0 1.49656e-19 $X=8.225 $Y=2.29
r36 12 16 4.57959 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=8.365 $Y=2.205
+ $X2=8.225 $Y2=2.205
r37 11 18 5.03363 $w=1.7e-07 $l=1.69926e-07 $layer=LI1_cond $X=9.545 $Y=2.205
+ $X2=9.71 $Y2=2.195
r38 11 12 76.984 $w=1.68e-07 $l=1.18e-06 $layer=LI1_cond $X=9.545 $Y=2.205
+ $X2=8.365 $Y2=2.205
r39 7 16 2.78046 $w=2.8e-07 $l=8.5e-08 $layer=LI1_cond $X=8.225 $Y=2.29
+ $X2=8.225 $Y2=2.205
r40 7 9 10.7013 $w=2.78e-07 $l=2.6e-07 $layer=LI1_cond $X=8.225 $Y=2.29
+ $X2=8.225 $Y2=2.55
r41 2 18 300 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=2 $X=9.56
+ $Y=2.12 $X2=9.71 $Y2=2.265
r42 1 16 600 $w=1.7e-07 $l=4.08167e-07 $layer=licon1_PDIFF $count=1 $X=8.1
+ $Y=1.865 $X2=8.25 $Y2=2.205
r43 1 9 600 $w=1.7e-07 $l=7.5629e-07 $layer=licon1_PDIFF $count=1 $X=8.1
+ $Y=1.865 $X2=8.25 $Y2=2.55
.ends

.subckt PM_SKY130_FD_SC_HS__SDFSTP_4%Q 1 2 3 4 15 17 19 21 22 23 27 31 33 35 39
+ 43 45 48
c84 35 0 2.92295e-20 $X=15.485 $Y=1.355
c85 21 0 2.40437e-20 $X=14.895 $Y=1.065
r86 45 48 2.9826 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=15.6 $Y=1.695 $X2=15.6
+ $Y2=1.61
r87 45 48 0.751593 $w=2.28e-07 $l=1.5e-08 $layer=LI1_cond $X=15.6 $Y=1.595
+ $X2=15.6 $Y2=1.61
r88 44 45 7.76646 $w=2.28e-07 $l=1.55e-07 $layer=LI1_cond $X=15.6 $Y=1.44
+ $X2=15.6 $Y2=1.595
r89 39 40 10.1275 $w=3.28e-07 $l=2.9e-07 $layer=LI1_cond $X=15.06 $Y=1.065
+ $X2=15.06 $Y2=1.355
r90 36 40 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=15.225 $Y=1.355
+ $X2=15.06 $Y2=1.355
r91 35 44 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=15.485 $Y=1.355
+ $X2=15.6 $Y2=1.44
r92 35 36 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=15.485 $Y=1.355
+ $X2=15.225 $Y2=1.355
r93 34 43 3.70735 $w=2.5e-07 $l=2.23495e-07 $layer=LI1_cond $X=15.195 $Y=1.695
+ $X2=15.11 $Y2=1.88
r94 33 45 4.03528 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=15.485 $Y=1.695
+ $X2=15.6 $Y2=1.695
r95 33 34 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=15.485 $Y=1.695
+ $X2=15.195 $Y2=1.695
r96 29 43 2.76166 $w=1.7e-07 $l=2.7e-07 $layer=LI1_cond $X=15.11 $Y=2.15
+ $X2=15.11 $Y2=1.88
r97 29 31 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=15.11 $Y=2.15
+ $X2=15.11 $Y2=2.4
r98 25 39 2.96841 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=15.06 $Y=0.98
+ $X2=15.06 $Y2=1.065
r99 25 27 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=15.06 $Y=0.98
+ $X2=15.06 $Y2=0.515
r100 24 38 3.1563 $w=3.3e-07 $l=1.4e-07 $layer=LI1_cond $X=14.325 $Y=1.985
+ $X2=14.185 $Y2=1.985
r101 23 43 3.70735 $w=2.5e-07 $l=1.41244e-07 $layer=LI1_cond $X=15.025 $Y=1.985
+ $X2=15.11 $Y2=1.88
r102 23 24 24.4458 $w=3.28e-07 $l=7e-07 $layer=LI1_cond $X=15.025 $Y=1.985
+ $X2=14.325 $Y2=1.985
r103 21 39 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=14.895 $Y=1.065
+ $X2=15.06 $Y2=1.065
r104 21 22 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=14.895 $Y=1.065
+ $X2=14.225 $Y2=1.065
r105 17 38 3.71993 $w=2.8e-07 $l=1.65e-07 $layer=LI1_cond $X=14.185 $Y=2.15
+ $X2=14.185 $Y2=1.985
r106 17 19 10.2897 $w=2.78e-07 $l=2.5e-07 $layer=LI1_cond $X=14.185 $Y=2.15
+ $X2=14.185 $Y2=2.4
r107 13 22 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=14.06 $Y=0.98
+ $X2=14.225 $Y2=1.065
r108 13 15 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=14.06 $Y=0.98
+ $X2=14.06 $Y2=0.515
r109 4 43 600 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=14.96
+ $Y=1.84 $X2=15.11 $Y2=1.985
r110 4 31 300 $w=1.7e-07 $l=6.30555e-07 $layer=licon1_PDIFF $count=2 $X=14.96
+ $Y=1.84 $X2=15.11 $Y2=2.4
r111 3 38 600 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=14.06
+ $Y=1.84 $X2=14.21 $Y2=1.985
r112 3 19 300 $w=1.7e-07 $l=6.30555e-07 $layer=licon1_PDIFF $count=2 $X=14.06
+ $Y=1.84 $X2=14.21 $Y2=2.4
r113 2 27 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=14.92
+ $Y=0.37 $X2=15.06 $Y2=0.515
r114 1 15 91 $w=1.7e-07 $l=2.88531e-07 $layer=licon1_NDIFF $count=2 $X=13.835
+ $Y=0.37 $X2=14.06 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__SDFSTP_4%VGND 1 2 3 4 5 6 7 8 9 10 33 37 39 43 47 51
+ 57 61 65 69 71 73 76 77 78 80 85 93 101 106 111 126 130 136 139 142 145 148
+ 151 154 157 161
c176 73 0 1.69241e-19 $X=15.56 $Y=0.515
r177 160 161 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=15.6 $Y=0
+ $X2=15.6 $Y2=0
r178 157 158 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=14.64 $Y=0
+ $X2=14.64 $Y2=0
r179 154 155 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.76 $Y=0
+ $X2=11.76 $Y2=0
r180 151 152 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=0
+ $X2=8.88 $Y2=0
r181 145 146 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6.48 $Y=0
+ $X2=6.48 $Y2=0
r182 142 143 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r183 140 143 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=0
+ $X2=3.6 $Y2=0
r184 139 140 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0
+ $X2=2.64 $Y2=0
r185 136 137 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0
+ $X2=0.72 $Y2=0
r186 134 161 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=15.12 $Y=0
+ $X2=15.6 $Y2=0
r187 134 158 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=15.12 $Y=0
+ $X2=14.64 $Y2=0
r188 133 134 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=15.12 $Y=0
+ $X2=15.12 $Y2=0
r189 131 157 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=14.725 $Y=0
+ $X2=14.56 $Y2=0
r190 131 133 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=14.725 $Y=0
+ $X2=15.12 $Y2=0
r191 130 160 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=15.395 $Y=0
+ $X2=15.617 $Y2=0
r192 130 133 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=15.395 $Y=0
+ $X2=15.12 $Y2=0
r193 129 158 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=14.16 $Y=0
+ $X2=14.64 $Y2=0
r194 128 129 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=14.16 $Y=0
+ $X2=14.16 $Y2=0
r195 126 157 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=14.395 $Y=0
+ $X2=14.56 $Y2=0
r196 126 128 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=14.395 $Y=0
+ $X2=14.16 $Y2=0
r197 125 129 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=13.2 $Y=0
+ $X2=14.16 $Y2=0
r198 124 125 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=13.2 $Y=0
+ $X2=13.2 $Y2=0
r199 122 125 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=12.24 $Y=0
+ $X2=13.2 $Y2=0
r200 122 155 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.24 $Y=0
+ $X2=11.76 $Y2=0
r201 121 124 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=12.24 $Y=0
+ $X2=13.2 $Y2=0
r202 121 122 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=12.24 $Y=0
+ $X2=12.24 $Y2=0
r203 119 154 11.2921 $w=1.7e-07 $l=2.5e-07 $layer=LI1_cond $X=12.15 $Y=0
+ $X2=11.9 $Y2=0
r204 119 121 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=12.15 $Y=0
+ $X2=12.24 $Y2=0
r205 118 155 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.28 $Y=0
+ $X2=11.76 $Y2=0
r206 117 118 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=11.28 $Y=0
+ $X2=11.28 $Y2=0
r207 115 118 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=9.36 $Y=0
+ $X2=11.28 $Y2=0
r208 115 152 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.36 $Y=0
+ $X2=8.88 $Y2=0
r209 114 117 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=9.36 $Y=0
+ $X2=11.28 $Y2=0
r210 114 115 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=9.36 $Y=0
+ $X2=9.36 $Y2=0
r211 112 151 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.12 $Y=0
+ $X2=8.955 $Y2=0
r212 112 114 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=9.12 $Y=0
+ $X2=9.36 $Y2=0
r213 111 154 11.2921 $w=1.7e-07 $l=2.5e-07 $layer=LI1_cond $X=11.65 $Y=0
+ $X2=11.9 $Y2=0
r214 111 117 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=11.65 $Y=0
+ $X2=11.28 $Y2=0
r215 110 152 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=0
+ $X2=8.88 $Y2=0
r216 109 110 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r217 107 148 13.3456 $w=1.7e-07 $l=3.35e-07 $layer=LI1_cond $X=8.26 $Y=0
+ $X2=7.925 $Y2=0
r218 107 109 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=8.26 $Y=0 $X2=8.4
+ $Y2=0
r219 106 151 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.79 $Y=0
+ $X2=8.955 $Y2=0
r220 106 109 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=8.79 $Y=0 $X2=8.4
+ $Y2=0
r221 105 146 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=7.44 $Y=0
+ $X2=6.48 $Y2=0
r222 104 105 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=7.44 $Y=0
+ $X2=7.44 $Y2=0
r223 102 145 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.54 $Y=0
+ $X2=6.375 $Y2=0
r224 102 104 58.7166 $w=1.68e-07 $l=9e-07 $layer=LI1_cond $X=6.54 $Y=0 $X2=7.44
+ $Y2=0
r225 101 148 13.3456 $w=1.7e-07 $l=3.35e-07 $layer=LI1_cond $X=7.59 $Y=0
+ $X2=7.925 $Y2=0
r226 101 104 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=7.59 $Y=0 $X2=7.44
+ $Y2=0
r227 100 146 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=0 $X2=6.48
+ $Y2=0
r228 99 100 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6 $Y=0 $X2=6
+ $Y2=0
r229 97 100 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=4.08 $Y=0 $X2=6
+ $Y2=0
r230 97 143 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=3.6
+ $Y2=0
r231 96 99 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=4.08 $Y=0 $X2=6
+ $Y2=0
r232 96 97 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.08 $Y=0
+ $X2=4.08 $Y2=0
r233 94 142 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.89 $Y=0
+ $X2=3.725 $Y2=0
r234 94 96 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=3.89 $Y=0 $X2=4.08
+ $Y2=0
r235 93 145 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.21 $Y=0
+ $X2=6.375 $Y2=0
r236 93 99 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=6.21 $Y=0 $X2=6
+ $Y2=0
r237 92 140 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0
+ $X2=2.64 $Y2=0
r238 91 92 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r239 89 92 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r240 89 137 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r241 88 91 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r242 88 89 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r243 86 136 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.945 $Y=0
+ $X2=0.78 $Y2=0
r244 86 88 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.945 $Y=0 $X2=1.2
+ $Y2=0
r245 85 139 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.45 $Y=0
+ $X2=2.615 $Y2=0
r246 85 91 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=2.45 $Y=0 $X2=2.16
+ $Y2=0
r247 83 137 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0
+ $X2=0.72 $Y2=0
r248 82 83 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r249 80 136 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.615 $Y=0
+ $X2=0.78 $Y2=0
r250 80 82 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=0.615 $Y=0
+ $X2=0.24 $Y2=0
r251 78 110 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=0 $X2=8.4
+ $Y2=0
r252 78 105 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=0
+ $X2=7.44 $Y2=0
r253 78 148 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=0 $X2=7.92
+ $Y2=0
r254 76 124 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=13.38 $Y=0
+ $X2=13.2 $Y2=0
r255 76 77 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=13.38 $Y=0
+ $X2=13.545 $Y2=0
r256 75 128 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=13.71 $Y=0
+ $X2=14.16 $Y2=0
r257 75 77 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=13.71 $Y=0
+ $X2=13.545 $Y2=0
r258 71 160 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=15.56 $Y=0.085
+ $X2=15.617 $Y2=0
r259 71 73 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=15.56 $Y=0.085
+ $X2=15.56 $Y2=0.515
r260 67 157 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=14.56 $Y=0.085
+ $X2=14.56 $Y2=0
r261 67 69 19.5566 $w=3.28e-07 $l=5.6e-07 $layer=LI1_cond $X=14.56 $Y=0.085
+ $X2=14.56 $Y2=0.645
r262 63 77 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=13.545 $Y=0.085
+ $X2=13.545 $Y2=0
r263 63 65 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=13.545 $Y=0.085
+ $X2=13.545 $Y2=0.515
r264 59 154 2.07448 $w=5e-07 $l=8.5e-08 $layer=LI1_cond $X=11.9 $Y=0.085
+ $X2=11.9 $Y2=0
r265 59 61 10.2863 $w=4.98e-07 $l=4.3e-07 $layer=LI1_cond $X=11.9 $Y=0.085
+ $X2=11.9 $Y2=0.515
r266 55 151 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.955 $Y=0.085
+ $X2=8.955 $Y2=0
r267 55 57 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=8.955 $Y=0.085
+ $X2=8.955 $Y2=0.515
r268 51 53 6.06965 $w=6.68e-07 $l=3.4e-07 $layer=LI1_cond $X=7.925 $Y=0.495
+ $X2=7.925 $Y2=0.835
r269 49 148 2.76849 $w=6.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.925 $Y=0.085
+ $X2=7.925 $Y2=0
r270 49 51 7.31929 $w=6.68e-07 $l=4.1e-07 $layer=LI1_cond $X=7.925 $Y=0.085
+ $X2=7.925 $Y2=0.495
r271 45 145 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.375 $Y=0.085
+ $X2=6.375 $Y2=0
r272 45 47 10.826 $w=3.28e-07 $l=3.1e-07 $layer=LI1_cond $X=6.375 $Y=0.085
+ $X2=6.375 $Y2=0.395
r273 41 142 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.725 $Y=0.085
+ $X2=3.725 $Y2=0
r274 41 43 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=3.725 $Y=0.085
+ $X2=3.725 $Y2=0.515
r275 40 139 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.78 $Y=0
+ $X2=2.615 $Y2=0
r276 39 142 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.56 $Y=0
+ $X2=3.725 $Y2=0
r277 39 40 50.8877 $w=1.68e-07 $l=7.8e-07 $layer=LI1_cond $X=3.56 $Y=0 $X2=2.78
+ $Y2=0
r278 35 139 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.615 $Y=0.085
+ $X2=2.615 $Y2=0
r279 35 37 16.0644 $w=3.28e-07 $l=4.6e-07 $layer=LI1_cond $X=2.615 $Y=0.085
+ $X2=2.615 $Y2=0.545
r280 31 136 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.78 $Y=0.085
+ $X2=0.78 $Y2=0
r281 31 33 16.0644 $w=3.28e-07 $l=4.6e-07 $layer=LI1_cond $X=0.78 $Y=0.085
+ $X2=0.78 $Y2=0.545
r282 10 73 91 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=2 $X=15.35
+ $Y=0.37 $X2=15.56 $Y2=0.515
r283 9 69 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=14.42
+ $Y=0.37 $X2=14.56 $Y2=0.645
r284 8 65 91 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=2 $X=13.335
+ $Y=0.37 $X2=13.545 $Y2=0.515
r285 7 61 182 $w=1.7e-07 $l=2.88531e-07 $layer=licon1_NDIFF $count=1 $X=11.675
+ $Y=0.37 $X2=11.9 $Y2=0.515
r286 6 57 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=8.815
+ $Y=0.37 $X2=8.955 $Y2=0.515
r287 5 53 121.333 $w=1.7e-07 $l=6.73498e-07 $layer=licon1_NDIFF $count=1
+ $X=7.615 $Y=0.37 $X2=8.095 $Y2=0.835
r288 5 51 121.333 $w=1.7e-07 $l=5.38888e-07 $layer=licon1_NDIFF $count=1
+ $X=7.615 $Y=0.37 $X2=8.095 $Y2=0.495
r289 4 47 182 $w=1.7e-07 $l=2.24944e-07 $layer=licon1_NDIFF $count=1 $X=6.155
+ $Y=0.405 $X2=6.375 $Y2=0.395
r290 3 43 91 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=2 $X=3.515
+ $Y=0.37 $X2=3.725 $Y2=0.515
r291 2 37 182 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_NDIFF $count=1 $X=2.475
+ $Y=0.37 $X2=2.615 $Y2=0.545
r292 1 33 182 $w=1.7e-07 $l=2.84341e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.37 $X2=0.78 $Y2=0.545
.ends

.subckt PM_SKY130_FD_SC_HS__SDFSTP_4%A_1677_74# 1 2 9 11 12 15
c36 9 0 1.22616e-19 $X=8.525 $Y=0.515
r37 13 15 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=9.945 $Y=1.11
+ $X2=9.945 $Y2=0.81
r38 11 13 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.86 $Y=1.195
+ $X2=9.945 $Y2=1.11
r39 11 12 81.5508 $w=1.68e-07 $l=1.25e-06 $layer=LI1_cond $X=9.86 $Y=1.195
+ $X2=8.61 $Y2=1.195
r40 7 12 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.525 $Y=1.11
+ $X2=8.61 $Y2=1.195
r41 7 9 38.8182 $w=1.68e-07 $l=5.95e-07 $layer=LI1_cond $X=8.525 $Y=1.11
+ $X2=8.525 $Y2=0.515
r42 2 15 182 $w=1.7e-07 $l=5.05173e-07 $layer=licon1_NDIFF $count=1 $X=9.805
+ $Y=0.37 $X2=9.945 $Y2=0.81
r43 1 9 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=8.385
+ $Y=0.37 $X2=8.525 $Y2=0.515
.ends

