* File: sky130_fd_sc_hs__xor3_1.pex.spice
* Created: Tue Sep  1 20:26:07 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HS__XOR3_1%A_84_108# 1 2 3 4 15 17 19 22 25 26 30 35 37
+ 38 40 43 45 46 51
r111 49 51 5.5876 $w=3.28e-07 $l=1.6e-07 $layer=LI1_cond $X=4.15 $Y=1.1 $X2=4.31
+ $Y2=1.1
r112 45 47 19.8947 $w=6.68e-07 $l=6.85e-07 $layer=LI1_cond $X=4.06 $Y=2.07
+ $X2=4.06 $Y2=2.755
r113 45 46 10.6117 $w=6.68e-07 $l=1.65e-07 $layer=LI1_cond $X=4.06 $Y=2.07
+ $X2=4.06 $Y2=1.905
r114 41 51 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.31 $Y=1.265
+ $X2=4.31 $Y2=1.1
r115 41 46 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=4.31 $Y=1.265
+ $X2=4.31 $Y2=1.905
r116 40 47 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=3.81 $Y=2.905
+ $X2=3.81 $Y2=2.755
r117 37 40 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.725 $Y=2.99
+ $X2=3.81 $Y2=2.905
r118 37 38 132.112 $w=1.68e-07 $l=2.025e-06 $layer=LI1_cond $X=3.725 $Y=2.99
+ $X2=1.7 $Y2=2.99
r119 33 43 3.70735 $w=2.5e-07 $l=1.7e-07 $layer=LI1_cond $X=1.54 $Y=1.92
+ $X2=1.37 $Y2=1.92
r120 33 35 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=1.54 $Y=1.92
+ $X2=1.54 $Y2=1.165
r121 30 32 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=1.535 $Y=2.105
+ $X2=1.535 $Y2=2.815
r122 28 38 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.535 $Y=2.905
+ $X2=1.7 $Y2=2.99
r123 28 32 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=1.535 $Y=2.905
+ $X2=1.535 $Y2=2.815
r124 27 43 3.70735 $w=2.5e-07 $l=2.38642e-07 $layer=LI1_cond $X=1.535 $Y=2.09
+ $X2=1.37 $Y2=1.92
r125 27 30 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=1.535 $Y=2.09
+ $X2=1.535 $Y2=2.105
r126 25 43 2.76166 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.37 $Y=2.005
+ $X2=1.37 $Y2=1.92
r127 25 26 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=1.37 $Y=2.005
+ $X2=0.75 $Y2=2.005
r128 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.585
+ $Y=1.635 $X2=0.585 $Y2=1.635
r129 20 26 7.72402 $w=1.7e-07 $l=2.01057e-07 $layer=LI1_cond $X=0.587 $Y=1.92
+ $X2=0.75 $Y2=2.005
r130 20 22 10.106 $w=3.23e-07 $l=2.85e-07 $layer=LI1_cond $X=0.587 $Y=1.92
+ $X2=0.587 $Y2=1.635
r131 17 23 52.2586 $w=2.99e-07 $l=2.85044e-07 $layer=POLY_cond $X=0.66 $Y=1.885
+ $X2=0.585 $Y2=1.635
r132 17 19 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=0.66 $Y=1.885
+ $X2=0.66 $Y2=2.46
r133 13 23 38.5562 $w=2.99e-07 $l=2.05122e-07 $layer=POLY_cond $X=0.495 $Y=1.47
+ $X2=0.585 $Y2=1.635
r134 13 15 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=0.495 $Y=1.47
+ $X2=0.495 $Y2=0.99
r135 4 45 300 $w=1.7e-07 $l=4.59238e-07 $layer=licon1_PDIFF $count=2 $X=3.43
+ $Y=1.895 $X2=3.81 $Y2=2.07
r136 3 32 600 $w=1.7e-07 $l=9.26971e-07 $layer=licon1_PDIFF $count=1 $X=1.385
+ $Y=1.96 $X2=1.535 $Y2=2.815
r137 3 30 300 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=2 $X=1.385
+ $Y=1.96 $X2=1.535 $Y2=2.105
r138 2 49 182 $w=1.7e-07 $l=6.10635e-07 $layer=licon1_NDIFF $count=1 $X=3.84
+ $Y=0.625 $X2=4.15 $Y2=1.1
r139 1 35 182 $w=1.7e-07 $l=5.60647e-07 $layer=licon1_NDIFF $count=1 $X=1.4
+ $Y=0.67 $X2=1.54 $Y2=1.165
.ends

.subckt PM_SKY130_FD_SC_HS__XOR3_1%A 1 3 4 6 7
r34 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.125
+ $Y=1.585 $X2=1.125 $Y2=1.585
r35 7 11 10.2833 $w=3.23e-07 $l=2.9e-07 $layer=LI1_cond $X=1.122 $Y=1.295
+ $X2=1.122 $Y2=1.585
r36 4 10 38.9663 $w=3.64e-07 $l=2.26164e-07 $layer=POLY_cond $X=1.325 $Y=1.42
+ $X2=1.18 $Y2=1.585
r37 4 6 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=1.325 $Y=1.42
+ $X2=1.325 $Y2=0.99
r38 1 10 56.8427 $w=3.64e-07 $l=3.59166e-07 $layer=POLY_cond $X=1.31 $Y=1.885
+ $X2=1.18 $Y2=1.585
r39 1 3 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=1.31 $Y=1.885
+ $X2=1.31 $Y2=2.46
.ends

.subckt PM_SKY130_FD_SC_HS__XOR3_1%A_452_288# 1 2 8 9 11 14 16 17 19 20 22 27 32
+ 34 35 36 40 43 50 51 53 55
c117 9 0 1.79271e-19 $X=2.35 $Y=1.885
r118 54 55 30.474 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=3.765 $Y=1.57
+ $X2=3.69 $Y2=1.57
r119 51 54 21.8577 $w=3.3e-07 $l=1.25e-07 $layer=POLY_cond $X=3.89 $Y=1.57
+ $X2=3.765 $Y2=1.57
r120 50 51 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.89
+ $Y=1.57 $X2=3.89 $Y2=1.57
r121 47 50 3.07318 $w=2.98e-07 $l=8e-08 $layer=LI1_cond $X=3.81 $Y=1.585
+ $X2=3.89 $Y2=1.585
r122 43 45 54.1497 $w=1.68e-07 $l=8.3e-07 $layer=LI1_cond $X=4.665 $Y=1.985
+ $X2=4.665 $Y2=2.815
r123 43 53 55.7807 $w=1.68e-07 $l=8.55e-07 $layer=LI1_cond $X=4.665 $Y=1.985
+ $X2=4.665 $Y2=1.13
r124 38 53 6.45221 $w=2.23e-07 $l=1.12e-07 $layer=LI1_cond $X=4.692 $Y=1.018
+ $X2=4.692 $Y2=1.13
r125 38 40 8.09271 $w=2.23e-07 $l=1.58e-07 $layer=LI1_cond $X=4.692 $Y=1.018
+ $X2=4.692 $Y2=0.86
r126 37 40 4.86587 $w=2.23e-07 $l=9.5e-08 $layer=LI1_cond $X=4.692 $Y=0.765
+ $X2=4.692 $Y2=0.86
r127 35 37 6.9898 $w=1.7e-07 $l=1.4854e-07 $layer=LI1_cond $X=4.58 $Y=0.68
+ $X2=4.692 $Y2=0.765
r128 35 36 44.6898 $w=1.68e-07 $l=6.85e-07 $layer=LI1_cond $X=4.58 $Y=0.68
+ $X2=3.895 $Y2=0.68
r129 34 47 4.061 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=3.81 $Y=1.435 $X2=3.81
+ $Y2=1.585
r130 33 36 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.81 $Y=0.765
+ $X2=3.895 $Y2=0.68
r131 33 34 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.81 $Y=0.765
+ $X2=3.81 $Y2=1.435
r132 25 54 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.765 $Y=1.405
+ $X2=3.765 $Y2=1.57
r133 25 27 235.872 $w=1.5e-07 $l=4.6e-07 $layer=POLY_cond $X=3.765 $Y=1.405
+ $X2=3.765 $Y2=0.945
r134 24 32 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=3.445 $Y=1.515
+ $X2=3.355 $Y2=1.515
r135 24 55 125.628 $w=1.5e-07 $l=2.45e-07 $layer=POLY_cond $X=3.445 $Y=1.515
+ $X2=3.69 $Y2=1.515
r136 20 22 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=3.355 $Y=1.82
+ $X2=3.355 $Y2=2.315
r137 19 20 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=3.355 $Y=1.73
+ $X2=3.355 $Y2=1.82
r138 18 32 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=3.355 $Y=1.59
+ $X2=3.355 $Y2=1.515
r139 18 19 54.4194 $w=1.8e-07 $l=1.4e-07 $layer=POLY_cond $X=3.355 $Y=1.59
+ $X2=3.355 $Y2=1.73
r140 17 31 38.4574 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.58 $Y=1.515
+ $X2=2.505 $Y2=1.515
r141 16 32 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=3.265 $Y=1.515
+ $X2=3.355 $Y2=1.515
r142 16 17 351.245 $w=1.5e-07 $l=6.85e-07 $layer=POLY_cond $X=3.265 $Y=1.515
+ $X2=2.58 $Y2=1.515
r143 12 31 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.505 $Y=1.44
+ $X2=2.505 $Y2=1.515
r144 12 14 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=2.505 $Y=1.44
+ $X2=2.505 $Y2=0.86
r145 9 11 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=2.35 $Y=1.885
+ $X2=2.35 $Y2=2.28
r146 8 9 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=2.35 $Y=1.795 $X2=2.35
+ $Y2=1.885
r147 7 31 79.4787 $w=1.5e-07 $l=1.55e-07 $layer=POLY_cond $X=2.35 $Y=1.515
+ $X2=2.505 $Y2=1.515
r148 7 8 79.6855 $w=1.8e-07 $l=2.05e-07 $layer=POLY_cond $X=2.35 $Y=1.59
+ $X2=2.35 $Y2=1.795
r149 2 45 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=4.52
+ $Y=1.84 $X2=4.665 $Y2=2.815
r150 2 43 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=4.52
+ $Y=1.84 $X2=4.665 $Y2=1.985
r151 1 40 182 $w=1.7e-07 $l=5.53399e-07 $layer=licon1_NDIFF $count=1 $X=4.585
+ $Y=0.37 $X2=4.72 $Y2=0.86
.ends

.subckt PM_SKY130_FD_SC_HS__XOR3_1%B 1 3 6 8 10 11 12 13 14 16 17 21 23 26 28 29
+ 31 33 36 38 40 41 42 43 48
c138 21 0 1.96802e-19 $X=3.175 $Y=0.75
c139 6 0 1.59849e-19 $X=2.005 $Y=0.75
r140 47 48 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.085
+ $Y=1.515 $X2=5.085 $Y2=1.515
r141 45 47 11.0102 $w=3.94e-07 $l=9e-08 $layer=POLY_cond $X=5.025 $Y=1.425
+ $X2=5.025 $Y2=1.515
r142 43 48 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=5.085 $Y=1.665
+ $X2=5.085 $Y2=1.515
r143 34 45 28.4597 $w=3.94e-07 $l=1.21861e-07 $layer=POLY_cond $X=4.935 $Y=1.35
+ $X2=5.025 $Y2=1.425
r144 34 36 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=4.935 $Y=1.35
+ $X2=4.935 $Y2=0.74
r145 31 47 49.8683 $w=3.94e-07 $l=3.10242e-07 $layer=POLY_cond $X=4.89 $Y=1.765
+ $X2=5.025 $Y2=1.515
r146 31 33 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=4.89 $Y=1.765
+ $X2=4.89 $Y2=2.4
r147 30 42 5.30422 $w=1.5e-07 $l=1.08e-07 $layer=POLY_cond $X=4.51 $Y=1.425
+ $X2=4.402 $Y2=1.425
r148 29 45 25.4929 $w=1.5e-07 $l=2.25e-07 $layer=POLY_cond $X=4.8 $Y=1.425
+ $X2=5.025 $Y2=1.425
r149 29 30 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=4.8 $Y=1.425
+ $X2=4.51 $Y2=1.425
r150 28 42 20.4101 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=4.435 $Y=1.35
+ $X2=4.402 $Y2=1.425
r151 27 28 561.479 $w=1.5e-07 $l=1.095e-06 $layer=POLY_cond $X=4.435 $Y=0.255
+ $X2=4.435 $Y2=1.35
r152 25 42 20.4101 $w=1.5e-07 $l=8.95824e-08 $layer=POLY_cond $X=4.37 $Y=1.5
+ $X2=4.402 $Y2=1.425
r153 25 26 807.606 $w=1.5e-07 $l=1.575e-06 $layer=POLY_cond $X=4.37 $Y=1.5
+ $X2=4.37 $Y2=3.075
r154 24 41 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.25 $Y=0.18
+ $X2=3.175 $Y2=0.18
r155 23 27 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.36 $Y=0.18
+ $X2=4.435 $Y2=0.255
r156 23 24 569.17 $w=1.5e-07 $l=1.11e-06 $layer=POLY_cond $X=4.36 $Y=0.18
+ $X2=3.25 $Y2=0.18
r157 19 41 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.175 $Y=0.255
+ $X2=3.175 $Y2=0.18
r158 19 21 253.819 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=3.175 $Y=0.255
+ $X2=3.175 $Y2=0.75
r159 18 40 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=2.91 $Y=3.15 $X2=2.82
+ $Y2=3.15
r160 17 26 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.295 $Y=3.15
+ $X2=4.37 $Y2=3.075
r161 17 18 710.181 $w=1.5e-07 $l=1.385e-06 $layer=POLY_cond $X=4.295 $Y=3.15
+ $X2=2.91 $Y2=3.15
r162 14 16 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=2.82 $Y=2.675
+ $X2=2.82 $Y2=2.28
r163 13 40 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=2.82 $Y=3.075
+ $X2=2.82 $Y2=3.15
r164 12 14 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=2.82 $Y=2.765
+ $X2=2.82 $Y2=2.675
r165 12 13 120.5 $w=1.8e-07 $l=3.1e-07 $layer=POLY_cond $X=2.82 $Y=2.765
+ $X2=2.82 $Y2=3.075
r166 10 41 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.1 $Y=0.18
+ $X2=3.175 $Y2=0.18
r167 10 11 523.021 $w=1.5e-07 $l=1.02e-06 $layer=POLY_cond $X=3.1 $Y=0.18
+ $X2=2.08 $Y2=0.18
r168 9 38 7.1379 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=1.935 $Y=3.15 $X2=1.845
+ $Y2=3.15
r169 8 40 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=2.73 $Y=3.15 $X2=2.82
+ $Y2=3.15
r170 8 9 407.649 $w=1.5e-07 $l=7.95e-07 $layer=POLY_cond $X=2.73 $Y=3.15
+ $X2=1.935 $Y2=3.15
r171 4 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.005 $Y=0.255
+ $X2=2.08 $Y2=0.18
r172 4 6 253.819 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=2.005 $Y=0.255
+ $X2=2.005 $Y2=0.75
r173 1 38 109.045 $w=1.8e-07 $l=2.75e-07 $layer=POLY_cond $X=1.845 $Y=2.875
+ $X2=1.845 $Y2=3.15
r174 1 3 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=1.845 $Y=2.875
+ $X2=1.845 $Y2=2.38
.ends

.subckt PM_SKY130_FD_SC_HS__XOR3_1%A_1157_298# 1 2 7 9 12 15 16 17 19 22 25 30
+ 36 38
c85 22 0 1.49313e-19 $X=7.9 $Y=0.63
c86 12 0 1.40824e-19 $X=6.155 $Y=0.925
r87 35 36 8.73063 $w=3.28e-07 $l=2.5e-07 $layer=LI1_cond $X=7.65 $Y=2.36 $X2=7.9
+ $Y2=2.36
r88 32 35 4.53993 $w=3.28e-07 $l=1.3e-07 $layer=LI1_cond $X=7.52 $Y=2.36
+ $X2=7.65 $Y2=2.36
r89 27 30 5.56352 $w=2.88e-07 $l=1.4e-07 $layer=LI1_cond $X=5.97 $Y=1.675
+ $X2=6.11 $Y2=1.675
r90 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.97
+ $Y=1.655 $X2=5.97 $Y2=1.655
r91 25 36 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.9 $Y=2.195 $X2=7.9
+ $Y2=2.36
r92 25 38 87.0963 $w=1.68e-07 $l=1.335e-06 $layer=LI1_cond $X=7.9 $Y=2.195
+ $X2=7.9 $Y2=0.86
r93 20 38 6.94937 $w=2.48e-07 $l=1.25e-07 $layer=LI1_cond $X=7.94 $Y=0.735
+ $X2=7.94 $Y2=0.86
r94 20 22 4.84026 $w=2.48e-07 $l=1.05e-07 $layer=LI1_cond $X=7.94 $Y=0.735
+ $X2=7.94 $Y2=0.63
r95 18 32 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.52 $Y=2.525
+ $X2=7.52 $Y2=2.36
r96 18 19 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=7.52 $Y=2.525
+ $X2=7.52 $Y2=2.905
r97 16 19 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.435 $Y=2.99
+ $X2=7.52 $Y2=2.905
r98 16 17 80.8984 $w=1.68e-07 $l=1.24e-06 $layer=LI1_cond $X=7.435 $Y=2.99
+ $X2=6.195 $Y2=2.99
r99 15 17 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.11 $Y=2.905
+ $X2=6.195 $Y2=2.99
r100 14 30 3.86198 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=6.11 $Y=1.82
+ $X2=6.11 $Y2=1.675
r101 14 15 70.7861 $w=1.68e-07 $l=1.085e-06 $layer=LI1_cond $X=6.11 $Y=1.82
+ $X2=6.11 $Y2=2.905
r102 10 28 39.3952 $w=3.9e-07 $l=2.27255e-07 $layer=POLY_cond $X=6.155 $Y=1.49
+ $X2=6.007 $Y2=1.655
r103 10 12 289.713 $w=1.5e-07 $l=5.65e-07 $layer=POLY_cond $X=6.155 $Y=1.49
+ $X2=6.155 $Y2=0.925
r104 7 28 49.9004 $w=3.9e-07 $l=2.53476e-07 $layer=POLY_cond $X=6 $Y=1.905
+ $X2=6.007 $Y2=1.655
r105 7 9 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=6 $Y=1.905 $X2=6
+ $Y2=2.4
r106 2 35 600 $w=1.7e-07 $l=5.84423e-07 $layer=licon1_PDIFF $count=1 $X=7.455
+ $Y=1.865 $X2=7.65 $Y2=2.36
r107 1 22 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=7.755
+ $Y=0.42 $X2=7.9 $Y2=0.63
.ends

.subckt PM_SKY130_FD_SC_HS__XOR3_1%C 1 3 4 6 7 10 11 13 14 16 19 22
r75 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.04
+ $Y=1.52 $X2=7.04 $Y2=1.52
r76 24 26 11.9176 $w=3.64e-07 $l=9e-08 $layer=POLY_cond $X=6.935 $Y=1.43
+ $X2=6.935 $Y2=1.52
r77 22 27 7.85757 $w=3.28e-07 $l=2.25e-07 $layer=LI1_cond $X=7.04 $Y=1.295
+ $X2=7.04 $Y2=1.52
r78 17 19 105.117 $w=1.5e-07 $l=2.05e-07 $layer=POLY_cond $X=7.91 $Y=0.99
+ $X2=8.115 $Y2=0.99
r79 14 19 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=8.115 $Y=0.915
+ $X2=8.115 $Y2=0.99
r80 14 16 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=8.115 $Y=0.915
+ $X2=8.115 $Y2=0.63
r81 11 21 103.4 $w=1.69e-07 $l=3.6e-07 $layer=POLY_cond $X=7.925 $Y=1.79
+ $X2=7.925 $Y2=1.43
r82 11 13 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=7.925 $Y=1.79
+ $X2=7.925 $Y2=2.185
r83 10 21 22.1159 $w=1.69e-07 $l=8.21584e-08 $layer=POLY_cond $X=7.91 $Y=1.355
+ $X2=7.925 $Y2=1.43
r84 9 17 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.91 $Y=1.065
+ $X2=7.91 $Y2=0.99
r85 9 10 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=7.91 $Y=1.065
+ $X2=7.91 $Y2=1.355
r86 8 24 23.572 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=7.205 $Y=1.43
+ $X2=6.935 $Y2=1.43
r87 7 21 5.66465 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=7.835 $Y=1.43 $X2=7.925
+ $Y2=1.43
r88 7 8 323.043 $w=1.5e-07 $l=6.3e-07 $layer=POLY_cond $X=7.835 $Y=1.43
+ $X2=7.205 $Y2=1.43
r89 4 24 27.0487 $w=3.64e-07 $l=1.32288e-07 $layer=POLY_cond $X=6.835 $Y=1.355
+ $X2=6.935 $Y2=1.43
r90 4 6 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=6.835 $Y=1.355
+ $X2=6.835 $Y2=0.925
r91 1 26 68.0982 $w=3.64e-07 $l=4.66396e-07 $layer=POLY_cond $X=6.755 $Y=1.905
+ $X2=6.935 $Y2=1.52
r92 1 3 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=6.755 $Y=1.905
+ $X2=6.755 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_HS__XOR3_1%A_1215_396# 1 2 7 9 12 16 20 22 23 26 29 34
c77 12 0 1.49313e-19 $X=8.625 $Y=0.79
r78 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.42
+ $Y=1.515 $X2=8.42 $Y2=1.515
r79 29 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=1.665 $X2=8.4
+ $Y2=1.665
r80 26 39 6.77715 $w=3.38e-07 $l=1.15e-07 $layer=LI1_cond $X=6.535 $Y=1.665
+ $X2=6.535 $Y2=1.55
r81 25 26 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=1.665
+ $X2=6.48 $Y2=1.665
r82 23 25 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.625 $Y=1.665
+ $X2=6.48 $Y2=1.665
r83 22 29 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=8.255 $Y=1.665
+ $X2=8.4 $Y2=1.665
r84 22 23 2.01732 $w=1.4e-07 $l=1.63e-06 $layer=MET1_cond $X=8.255 $Y=1.665
+ $X2=6.625 $Y2=1.665
r85 20 39 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=6.62 $Y=1.1 $X2=6.62
+ $Y2=1.55
r86 14 26 1.86425 $w=3.38e-07 $l=5.5e-08 $layer=LI1_cond $X=6.535 $Y=1.72
+ $X2=6.535 $Y2=1.665
r87 14 16 13.7276 $w=3.38e-07 $l=4.05e-07 $layer=LI1_cond $X=6.535 $Y=1.72
+ $X2=6.535 $Y2=2.125
r88 10 33 39.4323 $w=3.92e-07 $l=2.26164e-07 $layer=POLY_cond $X=8.625 $Y=1.35
+ $X2=8.48 $Y2=1.515
r89 10 12 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=8.625 $Y=1.35
+ $X2=8.625 $Y2=0.79
r90 7 33 49.8838 $w=3.92e-07 $l=3.10242e-07 $layer=POLY_cond $X=8.615 $Y=1.765
+ $X2=8.48 $Y2=1.515
r91 7 9 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=8.615 $Y=1.765
+ $X2=8.615 $Y2=2.4
r92 2 16 300 $w=1.7e-07 $l=5.22494e-07 $layer=licon1_PDIFF $count=2 $X=6.075
+ $Y=1.98 $X2=6.53 $Y2=2.125
r93 1 20 182 $w=1.7e-07 $l=6.61872e-07 $layer=licon1_NDIFF $count=1 $X=6.23
+ $Y=0.605 $X2=6.62 $Y2=1.1
.ends

.subckt PM_SKY130_FD_SC_HS__XOR3_1%A_27_134# 1 2 3 4 13 14 17 20 21 22 25 29 32
+ 35 37 38 40 41
r85 37 38 9.60999 $w=5.13e-07 $l=1.65e-07 $layer=LI1_cond $X=0.342 $Y=2.425
+ $X2=0.342 $Y2=2.26
r86 35 38 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.17 $Y=1.3 $X2=0.17
+ $Y2=2.26
r87 32 40 3.70735 $w=2.5e-07 $l=1.18427e-07 $layer=LI1_cond $X=2.675 $Y=1.26
+ $X2=2.595 $Y2=1.345
r88 32 41 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=2.675 $Y=1.26
+ $X2=2.675 $Y2=1.09
r89 27 41 7.14225 $w=2.58e-07 $l=1.3e-07 $layer=LI1_cond $X=2.72 $Y=0.96
+ $X2=2.72 $Y2=1.09
r90 27 29 4.43247 $w=2.58e-07 $l=1e-07 $layer=LI1_cond $X=2.72 $Y=0.96 $X2=2.72
+ $Y2=0.86
r91 23 40 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.595 $Y=1.43
+ $X2=2.595 $Y2=1.345
r92 23 25 27.0649 $w=3.28e-07 $l=7.75e-07 $layer=LI1_cond $X=2.595 $Y=1.43
+ $X2=2.595 $Y2=2.205
r93 21 40 2.76166 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.43 $Y=1.345
+ $X2=2.595 $Y2=1.345
r94 21 22 30.3369 $w=1.68e-07 $l=4.65e-07 $layer=LI1_cond $X=2.43 $Y=1.345
+ $X2=1.965 $Y2=1.345
r95 20 22 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.88 $Y=1.26
+ $X2=1.965 $Y2=1.345
r96 19 20 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=1.88 $Y=0.83
+ $X2=1.88 $Y2=1.26
r97 18 34 5.39736 $w=1.7e-07 $l=1.82483e-07 $layer=LI1_cond $X=0.445 $Y=0.745
+ $X2=0.265 $Y2=0.74
r98 17 19 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.795 $Y=0.745
+ $X2=1.88 $Y2=0.83
r99 17 18 88.0749 $w=1.68e-07 $l=1.35e-06 $layer=LI1_cond $X=1.795 $Y=0.745
+ $X2=0.445 $Y2=0.745
r100 14 35 8.99121 $w=3.58e-07 $l=1.8e-07 $layer=LI1_cond $X=0.265 $Y=1.12
+ $X2=0.265 $Y2=1.3
r101 13 34 2.62574 $w=3.6e-07 $l=9e-08 $layer=LI1_cond $X=0.265 $Y=0.83
+ $X2=0.265 $Y2=0.74
r102 13 14 9.28357 $w=3.58e-07 $l=2.9e-07 $layer=LI1_cond $X=0.265 $Y=0.83
+ $X2=0.265 $Y2=1.12
r103 4 25 600 $w=1.7e-07 $l=3.18865e-07 $layer=licon1_PDIFF $count=1 $X=2.425
+ $Y=1.96 $X2=2.595 $Y2=2.205
r104 3 37 300 $w=1.7e-07 $l=5.32588e-07 $layer=licon1_PDIFF $count=2 $X=0.29
+ $Y=1.96 $X2=0.435 $Y2=2.425
r105 2 29 182 $w=1.7e-07 $l=2.8801e-07 $layer=licon1_NDIFF $count=1 $X=2.58
+ $Y=0.65 $X2=2.765 $Y2=0.86
r106 1 34 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.67 $X2=0.28 $Y2=0.815
.ends

.subckt PM_SKY130_FD_SC_HS__XOR3_1%VPWR 1 2 3 12 16 22 27 28 29 35 42 52 53 56
+ 59
r74 59 60 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=3.33 $X2=8.4
+ $Y2=3.33
r75 56 57 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r76 53 60 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=3.33
+ $X2=8.4 $Y2=3.33
r77 52 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r78 50 59 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.555 $Y=3.33
+ $X2=8.39 $Y2=3.33
r79 50 52 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=8.555 $Y=3.33
+ $X2=8.88 $Y2=3.33
r80 49 60 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=3.33
+ $X2=8.4 $Y2=3.33
r81 48 49 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r82 46 49 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=7.92 $Y2=3.33
r83 46 57 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=5.04 $Y2=3.33
r84 45 48 156.578 $w=1.68e-07 $l=2.4e-06 $layer=LI1_cond $X=5.52 $Y=3.33
+ $X2=7.92 $Y2=3.33
r85 45 46 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r86 43 56 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.2 $Y=3.33
+ $X2=5.075 $Y2=3.33
r87 43 45 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=5.2 $Y=3.33 $X2=5.52
+ $Y2=3.33
r88 42 59 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.225 $Y=3.33
+ $X2=8.39 $Y2=3.33
r89 42 48 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=8.225 $Y=3.33
+ $X2=7.92 $Y2=3.33
r90 37 40 219.209 $w=1.68e-07 $l=3.36e-06 $layer=LI1_cond $X=1.2 $Y=3.33
+ $X2=4.56 $Y2=3.33
r91 37 38 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r92 35 56 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.95 $Y=3.33
+ $X2=5.075 $Y2=3.33
r93 35 40 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=4.95 $Y=3.33
+ $X2=4.56 $Y2=3.33
r94 33 38 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r95 32 33 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r96 29 57 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=5.04 $Y2=3.33
r97 29 38 0.936549 $w=4.9e-07 $l=3.36e-06 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=1.2 $Y2=3.33
r98 29 40 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r99 27 32 3.26203 $w=1.68e-07 $l=5e-08 $layer=LI1_cond $X=0.77 $Y=3.33 $X2=0.72
+ $Y2=3.33
r100 27 28 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.77 $Y=3.33
+ $X2=0.935 $Y2=3.33
r101 26 37 6.52406 $w=1.68e-07 $l=1e-07 $layer=LI1_cond $X=1.1 $Y=3.33 $X2=1.2
+ $Y2=3.33
r102 26 28 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.1 $Y=3.33
+ $X2=0.935 $Y2=3.33
r103 22 25 12.2229 $w=3.28e-07 $l=3.5e-07 $layer=LI1_cond $X=8.39 $Y=2.115
+ $X2=8.39 $Y2=2.465
r104 20 59 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.39 $Y=3.245
+ $X2=8.39 $Y2=3.33
r105 20 25 27.2396 $w=3.28e-07 $l=7.8e-07 $layer=LI1_cond $X=8.39 $Y=3.245
+ $X2=8.39 $Y2=2.465
r106 16 19 32.2684 $w=2.48e-07 $l=7e-07 $layer=LI1_cond $X=5.075 $Y=2.115
+ $X2=5.075 $Y2=2.815
r107 14 56 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.075 $Y=3.245
+ $X2=5.075 $Y2=3.33
r108 14 19 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=5.075 $Y=3.245
+ $X2=5.075 $Y2=2.815
r109 10 28 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.935 $Y=3.245
+ $X2=0.935 $Y2=3.33
r110 10 12 28.6365 $w=3.28e-07 $l=8.2e-07 $layer=LI1_cond $X=0.935 $Y=3.245
+ $X2=0.935 $Y2=2.425
r111 3 25 300 $w=1.7e-07 $l=7.70714e-07 $layer=licon1_PDIFF $count=2 $X=8
+ $Y=1.865 $X2=8.39 $Y2=2.465
r112 3 22 600 $w=1.7e-07 $l=4.996e-07 $layer=licon1_PDIFF $count=1 $X=8 $Y=1.865
+ $X2=8.39 $Y2=2.115
r113 2 19 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=4.965
+ $Y=1.84 $X2=5.115 $Y2=2.815
r114 2 16 400 $w=1.7e-07 $l=3.4187e-07 $layer=licon1_PDIFF $count=1 $X=4.965
+ $Y=1.84 $X2=5.115 $Y2=2.115
r115 1 12 300 $w=1.7e-07 $l=5.5608e-07 $layer=licon1_PDIFF $count=2 $X=0.735
+ $Y=1.96 $X2=0.935 $Y2=2.425
.ends

.subckt PM_SKY130_FD_SC_HS__XOR3_1%A_384_392# 1 2 3 4 15 17 18 22 23 24 26 27 28
+ 32 33 34 37 39 40 42
c125 15 0 1.79271e-19 $X=2.095 $Y=2.105
r126 41 42 93.2941 $w=1.68e-07 $l=1.43e-06 $layer=LI1_cond $X=7.56 $Y=0.425
+ $X2=7.56 $Y2=1.855
r127 39 42 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.475 $Y=1.94
+ $X2=7.56 $Y2=1.855
r128 39 40 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=7.475 $Y=1.94
+ $X2=7.205 $Y2=1.94
r129 35 40 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=7.04 $Y=2.025
+ $X2=7.205 $Y2=1.94
r130 35 37 3.49225 $w=3.28e-07 $l=1e-07 $layer=LI1_cond $X=7.04 $Y=2.025
+ $X2=7.04 $Y2=2.125
r131 33 41 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.475 $Y=0.34
+ $X2=7.56 $Y2=0.425
r132 33 34 94.5989 $w=1.68e-07 $l=1.45e-06 $layer=LI1_cond $X=7.475 $Y=0.34
+ $X2=6.025 $Y2=0.34
r133 30 32 2.30489 $w=2.48e-07 $l=5e-08 $layer=LI1_cond $X=5.9 $Y=0.85 $X2=5.9
+ $Y2=0.8
r134 29 34 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=5.9 $Y=0.425
+ $X2=6.025 $Y2=0.34
r135 29 32 17.2866 $w=2.48e-07 $l=3.75e-07 $layer=LI1_cond $X=5.9 $Y=0.425
+ $X2=5.9 $Y2=0.8
r136 27 30 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=5.775 $Y=0.935
+ $X2=5.9 $Y2=0.85
r137 27 28 41.1016 $w=1.68e-07 $l=6.3e-07 $layer=LI1_cond $X=5.775 $Y=0.935
+ $X2=5.145 $Y2=0.935
r138 26 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.06 $Y=0.85
+ $X2=5.145 $Y2=0.935
r139 25 26 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=5.06 $Y=0.425
+ $X2=5.06 $Y2=0.85
r140 23 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.975 $Y=0.34
+ $X2=5.06 $Y2=0.425
r141 23 24 92.6417 $w=1.68e-07 $l=1.42e-06 $layer=LI1_cond $X=4.975 $Y=0.34
+ $X2=3.555 $Y2=0.34
r142 20 22 129.829 $w=1.68e-07 $l=1.99e-06 $layer=LI1_cond $X=3.47 $Y=2.565
+ $X2=3.47 $Y2=0.575
r143 19 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.47 $Y=0.425
+ $X2=3.555 $Y2=0.34
r144 19 22 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=3.47 $Y=0.425
+ $X2=3.47 $Y2=0.575
r145 17 20 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.385 $Y=2.65
+ $X2=3.47 $Y2=2.565
r146 17 18 73.3957 $w=1.68e-07 $l=1.125e-06 $layer=LI1_cond $X=3.385 $Y=2.65
+ $X2=2.26 $Y2=2.65
r147 13 18 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.095 $Y=2.565
+ $X2=2.26 $Y2=2.65
r148 13 15 16.0644 $w=3.28e-07 $l=4.6e-07 $layer=LI1_cond $X=2.095 $Y=2.565
+ $X2=2.095 $Y2=2.105
r149 4 37 300 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_PDIFF $count=2 $X=6.83
+ $Y=1.98 $X2=7.04 $Y2=2.125
r150 3 15 300 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=2 $X=1.92
+ $Y=1.96 $X2=2.095 $Y2=2.105
r151 2 32 182 $w=1.7e-07 $l=2.53673e-07 $layer=licon1_NDIFF $count=1 $X=5.805
+ $Y=0.605 $X2=5.94 $Y2=0.8
r152 1 22 91 $w=1.7e-07 $l=2.83373e-07 $layer=licon1_NDIFF $count=2 $X=3.25
+ $Y=0.43 $X2=3.47 $Y2=0.575
.ends

.subckt PM_SKY130_FD_SC_HS__XOR3_1%A_416_86# 1 2 3 4 15 19 20 21 23 27 28 30 32
+ 38 41 42 44 45 48 51 52
c128 45 0 1.96802e-19 $X=3.265 $Y=1.665
c129 41 0 1.40824e-19 $X=7.095 $Y=0.76
c130 15 0 1.59849e-19 $X=2.22 $Y=0.575
r131 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=1.665
+ $X2=5.52 $Y2=1.665
r132 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=1.665
+ $X2=3.12 $Y2=1.665
r133 45 47 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.265 $Y=1.665
+ $X2=3.12 $Y2=1.665
r134 44 51 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.375 $Y=1.665
+ $X2=5.52 $Y2=1.665
r135 44 45 2.61138 $w=1.4e-07 $l=2.11e-06 $layer=MET1_cond $X=5.375 $Y=1.665
+ $X2=3.265 $Y2=1.665
r136 41 42 10.0337 $w=3.28e-07 $l=2.1e-07 $layer=LI1_cond $X=7.095 $Y=0.76
+ $X2=6.885 $Y2=0.76
r137 39 52 16.5011 $w=2.03e-07 $l=3.05e-07 $layer=LI1_cond $X=5.522 $Y=1.36
+ $X2=5.522 $Y2=1.665
r138 36 52 15.4191 $w=2.03e-07 $l=2.85e-07 $layer=LI1_cond $X=5.522 $Y=1.95
+ $X2=5.522 $Y2=1.665
r139 36 38 8.27032 $w=4.15e-07 $l=2.22542e-07 $layer=LI1_cond $X=5.522 $Y=1.95
+ $X2=5.63 $Y2=2.125
r140 35 48 68.5361 $w=1.93e-07 $l=1.205e-06 $layer=LI1_cond $X=3.117 $Y=0.46
+ $X2=3.117 $Y2=1.665
r141 34 48 11.9441 $w=1.93e-07 $l=2.1e-07 $layer=LI1_cond $X=3.117 $Y=1.875
+ $X2=3.117 $Y2=1.665
r142 32 42 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=6.365 $Y=0.68
+ $X2=6.885 $Y2=0.68
r143 29 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.28 $Y=0.765
+ $X2=6.365 $Y2=0.68
r144 29 30 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=6.28 $Y=0.765
+ $X2=6.28 $Y2=1.19
r145 28 39 6.89401 $w=1.7e-07 $l=1.39155e-07 $layer=LI1_cond $X=5.625 $Y=1.275
+ $X2=5.522 $Y2=1.36
r146 27 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.195 $Y=1.275
+ $X2=6.28 $Y2=1.19
r147 27 28 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=6.195 $Y=1.275
+ $X2=5.625 $Y2=1.275
r148 21 34 6.35106 $w=2.48e-07 $l=1.25e-07 $layer=LI1_cond $X=3.09 $Y=2 $X2=3.09
+ $Y2=1.875
r149 21 23 6.22319 $w=2.48e-07 $l=1.35e-07 $layer=LI1_cond $X=3.09 $Y=2 $X2=3.09
+ $Y2=2.135
r150 19 35 6.85817 $w=1.7e-07 $l=1.32868e-07 $layer=LI1_cond $X=3.02 $Y=0.375
+ $X2=3.117 $Y2=0.46
r151 19 20 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=3.02 $Y=0.375
+ $X2=2.385 $Y2=0.375
r152 15 17 16.1342 $w=2.48e-07 $l=3.5e-07 $layer=LI1_cond $X=2.26 $Y=0.575
+ $X2=2.26 $Y2=0.925
r153 13 20 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=2.26 $Y=0.46
+ $X2=2.385 $Y2=0.375
r154 13 15 5.30124 $w=2.48e-07 $l=1.15e-07 $layer=LI1_cond $X=2.26 $Y=0.46
+ $X2=2.26 $Y2=0.575
r155 4 38 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=5.545
+ $Y=1.98 $X2=5.69 $Y2=2.125
r156 3 23 600 $w=1.7e-07 $l=3.10403e-07 $layer=licon1_PDIFF $count=1 $X=2.895
+ $Y=1.96 $X2=3.13 $Y2=2.135
r157 2 41 182 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=1 $X=6.91
+ $Y=0.605 $X2=7.095 $Y2=0.76
r158 1 17 182 $w=1.7e-07 $l=5.60647e-07 $layer=licon1_NDIFF $count=1 $X=2.08
+ $Y=0.43 $X2=2.22 $Y2=0.925
r159 1 15 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=2.08
+ $Y=0.43 $X2=2.22 $Y2=0.575
.ends

.subckt PM_SKY130_FD_SC_HS__XOR3_1%X 1 2 7 8 9 10 11 12 13
r12 12 13 17.0562 $w=2.48e-07 $l=3.7e-07 $layer=LI1_cond $X=8.88 $Y=2.405
+ $X2=8.88 $Y2=2.775
r13 11 12 19.361 $w=2.48e-07 $l=4.2e-07 $layer=LI1_cond $X=8.88 $Y=1.985
+ $X2=8.88 $Y2=2.405
r14 10 11 14.7513 $w=2.48e-07 $l=3.2e-07 $layer=LI1_cond $X=8.88 $Y=1.665
+ $X2=8.88 $Y2=1.985
r15 9 10 17.0562 $w=2.48e-07 $l=3.7e-07 $layer=LI1_cond $X=8.88 $Y=1.295
+ $X2=8.88 $Y2=1.665
r16 8 9 17.0562 $w=2.48e-07 $l=3.7e-07 $layer=LI1_cond $X=8.88 $Y=0.925 $X2=8.88
+ $Y2=1.295
r17 7 8 17.0562 $w=2.48e-07 $l=3.7e-07 $layer=LI1_cond $X=8.88 $Y=0.555 $X2=8.88
+ $Y2=0.925
r18 2 13 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=8.69
+ $Y=1.84 $X2=8.84 $Y2=2.815
r19 2 11 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=8.69
+ $Y=1.84 $X2=8.84 $Y2=1.985
r20 1 7 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=8.7 $Y=0.42
+ $X2=8.84 $Y2=0.565
.ends

.subckt PM_SKY130_FD_SC_HS__XOR3_1%VGND 1 2 3 12 16 20 27 35 42 43 48 51 53 56
r71 56 57 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r72 53 54 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r73 50 51 12.4896 $w=5.73e-07 $l=2.85e-07 $layer=LI1_cond $X=0.91 $Y=0.202
+ $X2=1.195 $Y2=0.202
r74 46 50 3.95226 $w=5.73e-07 $l=1.9e-07 $layer=LI1_cond $X=0.72 $Y=0.202
+ $X2=0.91 $Y2=0.202
r75 46 48 8.53733 $w=5.73e-07 $l=9.5e-08 $layer=LI1_cond $X=0.72 $Y=0.202
+ $X2=0.625 $Y2=0.202
r76 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r77 43 57 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=0 $X2=8.4
+ $Y2=0
r78 42 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=0 $X2=8.88
+ $Y2=0
r79 40 56 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.575 $Y=0 $X2=8.41
+ $Y2=0
r80 40 42 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=8.575 $Y=0 $X2=8.88
+ $Y2=0
r81 39 57 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=0 $X2=8.4
+ $Y2=0
r82 39 54 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=7.92 $Y=0 $X2=5.52
+ $Y2=0
r83 38 39 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=7.92 $Y=0 $X2=7.92
+ $Y2=0
r84 36 53 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.565 $Y=0 $X2=5.44
+ $Y2=0
r85 36 38 153.642 $w=1.68e-07 $l=2.355e-06 $layer=LI1_cond $X=5.565 $Y=0
+ $X2=7.92 $Y2=0
r86 35 56 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.245 $Y=0 $X2=8.41
+ $Y2=0
r87 35 38 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=8.245 $Y=0 $X2=7.92
+ $Y2=0
r88 34 54 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=5.52
+ $Y2=0
r89 33 34 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=5.04 $Y=0
+ $X2=5.04 $Y2=0
r90 31 47 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r91 30 33 250.524 $w=1.68e-07 $l=3.84e-06 $layer=LI1_cond $X=1.2 $Y=0 $X2=5.04
+ $Y2=0
r92 30 51 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=1.2 $Y=0 $X2=1.195
+ $Y2=0
r93 30 31 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=1.2 $Y=0
+ $X2=1.2 $Y2=0
r94 27 53 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.315 $Y=0 $X2=5.44
+ $Y2=0
r95 27 33 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=5.315 $Y=0 $X2=5.04
+ $Y2=0
r96 25 47 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r97 24 48 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=0.24 $Y=0 $X2=0.625
+ $Y2=0
r98 24 25 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r99 20 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=5.04
+ $Y2=0
r100 20 31 0.936549 $w=4.9e-07 $l=3.36e-06 $layer=MET1_cond $X=4.56 $Y=0 $X2=1.2
+ $Y2=0
r101 16 18 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=8.41 $Y=0.565
+ $X2=8.41 $Y2=1.015
r102 14 56 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.41 $Y=0.085
+ $X2=8.41 $Y2=0
r103 14 16 16.7628 $w=3.28e-07 $l=4.8e-07 $layer=LI1_cond $X=8.41 $Y=0.085
+ $X2=8.41 $Y2=0.565
r104 10 53 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.44 $Y=0.085
+ $X2=5.44 $Y2=0
r105 10 12 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=5.44 $Y=0.085
+ $X2=5.44 $Y2=0.515
r106 3 18 182 $w=1.7e-07 $l=6.96366e-07 $layer=licon1_NDIFF $count=1 $X=8.19
+ $Y=0.42 $X2=8.41 $Y2=1.015
r107 3 16 182 $w=1.7e-07 $l=2.83373e-07 $layer=licon1_NDIFF $count=1 $X=8.19
+ $Y=0.42 $X2=8.41 $Y2=0.565
r108 2 12 182 $w=1.7e-07 $l=4.56782e-07 $layer=licon1_NDIFF $count=1 $X=5.01
+ $Y=0.37 $X2=5.4 $Y2=0.515
r109 1 50 182 $w=1.7e-07 $l=4.86133e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.67 $X2=0.91 $Y2=0.325
.ends

