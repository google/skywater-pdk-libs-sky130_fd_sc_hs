* File: sky130_fd_sc_hs__buf_16.pxi.spice
* Created: Tue Sep  1 19:56:37 2020
* 
x_PM_SKY130_FD_SC_HS__BUF_16%A_83_260# N_A_83_260#_M1002_d N_A_83_260#_M1011_d
+ N_A_83_260#_M1013_d N_A_83_260#_M1000_d N_A_83_260#_M1028_d
+ N_A_83_260#_M1036_d N_A_83_260#_c_216_n N_A_83_260#_M1001_g
+ N_A_83_260#_M1003_g N_A_83_260#_M1004_g N_A_83_260#_c_217_n
+ N_A_83_260#_M1007_g N_A_83_260#_M1008_g N_A_83_260#_c_218_n
+ N_A_83_260#_M1015_g N_A_83_260#_M1009_g N_A_83_260#_c_219_n
+ N_A_83_260#_M1017_g N_A_83_260#_M1010_g N_A_83_260#_c_220_n
+ N_A_83_260#_M1018_g N_A_83_260#_M1014_g N_A_83_260#_c_221_n
+ N_A_83_260#_M1020_g N_A_83_260#_M1016_g N_A_83_260#_c_222_n
+ N_A_83_260#_M1021_g N_A_83_260#_M1019_g N_A_83_260#_c_223_n
+ N_A_83_260#_M1022_g N_A_83_260#_M1023_g N_A_83_260#_c_224_n
+ N_A_83_260#_M1025_g N_A_83_260#_M1024_g N_A_83_260#_c_225_n
+ N_A_83_260#_M1026_g N_A_83_260#_M1032_g N_A_83_260#_c_226_n
+ N_A_83_260#_M1027_g N_A_83_260#_M1034_g N_A_83_260#_c_227_n
+ N_A_83_260#_M1029_g N_A_83_260#_M1035_g N_A_83_260#_c_228_n
+ N_A_83_260#_M1030_g N_A_83_260#_M1038_g N_A_83_260#_c_229_n
+ N_A_83_260#_M1033_g N_A_83_260#_c_230_n N_A_83_260#_M1037_g
+ N_A_83_260#_M1041_g N_A_83_260#_c_231_n N_A_83_260#_M1040_g
+ N_A_83_260#_M1042_g N_A_83_260#_c_198_n N_A_83_260#_c_418_p
+ N_A_83_260#_c_246_p N_A_83_260#_c_311_p N_A_83_260#_c_232_n
+ N_A_83_260#_c_199_n N_A_83_260#_c_200_n N_A_83_260#_c_258_p
+ N_A_83_260#_c_233_n N_A_83_260#_c_201_n N_A_83_260#_c_202_n
+ N_A_83_260#_c_270_p N_A_83_260#_c_277_p N_A_83_260#_c_234_n
+ N_A_83_260#_c_203_n N_A_83_260#_c_248_p N_A_83_260#_c_204_n
+ N_A_83_260#_c_266_p N_A_83_260#_c_205_n N_A_83_260#_c_206_n
+ N_A_83_260#_c_207_n N_A_83_260#_c_208_n N_A_83_260#_c_209_n
+ N_A_83_260#_c_210_n N_A_83_260#_c_211_n N_A_83_260#_c_212_n
+ N_A_83_260#_c_213_n N_A_83_260#_c_214_n N_A_83_260#_c_215_n
+ PM_SKY130_FD_SC_HS__BUF_16%A_83_260#
x_PM_SKY130_FD_SC_HS__BUF_16%A N_A_c_647_n N_A_M1000_g N_A_M1002_g N_A_M1005_g
+ N_A_c_648_n N_A_M1006_g N_A_M1011_g N_A_c_649_n N_A_M1028_g N_A_M1012_g
+ N_A_c_650_n N_A_M1031_g N_A_M1013_g N_A_c_651_n N_A_M1036_g N_A_c_652_n
+ N_A_M1039_g N_A_M1043_g A A A A A N_A_c_646_n PM_SKY130_FD_SC_HS__BUF_16%A
x_PM_SKY130_FD_SC_HS__BUF_16%VPWR N_VPWR_M1001_d N_VPWR_M1007_d N_VPWR_M1017_d
+ N_VPWR_M1020_d N_VPWR_M1022_d N_VPWR_M1026_d N_VPWR_M1029_d N_VPWR_M1033_d
+ N_VPWR_M1040_d N_VPWR_M1006_s N_VPWR_M1031_s N_VPWR_M1039_s N_VPWR_c_765_n
+ N_VPWR_c_766_n N_VPWR_c_767_n N_VPWR_c_768_n N_VPWR_c_769_n N_VPWR_c_770_n
+ N_VPWR_c_771_n N_VPWR_c_772_n N_VPWR_c_773_n N_VPWR_c_774_n N_VPWR_c_775_n
+ N_VPWR_c_776_n N_VPWR_c_777_n N_VPWR_c_778_n N_VPWR_c_779_n N_VPWR_c_780_n
+ N_VPWR_c_781_n N_VPWR_c_782_n N_VPWR_c_783_n N_VPWR_c_784_n N_VPWR_c_785_n
+ N_VPWR_c_786_n N_VPWR_c_787_n N_VPWR_c_788_n N_VPWR_c_789_n N_VPWR_c_790_n
+ N_VPWR_c_791_n N_VPWR_c_792_n N_VPWR_c_793_n N_VPWR_c_794_n N_VPWR_c_795_n
+ N_VPWR_c_796_n VPWR N_VPWR_c_797_n N_VPWR_c_798_n N_VPWR_c_799_n
+ N_VPWR_c_764_n PM_SKY130_FD_SC_HS__BUF_16%VPWR
x_PM_SKY130_FD_SC_HS__BUF_16%X N_X_M1003_d N_X_M1008_d N_X_M1010_d N_X_M1016_d
+ N_X_M1023_d N_X_M1032_d N_X_M1035_d N_X_M1041_d N_X_M1001_s N_X_M1015_s
+ N_X_M1018_s N_X_M1021_s N_X_M1025_s N_X_M1027_s N_X_M1030_s N_X_M1037_s
+ N_X_c_954_n N_X_c_955_n N_X_c_956_n N_X_c_971_n N_X_c_957_n N_X_c_958_n
+ N_X_c_959_n N_X_c_960_n N_X_c_961_n N_X_c_962_n N_X_c_972_n N_X_c_963_n
+ N_X_c_964_n N_X_c_965_n N_X_c_966_n X N_X_c_967_n N_X_c_968_n N_X_c_976_n
+ N_X_c_977_n N_X_c_978_n N_X_c_969_n N_X_c_980_n N_X_c_1091_n N_X_c_1118_n
+ N_X_c_970_n PM_SKY130_FD_SC_HS__BUF_16%X
x_PM_SKY130_FD_SC_HS__BUF_16%VGND N_VGND_M1003_s N_VGND_M1004_s N_VGND_M1009_s
+ N_VGND_M1014_s N_VGND_M1019_s N_VGND_M1024_s N_VGND_M1034_s N_VGND_M1038_s
+ N_VGND_M1042_s N_VGND_M1005_s N_VGND_M1012_s N_VGND_M1043_s N_VGND_c_1213_n
+ N_VGND_c_1214_n N_VGND_c_1215_n N_VGND_c_1216_n N_VGND_c_1217_n
+ N_VGND_c_1218_n N_VGND_c_1219_n N_VGND_c_1220_n N_VGND_c_1221_n
+ N_VGND_c_1222_n N_VGND_c_1223_n N_VGND_c_1224_n N_VGND_c_1225_n
+ N_VGND_c_1226_n N_VGND_c_1227_n N_VGND_c_1228_n N_VGND_c_1229_n
+ N_VGND_c_1230_n N_VGND_c_1231_n N_VGND_c_1232_n N_VGND_c_1233_n
+ N_VGND_c_1234_n N_VGND_c_1235_n N_VGND_c_1236_n N_VGND_c_1237_n VGND
+ N_VGND_c_1238_n N_VGND_c_1239_n N_VGND_c_1240_n N_VGND_c_1241_n
+ N_VGND_c_1242_n N_VGND_c_1243_n N_VGND_c_1244_n N_VGND_c_1245_n
+ N_VGND_c_1246_n N_VGND_c_1247_n N_VGND_c_1248_n
+ PM_SKY130_FD_SC_HS__BUF_16%VGND
cc_1 VNB N_A_83_260#_M1003_g 0.026031f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=0.74
cc_2 VNB N_A_83_260#_M1004_g 0.0204008f $X=-0.19 $Y=-0.245 $X2=0.94 $Y2=0.74
cc_3 VNB N_A_83_260#_M1008_g 0.0211569f $X=-0.19 $Y=-0.245 $X2=1.37 $Y2=0.74
cc_4 VNB N_A_83_260#_M1009_g 0.0211559f $X=-0.19 $Y=-0.245 $X2=1.8 $Y2=0.74
cc_5 VNB N_A_83_260#_M1010_g 0.0211579f $X=-0.19 $Y=-0.245 $X2=2.23 $Y2=0.74
cc_6 VNB N_A_83_260#_M1014_g 0.0203176f $X=-0.19 $Y=-0.245 $X2=2.66 $Y2=0.74
cc_7 VNB N_A_83_260#_M1016_g 0.0211668f $X=-0.19 $Y=-0.245 $X2=3.09 $Y2=0.74
cc_8 VNB N_A_83_260#_M1019_g 0.0203111f $X=-0.19 $Y=-0.245 $X2=3.52 $Y2=0.74
cc_9 VNB N_A_83_260#_M1023_g 0.0209859f $X=-0.19 $Y=-0.245 $X2=3.95 $Y2=0.74
cc_10 VNB N_A_83_260#_M1024_g 0.0219226f $X=-0.19 $Y=-0.245 $X2=4.38 $Y2=0.74
cc_11 VNB N_A_83_260#_M1032_g 0.022768f $X=-0.19 $Y=-0.245 $X2=4.95 $Y2=0.74
cc_12 VNB N_A_83_260#_M1034_g 0.0219411f $X=-0.19 $Y=-0.245 $X2=5.38 $Y2=0.74
cc_13 VNB N_A_83_260#_M1035_g 0.0225962f $X=-0.19 $Y=-0.245 $X2=5.95 $Y2=0.74
cc_14 VNB N_A_83_260#_M1038_g 0.0219225f $X=-0.19 $Y=-0.245 $X2=6.38 $Y2=0.74
cc_15 VNB N_A_83_260#_M1041_g 0.0219204f $X=-0.19 $Y=-0.245 $X2=6.95 $Y2=0.74
cc_16 VNB N_A_83_260#_M1042_g 0.0197121f $X=-0.19 $Y=-0.245 $X2=7.38 $Y2=0.74
cc_17 VNB N_A_83_260#_c_198_n 0.00373179f $X=-0.19 $Y=-0.245 $X2=7.94 $Y2=1.095
cc_18 VNB N_A_83_260#_c_199_n 0.00178908f $X=-0.19 $Y=-0.245 $X2=8.025 $Y2=0.515
cc_19 VNB N_A_83_260#_c_200_n 0.00324651f $X=-0.19 $Y=-0.245 $X2=8.8 $Y2=1.095
cc_20 VNB N_A_83_260#_c_201_n 0.00178908f $X=-0.19 $Y=-0.245 $X2=8.885 $Y2=0.515
cc_21 VNB N_A_83_260#_c_202_n 0.00616262f $X=-0.19 $Y=-0.245 $X2=9.695 $Y2=1.095
cc_22 VNB N_A_83_260#_c_203_n 0.00253445f $X=-0.19 $Y=-0.245 $X2=9.78 $Y2=0.515
cc_23 VNB N_A_83_260#_c_204_n 0.00127131f $X=-0.19 $Y=-0.245 $X2=8.025 $Y2=1.095
cc_24 VNB N_A_83_260#_c_205_n 0.00127131f $X=-0.19 $Y=-0.245 $X2=8.885 $Y2=1.095
cc_25 VNB N_A_83_260#_c_206_n 0.00137782f $X=-0.19 $Y=-0.245 $X2=7.505 $Y2=1.665
cc_26 VNB N_A_83_260#_c_207_n 0.00330716f $X=-0.19 $Y=-0.245 $X2=7.505 $Y2=1.665
cc_27 VNB N_A_83_260#_c_208_n 0.00103434f $X=-0.19 $Y=-0.245 $X2=1.15 $Y2=1.465
cc_28 VNB N_A_83_260#_c_209_n 0.00107044f $X=-0.19 $Y=-0.245 $X2=2.035 $Y2=1.465
cc_29 VNB N_A_83_260#_c_210_n 0.00100002f $X=-0.19 $Y=-0.245 $X2=2.995 $Y2=1.465
cc_30 VNB N_A_83_260#_c_211_n 0.00103148f $X=-0.19 $Y=-0.245 $X2=3.86 $Y2=1.465
cc_31 VNB N_A_83_260#_c_212_n 0.00227452f $X=-0.19 $Y=-0.245 $X2=4.72 $Y2=1.465
cc_32 VNB N_A_83_260#_c_213_n 0.0022469f $X=-0.19 $Y=-0.245 $X2=5.74 $Y2=1.465
cc_33 VNB N_A_83_260#_c_214_n 0.00233862f $X=-0.19 $Y=-0.245 $X2=6.665 $Y2=1.465
cc_34 VNB N_A_83_260#_c_215_n 0.470668f $X=-0.19 $Y=-0.245 $X2=7.305 $Y2=1.532
cc_35 VNB N_A_M1002_g 0.0227257f $X=-0.19 $Y=-0.245 $X2=9.68 $Y2=1.84
cc_36 VNB N_A_M1005_g 0.0224687f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_M1011_g 0.0224899f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_M1012_g 0.0230063f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=0.74
cc_39 VNB N_A_M1013_g 0.0246689f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=2.4
cc_40 VNB N_A_M1043_g 0.0327497f $X=-0.19 $Y=-0.245 $X2=1.8 $Y2=0.74
cc_41 VNB A 0.0168057f $X=-0.19 $Y=-0.245 $X2=2.23 $Y2=1.3
cc_42 VNB N_A_c_646_n 0.109956f $X=-0.19 $Y=-0.245 $X2=3.52 $Y2=0.74
cc_43 VNB N_VPWR_c_764_n 0.442315f $X=-0.19 $Y=-0.245 $X2=8.93 $Y2=2.115
cc_44 VNB N_X_c_954_n 0.00281054f $X=-0.19 $Y=-0.245 $X2=2.355 $Y2=1.765
cc_45 VNB N_X_c_955_n 0.00208122f $X=-0.19 $Y=-0.245 $X2=2.66 $Y2=0.74
cc_46 VNB N_X_c_956_n 0.00240191f $X=-0.19 $Y=-0.245 $X2=3.09 $Y2=1.3
cc_47 VNB N_X_c_957_n 0.00326079f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_X_c_958_n 0.00240191f $X=-0.19 $Y=-0.245 $X2=3.95 $Y2=1.3
cc_49 VNB N_X_c_959_n 0.00108974f $X=-0.19 $Y=-0.245 $X2=3.95 $Y2=0.74
cc_50 VNB N_X_c_960_n 0.00215522f $X=-0.19 $Y=-0.245 $X2=4.155 $Y2=1.765
cc_51 VNB N_X_c_961_n 9.52819e-19 $X=-0.19 $Y=-0.245 $X2=4.38 $Y2=0.74
cc_52 VNB N_X_c_962_n 0.00102081f $X=-0.19 $Y=-0.245 $X2=4.38 $Y2=0.74
cc_53 VNB N_X_c_963_n 0.00161278f $X=-0.19 $Y=-0.245 $X2=4.605 $Y2=1.765
cc_54 VNB N_X_c_964_n 0.00185376f $X=-0.19 $Y=-0.245 $X2=4.605 $Y2=2.4
cc_55 VNB N_X_c_965_n 8.00742e-19 $X=-0.19 $Y=-0.245 $X2=4.95 $Y2=0.74
cc_56 VNB N_X_c_966_n 6.01852e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_X_c_967_n 0.00381929f $X=-0.19 $Y=-0.245 $X2=5.38 $Y2=0.74
cc_58 VNB N_X_c_968_n 0.00583215f $X=-0.19 $Y=-0.245 $X2=5.955 $Y2=1.765
cc_59 VNB N_X_c_969_n 0.0016134f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_X_c_970_n 0.00174684f $X=-0.19 $Y=-0.245 $X2=8.885 $Y2=0.515
cc_61 VNB N_VGND_c_1213_n 0.0111565f $X=-0.19 $Y=-0.245 $X2=1.405 $Y2=1.765
cc_62 VNB N_VGND_c_1214_n 0.0498217f $X=-0.19 $Y=-0.245 $X2=1.405 $Y2=2.4
cc_63 VNB N_VGND_c_1215_n 0.00680404f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_VGND_c_1216_n 0.00938264f $X=-0.19 $Y=-0.245 $X2=2.23 $Y2=1.3
cc_65 VNB N_VGND_c_1217_n 0.00798157f $X=-0.19 $Y=-0.245 $X2=2.355 $Y2=1.765
cc_66 VNB N_VGND_c_1218_n 0.00928684f $X=-0.19 $Y=-0.245 $X2=2.66 $Y2=0.74
cc_67 VNB N_VGND_c_1219_n 0.0203336f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_VGND_c_1220_n 0.0104738f $X=-0.19 $Y=-0.245 $X2=3.09 $Y2=1.3
cc_69 VNB N_VGND_c_1221_n 0.0189682f $X=-0.19 $Y=-0.245 $X2=3.09 $Y2=0.74
cc_70 VNB N_VGND_c_1222_n 0.00830803f $X=-0.19 $Y=-0.245 $X2=3.255 $Y2=2.4
cc_71 VNB N_VGND_c_1223_n 0.0107583f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_VGND_c_1224_n 0.0169342f $X=-0.19 $Y=-0.245 $X2=3.705 $Y2=2.4
cc_73 VNB N_VGND_c_1225_n 0.002601f $X=-0.19 $Y=-0.245 $X2=3.95 $Y2=0.74
cc_74 VNB N_VGND_c_1226_n 0.00250542f $X=-0.19 $Y=-0.245 $X2=4.155 $Y2=2.4
cc_75 VNB N_VGND_c_1227_n 0.00498382f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_VGND_c_1228_n 0.0120272f $X=-0.19 $Y=-0.245 $X2=4.605 $Y2=2.4
cc_77 VNB N_VGND_c_1229_n 0.0417239f $X=-0.19 $Y=-0.245 $X2=4.95 $Y2=1.3
cc_78 VNB N_VGND_c_1230_n 0.0173714f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VNB N_VGND_c_1231_n 0.00394313f $X=-0.19 $Y=-0.245 $X2=5.055 $Y2=1.765
cc_80 VNB N_VGND_c_1232_n 0.019839f $X=-0.19 $Y=-0.245 $X2=5.055 $Y2=2.4
cc_81 VNB N_VGND_c_1233_n 0.00326991f $X=-0.19 $Y=-0.245 $X2=5.38 $Y2=1.3
cc_82 VNB N_VGND_c_1234_n 0.0198781f $X=-0.19 $Y=-0.245 $X2=5.38 $Y2=0.74
cc_83 VNB N_VGND_c_1235_n 0.00326991f $X=-0.19 $Y=-0.245 $X2=5.38 $Y2=0.74
cc_84 VNB N_VGND_c_1236_n 0.0186948f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_85 VNB N_VGND_c_1237_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=5.505 $Y2=1.765
cc_86 VNB N_VGND_c_1238_n 0.0172134f $X=-0.19 $Y=-0.245 $X2=5.95 $Y2=1.3
cc_87 VNB N_VGND_c_1239_n 0.0151736f $X=-0.19 $Y=-0.245 $X2=6.95 $Y2=0.74
cc_88 VNB N_VGND_c_1240_n 0.0151736f $X=-0.19 $Y=-0.245 $X2=7.38 $Y2=1.3
cc_89 VNB N_VGND_c_1241_n 0.018048f $X=-0.19 $Y=-0.245 $X2=7.59 $Y2=1.095
cc_90 VNB N_VGND_c_1242_n 0.0054847f $X=-0.19 $Y=-0.245 $X2=8.025 $Y2=0.515
cc_91 VNB N_VGND_c_1243_n 0.00528956f $X=-0.19 $Y=-0.245 $X2=8.11 $Y2=1.095
cc_92 VNB N_VGND_c_1244_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=8.93 $Y2=2.12
cc_93 VNB N_VGND_c_1245_n 0.00604233f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_94 VNB N_VGND_c_1246_n 0.00604233f $X=-0.19 $Y=-0.245 $X2=8.885 $Y2=0.515
cc_95 VNB N_VGND_c_1247_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=8.97 $Y2=1.095
cc_96 VNB N_VGND_c_1248_n 0.559056f $X=-0.19 $Y=-0.245 $X2=9.83 $Y2=2.815
cc_97 VPB N_A_83_260#_c_216_n 0.0174338f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.765
cc_98 VPB N_A_83_260#_c_217_n 0.0156243f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=1.765
cc_99 VPB N_A_83_260#_c_218_n 0.015236f $X=-0.19 $Y=1.66 $X2=1.405 $Y2=1.765
cc_100 VPB N_A_83_260#_c_219_n 0.0159493f $X=-0.19 $Y=1.66 $X2=1.855 $Y2=1.765
cc_101 VPB N_A_83_260#_c_220_n 0.0156164f $X=-0.19 $Y=1.66 $X2=2.355 $Y2=1.765
cc_102 VPB N_A_83_260#_c_221_n 0.0155721f $X=-0.19 $Y=1.66 $X2=2.805 $Y2=1.765
cc_103 VPB N_A_83_260#_c_222_n 0.0152217f $X=-0.19 $Y=1.66 $X2=3.255 $Y2=1.765
cc_104 VPB N_A_83_260#_c_223_n 0.0155751f $X=-0.19 $Y=1.66 $X2=3.705 $Y2=1.765
cc_105 VPB N_A_83_260#_c_224_n 0.0152378f $X=-0.19 $Y=1.66 $X2=4.155 $Y2=1.765
cc_106 VPB N_A_83_260#_c_225_n 0.0154838f $X=-0.19 $Y=1.66 $X2=4.605 $Y2=1.765
cc_107 VPB N_A_83_260#_c_226_n 0.0152381f $X=-0.19 $Y=1.66 $X2=5.055 $Y2=1.765
cc_108 VPB N_A_83_260#_c_227_n 0.0155744f $X=-0.19 $Y=1.66 $X2=5.505 $Y2=1.765
cc_109 VPB N_A_83_260#_c_228_n 0.0155725f $X=-0.19 $Y=1.66 $X2=5.955 $Y2=1.765
cc_110 VPB N_A_83_260#_c_229_n 0.0155387f $X=-0.19 $Y=1.66 $X2=6.405 $Y2=1.765
cc_111 VPB N_A_83_260#_c_230_n 0.0155725f $X=-0.19 $Y=1.66 $X2=6.855 $Y2=1.765
cc_112 VPB N_A_83_260#_c_231_n 0.0158479f $X=-0.19 $Y=1.66 $X2=7.305 $Y2=1.765
cc_113 VPB N_A_83_260#_c_232_n 0.00257348f $X=-0.19 $Y=1.66 $X2=8.03 $Y2=2.815
cc_114 VPB N_A_83_260#_c_233_n 0.00257348f $X=-0.19 $Y=1.66 $X2=8.93 $Y2=2.815
cc_115 VPB N_A_83_260#_c_234_n 0.00257348f $X=-0.19 $Y=1.66 $X2=9.83 $Y2=2.815
cc_116 VPB N_A_83_260#_c_206_n 0.0169336f $X=-0.19 $Y=1.66 $X2=7.505 $Y2=1.665
cc_117 VPB N_A_83_260#_c_207_n 0.0019053f $X=-0.19 $Y=1.66 $X2=7.505 $Y2=1.665
cc_118 VPB N_A_83_260#_c_208_n 0.00226633f $X=-0.19 $Y=1.66 $X2=1.15 $Y2=1.465
cc_119 VPB N_A_83_260#_c_209_n 0.00178272f $X=-0.19 $Y=1.66 $X2=2.035 $Y2=1.465
cc_120 VPB N_A_83_260#_c_210_n 0.00220169f $X=-0.19 $Y=1.66 $X2=2.995 $Y2=1.465
cc_121 VPB N_A_83_260#_c_211_n 0.00227704f $X=-0.19 $Y=1.66 $X2=3.86 $Y2=1.465
cc_122 VPB N_A_83_260#_c_212_n 0.00186064f $X=-0.19 $Y=1.66 $X2=4.72 $Y2=1.465
cc_123 VPB N_A_83_260#_c_213_n 0.00235875f $X=-0.19 $Y=1.66 $X2=5.74 $Y2=1.465
cc_124 VPB N_A_83_260#_c_214_n 0.00246f $X=-0.19 $Y=1.66 $X2=6.665 $Y2=1.465
cc_125 VPB N_A_83_260#_c_215_n 0.0956002f $X=-0.19 $Y=1.66 $X2=7.305 $Y2=1.532
cc_126 VPB N_A_c_647_n 0.016206f $X=-0.19 $Y=1.66 $X2=7.885 $Y2=0.37
cc_127 VPB N_A_c_648_n 0.0154919f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_128 VPB N_A_c_649_n 0.0155127f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.765
cc_129 VPB N_A_c_650_n 0.0155127f $X=-0.19 $Y=1.66 $X2=0.94 $Y2=1.3
cc_130 VPB N_A_c_651_n 0.0155127f $X=-0.19 $Y=1.66 $X2=1.37 $Y2=1.3
cc_131 VPB N_A_c_652_n 0.0179811f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_132 VPB A 0.0240837f $X=-0.19 $Y=1.66 $X2=2.23 $Y2=1.3
cc_133 VPB N_A_c_646_n 0.0746346f $X=-0.19 $Y=1.66 $X2=3.52 $Y2=0.74
cc_134 VPB N_VPWR_c_765_n 0.0106521f $X=-0.19 $Y=1.66 $X2=1.405 $Y2=1.765
cc_135 VPB N_VPWR_c_766_n 0.0645736f $X=-0.19 $Y=1.66 $X2=1.405 $Y2=2.4
cc_136 VPB N_VPWR_c_767_n 0.00800739f $X=-0.19 $Y=1.66 $X2=1.855 $Y2=2.4
cc_137 VPB N_VPWR_c_768_n 0.00893377f $X=-0.19 $Y=1.66 $X2=2.355 $Y2=1.765
cc_138 VPB N_VPWR_c_769_n 0.00800466f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_139 VPB N_VPWR_c_770_n 0.00800739f $X=-0.19 $Y=1.66 $X2=3.09 $Y2=0.74
cc_140 VPB N_VPWR_c_771_n 0.00799266f $X=-0.19 $Y=1.66 $X2=3.52 $Y2=0.74
cc_141 VPB N_VPWR_c_772_n 0.00800775f $X=-0.19 $Y=1.66 $X2=3.95 $Y2=1.3
cc_142 VPB N_VPWR_c_773_n 0.00800761f $X=-0.19 $Y=1.66 $X2=4.155 $Y2=2.4
cc_143 VPB N_VPWR_c_774_n 0.00886117f $X=-0.19 $Y=1.66 $X2=4.605 $Y2=2.4
cc_144 VPB N_VPWR_c_775_n 0.0196495f $X=-0.19 $Y=1.66 $X2=4.95 $Y2=1.3
cc_145 VPB N_VPWR_c_776_n 0.00799266f $X=-0.19 $Y=1.66 $X2=5.055 $Y2=1.765
cc_146 VPB N_VPWR_c_777_n 0.0206041f $X=-0.19 $Y=1.66 $X2=5.055 $Y2=2.4
cc_147 VPB N_VPWR_c_778_n 0.00799266f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_148 VPB N_VPWR_c_779_n 0.0106521f $X=-0.19 $Y=1.66 $X2=5.505 $Y2=2.4
cc_149 VPB N_VPWR_c_780_n 0.0498694f $X=-0.19 $Y=1.66 $X2=5.95 $Y2=1.3
cc_150 VPB N_VPWR_c_781_n 0.02119f $X=-0.19 $Y=1.66 $X2=5.955 $Y2=2.4
cc_151 VPB N_VPWR_c_782_n 0.00324402f $X=-0.19 $Y=1.66 $X2=5.955 $Y2=2.4
cc_152 VPB N_VPWR_c_783_n 0.0202353f $X=-0.19 $Y=1.66 $X2=6.38 $Y2=0.74
cc_153 VPB N_VPWR_c_784_n 0.0047828f $X=-0.19 $Y=1.66 $X2=6.38 $Y2=0.74
cc_154 VPB N_VPWR_c_785_n 0.0211509f $X=-0.19 $Y=1.66 $X2=6.405 $Y2=1.765
cc_155 VPB N_VPWR_c_786_n 0.00324402f $X=-0.19 $Y=1.66 $X2=6.405 $Y2=2.4
cc_156 VPB N_VPWR_c_787_n 0.02119f $X=-0.19 $Y=1.66 $X2=6.855 $Y2=1.765
cc_157 VPB N_VPWR_c_788_n 0.00324402f $X=-0.19 $Y=1.66 $X2=6.855 $Y2=2.4
cc_158 VPB N_VPWR_c_789_n 0.0206041f $X=-0.19 $Y=1.66 $X2=6.95 $Y2=1.3
cc_159 VPB N_VPWR_c_790_n 0.00324402f $X=-0.19 $Y=1.66 $X2=6.95 $Y2=0.74
cc_160 VPB N_VPWR_c_791_n 0.0208775f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_161 VPB N_VPWR_c_792_n 0.00324402f $X=-0.19 $Y=1.66 $X2=7.305 $Y2=1.765
cc_162 VPB N_VPWR_c_793_n 0.02106f $X=-0.19 $Y=1.66 $X2=7.305 $Y2=2.4
cc_163 VPB N_VPWR_c_794_n 0.00324402f $X=-0.19 $Y=1.66 $X2=7.38 $Y2=1.3
cc_164 VPB N_VPWR_c_795_n 0.0211119f $X=-0.19 $Y=1.66 $X2=7.38 $Y2=0.74
cc_165 VPB N_VPWR_c_796_n 0.0047828f $X=-0.19 $Y=1.66 $X2=7.38 $Y2=0.74
cc_166 VPB N_VPWR_c_797_n 0.0206041f $X=-0.19 $Y=1.66 $X2=9.665 $Y2=2.035
cc_167 VPB N_VPWR_c_798_n 0.00324402f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_168 VPB N_VPWR_c_799_n 0.00324402f $X=-0.19 $Y=1.66 $X2=8.03 $Y2=2.035
cc_169 VPB N_VPWR_c_764_n 0.137465f $X=-0.19 $Y=1.66 $X2=8.93 $Y2=2.115
cc_170 VPB N_X_c_971_n 0.00257348f $X=-0.19 $Y=1.66 $X2=3.255 $Y2=2.4
cc_171 VPB N_X_c_972_n 4.54153e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_172 VPB N_X_c_963_n 9.50018e-19 $X=-0.19 $Y=1.66 $X2=4.605 $Y2=1.765
cc_173 VPB N_X_c_967_n 0.00329612f $X=-0.19 $Y=1.66 $X2=5.38 $Y2=0.74
cc_174 VPB N_X_c_968_n 0.003249f $X=-0.19 $Y=1.66 $X2=5.955 $Y2=1.765
cc_175 VPB N_X_c_976_n 0.00321933f $X=-0.19 $Y=1.66 $X2=6.855 $Y2=1.765
cc_176 VPB N_X_c_977_n 0.00218493f $X=-0.19 $Y=1.66 $X2=7.305 $Y2=1.765
cc_177 VPB N_X_c_978_n 0.00357941f $X=-0.19 $Y=1.66 $X2=7.94 $Y2=1.095
cc_178 VPB N_X_c_969_n 0.00426681f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_179 VPB N_X_c_980_n 0.0032758f $X=-0.19 $Y=1.66 $X2=8.765 $Y2=2.035
cc_180 VPB N_X_c_970_n 0.00107279f $X=-0.19 $Y=1.66 $X2=8.885 $Y2=0.515
cc_181 N_A_83_260#_c_231_n N_A_c_647_n 0.0263543f $X=7.305 $Y=1.765 $X2=-0.19
+ $Y2=-0.245
cc_182 N_A_83_260#_c_246_p N_A_c_647_n 0.0132788f $X=7.865 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_183 N_A_83_260#_c_232_n N_A_c_647_n 0.0100846f $X=8.03 $Y=2.815 $X2=-0.19
+ $Y2=-0.245
cc_184 N_A_83_260#_c_248_p N_A_c_647_n 4.27055e-19 $X=8.03 $Y=2.115 $X2=-0.19
+ $Y2=-0.245
cc_185 N_A_83_260#_c_206_n N_A_c_647_n 3.16139e-19 $X=7.505 $Y=1.665 $X2=-0.19
+ $Y2=-0.245
cc_186 N_A_83_260#_c_207_n N_A_c_647_n 0.00386278f $X=7.505 $Y=1.665 $X2=-0.19
+ $Y2=-0.245
cc_187 N_A_83_260#_M1042_g N_A_M1002_g 0.0311726f $X=7.38 $Y=0.74 $X2=0 $Y2=0
cc_188 N_A_83_260#_c_198_n N_A_M1002_g 0.0142669f $X=7.94 $Y=1.095 $X2=0 $Y2=0
cc_189 N_A_83_260#_c_199_n N_A_M1002_g 3.92313e-19 $X=8.025 $Y=0.515 $X2=0 $Y2=0
cc_190 N_A_83_260#_c_207_n N_A_M1002_g 0.00360365f $X=7.505 $Y=1.665 $X2=0 $Y2=0
cc_191 N_A_83_260#_c_199_n N_A_M1005_g 3.92313e-19 $X=8.025 $Y=0.515 $X2=0 $Y2=0
cc_192 N_A_83_260#_c_200_n N_A_M1005_g 0.0130918f $X=8.8 $Y=1.095 $X2=0 $Y2=0
cc_193 N_A_83_260#_c_232_n N_A_c_648_n 0.0103431f $X=8.03 $Y=2.815 $X2=0 $Y2=0
cc_194 N_A_83_260#_c_258_p N_A_c_648_n 0.0120074f $X=8.765 $Y=2.035 $X2=0 $Y2=0
cc_195 N_A_83_260#_c_233_n N_A_c_648_n 6.45594e-19 $X=8.93 $Y=2.815 $X2=0 $Y2=0
cc_196 N_A_83_260#_c_248_p N_A_c_648_n 4.27055e-19 $X=8.03 $Y=2.115 $X2=0 $Y2=0
cc_197 N_A_83_260#_c_200_n N_A_M1011_g 0.0130918f $X=8.8 $Y=1.095 $X2=0 $Y2=0
cc_198 N_A_83_260#_c_201_n N_A_M1011_g 3.92313e-19 $X=8.885 $Y=0.515 $X2=0 $Y2=0
cc_199 N_A_83_260#_c_232_n N_A_c_649_n 6.45594e-19 $X=8.03 $Y=2.815 $X2=0 $Y2=0
cc_200 N_A_83_260#_c_258_p N_A_c_649_n 0.0120074f $X=8.765 $Y=2.035 $X2=0 $Y2=0
cc_201 N_A_83_260#_c_233_n N_A_c_649_n 0.0103431f $X=8.93 $Y=2.815 $X2=0 $Y2=0
cc_202 N_A_83_260#_c_266_p N_A_c_649_n 4.27055e-19 $X=8.93 $Y=2.115 $X2=0 $Y2=0
cc_203 N_A_83_260#_c_201_n N_A_M1012_g 3.92313e-19 $X=8.885 $Y=0.515 $X2=0 $Y2=0
cc_204 N_A_83_260#_c_202_n N_A_M1012_g 0.0132977f $X=9.695 $Y=1.095 $X2=0 $Y2=0
cc_205 N_A_83_260#_c_233_n N_A_c_650_n 0.0103431f $X=8.93 $Y=2.815 $X2=0 $Y2=0
cc_206 N_A_83_260#_c_270_p N_A_c_650_n 0.0120074f $X=9.665 $Y=2.035 $X2=0 $Y2=0
cc_207 N_A_83_260#_c_234_n N_A_c_650_n 6.45594e-19 $X=9.83 $Y=2.815 $X2=0 $Y2=0
cc_208 N_A_83_260#_c_266_p N_A_c_650_n 4.27055e-19 $X=8.93 $Y=2.115 $X2=0 $Y2=0
cc_209 N_A_83_260#_c_202_n N_A_M1013_g 0.0140368f $X=9.695 $Y=1.095 $X2=0 $Y2=0
cc_210 N_A_83_260#_c_203_n N_A_M1013_g 4.79998e-19 $X=9.78 $Y=0.515 $X2=0 $Y2=0
cc_211 N_A_83_260#_c_233_n N_A_c_651_n 6.45594e-19 $X=8.93 $Y=2.815 $X2=0 $Y2=0
cc_212 N_A_83_260#_c_270_p N_A_c_651_n 0.0120074f $X=9.665 $Y=2.035 $X2=0 $Y2=0
cc_213 N_A_83_260#_c_277_p N_A_c_651_n 4.27055e-19 $X=9.83 $Y=2.12 $X2=0 $Y2=0
cc_214 N_A_83_260#_c_234_n N_A_c_651_n 0.0103431f $X=9.83 $Y=2.815 $X2=0 $Y2=0
cc_215 N_A_83_260#_c_277_p N_A_c_652_n 0.00203651f $X=9.83 $Y=2.12 $X2=0 $Y2=0
cc_216 N_A_83_260#_c_234_n N_A_c_652_n 0.00960826f $X=9.83 $Y=2.815 $X2=0 $Y2=0
cc_217 N_A_83_260#_c_202_n N_A_M1043_g 0.00234945f $X=9.695 $Y=1.095 $X2=0 $Y2=0
cc_218 N_A_83_260#_c_203_n N_A_M1043_g 0.00349953f $X=9.78 $Y=0.515 $X2=0 $Y2=0
cc_219 N_A_83_260#_c_198_n A 0.0122081f $X=7.94 $Y=1.095 $X2=0 $Y2=0
cc_220 N_A_83_260#_c_246_p A 0.0065328f $X=7.865 $Y=2.035 $X2=0 $Y2=0
cc_221 N_A_83_260#_c_200_n A 0.0517342f $X=8.8 $Y=1.095 $X2=0 $Y2=0
cc_222 N_A_83_260#_c_258_p A 0.0393875f $X=8.765 $Y=2.035 $X2=0 $Y2=0
cc_223 N_A_83_260#_c_202_n A 0.0758934f $X=9.695 $Y=1.095 $X2=0 $Y2=0
cc_224 N_A_83_260#_c_270_p A 0.0393875f $X=9.665 $Y=2.035 $X2=0 $Y2=0
cc_225 N_A_83_260#_c_277_p A 0.0237598f $X=9.83 $Y=2.12 $X2=0 $Y2=0
cc_226 N_A_83_260#_c_248_p A 0.0237598f $X=8.03 $Y=2.115 $X2=0 $Y2=0
cc_227 N_A_83_260#_c_204_n A 0.0146029f $X=8.025 $Y=1.095 $X2=0 $Y2=0
cc_228 N_A_83_260#_c_266_p A 0.0237598f $X=8.93 $Y=2.115 $X2=0 $Y2=0
cc_229 N_A_83_260#_c_205_n A 0.0146029f $X=8.885 $Y=1.095 $X2=0 $Y2=0
cc_230 N_A_83_260#_c_206_n A 0.00817464f $X=7.505 $Y=1.665 $X2=0 $Y2=0
cc_231 N_A_83_260#_c_207_n A 0.029276f $X=7.505 $Y=1.665 $X2=0 $Y2=0
cc_232 N_A_83_260#_c_215_n A 2.51865e-19 $X=7.305 $Y=1.532 $X2=0 $Y2=0
cc_233 N_A_83_260#_c_198_n N_A_c_646_n 7.87309e-19 $X=7.94 $Y=1.095 $X2=0 $Y2=0
cc_234 N_A_83_260#_c_200_n N_A_c_646_n 0.00224206f $X=8.8 $Y=1.095 $X2=0 $Y2=0
cc_235 N_A_83_260#_c_258_p N_A_c_646_n 0.00130859f $X=8.765 $Y=2.035 $X2=0 $Y2=0
cc_236 N_A_83_260#_c_202_n N_A_c_646_n 0.00698704f $X=9.695 $Y=1.095 $X2=0 $Y2=0
cc_237 N_A_83_260#_c_270_p N_A_c_646_n 0.00131106f $X=9.665 $Y=2.035 $X2=0 $Y2=0
cc_238 N_A_83_260#_c_277_p N_A_c_646_n 0.00144657f $X=9.83 $Y=2.12 $X2=0 $Y2=0
cc_239 N_A_83_260#_c_248_p N_A_c_646_n 0.00144162f $X=8.03 $Y=2.115 $X2=0 $Y2=0
cc_240 N_A_83_260#_c_204_n N_A_c_646_n 0.00232957f $X=8.025 $Y=1.095 $X2=0 $Y2=0
cc_241 N_A_83_260#_c_266_p N_A_c_646_n 0.00144162f $X=8.93 $Y=2.115 $X2=0 $Y2=0
cc_242 N_A_83_260#_c_205_n N_A_c_646_n 0.00232957f $X=8.885 $Y=1.095 $X2=0 $Y2=0
cc_243 N_A_83_260#_c_206_n N_A_c_646_n 0.00475455f $X=7.505 $Y=1.665 $X2=0 $Y2=0
cc_244 N_A_83_260#_c_207_n N_A_c_646_n 0.00300854f $X=7.505 $Y=1.665 $X2=0 $Y2=0
cc_245 N_A_83_260#_c_215_n N_A_c_646_n 0.0191885f $X=7.305 $Y=1.532 $X2=0 $Y2=0
cc_246 N_A_83_260#_c_246_p N_VPWR_M1040_d 0.00251411f $X=7.865 $Y=2.035 $X2=0
+ $Y2=0
cc_247 N_A_83_260#_c_311_p N_VPWR_M1040_d 0.00305175f $X=7.59 $Y=2.035 $X2=0
+ $Y2=0
cc_248 N_A_83_260#_c_207_n N_VPWR_M1040_d 0.00192268f $X=7.505 $Y=1.665 $X2=0
+ $Y2=0
cc_249 N_A_83_260#_c_258_p N_VPWR_M1006_s 0.00408911f $X=8.765 $Y=2.035 $X2=0
+ $Y2=0
cc_250 N_A_83_260#_c_270_p N_VPWR_M1031_s 0.00408911f $X=9.665 $Y=2.035 $X2=0
+ $Y2=0
cc_251 N_A_83_260#_c_216_n N_VPWR_c_766_n 0.0100009f $X=0.505 $Y=1.765 $X2=0
+ $Y2=0
cc_252 N_A_83_260#_c_217_n N_VPWR_c_767_n 0.00688828f $X=0.955 $Y=1.765 $X2=0
+ $Y2=0
cc_253 N_A_83_260#_c_218_n N_VPWR_c_767_n 0.00580064f $X=1.405 $Y=1.765 $X2=0
+ $Y2=0
cc_254 N_A_83_260#_c_208_n N_VPWR_c_767_n 0.011185f $X=1.15 $Y=1.465 $X2=0 $Y2=0
cc_255 N_A_83_260#_c_215_n N_VPWR_c_767_n 7.65868e-19 $X=7.305 $Y=1.532 $X2=0
+ $Y2=0
cc_256 N_A_83_260#_c_219_n N_VPWR_c_768_n 0.00867391f $X=1.855 $Y=1.765 $X2=0
+ $Y2=0
cc_257 N_A_83_260#_c_220_n N_VPWR_c_768_n 0.00634247f $X=2.355 $Y=1.765 $X2=0
+ $Y2=0
cc_258 N_A_83_260#_c_206_n N_VPWR_c_768_n 4.79551e-19 $X=7.505 $Y=1.665 $X2=0
+ $Y2=0
cc_259 N_A_83_260#_c_209_n N_VPWR_c_768_n 0.0135207f $X=2.035 $Y=1.465 $X2=0
+ $Y2=0
cc_260 N_A_83_260#_c_215_n N_VPWR_c_768_n 0.00190937f $X=7.305 $Y=1.532 $X2=0
+ $Y2=0
cc_261 N_A_83_260#_c_221_n N_VPWR_c_769_n 0.00675646f $X=2.805 $Y=1.765 $X2=0
+ $Y2=0
cc_262 N_A_83_260#_c_222_n N_VPWR_c_769_n 0.0057301f $X=3.255 $Y=1.765 $X2=0
+ $Y2=0
cc_263 N_A_83_260#_c_210_n N_VPWR_c_769_n 0.011185f $X=2.995 $Y=1.465 $X2=0
+ $Y2=0
cc_264 N_A_83_260#_c_215_n N_VPWR_c_769_n 7.59789e-19 $X=7.305 $Y=1.532 $X2=0
+ $Y2=0
cc_265 N_A_83_260#_c_223_n N_VPWR_c_770_n 0.00688828f $X=3.705 $Y=1.765 $X2=0
+ $Y2=0
cc_266 N_A_83_260#_c_224_n N_VPWR_c_770_n 0.00580064f $X=4.155 $Y=1.765 $X2=0
+ $Y2=0
cc_267 N_A_83_260#_c_211_n N_VPWR_c_770_n 0.011185f $X=3.86 $Y=1.465 $X2=0 $Y2=0
cc_268 N_A_83_260#_c_215_n N_VPWR_c_770_n 7.59789e-19 $X=7.305 $Y=1.532 $X2=0
+ $Y2=0
cc_269 N_A_83_260#_c_225_n N_VPWR_c_771_n 0.00580064f $X=4.605 $Y=1.765 $X2=0
+ $Y2=0
cc_270 N_A_83_260#_c_226_n N_VPWR_c_771_n 0.00580064f $X=5.055 $Y=1.765 $X2=0
+ $Y2=0
cc_271 N_A_83_260#_c_206_n N_VPWR_c_771_n 4.48561e-19 $X=7.505 $Y=1.665 $X2=0
+ $Y2=0
cc_272 N_A_83_260#_c_212_n N_VPWR_c_771_n 0.0079227f $X=4.72 $Y=1.465 $X2=0
+ $Y2=0
cc_273 N_A_83_260#_c_215_n N_VPWR_c_771_n 0.00173834f $X=7.305 $Y=1.532 $X2=0
+ $Y2=0
cc_274 N_A_83_260#_c_227_n N_VPWR_c_772_n 0.00628588f $X=5.505 $Y=1.765 $X2=0
+ $Y2=0
cc_275 N_A_83_260#_c_228_n N_VPWR_c_772_n 0.0064218f $X=5.955 $Y=1.765 $X2=0
+ $Y2=0
cc_276 N_A_83_260#_c_213_n N_VPWR_c_772_n 0.011185f $X=5.74 $Y=1.465 $X2=0 $Y2=0
cc_277 N_A_83_260#_c_215_n N_VPWR_c_772_n 7.68239e-19 $X=7.305 $Y=1.532 $X2=0
+ $Y2=0
cc_278 N_A_83_260#_c_229_n N_VPWR_c_773_n 0.00601042f $X=6.405 $Y=1.765 $X2=0
+ $Y2=0
cc_279 N_A_83_260#_c_230_n N_VPWR_c_773_n 0.00669011f $X=6.855 $Y=1.765 $X2=0
+ $Y2=0
cc_280 N_A_83_260#_c_214_n N_VPWR_c_773_n 0.011185f $X=6.665 $Y=1.465 $X2=0
+ $Y2=0
cc_281 N_A_83_260#_c_215_n N_VPWR_c_773_n 7.70002e-19 $X=7.305 $Y=1.532 $X2=0
+ $Y2=0
cc_282 N_A_83_260#_c_231_n N_VPWR_c_774_n 0.00534288f $X=7.305 $Y=1.765 $X2=0
+ $Y2=0
cc_283 N_A_83_260#_c_246_p N_VPWR_c_774_n 0.00653467f $X=7.865 $Y=2.035 $X2=0
+ $Y2=0
cc_284 N_A_83_260#_c_311_p N_VPWR_c_774_n 0.0125073f $X=7.59 $Y=2.035 $X2=0
+ $Y2=0
cc_285 N_A_83_260#_c_232_n N_VPWR_c_774_n 0.0266484f $X=8.03 $Y=2.815 $X2=0
+ $Y2=0
cc_286 N_A_83_260#_c_206_n N_VPWR_c_774_n 7.55387e-19 $X=7.505 $Y=1.665 $X2=0
+ $Y2=0
cc_287 N_A_83_260#_c_232_n N_VPWR_c_775_n 0.014552f $X=8.03 $Y=2.815 $X2=0 $Y2=0
cc_288 N_A_83_260#_c_232_n N_VPWR_c_776_n 0.0449718f $X=8.03 $Y=2.815 $X2=0
+ $Y2=0
cc_289 N_A_83_260#_c_258_p N_VPWR_c_776_n 0.0136682f $X=8.765 $Y=2.035 $X2=0
+ $Y2=0
cc_290 N_A_83_260#_c_233_n N_VPWR_c_776_n 0.0449718f $X=8.93 $Y=2.815 $X2=0
+ $Y2=0
cc_291 N_A_83_260#_c_233_n N_VPWR_c_777_n 0.014552f $X=8.93 $Y=2.815 $X2=0 $Y2=0
cc_292 N_A_83_260#_c_233_n N_VPWR_c_778_n 0.0449718f $X=8.93 $Y=2.815 $X2=0
+ $Y2=0
cc_293 N_A_83_260#_c_270_p N_VPWR_c_778_n 0.0136682f $X=9.665 $Y=2.035 $X2=0
+ $Y2=0
cc_294 N_A_83_260#_c_234_n N_VPWR_c_778_n 0.0449718f $X=9.83 $Y=2.815 $X2=0
+ $Y2=0
cc_295 N_A_83_260#_c_277_p N_VPWR_c_780_n 0.0121024f $X=9.83 $Y=2.12 $X2=0 $Y2=0
cc_296 N_A_83_260#_c_234_n N_VPWR_c_780_n 0.0576605f $X=9.83 $Y=2.815 $X2=0
+ $Y2=0
cc_297 N_A_83_260#_c_216_n N_VPWR_c_781_n 0.00439937f $X=0.505 $Y=1.765 $X2=0
+ $Y2=0
cc_298 N_A_83_260#_c_217_n N_VPWR_c_781_n 0.00461464f $X=0.955 $Y=1.765 $X2=0
+ $Y2=0
cc_299 N_A_83_260#_c_218_n N_VPWR_c_783_n 0.00445602f $X=1.405 $Y=1.765 $X2=0
+ $Y2=0
cc_300 N_A_83_260#_c_219_n N_VPWR_c_783_n 0.00461464f $X=1.855 $Y=1.765 $X2=0
+ $Y2=0
cc_301 N_A_83_260#_c_220_n N_VPWR_c_785_n 0.00445602f $X=2.355 $Y=1.765 $X2=0
+ $Y2=0
cc_302 N_A_83_260#_c_221_n N_VPWR_c_785_n 0.00461464f $X=2.805 $Y=1.765 $X2=0
+ $Y2=0
cc_303 N_A_83_260#_c_222_n N_VPWR_c_787_n 0.00439937f $X=3.255 $Y=1.765 $X2=0
+ $Y2=0
cc_304 N_A_83_260#_c_223_n N_VPWR_c_787_n 0.00461464f $X=3.705 $Y=1.765 $X2=0
+ $Y2=0
cc_305 N_A_83_260#_c_224_n N_VPWR_c_789_n 0.00445602f $X=4.155 $Y=1.765 $X2=0
+ $Y2=0
cc_306 N_A_83_260#_c_225_n N_VPWR_c_789_n 0.00445602f $X=4.605 $Y=1.765 $X2=0
+ $Y2=0
cc_307 N_A_83_260#_c_226_n N_VPWR_c_791_n 0.00445602f $X=5.055 $Y=1.765 $X2=0
+ $Y2=0
cc_308 N_A_83_260#_c_227_n N_VPWR_c_791_n 0.00461464f $X=5.505 $Y=1.765 $X2=0
+ $Y2=0
cc_309 N_A_83_260#_c_228_n N_VPWR_c_793_n 0.00461464f $X=5.955 $Y=1.765 $X2=0
+ $Y2=0
cc_310 N_A_83_260#_c_229_n N_VPWR_c_793_n 0.00461464f $X=6.405 $Y=1.765 $X2=0
+ $Y2=0
cc_311 N_A_83_260#_c_230_n N_VPWR_c_795_n 0.00461464f $X=6.855 $Y=1.765 $X2=0
+ $Y2=0
cc_312 N_A_83_260#_c_231_n N_VPWR_c_795_n 0.00445602f $X=7.305 $Y=1.765 $X2=0
+ $Y2=0
cc_313 N_A_83_260#_c_234_n N_VPWR_c_797_n 0.014552f $X=9.83 $Y=2.815 $X2=0 $Y2=0
cc_314 N_A_83_260#_c_216_n N_VPWR_c_764_n 0.0084274f $X=0.505 $Y=1.765 $X2=0
+ $Y2=0
cc_315 N_A_83_260#_c_217_n N_VPWR_c_764_n 0.00908951f $X=0.955 $Y=1.765 $X2=0
+ $Y2=0
cc_316 N_A_83_260#_c_218_n N_VPWR_c_764_n 0.00857589f $X=1.405 $Y=1.765 $X2=0
+ $Y2=0
cc_317 N_A_83_260#_c_219_n N_VPWR_c_764_n 0.0090874f $X=1.855 $Y=1.765 $X2=0
+ $Y2=0
cc_318 N_A_83_260#_c_220_n N_VPWR_c_764_n 0.0085805f $X=2.355 $Y=1.765 $X2=0
+ $Y2=0
cc_319 N_A_83_260#_c_221_n N_VPWR_c_764_n 0.00908951f $X=2.805 $Y=1.765 $X2=0
+ $Y2=0
cc_320 N_A_83_260#_c_222_n N_VPWR_c_764_n 0.00839246f $X=3.255 $Y=1.765 $X2=0
+ $Y2=0
cc_321 N_A_83_260#_c_223_n N_VPWR_c_764_n 0.00908951f $X=3.705 $Y=1.765 $X2=0
+ $Y2=0
cc_322 N_A_83_260#_c_224_n N_VPWR_c_764_n 0.00857589f $X=4.155 $Y=1.765 $X2=0
+ $Y2=0
cc_323 N_A_83_260#_c_225_n N_VPWR_c_764_n 0.00857589f $X=4.605 $Y=1.765 $X2=0
+ $Y2=0
cc_324 N_A_83_260#_c_226_n N_VPWR_c_764_n 0.00857589f $X=5.055 $Y=1.765 $X2=0
+ $Y2=0
cc_325 N_A_83_260#_c_227_n N_VPWR_c_764_n 0.00908951f $X=5.505 $Y=1.765 $X2=0
+ $Y2=0
cc_326 N_A_83_260#_c_228_n N_VPWR_c_764_n 0.00908951f $X=5.955 $Y=1.765 $X2=0
+ $Y2=0
cc_327 N_A_83_260#_c_229_n N_VPWR_c_764_n 0.00908951f $X=6.405 $Y=1.765 $X2=0
+ $Y2=0
cc_328 N_A_83_260#_c_230_n N_VPWR_c_764_n 0.00908951f $X=6.855 $Y=1.765 $X2=0
+ $Y2=0
cc_329 N_A_83_260#_c_231_n N_VPWR_c_764_n 0.00858104f $X=7.305 $Y=1.765 $X2=0
+ $Y2=0
cc_330 N_A_83_260#_c_232_n N_VPWR_c_764_n 0.0119791f $X=8.03 $Y=2.815 $X2=0
+ $Y2=0
cc_331 N_A_83_260#_c_233_n N_VPWR_c_764_n 0.0119791f $X=8.93 $Y=2.815 $X2=0
+ $Y2=0
cc_332 N_A_83_260#_c_234_n N_VPWR_c_764_n 0.0119791f $X=9.83 $Y=2.815 $X2=0
+ $Y2=0
cc_333 N_A_83_260#_M1010_g N_X_c_954_n 0.00300705f $X=2.23 $Y=0.74 $X2=0 $Y2=0
cc_334 N_A_83_260#_M1014_g N_X_c_954_n 0.0116584f $X=2.66 $Y=0.74 $X2=0 $Y2=0
cc_335 N_A_83_260#_M1016_g N_X_c_954_n 7.51209e-19 $X=3.09 $Y=0.74 $X2=0 $Y2=0
cc_336 N_A_83_260#_M1016_g N_X_c_955_n 6.7859e-19 $X=3.09 $Y=0.74 $X2=0 $Y2=0
cc_337 N_A_83_260#_M1019_g N_X_c_955_n 0.00805893f $X=3.52 $Y=0.74 $X2=0 $Y2=0
cc_338 N_A_83_260#_M1023_g N_X_c_955_n 0.00107262f $X=3.95 $Y=0.74 $X2=0 $Y2=0
cc_339 N_A_83_260#_M1023_g N_X_c_956_n 0.00725398f $X=3.95 $Y=0.74 $X2=0 $Y2=0
cc_340 N_A_83_260#_M1024_g N_X_c_956_n 0.0099418f $X=4.38 $Y=0.74 $X2=0 $Y2=0
cc_341 N_A_83_260#_M1032_g N_X_c_956_n 7.58451e-19 $X=4.95 $Y=0.74 $X2=0 $Y2=0
cc_342 N_A_83_260#_c_224_n N_X_c_971_n 0.0100067f $X=4.155 $Y=1.765 $X2=0 $Y2=0
cc_343 N_A_83_260#_c_225_n N_X_c_971_n 0.0100067f $X=4.605 $Y=1.765 $X2=0 $Y2=0
cc_344 N_A_83_260#_M1032_g N_X_c_957_n 0.00326319f $X=4.95 $Y=0.74 $X2=0 $Y2=0
cc_345 N_A_83_260#_M1034_g N_X_c_957_n 0.0124415f $X=5.38 $Y=0.74 $X2=0 $Y2=0
cc_346 N_A_83_260#_M1035_g N_X_c_957_n 7.7473e-19 $X=5.95 $Y=0.74 $X2=0 $Y2=0
cc_347 N_A_83_260#_M1034_g N_X_c_958_n 4.33387e-19 $X=5.38 $Y=0.74 $X2=0 $Y2=0
cc_348 N_A_83_260#_M1035_g N_X_c_958_n 0.00752022f $X=5.95 $Y=0.74 $X2=0 $Y2=0
cc_349 N_A_83_260#_M1038_g N_X_c_958_n 0.00752022f $X=6.38 $Y=0.74 $X2=0 $Y2=0
cc_350 N_A_83_260#_M1041_g N_X_c_958_n 6.82839e-19 $X=6.95 $Y=0.74 $X2=0 $Y2=0
cc_351 N_A_83_260#_M1038_g N_X_c_959_n 5.36216e-19 $X=6.38 $Y=0.74 $X2=0 $Y2=0
cc_352 N_A_83_260#_M1041_g N_X_c_959_n 0.00618203f $X=6.95 $Y=0.74 $X2=0 $Y2=0
cc_353 N_A_83_260#_M1042_g N_X_c_959_n 0.00126597f $X=7.38 $Y=0.74 $X2=0 $Y2=0
cc_354 N_A_83_260#_c_418_p N_X_c_959_n 0.00454316f $X=7.59 $Y=1.095 $X2=0 $Y2=0
cc_355 N_A_83_260#_c_206_n N_X_c_959_n 2.22902e-19 $X=7.505 $Y=1.665 $X2=0 $Y2=0
cc_356 N_A_83_260#_c_207_n N_X_c_959_n 0.0144199f $X=7.505 $Y=1.665 $X2=0 $Y2=0
cc_357 N_A_83_260#_c_214_n N_X_c_959_n 0.00605471f $X=6.665 $Y=1.465 $X2=0 $Y2=0
cc_358 N_A_83_260#_c_215_n N_X_c_959_n 0.00673507f $X=7.305 $Y=1.532 $X2=0 $Y2=0
cc_359 N_A_83_260#_M1041_g N_X_c_960_n 0.00906114f $X=6.95 $Y=0.74 $X2=0 $Y2=0
cc_360 N_A_83_260#_M1042_g N_X_c_960_n 4.99876e-19 $X=7.38 $Y=0.74 $X2=0 $Y2=0
cc_361 N_A_83_260#_c_418_p N_X_c_960_n 0.00536506f $X=7.59 $Y=1.095 $X2=0 $Y2=0
cc_362 N_A_83_260#_M1014_g N_X_c_961_n 0.00706265f $X=2.66 $Y=0.74 $X2=0 $Y2=0
cc_363 N_A_83_260#_M1016_g N_X_c_961_n 4.00131e-19 $X=3.09 $Y=0.74 $X2=0 $Y2=0
cc_364 N_A_83_260#_c_206_n N_X_c_961_n 0.00315312f $X=7.505 $Y=1.665 $X2=0 $Y2=0
cc_365 N_A_83_260#_c_209_n N_X_c_961_n 0.00408163f $X=2.035 $Y=1.465 $X2=0 $Y2=0
cc_366 N_A_83_260#_c_210_n N_X_c_961_n 0.0337701f $X=2.995 $Y=1.465 $X2=0 $Y2=0
cc_367 N_A_83_260#_c_215_n N_X_c_961_n 0.00702624f $X=7.305 $Y=1.532 $X2=0 $Y2=0
cc_368 N_A_83_260#_M1019_g N_X_c_962_n 0.00157629f $X=3.52 $Y=0.74 $X2=0 $Y2=0
cc_369 N_A_83_260#_c_206_n N_X_c_962_n 0.00351265f $X=7.505 $Y=1.665 $X2=0 $Y2=0
cc_370 N_A_83_260#_c_215_n N_X_c_962_n 0.0026612f $X=7.305 $Y=1.532 $X2=0 $Y2=0
cc_371 N_A_83_260#_c_222_n N_X_c_972_n 0.00245312f $X=3.255 $Y=1.765 $X2=0 $Y2=0
cc_372 N_A_83_260#_c_223_n N_X_c_972_n 0.00623279f $X=3.705 $Y=1.765 $X2=0 $Y2=0
cc_373 N_A_83_260#_c_206_n N_X_c_972_n 0.00319451f $X=7.505 $Y=1.665 $X2=0 $Y2=0
cc_374 N_A_83_260#_c_215_n N_X_c_972_n 0.00331433f $X=7.305 $Y=1.532 $X2=0 $Y2=0
cc_375 N_A_83_260#_c_221_n N_X_c_963_n 9.26601e-19 $X=2.805 $Y=1.765 $X2=0 $Y2=0
cc_376 N_A_83_260#_M1016_g N_X_c_963_n 0.00237771f $X=3.09 $Y=0.74 $X2=0 $Y2=0
cc_377 N_A_83_260#_c_222_n N_X_c_963_n 0.00124811f $X=3.255 $Y=1.765 $X2=0 $Y2=0
cc_378 N_A_83_260#_M1019_g N_X_c_963_n 0.00419028f $X=3.52 $Y=0.74 $X2=0 $Y2=0
cc_379 N_A_83_260#_c_223_n N_X_c_963_n 9.19858e-19 $X=3.705 $Y=1.765 $X2=0 $Y2=0
cc_380 N_A_83_260#_c_206_n N_X_c_963_n 0.0207314f $X=7.505 $Y=1.665 $X2=0 $Y2=0
cc_381 N_A_83_260#_c_210_n N_X_c_963_n 0.03315f $X=2.995 $Y=1.465 $X2=0 $Y2=0
cc_382 N_A_83_260#_c_211_n N_X_c_963_n 0.0300775f $X=3.86 $Y=1.465 $X2=0 $Y2=0
cc_383 N_A_83_260#_c_215_n N_X_c_963_n 0.0211102f $X=7.305 $Y=1.532 $X2=0 $Y2=0
cc_384 N_A_83_260#_M1023_g N_X_c_964_n 0.00255654f $X=3.95 $Y=0.74 $X2=0 $Y2=0
cc_385 N_A_83_260#_M1024_g N_X_c_964_n 0.00291493f $X=4.38 $Y=0.74 $X2=0 $Y2=0
cc_386 N_A_83_260#_c_206_n N_X_c_964_n 0.00691749f $X=7.505 $Y=1.665 $X2=0 $Y2=0
cc_387 N_A_83_260#_c_211_n N_X_c_964_n 0.00354025f $X=3.86 $Y=1.465 $X2=0 $Y2=0
cc_388 N_A_83_260#_c_215_n N_X_c_964_n 0.00483855f $X=7.305 $Y=1.532 $X2=0 $Y2=0
cc_389 N_A_83_260#_M1034_g N_X_c_965_n 0.00742086f $X=5.38 $Y=0.74 $X2=0 $Y2=0
cc_390 N_A_83_260#_M1035_g N_X_c_965_n 3.38014e-19 $X=5.95 $Y=0.74 $X2=0 $Y2=0
cc_391 N_A_83_260#_c_206_n N_X_c_965_n 0.00369519f $X=7.505 $Y=1.665 $X2=0 $Y2=0
cc_392 N_A_83_260#_c_212_n N_X_c_965_n 0.00568676f $X=4.72 $Y=1.465 $X2=0 $Y2=0
cc_393 N_A_83_260#_c_213_n N_X_c_965_n 0.0341199f $X=5.74 $Y=1.465 $X2=0 $Y2=0
cc_394 N_A_83_260#_c_215_n N_X_c_965_n 0.0086822f $X=7.305 $Y=1.532 $X2=0 $Y2=0
cc_395 N_A_83_260#_M1035_g N_X_c_966_n 0.00345986f $X=5.95 $Y=0.74 $X2=0 $Y2=0
cc_396 N_A_83_260#_M1038_g N_X_c_966_n 0.00193058f $X=6.38 $Y=0.74 $X2=0 $Y2=0
cc_397 N_A_83_260#_c_206_n N_X_c_966_n 0.00223202f $X=7.505 $Y=1.665 $X2=0 $Y2=0
cc_398 N_A_83_260#_c_216_n N_X_c_967_n 0.0165427f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_399 N_A_83_260#_M1003_g N_X_c_967_n 0.018334f $X=0.51 $Y=0.74 $X2=0 $Y2=0
cc_400 N_A_83_260#_M1004_g N_X_c_967_n 0.00288964f $X=0.94 $Y=0.74 $X2=0 $Y2=0
cc_401 N_A_83_260#_c_217_n N_X_c_967_n 0.00689327f $X=0.955 $Y=1.765 $X2=0 $Y2=0
cc_402 N_A_83_260#_c_206_n N_X_c_967_n 0.0067013f $X=7.505 $Y=1.665 $X2=0 $Y2=0
cc_403 N_A_83_260#_c_208_n N_X_c_967_n 0.0330171f $X=1.15 $Y=1.465 $X2=0 $Y2=0
cc_404 N_A_83_260#_c_215_n N_X_c_967_n 0.0420067f $X=7.305 $Y=1.532 $X2=0 $Y2=0
cc_405 N_A_83_260#_c_217_n N_X_c_968_n 9.31623e-19 $X=0.955 $Y=1.765 $X2=0 $Y2=0
cc_406 N_A_83_260#_M1008_g N_X_c_968_n 0.00307196f $X=1.37 $Y=0.74 $X2=0 $Y2=0
cc_407 N_A_83_260#_c_218_n N_X_c_968_n 0.0145514f $X=1.405 $Y=1.765 $X2=0 $Y2=0
cc_408 N_A_83_260#_M1009_g N_X_c_968_n 0.00311337f $X=1.8 $Y=0.74 $X2=0 $Y2=0
cc_409 N_A_83_260#_c_219_n N_X_c_968_n 0.00856841f $X=1.855 $Y=1.765 $X2=0 $Y2=0
cc_410 N_A_83_260#_c_206_n N_X_c_968_n 0.0283165f $X=7.505 $Y=1.665 $X2=0 $Y2=0
cc_411 N_A_83_260#_c_208_n N_X_c_968_n 0.0338f $X=1.15 $Y=1.465 $X2=0 $Y2=0
cc_412 N_A_83_260#_c_209_n N_X_c_968_n 0.0336509f $X=2.035 $Y=1.465 $X2=0 $Y2=0
cc_413 N_A_83_260#_c_215_n N_X_c_968_n 0.0277364f $X=7.305 $Y=1.532 $X2=0 $Y2=0
cc_414 N_A_83_260#_c_219_n N_X_c_976_n 0.00131022f $X=1.855 $Y=1.765 $X2=0 $Y2=0
cc_415 N_A_83_260#_c_220_n N_X_c_976_n 0.0148683f $X=2.355 $Y=1.765 $X2=0 $Y2=0
cc_416 N_A_83_260#_c_221_n N_X_c_976_n 0.00183216f $X=2.805 $Y=1.765 $X2=0 $Y2=0
cc_417 N_A_83_260#_c_206_n N_X_c_976_n 0.0291691f $X=7.505 $Y=1.665 $X2=0 $Y2=0
cc_418 N_A_83_260#_c_209_n N_X_c_976_n 0.0214656f $X=2.035 $Y=1.465 $X2=0 $Y2=0
cc_419 N_A_83_260#_c_215_n N_X_c_976_n 0.0236446f $X=7.305 $Y=1.532 $X2=0 $Y2=0
cc_420 N_A_83_260#_c_222_n N_X_c_977_n 0.0110055f $X=3.255 $Y=1.765 $X2=0 $Y2=0
cc_421 N_A_83_260#_c_225_n N_X_c_978_n 0.00113175f $X=4.605 $Y=1.765 $X2=0 $Y2=0
cc_422 N_A_83_260#_c_226_n N_X_c_978_n 0.0144632f $X=5.055 $Y=1.765 $X2=0 $Y2=0
cc_423 N_A_83_260#_c_227_n N_X_c_978_n 0.00196959f $X=5.505 $Y=1.765 $X2=0 $Y2=0
cc_424 N_A_83_260#_c_206_n N_X_c_978_n 0.0324735f $X=7.505 $Y=1.665 $X2=0 $Y2=0
cc_425 N_A_83_260#_c_212_n N_X_c_978_n 0.0198131f $X=4.72 $Y=1.465 $X2=0 $Y2=0
cc_426 N_A_83_260#_c_215_n N_X_c_978_n 0.0245861f $X=7.305 $Y=1.532 $X2=0 $Y2=0
cc_427 N_A_83_260#_M1035_g N_X_c_969_n 0.00334296f $X=5.95 $Y=0.74 $X2=0 $Y2=0
cc_428 N_A_83_260#_c_228_n N_X_c_969_n 0.00192131f $X=5.955 $Y=1.765 $X2=0 $Y2=0
cc_429 N_A_83_260#_M1038_g N_X_c_969_n 0.0050051f $X=6.38 $Y=0.74 $X2=0 $Y2=0
cc_430 N_A_83_260#_c_229_n N_X_c_969_n 0.00145998f $X=6.405 $Y=1.765 $X2=0 $Y2=0
cc_431 N_A_83_260#_c_206_n N_X_c_969_n 0.0297651f $X=7.505 $Y=1.665 $X2=0 $Y2=0
cc_432 N_A_83_260#_c_213_n N_X_c_969_n 0.0338654f $X=5.74 $Y=1.465 $X2=0 $Y2=0
cc_433 N_A_83_260#_c_214_n N_X_c_969_n 0.0339281f $X=6.665 $Y=1.465 $X2=0 $Y2=0
cc_434 N_A_83_260#_c_215_n N_X_c_969_n 0.0289688f $X=7.305 $Y=1.532 $X2=0 $Y2=0
cc_435 N_A_83_260#_c_230_n N_X_c_980_n 0.00186241f $X=6.855 $Y=1.765 $X2=0 $Y2=0
cc_436 N_A_83_260#_c_231_n N_X_c_980_n 0.0143315f $X=7.305 $Y=1.765 $X2=0 $Y2=0
cc_437 N_A_83_260#_c_232_n N_X_c_980_n 0.00389261f $X=8.03 $Y=2.815 $X2=0 $Y2=0
cc_438 N_A_83_260#_c_206_n N_X_c_980_n 0.0291863f $X=7.505 $Y=1.665 $X2=0 $Y2=0
cc_439 N_A_83_260#_c_207_n N_X_c_980_n 0.0344742f $X=7.505 $Y=1.665 $X2=0 $Y2=0
cc_440 N_A_83_260#_c_214_n N_X_c_980_n 0.0277768f $X=6.665 $Y=1.465 $X2=0 $Y2=0
cc_441 N_A_83_260#_c_215_n N_X_c_980_n 0.0213283f $X=7.305 $Y=1.532 $X2=0 $Y2=0
cc_442 N_A_83_260#_c_217_n N_X_c_1091_n 0.0120167f $X=0.955 $Y=1.765 $X2=0 $Y2=0
cc_443 N_A_83_260#_c_218_n N_X_c_1091_n 0.00712255f $X=1.405 $Y=1.765 $X2=0
+ $Y2=0
cc_444 N_A_83_260#_c_219_n N_X_c_1091_n 0.00977814f $X=1.855 $Y=1.765 $X2=0
+ $Y2=0
cc_445 N_A_83_260#_c_220_n N_X_c_1091_n 0.00701001f $X=2.355 $Y=1.765 $X2=0
+ $Y2=0
cc_446 N_A_83_260#_c_221_n N_X_c_1091_n 0.00839781f $X=2.805 $Y=1.765 $X2=0
+ $Y2=0
cc_447 N_A_83_260#_c_222_n N_X_c_1091_n 0.00684285f $X=3.255 $Y=1.765 $X2=0
+ $Y2=0
cc_448 N_A_83_260#_c_223_n N_X_c_1091_n 0.00822149f $X=3.705 $Y=1.765 $X2=0
+ $Y2=0
cc_449 N_A_83_260#_c_224_n N_X_c_1091_n 0.00712255f $X=4.155 $Y=1.765 $X2=0
+ $Y2=0
cc_450 N_A_83_260#_c_225_n N_X_c_1091_n 0.00670462f $X=4.605 $Y=1.765 $X2=0
+ $Y2=0
cc_451 N_A_83_260#_c_226_n N_X_c_1091_n 0.00697331f $X=5.055 $Y=1.765 $X2=0
+ $Y2=0
cc_452 N_A_83_260#_c_227_n N_X_c_1091_n 0.00815687f $X=5.505 $Y=1.765 $X2=0
+ $Y2=0
cc_453 N_A_83_260#_c_228_n N_X_c_1091_n 0.00822823f $X=5.955 $Y=1.765 $X2=0
+ $Y2=0
cc_454 N_A_83_260#_c_229_n N_X_c_1091_n 0.00795077f $X=6.405 $Y=1.765 $X2=0
+ $Y2=0
cc_455 N_A_83_260#_c_230_n N_X_c_1091_n 0.0083639f $X=6.855 $Y=1.765 $X2=0 $Y2=0
cc_456 N_A_83_260#_c_231_n N_X_c_1091_n 0.00273259f $X=7.305 $Y=1.765 $X2=0
+ $Y2=0
cc_457 N_A_83_260#_c_311_p N_X_c_1091_n 0.00516877f $X=7.59 $Y=2.035 $X2=0 $Y2=0
cc_458 N_A_83_260#_c_232_n N_X_c_1091_n 6.0059e-19 $X=8.03 $Y=2.815 $X2=0 $Y2=0
cc_459 N_A_83_260#_c_206_n N_X_c_1091_n 0.612349f $X=7.505 $Y=1.665 $X2=0 $Y2=0
cc_460 N_A_83_260#_c_207_n N_X_c_1091_n 8.80153e-19 $X=7.505 $Y=1.665 $X2=0
+ $Y2=0
cc_461 N_A_83_260#_c_208_n N_X_c_1091_n 0.00210155f $X=1.15 $Y=1.465 $X2=0 $Y2=0
cc_462 N_A_83_260#_c_209_n N_X_c_1091_n 0.00168006f $X=2.035 $Y=1.465 $X2=0
+ $Y2=0
cc_463 N_A_83_260#_c_210_n N_X_c_1091_n 0.00188729f $X=2.995 $Y=1.465 $X2=0
+ $Y2=0
cc_464 N_A_83_260#_c_211_n N_X_c_1091_n 0.00322453f $X=3.86 $Y=1.465 $X2=0 $Y2=0
cc_465 N_A_83_260#_c_212_n N_X_c_1091_n 0.00291335f $X=4.72 $Y=1.465 $X2=0 $Y2=0
cc_466 N_A_83_260#_c_213_n N_X_c_1091_n 0.00176418f $X=5.74 $Y=1.465 $X2=0 $Y2=0
cc_467 N_A_83_260#_c_214_n N_X_c_1091_n 0.00195696f $X=6.665 $Y=1.465 $X2=0
+ $Y2=0
cc_468 N_A_83_260#_c_215_n N_X_c_1091_n 0.00498224f $X=7.305 $Y=1.532 $X2=0
+ $Y2=0
cc_469 N_A_83_260#_c_224_n N_X_c_1118_n 0.00167853f $X=4.155 $Y=1.765 $X2=0
+ $Y2=0
cc_470 N_A_83_260#_c_225_n N_X_c_1118_n 0.00183229f $X=4.605 $Y=1.765 $X2=0
+ $Y2=0
cc_471 N_A_83_260#_c_226_n N_X_c_1118_n 5.42377e-19 $X=5.055 $Y=1.765 $X2=0
+ $Y2=0
cc_472 N_A_83_260#_c_206_n N_X_c_1118_n 0.00540615f $X=7.505 $Y=1.665 $X2=0
+ $Y2=0
cc_473 N_A_83_260#_c_215_n N_X_c_1118_n 0.00369434f $X=7.305 $Y=1.532 $X2=0
+ $Y2=0
cc_474 N_A_83_260#_c_223_n N_X_c_970_n 0.00100346f $X=3.705 $Y=1.765 $X2=0 $Y2=0
cc_475 N_A_83_260#_M1023_g N_X_c_970_n 0.00341074f $X=3.95 $Y=0.74 $X2=0 $Y2=0
cc_476 N_A_83_260#_c_224_n N_X_c_970_n 0.00281847f $X=4.155 $Y=1.765 $X2=0 $Y2=0
cc_477 N_A_83_260#_M1024_g N_X_c_970_n 0.00497263f $X=4.38 $Y=0.74 $X2=0 $Y2=0
cc_478 N_A_83_260#_c_225_n N_X_c_970_n 0.00243082f $X=4.605 $Y=1.765 $X2=0 $Y2=0
cc_479 N_A_83_260#_c_206_n N_X_c_970_n 0.0204733f $X=7.505 $Y=1.665 $X2=0 $Y2=0
cc_480 N_A_83_260#_c_211_n N_X_c_970_n 0.0337669f $X=3.86 $Y=1.465 $X2=0 $Y2=0
cc_481 N_A_83_260#_c_212_n N_X_c_970_n 0.0318624f $X=4.72 $Y=1.465 $X2=0 $Y2=0
cc_482 N_A_83_260#_c_215_n N_X_c_970_n 0.019992f $X=7.305 $Y=1.532 $X2=0 $Y2=0
cc_483 N_A_83_260#_c_198_n N_VGND_M1042_s 9.24827e-19 $X=7.94 $Y=1.095 $X2=0
+ $Y2=0
cc_484 N_A_83_260#_c_418_p N_VGND_M1042_s 8.63167e-19 $X=7.59 $Y=1.095 $X2=0
+ $Y2=0
cc_485 N_A_83_260#_c_200_n N_VGND_M1005_s 0.00176461f $X=8.8 $Y=1.095 $X2=0
+ $Y2=0
cc_486 N_A_83_260#_c_202_n N_VGND_M1012_s 0.00213667f $X=9.695 $Y=1.095 $X2=0
+ $Y2=0
cc_487 N_A_83_260#_M1003_g N_VGND_c_1214_n 0.00511162f $X=0.51 $Y=0.74 $X2=0
+ $Y2=0
cc_488 N_A_83_260#_M1003_g N_VGND_c_1215_n 6.09578e-19 $X=0.51 $Y=0.74 $X2=0
+ $Y2=0
cc_489 N_A_83_260#_M1004_g N_VGND_c_1215_n 0.0131166f $X=0.94 $Y=0.74 $X2=0
+ $Y2=0
cc_490 N_A_83_260#_M1008_g N_VGND_c_1215_n 0.00231293f $X=1.37 $Y=0.74 $X2=0
+ $Y2=0
cc_491 N_A_83_260#_c_206_n N_VGND_c_1215_n 0.00144039f $X=7.505 $Y=1.665 $X2=0
+ $Y2=0
cc_492 N_A_83_260#_c_208_n N_VGND_c_1215_n 0.0241312f $X=1.15 $Y=1.465 $X2=0
+ $Y2=0
cc_493 N_A_83_260#_c_215_n N_VGND_c_1215_n 7.91474e-19 $X=7.305 $Y=1.532 $X2=0
+ $Y2=0
cc_494 N_A_83_260#_M1009_g N_VGND_c_1216_n 0.00216549f $X=1.8 $Y=0.74 $X2=0
+ $Y2=0
cc_495 N_A_83_260#_M1010_g N_VGND_c_1216_n 0.00335886f $X=2.23 $Y=0.74 $X2=0
+ $Y2=0
cc_496 N_A_83_260#_c_206_n N_VGND_c_1216_n 0.00100477f $X=7.505 $Y=1.665 $X2=0
+ $Y2=0
cc_497 N_A_83_260#_c_209_n N_VGND_c_1216_n 0.0167867f $X=2.035 $Y=1.465 $X2=0
+ $Y2=0
cc_498 N_A_83_260#_c_215_n N_VGND_c_1216_n 7.91474e-19 $X=7.305 $Y=1.532 $X2=0
+ $Y2=0
cc_499 N_A_83_260#_M1014_g N_VGND_c_1217_n 0.0027473f $X=2.66 $Y=0.74 $X2=0
+ $Y2=0
cc_500 N_A_83_260#_M1016_g N_VGND_c_1217_n 0.00276906f $X=3.09 $Y=0.74 $X2=0
+ $Y2=0
cc_501 N_A_83_260#_c_206_n N_VGND_c_1217_n 0.0025197f $X=7.505 $Y=1.665 $X2=0
+ $Y2=0
cc_502 N_A_83_260#_c_210_n N_VGND_c_1217_n 0.00578402f $X=2.995 $Y=1.465 $X2=0
+ $Y2=0
cc_503 N_A_83_260#_c_215_n N_VGND_c_1217_n 0.00148272f $X=7.305 $Y=1.532 $X2=0
+ $Y2=0
cc_504 N_A_83_260#_M1019_g N_VGND_c_1218_n 0.00321813f $X=3.52 $Y=0.74 $X2=0
+ $Y2=0
cc_505 N_A_83_260#_M1023_g N_VGND_c_1218_n 0.00322379f $X=3.95 $Y=0.74 $X2=0
+ $Y2=0
cc_506 N_A_83_260#_c_206_n N_VGND_c_1218_n 8.11739e-19 $X=7.505 $Y=1.665 $X2=0
+ $Y2=0
cc_507 N_A_83_260#_c_211_n N_VGND_c_1218_n 0.0134172f $X=3.86 $Y=1.465 $X2=0
+ $Y2=0
cc_508 N_A_83_260#_c_215_n N_VGND_c_1218_n 7.8229e-19 $X=7.305 $Y=1.532 $X2=0
+ $Y2=0
cc_509 N_A_83_260#_M1023_g N_VGND_c_1219_n 0.00434272f $X=3.95 $Y=0.74 $X2=0
+ $Y2=0
cc_510 N_A_83_260#_M1024_g N_VGND_c_1219_n 0.00371957f $X=4.38 $Y=0.74 $X2=0
+ $Y2=0
cc_511 N_A_83_260#_M1024_g N_VGND_c_1220_n 0.00931981f $X=4.38 $Y=0.74 $X2=0
+ $Y2=0
cc_512 N_A_83_260#_M1032_g N_VGND_c_1220_n 0.00663936f $X=4.95 $Y=0.74 $X2=0
+ $Y2=0
cc_513 N_A_83_260#_c_206_n N_VGND_c_1220_n 0.00135125f $X=7.505 $Y=1.665 $X2=0
+ $Y2=0
cc_514 N_A_83_260#_c_212_n N_VGND_c_1220_n 0.0224942f $X=4.72 $Y=1.465 $X2=0
+ $Y2=0
cc_515 N_A_83_260#_c_215_n N_VGND_c_1220_n 0.00180013f $X=7.305 $Y=1.532 $X2=0
+ $Y2=0
cc_516 N_A_83_260#_M1032_g N_VGND_c_1221_n 0.00461464f $X=4.95 $Y=0.74 $X2=0
+ $Y2=0
cc_517 N_A_83_260#_M1034_g N_VGND_c_1221_n 0.00434272f $X=5.38 $Y=0.74 $X2=0
+ $Y2=0
cc_518 N_A_83_260#_M1034_g N_VGND_c_1222_n 0.00602841f $X=5.38 $Y=0.74 $X2=0
+ $Y2=0
cc_519 N_A_83_260#_M1035_g N_VGND_c_1222_n 0.00602841f $X=5.95 $Y=0.74 $X2=0
+ $Y2=0
cc_520 N_A_83_260#_c_206_n N_VGND_c_1222_n 0.00419098f $X=7.505 $Y=1.665 $X2=0
+ $Y2=0
cc_521 N_A_83_260#_c_213_n N_VGND_c_1222_n 0.0133056f $X=5.74 $Y=1.465 $X2=0
+ $Y2=0
cc_522 N_A_83_260#_c_215_n N_VGND_c_1222_n 0.00310051f $X=7.305 $Y=1.532 $X2=0
+ $Y2=0
cc_523 N_A_83_260#_M1038_g N_VGND_c_1223_n 0.00666821f $X=6.38 $Y=0.74 $X2=0
+ $Y2=0
cc_524 N_A_83_260#_M1041_g N_VGND_c_1223_n 0.00657867f $X=6.95 $Y=0.74 $X2=0
+ $Y2=0
cc_525 N_A_83_260#_c_206_n N_VGND_c_1223_n 0.00231384f $X=7.505 $Y=1.665 $X2=0
+ $Y2=0
cc_526 N_A_83_260#_c_214_n N_VGND_c_1223_n 0.0254679f $X=6.665 $Y=1.465 $X2=0
+ $Y2=0
cc_527 N_A_83_260#_c_215_n N_VGND_c_1223_n 0.00189844f $X=7.305 $Y=1.532 $X2=0
+ $Y2=0
cc_528 N_A_83_260#_M1041_g N_VGND_c_1224_n 0.00434272f $X=6.95 $Y=0.74 $X2=0
+ $Y2=0
cc_529 N_A_83_260#_M1042_g N_VGND_c_1224_n 0.00383152f $X=7.38 $Y=0.74 $X2=0
+ $Y2=0
cc_530 N_A_83_260#_M1041_g N_VGND_c_1225_n 5.17822e-19 $X=6.95 $Y=0.74 $X2=0
+ $Y2=0
cc_531 N_A_83_260#_M1042_g N_VGND_c_1225_n 0.0107288f $X=7.38 $Y=0.74 $X2=0
+ $Y2=0
cc_532 N_A_83_260#_c_198_n N_VGND_c_1225_n 0.00890916f $X=7.94 $Y=1.095 $X2=0
+ $Y2=0
cc_533 N_A_83_260#_c_418_p N_VGND_c_1225_n 0.00902191f $X=7.59 $Y=1.095 $X2=0
+ $Y2=0
cc_534 N_A_83_260#_c_199_n N_VGND_c_1225_n 0.0182488f $X=8.025 $Y=0.515 $X2=0
+ $Y2=0
cc_535 N_A_83_260#_c_199_n N_VGND_c_1226_n 0.0182488f $X=8.025 $Y=0.515 $X2=0
+ $Y2=0
cc_536 N_A_83_260#_c_200_n N_VGND_c_1226_n 0.0170777f $X=8.8 $Y=1.095 $X2=0
+ $Y2=0
cc_537 N_A_83_260#_c_201_n N_VGND_c_1226_n 0.0182488f $X=8.885 $Y=0.515 $X2=0
+ $Y2=0
cc_538 N_A_83_260#_c_201_n N_VGND_c_1227_n 0.0182488f $X=8.885 $Y=0.515 $X2=0
+ $Y2=0
cc_539 N_A_83_260#_c_202_n N_VGND_c_1227_n 0.0181391f $X=9.695 $Y=1.095 $X2=0
+ $Y2=0
cc_540 N_A_83_260#_c_203_n N_VGND_c_1227_n 0.00131301f $X=9.78 $Y=0.515 $X2=0
+ $Y2=0
cc_541 N_A_83_260#_c_202_n N_VGND_c_1229_n 0.00540984f $X=9.695 $Y=1.095 $X2=0
+ $Y2=0
cc_542 N_A_83_260#_c_203_n N_VGND_c_1229_n 0.0255227f $X=9.78 $Y=0.515 $X2=0
+ $Y2=0
cc_543 N_A_83_260#_M1008_g N_VGND_c_1230_n 0.00461464f $X=1.37 $Y=0.74 $X2=0
+ $Y2=0
cc_544 N_A_83_260#_M1009_g N_VGND_c_1230_n 0.00461464f $X=1.8 $Y=0.74 $X2=0
+ $Y2=0
cc_545 N_A_83_260#_M1010_g N_VGND_c_1232_n 0.00461464f $X=2.23 $Y=0.74 $X2=0
+ $Y2=0
cc_546 N_A_83_260#_M1014_g N_VGND_c_1232_n 0.00434272f $X=2.66 $Y=0.74 $X2=0
+ $Y2=0
cc_547 N_A_83_260#_M1016_g N_VGND_c_1234_n 0.00461464f $X=3.09 $Y=0.74 $X2=0
+ $Y2=0
cc_548 N_A_83_260#_M1019_g N_VGND_c_1234_n 0.00422942f $X=3.52 $Y=0.74 $X2=0
+ $Y2=0
cc_549 N_A_83_260#_M1035_g N_VGND_c_1236_n 0.00434272f $X=5.95 $Y=0.74 $X2=0
+ $Y2=0
cc_550 N_A_83_260#_M1038_g N_VGND_c_1236_n 0.00434272f $X=6.38 $Y=0.74 $X2=0
+ $Y2=0
cc_551 N_A_83_260#_M1003_g N_VGND_c_1238_n 0.00434272f $X=0.51 $Y=0.74 $X2=0
+ $Y2=0
cc_552 N_A_83_260#_M1004_g N_VGND_c_1238_n 0.00383152f $X=0.94 $Y=0.74 $X2=0
+ $Y2=0
cc_553 N_A_83_260#_c_199_n N_VGND_c_1239_n 0.00749631f $X=8.025 $Y=0.515 $X2=0
+ $Y2=0
cc_554 N_A_83_260#_c_201_n N_VGND_c_1240_n 0.00749631f $X=8.885 $Y=0.515 $X2=0
+ $Y2=0
cc_555 N_A_83_260#_c_203_n N_VGND_c_1241_n 0.011066f $X=9.78 $Y=0.515 $X2=0
+ $Y2=0
cc_556 N_A_83_260#_M1003_g N_VGND_c_1248_n 0.00823992f $X=0.51 $Y=0.74 $X2=0
+ $Y2=0
cc_557 N_A_83_260#_M1004_g N_VGND_c_1248_n 0.0075754f $X=0.94 $Y=0.74 $X2=0
+ $Y2=0
cc_558 N_A_83_260#_M1008_g N_VGND_c_1248_n 0.00907324f $X=1.37 $Y=0.74 $X2=0
+ $Y2=0
cc_559 N_A_83_260#_M1009_g N_VGND_c_1248_n 0.00907549f $X=1.8 $Y=0.74 $X2=0
+ $Y2=0
cc_560 N_A_83_260#_M1010_g N_VGND_c_1248_n 0.00908333f $X=2.23 $Y=0.74 $X2=0
+ $Y2=0
cc_561 N_A_83_260#_M1014_g N_VGND_c_1248_n 0.00820284f $X=2.66 $Y=0.74 $X2=0
+ $Y2=0
cc_562 N_A_83_260#_M1016_g N_VGND_c_1248_n 0.00908333f $X=3.09 $Y=0.74 $X2=0
+ $Y2=0
cc_563 N_A_83_260#_M1019_g N_VGND_c_1248_n 0.00783597f $X=3.52 $Y=0.74 $X2=0
+ $Y2=0
cc_564 N_A_83_260#_M1023_g N_VGND_c_1248_n 0.00820284f $X=3.95 $Y=0.74 $X2=0
+ $Y2=0
cc_565 N_A_83_260#_M1024_g N_VGND_c_1248_n 0.00620726f $X=4.38 $Y=0.74 $X2=0
+ $Y2=0
cc_566 N_A_83_260#_M1032_g N_VGND_c_1248_n 0.00909342f $X=4.95 $Y=0.74 $X2=0
+ $Y2=0
cc_567 N_A_83_260#_M1034_g N_VGND_c_1248_n 0.00821294f $X=5.38 $Y=0.74 $X2=0
+ $Y2=0
cc_568 N_A_83_260#_M1035_g N_VGND_c_1248_n 0.00821294f $X=5.95 $Y=0.74 $X2=0
+ $Y2=0
cc_569 N_A_83_260#_M1038_g N_VGND_c_1248_n 0.00821294f $X=6.38 $Y=0.74 $X2=0
+ $Y2=0
cc_570 N_A_83_260#_M1041_g N_VGND_c_1248_n 0.00821294f $X=6.95 $Y=0.74 $X2=0
+ $Y2=0
cc_571 N_A_83_260#_M1042_g N_VGND_c_1248_n 0.0075754f $X=7.38 $Y=0.74 $X2=0
+ $Y2=0
cc_572 N_A_83_260#_c_199_n N_VGND_c_1248_n 0.0062048f $X=8.025 $Y=0.515 $X2=0
+ $Y2=0
cc_573 N_A_83_260#_c_201_n N_VGND_c_1248_n 0.0062048f $X=8.885 $Y=0.515 $X2=0
+ $Y2=0
cc_574 N_A_83_260#_c_203_n N_VGND_c_1248_n 0.00915947f $X=9.78 $Y=0.515 $X2=0
+ $Y2=0
cc_575 N_A_c_647_n N_VPWR_c_774_n 0.00671059f $X=7.805 $Y=1.765 $X2=0 $Y2=0
cc_576 N_A_c_647_n N_VPWR_c_775_n 0.00445602f $X=7.805 $Y=1.765 $X2=0 $Y2=0
cc_577 N_A_c_648_n N_VPWR_c_775_n 0.00445602f $X=8.255 $Y=1.765 $X2=0 $Y2=0
cc_578 N_A_c_648_n N_VPWR_c_776_n 0.00486623f $X=8.255 $Y=1.765 $X2=0 $Y2=0
cc_579 N_A_c_649_n N_VPWR_c_776_n 0.00486623f $X=8.705 $Y=1.765 $X2=0 $Y2=0
cc_580 N_A_c_649_n N_VPWR_c_777_n 0.00445602f $X=8.705 $Y=1.765 $X2=0 $Y2=0
cc_581 N_A_c_650_n N_VPWR_c_777_n 0.00445602f $X=9.155 $Y=1.765 $X2=0 $Y2=0
cc_582 N_A_c_650_n N_VPWR_c_778_n 0.00486623f $X=9.155 $Y=1.765 $X2=0 $Y2=0
cc_583 N_A_c_651_n N_VPWR_c_778_n 0.00486623f $X=9.605 $Y=1.765 $X2=0 $Y2=0
cc_584 N_A_c_652_n N_VPWR_c_780_n 0.00831454f $X=10.055 $Y=1.765 $X2=0 $Y2=0
cc_585 A N_VPWR_c_780_n 0.0211447f $X=10.235 $Y=1.58 $X2=0 $Y2=0
cc_586 N_A_c_651_n N_VPWR_c_797_n 0.00445602f $X=9.605 $Y=1.765 $X2=0 $Y2=0
cc_587 N_A_c_652_n N_VPWR_c_797_n 0.00445602f $X=10.055 $Y=1.765 $X2=0 $Y2=0
cc_588 N_A_c_647_n N_VPWR_c_764_n 0.00857432f $X=7.805 $Y=1.765 $X2=0 $Y2=0
cc_589 N_A_c_648_n N_VPWR_c_764_n 0.00857589f $X=8.255 $Y=1.765 $X2=0 $Y2=0
cc_590 N_A_c_649_n N_VPWR_c_764_n 0.00857589f $X=8.705 $Y=1.765 $X2=0 $Y2=0
cc_591 N_A_c_650_n N_VPWR_c_764_n 0.00857589f $X=9.155 $Y=1.765 $X2=0 $Y2=0
cc_592 N_A_c_651_n N_VPWR_c_764_n 0.00857589f $X=9.605 $Y=1.765 $X2=0 $Y2=0
cc_593 N_A_c_652_n N_VPWR_c_764_n 0.00861084f $X=10.055 $Y=1.765 $X2=0 $Y2=0
cc_594 N_A_c_647_n N_X_c_980_n 9.59128e-19 $X=7.805 $Y=1.765 $X2=0 $Y2=0
cc_595 N_A_M1002_g N_VGND_c_1225_n 0.010609f $X=7.81 $Y=0.74 $X2=0 $Y2=0
cc_596 N_A_M1005_g N_VGND_c_1225_n 4.71636e-19 $X=8.24 $Y=0.74 $X2=0 $Y2=0
cc_597 N_A_M1002_g N_VGND_c_1226_n 4.71636e-19 $X=7.81 $Y=0.74 $X2=0 $Y2=0
cc_598 N_A_M1005_g N_VGND_c_1226_n 0.0106755f $X=8.24 $Y=0.74 $X2=0 $Y2=0
cc_599 N_A_M1011_g N_VGND_c_1226_n 0.0106755f $X=8.67 $Y=0.74 $X2=0 $Y2=0
cc_600 N_A_M1012_g N_VGND_c_1226_n 4.71636e-19 $X=9.1 $Y=0.74 $X2=0 $Y2=0
cc_601 N_A_M1011_g N_VGND_c_1227_n 4.71636e-19 $X=8.67 $Y=0.74 $X2=0 $Y2=0
cc_602 N_A_M1012_g N_VGND_c_1227_n 0.0105121f $X=9.1 $Y=0.74 $X2=0 $Y2=0
cc_603 N_A_M1013_g N_VGND_c_1227_n 0.0024857f $X=9.565 $Y=0.74 $X2=0 $Y2=0
cc_604 N_A_M1013_g N_VGND_c_1229_n 5.35525e-19 $X=9.565 $Y=0.74 $X2=0 $Y2=0
cc_605 N_A_M1043_g N_VGND_c_1229_n 0.015186f $X=10.065 $Y=0.74 $X2=0 $Y2=0
cc_606 A N_VGND_c_1229_n 0.023753f $X=10.235 $Y=1.58 $X2=0 $Y2=0
cc_607 N_A_M1002_g N_VGND_c_1239_n 0.00383152f $X=7.81 $Y=0.74 $X2=0 $Y2=0
cc_608 N_A_M1005_g N_VGND_c_1239_n 0.00383152f $X=8.24 $Y=0.74 $X2=0 $Y2=0
cc_609 N_A_M1011_g N_VGND_c_1240_n 0.00383152f $X=8.67 $Y=0.74 $X2=0 $Y2=0
cc_610 N_A_M1012_g N_VGND_c_1240_n 0.00383152f $X=9.1 $Y=0.74 $X2=0 $Y2=0
cc_611 N_A_M1013_g N_VGND_c_1241_n 0.00461464f $X=9.565 $Y=0.74 $X2=0 $Y2=0
cc_612 N_A_M1043_g N_VGND_c_1241_n 0.00383152f $X=10.065 $Y=0.74 $X2=0 $Y2=0
cc_613 N_A_M1002_g N_VGND_c_1248_n 0.0075754f $X=7.81 $Y=0.74 $X2=0 $Y2=0
cc_614 N_A_M1005_g N_VGND_c_1248_n 0.0075754f $X=8.24 $Y=0.74 $X2=0 $Y2=0
cc_615 N_A_M1011_g N_VGND_c_1248_n 0.0075754f $X=8.67 $Y=0.74 $X2=0 $Y2=0
cc_616 N_A_M1012_g N_VGND_c_1248_n 0.0075754f $X=9.1 $Y=0.74 $X2=0 $Y2=0
cc_617 N_A_M1013_g N_VGND_c_1248_n 0.00908323f $X=9.565 $Y=0.74 $X2=0 $Y2=0
cc_618 N_A_M1043_g N_VGND_c_1248_n 0.00758198f $X=10.065 $Y=0.74 $X2=0 $Y2=0
cc_619 N_VPWR_c_789_n N_X_c_971_n 0.014552f $X=4.745 $Y=3.33 $X2=0 $Y2=0
cc_620 N_VPWR_c_764_n N_X_c_971_n 0.0119791f $X=10.32 $Y=3.33 $X2=0 $Y2=0
cc_621 N_VPWR_c_766_n N_X_c_967_n 0.0761208f $X=0.28 $Y=1.985 $X2=0 $Y2=0
cc_622 N_VPWR_c_767_n N_X_c_967_n 0.0507192f $X=1.18 $Y=2.13 $X2=0 $Y2=0
cc_623 N_VPWR_c_781_n N_X_c_967_n 0.0112323f $X=1.095 $Y=3.33 $X2=0 $Y2=0
cc_624 N_VPWR_c_764_n N_X_c_967_n 0.00925249f $X=10.32 $Y=3.33 $X2=0 $Y2=0
cc_625 N_VPWR_c_767_n N_X_c_968_n 0.0634465f $X=1.18 $Y=2.13 $X2=0 $Y2=0
cc_626 N_VPWR_c_768_n N_X_c_968_n 0.0317846f $X=2.13 $Y=2.13 $X2=0 $Y2=0
cc_627 N_VPWR_c_783_n N_X_c_968_n 0.0112472f $X=1.965 $Y=3.33 $X2=0 $Y2=0
cc_628 N_VPWR_c_764_n N_X_c_968_n 0.00927661f $X=10.32 $Y=3.33 $X2=0 $Y2=0
cc_629 N_VPWR_c_768_n N_X_c_976_n 0.0651544f $X=2.13 $Y=2.13 $X2=0 $Y2=0
cc_630 N_VPWR_c_769_n N_X_c_976_n 0.0280596f $X=3.03 $Y=2.13 $X2=0 $Y2=0
cc_631 N_VPWR_c_785_n N_X_c_976_n 0.0114703f $X=2.945 $Y=3.33 $X2=0 $Y2=0
cc_632 N_VPWR_c_764_n N_X_c_976_n 0.00946127f $X=10.32 $Y=3.33 $X2=0 $Y2=0
cc_633 N_VPWR_c_769_n N_X_c_977_n 0.0647726f $X=3.03 $Y=2.13 $X2=0 $Y2=0
cc_634 N_VPWR_c_770_n N_X_c_977_n 0.0507192f $X=3.93 $Y=2.13 $X2=0 $Y2=0
cc_635 N_VPWR_c_787_n N_X_c_977_n 0.0112323f $X=3.845 $Y=3.33 $X2=0 $Y2=0
cc_636 N_VPWR_c_764_n N_X_c_977_n 0.00925249f $X=10.32 $Y=3.33 $X2=0 $Y2=0
cc_637 N_VPWR_c_771_n N_X_c_978_n 0.0640463f $X=4.83 $Y=2.13 $X2=0 $Y2=0
cc_638 N_VPWR_c_772_n N_X_c_978_n 0.0313576f $X=5.73 $Y=2.13 $X2=0 $Y2=0
cc_639 N_VPWR_c_791_n N_X_c_978_n 0.0130321f $X=5.645 $Y=3.33 $X2=0 $Y2=0
cc_640 N_VPWR_c_764_n N_X_c_978_n 0.0107539f $X=10.32 $Y=3.33 $X2=0 $Y2=0
cc_641 N_VPWR_c_772_n N_X_c_969_n 0.0303219f $X=5.73 $Y=2.13 $X2=0 $Y2=0
cc_642 N_VPWR_c_773_n N_X_c_969_n 0.0622757f $X=6.63 $Y=2.13 $X2=0 $Y2=0
cc_643 N_VPWR_c_793_n N_X_c_969_n 0.0119584f $X=6.545 $Y=3.33 $X2=0 $Y2=0
cc_644 N_VPWR_c_764_n N_X_c_969_n 0.00989813f $X=10.32 $Y=3.33 $X2=0 $Y2=0
cc_645 N_VPWR_c_773_n N_X_c_980_n 0.0284839f $X=6.63 $Y=2.13 $X2=0 $Y2=0
cc_646 N_VPWR_c_774_n N_X_c_980_n 0.0455435f $X=7.53 $Y=2.455 $X2=0 $Y2=0
cc_647 N_VPWR_c_795_n N_X_c_980_n 0.0116935f $X=7.445 $Y=3.33 $X2=0 $Y2=0
cc_648 N_VPWR_c_764_n N_X_c_980_n 0.00964594f $X=10.32 $Y=3.33 $X2=0 $Y2=0
cc_649 N_VPWR_M1007_d N_X_c_1091_n 0.00655748f $X=1.03 $Y=1.84 $X2=0 $Y2=0
cc_650 N_VPWR_M1017_d N_X_c_1091_n 0.00571508f $X=1.93 $Y=1.84 $X2=0 $Y2=0
cc_651 N_VPWR_M1020_d N_X_c_1091_n 0.0065703f $X=2.88 $Y=1.84 $X2=0 $Y2=0
cc_652 N_VPWR_M1022_d N_X_c_1091_n 0.00655491f $X=3.78 $Y=1.84 $X2=0 $Y2=0
cc_653 N_VPWR_M1026_d N_X_c_1091_n 0.00676008f $X=4.68 $Y=1.84 $X2=0 $Y2=0
cc_654 N_VPWR_M1029_d N_X_c_1091_n 0.00646217f $X=5.58 $Y=1.84 $X2=0 $Y2=0
cc_655 N_VPWR_M1033_d N_X_c_1091_n 0.00651901f $X=6.48 $Y=1.84 $X2=0 $Y2=0
cc_656 N_VPWR_c_766_n N_X_c_1091_n 0.00164279f $X=0.28 $Y=1.985 $X2=0 $Y2=0
cc_657 N_VPWR_c_767_n N_X_c_1091_n 0.0180973f $X=1.18 $Y=2.13 $X2=0 $Y2=0
cc_658 N_VPWR_c_768_n N_X_c_1091_n 0.0249156f $X=2.13 $Y=2.13 $X2=0 $Y2=0
cc_659 N_VPWR_c_769_n N_X_c_1091_n 0.0179781f $X=3.03 $Y=2.13 $X2=0 $Y2=0
cc_660 N_VPWR_c_770_n N_X_c_1091_n 0.0180973f $X=3.93 $Y=2.13 $X2=0 $Y2=0
cc_661 N_VPWR_c_771_n N_X_c_1091_n 0.0181811f $X=4.83 $Y=2.13 $X2=0 $Y2=0
cc_662 N_VPWR_c_772_n N_X_c_1091_n 0.0181266f $X=5.73 $Y=2.13 $X2=0 $Y2=0
cc_663 N_VPWR_c_773_n N_X_c_1091_n 0.0181154f $X=6.63 $Y=2.13 $X2=0 $Y2=0
cc_664 N_VPWR_c_770_n N_X_c_1118_n 0.0644893f $X=3.93 $Y=2.13 $X2=0 $Y2=0
cc_665 N_VPWR_c_771_n N_X_c_1118_n 0.0644893f $X=4.83 $Y=2.13 $X2=0 $Y2=0
cc_666 N_X_c_967_n N_VGND_c_1214_n 0.0283292f $X=0.725 $Y=0.515 $X2=0 $Y2=0
cc_667 N_X_c_967_n N_VGND_c_1215_n 0.0295974f $X=0.725 $Y=0.515 $X2=0 $Y2=0
cc_668 N_X_c_968_n N_VGND_c_1215_n 0.00295309f $X=1.585 $Y=0.515 $X2=0 $Y2=0
cc_669 N_X_c_954_n N_VGND_c_1216_n 0.00232335f $X=2.445 $Y=0.515 $X2=0 $Y2=0
cc_670 N_X_c_968_n N_VGND_c_1216_n 0.00293065f $X=1.585 $Y=0.515 $X2=0 $Y2=0
cc_671 N_X_c_954_n N_VGND_c_1217_n 0.0237333f $X=2.445 $Y=0.515 $X2=0 $Y2=0
cc_672 N_X_c_955_n N_VGND_c_1217_n 0.00109788f $X=3.305 $Y=0.515 $X2=0 $Y2=0
cc_673 N_X_c_955_n N_VGND_c_1218_n 0.0296111f $X=3.305 $Y=0.515 $X2=0 $Y2=0
cc_674 N_X_c_956_n N_VGND_c_1218_n 0.02996f $X=4.165 $Y=0.515 $X2=0 $Y2=0
cc_675 N_X_c_956_n N_VGND_c_1219_n 0.0167819f $X=4.165 $Y=0.515 $X2=0 $Y2=0
cc_676 N_X_c_956_n N_VGND_c_1220_n 0.0604257f $X=4.165 $Y=0.515 $X2=0 $Y2=0
cc_677 N_X_c_957_n N_VGND_c_1220_n 0.0027108f $X=5.165 $Y=0.515 $X2=0 $Y2=0
cc_678 N_X_c_957_n N_VGND_c_1221_n 0.0130022f $X=5.165 $Y=0.515 $X2=0 $Y2=0
cc_679 N_X_c_957_n N_VGND_c_1222_n 0.0260557f $X=5.165 $Y=0.515 $X2=0 $Y2=0
cc_680 N_X_c_958_n N_VGND_c_1222_n 0.0264558f $X=6.165 $Y=0.515 $X2=0 $Y2=0
cc_681 N_X_c_958_n N_VGND_c_1223_n 0.0308109f $X=6.165 $Y=0.515 $X2=0 $Y2=0
cc_682 N_X_c_959_n N_VGND_c_1223_n 3.89769e-19 $X=7.125 $Y=1.125 $X2=0 $Y2=0
cc_683 N_X_c_960_n N_VGND_c_1223_n 0.0292056f $X=7.165 $Y=0.515 $X2=0 $Y2=0
cc_684 N_X_c_960_n N_VGND_c_1224_n 0.0109942f $X=7.165 $Y=0.515 $X2=0 $Y2=0
cc_685 N_X_c_960_n N_VGND_c_1225_n 0.0182902f $X=7.165 $Y=0.515 $X2=0 $Y2=0
cc_686 N_X_c_968_n N_VGND_c_1230_n 0.0112891f $X=1.585 $Y=0.515 $X2=0 $Y2=0
cc_687 N_X_c_954_n N_VGND_c_1232_n 0.0116636f $X=2.445 $Y=0.515 $X2=0 $Y2=0
cc_688 N_X_c_955_n N_VGND_c_1234_n 0.0114106f $X=3.305 $Y=0.515 $X2=0 $Y2=0
cc_689 N_X_c_958_n N_VGND_c_1236_n 0.0144922f $X=6.165 $Y=0.515 $X2=0 $Y2=0
cc_690 N_X_c_967_n N_VGND_c_1238_n 0.0112174f $X=0.725 $Y=0.515 $X2=0 $Y2=0
cc_691 N_X_c_954_n N_VGND_c_1248_n 0.00959771f $X=2.445 $Y=0.515 $X2=0 $Y2=0
cc_692 N_X_c_955_n N_VGND_c_1248_n 0.00936481f $X=3.305 $Y=0.515 $X2=0 $Y2=0
cc_693 N_X_c_956_n N_VGND_c_1248_n 0.0136487f $X=4.165 $Y=0.515 $X2=0 $Y2=0
cc_694 N_X_c_957_n N_VGND_c_1248_n 0.0107057f $X=5.165 $Y=0.515 $X2=0 $Y2=0
cc_695 N_X_c_958_n N_VGND_c_1248_n 0.0118826f $X=6.165 $Y=0.515 $X2=0 $Y2=0
cc_696 N_X_c_960_n N_VGND_c_1248_n 0.00904371f $X=7.165 $Y=0.515 $X2=0 $Y2=0
cc_697 N_X_c_967_n N_VGND_c_1248_n 0.00922837f $X=0.725 $Y=0.515 $X2=0 $Y2=0
cc_698 N_X_c_968_n N_VGND_c_1248_n 0.00934413f $X=1.585 $Y=0.515 $X2=0 $Y2=0
