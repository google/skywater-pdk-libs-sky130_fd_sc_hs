* File: sky130_fd_sc_hs__dfsbp_2.pex.spice
* Created: Thu Aug 27 20:39:11 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HS__DFSBP_2%D 2 4 7 9 11 12 13 17 18 21
c35 18 0 8.44909e-20 $X=0.64 $Y=1.145
r36 21 23 39.7991 $w=3.9e-07 $l=1.65e-07 $layer=POLY_cond $X=0.61 $Y=1.825
+ $X2=0.61 $Y2=1.99
r37 21 22 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=0.64
+ $Y=1.825 $X2=0.64 $Y2=1.825
r38 17 19 45.456 $w=3.9e-07 $l=1.65e-07 $layer=POLY_cond $X=0.61 $Y=1.145
+ $X2=0.61 $Y2=0.98
r39 17 18 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=0.64
+ $Y=1.145 $X2=0.64 $Y2=1.145
r40 13 22 5.5876 $w=3.28e-07 $l=1.6e-07 $layer=LI1_cond $X=0.64 $Y=1.665
+ $X2=0.64 $Y2=1.825
r41 12 13 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=0.64 $Y=1.295
+ $X2=0.64 $Y2=1.665
r42 12 18 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=0.64 $Y=1.295
+ $X2=0.64 $Y2=1.145
r43 9 11 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=0.505 $Y=2.465
+ $X2=0.505 $Y2=2.75
r44 7 19 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=0.495 $Y=0.58 $X2=0.495
+ $Y2=0.98
r45 4 9 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=0.505 $Y=2.375 $X2=0.505
+ $Y2=2.465
r46 4 23 149.653 $w=1.8e-07 $l=3.85e-07 $layer=POLY_cond $X=0.505 $Y=2.375
+ $X2=0.505 $Y2=1.99
r47 2 21 4.27811 $w=3.9e-07 $l=3e-08 $layer=POLY_cond $X=0.61 $Y=1.795 $X2=0.61
+ $Y2=1.825
r48 1 17 4.27811 $w=3.9e-07 $l=3e-08 $layer=POLY_cond $X=0.61 $Y=1.175 $X2=0.61
+ $Y2=1.145
r49 1 2 88.4142 $w=3.9e-07 $l=6.2e-07 $layer=POLY_cond $X=0.61 $Y=1.175 $X2=0.61
+ $Y2=1.795
.ends

.subckt PM_SKY130_FD_SC_HS__DFSBP_2%CLK 1 3 4 6 7
c33 4 0 2.24304e-19 $X=1.515 $Y=1.715
r34 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.465
+ $Y=1.385 $X2=1.465 $Y2=1.385
r35 7 11 6.69663 $w=3.68e-07 $l=2.15e-07 $layer=LI1_cond $X=1.68 $Y=1.365
+ $X2=1.465 $Y2=1.365
r36 4 10 67.1335 $w=2.8e-07 $l=3.54119e-07 $layer=POLY_cond $X=1.515 $Y=1.715
+ $X2=1.465 $Y2=1.385
r37 4 6 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.515 $Y=1.715
+ $X2=1.515 $Y2=2.35
r38 1 10 38.7299 $w=2.8e-07 $l=1.74714e-07 $layer=POLY_cond $X=1.485 $Y=1.22
+ $X2=1.465 $Y2=1.385
r39 1 3 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.485 $Y=1.22 $X2=1.485
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HS__DFSBP_2%A_398_74# 1 2 7 8 9 11 12 16 20 21 23 26 30
+ 32 33 34 35 38 45 46 49 50 53 54 55 57 58 59 61 63 64 65 68 69 73 74 77 79 86
c275 77 0 2.30667e-19 $X=7.415 $Y=2.185
c276 74 0 8.86437e-20 $X=6.71 $Y=1.285
c277 59 0 1.18171e-19 $X=5.53 $Y=2.275
c278 58 0 1.74055e-19 $X=6.33 $Y=2.275
r279 77 79 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=7.415 $Y=2.185
+ $X2=7.415 $Y2=2.02
r280 77 78 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.415
+ $Y=2.185 $X2=7.415 $Y2=2.185
r281 74 86 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.71 $Y=1.285
+ $X2=6.71 $Y2=1.12
r282 73 74 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.71
+ $Y=1.285 $X2=6.71 $Y2=1.285
r283 70 73 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=6.415 $Y=1.285
+ $X2=6.71 $Y2=1.285
r284 66 79 102.428 $w=1.68e-07 $l=1.57e-06 $layer=LI1_cond $X=7.47 $Y=0.45
+ $X2=7.47 $Y2=2.02
r285 64 66 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.385 $Y=0.365
+ $X2=7.47 $Y2=0.45
r286 64 65 57.738 $w=1.68e-07 $l=8.85e-07 $layer=LI1_cond $X=7.385 $Y=0.365
+ $X2=6.5 $Y2=0.365
r287 62 70 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.415 $Y=1.45
+ $X2=6.415 $Y2=1.285
r288 62 63 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=6.415 $Y=1.45
+ $X2=6.415 $Y2=2.19
r289 61 70 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.415 $Y=1.12
+ $X2=6.415 $Y2=1.285
r290 60 65 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.415 $Y=0.45
+ $X2=6.5 $Y2=0.365
r291 60 61 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=6.415 $Y=0.45
+ $X2=6.415 $Y2=1.12
r292 58 63 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.33 $Y=2.275
+ $X2=6.415 $Y2=2.19
r293 58 59 52.1925 $w=1.68e-07 $l=8e-07 $layer=LI1_cond $X=6.33 $Y=2.275
+ $X2=5.53 $Y2=2.275
r294 56 59 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.445 $Y=2.36
+ $X2=5.53 $Y2=2.275
r295 56 57 35.5561 $w=1.68e-07 $l=5.45e-07 $layer=LI1_cond $X=5.445 $Y=2.36
+ $X2=5.445 $Y2=2.905
r296 54 57 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.36 $Y=2.99
+ $X2=5.445 $Y2=2.905
r297 54 55 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.36 $Y=2.99
+ $X2=4.69 $Y2=2.99
r298 53 55 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.605 $Y=2.905
+ $X2=4.69 $Y2=2.99
r299 52 53 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=4.605 $Y=2.565
+ $X2=4.605 $Y2=2.905
r300 51 69 2.28545 $w=1.7e-07 $l=1.1e-07 $layer=LI1_cond $X=3.845 $Y=2.48
+ $X2=3.735 $Y2=2.48
r301 50 52 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.52 $Y=2.48
+ $X2=4.605 $Y2=2.565
r302 50 51 44.0374 $w=1.68e-07 $l=6.75e-07 $layer=LI1_cond $X=4.52 $Y=2.48
+ $X2=3.845 $Y2=2.48
r303 48 69 4.14756 $w=2.2e-07 $l=8.5e-08 $layer=LI1_cond $X=3.735 $Y=2.565
+ $X2=3.735 $Y2=2.48
r304 48 49 17.8105 $w=2.18e-07 $l=3.4e-07 $layer=LI1_cond $X=3.735 $Y=2.565
+ $X2=3.735 $Y2=2.905
r305 46 82 27.1035 $w=3.3e-07 $l=1.55e-07 $layer=POLY_cond $X=3.735 $Y=1.6
+ $X2=3.58 $Y2=1.6
r306 45 46 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.735
+ $Y=1.6 $X2=3.735 $Y2=1.6
r307 43 69 4.14756 $w=2.2e-07 $l=8.5e-08 $layer=LI1_cond $X=3.735 $Y=2.395
+ $X2=3.735 $Y2=2.48
r308 43 45 41.6451 $w=2.18e-07 $l=7.95e-07 $layer=LI1_cond $X=3.735 $Y=2.395
+ $X2=3.735 $Y2=1.6
r309 41 68 65.8931 $w=1.68e-07 $l=1.01e-06 $layer=LI1_cond $X=3.025 $Y=0.425
+ $X2=3.025 $Y2=1.435
r310 38 68 8.30336 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=2.95 $Y=1.6
+ $X2=2.95 $Y2=1.435
r311 38 39 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.95
+ $Y=1.6 $X2=2.95 $Y2=1.6
r312 34 49 6.96323 $w=1.7e-07 $l=1.46458e-07 $layer=LI1_cond $X=3.625 $Y=2.99
+ $X2=3.735 $Y2=2.905
r313 34 35 88.0749 $w=1.68e-07 $l=1.35e-06 $layer=LI1_cond $X=3.625 $Y=2.99
+ $X2=2.275 $Y2=2.99
r314 32 41 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.94 $Y=0.34
+ $X2=3.025 $Y2=0.425
r315 32 33 47.2995 $w=1.68e-07 $l=7.25e-07 $layer=LI1_cond $X=2.94 $Y=0.34
+ $X2=2.215 $Y2=0.34
r316 28 35 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.19 $Y=2.905
+ $X2=2.275 $Y2=2.99
r317 28 30 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=2.19 $Y=2.905
+ $X2=2.19 $Y2=2.665
r318 24 33 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.13 $Y=0.425
+ $X2=2.215 $Y2=0.34
r319 24 26 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=2.13 $Y=0.425
+ $X2=2.13 $Y2=0.515
r320 21 78 55.8714 $w=3.2e-07 $l=3.24037e-07 $layer=POLY_cond $X=7.53 $Y=2.465
+ $X2=7.435 $Y2=2.185
r321 21 23 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=7.53 $Y=2.465
+ $X2=7.53 $Y2=2.75
r322 20 86 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=6.62 $Y=0.69
+ $X2=6.62 $Y2=1.12
r323 14 82 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.58 $Y=1.435
+ $X2=3.58 $Y2=1.6
r324 14 16 379.447 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=3.58 $Y=1.435
+ $X2=3.58 $Y2=0.695
r325 13 39 13.4654 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.115 $Y=1.6
+ $X2=2.95 $Y2=1.6
r326 12 82 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=3.505 $Y=1.6
+ $X2=3.58 $Y2=1.6
r327 12 13 68.1959 $w=3.3e-07 $l=3.9e-07 $layer=POLY_cond $X=3.505 $Y=1.6
+ $X2=3.115 $Y2=1.6
r328 9 11 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=3.005 $Y=2.24
+ $X2=3.005 $Y2=2.525
r329 8 9 55.1908 $w=2.62e-07 $l=3.26343e-07 $layer=POLY_cond $X=2.95 $Y=1.94
+ $X2=3.005 $Y2=2.24
r330 7 39 13.4654 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.95 $Y=1.765
+ $X2=2.95 $Y2=1.6
r331 7 8 30.6007 $w=3.3e-07 $l=1.75e-07 $layer=POLY_cond $X=2.95 $Y=1.765
+ $X2=2.95 $Y2=1.94
r332 2 30 600 $w=1.7e-07 $l=9.47035e-07 $layer=licon1_PDIFF $count=1 $X=2.04
+ $Y=1.79 $X2=2.19 $Y2=2.665
r333 1 26 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.99
+ $Y=0.37 $X2=2.13 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__DFSBP_2%A_757_401# 1 2 7 9 10 12 13 15 16 19 21 24
+ 25 30 34 38
c92 24 0 1.10712e-19 $X=4.305 $Y=1.99
c93 7 0 4.67629e-20 $X=3.875 $Y=2.24
r94 38 44 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=4.37 $Y=1.825
+ $X2=4.37 $Y2=1.345
r95 34 36 16.7582 $w=2.73e-07 $l=3.75e-07 $layer=LI1_cond $X=5.025 $Y=2.14
+ $X2=5.025 $Y2=2.515
r96 33 44 46.255 $w=3.35e-07 $l=1.65e-07 $layer=POLY_cond $X=4.462 $Y=1.18
+ $X2=4.462 $Y2=1.345
r97 32 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.465
+ $Y=1.18 $X2=4.465 $Y2=1.18
r98 30 32 18.866 $w=3.88e-07 $l=6.71714e-07 $layer=LI1_cond $X=4.617 $Y=0.58
+ $X2=4.465 $Y2=1.18
r99 25 39 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=4.305 $Y=1.99
+ $X2=4.305 $Y2=2.08
r100 25 38 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.305 $Y=1.99
+ $X2=4.305 $Y2=1.825
r101 24 27 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=4.305 $Y=1.99
+ $X2=4.305 $Y2=2.14
r102 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.305
+ $Y=1.99 $X2=4.305 $Y2=1.99
r103 22 27 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.47 $Y=2.14
+ $X2=4.305 $Y2=2.14
r104 21 34 3.50848 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.86 $Y=2.14
+ $X2=5.025 $Y2=2.14
r105 21 22 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=4.86 $Y=2.14
+ $X2=4.47 $Y2=2.14
r106 15 33 15.5026 $w=3.35e-07 $l=9e-08 $layer=POLY_cond $X=4.462 $Y=1.09
+ $X2=4.462 $Y2=1.18
r107 15 16 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=4.295 $Y=1.09
+ $X2=4.015 $Y2=1.09
r108 14 19 7.1379 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=3.965 $Y=2.08
+ $X2=3.875 $Y2=2.08
r109 13 39 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.14 $Y=2.08
+ $X2=4.305 $Y2=2.08
r110 13 14 89.734 $w=1.5e-07 $l=1.75e-07 $layer=POLY_cond $X=4.14 $Y=2.08
+ $X2=3.965 $Y2=2.08
r111 10 16 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.94 $Y=1.015
+ $X2=4.015 $Y2=1.09
r112 10 12 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=3.94 $Y=1.015
+ $X2=3.94 $Y2=0.695
r113 7 19 64.3434 $w=1.8e-07 $l=1.6e-07 $layer=POLY_cond $X=3.875 $Y=2.24
+ $X2=3.875 $Y2=2.08
r114 7 9 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=3.875 $Y=2.24
+ $X2=3.875 $Y2=2.525
r115 2 36 600 $w=1.7e-07 $l=2.64575e-07 $layer=licon1_PDIFF $count=1 $X=4.875
+ $Y=2.315 $X2=5.025 $Y2=2.515
r116 1 30 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=4.57
+ $Y=0.37 $X2=4.715 $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_HS__DFSBP_2%A_595_97# 1 2 8 9 11 14 16 19 20 22 23 25 26
+ 29 32 34 35 38 39 40 46 48 49 50 55 58 60 65
c171 58 0 8.86437e-20 $X=5.75 $Y=1.285
c172 55 0 2.29347e-19 $X=4.85 $Y=1.72
c173 48 0 1.55885e-19 $X=3.405 $Y=0.925
c174 34 0 4.67629e-20 $X=3.37 $Y=2.295
c175 9 0 1.18171e-19 $X=4.8 $Y=2.24
r176 59 65 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=5.75 $Y=1.285
+ $X2=5.75 $Y2=1.195
r177 58 60 8.51388 $w=2.88e-07 $l=1.65e-07 $layer=LI1_cond $X=5.75 $Y=1.265
+ $X2=5.585 $Y2=1.265
r178 58 59 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.75
+ $Y=1.285 $X2=5.75 $Y2=1.285
r179 55 64 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.85 $Y=1.72
+ $X2=4.85 $Y2=1.885
r180 55 63 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.85 $Y=1.72
+ $X2=4.85 $Y2=1.555
r181 54 55 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.85
+ $Y=1.72 $X2=4.85 $Y2=1.72
r182 44 46 3.66686 $w=4.38e-07 $l=1.4e-07 $layer=LI1_cond $X=3.23 $Y=2.515
+ $X2=3.37 $Y2=2.515
r183 42 50 3.33486 $w=1.7e-07 $l=1.33e-07 $layer=LI1_cond $X=5.015 $Y=1.325
+ $X2=4.882 $Y2=1.325
r184 42 60 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=5.015 $Y=1.325
+ $X2=5.585 $Y2=1.325
r185 39 54 5.21861 $w=2.63e-07 $l=1.2e-07 $layer=LI1_cond $X=4.882 $Y=1.6
+ $X2=4.882 $Y2=1.72
r186 39 50 11.9593 $w=2.63e-07 $l=2.75e-07 $layer=LI1_cond $X=4.882 $Y=1.6
+ $X2=4.882 $Y2=1.325
r187 39 40 36.861 $w=1.68e-07 $l=5.65e-07 $layer=LI1_cond $X=4.75 $Y=1.6
+ $X2=4.185 $Y2=1.6
r188 38 40 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.1 $Y=1.515
+ $X2=4.185 $Y2=1.6
r189 37 38 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=4.1 $Y=1.265
+ $X2=4.1 $Y2=1.515
r190 36 49 2.06925 $w=1.7e-07 $l=1.23e-07 $layer=LI1_cond $X=3.53 $Y=1.18
+ $X2=3.407 $Y2=1.18
r191 35 37 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.015 $Y=1.18
+ $X2=4.1 $Y2=1.265
r192 35 36 31.6417 $w=1.68e-07 $l=4.85e-07 $layer=LI1_cond $X=4.015 $Y=1.18
+ $X2=3.53 $Y2=1.18
r193 34 46 6.36164 $w=1.7e-07 $l=2.2e-07 $layer=LI1_cond $X=3.37 $Y=2.295
+ $X2=3.37 $Y2=2.515
r194 33 49 4.36305 $w=2.07e-07 $l=1.01833e-07 $layer=LI1_cond $X=3.37 $Y=1.265
+ $X2=3.407 $Y2=1.18
r195 33 34 67.1979 $w=1.68e-07 $l=1.03e-06 $layer=LI1_cond $X=3.37 $Y=1.265
+ $X2=3.37 $Y2=2.295
r196 32 49 4.36305 $w=2.07e-07 $l=8.5e-08 $layer=LI1_cond $X=3.407 $Y=1.095
+ $X2=3.407 $Y2=1.18
r197 32 48 7.99654 $w=2.43e-07 $l=1.7e-07 $layer=LI1_cond $X=3.407 $Y=1.095
+ $X2=3.407 $Y2=0.925
r198 27 48 5.76222 $w=2.48e-07 $l=1.25e-07 $layer=LI1_cond $X=3.405 $Y=0.8
+ $X2=3.405 $Y2=0.925
r199 27 29 4.84026 $w=2.48e-07 $l=1.05e-07 $layer=LI1_cond $X=3.405 $Y=0.8
+ $X2=3.405 $Y2=0.695
r200 23 26 18.8402 $w=1.65e-07 $l=8.21584e-08 $layer=POLY_cond $X=6.23 $Y=1.12
+ $X2=6.215 $Y2=1.195
r201 23 25 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=6.23 $Y=1.12
+ $X2=6.23 $Y2=0.69
r202 20 22 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=6.215 $Y=1.63
+ $X2=6.215 $Y2=2.205
r203 19 20 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=6.215 $Y=1.54
+ $X2=6.215 $Y2=1.63
r204 18 26 18.8402 $w=1.65e-07 $l=7.5e-08 $layer=POLY_cond $X=6.215 $Y=1.27
+ $X2=6.215 $Y2=1.195
r205 18 19 104.952 $w=1.8e-07 $l=2.7e-07 $layer=POLY_cond $X=6.215 $Y=1.27
+ $X2=6.215 $Y2=1.54
r206 17 65 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.915 $Y=1.195
+ $X2=5.75 $Y2=1.195
r207 16 26 6.66866 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=6.125 $Y=1.195
+ $X2=6.215 $Y2=1.195
r208 16 17 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=6.125 $Y=1.195
+ $X2=5.915 $Y2=1.195
r209 14 63 499.947 $w=1.5e-07 $l=9.75e-07 $layer=POLY_cond $X=4.93 $Y=0.58
+ $X2=4.93 $Y2=1.555
r210 9 11 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=4.8 $Y=2.24 $X2=4.8
+ $Y2=2.525
r211 8 9 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=4.8 $Y=2.15 $X2=4.8
+ $Y2=2.24
r212 8 64 103.008 $w=1.8e-07 $l=2.65e-07 $layer=POLY_cond $X=4.8 $Y=2.15 $X2=4.8
+ $Y2=1.885
r213 2 44 600 $w=1.7e-07 $l=2.64575e-07 $layer=licon1_PDIFF $count=1 $X=3.08
+ $Y=2.315 $X2=3.23 $Y2=2.515
r214 1 29 182 $w=1.7e-07 $l=4.83735e-07 $layer=licon1_NDIFF $count=1 $X=2.975
+ $Y=0.485 $X2=3.365 $Y2=0.695
.ends

.subckt PM_SKY130_FD_SC_HS__DFSBP_2%SET_B 3 5 6 8 9 11 12 13 15 16 18 19 20 21
+ 22 25 27 32 36
c124 22 0 1.18634e-19 $X=5.665 $Y=1.665
c125 6 0 1.74055e-19 $X=5.315 $Y=2.24
r126 36 45 10.3882 $w=3.53e-07 $l=3.2e-07 $layer=LI1_cond $X=8.462 $Y=1.345
+ $X2=8.462 $Y2=1.665
r127 35 37 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=8.475 $Y=1.345
+ $X2=8.475 $Y2=1.51
r128 35 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.475
+ $Y=1.345 $X2=8.475 $Y2=1.345
r129 32 35 31.475 $w=3.3e-07 $l=1.8e-07 $layer=POLY_cond $X=8.475 $Y=1.165
+ $X2=8.475 $Y2=1.345
r130 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.39
+ $Y=1.855 $X2=5.39 $Y2=1.855
r131 27 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=1.665
+ $X2=8.4 $Y2=1.665
r132 25 31 5.34059 $w=4.08e-07 $l=1.9e-07 $layer=LI1_cond $X=5.43 $Y=1.665
+ $X2=5.43 $Y2=1.855
r133 24 25 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=1.665
+ $X2=5.52 $Y2=1.665
r134 22 24 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.665 $Y=1.665
+ $X2=5.52 $Y2=1.665
r135 21 27 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=8.255 $Y=1.665
+ $X2=8.4 $Y2=1.665
r136 21 22 3.20544 $w=1.4e-07 $l=2.59e-06 $layer=MET1_cond $X=8.255 $Y=1.665
+ $X2=5.665 $Y2=1.665
r137 19 20 69.5192 $w=1.6e-07 $l=1.5e-07 $layer=POLY_cond $X=5.295 $Y=0.865
+ $X2=5.295 $Y2=1.015
r138 16 18 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=8.4 $Y=2.465 $X2=8.4
+ $Y2=2.75
r139 15 16 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=8.4 $Y=2.375 $X2=8.4
+ $Y2=2.465
r140 15 37 336.234 $w=1.8e-07 $l=8.65e-07 $layer=POLY_cond $X=8.4 $Y=2.375
+ $X2=8.4 $Y2=1.51
r141 12 32 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.31 $Y=1.165
+ $X2=8.475 $Y2=1.165
r142 12 13 135.883 $w=1.5e-07 $l=2.65e-07 $layer=POLY_cond $X=8.31 $Y=1.165
+ $X2=8.045 $Y2=1.165
r143 9 13 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=7.97 $Y=1.09
+ $X2=8.045 $Y2=1.165
r144 9 11 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=7.97 $Y=1.09
+ $X2=7.97 $Y2=0.8
r145 6 30 78.1767 $w=2.7e-07 $l=4.20833e-07 $layer=POLY_cond $X=5.315 $Y=2.24
+ $X2=5.39 $Y2=1.855
r146 6 8 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=5.315 $Y=2.24
+ $X2=5.315 $Y2=2.525
r147 5 30 38.9026 $w=2.7e-07 $l=2.05122e-07 $layer=POLY_cond $X=5.3 $Y=1.69
+ $X2=5.39 $Y2=1.855
r148 5 20 346.117 $w=1.5e-07 $l=6.75e-07 $layer=POLY_cond $X=5.3 $Y=1.69 $X2=5.3
+ $Y2=1.015
r149 3 19 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=5.29 $Y=0.58 $X2=5.29
+ $Y2=0.865
.ends

.subckt PM_SKY130_FD_SC_HS__DFSBP_2%A_225_74# 1 2 9 11 13 15 16 18 19 22 24 25
+ 26 28 29 34 35 36 39 43 46 47 49 50 51 54 58 62 65
c189 54 0 2.99812e-20 $X=1.945 $Y=1.805
c190 35 0 1.08117e-19 $X=7.115 $Y=1.735
r191 62 64 17.8607 $w=4.58e-07 $l=4.95e-07 $layer=LI1_cond $X=1.205 $Y=0.515
+ $X2=1.205 $Y2=1.01
r192 58 59 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.11
+ $Y=1.465 $X2=2.11 $Y2=1.465
r193 56 58 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=2.11 $Y=1.72
+ $X2=2.11 $Y2=1.465
r194 54 56 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.945 $Y=1.805
+ $X2=2.11 $Y2=1.72
r195 54 65 31.9679 $w=1.68e-07 $l=4.9e-07 $layer=LI1_cond $X=1.945 $Y=1.805
+ $X2=1.455 $Y2=1.805
r196 51 53 5.57014 $w=2.98e-07 $l=1.45e-07 $layer=LI1_cond $X=1.145 $Y=1.87
+ $X2=1.29 $Y2=1.87
r197 50 65 7.90841 $w=2.98e-07 $l=1.5e-07 $layer=LI1_cond $X=1.305 $Y=1.87
+ $X2=1.455 $Y2=1.87
r198 50 53 0.576222 $w=2.98e-07 $l=1.5e-08 $layer=LI1_cond $X=1.305 $Y=1.87
+ $X2=1.29 $Y2=1.87
r199 49 51 7.51767 $w=3e-07 $l=1.8775e-07 $layer=LI1_cond $X=1.06 $Y=1.72
+ $X2=1.145 $Y2=1.87
r200 49 64 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=1.06 $Y=1.72
+ $X2=1.06 $Y2=1.01
r201 46 59 52.4584 $w=3.3e-07 $l=3e-07 $layer=POLY_cond $X=2.41 $Y=1.465
+ $X2=2.11 $Y2=1.465
r202 43 46 176.904 $w=1.5e-07 $l=3.45e-07 $layer=POLY_cond $X=2.485 $Y=1.12
+ $X2=2.485 $Y2=1.465
r203 42 59 9.61737 $w=3.3e-07 $l=5.5e-08 $layer=POLY_cond $X=2.055 $Y=1.465
+ $X2=2.11 $Y2=1.465
r204 37 39 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=7.19 $Y=1.66
+ $X2=7.19 $Y2=0.8
r205 35 37 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=7.115 $Y=1.735
+ $X2=7.19 $Y2=1.66
r206 35 36 156.394 $w=1.5e-07 $l=3.05e-07 $layer=POLY_cond $X=7.115 $Y=1.735
+ $X2=6.81 $Y2=1.735
r207 32 34 294.84 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=6.72 $Y=3.035
+ $X2=6.72 $Y2=2.46
r208 31 36 26.9307 $w=1.5e-07 $l=1.89737e-07 $layer=POLY_cond $X=6.72 $Y=1.885
+ $X2=6.81 $Y2=1.735
r209 31 34 294.84 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=6.72 $Y=1.885
+ $X2=6.72 $Y2=2.46
r210 30 47 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=3.545 $Y=3.15
+ $X2=3.455 $Y2=3.15
r211 29 32 26.9307 $w=1.5e-07 $l=1.53542e-07 $layer=POLY_cond $X=6.63 $Y=3.15
+ $X2=6.72 $Y2=3.035
r212 29 30 1581.88 $w=1.5e-07 $l=3.085e-06 $layer=POLY_cond $X=6.63 $Y=3.15
+ $X2=3.545 $Y2=3.15
r213 26 28 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=3.455 $Y=2.81
+ $X2=3.455 $Y2=2.525
r214 25 47 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=3.455 $Y=3.075
+ $X2=3.455 $Y2=3.15
r215 24 26 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=3.455 $Y=2.9
+ $X2=3.455 $Y2=2.81
r216 24 25 68.0242 $w=1.8e-07 $l=1.75e-07 $layer=POLY_cond $X=3.455 $Y=2.9
+ $X2=3.455 $Y2=3.075
r217 20 22 179.468 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=2.9 $Y=1.045
+ $X2=2.9 $Y2=0.695
r218 18 47 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=3.365 $Y=3.15
+ $X2=3.455 $Y2=3.15
r219 18 19 412.777 $w=1.5e-07 $l=8.05e-07 $layer=POLY_cond $X=3.365 $Y=3.15
+ $X2=2.56 $Y2=3.15
r220 17 43 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.56 $Y=1.12
+ $X2=2.485 $Y2=1.12
r221 16 20 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.825 $Y=1.12
+ $X2=2.9 $Y2=1.045
r222 16 17 135.883 $w=1.5e-07 $l=2.65e-07 $layer=POLY_cond $X=2.825 $Y=1.12
+ $X2=2.56 $Y2=1.12
r223 15 19 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.485 $Y=3.075
+ $X2=2.56 $Y2=3.15
r224 14 46 84.6064 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.485 $Y=1.63
+ $X2=2.485 $Y2=1.465
r225 14 15 740.947 $w=1.5e-07 $l=1.445e-06 $layer=POLY_cond $X=2.485 $Y=1.63
+ $X2=2.485 $Y2=3.075
r226 11 42 61.9504 $w=2.07e-07 $l=2.58844e-07 $layer=POLY_cond $X=1.965 $Y=1.715
+ $X2=1.947 $Y2=1.465
r227 11 13 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.965 $Y=1.715
+ $X2=1.965 $Y2=2.35
r228 7 42 42.1581 $w=2.07e-07 $l=1.80291e-07 $layer=POLY_cond $X=1.915 $Y=1.3
+ $X2=1.947 $Y2=1.465
r229 7 9 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=1.915 $Y=1.3
+ $X2=1.915 $Y2=0.74
r230 2 53 600 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=1.145
+ $Y=1.79 $X2=1.29 $Y2=1.935
r231 1 62 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=1.125
+ $Y=0.37 $X2=1.27 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__DFSBP_2%A_1501_92# 1 2 9 12 13 15 18 19 21 22 23 25
+ 28 29 35
c108 23 0 1.4228e-19 $X=9.74 $Y=2.375
c109 19 0 2.30361e-19 $X=7.89 $Y=1.615
r110 37 38 5.93683 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=9.27 $Y=0.925
+ $X2=9.27 $Y2=1.095
r111 35 37 4.36531 $w=3.28e-07 $l=1.25e-07 $layer=LI1_cond $X=9.27 $Y=0.8
+ $X2=9.27 $Y2=0.925
r112 29 32 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=9.18 $Y=2.375 $X2=9.18
+ $Y2=2.455
r113 27 28 72.4171 $w=1.68e-07 $l=1.11e-06 $layer=LI1_cond $X=9.825 $Y=1.18
+ $X2=9.825 $Y2=2.29
r114 26 38 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.435 $Y=1.095
+ $X2=9.27 $Y2=1.095
r115 25 27 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.74 $Y=1.095
+ $X2=9.825 $Y2=1.18
r116 25 26 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=9.74 $Y=1.095
+ $X2=9.435 $Y2=1.095
r117 24 29 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.345 $Y=2.375
+ $X2=9.18 $Y2=2.375
r118 23 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.74 $Y=2.375
+ $X2=9.825 $Y2=2.29
r119 23 24 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=9.74 $Y=2.375
+ $X2=9.345 $Y2=2.375
r120 21 37 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.105 $Y=0.925
+ $X2=9.27 $Y2=0.925
r121 21 22 68.5027 $w=1.68e-07 $l=1.05e-06 $layer=LI1_cond $X=9.105 $Y=0.925
+ $X2=8.055 $Y2=0.925
r122 19 42 11.2093 $w=2.58e-07 $l=6e-08 $layer=POLY_cond $X=7.89 $Y=1.615
+ $X2=7.95 $Y2=1.615
r123 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.89
+ $Y=1.615 $X2=7.89 $Y2=1.615
r124 16 22 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=7.89 $Y=1.01
+ $X2=8.055 $Y2=0.925
r125 16 18 21.1281 $w=3.28e-07 $l=6.05e-07 $layer=LI1_cond $X=7.89 $Y=1.01
+ $X2=7.89 $Y2=1.615
r126 13 15 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=7.95 $Y=2.465
+ $X2=7.95 $Y2=2.75
r127 12 13 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=7.95 $Y=2.375
+ $X2=7.95 $Y2=2.465
r128 11 42 11.2427 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=7.95 $Y=1.78
+ $X2=7.95 $Y2=1.615
r129 11 12 231.282 $w=1.8e-07 $l=5.95e-07 $layer=POLY_cond $X=7.95 $Y=1.78
+ $X2=7.95 $Y2=2.375
r130 7 19 57.9147 $w=2.58e-07 $l=3.83732e-07 $layer=POLY_cond $X=7.58 $Y=1.45
+ $X2=7.89 $Y2=1.615
r131 7 9 333.298 $w=1.5e-07 $l=6.5e-07 $layer=POLY_cond $X=7.58 $Y=1.45 $X2=7.58
+ $Y2=0.8
r132 2 32 600 $w=1.7e-07 $l=6.83667e-07 $layer=licon1_PDIFF $count=1 $X=9.035
+ $Y=1.84 $X2=9.18 $Y2=2.455
r133 1 35 182 $w=1.7e-07 $l=3.07571e-07 $layer=licon1_NDIFF $count=1 $X=9.05
+ $Y=0.59 $X2=9.27 $Y2=0.8
.ends

.subckt PM_SKY130_FD_SC_HS__DFSBP_2%A_1339_74# 1 2 3 12 14 15 16 18 19 21 23 26
+ 28 30 33 35 36 39 41 43 48 49 56 58 61 63 65 69 75 76 77 80
c194 61 0 1.07812e-19 $X=8.46 $Y=2.215
c195 48 0 8.81429e-20 $X=11.475 $Y=1.557
c196 14 0 1.4228e-19 $X=9.395 $Y=1.515
r197 79 80 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=9.405
+ $Y=1.515 $X2=9.405 $Y2=1.515
r198 76 77 9.81721 $w=5.28e-07 $l=1.7e-07 $layer=LI1_cond $X=7.75 $Y=2.3
+ $X2=7.92 $Y2=2.3
r199 75 76 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=7.47 $Y=2.565
+ $X2=7.75 $Y2=2.565
r200 74 75 9.51712 $w=4.98e-07 $l=1.65e-07 $layer=LI1_cond $X=7.305 $Y=2.73
+ $X2=7.47 $Y2=2.73
r201 71 74 9.56863 $w=4.98e-07 $l=4e-07 $layer=LI1_cond $X=6.905 $Y=2.73
+ $X2=7.305 $Y2=2.73
r202 63 65 9.42908 $w=3.28e-07 $l=2.7e-07 $layer=LI1_cond $X=8.625 $Y=2.48
+ $X2=8.625 $Y2=2.75
r203 61 63 7.87997 $w=6.27e-07 $l=3.37565e-07 $layer=LI1_cond $X=8.46 $Y=2.215
+ $X2=8.625 $Y2=2.48
r204 61 79 13.6204 $w=6.27e-07 $l=9.37283e-07 $layer=LI1_cond $X=8.46 $Y=2.215
+ $X2=9.015 $Y2=1.515
r205 61 77 12.1865 $w=5.28e-07 $l=5.4e-07 $layer=LI1_cond $X=8.46 $Y=2.215
+ $X2=7.92 $Y2=2.215
r206 58 69 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.13 $Y=1.68
+ $X2=7.13 $Y2=1.765
r207 57 58 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=7.13 $Y=0.95
+ $X2=7.13 $Y2=1.68
r208 54 71 4.80115 $w=2.5e-07 $l=2.5e-07 $layer=LI1_cond $X=6.905 $Y=2.48
+ $X2=6.905 $Y2=2.73
r209 54 56 15.9037 $w=2.48e-07 $l=3.45e-07 $layer=LI1_cond $X=6.905 $Y=2.48
+ $X2=6.905 $Y2=2.135
r210 53 69 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=6.905 $Y=1.765
+ $X2=7.13 $Y2=1.765
r211 53 56 13.1378 $w=2.48e-07 $l=2.85e-07 $layer=LI1_cond $X=6.905 $Y=1.85
+ $X2=6.905 $Y2=2.135
r212 49 57 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=7.045 $Y=0.785
+ $X2=7.13 $Y2=0.95
r213 49 51 4.88915 $w=3.28e-07 $l=1.4e-07 $layer=LI1_cond $X=7.045 $Y=0.785
+ $X2=6.905 $Y2=0.785
r214 46 47 0.67507 $w=3.57e-07 $l=5e-09 $layer=POLY_cond $X=10.47 $Y=1.557
+ $X2=10.475 $Y2=1.557
r215 45 46 57.381 $w=3.57e-07 $l=4.25e-07 $layer=POLY_cond $X=10.045 $Y=1.557
+ $X2=10.47 $Y2=1.557
r216 44 45 3.37535 $w=3.57e-07 $l=2.5e-08 $layer=POLY_cond $X=10.02 $Y=1.557
+ $X2=10.045 $Y2=1.557
r217 41 48 33.0931 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=11.475 $Y=1.765
+ $X2=11.475 $Y2=1.557
r218 41 43 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=11.475 $Y=1.765
+ $X2=11.475 $Y2=2.34
r219 37 48 33.0931 $w=1.5e-07 $l=2.11941e-07 $layer=POLY_cond $X=11.465 $Y=1.35
+ $X2=11.475 $Y2=1.557
r220 37 39 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=11.465 $Y=1.35
+ $X2=11.465 $Y2=0.69
r221 36 47 13.8507 $w=3.57e-07 $l=1.13666e-07 $layer=POLY_cond $X=10.56 $Y=1.49
+ $X2=10.475 $Y2=1.557
r222 35 48 3.06035 $w=2.8e-07 $l=1.1887e-07 $layer=POLY_cond $X=11.385 $Y=1.49
+ $X2=11.475 $Y2=1.557
r223 35 36 176.747 $w=2.8e-07 $l=8.25e-07 $layer=POLY_cond $X=11.385 $Y=1.49
+ $X2=10.56 $Y2=1.49
r224 31 47 23.1043 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=10.475 $Y=1.35
+ $X2=10.475 $Y2=1.557
r225 31 33 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=10.475 $Y=1.35
+ $X2=10.475 $Y2=0.74
r226 28 46 23.1043 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=10.47 $Y=1.765
+ $X2=10.47 $Y2=1.557
r227 28 30 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=10.47 $Y=1.765
+ $X2=10.47 $Y2=2.4
r228 24 45 23.1043 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=10.045 $Y=1.35
+ $X2=10.045 $Y2=1.557
r229 24 26 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=10.045 $Y=1.35
+ $X2=10.045 $Y2=0.74
r230 21 44 23.1043 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=10.02 $Y=1.765
+ $X2=10.02 $Y2=1.557
r231 21 23 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=10.02 $Y=1.765
+ $X2=10.02 $Y2=2.4
r232 20 80 10.9339 $w=3.05e-07 $l=1.1887e-07 $layer=POLY_cond $X=9.575 $Y=1.49
+ $X2=9.485 $Y2=1.557
r233 19 44 14.5258 $w=3.57e-07 $l=1.1887e-07 $layer=POLY_cond $X=9.93 $Y=1.49
+ $X2=10.02 $Y2=1.557
r234 19 20 76.0548 $w=2.8e-07 $l=3.55e-07 $layer=POLY_cond $X=9.93 $Y=1.49
+ $X2=9.575 $Y2=1.49
r235 16 80 15.748 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=9.485 $Y=1.765
+ $X2=9.485 $Y2=1.557
r236 16 18 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=9.485 $Y=1.765
+ $X2=9.485 $Y2=2.05
r237 14 80 10.9339 $w=3.05e-07 $l=1.08995e-07 $layer=POLY_cond $X=9.395 $Y=1.515
+ $X2=9.485 $Y2=1.557
r238 14 15 60.3271 $w=3.3e-07 $l=3.45e-07 $layer=POLY_cond $X=9.395 $Y=1.515
+ $X2=9.05 $Y2=1.515
r239 10 15 32.1775 $w=3.3e-07 $l=1.98997e-07 $layer=POLY_cond $X=8.975 $Y=1.35
+ $X2=9.05 $Y2=1.515
r240 10 12 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=8.975 $Y=1.35
+ $X2=8.975 $Y2=0.8
r241 3 65 600 $w=1.7e-07 $l=2.74955e-07 $layer=licon1_PDIFF $count=1 $X=8.475
+ $Y=2.54 $X2=8.625 $Y2=2.75
r242 2 74 300 $w=1.7e-07 $l=1.08031e-06 $layer=licon1_PDIFF $count=2 $X=6.795
+ $Y=1.96 $X2=7.305 $Y2=2.815
r243 2 56 300 $w=1.7e-07 $l=2.38485e-07 $layer=licon1_PDIFF $count=2 $X=6.795
+ $Y=1.96 $X2=6.945 $Y2=2.135
r244 1 51 182 $w=1.7e-07 $l=5.09289e-07 $layer=licon1_NDIFF $count=1 $X=6.695
+ $Y=0.37 $X2=6.905 $Y2=0.785
.ends

.subckt PM_SKY130_FD_SC_HS__DFSBP_2%A_2221_74# 1 2 7 9 12 14 16 19 23 27 33 36
+ 40
c71 7 0 1.00299e-19 $X=12.005 $Y=1.765
r72 40 41 1.22646 $w=3.93e-07 $l=1e-08 $layer=POLY_cond $X=12.455 $Y=1.532
+ $X2=12.465 $Y2=1.532
r73 39 40 51.5115 $w=3.93e-07 $l=4.2e-07 $layer=POLY_cond $X=12.035 $Y=1.532
+ $X2=12.455 $Y2=1.532
r74 38 39 3.67939 $w=3.93e-07 $l=3e-08 $layer=POLY_cond $X=12.005 $Y=1.532
+ $X2=12.035 $Y2=1.532
r75 34 38 7.97201 $w=3.93e-07 $l=6.5e-08 $layer=POLY_cond $X=11.94 $Y=1.532
+ $X2=12.005 $Y2=1.532
r76 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=11.94
+ $Y=1.465 $X2=11.94 $Y2=1.465
r77 31 36 1.34256 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=11.415 $Y=1.465
+ $X2=11.25 $Y2=1.465
r78 31 33 18.3343 $w=3.28e-07 $l=5.25e-07 $layer=LI1_cond $X=11.415 $Y=1.465
+ $X2=11.94 $Y2=1.465
r79 27 29 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=11.25 $Y=1.985
+ $X2=11.25 $Y2=2.695
r80 25 36 5.16603 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=11.25 $Y=1.63
+ $X2=11.25 $Y2=1.465
r81 25 27 12.3975 $w=3.28e-07 $l=3.55e-07 $layer=LI1_cond $X=11.25 $Y=1.63
+ $X2=11.25 $Y2=1.985
r82 21 36 5.16603 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=11.25 $Y=1.3
+ $X2=11.25 $Y2=1.465
r83 21 23 27.4142 $w=3.28e-07 $l=7.85e-07 $layer=LI1_cond $X=11.25 $Y=1.3
+ $X2=11.25 $Y2=0.515
r84 17 41 25.4309 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=12.465 $Y=1.3
+ $X2=12.465 $Y2=1.532
r85 17 19 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=12.465 $Y=1.3
+ $X2=12.465 $Y2=0.74
r86 14 40 25.4309 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=12.455 $Y=1.765
+ $X2=12.455 $Y2=1.532
r87 14 16 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=12.455 $Y=1.765
+ $X2=12.455 $Y2=2.4
r88 10 39 25.4309 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=12.035 $Y=1.3
+ $X2=12.035 $Y2=1.532
r89 10 12 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=12.035 $Y=1.3
+ $X2=12.035 $Y2=0.74
r90 7 38 25.4309 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=12.005 $Y=1.765
+ $X2=12.005 $Y2=1.532
r91 7 9 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=12.005 $Y=1.765
+ $X2=12.005 $Y2=2.4
r92 2 29 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=11.105
+ $Y=1.84 $X2=11.25 $Y2=2.695
r93 2 27 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=11.105
+ $Y=1.84 $X2=11.25 $Y2=1.985
r94 1 23 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=11.105
+ $Y=0.37 $X2=11.25 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__DFSBP_2%A_27_74# 1 2 3 4 15 18 21 23 25 28 29 30 31
+ 38
r70 35 38 5.41299 $w=3.28e-07 $l=1.55e-07 $layer=LI1_cond $X=2.53 $Y=0.76
+ $X2=2.685 $Y2=0.76
r71 31 33 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=1.71 $Y=2.145
+ $X2=1.71 $Y2=2.275
r72 27 35 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.53 $Y=0.925
+ $X2=2.53 $Y2=0.76
r73 27 28 74.0481 $w=1.68e-07 $l=1.135e-06 $layer=LI1_cond $X=2.53 $Y=0.925
+ $X2=2.53 $Y2=2.06
r74 26 31 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.795 $Y=2.145
+ $X2=1.71 $Y2=2.145
r75 25 42 13.5964 $w=3.32e-07 $l=4.63249e-07 $layer=LI1_cond $X=2.445 $Y=2.145
+ $X2=2.655 $Y2=2.515
r76 25 28 6.01991 $w=3.32e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.445 $Y=2.145
+ $X2=2.53 $Y2=2.06
r77 25 26 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=2.445 $Y=2.145
+ $X2=1.795 $Y2=2.145
r78 24 30 2.11342 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.365 $Y=2.275
+ $X2=0.24 $Y2=2.275
r79 23 33 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.625 $Y=2.275
+ $X2=1.71 $Y2=2.275
r80 23 24 82.2032 $w=1.68e-07 $l=1.26e-06 $layer=LI1_cond $X=1.625 $Y=2.275
+ $X2=0.365 $Y2=2.275
r81 19 30 4.3182 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=0.24 $Y=2.36 $X2=0.24
+ $Y2=2.275
r82 19 21 17.9781 $w=2.48e-07 $l=3.9e-07 $layer=LI1_cond $X=0.24 $Y=2.36
+ $X2=0.24 $Y2=2.75
r83 18 30 4.3182 $w=2.1e-07 $l=1.03078e-07 $layer=LI1_cond $X=0.2 $Y=2.19
+ $X2=0.24 $Y2=2.275
r84 18 29 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=0.2 $Y=2.19 $X2=0.2
+ $Y2=0.81
r85 13 29 6.94937 $w=2.48e-07 $l=1.25e-07 $layer=LI1_cond $X=0.24 $Y=0.685
+ $X2=0.24 $Y2=0.81
r86 13 15 4.84026 $w=2.48e-07 $l=1.05e-07 $layer=LI1_cond $X=0.24 $Y=0.685
+ $X2=0.24 $Y2=0.58
r87 4 42 600 $w=1.7e-07 $l=2.62678e-07 $layer=licon1_PDIFF $count=1 $X=2.635
+ $Y=2.315 $X2=2.78 $Y2=2.515
r88 3 21 600 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.54 $X2=0.28 $Y2=2.75
r89 2 38 182 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_NDIFF $count=1 $X=2.54
+ $Y=0.485 $X2=2.685 $Y2=0.76
r90 1 15 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_HS__DFSBP_2%VPWR 1 2 3 4 5 6 7 8 9 30 34 38 42 46 50 54
+ 60 64 66 71 72 74 75 76 78 83 88 93 105 116 120 126 129 132 135 138 141 145
c146 34 0 2.99812e-20 $X=1.74 $Y=2.73
r147 144 145 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.72 $Y=3.33
+ $X2=12.72 $Y2=3.33
r148 141 142 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.76 $Y=3.33
+ $X2=11.76 $Y2=3.33
r149 138 139 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.84 $Y=3.33
+ $X2=9.84 $Y2=3.33
r150 135 136 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r151 132 133 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r152 129 130 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r153 126 127 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r154 124 145 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.24 $Y=3.33
+ $X2=12.72 $Y2=3.33
r155 124 142 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.24 $Y=3.33
+ $X2=11.76 $Y2=3.33
r156 123 124 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.24 $Y=3.33
+ $X2=12.24 $Y2=3.33
r157 121 141 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=11.865 $Y=3.33
+ $X2=11.74 $Y2=3.33
r158 121 123 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=11.865 $Y=3.33
+ $X2=12.24 $Y2=3.33
r159 120 144 4.01252 $w=1.7e-07 $l=1.82e-07 $layer=LI1_cond $X=12.595 $Y=3.33
+ $X2=12.777 $Y2=3.33
r160 120 123 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=12.595 $Y=3.33
+ $X2=12.24 $Y2=3.33
r161 119 142 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.28 $Y=3.33
+ $X2=11.76 $Y2=3.33
r162 118 119 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=11.28 $Y=3.33
+ $X2=11.28 $Y2=3.33
r163 116 141 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=11.615 $Y=3.33
+ $X2=11.74 $Y2=3.33
r164 116 118 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=11.615 $Y=3.33
+ $X2=11.28 $Y2=3.33
r165 115 119 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=10.32 $Y=3.33
+ $X2=11.28 $Y2=3.33
r166 115 139 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.32 $Y=3.33
+ $X2=9.84 $Y2=3.33
r167 114 115 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.32 $Y=3.33
+ $X2=10.32 $Y2=3.33
r168 112 138 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.96 $Y=3.33
+ $X2=9.795 $Y2=3.33
r169 112 114 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=9.96 $Y=3.33
+ $X2=10.32 $Y2=3.33
r170 111 139 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.36 $Y=3.33
+ $X2=9.84 $Y2=3.33
r171 110 111 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=9.36 $Y=3.33
+ $X2=9.36 $Y2=3.33
r172 108 111 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=8.4 $Y=3.33
+ $X2=9.36 $Y2=3.33
r173 107 110 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=8.4 $Y=3.33
+ $X2=9.36 $Y2=3.33
r174 107 108 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=8.4 $Y=3.33
+ $X2=8.4 $Y2=3.33
r175 105 138 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.63 $Y=3.33
+ $X2=9.795 $Y2=3.33
r176 105 110 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=9.63 $Y=3.33
+ $X2=9.36 $Y2=3.33
r177 104 108 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=3.33
+ $X2=8.4 $Y2=3.33
r178 103 104 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r179 101 135 9.31531 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=6.07 $Y=3.33
+ $X2=5.885 $Y2=3.33
r180 101 103 120.695 $w=1.68e-07 $l=1.85e-06 $layer=LI1_cond $X=6.07 $Y=3.33
+ $X2=7.92 $Y2=3.33
r181 100 136 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=6 $Y2=3.33
r182 99 100 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r183 97 100 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=5.52 $Y2=3.33
r184 97 133 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=4.08 $Y2=3.33
r185 96 99 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=4.56 $Y=3.33
+ $X2=5.52 $Y2=3.33
r186 96 97 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r187 94 132 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.35 $Y=3.33
+ $X2=4.185 $Y2=3.33
r188 94 96 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=4.35 $Y=3.33
+ $X2=4.56 $Y2=3.33
r189 93 135 9.31531 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=5.7 $Y=3.33
+ $X2=5.885 $Y2=3.33
r190 93 99 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=5.7 $Y=3.33
+ $X2=5.52 $Y2=3.33
r191 92 133 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=4.08 $Y2=3.33
r192 92 130 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.68 $Y2=3.33
r193 91 92 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r194 89 129 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.905 $Y=3.33
+ $X2=1.74 $Y2=3.33
r195 89 91 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=1.905 $Y=3.33
+ $X2=2.16 $Y2=3.33
r196 88 132 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.02 $Y=3.33
+ $X2=4.185 $Y2=3.33
r197 88 91 121.348 $w=1.68e-07 $l=1.86e-06 $layer=LI1_cond $X=4.02 $Y=3.33
+ $X2=2.16 $Y2=3.33
r198 87 130 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=1.68 $Y2=3.33
r199 87 127 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r200 86 87 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r201 84 126 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.895 $Y=3.33
+ $X2=0.73 $Y2=3.33
r202 84 86 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.895 $Y=3.33
+ $X2=1.2 $Y2=3.33
r203 83 129 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.575 $Y=3.33
+ $X2=1.74 $Y2=3.33
r204 83 86 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=1.575 $Y=3.33
+ $X2=1.2 $Y2=3.33
r205 81 127 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r206 80 81 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r207 78 126 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.565 $Y=3.33
+ $X2=0.73 $Y2=3.33
r208 78 80 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.565 $Y=3.33
+ $X2=0.24 $Y2=3.33
r209 76 104 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=7.92 $Y2=3.33
r210 76 136 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=6 $Y2=3.33
r211 74 114 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=10.605 $Y=3.33
+ $X2=10.32 $Y2=3.33
r212 74 75 7.13466 $w=1.7e-07 $l=1.27e-07 $layer=LI1_cond $X=10.605 $Y=3.33
+ $X2=10.732 $Y2=3.33
r213 73 118 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=10.86 $Y=3.33
+ $X2=11.28 $Y2=3.33
r214 73 75 7.13466 $w=1.7e-07 $l=1.28e-07 $layer=LI1_cond $X=10.86 $Y=3.33
+ $X2=10.732 $Y2=3.33
r215 71 103 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=8.09 $Y=3.33
+ $X2=7.92 $Y2=3.33
r216 71 72 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.09 $Y=3.33
+ $X2=8.175 $Y2=3.33
r217 70 107 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=8.26 $Y=3.33
+ $X2=8.4 $Y2=3.33
r218 70 72 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.26 $Y=3.33
+ $X2=8.175 $Y2=3.33
r219 66 69 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=12.72 $Y=1.985
+ $X2=12.72 $Y2=2.815
r220 64 144 3.13065 $w=2.5e-07 $l=1.09864e-07 $layer=LI1_cond $X=12.72 $Y=3.245
+ $X2=12.777 $Y2=3.33
r221 64 69 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=12.72 $Y=3.245
+ $X2=12.72 $Y2=2.815
r222 60 63 32.7294 $w=2.48e-07 $l=7.1e-07 $layer=LI1_cond $X=11.74 $Y=1.985
+ $X2=11.74 $Y2=2.695
r223 58 141 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=11.74 $Y=3.245
+ $X2=11.74 $Y2=3.33
r224 58 63 25.3537 $w=2.48e-07 $l=5.5e-07 $layer=LI1_cond $X=11.74 $Y=3.245
+ $X2=11.74 $Y2=2.695
r225 54 57 37.059 $w=2.53e-07 $l=8.2e-07 $layer=LI1_cond $X=10.732 $Y=1.985
+ $X2=10.732 $Y2=2.805
r226 52 75 0.067832 $w=2.55e-07 $l=8.5e-08 $layer=LI1_cond $X=10.732 $Y=3.245
+ $X2=10.732 $Y2=3.33
r227 52 57 19.8853 $w=2.53e-07 $l=4.4e-07 $layer=LI1_cond $X=10.732 $Y=3.245
+ $X2=10.732 $Y2=2.805
r228 48 138 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.795 $Y=3.245
+ $X2=9.795 $Y2=3.33
r229 48 50 15.3659 $w=3.28e-07 $l=4.4e-07 $layer=LI1_cond $X=9.795 $Y=3.245
+ $X2=9.795 $Y2=2.805
r230 44 72 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.175 $Y=3.245
+ $X2=8.175 $Y2=3.33
r231 44 46 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=8.175 $Y=3.245
+ $X2=8.175 $Y2=2.815
r232 40 135 1.24149 $w=3.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.885 $Y=3.245
+ $X2=5.885 $Y2=3.33
r233 40 42 17.1309 $w=3.68e-07 $l=5.5e-07 $layer=LI1_cond $X=5.885 $Y=3.245
+ $X2=5.885 $Y2=2.695
r234 36 132 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.185 $Y=3.245
+ $X2=4.185 $Y2=3.33
r235 36 38 14.8421 $w=3.28e-07 $l=4.25e-07 $layer=LI1_cond $X=4.185 $Y=3.245
+ $X2=4.185 $Y2=2.82
r236 32 129 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.74 $Y=3.245
+ $X2=1.74 $Y2=3.33
r237 32 34 17.9851 $w=3.28e-07 $l=5.15e-07 $layer=LI1_cond $X=1.74 $Y=3.245
+ $X2=1.74 $Y2=2.73
r238 28 126 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.73 $Y=3.245
+ $X2=0.73 $Y2=3.33
r239 28 30 17.112 $w=3.28e-07 $l=4.9e-07 $layer=LI1_cond $X=0.73 $Y=3.245
+ $X2=0.73 $Y2=2.755
r240 9 69 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=12.53
+ $Y=1.84 $X2=12.68 $Y2=2.815
r241 9 66 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=12.53
+ $Y=1.84 $X2=12.68 $Y2=1.985
r242 8 63 400 $w=1.7e-07 $l=9.63159e-07 $layer=licon1_PDIFF $count=1 $X=11.55
+ $Y=1.84 $X2=11.78 $Y2=2.695
r243 8 60 400 $w=1.7e-07 $l=2.93684e-07 $layer=licon1_PDIFF $count=1 $X=11.55
+ $Y=1.84 $X2=11.78 $Y2=1.985
r244 7 57 400 $w=1.7e-07 $l=1.03729e-06 $layer=licon1_PDIFF $count=1 $X=10.545
+ $Y=1.84 $X2=10.695 $Y2=2.805
r245 7 54 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=10.545
+ $Y=1.84 $X2=10.695 $Y2=1.985
r246 6 50 600 $w=1.7e-07 $l=1.0761e-06 $layer=licon1_PDIFF $count=1 $X=9.56
+ $Y=1.84 $X2=9.795 $Y2=2.805
r247 5 46 600 $w=1.7e-07 $l=3.4187e-07 $layer=licon1_PDIFF $count=1 $X=8.025
+ $Y=2.54 $X2=8.175 $Y2=2.815
r248 4 42 600 $w=1.7e-07 $l=6.58122e-07 $layer=licon1_PDIFF $count=1 $X=5.39
+ $Y=2.315 $X2=5.885 $Y2=2.695
r249 3 38 600 $w=1.7e-07 $l=6.1131e-07 $layer=licon1_PDIFF $count=1 $X=3.95
+ $Y=2.315 $X2=4.185 $Y2=2.82
r250 2 34 600 $w=1.7e-07 $l=1.01223e-06 $layer=licon1_PDIFF $count=1 $X=1.59
+ $Y=1.79 $X2=1.74 $Y2=2.73
r251 1 30 600 $w=1.7e-07 $l=2.80134e-07 $layer=licon1_PDIFF $count=1 $X=0.58
+ $Y=2.54 $X2=0.73 $Y2=2.755
.ends

.subckt PM_SKY130_FD_SC_HS__DFSBP_2%Q_N 1 2 7 8 9 10 11 32
r27 29 32 0.491205 $w=3.03e-07 $l=1.3e-08 $layer=LI1_cond $X=10.282 $Y=1.972
+ $X2=10.282 $Y2=1.985
r28 11 29 0.415635 $w=3.03e-07 $l=1.1e-08 $layer=LI1_cond $X=10.282 $Y=1.961
+ $X2=10.282 $Y2=1.972
r29 11 38 5.61139 $w=3.03e-07 $l=1.41e-07 $layer=LI1_cond $X=10.282 $Y=1.961
+ $X2=10.282 $Y2=1.82
r30 11 35 28.6788 $w=3.03e-07 $l=7.59e-07 $layer=LI1_cond $X=10.282 $Y=2.046
+ $X2=10.282 $Y2=2.805
r31 11 32 2.30489 $w=3.03e-07 $l=6.1e-08 $layer=LI1_cond $X=10.282 $Y=2.046
+ $X2=10.282 $Y2=1.985
r32 10 38 6.87033 $w=2.58e-07 $l=1.55e-07 $layer=LI1_cond $X=10.305 $Y=1.665
+ $X2=10.305 $Y2=1.82
r33 9 10 16.4002 $w=2.58e-07 $l=3.7e-07 $layer=LI1_cond $X=10.305 $Y=1.295
+ $X2=10.305 $Y2=1.665
r34 8 9 16.4002 $w=2.58e-07 $l=3.7e-07 $layer=LI1_cond $X=10.305 $Y=0.925
+ $X2=10.305 $Y2=1.295
r35 7 8 18.1731 $w=2.58e-07 $l=4.1e-07 $layer=LI1_cond $X=10.305 $Y=0.515
+ $X2=10.305 $Y2=0.925
r36 2 35 400 $w=1.7e-07 $l=1.03729e-06 $layer=licon1_PDIFF $count=1 $X=10.095
+ $Y=1.84 $X2=10.245 $Y2=2.805
r37 2 32 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=10.095
+ $Y=1.84 $X2=10.245 $Y2=1.985
r38 1 7 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=10.12
+ $Y=0.37 $X2=10.26 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__DFSBP_2%Q 1 2 9 14 15 16 17 28
c32 15 0 1.88442e-19 $X=12.245 $Y=1.82
r33 21 28 1.18634 $w=3.38e-07 $l=3.5e-08 $layer=LI1_cond $X=12.255 $Y=0.96
+ $X2=12.255 $Y2=0.925
r34 17 30 7.79401 $w=3.38e-07 $l=1.45e-07 $layer=LI1_cond $X=12.255 $Y=0.985
+ $X2=12.255 $Y2=1.13
r35 17 21 0.847385 $w=3.38e-07 $l=2.5e-08 $layer=LI1_cond $X=12.255 $Y=0.985
+ $X2=12.255 $Y2=0.96
r36 17 28 0.847385 $w=3.38e-07 $l=2.5e-08 $layer=LI1_cond $X=12.255 $Y=0.9
+ $X2=12.255 $Y2=0.925
r37 16 17 13.0497 $w=3.38e-07 $l=3.85e-07 $layer=LI1_cond $X=12.255 $Y=0.515
+ $X2=12.255 $Y2=0.9
r38 15 30 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=12.34 $Y=1.82
+ $X2=12.34 $Y2=1.13
r39 14 15 8.51103 $w=3.58e-07 $l=1.65e-07 $layer=LI1_cond $X=12.245 $Y=1.985
+ $X2=12.245 $Y2=1.82
r40 7 14 0.480185 $w=3.58e-07 $l=1.5e-08 $layer=LI1_cond $X=12.245 $Y=2
+ $X2=12.245 $Y2=1.985
r41 7 9 26.09 $w=3.58e-07 $l=8.15e-07 $layer=LI1_cond $X=12.245 $Y=2 $X2=12.245
+ $Y2=2.815
r42 2 14 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=12.08
+ $Y=1.84 $X2=12.23 $Y2=1.985
r43 2 9 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=12.08
+ $Y=1.84 $X2=12.23 $Y2=2.815
r44 1 16 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=12.11
+ $Y=0.37 $X2=12.25 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__DFSBP_2%VGND 1 2 3 4 5 6 7 8 9 30 32 36 40 44 48 52
+ 54 56 59 60 61 63 68 89 98 102 108 111 114 119 125 129 132 134 137 141
c142 36 0 1.39813e-19 $X=1.7 $Y=0.505
r143 140 141 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.72 $Y=0
+ $X2=12.72 $Y2=0
r144 137 138 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.76 $Y=0
+ $X2=11.76 $Y2=0
r145 134 135 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.84 $Y=0
+ $X2=9.84 $Y2=0
r146 131 132 11.1544 $w=7.53e-07 $l=1.65e-07 $layer=LI1_cond $X=8.68 $Y=0.292
+ $X2=8.845 $Y2=0.292
r147 127 131 4.43579 $w=7.53e-07 $l=2.8e-07 $layer=LI1_cond $X=8.4 $Y=0.292
+ $X2=8.68 $Y2=0.292
r148 127 129 13.2931 $w=7.53e-07 $l=3e-07 $layer=LI1_cond $X=8.4 $Y=0.292
+ $X2=8.1 $Y2=0.292
r149 127 128 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r150 123 125 11.1389 $w=7.63e-07 $l=1.6e-07 $layer=LI1_cond $X=6 $Y=0.297
+ $X2=6.16 $Y2=0.297
r151 123 124 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=0 $X2=6
+ $Y2=0
r152 121 123 0.0781751 $w=7.63e-07 $l=5e-09 $layer=LI1_cond $X=5.995 $Y=0.297
+ $X2=6 $Y2=0.297
r153 118 124 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=6
+ $Y2=0
r154 117 121 7.42663 $w=7.63e-07 $l=4.75e-07 $layer=LI1_cond $X=5.52 $Y=0.297
+ $X2=5.995 $Y2=0.297
r155 117 119 11.4516 $w=7.63e-07 $l=1.8e-07 $layer=LI1_cond $X=5.52 $Y=0.297
+ $X2=5.34 $Y2=0.297
r156 117 118 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=0
+ $X2=5.52 $Y2=0
r157 114 115 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=0
+ $X2=4.08 $Y2=0
r158 111 112 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=0
+ $X2=1.68 $Y2=0
r159 109 112 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=0
+ $X2=1.68 $Y2=0
r160 108 109 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.72 $Y=0
+ $X2=0.72 $Y2=0
r161 106 141 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.24 $Y=0
+ $X2=12.72 $Y2=0
r162 106 138 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.24 $Y=0
+ $X2=11.76 $Y2=0
r163 105 106 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.24 $Y=0
+ $X2=12.24 $Y2=0
r164 103 137 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.915 $Y=0
+ $X2=11.75 $Y2=0
r165 103 105 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=11.915 $Y=0
+ $X2=12.24 $Y2=0
r166 102 140 4.01252 $w=1.7e-07 $l=1.82e-07 $layer=LI1_cond $X=12.595 $Y=0
+ $X2=12.777 $Y2=0
r167 102 105 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=12.595 $Y=0
+ $X2=12.24 $Y2=0
r168 101 138 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.28 $Y=0
+ $X2=11.76 $Y2=0
r169 100 101 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=11.28 $Y=0
+ $X2=11.28 $Y2=0
r170 98 137 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.585 $Y=0
+ $X2=11.75 $Y2=0
r171 98 100 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=11.585 $Y=0
+ $X2=11.28 $Y2=0
r172 97 101 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=10.32 $Y=0
+ $X2=11.28 $Y2=0
r173 97 135 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.32 $Y=0
+ $X2=9.84 $Y2=0
r174 96 97 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.32 $Y=0
+ $X2=10.32 $Y2=0
r175 94 134 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.995 $Y=0
+ $X2=9.83 $Y2=0
r176 94 96 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=9.995 $Y=0
+ $X2=10.32 $Y2=0
r177 93 135 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.36 $Y=0
+ $X2=9.84 $Y2=0
r178 93 128 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=9.36 $Y=0 $X2=8.4
+ $Y2=0
r179 92 132 33.5989 $w=1.68e-07 $l=5.15e-07 $layer=LI1_cond $X=9.36 $Y=0
+ $X2=8.845 $Y2=0
r180 92 93 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.36 $Y=0 $X2=9.36
+ $Y2=0
r181 89 134 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.665 $Y=0
+ $X2=9.83 $Y2=0
r182 89 92 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=9.665 $Y=0
+ $X2=9.36 $Y2=0
r183 88 128 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=0 $X2=8.4
+ $Y2=0
r184 87 129 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=7.92 $Y=0 $X2=8.1
+ $Y2=0
r185 87 88 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.92 $Y=0 $X2=7.92
+ $Y2=0
r186 84 87 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=6.48 $Y=0 $X2=7.92
+ $Y2=0
r187 84 125 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=6.48 $Y=0 $X2=6.16
+ $Y2=0
r188 80 118 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=0
+ $X2=5.52 $Y2=0
r189 80 115 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.04 $Y=0
+ $X2=4.08 $Y2=0
r190 79 119 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=5.04 $Y=0 $X2=5.34
+ $Y2=0
r191 79 80 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r192 77 114 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.24 $Y=0
+ $X2=4.115 $Y2=0
r193 77 79 52.1925 $w=1.68e-07 $l=8e-07 $layer=LI1_cond $X=4.24 $Y=0 $X2=5.04
+ $Y2=0
r194 75 115 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.08
+ $Y2=0
r195 74 75 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r196 72 75 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=2.16 $Y=0 $X2=3.6
+ $Y2=0
r197 72 112 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0
+ $X2=1.68 $Y2=0
r198 71 74 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=2.16 $Y=0 $X2=3.6
+ $Y2=0
r199 71 72 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r200 69 111 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.865 $Y=0
+ $X2=1.735 $Y2=0
r201 69 71 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=1.865 $Y=0 $X2=2.16
+ $Y2=0
r202 68 114 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.99 $Y=0
+ $X2=4.115 $Y2=0
r203 68 74 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=3.99 $Y=0 $X2=3.6
+ $Y2=0
r204 66 109 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0
+ $X2=0.72 $Y2=0
r205 65 66 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r206 63 108 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.545 $Y=0
+ $X2=0.67 $Y2=0
r207 63 65 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.545 $Y=0
+ $X2=0.24 $Y2=0
r208 61 88 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=6.48 $Y=0
+ $X2=7.92 $Y2=0
r209 61 124 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=0 $X2=6
+ $Y2=0
r210 61 84 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.48 $Y=0 $X2=6.48
+ $Y2=0
r211 59 96 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=10.605 $Y=0
+ $X2=10.32 $Y2=0
r212 59 60 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=10.605 $Y=0
+ $X2=10.73 $Y2=0
r213 58 100 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=10.855 $Y=0
+ $X2=11.28 $Y2=0
r214 58 60 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=10.855 $Y=0
+ $X2=10.73 $Y2=0
r215 54 140 3.13065 $w=2.5e-07 $l=1.09864e-07 $layer=LI1_cond $X=12.72 $Y=0.085
+ $X2=12.777 $Y2=0
r216 54 56 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=12.72 $Y=0.085
+ $X2=12.72 $Y2=0.515
r217 50 137 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=11.75 $Y=0.085
+ $X2=11.75 $Y2=0
r218 50 52 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=11.75 $Y=0.085
+ $X2=11.75 $Y2=0.515
r219 46 60 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=10.73 $Y=0.085
+ $X2=10.73 $Y2=0
r220 46 48 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=10.73 $Y=0.085
+ $X2=10.73 $Y2=0.515
r221 42 134 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.83 $Y=0.085
+ $X2=9.83 $Y2=0
r222 42 44 20.6043 $w=3.28e-07 $l=5.9e-07 $layer=LI1_cond $X=9.83 $Y=0.085
+ $X2=9.83 $Y2=0.675
r223 38 114 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.115 $Y=0.085
+ $X2=4.115 $Y2=0
r224 38 40 26.2757 $w=2.48e-07 $l=5.7e-07 $layer=LI1_cond $X=4.115 $Y=0.085
+ $X2=4.115 $Y2=0.655
r225 34 111 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=1.735 $Y=0.085
+ $X2=1.735 $Y2=0
r226 34 36 18.6164 $w=2.58e-07 $l=4.2e-07 $layer=LI1_cond $X=1.735 $Y=0.085
+ $X2=1.735 $Y2=0.505
r227 33 108 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.795 $Y=0
+ $X2=0.67 $Y2=0
r228 32 111 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.605 $Y=0
+ $X2=1.735 $Y2=0
r229 32 33 52.8449 $w=1.68e-07 $l=8.1e-07 $layer=LI1_cond $X=1.605 $Y=0
+ $X2=0.795 $Y2=0
r230 28 108 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.67 $Y=0.085
+ $X2=0.67 $Y2=0
r231 28 30 22.8184 $w=2.48e-07 $l=4.95e-07 $layer=LI1_cond $X=0.67 $Y=0.085
+ $X2=0.67 $Y2=0.58
r232 9 56 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=12.54
+ $Y=0.37 $X2=12.68 $Y2=0.515
r233 8 52 91 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=2 $X=11.54
+ $Y=0.37 $X2=11.75 $Y2=0.515
r234 7 48 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=10.55
+ $Y=0.37 $X2=10.69 $Y2=0.515
r235 6 44 182 $w=1.7e-07 $l=3.70473e-07 $layer=licon1_NDIFF $count=1 $X=9.685
+ $Y=0.37 $X2=9.83 $Y2=0.675
r236 5 131 91 $w=1.7e-07 $l=6.76166e-07 $layer=licon1_NDIFF $count=2 $X=8.045
+ $Y=0.59 $X2=8.68 $Y2=0.505
r237 4 121 91 $w=1.7e-07 $l=6.98749e-07 $layer=licon1_NDIFF $count=2 $X=5.365
+ $Y=0.37 $X2=5.995 $Y2=0.515
r238 3 40 182 $w=1.7e-07 $l=2.29565e-07 $layer=licon1_NDIFF $count=1 $X=4.015
+ $Y=0.485 $X2=4.155 $Y2=0.655
r239 2 36 91 $w=1.7e-07 $l=1.96214e-07 $layer=licon1_NDIFF $count=2 $X=1.56
+ $Y=0.37 $X2=1.7 $Y2=0.505
r240 1 30 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.37 $X2=0.71 $Y2=0.58
.ends

