* File: sky130_fd_sc_hs__dlclkp_4.spice
* Created: Tue Sep  1 20:01:33 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hs__dlclkp_4.pex.spice"
.subckt sky130_fd_sc_hs__dlclkp_4  VNB VPB GATE CLK VPWR GCLK VGND
* 
* VGND	VGND
* GCLK	GCLK
* VPWR	VPWR
* CLK	CLK
* GATE	GATE
* VPB	VPB
* VNB	VNB
MM1021 N_VGND_M1021_d N_A_84_48#_M1021_g N_A_27_74#_M1021_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.258437 AS=0.2109 PD=1.55507 PS=2.05 NRD=4.044 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75001.8 A=0.111 P=1.78 MULT=1
MM1017 A_286_80# N_GATE_M1017_g N_VGND_M1021_d VNB NLOWVT L=0.15 W=0.64
+ AD=0.0768 AS=0.223513 PD=0.88 PS=1.34493 NRD=12.18 NRS=75.936 M=1 R=4.26667
+ SA=75001.1 SB=75001.2 A=0.096 P=1.58 MULT=1
MM1018 N_A_84_48#_M1018_d N_A_334_54#_M1018_g A_286_80# VNB NLOWVT L=0.15 W=0.64
+ AD=0.156196 AS=0.0768 PD=1.35849 PS=0.88 NRD=18.744 NRS=12.18 M=1 R=4.26667
+ SA=75001.5 SB=75000.8 A=0.096 P=1.58 MULT=1
MM1012 A_491_124# N_A_334_338#_M1012_g N_A_84_48#_M1018_d VNB NLOWVT L=0.15
+ W=0.42 AD=0.118875 AS=0.102504 PD=1.195 PS=0.891509 NRD=65.148 NRS=30 M=1
+ R=2.8 SA=75002.1 SB=75000.5 A=0.063 P=1.14 MULT=1
MM1000 N_VGND_M1000_d N_A_27_74#_M1000_g A_491_124# VNB NLOWVT L=0.15 W=0.42
+ AD=0.11894 AS=0.118875 PD=0.945 PS=1.195 NRD=65.196 NRS=65.148 M=1 R=2.8
+ SA=75000.8 SB=75000.9 A=0.063 P=1.14 MULT=1
MM1025 N_A_334_338#_M1025_d N_A_334_54#_M1025_g N_VGND_M1000_d VNB NLOWVT L=0.15
+ W=0.74 AD=0.2675 AS=0.20956 PD=2.66 PS=1.665 NRD=49.692 NRS=0 M=1 R=4.93333
+ SA=75001 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1019 N_VGND_M1019_d N_CLK_M1019_g N_A_334_54#_M1019_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.2333 PD=1.02 PS=2.19 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75000.2
+ SB=75001 A=0.111 P=1.78 MULT=1
MM1005 A_1047_74# N_CLK_M1005_g N_VGND_M1019_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.0888 AS=0.1036 PD=0.98 PS=1.02 NRD=10.536 NRS=0 M=1 R=4.93333 SA=75000.7
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1023 N_A_1044_368#_M1023_d N_A_27_74#_M1023_g A_1047_74# VNB NLOWVT L=0.15
+ W=0.74 AD=0.2109 AS=0.0888 PD=2.05 PS=0.98 NRD=0 NRS=10.536 M=1 R=4.93333
+ SA=75001.1 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1006 N_GCLK_M1006_d N_A_1044_368#_M1006_g N_VGND_M1006_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.2977 PD=1.02 PS=2.9 NRD=0 NRS=56.316 M=1 R=4.93333
+ SA=75000.2 SB=75001.6 A=0.111 P=1.78 MULT=1
MM1008 N_GCLK_M1006_d N_A_1044_368#_M1008_g N_VGND_M1008_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.1295 PD=1.02 PS=1.09 NRD=0 NRS=11.34 M=1 R=4.93333
+ SA=75000.6 SB=75001.1 A=0.111 P=1.78 MULT=1
MM1013 N_GCLK_M1013_d N_A_1044_368#_M1013_g N_VGND_M1008_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.1295 PD=1.02 PS=1.09 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75001.1 SB=75000.6 A=0.111 P=1.78 MULT=1
MM1015 N_GCLK_M1013_d N_A_1044_368#_M1015_g N_VGND_M1015_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.2109 PD=1.02 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75001.6 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1011 N_VPWR_M1011_d N_A_84_48#_M1011_g N_A_27_74#_M1011_s VPB PSHORT L=0.15
+ W=1.12 AD=0.328498 AS=0.3304 PD=1.80679 PS=2.83 NRD=26.3783 NRS=1.7533 M=1
+ R=7.46667 SA=75000.2 SB=75001.9 A=0.168 P=2.54 MULT=1
MM1002 A_283_392# N_GATE_M1002_g N_VPWR_M1011_d VPB PSHORT L=0.15 W=1 AD=0.135
+ AS=0.293302 PD=1.27 PS=1.61321 NRD=15.7403 NRS=31.5003 M=1 R=6.66667 SA=75001
+ SB=75001.4 A=0.15 P=2.3 MULT=1
MM1009 N_A_84_48#_M1009_d N_A_334_338#_M1009_g A_283_392# VPB PSHORT L=0.15 W=1
+ AD=0.296056 AS=0.135 PD=2.30282 PS=1.27 NRD=34.4553 NRS=15.7403 M=1 R=6.66667
+ SA=75001.4 SB=75001 A=0.15 P=2.3 MULT=1
MM1003 A_524_508# N_A_334_54#_M1003_g N_A_84_48#_M1009_d VPB PSHORT L=0.15
+ W=0.42 AD=0.0567 AS=0.124344 PD=0.69 PS=0.967183 NRD=37.5088 NRS=84.4145 M=1
+ R=2.8 SA=75002.2 SB=75001.3 A=0.063 P=1.14 MULT=1
MM1010 N_VPWR_M1010_d N_A_27_74#_M1010_g A_524_508# VPB PSHORT L=0.15 W=0.42
+ AD=0.1232 AS=0.0567 PD=1.01333 PS=0.69 NRD=46.886 NRS=37.5088 M=1 R=2.8
+ SA=75002.6 SB=75000.8 A=0.063 P=1.14 MULT=1
MM1004 N_A_334_338#_M1004_d N_A_334_54#_M1004_g N_VPWR_M1010_d VPB PSHORT L=0.15
+ W=0.84 AD=0.2478 AS=0.2464 PD=2.27 PS=2.02667 NRD=0 NRS=55.8889 M=1 R=5.6
+ SA=75001.7 SB=75000.2 A=0.126 P=1.98 MULT=1
MM1016 N_VPWR_M1016_d N_CLK_M1016_g N_A_334_54#_M1016_s VPB PSHORT L=0.15 W=0.84
+ AD=0.1812 AS=0.2478 PD=1.30286 PS=2.27 NRD=22.261 NRS=2.3443 M=1 R=5.6
+ SA=75000.2 SB=75003.8 A=0.126 P=1.98 MULT=1
MM1014 N_A_1044_368#_M1014_d N_CLK_M1014_g N_VPWR_M1016_d VPB PSHORT L=0.15
+ W=1.12 AD=0.1876 AS=0.2416 PD=1.455 PS=1.73714 NRD=7.8997 NRS=4.3931 M=1
+ R=7.46667 SA=75000.6 SB=75003.2 A=0.168 P=2.54 MULT=1
MM1007 N_VPWR_M1007_d N_A_27_74#_M1007_g N_A_1044_368#_M1014_d VPB PSHORT L=0.15
+ W=1.12 AD=0.5348 AS=0.1876 PD=2.075 PS=1.455 NRD=10.5395 NRS=1.7533 M=1
+ R=7.46667 SA=75001.1 SB=75002.7 A=0.168 P=2.54 MULT=1
MM1001 N_VPWR_M1007_d N_A_1044_368#_M1001_g N_GCLK_M1001_s VPB PSHORT L=0.15
+ W=1.12 AD=0.5348 AS=0.1764 PD=2.075 PS=1.435 NRD=10.5395 NRS=1.7533 M=1
+ R=7.46667 SA=75002.2 SB=75001.6 A=0.168 P=2.54 MULT=1
MM1020 N_VPWR_M1020_d N_A_1044_368#_M1020_g N_GCLK_M1001_s VPB PSHORT L=0.15
+ W=1.12 AD=0.1876 AS=0.1764 PD=1.455 PS=1.435 NRD=7.8997 NRS=4.3931 M=1
+ R=7.46667 SA=75002.7 SB=75001.2 A=0.168 P=2.54 MULT=1
MM1022 N_VPWR_M1020_d N_A_1044_368#_M1022_g N_GCLK_M1022_s VPB PSHORT L=0.15
+ W=1.12 AD=0.1876 AS=0.168 PD=1.455 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75003.2 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1024 N_VPWR_M1024_d N_A_1044_368#_M1024_g N_GCLK_M1022_s VPB PSHORT L=0.15
+ W=1.12 AD=0.3304 AS=0.168 PD=2.83 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75003.6 SB=75000.2 A=0.168 P=2.54 MULT=1
DX26_noxref VNB VPB NWDIODE A=16.3897 P=22.3
*
.include "sky130_fd_sc_hs__dlclkp_4.pxi.spice"
*
.ends
*
*
