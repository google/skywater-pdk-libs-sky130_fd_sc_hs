* File: sky130_fd_sc_hs__bufbuf_8.spice
* Created: Tue Sep  1 19:57:12 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hs__bufbuf_8.pex.spice"
.subckt sky130_fd_sc_hs__bufbuf_8  VNB VPB A VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A	A
* VPB	VPB
* VNB	VNB
MM1020 N_VGND_M1020_d N_A_M1020_g N_A_27_112#_M1020_s VNB NLOWVT L=0.15 W=0.55
+ AD=0.129591 AS=0.15675 PD=0.997674 PS=1.67 NRD=17.448 NRS=0 M=1 R=3.66667
+ SA=75000.2 SB=75000.8 A=0.0825 P=1.4 MULT=1
MM1017 N_A_221_368#_M1017_d N_A_27_112#_M1017_g N_VGND_M1020_d VNB NLOWVT L=0.15
+ W=0.74 AD=0.2109 AS=0.174359 PD=2.05 PS=1.34233 NRD=0 NRS=11.34 M=1 R=4.93333
+ SA=75000.7 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1005 N_A_334_368#_M1005_d N_A_221_368#_M1005_g N_VGND_M1005_s VNB NLOWVT
+ L=0.15 W=0.74 AD=0.2109 AS=0.1036 PD=2.05 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75004.8 A=0.111 P=1.78 MULT=1
MM1018 N_A_334_368#_M1018_d N_A_221_368#_M1018_g N_VGND_M1005_s VNB NLOWVT
+ L=0.15 W=0.74 AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.6 SB=75004.4 A=0.111 P=1.78 MULT=1
MM1024 N_A_334_368#_M1018_d N_A_221_368#_M1024_g N_VGND_M1024_s VNB NLOWVT
+ L=0.15 W=0.74 AD=0.1036 AS=0.1295 PD=1.02 PS=1.09 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75001.1 SB=75004 A=0.111 P=1.78 MULT=1
MM1000 N_VGND_M1024_s N_A_334_368#_M1000_g N_X_M1000_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1295 AS=0.1036 PD=1.09 PS=1.02 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75001.6
+ SB=75003.5 A=0.111 P=1.78 MULT=1
MM1002 N_VGND_M1002_d N_A_334_368#_M1002_g N_X_M1000_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1295 AS=0.1036 PD=1.09 PS=1.02 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75002
+ SB=75003.1 A=0.111 P=1.78 MULT=1
MM1007 N_VGND_M1002_d N_A_334_368#_M1007_g N_X_M1007_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1295 AS=0.1036 PD=1.09 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75002.5
+ SB=75002.6 A=0.111 P=1.78 MULT=1
MM1010 N_VGND_M1010_d N_A_334_368#_M1010_g N_X_M1007_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75002.9
+ SB=75002.1 A=0.111 P=1.78 MULT=1
MM1014 N_VGND_M1010_d N_A_334_368#_M1014_g N_X_M1014_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1258 PD=1.02 PS=1.08 NRD=0 NRS=4.86 M=1 R=4.93333 SA=75003.4
+ SB=75001.7 A=0.111 P=1.78 MULT=1
MM1015 N_VGND_M1015_d N_A_334_368#_M1015_g N_X_M1014_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1295 AS=0.1258 PD=1.09 PS=1.08 NRD=0 NRS=4.86 M=1 R=4.93333 SA=75003.8
+ SB=75001.2 A=0.111 P=1.78 MULT=1
MM1023 N_VGND_M1015_d N_A_334_368#_M1023_g N_X_M1023_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1295 AS=0.1036 PD=1.09 PS=1.02 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75004.4
+ SB=75000.7 A=0.111 P=1.78 MULT=1
MM1025 N_VGND_M1025_d N_A_334_368#_M1025_g N_X_M1023_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.25955 AS=0.1036 PD=2.19 PS=1.02 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75004.8
+ SB=75000.3 A=0.111 P=1.78 MULT=1
MM1021 N_VPWR_M1021_d N_A_M1021_g N_A_27_112#_M1021_s VPB PSHORT L=0.15 W=0.84
+ AD=0.1668 AS=0.2478 PD=1.28143 PS=2.27 NRD=4.6886 NRS=2.3443 M=1 R=5.6
+ SA=75000.2 SB=75000.7 A=0.126 P=1.98 MULT=1
MM1022 N_A_221_368#_M1022_d N_A_27_112#_M1022_g N_VPWR_M1021_d VPB PSHORT L=0.15
+ W=1.12 AD=0.3304 AS=0.2224 PD=2.83 PS=1.70857 NRD=1.7533 NRS=13.1793 M=1
+ R=7.46667 SA=75000.6 SB=75000.2 A=0.168 P=2.54 MULT=1
MM1001 N_VPWR_M1001_d N_A_221_368#_M1001_g N_A_334_368#_M1001_s VPB PSHORT
+ L=0.15 W=1.12 AD=0.168 AS=0.3304 PD=1.42 PS=2.83 NRD=1.7533 NRS=1.7533 M=1
+ R=7.46667 SA=75000.2 SB=75004.8 A=0.168 P=2.54 MULT=1
MM1003 N_VPWR_M1001_d N_A_221_368#_M1003_g N_A_334_368#_M1003_s VPB PSHORT
+ L=0.15 W=1.12 AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1
+ R=7.46667 SA=75000.7 SB=75004.4 A=0.168 P=2.54 MULT=1
MM1008 N_VPWR_M1008_d N_A_221_368#_M1008_g N_A_334_368#_M1003_s VPB PSHORT
+ L=0.15 W=1.12 AD=0.196 AS=0.168 PD=1.47 PS=1.42 NRD=10.5395 NRS=1.7533 M=1
+ R=7.46667 SA=75001.1 SB=75003.9 A=0.168 P=2.54 MULT=1
MM1004 N_VPWR_M1008_d N_A_334_368#_M1004_g N_X_M1004_s VPB PSHORT L=0.15 W=1.12
+ AD=0.196 AS=0.196 PD=1.47 PS=1.47 NRD=1.7533 NRS=10.5395 M=1 R=7.46667
+ SA=75001.6 SB=75003.4 A=0.168 P=2.54 MULT=1
MM1006 N_VPWR_M1006_d N_A_334_368#_M1006_g N_X_M1004_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.196 PD=1.42 PS=1.47 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75002.1 SB=75002.9 A=0.168 P=2.54 MULT=1
MM1009 N_VPWR_M1006_d N_A_334_368#_M1009_g N_X_M1009_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75002.6 SB=75002.5 A=0.168 P=2.54 MULT=1
MM1011 N_VPWR_M1011_d N_A_334_368#_M1011_g N_X_M1009_s VPB PSHORT L=0.15 W=1.12
+ AD=0.1708 AS=0.168 PD=1.425 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75003 SB=75002 A=0.168 P=2.54 MULT=1
MM1012 N_VPWR_M1011_d N_A_334_368#_M1012_g N_X_M1012_s VPB PSHORT L=0.15 W=1.12
+ AD=0.1708 AS=0.168 PD=1.425 PS=1.42 NRD=2.6201 NRS=1.7533 M=1 R=7.46667
+ SA=75003.5 SB=75001.6 A=0.168 P=2.54 MULT=1
MM1013 N_VPWR_M1013_d N_A_334_368#_M1013_g N_X_M1012_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75003.9 SB=75001.1 A=0.168 P=2.54 MULT=1
MM1016 N_VPWR_M1013_d N_A_334_368#_M1016_g N_X_M1016_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75004.4 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1019 N_VPWR_M1019_d N_A_334_368#_M1019_g N_X_M1016_s VPB PSHORT L=0.15 W=1.12
+ AD=0.3136 AS=0.168 PD=2.8 PS=1.42 NRD=2.6201 NRS=1.7533 M=1 R=7.46667
+ SA=75004.8 SB=75000.2 A=0.168 P=2.54 MULT=1
DX26_noxref VNB VPB NWDIODE A=14.0988 P=18.88
*
.include "sky130_fd_sc_hs__bufbuf_8.pxi.spice"
*
.ends
*
*
