* File: sky130_fd_sc_hs__einvn_2.pex.spice
* Created: Tue Sep  1 20:04:39 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HS__EINVN_2%A_115_464# 1 2 7 11 13 17 19 22 25 29 32 36
+ 39
c61 17 0 2.14956e-19 $X=1.945 $Y=0.74
c62 13 0 2.02228e-20 $X=1.87 $Y=1.395
r63 37 39 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=0.995 $Y=1.485
+ $X2=0.995 $Y2=1.395
r64 36 37 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.995
+ $Y=1.485 $X2=0.995 $Y2=1.485
r65 33 36 6.63528 $w=3.28e-07 $l=1.9e-07 $layer=LI1_cond $X=0.805 $Y=1.485
+ $X2=0.995 $Y2=1.485
r66 29 31 10.7321 $w=3.28e-07 $l=2.3e-07 $layer=LI1_cond $X=0.725 $Y=0.58
+ $X2=0.725 $Y2=0.81
r67 26 33 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.805 $Y=1.65
+ $X2=0.805 $Y2=1.485
r68 26 32 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=0.805 $Y=1.65
+ $X2=0.805 $Y2=2.3
r69 25 33 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.805 $Y=1.32
+ $X2=0.805 $Y2=1.485
r70 25 31 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=0.805 $Y=1.32
+ $X2=0.805 $Y2=0.81
r71 22 32 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=0.725 $Y=2.465
+ $X2=0.725 $Y2=2.3
r72 15 17 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=1.945 $Y=1.32
+ $X2=1.945 $Y2=0.74
r73 14 19 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.59 $Y=1.395
+ $X2=1.515 $Y2=1.395
r74 13 15 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.87 $Y=1.395
+ $X2=1.945 $Y2=1.32
r75 13 14 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=1.87 $Y=1.395
+ $X2=1.59 $Y2=1.395
r76 9 19 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.515 $Y=1.32
+ $X2=1.515 $Y2=1.395
r77 9 11 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=1.515 $Y=1.32
+ $X2=1.515 $Y2=0.74
r78 8 39 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.16 $Y=1.395
+ $X2=0.995 $Y2=1.395
r79 7 19 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.44 $Y=1.395
+ $X2=1.515 $Y2=1.395
r80 7 8 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=1.44 $Y=1.395 $X2=1.16
+ $Y2=1.395
r81 2 22 300 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=2 $X=0.575
+ $Y=2.32 $X2=0.725 $Y2=2.465
r82 1 29 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=0.585
+ $Y=0.37 $X2=0.725 $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_HS__EINVN_2%TE_B 2 3 6 9 11 12 13 15 16 18 20 21 22 23
+ 27 28
r65 31 32 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=0.385
+ $Y=1.965 $X2=0.385 $Y2=1.965
r66 27 29 46.6671 $w=3.65e-07 $l=1.65e-07 $layer=POLY_cond $X=0.402 $Y=1.285
+ $X2=0.402 $Y2=1.12
r67 27 28 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=0.385
+ $Y=1.285 $X2=0.385 $Y2=1.285
r68 23 32 8.13489 $w=4.23e-07 $l=3e-07 $layer=LI1_cond $X=0.337 $Y=1.665
+ $X2=0.337 $Y2=1.965
r69 22 23 10.033 $w=4.23e-07 $l=3.7e-07 $layer=LI1_cond $X=0.337 $Y=1.295
+ $X2=0.337 $Y2=1.665
r70 22 28 0.271163 $w=4.23e-07 $l=1e-08 $layer=LI1_cond $X=0.337 $Y=1.295
+ $X2=0.337 $Y2=1.285
r71 18 20 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.955 $Y=3.035
+ $X2=1.955 $Y2=2.4
r72 17 21 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.58 $Y=3.11
+ $X2=1.505 $Y2=3.11
r73 16 18 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.88 $Y=3.11
+ $X2=1.955 $Y2=3.035
r74 16 17 153.83 $w=1.5e-07 $l=3e-07 $layer=POLY_cond $X=1.88 $Y=3.11 $X2=1.58
+ $Y2=3.11
r75 13 21 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.505 $Y=3.035
+ $X2=1.505 $Y2=3.11
r76 13 15 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.505 $Y=3.035
+ $X2=1.505 $Y2=2.4
r77 11 21 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.43 $Y=3.11
+ $X2=1.505 $Y2=3.11
r78 11 12 438.415 $w=1.5e-07 $l=8.55e-07 $layer=POLY_cond $X=1.43 $Y=3.11
+ $X2=0.575 $Y2=3.11
r79 9 29 276.894 $w=1.5e-07 $l=5.4e-07 $layer=POLY_cond $X=0.51 $Y=0.58 $X2=0.51
+ $Y2=1.12
r80 4 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.5 $Y=3.035
+ $X2=0.575 $Y2=3.11
r81 4 6 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=0.5 $Y=3.035 $X2=0.5
+ $Y2=2.64
r82 3 31 57.6553 $w=2.91e-07 $l=3.25331e-07 $layer=POLY_cond $X=0.5 $Y=2.245
+ $X2=0.402 $Y2=1.965
r83 3 6 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=0.5 $Y=2.245 $X2=0.5
+ $Y2=2.64
r84 2 31 4.36393 $w=3.65e-07 $l=1.7e-08 $layer=POLY_cond $X=0.402 $Y=1.948
+ $X2=0.402 $Y2=1.965
r85 1 27 2.68759 $w=3.65e-07 $l=1.7e-08 $layer=POLY_cond $X=0.402 $Y=1.302
+ $X2=0.402 $Y2=1.285
r86 1 2 102.129 $w=3.65e-07 $l=6.46e-07 $layer=POLY_cond $X=0.402 $Y=1.302
+ $X2=0.402 $Y2=1.948
.ends

.subckt PM_SKY130_FD_SC_HS__EINVN_2%A 1 3 5 6 8 9 11 13 14 16 17 18 19
c50 6 0 2.66534e-19 $X=2.405 $Y=1.765
r51 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.09
+ $Y=1.385 $X2=3.09 $Y2=1.385
r52 22 24 11.2675 $w=3.85e-07 $l=9e-08 $layer=POLY_cond $X=2.995 $Y=1.295
+ $X2=2.995 $Y2=1.385
r53 19 25 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=3.09 $Y=1.295 $X2=3.09
+ $Y2=1.385
r54 18 19 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=3.09 $Y=0.925
+ $X2=3.09 $Y2=1.295
r55 14 24 66.2218 $w=3.85e-07 $l=4.44522e-07 $layer=POLY_cond $X=2.855 $Y=1.765
+ $X2=2.995 $Y2=1.385
r56 14 16 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.855 $Y=1.765
+ $X2=2.855 $Y2=2.4
r57 11 22 28.0374 $w=3.85e-07 $l=2.19317e-07 $layer=POLY_cond $X=2.81 $Y=1.22
+ $X2=2.995 $Y2=1.295
r58 11 13 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=2.81 $Y=1.22 $X2=2.81
+ $Y2=0.74
r59 10 17 6.66866 $w=1.5e-07 $l=9.8e-08 $layer=POLY_cond $X=2.495 $Y=1.295
+ $X2=2.397 $Y2=1.295
r60 9 22 24.9301 $w=1.5e-07 $l=2.6e-07 $layer=POLY_cond $X=2.735 $Y=1.295
+ $X2=2.995 $Y2=1.295
r61 9 10 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=2.735 $Y=1.295
+ $X2=2.495 $Y2=1.295
r62 6 8 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.405 $Y=1.765
+ $X2=2.405 $Y2=2.4
r63 5 6 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=2.405 $Y=1.675 $X2=2.405
+ $Y2=1.765
r64 4 17 18.8402 $w=1.65e-07 $l=7.88987e-08 $layer=POLY_cond $X=2.405 $Y=1.37
+ $X2=2.397 $Y2=1.295
r65 4 5 118.556 $w=1.8e-07 $l=3.05e-07 $layer=POLY_cond $X=2.405 $Y=1.37
+ $X2=2.405 $Y2=1.675
r66 1 17 18.8402 $w=1.65e-07 $l=8.52936e-08 $layer=POLY_cond $X=2.375 $Y=1.22
+ $X2=2.397 $Y2=1.295
r67 1 3 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=2.375 $Y=1.22 $X2=2.375
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HS__EINVN_2%VPWR 1 2 7 9 13 15 17 27 28 34
c39 13 0 9.65954e-20 $X=1.73 $Y=2.325
r40 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r41 27 28 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r42 25 28 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=3.12 $Y2=3.33
r43 24 27 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=2.16 $Y=3.33 $X2=3.12
+ $Y2=3.33
r44 24 25 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r45 22 34 6.70225 $w=1.7e-07 $l=1.18e-07 $layer=LI1_cond $X=1.815 $Y=3.33
+ $X2=1.697 $Y2=3.33
r46 22 24 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.815 $Y=3.33
+ $X2=2.16 $Y2=3.33
r47 21 32 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.24 $Y2=3.33
r48 20 21 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r49 18 31 4.01803 $w=1.7e-07 $l=1.8e-07 $layer=LI1_cond $X=0.36 $Y=3.33 $X2=0.18
+ $Y2=3.33
r50 18 20 54.8021 $w=1.68e-07 $l=8.4e-07 $layer=LI1_cond $X=0.36 $Y=3.33 $X2=1.2
+ $Y2=3.33
r51 17 34 6.70225 $w=1.7e-07 $l=1.17e-07 $layer=LI1_cond $X=1.58 $Y=3.33
+ $X2=1.697 $Y2=3.33
r52 17 20 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=1.58 $Y=3.33 $X2=1.2
+ $Y2=3.33
r53 15 25 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r54 15 21 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r55 15 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r56 11 34 0.207053 $w=2.35e-07 $l=8.5e-08 $layer=LI1_cond $X=1.697 $Y=3.245
+ $X2=1.697 $Y2=3.33
r57 11 13 45.1169 $w=2.33e-07 $l=9.2e-07 $layer=LI1_cond $X=1.697 $Y=3.245
+ $X2=1.697 $Y2=2.325
r58 7 31 3.12513 $w=2.5e-07 $l=1.09087e-07 $layer=LI1_cond $X=0.235 $Y=3.245
+ $X2=0.18 $Y2=3.33
r59 7 9 35.9562 $w=2.48e-07 $l=7.8e-07 $layer=LI1_cond $X=0.235 $Y=3.245
+ $X2=0.235 $Y2=2.465
r60 2 13 300 $w=1.7e-07 $l=5.54955e-07 $layer=licon1_PDIFF $count=2 $X=1.58
+ $Y=1.84 $X2=1.73 $Y2=2.325
r61 1 9 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=2.32 $X2=0.275 $Y2=2.465
.ends

.subckt PM_SKY130_FD_SC_HS__EINVN_2%A_227_368# 1 2 3 10 12 14 16 19 20 21 24
c48 16 0 1.90161e-19 $X=2.155 $Y=1.99
r49 24 27 34.1617 $w=2.78e-07 $l=8.3e-07 $layer=LI1_cond $X=3.105 $Y=1.985
+ $X2=3.105 $Y2=2.815
r50 22 27 3.70428 $w=2.78e-07 $l=9e-08 $layer=LI1_cond $X=3.105 $Y=2.905
+ $X2=3.105 $Y2=2.815
r51 20 22 7.36005 $w=1.7e-07 $l=1.77482e-07 $layer=LI1_cond $X=2.965 $Y=2.99
+ $X2=3.105 $Y2=2.905
r52 20 21 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.965 $Y=2.99
+ $X2=2.295 $Y2=2.99
r53 17 21 7.36005 $w=1.7e-07 $l=1.77482e-07 $layer=LI1_cond $X=2.155 $Y=2.905
+ $X2=2.295 $Y2=2.99
r54 17 19 3.70428 $w=2.78e-07 $l=9e-08 $layer=LI1_cond $X=2.155 $Y=2.905
+ $X2=2.155 $Y2=2.815
r55 16 31 2.78046 $w=2.8e-07 $l=8.5e-08 $layer=LI1_cond $X=2.155 $Y=1.99
+ $X2=2.155 $Y2=1.905
r56 16 19 33.9559 $w=2.78e-07 $l=8.25e-07 $layer=LI1_cond $X=2.155 $Y=1.99
+ $X2=2.155 $Y2=2.815
r57 15 29 4.64039 $w=1.7e-07 $l=1.43e-07 $layer=LI1_cond $X=1.4 $Y=1.905
+ $X2=1.257 $Y2=1.905
r58 14 31 4.57959 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=2.015 $Y=1.905
+ $X2=2.155 $Y2=1.905
r59 14 15 40.123 $w=1.68e-07 $l=6.15e-07 $layer=LI1_cond $X=2.015 $Y=1.905
+ $X2=1.4 $Y2=1.905
r60 10 29 2.75828 $w=2.85e-07 $l=8.5e-08 $layer=LI1_cond $X=1.257 $Y=1.99
+ $X2=1.257 $Y2=1.905
r61 10 12 33.3602 $w=2.83e-07 $l=8.25e-07 $layer=LI1_cond $X=1.257 $Y=1.99
+ $X2=1.257 $Y2=2.815
r62 3 27 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=2.93
+ $Y=1.84 $X2=3.08 $Y2=2.815
r63 3 24 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=2.93
+ $Y=1.84 $X2=3.08 $Y2=1.985
r64 2 31 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=2.03
+ $Y=1.84 $X2=2.18 $Y2=1.985
r65 2 19 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=2.03
+ $Y=1.84 $X2=2.18 $Y2=2.815
r66 1 29 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=1.135
+ $Y=1.84 $X2=1.28 $Y2=1.985
r67 1 12 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=1.135
+ $Y=1.84 $X2=1.28 $Y2=2.815
.ends

.subckt PM_SKY130_FD_SC_HS__EINVN_2%Z 1 2 7 8 9 10 24
c29 7 0 5.33156e-20 $X=2.64 $Y=0.925
r30 22 24 1.74613 $w=3.28e-07 $l=5e-08 $layer=LI1_cond $X=2.63 $Y=1.985 $X2=2.63
+ $Y2=2.035
r31 10 22 0.628605 $w=3.28e-07 $l=1.8e-08 $layer=LI1_cond $X=2.63 $Y=1.967
+ $X2=2.63 $Y2=1.985
r32 10 35 5.33231 $w=3.28e-07 $l=1.47e-07 $layer=LI1_cond $X=2.63 $Y=1.967
+ $X2=2.63 $Y2=1.82
r33 10 27 20.8837 $w=3.28e-07 $l=5.98e-07 $layer=LI1_cond $X=2.63 $Y=2.052
+ $X2=2.63 $Y2=2.65
r34 10 24 0.593683 $w=3.28e-07 $l=1.7e-08 $layer=LI1_cond $X=2.63 $Y=2.052
+ $X2=2.63 $Y2=2.035
r35 9 35 6.15961 $w=2.88e-07 $l=1.55e-07 $layer=LI1_cond $X=2.61 $Y=1.665
+ $X2=2.61 $Y2=1.82
r36 8 9 14.7036 $w=2.88e-07 $l=3.7e-07 $layer=LI1_cond $X=2.61 $Y=1.295 $X2=2.61
+ $Y2=1.665
r37 8 33 6.557 $w=2.88e-07 $l=1.65e-07 $layer=LI1_cond $X=2.61 $Y=1.295 $X2=2.61
+ $Y2=1.13
r38 7 33 7.88165 $w=3.28e-07 $l=2.2e-07 $layer=LI1_cond $X=2.59 $Y=0.91 $X2=2.59
+ $Y2=1.13
r39 2 10 400 $w=1.7e-07 $l=2.04939e-07 $layer=licon1_PDIFF $count=1 $X=2.48
+ $Y=1.84 $X2=2.63 $Y2=1.97
r40 2 27 400 $w=1.7e-07 $l=8.81816e-07 $layer=licon1_PDIFF $count=1 $X=2.48
+ $Y=1.84 $X2=2.63 $Y2=2.65
r41 1 7 182 $w=1.7e-07 $l=6.0597e-07 $layer=licon1_NDIFF $count=1 $X=2.45
+ $Y=0.37 $X2=2.59 $Y2=0.91
.ends

.subckt PM_SKY130_FD_SC_HS__EINVN_2%VGND 1 2 7 9 13 15 17 27 28 34
r37 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r38 27 28 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r39 25 28 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=3.12
+ $Y2=0
r40 24 27 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=2.16 $Y=0 $X2=3.12
+ $Y2=0
r41 24 25 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r42 22 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.895 $Y=0 $X2=1.73
+ $Y2=0
r43 22 24 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=1.895 $Y=0 $X2=2.16
+ $Y2=0
r44 21 32 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.24
+ $Y2=0
r45 20 21 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r46 18 31 3.99177 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.38 $Y=0 $X2=0.19
+ $Y2=0
r47 18 20 53.4973 $w=1.68e-07 $l=8.2e-07 $layer=LI1_cond $X=0.38 $Y=0 $X2=1.2
+ $Y2=0
r48 17 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.565 $Y=0 $X2=1.73
+ $Y2=0
r49 17 20 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=1.565 $Y=0 $X2=1.2
+ $Y2=0
r50 15 25 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r51 15 21 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r52 15 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r53 11 34 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.73 $Y=0.085
+ $X2=1.73 $Y2=0
r54 11 13 18.3343 $w=3.28e-07 $l=5.25e-07 $layer=LI1_cond $X=1.73 $Y=0.085
+ $X2=1.73 $Y2=0.61
r55 7 31 3.1514 $w=2.5e-07 $l=1.12916e-07 $layer=LI1_cond $X=0.255 $Y=0.085
+ $X2=0.19 $Y2=0
r56 7 9 22.8184 $w=2.48e-07 $l=4.95e-07 $layer=LI1_cond $X=0.255 $Y=0.085
+ $X2=0.255 $Y2=0.58
r57 2 13 182 $w=1.7e-07 $l=3.01993e-07 $layer=licon1_NDIFF $count=1 $X=1.59
+ $Y=0.37 $X2=1.73 $Y2=0.61
r58 1 9 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=0.15
+ $Y=0.37 $X2=0.295 $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_HS__EINVN_2%A_231_74# 1 2 3 12 14 15 16 22
c42 16 0 1.6164e-19 $X=2.16 $Y=0.6
r43 20 25 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.245 $Y=0.475
+ $X2=2.16 $Y2=0.475
r44 20 22 35.9562 $w=2.48e-07 $l=7.8e-07 $layer=LI1_cond $X=2.245 $Y=0.475
+ $X2=3.025 $Y2=0.475
r45 17 19 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=2.16 $Y=0.98
+ $X2=2.16 $Y2=0.965
r46 16 25 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.16 $Y=0.6 $X2=2.16
+ $Y2=0.475
r47 16 19 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=2.16 $Y=0.6
+ $X2=2.16 $Y2=0.965
r48 14 17 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.075 $Y=1.065
+ $X2=2.16 $Y2=0.98
r49 14 15 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=2.075 $Y=1.065
+ $X2=1.385 $Y2=1.065
r50 10 15 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.26 $Y=0.98
+ $X2=1.385 $Y2=1.065
r51 10 12 21.4354 $w=2.48e-07 $l=4.65e-07 $layer=LI1_cond $X=1.26 $Y=0.98
+ $X2=1.26 $Y2=0.515
r52 3 22 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=2.885
+ $Y=0.37 $X2=3.025 $Y2=0.515
r53 2 25 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=2.02
+ $Y=0.37 $X2=2.16 $Y2=0.515
r54 2 19 182 $w=1.7e-07 $l=6.61306e-07 $layer=licon1_NDIFF $count=1 $X=2.02
+ $Y=0.37 $X2=2.16 $Y2=0.965
r55 1 12 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=1.155
+ $Y=0.37 $X2=1.3 $Y2=0.515
.ends

