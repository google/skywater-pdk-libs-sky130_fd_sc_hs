* File: sky130_fd_sc_hs__buf_2.pex.spice
* Created: Tue Sep  1 19:56:48 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HS__BUF_2%A_21_260# 1 2 7 9 12 16 18 20 21 24 28 29 30
+ 31 33 34 35 36 40 44 48 51 53 54
r95 51 52 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.61
+ $Y=1.465 $X2=0.61 $Y2=1.465
r96 46 48 13.7944 $w=3.28e-07 $l=3.95e-07 $layer=LI1_cond $X=2.12 $Y=1.01
+ $X2=2.12 $Y2=0.615
r97 42 54 2.70057 $w=3.55e-07 $l=8.5e-08 $layer=LI1_cond $X=2.107 $Y=2.49
+ $X2=2.107 $Y2=2.405
r98 42 44 7.30422 $w=3.53e-07 $l=2.25e-07 $layer=LI1_cond $X=2.107 $Y=2.49
+ $X2=2.107 $Y2=2.715
r99 38 54 2.70057 $w=3.55e-07 $l=8.5e-08 $layer=LI1_cond $X=2.107 $Y=2.32
+ $X2=2.107 $Y2=2.405
r100 38 40 9.25201 $w=3.53e-07 $l=2.85e-07 $layer=LI1_cond $X=2.107 $Y=2.32
+ $X2=2.107 $Y2=2.035
r101 37 53 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.655 $Y=2.405
+ $X2=1.57 $Y2=2.405
r102 36 54 4.08752 $w=1.7e-07 $l=1.77e-07 $layer=LI1_cond $X=1.93 $Y=2.405
+ $X2=2.107 $Y2=2.405
r103 36 37 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=1.93 $Y=2.405
+ $X2=1.655 $Y2=2.405
r104 34 46 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.955 $Y=1.095
+ $X2=2.12 $Y2=1.01
r105 34 35 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=1.955 $Y=1.095
+ $X2=1.655 $Y2=1.095
r106 33 53 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.57 $Y=2.32
+ $X2=1.57 $Y2=2.405
r107 32 35 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.57 $Y=1.18
+ $X2=1.655 $Y2=1.095
r108 32 33 74.3743 $w=1.68e-07 $l=1.14e-06 $layer=LI1_cond $X=1.57 $Y=1.18
+ $X2=1.57 $Y2=2.32
r109 30 53 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.485 $Y=2.405
+ $X2=1.57 $Y2=2.405
r110 30 31 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=1.485 $Y=2.405
+ $X2=0.775 $Y2=2.405
r111 29 31 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.69 $Y=2.32
+ $X2=0.775 $Y2=2.405
r112 28 51 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.69 $Y=1.63
+ $X2=0.69 $Y2=1.465
r113 28 29 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=0.69 $Y=1.63
+ $X2=0.69 $Y2=2.32
r114 24 25 1.202 $w=4.01e-07 $l=1e-08 $layer=POLY_cond $X=1.325 $Y=1.532
+ $X2=1.335 $Y2=1.532
r115 23 24 51.6858 $w=4.01e-07 $l=4.3e-07 $layer=POLY_cond $X=0.895 $Y=1.532
+ $X2=1.325 $Y2=1.532
r116 22 23 1.202 $w=4.01e-07 $l=1e-08 $layer=POLY_cond $X=0.885 $Y=1.532
+ $X2=0.895 $Y2=1.532
r117 21 52 32.3493 $w=3.3e-07 $l=1.85e-07 $layer=POLY_cond $X=0.795 $Y=1.465
+ $X2=0.61 $Y2=1.465
r118 21 22 12.4716 $w=4.01e-07 $l=1.1887e-07 $layer=POLY_cond $X=0.795 $Y=1.465
+ $X2=0.885 $Y2=1.532
r119 18 25 25.923 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=1.335 $Y=1.765
+ $X2=1.335 $Y2=1.532
r120 18 20 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.335 $Y=1.765
+ $X2=1.335 $Y2=2.4
r121 14 24 25.923 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=1.325 $Y=1.3
+ $X2=1.325 $Y2=1.532
r122 14 16 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=1.325 $Y=1.3
+ $X2=1.325 $Y2=0.74
r123 10 23 25.923 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=0.895 $Y=1.3
+ $X2=0.895 $Y2=1.532
r124 10 12 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=0.895 $Y=1.3
+ $X2=0.895 $Y2=0.74
r125 7 22 25.923 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=0.885 $Y=1.765
+ $X2=0.885 $Y2=1.532
r126 7 9 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.885 $Y=1.765
+ $X2=0.885 $Y2=2.4
r127 2 44 400 $w=1.7e-07 $l=9.51643e-07 $layer=licon1_PDIFF $count=1 $X=1.945
+ $Y=1.84 $X2=2.105 $Y2=2.715
r128 2 40 400 $w=1.7e-07 $l=2.63106e-07 $layer=licon1_PDIFF $count=1 $X=1.945
+ $Y=1.84 $X2=2.105 $Y2=2.035
r129 1 48 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.98
+ $Y=0.47 $X2=2.12 $Y2=0.615
.ends

.subckt PM_SKY130_FD_SC_HS__BUF_2%A 1 3 6 8
r28 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.99
+ $Y=1.515 $X2=1.99 $Y2=1.515
r29 8 12 4.55617 $w=4.28e-07 $l=1.7e-07 $layer=LI1_cond $X=2.16 $Y=1.565
+ $X2=1.99 $Y2=1.565
r30 4 11 38.6365 $w=3.35e-07 $l=1.93533e-07 $layer=POLY_cond $X=1.905 $Y=1.35
+ $X2=1.967 $Y2=1.515
r31 4 6 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=1.905 $Y=1.35
+ $X2=1.905 $Y2=0.79
r32 1 11 50.8664 $w=3.35e-07 $l=2.94534e-07 $layer=POLY_cond $X=1.87 $Y=1.765
+ $X2=1.967 $Y2=1.515
r33 1 3 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=1.87 $Y=1.765
+ $X2=1.87 $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_HS__BUF_2%VPWR 1 2 9 13 16 17 18 20 25 26
r42 33 34 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r43 31 33 1.20395 $w=6.08e-07 $l=6e-08 $layer=LI1_cond $X=0.66 $Y=3.075 $X2=0.72
+ $Y2=3.075
r44 29 31 7.88586 $w=6.08e-07 $l=3.93e-07 $layer=LI1_cond $X=0.267 $Y=3.075
+ $X2=0.66 $Y2=3.075
r45 25 26 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r46 20 33 9.20845 $w=6.08e-07 $l=3.02985e-07 $layer=LI1_cond $X=0.825 $Y=3.33
+ $X2=0.72 $Y2=3.075
r47 20 22 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=0.825 $Y=3.33
+ $X2=1.2 $Y2=3.33
r48 18 26 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.16 $Y2=3.33
r49 18 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r50 18 22 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r51 16 22 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=1.395 $Y=3.33
+ $X2=1.2 $Y2=3.33
r52 16 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.395 $Y=3.33
+ $X2=1.56 $Y2=3.33
r53 15 25 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=1.725 $Y=3.33
+ $X2=2.16 $Y2=3.33
r54 15 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.725 $Y=3.33
+ $X2=1.56 $Y2=3.33
r55 11 17 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.56 $Y=3.245
+ $X2=1.56 $Y2=3.33
r56 11 13 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=1.56 $Y=3.245
+ $X2=1.56 $Y2=2.78
r57 7 29 4.79164 $w=3.05e-07 $l=3.4e-07 $layer=LI1_cond $X=0.267 $Y=2.735
+ $X2=0.267 $Y2=3.075
r58 7 9 28.3388 $w=3.03e-07 $l=7.5e-07 $layer=LI1_cond $X=0.267 $Y=2.735
+ $X2=0.267 $Y2=1.985
r59 2 13 600 $w=1.7e-07 $l=1.01223e-06 $layer=licon1_PDIFF $count=1 $X=1.41
+ $Y=1.84 $X2=1.56 $Y2=2.78
r60 1 31 600 $w=1.7e-07 $l=1.21445e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.66 $Y2=2.82
r61 1 29 600 $w=1.7e-07 $l=1.05e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.82
r62 1 9 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HS__BUF_2%X 1 2 9 11 12 13 30
r19 18 30 2.1803 $w=3.68e-07 $l=7e-08 $layer=LI1_cond $X=1.13 $Y=1.365 $X2=1.13
+ $Y2=1.295
r20 13 23 1.55736 $w=3.68e-07 $l=5e-08 $layer=LI1_cond $X=1.13 $Y=2.035 $X2=1.13
+ $Y2=1.985
r21 12 23 9.96707 $w=3.68e-07 $l=3.2e-07 $layer=LI1_cond $X=1.13 $Y=1.665
+ $X2=1.13 $Y2=1.985
r22 11 30 0.249177 $w=3.68e-07 $l=8e-09 $layer=LI1_cond $X=1.13 $Y=1.287
+ $X2=1.13 $Y2=1.295
r23 11 28 3.49432 $w=3.68e-07 $l=1.07e-07 $layer=LI1_cond $X=1.13 $Y=1.287
+ $X2=1.13 $Y2=1.18
r24 11 12 9.1261 $w=3.68e-07 $l=2.93e-07 $layer=LI1_cond $X=1.13 $Y=1.372
+ $X2=1.13 $Y2=1.665
r25 11 18 0.21803 $w=3.68e-07 $l=7e-09 $layer=LI1_cond $X=1.13 $Y=1.372 $X2=1.13
+ $Y2=1.365
r26 9 28 23.2235 $w=3.28e-07 $l=6.65e-07 $layer=LI1_cond $X=1.11 $Y=0.515
+ $X2=1.11 $Y2=1.18
r27 2 23 600 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=0.96
+ $Y=1.84 $X2=1.11 $Y2=1.985
r28 1 9 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=0.97
+ $Y=0.37 $X2=1.11 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__BUF_2%VGND 1 2 9 13 16 17 18 24 30 31 34
r31 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r32 31 35 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.68
+ $Y2=0
r33 30 31 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r34 28 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.775 $Y=0 $X2=1.61
+ $Y2=0
r35 28 30 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=1.775 $Y=0 $X2=2.16
+ $Y2=0
r36 24 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.445 $Y=0 $X2=1.61
+ $Y2=0
r37 24 26 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=1.445 $Y=0 $X2=1.2
+ $Y2=0
r38 21 22 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r39 18 35 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=1.68
+ $Y2=0
r40 18 22 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.24
+ $Y2=0
r41 18 26 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r42 16 21 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=0.515 $Y=0 $X2=0.24
+ $Y2=0
r43 16 17 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.515 $Y=0 $X2=0.64
+ $Y2=0
r44 15 26 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=0.765 $Y=0 $X2=1.2
+ $Y2=0
r45 15 17 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.765 $Y=0 $X2=0.64
+ $Y2=0
r46 11 34 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.61 $Y=0.085
+ $X2=1.61 $Y2=0
r47 11 13 20.6043 $w=3.28e-07 $l=5.9e-07 $layer=LI1_cond $X=1.61 $Y=0.085
+ $X2=1.61 $Y2=0.675
r48 7 17 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.64 $Y=0.085
+ $X2=0.64 $Y2=0
r49 7 9 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=0.64 $Y=0.085 $X2=0.64
+ $Y2=0.515
r50 2 13 182 $w=1.7e-07 $l=3.96327e-07 $layer=licon1_NDIFF $count=1 $X=1.4
+ $Y=0.37 $X2=1.61 $Y2=0.675
r51 1 9 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.535
+ $Y=0.37 $X2=0.68 $Y2=0.515
.ends

