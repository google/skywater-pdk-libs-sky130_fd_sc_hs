* File: sky130_fd_sc_hs__a22o_2.pex.spice
* Created: Thu Aug 27 20:26:58 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HS__A22O_2%A_81_48# 1 2 7 9 10 12 13 15 16 18 22 23 24
+ 25 26 29 34 35 36 38
c78 23 0 1.25043e-19 $X=2 $Y=1.095
c79 16 0 5.41976e-20 $X=1.325 $Y=1.765
r80 40 41 4.15517 $w=4.06e-07 $l=3.5e-08 $layer=POLY_cond $X=0.875 $Y=1.492
+ $X2=0.91 $Y2=1.492
r81 39 40 46.8941 $w=4.06e-07 $l=3.95e-07 $layer=POLY_cond $X=0.48 $Y=1.492
+ $X2=0.875 $Y2=1.492
r82 35 43 8.90394 $w=4.06e-07 $l=7.5e-08 $layer=POLY_cond $X=1.25 $Y=1.492
+ $X2=1.325 $Y2=1.492
r83 35 41 40.3645 $w=4.06e-07 $l=3.4e-07 $layer=POLY_cond $X=1.25 $Y=1.492
+ $X2=0.91 $Y2=1.492
r84 34 36 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=1.25 $Y=1.385
+ $X2=1.25 $Y2=1.55
r85 34 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.25
+ $Y=1.385 $X2=1.25 $Y2=1.385
r86 27 29 8.73063 $w=3.28e-07 $l=2.5e-07 $layer=LI1_cond $X=2.165 $Y=1.01
+ $X2=2.165 $Y2=0.76
r87 25 38 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.455 $Y=2.035
+ $X2=2.58 $Y2=2.035
r88 25 26 67.8503 $w=1.68e-07 $l=1.04e-06 $layer=LI1_cond $X=2.455 $Y=2.035
+ $X2=1.415 $Y2=2.035
r89 23 27 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2 $Y=1.095
+ $X2=2.165 $Y2=1.01
r90 23 24 38.1658 $w=1.68e-07 $l=5.85e-07 $layer=LI1_cond $X=2 $Y=1.095
+ $X2=1.415 $Y2=1.095
r91 22 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.33 $Y=1.95
+ $X2=1.415 $Y2=2.035
r92 22 36 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=1.33 $Y=1.95 $X2=1.33
+ $Y2=1.55
r93 19 24 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.25 $Y=1.18
+ $X2=1.415 $Y2=1.095
r94 19 34 7.15912 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=1.25 $Y=1.18
+ $X2=1.25 $Y2=1.385
r95 16 43 26.2263 $w=1.5e-07 $l=2.73e-07 $layer=POLY_cond $X=1.325 $Y=1.765
+ $X2=1.325 $Y2=1.492
r96 16 18 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.325 $Y=1.765
+ $X2=1.325 $Y2=2.4
r97 13 41 26.2263 $w=1.5e-07 $l=2.72e-07 $layer=POLY_cond $X=0.91 $Y=1.22
+ $X2=0.91 $Y2=1.492
r98 13 15 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=0.91 $Y=1.22 $X2=0.91
+ $Y2=0.74
r99 10 40 26.2263 $w=1.5e-07 $l=2.73e-07 $layer=POLY_cond $X=0.875 $Y=1.765
+ $X2=0.875 $Y2=1.492
r100 10 12 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.875 $Y=1.765
+ $X2=0.875 $Y2=2.4
r101 7 39 26.2263 $w=1.5e-07 $l=2.72e-07 $layer=POLY_cond $X=0.48 $Y=1.22
+ $X2=0.48 $Y2=1.492
r102 7 9 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=0.48 $Y=1.22 $X2=0.48
+ $Y2=0.74
r103 2 38 300 $w=1.7e-07 $l=3.4187e-07 $layer=licon1_PDIFF $count=2 $X=2.39
+ $Y=1.84 $X2=2.54 $Y2=2.115
r104 1 29 182 $w=1.7e-07 $l=4.83735e-07 $layer=licon1_NDIFF $count=1 $X=1.955
+ $Y=0.37 $X2=2.165 $Y2=0.76
.ends

.subckt PM_SKY130_FD_SC_HS__A22O_2%A1 1 3 6 8 12
c34 12 0 5.41976e-20 $X=1.79 $Y=1.515
r35 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.79
+ $Y=1.515 $X2=1.79 $Y2=1.515
r36 8 12 5.40208 $w=3.18e-07 $l=1.5e-07 $layer=LI1_cond $X=1.745 $Y=1.665
+ $X2=1.745 $Y2=1.515
r37 4 11 38.5562 $w=2.99e-07 $l=2.05122e-07 $layer=POLY_cond $X=1.88 $Y=1.35
+ $X2=1.79 $Y2=1.515
r38 4 6 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.88 $Y=1.35 $X2=1.88
+ $Y2=0.74
r39 1 11 52.2586 $w=2.99e-07 $l=2.85044e-07 $layer=POLY_cond $X=1.865 $Y=1.765
+ $X2=1.79 $Y2=1.515
r40 1 3 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=1.865 $Y=1.765
+ $X2=1.865 $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_HS__A22O_2%B1 1 3 6 8 12
r33 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.33
+ $Y=1.515 $X2=2.33 $Y2=1.515
r34 8 12 4.55617 $w=4.28e-07 $l=1.7e-07 $layer=LI1_cond $X=2.16 $Y=1.565
+ $X2=2.33 $Y2=1.565
r35 4 11 38.5562 $w=2.99e-07 $l=1.88348e-07 $layer=POLY_cond $X=2.38 $Y=1.35
+ $X2=2.33 $Y2=1.515
r36 4 6 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.38 $Y=1.35 $X2=2.38
+ $Y2=0.74
r37 1 11 52.2586 $w=2.99e-07 $l=2.57391e-07 $layer=POLY_cond $X=2.315 $Y=1.765
+ $X2=2.33 $Y2=1.515
r38 1 3 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=2.315 $Y=1.765
+ $X2=2.315 $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_HS__A22O_2%B2 3 5 7 8
c29 3 0 1.25043e-19 $X=2.78 $Y=0.74
r30 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.87
+ $Y=1.515 $X2=2.87 $Y2=1.515
r31 8 12 6.70025 $w=4.28e-07 $l=2.5e-07 $layer=LI1_cond $X=3.12 $Y=1.565
+ $X2=2.87 $Y2=1.565
r32 5 11 52.2586 $w=2.99e-07 $l=2.76134e-07 $layer=POLY_cond $X=2.815 $Y=1.765
+ $X2=2.87 $Y2=1.515
r33 5 7 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=2.815 $Y=1.765
+ $X2=2.815 $Y2=2.34
r34 1 11 38.5562 $w=2.99e-07 $l=2.05122e-07 $layer=POLY_cond $X=2.78 $Y=1.35
+ $X2=2.87 $Y2=1.515
r35 1 3 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.78 $Y=1.35 $X2=2.78
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HS__A22O_2%A2 3 5 7 8 12
r23 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.57
+ $Y=1.515 $X2=3.57 $Y2=1.515
r24 8 12 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=3.57 $Y=1.665
+ $X2=3.57 $Y2=1.515
r25 5 11 49.7466 $w=4.26e-07 $l=3.18198e-07 $layer=POLY_cond $X=3.335 $Y=1.765
+ $X2=3.49 $Y2=1.515
r26 5 7 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=3.335 $Y=1.765
+ $X2=3.335 $Y2=2.34
r27 1 11 40.1292 $w=4.26e-07 $l=2.38642e-07 $layer=POLY_cond $X=3.32 $Y=1.35
+ $X2=3.49 $Y2=1.515
r28 1 3 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=3.32 $Y=1.35 $X2=3.32
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HS__A22O_2%VPWR 1 2 3 12 16 18 20 23 24 25 31 35 41 45
r46 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r47 41 42 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r48 39 45 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=3.6 $Y2=3.33
r49 38 39 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r50 36 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.715 $Y=3.33
+ $X2=1.55 $Y2=3.33
r51 36 38 91.6631 $w=1.68e-07 $l=1.405e-06 $layer=LI1_cond $X=1.715 $Y=3.33
+ $X2=3.12 $Y2=3.33
r52 35 44 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=3.395 $Y=3.33
+ $X2=3.617 $Y2=3.33
r53 35 38 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=3.395 $Y=3.33
+ $X2=3.12 $Y2=3.33
r54 34 42 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=1.68 $Y2=3.33
r55 33 34 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r56 31 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.385 $Y=3.33
+ $X2=1.55 $Y2=3.33
r57 31 33 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=1.385 $Y=3.33
+ $X2=1.2 $Y2=3.33
r58 29 34 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=1.2 $Y2=3.33
r59 28 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r60 25 39 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=3.12 $Y2=3.33
r61 25 42 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=1.68 $Y2=3.33
r62 23 28 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=0.485 $Y=3.33
+ $X2=0.24 $Y2=3.33
r63 23 24 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.485 $Y=3.33
+ $X2=0.61 $Y2=3.33
r64 22 33 30.3369 $w=1.68e-07 $l=4.65e-07 $layer=LI1_cond $X=0.735 $Y=3.33
+ $X2=1.2 $Y2=3.33
r65 22 24 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.735 $Y=3.33
+ $X2=0.61 $Y2=3.33
r66 18 44 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=3.56 $Y=3.245
+ $X2=3.617 $Y2=3.33
r67 18 20 39.4624 $w=3.28e-07 $l=1.13e-06 $layer=LI1_cond $X=3.56 $Y=3.245
+ $X2=3.56 $Y2=2.115
r68 14 41 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.55 $Y=3.245
+ $X2=1.55 $Y2=3.33
r69 14 16 30.3826 $w=3.28e-07 $l=8.7e-07 $layer=LI1_cond $X=1.55 $Y=3.245
+ $X2=1.55 $Y2=2.375
r70 10 24 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.61 $Y=3.245
+ $X2=0.61 $Y2=3.33
r71 10 12 47.0197 $w=2.48e-07 $l=1.02e-06 $layer=LI1_cond $X=0.61 $Y=3.245
+ $X2=0.61 $Y2=2.225
r72 3 20 300 $w=1.7e-07 $l=3.4187e-07 $layer=licon1_PDIFF $count=2 $X=3.41
+ $Y=1.84 $X2=3.56 $Y2=2.115
r73 2 16 300 $w=1.7e-07 $l=6.05372e-07 $layer=licon1_PDIFF $count=2 $X=1.4
+ $Y=1.84 $X2=1.55 $Y2=2.375
r74 1 12 300 $w=1.7e-07 $l=4.43114e-07 $layer=licon1_PDIFF $count=2 $X=0.525
+ $Y=1.84 $X2=0.65 $Y2=2.225
.ends

.subckt PM_SKY130_FD_SC_HS__A22O_2%X 1 2 9 11 13 14 15 16 17 34 38
r29 23 34 1.92074 $w=3.28e-07 $l=5.5e-08 $layer=LI1_cond $X=0.695 $Y=1.72
+ $X2=0.695 $Y2=1.665
r30 17 38 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=0.72 $Y=1.805
+ $X2=0.99 $Y2=1.805
r31 17 23 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=0.72 $Y=1.805
+ $X2=0.695 $Y2=1.805
r32 17 34 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=0.695 $Y=1.65
+ $X2=0.695 $Y2=1.665
r33 16 17 12.3975 $w=3.28e-07 $l=3.55e-07 $layer=LI1_cond $X=0.695 $Y=1.295
+ $X2=0.695 $Y2=1.65
r34 15 16 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=0.695 $Y=0.925
+ $X2=0.695 $Y2=1.295
r35 14 15 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=0.695 $Y=0.515
+ $X2=0.695 $Y2=0.925
r36 9 13 7.52792 $w=2.78e-07 $l=1.4e-07 $layer=LI1_cond $X=1.045 $Y=2.43
+ $X2=1.045 $Y2=2.29
r37 9 11 1.02897 $w=2.78e-07 $l=2.5e-08 $layer=LI1_cond $X=1.045 $Y=2.43
+ $X2=1.045 $Y2=2.455
r38 7 38 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.99 $Y=1.89 $X2=0.99
+ $Y2=1.805
r39 7 13 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=0.99 $Y=1.89 $X2=0.99
+ $Y2=2.29
r40 2 11 300 $w=1.7e-07 $l=6.85912e-07 $layer=licon1_PDIFF $count=2 $X=0.95
+ $Y=1.84 $X2=1.1 $Y2=2.455
r41 1 14 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=0.555
+ $Y=0.37 $X2=0.695 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__A22O_2%A_388_368# 1 2 9 11 12 15
r28 15 18 22.3903 $w=3.48e-07 $l=6.8e-07 $layer=LI1_cond $X=3.05 $Y=2.035
+ $X2=3.05 $Y2=2.715
r29 13 18 6.25612 $w=3.48e-07 $l=1.9e-07 $layer=LI1_cond $X=3.05 $Y=2.905
+ $X2=3.05 $Y2=2.715
r30 11 13 7.93686 $w=1.7e-07 $l=2.13307e-07 $layer=LI1_cond $X=2.875 $Y=2.99
+ $X2=3.05 $Y2=2.905
r31 11 12 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=2.875 $Y=2.99
+ $X2=2.255 $Y2=2.99
r32 7 12 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.09 $Y=2.905
+ $X2=2.255 $Y2=2.99
r33 7 9 18.5089 $w=3.28e-07 $l=5.3e-07 $layer=LI1_cond $X=2.09 $Y=2.905 $X2=2.09
+ $Y2=2.375
r34 2 18 400 $w=1.7e-07 $l=9.51643e-07 $layer=licon1_PDIFF $count=1 $X=2.89
+ $Y=1.84 $X2=3.05 $Y2=2.715
r35 2 15 400 $w=1.7e-07 $l=2.63106e-07 $layer=licon1_PDIFF $count=1 $X=2.89
+ $Y=1.84 $X2=3.05 $Y2=2.035
r36 1 9 300 $w=1.7e-07 $l=6.05372e-07 $layer=licon1_PDIFF $count=2 $X=1.94
+ $Y=1.84 $X2=2.09 $Y2=2.375
.ends

.subckt PM_SKY130_FD_SC_HS__A22O_2%VGND 1 2 3 10 12 16 20 23 24 25 27 40 41 47
r46 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r47 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r48 40 41 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r49 38 41 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.6
+ $Y2=0
r50 37 38 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r51 35 48 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r52 34 37 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.68 $Y=0 $X2=2.64
+ $Y2=0
r53 34 35 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r54 32 47 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.29 $Y=0 $X2=1.165
+ $Y2=0
r55 32 34 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=1.29 $Y=0 $X2=1.68
+ $Y2=0
r56 31 48 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r57 31 45 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r58 30 31 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r59 28 44 4.03243 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=0.35 $Y=0 $X2=0.175
+ $Y2=0
r60 28 30 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.35 $Y=0 $X2=0.72
+ $Y2=0
r61 27 47 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.04 $Y=0 $X2=1.165
+ $Y2=0
r62 27 30 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=1.04 $Y=0 $X2=0.72
+ $Y2=0
r63 25 38 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=2.64
+ $Y2=0
r64 25 35 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=1.68
+ $Y2=0
r65 23 37 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=2.87 $Y=0 $X2=2.64
+ $Y2=0
r66 23 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.87 $Y=0 $X2=3.035
+ $Y2=0
r67 22 40 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=3.2 $Y=0 $X2=3.6 $Y2=0
r68 22 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.2 $Y=0 $X2=3.035
+ $Y2=0
r69 18 24 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.035 $Y=0.085
+ $X2=3.035 $Y2=0
r70 18 20 20.6043 $w=3.28e-07 $l=5.9e-07 $layer=LI1_cond $X=3.035 $Y=0.085
+ $X2=3.035 $Y2=0.675
r71 14 47 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.165 $Y=0.085
+ $X2=1.165 $Y2=0
r72 14 16 27.1977 $w=2.48e-07 $l=5.9e-07 $layer=LI1_cond $X=1.165 $Y=0.085
+ $X2=1.165 $Y2=0.675
r73 10 44 3.11073 $w=2.5e-07 $l=1.07121e-07 $layer=LI1_cond $X=0.225 $Y=0.085
+ $X2=0.175 $Y2=0
r74 10 12 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=0.225 $Y=0.085
+ $X2=0.225 $Y2=0.515
r75 3 20 182 $w=1.7e-07 $l=3.8461e-07 $layer=licon1_NDIFF $count=1 $X=2.855
+ $Y=0.37 $X2=3.035 $Y2=0.675
r76 2 16 182 $w=1.7e-07 $l=3.68409e-07 $layer=licon1_NDIFF $count=1 $X=0.985
+ $Y=0.37 $X2=1.125 $Y2=0.675
r77 1 12 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.14
+ $Y=0.37 $X2=0.265 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__A22O_2%A_304_74# 1 2 9 11 12 14 15 16 19
c40 16 0 7.19554e-20 $X=2.67 $Y=1.095
c41 11 0 3.95755e-20 $X=2.5 $Y=0.34
r42 17 19 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=3.535 $Y=1.01
+ $X2=3.535 $Y2=0.515
r43 15 17 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.37 $Y=1.095
+ $X2=3.535 $Y2=1.01
r44 15 16 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=3.37 $Y=1.095 $X2=2.67
+ $Y2=1.095
r45 14 16 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.585 $Y=1.01
+ $X2=2.67 $Y2=1.095
r46 13 14 38.1658 $w=1.68e-07 $l=5.85e-07 $layer=LI1_cond $X=2.585 $Y=0.425
+ $X2=2.585 $Y2=1.01
r47 11 13 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.5 $Y=0.34
+ $X2=2.585 $Y2=0.425
r48 11 12 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.5 $Y=0.34 $X2=1.83
+ $Y2=0.34
r49 7 12 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.665 $Y=0.425
+ $X2=1.83 $Y2=0.34
r50 7 9 8.73063 $w=3.28e-07 $l=2.5e-07 $layer=LI1_cond $X=1.665 $Y=0.425
+ $X2=1.665 $Y2=0.675
r51 2 19 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.395
+ $Y=0.37 $X2=3.535 $Y2=0.515
r52 1 9 182 $w=1.7e-07 $l=3.70473e-07 $layer=licon1_NDIFF $count=1 $X=1.52
+ $Y=0.37 $X2=1.665 $Y2=0.675
.ends

