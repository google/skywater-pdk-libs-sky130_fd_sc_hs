* File: sky130_fd_sc_hs__nor2b_4.pex.spice
* Created: Tue Sep  1 20:11:20 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HS__NOR2B_4%A 2 3 5 7 8 10 12 13 15 16 18 19 21 22 24 25
+ 26 29 30 32 33 39
c112 19 0 6.85393e-20 $X=3.705 $Y=1.765
r113 39 41 16.3138 $w=3.25e-07 $l=1.1e-07 $layer=POLY_cond $X=1.295 $Y=1.175
+ $X2=1.405 $Y2=1.175
r114 39 40 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.295
+ $Y=1.175 $X2=1.295 $Y2=1.175
r115 37 39 50.4246 $w=3.25e-07 $l=3.4e-07 $layer=POLY_cond $X=0.955 $Y=1.175
+ $X2=1.295 $Y2=1.175
r116 36 37 66.7385 $w=3.25e-07 $l=4.5e-07 $layer=POLY_cond $X=0.505 $Y=1.175
+ $X2=0.955 $Y2=1.175
r117 33 40 12.3931 $w=3.79e-07 $l=3.85e-07 $layer=LI1_cond $X=1.68 $Y=1.21
+ $X2=1.295 $Y2=1.21
r118 32 40 3.05805 $w=3.79e-07 $l=9.5e-08 $layer=LI1_cond $X=1.2 $Y=1.21
+ $X2=1.295 $Y2=1.21
r119 30 45 18.4294 $w=3.4e-07 $l=1.3e-07 $layer=POLY_cond $X=3.81 $Y=1.492
+ $X2=3.94 $Y2=1.492
r120 30 43 14.8853 $w=3.4e-07 $l=1.05e-07 $layer=POLY_cond $X=3.81 $Y=1.492
+ $X2=3.705 $Y2=1.492
r121 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.81
+ $Y=1.385 $X2=3.81 $Y2=1.385
r122 27 29 7.15912 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=3.81 $Y=1.18
+ $X2=3.81 $Y2=1.385
r123 26 33 7.46052 $w=3.79e-07 $l=1.62635e-07 $layer=LI1_cond $X=1.795 $Y=1.095
+ $X2=1.68 $Y2=1.21
r124 25 27 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.645 $Y=1.095
+ $X2=3.81 $Y2=1.18
r125 25 26 120.695 $w=1.68e-07 $l=1.85e-06 $layer=LI1_cond $X=3.645 $Y=1.095
+ $X2=1.795 $Y2=1.095
r126 22 45 21.9347 $w=1.5e-07 $l=2.72e-07 $layer=POLY_cond $X=3.94 $Y=1.22
+ $X2=3.94 $Y2=1.492
r127 22 24 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=3.94 $Y=1.22
+ $X2=3.94 $Y2=0.74
r128 19 43 21.9347 $w=1.5e-07 $l=2.73e-07 $layer=POLY_cond $X=3.705 $Y=1.765
+ $X2=3.705 $Y2=1.492
r129 19 21 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.705 $Y=1.765
+ $X2=3.705 $Y2=2.4
r130 16 43 27.6441 $w=3.4e-07 $l=3.56404e-07 $layer=POLY_cond $X=3.51 $Y=1.22
+ $X2=3.705 $Y2=1.492
r131 16 18 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=3.51 $Y=1.22
+ $X2=3.51 $Y2=0.74
r132 13 15 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.405 $Y=1.765
+ $X2=1.405 $Y2=2.4
r133 12 13 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=1.405 $Y=1.675
+ $X2=1.405 $Y2=1.765
r134 11 41 16.5763 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.405 $Y=1.34
+ $X2=1.405 $Y2=1.175
r135 11 12 130.218 $w=1.8e-07 $l=3.35e-07 $layer=POLY_cond $X=1.405 $Y=1.34
+ $X2=1.405 $Y2=1.675
r136 8 10 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.955 $Y=1.765
+ $X2=0.955 $Y2=2.4
r137 7 8 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=0.955 $Y=1.675
+ $X2=0.955 $Y2=1.765
r138 6 37 16.5763 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=0.955 $Y=1.34
+ $X2=0.955 $Y2=1.175
r139 6 7 130.218 $w=1.8e-07 $l=3.35e-07 $layer=POLY_cond $X=0.955 $Y=1.34
+ $X2=0.955 $Y2=1.675
r140 3 5 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.505 $Y=1.765
+ $X2=0.505 $Y2=2.4
r141 2 3 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=0.505 $Y=1.675
+ $X2=0.505 $Y2=1.765
r142 1 36 16.5763 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=0.505 $Y=1.34
+ $X2=0.505 $Y2=1.175
r143 1 2 130.218 $w=1.8e-07 $l=3.35e-07 $layer=POLY_cond $X=0.505 $Y=1.34
+ $X2=0.505 $Y2=1.675
.ends

.subckt PM_SKY130_FD_SC_HS__NOR2B_4%A_353_323# 1 2 7 9 10 12 13 15 16 18 19 21
+ 22 24 25 30 34 37 41 48
c105 25 0 6.85393e-20 $X=3.055 $Y=1.515
r106 54 55 31.7636 $w=4.78e-07 $l=3.15e-07 $layer=POLY_cond $X=2.44 $Y=1.495
+ $X2=2.755 $Y2=1.495
r107 51 52 29.7469 $w=4.78e-07 $l=2.95e-07 $layer=POLY_cond $X=2.01 $Y=1.495
+ $X2=2.305 $Y2=1.495
r108 45 48 9.083 $w=6.63e-07 $l=5.05e-07 $layer=LI1_cond $X=4.495 $Y=0.677 $X2=5
+ $Y2=0.677
r109 41 57 14.6213 $w=4.78e-07 $l=1.45e-07 $layer=POLY_cond $X=3.06 $Y=1.495
+ $X2=3.205 $Y2=1.495
r110 41 55 30.7552 $w=4.78e-07 $l=3.05e-07 $layer=POLY_cond $X=3.06 $Y=1.495
+ $X2=2.755 $Y2=1.495
r111 37 44 5.48801 $w=2.67e-07 $l=9.44722e-08 $layer=LI1_cond $X=4.495 $Y=1.72
+ $X2=4.515 $Y2=1.805
r112 36 45 8.98481 $w=1.7e-07 $l=3.33e-07 $layer=LI1_cond $X=4.495 $Y=1.01
+ $X2=4.495 $Y2=0.677
r113 36 37 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=4.495 $Y=1.01
+ $X2=4.495 $Y2=1.72
r114 34 44 13.6046 $w=3.3e-07 $l=3.55e-07 $layer=LI1_cond $X=4.515 $Y=2.16
+ $X2=4.515 $Y2=1.805
r115 31 42 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.225 $Y=1.805
+ $X2=3.14 $Y2=1.805
r116 30 44 3.37873 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.35 $Y=1.805
+ $X2=4.515 $Y2=1.805
r117 30 31 73.3957 $w=1.68e-07 $l=1.125e-06 $layer=LI1_cond $X=4.35 $Y=1.805
+ $X2=3.225 $Y2=1.805
r118 28 54 6.05021 $w=4.78e-07 $l=6e-08 $layer=POLY_cond $X=2.38 $Y=1.495
+ $X2=2.44 $Y2=1.495
r119 28 52 7.56276 $w=4.78e-07 $l=7.5e-08 $layer=POLY_cond $X=2.38 $Y=1.495
+ $X2=2.305 $Y2=1.495
r120 27 28 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=2.38
+ $Y=1.515 $X2=2.38 $Y2=1.515
r121 25 42 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=3.14 $Y=1.515
+ $X2=3.14 $Y2=1.805
r122 25 41 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=3.06
+ $Y=1.515 $X2=3.06 $Y2=1.515
r123 25 27 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=3.055 $Y=1.515
+ $X2=2.38 $Y2=1.515
r124 22 57 30.2749 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=3.205 $Y=1.765
+ $X2=3.205 $Y2=1.495
r125 22 24 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.205 $Y=1.765
+ $X2=3.205 $Y2=2.4
r126 19 55 30.2749 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=2.755 $Y=1.765
+ $X2=2.755 $Y2=1.495
r127 19 21 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.755 $Y=1.765
+ $X2=2.755 $Y2=2.4
r128 16 54 30.2749 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=2.44 $Y=1.225
+ $X2=2.44 $Y2=1.495
r129 16 18 155.847 $w=1.5e-07 $l=4.85e-07 $layer=POLY_cond $X=2.44 $Y=1.225
+ $X2=2.44 $Y2=0.74
r130 13 52 30.2749 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=2.305 $Y=1.765
+ $X2=2.305 $Y2=1.495
r131 13 15 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.305 $Y=1.765
+ $X2=2.305 $Y2=2.4
r132 10 51 30.2749 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=2.01 $Y=1.225
+ $X2=2.01 $Y2=1.495
r133 10 12 155.847 $w=1.5e-07 $l=4.85e-07 $layer=POLY_cond $X=2.01 $Y=1.225
+ $X2=2.01 $Y2=0.74
r134 7 51 15.6297 $w=4.78e-07 $l=3.38748e-07 $layer=POLY_cond $X=1.855 $Y=1.765
+ $X2=2.01 $Y2=1.495
r135 7 9 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.855 $Y=1.765
+ $X2=1.855 $Y2=2.4
r136 2 34 300 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=2 $X=4.365
+ $Y=2.015 $X2=4.515 $Y2=2.16
r137 1 48 45.5 $w=1.7e-07 $l=6.1883e-07 $layer=licon1_NDIFF $count=4 $X=4.445
+ $Y=0.37 $X2=5 $Y2=0.505
.ends

.subckt PM_SKY130_FD_SC_HS__NOR2B_4%B_N 1 3 6 8 10 11 12 17
r35 19 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.895
+ $Y=1.66 $X2=4.895 $Y2=1.66
r36 17 19 18.1335 $w=4.12e-07 $l=1.55e-07 $layer=POLY_cond $X=4.74 $Y=1.717
+ $X2=4.895 $Y2=1.717
r37 16 17 43.2864 $w=4.12e-07 $l=3.7e-07 $layer=POLY_cond $X=4.37 $Y=1.717
+ $X2=4.74 $Y2=1.717
r38 12 20 0.142277 $w=4.03e-07 $l=5e-09 $layer=LI1_cond $X=4.952 $Y=1.665
+ $X2=4.952 $Y2=1.66
r39 11 20 10.3862 $w=4.03e-07 $l=3.65e-07 $layer=LI1_cond $X=4.952 $Y=1.295
+ $X2=4.952 $Y2=1.66
r40 8 17 26.5862 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=4.74 $Y=1.94
+ $X2=4.74 $Y2=1.717
r41 8 10 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=4.74 $Y=1.94 $X2=4.74
+ $Y2=2.435
r42 4 16 26.5862 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=4.37 $Y=1.495
+ $X2=4.37 $Y2=1.717
r43 4 6 387.138 $w=1.5e-07 $l=7.55e-07 $layer=POLY_cond $X=4.37 $Y=1.495
+ $X2=4.37 $Y2=0.74
r44 1 16 9.35922 $w=4.12e-07 $l=2.5994e-07 $layer=POLY_cond $X=4.29 $Y=1.94
+ $X2=4.37 $Y2=1.717
r45 1 3 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=4.29 $Y=1.94 $X2=4.29
+ $Y2=2.435
.ends

.subckt PM_SKY130_FD_SC_HS__NOR2B_4%VPWR 1 2 3 4 13 15 21 25 29 31 34 35 36 38
+ 47 55 59
r67 58 59 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r68 55 56 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r69 52 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r70 50 59 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=5.04 $Y2=3.33
r71 49 50 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r72 47 58 3.96842 $w=1.7e-07 $l=2e-07 $layer=LI1_cond $X=4.88 $Y=3.33 $X2=5.08
+ $Y2=3.33
r73 47 49 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=4.88 $Y=3.33 $X2=4.56
+ $Y2=3.33
r74 46 50 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.56 $Y2=3.33
r75 45 46 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r76 43 55 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.265 $Y=3.33
+ $X2=1.18 $Y2=3.33
r77 43 45 152.337 $w=1.68e-07 $l=2.335e-06 $layer=LI1_cond $X=1.265 $Y=3.33
+ $X2=3.6 $Y2=3.33
r78 42 56 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r79 42 53 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r80 41 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r81 39 52 4.00981 $w=1.7e-07 $l=1.83e-07 $layer=LI1_cond $X=0.365 $Y=3.33
+ $X2=0.182 $Y2=3.33
r82 39 41 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=0.365 $Y=3.33
+ $X2=0.72 $Y2=3.33
r83 38 55 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.095 $Y=3.33
+ $X2=1.18 $Y2=3.33
r84 38 41 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=1.095 $Y=3.33
+ $X2=0.72 $Y2=3.33
r85 36 46 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.6 $Y2=3.33
r86 36 56 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=1.2 $Y2=3.33
r87 34 45 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=3.815 $Y=3.33
+ $X2=3.6 $Y2=3.33
r88 34 35 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.815 $Y=3.33
+ $X2=3.98 $Y2=3.33
r89 33 49 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=4.145 $Y=3.33
+ $X2=4.56 $Y2=3.33
r90 33 35 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.145 $Y=3.33
+ $X2=3.98 $Y2=3.33
r91 29 58 3.17474 $w=2.5e-07 $l=1.16619e-07 $layer=LI1_cond $X=5.005 $Y=3.245
+ $X2=5.08 $Y2=3.33
r92 29 31 50.016 $w=2.48e-07 $l=1.085e-06 $layer=LI1_cond $X=5.005 $Y=3.245
+ $X2=5.005 $Y2=2.16
r93 25 28 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=3.98 $Y=2.145
+ $X2=3.98 $Y2=2.825
r94 23 35 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.98 $Y=3.245
+ $X2=3.98 $Y2=3.33
r95 23 28 14.6675 $w=3.28e-07 $l=4.2e-07 $layer=LI1_cond $X=3.98 $Y=3.245
+ $X2=3.98 $Y2=2.825
r96 19 55 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.18 $Y=3.245
+ $X2=1.18 $Y2=3.33
r97 19 21 53.4973 $w=1.68e-07 $l=8.2e-07 $layer=LI1_cond $X=1.18 $Y=3.245
+ $X2=1.18 $Y2=2.425
r98 15 18 36.8782 $w=2.48e-07 $l=8e-07 $layer=LI1_cond $X=0.24 $Y=2.015 $X2=0.24
+ $Y2=2.815
r99 13 52 3.13335 $w=2.5e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.24 $Y=3.245
+ $X2=0.182 $Y2=3.33
r100 13 18 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=0.24 $Y=3.245
+ $X2=0.24 $Y2=2.815
r101 4 31 300 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=2 $X=4.815
+ $Y=2.015 $X2=4.965 $Y2=2.16
r102 3 28 600 $w=1.7e-07 $l=1.08038e-06 $layer=licon1_PDIFF $count=1 $X=3.78
+ $Y=1.84 $X2=3.98 $Y2=2.825
r103 3 25 300 $w=1.7e-07 $l=3.9246e-07 $layer=licon1_PDIFF $count=2 $X=3.78
+ $Y=1.84 $X2=3.98 $Y2=2.145
r104 2 21 300 $w=1.7e-07 $l=6.55725e-07 $layer=licon1_PDIFF $count=2 $X=1.03
+ $Y=1.84 $X2=1.18 $Y2=2.425
r105 1 18 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.815
r106 1 15 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.015
.ends

.subckt PM_SKY130_FD_SC_HS__NOR2B_4%A_116_368# 1 2 3 4 13 15 17 19 22 23 24 27
+ 29 33 41
r64 33 36 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=3.48 $Y=2.145
+ $X2=3.48 $Y2=2.825
r65 31 36 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=3.48 $Y=2.905 $X2=3.48
+ $Y2=2.825
r66 30 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.695 $Y=2.99
+ $X2=2.53 $Y2=2.99
r67 29 31 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.315 $Y=2.99
+ $X2=3.48 $Y2=2.905
r68 29 30 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=3.315 $Y=2.99
+ $X2=2.695 $Y2=2.99
r69 25 41 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.53 $Y=2.905
+ $X2=2.53 $Y2=2.99
r70 25 27 14.6675 $w=3.28e-07 $l=4.2e-07 $layer=LI1_cond $X=2.53 $Y=2.905
+ $X2=2.53 $Y2=2.485
r71 23 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.365 $Y=2.99
+ $X2=2.53 $Y2=2.99
r72 23 24 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=2.365 $Y=2.99
+ $X2=1.715 $Y2=2.99
r73 20 24 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.59 $Y=2.905
+ $X2=1.715 $Y2=2.99
r74 20 22 4.14879 $w=2.48e-07 $l=9e-08 $layer=LI1_cond $X=1.59 $Y=2.905 $X2=1.59
+ $Y2=2.815
r75 19 40 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.59 $Y=2.09 $X2=1.59
+ $Y2=2.005
r76 19 22 33.4208 $w=2.48e-07 $l=7.25e-07 $layer=LI1_cond $X=1.59 $Y=2.09
+ $X2=1.59 $Y2=2.815
r77 18 38 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.895 $Y=2.005
+ $X2=0.73 $Y2=2.005
r78 17 40 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.465 $Y=2.005
+ $X2=1.59 $Y2=2.005
r79 17 18 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=1.465 $Y=2.005
+ $X2=0.895 $Y2=2.005
r80 13 38 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.73 $Y=2.09 $X2=0.73
+ $Y2=2.005
r81 13 15 25.3188 $w=3.28e-07 $l=7.25e-07 $layer=LI1_cond $X=0.73 $Y=2.09
+ $X2=0.73 $Y2=2.815
r82 4 36 400 $w=1.7e-07 $l=1.08038e-06 $layer=licon1_PDIFF $count=1 $X=3.28
+ $Y=1.84 $X2=3.48 $Y2=2.825
r83 4 33 400 $w=1.7e-07 $l=3.9246e-07 $layer=licon1_PDIFF $count=1 $X=3.28
+ $Y=1.84 $X2=3.48 $Y2=2.145
r84 3 27 300 $w=1.7e-07 $l=7.16083e-07 $layer=licon1_PDIFF $count=2 $X=2.38
+ $Y=1.84 $X2=2.53 $Y2=2.485
r85 2 40 400 $w=1.7e-07 $l=3.11087e-07 $layer=licon1_PDIFF $count=1 $X=1.48
+ $Y=1.84 $X2=1.63 $Y2=2.085
r86 2 22 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=1.48
+ $Y=1.84 $X2=1.63 $Y2=2.815
r87 1 38 400 $w=1.7e-07 $l=3.11087e-07 $layer=licon1_PDIFF $count=1 $X=0.58
+ $Y=1.84 $X2=0.73 $Y2=2.085
r88 1 15 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=0.58
+ $Y=1.84 $X2=0.73 $Y2=2.815
.ends

.subckt PM_SKY130_FD_SC_HS__NOR2B_4%Y 1 2 3 4 14 17 19 21 23 25 27 29 31 32 39
+ 40 44 48 49 60
r96 49 64 16.8321 $w=1.87e-07 $l=2.58e-07 $layer=LI1_cond $X=0.24 $Y=1.337
+ $X2=0.24 $Y2=1.595
r97 49 60 2.74011 $w=1.87e-07 $l=4.2e-08 $layer=LI1_cond $X=0.24 $Y=1.337
+ $X2=0.24 $Y2=1.295
r98 49 60 2.15457 $w=2.28e-07 $l=4.3e-08 $layer=LI1_cond $X=0.24 $Y=1.252
+ $X2=0.24 $Y2=1.295
r99 48 49 16.3847 $w=2.28e-07 $l=3.27e-07 $layer=LI1_cond $X=0.24 $Y=0.925
+ $X2=0.24 $Y2=1.252
r100 44 46 3.68782 $w=2.48e-07 $l=8e-08 $layer=LI1_cond $X=3.685 $Y=0.675
+ $X2=3.685 $Y2=0.755
r101 38 40 8.46729 $w=3.08e-07 $l=1.65e-07 $layer=LI1_cond $X=2.225 $Y=0.685
+ $X2=2.39 $Y2=0.685
r102 38 39 8.46729 $w=3.08e-07 $l=1.65e-07 $layer=LI1_cond $X=2.225 $Y=0.685
+ $X2=2.06 $Y2=0.685
r103 35 36 6.77778 $w=2.34e-07 $l=1.3e-07 $layer=LI1_cond $X=2.025 $Y=2.015
+ $X2=2.025 $Y2=2.145
r104 33 35 18.2479 $w=2.34e-07 $l=3.5e-07 $layer=LI1_cond $X=2.025 $Y=1.665
+ $X2=2.025 $Y2=2.015
r105 31 32 8.16314 $w=2.38e-07 $l=1.7e-07 $layer=LI1_cond $X=0.535 $Y=1.63
+ $X2=0.705 $Y2=1.63
r106 27 42 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.02 $Y=2.23
+ $X2=3.02 $Y2=2.145
r107 27 29 15.6732 $w=2.48e-07 $l=3.4e-07 $layer=LI1_cond $X=3.02 $Y=2.23
+ $X2=3.02 $Y2=2.57
r108 25 46 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.56 $Y=0.755
+ $X2=3.685 $Y2=0.755
r109 25 40 76.3316 $w=1.68e-07 $l=1.17e-06 $layer=LI1_cond $X=3.56 $Y=0.755
+ $X2=2.39 $Y2=0.755
r110 24 36 2.60974 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=2.165 $Y=2.145
+ $X2=2.025 $Y2=2.145
r111 23 42 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.895 $Y=2.145
+ $X2=3.02 $Y2=2.145
r112 23 24 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=2.895 $Y=2.145
+ $X2=2.165 $Y2=2.145
r113 19 36 4.06873 $w=2.8e-07 $l=8.5e-08 $layer=LI1_cond $X=2.025 $Y=2.23
+ $X2=2.025 $Y2=2.145
r114 19 21 13.994 $w=2.78e-07 $l=3.4e-07 $layer=LI1_cond $X=2.025 $Y=2.23
+ $X2=2.025 $Y2=2.57
r115 17 33 2.60974 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=1.885 $Y=1.665
+ $X2=2.025 $Y2=1.665
r116 17 32 76.984 $w=1.68e-07 $l=1.18e-06 $layer=LI1_cond $X=1.885 $Y=1.665
+ $X2=0.705 $Y2=1.665
r117 16 64 1.29116 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=0.355 $Y=1.595
+ $X2=0.24 $Y2=1.595
r118 16 31 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=0.355 $Y=1.595
+ $X2=0.535 $Y2=1.595
r119 14 48 8.37092 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=0.355 $Y=0.755
+ $X2=0.24 $Y2=0.84
r120 14 39 111.235 $w=1.68e-07 $l=1.705e-06 $layer=LI1_cond $X=0.355 $Y=0.755
+ $X2=2.06 $Y2=0.755
r121 4 42 600 $w=1.7e-07 $l=3.72525e-07 $layer=licon1_PDIFF $count=1 $X=2.83
+ $Y=1.84 $X2=2.98 $Y2=2.145
r122 4 29 600 $w=1.7e-07 $l=8.01499e-07 $layer=licon1_PDIFF $count=1 $X=2.83
+ $Y=1.84 $X2=2.98 $Y2=2.57
r123 3 35 600 $w=1.7e-07 $l=2.38485e-07 $layer=licon1_PDIFF $count=1 $X=1.93
+ $Y=1.84 $X2=2.08 $Y2=2.015
r124 3 21 600 $w=1.7e-07 $l=8.01499e-07 $layer=licon1_PDIFF $count=1 $X=1.93
+ $Y=1.84 $X2=2.08 $Y2=2.57
r125 2 44 182 $w=1.7e-07 $l=3.68409e-07 $layer=licon1_NDIFF $count=1 $X=3.585
+ $Y=0.37 $X2=3.725 $Y2=0.675
r126 1 38 182 $w=1.7e-07 $l=3.68409e-07 $layer=licon1_NDIFF $count=1 $X=2.085
+ $Y=0.37 $X2=2.225 $Y2=0.675
.ends

.subckt PM_SKY130_FD_SC_HS__NOR2B_4%VGND 1 2 3 12 18 20 22 30 37 38 41 46 52 54
r48 54 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r49 51 52 10.0584 $w=5.83e-07 $l=1.65e-07 $layer=LI1_cond $X=3.215 $Y=0.207
+ $X2=3.38 $Y2=0.207
r50 48 51 1.94235 $w=5.83e-07 $l=9.5e-08 $layer=LI1_cond $X=3.12 $Y=0.207
+ $X2=3.215 $Y2=0.207
r51 48 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r52 44 48 9.81398 $w=5.83e-07 $l=4.8e-07 $layer=LI1_cond $X=2.64 $Y=0.207
+ $X2=3.12 $Y2=0.207
r53 44 46 8.11604 $w=5.83e-07 $l=7e-08 $layer=LI1_cond $X=2.64 $Y=0.207 $X2=2.57
+ $Y2=0.207
r54 41 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r55 38 55 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=4.08
+ $Y2=0
r56 37 38 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r57 35 54 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.24 $Y=0 $X2=4.115
+ $Y2=0
r58 35 37 52.1925 $w=1.68e-07 $l=8e-07 $layer=LI1_cond $X=4.24 $Y=0 $X2=5.04
+ $Y2=0
r59 34 55 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.08
+ $Y2=0
r60 34 49 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=3.12
+ $Y2=0
r61 33 52 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=3.6 $Y=0 $X2=3.38
+ $Y2=0
r62 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r63 30 54 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.99 $Y=0 $X2=4.115
+ $Y2=0
r64 30 33 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=3.99 $Y=0 $X2=3.6
+ $Y2=0
r65 29 42 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=1.68
+ $Y2=0
r66 28 29 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r67 25 29 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=1.2
+ $Y2=0
r68 24 28 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.24 $Y=0 $X2=1.2
+ $Y2=0
r69 24 25 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r70 22 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.55 $Y=0 $X2=1.715
+ $Y2=0
r71 22 28 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=1.55 $Y=0 $X2=1.2
+ $Y2=0
r72 20 49 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r73 20 42 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=1.68
+ $Y2=0
r74 20 44 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r75 16 54 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.115 $Y=0.085
+ $X2=4.115 $Y2=0
r76 16 18 27.1977 $w=2.48e-07 $l=5.9e-07 $layer=LI1_cond $X=4.115 $Y=0.085
+ $X2=4.115 $Y2=0.675
r77 15 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.88 $Y=0 $X2=1.715
+ $Y2=0
r78 15 46 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.88 $Y=0 $X2=2.57
+ $Y2=0
r79 10 41 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.715 $Y=0.085
+ $X2=1.715 $Y2=0
r80 10 12 8.73063 $w=3.28e-07 $l=2.5e-07 $layer=LI1_cond $X=1.715 $Y=0.085
+ $X2=1.715 $Y2=0.335
r81 3 18 182 $w=1.7e-07 $l=3.68409e-07 $layer=licon1_NDIFF $count=1 $X=4.015
+ $Y=0.37 $X2=4.155 $Y2=0.675
r82 2 51 91 $w=1.7e-07 $l=7.17287e-07 $layer=licon1_NDIFF $count=2 $X=2.515
+ $Y=0.37 $X2=3.215 $Y2=0.335
r83 1 12 182 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=1 $X=1.57
+ $Y=0.19 $X2=1.715 $Y2=0.335
.ends

