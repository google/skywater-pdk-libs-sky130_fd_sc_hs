* File: sky130_fd_sc_hs__a2bb2o_2.spice
* Created: Thu Aug 27 20:27:45 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hs__a2bb2o_2.pex.spice"
.subckt sky130_fd_sc_hs__a2bb2o_2  VNB VPB B1 B2 A2_N A1_N VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A1_N	A1_N
* A2_N	A2_N
* B2	B2
* B1	B1
* VPB	VPB
* VNB	VNB
MM1008 A_149_74# N_B1_M1008_g N_VGND_M1008_s VNB NLOWVT L=0.15 W=0.74 AD=0.0777
+ AS=0.2109 PD=0.95 PS=2.05 NRD=8.1 NRS=0 M=1 R=4.93333 SA=75000.2 SB=75002.9
+ A=0.111 P=1.78 MULT=1
MM1001 N_A_221_74#_M1001_d N_B2_M1001_g A_149_74# VNB NLOWVT L=0.15 W=0.74
+ AD=0.1443 AS=0.0777 PD=1.13 PS=0.95 NRD=8.916 NRS=8.1 M=1 R=4.93333 SA=75000.6
+ SB=75002.5 A=0.111 P=1.78 MULT=1
MM1007 N_VGND_M1007_d N_A_293_333#_M1007_g N_A_221_74#_M1001_d VNB NLOWVT L=0.15
+ W=0.74 AD=0.295426 AS=0.1443 PD=1.82419 PS=1.13 NRD=4.86 NRS=8.916 M=1
+ R=4.93333 SA=75001.1 SB=75002 A=0.111 P=1.78 MULT=1
MM1006 N_A_293_333#_M1006_d N_A2_N_M1006_g N_VGND_M1007_d VNB NLOWVT L=0.15
+ W=0.55 AD=0.077 AS=0.219574 PD=0.83 PS=1.35581 NRD=0 NRS=0 M=1 R=3.66667
+ SA=75002.1 SB=75001.6 A=0.0825 P=1.4 MULT=1
MM1010 N_VGND_M1010_d N_A1_N_M1010_g N_A_293_333#_M1006_d VNB NLOWVT L=0.15
+ W=0.55 AD=0.111705 AS=0.077 PD=0.963566 PS=0.83 NRD=1.08 NRS=0 M=1 R=3.66667
+ SA=75002.5 SB=75001.2 A=0.0825 P=1.4 MULT=1
MM1000 N_X_M1000_d N_A_221_74#_M1000_g N_VGND_M1010_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.150295 PD=1.02 PS=1.29643 NRD=0 NRS=17.016 M=1 R=4.93333
+ SA=75002.3 SB=75000.6 A=0.111 P=1.78 MULT=1
MM1009 N_X_M1000_d N_A_221_74#_M1009_g N_VGND_M1009_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1961 PD=1.02 PS=2.01 NRD=0 NRS=0 M=1 R=4.93333 SA=75002.8
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1011 N_VPWR_M1011_d N_B1_M1011_g N_A_61_392#_M1011_s VPB PSHORT L=0.15 W=1
+ AD=0.15 AS=0.275 PD=1.3 PS=2.55 NRD=1.9503 NRS=1.9503 M=1 R=6.66667 SA=75000.2
+ SB=75001.1 A=0.15 P=2.3 MULT=1
MM1012 N_A_61_392#_M1012_d N_B2_M1012_g N_VPWR_M1011_d VPB PSHORT L=0.15 W=1
+ AD=0.15 AS=0.15 PD=1.3 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=6.66667 SA=75000.6
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1002 N_A_221_74#_M1002_d N_A_293_333#_M1002_g N_A_61_392#_M1012_d VPB PSHORT
+ L=0.15 W=1 AD=0.275 AS=0.15 PD=2.55 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=6.66667
+ SA=75001.1 SB=75000.2 A=0.15 P=2.3 MULT=1
MM1003 A_546_378# N_A2_N_M1003_g N_A_293_333#_M1003_s VPB PSHORT L=0.15 W=1
+ AD=0.12 AS=0.275 PD=1.24 PS=2.55 NRD=12.7853 NRS=1.9503 M=1 R=6.66667
+ SA=75000.2 SB=75001.5 A=0.15 P=2.3 MULT=1
MM1013 N_VPWR_M1013_d N_A1_N_M1013_g A_546_378# VPB PSHORT L=0.15 W=1
+ AD=0.184811 AS=0.12 PD=1.39623 PS=1.24 NRD=7.8603 NRS=12.7853 M=1 R=6.66667
+ SA=75000.6 SB=75001.2 A=0.15 P=2.3 MULT=1
MM1004 N_X_M1004_d N_A_221_74#_M1004_g N_VPWR_M1013_d VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.206989 PD=1.42 PS=1.56377 NRD=1.7533 NRS=7.0329 M=1 R=7.46667
+ SA=75001 SB=75000.6 A=0.168 P=2.54 MULT=1
MM1005 N_X_M1004_d N_A_221_74#_M1005_g N_VPWR_M1005_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.308 PD=1.42 PS=2.79 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.5 SB=75000.2 A=0.168 P=2.54 MULT=1
DX14_noxref VNB VPB NWDIODE A=9.6348 P=14.08
c_519 A_546_378# 0 4.64943e-20 $X=2.73 $Y=1.89
*
.include "sky130_fd_sc_hs__a2bb2o_2.pxi.spice"
*
.ends
*
*
