* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hs__dfxtp_4 CLK D VGND VNB VPB VPWR Q
M1000 VGND a_1226_296# Q VNB nlowvt w=740000u l=150000u
+  ad=1.88282e+12p pd=1.54e+07u as=4.44e+11p ps=4.16e+06u
M1001 Q a_1226_296# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1002 VPWR a_696_458# a_651_503# VPB pshort w=420000u l=150000u
+  ad=2.4029e+12p pd=1.958e+07u as=1.008e+11p ps=1.32e+06u
M1003 a_696_458# a_544_485# VPWR VPB pshort w=840000u l=150000u
+  ad=4.452e+11p pd=2.74e+06u as=0p ps=0u
M1004 Q a_1226_296# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_696_458# a_544_485# VGND VNB nlowvt w=550000u l=150000u
+  ad=1.98e+11p pd=1.97e+06u as=0p ps=0u
M1006 VPWR a_1226_296# a_1141_508# VPB pshort w=420000u l=150000u
+  ad=0p pd=0u as=1.995e+11p ps=1.79e+06u
M1007 Q a_1226_296# VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=6.72e+11p pd=5.68e+06u as=0p ps=0u
M1008 VPWR a_1226_296# Q VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 Q a_1226_296# VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_437_503# D VPWR VPB pshort w=420000u l=150000u
+  ad=1.7745e+11p pd=1.79e+06u as=0p ps=0u
M1011 VPWR a_1226_296# Q VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VGND a_696_458# a_735_102# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=8.82e+10p ps=1.26e+06u
M1013 VGND a_1226_296# Q VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_206_368# a_27_74# VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=3.304e+11p pd=2.83e+06u as=0p ps=0u
M1015 VPWR CLK a_27_74# VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=3.304e+11p ps=2.83e+06u
M1016 VGND a_1226_296# a_1178_124# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.323e+11p ps=1.47e+06u
M1017 a_735_102# a_206_368# a_544_485# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.51375e+11p ps=1.66e+06u
M1018 a_437_503# D VGND VNB nlowvt w=420000u l=150000u
+  ad=1.176e+11p pd=1.4e+06u as=0p ps=0u
M1019 a_544_485# a_206_368# a_437_503# VPB pshort w=420000u l=150000u
+  ad=1.7745e+11p pd=1.79e+06u as=0p ps=0u
M1020 a_651_503# a_27_74# a_544_485# VPB pshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_1141_508# a_206_368# a_1034_424# VPB pshort w=420000u l=150000u
+  ad=0p pd=0u as=2.856e+11p ps=2.45e+06u
M1022 a_544_485# a_27_74# a_437_503# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_1034_424# a_206_368# a_696_458# VNB nlowvt w=550000u l=150000u
+  ad=2.152e+11p pd=1.97e+06u as=0p ps=0u
M1024 a_206_368# a_27_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.516e+11p pd=2.16e+06u as=0p ps=0u
M1025 a_1226_296# a_1034_424# VPWR VPB pshort w=840000u l=150000u
+  ad=2.52e+11p pd=2.28e+06u as=0p ps=0u
M1026 VGND a_1034_424# a_1226_296# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1027 VGND CLK a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1028 a_1034_424# a_27_74# a_696_458# VPB pshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1029 VPWR a_1034_424# a_1226_296# VPB pshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1030 a_1178_124# a_27_74# a_1034_424# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
