* File: sky130_fd_sc_hs__a221oi_4.pex.spice
* Created: Tue Sep  1 19:50:37 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HS__A221OI_4%C1 1 3 6 8 10 13 15 17 20 22 24 27 29 30 31
+ 46 47
r82 47 48 8.62916 $w=3.91e-07 $l=7e-08 $layer=POLY_cond $X=1.845 $Y=1.542
+ $X2=1.915 $Y2=1.542
r83 45 47 16.6419 $w=3.91e-07 $l=1.35e-07 $layer=POLY_cond $X=1.71 $Y=1.542
+ $X2=1.845 $Y2=1.542
r84 45 46 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.71
+ $Y=1.515 $X2=1.71 $Y2=1.515
r85 43 45 27.7366 $w=3.91e-07 $l=2.25e-07 $layer=POLY_cond $X=1.485 $Y=1.542
+ $X2=1.71 $Y2=1.542
r86 42 43 11.0946 $w=3.91e-07 $l=9e-08 $layer=POLY_cond $X=1.395 $Y=1.542
+ $X2=1.485 $Y2=1.542
r87 41 42 41.913 $w=3.91e-07 $l=3.4e-07 $layer=POLY_cond $X=1.055 $Y=1.542
+ $X2=1.395 $Y2=1.542
r88 40 41 13.5601 $w=3.91e-07 $l=1.1e-07 $layer=POLY_cond $X=0.945 $Y=1.542
+ $X2=1.055 $Y2=1.542
r89 38 40 31.4348 $w=3.91e-07 $l=2.55e-07 $layer=POLY_cond $X=0.69 $Y=1.542
+ $X2=0.945 $Y2=1.542
r90 38 39 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.69
+ $Y=1.515 $X2=0.69 $Y2=1.515
r91 36 38 8.01279 $w=3.91e-07 $l=6.5e-08 $layer=POLY_cond $X=0.625 $Y=1.542
+ $X2=0.69 $Y2=1.542
r92 35 36 16.0256 $w=3.91e-07 $l=1.3e-07 $layer=POLY_cond $X=0.495 $Y=1.542
+ $X2=0.625 $Y2=1.542
r93 31 46 0.80403 $w=4.28e-07 $l=3e-08 $layer=LI1_cond $X=1.68 $Y=1.565 $X2=1.71
+ $Y2=1.565
r94 30 31 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=1.2 $Y=1.565
+ $X2=1.68 $Y2=1.565
r95 29 30 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=0.72 $Y=1.565
+ $X2=1.2 $Y2=1.565
r96 29 39 0.80403 $w=4.28e-07 $l=3e-08 $layer=LI1_cond $X=0.72 $Y=1.565 $X2=0.69
+ $Y2=1.565
r97 25 48 25.3065 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=1.915 $Y=1.32
+ $X2=1.915 $Y2=1.542
r98 25 27 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=1.915 $Y=1.32
+ $X2=1.915 $Y2=0.74
r99 22 47 25.3065 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=1.845 $Y=1.765
+ $X2=1.845 $Y2=1.542
r100 22 24 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.845 $Y=1.765
+ $X2=1.845 $Y2=2.4
r101 18 43 25.3065 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=1.485 $Y=1.32
+ $X2=1.485 $Y2=1.542
r102 18 20 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=1.485 $Y=1.32
+ $X2=1.485 $Y2=0.74
r103 15 42 25.3065 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=1.395 $Y=1.765
+ $X2=1.395 $Y2=1.542
r104 15 17 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.395 $Y=1.765
+ $X2=1.395 $Y2=2.4
r105 11 41 25.3065 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=1.055 $Y=1.32
+ $X2=1.055 $Y2=1.542
r106 11 13 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=1.055 $Y=1.32
+ $X2=1.055 $Y2=0.74
r107 8 40 25.3065 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=0.945 $Y=1.765
+ $X2=0.945 $Y2=1.542
r108 8 10 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.945 $Y=1.765
+ $X2=0.945 $Y2=2.4
r109 4 36 25.3065 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=0.625 $Y=1.32
+ $X2=0.625 $Y2=1.542
r110 4 6 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=0.625 $Y=1.32
+ $X2=0.625 $Y2=0.74
r111 1 35 25.3065 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=0.495 $Y=1.765
+ $X2=0.495 $Y2=1.542
r112 1 3 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.495 $Y=1.765
+ $X2=0.495 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_HS__A221OI_4%A2 1 3 6 10 12 14 17 19 21 24 26 28 29 30
+ 31 32 33 53 54
r84 54 55 7.24317 $w=3.66e-07 $l=5.5e-08 $layer=POLY_cond $X=4.3 $Y=1.557
+ $X2=4.355 $Y2=1.557
r85 52 54 26.3388 $w=3.66e-07 $l=2e-07 $layer=POLY_cond $X=4.1 $Y=1.557 $X2=4.3
+ $Y2=1.557
r86 52 53 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.1
+ $Y=1.515 $X2=4.1 $Y2=1.515
r87 50 52 25.6803 $w=3.66e-07 $l=1.95e-07 $layer=POLY_cond $X=3.905 $Y=1.557
+ $X2=4.1 $Y2=1.557
r88 49 50 4.60929 $w=3.66e-07 $l=3.5e-08 $layer=POLY_cond $X=3.87 $Y=1.557
+ $X2=3.905 $Y2=1.557
r89 47 49 14.4863 $w=3.66e-07 $l=1.1e-07 $layer=POLY_cond $X=3.76 $Y=1.557
+ $X2=3.87 $Y2=1.557
r90 47 48 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.76
+ $Y=1.515 $X2=3.76 $Y2=1.515
r91 45 47 40.1667 $w=3.66e-07 $l=3.05e-07 $layer=POLY_cond $X=3.455 $Y=1.557
+ $X2=3.76 $Y2=1.557
r92 44 45 1.97541 $w=3.66e-07 $l=1.5e-08 $layer=POLY_cond $X=3.44 $Y=1.557
+ $X2=3.455 $Y2=1.557
r93 42 44 2.63388 $w=3.66e-07 $l=2e-08 $layer=POLY_cond $X=3.42 $Y=1.557
+ $X2=3.44 $Y2=1.557
r94 42 43 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.42
+ $Y=1.515 $X2=3.42 $Y2=1.515
r95 40 42 53.9945 $w=3.66e-07 $l=4.1e-07 $layer=POLY_cond $X=3.01 $Y=1.557
+ $X2=3.42 $Y2=1.557
r96 39 40 0.65847 $w=3.66e-07 $l=5e-09 $layer=POLY_cond $X=3.005 $Y=1.557
+ $X2=3.01 $Y2=1.557
r97 33 53 0.658539 $w=3.48e-07 $l=2e-08 $layer=LI1_cond $X=4.08 $Y=1.605 $X2=4.1
+ $Y2=1.605
r98 33 48 10.5366 $w=3.48e-07 $l=3.2e-07 $layer=LI1_cond $X=4.08 $Y=1.605
+ $X2=3.76 $Y2=1.605
r99 32 48 5.26831 $w=3.48e-07 $l=1.6e-07 $layer=LI1_cond $X=3.6 $Y=1.605
+ $X2=3.76 $Y2=1.605
r100 32 43 5.92685 $w=3.48e-07 $l=1.8e-07 $layer=LI1_cond $X=3.6 $Y=1.605
+ $X2=3.42 $Y2=1.605
r101 31 43 9.87808 $w=3.48e-07 $l=3e-07 $layer=LI1_cond $X=3.12 $Y=1.605
+ $X2=3.42 $Y2=1.605
r102 30 31 15.8049 $w=3.48e-07 $l=4.8e-07 $layer=LI1_cond $X=2.64 $Y=1.605
+ $X2=3.12 $Y2=1.605
r103 29 30 15.8049 $w=3.48e-07 $l=4.8e-07 $layer=LI1_cond $X=2.16 $Y=1.605
+ $X2=2.64 $Y2=1.605
r104 26 55 23.7042 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=4.355 $Y=1.765
+ $X2=4.355 $Y2=1.557
r105 26 28 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=4.355 $Y=1.765
+ $X2=4.355 $Y2=2.4
r106 22 54 23.7042 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.3 $Y=1.35
+ $X2=4.3 $Y2=1.557
r107 22 24 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=4.3 $Y=1.35 $X2=4.3
+ $Y2=0.74
r108 19 50 23.7042 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=3.905 $Y=1.765
+ $X2=3.905 $Y2=1.557
r109 19 21 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.905 $Y=1.765
+ $X2=3.905 $Y2=2.4
r110 15 49 23.7042 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.87 $Y=1.35
+ $X2=3.87 $Y2=1.557
r111 15 17 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=3.87 $Y=1.35
+ $X2=3.87 $Y2=0.74
r112 12 45 23.7042 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=3.455 $Y=1.765
+ $X2=3.455 $Y2=1.557
r113 12 14 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.455 $Y=1.765
+ $X2=3.455 $Y2=2.4
r114 8 44 23.7042 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.44 $Y=1.35
+ $X2=3.44 $Y2=1.557
r115 8 10 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=3.44 $Y=1.35
+ $X2=3.44 $Y2=0.74
r116 4 40 23.7042 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.01 $Y=1.35
+ $X2=3.01 $Y2=1.557
r117 4 6 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=3.01 $Y=1.35 $X2=3.01
+ $Y2=0.74
r118 1 39 23.7042 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=3.005 $Y=1.765
+ $X2=3.005 $Y2=1.557
r119 1 3 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.005 $Y=1.765
+ $X2=3.005 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_HS__A221OI_4%A1 3 5 7 10 12 14 17 19 21 24 26 28 29 30
+ 31 32 51
c98 32 0 1.32887e-19 $X=6 $Y=1.665
c99 19 0 1.00303e-20 $X=5.705 $Y=1.765
r100 51 52 43.8728 $w=4.01e-07 $l=3.65e-07 $layer=POLY_cond $X=6.02 $Y=1.542
+ $X2=6.385 $Y2=1.542
r101 49 51 8.41397 $w=4.01e-07 $l=7e-08 $layer=POLY_cond $X=5.95 $Y=1.542
+ $X2=6.02 $Y2=1.542
r102 49 50 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.95
+ $Y=1.515 $X2=5.95 $Y2=1.515
r103 47 49 29.4489 $w=4.01e-07 $l=2.45e-07 $layer=POLY_cond $X=5.705 $Y=1.542
+ $X2=5.95 $Y2=1.542
r104 46 47 13.8229 $w=4.01e-07 $l=1.15e-07 $layer=POLY_cond $X=5.59 $Y=1.542
+ $X2=5.705 $Y2=1.542
r105 44 46 10.818 $w=4.01e-07 $l=9e-08 $layer=POLY_cond $X=5.5 $Y=1.542 $X2=5.59
+ $Y2=1.542
r106 44 45 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.5
+ $Y=1.515 $X2=5.5 $Y2=1.515
r107 42 44 29.4489 $w=4.01e-07 $l=2.45e-07 $layer=POLY_cond $X=5.255 $Y=1.542
+ $X2=5.5 $Y2=1.542
r108 41 45 11.1952 $w=3.48e-07 $l=3.4e-07 $layer=LI1_cond $X=5.16 $Y=1.605
+ $X2=5.5 $Y2=1.605
r109 40 42 11.419 $w=4.01e-07 $l=9.5e-08 $layer=POLY_cond $X=5.16 $Y=1.542
+ $X2=5.255 $Y2=1.542
r110 40 41 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.16
+ $Y=1.515 $X2=5.16 $Y2=1.515
r111 38 40 42.6708 $w=4.01e-07 $l=3.55e-07 $layer=POLY_cond $X=4.805 $Y=1.542
+ $X2=5.16 $Y2=1.542
r112 37 38 9.01496 $w=4.01e-07 $l=7.5e-08 $layer=POLY_cond $X=4.73 $Y=1.542
+ $X2=4.805 $Y2=1.542
r113 32 50 1.64635 $w=3.48e-07 $l=5e-08 $layer=LI1_cond $X=6 $Y=1.605 $X2=5.95
+ $Y2=1.605
r114 31 50 14.1586 $w=3.48e-07 $l=4.3e-07 $layer=LI1_cond $X=5.52 $Y=1.605
+ $X2=5.95 $Y2=1.605
r115 31 45 0.658539 $w=3.48e-07 $l=2e-08 $layer=LI1_cond $X=5.52 $Y=1.605
+ $X2=5.5 $Y2=1.605
r116 30 41 3.95123 $w=3.48e-07 $l=1.2e-07 $layer=LI1_cond $X=5.04 $Y=1.605
+ $X2=5.16 $Y2=1.605
r117 29 30 15.8049 $w=3.48e-07 $l=4.8e-07 $layer=LI1_cond $X=4.56 $Y=1.605
+ $X2=5.04 $Y2=1.605
r118 26 52 25.923 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=6.385 $Y=1.765
+ $X2=6.385 $Y2=1.542
r119 26 28 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=6.385 $Y=1.765
+ $X2=6.385 $Y2=2.4
r120 22 51 25.923 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=6.02 $Y=1.32
+ $X2=6.02 $Y2=1.542
r121 22 24 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=6.02 $Y=1.32
+ $X2=6.02 $Y2=0.74
r122 19 47 25.923 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=5.705 $Y=1.765
+ $X2=5.705 $Y2=1.542
r123 19 21 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=5.705 $Y=1.765
+ $X2=5.705 $Y2=2.4
r124 15 46 25.923 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=5.59 $Y=1.32
+ $X2=5.59 $Y2=1.542
r125 15 17 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=5.59 $Y=1.32
+ $X2=5.59 $Y2=0.74
r126 12 42 25.923 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=5.255 $Y=1.765
+ $X2=5.255 $Y2=1.542
r127 12 14 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=5.255 $Y=1.765
+ $X2=5.255 $Y2=2.4
r128 8 40 25.923 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=5.16 $Y=1.32
+ $X2=5.16 $Y2=1.542
r129 8 10 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=5.16 $Y=1.32
+ $X2=5.16 $Y2=0.74
r130 5 38 25.923 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=4.805 $Y=1.765
+ $X2=4.805 $Y2=1.542
r131 5 7 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=4.805 $Y=1.765
+ $X2=4.805 $Y2=2.4
r132 1 37 25.923 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=4.73 $Y=1.32
+ $X2=4.73 $Y2=1.542
r133 1 3 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=4.73 $Y=1.32 $X2=4.73
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HS__A221OI_4%B1 1 3 6 8 10 13 15 17 20 22 24 27 29 30 31
+ 32 49 50 56 58 67
c88 67 0 1.00303e-20 $X=6.73 $Y=1.565
c89 50 0 2.78543e-19 $X=8.185 $Y=1.557
c90 22 0 1.25478e-19 $X=8.185 $Y=1.765
r91 56 58 0.402015 $w=4.28e-07 $l=1.5e-08 $layer=LI1_cond $X=6.945 $Y=1.565
+ $X2=6.96 $Y2=1.565
r92 50 51 10.0139 $w=3.61e-07 $l=7.5e-08 $layer=POLY_cond $X=8.185 $Y=1.557
+ $X2=8.26 $Y2=1.557
r93 48 50 34.0471 $w=3.61e-07 $l=2.55e-07 $layer=POLY_cond $X=7.93 $Y=1.557
+ $X2=8.185 $Y2=1.557
r94 48 49 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=7.93
+ $Y=1.515 $X2=7.93 $Y2=1.515
r95 46 48 13.3518 $w=3.61e-07 $l=1e-07 $layer=POLY_cond $X=7.83 $Y=1.557
+ $X2=7.93 $Y2=1.557
r96 45 46 12.6842 $w=3.61e-07 $l=9.5e-08 $layer=POLY_cond $X=7.735 $Y=1.557
+ $X2=7.83 $Y2=1.557
r97 44 45 44.7285 $w=3.61e-07 $l=3.35e-07 $layer=POLY_cond $X=7.4 $Y=1.557
+ $X2=7.735 $Y2=1.557
r98 43 44 15.3546 $w=3.61e-07 $l=1.15e-07 $layer=POLY_cond $X=7.285 $Y=1.557
+ $X2=7.4 $Y2=1.557
r99 42 43 42.0582 $w=3.61e-07 $l=3.15e-07 $layer=POLY_cond $X=6.97 $Y=1.557
+ $X2=7.285 $Y2=1.557
r100 40 42 8.01108 $w=3.61e-07 $l=6e-08 $layer=POLY_cond $X=6.91 $Y=1.557
+ $X2=6.97 $Y2=1.557
r101 38 40 10.0139 $w=3.61e-07 $l=7.5e-08 $layer=POLY_cond $X=6.835 $Y=1.557
+ $X2=6.91 $Y2=1.557
r102 32 49 0.26801 $w=4.28e-07 $l=1e-08 $layer=LI1_cond $X=7.92 $Y=1.565
+ $X2=7.93 $Y2=1.565
r103 31 32 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=7.44 $Y=1.565
+ $X2=7.92 $Y2=1.565
r104 30 56 0.938035 $w=4.28e-07 $l=3.5e-08 $layer=LI1_cond $X=6.91 $Y=1.565
+ $X2=6.945 $Y2=1.565
r105 30 67 5.25701 $w=4.28e-07 $l=1.8e-07 $layer=LI1_cond $X=6.91 $Y=1.565
+ $X2=6.73 $Y2=1.565
r106 30 31 11.9264 $w=4.28e-07 $l=4.45e-07 $layer=LI1_cond $X=6.995 $Y=1.565
+ $X2=7.44 $Y2=1.565
r107 30 58 0.938035 $w=4.28e-07 $l=3.5e-08 $layer=LI1_cond $X=6.995 $Y=1.565
+ $X2=6.96 $Y2=1.565
r108 30 40 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.91
+ $Y=1.515 $X2=6.91 $Y2=1.515
r109 29 67 8.23174 $w=3.48e-07 $l=2.5e-07 $layer=LI1_cond $X=6.48 $Y=1.605
+ $X2=6.73 $Y2=1.605
r110 25 51 23.3725 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=8.26 $Y=1.35
+ $X2=8.26 $Y2=1.557
r111 25 27 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=8.26 $Y=1.35
+ $X2=8.26 $Y2=0.74
r112 22 50 23.3725 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=8.185 $Y=1.765
+ $X2=8.185 $Y2=1.557
r113 22 24 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=8.185 $Y=1.765
+ $X2=8.185 $Y2=2.4
r114 18 46 23.3725 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=7.83 $Y=1.35
+ $X2=7.83 $Y2=1.557
r115 18 20 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=7.83 $Y=1.35
+ $X2=7.83 $Y2=0.74
r116 15 45 23.3725 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=7.735 $Y=1.765
+ $X2=7.735 $Y2=1.557
r117 15 17 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=7.735 $Y=1.765
+ $X2=7.735 $Y2=2.4
r118 11 44 23.3725 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=7.4 $Y=1.35
+ $X2=7.4 $Y2=1.557
r119 11 13 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=7.4 $Y=1.35 $X2=7.4
+ $Y2=0.74
r120 8 43 23.3725 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=7.285 $Y=1.765
+ $X2=7.285 $Y2=1.557
r121 8 10 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=7.285 $Y=1.765
+ $X2=7.285 $Y2=2.4
r122 4 42 23.3725 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=6.97 $Y=1.35
+ $X2=6.97 $Y2=1.557
r123 4 6 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=6.97 $Y=1.35 $X2=6.97
+ $Y2=0.74
r124 1 38 23.3725 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=6.835 $Y=1.765
+ $X2=6.835 $Y2=1.557
r125 1 3 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=6.835 $Y=1.765
+ $X2=6.835 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_HS__A221OI_4%B2 1 3 6 8 10 13 15 17 20 24 26 28 29 30 31
+ 32 49
c77 32 0 1.25478e-19 $X=9.84 $Y=1.665
c78 6 0 2.41835e-19 $X=8.69 $Y=0.74
r79 49 50 0.654891 $w=3.68e-07 $l=5e-09 $layer=POLY_cond $X=9.98 $Y=1.557
+ $X2=9.985 $Y2=1.557
r80 47 49 32.7446 $w=3.68e-07 $l=2.5e-07 $layer=POLY_cond $X=9.73 $Y=1.557
+ $X2=9.98 $Y2=1.557
r81 47 48 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=9.73
+ $Y=1.515 $X2=9.73 $Y2=1.515
r82 45 47 23.5761 $w=3.68e-07 $l=1.8e-07 $layer=POLY_cond $X=9.55 $Y=1.557
+ $X2=9.73 $Y2=1.557
r83 44 45 1.96467 $w=3.68e-07 $l=1.5e-08 $layer=POLY_cond $X=9.535 $Y=1.557
+ $X2=9.55 $Y2=1.557
r84 43 44 54.356 $w=3.68e-07 $l=4.15e-07 $layer=POLY_cond $X=9.12 $Y=1.557
+ $X2=9.535 $Y2=1.557
r85 42 43 4.58424 $w=3.68e-07 $l=3.5e-08 $layer=POLY_cond $X=9.085 $Y=1.557
+ $X2=9.12 $Y2=1.557
r86 40 42 49.1168 $w=3.68e-07 $l=3.75e-07 $layer=POLY_cond $X=8.71 $Y=1.557
+ $X2=9.085 $Y2=1.557
r87 40 41 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=8.71
+ $Y=1.515 $X2=8.71 $Y2=1.515
r88 38 40 2.61957 $w=3.68e-07 $l=2e-08 $layer=POLY_cond $X=8.69 $Y=1.557
+ $X2=8.71 $Y2=1.557
r89 37 38 7.2038 $w=3.68e-07 $l=5.5e-08 $layer=POLY_cond $X=8.635 $Y=1.557
+ $X2=8.69 $Y2=1.557
r90 32 48 2.94811 $w=4.28e-07 $l=1.1e-07 $layer=LI1_cond $X=9.84 $Y=1.565
+ $X2=9.73 $Y2=1.565
r91 31 48 9.91637 $w=4.28e-07 $l=3.7e-07 $layer=LI1_cond $X=9.36 $Y=1.565
+ $X2=9.73 $Y2=1.565
r92 30 31 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=8.88 $Y=1.565
+ $X2=9.36 $Y2=1.565
r93 30 41 4.55617 $w=4.28e-07 $l=1.7e-07 $layer=LI1_cond $X=8.88 $Y=1.565
+ $X2=8.71 $Y2=1.565
r94 29 41 8.30831 $w=4.28e-07 $l=3.1e-07 $layer=LI1_cond $X=8.4 $Y=1.565
+ $X2=8.71 $Y2=1.565
r95 26 50 23.8357 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=9.985 $Y=1.765
+ $X2=9.985 $Y2=1.557
r96 26 28 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=9.985 $Y=1.765
+ $X2=9.985 $Y2=2.4
r97 22 49 23.8357 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=9.98 $Y=1.35
+ $X2=9.98 $Y2=1.557
r98 22 24 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=9.98 $Y=1.35
+ $X2=9.98 $Y2=0.74
r99 18 45 23.8357 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=9.55 $Y=1.35
+ $X2=9.55 $Y2=1.557
r100 18 20 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=9.55 $Y=1.35
+ $X2=9.55 $Y2=0.74
r101 15 44 23.8357 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=9.535 $Y=1.765
+ $X2=9.535 $Y2=1.557
r102 15 17 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=9.535 $Y=1.765
+ $X2=9.535 $Y2=2.4
r103 11 43 23.8357 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=9.12 $Y=1.35
+ $X2=9.12 $Y2=1.557
r104 11 13 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=9.12 $Y=1.35
+ $X2=9.12 $Y2=0.74
r105 8 42 23.8357 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=9.085 $Y=1.765
+ $X2=9.085 $Y2=1.557
r106 8 10 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=9.085 $Y=1.765
+ $X2=9.085 $Y2=2.4
r107 4 38 23.8357 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=8.69 $Y=1.35
+ $X2=8.69 $Y2=1.557
r108 4 6 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=8.69 $Y=1.35 $X2=8.69
+ $Y2=0.74
r109 1 37 23.8357 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=8.635 $Y=1.765
+ $X2=8.635 $Y2=1.557
r110 1 3 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=8.635 $Y=1.765
+ $X2=8.635 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_HS__A221OI_4%Y 1 2 3 4 5 6 7 8 9 10 31 32 33 37 41 43 45
+ 49 53 55 59 61 65 74 75 76 77 78 79 80 82 83 85 86 87 88 89 90 91 102 121
c162 82 0 8.01953e-20 $X=8.045 $Y=0.95
r163 108 121 2.39067 $w=4.05e-07 $l=1.14782e-07 $layer=LI1_cond $X=0.23 $Y=1.18
+ $X2=0.3 $Y2=1.095
r164 90 91 17.0562 $w=2.48e-07 $l=3.7e-07 $layer=LI1_cond $X=0.23 $Y=2.405
+ $X2=0.23 $Y2=2.775
r165 89 90 19.361 $w=2.48e-07 $l=4.2e-07 $layer=LI1_cond $X=0.23 $Y=1.985
+ $X2=0.23 $Y2=2.405
r166 88 89 14.7513 $w=2.48e-07 $l=3.2e-07 $layer=LI1_cond $X=0.23 $Y=1.665
+ $X2=0.23 $Y2=1.985
r167 87 88 17.0562 $w=2.48e-07 $l=3.7e-07 $layer=LI1_cond $X=0.23 $Y=1.295
+ $X2=0.23 $Y2=1.665
r168 87 108 5.30124 $w=2.48e-07 $l=1.15e-07 $layer=LI1_cond $X=0.23 $Y=1.295
+ $X2=0.23 $Y2=1.18
r169 86 121 2.39067 $w=4.05e-07 $l=1.11018e-07 $layer=LI1_cond $X=0.24 $Y=1.01
+ $X2=0.3 $Y2=1.095
r170 85 86 10.9334 $w=3.88e-07 $l=3.7e-07 $layer=LI1_cond $X=0.3 $Y=0.555
+ $X2=0.3 $Y2=0.925
r171 85 102 1.18199 $w=3.88e-07 $l=4e-08 $layer=LI1_cond $X=0.3 $Y=0.555 $X2=0.3
+ $Y2=0.515
r172 82 83 4.12636 $w=4.08e-07 $l=1.3e-07 $layer=LI1_cond $X=8.045 $Y=0.975
+ $X2=7.915 $Y2=0.975
r173 79 80 8.63679 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=6.36 $Y=1.055
+ $X2=6.53 $Y2=1.055
r174 73 91 5.9927 $w=2.48e-07 $l=1.3e-07 $layer=LI1_cond $X=0.23 $Y=2.905
+ $X2=0.23 $Y2=2.775
r175 72 83 25.4934 $w=3.28e-07 $l=7.3e-07 $layer=LI1_cond $X=7.185 $Y=1.015
+ $X2=7.915 $Y2=1.015
r176 72 80 22.8742 $w=3.28e-07 $l=6.55e-07 $layer=LI1_cond $X=7.185 $Y=1.015
+ $X2=6.53 $Y2=1.015
r177 68 78 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=5.9 $Y=1.175
+ $X2=5.805 $Y2=1.175
r178 68 79 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=5.9 $Y=1.175
+ $X2=6.36 $Y2=1.175
r179 63 78 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=5.805 $Y=1.09
+ $X2=5.805 $Y2=1.175
r180 63 65 16.6364 $w=1.88e-07 $l=2.85e-07 $layer=LI1_cond $X=5.805 $Y=1.09
+ $X2=5.805 $Y2=0.805
r181 62 77 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=5.04 $Y=1.175
+ $X2=4.945 $Y2=1.175
r182 61 78 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=5.71 $Y=1.175
+ $X2=5.805 $Y2=1.175
r183 61 62 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.71 $Y=1.175
+ $X2=5.04 $Y2=1.175
r184 57 77 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=4.945 $Y=1.09
+ $X2=4.945 $Y2=1.175
r185 57 59 16.6364 $w=1.88e-07 $l=2.85e-07 $layer=LI1_cond $X=4.945 $Y=1.09
+ $X2=4.945 $Y2=0.805
r186 56 76 7.02821 $w=1.7e-07 $l=1.43614e-07 $layer=LI1_cond $X=2.295 $Y=1.175
+ $X2=2.17 $Y2=1.135
r187 55 77 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=4.85 $Y=1.175
+ $X2=4.945 $Y2=1.175
r188 55 56 166.69 $w=1.68e-07 $l=2.555e-06 $layer=LI1_cond $X=4.85 $Y=1.175
+ $X2=2.295 $Y2=1.175
r189 51 76 0.00168595 $w=2.5e-07 $l=1.25e-07 $layer=LI1_cond $X=2.17 $Y=1.01
+ $X2=2.17 $Y2=1.135
r190 51 53 22.8184 $w=2.48e-07 $l=4.95e-07 $layer=LI1_cond $X=2.17 $Y=1.01
+ $X2=2.17 $Y2=0.515
r191 47 49 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=2.07 $Y=2.905
+ $X2=2.07 $Y2=2.41
r192 46 75 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.355 $Y=1.095
+ $X2=1.27 $Y2=1.095
r193 45 76 7.02821 $w=1.7e-07 $l=1.43614e-07 $layer=LI1_cond $X=2.045 $Y=1.095
+ $X2=2.17 $Y2=1.135
r194 45 46 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=2.045 $Y=1.095
+ $X2=1.355 $Y2=1.095
r195 44 74 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.335 $Y=2.99
+ $X2=1.17 $Y2=2.99
r196 43 47 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.905 $Y=2.99
+ $X2=2.07 $Y2=2.905
r197 43 44 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=1.905 $Y=2.99
+ $X2=1.335 $Y2=2.99
r198 39 75 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.27 $Y=1.01
+ $X2=1.27 $Y2=1.095
r199 39 41 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=1.27 $Y=1.01
+ $X2=1.27 $Y2=0.515
r200 35 74 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.17 $Y=2.905
+ $X2=1.17 $Y2=2.99
r201 35 37 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=1.17 $Y=2.905
+ $X2=1.17 $Y2=2.41
r202 34 121 4.59089 $w=1.7e-07 $l=1.95e-07 $layer=LI1_cond $X=0.495 $Y=1.095
+ $X2=0.3 $Y2=1.095
r203 33 75 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.185 $Y=1.095
+ $X2=1.27 $Y2=1.095
r204 33 34 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.185 $Y=1.095
+ $X2=0.495 $Y2=1.095
r205 32 73 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.355 $Y=2.99
+ $X2=0.23 $Y2=2.905
r206 31 74 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.005 $Y=2.99
+ $X2=1.17 $Y2=2.99
r207 31 32 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=1.005 $Y=2.99
+ $X2=0.355 $Y2=2.99
r208 10 49 300 $w=1.7e-07 $l=6.40625e-07 $layer=licon1_PDIFF $count=2 $X=1.92
+ $Y=1.84 $X2=2.07 $Y2=2.41
r209 9 37 300 $w=1.7e-07 $l=6.40625e-07 $layer=licon1_PDIFF $count=2 $X=1.02
+ $Y=1.84 $X2=1.17 $Y2=2.41
r210 8 91 400 $w=1.7e-07 $l=1.03562e-06 $layer=licon1_PDIFF $count=1 $X=0.145
+ $Y=1.84 $X2=0.27 $Y2=2.815
r211 8 89 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.145
+ $Y=1.84 $X2=0.27 $Y2=1.985
r212 7 82 182 $w=1.7e-07 $l=6.4622e-07 $layer=licon1_NDIFF $count=1 $X=7.905
+ $Y=0.37 $X2=8.045 $Y2=0.95
r213 6 72 182 $w=1.7e-07 $l=6.4622e-07 $layer=licon1_NDIFF $count=1 $X=7.045
+ $Y=0.37 $X2=7.185 $Y2=0.95
r214 5 65 182 $w=1.7e-07 $l=5.00125e-07 $layer=licon1_NDIFF $count=1 $X=5.665
+ $Y=0.37 $X2=5.805 $Y2=0.805
r215 4 59 182 $w=1.7e-07 $l=5.00125e-07 $layer=licon1_NDIFF $count=1 $X=4.805
+ $Y=0.37 $X2=4.945 $Y2=0.805
r216 3 53 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.99
+ $Y=0.37 $X2=2.13 $Y2=0.515
r217 2 41 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.13
+ $Y=0.37 $X2=1.27 $Y2=0.515
r218 1 102 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.285
+ $Y=0.37 $X2=0.41 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__A221OI_4%A_114_368# 1 2 3 4 5 6 19 21 23 27 29 33 37
+ 41 48 50 52 54 56
c105 37 0 1.45655e-19 $X=8.695 $Y=2.035
r106 42 54 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.025 $Y=2.035
+ $X2=8.86 $Y2=2.035
r107 41 56 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.595 $Y=2.035
+ $X2=9.76 $Y2=2.035
r108 41 42 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=9.595 $Y=2.035
+ $X2=9.025 $Y2=2.035
r109 38 52 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.125 $Y=2.035
+ $X2=7.96 $Y2=2.035
r110 37 54 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.695 $Y=2.035
+ $X2=8.86 $Y2=2.035
r111 37 38 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=8.695 $Y=2.035
+ $X2=8.125 $Y2=2.035
r112 34 50 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.225 $Y=2.035
+ $X2=7.06 $Y2=2.035
r113 33 52 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.795 $Y=2.035
+ $X2=7.96 $Y2=2.035
r114 33 34 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=7.795 $Y=2.035
+ $X2=7.225 $Y2=2.035
r115 30 48 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=1.735 $Y=2.035
+ $X2=1.62 $Y2=2.035
r116 29 50 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.895 $Y=2.035
+ $X2=7.06 $Y2=2.035
r117 29 30 336.642 $w=1.68e-07 $l=5.16e-06 $layer=LI1_cond $X=6.895 $Y=2.035
+ $X2=1.735 $Y2=2.035
r118 25 48 0.280307 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.62 $Y=2.12
+ $X2=1.62 $Y2=2.035
r119 25 27 22.5478 $w=2.28e-07 $l=4.5e-07 $layer=LI1_cond $X=1.62 $Y=2.12
+ $X2=1.62 $Y2=2.57
r120 24 46 4.57959 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=0.835 $Y=2.035
+ $X2=0.695 $Y2=2.035
r121 23 48 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=1.505 $Y=2.035
+ $X2=1.62 $Y2=2.035
r122 23 24 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.505 $Y=2.035
+ $X2=0.835 $Y2=2.035
r123 19 46 2.78046 $w=2.8e-07 $l=8.5e-08 $layer=LI1_cond $X=0.695 $Y=2.12
+ $X2=0.695 $Y2=2.035
r124 19 21 18.5214 $w=2.78e-07 $l=4.5e-07 $layer=LI1_cond $X=0.695 $Y=2.12
+ $X2=0.695 $Y2=2.57
r125 6 56 300 $w=1.7e-07 $l=2.59374e-07 $layer=licon1_PDIFF $count=2 $X=9.61
+ $Y=1.84 $X2=9.76 $Y2=2.035
r126 5 54 300 $w=1.7e-07 $l=2.59374e-07 $layer=licon1_PDIFF $count=2 $X=8.71
+ $Y=1.84 $X2=8.86 $Y2=2.035
r127 4 52 300 $w=1.7e-07 $l=2.59374e-07 $layer=licon1_PDIFF $count=2 $X=7.81
+ $Y=1.84 $X2=7.96 $Y2=2.035
r128 3 50 300 $w=1.7e-07 $l=2.59374e-07 $layer=licon1_PDIFF $count=2 $X=6.91
+ $Y=1.84 $X2=7.06 $Y2=2.035
r129 2 48 600 $w=1.7e-07 $l=2.59374e-07 $layer=licon1_PDIFF $count=1 $X=1.47
+ $Y=1.84 $X2=1.62 $Y2=2.035
r130 2 27 600 $w=1.7e-07 $l=8.01499e-07 $layer=licon1_PDIFF $count=1 $X=1.47
+ $Y=1.84 $X2=1.62 $Y2=2.57
r131 1 46 600 $w=1.7e-07 $l=2.59374e-07 $layer=licon1_PDIFF $count=1 $X=0.57
+ $Y=1.84 $X2=0.72 $Y2=2.035
r132 1 21 600 $w=1.7e-07 $l=8.01499e-07 $layer=licon1_PDIFF $count=1 $X=0.57
+ $Y=1.84 $X2=0.72 $Y2=2.57
.ends

.subckt PM_SKY130_FD_SC_HS__A221OI_4%A_531_368# 1 2 3 4 5 6 7 8 9 30 34 38 42 44
+ 45 46 47 50 52 56 58 62 64 68 73 75 77 79 82 83 84
r121 68 71 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=10.25 $Y=1.985
+ $X2=10.25 $Y2=2.815
r122 66 71 4.14879 $w=2.48e-07 $l=9e-08 $layer=LI1_cond $X=10.25 $Y=2.905
+ $X2=10.25 $Y2=2.815
r123 65 84 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=9.425 $Y=2.99
+ $X2=9.31 $Y2=2.99
r124 64 66 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=10.125 $Y=2.99
+ $X2=10.25 $Y2=2.905
r125 64 65 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=10.125 $Y=2.99
+ $X2=9.425 $Y2=2.99
r126 60 84 0.280307 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.31 $Y=2.905
+ $X2=9.31 $Y2=2.99
r127 60 62 22.5478 $w=2.28e-07 $l=4.5e-07 $layer=LI1_cond $X=9.31 $Y=2.905
+ $X2=9.31 $Y2=2.455
r128 59 83 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=8.525 $Y=2.99
+ $X2=8.41 $Y2=2.99
r129 58 84 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=9.195 $Y=2.99
+ $X2=9.31 $Y2=2.99
r130 58 59 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=9.195 $Y=2.99
+ $X2=8.525 $Y2=2.99
r131 54 83 0.280307 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.41 $Y=2.905
+ $X2=8.41 $Y2=2.99
r132 54 56 22.5478 $w=2.28e-07 $l=4.5e-07 $layer=LI1_cond $X=8.41 $Y=2.905
+ $X2=8.41 $Y2=2.455
r133 53 82 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=7.625 $Y=2.99
+ $X2=7.51 $Y2=2.99
r134 52 83 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=8.295 $Y=2.99
+ $X2=8.41 $Y2=2.99
r135 52 53 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=8.295 $Y=2.99
+ $X2=7.625 $Y2=2.99
r136 48 82 0.280307 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.51 $Y=2.905
+ $X2=7.51 $Y2=2.99
r137 48 50 22.5478 $w=2.28e-07 $l=4.5e-07 $layer=LI1_cond $X=7.51 $Y=2.905
+ $X2=7.51 $Y2=2.455
r138 46 82 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=7.395 $Y=2.99
+ $X2=7.51 $Y2=2.99
r139 46 47 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=7.395 $Y=2.99
+ $X2=6.725 $Y2=2.99
r140 45 47 7.36005 $w=1.7e-07 $l=1.77482e-07 $layer=LI1_cond $X=6.585 $Y=2.905
+ $X2=6.725 $Y2=2.99
r141 44 81 2.78046 $w=2.8e-07 $l=8.5e-08 $layer=LI1_cond $X=6.585 $Y=2.46
+ $X2=6.585 $Y2=2.375
r142 44 45 18.3156 $w=2.78e-07 $l=4.45e-07 $layer=LI1_cond $X=6.585 $Y=2.46
+ $X2=6.585 $Y2=2.905
r143 43 79 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.645 $Y=2.375
+ $X2=5.48 $Y2=2.375
r144 42 81 4.57959 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=6.445 $Y=2.375
+ $X2=6.585 $Y2=2.375
r145 42 43 52.1925 $w=1.68e-07 $l=8e-07 $layer=LI1_cond $X=6.445 $Y=2.375
+ $X2=5.645 $Y2=2.375
r146 39 77 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.745 $Y=2.375
+ $X2=4.58 $Y2=2.375
r147 38 79 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.315 $Y=2.375
+ $X2=5.48 $Y2=2.375
r148 38 39 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=5.315 $Y=2.375
+ $X2=4.745 $Y2=2.375
r149 35 75 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.845 $Y=2.375
+ $X2=3.68 $Y2=2.375
r150 34 77 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.415 $Y=2.375
+ $X2=4.58 $Y2=2.375
r151 34 35 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=4.415 $Y=2.375
+ $X2=3.845 $Y2=2.375
r152 31 73 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.945 $Y=2.375
+ $X2=2.78 $Y2=2.375
r153 30 75 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.515 $Y=2.375
+ $X2=3.68 $Y2=2.375
r154 30 31 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=3.515 $Y=2.375
+ $X2=2.945 $Y2=2.375
r155 9 71 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=10.06
+ $Y=1.84 $X2=10.21 $Y2=2.815
r156 9 68 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=10.06
+ $Y=1.84 $X2=10.21 $Y2=1.985
r157 8 62 300 $w=1.7e-07 $l=6.85912e-07 $layer=licon1_PDIFF $count=2 $X=9.16
+ $Y=1.84 $X2=9.31 $Y2=2.455
r158 7 56 300 $w=1.7e-07 $l=6.85912e-07 $layer=licon1_PDIFF $count=2 $X=8.26
+ $Y=1.84 $X2=8.41 $Y2=2.455
r159 6 50 300 $w=1.7e-07 $l=6.85912e-07 $layer=licon1_PDIFF $count=2 $X=7.36
+ $Y=1.84 $X2=7.51 $Y2=2.455
r160 5 81 300 $w=1.7e-07 $l=6.85912e-07 $layer=licon1_PDIFF $count=2 $X=6.46
+ $Y=1.84 $X2=6.61 $Y2=2.455
r161 4 79 300 $w=1.7e-07 $l=6.30555e-07 $layer=licon1_PDIFF $count=2 $X=5.33
+ $Y=1.84 $X2=5.48 $Y2=2.4
r162 3 77 300 $w=1.7e-07 $l=6.30555e-07 $layer=licon1_PDIFF $count=2 $X=4.43
+ $Y=1.84 $X2=4.58 $Y2=2.4
r163 2 75 300 $w=1.7e-07 $l=6.30555e-07 $layer=licon1_PDIFF $count=2 $X=3.53
+ $Y=1.84 $X2=3.68 $Y2=2.4
r164 1 73 300 $w=1.7e-07 $l=6.19354e-07 $layer=licon1_PDIFF $count=2 $X=2.655
+ $Y=1.84 $X2=2.78 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_HS__A221OI_4%VPWR 1 2 3 4 15 17 21 25 29 31 32 34 35 36
+ 49 58 59 62 65
r115 65 66 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r116 62 63 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r117 58 59 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=10.32 $Y=3.33
+ $X2=10.32 $Y2=3.33
r118 56 59 1.07034 $w=4.9e-07 $l=3.84e-06 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=10.32 $Y2=3.33
r119 56 66 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=3.33 $X2=6
+ $Y2=3.33
r120 55 58 250.524 $w=1.68e-07 $l=3.84e-06 $layer=LI1_cond $X=6.48 $Y=3.33
+ $X2=10.32 $Y2=3.33
r121 55 56 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r122 53 65 10.7288 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=6.275 $Y=3.33
+ $X2=6.045 $Y2=3.33
r123 53 55 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=6.275 $Y=3.33
+ $X2=6.48 $Y2=3.33
r124 52 66 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=3.33 $X2=6
+ $Y2=3.33
r125 51 52 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r126 49 65 10.7288 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=5.815 $Y=3.33
+ $X2=6.045 $Y2=3.33
r127 49 51 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=5.815 $Y=3.33
+ $X2=5.52 $Y2=3.33
r128 48 63 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=4.08 $Y2=3.33
r129 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r130 45 62 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.215 $Y=3.33
+ $X2=4.13 $Y2=3.33
r131 45 47 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=4.215 $Y=3.33
+ $X2=4.56 $Y2=3.33
r132 44 63 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=4.08 $Y2=3.33
r133 43 44 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r134 40 44 0.802756 $w=4.9e-07 $l=2.88e-06 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=3.12 $Y2=3.33
r135 39 43 187.893 $w=1.68e-07 $l=2.88e-06 $layer=LI1_cond $X=0.24 $Y=3.33
+ $X2=3.12 $Y2=3.33
r136 39 40 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r137 36 52 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=5.28 $Y=3.33
+ $X2=5.52 $Y2=3.33
r138 36 48 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=5.28 $Y=3.33
+ $X2=4.56 $Y2=3.33
r139 34 47 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=4.945 $Y=3.33
+ $X2=4.56 $Y2=3.33
r140 34 35 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.945 $Y=3.33
+ $X2=5.03 $Y2=3.33
r141 33 51 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=5.115 $Y=3.33
+ $X2=5.52 $Y2=3.33
r142 33 35 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.115 $Y=3.33
+ $X2=5.03 $Y2=3.33
r143 31 43 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=3.145 $Y=3.33
+ $X2=3.12 $Y2=3.33
r144 31 32 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.145 $Y=3.33
+ $X2=3.23 $Y2=3.33
r145 27 65 1.85547 $w=4.6e-07 $l=8.5e-08 $layer=LI1_cond $X=6.045 $Y=3.245
+ $X2=6.045 $Y2=3.33
r146 27 29 11.4408 $w=4.58e-07 $l=4.4e-07 $layer=LI1_cond $X=6.045 $Y=3.245
+ $X2=6.045 $Y2=2.805
r147 23 35 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.03 $Y=3.245
+ $X2=5.03 $Y2=3.33
r148 23 25 28.7059 $w=1.68e-07 $l=4.4e-07 $layer=LI1_cond $X=5.03 $Y=3.245
+ $X2=5.03 $Y2=2.805
r149 19 62 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.13 $Y=3.245
+ $X2=4.13 $Y2=3.33
r150 19 21 28.7059 $w=1.68e-07 $l=4.4e-07 $layer=LI1_cond $X=4.13 $Y=3.245
+ $X2=4.13 $Y2=2.805
r151 18 32 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.315 $Y=3.33
+ $X2=3.23 $Y2=3.33
r152 17 62 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.045 $Y=3.33
+ $X2=4.13 $Y2=3.33
r153 17 18 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=4.045 $Y=3.33
+ $X2=3.315 $Y2=3.33
r154 13 32 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.23 $Y=3.245
+ $X2=3.23 $Y2=3.33
r155 13 15 28.7059 $w=1.68e-07 $l=4.4e-07 $layer=LI1_cond $X=3.23 $Y=3.245
+ $X2=3.23 $Y2=2.805
r156 4 29 600 $w=1.7e-07 $l=1.08947e-06 $layer=licon1_PDIFF $count=1 $X=5.78
+ $Y=1.84 $X2=6.045 $Y2=2.805
r157 3 25 600 $w=1.7e-07 $l=1.03729e-06 $layer=licon1_PDIFF $count=1 $X=4.88
+ $Y=1.84 $X2=5.03 $Y2=2.805
r158 2 21 600 $w=1.7e-07 $l=1.03729e-06 $layer=licon1_PDIFF $count=1 $X=3.98
+ $Y=1.84 $X2=4.13 $Y2=2.805
r159 1 15 600 $w=1.7e-07 $l=1.03729e-06 $layer=licon1_PDIFF $count=1 $X=3.08
+ $Y=1.84 $X2=3.23 $Y2=2.805
.ends

.subckt PM_SKY130_FD_SC_HS__A221OI_4%VGND 1 2 3 4 5 6 23 27 31 35 39 43 45 47 52
+ 57 62 70 77 78 81 84 87 90 93 96
r140 96 97 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.84 $Y=0 $X2=9.84
+ $Y2=0
r141 93 94 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=0 $X2=8.88
+ $Y2=0
r142 90 91 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r143 87 88 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r144 84 85 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r145 81 82 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r146 78 97 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.32 $Y=0
+ $X2=9.84 $Y2=0
r147 77 78 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.32 $Y=0
+ $X2=10.32 $Y2=0
r148 75 96 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.93 $Y=0 $X2=9.765
+ $Y2=0
r149 75 77 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=9.93 $Y=0 $X2=10.32
+ $Y2=0
r150 74 97 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.36 $Y=0 $X2=9.84
+ $Y2=0
r151 74 94 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.36 $Y=0 $X2=8.88
+ $Y2=0
r152 73 74 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.36 $Y=0 $X2=9.36
+ $Y2=0
r153 71 93 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.07 $Y=0 $X2=8.905
+ $Y2=0
r154 71 73 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=9.07 $Y=0 $X2=9.36
+ $Y2=0
r155 70 96 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.6 $Y=0 $X2=9.765
+ $Y2=0
r156 70 73 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=9.6 $Y=0 $X2=9.36
+ $Y2=0
r157 69 94 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=0 $X2=8.88
+ $Y2=0
r158 68 69 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=8.4 $Y=0
+ $X2=8.4 $Y2=0
r159 66 91 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=4.08
+ $Y2=0
r160 65 68 250.524 $w=1.68e-07 $l=3.84e-06 $layer=LI1_cond $X=4.56 $Y=0 $X2=8.4
+ $Y2=0
r161 65 66 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=4.56 $Y=0
+ $X2=4.56 $Y2=0
r162 63 90 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.25 $Y=0 $X2=4.085
+ $Y2=0
r163 63 65 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=4.25 $Y=0 $X2=4.56
+ $Y2=0
r164 62 93 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.74 $Y=0 $X2=8.905
+ $Y2=0
r165 62 68 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=8.74 $Y=0 $X2=8.4
+ $Y2=0
r166 61 91 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.08
+ $Y2=0
r167 61 88 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=3.12
+ $Y2=0
r168 60 61 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r169 58 87 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.39 $Y=0 $X2=3.225
+ $Y2=0
r170 58 60 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=3.39 $Y=0 $X2=3.6
+ $Y2=0
r171 57 90 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.92 $Y=0 $X2=4.085
+ $Y2=0
r172 57 60 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=3.92 $Y=0 $X2=3.6
+ $Y2=0
r173 56 88 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=3.12
+ $Y2=0
r174 56 85 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.68
+ $Y2=0
r175 55 56 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r176 53 84 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.865 $Y=0 $X2=1.7
+ $Y2=0
r177 53 55 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=1.865 $Y=0 $X2=2.16
+ $Y2=0
r178 52 87 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.06 $Y=0 $X2=3.225
+ $Y2=0
r179 52 55 58.7166 $w=1.68e-07 $l=9e-07 $layer=LI1_cond $X=3.06 $Y=0 $X2=2.16
+ $Y2=0
r180 51 85 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=1.68
+ $Y2=0
r181 51 82 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r182 50 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r183 48 81 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.005 $Y=0 $X2=0.84
+ $Y2=0
r184 48 50 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=1.005 $Y=0 $X2=1.2
+ $Y2=0
r185 47 84 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.535 $Y=0 $X2=1.7
+ $Y2=0
r186 47 50 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=1.535 $Y=0 $X2=1.2
+ $Y2=0
r187 45 69 0.869652 $w=4.9e-07 $l=3.12e-06 $layer=MET1_cond $X=5.28 $Y=0 $X2=8.4
+ $Y2=0
r188 45 66 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=5.28 $Y=0 $X2=4.56
+ $Y2=0
r189 41 96 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.765 $Y=0.085
+ $X2=9.765 $Y2=0
r190 41 43 20.6043 $w=3.28e-07 $l=5.9e-07 $layer=LI1_cond $X=9.765 $Y=0.085
+ $X2=9.765 $Y2=0.675
r191 37 93 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.905 $Y=0.085
+ $X2=8.905 $Y2=0
r192 37 39 20.6043 $w=3.28e-07 $l=5.9e-07 $layer=LI1_cond $X=8.905 $Y=0.085
+ $X2=8.905 $Y2=0.675
r193 33 90 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.085 $Y=0.085
+ $X2=4.085 $Y2=0
r194 33 35 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=4.085 $Y=0.085
+ $X2=4.085 $Y2=0.495
r195 29 87 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.225 $Y=0.085
+ $X2=3.225 $Y2=0
r196 29 31 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=3.225 $Y=0.085
+ $X2=3.225 $Y2=0.495
r197 25 84 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.7 $Y=0.085 $X2=1.7
+ $Y2=0
r198 25 27 20.6043 $w=3.28e-07 $l=5.9e-07 $layer=LI1_cond $X=1.7 $Y=0.085
+ $X2=1.7 $Y2=0.675
r199 21 81 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.84 $Y=0.085
+ $X2=0.84 $Y2=0
r200 21 23 20.6043 $w=3.28e-07 $l=5.9e-07 $layer=LI1_cond $X=0.84 $Y=0.085
+ $X2=0.84 $Y2=0.675
r201 6 43 182 $w=1.7e-07 $l=3.68409e-07 $layer=licon1_NDIFF $count=1 $X=9.625
+ $Y=0.37 $X2=9.765 $Y2=0.675
r202 5 39 182 $w=1.7e-07 $l=3.68409e-07 $layer=licon1_NDIFF $count=1 $X=8.765
+ $Y=0.37 $X2=8.905 $Y2=0.675
r203 4 35 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=3.945
+ $Y=0.37 $X2=4.085 $Y2=0.495
r204 3 31 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=3.085
+ $Y=0.37 $X2=3.225 $Y2=0.495
r205 2 27 182 $w=1.7e-07 $l=3.68409e-07 $layer=licon1_NDIFF $count=1 $X=1.56
+ $Y=0.37 $X2=1.7 $Y2=0.675
r206 1 23 182 $w=1.7e-07 $l=3.68409e-07 $layer=licon1_NDIFF $count=1 $X=0.7
+ $Y=0.37 $X2=0.84 $Y2=0.675
.ends

.subckt PM_SKY130_FD_SC_HS__A221OI_4%A_534_74# 1 2 3 4 5 18 20 21 24 26 29 31 32
+ 33 36 38 40 43 44
r86 44 47 4.53993 $w=3.28e-07 $l=1.3e-07 $layer=LI1_cond $X=6.235 $Y=0.385
+ $X2=6.235 $Y2=0.515
r87 39 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.54 $Y=0.385
+ $X2=5.375 $Y2=0.385
r88 38 44 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.07 $Y=0.385
+ $X2=6.235 $Y2=0.385
r89 38 39 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=6.07 $Y=0.385
+ $X2=5.54 $Y2=0.385
r90 34 43 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.375 $Y=0.47
+ $X2=5.375 $Y2=0.385
r91 34 36 0.873063 $w=3.28e-07 $l=2.5e-08 $layer=LI1_cond $X=5.375 $Y=0.47
+ $X2=5.375 $Y2=0.495
r92 32 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.21 $Y=0.385
+ $X2=5.375 $Y2=0.385
r93 32 33 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=5.21 $Y=0.385
+ $X2=4.68 $Y2=0.385
r94 29 42 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.555 $Y=0.75
+ $X2=4.555 $Y2=0.835
r95 29 31 11.7549 $w=2.48e-07 $l=2.55e-07 $layer=LI1_cond $X=4.555 $Y=0.75
+ $X2=4.555 $Y2=0.495
r96 28 33 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=4.555 $Y=0.47
+ $X2=4.68 $Y2=0.385
r97 28 31 1.15244 $w=2.48e-07 $l=2.5e-08 $layer=LI1_cond $X=4.555 $Y=0.47
+ $X2=4.555 $Y2=0.495
r98 27 40 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.74 $Y=0.835
+ $X2=3.655 $Y2=0.835
r99 26 42 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.43 $Y=0.835
+ $X2=4.555 $Y2=0.835
r100 26 27 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=4.43 $Y=0.835
+ $X2=3.74 $Y2=0.835
r101 22 40 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.655 $Y=0.75
+ $X2=3.655 $Y2=0.835
r102 22 24 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=3.655 $Y=0.75
+ $X2=3.655 $Y2=0.635
r103 20 40 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.57 $Y=0.835
+ $X2=3.655 $Y2=0.835
r104 20 21 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=3.57 $Y=0.835
+ $X2=2.88 $Y2=0.835
r105 16 21 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=2.755 $Y=0.75
+ $X2=2.88 $Y2=0.835
r106 16 18 5.30124 $w=2.48e-07 $l=1.15e-07 $layer=LI1_cond $X=2.755 $Y=0.75
+ $X2=2.755 $Y2=0.635
r107 5 47 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=6.095
+ $Y=0.37 $X2=6.235 $Y2=0.515
r108 4 36 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=5.235
+ $Y=0.37 $X2=5.375 $Y2=0.495
r109 3 42 182 $w=1.7e-07 $l=5.30401e-07 $layer=licon1_NDIFF $count=1 $X=4.375
+ $Y=0.37 $X2=4.515 $Y2=0.835
r110 3 31 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=4.375
+ $Y=0.37 $X2=4.515 $Y2=0.495
r111 2 24 182 $w=1.7e-07 $l=3.27605e-07 $layer=licon1_NDIFF $count=1 $X=3.515
+ $Y=0.37 $X2=3.655 $Y2=0.635
r112 1 18 182 $w=1.7e-07 $l=3.21481e-07 $layer=licon1_NDIFF $count=1 $X=2.67
+ $Y=0.37 $X2=2.795 $Y2=0.635
.ends

.subckt PM_SKY130_FD_SC_HS__A221OI_4%A_1326_74# 1 2 3 4 5 18 20 24 25 28 30 34
+ 39 42 43 46
c64 20 0 1.6164e-19 $X=8.475 $Y=0.6
r65 41 43 5.24459 $w=3.28e-07 $l=1.3e-07 $layer=LI1_cond $X=7.615 $Y=0.515
+ $X2=7.745 $Y2=0.515
r66 41 42 6.46688 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=7.615 $Y=0.515
+ $X2=7.45 $Y2=0.515
r67 39 42 24.4318 $w=2.48e-07 $l=5.3e-07 $layer=LI1_cond $X=6.92 $Y=0.475
+ $X2=7.45 $Y2=0.475
r68 37 39 6.46688 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=6.755 $Y=0.515
+ $X2=6.92 $Y2=0.515
r69 32 34 22.8184 $w=2.48e-07 $l=4.95e-07 $layer=LI1_cond $X=10.235 $Y=1.01
+ $X2=10.235 $Y2=0.515
r70 31 46 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.42 $Y=1.095
+ $X2=9.335 $Y2=1.095
r71 30 32 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=10.11 $Y=1.095
+ $X2=10.235 $Y2=1.01
r72 30 31 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=10.11 $Y=1.095
+ $X2=9.42 $Y2=1.095
r73 26 46 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.335 $Y=1.01
+ $X2=9.335 $Y2=1.095
r74 26 28 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=9.335 $Y=1.01
+ $X2=9.335 $Y2=0.515
r75 24 46 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.25 $Y=1.095
+ $X2=9.335 $Y2=1.095
r76 24 25 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=9.25 $Y=1.095
+ $X2=8.56 $Y2=1.095
r77 21 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.475 $Y=1.01
+ $X2=8.56 $Y2=1.095
r78 21 23 2.93583 $w=1.68e-07 $l=4.5e-08 $layer=LI1_cond $X=8.475 $Y=1.01
+ $X2=8.475 $Y2=0.965
r79 20 45 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.475 $Y=0.6
+ $X2=8.475 $Y2=0.475
r80 20 23 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=8.475 $Y=0.6
+ $X2=8.475 $Y2=0.965
r81 18 45 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=8.39 $Y=0.475
+ $X2=8.475 $Y2=0.475
r82 18 43 29.733 $w=2.48e-07 $l=6.45e-07 $layer=LI1_cond $X=8.39 $Y=0.475
+ $X2=7.745 $Y2=0.475
r83 5 34 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=10.055
+ $Y=0.37 $X2=10.195 $Y2=0.515
r84 4 28 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=9.195
+ $Y=0.37 $X2=9.335 $Y2=0.515
r85 3 45 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=8.335
+ $Y=0.37 $X2=8.475 $Y2=0.515
r86 3 23 182 $w=1.7e-07 $l=6.61306e-07 $layer=licon1_NDIFF $count=1 $X=8.335
+ $Y=0.37 $X2=8.475 $Y2=0.965
r87 2 41 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=7.475
+ $Y=0.37 $X2=7.615 $Y2=0.515
r88 1 37 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=6.63
+ $Y=0.37 $X2=6.755 $Y2=0.515
.ends

