# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_hs__dlxtp_1
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_hs__dlxtp_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  7.680000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.208500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.180000 0.595000 1.850000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.541300 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.230000 1.820000 7.595000 2.980000 ;
        RECT 7.235000 0.390000 7.595000 1.150000 ;
        RECT 7.425000 1.150000 7.595000 1.820000 ;
    END
  END Q
  PIN GATE
    ANTENNAGATEAREA  0.237000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 6.365000 1.350000 6.715000 1.780000 ;
    END
  END GATE
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 7.680000 0.085000 ;
        RECT 0.115000  0.085000 0.445000 1.010000 ;
        RECT 1.675000  0.085000 2.005000 1.185000 ;
        RECT 4.995000  0.085000 5.325000 0.410000 ;
        RECT 6.590000  0.085000 7.055000 0.410000 ;
      LAYER mcon ;
        RECT 0.155000 -0.085000 0.325000 0.085000 ;
        RECT 0.635000 -0.085000 0.805000 0.085000 ;
        RECT 1.115000 -0.085000 1.285000 0.085000 ;
        RECT 1.595000 -0.085000 1.765000 0.085000 ;
        RECT 2.075000 -0.085000 2.245000 0.085000 ;
        RECT 2.555000 -0.085000 2.725000 0.085000 ;
        RECT 3.035000 -0.085000 3.205000 0.085000 ;
        RECT 3.515000 -0.085000 3.685000 0.085000 ;
        RECT 3.995000 -0.085000 4.165000 0.085000 ;
        RECT 4.475000 -0.085000 4.645000 0.085000 ;
        RECT 4.955000 -0.085000 5.125000 0.085000 ;
        RECT 5.435000 -0.085000 5.605000 0.085000 ;
        RECT 5.915000 -0.085000 6.085000 0.085000 ;
        RECT 6.395000 -0.085000 6.565000 0.085000 ;
        RECT 6.875000 -0.085000 7.045000 0.085000 ;
        RECT 7.355000 -0.085000 7.525000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.245000 7.680000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 3.245000 7.680000 3.415000 ;
        RECT 0.115000 2.100000 0.445000 3.245000 ;
        RECT 1.660000 2.955000 1.995000 3.245000 ;
        RECT 4.840000 2.845000 5.170000 3.245000 ;
        RECT 6.730000 1.950000 7.060000 3.245000 ;
      LAYER mcon ;
        RECT 0.155000 3.245000 0.325000 3.415000 ;
        RECT 0.635000 3.245000 0.805000 3.415000 ;
        RECT 1.115000 3.245000 1.285000 3.415000 ;
        RECT 1.595000 3.245000 1.765000 3.415000 ;
        RECT 2.075000 3.245000 2.245000 3.415000 ;
        RECT 2.555000 3.245000 2.725000 3.415000 ;
        RECT 3.035000 3.245000 3.205000 3.415000 ;
        RECT 3.515000 3.245000 3.685000 3.415000 ;
        RECT 3.995000 3.245000 4.165000 3.415000 ;
        RECT 4.475000 3.245000 4.645000 3.415000 ;
        RECT 4.955000 3.245000 5.125000 3.415000 ;
        RECT 5.435000 3.245000 5.605000 3.415000 ;
        RECT 5.915000 3.245000 6.085000 3.415000 ;
        RECT 6.395000 3.245000 6.565000 3.415000 ;
        RECT 6.875000 3.245000 7.045000 3.415000 ;
        RECT 7.355000 3.245000 7.525000 3.415000 ;
      LAYER met1 ;
        RECT 0.000000 3.085000 7.680000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.615000 0.420000 0.945000 1.010000 ;
      RECT 0.645000 2.100000 0.945000 2.980000 ;
      RECT 0.775000 1.010000 0.945000 1.100000 ;
      RECT 0.775000 1.100000 1.165000 1.770000 ;
      RECT 0.775000 1.770000 0.945000 2.100000 ;
      RECT 1.125000 1.940000 1.455000 2.615000 ;
      RECT 1.125000 2.615000 2.335000 2.735000 ;
      RECT 1.125000 2.735000 2.970000 2.785000 ;
      RECT 1.125000 2.785000 1.455000 2.980000 ;
      RECT 1.175000 0.405000 1.505000 0.930000 ;
      RECT 1.335000 0.930000 1.505000 1.355000 ;
      RECT 1.335000 1.355000 2.345000 1.525000 ;
      RECT 2.080000 1.940000 2.330000 2.275000 ;
      RECT 2.080000 2.275000 2.675000 2.395000 ;
      RECT 2.080000 2.395000 3.310000 2.445000 ;
      RECT 2.165000 2.785000 2.970000 2.985000 ;
      RECT 2.175000 0.255000 4.815000 0.425000 ;
      RECT 2.175000 0.425000 2.505000 0.585000 ;
      RECT 2.175000 0.755000 3.895000 0.765000 ;
      RECT 2.175000 0.765000 2.845000 0.925000 ;
      RECT 2.175000 0.925000 2.345000 1.355000 ;
      RECT 2.505000 2.445000 3.310000 2.565000 ;
      RECT 2.515000 1.095000 4.395000 1.105000 ;
      RECT 2.515000 1.105000 3.355000 1.265000 ;
      RECT 2.515000 1.265000 2.685000 1.935000 ;
      RECT 2.515000 1.935000 3.015000 2.055000 ;
      RECT 2.515000 2.055000 3.420000 2.105000 ;
      RECT 2.675000 0.595000 3.895000 0.755000 ;
      RECT 2.845000 2.105000 3.420000 2.225000 ;
      RECT 2.855000 1.435000 3.355000 1.715000 ;
      RECT 2.855000 1.715000 3.760000 1.765000 ;
      RECT 3.015000 0.935000 4.395000 1.095000 ;
      RECT 3.140000 2.565000 3.310000 2.845000 ;
      RECT 3.140000 2.845000 4.040000 3.015000 ;
      RECT 3.185000 1.765000 3.760000 1.885000 ;
      RECT 3.525000 1.275000 4.100000 1.545000 ;
      RECT 3.590000 1.885000 3.760000 2.505000 ;
      RECT 3.590000 2.505000 6.525000 2.675000 ;
      RECT 3.930000 1.545000 4.100000 2.165000 ;
      RECT 3.930000 2.165000 5.625000 2.335000 ;
      RECT 4.065000 0.775000 4.395000 0.935000 ;
      RECT 4.270000 1.665000 4.815000 1.995000 ;
      RECT 4.565000 0.425000 4.815000 0.580000 ;
      RECT 4.565000 0.580000 7.065000 0.750000 ;
      RECT 4.565000 0.750000 4.815000 1.665000 ;
      RECT 5.340000 2.675000 6.525000 2.700000 ;
      RECT 5.375000 0.920000 5.835000 1.170000 ;
      RECT 5.375000 1.170000 5.625000 2.165000 ;
      RECT 5.845000 1.350000 6.175000 1.950000 ;
      RECT 5.845000 1.950000 6.525000 2.505000 ;
      RECT 6.005000 0.920000 6.410000 1.170000 ;
      RECT 6.005000 1.170000 6.175000 1.350000 ;
      RECT 6.895000 0.750000 7.065000 1.320000 ;
      RECT 6.895000 1.320000 7.255000 1.650000 ;
  END
END sky130_fd_sc_hs__dlxtp_1
