* File: sky130_fd_sc_hs__o41ai_4.pex.spice
* Created: Tue Sep  1 20:19:41 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HS__O41AI_4%B1 1 3 4 6 7 9 10 12 13 15 16 17 18 20 21 22
+ 33
c67 13 0 6.95413e-20 $X=1.355 $Y=1.185
c68 7 0 6.95413e-20 $X=0.925 $Y=1.185
r69 32 34 9.58886 $w=3.77e-07 $l=7.5e-08 $layer=POLY_cond $X=0.98 $Y=1.475
+ $X2=1.055 $Y2=1.475
r70 32 33 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=0.98
+ $Y=1.385 $X2=0.98 $Y2=1.385
r71 30 32 7.03183 $w=3.77e-07 $l=5.5e-08 $layer=POLY_cond $X=0.925 $Y=1.475
+ $X2=0.98 $Y2=1.475
r72 29 30 53.6976 $w=3.77e-07 $l=4.2e-07 $layer=POLY_cond $X=0.505 $Y=1.475
+ $X2=0.925 $Y2=1.475
r73 28 29 1.27851 $w=3.77e-07 $l=1e-08 $layer=POLY_cond $X=0.495 $Y=1.475
+ $X2=0.505 $Y2=1.475
r74 26 28 24.931 $w=3.77e-07 $l=1.95e-07 $layer=POLY_cond $X=0.3 $Y=1.475
+ $X2=0.495 $Y2=1.475
r75 26 27 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=0.3
+ $Y=1.385 $X2=0.3 $Y2=1.385
r76 22 33 8.09825 $w=3.68e-07 $l=2.6e-07 $layer=LI1_cond $X=0.72 $Y=1.365
+ $X2=0.98 $Y2=1.365
r77 22 27 13.0818 $w=3.68e-07 $l=4.2e-07 $layer=LI1_cond $X=0.72 $Y=1.365
+ $X2=0.3 $Y2=1.365
r78 21 27 1.86883 $w=3.68e-07 $l=6e-08 $layer=LI1_cond $X=0.24 $Y=1.365 $X2=0.3
+ $Y2=1.365
r79 18 20 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=1.855 $Y=1.185
+ $X2=1.855 $Y2=0.74
r80 16 18 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.78 $Y=1.26
+ $X2=1.855 $Y2=1.185
r81 16 17 179.468 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=1.78 $Y=1.26
+ $X2=1.43 $Y2=1.26
r82 13 17 27.6612 $w=3.77e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.355 $Y=1.185
+ $X2=1.43 $Y2=1.26
r83 13 34 38.3554 $w=3.77e-07 $l=4.20714e-07 $layer=POLY_cond $X=1.355 $Y=1.185
+ $X2=1.055 $Y2=1.475
r84 13 15 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=1.355 $Y=1.185
+ $X2=1.355 $Y2=0.74
r85 10 34 24.4204 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=1.055 $Y=1.765
+ $X2=1.055 $Y2=1.475
r86 10 12 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.055 $Y=1.765
+ $X2=1.055 $Y2=2.4
r87 7 30 24.4204 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=0.925 $Y=1.185
+ $X2=0.925 $Y2=1.475
r88 7 9 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=0.925 $Y=1.185
+ $X2=0.925 $Y2=0.74
r89 4 29 24.4204 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=0.505 $Y=1.765
+ $X2=0.505 $Y2=1.475
r90 4 6 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.505 $Y=1.765
+ $X2=0.505 $Y2=2.4
r91 1 28 24.4204 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=0.495 $Y=1.185
+ $X2=0.495 $Y2=1.475
r92 1 3 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=0.495 $Y=1.185
+ $X2=0.495 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HS__O41AI_4%A4 1 3 4 6 7 9 10 12 13 15 16 18 19 21 22 23
+ 24 26 27 28 40
c88 24 0 3.37137e-19 $X=3.97 $Y=1.185
c89 23 0 1.72039e-20 $X=3.615 $Y=1.26
c90 22 0 7.05393e-20 $X=3.895 $Y=1.26
c91 19 0 1.95112e-19 $X=3.54 $Y=1.185
c92 4 0 1.05859e-19 $X=2.355 $Y=1.185
r93 41 42 32.5276 $w=4.89e-07 $l=3.3e-07 $layer=POLY_cond $X=3.085 $Y=1.475
+ $X2=3.415 $Y2=1.475
r94 39 41 8.87117 $w=4.89e-07 $l=9e-08 $layer=POLY_cond $X=2.995 $Y=1.475
+ $X2=3.085 $Y2=1.475
r95 39 40 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.995
+ $Y=1.385 $X2=2.995 $Y2=1.385
r96 37 39 2.95706 $w=4.89e-07 $l=3e-08 $layer=POLY_cond $X=2.965 $Y=1.475
+ $X2=2.995 $Y2=1.475
r97 36 37 44.3558 $w=4.89e-07 $l=4.5e-07 $layer=POLY_cond $X=2.515 $Y=1.475
+ $X2=2.965 $Y2=1.475
r98 35 36 15.771 $w=4.89e-07 $l=1.6e-07 $layer=POLY_cond $X=2.355 $Y=1.475
+ $X2=2.515 $Y2=1.475
r99 33 35 3.94274 $w=4.89e-07 $l=4e-08 $layer=POLY_cond $X=2.315 $Y=1.475
+ $X2=2.355 $Y2=1.475
r100 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.315
+ $Y=1.385 $X2=2.315 $Y2=1.385
r101 28 40 11.0572 $w=3.68e-07 $l=3.55e-07 $layer=LI1_cond $X=2.64 $Y=1.365
+ $X2=2.995 $Y2=1.365
r102 28 34 10.1228 $w=3.68e-07 $l=3.25e-07 $layer=LI1_cond $X=2.64 $Y=1.365
+ $X2=2.315 $Y2=1.365
r103 27 34 4.8278 $w=3.68e-07 $l=1.55e-07 $layer=LI1_cond $X=2.16 $Y=1.365
+ $X2=2.315 $Y2=1.365
r104 24 26 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=3.97 $Y=1.185
+ $X2=3.97 $Y2=0.74
r105 22 24 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.895 $Y=1.26
+ $X2=3.97 $Y2=1.185
r106 22 23 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=3.895 $Y=1.26
+ $X2=3.615 $Y2=1.26
r107 19 23 32.7723 $w=4.89e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.54 $Y=1.185
+ $X2=3.615 $Y2=1.26
r108 19 42 12.3211 $w=4.89e-07 $l=3.46915e-07 $layer=POLY_cond $X=3.54 $Y=1.185
+ $X2=3.415 $Y2=1.475
r109 19 21 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=3.54 $Y=1.185
+ $X2=3.54 $Y2=0.74
r110 16 42 30.8469 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=3.415 $Y=1.765
+ $X2=3.415 $Y2=1.475
r111 16 18 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.415 $Y=1.765
+ $X2=3.415 $Y2=2.4
r112 13 41 30.8469 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=3.085 $Y=1.185
+ $X2=3.085 $Y2=1.475
r113 13 15 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=3.085 $Y=1.185
+ $X2=3.085 $Y2=0.74
r114 10 37 30.8469 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=2.965 $Y=1.765
+ $X2=2.965 $Y2=1.475
r115 10 12 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.965 $Y=1.765
+ $X2=2.965 $Y2=2.4
r116 7 36 30.8469 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=2.515 $Y=1.765
+ $X2=2.515 $Y2=1.475
r117 7 9 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.515 $Y=1.765
+ $X2=2.515 $Y2=2.4
r118 4 35 30.8469 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=2.355 $Y=1.185
+ $X2=2.355 $Y2=1.475
r119 4 6 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=2.355 $Y=1.185
+ $X2=2.355 $Y2=0.74
r120 1 33 24.6421 $w=4.89e-07 $l=3.95727e-07 $layer=POLY_cond $X=2.065 $Y=1.765
+ $X2=2.315 $Y2=1.475
r121 1 3 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.065 $Y=1.765
+ $X2=2.065 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_HS__O41AI_4%A3 1 3 4 5 6 8 9 11 12 14 15 17 18 20 21 23
+ 24 26 27 28 29 30 44
c104 30 0 1.39749e-19 $X=6 $Y=1.295
c105 5 0 1.32046e-19 $X=3.955 $Y=1.65
r106 44 45 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.58
+ $Y=1.385 $X2=5.58 $Y2=1.385
r107 42 44 27.0179 $w=4.46e-07 $l=2.5e-07 $layer=POLY_cond $X=5.33 $Y=1.492
+ $X2=5.58 $Y2=1.492
r108 41 42 1.62108 $w=4.46e-07 $l=1.5e-08 $layer=POLY_cond $X=5.315 $Y=1.492
+ $X2=5.33 $Y2=1.492
r109 39 41 44.8498 $w=4.46e-07 $l=4.15e-07 $layer=POLY_cond $X=4.9 $Y=1.492
+ $X2=5.315 $Y2=1.492
r110 39 40 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.9
+ $Y=1.385 $X2=4.9 $Y2=1.385
r111 37 39 3.78251 $w=4.46e-07 $l=3.5e-08 $layer=POLY_cond $X=4.865 $Y=1.492
+ $X2=4.9 $Y2=1.492
r112 36 37 48.6323 $w=4.46e-07 $l=4.5e-07 $layer=POLY_cond $X=4.415 $Y=1.492
+ $X2=4.865 $Y2=1.492
r113 35 36 1.62108 $w=4.46e-07 $l=1.5e-08 $layer=POLY_cond $X=4.4 $Y=1.492
+ $X2=4.415 $Y2=1.492
r114 30 45 13.0818 $w=3.68e-07 $l=4.2e-07 $layer=LI1_cond $X=6 $Y=1.365 $X2=5.58
+ $Y2=1.365
r115 29 45 1.86883 $w=3.68e-07 $l=6e-08 $layer=LI1_cond $X=5.52 $Y=1.365
+ $X2=5.58 $Y2=1.365
r116 28 29 14.9506 $w=3.68e-07 $l=4.8e-07 $layer=LI1_cond $X=5.04 $Y=1.365
+ $X2=5.52 $Y2=1.365
r117 28 40 4.3606 $w=3.68e-07 $l=1.4e-07 $layer=LI1_cond $X=5.04 $Y=1.365
+ $X2=4.9 $Y2=1.365
r118 27 40 10.59 $w=3.68e-07 $l=3.4e-07 $layer=LI1_cond $X=4.56 $Y=1.365 $X2=4.9
+ $Y2=1.365
r119 24 44 27.0179 $w=4.46e-07 $l=3.76808e-07 $layer=POLY_cond $X=5.83 $Y=1.22
+ $X2=5.58 $Y2=1.492
r120 24 26 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=5.83 $Y=1.22
+ $X2=5.83 $Y2=0.74
r121 21 42 28.5447 $w=1.5e-07 $l=2.72e-07 $layer=POLY_cond $X=5.33 $Y=1.22
+ $X2=5.33 $Y2=1.492
r122 21 23 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=5.33 $Y=1.22
+ $X2=5.33 $Y2=0.74
r123 18 41 28.5447 $w=1.5e-07 $l=2.73e-07 $layer=POLY_cond $X=5.315 $Y=1.765
+ $X2=5.315 $Y2=1.492
r124 18 20 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=5.315 $Y=1.765
+ $X2=5.315 $Y2=2.4
r125 15 39 28.5447 $w=1.5e-07 $l=2.72e-07 $layer=POLY_cond $X=4.9 $Y=1.22
+ $X2=4.9 $Y2=1.492
r126 15 17 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=4.9 $Y=1.22 $X2=4.9
+ $Y2=0.74
r127 12 37 28.5447 $w=1.5e-07 $l=2.73e-07 $layer=POLY_cond $X=4.865 $Y=1.765
+ $X2=4.865 $Y2=1.492
r128 12 14 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=4.865 $Y=1.765
+ $X2=4.865 $Y2=2.4
r129 9 36 28.5447 $w=1.5e-07 $l=2.73e-07 $layer=POLY_cond $X=4.415 $Y=1.765
+ $X2=4.415 $Y2=1.492
r130 9 11 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=4.415 $Y=1.765
+ $X2=4.415 $Y2=2.4
r131 6 35 28.5447 $w=1.5e-07 $l=2.72e-07 $layer=POLY_cond $X=4.4 $Y=1.22 $X2=4.4
+ $Y2=1.492
r132 6 8 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=4.4 $Y=1.22 $X2=4.4
+ $Y2=0.74
r133 4 35 30.8594 $w=4.46e-07 $l=1.9187e-07 $layer=POLY_cond $X=4.325 $Y=1.65
+ $X2=4.4 $Y2=1.492
r134 4 5 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=4.325 $Y=1.65
+ $X2=3.955 $Y2=1.65
r135 1 5 26.9307 $w=1.5e-07 $l=1.53542e-07 $layer=POLY_cond $X=3.865 $Y=1.765
+ $X2=3.955 $Y2=1.65
r136 1 3 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.865 $Y=1.765
+ $X2=3.865 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_HS__O41AI_4%A2 1 3 4 6 7 9 10 12 13 15 16 18 19 21 22 24
+ 25 26 27 28 45
c95 22 0 4.41485e-20 $X=7.675 $Y=1.765
c96 16 0 6.88708e-20 $X=7.225 $Y=1.765
r97 45 46 2.25761 $w=4.27e-07 $l=2e-08 $layer=POLY_cond $X=7.655 $Y=1.492
+ $X2=7.675 $Y2=1.492
r98 43 45 11.8525 $w=4.27e-07 $l=1.05e-07 $layer=POLY_cond $X=7.55 $Y=1.492
+ $X2=7.655 $Y2=1.492
r99 43 44 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=7.55
+ $Y=1.385 $X2=7.55 $Y2=1.385
r100 41 43 36.6862 $w=4.27e-07 $l=3.25e-07 $layer=POLY_cond $X=7.225 $Y=1.492
+ $X2=7.55 $Y2=1.492
r101 40 41 3.95082 $w=4.27e-07 $l=3.5e-08 $layer=POLY_cond $X=7.19 $Y=1.492
+ $X2=7.225 $Y2=1.492
r102 39 40 46.8454 $w=4.27e-07 $l=4.15e-07 $layer=POLY_cond $X=6.775 $Y=1.492
+ $X2=7.19 $Y2=1.492
r103 38 39 1.69321 $w=4.27e-07 $l=1.5e-08 $layer=POLY_cond $X=6.76 $Y=1.492
+ $X2=6.775 $Y2=1.492
r104 36 38 25.9625 $w=4.27e-07 $l=2.3e-07 $layer=POLY_cond $X=6.53 $Y=1.492
+ $X2=6.76 $Y2=1.492
r105 36 37 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.53
+ $Y=1.385 $X2=6.53 $Y2=1.385
r106 34 36 23.1405 $w=4.27e-07 $l=2.05e-07 $layer=POLY_cond $X=6.325 $Y=1.492
+ $X2=6.53 $Y2=1.492
r107 33 34 7.33724 $w=4.27e-07 $l=6.5e-08 $layer=POLY_cond $X=6.26 $Y=1.492
+ $X2=6.325 $Y2=1.492
r108 28 44 11.5244 $w=3.68e-07 $l=3.7e-07 $layer=LI1_cond $X=7.92 $Y=1.365
+ $X2=7.55 $Y2=1.365
r109 27 44 3.42618 $w=3.68e-07 $l=1.1e-07 $layer=LI1_cond $X=7.44 $Y=1.365
+ $X2=7.55 $Y2=1.365
r110 26 27 14.9506 $w=3.68e-07 $l=4.8e-07 $layer=LI1_cond $X=6.96 $Y=1.365
+ $X2=7.44 $Y2=1.365
r111 26 37 13.3933 $w=3.68e-07 $l=4.3e-07 $layer=LI1_cond $X=6.96 $Y=1.365
+ $X2=6.53 $Y2=1.365
r112 25 37 1.55736 $w=3.68e-07 $l=5e-08 $layer=LI1_cond $X=6.48 $Y=1.365
+ $X2=6.53 $Y2=1.365
r113 22 46 27.4666 $w=1.5e-07 $l=2.73e-07 $layer=POLY_cond $X=7.675 $Y=1.765
+ $X2=7.675 $Y2=1.492
r114 22 24 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=7.675 $Y=1.765
+ $X2=7.675 $Y2=2.4
r115 19 45 27.4666 $w=1.5e-07 $l=2.72e-07 $layer=POLY_cond $X=7.655 $Y=1.22
+ $X2=7.655 $Y2=1.492
r116 19 21 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=7.655 $Y=1.22
+ $X2=7.655 $Y2=0.74
r117 16 41 27.4666 $w=1.5e-07 $l=2.73e-07 $layer=POLY_cond $X=7.225 $Y=1.765
+ $X2=7.225 $Y2=1.492
r118 16 18 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=7.225 $Y=1.765
+ $X2=7.225 $Y2=2.4
r119 13 40 27.4666 $w=1.5e-07 $l=2.72e-07 $layer=POLY_cond $X=7.19 $Y=1.22
+ $X2=7.19 $Y2=1.492
r120 13 15 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=7.19 $Y=1.22
+ $X2=7.19 $Y2=0.74
r121 10 39 27.4666 $w=1.5e-07 $l=2.73e-07 $layer=POLY_cond $X=6.775 $Y=1.765
+ $X2=6.775 $Y2=1.492
r122 10 12 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=6.775 $Y=1.765
+ $X2=6.775 $Y2=2.4
r123 7 38 27.4666 $w=1.5e-07 $l=2.72e-07 $layer=POLY_cond $X=6.76 $Y=1.22
+ $X2=6.76 $Y2=1.492
r124 7 9 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=6.76 $Y=1.22 $X2=6.76
+ $Y2=0.74
r125 4 34 27.4666 $w=1.5e-07 $l=2.73e-07 $layer=POLY_cond $X=6.325 $Y=1.765
+ $X2=6.325 $Y2=1.492
r126 4 6 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=6.325 $Y=1.765
+ $X2=6.325 $Y2=2.4
r127 1 33 27.4666 $w=1.5e-07 $l=2.72e-07 $layer=POLY_cond $X=6.26 $Y=1.22
+ $X2=6.26 $Y2=1.492
r128 1 3 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=6.26 $Y=1.22 $X2=6.26
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HS__O41AI_4%A1 1 3 4 6 7 9 10 12 13 15 16 18 19 21 22 24
+ 25 26 27 28 45
r78 45 46 1.15311 $w=4.18e-07 $l=1e-08 $layer=POLY_cond $X=9.575 $Y=1.492
+ $X2=9.585 $Y2=1.492
r79 43 45 12.1077 $w=4.18e-07 $l=1.05e-07 $layer=POLY_cond $X=9.47 $Y=1.492
+ $X2=9.575 $Y2=1.492
r80 43 44 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=9.47
+ $Y=1.385 $X2=9.47 $Y2=1.385
r81 41 43 44.3947 $w=4.18e-07 $l=3.85e-07 $layer=POLY_cond $X=9.085 $Y=1.492
+ $X2=9.47 $Y2=1.492
r82 40 41 1.15311 $w=4.18e-07 $l=1e-08 $layer=POLY_cond $X=9.075 $Y=1.492
+ $X2=9.085 $Y2=1.492
r83 38 40 32.8636 $w=4.18e-07 $l=2.85e-07 $layer=POLY_cond $X=8.79 $Y=1.492
+ $X2=9.075 $Y2=1.492
r84 38 39 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=8.79
+ $Y=1.385 $X2=8.79 $Y2=1.385
r85 36 38 15.567 $w=4.18e-07 $l=1.35e-07 $layer=POLY_cond $X=8.655 $Y=1.492
+ $X2=8.79 $Y2=1.492
r86 35 36 3.45933 $w=4.18e-07 $l=3e-08 $layer=POLY_cond $X=8.625 $Y=1.492
+ $X2=8.655 $Y2=1.492
r87 34 35 55.9258 $w=4.18e-07 $l=4.85e-07 $layer=POLY_cond $X=8.14 $Y=1.492
+ $X2=8.625 $Y2=1.492
r88 33 34 1.72967 $w=4.18e-07 $l=1.5e-08 $layer=POLY_cond $X=8.125 $Y=1.492
+ $X2=8.14 $Y2=1.492
r89 28 44 11.5244 $w=3.68e-07 $l=3.7e-07 $layer=LI1_cond $X=9.84 $Y=1.365
+ $X2=9.47 $Y2=1.365
r90 27 44 3.42618 $w=3.68e-07 $l=1.1e-07 $layer=LI1_cond $X=9.36 $Y=1.365
+ $X2=9.47 $Y2=1.365
r91 26 27 14.9506 $w=3.68e-07 $l=4.8e-07 $layer=LI1_cond $X=8.88 $Y=1.365
+ $X2=9.36 $Y2=1.365
r92 26 39 2.80324 $w=3.68e-07 $l=9e-08 $layer=LI1_cond $X=8.88 $Y=1.365 $X2=8.79
+ $Y2=1.365
r93 25 39 12.1474 $w=3.68e-07 $l=3.9e-07 $layer=LI1_cond $X=8.4 $Y=1.365
+ $X2=8.79 $Y2=1.365
r94 22 46 26.9416 $w=1.5e-07 $l=2.72e-07 $layer=POLY_cond $X=9.585 $Y=1.22
+ $X2=9.585 $Y2=1.492
r95 22 24 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=9.585 $Y=1.22
+ $X2=9.585 $Y2=0.74
r96 19 45 26.9416 $w=1.5e-07 $l=2.73e-07 $layer=POLY_cond $X=9.575 $Y=1.765
+ $X2=9.575 $Y2=1.492
r97 19 21 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=9.575 $Y=1.765
+ $X2=9.575 $Y2=2.4
r98 16 41 26.9416 $w=1.5e-07 $l=2.72e-07 $layer=POLY_cond $X=9.085 $Y=1.22
+ $X2=9.085 $Y2=1.492
r99 16 18 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=9.085 $Y=1.22
+ $X2=9.085 $Y2=0.74
r100 13 40 26.9416 $w=1.5e-07 $l=2.73e-07 $layer=POLY_cond $X=9.075 $Y=1.765
+ $X2=9.075 $Y2=1.492
r101 13 15 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=9.075 $Y=1.765
+ $X2=9.075 $Y2=2.4
r102 10 36 26.9416 $w=1.5e-07 $l=2.72e-07 $layer=POLY_cond $X=8.655 $Y=1.22
+ $X2=8.655 $Y2=1.492
r103 10 12 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=8.655 $Y=1.22
+ $X2=8.655 $Y2=0.74
r104 7 35 26.9416 $w=1.5e-07 $l=2.73e-07 $layer=POLY_cond $X=8.625 $Y=1.765
+ $X2=8.625 $Y2=1.492
r105 7 9 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=8.625 $Y=1.765
+ $X2=8.625 $Y2=2.4
r106 4 34 26.9416 $w=1.5e-07 $l=2.72e-07 $layer=POLY_cond $X=8.14 $Y=1.22
+ $X2=8.14 $Y2=1.492
r107 4 6 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=8.14 $Y=1.22 $X2=8.14
+ $Y2=0.74
r108 1 33 26.9416 $w=1.5e-07 $l=2.73e-07 $layer=POLY_cond $X=8.125 $Y=1.765
+ $X2=8.125 $Y2=1.492
r109 1 3 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=8.125 $Y=1.765
+ $X2=8.125 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_HS__O41AI_4%VPWR 1 2 3 4 13 15 21 25 29 31 33 38 46 53
+ 54 60 63 66
r107 66 67 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.36 $Y=3.33
+ $X2=9.36 $Y2=3.33
r108 63 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=3.33 $X2=8.4
+ $Y2=3.33
r109 60 61 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r110 57 58 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r111 54 67 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.84 $Y=3.33
+ $X2=9.36 $Y2=3.33
r112 53 54 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.84 $Y=3.33
+ $X2=9.84 $Y2=3.33
r113 51 66 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.515 $Y=3.33
+ $X2=9.35 $Y2=3.33
r114 51 53 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=9.515 $Y=3.33
+ $X2=9.84 $Y2=3.33
r115 50 67 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=3.33
+ $X2=9.36 $Y2=3.33
r116 50 64 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=3.33
+ $X2=8.4 $Y2=3.33
r117 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r118 47 63 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.515 $Y=3.33
+ $X2=8.35 $Y2=3.33
r119 47 49 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=8.515 $Y=3.33
+ $X2=8.88 $Y2=3.33
r120 46 66 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.185 $Y=3.33
+ $X2=9.35 $Y2=3.33
r121 46 49 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=9.185 $Y=3.33
+ $X2=8.88 $Y2=3.33
r122 45 64 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=3.33
+ $X2=8.4 $Y2=3.33
r123 44 45 1.32857 $w=1.7e-07 $l=1.19e-06 $layer=mcon $count=7 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r124 42 61 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r125 41 44 407.102 $w=1.68e-07 $l=6.24e-06 $layer=LI1_cond $X=1.68 $Y=3.33
+ $X2=7.92 $Y2=3.33
r126 41 42 1.32857 $w=1.7e-07 $l=1.19e-06 $layer=mcon $count=7 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r127 39 60 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.445 $Y=3.33
+ $X2=1.28 $Y2=3.33
r128 39 41 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=1.445 $Y=3.33
+ $X2=1.68 $Y2=3.33
r129 38 63 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.185 $Y=3.33
+ $X2=8.35 $Y2=3.33
r130 38 44 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=8.185 $Y=3.33
+ $X2=7.92 $Y2=3.33
r131 37 61 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r132 37 58 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r133 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r134 34 57 4.73185 $w=1.7e-07 $l=2.23e-07 $layer=LI1_cond $X=0.445 $Y=3.33
+ $X2=0.222 $Y2=3.33
r135 34 36 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=0.445 $Y=3.33
+ $X2=0.72 $Y2=3.33
r136 33 60 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.115 $Y=3.33
+ $X2=1.28 $Y2=3.33
r137 33 36 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=1.115 $Y=3.33
+ $X2=0.72 $Y2=3.33
r138 31 45 0.802756 $w=4.9e-07 $l=2.88e-06 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=7.92 $Y2=3.33
r139 31 42 0.936549 $w=4.9e-07 $l=3.36e-06 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=1.68 $Y2=3.33
r140 27 66 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.35 $Y=3.245
+ $X2=9.35 $Y2=3.33
r141 27 29 35.621 $w=3.28e-07 $l=1.02e-06 $layer=LI1_cond $X=9.35 $Y=3.245
+ $X2=9.35 $Y2=2.225
r142 23 63 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.35 $Y=3.245
+ $X2=8.35 $Y2=3.33
r143 23 25 35.621 $w=3.28e-07 $l=1.02e-06 $layer=LI1_cond $X=8.35 $Y=3.245
+ $X2=8.35 $Y2=2.225
r144 19 60 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.28 $Y=3.245
+ $X2=1.28 $Y2=3.33
r145 19 21 35.621 $w=3.28e-07 $l=1.02e-06 $layer=LI1_cond $X=1.28 $Y=3.245
+ $X2=1.28 $Y2=2.225
r146 15 18 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=0.28 $Y=1.985
+ $X2=0.28 $Y2=2.815
r147 13 57 3.03433 $w=3.3e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.28 $Y=3.245
+ $X2=0.222 $Y2=3.33
r148 13 18 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=0.28 $Y=3.245
+ $X2=0.28 $Y2=2.815
r149 4 29 300 $w=1.7e-07 $l=4.74579e-07 $layer=licon1_PDIFF $count=2 $X=9.15
+ $Y=1.84 $X2=9.35 $Y2=2.225
r150 3 25 300 $w=1.7e-07 $l=4.53845e-07 $layer=licon1_PDIFF $count=2 $X=8.2
+ $Y=1.84 $X2=8.35 $Y2=2.225
r151 2 21 300 $w=1.7e-07 $l=4.53845e-07 $layer=licon1_PDIFF $count=2 $X=1.13
+ $Y=1.84 $X2=1.28 $Y2=2.225
r152 1 18 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.815
r153 1 15 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HS__O41AI_4%Y 1 2 3 4 5 18 22 24 25 26 27 28 32 34 36 39
+ 45 48 49 50 54
c72 34 0 1.32046e-19 $X=3.19 $Y=2.15
c73 26 0 1.05859e-19 $X=1.64 $Y=1.01
r74 50 54 2.84726 $w=4.3e-07 $l=1.4e-07 $layer=LI1_cond $X=3.19 $Y=1.935
+ $X2=3.05 $Y2=1.935
r75 50 54 0.214408 $w=4.28e-07 $l=8e-09 $layer=LI1_cond $X=3.042 $Y=1.935
+ $X2=3.05 $Y2=1.935
r76 49 50 10.774 $w=4.28e-07 $l=4.02e-07 $layer=LI1_cond $X=2.64 $Y=1.935
+ $X2=3.042 $Y2=1.935
r77 46 49 5.62821 $w=4.28e-07 $l=2.1e-07 $layer=LI1_cond $X=2.43 $Y=1.935
+ $X2=2.64 $Y2=1.935
r78 46 48 4.87592 $w=3e-07 $l=1.4e-07 $layer=LI1_cond $X=2.43 $Y=1.935 $X2=2.29
+ $Y2=1.935
r79 39 41 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=0.71 $Y=0.8
+ $X2=0.71 $Y2=0.925
r80 34 50 4.37257 $w=2.8e-07 $l=2.15e-07 $layer=LI1_cond $X=3.19 $Y=2.15
+ $X2=3.19 $Y2=1.935
r81 34 36 17.2866 $w=2.78e-07 $l=4.2e-07 $layer=LI1_cond $X=3.19 $Y=2.15
+ $X2=3.19 $Y2=2.57
r82 30 48 1.59214 $w=2.8e-07 $l=2.15e-07 $layer=LI1_cond $X=2.29 $Y=2.15
+ $X2=2.29 $Y2=1.935
r83 30 32 17.2866 $w=2.78e-07 $l=4.2e-07 $layer=LI1_cond $X=2.29 $Y=2.15
+ $X2=2.29 $Y2=2.57
r84 29 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.805 $Y=1.805
+ $X2=1.64 $Y2=1.805
r85 28 48 4.87592 $w=3e-07 $l=1.94422e-07 $layer=LI1_cond $X=2.15 $Y=1.805
+ $X2=2.29 $Y2=1.935
r86 28 29 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=2.15 $Y=1.805
+ $X2=1.805 $Y2=1.805
r87 27 45 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.64 $Y=1.72 $X2=1.64
+ $Y2=1.805
r88 26 44 3.25678 $w=3.3e-07 $l=2.08e-07 $layer=LI1_cond $X=1.64 $Y=1.01
+ $X2=1.64 $Y2=0.802
r89 26 27 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=1.64 $Y=1.01 $X2=1.64
+ $Y2=1.72
r90 24 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.475 $Y=1.805
+ $X2=1.64 $Y2=1.805
r91 24 25 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=1.475 $Y=1.805
+ $X2=0.945 $Y2=1.805
r92 23 41 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.795 $Y=0.925
+ $X2=0.71 $Y2=0.925
r93 22 44 4.50939 $w=1.7e-07 $l=2.17991e-07 $layer=LI1_cond $X=1.475 $Y=0.925
+ $X2=1.64 $Y2=0.802
r94 22 23 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.475 $Y=0.925
+ $X2=0.795 $Y2=0.925
r95 18 20 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=0.78 $Y=1.985
+ $X2=0.78 $Y2=2.815
r96 16 25 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.78 $Y=1.89
+ $X2=0.945 $Y2=1.805
r97 16 18 3.31764 $w=3.28e-07 $l=9.5e-08 $layer=LI1_cond $X=0.78 $Y=1.89
+ $X2=0.78 $Y2=1.985
r98 5 50 600 $w=1.7e-07 $l=2.03101e-07 $layer=licon1_PDIFF $count=1 $X=3.04
+ $Y=1.84 $X2=3.19 $Y2=1.965
r99 5 36 600 $w=1.7e-07 $l=8.01499e-07 $layer=licon1_PDIFF $count=1 $X=3.04
+ $Y=1.84 $X2=3.19 $Y2=2.57
r100 4 48 600 $w=1.7e-07 $l=2.03101e-07 $layer=licon1_PDIFF $count=1 $X=2.14
+ $Y=1.84 $X2=2.29 $Y2=1.965
r101 4 32 600 $w=1.7e-07 $l=8.01499e-07 $layer=licon1_PDIFF $count=1 $X=2.14
+ $Y=1.84 $X2=2.29 $Y2=2.57
r102 3 20 400 $w=1.7e-07 $l=1.07034e-06 $layer=licon1_PDIFF $count=1 $X=0.58
+ $Y=1.84 $X2=0.78 $Y2=2.815
r103 3 18 400 $w=1.7e-07 $l=2.62678e-07 $layer=licon1_PDIFF $count=1 $X=0.58
+ $Y=1.84 $X2=0.78 $Y2=1.985
r104 2 44 182 $w=1.7e-07 $l=5.85662e-07 $layer=licon1_NDIFF $count=1 $X=1.43
+ $Y=0.37 $X2=1.64 $Y2=0.86
r105 1 39 182 $w=1.7e-07 $l=4.95076e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.37 $X2=0.71 $Y2=0.8
.ends

.subckt PM_SKY130_FD_SC_HS__O41AI_4%A_339_368# 1 2 3 4 5 18 20 21 24 26 30 34 38
+ 40 44 46 47 48
c81 30 0 1.08401e-20 $X=3.64 $Y=1.965
r82 42 44 26.5411 $w=3.28e-07 $l=7.6e-07 $layer=LI1_cond $X=5.54 $Y=2.905
+ $X2=5.54 $Y2=2.145
r83 41 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.805 $Y=2.99
+ $X2=4.64 $Y2=2.99
r84 40 42 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=5.375 $Y=2.99
+ $X2=5.54 $Y2=2.905
r85 40 41 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=5.375 $Y=2.99
+ $X2=4.805 $Y2=2.99
r86 36 48 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.64 $Y=2.905
+ $X2=4.64 $Y2=2.99
r87 36 38 26.5411 $w=3.28e-07 $l=7.6e-07 $layer=LI1_cond $X=4.64 $Y=2.905
+ $X2=4.64 $Y2=2.145
r88 35 47 8.14251 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=3.805 $Y=2.99
+ $X2=3.652 $Y2=2.99
r89 34 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.475 $Y=2.99
+ $X2=4.64 $Y2=2.99
r90 34 35 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.475 $Y=2.99
+ $X2=3.805 $Y2=2.99
r91 30 33 32.873 $w=3.03e-07 $l=8.7e-07 $layer=LI1_cond $X=3.652 $Y=1.965
+ $X2=3.652 $Y2=2.835
r92 28 47 0.649941 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=3.652 $Y=2.905
+ $X2=3.652 $Y2=2.99
r93 28 33 2.64495 $w=3.03e-07 $l=7e-08 $layer=LI1_cond $X=3.652 $Y=2.905
+ $X2=3.652 $Y2=2.835
r94 27 46 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=2.88 $Y=2.99 $X2=2.74
+ $Y2=2.99
r95 26 47 8.14251 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=3.5 $Y=2.99
+ $X2=3.652 $Y2=2.99
r96 26 27 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=3.5 $Y=2.99 $X2=2.88
+ $Y2=2.99
r97 22 46 0.375625 $w=2.8e-07 $l=8.5e-08 $layer=LI1_cond $X=2.74 $Y=2.905
+ $X2=2.74 $Y2=2.99
r98 22 24 17.2866 $w=2.78e-07 $l=4.2e-07 $layer=LI1_cond $X=2.74 $Y=2.905
+ $X2=2.74 $Y2=2.485
r99 20 46 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=2.6 $Y=2.99 $X2=2.74
+ $Y2=2.99
r100 20 21 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=2.6 $Y=2.99
+ $X2=1.98 $Y2=2.99
r101 16 21 7.55824 $w=1.7e-07 $l=1.90825e-07 $layer=LI1_cond $X=1.827 $Y=2.905
+ $X2=1.98 $Y2=2.99
r102 16 18 25.6938 $w=3.03e-07 $l=6.8e-07 $layer=LI1_cond $X=1.827 $Y=2.905
+ $X2=1.827 $Y2=2.225
r103 5 44 300 $w=1.7e-07 $l=3.72525e-07 $layer=licon1_PDIFF $count=2 $X=5.39
+ $Y=1.84 $X2=5.54 $Y2=2.145
r104 4 38 300 $w=1.7e-07 $l=3.72525e-07 $layer=licon1_PDIFF $count=2 $X=4.49
+ $Y=1.84 $X2=4.64 $Y2=2.145
r105 3 33 400 $w=1.7e-07 $l=1.06737e-06 $layer=licon1_PDIFF $count=1 $X=3.49
+ $Y=1.84 $X2=3.64 $Y2=2.835
r106 3 30 400 $w=1.7e-07 $l=2.03101e-07 $layer=licon1_PDIFF $count=1 $X=3.49
+ $Y=1.84 $X2=3.64 $Y2=1.965
r107 2 24 300 $w=1.7e-07 $l=7.16083e-07 $layer=licon1_PDIFF $count=2 $X=2.59
+ $Y=1.84 $X2=2.74 $Y2=2.485
r108 1 18 300 $w=1.7e-07 $l=4.51719e-07 $layer=licon1_PDIFF $count=2 $X=1.695
+ $Y=1.84 $X2=1.84 $Y2=2.225
.ends

.subckt PM_SKY130_FD_SC_HS__O41AI_4%A_788_368# 1 2 3 4 15 17 18 21 23 27 29 33
+ 35 36
c47 18 0 7.69031e-20 $X=4.305 $Y=1.805
r48 31 33 7.76646 $w=2.28e-07 $l=1.55e-07 $layer=LI1_cond $X=7.45 $Y=1.89
+ $X2=7.45 $Y2=2.045
r49 30 36 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=6.665 $Y=1.805
+ $X2=6.55 $Y2=1.805
r50 29 31 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=7.335 $Y=1.805
+ $X2=7.45 $Y2=1.89
r51 29 30 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=7.335 $Y=1.805
+ $X2=6.665 $Y2=1.805
r52 25 36 0.280307 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.55 $Y=1.89
+ $X2=6.55 $Y2=1.805
r53 25 27 3.75797 $w=2.28e-07 $l=7.5e-08 $layer=LI1_cond $X=6.55 $Y=1.89
+ $X2=6.55 $Y2=1.965
r54 24 35 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=5.205 $Y=1.805
+ $X2=5.09 $Y2=1.805
r55 23 36 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=6.435 $Y=1.805
+ $X2=6.55 $Y2=1.805
r56 23 24 80.246 $w=1.68e-07 $l=1.23e-06 $layer=LI1_cond $X=6.435 $Y=1.805
+ $X2=5.205 $Y2=1.805
r57 19 35 0.280307 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.09 $Y=1.89
+ $X2=5.09 $Y2=1.805
r58 19 21 3.75797 $w=2.28e-07 $l=7.5e-08 $layer=LI1_cond $X=5.09 $Y=1.89
+ $X2=5.09 $Y2=1.965
r59 17 35 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=4.975 $Y=1.805
+ $X2=5.09 $Y2=1.805
r60 17 18 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.975 $Y=1.805
+ $X2=4.305 $Y2=1.805
r61 13 18 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.14 $Y=1.89
+ $X2=4.305 $Y2=1.805
r62 13 15 5.41299 $w=3.28e-07 $l=1.55e-07 $layer=LI1_cond $X=4.14 $Y=1.89
+ $X2=4.14 $Y2=2.045
r63 4 33 300 $w=1.7e-07 $l=2.69768e-07 $layer=licon1_PDIFF $count=2 $X=7.3
+ $Y=1.84 $X2=7.45 $Y2=2.045
r64 3 27 300 $w=1.7e-07 $l=2.03101e-07 $layer=licon1_PDIFF $count=2 $X=6.4
+ $Y=1.84 $X2=6.55 $Y2=1.965
r65 2 21 300 $w=1.7e-07 $l=2.03101e-07 $layer=licon1_PDIFF $count=2 $X=4.94
+ $Y=1.84 $X2=5.09 $Y2=1.965
r66 1 15 300 $w=1.7e-07 $l=2.88141e-07 $layer=licon1_PDIFF $count=2 $X=3.94
+ $Y=1.84 $X2=4.14 $Y2=2.045
.ends

.subckt PM_SKY130_FD_SC_HS__O41AI_4%A_1191_368# 1 2 3 4 5 18 20 21 24 26 31 34
+ 35 38 42 46 50 51
c82 50 0 4.41485e-20 $X=7 $Y=2.982
c83 35 0 6.88708e-20 $X=8.015 $Y=1.805
r84 46 48 35.8081 $w=2.78e-07 $l=8.7e-07 $layer=LI1_cond $X=9.825 $Y=1.965
+ $X2=9.825 $Y2=2.835
r85 44 46 3.0869 $w=2.78e-07 $l=7.5e-08 $layer=LI1_cond $X=9.825 $Y=1.89
+ $X2=9.825 $Y2=1.965
r86 43 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.015 $Y=1.805
+ $X2=8.85 $Y2=1.805
r87 42 44 7.36005 $w=1.7e-07 $l=1.77482e-07 $layer=LI1_cond $X=9.685 $Y=1.805
+ $X2=9.825 $Y2=1.89
r88 42 43 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=9.685 $Y=1.805
+ $X2=9.015 $Y2=1.805
r89 38 40 30.3826 $w=3.28e-07 $l=8.7e-07 $layer=LI1_cond $X=8.85 $Y=1.965
+ $X2=8.85 $Y2=2.835
r90 36 51 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.85 $Y=1.89 $X2=8.85
+ $Y2=1.805
r91 36 38 2.61919 $w=3.28e-07 $l=7.5e-08 $layer=LI1_cond $X=8.85 $Y=1.89
+ $X2=8.85 $Y2=1.965
r92 34 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.685 $Y=1.805
+ $X2=8.85 $Y2=1.805
r93 34 35 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=8.685 $Y=1.805
+ $X2=8.015 $Y2=1.805
r94 31 33 35.8081 $w=2.78e-07 $l=8.7e-07 $layer=LI1_cond $X=7.875 $Y=1.965
+ $X2=7.875 $Y2=2.835
r95 29 33 2.88111 $w=2.78e-07 $l=7e-08 $layer=LI1_cond $X=7.875 $Y=2.905
+ $X2=7.875 $Y2=2.835
r96 28 35 7.36005 $w=1.7e-07 $l=1.77482e-07 $layer=LI1_cond $X=7.875 $Y=1.89
+ $X2=8.015 $Y2=1.805
r97 28 31 3.0869 $w=2.78e-07 $l=7.5e-08 $layer=LI1_cond $X=7.875 $Y=1.89
+ $X2=7.875 $Y2=1.965
r98 27 50 8.35232 $w=1.77e-07 $l=1.68953e-07 $layer=LI1_cond $X=7.165 $Y=2.99
+ $X2=7 $Y2=2.982
r99 26 29 7.36005 $w=1.7e-07 $l=1.77482e-07 $layer=LI1_cond $X=7.735 $Y=2.99
+ $X2=7.875 $Y2=2.905
r100 26 27 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=7.735 $Y=2.99
+ $X2=7.165 $Y2=2.99
r101 22 50 0.762005 $w=3.3e-07 $l=9.2e-08 $layer=LI1_cond $X=7 $Y=2.89 $X2=7
+ $Y2=2.982
r102 22 24 26.0173 $w=3.28e-07 $l=7.45e-07 $layer=LI1_cond $X=7 $Y=2.89 $X2=7
+ $Y2=2.145
r103 20 50 8.35232 $w=1.77e-07 $l=1.65e-07 $layer=LI1_cond $X=6.835 $Y=2.982
+ $X2=7 $Y2=2.982
r104 20 21 34.172 $w=1.83e-07 $l=5.7e-07 $layer=LI1_cond $X=6.835 $Y=2.982
+ $X2=6.265 $Y2=2.982
r105 16 21 7.54394 $w=1.85e-07 $l=2.05925e-07 $layer=LI1_cond $X=6.1 $Y=2.89
+ $X2=6.265 $Y2=2.982
r106 16 18 26.0173 $w=3.28e-07 $l=7.45e-07 $layer=LI1_cond $X=6.1 $Y=2.89
+ $X2=6.1 $Y2=2.145
r107 5 48 400 $w=1.7e-07 $l=1.06737e-06 $layer=licon1_PDIFF $count=1 $X=9.65
+ $Y=1.84 $X2=9.8 $Y2=2.835
r108 5 46 400 $w=1.7e-07 $l=2.03101e-07 $layer=licon1_PDIFF $count=1 $X=9.65
+ $Y=1.84 $X2=9.8 $Y2=1.965
r109 4 40 400 $w=1.7e-07 $l=1.06737e-06 $layer=licon1_PDIFF $count=1 $X=8.7
+ $Y=1.84 $X2=8.85 $Y2=2.835
r110 4 38 400 $w=1.7e-07 $l=2.03101e-07 $layer=licon1_PDIFF $count=1 $X=8.7
+ $Y=1.84 $X2=8.85 $Y2=1.965
r111 3 33 400 $w=1.7e-07 $l=1.06737e-06 $layer=licon1_PDIFF $count=1 $X=7.75
+ $Y=1.84 $X2=7.9 $Y2=2.835
r112 3 31 400 $w=1.7e-07 $l=2.03101e-07 $layer=licon1_PDIFF $count=1 $X=7.75
+ $Y=1.84 $X2=7.9 $Y2=1.965
r113 2 24 300 $w=1.7e-07 $l=3.72525e-07 $layer=licon1_PDIFF $count=2 $X=6.85
+ $Y=1.84 $X2=7 $Y2=2.145
r114 1 18 300 $w=1.7e-07 $l=3.70473e-07 $layer=licon1_PDIFF $count=2 $X=5.955
+ $Y=1.84 $X2=6.1 $Y2=2.145
.ends

.subckt PM_SKY130_FD_SC_HS__O41AI_4%A_27_74# 1 2 3 4 5 6 7 8 9 10 11 36 38 39 40
+ 45 46 47 50 53 54 55 58 61 62 66 68 72 74 78 80 84 86 90 92 94 96 98 103 104
+ 106 108 110 112 113
c190 61 0 1.95112e-19 $X=4.105 $Y=1.3
c191 53 0 1.97387e-19 $X=3.415 $Y=1.3
c192 40 0 6.95413e-20 $X=1.975 $Y=0.34
c193 38 0 6.95413e-20 $X=0.975 $Y=0.34
r194 98 101 7.33373 $w=3.28e-07 $l=2.1e-07 $layer=LI1_cond $X=1.14 $Y=0.34
+ $X2=1.14 $Y2=0.55
r195 94 115 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=9.84 $Y=0.84
+ $X2=9.84 $Y2=0.925
r196 94 96 14.9818 $w=2.48e-07 $l=3.25e-07 $layer=LI1_cond $X=9.84 $Y=0.84
+ $X2=9.84 $Y2=0.515
r197 93 113 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.035 $Y=0.925
+ $X2=8.87 $Y2=0.925
r198 92 115 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=9.715 $Y=0.925
+ $X2=9.84 $Y2=0.925
r199 92 93 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=9.715 $Y=0.925
+ $X2=9.035 $Y2=0.925
r200 88 113 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.87 $Y=0.84
+ $X2=8.87 $Y2=0.925
r201 88 90 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=8.87 $Y=0.84
+ $X2=8.87 $Y2=0.515
r202 87 112 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.035 $Y=0.925
+ $X2=7.91 $Y2=0.925
r203 86 113 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.705 $Y=0.925
+ $X2=8.87 $Y2=0.925
r204 86 87 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=8.705 $Y=0.925
+ $X2=8.035 $Y2=0.925
r205 82 112 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=7.91 $Y=0.84
+ $X2=7.91 $Y2=0.925
r206 82 84 14.9818 $w=2.48e-07 $l=3.25e-07 $layer=LI1_cond $X=7.91 $Y=0.84
+ $X2=7.91 $Y2=0.515
r207 81 110 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.06 $Y=0.925
+ $X2=6.975 $Y2=0.925
r208 80 112 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.785 $Y=0.925
+ $X2=7.91 $Y2=0.925
r209 80 81 47.2995 $w=1.68e-07 $l=7.25e-07 $layer=LI1_cond $X=7.785 $Y=0.925
+ $X2=7.06 $Y2=0.925
r210 76 110 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.975 $Y=0.84
+ $X2=6.975 $Y2=0.925
r211 76 78 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=6.975 $Y=0.84
+ $X2=6.975 $Y2=0.515
r212 75 108 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.21 $Y=0.925
+ $X2=6.085 $Y2=0.925
r213 74 110 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.89 $Y=0.925
+ $X2=6.975 $Y2=0.925
r214 74 75 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=6.89 $Y=0.925
+ $X2=6.21 $Y2=0.925
r215 70 108 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.085 $Y=0.84
+ $X2=6.085 $Y2=0.925
r216 70 72 14.9818 $w=2.48e-07 $l=3.25e-07 $layer=LI1_cond $X=6.085 $Y=0.84
+ $X2=6.085 $Y2=0.515
r217 69 106 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.28 $Y=0.925
+ $X2=5.155 $Y2=0.925
r218 68 108 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.96 $Y=0.925
+ $X2=6.085 $Y2=0.925
r219 68 69 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=5.96 $Y=0.925
+ $X2=5.28 $Y2=0.925
r220 64 106 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.155 $Y=0.84
+ $X2=5.155 $Y2=0.925
r221 64 66 14.9818 $w=2.48e-07 $l=3.25e-07 $layer=LI1_cond $X=5.155 $Y=0.84
+ $X2=5.155 $Y2=0.515
r222 63 104 2.76166 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.35 $Y=0.925
+ $X2=4.185 $Y2=0.925
r223 62 106 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.03 $Y=0.925
+ $X2=5.155 $Y2=0.925
r224 62 63 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=5.03 $Y=0.925
+ $X2=4.35 $Y2=0.925
r225 60 104 3.70735 $w=2.5e-07 $l=1.18427e-07 $layer=LI1_cond $X=4.105 $Y=1.01
+ $X2=4.185 $Y2=0.925
r226 60 61 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=4.105 $Y=1.01
+ $X2=4.105 $Y2=1.3
r227 56 104 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.185 $Y=0.84
+ $X2=4.185 $Y2=0.925
r228 56 58 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=4.185 $Y=0.84
+ $X2=4.185 $Y2=0.515
r229 54 61 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.02 $Y=1.385
+ $X2=4.105 $Y2=1.3
r230 54 55 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=4.02 $Y=1.385
+ $X2=3.5 $Y2=1.385
r231 53 55 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.415 $Y=1.3
+ $X2=3.5 $Y2=1.385
r232 52 103 3.64284 $w=2.55e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.415 $Y=1.01
+ $X2=3.33 $Y2=0.925
r233 52 53 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=3.415 $Y=1.01
+ $X2=3.415 $Y2=1.3
r234 48 103 3.64284 $w=2.55e-07 $l=8.5e-08 $layer=LI1_cond $X=3.33 $Y=0.84
+ $X2=3.33 $Y2=0.925
r235 48 50 11.016 $w=3.38e-07 $l=3.25e-07 $layer=LI1_cond $X=3.33 $Y=0.84
+ $X2=3.33 $Y2=0.515
r236 46 103 2.83584 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=3.16 $Y=0.925
+ $X2=3.33 $Y2=0.925
r237 46 47 55.7807 $w=1.68e-07 $l=8.55e-07 $layer=LI1_cond $X=3.16 $Y=0.925
+ $X2=2.305 $Y2=0.925
r238 43 47 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.14 $Y=0.84
+ $X2=2.305 $Y2=0.925
r239 43 45 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=2.14 $Y=0.84
+ $X2=2.14 $Y2=0.515
r240 42 45 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=2.14 $Y=0.425
+ $X2=2.14 $Y2=0.515
r241 41 98 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.305 $Y=0.34
+ $X2=1.14 $Y2=0.34
r242 40 42 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.975 $Y=0.34
+ $X2=2.14 $Y2=0.425
r243 40 41 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.975 $Y=0.34
+ $X2=1.305 $Y2=0.34
r244 38 98 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.975 $Y=0.34
+ $X2=1.14 $Y2=0.34
r245 38 39 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=0.975 $Y=0.34
+ $X2=0.445 $Y2=0.34
r246 34 39 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.28 $Y=0.425
+ $X2=0.445 $Y2=0.34
r247 34 36 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=0.28 $Y=0.425
+ $X2=0.28 $Y2=0.515
r248 11 115 182 $w=1.7e-07 $l=6.21068e-07 $layer=licon1_NDIFF $count=1 $X=9.66
+ $Y=0.37 $X2=9.8 $Y2=0.925
r249 11 96 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=9.66
+ $Y=0.37 $X2=9.8 $Y2=0.515
r250 10 90 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=8.73
+ $Y=0.37 $X2=8.87 $Y2=0.515
r251 9 112 182 $w=1.7e-07 $l=6.21068e-07 $layer=licon1_NDIFF $count=1 $X=7.73
+ $Y=0.37 $X2=7.87 $Y2=0.925
r252 9 84 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=7.73
+ $Y=0.37 $X2=7.87 $Y2=0.515
r253 8 110 182 $w=1.7e-07 $l=6.21068e-07 $layer=licon1_NDIFF $count=1 $X=6.835
+ $Y=0.37 $X2=6.975 $Y2=0.925
r254 8 78 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=6.835
+ $Y=0.37 $X2=6.975 $Y2=0.515
r255 7 108 182 $w=1.7e-07 $l=6.21068e-07 $layer=licon1_NDIFF $count=1 $X=5.905
+ $Y=0.37 $X2=6.045 $Y2=0.925
r256 7 72 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=5.905
+ $Y=0.37 $X2=6.045 $Y2=0.515
r257 6 106 182 $w=1.7e-07 $l=6.21068e-07 $layer=licon1_NDIFF $count=1 $X=4.975
+ $Y=0.37 $X2=5.115 $Y2=0.925
r258 6 66 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=4.975
+ $Y=0.37 $X2=5.115 $Y2=0.515
r259 5 58 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=4.045
+ $Y=0.37 $X2=4.185 $Y2=0.515
r260 4 50 91 $w=1.7e-07 $l=2.26164e-07 $layer=licon1_NDIFF $count=2 $X=3.16
+ $Y=0.37 $X2=3.325 $Y2=0.515
r261 3 45 91 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=2 $X=1.93
+ $Y=0.37 $X2=2.14 $Y2=0.515
r262 2 101 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=1 $Y=0.37
+ $X2=1.14 $Y2=0.55
r263 1 36 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__O41AI_4%VGND 1 2 3 4 5 6 7 8 27 29 33 35 39 43 47 51
+ 55 57 58 59 61 73 78 83 88 95 96 106 109 112 115 118 121
r149 121 122 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.36 $Y=0
+ $X2=9.36 $Y2=0
r150 118 119 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r151 115 116 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=0
+ $X2=7.44 $Y2=0
r152 112 113 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=0
+ $X2=6.48 $Y2=0
r153 109 110 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.52 $Y=0
+ $X2=5.52 $Y2=0
r154 106 107 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=0
+ $X2=4.56 $Y2=0
r155 96 122 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.84 $Y=0
+ $X2=9.36 $Y2=0
r156 95 96 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.84 $Y=0 $X2=9.84
+ $Y2=0
r157 93 121 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.535 $Y=0
+ $X2=9.37 $Y2=0
r158 93 95 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=9.535 $Y=0
+ $X2=9.84 $Y2=0
r159 92 122 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=0
+ $X2=9.36 $Y2=0
r160 92 119 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=0 $X2=8.4
+ $Y2=0
r161 91 92 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=0 $X2=8.88
+ $Y2=0
r162 89 118 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.535 $Y=0
+ $X2=8.37 $Y2=0
r163 89 91 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=8.535 $Y=0 $X2=8.88
+ $Y2=0
r164 88 121 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.205 $Y=0
+ $X2=9.37 $Y2=0
r165 88 91 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=9.205 $Y=0
+ $X2=8.88 $Y2=0
r166 87 119 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=0 $X2=8.4
+ $Y2=0
r167 87 116 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=0
+ $X2=7.44 $Y2=0
r168 86 87 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=0 $X2=7.92
+ $Y2=0
r169 84 115 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.57 $Y=0
+ $X2=7.405 $Y2=0
r170 84 86 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=7.57 $Y=0 $X2=7.92
+ $Y2=0
r171 83 118 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.205 $Y=0
+ $X2=8.37 $Y2=0
r172 83 86 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=8.205 $Y=0
+ $X2=7.92 $Y2=0
r173 82 116 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=0
+ $X2=7.44 $Y2=0
r174 82 113 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=0
+ $X2=6.48 $Y2=0
r175 81 82 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=0 $X2=6.96
+ $Y2=0
r176 79 112 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.71 $Y=0
+ $X2=6.545 $Y2=0
r177 79 81 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=6.71 $Y=0 $X2=6.96
+ $Y2=0
r178 78 115 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.24 $Y=0
+ $X2=7.405 $Y2=0
r179 78 81 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=7.24 $Y=0 $X2=6.96
+ $Y2=0
r180 77 113 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=0 $X2=6.48
+ $Y2=0
r181 77 110 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=0 $X2=5.52
+ $Y2=0
r182 76 77 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=0 $X2=6 $Y2=0
r183 74 109 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.78 $Y=0
+ $X2=5.615 $Y2=0
r184 74 76 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=5.78 $Y=0 $X2=6
+ $Y2=0
r185 73 112 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.38 $Y=0
+ $X2=6.545 $Y2=0
r186 73 76 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=6.38 $Y=0 $X2=6
+ $Y2=0
r187 72 107 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.56
+ $Y2=0
r188 72 101 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=2.64
+ $Y2=0
r189 71 72 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r190 69 71 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=2.99 $Y=0 $X2=3.6
+ $Y2=0
r191 68 101 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0
+ $X2=2.64 $Y2=0
r192 67 68 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.16 $Y=0
+ $X2=2.16 $Y2=0
r193 64 68 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=0.24 $Y=0
+ $X2=2.16 $Y2=0
r194 63 67 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=0.24 $Y=0 $X2=2.16
+ $Y2=0
r195 63 64 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.24 $Y=0
+ $X2=0.24 $Y2=0
r196 61 103 11.9608 $w=5.13e-07 $l=5.15e-07 $layer=LI1_cond $X=2.732 $Y=0
+ $X2=2.732 $Y2=0.515
r197 61 69 7.34265 $w=1.7e-07 $l=2.58e-07 $layer=LI1_cond $X=2.732 $Y=0 $X2=2.99
+ $Y2=0
r198 61 101 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r199 61 67 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=2.475 $Y=0
+ $X2=2.16 $Y2=0
r200 59 110 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=0
+ $X2=5.52 $Y2=0
r201 59 107 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=0
+ $X2=4.56 $Y2=0
r202 57 71 4.56684 $w=1.68e-07 $l=7e-08 $layer=LI1_cond $X=3.67 $Y=0 $X2=3.6
+ $Y2=0
r203 57 58 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.67 $Y=0 $X2=3.755
+ $Y2=0
r204 53 121 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.37 $Y=0.085
+ $X2=9.37 $Y2=0
r205 53 55 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=9.37 $Y=0.085
+ $X2=9.37 $Y2=0.55
r206 49 118 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.37 $Y=0.085
+ $X2=8.37 $Y2=0
r207 49 51 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=8.37 $Y=0.085
+ $X2=8.37 $Y2=0.55
r208 45 115 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.405 $Y=0.085
+ $X2=7.405 $Y2=0
r209 45 47 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=7.405 $Y=0.085
+ $X2=7.405 $Y2=0.55
r210 41 112 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.545 $Y=0.085
+ $X2=6.545 $Y2=0
r211 41 43 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=6.545 $Y=0.085
+ $X2=6.545 $Y2=0.55
r212 37 109 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.615 $Y=0.085
+ $X2=5.615 $Y2=0
r213 37 39 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=5.615 $Y=0.085
+ $X2=5.615 $Y2=0.55
r214 36 106 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.85 $Y=0
+ $X2=4.685 $Y2=0
r215 35 109 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.45 $Y=0
+ $X2=5.615 $Y2=0
r216 35 36 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=5.45 $Y=0 $X2=4.85
+ $Y2=0
r217 31 106 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.685 $Y=0.085
+ $X2=4.685 $Y2=0
r218 31 33 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=4.685 $Y=0.085
+ $X2=4.685 $Y2=0.55
r219 30 58 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.84 $Y=0 $X2=3.755
+ $Y2=0
r220 29 106 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.52 $Y=0
+ $X2=4.685 $Y2=0
r221 29 30 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=4.52 $Y=0 $X2=3.84
+ $Y2=0
r222 25 58 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.755 $Y=0.085
+ $X2=3.755 $Y2=0
r223 25 27 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=3.755 $Y=0.085
+ $X2=3.755 $Y2=0.515
r224 8 55 182 $w=1.7e-07 $l=2.86182e-07 $layer=licon1_NDIFF $count=1 $X=9.16
+ $Y=0.37 $X2=9.37 $Y2=0.55
r225 7 51 182 $w=1.7e-07 $l=2.45561e-07 $layer=licon1_NDIFF $count=1 $X=8.215
+ $Y=0.37 $X2=8.37 $Y2=0.55
r226 6 47 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=7.265
+ $Y=0.37 $X2=7.405 $Y2=0.55
r227 5 43 182 $w=1.7e-07 $l=2.86182e-07 $layer=licon1_NDIFF $count=1 $X=6.335
+ $Y=0.37 $X2=6.545 $Y2=0.55
r228 4 39 182 $w=1.7e-07 $l=2.86182e-07 $layer=licon1_NDIFF $count=1 $X=5.405
+ $Y=0.37 $X2=5.615 $Y2=0.55
r229 3 33 182 $w=1.7e-07 $l=2.86182e-07 $layer=licon1_NDIFF $count=1 $X=4.475
+ $Y=0.37 $X2=4.685 $Y2=0.55
r230 2 27 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.615
+ $Y=0.37 $X2=3.755 $Y2=0.515
r231 1 103 182 $w=1.7e-07 $l=3.65377e-07 $layer=licon1_NDIFF $count=1 $X=2.43
+ $Y=0.37 $X2=2.73 $Y2=0.515
.ends

