* File: sky130_fd_sc_hs__dlclkp_1.pex.spice
* Created: Tue Sep  1 20:01:21 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HS__DLCLKP_1%A_83_260# 1 2 9 11 13 14 15 16 18 19 21 23
+ 24 26 28 30
c84 11 0 1.96644e-19 $X=0.505 $Y=1.765
r85 34 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.6
+ $Y=1.465 $X2=0.6 $Y2=1.465
r86 28 30 15.1913 $w=3.28e-07 $l=4.35e-07 $layer=LI1_cond $X=1.555 $Y=2.715
+ $X2=1.99 $Y2=2.715
r87 24 26 14.8421 $w=3.28e-07 $l=4.25e-07 $layer=LI1_cond $X=1.555 $Y=0.815
+ $X2=1.98 $Y2=0.815
r88 23 28 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.47 $Y=2.55
+ $X2=1.555 $Y2=2.715
r89 22 23 26.7487 $w=1.68e-07 $l=4.1e-07 $layer=LI1_cond $X=1.47 $Y=2.14
+ $X2=1.47 $Y2=2.55
r90 20 24 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.47 $Y=0.98
+ $X2=1.555 $Y2=0.815
r91 20 21 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=1.47 $Y=0.98 $X2=1.47
+ $Y2=1.13
r92 18 22 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.385 $Y=2.055
+ $X2=1.47 $Y2=2.14
r93 18 19 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=1.385 $Y=2.055
+ $X2=0.785 $Y2=2.055
r94 17 34 10.5903 $w=2.88e-07 $l=3.2596e-07 $layer=LI1_cond $X=0.785 $Y=1.215
+ $X2=0.61 $Y2=1.465
r95 16 21 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.385 $Y=1.215
+ $X2=1.47 $Y2=1.13
r96 16 17 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=1.385 $Y=1.215
+ $X2=0.785 $Y2=1.215
r97 15 19 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.7 $Y=1.97
+ $X2=0.785 $Y2=2.055
r98 14 34 9.02084 $w=2.88e-07 $l=2.05122e-07 $layer=LI1_cond $X=0.7 $Y=1.63
+ $X2=0.61 $Y2=1.465
r99 14 15 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=0.7 $Y=1.63 $X2=0.7
+ $Y2=1.97
r100 11 35 60.2419 $w=3e-07 $l=3.39853e-07 $layer=POLY_cond $X=0.505 $Y=1.765
+ $X2=0.59 $Y2=1.465
r101 11 13 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.505 $Y=1.765
+ $X2=0.505 $Y2=2.4
r102 7 35 38.5519 $w=3e-07 $l=2.07123e-07 $layer=POLY_cond $X=0.495 $Y=1.3
+ $X2=0.59 $Y2=1.465
r103 7 9 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=0.495 $Y=1.3
+ $X2=0.495 $Y2=0.74
r104 2 30 600 $w=1.7e-07 $l=8.83982e-07 $layer=licon1_PDIFF $count=1 $X=1.71
+ $Y=1.96 $X2=1.99 $Y2=2.715
r105 1 26 182 $w=1.7e-07 $l=5.27304e-07 $layer=licon1_NDIFF $count=1 $X=1.725
+ $Y=0.4 $X2=1.98 $Y2=0.815
.ends

.subckt PM_SKY130_FD_SC_HS__DLCLKP_1%GATE 1 3 6 8
c39 8 0 2.38625e-19 $X=1.2 $Y=1.665
c40 1 0 1.10289e-19 $X=1.215 $Y=1.885
r41 8 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.17
+ $Y=1.635 $X2=1.17 $Y2=1.635
r42 4 11 38.5562 $w=2.99e-07 $l=2.05122e-07 $layer=POLY_cond $X=1.26 $Y=1.47
+ $X2=1.17 $Y2=1.635
r43 4 6 384.574 $w=1.5e-07 $l=7.5e-07 $layer=POLY_cond $X=1.26 $Y=1.47 $X2=1.26
+ $Y2=0.72
r44 1 11 52.2586 $w=2.99e-07 $l=2.7157e-07 $layer=POLY_cond $X=1.215 $Y=1.885
+ $X2=1.17 $Y2=1.635
r45 1 3 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=1.215 $Y=1.885
+ $X2=1.215 $Y2=2.46
.ends

.subckt PM_SKY130_FD_SC_HS__DLCLKP_1%A_315_54# 1 2 7 9 10 12 13 15 18 22 23 25
+ 26 31 32 36 38 41 45 48
c115 38 0 1.99284e-19 $X=4.102 $Y=2.102
c116 26 0 1.78419e-19 $X=1.995 $Y=2.215
c117 23 0 4.19812e-20 $X=1.83 $Y=1.315
c118 18 0 1.44503e-20 $X=3.335 $Y=0.995
c119 7 0 1.29101e-19 $X=1.65 $Y=1.15
r120 45 46 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.27
+ $Y=1.665 $X2=3.27 $Y2=1.665
r121 42 45 5.41299 $w=3.28e-07 $l=1.55e-07 $layer=LI1_cond $X=3.115 $Y=1.665
+ $X2=3.27 $Y2=1.665
r122 39 41 10.2439 $w=3.13e-07 $l=2.8e-07 $layer=LI1_cond $X=4.102 $Y=2.39
+ $X2=4.102 $Y2=2.11
r123 38 49 6.12936 $w=3.13e-07 $l=1.57e-07 $layer=LI1_cond $X=4.102 $Y=2.102
+ $X2=4.102 $Y2=1.945
r124 38 41 0.292684 $w=3.13e-07 $l=8e-09 $layer=LI1_cond $X=4.102 $Y=2.102
+ $X2=4.102 $Y2=2.11
r125 36 49 32.1354 $w=2.58e-07 $l=7.25e-07 $layer=LI1_cond $X=4.075 $Y=1.22
+ $X2=4.075 $Y2=1.945
r126 33 48 3.70735 $w=2.5e-07 $l=2.08207e-07 $layer=LI1_cond $X=3.2 $Y=2.475
+ $X2=3.115 $Y2=2.305
r127 32 39 7.64049 $w=1.7e-07 $l=1.94921e-07 $layer=LI1_cond $X=3.945 $Y=2.475
+ $X2=4.102 $Y2=2.39
r128 32 33 48.6043 $w=1.68e-07 $l=7.45e-07 $layer=LI1_cond $X=3.945 $Y=2.475
+ $X2=3.2 $Y2=2.475
r129 31 48 2.76166 $w=1.7e-07 $l=2.55e-07 $layer=LI1_cond $X=3.115 $Y=2.05
+ $X2=3.115 $Y2=2.305
r130 30 42 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.115 $Y=1.83
+ $X2=3.115 $Y2=1.665
r131 30 31 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=3.115 $Y=1.83
+ $X2=3.115 $Y2=2.05
r132 28 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.3
+ $Y=2.215 $X2=2.3 $Y2=2.215
r133 26 28 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=1.995 $Y=2.215
+ $X2=2.3 $Y2=2.215
r134 25 48 3.70735 $w=2.5e-07 $l=1.25499e-07 $layer=LI1_cond $X=3.03 $Y=2.215
+ $X2=3.115 $Y2=2.305
r135 25 28 25.4934 $w=3.28e-07 $l=7.3e-07 $layer=LI1_cond $X=3.03 $Y=2.215
+ $X2=2.3 $Y2=2.215
r136 23 50 31.475 $w=3.3e-07 $l=1.8e-07 $layer=POLY_cond $X=1.83 $Y=1.315
+ $X2=1.65 $Y2=1.315
r137 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.83
+ $Y=1.315 $X2=1.83 $Y2=1.315
r138 20 26 6.90553 $w=3.3e-07 $l=2.22486e-07 $layer=LI1_cond $X=1.86 $Y=2.05
+ $X2=1.995 $Y2=2.215
r139 20 22 31.3721 $w=2.68e-07 $l=7.35e-07 $layer=LI1_cond $X=1.86 $Y=2.05
+ $X2=1.86 $Y2=1.315
r140 16 46 38.5562 $w=2.99e-07 $l=1.94808e-07 $layer=POLY_cond $X=3.335 $Y=1.5
+ $X2=3.27 $Y2=1.665
r141 16 18 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=3.335 $Y=1.5
+ $X2=3.335 $Y2=0.995
r142 13 46 52.2586 $w=2.99e-07 $l=2.69258e-07 $layer=POLY_cond $X=3.31 $Y=1.915
+ $X2=3.27 $Y2=1.665
r143 13 15 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=3.31 $Y=1.915
+ $X2=3.31 $Y2=2.41
r144 10 29 52.2586 $w=2.99e-07 $l=2.7157e-07 $layer=POLY_cond $X=2.345 $Y=2.465
+ $X2=2.3 $Y2=2.215
r145 10 12 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=2.345 $Y=2.465
+ $X2=2.345 $Y2=2.75
r146 7 50 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.65 $Y=1.15
+ $X2=1.65 $Y2=1.315
r147 7 9 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=1.65 $Y=1.15 $X2=1.65
+ $Y2=0.72
r148 2 41 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=3.95
+ $Y=1.965 $X2=4.095 $Y2=2.11
r149 1 36 182 $w=1.7e-07 $l=6.65789e-07 $layer=licon1_NDIFF $count=1 $X=3.965
+ $Y=0.625 $X2=4.115 $Y2=1.22
.ends

.subckt PM_SKY130_FD_SC_HS__DLCLKP_1%A_309_338# 1 2 7 9 10 11 14 18 19 21 22 25
+ 28 32 34
c77 32 0 1.14189e-19 $X=3.69 $Y=2.135
c78 28 0 1.80935e-19 $X=3.69 $Y=2.05
c79 14 0 1.23395e-19 $X=2.31 $Y=0.83
r80 30 32 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=3.535 $Y=2.135
+ $X2=3.69 $Y2=2.135
r81 28 32 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.69 $Y=2.05
+ $X2=3.69 $Y2=2.135
r82 27 34 3.84343 $w=2.4e-07 $l=1.14782e-07 $layer=LI1_cond $X=3.69 $Y=1.33
+ $X2=3.62 $Y2=1.245
r83 27 28 46.9733 $w=1.68e-07 $l=7.2e-07 $layer=LI1_cond $X=3.69 $Y=1.33
+ $X2=3.69 $Y2=2.05
r84 23 34 3.84343 $w=2.4e-07 $l=8.5e-08 $layer=LI1_cond $X=3.62 $Y=1.16 $X2=3.62
+ $Y2=1.245
r85 23 25 14.4985 $w=3.08e-07 $l=3.9e-07 $layer=LI1_cond $X=3.62 $Y=1.16
+ $X2=3.62 $Y2=0.77
r86 21 34 2.60907 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=3.465 $Y=1.245
+ $X2=3.62 $Y2=1.245
r87 21 22 60.6738 $w=1.68e-07 $l=9.3e-07 $layer=LI1_cond $X=3.465 $Y=1.245
+ $X2=2.535 $Y2=1.245
r88 19 37 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=2.37 $Y=1.675 $X2=2.37
+ $Y2=1.765
r89 19 36 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.37 $Y=1.675
+ $X2=2.37 $Y2=1.51
r90 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.37
+ $Y=1.675 $X2=2.37 $Y2=1.675
r91 16 22 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.37 $Y=1.33
+ $X2=2.535 $Y2=1.245
r92 16 18 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=2.37 $Y=1.33
+ $X2=2.37 $Y2=1.675
r93 14 36 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=2.31 $Y=0.83
+ $X2=2.31 $Y2=1.51
r94 10 37 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.205 $Y=1.765
+ $X2=2.37 $Y2=1.765
r95 10 11 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=2.205 $Y=1.765
+ $X2=1.725 $Y2=1.765
r96 7 11 26.9307 $w=1.5e-07 $l=1.58745e-07 $layer=POLY_cond $X=1.635 $Y=1.885
+ $X2=1.725 $Y2=1.765
r97 7 9 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=1.635 $Y=1.885
+ $X2=1.635 $Y2=2.46
r98 2 30 600 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=3.385
+ $Y=1.99 $X2=3.535 $Y2=2.135
r99 1 25 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.41
+ $Y=0.625 $X2=3.55 $Y2=0.77
.ends

.subckt PM_SKY130_FD_SC_HS__DLCLKP_1%CLK 1 3 4 6 9 11 13 14 15 23
c47 23 0 1.11691e-19 $X=4.845 $Y=1.682
c48 15 0 1.36678e-19 $X=5.04 $Y=1.665
c49 11 0 1.99284e-19 $X=4.86 $Y=1.89
c50 1 0 1.80935e-19 $X=4.32 $Y=1.89
r51 23 24 1.81203 $w=3.99e-07 $l=1.5e-08 $layer=POLY_cond $X=4.845 $Y=1.682
+ $X2=4.86 $Y2=1.682
r52 21 23 10.8722 $w=3.99e-07 $l=9e-08 $layer=POLY_cond $X=4.755 $Y=1.682
+ $X2=4.845 $Y2=1.682
r53 21 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.755
+ $Y=1.64 $X2=4.755 $Y2=1.64
r54 19 21 50.7368 $w=3.99e-07 $l=4.2e-07 $layer=POLY_cond $X=4.335 $Y=1.682
+ $X2=4.755 $Y2=1.682
r55 18 19 1.81203 $w=3.99e-07 $l=1.5e-08 $layer=POLY_cond $X=4.32 $Y=1.682
+ $X2=4.335 $Y2=1.682
r56 15 22 9.95292 $w=3.28e-07 $l=2.85e-07 $layer=LI1_cond $X=5.04 $Y=1.64
+ $X2=4.755 $Y2=1.64
r57 14 22 6.80989 $w=3.28e-07 $l=1.95e-07 $layer=LI1_cond $X=4.56 $Y=1.64
+ $X2=4.755 $Y2=1.64
r58 11 24 25.8008 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=4.86 $Y=1.89
+ $X2=4.86 $Y2=1.682
r59 11 13 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=4.86 $Y=1.89
+ $X2=4.86 $Y2=2.385
r60 7 23 25.8008 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.845 $Y=1.475
+ $X2=4.845 $Y2=1.682
r61 7 9 271.766 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=4.845 $Y=1.475
+ $X2=4.845 $Y2=0.945
r62 4 19 25.8008 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.335 $Y=1.475
+ $X2=4.335 $Y2=1.682
r63 4 6 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=4.335 $Y=1.475
+ $X2=4.335 $Y2=0.995
r64 1 18 25.8008 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=4.32 $Y=1.89
+ $X2=4.32 $Y2=1.682
r65 1 3 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=4.32 $Y=1.89 $X2=4.32
+ $Y2=2.385
.ends

.subckt PM_SKY130_FD_SC_HS__DLCLKP_1%A_27_74# 1 2 10 12 13 15 18 23 25 26 28 31
+ 33 34 36 39 45 47 50 52 53 56 57 59 61 63
c140 59 0 1.37846e-19 $X=2.79 $Y=0.345
c141 56 0 1.10289e-19 $X=0.28 $Y=1.985
c142 47 0 1.29101e-19 $X=1.045 $Y=0.875
c143 36 0 1.36678e-19 $X=5.285 $Y=1.49
c144 33 0 1.14189e-19 $X=2.785 $Y=2.08
r145 60 66 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.79 $Y=0.345
+ $X2=2.79 $Y2=0.51
r146 60 63 28.8521 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.79 $Y=0.345
+ $X2=2.79 $Y2=0.18
r147 59 61 8.74048 $w=2.53e-07 $l=1.65e-07 $layer=LI1_cond $X=2.79 $Y=0.382
+ $X2=2.625 $Y2=0.382
r148 59 60 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.79
+ $Y=0.345 $X2=2.79 $Y2=0.345
r149 56 57 8.48848 $w=3.48e-07 $l=1.65e-07 $layer=LI1_cond $X=0.27 $Y=1.985
+ $X2=0.27 $Y2=1.82
r150 54 57 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=0.18 $Y=1.13
+ $X2=0.18 $Y2=1.82
r151 53 54 11.4519 $w=3.48e-07 $l=2.55e-07 $layer=LI1_cond $X=0.27 $Y=0.875
+ $X2=0.27 $Y2=1.13
r152 52 61 91.9893 $w=1.68e-07 $l=1.41e-06 $layer=LI1_cond $X=1.215 $Y=0.34
+ $X2=2.625 $Y2=0.34
r153 49 52 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.13 $Y=0.425
+ $X2=1.215 $Y2=0.34
r154 49 50 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=1.13 $Y=0.425
+ $X2=1.13 $Y2=0.79
r155 48 53 4.974 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=0.445 $Y=0.875
+ $X2=0.27 $Y2=0.875
r156 47 50 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.045 $Y=0.875
+ $X2=1.13 $Y2=0.79
r157 47 48 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=1.045 $Y=0.875
+ $X2=0.445 $Y2=0.875
r158 43 56 0.329269 $w=3.48e-07 $l=1e-08 $layer=LI1_cond $X=0.27 $Y=1.995
+ $X2=0.27 $Y2=1.985
r159 43 45 27.0001 $w=3.48e-07 $l=8.2e-07 $layer=LI1_cond $X=0.27 $Y=1.995
+ $X2=0.27 $Y2=2.815
r160 37 53 2.79879 $w=3.48e-07 $l=8.5e-08 $layer=LI1_cond $X=0.27 $Y=0.79
+ $X2=0.27 $Y2=0.875
r161 37 39 9.05491 $w=3.48e-07 $l=2.75e-07 $layer=LI1_cond $X=0.27 $Y=0.79
+ $X2=0.27 $Y2=0.515
r162 35 36 60.4563 $w=1.8e-07 $l=1.5e-07 $layer=POLY_cond $X=5.285 $Y=1.34
+ $X2=5.285 $Y2=1.49
r163 33 34 60.4563 $w=1.8e-07 $l=1.5e-07 $layer=POLY_cond $X=2.785 $Y=2.08
+ $X2=2.785 $Y2=2.23
r164 29 31 61.5319 $w=1.5e-07 $l=1.2e-07 $layer=POLY_cond $X=2.7 $Y=1.19
+ $X2=2.82 $Y2=1.19
r165 26 28 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=5.32 $Y=1.89
+ $X2=5.32 $Y2=2.385
r166 25 26 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=5.32 $Y=1.8 $X2=5.32
+ $Y2=1.89
r167 25 36 120.5 $w=1.8e-07 $l=3.1e-07 $layer=POLY_cond $X=5.32 $Y=1.8 $X2=5.32
+ $Y2=1.49
r168 23 35 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=5.235 $Y=0.945
+ $X2=5.235 $Y2=1.34
r169 20 23 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=5.235 $Y=0.255
+ $X2=5.235 $Y2=0.945
r170 19 63 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.955 $Y=0.18
+ $X2=2.79 $Y2=0.18
r171 18 20 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.16 $Y=0.18
+ $X2=5.235 $Y2=0.255
r172 18 19 1130.65 $w=1.5e-07 $l=2.205e-06 $layer=POLY_cond $X=5.16 $Y=0.18
+ $X2=2.955 $Y2=0.18
r173 16 31 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.82 $Y=1.265
+ $X2=2.82 $Y2=1.19
r174 16 33 417.904 $w=1.5e-07 $l=8.15e-07 $layer=POLY_cond $X=2.82 $Y=1.265
+ $X2=2.82 $Y2=2.08
r175 13 15 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=2.765 $Y=2.465
+ $X2=2.765 $Y2=2.75
r176 12 13 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=2.765 $Y=2.375
+ $X2=2.765 $Y2=2.465
r177 12 34 56.3629 $w=1.8e-07 $l=1.45e-07 $layer=POLY_cond $X=2.765 $Y=2.375
+ $X2=2.765 $Y2=2.23
r178 10 66 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.7 $Y=0.83 $X2=2.7
+ $Y2=0.51
r179 8 29 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.7 $Y=1.115 $X2=2.7
+ $Y2=1.19
r180 8 10 146.138 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=2.7 $Y=1.115
+ $X2=2.7 $Y2=0.83
r181 2 56 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=1.985
r182 2 45 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.815
r183 1 39 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__DLCLKP_1%A_987_393# 1 2 7 9 12 15 20 23 26 30 32 34
c64 34 0 1.11691e-19 $X=5.285 $Y=1.12
r65 30 32 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=5.095 $Y=2.06
+ $X2=5.45 $Y2=2.06
r66 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.87
+ $Y=1.465 $X2=5.87 $Y2=1.465
r67 24 34 0.364692 $w=3.3e-07 $l=4.82571e-07 $layer=LI1_cond $X=5.615 $Y=1.465
+ $X2=5.285 $Y2=1.12
r68 24 26 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=5.615 $Y=1.465
+ $X2=5.87 $Y2=1.465
r69 23 32 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.45 $Y=1.975
+ $X2=5.45 $Y2=2.06
r70 22 34 6.46576 $w=2.5e-07 $l=5.86728e-07 $layer=LI1_cond $X=5.45 $Y=1.63
+ $X2=5.285 $Y2=1.12
r71 22 23 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=5.45 $Y=1.63
+ $X2=5.45 $Y2=1.975
r72 18 34 6.46576 $w=2.5e-07 $l=1.65e-07 $layer=LI1_cond $X=5.45 $Y=1.12
+ $X2=5.285 $Y2=1.12
r73 18 20 12.2229 $w=3.28e-07 $l=3.5e-07 $layer=LI1_cond $X=5.45 $Y=1.12
+ $X2=5.45 $Y2=0.77
r74 15 27 32.3493 $w=3.3e-07 $l=1.85e-07 $layer=POLY_cond $X=6.055 $Y=1.465
+ $X2=5.87 $Y2=1.465
r75 10 15 42.8856 $w=2e-07 $l=1.8747e-07 $layer=POLY_cond $X=6.225 $Y=1.3
+ $X2=6.177 $Y2=1.465
r76 10 12 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=6.225 $Y=1.3
+ $X2=6.225 $Y2=0.74
r77 7 15 75.4206 $w=2e-07 $l=3.15595e-07 $layer=POLY_cond $X=6.145 $Y=1.765
+ $X2=6.177 $Y2=1.465
r78 7 9 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=6.145 $Y=1.765
+ $X2=6.145 $Y2=2.4
r79 2 30 300 $w=1.7e-07 $l=2.42126e-07 $layer=licon1_PDIFF $count=2 $X=4.935
+ $Y=1.965 $X2=5.095 $Y2=2.14
r80 1 20 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=5.31
+ $Y=0.625 $X2=5.45 $Y2=0.77
.ends

.subckt PM_SKY130_FD_SC_HS__DLCLKP_1%VPWR 1 2 3 4 15 19 23 27 32 33 34 36 41 49
+ 59 60 63 66 69
r83 69 70 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r84 66 67 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r85 63 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r86 59 60 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r87 57 60 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=6.48 $Y2=3.33
r88 57 70 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=4.56 $Y2=3.33
r89 56 57 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r90 54 69 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.76 $Y=3.33
+ $X2=4.595 $Y2=3.33
r91 54 56 49.5829 $w=1.68e-07 $l=7.6e-07 $layer=LI1_cond $X=4.76 $Y=3.33
+ $X2=5.52 $Y2=3.33
r92 53 70 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=4.56 $Y2=3.33
r93 52 53 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r94 50 66 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.165 $Y=3.33 $X2=3
+ $Y2=3.33
r95 50 52 59.6952 $w=1.68e-07 $l=9.15e-07 $layer=LI1_cond $X=3.165 $Y=3.33
+ $X2=4.08 $Y2=3.33
r96 49 69 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.43 $Y=3.33
+ $X2=4.595 $Y2=3.33
r97 49 52 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=4.43 $Y=3.33
+ $X2=4.08 $Y2=3.33
r98 48 67 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r99 47 48 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r100 45 48 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.64 $Y2=3.33
r101 45 64 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r102 44 47 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.2 $Y=3.33
+ $X2=2.64 $Y2=3.33
r103 44 45 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r104 42 63 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.945 $Y=3.33
+ $X2=0.78 $Y2=3.33
r105 42 44 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.945 $Y=3.33
+ $X2=1.2 $Y2=3.33
r106 41 66 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.835 $Y=3.33 $X2=3
+ $Y2=3.33
r107 41 47 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=2.835 $Y=3.33
+ $X2=2.64 $Y2=3.33
r108 39 64 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r109 38 39 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r110 36 63 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.615 $Y=3.33
+ $X2=0.78 $Y2=3.33
r111 36 38 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=0.615 $Y=3.33
+ $X2=0.24 $Y2=3.33
r112 34 53 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=3.36 $Y=3.33
+ $X2=4.08 $Y2=3.33
r113 34 67 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=3.36 $Y=3.33
+ $X2=3.12 $Y2=3.33
r114 32 56 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=5.705 $Y=3.33
+ $X2=5.52 $Y2=3.33
r115 32 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.705 $Y=3.33
+ $X2=5.87 $Y2=3.33
r116 31 59 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=6.035 $Y=3.33
+ $X2=6.48 $Y2=3.33
r117 31 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.035 $Y=3.33
+ $X2=5.87 $Y2=3.33
r118 27 30 24.6204 $w=3.28e-07 $l=7.05e-07 $layer=LI1_cond $X=5.87 $Y=2.11
+ $X2=5.87 $Y2=2.815
r119 25 33 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.87 $Y=3.245
+ $X2=5.87 $Y2=3.33
r120 25 30 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=5.87 $Y=3.245
+ $X2=5.87 $Y2=2.815
r121 21 69 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.595 $Y=3.245
+ $X2=4.595 $Y2=3.33
r122 21 23 38.5894 $w=3.28e-07 $l=1.105e-06 $layer=LI1_cond $X=4.595 $Y=3.245
+ $X2=4.595 $Y2=2.14
r123 17 66 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3 $Y=3.245 $X2=3
+ $Y2=3.33
r124 17 19 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=3 $Y=3.245 $X2=3
+ $Y2=2.815
r125 13 63 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.78 $Y=3.245
+ $X2=0.78 $Y2=3.33
r126 13 15 26.8903 $w=3.28e-07 $l=7.7e-07 $layer=LI1_cond $X=0.78 $Y=3.245
+ $X2=0.78 $Y2=2.475
r127 4 30 600 $w=1.7e-07 $l=1.06125e-06 $layer=licon1_PDIFF $count=1 $X=5.395
+ $Y=1.965 $X2=5.87 $Y2=2.815
r128 4 27 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=5.395
+ $Y=1.965 $X2=5.87 $Y2=2.11
r129 3 23 300 $w=1.7e-07 $l=2.73861e-07 $layer=licon1_PDIFF $count=2 $X=4.395
+ $Y=1.965 $X2=4.595 $Y2=2.14
r130 2 19 600 $w=1.7e-07 $l=3.45868e-07 $layer=licon1_PDIFF $count=1 $X=2.84
+ $Y=2.54 $X2=3 $Y2=2.815
r131 1 15 300 $w=1.7e-07 $l=7.28166e-07 $layer=licon1_PDIFF $count=2 $X=0.58
+ $Y=1.84 $X2=0.78 $Y2=2.475
.ends

.subckt PM_SKY130_FD_SC_HS__DLCLKP_1%GCLK 1 2 9 11 12 13 14 22
r18 14 31 1.15244 $w=3.98e-07 $l=4e-08 $layer=LI1_cond $X=6.405 $Y=2.775
+ $X2=6.405 $Y2=2.815
r19 13 14 10.6601 $w=3.98e-07 $l=3.7e-07 $layer=LI1_cond $X=6.405 $Y=2.405
+ $X2=6.405 $Y2=2.775
r20 12 13 10.6601 $w=3.98e-07 $l=3.7e-07 $layer=LI1_cond $X=6.405 $Y=2.035
+ $X2=6.405 $Y2=2.405
r21 12 22 1.44055 $w=3.98e-07 $l=5e-08 $layer=LI1_cond $X=6.405 $Y=2.035
+ $X2=6.405 $Y2=1.985
r22 11 34 3.70031 $w=3.98e-07 $l=1.15e-07 $layer=LI1_cond $X=6.405 $Y=1.665
+ $X2=6.405 $Y2=1.55
r23 11 22 6.00917 $w=5.68e-07 $l=2.35e-07 $layer=LI1_cond $X=6.405 $Y=1.75
+ $X2=6.405 $Y2=1.985
r24 9 34 36.1448 $w=3.28e-07 $l=1.035e-06 $layer=LI1_cond $X=6.44 $Y=0.515
+ $X2=6.44 $Y2=1.55
r25 2 31 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=6.22
+ $Y=1.84 $X2=6.37 $Y2=2.815
r26 2 22 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=6.22
+ $Y=1.84 $X2=6.37 $Y2=1.985
r27 1 9 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=6.3 $Y=0.37
+ $X2=6.44 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__DLCLKP_1%VGND 1 2 3 4 15 17 22 25 29 32 33 34 36 48
+ 52 59 60 63 66 69
r83 69 70 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=0 $X2=6 $Y2=0
r84 66 67 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r85 63 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r86 60 70 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=0 $X2=6
+ $Y2=0
r87 59 60 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=0 $X2=6.48
+ $Y2=0
r88 57 69 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.095 $Y=0 $X2=5.97
+ $Y2=0
r89 57 59 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=6.095 $Y=0 $X2=6.48
+ $Y2=0
r90 56 70 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=6
+ $Y2=0
r91 56 67 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=4.56
+ $Y2=0
r92 55 56 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r93 53 66 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.715 $Y=0 $X2=4.55
+ $Y2=0
r94 53 55 52.5187 $w=1.68e-07 $l=8.05e-07 $layer=LI1_cond $X=4.715 $Y=0 $X2=5.52
+ $Y2=0
r95 52 69 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.845 $Y=0 $X2=5.97
+ $Y2=0
r96 52 55 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=5.845 $Y=0 $X2=5.52
+ $Y2=0
r97 51 67 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=4.56
+ $Y2=0
r98 50 51 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r99 48 66 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.385 $Y=0 $X2=4.55
+ $Y2=0
r100 48 50 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=4.385 $Y=0
+ $X2=4.08 $Y2=0
r101 46 47 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.12 $Y=0
+ $X2=3.12 $Y2=0
r102 44 47 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=1.2 $Y=0 $X2=3.12
+ $Y2=0
r103 44 64 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r104 43 46 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=1.2 $Y=0 $X2=3.12
+ $Y2=0
r105 43 44 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r106 41 63 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.875 $Y=0 $X2=0.75
+ $Y2=0
r107 41 43 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.875 $Y=0 $X2=1.2
+ $Y2=0
r108 39 64 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r109 38 39 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r110 36 63 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.625 $Y=0 $X2=0.75
+ $Y2=0
r111 36 38 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=0.625 $Y=0
+ $X2=0.24 $Y2=0
r112 34 51 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=3.36 $Y=0 $X2=4.08
+ $Y2=0
r113 34 47 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=3.36 $Y=0
+ $X2=3.12 $Y2=0
r114 32 46 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=3.125 $Y=0 $X2=3.12
+ $Y2=0
r115 32 33 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.125 $Y=0 $X2=3.21
+ $Y2=0
r116 31 50 51.2139 $w=1.68e-07 $l=7.85e-07 $layer=LI1_cond $X=3.295 $Y=0
+ $X2=4.08 $Y2=0
r117 31 33 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.295 $Y=0 $X2=3.21
+ $Y2=0
r118 27 69 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.97 $Y=0.085
+ $X2=5.97 $Y2=0
r119 27 29 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=5.97 $Y=0.085
+ $X2=5.97 $Y2=0.515
r120 23 66 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.55 $Y=0.085
+ $X2=4.55 $Y2=0
r121 23 25 23.9219 $w=3.28e-07 $l=6.85e-07 $layer=LI1_cond $X=4.55 $Y=0.085
+ $X2=4.55 $Y2=0.77
r122 21 33 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.21 $Y=0.085
+ $X2=3.21 $Y2=0
r123 21 22 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=3.21 $Y=0.085
+ $X2=3.21 $Y2=0.685
r124 17 22 7.14316 $w=2.5e-07 $l=1.62019e-07 $layer=LI1_cond $X=3.125 $Y=0.81
+ $X2=3.21 $Y2=0.685
r125 17 19 5.07075 $w=2.48e-07 $l=1.1e-07 $layer=LI1_cond $X=3.125 $Y=0.81
+ $X2=3.015 $Y2=0.81
r126 13 63 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.75 $Y=0.085
+ $X2=0.75 $Y2=0
r127 13 15 17.0562 $w=2.48e-07 $l=3.7e-07 $layer=LI1_cond $X=0.75 $Y=0.085
+ $X2=0.75 $Y2=0.455
r128 4 29 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=5.865
+ $Y=0.37 $X2=6.01 $Y2=0.515
r129 3 25 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=4.41
+ $Y=0.625 $X2=4.55 $Y2=0.77
r130 2 19 182 $w=1.7e-07 $l=3.05941e-07 $layer=licon1_NDIFF $count=1 $X=2.775
+ $Y=0.62 $X2=3.015 $Y2=0.77
r131 1 15 182 $w=1.7e-07 $l=2.59037e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.37 $X2=0.79 $Y2=0.455
.ends

