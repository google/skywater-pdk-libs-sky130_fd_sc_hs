# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_hs__edfxbp_1
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_hs__edfxbp_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  14.40000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425000 0.980000 0.835000 1.990000 ;
    END
  END D
  PIN DE
    ANTENNAGATEAREA  0.285000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.565000 1.450000 1.905000 1.780000 ;
    END
  END DE
  PIN Q
    ANTENNADIFFAREA  0.541300 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 12.765000 0.620000 13.095000 1.000000 ;
        RECT 12.925000 1.000000 13.095000 1.820000 ;
        RECT 12.925000 1.820000 13.340000 2.980000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.541300 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 13.955000 0.370000 14.315000 1.150000 ;
        RECT 13.990000 1.820000 14.315000 2.980000 ;
        RECT 14.145000 1.150000 14.315000 1.820000 ;
    END
  END Q_N
  PIN CLK
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 3.715000 1.180000 4.385000 1.550000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT  0.000000 -0.085000 14.400000 0.085000 ;
        RECT  1.090000  0.085000  1.420000 0.810000 ;
        RECT  2.170000  0.085000  2.500000 0.810000 ;
        RECT  3.715000  0.085000  3.885000 1.010000 ;
        RECT  4.585000  0.085000  4.915000 0.670000 ;
        RECT  7.220000  0.085000  7.470000 0.795000 ;
        RECT  8.660000  0.085000  8.910000 0.770000 ;
        RECT 11.655000  0.085000 11.985000 0.985000 ;
        RECT 13.605000  0.085000 13.775000 1.150000 ;
      LAYER mcon ;
        RECT  0.155000 -0.085000  0.325000 0.085000 ;
        RECT  0.635000 -0.085000  0.805000 0.085000 ;
        RECT  1.115000 -0.085000  1.285000 0.085000 ;
        RECT  1.595000 -0.085000  1.765000 0.085000 ;
        RECT  2.075000 -0.085000  2.245000 0.085000 ;
        RECT  2.555000 -0.085000  2.725000 0.085000 ;
        RECT  3.035000 -0.085000  3.205000 0.085000 ;
        RECT  3.515000 -0.085000  3.685000 0.085000 ;
        RECT  3.995000 -0.085000  4.165000 0.085000 ;
        RECT  4.475000 -0.085000  4.645000 0.085000 ;
        RECT  4.955000 -0.085000  5.125000 0.085000 ;
        RECT  5.435000 -0.085000  5.605000 0.085000 ;
        RECT  5.915000 -0.085000  6.085000 0.085000 ;
        RECT  6.395000 -0.085000  6.565000 0.085000 ;
        RECT  6.875000 -0.085000  7.045000 0.085000 ;
        RECT  7.355000 -0.085000  7.525000 0.085000 ;
        RECT  7.835000 -0.085000  8.005000 0.085000 ;
        RECT  8.315000 -0.085000  8.485000 0.085000 ;
        RECT  8.795000 -0.085000  8.965000 0.085000 ;
        RECT  9.275000 -0.085000  9.445000 0.085000 ;
        RECT  9.755000 -0.085000  9.925000 0.085000 ;
        RECT 10.235000 -0.085000 10.405000 0.085000 ;
        RECT 10.715000 -0.085000 10.885000 0.085000 ;
        RECT 11.195000 -0.085000 11.365000 0.085000 ;
        RECT 11.675000 -0.085000 11.845000 0.085000 ;
        RECT 12.155000 -0.085000 12.325000 0.085000 ;
        RECT 12.635000 -0.085000 12.805000 0.085000 ;
        RECT 13.115000 -0.085000 13.285000 0.085000 ;
        RECT 13.595000 -0.085000 13.765000 0.085000 ;
        RECT 14.075000 -0.085000 14.245000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.245000 14.400000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT  0.000000 3.245000 14.400000 3.415000 ;
        RECT  0.955000 2.630000  1.205000 3.245000 ;
        RECT  2.395000 2.630000  2.645000 3.245000 ;
        RECT  3.715000 2.650000  4.045000 3.245000 ;
        RECT  5.105000 2.650000  5.435000 3.245000 ;
        RECT  7.695000 2.885000  8.025000 3.245000 ;
        RECT  9.575000 1.960000  9.905000 3.245000 ;
        RECT 11.495000 2.325000 12.280000 3.245000 ;
        RECT 13.540000 1.820000 13.790000 3.245000 ;
      LAYER mcon ;
        RECT  0.155000 3.245000  0.325000 3.415000 ;
        RECT  0.635000 3.245000  0.805000 3.415000 ;
        RECT  1.115000 3.245000  1.285000 3.415000 ;
        RECT  1.595000 3.245000  1.765000 3.415000 ;
        RECT  2.075000 3.245000  2.245000 3.415000 ;
        RECT  2.555000 3.245000  2.725000 3.415000 ;
        RECT  3.035000 3.245000  3.205000 3.415000 ;
        RECT  3.515000 3.245000  3.685000 3.415000 ;
        RECT  3.995000 3.245000  4.165000 3.415000 ;
        RECT  4.475000 3.245000  4.645000 3.415000 ;
        RECT  4.955000 3.245000  5.125000 3.415000 ;
        RECT  5.435000 3.245000  5.605000 3.415000 ;
        RECT  5.915000 3.245000  6.085000 3.415000 ;
        RECT  6.395000 3.245000  6.565000 3.415000 ;
        RECT  6.875000 3.245000  7.045000 3.415000 ;
        RECT  7.355000 3.245000  7.525000 3.415000 ;
        RECT  7.835000 3.245000  8.005000 3.415000 ;
        RECT  8.315000 3.245000  8.485000 3.415000 ;
        RECT  8.795000 3.245000  8.965000 3.415000 ;
        RECT  9.275000 3.245000  9.445000 3.415000 ;
        RECT  9.755000 3.245000  9.925000 3.415000 ;
        RECT 10.235000 3.245000 10.405000 3.415000 ;
        RECT 10.715000 3.245000 10.885000 3.415000 ;
        RECT 11.195000 3.245000 11.365000 3.415000 ;
        RECT 11.675000 3.245000 11.845000 3.415000 ;
        RECT 12.155000 3.245000 12.325000 3.415000 ;
        RECT 12.635000 3.245000 12.805000 3.415000 ;
        RECT 13.115000 3.245000 13.285000 3.415000 ;
        RECT 13.595000 3.245000 13.765000 3.415000 ;
        RECT 14.075000 3.245000 14.245000 3.415000 ;
      LAYER met1 ;
        RECT 0.000000 3.085000 14.400000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.085000 0.420000  0.600000 0.750000 ;
      RECT  0.085000 0.750000  0.255000 2.290000 ;
      RECT  0.085000 2.290000  1.545000 2.460000 ;
      RECT  0.085000 2.460000  0.445000 2.980000 ;
      RECT  1.005000 1.110000  2.000000 1.280000 ;
      RECT  1.005000 1.280000  1.335000 1.950000 ;
      RECT  1.005000 1.950000  2.665000 2.120000 ;
      RECT  1.375000 2.460000  1.545000 2.905000 ;
      RECT  1.375000 2.905000  2.225000 3.075000 ;
      RECT  1.650000 0.480000  2.000000 1.110000 ;
      RECT  1.715000 2.120000  1.885000 2.735000 ;
      RECT  2.055000 2.290000  3.545000 2.310000 ;
      RECT  2.055000 2.310000  5.775000 2.460000 ;
      RECT  2.055000 2.460000  2.225000 2.905000 ;
      RECT  2.335000 0.980000  2.665000 1.950000 ;
      RECT  2.875000 0.980000  3.205000 1.990000 ;
      RECT  3.000000 0.350000  3.545000 0.810000 ;
      RECT  3.155000 2.460000  5.775000 2.480000 ;
      RECT  3.155000 2.480000  3.545000 2.960000 ;
      RECT  3.375000 0.810000  3.545000 2.290000 ;
      RECT  4.065000 0.350000  4.395000 0.840000 ;
      RECT  4.065000 0.840000  4.725000 1.010000 ;
      RECT  4.165000 1.810000  4.965000 2.140000 ;
      RECT  4.555000 1.010000  4.725000 1.810000 ;
      RECT  5.095000 0.255000  6.885000 0.425000 ;
      RECT  5.095000 0.425000  5.345000 1.130000 ;
      RECT  5.215000 1.300000  5.785000 1.470000 ;
      RECT  5.215000 1.470000  5.385000 2.310000 ;
      RECT  5.535000 0.595000  5.785000 1.300000 ;
      RECT  5.555000 1.810000  6.125000 1.970000 ;
      RECT  5.555000 1.970000  6.355000 2.140000 ;
      RECT  5.605000 2.480000  5.775000 2.890000 ;
      RECT  5.605000 2.890000  6.445000 3.060000 ;
      RECT  5.955000 0.425000  6.125000 1.810000 ;
      RECT  5.955000 2.140000  6.355000 2.380000 ;
      RECT  6.295000 0.595000  6.465000 1.515000 ;
      RECT  6.295000 1.515000  6.720000 1.685000 ;
      RECT  6.550000 1.685000  6.720000 1.740000 ;
      RECT  6.550000 1.740000  8.260000 1.910000 ;
      RECT  6.550000 1.910000  6.720000 2.550000 ;
      RECT  6.550000 2.550000  6.980000 2.720000 ;
      RECT  6.635000 0.425000  6.885000 0.965000 ;
      RECT  6.635000 0.965000  7.810000 1.135000 ;
      RECT  6.635000 1.135000  6.885000 1.345000 ;
      RECT  6.650000 2.720000  6.980000 2.980000 ;
      RECT  6.890000 2.080000  7.320000 2.380000 ;
      RECT  7.150000 2.380000  7.320000 2.545000 ;
      RECT  7.150000 2.545000  8.365000 2.715000 ;
      RECT  7.205000 1.305000  9.030000 1.475000 ;
      RECT  7.205000 1.475000  7.535000 1.570000 ;
      RECT  7.640000 0.255000  8.490000 0.425000 ;
      RECT  7.640000 0.425000  7.810000 0.965000 ;
      RECT  7.930000 1.645000  8.260000 1.740000 ;
      RECT  7.930000 1.910000  8.260000 1.955000 ;
      RECT  7.980000 0.595000  8.150000 1.305000 ;
      RECT  8.195000 2.715000  8.365000 2.755000 ;
      RECT  8.195000 2.755000  9.405000 2.925000 ;
      RECT  8.230000 2.125000  9.030000 2.375000 ;
      RECT  8.320000 0.425000  8.490000 0.965000 ;
      RECT  8.320000 0.965000  9.370000 1.120000 ;
      RECT  8.320000 1.120000 11.105000 1.135000 ;
      RECT  8.700000 1.475000  9.030000 2.125000 ;
      RECT  8.700000 2.375000  9.030000 2.585000 ;
      RECT  9.200000 1.135000 11.105000 1.290000 ;
      RECT  9.200000 1.290000 10.085000 1.450000 ;
      RECT  9.235000 1.620000 10.625000 1.790000 ;
      RECT  9.235000 1.790000  9.405000 2.755000 ;
      RECT  9.540000 0.620000 11.445000 0.950000 ;
      RECT 10.295000 1.460000 10.625000 1.620000 ;
      RECT 10.445000 1.985000 11.445000 2.155000 ;
      RECT 10.445000 2.155000 10.775000 2.980000 ;
      RECT 10.835000 1.290000 11.105000 1.800000 ;
      RECT 11.275000 0.950000 11.445000 1.155000 ;
      RECT 11.275000 1.155000 11.985000 1.485000 ;
      RECT 11.275000 1.485000 11.445000 1.985000 ;
      RECT 11.615000 1.725000 12.485000 1.805000 ;
      RECT 11.615000 1.805000 12.700000 2.120000 ;
      RECT 12.155000 0.255000 13.435000 0.425000 ;
      RECT 12.155000 0.425000 12.485000 1.725000 ;
      RECT 12.450000 2.120000 12.700000 2.845000 ;
      RECT 13.265000 0.425000 13.435000 1.320000 ;
      RECT 13.265000 1.320000 13.975000 1.650000 ;
    LAYER mcon ;
      RECT  3.035000 1.580000  3.205000 1.750000 ;
      RECT 12.155000 1.580000 12.325000 1.750000 ;
    LAYER met1 ;
      RECT  2.975000 1.550000  3.265000 1.595000 ;
      RECT  2.975000 1.595000 12.385000 1.735000 ;
      RECT  2.975000 1.735000  3.265000 1.780000 ;
      RECT 12.095000 1.550000 12.385000 1.595000 ;
      RECT 12.095000 1.735000 12.385000 1.780000 ;
  END
END sky130_fd_sc_hs__edfxbp_1
