# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_hs__a222oi_2
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_hs__a222oi_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  6.720000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.685000 1.450000 5.115000 1.780000 ;
        RECT 4.945000 1.780000 5.115000 1.950000 ;
        RECT 4.945000 1.950000 6.055000 2.120000 ;
        RECT 5.885000 1.450000 6.455000 1.780000 ;
        RECT 5.885000 1.780000 6.055000 1.950000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.305000 1.450000 5.635000 1.780000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.675000 1.470000 3.235000 1.800000 ;
        RECT 3.065000 1.800000 3.235000 1.950000 ;
        RECT 3.065000 1.950000 4.275000 2.120000 ;
        RECT 4.105000 1.450000 4.475000 1.780000 ;
        RECT 4.105000 1.780000 4.275000 1.950000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.405000 1.260000 3.735000 1.780000 ;
    END
  END B2
  PIN C1
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.005000 1.165000 1.335000 1.495000 ;
    END
  END C1
  PIN C2
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425000 1.165000 0.835000 1.495000 ;
        RECT 0.605000 1.495000 0.835000 1.665000 ;
        RECT 0.605000 1.665000 2.125000 1.835000 ;
        RECT 1.795000 1.130000 2.125000 1.665000 ;
    END
  END C2
  PIN Y
    ANTENNADIFFAREA  1.693200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.825000 1.420000 0.995000 ;
        RECT 0.085000 0.995000 0.255000 1.920000 ;
        RECT 0.085000 1.920000 0.365000 2.005000 ;
        RECT 0.085000 2.005000 2.465000 2.175000 ;
        RECT 0.085000 2.175000 0.365000 2.980000 ;
        RECT 1.065000 2.175000 1.325000 2.735000 ;
        RECT 1.090000 0.780000 1.420000 0.825000 ;
        RECT 1.995000 2.175000 2.465000 2.735000 ;
        RECT 2.295000 1.130000 2.840000 1.300000 ;
        RECT 2.295000 1.300000 2.465000 2.005000 ;
        RECT 2.510000 0.350000 2.840000 0.920000 ;
        RECT 2.510000 0.920000 4.715000 1.090000 ;
        RECT 2.510000 1.090000 2.840000 1.130000 ;
        RECT 4.450000 0.350000 4.715000 0.920000 ;
        RECT 4.450000 1.090000 4.715000 1.110000 ;
        RECT 4.450000 1.110000 6.580000 1.280000 ;
        RECT 6.320000 0.350000 6.580000 1.110000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 6.720000 0.085000 ;
        RECT 0.115000  0.085000 0.480000 0.655000 ;
        RECT 1.950000  0.085000 2.280000 0.940000 ;
        RECT 3.450000  0.085000 3.840000 0.410000 ;
        RECT 5.385000  0.085000 5.715000 0.600000 ;
      LAYER mcon ;
        RECT 0.155000 -0.085000 0.325000 0.085000 ;
        RECT 0.635000 -0.085000 0.805000 0.085000 ;
        RECT 1.115000 -0.085000 1.285000 0.085000 ;
        RECT 1.595000 -0.085000 1.765000 0.085000 ;
        RECT 2.075000 -0.085000 2.245000 0.085000 ;
        RECT 2.555000 -0.085000 2.725000 0.085000 ;
        RECT 3.035000 -0.085000 3.205000 0.085000 ;
        RECT 3.515000 -0.085000 3.685000 0.085000 ;
        RECT 3.995000 -0.085000 4.165000 0.085000 ;
        RECT 4.475000 -0.085000 4.645000 0.085000 ;
        RECT 4.955000 -0.085000 5.125000 0.085000 ;
        RECT 5.435000 -0.085000 5.605000 0.085000 ;
        RECT 5.915000 -0.085000 6.085000 0.085000 ;
        RECT 6.395000 -0.085000 6.565000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.245000 6.720000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 3.245000 6.720000 3.415000 ;
        RECT 4.895000 2.650000 5.255000 3.245000 ;
        RECT 5.825000 2.650000 6.155000 3.245000 ;
      LAYER mcon ;
        RECT 0.155000 3.245000 0.325000 3.415000 ;
        RECT 0.635000 3.245000 0.805000 3.415000 ;
        RECT 1.115000 3.245000 1.285000 3.415000 ;
        RECT 1.595000 3.245000 1.765000 3.415000 ;
        RECT 2.075000 3.245000 2.245000 3.415000 ;
        RECT 2.555000 3.245000 2.725000 3.415000 ;
        RECT 3.035000 3.245000 3.205000 3.415000 ;
        RECT 3.515000 3.245000 3.685000 3.415000 ;
        RECT 3.995000 3.245000 4.165000 3.415000 ;
        RECT 4.475000 3.245000 4.645000 3.415000 ;
        RECT 4.955000 3.245000 5.125000 3.415000 ;
        RECT 5.435000 3.245000 5.605000 3.415000 ;
        RECT 5.915000 3.245000 6.085000 3.415000 ;
        RECT 6.395000 3.245000 6.565000 3.415000 ;
      LAYER met1 ;
        RECT 0.000000 3.085000 6.720000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.565000 2.345000 0.895000 2.905000 ;
      RECT 0.565000 2.905000 4.325000 2.980000 ;
      RECT 0.565000 2.980000 3.335000 3.075000 ;
      RECT 0.660000 0.350000 1.780000 0.610000 ;
      RECT 1.495000 2.345000 1.825000 2.905000 ;
      RECT 1.590000 0.610000 1.780000 0.885000 ;
      RECT 2.635000 1.970000 2.805000 2.290000 ;
      RECT 2.635000 2.290000 6.605000 2.460000 ;
      RECT 2.635000 2.460000 2.805000 2.735000 ;
      RECT 3.005000 2.630000 3.335000 2.650000 ;
      RECT 3.005000 2.650000 4.325000 2.905000 ;
      RECT 3.020000 0.350000 3.270000 0.580000 ;
      RECT 3.020000 0.580000 4.270000 0.750000 ;
      RECT 4.020000 0.350000 4.270000 0.580000 ;
      RECT 4.445000 1.950000 4.775000 2.290000 ;
      RECT 4.500000 2.460000 6.605000 2.480000 ;
      RECT 4.500000 2.480000 4.715000 2.980000 ;
      RECT 4.885000 0.350000 5.215000 0.770000 ;
      RECT 4.885000 0.770000 6.150000 0.940000 ;
      RECT 5.425000 2.480000 5.655000 2.980000 ;
      RECT 5.900000 0.330000 6.150000 0.770000 ;
      RECT 6.275000 1.950000 6.605000 2.290000 ;
      RECT 6.335000 2.480000 6.605000 3.000000 ;
  END
END sky130_fd_sc_hs__a222oi_2
