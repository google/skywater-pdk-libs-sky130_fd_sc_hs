* File: sky130_fd_sc_hs__sdfxbp_1.pex.spice
* Created: Tue Sep  1 20:23:29 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HS__SDFXBP_1%A_31_74# 1 2 9 11 13 14 16 19 21 22 24 33
c84 22 0 1.68868e-19 $X=0.915 $Y=2.04
r85 33 36 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=2.005 $Y=1.96 $X2=2.005
+ $Y2=2.04
r86 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.005
+ $Y=1.96 $X2=2.005 $Y2=1.96
r87 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.75
+ $Y=1.69 $X2=0.75 $Y2=1.69
r88 24 26 10.2392 $w=3.78e-07 $l=2.2e-07 $layer=LI1_cond $X=0.275 $Y=0.565
+ $X2=0.275 $Y2=0.785
r89 22 30 9.09243 $w=3.85e-07 $l=2.85832e-07 $layer=LI1_cond $X=0.915 $Y=2.04
+ $X2=0.75 $Y2=1.825
r90 21 36 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.84 $Y=2.04
+ $X2=2.005 $Y2=2.04
r91 21 22 60.3476 $w=1.68e-07 $l=9.25e-07 $layer=LI1_cond $X=1.84 $Y=2.04
+ $X2=0.915 $Y2=2.04
r92 17 30 14.0379 $w=3.85e-07 $l=4.43e-07 $layer=LI1_cond $X=0.307 $Y=1.825
+ $X2=0.75 $Y2=1.825
r93 17 27 4.3413 $w=3.85e-07 $l=1.37e-07 $layer=LI1_cond $X=0.307 $Y=1.825
+ $X2=0.17 $Y2=1.825
r94 17 19 15.7975 $w=4.43e-07 $l=6.1e-07 $layer=LI1_cond $X=0.307 $Y=1.855
+ $X2=0.307 $Y2=2.465
r95 16 27 5.54671 $w=1.7e-07 $l=3e-07 $layer=LI1_cond $X=0.17 $Y=1.525 $X2=0.17
+ $Y2=1.825
r96 16 26 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=0.17 $Y=1.525
+ $X2=0.17 $Y2=0.785
r97 14 31 33.2236 $w=3.3e-07 $l=1.9e-07 $layer=POLY_cond $X=0.94 $Y=1.69
+ $X2=0.75 $Y2=1.69
r98 11 34 58.5605 $w=2.9e-07 $l=3.06676e-07 $layer=POLY_cond $X=1.96 $Y=2.245
+ $X2=2.005 $Y2=1.96
r99 11 13 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=1.96 $Y=2.245
+ $X2=1.96 $Y2=2.64
r100 7 14 32.1775 $w=3.3e-07 $l=1.98997e-07 $layer=POLY_cond $X=1.015 $Y=1.525
+ $X2=0.94 $Y2=1.69
r101 7 9 484.564 $w=1.5e-07 $l=9.45e-07 $layer=POLY_cond $X=1.015 $Y=1.525
+ $X2=1.015 $Y2=0.58
r102 2 19 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=0.22
+ $Y=2.32 $X2=0.365 $Y2=2.465
r103 1 24 182 $w=1.7e-07 $l=2.57488e-07 $layer=licon1_NDIFF $count=1 $X=0.155
+ $Y=0.37 $X2=0.3 $Y2=0.565
.ends

.subckt PM_SKY130_FD_SC_HS__SDFXBP_1%SCE 2 3 4 7 9 11 12 14 16 17 19 20 26 29 33
+ 35 38
r80 32 35 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=1.885 $Y=1.065
+ $X2=2.095 $Y2=1.065
r81 32 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.885
+ $Y=1.065 $X2=1.885 $Y2=1.065
r82 26 33 5.16202 $w=4.73e-07 $l=2.05e-07 $layer=LI1_cond $X=1.68 $Y=1.047
+ $X2=1.885 $Y2=1.047
r83 26 38 4.02225 $w=4.73e-07 $l=1.15e-07 $layer=LI1_cond $X=1.68 $Y=1.047
+ $X2=1.565 $Y2=1.047
r84 24 29 9.23372 $w=2.61e-07 $l=5e-08 $layer=POLY_cond $X=0.565 $Y=1.12
+ $X2=0.515 $Y2=1.12
r85 23 38 34.9225 $w=3.28e-07 $l=1e-06 $layer=LI1_cond $X=0.565 $Y=1.12
+ $X2=1.565 $Y2=1.12
r86 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.565
+ $Y=1.12 $X2=0.565 $Y2=1.12
r87 17 35 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.095 $Y=0.9
+ $X2=2.095 $Y2=1.065
r88 17 19 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.095 $Y=0.9
+ $X2=2.095 $Y2=0.58
r89 14 16 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=1.09 $Y=2.245
+ $X2=1.09 $Y2=2.64
r90 13 20 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.665 $Y=2.17
+ $X2=0.59 $Y2=2.17
r91 12 14 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.015 $Y=2.17
+ $X2=1.09 $Y2=2.245
r92 12 13 179.468 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=1.015 $Y=2.17
+ $X2=0.665 $Y2=2.17
r93 9 20 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.59 $Y=2.245
+ $X2=0.59 $Y2=2.17
r94 9 11 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=0.59 $Y=2.245
+ $X2=0.59 $Y2=2.64
r95 5 29 15.717 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.515 $Y=0.955
+ $X2=0.515 $Y2=1.12
r96 5 7 192.287 $w=1.5e-07 $l=3.75e-07 $layer=POLY_cond $X=0.515 $Y=0.955
+ $X2=0.515 $Y2=0.58
r97 3 20 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.515 $Y=2.17
+ $X2=0.59 $Y2=2.17
r98 3 4 87.1702 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=0.515 $Y=2.17
+ $X2=0.345 $Y2=2.17
r99 2 4 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.27 $Y=2.095
+ $X2=0.345 $Y2=2.17
r100 1 29 45.2452 $w=2.61e-07 $l=3.16938e-07 $layer=POLY_cond $X=0.27 $Y=1.285
+ $X2=0.515 $Y2=1.12
r101 1 2 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=0.27 $Y=1.285 $X2=0.27
+ $Y2=2.095
.ends

.subckt PM_SKY130_FD_SC_HS__SDFXBP_1%D 3 6 7 9 10 13 14
c37 13 0 1.68868e-19 $X=1.465 $Y=1.62
r38 13 16 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.465 $Y=1.62
+ $X2=1.465 $Y2=1.785
r39 13 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.465 $Y=1.62
+ $X2=1.465 $Y2=1.455
r40 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.465
+ $Y=1.62 $X2=1.465 $Y2=1.62
r41 10 14 9.25447 $w=3.28e-07 $l=2.65e-07 $layer=LI1_cond $X=1.2 $Y=1.62
+ $X2=1.465 $Y2=1.62
r42 7 9 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=1.51 $Y=2.245
+ $X2=1.51 $Y2=2.64
r43 6 7 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=1.51 $Y=2.155 $X2=1.51
+ $Y2=2.245
r44 6 16 143.823 $w=1.8e-07 $l=3.7e-07 $layer=POLY_cond $X=1.51 $Y=2.155
+ $X2=1.51 $Y2=1.785
r45 3 15 448.67 $w=1.5e-07 $l=8.75e-07 $layer=POLY_cond $X=1.405 $Y=0.58
+ $X2=1.405 $Y2=1.455
.ends

.subckt PM_SKY130_FD_SC_HS__SDFXBP_1%SCD 3 6 7 9 10 11 15
c44 15 0 6.03804e-20 $X=2.545 $Y=1.775
c45 3 0 8.79478e-20 $X=2.485 $Y=0.58
r46 15 18 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.545 $Y=1.775
+ $X2=2.545 $Y2=1.94
r47 15 17 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.545 $Y=1.775
+ $X2=2.545 $Y2=1.61
r48 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.545
+ $Y=1.775 $X2=2.545 $Y2=1.775
r49 11 16 8.68508 $w=3.43e-07 $l=2.6e-07 $layer=LI1_cond $X=2.552 $Y=2.035
+ $X2=2.552 $Y2=1.775
r50 10 16 3.67446 $w=3.43e-07 $l=1.1e-07 $layer=LI1_cond $X=2.552 $Y=1.665
+ $X2=2.552 $Y2=1.775
r51 7 9 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=2.5 $Y=2.245 $X2=2.5
+ $Y2=2.64
r52 6 7 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=2.5 $Y=2.155 $X2=2.5
+ $Y2=2.245
r53 6 18 83.5726 $w=1.8e-07 $l=2.15e-07 $layer=POLY_cond $X=2.5 $Y=2.155 $X2=2.5
+ $Y2=1.94
r54 3 17 528.149 $w=1.5e-07 $l=1.03e-06 $layer=POLY_cond $X=2.485 $Y=0.58
+ $X2=2.485 $Y2=1.61
.ends

.subckt PM_SKY130_FD_SC_HS__SDFXBP_1%CLK 1 3 4 6 7 10
c43 7 0 8.79478e-20 $X=3.6 $Y=1.295
c44 4 0 6.57996e-20 $X=3.21 $Y=1.765
r45 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.4
+ $Y=1.385 $X2=3.4 $Y2=1.385
r46 10 12 27.6677 $w=3.31e-07 $l=1.9e-07 $layer=POLY_cond $X=3.21 $Y=1.492
+ $X2=3.4 $Y2=1.492
r47 7 13 6.22942 $w=3.68e-07 $l=2e-07 $layer=LI1_cond $X=3.6 $Y=1.365 $X2=3.4
+ $Y2=1.365
r48 4 10 21.295 $w=1.5e-07 $l=2.73e-07 $layer=POLY_cond $X=3.21 $Y=1.765
+ $X2=3.21 $Y2=1.492
r49 4 6 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.21 $Y=1.765
+ $X2=3.21 $Y2=2.4
r50 1 10 32.7644 $w=3.31e-07 $l=3.67674e-07 $layer=POLY_cond $X=2.985 $Y=1.22
+ $X2=3.21 $Y2=1.492
r51 1 3 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=2.985 $Y=1.22 $X2=2.985
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HS__SDFXBP_1%A_828_74# 1 2 7 9 10 12 15 18 19 21 24 25
+ 28 30 31 33 34 37 40 41 43 46 47 48 55 56 61 62 64 65 67 68 69 72 73
c205 68 0 1.71252e-20 $X=7.615 $Y=1.255
c206 62 0 2.55557e-20 $X=5.075 $Y=2.155
c207 56 0 1.07508e-19 $X=8.515 $Y=1.52
c208 55 0 8.08518e-20 $X=8.515 $Y=1.52
c209 37 0 1.67448e-19 $X=5.892 $Y=0.69
c210 25 0 1.8865e-19 $X=8.395 $Y=2.17
c211 24 0 1.40714e-19 $X=8.395 $Y=2.02
r212 72 73 8.96645 $w=2.53e-07 $l=1.7e-07 $layer=LI1_cond $X=8.05 $Y=1.43
+ $X2=8.22 $Y2=1.43
r213 68 81 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=7.615 $Y=1.255
+ $X2=7.615 $Y2=1.09
r214 67 70 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=7.695 $Y=1.255
+ $X2=7.695 $Y2=1.335
r215 67 69 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=7.695 $Y=1.255
+ $X2=7.695 $Y2=1.09
r216 67 68 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.615
+ $Y=1.255 $X2=7.615 $Y2=1.255
r217 62 75 50.9155 $w=2.84e-07 $l=3e-07 $layer=POLY_cond $X=5.075 $Y=2.197
+ $X2=5.375 $Y2=2.197
r218 61 63 2.28037 $w=4.28e-07 $l=8e-08 $layer=LI1_cond $X=5.075 $Y=2.05
+ $X2=5.155 $Y2=2.05
r219 61 62 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.075
+ $Y=2.155 $X2=5.075 $Y2=2.155
r220 59 61 12.9696 $w=4.28e-07 $l=4.55e-07 $layer=LI1_cond $X=4.62 $Y=2.05
+ $X2=5.075 $Y2=2.05
r221 56 85 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=8.515 $Y=1.52
+ $X2=8.515 $Y2=1.685
r222 55 73 13.3322 $w=2.53e-07 $l=2.95e-07 $layer=LI1_cond $X=8.515 $Y=1.482
+ $X2=8.22 $Y2=1.482
r223 55 56 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.515
+ $Y=1.52 $X2=8.515 $Y2=1.52
r224 52 70 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.86 $Y=1.335
+ $X2=7.695 $Y2=1.335
r225 52 72 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=7.86 $Y=1.335
+ $X2=8.05 $Y2=1.335
r226 49 69 43.385 $w=1.68e-07 $l=6.65e-07 $layer=LI1_cond $X=7.775 $Y=0.425
+ $X2=7.775 $Y2=1.09
r227 47 49 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.69 $Y=0.34
+ $X2=7.775 $Y2=0.425
r228 47 48 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=7.69 $Y=0.34
+ $X2=7.02 $Y2=0.34
r229 45 48 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.935 $Y=0.425
+ $X2=7.02 $Y2=0.34
r230 45 46 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=6.935 $Y=0.425
+ $X2=6.935 $Y2=0.69
r231 44 65 3.25423 $w=1.7e-07 $l=1.43e-07 $layer=LI1_cond $X=6.035 $Y=0.775
+ $X2=5.892 $Y2=0.775
r232 43 46 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.85 $Y=0.775
+ $X2=6.935 $Y2=0.69
r233 43 44 53.1711 $w=1.68e-07 $l=8.15e-07 $layer=LI1_cond $X=6.85 $Y=0.775
+ $X2=6.035 $Y2=0.775
r234 41 76 27.9778 $w=3.3e-07 $l=1.6e-07 $layer=POLY_cond $X=5.87 $Y=1.195
+ $X2=5.71 $Y2=1.195
r235 40 41 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.87
+ $Y=1.195 $X2=5.87 $Y2=1.195
r236 38 65 3.29812 $w=2.85e-07 $l=8.5e-08 $layer=LI1_cond $X=5.892 $Y=0.86
+ $X2=5.892 $Y2=0.775
r237 38 40 13.5463 $w=2.83e-07 $l=3.35e-07 $layer=LI1_cond $X=5.892 $Y=0.86
+ $X2=5.892 $Y2=1.195
r238 37 65 3.29812 $w=2.85e-07 $l=8.5e-08 $layer=LI1_cond $X=5.892 $Y=0.69
+ $X2=5.892 $Y2=0.775
r239 36 37 10.7157 $w=2.83e-07 $l=2.65e-07 $layer=LI1_cond $X=5.892 $Y=0.425
+ $X2=5.892 $Y2=0.69
r240 35 64 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.24 $Y=0.34
+ $X2=5.155 $Y2=0.34
r241 34 36 7.39867 $w=1.7e-07 $l=1.79538e-07 $layer=LI1_cond $X=5.75 $Y=0.34
+ $X2=5.892 $Y2=0.425
r242 34 35 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=5.75 $Y=0.34
+ $X2=5.24 $Y2=0.34
r243 33 63 6.19161 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=5.155 $Y=1.82
+ $X2=5.155 $Y2=2.05
r244 32 64 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.155 $Y=0.425
+ $X2=5.155 $Y2=0.34
r245 32 33 91.0107 $w=1.68e-07 $l=1.395e-06 $layer=LI1_cond $X=5.155 $Y=0.425
+ $X2=5.155 $Y2=1.82
r246 30 64 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.07 $Y=0.34
+ $X2=5.155 $Y2=0.34
r247 30 31 40.7754 $w=1.68e-07 $l=6.25e-07 $layer=LI1_cond $X=5.07 $Y=0.34
+ $X2=4.445 $Y2=0.34
r248 26 31 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=4.32 $Y=0.425
+ $X2=4.445 $Y2=0.34
r249 26 28 4.14879 $w=2.48e-07 $l=9e-08 $layer=LI1_cond $X=4.32 $Y=0.425
+ $X2=4.32 $Y2=0.515
r250 24 25 60.4563 $w=1.8e-07 $l=1.5e-07 $layer=POLY_cond $X=8.395 $Y=2.02
+ $X2=8.395 $Y2=2.17
r251 24 85 171.777 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=8.425 $Y=2.02
+ $X2=8.425 $Y2=1.685
r252 19 21 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=8.38 $Y=2.465
+ $X2=8.38 $Y2=2.75
r253 18 19 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=8.38 $Y=2.375
+ $X2=8.38 $Y2=2.465
r254 18 25 79.6855 $w=1.8e-07 $l=2.05e-07 $layer=POLY_cond $X=8.38 $Y=2.375
+ $X2=8.38 $Y2=2.17
r255 15 81 228.181 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=7.57 $Y=0.645
+ $X2=7.57 $Y2=1.09
r256 10 76 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.71 $Y=1.03
+ $X2=5.71 $Y2=1.195
r257 10 12 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=5.71 $Y=1.03
+ $X2=5.71 $Y2=0.71
r258 7 75 17.6835 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=5.375 $Y=2.405
+ $X2=5.375 $Y2=2.197
r259 7 9 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=5.375 $Y=2.405
+ $X2=5.375 $Y2=2.69
r260 2 59 600 $w=1.7e-07 $l=2.43721e-07 $layer=licon1_PDIFF $count=1 $X=4.47
+ $Y=1.84 $X2=4.62 $Y2=2.02
r261 1 28 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=4.14
+ $Y=0.37 $X2=4.28 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__SDFXBP_1%A_612_74# 1 2 9 11 13 15 16 20 22 25 26 28
+ 29 31 33 36 38 39 42 46 48 49 50 55 56 58 59 60 62 63 72 75 85
c215 75 0 1.40714e-19 $X=7.72 $Y=1.795
c216 72 0 2.55557e-20 $X=6.02 $Y=2.035
c217 50 0 6.57996e-20 $X=3.855 $Y=1.905
c218 42 0 5.43913e-20 $X=8.33 $Y=1.04
c219 20 0 1.67448e-19 $X=5.03 $Y=0.71
r220 76 85 20.5631 $w=2.93e-07 $l=1.25e-07 $layer=POLY_cond $X=7.72 $Y=1.837
+ $X2=7.845 $Y2=1.837
r221 75 78 8.46257 $w=3.13e-07 $l=1.65e-07 $layer=LI1_cond $X=7.722 $Y=1.795
+ $X2=7.722 $Y2=1.96
r222 75 76 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.72
+ $Y=1.795 $X2=7.72 $Y2=1.795
r223 69 72 6.28605 $w=3.28e-07 $l=1.8e-07 $layer=LI1_cond $X=5.84 $Y=2.035
+ $X2=6.02 $Y2=2.035
r224 69 70 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.84
+ $Y=2.035 $X2=5.84 $Y2=2.035
r225 63 66 4.01609 $w=3.28e-07 $l=1.15e-07 $layer=LI1_cond $X=3.435 $Y=1.905
+ $X2=3.435 $Y2=2.02
r226 62 78 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=7.65 $Y=2.52
+ $X2=7.65 $Y2=1.96
r227 59 62 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.565 $Y=2.605
+ $X2=7.65 $Y2=2.52
r228 59 60 95.2513 $w=1.68e-07 $l=1.46e-06 $layer=LI1_cond $X=7.565 $Y=2.605
+ $X2=6.105 $Y2=2.605
r229 58 60 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.02 $Y=2.52
+ $X2=6.105 $Y2=2.605
r230 57 72 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.02 $Y=2.2
+ $X2=6.02 $Y2=2.035
r231 57 58 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=6.02 $Y=2.2 $X2=6.02
+ $Y2=2.52
r232 56 81 25.295 $w=3.65e-07 $l=1.6e-07 $layer=POLY_cond $X=3.957 $Y=1.515
+ $X2=3.957 $Y2=1.675
r233 56 80 46.6671 $w=3.65e-07 $l=1.65e-07 $layer=POLY_cond $X=3.957 $Y=1.515
+ $X2=3.957 $Y2=1.35
r234 55 56 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.94
+ $Y=1.515 $X2=3.94 $Y2=1.515
r235 53 55 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=3.94 $Y=1.82
+ $X2=3.94 $Y2=1.515
r236 52 55 32.9465 $w=1.68e-07 $l=5.05e-07 $layer=LI1_cond $X=3.94 $Y=1.01
+ $X2=3.94 $Y2=1.515
r237 51 63 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.6 $Y=1.905
+ $X2=3.435 $Y2=1.905
r238 50 53 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.855 $Y=1.905
+ $X2=3.94 $Y2=1.82
r239 50 51 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=3.855 $Y=1.905
+ $X2=3.6 $Y2=1.905
r240 48 52 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.855 $Y=0.925
+ $X2=3.94 $Y2=1.01
r241 48 49 31.9679 $w=1.68e-07 $l=4.9e-07 $layer=LI1_cond $X=3.855 $Y=0.925
+ $X2=3.365 $Y2=0.925
r242 44 49 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.2 $Y=0.84
+ $X2=3.365 $Y2=0.925
r243 44 46 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=3.2 $Y=0.84
+ $X2=3.2 $Y2=0.515
r244 40 42 135.883 $w=1.5e-07 $l=2.65e-07 $layer=POLY_cond $X=8.065 $Y=1.04
+ $X2=8.33 $Y2=1.04
r245 34 42 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=8.33 $Y=0.965
+ $X2=8.33 $Y2=1.04
r246 34 36 197.415 $w=1.5e-07 $l=3.85e-07 $layer=POLY_cond $X=8.33 $Y=0.965
+ $X2=8.33 $Y2=0.58
r247 33 85 36.1911 $w=2.93e-07 $l=3.06496e-07 $layer=POLY_cond $X=8.065 $Y=1.63
+ $X2=7.845 $Y2=1.837
r248 32 40 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=8.065 $Y=1.115
+ $X2=8.065 $Y2=1.04
r249 32 33 264.074 $w=1.5e-07 $l=5.15e-07 $layer=POLY_cond $X=8.065 $Y=1.115
+ $X2=8.065 $Y2=1.63
r250 29 85 18.414 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=7.845 $Y=2.045
+ $X2=7.845 $Y2=1.837
r251 29 31 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=7.845 $Y=2.045
+ $X2=7.845 $Y2=2.54
r252 26 70 79.7845 $w=2.46e-07 $l=3.77425e-07 $layer=POLY_cond $X=5.825 $Y=2.405
+ $X2=5.84 $Y2=2.035
r253 26 28 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=5.825 $Y=2.405
+ $X2=5.825 $Y2=2.69
r254 25 70 3.22709 $w=3.3e-07 $l=8.75758e-08 $layer=POLY_cond $X=5.84 $Y=2.035
+ $X2=5.84 $Y2=2.035
r255 24 25 49.8355 $w=3.3e-07 $l=2.85e-07 $layer=POLY_cond $X=5.84 $Y=1.75
+ $X2=5.84 $Y2=2.035
r256 23 39 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.105 $Y=1.675
+ $X2=5.03 $Y2=1.675
r257 22 24 32.1775 $w=1.5e-07 $l=1.98997e-07 $layer=POLY_cond $X=5.675 $Y=1.675
+ $X2=5.84 $Y2=1.75
r258 22 23 292.277 $w=1.5e-07 $l=5.7e-07 $layer=POLY_cond $X=5.675 $Y=1.675
+ $X2=5.105 $Y2=1.675
r259 18 39 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.03 $Y=1.6
+ $X2=5.03 $Y2=1.675
r260 18 20 456.362 $w=1.5e-07 $l=8.9e-07 $layer=POLY_cond $X=5.03 $Y=1.6
+ $X2=5.03 $Y2=0.71
r261 17 38 20.4101 $w=1.5e-07 $l=9.34345e-08 $layer=POLY_cond $X=4.485 $Y=1.675
+ $X2=4.395 $Y2=1.682
r262 16 39 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.955 $Y=1.675
+ $X2=5.03 $Y2=1.675
r263 16 17 241 $w=1.5e-07 $l=4.7e-07 $layer=POLY_cond $X=4.955 $Y=1.675
+ $X2=4.485 $Y2=1.675
r264 13 38 5.30422 $w=1.5e-07 $l=8.3e-08 $layer=POLY_cond $X=4.395 $Y=1.765
+ $X2=4.395 $Y2=1.682
r265 13 15 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=4.395 $Y=1.765
+ $X2=4.395 $Y2=2.4
r266 12 81 23.6381 $w=1.5e-07 $l=1.83e-07 $layer=POLY_cond $X=4.14 $Y=1.675
+ $X2=3.957 $Y2=1.675
r267 11 38 20.4101 $w=1.5e-07 $l=9.34345e-08 $layer=POLY_cond $X=4.305 $Y=1.675
+ $X2=4.395 $Y2=1.682
r268 11 12 84.6064 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.305 $Y=1.675
+ $X2=4.14 $Y2=1.675
r269 9 80 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=4.065 $Y=0.74
+ $X2=4.065 $Y2=1.35
r270 2 66 600 $w=1.7e-07 $l=2.43721e-07 $layer=licon1_PDIFF $count=1 $X=3.285
+ $Y=1.84 $X2=3.435 $Y2=2.02
r271 1 46 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.06
+ $Y=0.37 $X2=3.2 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__SDFXBP_1%A_1243_398# 1 2 7 8 9 11 14 17 18 21 23 24
+ 28 34
c77 17 0 1.47351e-19 $X=6.305 $Y=1.99
r78 26 28 3.91831 $w=2.48e-07 $l=8.5e-08 $layer=LI1_cond $X=7.19 $Y=2.225
+ $X2=7.275 $Y2=2.225
r79 24 28 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.275 $Y=2.1
+ $X2=7.275 $Y2=2.225
r80 23 24 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=7.275 $Y=1.36
+ $X2=7.275 $Y2=2.1
r81 21 35 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.41 $Y=1.195
+ $X2=6.41 $Y2=1.36
r82 21 34 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.41 $Y=1.195
+ $X2=6.41 $Y2=1.03
r83 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.41
+ $Y=1.195 $X2=6.41 $Y2=1.195
r84 18 23 9.48765 $w=2.37e-07 $l=2.0106e-07 $layer=LI1_cond $X=7.355 $Y=1.195
+ $X2=7.275 $Y2=1.36
r85 18 31 24.7089 $w=2.37e-07 $l=4.8e-07 $layer=LI1_cond $X=7.355 $Y=1.195
+ $X2=7.355 $Y2=0.715
r86 18 20 27.2396 $w=3.28e-07 $l=7.8e-07 $layer=LI1_cond $X=7.19 $Y=1.195
+ $X2=6.41 $Y2=1.195
r87 17 35 323.043 $w=1.5e-07 $l=6.3e-07 $layer=POLY_cond $X=6.32 $Y=1.99
+ $X2=6.32 $Y2=1.36
r88 14 34 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=6.32 $Y=0.71
+ $X2=6.32 $Y2=1.03
r89 9 11 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=6.305 $Y=2.405
+ $X2=6.305 $Y2=2.69
r90 8 9 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=6.305 $Y=2.315 $X2=6.305
+ $Y2=2.405
r91 7 17 37.1337 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=6.305 $Y=2.08 $X2=6.305
+ $Y2=1.99
r92 7 8 91.3468 $w=1.8e-07 $l=2.35e-07 $layer=POLY_cond $X=6.305 $Y=2.08
+ $X2=6.305 $Y2=2.315
r93 2 26 600 $w=1.7e-07 $l=2.5229e-07 $layer=licon1_PDIFF $count=1 $X=7 $Y=2.12
+ $X2=7.19 $Y2=2.265
r94 1 31 182 $w=1.7e-07 $l=4.11157e-07 $layer=licon1_NDIFF $count=1 $X=7.21
+ $Y=0.37 $X2=7.355 $Y2=0.715
.ends

.subckt PM_SKY130_FD_SC_HS__SDFXBP_1%A_1021_100# 1 2 7 9 12 16 20 22 24 25 27
c80 25 0 1.47351e-19 $X=5.587 $Y=2.46
r81 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.855
+ $Y=1.765 $X2=6.855 $Y2=1.765
r82 27 30 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=6.855 $Y=1.615
+ $X2=6.855 $Y2=1.765
r83 24 25 10.6092 $w=3.53e-07 $l=2.3e-07 $layer=LI1_cond $X=5.587 $Y=2.69
+ $X2=5.587 $Y2=2.46
r84 21 22 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.58 $Y=1.615
+ $X2=5.495 $Y2=1.615
r85 20 27 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.69 $Y=1.615
+ $X2=6.855 $Y2=1.615
r86 20 21 72.4171 $w=1.68e-07 $l=1.11e-06 $layer=LI1_cond $X=6.69 $Y=1.615
+ $X2=5.58 $Y2=1.615
r87 18 22 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.495 $Y=1.7
+ $X2=5.495 $Y2=1.615
r88 18 25 49.5829 $w=1.68e-07 $l=7.6e-07 $layer=LI1_cond $X=5.495 $Y=1.7
+ $X2=5.495 $Y2=2.46
r89 14 22 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.495 $Y=1.53
+ $X2=5.495 $Y2=1.615
r90 14 16 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=5.495 $Y=1.53
+ $X2=5.495 $Y2=0.765
r91 10 31 40.2632 $w=4.32e-07 $l=2.5446e-07 $layer=POLY_cond $X=7.135 $Y=1.6
+ $X2=6.95 $Y2=1.765
r92 10 12 489.691 $w=1.5e-07 $l=9.55e-07 $layer=POLY_cond $X=7.135 $Y=1.6
+ $X2=7.135 $Y2=0.645
r93 7 31 53.0942 $w=4.32e-07 $l=2.92233e-07 $layer=POLY_cond $X=6.925 $Y=2.045
+ $X2=6.95 $Y2=1.765
r94 7 9 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=6.925 $Y=2.045
+ $X2=6.925 $Y2=2.54
r95 2 24 600 $w=1.7e-07 $l=2.74955e-07 $layer=licon1_PDIFF $count=1 $X=5.45
+ $Y=2.48 $X2=5.6 $Y2=2.69
r96 1 16 182 $w=1.7e-07 $l=5.05421e-07 $layer=licon1_NDIFF $count=1 $X=5.105
+ $Y=0.5 $X2=5.495 $Y2=0.765
.ends

.subckt PM_SKY130_FD_SC_HS__SDFXBP_1%A_1723_48# 1 2 9 11 13 15 16 20 22 24 25 29
+ 35 38 40 41 42 43 48 53 56 61 64 66 67 69
c140 67 0 1.65961e-19 $X=9.775 $Y=1.94
c141 43 0 1.8865e-19 $X=9.6 $Y=2.235
c142 38 0 8.08518e-20 $X=8.965 $Y=1.07
c143 9 0 3.89393e-20 $X=8.69 $Y=0.58
r144 66 68 4.2805 $w=3.48e-07 $l=1.3e-07 $layer=LI1_cond $X=9.775 $Y=2.105
+ $X2=9.775 $Y2=2.235
r145 66 67 8.48848 $w=3.48e-07 $l=1.65e-07 $layer=LI1_cond $X=9.775 $Y=2.105
+ $X2=9.775 $Y2=1.94
r146 59 69 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.95 $Y=1.485
+ $X2=9.865 $Y2=1.485
r147 59 61 16.0644 $w=3.28e-07 $l=4.6e-07 $layer=LI1_cond $X=9.95 $Y=1.485
+ $X2=10.41 $Y2=1.485
r148 57 69 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.865 $Y=1.65
+ $X2=9.865 $Y2=1.485
r149 57 67 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=9.865 $Y=1.65
+ $X2=9.865 $Y2=1.94
r150 56 69 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.865 $Y=1.32
+ $X2=9.865 $Y2=1.485
r151 56 64 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=9.865 $Y=1.32
+ $X2=9.865 $Y2=0.93
r152 51 68 3.7866 $w=3.48e-07 $l=1.15e-07 $layer=LI1_cond $X=9.775 $Y=2.35
+ $X2=9.775 $Y2=2.235
r153 51 53 15.311 $w=3.48e-07 $l=4.65e-07 $layer=LI1_cond $X=9.775 $Y=2.35
+ $X2=9.775 $Y2=2.815
r154 48 64 8.99121 $w=3.58e-07 $l=1.8e-07 $layer=LI1_cond $X=9.77 $Y=0.75
+ $X2=9.77 $Y2=0.93
r155 48 50 3.72778 $w=3.6e-07 $l=1.1e-07 $layer=LI1_cond $X=9.77 $Y=0.75
+ $X2=9.77 $Y2=0.64
r156 45 46 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.875
+ $Y=2.215 $X2=8.875 $Y2=2.215
r157 43 68 3.19443 $w=2.3e-07 $l=1.75e-07 $layer=LI1_cond $X=9.6 $Y=2.235
+ $X2=9.775 $Y2=2.235
r158 43 45 36.327 $w=2.28e-07 $l=7.25e-07 $layer=LI1_cond $X=9.6 $Y=2.235
+ $X2=8.875 $Y2=2.235
r159 41 42 48.5235 $w=2.05e-07 $l=1.5e-07 $layer=POLY_cond $X=11.467 $Y=1.79
+ $X2=11.467 $Y2=1.94
r160 36 38 141.011 $w=1.5e-07 $l=2.75e-07 $layer=POLY_cond $X=8.69 $Y=1.07
+ $X2=8.965 $Y2=1.07
r161 35 42 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=11.48 $Y=2.435
+ $X2=11.48 $Y2=1.94
r162 31 40 32.2453 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=11.44 $Y=1.59
+ $X2=11.44 $Y2=1.455
r163 31 41 102.553 $w=1.5e-07 $l=2e-07 $layer=POLY_cond $X=11.44 $Y=1.59
+ $X2=11.44 $Y2=1.79
r164 27 40 32.2453 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=11.44 $Y=1.32
+ $X2=11.44 $Y2=1.455
r165 27 29 271.766 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=11.44 $Y=1.32
+ $X2=11.44 $Y2=0.79
r166 25 40 2.60871 $w=2.7e-07 $l=7.5e-08 $layer=POLY_cond $X=11.365 $Y=1.455
+ $X2=11.44 $Y2=1.455
r167 25 26 169.963 $w=2.7e-07 $l=7.65e-07 $layer=POLY_cond $X=11.365 $Y=1.455
+ $X2=10.6 $Y2=1.455
r168 22 24 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=10.51 $Y=1.765
+ $X2=10.51 $Y2=2.4
r169 18 26 34.8256 $w=2.13e-07 $l=1.52381e-07 $layer=POLY_cond $X=10.45 $Y=1.32
+ $X2=10.487 $Y2=1.455
r170 18 20 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=10.45 $Y=1.32
+ $X2=10.45 $Y2=0.74
r171 16 22 67.6378 $w=2.13e-07 $l=2.91273e-07 $layer=POLY_cond $X=10.487
+ $Y=1.485 $X2=10.51 $Y2=1.765
r172 16 26 6.78873 $w=2.13e-07 $l=3e-08 $layer=POLY_cond $X=10.487 $Y=1.485
+ $X2=10.487 $Y2=1.455
r173 16 61 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=10.41
+ $Y=1.485 $X2=10.41 $Y2=1.485
r174 15 46 38.5562 $w=2.99e-07 $l=2.05122e-07 $layer=POLY_cond $X=8.965 $Y=2.05
+ $X2=8.875 $Y2=2.215
r175 14 38 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=8.965 $Y=1.145
+ $X2=8.965 $Y2=1.07
r176 14 15 464.053 $w=1.5e-07 $l=9.05e-07 $layer=POLY_cond $X=8.965 $Y=1.145
+ $X2=8.965 $Y2=2.05
r177 11 46 52.2586 $w=2.99e-07 $l=2.85044e-07 $layer=POLY_cond $X=8.8 $Y=2.465
+ $X2=8.875 $Y2=2.215
r178 11 13 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=8.8 $Y=2.465 $X2=8.8
+ $Y2=2.75
r179 7 36 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=8.69 $Y=0.995
+ $X2=8.69 $Y2=1.07
r180 7 9 212.798 $w=1.5e-07 $l=4.15e-07 $layer=POLY_cond $X=8.69 $Y=0.995
+ $X2=8.69 $Y2=0.58
r181 2 66 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=9.615
+ $Y=1.96 $X2=9.765 $Y2=2.105
r182 2 53 400 $w=1.7e-07 $l=9.26971e-07 $layer=licon1_PDIFF $count=1 $X=9.615
+ $Y=1.96 $X2=9.765 $Y2=2.815
r183 1 50 182 $w=1.7e-07 $l=3.32716e-07 $layer=licon1_NDIFF $count=1 $X=9.535
+ $Y=0.37 $X2=9.675 $Y2=0.64
.ends

.subckt PM_SKY130_FD_SC_HS__SDFXBP_1%A_1529_74# 1 2 8 11 13 15 18 20 24 25 27 28
+ 29 31 32 36 40 42 46 47
c123 42 0 9.33306e-20 $X=8.935 $Y=1.065
c124 40 0 1.07508e-19 $X=8.475 $Y=0.58
c125 29 0 1.71252e-20 $X=8.56 $Y=1.065
r126 47 49 46.4315 $w=3.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.455 $Y=1.265
+ $X2=9.455 $Y2=1.1
r127 46 47 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=9.445
+ $Y=1.265 $X2=9.445 $Y2=1.265
r128 42 44 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=8.935 $Y=1.065
+ $X2=8.935 $Y2=1.185
r129 38 40 9.36061 $w=4.58e-07 $l=3.6e-07 $layer=LI1_cond $X=8.115 $Y=0.58
+ $X2=8.475 $Y2=0.58
r130 33 44 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.02 $Y=1.185
+ $X2=8.935 $Y2=1.185
r131 32 46 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.28 $Y=1.185
+ $X2=9.445 $Y2=1.185
r132 32 33 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=9.28 $Y=1.185
+ $X2=9.02 $Y2=1.185
r133 30 44 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=8.935 $Y=1.27
+ $X2=8.935 $Y2=1.185
r134 30 31 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=8.935 $Y=1.27
+ $X2=8.935 $Y2=1.78
r135 28 42 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.85 $Y=1.065
+ $X2=8.935 $Y2=1.065
r136 28 29 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=8.85 $Y=1.065
+ $X2=8.56 $Y2=1.065
r137 27 29 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.475 $Y=0.98
+ $X2=8.56 $Y2=1.065
r138 26 40 6.6364 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=8.475 $Y=0.81
+ $X2=8.475 $Y2=0.58
r139 26 27 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=8.475 $Y=0.81
+ $X2=8.475 $Y2=0.98
r140 24 31 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.85 $Y=1.865
+ $X2=8.935 $Y2=1.78
r141 24 25 40.123 $w=1.68e-07 $l=6.15e-07 $layer=LI1_cond $X=8.85 $Y=1.865
+ $X2=8.235 $Y2=1.865
r142 22 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.15 $Y=1.95
+ $X2=8.235 $Y2=1.865
r143 22 36 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=8.15 $Y=1.95
+ $X2=8.15 $Y2=2.13
r144 18 36 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=8.07 $Y=2.295
+ $X2=8.07 $Y2=2.13
r145 18 20 18.1597 $w=3.28e-07 $l=5.2e-07 $layer=LI1_cond $X=8.07 $Y=2.295
+ $X2=8.07 $Y2=2.815
r146 13 15 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=9.54 $Y=1.885
+ $X2=9.54 $Y2=2.46
r147 11 49 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=9.46 $Y=0.645
+ $X2=9.46 $Y2=1.1
r148 8 13 49.5674 $w=2.82e-07 $l=3.29773e-07 $layer=POLY_cond $X=9.455 $Y=1.595
+ $X2=9.54 $Y2=1.885
r149 7 47 1.64869 $w=3.5e-07 $l=1e-08 $layer=POLY_cond $X=9.455 $Y=1.275
+ $X2=9.455 $Y2=1.265
r150 7 8 52.7581 $w=3.5e-07 $l=3.2e-07 $layer=POLY_cond $X=9.455 $Y=1.275
+ $X2=9.455 $Y2=1.595
r151 2 20 600 $w=1.7e-07 $l=7.66339e-07 $layer=licon1_PDIFF $count=1 $X=7.92
+ $Y=2.12 $X2=8.07 $Y2=2.815
r152 2 18 600 $w=1.7e-07 $l=2.38485e-07 $layer=licon1_PDIFF $count=1 $X=7.92
+ $Y=2.12 $X2=8.07 $Y2=2.295
r153 1 38 182 $w=1.7e-07 $l=5.65332e-07 $layer=licon1_NDIFF $count=1 $X=7.645
+ $Y=0.37 $X2=8.115 $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_HS__SDFXBP_1%A_2216_94# 1 2 7 9 10 12 15 19 23 26
r46 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=11.89
+ $Y=1.385 $X2=11.89 $Y2=1.385
r47 21 26 0.153733 $w=3.3e-07 $l=1.25e-07 $layer=LI1_cond $X=11.34 $Y=1.385
+ $X2=11.215 $Y2=1.385
r48 21 23 19.2074 $w=3.28e-07 $l=5.5e-07 $layer=LI1_cond $X=11.34 $Y=1.385
+ $X2=11.89 $Y2=1.385
r49 17 26 6.7841 $w=2.35e-07 $l=1.65e-07 $layer=LI1_cond $X=11.215 $Y=1.55
+ $X2=11.215 $Y2=1.385
r50 17 19 28.1196 $w=2.48e-07 $l=6.1e-07 $layer=LI1_cond $X=11.215 $Y=1.55
+ $X2=11.215 $Y2=2.16
r51 13 26 6.7841 $w=2.35e-07 $l=1.72337e-07 $layer=LI1_cond $X=11.2 $Y=1.22
+ $X2=11.215 $Y2=1.385
r52 13 15 20.1678 $w=2.18e-07 $l=3.85e-07 $layer=LI1_cond $X=11.2 $Y=1.22
+ $X2=11.2 $Y2=0.835
r53 10 24 76.8038 $w=2.73e-07 $l=4.20357e-07 $layer=POLY_cond $X=11.985 $Y=1.765
+ $X2=11.9 $Y2=1.385
r54 10 12 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=11.985 $Y=1.765
+ $X2=11.985 $Y2=2.4
r55 7 24 38.8441 $w=2.73e-07 $l=2.03101e-07 $layer=POLY_cond $X=11.985 $Y=1.22
+ $X2=11.9 $Y2=1.385
r56 7 9 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=11.985 $Y=1.22
+ $X2=11.985 $Y2=0.74
r57 2 19 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=11.13
+ $Y=2.015 $X2=11.255 $Y2=2.16
r58 1 15 182 $w=1.7e-07 $l=4.31451e-07 $layer=licon1_NDIFF $count=1 $X=11.08
+ $Y=0.47 $X2=11.225 $Y2=0.835
.ends

.subckt PM_SKY130_FD_SC_HS__SDFXBP_1%VPWR 1 2 3 4 5 6 7 26 30 34 38 42 48 50 52
+ 57 62 67 72 77 84 85 88 91 98 101 104 107 110
r140 110 111 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.76 $Y=3.33
+ $X2=11.76 $Y2=3.33
r141 107 108 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.32 $Y=3.33
+ $X2=10.32 $Y2=3.33
r142 104 105 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r143 101 102 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r144 98 99 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r145 94 95 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r146 91 94 10.4403 $w=5.88e-07 $l=5.15e-07 $layer=LI1_cond $X=2.855 $Y=2.815
+ $X2=2.855 $Y2=3.33
r147 88 89 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r148 85 111 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.24 $Y=3.33
+ $X2=11.76 $Y2=3.33
r149 84 85 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.24 $Y=3.33
+ $X2=12.24 $Y2=3.33
r150 82 110 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.87 $Y=3.33
+ $X2=11.705 $Y2=3.33
r151 82 84 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=11.87 $Y=3.33
+ $X2=12.24 $Y2=3.33
r152 81 111 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.28 $Y=3.33
+ $X2=11.76 $Y2=3.33
r153 81 108 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=11.28 $Y=3.33
+ $X2=10.32 $Y2=3.33
r154 80 81 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=11.28 $Y=3.33
+ $X2=11.28 $Y2=3.33
r155 78 107 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.45 $Y=3.33
+ $X2=10.285 $Y2=3.33
r156 78 80 54.1497 $w=1.68e-07 $l=8.3e-07 $layer=LI1_cond $X=10.45 $Y=3.33
+ $X2=11.28 $Y2=3.33
r157 77 110 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.54 $Y=3.33
+ $X2=11.705 $Y2=3.33
r158 77 80 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=11.54 $Y=3.33
+ $X2=11.28 $Y2=3.33
r159 76 108 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.84 $Y=3.33
+ $X2=10.32 $Y2=3.33
r160 76 105 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=9.84 $Y=3.33
+ $X2=8.88 $Y2=3.33
r161 75 76 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.84 $Y=3.33
+ $X2=9.84 $Y2=3.33
r162 73 104 12.1981 $w=1.7e-07 $l=2.85e-07 $layer=LI1_cond $X=9.43 $Y=3.33
+ $X2=9.145 $Y2=3.33
r163 73 75 26.7487 $w=1.68e-07 $l=4.1e-07 $layer=LI1_cond $X=9.43 $Y=3.33
+ $X2=9.84 $Y2=3.33
r164 72 107 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.12 $Y=3.33
+ $X2=10.285 $Y2=3.33
r165 72 75 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=10.12 $Y=3.33
+ $X2=9.84 $Y2=3.33
r166 71 105 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=8.88 $Y2=3.33
r167 71 102 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=6.48 $Y2=3.33
r168 70 71 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r169 68 101 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.78 $Y=3.33
+ $X2=6.615 $Y2=3.33
r170 68 70 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=6.78 $Y=3.33
+ $X2=6.96 $Y2=3.33
r171 67 104 12.1981 $w=1.7e-07 $l=2.85e-07 $layer=LI1_cond $X=8.86 $Y=3.33
+ $X2=9.145 $Y2=3.33
r172 67 70 123.957 $w=1.68e-07 $l=1.9e-06 $layer=LI1_cond $X=8.86 $Y=3.33
+ $X2=6.96 $Y2=3.33
r173 66 99 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=4.08 $Y2=3.33
r174 65 66 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r175 63 98 11.3601 $w=1.7e-07 $l=2.53e-07 $layer=LI1_cond $X=4.335 $Y=3.33
+ $X2=4.082 $Y2=3.33
r176 63 65 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=4.335 $Y=3.33
+ $X2=4.56 $Y2=3.33
r177 62 101 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.45 $Y=3.33
+ $X2=6.615 $Y2=3.33
r178 62 65 123.305 $w=1.68e-07 $l=1.89e-06 $layer=LI1_cond $X=6.45 $Y=3.33
+ $X2=4.56 $Y2=3.33
r179 61 99 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.08 $Y2=3.33
r180 61 95 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=2.64 $Y2=3.33
r181 60 61 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r182 58 94 8.20854 $w=1.7e-07 $l=2.95e-07 $layer=LI1_cond $X=3.15 $Y=3.33
+ $X2=2.855 $Y2=3.33
r183 58 60 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=3.15 $Y=3.33
+ $X2=3.6 $Y2=3.33
r184 57 98 11.3601 $w=1.7e-07 $l=2.52e-07 $layer=LI1_cond $X=3.83 $Y=3.33
+ $X2=4.082 $Y2=3.33
r185 57 60 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=3.83 $Y=3.33
+ $X2=3.6 $Y2=3.33
r186 56 95 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.64 $Y2=3.33
r187 56 89 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r188 55 56 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r189 53 88 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.03 $Y=3.33
+ $X2=0.865 $Y2=3.33
r190 53 55 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=1.03 $Y=3.33
+ $X2=1.2 $Y2=3.33
r191 52 94 8.20854 $w=1.7e-07 $l=2.95e-07 $layer=LI1_cond $X=2.56 $Y=3.33
+ $X2=2.855 $Y2=3.33
r192 52 55 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=2.56 $Y=3.33
+ $X2=1.2 $Y2=3.33
r193 50 102 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=6.24 $Y=3.33
+ $X2=6.48 $Y2=3.33
r194 50 66 0.468274 $w=4.9e-07 $l=1.68e-06 $layer=MET1_cond $X=6.24 $Y=3.33
+ $X2=4.56 $Y2=3.33
r195 46 110 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=11.705 $Y=3.245
+ $X2=11.705 $Y2=3.33
r196 46 48 37.8909 $w=3.28e-07 $l=1.085e-06 $layer=LI1_cond $X=11.705 $Y=3.245
+ $X2=11.705 $Y2=2.16
r197 42 45 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=10.285 $Y=1.985
+ $X2=10.285 $Y2=2.815
r198 40 107 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=10.285 $Y=3.245
+ $X2=10.285 $Y2=3.33
r199 40 45 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=10.285 $Y=3.245
+ $X2=10.285 $Y2=2.815
r200 36 104 2.39972 $w=5.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.145 $Y=3.245
+ $X2=9.145 $Y2=3.33
r201 36 38 9.02305 $w=5.68e-07 $l=4.3e-07 $layer=LI1_cond $X=9.145 $Y=3.245
+ $X2=9.145 $Y2=2.815
r202 32 101 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.615 $Y=3.245
+ $X2=6.615 $Y2=3.33
r203 32 34 7.68295 $w=3.28e-07 $l=2.2e-07 $layer=LI1_cond $X=6.615 $Y=3.245
+ $X2=6.615 $Y2=3.025
r204 28 98 2.09999 $w=5.05e-07 $l=8.5e-08 $layer=LI1_cond $X=4.082 $Y=3.245
+ $X2=4.082 $Y2=3.33
r205 28 30 10.1844 $w=5.03e-07 $l=4.3e-07 $layer=LI1_cond $X=4.082 $Y=3.245
+ $X2=4.082 $Y2=2.815
r206 24 88 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.865 $Y=3.245
+ $X2=0.865 $Y2=3.33
r207 24 26 27.2396 $w=3.28e-07 $l=7.8e-07 $layer=LI1_cond $X=0.865 $Y=3.245
+ $X2=0.865 $Y2=2.465
r208 7 48 300 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=2 $X=11.555
+ $Y=2.015 $X2=11.705 $Y2=2.16
r209 6 45 400 $w=1.7e-07 $l=1.03562e-06 $layer=licon1_PDIFF $count=1 $X=10.16
+ $Y=1.84 $X2=10.285 $Y2=2.815
r210 6 42 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=10.16
+ $Y=1.84 $X2=10.285 $Y2=1.985
r211 5 38 600 $w=1.7e-07 $l=3.995e-07 $layer=licon1_PDIFF $count=1 $X=8.875
+ $Y=2.54 $X2=9.16 $Y2=2.815
r212 4 34 600 $w=1.7e-07 $l=6.51997e-07 $layer=licon1_PDIFF $count=1 $X=6.38
+ $Y=2.48 $X2=6.615 $Y2=3.025
r213 3 30 600 $w=1.7e-07 $l=1.08392e-06 $layer=licon1_PDIFF $count=1 $X=3.85
+ $Y=1.84 $X2=4.08 $Y2=2.815
r214 2 91 600 $w=1.7e-07 $l=6.19375e-07 $layer=licon1_PDIFF $count=1 $X=2.575
+ $Y=2.32 $X2=2.855 $Y2=2.815
r215 1 26 300 $w=1.7e-07 $l=2.62678e-07 $layer=licon1_PDIFF $count=2 $X=0.665
+ $Y=2.32 $X2=0.865 $Y2=2.465
.ends

.subckt PM_SKY130_FD_SC_HS__SDFXBP_1%A_296_74# 1 2 3 4 13 19 22 23 24 26 27 30
+ 31 32 35 37 38 41 44 45
c131 24 0 6.03804e-20 $X=2.39 $Y=1.265
c132 22 0 2.47416e-20 $X=2.305 $Y=1.18
r133 39 41 2.76586 $w=2.48e-07 $l=6e-08 $layer=LI1_cond $X=5.11 $Y=2.63 $X2=5.11
+ $Y2=2.69
r134 38 46 25.0585 $w=1.94e-07 $l=4.12129e-07 $layer=LI1_cond $X=4.675 $Y=2.545
+ $X2=4.28 $Y2=2.51
r135 37 39 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=4.985 $Y=2.545
+ $X2=5.11 $Y2=2.63
r136 37 38 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=4.985 $Y=2.545
+ $X2=4.675 $Y2=2.545
r137 33 35 32.9599 $w=2.48e-07 $l=7.15e-07 $layer=LI1_cond $X=4.775 $Y=1.48
+ $X2=4.775 $Y2=0.765
r138 31 33 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=4.65 $Y=1.565
+ $X2=4.775 $Y2=1.48
r139 31 32 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=4.65 $Y=1.565
+ $X2=4.365 $Y2=1.565
r140 30 46 1.50975 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=4.28 $Y=2.39
+ $X2=4.28 $Y2=2.51
r141 29 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.28 $Y=1.65
+ $X2=4.365 $Y2=1.565
r142 29 30 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=4.28 $Y=1.65
+ $X2=4.28 $Y2=2.39
r143 28 45 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.065 $Y=2.475
+ $X2=2.98 $Y2=2.475
r144 27 46 5.56362 $w=1.94e-07 $l=1.00995e-07 $layer=LI1_cond $X=4.195 $Y=2.475
+ $X2=4.28 $Y2=2.51
r145 27 28 73.7219 $w=1.68e-07 $l=1.13e-06 $layer=LI1_cond $X=4.195 $Y=2.475
+ $X2=3.065 $Y2=2.475
r146 26 45 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.98 $Y=2.39
+ $X2=2.98 $Y2=2.475
r147 25 26 67.8503 $w=1.68e-07 $l=1.04e-06 $layer=LI1_cond $X=2.98 $Y=1.35
+ $X2=2.98 $Y2=2.39
r148 23 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.895 $Y=1.265
+ $X2=2.98 $Y2=1.35
r149 23 24 32.9465 $w=1.68e-07 $l=5.05e-07 $layer=LI1_cond $X=2.895 $Y=1.265
+ $X2=2.39 $Y2=1.265
r150 22 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.305 $Y=1.18
+ $X2=2.39 $Y2=1.265
r151 21 22 35.2299 $w=1.68e-07 $l=5.4e-07 $layer=LI1_cond $X=2.305 $Y=0.64
+ $X2=2.305 $Y2=1.18
r152 20 44 4.79676 $w=1.7e-07 $l=1.86145e-07 $layer=LI1_cond $X=1.9 $Y=2.475
+ $X2=1.735 $Y2=2.43
r153 19 45 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.895 $Y=2.475
+ $X2=2.98 $Y2=2.475
r154 19 20 64.9144 $w=1.68e-07 $l=9.95e-07 $layer=LI1_cond $X=2.895 $Y=2.475
+ $X2=1.9 $Y2=2.475
r155 13 21 7.14316 $w=2.5e-07 $l=1.62019e-07 $layer=LI1_cond $X=2.22 $Y=0.515
+ $X2=2.305 $Y2=0.64
r156 13 15 21.6659 $w=2.48e-07 $l=4.7e-07 $layer=LI1_cond $X=2.22 $Y=0.515
+ $X2=1.75 $Y2=0.515
r157 4 41 600 $w=1.7e-07 $l=2.67208e-07 $layer=licon1_PDIFF $count=1 $X=5.02
+ $Y=2.48 $X2=5.15 $Y2=2.69
r158 3 44 300 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=2 $X=1.585
+ $Y=2.32 $X2=1.735 $Y2=2.465
r159 2 35 182 $w=1.7e-07 $l=3.25576e-07 $layer=licon1_NDIFF $count=1 $X=4.68
+ $Y=0.5 $X2=4.815 $Y2=0.765
r160 1 15 182 $w=1.7e-07 $l=3.505e-07 $layer=licon1_NDIFF $count=1 $X=1.48
+ $Y=0.37 $X2=1.75 $Y2=0.555
.ends

.subckt PM_SKY130_FD_SC_HS__SDFXBP_1%Q 1 2 7 9 15 16 17 23 29
r30 21 29 0.0555394 $w=4.13e-07 $l=2e-09 $layer=LI1_cond $X=10.707 $Y=0.923
+ $X2=10.707 $Y2=0.925
r31 17 31 8.68557 $w=4.13e-07 $l=1.64e-07 $layer=LI1_cond $X=10.707 $Y=0.966
+ $X2=10.707 $Y2=1.13
r32 17 29 1.13856 $w=4.13e-07 $l=4.1e-08 $layer=LI1_cond $X=10.707 $Y=0.966
+ $X2=10.707 $Y2=0.925
r33 17 21 1.16633 $w=4.13e-07 $l=4.2e-08 $layer=LI1_cond $X=10.707 $Y=0.881
+ $X2=10.707 $Y2=0.923
r34 16 17 9.05293 $w=4.13e-07 $l=3.26e-07 $layer=LI1_cond $X=10.707 $Y=0.555
+ $X2=10.707 $Y2=0.881
r35 16 23 1.11079 $w=4.13e-07 $l=4e-08 $layer=LI1_cond $X=10.707 $Y=0.555
+ $X2=10.707 $Y2=0.515
r36 15 31 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=10.83 $Y=1.82
+ $X2=10.83 $Y2=1.13
r37 9 11 36.0954 $w=2.63e-07 $l=8.3e-07 $layer=LI1_cond $X=10.782 $Y=1.985
+ $X2=10.782 $Y2=2.815
r38 7 15 7.21712 $w=2.63e-07 $l=1.32e-07 $layer=LI1_cond $X=10.782 $Y=1.952
+ $X2=10.782 $Y2=1.82
r39 7 9 1.43512 $w=2.63e-07 $l=3.3e-08 $layer=LI1_cond $X=10.782 $Y=1.952
+ $X2=10.782 $Y2=1.985
r40 2 11 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=10.585
+ $Y=1.84 $X2=10.735 $Y2=2.815
r41 2 9 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=10.585
+ $Y=1.84 $X2=10.735 $Y2=1.985
r42 1 23 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=10.525
+ $Y=0.37 $X2=10.665 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__SDFXBP_1%Q_N 1 2 7 8 9 10 11 12 13 38 47
r19 23 47 1.52529 $w=3.38e-07 $l=4.5e-08 $layer=LI1_cond $X=12.205 $Y=0.88
+ $X2=12.205 $Y2=0.925
r20 12 13 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=12.21 $Y=2.405
+ $X2=12.21 $Y2=2.775
r21 11 38 0.628605 $w=3.28e-07 $l=1.8e-08 $layer=LI1_cond $X=12.21 $Y=1.967
+ $X2=12.21 $Y2=1.985
r22 11 51 6.4171 $w=3.28e-07 $l=1.47e-07 $layer=LI1_cond $X=12.21 $Y=1.967
+ $X2=12.21 $Y2=1.82
r23 11 12 12.3276 $w=3.28e-07 $l=3.53e-07 $layer=LI1_cond $X=12.21 $Y=2.052
+ $X2=12.21 $Y2=2.405
r24 11 38 2.33981 $w=3.28e-07 $l=6.7e-08 $layer=LI1_cond $X=12.21 $Y=2.052
+ $X2=12.21 $Y2=1.985
r25 10 51 8.11948 $w=2.18e-07 $l=1.55e-07 $layer=LI1_cond $X=12.265 $Y=1.665
+ $X2=12.265 $Y2=1.82
r26 9 10 19.382 $w=2.18e-07 $l=3.7e-07 $layer=LI1_cond $X=12.265 $Y=1.295
+ $X2=12.265 $Y2=1.665
r27 9 49 12.834 $w=2.18e-07 $l=2.45e-07 $layer=LI1_cond $X=12.265 $Y=1.295
+ $X2=12.265 $Y2=1.05
r28 8 49 4.99175 $w=3.38e-07 $l=1.05e-07 $layer=LI1_cond $X=12.205 $Y=0.945
+ $X2=12.205 $Y2=1.05
r29 8 47 0.677908 $w=3.38e-07 $l=2e-08 $layer=LI1_cond $X=12.205 $Y=0.945
+ $X2=12.205 $Y2=0.925
r30 8 23 0.677908 $w=3.38e-07 $l=2e-08 $layer=LI1_cond $X=12.205 $Y=0.86
+ $X2=12.205 $Y2=0.88
r31 7 8 11.6939 $w=3.38e-07 $l=3.45e-07 $layer=LI1_cond $X=12.205 $Y=0.515
+ $X2=12.205 $Y2=0.86
r32 2 13 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=12.06
+ $Y=1.84 $X2=12.21 $Y2=2.815
r33 2 38 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=12.06
+ $Y=1.84 $X2=12.21 $Y2=1.985
r34 1 7 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=12.06
+ $Y=0.37 $X2=12.2 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__SDFXBP_1%VGND 1 2 3 4 5 6 7 24 28 30 34 38 42 46 50
+ 55 56 57 59 64 69 74 86 95 96 99 102 105 108 111 114
r142 114 115 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.76 $Y=0
+ $X2=11.76 $Y2=0
r143 111 112 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=0
+ $X2=8.88 $Y2=0
r144 108 109 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=6.48 $Y=0
+ $X2=6.48 $Y2=0
r145 105 106 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r146 103 106 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=0
+ $X2=3.6 $Y2=0
r147 102 103 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0
+ $X2=2.64 $Y2=0
r148 99 100 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r149 96 115 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.24 $Y=0
+ $X2=11.76 $Y2=0
r150 95 96 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.24 $Y=0
+ $X2=12.24 $Y2=0
r151 93 114 9.39981 $w=1.7e-07 $l=1.88e-07 $layer=LI1_cond $X=11.865 $Y=0
+ $X2=11.677 $Y2=0
r152 93 95 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=11.865 $Y=0
+ $X2=12.24 $Y2=0
r153 92 115 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.28 $Y=0
+ $X2=11.76 $Y2=0
r154 91 92 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=11.28 $Y=0
+ $X2=11.28 $Y2=0
r155 89 92 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=10.32 $Y=0
+ $X2=11.28 $Y2=0
r156 88 91 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=10.32 $Y=0 $X2=11.28
+ $Y2=0
r157 88 89 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=10.32 $Y=0
+ $X2=10.32 $Y2=0
r158 86 114 9.39981 $w=1.7e-07 $l=1.87e-07 $layer=LI1_cond $X=11.49 $Y=0
+ $X2=11.677 $Y2=0
r159 86 91 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=11.49 $Y=0
+ $X2=11.28 $Y2=0
r160 85 89 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.84 $Y=0
+ $X2=10.32 $Y2=0
r161 85 112 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=9.84 $Y=0
+ $X2=8.88 $Y2=0
r162 84 85 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.84 $Y=0 $X2=9.84
+ $Y2=0
r163 82 111 13.3456 $w=1.7e-07 $l=3.35e-07 $layer=LI1_cond $X=9.41 $Y=0
+ $X2=9.075 $Y2=0
r164 82 84 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=9.41 $Y=0 $X2=9.84
+ $Y2=0
r165 81 112 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=0 $X2=8.88
+ $Y2=0
r166 80 81 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r167 78 81 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=6.96 $Y=0 $X2=8.4
+ $Y2=0
r168 78 109 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=0
+ $X2=6.48 $Y2=0
r169 77 80 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=6.96 $Y=0 $X2=8.4
+ $Y2=0
r170 77 78 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.96 $Y=0 $X2=6.96
+ $Y2=0
r171 75 108 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.68 $Y=0
+ $X2=6.555 $Y2=0
r172 75 77 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=6.68 $Y=0 $X2=6.96
+ $Y2=0
r173 74 111 13.3456 $w=1.7e-07 $l=3.35e-07 $layer=LI1_cond $X=8.74 $Y=0
+ $X2=9.075 $Y2=0
r174 74 80 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=8.74 $Y=0 $X2=8.4
+ $Y2=0
r175 73 106 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=3.6
+ $Y2=0
r176 72 73 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r177 70 105 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=3.935 $Y=0
+ $X2=3.765 $Y2=0
r178 70 72 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=3.935 $Y=0
+ $X2=4.08 $Y2=0
r179 69 108 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.43 $Y=0
+ $X2=6.555 $Y2=0
r180 69 72 153.316 $w=1.68e-07 $l=2.35e-06 $layer=LI1_cond $X=6.43 $Y=0 $X2=4.08
+ $Y2=0
r181 68 103 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=1.2 $Y=0
+ $X2=2.64 $Y2=0
r182 68 100 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r183 67 68 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r184 65 99 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.965 $Y=0 $X2=0.8
+ $Y2=0
r185 65 67 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=0.965 $Y=0 $X2=1.2
+ $Y2=0
r186 64 102 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.615 $Y=0
+ $X2=2.74 $Y2=0
r187 64 67 92.3155 $w=1.68e-07 $l=1.415e-06 $layer=LI1_cond $X=2.615 $Y=0
+ $X2=1.2 $Y2=0
r188 62 100 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0
+ $X2=0.72 $Y2=0
r189 61 62 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r190 59 99 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.635 $Y=0 $X2=0.8
+ $Y2=0
r191 59 61 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=0.635 $Y=0
+ $X2=0.24 $Y2=0
r192 57 109 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=6.24 $Y=0
+ $X2=6.48 $Y2=0
r193 57 73 0.602067 $w=4.9e-07 $l=2.16e-06 $layer=MET1_cond $X=6.24 $Y=0
+ $X2=4.08 $Y2=0
r194 56 88 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.235 $Y=0
+ $X2=10.32 $Y2=0
r195 55 84 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=10.15 $Y=0 $X2=9.84
+ $Y2=0
r196 55 56 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.15 $Y=0
+ $X2=10.235 $Y2=0
r197 50 52 12.2927 $w=3.73e-07 $l=4e-07 $layer=LI1_cond $X=11.677 $Y=0.515
+ $X2=11.677 $Y2=0.915
r198 48 114 1.28102 $w=3.75e-07 $l=8.5e-08 $layer=LI1_cond $X=11.677 $Y=0.085
+ $X2=11.677 $Y2=0
r199 48 50 13.2147 $w=3.73e-07 $l=4.3e-07 $layer=LI1_cond $X=11.677 $Y=0.085
+ $X2=11.677 $Y2=0.515
r200 44 56 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.235 $Y=0.085
+ $X2=10.235 $Y2=0
r201 44 46 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=10.235 $Y=0.085
+ $X2=10.235 $Y2=0.515
r202 40 111 2.76849 $w=6.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.075 $Y=0.085
+ $X2=9.075 $Y2=0
r203 40 42 8.8367 $w=6.68e-07 $l=4.95e-07 $layer=LI1_cond $X=9.075 $Y=0.085
+ $X2=9.075 $Y2=0.58
r204 36 108 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.555 $Y=0.085
+ $X2=6.555 $Y2=0
r205 36 38 12.4464 $w=2.48e-07 $l=2.7e-07 $layer=LI1_cond $X=6.555 $Y=0.085
+ $X2=6.555 $Y2=0.355
r206 32 105 0.987631 $w=3.4e-07 $l=8.5e-08 $layer=LI1_cond $X=3.765 $Y=0.085
+ $X2=3.765 $Y2=0
r207 32 34 14.2361 $w=3.38e-07 $l=4.2e-07 $layer=LI1_cond $X=3.765 $Y=0.085
+ $X2=3.765 $Y2=0.505
r208 31 102 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.865 $Y=0
+ $X2=2.74 $Y2=0
r209 30 105 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=3.595 $Y=0
+ $X2=3.765 $Y2=0
r210 30 31 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=3.595 $Y=0
+ $X2=2.865 $Y2=0
r211 26 102 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.74 $Y=0.085
+ $X2=2.74 $Y2=0
r212 26 28 22.8184 $w=2.48e-07 $l=4.95e-07 $layer=LI1_cond $X=2.74 $Y=0.085
+ $X2=2.74 $Y2=0.58
r213 22 99 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.8 $Y=0.085 $X2=0.8
+ $Y2=0
r214 22 24 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=0.8 $Y=0.085
+ $X2=0.8 $Y2=0.58
r215 7 52 182 $w=1.7e-07 $l=5.18869e-07 $layer=licon1_NDIFF $count=1 $X=11.515
+ $Y=0.47 $X2=11.675 $Y2=0.915
r216 7 50 182 $w=1.7e-07 $l=2.56515e-07 $layer=licon1_NDIFF $count=1 $X=11.515
+ $Y=0.47 $X2=11.75 $Y2=0.515
r217 6 46 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=10.09
+ $Y=0.37 $X2=10.235 $Y2=0.515
r218 5 42 91 $w=1.7e-07 $l=5.755e-07 $layer=licon1_NDIFF $count=2 $X=8.765
+ $Y=0.37 $X2=9.245 $Y2=0.58
r219 4 38 182 $w=1.7e-07 $l=2.62678e-07 $layer=licon1_NDIFF $count=1 $X=6.395
+ $Y=0.5 $X2=6.595 $Y2=0.355
r220 3 34 182 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_NDIFF $count=1 $X=3.615
+ $Y=0.36 $X2=3.765 $Y2=0.505
r221 2 28 182 $w=1.7e-07 $l=2.86182e-07 $layer=licon1_NDIFF $count=1 $X=2.56
+ $Y=0.37 $X2=2.74 $Y2=0.58
r222 1 24 182 $w=1.7e-07 $l=2.96985e-07 $layer=licon1_NDIFF $count=1 $X=0.59
+ $Y=0.37 $X2=0.8 $Y2=0.58
.ends

