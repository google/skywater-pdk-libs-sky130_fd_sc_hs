* File: sky130_fd_sc_hs__and2b_1.pxi.spice
* Created: Thu Aug 27 20:31:53 2020
* 
x_PM_SKY130_FD_SC_HS__AND2B_1%A_N N_A_N_M1007_g N_A_N_c_62_n N_A_N_c_66_n
+ N_A_N_M1002_g A_N A_N N_A_N_c_63_n N_A_N_c_64_n
+ PM_SKY130_FD_SC_HS__AND2B_1%A_N
x_PM_SKY130_FD_SC_HS__AND2B_1%A_27_74# N_A_27_74#_M1007_s N_A_27_74#_M1002_s
+ N_A_27_74#_c_97_n N_A_27_74#_c_98_n N_A_27_74#_c_107_n N_A_27_74#_M1003_g
+ N_A_27_74#_c_99_n N_A_27_74#_M1001_g N_A_27_74#_c_100_n N_A_27_74#_c_101_n
+ N_A_27_74#_c_108_n N_A_27_74#_c_102_n N_A_27_74#_c_103_n N_A_27_74#_c_122_n
+ N_A_27_74#_c_104_n N_A_27_74#_c_105_n PM_SKY130_FD_SC_HS__AND2B_1%A_27_74#
x_PM_SKY130_FD_SC_HS__AND2B_1%B N_B_M1000_g N_B_c_166_n N_B_M1005_g B
+ N_B_c_167_n PM_SKY130_FD_SC_HS__AND2B_1%B
x_PM_SKY130_FD_SC_HS__AND2B_1%A_266_98# N_A_266_98#_M1001_s N_A_266_98#_M1003_d
+ N_A_266_98#_c_199_n N_A_266_98#_M1006_g N_A_266_98#_M1004_g
+ N_A_266_98#_c_201_n N_A_266_98#_c_202_n N_A_266_98#_c_203_n
+ N_A_266_98#_c_204_n N_A_266_98#_c_208_n N_A_266_98#_c_205_n
+ N_A_266_98#_c_206_n PM_SKY130_FD_SC_HS__AND2B_1%A_266_98#
x_PM_SKY130_FD_SC_HS__AND2B_1%VPWR N_VPWR_M1002_d N_VPWR_M1005_d N_VPWR_c_273_n
+ N_VPWR_c_274_n N_VPWR_c_275_n N_VPWR_c_276_n N_VPWR_c_277_n N_VPWR_c_278_n
+ VPWR N_VPWR_c_279_n N_VPWR_c_272_n PM_SKY130_FD_SC_HS__AND2B_1%VPWR
x_PM_SKY130_FD_SC_HS__AND2B_1%X N_X_M1004_d N_X_M1006_d N_X_c_310_n N_X_c_311_n
+ X X X N_X_c_314_n N_X_c_312_n X PM_SKY130_FD_SC_HS__AND2B_1%X
x_PM_SKY130_FD_SC_HS__AND2B_1%VGND N_VGND_M1007_d N_VGND_M1000_d N_VGND_c_333_n
+ N_VGND_c_334_n VGND N_VGND_c_335_n N_VGND_c_336_n N_VGND_c_337_n
+ N_VGND_c_338_n N_VGND_c_339_n N_VGND_c_340_n PM_SKY130_FD_SC_HS__AND2B_1%VGND
cc_1 VNB N_A_N_M1007_g 0.0473335f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.645
cc_2 VNB N_A_N_c_62_n 0.0192462f $X=-0.19 $Y=-0.245 $X2=1.135 $Y2=1.675
cc_3 VNB N_A_N_c_63_n 0.0323686f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.515
cc_4 VNB N_A_N_c_64_n 0.0146719f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.515
cc_5 VNB N_A_27_74#_c_97_n 0.0332487f $X=-0.19 $Y=-0.245 $X2=1.225 $Y2=1.765
cc_6 VNB N_A_27_74#_c_98_n 0.016924f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_7 VNB N_A_27_74#_c_99_n 0.016514f $X=-0.19 $Y=-0.245 $X2=0.395 $Y2=1.515
cc_8 VNB N_A_27_74#_c_100_n 0.00534155f $X=-0.19 $Y=-0.245 $X2=0.395 $Y2=1.35
cc_9 VNB N_A_27_74#_c_101_n 0.0280542f $X=-0.19 $Y=-0.245 $X2=0.337 $Y2=1.515
cc_10 VNB N_A_27_74#_c_102_n 0.0167838f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_27_74#_c_103_n 0.0102182f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_27_74#_c_104_n 0.0043967f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_27_74#_c_105_n 0.033482f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_B_M1000_g 0.0247191f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.645
cc_15 VNB N_B_c_166_n 0.029118f $X=-0.19 $Y=-0.245 $X2=1.135 $Y2=1.675
cc_16 VNB N_B_c_167_n 0.00215995f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_266_98#_c_199_n 0.0367215f $X=-0.19 $Y=-0.245 $X2=1.225 $Y2=1.765
cc_18 VNB N_A_266_98#_M1004_g 0.028553f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_266_98#_c_201_n 0.0134821f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.515
cc_20 VNB N_A_266_98#_c_202_n 0.0129986f $X=-0.19 $Y=-0.245 $X2=0.337 $Y2=1.665
cc_21 VNB N_A_266_98#_c_203_n 0.0054423f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_266_98#_c_204_n 0.00336141f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_266_98#_c_205_n 0.00401614f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_266_98#_c_206_n 0.00245262f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_VPWR_c_272_n 0.143779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_X_c_310_n 0.026297f $X=-0.19 $Y=-0.245 $X2=1.225 $Y2=2.26
cc_27 VNB N_X_c_311_n 0.00881925f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_X_c_312_n 0.023581f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_333_n 0.0189444f $X=-0.19 $Y=-0.245 $X2=1.225 $Y2=2.26
cc_30 VNB N_VGND_c_334_n 0.0166279f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_335_n 0.0191515f $X=-0.19 $Y=-0.245 $X2=0.395 $Y2=1.675
cc_32 VNB N_VGND_c_336_n 0.0356214f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_337_n 0.0191749f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_338_n 0.232503f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_339_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_340_n 0.0118294f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VPB N_A_N_c_62_n 0.0271915f $X=-0.19 $Y=1.66 $X2=1.135 $Y2=1.675
cc_38 VPB N_A_N_c_66_n 0.0196782f $X=-0.19 $Y=1.66 $X2=1.225 $Y2=1.765
cc_39 VPB N_A_N_c_63_n 0.0160383f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.515
cc_40 VPB N_A_N_c_64_n 0.0197858f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.515
cc_41 VPB N_A_27_74#_c_98_n 6.93665e-19 $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_42 VPB N_A_27_74#_c_107_n 0.02128f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.95
cc_43 VPB N_A_27_74#_c_108_n 0.0143702f $X=-0.19 $Y=1.66 $X2=0.337 $Y2=1.665
cc_44 VPB N_A_27_74#_c_104_n 0.00159553f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_45 VPB N_B_c_166_n 0.0289588f $X=-0.19 $Y=1.66 $X2=1.135 $Y2=1.675
cc_46 VPB N_B_c_167_n 0.00489452f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_47 VPB N_A_266_98#_c_199_n 0.029602f $X=-0.19 $Y=1.66 $X2=1.225 $Y2=1.765
cc_48 VPB N_A_266_98#_c_208_n 0.00394633f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_49 VPB N_A_266_98#_c_205_n 0.00129478f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_50 VPB N_VPWR_c_273_n 0.0311212f $X=-0.19 $Y=1.66 $X2=1.225 $Y2=2.26
cc_51 VPB N_VPWR_c_274_n 0.0202787f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_52 VPB N_VPWR_c_275_n 0.0413121f $X=-0.19 $Y=1.66 $X2=0.395 $Y2=1.675
cc_53 VPB N_VPWR_c_276_n 0.00324402f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_54 VPB N_VPWR_c_277_n 0.0217159f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_55 VPB N_VPWR_c_278_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0.337 $Y2=1.665
cc_56 VPB N_VPWR_c_279_n 0.0225548f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_57 VPB N_VPWR_c_272_n 0.0820446f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_58 VPB X 0.0458336f $X=-0.19 $Y=1.66 $X2=0.395 $Y2=1.515
cc_59 VPB N_X_c_314_n 0.0142631f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_60 VPB N_X_c_312_n 0.00786764f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_61 N_A_N_c_64_n N_A_27_74#_M1002_s 0.0133535f $X=0.385 $Y=1.515 $X2=0 $Y2=0
cc_62 N_A_N_c_62_n N_A_27_74#_c_98_n 0.00796509f $X=1.135 $Y=1.675 $X2=0 $Y2=0
cc_63 N_A_N_c_66_n N_A_27_74#_c_107_n 0.0118449f $X=1.225 $Y=1.765 $X2=0 $Y2=0
cc_64 N_A_N_M1007_g N_A_27_74#_c_101_n 0.0182367f $X=0.495 $Y=0.645 $X2=0 $Y2=0
cc_65 N_A_N_c_63_n N_A_27_74#_c_108_n 0.00752285f $X=0.385 $Y=1.515 $X2=0 $Y2=0
cc_66 N_A_N_c_64_n N_A_27_74#_c_108_n 0.036054f $X=0.385 $Y=1.515 $X2=0 $Y2=0
cc_67 N_A_N_M1007_g N_A_27_74#_c_102_n 0.0116944f $X=0.495 $Y=0.645 $X2=0 $Y2=0
cc_68 N_A_N_c_62_n N_A_27_74#_c_102_n 0.00628292f $X=1.135 $Y=1.675 $X2=0 $Y2=0
cc_69 N_A_N_c_64_n N_A_27_74#_c_102_n 0.00788818f $X=0.385 $Y=1.515 $X2=0 $Y2=0
cc_70 N_A_N_M1007_g N_A_27_74#_c_103_n 0.00419608f $X=0.495 $Y=0.645 $X2=0 $Y2=0
cc_71 N_A_N_c_63_n N_A_27_74#_c_103_n 0.00157825f $X=0.385 $Y=1.515 $X2=0 $Y2=0
cc_72 N_A_N_c_64_n N_A_27_74#_c_103_n 0.0287548f $X=0.385 $Y=1.515 $X2=0 $Y2=0
cc_73 N_A_N_c_66_n N_A_27_74#_c_122_n 0.00429418f $X=1.225 $Y=1.765 $X2=0 $Y2=0
cc_74 N_A_N_M1007_g N_A_27_74#_c_104_n 0.00113276f $X=0.495 $Y=0.645 $X2=0 $Y2=0
cc_75 N_A_N_c_62_n N_A_27_74#_c_104_n 0.0214709f $X=1.135 $Y=1.675 $X2=0 $Y2=0
cc_76 N_A_N_c_66_n N_A_27_74#_c_104_n 0.0111792f $X=1.225 $Y=1.765 $X2=0 $Y2=0
cc_77 N_A_N_c_63_n N_A_27_74#_c_104_n 0.00535237f $X=0.385 $Y=1.515 $X2=0 $Y2=0
cc_78 N_A_N_c_64_n N_A_27_74#_c_104_n 0.0470333f $X=0.385 $Y=1.515 $X2=0 $Y2=0
cc_79 N_A_N_M1007_g N_A_27_74#_c_105_n 0.018827f $X=0.495 $Y=0.645 $X2=0 $Y2=0
cc_80 N_A_N_c_62_n N_A_27_74#_c_105_n 0.0294207f $X=1.135 $Y=1.675 $X2=0 $Y2=0
cc_81 N_A_N_c_62_n N_A_266_98#_c_205_n 6.37275e-19 $X=1.135 $Y=1.675 $X2=0 $Y2=0
cc_82 N_A_N_c_66_n N_A_266_98#_c_205_n 4.18137e-19 $X=1.225 $Y=1.765 $X2=0 $Y2=0
cc_83 N_A_N_c_66_n N_VPWR_c_273_n 0.00725845f $X=1.225 $Y=1.765 $X2=0 $Y2=0
cc_84 N_A_N_c_66_n N_VPWR_c_275_n 0.00393546f $X=1.225 $Y=1.765 $X2=0 $Y2=0
cc_85 N_A_N_c_66_n N_VPWR_c_272_n 0.00462577f $X=1.225 $Y=1.765 $X2=0 $Y2=0
cc_86 N_A_N_M1007_g N_VGND_c_333_n 0.0141934f $X=0.495 $Y=0.645 $X2=0 $Y2=0
cc_87 N_A_N_M1007_g N_VGND_c_335_n 0.00434272f $X=0.495 $Y=0.645 $X2=0 $Y2=0
cc_88 N_A_N_M1007_g N_VGND_c_338_n 0.00828717f $X=0.495 $Y=0.645 $X2=0 $Y2=0
cc_89 N_A_27_74#_c_99_n N_B_M1000_g 0.0339588f $X=1.69 $Y=1.21 $X2=0 $Y2=0
cc_90 N_A_27_74#_c_98_n N_B_c_166_n 0.0339588f $X=1.675 $Y=1.675 $X2=0 $Y2=0
cc_91 N_A_27_74#_c_107_n N_B_c_166_n 0.0157645f $X=1.675 $Y=1.765 $X2=0 $Y2=0
cc_92 N_A_27_74#_c_100_n N_B_c_167_n 4.08878e-19 $X=1.675 $Y=1.285 $X2=0 $Y2=0
cc_93 N_A_27_74#_c_99_n N_A_266_98#_c_201_n 0.00940974f $X=1.69 $Y=1.21 $X2=0
+ $Y2=0
cc_94 N_A_27_74#_c_97_n N_A_266_98#_c_203_n 0.0101577f $X=1.585 $Y=1.285 $X2=0
+ $Y2=0
cc_95 N_A_27_74#_c_99_n N_A_266_98#_c_203_n 0.0140365f $X=1.69 $Y=1.21 $X2=0
+ $Y2=0
cc_96 N_A_27_74#_c_102_n N_A_266_98#_c_203_n 0.0124833f $X=0.81 $Y=1.095 $X2=0
+ $Y2=0
cc_97 N_A_27_74#_c_105_n N_A_266_98#_c_203_n 5.41958e-19 $X=0.975 $Y=1.195 $X2=0
+ $Y2=0
cc_98 N_A_27_74#_c_107_n N_A_266_98#_c_208_n 0.0099463f $X=1.675 $Y=1.765 $X2=0
+ $Y2=0
cc_99 N_A_27_74#_c_98_n N_A_266_98#_c_205_n 0.00887025f $X=1.675 $Y=1.675 $X2=0
+ $Y2=0
cc_100 N_A_27_74#_c_107_n N_A_266_98#_c_205_n 0.00649341f $X=1.675 $Y=1.765
+ $X2=0 $Y2=0
cc_101 N_A_27_74#_c_99_n N_A_266_98#_c_205_n 0.00176326f $X=1.69 $Y=1.21 $X2=0
+ $Y2=0
cc_102 N_A_27_74#_c_100_n N_A_266_98#_c_205_n 0.00560709f $X=1.675 $Y=1.285
+ $X2=0 $Y2=0
cc_103 N_A_27_74#_c_102_n N_A_266_98#_c_205_n 8.47818e-19 $X=0.81 $Y=1.095 $X2=0
+ $Y2=0
cc_104 N_A_27_74#_c_104_n N_A_266_98#_c_205_n 0.018139f $X=0.975 $Y=1.195 $X2=0
+ $Y2=0
cc_105 N_A_27_74#_c_97_n N_VPWR_c_273_n 0.00310442f $X=1.585 $Y=1.285 $X2=0
+ $Y2=0
cc_106 N_A_27_74#_c_107_n N_VPWR_c_273_n 0.00589047f $X=1.675 $Y=1.765 $X2=0
+ $Y2=0
cc_107 N_A_27_74#_c_122_n N_VPWR_c_273_n 0.0228589f $X=0.975 $Y=2.32 $X2=0 $Y2=0
cc_108 N_A_27_74#_c_104_n N_VPWR_c_273_n 0.0154361f $X=0.975 $Y=1.195 $X2=0
+ $Y2=0
cc_109 N_A_27_74#_c_108_n N_VPWR_c_275_n 0.0115433f $X=0.81 $Y=2.485 $X2=0 $Y2=0
cc_110 N_A_27_74#_c_122_n N_VPWR_c_275_n 0.00567516f $X=0.975 $Y=2.32 $X2=0
+ $Y2=0
cc_111 N_A_27_74#_c_107_n N_VPWR_c_277_n 0.00375627f $X=1.675 $Y=1.765 $X2=0
+ $Y2=0
cc_112 N_A_27_74#_c_107_n N_VPWR_c_272_n 0.00462577f $X=1.675 $Y=1.765 $X2=0
+ $Y2=0
cc_113 N_A_27_74#_c_108_n N_VPWR_c_272_n 0.0197081f $X=0.81 $Y=2.485 $X2=0 $Y2=0
cc_114 N_A_27_74#_c_122_n N_VPWR_c_272_n 0.0103466f $X=0.975 $Y=2.32 $X2=0 $Y2=0
cc_115 N_A_27_74#_c_99_n N_VGND_c_333_n 0.0032597f $X=1.69 $Y=1.21 $X2=0 $Y2=0
cc_116 N_A_27_74#_c_101_n N_VGND_c_333_n 0.0191765f $X=0.28 $Y=0.645 $X2=0 $Y2=0
cc_117 N_A_27_74#_c_102_n N_VGND_c_333_n 0.027862f $X=0.81 $Y=1.095 $X2=0 $Y2=0
cc_118 N_A_27_74#_c_105_n N_VGND_c_333_n 0.00100291f $X=0.975 $Y=1.195 $X2=0
+ $Y2=0
cc_119 N_A_27_74#_c_99_n N_VGND_c_334_n 0.0014983f $X=1.69 $Y=1.21 $X2=0 $Y2=0
cc_120 N_A_27_74#_c_101_n N_VGND_c_335_n 0.0145639f $X=0.28 $Y=0.645 $X2=0 $Y2=0
cc_121 N_A_27_74#_c_99_n N_VGND_c_336_n 0.00473385f $X=1.69 $Y=1.21 $X2=0 $Y2=0
cc_122 N_A_27_74#_c_99_n N_VGND_c_338_n 0.00508379f $X=1.69 $Y=1.21 $X2=0 $Y2=0
cc_123 N_A_27_74#_c_101_n N_VGND_c_338_n 0.0119984f $X=0.28 $Y=0.645 $X2=0 $Y2=0
cc_124 N_B_M1000_g N_A_266_98#_c_199_n 7.12296e-19 $X=2.08 $Y=0.81 $X2=0 $Y2=0
cc_125 N_B_c_166_n N_A_266_98#_c_199_n 0.0437166f $X=2.125 $Y=1.765 $X2=0 $Y2=0
cc_126 N_B_c_167_n N_A_266_98#_c_199_n 0.00283767f $X=2.21 $Y=1.515 $X2=0 $Y2=0
cc_127 N_B_M1000_g N_A_266_98#_M1004_g 0.00824273f $X=2.08 $Y=0.81 $X2=0 $Y2=0
cc_128 N_B_M1000_g N_A_266_98#_c_201_n 0.00180506f $X=2.08 $Y=0.81 $X2=0 $Y2=0
cc_129 N_B_M1000_g N_A_266_98#_c_202_n 0.0163783f $X=2.08 $Y=0.81 $X2=0 $Y2=0
cc_130 N_B_c_166_n N_A_266_98#_c_202_n 0.00148677f $X=2.125 $Y=1.765 $X2=0 $Y2=0
cc_131 N_B_c_167_n N_A_266_98#_c_202_n 0.0219406f $X=2.21 $Y=1.515 $X2=0 $Y2=0
cc_132 N_B_M1000_g N_A_266_98#_c_204_n 0.00297924f $X=2.08 $Y=0.81 $X2=0 $Y2=0
cc_133 N_B_c_166_n N_A_266_98#_c_208_n 0.0088849f $X=2.125 $Y=1.765 $X2=0 $Y2=0
cc_134 N_B_c_167_n N_A_266_98#_c_208_n 0.00127779f $X=2.21 $Y=1.515 $X2=0 $Y2=0
cc_135 N_B_M1000_g N_A_266_98#_c_205_n 0.00630861f $X=2.08 $Y=0.81 $X2=0 $Y2=0
cc_136 N_B_c_166_n N_A_266_98#_c_205_n 0.00393624f $X=2.125 $Y=1.765 $X2=0 $Y2=0
cc_137 N_B_c_167_n N_A_266_98#_c_205_n 0.0323775f $X=2.21 $Y=1.515 $X2=0 $Y2=0
cc_138 N_B_M1000_g N_A_266_98#_c_206_n 5.40545e-19 $X=2.08 $Y=0.81 $X2=0 $Y2=0
cc_139 N_B_c_166_n N_A_266_98#_c_206_n 0.00173367f $X=2.125 $Y=1.765 $X2=0 $Y2=0
cc_140 N_B_c_167_n N_A_266_98#_c_206_n 0.0210902f $X=2.21 $Y=1.515 $X2=0 $Y2=0
cc_141 N_B_c_166_n N_VPWR_c_274_n 0.0110134f $X=2.125 $Y=1.765 $X2=0 $Y2=0
cc_142 N_B_c_167_n N_VPWR_c_274_n 0.00914737f $X=2.21 $Y=1.515 $X2=0 $Y2=0
cc_143 N_B_c_166_n N_VPWR_c_277_n 0.00393873f $X=2.125 $Y=1.765 $X2=0 $Y2=0
cc_144 N_B_c_166_n N_VPWR_c_272_n 0.00462577f $X=2.125 $Y=1.765 $X2=0 $Y2=0
cc_145 N_B_c_166_n N_X_c_314_n 7.36066e-19 $X=2.125 $Y=1.765 $X2=0 $Y2=0
cc_146 N_B_M1000_g N_VGND_c_334_n 0.0110841f $X=2.08 $Y=0.81 $X2=0 $Y2=0
cc_147 N_B_M1000_g N_VGND_c_336_n 0.00410575f $X=2.08 $Y=0.81 $X2=0 $Y2=0
cc_148 N_B_M1000_g N_VGND_c_338_n 0.00427039f $X=2.08 $Y=0.81 $X2=0 $Y2=0
cc_149 N_A_266_98#_c_203_n N_VPWR_c_273_n 0.00536405f $X=1.875 $Y=1.065 $X2=0
+ $Y2=0
cc_150 N_A_266_98#_c_205_n N_VPWR_c_273_n 0.0648615f $X=1.885 $Y=1.95 $X2=0
+ $Y2=0
cc_151 N_A_266_98#_c_199_n N_VPWR_c_274_n 0.0135717f $X=2.71 $Y=1.765 $X2=0
+ $Y2=0
cc_152 N_A_266_98#_c_208_n N_VPWR_c_274_n 0.0507312f $X=1.9 $Y=2.115 $X2=0 $Y2=0
cc_153 N_A_266_98#_c_206_n N_VPWR_c_274_n 7.04423e-19 $X=2.75 $Y=1.485 $X2=0
+ $Y2=0
cc_154 N_A_266_98#_c_208_n N_VPWR_c_277_n 0.00719065f $X=1.9 $Y=2.115 $X2=0
+ $Y2=0
cc_155 N_A_266_98#_c_199_n N_VPWR_c_279_n 0.00445602f $X=2.71 $Y=1.765 $X2=0
+ $Y2=0
cc_156 N_A_266_98#_c_199_n N_VPWR_c_272_n 0.00865604f $X=2.71 $Y=1.765 $X2=0
+ $Y2=0
cc_157 N_A_266_98#_c_208_n N_VPWR_c_272_n 0.010834f $X=1.9 $Y=2.115 $X2=0 $Y2=0
cc_158 N_A_266_98#_M1004_g N_X_c_310_n 0.0138984f $X=2.865 $Y=0.76 $X2=0 $Y2=0
cc_159 N_A_266_98#_M1004_g N_X_c_311_n 0.00281566f $X=2.865 $Y=0.76 $X2=0 $Y2=0
cc_160 N_A_266_98#_c_202_n N_X_c_311_n 0.00732422f $X=2.575 $Y=1.065 $X2=0 $Y2=0
cc_161 N_A_266_98#_c_199_n X 0.0105773f $X=2.71 $Y=1.765 $X2=0 $Y2=0
cc_162 N_A_266_98#_c_199_n N_X_c_314_n 0.00885445f $X=2.71 $Y=1.765 $X2=0 $Y2=0
cc_163 N_A_266_98#_c_206_n N_X_c_314_n 0.0120807f $X=2.75 $Y=1.485 $X2=0 $Y2=0
cc_164 N_A_266_98#_c_199_n N_X_c_312_n 0.00368867f $X=2.71 $Y=1.765 $X2=0 $Y2=0
cc_165 N_A_266_98#_M1004_g N_X_c_312_n 0.0103424f $X=2.865 $Y=0.76 $X2=0 $Y2=0
cc_166 N_A_266_98#_c_204_n N_X_c_312_n 0.00557533f $X=2.66 $Y=1.32 $X2=0 $Y2=0
cc_167 N_A_266_98#_c_206_n N_X_c_312_n 0.0248284f $X=2.75 $Y=1.485 $X2=0 $Y2=0
cc_168 N_A_266_98#_c_202_n N_VGND_M1000_d 0.00883207f $X=2.575 $Y=1.065 $X2=0
+ $Y2=0
cc_169 N_A_266_98#_c_201_n N_VGND_c_333_n 0.0181686f $X=1.475 $Y=0.635 $X2=0
+ $Y2=0
cc_170 N_A_266_98#_c_199_n N_VGND_c_334_n 5.91326e-19 $X=2.71 $Y=1.765 $X2=0
+ $Y2=0
cc_171 N_A_266_98#_M1004_g N_VGND_c_334_n 0.00570254f $X=2.865 $Y=0.76 $X2=0
+ $Y2=0
cc_172 N_A_266_98#_c_201_n N_VGND_c_334_n 0.0113091f $X=1.475 $Y=0.635 $X2=0
+ $Y2=0
cc_173 N_A_266_98#_c_202_n N_VGND_c_334_n 0.0448368f $X=2.575 $Y=1.065 $X2=0
+ $Y2=0
cc_174 N_A_266_98#_c_201_n N_VGND_c_336_n 0.00957354f $X=1.475 $Y=0.635 $X2=0
+ $Y2=0
cc_175 N_A_266_98#_M1004_g N_VGND_c_337_n 0.00537471f $X=2.865 $Y=0.76 $X2=0
+ $Y2=0
cc_176 N_A_266_98#_M1004_g N_VGND_c_338_n 0.00539454f $X=2.865 $Y=0.76 $X2=0
+ $Y2=0
cc_177 N_A_266_98#_c_201_n N_VGND_c_338_n 0.0110524f $X=1.475 $Y=0.635 $X2=0
+ $Y2=0
cc_178 N_A_266_98#_c_202_n A_353_98# 0.0027472f $X=2.575 $Y=1.065 $X2=-0.19
+ $Y2=-0.245
cc_179 N_A_266_98#_c_203_n A_353_98# 0.00202224f $X=1.875 $Y=1.065 $X2=-0.19
+ $Y2=-0.245
cc_180 N_VPWR_c_279_n X 0.0215101f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_181 N_VPWR_c_272_n X 0.0177713f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_182 N_VPWR_c_274_n N_X_c_314_n 0.0417431f $X=2.435 $Y=2.045 $X2=0 $Y2=0
cc_183 N_X_c_310_n N_VGND_c_334_n 0.0174539f $X=3.08 $Y=0.535 $X2=0 $Y2=0
cc_184 N_X_c_310_n N_VGND_c_337_n 0.0138903f $X=3.08 $Y=0.535 $X2=0 $Y2=0
cc_185 N_X_c_310_n N_VGND_c_338_n 0.0123115f $X=3.08 $Y=0.535 $X2=0 $Y2=0
