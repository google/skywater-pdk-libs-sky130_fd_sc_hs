* File: sky130_fd_sc_hs__a32o_1.pex.spice
* Created: Thu Aug 27 20:29:56 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HS__A32O_1%A_84_48# 1 2 9 11 13 15 17 18 22 27 31 32
r83 31 32 17.1863 $w=5.88e-07 $l=5.15e-07 $layer=LI1_cond $X=2.715 $Y=0.725
+ $X2=2.2 $Y2=0.725
r84 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.59
+ $Y=1.465 $X2=0.59 $Y2=1.465
r85 22 24 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=3.06 $Y=1.97
+ $X2=3.06 $Y2=2.65
r86 20 22 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=3.06 $Y=1.89 $X2=3.06
+ $Y2=1.97
r87 19 27 14.7616 $w=2.81e-07 $l=4.22493e-07 $layer=LI1_cond $X=0.795 $Y=1.805
+ $X2=0.61 $Y2=1.465
r88 18 20 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.895 $Y=1.805
+ $X2=3.06 $Y2=1.89
r89 18 19 137.005 $w=1.68e-07 $l=2.1e-06 $layer=LI1_cond $X=2.895 $Y=1.805
+ $X2=0.795 $Y2=1.805
r90 17 32 91.6631 $w=1.68e-07 $l=1.405e-06 $layer=LI1_cond $X=0.795 $Y=0.935
+ $X2=2.2 $Y2=0.935
r91 15 27 9.05323 $w=2.81e-07 $l=2.09105e-07 $layer=LI1_cond $X=0.71 $Y=1.3
+ $X2=0.61 $Y2=1.465
r92 14 17 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.71 $Y=1.02
+ $X2=0.795 $Y2=0.935
r93 14 15 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=0.71 $Y=1.02
+ $X2=0.71 $Y2=1.3
r94 11 28 61.0536 $w=2.9e-07 $l=3.34066e-07 $layer=POLY_cond $X=0.515 $Y=1.765
+ $X2=0.587 $Y2=1.465
r95 11 13 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.515 $Y=1.765
+ $X2=0.515 $Y2=2.4
r96 7 28 38.6157 $w=2.9e-07 $l=2.05925e-07 $layer=POLY_cond $X=0.495 $Y=1.3
+ $X2=0.587 $Y2=1.465
r97 7 9 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=0.495 $Y=1.3 $X2=0.495
+ $Y2=0.74
r98 2 24 400 $w=1.7e-07 $l=9.04489e-07 $layer=licon1_PDIFF $count=1 $X=2.86
+ $Y=1.84 $X2=3.06 $Y2=2.65
r99 2 22 400 $w=1.7e-07 $l=2.56905e-07 $layer=licon1_PDIFF $count=1 $X=2.86
+ $Y=1.84 $X2=3.06 $Y2=1.97
r100 1 31 45.5 $w=1.7e-07 $l=5.48954e-07 $layer=licon1_NDIFF $count=4 $X=2.225
+ $Y=0.47 $X2=2.715 $Y2=0.595
.ends

.subckt PM_SKY130_FD_SC_HS__A32O_1%A3 1 3 4 6 7
c31 7 0 9.8332e-20 $X=1.2 $Y=1.295
c32 4 0 9.95713e-20 $X=1.22 $Y=1.22
r33 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.13
+ $Y=1.385 $X2=1.13 $Y2=1.385
r34 7 11 2.96342 $w=3.48e-07 $l=9e-08 $layer=LI1_cond $X=1.14 $Y=1.295 $X2=1.14
+ $Y2=1.385
r35 4 10 38.9026 $w=2.7e-07 $l=2.05122e-07 $layer=POLY_cond $X=1.22 $Y=1.22
+ $X2=1.13 $Y2=1.385
r36 4 6 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=1.22 $Y=1.22 $X2=1.22
+ $Y2=0.79
r37 1 10 77.2841 $w=2.7e-07 $l=3.87427e-07 $layer=POLY_cond $X=1.145 $Y=1.765
+ $X2=1.13 $Y2=1.385
r38 1 3 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=1.145 $Y=1.765
+ $X2=1.145 $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_HS__A32O_1%A2 1 3 4 6 7
c27 7 0 2.09874e-19 $X=1.68 $Y=1.295
c28 4 0 1.83337e-19 $X=1.61 $Y=1.22
r29 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.67
+ $Y=1.385 $X2=1.67 $Y2=1.385
r30 7 11 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=1.67 $Y=1.295 $X2=1.67
+ $Y2=1.385
r31 4 10 38.9026 $w=2.7e-07 $l=1.92678e-07 $layer=POLY_cond $X=1.61 $Y=1.22
+ $X2=1.67 $Y2=1.385
r32 4 6 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=1.61 $Y=1.22 $X2=1.61
+ $Y2=0.79
r33 1 10 77.2841 $w=2.7e-07 $l=4.15812e-07 $layer=POLY_cond $X=1.595 $Y=1.765
+ $X2=1.67 $Y2=1.385
r34 1 3 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=1.595 $Y=1.765
+ $X2=1.595 $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_HS__A32O_1%A1 1 3 4 6 7
c29 7 0 1.47811e-19 $X=2.16 $Y=1.295
c30 1 0 2.02667e-19 $X=2.15 $Y=1.22
r31 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.21
+ $Y=1.385 $X2=2.21 $Y2=1.385
r32 7 11 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=2.21 $Y=1.295 $X2=2.21
+ $Y2=1.385
r33 4 10 72.9766 $w=3.01e-07 $l=4.27083e-07 $layer=POLY_cond $X=2.335 $Y=1.765
+ $X2=2.235 $Y2=1.385
r34 4 6 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=2.335 $Y=1.765
+ $X2=2.335 $Y2=2.34
r35 1 10 38.5481 $w=3.01e-07 $l=2.03101e-07 $layer=POLY_cond $X=2.15 $Y=1.22
+ $X2=2.235 $Y2=1.385
r36 1 3 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=2.15 $Y=1.22 $X2=2.15
+ $Y2=0.79
.ends

.subckt PM_SKY130_FD_SC_HS__A32O_1%B1 1 3 4 6 7 11
c28 11 0 9.23649e-20 $X=2.84 $Y=1.385
c29 4 0 6.28053e-20 $X=2.93 $Y=1.22
r30 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.84
+ $Y=1.385 $X2=2.84 $Y2=1.385
r31 7 11 6.40246 $w=3.58e-07 $l=2e-07 $layer=LI1_cond $X=2.64 $Y=1.37 $X2=2.84
+ $Y2=1.37
r32 4 10 38.9026 $w=2.7e-07 $l=2.05122e-07 $layer=POLY_cond $X=2.93 $Y=1.22
+ $X2=2.84 $Y2=1.385
r33 4 6 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=2.93 $Y=1.22 $X2=2.93
+ $Y2=0.79
r34 1 10 77.2841 $w=2.7e-07 $l=4.06571e-07 $layer=POLY_cond $X=2.785 $Y=1.765
+ $X2=2.84 $Y2=1.385
r35 1 3 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=2.785 $Y=1.765
+ $X2=2.785 $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_HS__A32O_1%B2 1 3 4 6 7
r21 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.455
+ $Y=1.385 $X2=3.455 $Y2=1.385
r22 7 11 4.91483 $w=3.38e-07 $l=1.45e-07 $layer=LI1_cond $X=3.6 $Y=1.38
+ $X2=3.455 $Y2=1.38
r23 4 10 73.3362 $w=2.98e-07 $l=4.25746e-07 $layer=POLY_cond $X=3.335 $Y=1.765
+ $X2=3.432 $Y2=1.385
r24 4 6 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=3.335 $Y=1.765
+ $X2=3.335 $Y2=2.34
r25 1 10 38.561 $w=2.98e-07 $l=2.13787e-07 $layer=POLY_cond $X=3.32 $Y=1.22
+ $X2=3.432 $Y2=1.385
r26 1 3 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=3.32 $Y=1.22 $X2=3.32
+ $Y2=0.79
.ends

.subckt PM_SKY130_FD_SC_HS__A32O_1%X 1 2 11 14 15 16 17 28
r24 21 28 0.800308 $w=3.58e-07 $l=2.5e-08 $layer=LI1_cond $X=0.265 $Y=0.95
+ $X2=0.265 $Y2=0.925
r25 17 30 8.03084 $w=3.58e-07 $l=1.5e-07 $layer=LI1_cond $X=0.265 $Y=0.98
+ $X2=0.265 $Y2=1.13
r26 17 21 0.960369 $w=3.58e-07 $l=3e-08 $layer=LI1_cond $X=0.265 $Y=0.98
+ $X2=0.265 $Y2=0.95
r27 17 28 0.960369 $w=3.58e-07 $l=3e-08 $layer=LI1_cond $X=0.265 $Y=0.895
+ $X2=0.265 $Y2=0.925
r28 16 17 12.1647 $w=3.58e-07 $l=3.8e-07 $layer=LI1_cond $X=0.265 $Y=0.515
+ $X2=0.265 $Y2=0.895
r29 15 30 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=0.17 $Y=1.82 $X2=0.17
+ $Y2=1.13
r30 14 15 8.53881 $w=3.68e-07 $l=1.65e-07 $layer=LI1_cond $X=0.27 $Y=1.985
+ $X2=0.27 $Y2=1.82
r31 9 14 0.622942 $w=3.68e-07 $l=2e-08 $layer=LI1_cond $X=0.27 $Y=2.005 $X2=0.27
+ $Y2=1.985
r32 9 11 25.2292 $w=3.68e-07 $l=8.1e-07 $layer=LI1_cond $X=0.27 $Y=2.005
+ $X2=0.27 $Y2=2.815
r33 2 14 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.145
+ $Y=1.84 $X2=0.29 $Y2=1.985
r34 2 11 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=0.145
+ $Y=1.84 $X2=0.29 $Y2=2.815
r35 1 16 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__A32O_1%VPWR 1 2 9 15 18 19 20 22 35 36 39
r43 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r44 35 36 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r45 33 36 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=3.6 $Y2=3.33
r46 32 35 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=2.16 $Y=3.33
+ $X2=3.6 $Y2=3.33
r47 32 33 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r48 30 40 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=0.72 $Y2=3.33
r49 29 30 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r50 27 39 9.6488 $w=1.7e-07 $l=1.95e-07 $layer=LI1_cond $X=1.015 $Y=3.33
+ $X2=0.82 $Y2=3.33
r51 27 29 43.385 $w=1.68e-07 $l=6.65e-07 $layer=LI1_cond $X=1.015 $Y=3.33
+ $X2=1.68 $Y2=3.33
r52 25 40 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r53 24 25 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r54 22 39 9.6488 $w=1.7e-07 $l=1.95e-07 $layer=LI1_cond $X=0.625 $Y=3.33
+ $X2=0.82 $Y2=3.33
r55 22 24 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=0.625 $Y=3.33
+ $X2=0.24 $Y2=3.33
r56 20 33 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=2.16 $Y2=3.33
r57 20 30 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=1.68 $Y2=3.33
r58 18 29 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=1.8 $Y=3.33 $X2=1.68
+ $Y2=3.33
r59 18 19 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.8 $Y=3.33
+ $X2=1.965 $Y2=3.33
r60 17 32 1.95722 $w=1.68e-07 $l=3e-08 $layer=LI1_cond $X=2.13 $Y=3.33 $X2=2.16
+ $Y2=3.33
r61 17 19 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.13 $Y=3.33
+ $X2=1.965 $Y2=3.33
r62 13 19 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.965 $Y=3.245
+ $X2=1.965 $Y2=3.33
r63 13 15 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=1.965 $Y=3.245
+ $X2=1.965 $Y2=2.565
r64 9 12 17.4344 $w=3.88e-07 $l=5.9e-07 $layer=LI1_cond $X=0.82 $Y=2.225
+ $X2=0.82 $Y2=2.815
r65 7 39 1.39532 $w=3.9e-07 $l=8.5e-08 $layer=LI1_cond $X=0.82 $Y=3.245 $X2=0.82
+ $Y2=3.33
r66 7 12 12.7064 $w=3.88e-07 $l=4.3e-07 $layer=LI1_cond $X=0.82 $Y=3.245
+ $X2=0.82 $Y2=2.815
r67 2 15 600 $w=1.7e-07 $l=8.59942e-07 $layer=licon1_PDIFF $count=1 $X=1.67
+ $Y=1.84 $X2=1.965 $Y2=2.565
r68 1 12 600 $w=1.7e-07 $l=1.07034e-06 $layer=licon1_PDIFF $count=1 $X=0.59
+ $Y=1.84 $X2=0.79 $Y2=2.815
r69 1 9 600 $w=1.7e-07 $l=4.98322e-07 $layer=licon1_PDIFF $count=1 $X=0.59
+ $Y=1.84 $X2=0.85 $Y2=2.225
.ends

.subckt PM_SKY130_FD_SC_HS__A32O_1%A_244_368# 1 2 3 12 14 15 16 17 20 25
r39 20 23 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=3.56 $Y=1.985
+ $X2=3.56 $Y2=2.695
r40 18 23 7.33373 $w=3.28e-07 $l=2.1e-07 $layer=LI1_cond $X=3.56 $Y=2.905
+ $X2=3.56 $Y2=2.695
r41 16 18 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.395 $Y=2.99
+ $X2=3.56 $Y2=2.905
r42 16 17 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.395 $Y=2.99
+ $X2=2.725 $Y2=2.99
r43 15 17 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.56 $Y=2.905
+ $X2=2.725 $Y2=2.99
r44 14 27 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.56 $Y=2.23 $X2=2.56
+ $Y2=2.145
r45 14 15 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=2.56 $Y=2.23
+ $X2=2.56 $Y2=2.905
r46 13 25 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.535 $Y=2.145
+ $X2=1.37 $Y2=2.145
r47 12 27 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.395 $Y=2.145
+ $X2=2.56 $Y2=2.145
r48 12 13 56.107 $w=1.68e-07 $l=8.6e-07 $layer=LI1_cond $X=2.395 $Y=2.145
+ $X2=1.535 $Y2=2.145
r49 3 23 400 $w=1.7e-07 $l=9.26971e-07 $layer=licon1_PDIFF $count=1 $X=3.41
+ $Y=1.84 $X2=3.56 $Y2=2.695
r50 3 20 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=3.41
+ $Y=1.84 $X2=3.56 $Y2=1.985
r51 2 27 300 $w=1.7e-07 $l=4.08167e-07 $layer=licon1_PDIFF $count=2 $X=2.41
+ $Y=1.84 $X2=2.56 $Y2=2.18
r52 1 25 300 $w=1.7e-07 $l=4.08167e-07 $layer=licon1_PDIFF $count=2 $X=1.22
+ $Y=1.84 $X2=1.37 $Y2=2.18
.ends

.subckt PM_SKY130_FD_SC_HS__A32O_1%VGND 1 2 11 13 15 17 19 28 32
r38 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r39 28 29 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r40 26 32 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=3.6
+ $Y2=0
r41 25 26 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r42 23 29 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r43 22 25 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=1.2 $Y=0 $X2=3.12
+ $Y2=0
r44 22 23 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r45 20 28 9.81116 $w=1.7e-07 $l=2e-07 $layer=LI1_cond $X=1.05 $Y=0 $X2=0.85
+ $Y2=0
r46 20 22 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=1.05 $Y=0 $X2=1.2
+ $Y2=0
r47 19 31 4.67962 $w=1.7e-07 $l=2.35e-07 $layer=LI1_cond $X=3.37 $Y=0 $X2=3.605
+ $Y2=0
r48 19 25 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=3.37 $Y=0 $X2=3.12
+ $Y2=0
r49 17 26 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=1.92 $Y=0 $X2=3.12
+ $Y2=0
r50 17 23 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=1.2
+ $Y2=0
r51 13 31 3.08656 $w=3.3e-07 $l=1.14782e-07 $layer=LI1_cond $X=3.535 $Y=0.085
+ $X2=3.605 $Y2=0
r52 13 15 18.5089 $w=3.28e-07 $l=5.3e-07 $layer=LI1_cond $X=3.535 $Y=0.085
+ $X2=3.535 $Y2=0.615
r53 9 28 1.46811 $w=4e-07 $l=8.5e-08 $layer=LI1_cond $X=0.85 $Y=0.085 $X2=0.85
+ $Y2=0
r54 9 11 13.2531 $w=3.98e-07 $l=4.6e-07 $layer=LI1_cond $X=0.85 $Y=0.085
+ $X2=0.85 $Y2=0.545
r55 2 15 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.395
+ $Y=0.47 $X2=3.535 $Y2=0.615
r56 1 11 182 $w=1.7e-07 $l=3.56931e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.37 $X2=0.85 $Y2=0.545
.ends

