* NGSPICE file created from sky130_fd_sc_hs__a2bb2o_4.ext - technology: sky130A

.subckt sky130_fd_sc_hs__a2bb2o_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
M1000 VPWR a_162_48# X VPB pshort w=1.12e+06u l=150000u
+  ad=1.6808e+12p pd=1.385e+07u as=6.72e+11p ps=5.68e+06u
M1001 a_586_94# A2_N a_583_368# VPB pshort w=1.12e+06u l=150000u
+  ad=3.08e+11p pd=2.79e+06u as=2.688e+11p ps=2.72e+06u
M1002 VGND a_162_48# X VNB nlowvt w=740000u l=150000u
+  ad=1.6403e+12p pd=1.199e+07u as=4.144e+11p ps=4.08e+06u
M1003 a_1009_74# B2 a_162_48# VNB nlowvt w=640000u l=150000u
+  ad=5.184e+11p pd=5.46e+06u as=3.753e+11p ps=3.85e+06u
M1004 a_583_368# A1_N VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_162_48# a_586_94# a_820_392# VPB pshort w=1e+06u l=150000u
+  ad=3e+11p pd=2.6e+06u as=1.15e+12p ps=1.03e+07u
M1006 a_1009_74# B1 VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 X a_162_48# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VGND B1 a_1009_74# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_820_392# a_586_94# a_162_48# VPB pshort w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 X a_162_48# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_162_48# B2 a_1009_74# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_586_94# A1_N VGND VNB nlowvt w=640000u l=150000u
+  ad=1.792e+11p pd=1.84e+06u as=0p ps=0u
M1013 a_162_48# a_586_94# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 VPWR B2 a_820_392# VPB pshort w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 X a_162_48# VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_820_392# B2 VPWR VPB pshort w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 VGND a_162_48# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 VPWR a_162_48# X VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VPWR B1 a_820_392# VPB pshort w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 VGND A2_N a_586_94# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 X a_162_48# VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_820_392# B1 VPWR VPB pshort w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

