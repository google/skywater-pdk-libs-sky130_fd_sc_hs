# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_hs__bufbuf_8
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_hs__bufbuf_8 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  7.200000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.208500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.350000 0.570000 1.780000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  2.273200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.475000 0.350000 3.805000 0.880000 ;
        RECT 3.475000 0.880000 6.585000 1.130000 ;
        RECT 3.565000 1.800000 6.555000 1.970000 ;
        RECT 3.565000 1.970000 3.830000 2.980000 ;
        RECT 4.495000 1.970000 4.745000 2.980000 ;
        RECT 5.385000 1.970000 5.655000 2.980000 ;
        RECT 6.255000 0.350000 6.585000 0.880000 ;
        RECT 6.255000 1.130000 6.585000 1.270000 ;
        RECT 6.255000 1.270000 7.075000 1.780000 ;
        RECT 6.255000 1.780000 6.555000 1.800000 ;
        RECT 6.285000 1.970000 6.555000 2.980000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 7.200000 0.085000 ;
        RECT 0.625000  0.085000 0.955000 0.840000 ;
        RECT 2.115000  0.085000 2.445000 0.710000 ;
        RECT 2.975000  0.085000 3.305000 0.710000 ;
        RECT 3.975000  0.085000 4.305000 0.710000 ;
        RECT 4.835000  0.085000 5.165000 0.710000 ;
        RECT 5.755000  0.085000 6.085000 0.710000 ;
        RECT 6.755000  0.085000 7.085000 1.100000 ;
      LAYER mcon ;
        RECT 0.155000 -0.085000 0.325000 0.085000 ;
        RECT 0.635000 -0.085000 0.805000 0.085000 ;
        RECT 1.115000 -0.085000 1.285000 0.085000 ;
        RECT 1.595000 -0.085000 1.765000 0.085000 ;
        RECT 2.075000 -0.085000 2.245000 0.085000 ;
        RECT 2.555000 -0.085000 2.725000 0.085000 ;
        RECT 3.035000 -0.085000 3.205000 0.085000 ;
        RECT 3.515000 -0.085000 3.685000 0.085000 ;
        RECT 3.995000 -0.085000 4.165000 0.085000 ;
        RECT 4.475000 -0.085000 4.645000 0.085000 ;
        RECT 4.955000 -0.085000 5.125000 0.085000 ;
        RECT 5.435000 -0.085000 5.605000 0.085000 ;
        RECT 5.915000 -0.085000 6.085000 0.085000 ;
        RECT 6.395000 -0.085000 6.565000 0.085000 ;
        RECT 6.875000 -0.085000 7.045000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.245000 7.200000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 3.245000 7.200000 3.415000 ;
        RECT 0.565000 2.370000 0.920000 3.245000 ;
        RECT 2.150000 2.160000 2.380000 3.245000 ;
        RECT 3.050000 1.820000 3.380000 3.245000 ;
        RECT 4.035000 2.140000 4.290000 3.245000 ;
        RECT 4.930000 2.140000 5.205000 3.245000 ;
        RECT 5.835000 2.140000 6.105000 3.245000 ;
        RECT 6.735000 1.950000 7.040000 3.245000 ;
      LAYER mcon ;
        RECT 0.155000 3.245000 0.325000 3.415000 ;
        RECT 0.635000 3.245000 0.805000 3.415000 ;
        RECT 1.115000 3.245000 1.285000 3.415000 ;
        RECT 1.595000 3.245000 1.765000 3.415000 ;
        RECT 2.075000 3.245000 2.245000 3.415000 ;
        RECT 2.555000 3.245000 2.725000 3.415000 ;
        RECT 3.035000 3.245000 3.205000 3.415000 ;
        RECT 3.515000 3.245000 3.685000 3.415000 ;
        RECT 3.995000 3.245000 4.165000 3.415000 ;
        RECT 4.475000 3.245000 4.645000 3.415000 ;
        RECT 4.955000 3.245000 5.125000 3.415000 ;
        RECT 5.435000 3.245000 5.605000 3.415000 ;
        RECT 5.915000 3.245000 6.085000 3.415000 ;
        RECT 6.395000 3.245000 6.565000 3.415000 ;
        RECT 6.875000 3.245000 7.045000 3.415000 ;
      LAYER met1 ;
        RECT 0.000000 3.085000 7.200000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.115000 0.540000 0.445000 1.010000 ;
      RECT 0.115000 1.010000 0.920000 1.180000 ;
      RECT 0.115000 1.950000 0.920000 2.200000 ;
      RECT 0.115000 2.200000 0.380000 2.700000 ;
      RECT 0.750000 1.180000 0.920000 1.300000 ;
      RECT 0.750000 1.300000 1.140000 1.630000 ;
      RECT 0.750000 1.630000 0.920000 1.950000 ;
      RECT 1.090000 1.820000 1.480000 2.980000 ;
      RECT 1.125000 0.350000 1.480000 1.130000 ;
      RECT 1.310000 1.130000 1.480000 1.300000 ;
      RECT 1.310000 1.300000 2.500000 1.630000 ;
      RECT 1.310000 1.630000 1.480000 1.820000 ;
      RECT 1.650000 1.820000 2.880000 1.990000 ;
      RECT 1.650000 1.990000 1.980000 2.980000 ;
      RECT 1.685000 0.350000 1.935000 0.880000 ;
      RECT 1.685000 0.880000 3.125000 1.130000 ;
      RECT 2.550000 1.990000 2.880000 2.980000 ;
      RECT 2.670000 1.130000 3.125000 1.300000 ;
      RECT 2.670000 1.300000 6.020000 1.630000 ;
      RECT 2.670000 1.630000 2.880000 1.820000 ;
  END
END sky130_fd_sc_hs__bufbuf_8
