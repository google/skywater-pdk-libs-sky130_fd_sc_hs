* File: sky130_fd_sc_hs__o21bai_1.spice
* Created: Tue Sep  1 20:15:08 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hs__o21bai_1.pex.spice"
.subckt sky130_fd_sc_hs__o21bai_1  VNB VPB B1_N A2 A1 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A1	A1
* A2	A2
* B1_N	B1_N
* VPB	VPB
* VNB	VNB
MM1001 N_VGND_M1001_d N_B1_N_M1001_g N_A_27_74#_M1001_s VNB NLOWVT L=0.15 W=0.55
+ AD=0.15125 AS=0.154 PD=1.65 PS=1.66 NRD=0 NRS=0 M=1 R=3.66667 SA=75000.2
+ SB=75000.2 A=0.0825 P=1.4 MULT=1
MM1003 N_A_308_74#_M1003_d N_A_27_74#_M1003_g N_Y_M1003_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1221 AS=0.2072 PD=1.07 PS=2.04 NRD=8.1 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75001.1 A=0.111 P=1.78 MULT=1
MM1004 N_VGND_M1004_d N_A2_M1004_g N_A_308_74#_M1003_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.1073 AS=0.1221 PD=1.03 PS=1.07 NRD=0.804 NRS=0 M=1 R=4.93333 SA=75000.7
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1002 N_A_308_74#_M1002_d N_A1_M1002_g N_VGND_M1004_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.1073 PD=2.05 PS=1.03 NRD=0 NRS=0.804 M=1 R=4.93333 SA=75001.1
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1000 N_VPWR_M1000_d N_B1_N_M1000_g N_A_27_74#_M1000_s VPB PSHORT L=0.15 W=0.84
+ AD=0.3108 AS=0.2478 PD=1.62429 PS=2.27 NRD=14.0658 NRS=2.3443 M=1 R=5.6
+ SA=75000.2 SB=75002.1 A=0.126 P=1.98 MULT=1
MM1005 N_Y_M1005_d N_A_27_74#_M1005_g N_VPWR_M1000_d VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.4144 PD=1.42 PS=2.16571 NRD=1.7533 NRS=16.7056 M=1 R=7.46667
+ SA=75000.9 SB=75001.1 A=0.168 P=2.54 MULT=1
MM1007 A_395_368# N_A2_M1007_g N_Y_M1005_d VPB PSHORT L=0.15 W=1.12 AD=0.1848
+ AS=0.168 PD=1.45 PS=1.42 NRD=19.3454 NRS=1.7533 M=1 R=7.46667 SA=75001.4
+ SB=75000.7 A=0.168 P=2.54 MULT=1
MM1006 N_VPWR_M1006_d N_A1_M1006_g A_395_368# VPB PSHORT L=0.15 W=1.12 AD=0.3248
+ AS=0.1848 PD=2.82 PS=1.45 NRD=1.7533 NRS=19.3454 M=1 R=7.46667 SA=75001.8
+ SB=75000.2 A=0.168 P=2.54 MULT=1
DX8_noxref VNB VPB NWDIODE A=6.0636 P=10.24
*
.include "sky130_fd_sc_hs__o21bai_1.pxi.spice"
*
.ends
*
*
