* File: sky130_fd_sc_hs__a2111o_1.spice
* Created: Tue Sep  1 19:47:49 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hs__a2111o_1.pex.spice"
.subckt sky130_fd_sc_hs__a2111o_1  VNB VPB A1 A2 B1 C1 D1 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* D1	D1
* C1	C1
* B1	B1
* A2	A2
* A1	A1
* VPB	VPB
* VNB	VNB
MM1001 A_168_136# N_A1_M1001_g N_A_85_136#_M1001_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.0672 AS=0.1696 PD=0.85 PS=1.81 NRD=9.372 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75002.1 A=0.096 P=1.58 MULT=1
MM1003 N_VGND_M1003_d N_A2_M1003_g A_168_136# VNB NLOWVT L=0.15 W=0.64 AD=0.1248
+ AS=0.0672 PD=1.03 PS=0.85 NRD=0 NRS=9.372 M=1 R=4.26667 SA=75000.6 SB=75001.8
+ A=0.096 P=1.58 MULT=1
MM1004 N_A_85_136#_M1004_d N_B1_M1004_g N_VGND_M1003_d VNB NLOWVT L=0.15 W=0.64
+ AD=0.0896 AS=0.1248 PD=0.92 PS=1.03 NRD=0 NRS=20.616 M=1 R=4.26667 SA=75001.1
+ SB=75001.2 A=0.096 P=1.58 MULT=1
MM1005 N_VGND_M1005_d N_C1_M1005_g N_A_85_136#_M1004_d VNB NLOWVT L=0.15 W=0.64
+ AD=0.1504 AS=0.0896 PD=1.11 PS=0.92 NRD=35.616 NRS=0 M=1 R=4.26667 SA=75001.5
+ SB=75000.8 A=0.096 P=1.58 MULT=1
MM1002 N_A_85_136#_M1002_d N_D1_M1002_g N_VGND_M1005_d VNB NLOWVT L=0.15 W=0.64
+ AD=0.1696 AS=0.1504 PD=1.81 PS=1.11 NRD=0 NRS=0 M=1 R=4.26667 SA=75002.1
+ SB=75000.2 A=0.096 P=1.58 MULT=1
MM1008 N_X_M1008_d N_A_85_136#_M1008_g N_VGND_M1008_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1961 AS=0.1961 PD=2.01 PS=2.01 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1010 N_VPWR_M1010_d N_A1_M1010_g N_A_80_392#_M1010_s VPB PSHORT L=0.15 W=1
+ AD=0.17 AS=0.275 PD=1.34 PS=2.55 NRD=5.8903 NRS=1.9503 M=1 R=6.66667
+ SA=75000.2 SB=75001.9 A=0.15 P=2.3 MULT=1
MM1006 N_A_80_392#_M1006_d N_A2_M1006_g N_VPWR_M1010_d VPB PSHORT L=0.15 W=1
+ AD=0.15 AS=0.17 PD=1.3 PS=1.34 NRD=1.9503 NRS=5.8903 M=1 R=6.66667 SA=75000.7
+ SB=75001.4 A=0.15 P=2.3 MULT=1
MM1007 A_353_392# N_B1_M1007_g N_A_80_392#_M1006_d VPB PSHORT L=0.15 W=1 AD=0.12
+ AS=0.15 PD=1.24 PS=1.3 NRD=12.7853 NRS=1.9503 M=1 R=6.66667 SA=75001.1
+ SB=75001 A=0.15 P=2.3 MULT=1
MM1000 A_431_392# N_C1_M1000_g A_353_392# VPB PSHORT L=0.15 W=1 AD=0.12 AS=0.12
+ PD=1.24 PS=1.24 NRD=12.7853 NRS=12.7853 M=1 R=6.66667 SA=75001.5 SB=75000.6
+ A=0.15 P=2.3 MULT=1
MM1009 N_A_85_136#_M1009_d N_D1_M1009_g A_431_392# VPB PSHORT L=0.15 W=1
+ AD=0.275 AS=0.12 PD=2.55 PS=1.24 NRD=1.9503 NRS=12.7853 M=1 R=6.66667
+ SA=75001.9 SB=75000.2 A=0.15 P=2.3 MULT=1
MM1011 N_X_M1011_d N_A_85_136#_M1011_g N_VPWR_M1011_s VPB PSHORT L=0.15 W=1.12
+ AD=0.308 AS=0.308 PD=2.79 PS=2.79 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75000.2 A=0.168 P=2.54 MULT=1
DX12_noxref VNB VPB NWDIODE A=8.742 P=13.12
*
.include "sky130_fd_sc_hs__a2111o_1.pxi.spice"
*
.ends
*
*
