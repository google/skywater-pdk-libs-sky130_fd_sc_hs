# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_sc_hs__a31oi_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__a31oi_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  8.640000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  1.116000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.925000 1.350000 6.115000 1.780000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  1.116000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.415000 1.350000 4.195000 1.780000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  1.116000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.350000 1.745000 1.780000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.894000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.365000 1.350000 8.515000 1.780000 ;
    END
  END B1
  PIN Y
    ANTENNADIFFAREA  1.621350 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.350000 0.770000 4.685000 0.965000 ;
        RECT 4.350000 0.965000 5.840000 1.010000 ;
        RECT 4.350000 1.010000 8.525000 1.130000 ;
        RECT 4.445000 1.130000 8.525000 1.180000 ;
        RECT 4.445000 1.180000 4.690000 1.950000 ;
        RECT 4.445000 1.950000 8.075000 2.120000 ;
        RECT 5.510000 0.595000 5.840000 0.965000 ;
        RECT 6.510000 0.350000 6.840000 1.010000 ;
        RECT 6.845000 2.120000 7.175000 2.735000 ;
        RECT 7.745000 2.120000 8.075000 2.735000 ;
        RECT 8.195000 0.350000 8.525000 1.010000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 8.640000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.000000 0.000000 8.640000 0.245000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.660000 8.830000 3.520000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 8.640000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 8.640000 0.085000 ;
      RECT 0.000000  3.245000 8.640000 3.415000 ;
      RECT 0.115000  1.950000 4.195000 2.120000 ;
      RECT 0.115000  2.120000 0.395000 2.980000 ;
      RECT 0.130000  0.350000 0.380000 1.010000 ;
      RECT 0.130000  1.010000 4.120000 1.180000 ;
      RECT 0.560000  0.085000 0.890000 0.840000 ;
      RECT 0.565000  2.290000 0.895000 3.245000 ;
      RECT 1.065000  2.120000 1.295000 2.935000 ;
      RECT 1.070000  0.350000 1.240000 1.010000 ;
      RECT 1.420000  0.085000 1.750000 0.840000 ;
      RECT 1.465000  2.290000 1.795000 3.245000 ;
      RECT 1.915000  1.820000 2.245000 1.950000 ;
      RECT 1.920000  0.330000 2.170000 1.010000 ;
      RECT 1.965000  2.120000 3.195000 2.150000 ;
      RECT 1.965000  2.150000 2.195000 2.950000 ;
      RECT 2.350000  0.255000 6.340000 0.425000 ;
      RECT 2.350000  0.425000 2.655000 0.840000 ;
      RECT 2.365000  2.320000 2.695000 3.245000 ;
      RECT 2.825000  0.595000 3.120000 1.010000 ;
      RECT 2.865000  2.150000 3.195000 2.980000 ;
      RECT 3.290000  0.425000 3.620000 0.840000 ;
      RECT 3.365000  2.290000 3.695000 3.245000 ;
      RECT 3.790000  0.595000 4.120000 1.010000 ;
      RECT 3.865000  2.120000 4.195000 2.290000 ;
      RECT 3.865000  2.290000 6.675000 2.460000 ;
      RECT 3.865000  2.460000 4.195000 2.980000 ;
      RECT 4.365000  2.630000 4.695000 3.245000 ;
      RECT 4.865000  2.460000 5.675000 2.930000 ;
      RECT 4.935000  0.425000 5.265000 0.795000 ;
      RECT 5.845000  2.630000 6.175000 3.245000 ;
      RECT 6.010000  0.425000 6.340000 0.840000 ;
      RECT 6.345000  2.460000 6.675000 2.905000 ;
      RECT 6.345000  2.905000 8.525000 3.075000 ;
      RECT 7.010000  0.085000 8.025000 0.840000 ;
      RECT 7.375000  2.290000 7.575000 2.905000 ;
      RECT 8.255000  1.950000 8.525000 2.905000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
      RECT 7.835000 -0.085000 8.005000 0.085000 ;
      RECT 7.835000  3.245000 8.005000 3.415000 ;
      RECT 8.315000 -0.085000 8.485000 0.085000 ;
      RECT 8.315000  3.245000 8.485000 3.415000 ;
  END
END sky130_fd_sc_hs__a31oi_4
END LIBRARY
