* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hs__dlymetal6s6s_1 A VGND VNB VPB VPWR X
M1000 VGND a_497_74# a_604_138# VNB nlowvt w=420000u l=150000u
+  ad=6.828e+11p pd=6.48e+06u as=1.113e+11p ps=1.37e+06u
M1001 a_497_74# a_316_138# VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=3.08e+11p pd=2.79e+06u as=1.043e+12p ps=8.92e+06u
M1002 a_209_74# a_28_138# VGND VNB nlowvt w=740000u l=150000u
+  ad=1.961e+11p pd=2.01e+06u as=0p ps=0u
M1003 VPWR a_497_74# a_604_138# VPB pshort w=420000u l=150000u
+  ad=0p pd=0u as=1.155e+11p ps=1.39e+06u
M1004 VPWR A a_28_138# VPB pshort w=420000u l=150000u
+  ad=0p pd=0u as=1.155e+11p ps=1.39e+06u
M1005 X a_604_138# VGND VNB nlowvt w=740000u l=150000u
+  ad=1.961e+11p pd=2.01e+06u as=0p ps=0u
M1006 VGND A a_28_138# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1007 a_209_74# a_28_138# VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=3.08e+11p pd=2.79e+06u as=0p ps=0u
M1008 VGND a_209_74# a_316_138# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1009 X a_604_138# VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=3.08e+11p pd=2.79e+06u as=0p ps=0u
M1010 a_497_74# a_316_138# VGND VNB nlowvt w=740000u l=150000u
+  ad=1.961e+11p pd=2.01e+06u as=0p ps=0u
M1011 VPWR a_209_74# a_316_138# VPB pshort w=420000u l=150000u
+  ad=0p pd=0u as=1.155e+11p ps=1.39e+06u
.ends
