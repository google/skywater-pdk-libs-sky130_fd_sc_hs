* File: sky130_fd_sc_hs__sdfxtp_4.spice
* Created: Thu Aug 27 21:10:23 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hs__sdfxtp_4.pex.spice"
.subckt sky130_fd_sc_hs__sdfxtp_4  VNB VPB SCE D SCD CLK VPWR Q VGND
* 
* VGND	VGND
* Q	Q
* VPWR	VPWR
* CLK	CLK
* SCD	SCD
* D	D
* SCE	SCE
* VPB	VPB
* VNB	VNB
MM1037 N_VGND_M1037_d N_SCE_M1037_g N_A_36_74#_M1037_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.0735 AS=0.1197 PD=0.77 PS=1.41 NRD=19.992 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75002.7 A=0.063 P=1.14 MULT=1
MM1023 A_223_74# N_A_36_74#_M1023_g N_VGND_M1037_d VNB NLOWVT L=0.15 W=0.42
+ AD=0.0504 AS=0.0735 PD=0.66 PS=0.77 NRD=18.564 NRS=0 M=1 R=2.8 SA=75000.7
+ SB=75002.2 A=0.063 P=1.14 MULT=1
MM1024 N_A_301_74#_M1024_d N_D_M1024_g A_223_74# VNB NLOWVT L=0.15 W=0.42
+ AD=0.12705 AS=0.0504 PD=1.025 PS=0.66 NRD=45.708 NRS=18.564 M=1 R=2.8
+ SA=75001.1 SB=75001.9 A=0.063 P=1.14 MULT=1
MM1008 A_452_74# N_SCE_M1008_g N_A_301_74#_M1024_d VNB NLOWVT L=0.15 W=0.42
+ AD=0.0504 AS=0.12705 PD=0.66 PS=1.025 NRD=18.564 NRS=47.136 M=1 R=2.8
+ SA=75001.9 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1005 N_VGND_M1005_d N_SCD_M1005_g A_452_74# VNB NLOWVT L=0.15 W=0.42
+ AD=0.0821897 AS=0.0504 PD=0.78931 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8
+ SA=75002.2 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1002 N_A_630_74#_M1002_d N_CLK_M1002_g N_VGND_M1005_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.14481 PD=2.05 PS=1.39069 NRD=0 NRS=11.34 M=1 R=4.93333
+ SA=75001.6 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1020 N_A_828_74#_M1020_d N_A_630_74#_M1020_g N_VGND_M1020_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.2109 AS=0.2109 PD=2.05 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1027 N_A_1026_100#_M1027_d N_A_630_74#_M1027_g N_A_301_74#_M1027_s VNB NLOWVT
+ L=0.15 W=0.42 AD=0.1113 AS=0.1197 PD=0.95 PS=1.41 NRD=71.424 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75004 A=0.063 P=1.14 MULT=1
MM1012 A_1162_100# N_A_828_74#_M1012_g N_A_1026_100#_M1027_d VNB NLOWVT L=0.15
+ W=0.42 AD=0.09975 AS=0.1113 PD=0.895 PS=0.95 NRD=52.14 NRS=0 M=1 R=2.8
+ SA=75000.9 SB=75003.3 A=0.063 P=1.14 MULT=1
MM1035 N_VGND_M1035_d N_A_1257_74#_M1035_g A_1162_100# VNB NLOWVT L=0.15 W=0.42
+ AD=0.179149 AS=0.09975 PD=1.14309 PS=0.895 NRD=24.276 NRS=52.14 M=1 R=2.8
+ SA=75001.5 SB=75002.7 A=0.063 P=1.14 MULT=1
MM1036 N_A_1257_74#_M1036_d N_A_1026_100#_M1036_g N_VGND_M1035_d VNB NLOWVT
+ L=0.15 W=0.55 AD=0.11825 AS=0.234601 PD=0.98 PS=1.49691 NRD=13.08 NRS=89.448
+ M=1 R=3.66667 SA=75002 SB=75001.9 A=0.0825 P=1.4 MULT=1
MM1032 N_A_1587_74#_M1032_d N_A_828_74#_M1032_g N_A_1257_74#_M1036_d VNB NLOWVT
+ L=0.15 W=0.55 AD=0.226804 AS=0.11825 PD=1.46856 PS=0.98 NRD=84 NRS=19.632 M=1
+ R=3.66667 SA=75002.6 SB=75001.3 A=0.0825 P=1.4 MULT=1
MM1018 A_1766_74# N_A_630_74#_M1018_g N_A_1587_74#_M1032_d VNB NLOWVT L=0.15
+ W=0.42 AD=0.0504 AS=0.173196 PD=0.66 PS=1.12144 NRD=18.564 NRS=22.848 M=1
+ R=2.8 SA=75003.3 SB=75000.6 A=0.063 P=1.14 MULT=1
MM1016 N_VGND_M1016_d N_A_1814_48#_M1016_g A_1766_74# VNB NLOWVT L=0.15 W=0.42
+ AD=0.1197 AS=0.0504 PD=1.41 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75003.7
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1029 N_VGND_M1029_d N_A_1587_74#_M1029_g N_A_1814_48#_M1029_s VNB NLOWVT
+ L=0.15 W=0.74 AD=0.12025 AS=0.2109 PD=1.065 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75002.1 A=0.111 P=1.78 MULT=1
MM1004 N_VGND_M1029_d N_A_1814_48#_M1004_g N_Q_M1004_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.12025 AS=0.13505 PD=1.065 PS=1.105 NRD=7.296 NRS=13.776 M=1 R=4.93333
+ SA=75000.7 SB=75001.6 A=0.111 P=1.78 MULT=1
MM1015 N_VGND_M1015_d N_A_1814_48#_M1015_g N_Q_M1004_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.13505 PD=1.02 PS=1.105 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.2
+ SB=75001.1 A=0.111 P=1.78 MULT=1
MM1017 N_VGND_M1015_d N_A_1814_48#_M1017_g N_Q_M1017_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.6
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1030 N_VGND_M1030_d N_A_1814_48#_M1030_g N_Q_M1017_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.1036 PD=2.05 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75002.1
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1025 N_VPWR_M1025_d N_SCE_M1025_g N_A_36_74#_M1025_s VPB PSHORT L=0.15 W=0.64
+ AD=0.112 AS=0.1888 PD=0.99 PS=1.87 NRD=18.4589 NRS=3.0732 M=1 R=4.26667
+ SA=75000.2 SB=75002.9 A=0.096 P=1.58 MULT=1
MM1026 A_238_464# N_SCE_M1026_g N_VPWR_M1025_d VPB PSHORT L=0.15 W=0.64
+ AD=0.0864 AS=0.112 PD=0.91 PS=0.99 NRD=24.625 NRS=3.0732 M=1 R=4.26667
+ SA=75000.7 SB=75002.4 A=0.096 P=1.58 MULT=1
MM1006 N_A_301_74#_M1006_d N_D_M1006_g A_238_464# VPB PSHORT L=0.15 W=0.64
+ AD=0.096 AS=0.0864 PD=0.94 PS=0.91 NRD=3.0732 NRS=24.625 M=1 R=4.26667
+ SA=75001.1 SB=75001.9 A=0.096 P=1.58 MULT=1
MM1011 A_412_464# N_A_36_74#_M1011_g N_A_301_74#_M1006_d VPB PSHORT L=0.15
+ W=0.64 AD=0.1248 AS=0.096 PD=1.03 PS=0.94 NRD=43.0839 NRS=3.0732 M=1 R=4.26667
+ SA=75001.6 SB=75001.5 A=0.096 P=1.58 MULT=1
MM1028 N_VPWR_M1028_d N_SCD_M1028_g A_412_464# VPB PSHORT L=0.15 W=0.64
+ AD=0.183564 AS=0.1248 PD=1.24364 PS=1.03 NRD=47.6937 NRS=43.0839 M=1 R=4.26667
+ SA=75002.1 SB=75001 A=0.096 P=1.58 MULT=1
MM1013 N_A_630_74#_M1013_d N_CLK_M1013_g N_VPWR_M1028_d VPB PSHORT L=0.15 W=1.12
+ AD=0.3304 AS=0.321236 PD=2.83 PS=2.17636 NRD=1.7533 NRS=27.2451 M=1 R=7.46667
+ SA=75001.7 SB=75000.2 A=0.168 P=2.54 MULT=1
MM1007 N_A_828_74#_M1007_d N_A_630_74#_M1007_g N_VPWR_M1007_s VPB PSHORT L=0.15
+ W=1.12 AD=0.3304 AS=0.6216 PD=2.83 PS=3.35 NRD=1.7533 NRS=24.625 M=1 R=7.46667
+ SA=75000.5 SB=75000.2 A=0.168 P=2.54 MULT=1
MM1014 N_A_1026_100#_M1014_d N_A_828_74#_M1014_g N_A_301_74#_M1014_s VPB PSHORT
+ L=0.15 W=0.42 AD=0.063 AS=0.1239 PD=0.72 PS=1.43 NRD=4.6886 NRS=4.6886 M=1
+ R=2.8 SA=75000.2 SB=75005.3 A=0.063 P=1.14 MULT=1
MM1019 A_1214_506# N_A_630_74#_M1019_g N_A_1026_100#_M1014_d VPB PSHORT L=0.15
+ W=0.42 AD=0.0819 AS=0.063 PD=0.81 PS=0.72 NRD=65.6601 NRS=4.6886 M=1 R=2.8
+ SA=75000.7 SB=75004.9 A=0.063 P=1.14 MULT=1
MM1033 N_VPWR_M1033_d N_A_1257_74#_M1033_g A_1214_506# VPB PSHORT L=0.15 W=0.42
+ AD=0.123392 AS=0.0819 PD=1.01333 PS=0.81 NRD=46.886 NRS=65.6601 M=1 R=2.8
+ SA=75001.2 SB=75004.3 A=0.063 P=1.14 MULT=1
MM1009 N_A_1257_74#_M1009_d N_A_1026_100#_M1009_g N_VPWR_M1033_d VPB PSHORT
+ L=0.15 W=0.84 AD=0.378 AS=0.246783 PD=1.74 PS=2.02667 NRD=7.0329 NRS=55.9874
+ M=1 R=5.6 SA=75001 SB=75003.2 A=0.126 P=1.98 MULT=1
MM1003 N_A_1587_74#_M1003_d N_A_630_74#_M1003_g N_A_1257_74#_M1009_d VPB PSHORT
+ L=0.15 W=0.84 AD=0.1932 AS=0.378 PD=1.64 PS=1.74 NRD=3.5066 NRS=118.417 M=1
+ R=5.6 SA=75002.1 SB=75002.1 A=0.126 P=1.98 MULT=1
MM1010 A_1764_476# N_A_828_74#_M1010_g N_A_1587_74#_M1003_d VPB PSHORT L=0.15
+ W=0.42 AD=0.0567 AS=0.0966 PD=0.69 PS=0.82 NRD=37.5088 NRS=44.5417 M=1 R=2.8
+ SA=75002.8 SB=75003.5 A=0.063 P=1.14 MULT=1
MM1021 N_VPWR_M1021_d N_A_1814_48#_M1021_g A_1764_476# VPB PSHORT L=0.15 W=0.42
+ AD=0.0868 AS=0.0567 PD=0.796667 PS=0.69 NRD=4.6886 NRS=37.5088 M=1 R=2.8
+ SA=75003.3 SB=75003 A=0.063 P=1.14 MULT=1
MM1022 N_VPWR_M1021_d N_A_1587_74#_M1022_g N_A_1814_48#_M1022_s VPB PSHORT
+ L=0.15 W=0.84 AD=0.1736 AS=0.126 PD=1.59333 PS=1.14 NRD=15.2281 NRS=2.3443 M=1
+ R=5.6 SA=75002 SB=75002.5 A=0.126 P=1.98 MULT=1
MM1038 N_VPWR_M1038_d N_A_1587_74#_M1038_g N_A_1814_48#_M1022_s VPB PSHORT
+ L=0.15 W=0.84 AD=0.1596 AS=0.126 PD=1.26429 PS=1.14 NRD=12.8838 NRS=2.3443 M=1
+ R=5.6 SA=75002.4 SB=75002.1 A=0.126 P=1.98 MULT=1
MM1000 N_Q_M1000_d N_A_1814_48#_M1000_g N_VPWR_M1038_d VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.2128 PD=1.42 PS=1.68571 NRD=1.7533 NRS=3.5066 M=1 R=7.46667
+ SA=75002.2 SB=75001.6 A=0.168 P=2.54 MULT=1
MM1001 N_Q_M1000_d N_A_1814_48#_M1001_g N_VPWR_M1001_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75002.7 SB=75001.1 A=0.168 P=2.54 MULT=1
MM1031 N_Q_M1031_d N_A_1814_48#_M1031_g N_VPWR_M1001_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75003.1 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1034 N_Q_M1031_d N_A_1814_48#_M1034_g N_VPWR_M1034_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.3304 PD=1.42 PS=2.83 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75003.6 SB=75000.2 A=0.168 P=2.54 MULT=1
DX39_noxref VNB VPB NWDIODE A=23.9196 P=29.44
c_139 VNB 0 1.73925e-19 $X=0 $Y=0
c_247 VPB 0 3.03227e-19 $X=0 $Y=3.085
*
.include "sky130_fd_sc_hs__sdfxtp_4.pxi.spice"
*
.ends
*
*
