* File: sky130_fd_sc_hs__buf_4.spice
* Created: Thu Aug 27 20:34:35 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hs__buf_4.pex.spice"
.subckt sky130_fd_sc_hs__buf_4  VNB VPB A VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A	A
* VPB	VPB
* VNB	VNB
MM1000 N_VGND_M1000_d N_A_86_260#_M1000_g N_X_M1000_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.2627 AS=0.1036 PD=2.19 PS=1.02 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75000.3
+ SB=75002.5 A=0.111 P=1.78 MULT=1
MM1001 N_VGND_M1001_d N_A_86_260#_M1001_g N_X_M1000_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1554 AS=0.1036 PD=1.16 PS=1.02 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75000.7
+ SB=75002.1 A=0.111 P=1.78 MULT=1
MM1002 N_VGND_M1001_d N_A_86_260#_M1002_g N_X_M1002_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1554 AS=0.1036 PD=1.16 PS=1.02 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75001.3
+ SB=75001.5 A=0.111 P=1.78 MULT=1
MM1008 N_VGND_M1008_d N_A_86_260#_M1008_g N_X_M1002_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.2664 AS=0.1036 PD=1.46 PS=1.02 NRD=35.664 NRS=0 M=1 R=4.93333 SA=75001.7
+ SB=75001.1 A=0.111 P=1.78 MULT=1
MM1004 N_A_86_260#_M1004_d N_A_M1004_g N_VGND_M1008_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.2664 PD=2.05 PS=1.46 NRD=0 NRS=35.664 M=1 R=4.93333 SA=75002.6
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1006 N_X_M1006_d N_A_86_260#_M1006_g N_VPWR_M1006_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.3304 PD=1.42 PS=2.83 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75002.3 A=0.168 P=2.54 MULT=1
MM1007 N_X_M1006_d N_A_86_260#_M1007_g N_VPWR_M1007_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.7 SB=75001.9 A=0.168 P=2.54 MULT=1
MM1009 N_X_M1009_d N_A_86_260#_M1009_g N_VPWR_M1007_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.1 SB=75001.4 A=0.168 P=2.54 MULT=1
MM1010 N_X_M1009_d N_A_86_260#_M1010_g N_VPWR_M1010_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.232 PD=1.42 PS=1.72 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.6 SB=75001 A=0.168 P=2.54 MULT=1
MM1003 N_A_86_260#_M1003_d N_A_M1003_g N_VPWR_M1010_s VPB PSHORT L=0.15 W=0.84
+ AD=0.126 AS=0.174 PD=1.14 PS=1.29 NRD=2.3443 NRS=22.261 M=1 R=5.6 SA=75002.1
+ SB=75000.7 A=0.126 P=1.98 MULT=1
MM1005 N_A_86_260#_M1003_d N_A_M1005_g N_VPWR_M1005_s VPB PSHORT L=0.15 W=0.84
+ AD=0.126 AS=0.2478 PD=1.14 PS=2.27 NRD=2.3443 NRS=2.3443 M=1 R=5.6 SA=75002.6
+ SB=75000.2 A=0.126 P=1.98 MULT=1
DX11_noxref VNB VPB NWDIODE A=6.9564 P=11.2
c_33 VNB 0 1.88724e-19 $X=0 $Y=0
*
.include "sky130_fd_sc_hs__buf_4.pxi.spice"
*
.ends
*
*
