* File: sky130_fd_sc_hs__a2bb2o_2.pex.spice
* Created: Thu Aug 27 20:27:45 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HS__A2BB2O_2%B1 2 3 5 6 8 9 10 11
c29 11 0 1.52931e-19 $X=0.24 $Y=1.295
r30 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.27
+ $Y=1.385 $X2=0.27 $Y2=1.385
r31 11 15 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=0.27 $Y=1.295 $X2=0.27
+ $Y2=1.385
r32 9 14 51.5841 $w=3.3e-07 $l=2.95e-07 $layer=POLY_cond $X=0.565 $Y=1.385
+ $X2=0.27 $Y2=1.385
r33 9 10 3.90195 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=0.565 $Y=1.385
+ $X2=0.655 $Y2=1.385
r34 6 10 34.7346 $w=1.65e-07 $l=1.72337e-07 $layer=POLY_cond $X=0.67 $Y=1.22
+ $X2=0.655 $Y2=1.385
r35 6 8 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=0.67 $Y=1.22 $X2=0.67
+ $Y2=0.74
r36 3 5 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=0.655 $Y=1.885
+ $X2=0.655 $Y2=2.46
r37 2 3 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=0.655 $Y=1.795 $X2=0.655
+ $Y2=1.885
r38 1 10 34.7346 $w=1.65e-07 $l=1.65e-07 $layer=POLY_cond $X=0.655 $Y=1.55
+ $X2=0.655 $Y2=1.385
r39 1 2 95.2339 $w=1.8e-07 $l=2.45e-07 $layer=POLY_cond $X=0.655 $Y=1.55
+ $X2=0.655 $Y2=1.795
.ends

.subckt PM_SKY130_FD_SC_HS__A2BB2O_2%B2 3 5 6 8 9 10 14 16
c42 14 0 2.2036e-19 $X=1.12 $Y=1.385
c43 10 0 3.17462e-20 $X=1.2 $Y=1.295
r44 14 17 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.12 $Y=1.385
+ $X2=1.12 $Y2=1.55
r45 14 16 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.12 $Y=1.385
+ $X2=1.12 $Y2=1.22
r46 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.12
+ $Y=1.385 $X2=1.12 $Y2=1.385
r47 10 15 2.49177 $w=3.68e-07 $l=8e-08 $layer=LI1_cond $X=1.2 $Y=1.365 $X2=1.12
+ $Y2=1.365
r48 9 15 12.4588 $w=3.68e-07 $l=4e-07 $layer=LI1_cond $X=0.72 $Y=1.365 $X2=1.12
+ $Y2=1.365
r49 6 8 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=1.105 $Y=1.885
+ $X2=1.105 $Y2=2.46
r50 5 6 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=1.105 $Y=1.795 $X2=1.105
+ $Y2=1.885
r51 5 17 95.2339 $w=1.8e-07 $l=2.45e-07 $layer=POLY_cond $X=1.105 $Y=1.795
+ $X2=1.105 $Y2=1.55
r52 3 16 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.03 $Y=0.74 $X2=1.03
+ $Y2=1.22
.ends

.subckt PM_SKY130_FD_SC_HS__A2BB2O_2%A_293_333# 1 2 7 9 10 12 18 19 20 21 22 24
+ 28
c78 22 0 1.59253e-19 $X=2.422 $Y=1.85
c79 18 0 9.91756e-20 $X=2.01 $Y=1.385
r80 26 28 12.0152 $w=1.78e-07 $l=1.95e-07 $layer=LI1_cond $X=2.78 $Y=0.84
+ $X2=2.78 $Y2=0.645
r81 22 24 7.3171 $w=3.13e-07 $l=2e-07 $layer=LI1_cond $X=2.422 $Y=1.85 $X2=2.422
+ $Y2=2.05
r82 20 26 6.82373 $w=1.7e-07 $l=1.25499e-07 $layer=LI1_cond $X=2.69 $Y=0.925
+ $X2=2.78 $Y2=0.84
r83 20 21 33.5989 $w=1.68e-07 $l=5.15e-07 $layer=LI1_cond $X=2.69 $Y=0.925
+ $X2=2.175 $Y2=0.925
r84 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.01
+ $Y=1.385 $X2=2.01 $Y2=1.385
r85 16 22 24.2695 $w=1.68e-07 $l=3.72e-07 $layer=LI1_cond $X=2.05 $Y=1.765
+ $X2=2.422 $Y2=1.765
r86 16 18 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=2.05 $Y=1.68
+ $X2=2.05 $Y2=1.385
r87 15 21 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=2.05 $Y=1.01
+ $X2=2.175 $Y2=0.925
r88 15 18 17.2866 $w=2.48e-07 $l=3.75e-07 $layer=LI1_cond $X=2.05 $Y=1.01
+ $X2=2.05 $Y2=1.385
r89 14 19 63.8244 $w=3.3e-07 $l=3.65e-07 $layer=POLY_cond $X=1.645 $Y=1.385
+ $X2=2.01 $Y2=1.385
r90 10 14 50.2292 $w=1.59e-07 $l=1.72337e-07 $layer=POLY_cond $X=1.57 $Y=1.22
+ $X2=1.555 $Y2=1.385
r91 10 12 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.57 $Y=1.22 $X2=1.57
+ $Y2=0.74
r92 7 14 151.783 $w=1.59e-07 $l=5e-07 $layer=POLY_cond $X=1.555 $Y=1.885
+ $X2=1.555 $Y2=1.385
r93 7 9 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=1.555 $Y=1.885
+ $X2=1.555 $Y2=2.46
r94 2 24 300 $w=1.7e-07 $l=2.13542e-07 $layer=licon1_PDIFF $count=2 $X=2.305
+ $Y=1.89 $X2=2.43 $Y2=2.05
r95 1 28 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=2.645
+ $Y=0.37 $X2=2.785 $Y2=0.645
.ends

.subckt PM_SKY130_FD_SC_HS__A2BB2O_2%A2_N 3 7 9 10 11 14
r41 14 17 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.55 $Y=1.345
+ $X2=2.55 $Y2=1.51
r42 14 16 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.55 $Y=1.345
+ $X2=2.55 $Y2=1.18
r43 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.55
+ $Y=1.345 $X2=2.55 $Y2=1.345
r44 11 15 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=2.64 $Y=1.345 $X2=2.55
+ $Y2=1.345
r45 10 17 76.9149 $w=1.5e-07 $l=1.5e-07 $layer=POLY_cond $X=2.64 $Y=1.66
+ $X2=2.64 $Y2=1.51
r46 7 10 60.25 $w=1.8e-07 $l=1.55e-07 $layer=POLY_cond $X=2.655 $Y=1.815
+ $X2=2.655 $Y2=1.66
r47 7 9 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=2.655 $Y=1.815
+ $X2=2.655 $Y2=2.39
r48 3 16 274.33 $w=1.5e-07 $l=5.35e-07 $layer=POLY_cond $X=2.57 $Y=0.645
+ $X2=2.57 $Y2=1.18
.ends

.subckt PM_SKY130_FD_SC_HS__A2BB2O_2%A1_N 3 6 7 9 10 11 12 17
c47 7 0 3.18369e-20 $X=3.045 $Y=1.815
c48 6 0 1.27416e-19 $X=3.045 $Y=1.725
r49 17 20 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.09 $Y=1.385
+ $X2=3.09 $Y2=1.55
r50 17 19 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.09 $Y=1.385
+ $X2=3.09 $Y2=1.22
r51 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.09
+ $Y=1.385 $X2=3.09 $Y2=1.385
r52 11 12 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=3.09 $Y=1.665
+ $X2=3.09 $Y2=2.035
r53 11 18 9.7783 $w=3.28e-07 $l=2.8e-07 $layer=LI1_cond $X=3.09 $Y=1.665
+ $X2=3.09 $Y2=1.385
r54 10 18 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=3.09 $Y=1.295 $X2=3.09
+ $Y2=1.385
r55 7 9 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=3.045 $Y=1.815
+ $X2=3.045 $Y2=2.39
r56 6 7 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=3.045 $Y=1.725 $X2=3.045
+ $Y2=1.815
r57 6 20 68.0242 $w=1.8e-07 $l=1.75e-07 $layer=POLY_cond $X=3.045 $Y=1.725
+ $X2=3.045 $Y2=1.55
r58 3 19 294.84 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=3 $Y=0.645 $X2=3
+ $Y2=1.22
.ends

.subckt PM_SKY130_FD_SC_HS__A2BB2O_2%A_221_74# 1 2 9 11 13 14 18 20 22 23 27 30
+ 34 35 39 40 43 47 50 53 54 58
c112 38 0 4.64943e-20 $X=2.835 $Y=2.81
r113 57 58 4.69916 $w=3.59e-07 $l=3.5e-08 $layer=POLY_cond $X=3.97 $Y=1.557
+ $X2=4.005 $Y2=1.557
r114 53 54 5.95004 $w=3.58e-07 $l=8.5e-08 $layer=LI1_cond $X=1.765 $Y=2.105
+ $X2=1.765 $Y2=2.02
r115 48 50 6.52406 $w=1.68e-07 $l=1e-07 $layer=LI1_cond $X=1.57 $Y=1.465
+ $X2=1.67 $Y2=1.465
r116 46 47 8.79167 $w=3.98e-07 $l=1.7e-07 $layer=LI1_cond $X=1.367 $Y=0.84
+ $X2=1.367 $Y2=1.01
r117 44 58 33.5655 $w=3.59e-07 $l=2.5e-07 $layer=POLY_cond $X=4.255 $Y=1.557
+ $X2=4.005 $Y2=1.557
r118 43 44 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.255
+ $Y=1.515 $X2=4.255 $Y2=1.515
r119 41 43 24.4136 $w=3.78e-07 $l=8.05e-07 $layer=LI1_cond $X=4.28 $Y=2.32
+ $X2=4.28 $Y2=1.515
r120 39 41 8.19669 $w=1.7e-07 $l=2.28583e-07 $layer=LI1_cond $X=4.09 $Y=2.405
+ $X2=4.28 $Y2=2.32
r121 39 40 76.3316 $w=1.68e-07 $l=1.17e-06 $layer=LI1_cond $X=4.09 $Y=2.405
+ $X2=2.92 $Y2=2.405
r122 37 40 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.835 $Y=2.49
+ $X2=2.92 $Y2=2.405
r123 37 38 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=2.835 $Y=2.49
+ $X2=2.835 $Y2=2.81
r124 36 56 5.44966 $w=1.7e-07 $l=1.8e-07 $layer=LI1_cond $X=1.945 $Y=2.895
+ $X2=1.765 $Y2=2.895
r125 35 38 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.75 $Y=2.895
+ $X2=2.835 $Y2=2.81
r126 35 36 52.5187 $w=1.68e-07 $l=8.05e-07 $layer=LI1_cond $X=2.75 $Y=2.895
+ $X2=1.945 $Y2=2.895
r127 34 56 2.57345 $w=3.6e-07 $l=8.5e-08 $layer=LI1_cond $X=1.765 $Y=2.81
+ $X2=1.765 $Y2=2.895
r128 33 53 3.04117 $w=3.58e-07 $l=9.5e-08 $layer=LI1_cond $X=1.765 $Y=2.2
+ $X2=1.765 $Y2=2.105
r129 33 34 19.5275 $w=3.58e-07 $l=6.1e-07 $layer=LI1_cond $X=1.765 $Y=2.2
+ $X2=1.765 $Y2=2.81
r130 31 50 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.67 $Y=1.55
+ $X2=1.67 $Y2=1.465
r131 31 54 30.6631 $w=1.68e-07 $l=4.7e-07 $layer=LI1_cond $X=1.67 $Y=1.55
+ $X2=1.67 $Y2=2.02
r132 30 48 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.57 $Y=1.38
+ $X2=1.57 $Y2=1.465
r133 30 47 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=1.57 $Y=1.38
+ $X2=1.57 $Y2=1.01
r134 27 46 9.93982 $w=3.98e-07 $l=3.45e-07 $layer=LI1_cond $X=1.28 $Y=0.495
+ $X2=1.28 $Y2=0.84
r135 23 24 31.303 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=3.555 $Y=1.605
+ $X2=3.555 $Y2=1.53
r136 20 58 23.2387 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=4.005 $Y=1.765
+ $X2=4.005 $Y2=1.557
r137 20 22 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=4.005 $Y=1.765
+ $X2=4.005 $Y2=2.4
r138 16 57 23.2387 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.97 $Y=1.35
+ $X2=3.97 $Y2=1.557
r139 16 18 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=3.97 $Y=1.35
+ $X2=3.97 $Y2=0.74
r140 15 23 7.1379 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=3.645 $Y=1.605
+ $X2=3.555 $Y2=1.605
r141 14 57 26.8132 $w=3.59e-07 $l=9.60469e-08 $layer=POLY_cond $X=3.895 $Y=1.605
+ $X2=3.97 $Y2=1.557
r142 14 15 128.191 $w=1.5e-07 $l=2.5e-07 $layer=POLY_cond $X=3.895 $Y=1.605
+ $X2=3.645 $Y2=1.605
r143 11 23 64.3434 $w=1.8e-07 $l=1.6e-07 $layer=POLY_cond $X=3.555 $Y=1.765
+ $X2=3.555 $Y2=1.605
r144 11 13 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.555 $Y=1.765
+ $X2=3.555 $Y2=2.4
r145 9 24 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=3.54 $Y=0.74
+ $X2=3.54 $Y2=1.53
r146 2 56 400 $w=1.7e-07 $l=9.26971e-07 $layer=licon1_PDIFF $count=1 $X=1.63
+ $Y=1.96 $X2=1.78 $Y2=2.815
r147 2 53 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=1.63
+ $Y=1.96 $X2=1.78 $Y2=2.105
r148 1 27 91 $w=1.7e-07 $l=2.498e-07 $layer=licon1_NDIFF $count=2 $X=1.105
+ $Y=0.37 $X2=1.3 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_HS__A2BB2O_2%A_61_392# 1 2 9 13 14 17
r27 17 19 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=1.33 $Y=2.105
+ $X2=1.33 $Y2=2.815
r28 15 17 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=1.33 $Y=1.89
+ $X2=1.33 $Y2=2.105
r29 13 15 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.245 $Y=1.805
+ $X2=1.33 $Y2=1.89
r30 13 14 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=1.245 $Y=1.805
+ $X2=0.515 $Y2=1.805
r31 9 11 32.7294 $w=2.48e-07 $l=7.1e-07 $layer=LI1_cond $X=0.39 $Y=2.105
+ $X2=0.39 $Y2=2.815
r32 7 14 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.39 $Y=1.89
+ $X2=0.515 $Y2=1.805
r33 7 9 9.91101 $w=2.48e-07 $l=2.15e-07 $layer=LI1_cond $X=0.39 $Y=1.89 $X2=0.39
+ $Y2=2.105
r34 2 19 400 $w=1.7e-07 $l=9.26971e-07 $layer=licon1_PDIFF $count=1 $X=1.18
+ $Y=1.96 $X2=1.33 $Y2=2.815
r35 2 17 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=1.18
+ $Y=1.96 $X2=1.33 $Y2=2.105
r36 1 11 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=0.305
+ $Y=1.96 $X2=0.43 $Y2=2.815
r37 1 9 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.305
+ $Y=1.96 $X2=0.43 $Y2=2.105
.ends

.subckt PM_SKY130_FD_SC_HS__A2BB2O_2%VPWR 1 2 3 14 18 20 24 26 28 35 36 39 42 45
r53 45 46 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r54 43 46 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=4.08 $Y2=3.33
r55 42 43 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r56 39 40 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r57 36 46 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=4.08 $Y2=3.33
r58 35 36 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r59 33 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.395 $Y=3.33
+ $X2=4.23 $Y2=3.33
r60 33 35 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=4.395 $Y=3.33
+ $X2=4.56 $Y2=3.33
r61 32 40 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r62 31 32 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r63 29 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.045 $Y=3.33
+ $X2=0.88 $Y2=3.33
r64 29 31 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=1.045 $Y=3.33
+ $X2=1.2 $Y2=3.33
r65 28 42 9.6488 $w=1.7e-07 $l=1.95e-07 $layer=LI1_cond $X=3.105 $Y=3.33 $X2=3.3
+ $Y2=3.33
r66 28 31 124.283 $w=1.68e-07 $l=1.905e-06 $layer=LI1_cond $X=3.105 $Y=3.33
+ $X2=1.2 $Y2=3.33
r67 26 43 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=2.4 $Y=3.33
+ $X2=3.12 $Y2=3.33
r68 26 32 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=2.4 $Y=3.33 $X2=1.2
+ $Y2=3.33
r69 22 45 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.23 $Y=3.245
+ $X2=4.23 $Y2=3.33
r70 22 24 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=4.23 $Y=3.245
+ $X2=4.23 $Y2=2.78
r71 21 42 9.6488 $w=1.7e-07 $l=1.95e-07 $layer=LI1_cond $X=3.495 $Y=3.33 $X2=3.3
+ $Y2=3.33
r72 20 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.065 $Y=3.33
+ $X2=4.23 $Y2=3.33
r73 20 21 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=4.065 $Y=3.33
+ $X2=3.495 $Y2=3.33
r74 16 42 1.39532 $w=3.9e-07 $l=8.5e-08 $layer=LI1_cond $X=3.3 $Y=3.245 $X2=3.3
+ $Y2=3.33
r75 16 18 14.7749 $w=3.88e-07 $l=5e-07 $layer=LI1_cond $X=3.3 $Y=3.245 $X2=3.3
+ $Y2=2.745
r76 12 39 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.88 $Y=3.245
+ $X2=0.88 $Y2=3.33
r77 12 14 35.621 $w=3.28e-07 $l=1.02e-06 $layer=LI1_cond $X=0.88 $Y=3.245
+ $X2=0.88 $Y2=2.225
r78 3 24 600 $w=1.7e-07 $l=1.01223e-06 $layer=licon1_PDIFF $count=1 $X=4.08
+ $Y=1.84 $X2=4.23 $Y2=2.78
r79 2 18 600 $w=1.7e-07 $l=9.40705e-07 $layer=licon1_PDIFF $count=1 $X=3.12
+ $Y=1.89 $X2=3.3 $Y2=2.745
r80 1 14 300 $w=1.7e-07 $l=3.31625e-07 $layer=licon1_PDIFF $count=2 $X=0.73
+ $Y=1.96 $X2=0.88 $Y2=2.225
.ends

.subckt PM_SKY130_FD_SC_HS__A2BB2O_2%X 1 2 7 8 9 10 11 18
r22 11 29 1.32465 $w=4.33e-07 $l=5e-08 $layer=LI1_cond $X=3.702 $Y=2.035
+ $X2=3.702 $Y2=1.985
r23 10 29 8.47774 $w=4.33e-07 $l=3.2e-07 $layer=LI1_cond $X=3.702 $Y=1.665
+ $X2=3.702 $Y2=1.985
r24 9 10 9.80239 $w=4.33e-07 $l=3.7e-07 $layer=LI1_cond $X=3.702 $Y=1.295
+ $X2=3.702 $Y2=1.665
r25 8 9 9.80239 $w=4.33e-07 $l=3.7e-07 $layer=LI1_cond $X=3.702 $Y=0.925
+ $X2=3.702 $Y2=1.295
r26 7 8 9.80239 $w=4.33e-07 $l=3.7e-07 $layer=LI1_cond $X=3.702 $Y=0.555
+ $X2=3.702 $Y2=0.925
r27 7 18 1.05972 $w=4.33e-07 $l=4e-08 $layer=LI1_cond $X=3.702 $Y=0.555
+ $X2=3.702 $Y2=0.515
r28 2 29 600 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=3.63
+ $Y=1.84 $X2=3.78 $Y2=1.985
r29 1 18 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.615
+ $Y=0.37 $X2=3.755 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__A2BB2O_2%VGND 1 2 3 4 15 17 21 25 28 29 31 32 33 47
+ 48 53 59 61
r64 61 62 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r65 58 59 11.1544 $w=7.53e-07 $l=1.65e-07 $layer=LI1_cond $X=2.355 $Y=0.292
+ $X2=2.52 $Y2=0.292
r66 55 58 3.08921 $w=7.53e-07 $l=1.95e-07 $layer=LI1_cond $X=2.16 $Y=0.292
+ $X2=2.355 $Y2=0.292
r67 55 56 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r68 52 56 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r69 51 55 7.60421 $w=7.53e-07 $l=4.8e-07 $layer=LI1_cond $X=1.68 $Y=0.292
+ $X2=2.16 $Y2=0.292
r70 51 53 9.01574 $w=7.53e-07 $l=3e-08 $layer=LI1_cond $X=1.68 $Y=0.292 $X2=1.65
+ $Y2=0.292
r71 51 52 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r72 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r73 45 48 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=4.56
+ $Y2=0
r74 45 62 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=3.12
+ $Y2=0
r75 44 45 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r76 42 61 7.34436 $w=1.7e-07 $l=1.33e-07 $layer=LI1_cond $X=3.315 $Y=0 $X2=3.182
+ $Y2=0
r77 42 44 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=3.315 $Y=0 $X2=4.08
+ $Y2=0
r78 41 52 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r79 40 53 60.6738 $w=1.68e-07 $l=9.3e-07 $layer=LI1_cond $X=0.72 $Y=0 $X2=1.65
+ $Y2=0
r80 40 41 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r81 37 41 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r82 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r83 33 62 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=2.4 $Y=0 $X2=3.12
+ $Y2=0
r84 33 56 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.4 $Y=0 $X2=2.16
+ $Y2=0
r85 31 44 1.30481 $w=1.68e-07 $l=2e-08 $layer=LI1_cond $X=4.1 $Y=0 $X2=4.08
+ $Y2=0
r86 31 32 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.1 $Y=0 $X2=4.225
+ $Y2=0
r87 30 47 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=4.35 $Y=0 $X2=4.56
+ $Y2=0
r88 30 32 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.35 $Y=0 $X2=4.225
+ $Y2=0
r89 28 36 3.58824 $w=1.7e-07 $l=5e-08 $layer=LI1_cond $X=0.29 $Y=0 $X2=0.24
+ $Y2=0
r90 28 29 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.29 $Y=0 $X2=0.455
+ $Y2=0
r91 27 40 6.52406 $w=1.68e-07 $l=1e-07 $layer=LI1_cond $X=0.62 $Y=0 $X2=0.72
+ $Y2=0
r92 27 29 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.62 $Y=0 $X2=0.455
+ $Y2=0
r93 23 32 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.225 $Y=0.085
+ $X2=4.225 $Y2=0
r94 23 25 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=4.225 $Y=0.085
+ $X2=4.225 $Y2=0.515
r95 19 61 0.195364 $w=2.65e-07 $l=8.5e-08 $layer=LI1_cond $X=3.182 $Y=0.085
+ $X2=3.182 $Y2=0
r96 19 21 24.3535 $w=2.63e-07 $l=5.6e-07 $layer=LI1_cond $X=3.182 $Y=0.085
+ $X2=3.182 $Y2=0.645
r97 17 61 7.34436 $w=1.7e-07 $l=1.32e-07 $layer=LI1_cond $X=3.05 $Y=0 $X2=3.182
+ $Y2=0
r98 17 59 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=3.05 $Y=0 $X2=2.52
+ $Y2=0
r99 13 29 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.455 $Y=0.085
+ $X2=0.455 $Y2=0
r100 13 15 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=0.455 $Y=0.085
+ $X2=0.455 $Y2=0.515
r101 4 25 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=4.045
+ $Y=0.37 $X2=4.185 $Y2=0.515
r102 3 21 182 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_NDIFF $count=1 $X=3.075
+ $Y=0.37 $X2=3.22 $Y2=0.645
r103 2 58 91 $w=1.7e-07 $l=7.94921e-07 $layer=licon1_NDIFF $count=2 $X=1.645
+ $Y=0.37 $X2=2.355 $Y2=0.55
r104 1 15 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.31
+ $Y=0.37 $X2=0.455 $Y2=0.515
.ends

