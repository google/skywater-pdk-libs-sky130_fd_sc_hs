* NGSPICE file created from sky130_fd_sc_hs__dlrtp_4.ext - technology: sky130A

.subckt sky130_fd_sc_hs__dlrtp_4 D GATE RESET_B VGND VNB VPB VPWR Q
M1000 a_938_74# a_640_74# a_797_48# VNB nlowvt w=640000u l=150000u
+  ad=5.44e+11p pd=5.54e+06u as=1.824e+11p ps=1.85e+06u
M1001 a_559_74# a_27_126# VGND VNB nlowvt w=640000u l=150000u
+  ad=1.632e+11p pd=1.79e+06u as=1.6158e+12p ps=1.463e+07u
M1002 a_755_74# a_240_394# a_640_74# VNB nlowvt w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=2.555e+11p ps=2.13e+06u
M1003 VPWR a_797_48# a_747_508# VPB pshort w=420000u l=150000u
+  ad=2.7109e+12p pd=2.052e+07u as=1.995e+11p ps=1.79e+06u
M1004 a_240_394# GATE VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1005 a_747_508# a_364_120# a_640_74# VPB pshort w=420000u l=150000u
+  ad=0p pd=0u as=3.328e+11p ps=2.77e+06u
M1006 a_797_48# a_640_74# a_938_74# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_240_394# GATE VPWR VPB pshort w=840000u l=150000u
+  ad=2.94e+11p pd=2.38e+06u as=0p ps=0u
M1008 a_640_74# a_240_394# a_562_392# VPB pshort w=1e+06u l=150000u
+  ad=0p pd=0u as=2.4e+11p ps=2.48e+06u
M1009 VPWR D a_27_126# VPB pshort w=840000u l=150000u
+  ad=0p pd=0u as=2.478e+11p ps=2.27e+06u
M1010 Q a_797_48# VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=7.504e+11p pd=5.82e+06u as=0p ps=0u
M1011 Q a_797_48# VGND VNB nlowvt w=740000u l=150000u
+  ad=4.144e+11p pd=4.08e+06u as=0p ps=0u
M1012 VPWR a_797_48# Q VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 Q a_797_48# VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 VPWR a_797_48# Q VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 Q a_797_48# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VPWR a_240_394# a_364_120# VPB pshort w=840000u l=150000u
+  ad=0p pd=0u as=2.478e+11p ps=2.27e+06u
M1017 a_797_48# a_640_74# VPWR VPB pshort w=840000u l=150000u
+  ad=5.46e+11p pd=4.66e+06u as=0p ps=0u
M1018 a_562_392# a_27_126# VPWR VPB pshort w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VGND D a_27_126# VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=1.5675e+11p ps=1.67e+06u
M1020 VGND RESET_B a_938_74# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_797_48# RESET_B VPWR VPB pshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 VPWR RESET_B a_797_48# VPB pshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 VGND a_797_48# Q VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 VGND a_240_394# a_364_120# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.294e+11p ps=2.1e+06u
M1025 VPWR a_640_74# a_797_48# VPB pshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 VGND a_797_48# a_755_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 a_640_74# a_364_120# a_559_74# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1028 a_938_74# RESET_B VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1029 VGND a_797_48# Q VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

