* File: sky130_fd_sc_hs__a31o_2.spice
* Created: Thu Aug 27 20:29:15 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hs__a31o_2.pex.spice"
.subckt sky130_fd_sc_hs__a31o_2  VNB VPB A3 A2 A1 B1 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* B1	B1
* A1	A1
* A2	A2
* A3	A3
* VPB	VPB
* VNB	VNB
MM1005 N_VGND_M1005_d N_A_97_296#_M1005_g N_X_M1005_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.2627 AS=0.1036 PD=2.19 PS=1.02 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75000.3
+ SB=75003 A=0.111 P=1.78 MULT=1
MM1006 N_VGND_M1006_d N_A_97_296#_M1006_g N_X_M1005_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.23495 AS=0.1036 PD=1.375 PS=1.02 NRD=2.424 NRS=0 M=1 R=4.93333 SA=75000.7
+ SB=75002.5 A=0.111 P=1.78 MULT=1
MM1002 A_371_74# N_A3_M1002_g N_VGND_M1006_d VNB NLOWVT L=0.15 W=0.74 AD=0.0888
+ AS=0.23495 PD=0.98 PS=1.375 NRD=10.536 NRS=0 M=1 R=4.93333 SA=75001.5
+ SB=75001.7 A=0.111 P=1.78 MULT=1
MM1004 A_449_74# N_A2_M1004_g A_371_74# VNB NLOWVT L=0.15 W=0.74 AD=0.1554
+ AS=0.0888 PD=1.16 PS=0.98 NRD=25.128 NRS=10.536 M=1 R=4.93333 SA=75001.9
+ SB=75001.4 A=0.111 P=1.78 MULT=1
MM1007 N_A_97_296#_M1007_d N_A1_M1007_g A_449_74# VNB NLOWVT L=0.15 W=0.74
+ AD=0.1554 AS=0.1554 PD=1.16 PS=1.16 NRD=9.72 NRS=25.128 M=1 R=4.93333
+ SA=75002.5 SB=75000.8 A=0.111 P=1.78 MULT=1
MM1000 N_VGND_M1000_d N_B1_M1000_g N_A_97_296#_M1007_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.1554 PD=2.05 PS=1.16 NRD=0 NRS=12.972 M=1 R=4.93333 SA=75003
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1008 N_X_M1008_d N_A_97_296#_M1008_g N_VPWR_M1008_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.3304 PD=1.42 PS=2.83 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75002.7 A=0.168 P=2.54 MULT=1
MM1009 N_X_M1008_d N_A_97_296#_M1009_g N_VPWR_M1009_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.323743 PD=1.42 PS=1.77509 NRD=1.7533 NRS=17.2769 M=1 R=7.46667
+ SA=75000.7 SB=75002.3 A=0.168 P=2.54 MULT=1
MM1010 N_A_362_368#_M1010_d N_A3_M1010_g N_VPWR_M1009_s VPB PSHORT L=0.15 W=1
+ AD=0.15 AS=0.289057 PD=1.3 PS=1.58491 NRD=1.9503 NRS=36.1101 M=1 R=6.66667
+ SA=75001.4 SB=75001.8 A=0.15 P=2.3 MULT=1
MM1011 N_VPWR_M1011_d N_A2_M1011_g N_A_362_368#_M1010_d VPB PSHORT L=0.15 W=1
+ AD=0.245 AS=0.15 PD=1.49 PS=1.3 NRD=22.6353 NRS=1.9503 M=1 R=6.66667
+ SA=75001.8 SB=75001.4 A=0.15 P=2.3 MULT=1
MM1003 N_A_362_368#_M1003_d N_A1_M1003_g N_VPWR_M1011_d VPB PSHORT L=0.15 W=1
+ AD=0.175 AS=0.245 PD=1.35 PS=1.49 NRD=1.9503 NRS=18.715 M=1 R=6.66667
+ SA=75002.5 SB=75000.7 A=0.15 P=2.3 MULT=1
MM1001 N_A_97_296#_M1001_d N_B1_M1001_g N_A_362_368#_M1003_d VPB PSHORT L=0.15
+ W=1 AD=0.305 AS=0.175 PD=2.61 PS=1.35 NRD=2.9353 NRS=11.8003 M=1 R=6.66667
+ SA=75003 SB=75000.2 A=0.15 P=2.3 MULT=1
DX12_noxref VNB VPB NWDIODE A=7.8492 P=12.16
*
.include "sky130_fd_sc_hs__a31o_2.pxi.spice"
*
.ends
*
*
