* File: sky130_fd_sc_hs__fah_1.spice
* Created: Tue Sep  1 20:05:39 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hs__fah_1.pex.spice"
.subckt sky130_fd_sc_hs__fah_1  VNB VPB CI B A SUM VPWR COUT VGND
* 
* VGND	VGND
* COUT	COUT
* VPWR	VPWR
* SUM	SUM
* A	A
* B	B
* CI	CI
* VPB	VPB
* VNB	VNB
MM1029 N_VGND_M1029_d N_A_83_21#_M1029_g N_SUM_M1029_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.206342 AS=0.2072 PD=1.51217 PS=2.04 NRD=36.288 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75000.8 A=0.111 P=1.78 MULT=1
MM1010 N_A_231_132#_M1010_d N_CI_M1010_g N_VGND_M1029_d VNB NLOWVT L=0.15 W=0.64
+ AD=0.2016 AS=0.178458 PD=1.91 PS=1.30783 NRD=2.808 NRS=41.964 M=1 R=4.26667
+ SA=75000.8 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1006 N_VGND_M1006_d N_A_410_58#_M1006_g N_COUT_M1006_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.313857 AS=0.2072 PD=1.72667 PS=2.04 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75001.2 A=0.111 P=1.78 MULT=1
MM1028 N_A_644_104#_M1028_d N_A_231_132#_M1028_g N_VGND_M1006_d VNB NLOWVT
+ L=0.15 W=0.64 AD=0.23505 AS=0.271443 PD=2.02 PS=1.49333 NRD=14.988 NRS=111.552
+ M=1 R=4.26667 SA=75001.2 SB=75000.3 A=0.096 P=1.58 MULT=1
MM1000 N_A_410_58#_M1000_d N_A_811_379#_M1000_g N_A_879_55#_M1000_s VNB NLOWVT
+ L=0.15 W=0.64 AD=0.131975 AS=0.28315 PD=1.205 PS=3.17 NRD=0 NRS=72.636 M=1
+ R=4.26667 SA=75000.2 SB=75001.1 A=0.096 P=1.58 MULT=1
MM1012 N_A_231_132#_M1012_d N_A_1023_379#_M1012_g N_A_410_58#_M1000_d VNB NLOWVT
+ L=0.15 W=0.64 AD=0.0896 AS=0.131975 PD=0.92 PS=1.205 NRD=0 NRS=14.988 M=1
+ R=4.26667 SA=75000.5 SB=75001.1 A=0.096 P=1.58 MULT=1
MM1001 N_A_83_21#_M1001_d N_A_811_379#_M1001_g N_A_231_132#_M1012_d VNB NLOWVT
+ L=0.15 W=0.64 AD=0.11875 AS=0.0896 PD=1.08 PS=0.92 NRD=13.116 NRS=0 M=1
+ R=4.26667 SA=75000.9 SB=75000.6 A=0.096 P=1.58 MULT=1
MM1020 N_A_644_104#_M1020_d N_A_1023_379#_M1020_g N_A_83_21#_M1001_d VNB NLOWVT
+ L=0.15 W=0.64 AD=0.1824 AS=0.11875 PD=1.85 PS=1.08 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75001.2 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1026 N_VGND_M1026_d N_B_M1026_g N_A_879_55#_M1026_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.3136 AS=0.2109 PD=2.51 PS=2.05 NRD=13.776 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75000.3 A=0.111 P=1.78 MULT=1
MM1004 N_A_1023_379#_M1004_d N_A_879_55#_M1004_g N_A_1660_374#_M1004_s VNB
+ NLOWVT L=0.15 W=0.64 AD=0.24825 AS=0.2568 PD=1.49 PS=2.17 NRD=62.412
+ NRS=15.936 M=1 R=4.26667 SA=75000.3 SB=75003.3 A=0.096 P=1.58 MULT=1
MM1030 N_A_1849_374#_M1030_d N_B_M1030_g N_A_1023_379#_M1004_d VNB NLOWVT L=0.15
+ W=0.64 AD=0.1524 AS=0.24825 PD=1.16 PS=1.49 NRD=15.936 NRS=62.412 M=1
+ R=4.26667 SA=75001 SB=75002.6 A=0.096 P=1.58 MULT=1
MM1002 N_A_811_379#_M1002_d N_A_879_55#_M1002_g N_A_1849_374#_M1030_d VNB NLOWVT
+ L=0.15 W=0.64 AD=0.3264 AS=0.1524 PD=1.66 PS=1.16 NRD=61.872 NRS=15.936 M=1
+ R=4.26667 SA=75001.6 SB=75002 A=0.096 P=1.58 MULT=1
MM1027 N_A_1660_374#_M1027_d N_B_M1027_g N_A_811_379#_M1002_d VNB NLOWVT L=0.15
+ W=0.64 AD=0.12007 AS=0.3264 PD=1.02029 PS=1.66 NRD=15.468 NRS=76.872 M=1
+ R=4.26667 SA=75002.8 SB=75000.8 A=0.096 P=1.58 MULT=1
MM1025 N_VGND_M1025_d N_A_2342_48#_M1025_g N_A_1660_374#_M1027_d VNB NLOWVT
+ L=0.15 W=0.74 AD=0.2875 AS=0.13883 PD=2.33 PS=1.17971 NRD=13.776 NRS=0 M=1
+ R=4.93333 SA=75002.9 SB=75000.3 A=0.111 P=1.78 MULT=1
MM1014 N_VGND_M1014_d N_A_M1014_g N_A_1849_374#_M1014_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.1216 AS=0.208 PD=1.02 PS=1.93 NRD=5.616 NRS=7.488 M=1 R=4.26667
+ SA=75000.2 SB=75000.7 A=0.096 P=1.58 MULT=1
MM1011 N_A_2342_48#_M1011_d N_A_M1011_g N_VGND_M1014_d VNB NLOWVT L=0.15 W=0.64
+ AD=0.1824 AS=0.1216 PD=1.85 PS=1.02 NRD=0 NRS=13.116 M=1 R=4.26667 SA=75000.8
+ SB=75000.2 A=0.096 P=1.58 MULT=1
MM1021 N_VPWR_M1021_d N_A_83_21#_M1021_g N_SUM_M1021_s VPB PSHORT L=0.15 W=1.12
+ AD=0.298226 AS=0.3304 PD=1.7434 PS=2.83 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75000.8 A=0.168 P=2.54 MULT=1
MM1022 N_A_231_132#_M1022_d N_CI_M1022_g N_VPWR_M1021_d VPB PSHORT L=0.15 W=1
+ AD=0.295 AS=0.266274 PD=2.59 PS=1.5566 NRD=1.9503 NRS=47.7528 M=1 R=6.66667
+ SA=75000.9 SB=75000.2 A=0.15 P=2.3 MULT=1
MM1015 N_VPWR_M1015_d N_A_410_58#_M1015_g N_COUT_M1015_s VPB PSHORT L=0.15
+ W=1.12 AD=0.322964 AS=0.46765 PD=1.95472 PS=3.29 NRD=41.0351 NRS=17.5724 M=1
+ R=7.46667 SA=75000.3 SB=75003.4 A=0.168 P=2.54 MULT=1
MM1024 N_A_644_104#_M1024_d N_A_231_132#_M1024_g N_VPWR_M1015_d VPB PSHORT
+ L=0.15 W=1 AD=0.303655 AS=0.288361 PD=1.77717 PS=1.74528 NRD=18.715
+ NRS=45.9601 M=1 R=6.66667 SA=75000.9 SB=75003.1 A=0.15 P=2.3 MULT=1
MM1023 N_A_83_21#_M1023_d N_A_811_379#_M1023_g N_A_644_104#_M1024_d VPB PSHORT
+ L=0.15 W=0.84 AD=0.3822 AS=0.25507 PD=1.75 PS=1.49283 NRD=2.3443 NRS=58.312
+ M=1 R=5.6 SA=75001.5 SB=75003.1 A=0.126 P=1.98 MULT=1
MM1005 N_A_231_132#_M1005_d N_A_1023_379#_M1005_g N_A_83_21#_M1023_d VPB PSHORT
+ L=0.15 W=0.84 AD=0.406612 AS=0.3822 PD=2.01 PS=1.75 NRD=2.3443 NRS=145.386 M=1
+ R=5.6 SA=75002.6 SB=75002.1 A=0.126 P=1.98 MULT=1
MM1017 N_A_410_58#_M1017_d N_A_811_379#_M1017_g N_A_231_132#_M1005_d VPB PSHORT
+ L=0.15 W=0.84 AD=0.2541 AS=0.406612 PD=1.445 PS=2.01 NRD=2.3443 NRS=100.608
+ M=1 R=5.6 SA=75002.7 SB=75001.6 A=0.126 P=1.98 MULT=1
MM1003 N_A_879_55#_M1003_d N_A_1023_379#_M1003_g N_A_410_58#_M1017_d VPB PSHORT
+ L=0.15 W=0.84 AD=0.172971 AS=0.2541 PD=1.29 PS=1.445 NRD=22.655 NRS=73.8553
+ M=1 R=5.6 SA=75003.4 SB=75000.8 A=0.126 P=1.98 MULT=1
MM1031 N_VPWR_M1031_d N_B_M1031_g N_A_879_55#_M1003_d VPB PSHORT L=0.15 W=1.12
+ AD=0.3864 AS=0.230629 PD=2.93 PS=1.72 NRD=10.5395 NRS=1.7533 M=1 R=7.46667
+ SA=75003 SB=75000.3 A=0.168 P=2.54 MULT=1
MM1018 N_A_811_379#_M1018_d N_A_879_55#_M1018_g N_A_1660_374#_M1018_s VPB PSHORT
+ L=0.15 W=0.84 AD=0.147 AS=0.2478 PD=1.19 PS=2.27 NRD=14.0658 NRS=2.3443 M=1
+ R=5.6 SA=75000.2 SB=75003.4 A=0.126 P=1.98 MULT=1
MM1019 N_A_1849_374#_M1019_d N_B_M1019_g N_A_811_379#_M1018_d VPB PSHORT L=0.15
+ W=0.84 AD=0.660675 AS=0.147 PD=2.395 PS=1.19 NRD=22.261 NRS=2.3443 M=1 R=5.6
+ SA=75000.7 SB=75002.9 A=0.126 P=1.98 MULT=1
MM1013 N_A_1023_379#_M1013_d N_A_879_55#_M1013_g N_A_1849_374#_M1019_d VPB
+ PSHORT L=0.15 W=0.84 AD=0.126 AS=0.660675 PD=1.14 PS=2.395 NRD=2.3443
+ NRS=75.0373 M=1 R=5.6 SA=75002.4 SB=75001.3 A=0.126 P=1.98 MULT=1
MM1016 N_A_1660_374#_M1016_d N_B_M1016_g N_A_1023_379#_M1013_d VPB PSHORT L=0.15
+ W=0.84 AD=0.1596 AS=0.126 PD=1.26429 PS=1.14 NRD=8.1952 NRS=2.3443 M=1 R=5.6
+ SA=75002.8 SB=75000.8 A=0.126 P=1.98 MULT=1
MM1007 N_VPWR_M1007_d N_A_2342_48#_M1007_g N_A_1660_374#_M1016_d VPB PSHORT
+ L=0.15 W=1.12 AD=0.4851 AS=0.2128 PD=3.31 PS=1.68571 NRD=17.8679 NRS=7.0329
+ M=1 R=7.46667 SA=75002.5 SB=75000.3 A=0.168 P=2.54 MULT=1
MM1009 N_VPWR_M1009_d N_A_M1009_g N_A_1849_374#_M1009_s VPB PSHORT L=0.15 W=1
+ AD=0.175 AS=0.295 PD=1.35 PS=2.59 NRD=1.9503 NRS=1.9503 M=1 R=6.66667
+ SA=75000.2 SB=75000.7 A=0.15 P=2.3 MULT=1
MM1008 N_A_2342_48#_M1008_d N_A_M1008_g N_VPWR_M1009_d VPB PSHORT L=0.15 W=1
+ AD=0.3 AS=0.175 PD=2.6 PS=1.35 NRD=1.9503 NRS=11.8003 M=1 R=6.66667 SA=75000.7
+ SB=75000.2 A=0.15 P=2.3 MULT=1
DX32_noxref VNB VPB NWDIODE A=26.8204 P=33.14
*
.include "sky130_fd_sc_hs__fah_1.pxi.spice"
*
.ends
*
*
