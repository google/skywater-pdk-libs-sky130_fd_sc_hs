* File: sky130_fd_sc_hs__fahcin_1.pxi.spice
* Created: Thu Aug 27 20:46:36 2020
* 
x_PM_SKY130_FD_SC_HS__FAHCIN_1%A N_A_M1017_g N_A_c_238_n N_A_M1005_g A
+ N_A_c_239_n PM_SKY130_FD_SC_HS__FAHCIN_1%A
x_PM_SKY130_FD_SC_HS__FAHCIN_1%A_28_74# N_A_28_74#_M1017_s N_A_28_74#_M1014_d
+ N_A_28_74#_M1005_s N_A_28_74#_M1021_d N_A_28_74#_c_267_n N_A_28_74#_M1000_g
+ N_A_28_74#_M1008_g N_A_28_74#_c_269_n N_A_28_74#_c_270_n N_A_28_74#_c_271_n
+ N_A_28_74#_c_272_n N_A_28_74#_c_279_n N_A_28_74#_c_273_n N_A_28_74#_c_280_n
+ N_A_28_74#_c_281_n N_A_28_74#_c_274_n N_A_28_74#_c_275_n N_A_28_74#_c_302_p
+ N_A_28_74#_c_282_n N_A_28_74#_c_276_n PM_SKY130_FD_SC_HS__FAHCIN_1%A_28_74#
x_PM_SKY130_FD_SC_HS__FAHCIN_1%A_492_48# N_A_492_48#_M1015_s N_A_492_48#_M1007_s
+ N_A_492_48#_M1014_g N_A_492_48#_c_388_n N_A_492_48#_c_389_n
+ N_A_492_48#_M1011_g N_A_492_48#_c_373_n N_A_492_48#_c_374_n
+ N_A_492_48#_M1021_g N_A_492_48#_M1025_g N_A_492_48#_c_376_n
+ N_A_492_48#_M1012_g N_A_492_48#_M1027_g N_A_492_48#_c_378_n
+ N_A_492_48#_c_379_n N_A_492_48#_c_380_n N_A_492_48#_c_381_n
+ N_A_492_48#_c_382_n N_A_492_48#_c_394_n N_A_492_48#_c_440_p
+ N_A_492_48#_c_383_n N_A_492_48#_c_384_n N_A_492_48#_c_385_n
+ N_A_492_48#_c_397_n N_A_492_48#_c_386_n N_A_492_48#_c_387_n
+ PM_SKY130_FD_SC_HS__FAHCIN_1%A_492_48#
x_PM_SKY130_FD_SC_HS__FAHCIN_1%B N_B_c_543_n N_B_M1006_g N_B_c_555_n N_B_M1029_g
+ N_B_c_544_n N_B_c_545_n N_B_c_556_n N_B_c_557_n N_B_c_558_n N_B_c_559_n
+ N_B_c_560_n N_B_M1016_g N_B_M1031_g N_B_c_547_n N_B_c_561_n N_B_c_548_n
+ N_B_c_549_n N_B_c_563_n N_B_M1007_g N_B_M1015_g N_B_c_564_n N_B_c_550_n
+ N_B_c_551_n N_B_c_552_n N_B_c_553_n B PM_SKY130_FD_SC_HS__FAHCIN_1%B
x_PM_SKY130_FD_SC_HS__FAHCIN_1%A_608_74# N_A_608_74#_M1006_d N_A_608_74#_M1029_d
+ N_A_608_74#_c_685_n N_A_608_74#_M1030_g N_A_608_74#_c_686_n
+ N_A_608_74#_M1023_g N_A_608_74#_M1018_g N_A_608_74#_c_688_n
+ N_A_608_74#_c_689_n N_A_608_74#_c_704_n N_A_608_74#_M1024_g
+ N_A_608_74#_c_690_n N_A_608_74#_c_705_n N_A_608_74#_c_691_n
+ N_A_608_74#_c_707_n N_A_608_74#_c_708_n N_A_608_74#_c_709_n
+ N_A_608_74#_c_710_n N_A_608_74#_c_741_n N_A_608_74#_c_742_n
+ N_A_608_74#_c_711_n N_A_608_74#_c_712_n N_A_608_74#_c_713_n
+ N_A_608_74#_c_714_n N_A_608_74#_c_715_n N_A_608_74#_c_692_n
+ N_A_608_74#_c_717_n N_A_608_74#_c_718_n N_A_608_74#_c_693_n
+ N_A_608_74#_c_694_n N_A_608_74#_c_695_n N_A_608_74#_c_696_n
+ N_A_608_74#_c_697_n N_A_608_74#_c_698_n N_A_608_74#_c_720_n
+ N_A_608_74#_c_801_p N_A_608_74#_c_699_n N_A_608_74#_c_700_n
+ N_A_608_74#_c_722_n N_A_608_74#_c_701_n PM_SKY130_FD_SC_HS__FAHCIN_1%A_608_74#
x_PM_SKY130_FD_SC_HS__FAHCIN_1%A_430_418# N_A_430_418#_M1014_s
+ N_A_430_418#_M1031_d N_A_430_418#_M1011_s N_A_430_418#_M1016_d
+ N_A_430_418#_c_950_n N_A_430_418#_M1002_g N_A_430_418#_c_951_n
+ N_A_430_418#_c_952_n N_A_430_418#_c_960_n N_A_430_418#_c_961_n
+ N_A_430_418#_c_962_n N_A_430_418#_M1026_g N_A_430_418#_c_953_n
+ N_A_430_418#_M1028_g N_A_430_418#_c_954_n N_A_430_418#_M1009_g
+ N_A_430_418#_c_955_n N_A_430_418#_c_956_n N_A_430_418#_c_966_n
+ N_A_430_418#_c_967_n N_A_430_418#_c_968_n N_A_430_418#_c_969_n
+ N_A_430_418#_c_970_n N_A_430_418#_c_971_n N_A_430_418#_c_972_n
+ N_A_430_418#_c_973_n N_A_430_418#_c_974_n N_A_430_418#_c_1077_p
+ N_A_430_418#_c_957_n N_A_430_418#_c_958_n N_A_430_418#_c_959_n
+ PM_SKY130_FD_SC_HS__FAHCIN_1%A_430_418#
x_PM_SKY130_FD_SC_HS__FAHCIN_1%CIN N_CIN_c_1167_n N_CIN_M1004_g N_CIN_c_1163_n
+ N_CIN_M1019_g N_CIN_c_1168_n N_CIN_M1010_g N_CIN_c_1164_n N_CIN_M1003_g CIN
+ N_CIN_c_1166_n PM_SKY130_FD_SC_HS__FAHCIN_1%CIN
x_PM_SKY130_FD_SC_HS__FAHCIN_1%A_1854_368# N_A_1854_368#_M1003_d
+ N_A_1854_368#_M1010_d N_A_1854_368#_M1028_d N_A_1854_368#_c_1222_n
+ N_A_1854_368#_M1001_g N_A_1854_368#_c_1227_n N_A_1854_368#_M1013_g
+ N_A_1854_368#_c_1228_n N_A_1854_368#_c_1239_n N_A_1854_368#_c_1229_n
+ N_A_1854_368#_c_1230_n N_A_1854_368#_c_1231_n N_A_1854_368#_c_1232_n
+ N_A_1854_368#_c_1223_n N_A_1854_368#_c_1224_n N_A_1854_368#_c_1234_n
+ N_A_1854_368#_c_1235_n N_A_1854_368#_c_1225_n N_A_1854_368#_c_1226_n
+ PM_SKY130_FD_SC_HS__FAHCIN_1%A_1854_368#
x_PM_SKY130_FD_SC_HS__FAHCIN_1%A_2004_136# N_A_2004_136#_M1018_d
+ N_A_2004_136#_M1024_d N_A_2004_136#_c_1317_n N_A_2004_136#_M1022_g
+ N_A_2004_136#_c_1318_n N_A_2004_136#_M1020_g N_A_2004_136#_c_1319_n
+ N_A_2004_136#_c_1320_n N_A_2004_136#_c_1321_n N_A_2004_136#_c_1322_n
+ N_A_2004_136#_c_1323_n N_A_2004_136#_c_1360_n N_A_2004_136#_c_1362_n
+ N_A_2004_136#_c_1324_n N_A_2004_136#_c_1336_n
+ PM_SKY130_FD_SC_HS__FAHCIN_1%A_2004_136#
x_PM_SKY130_FD_SC_HS__FAHCIN_1%VPWR N_VPWR_M1005_d N_VPWR_M1007_d N_VPWR_M1004_d
+ N_VPWR_M1013_d N_VPWR_c_1401_n N_VPWR_c_1402_n N_VPWR_c_1403_n N_VPWR_c_1404_n
+ N_VPWR_c_1405_n N_VPWR_c_1406_n VPWR N_VPWR_c_1407_n N_VPWR_c_1408_n
+ N_VPWR_c_1409_n N_VPWR_c_1410_n N_VPWR_c_1400_n N_VPWR_c_1412_n
+ N_VPWR_c_1413_n N_VPWR_c_1414_n PM_SKY130_FD_SC_HS__FAHCIN_1%VPWR
x_PM_SKY130_FD_SC_HS__FAHCIN_1%A_256_368# N_A_256_368#_M1008_d
+ N_A_256_368#_M1025_d N_A_256_368#_M1000_d N_A_256_368#_M1011_d
+ N_A_256_368#_c_1505_n N_A_256_368#_c_1506_n N_A_256_368#_c_1507_n
+ N_A_256_368#_c_1508_n N_A_256_368#_c_1516_n N_A_256_368#_c_1550_n
+ N_A_256_368#_c_1534_n N_A_256_368#_c_1499_n N_A_256_368#_c_1517_n
+ N_A_256_368#_c_1500_n N_A_256_368#_c_1509_n N_A_256_368#_c_1501_n
+ N_A_256_368#_c_1502_n N_A_256_368#_c_1503_n N_A_256_368#_c_1504_n
+ PM_SKY130_FD_SC_HS__FAHCIN_1%A_256_368#
x_PM_SKY130_FD_SC_HS__FAHCIN_1%A_1197_368# N_A_1197_368#_M1027_d
+ N_A_1197_368#_M1012_d N_A_1197_368#_c_1593_n N_A_1197_368#_c_1596_n
+ N_A_1197_368#_c_1594_n N_A_1197_368#_c_1595_n
+ PM_SKY130_FD_SC_HS__FAHCIN_1%A_1197_368#
x_PM_SKY130_FD_SC_HS__FAHCIN_1%COUT N_COUT_M1002_d N_COUT_M1030_d
+ N_COUT_c_1630_n N_COUT_c_1643_n N_COUT_c_1631_n COUT COUT
+ PM_SKY130_FD_SC_HS__FAHCIN_1%COUT
x_PM_SKY130_FD_SC_HS__FAHCIN_1%A_1595_400# N_A_1595_400#_M1023_d
+ N_A_1595_400#_M1026_d N_A_1595_400#_c_1680_n N_A_1595_400#_c_1685_n
+ N_A_1595_400#_c_1677_n N_A_1595_400#_c_1678_n N_A_1595_400#_c_1679_n
+ PM_SKY130_FD_SC_HS__FAHCIN_1%A_1595_400#
x_PM_SKY130_FD_SC_HS__FAHCIN_1%A_1967_384# N_A_1967_384#_M1009_d
+ N_A_1967_384#_M1024_s N_A_1967_384#_M1013_s N_A_1967_384#_c_1729_n
+ N_A_1967_384#_c_1708_n N_A_1967_384#_c_1709_n N_A_1967_384#_c_1706_n
+ N_A_1967_384#_c_1723_n N_A_1967_384#_c_1710_n N_A_1967_384#_c_1711_n
+ N_A_1967_384#_c_1707_n PM_SKY130_FD_SC_HS__FAHCIN_1%A_1967_384#
x_PM_SKY130_FD_SC_HS__FAHCIN_1%SUM N_SUM_M1020_d N_SUM_M1022_d SUM SUM SUM SUM
+ SUM SUM SUM PM_SKY130_FD_SC_HS__FAHCIN_1%SUM
x_PM_SKY130_FD_SC_HS__FAHCIN_1%VGND N_VGND_M1017_d N_VGND_M1015_d N_VGND_M1019_d
+ N_VGND_M1001_d N_VGND_c_1770_n N_VGND_c_1771_n N_VGND_c_1772_n N_VGND_c_1773_n
+ VGND N_VGND_c_1774_n N_VGND_c_1775_n N_VGND_c_1776_n N_VGND_c_1777_n
+ N_VGND_c_1778_n N_VGND_c_1779_n N_VGND_c_1780_n N_VGND_c_1781_n
+ N_VGND_c_1782_n N_VGND_c_1783_n PM_SKY130_FD_SC_HS__FAHCIN_1%VGND
cc_1 VNB N_A_M1017_g 0.0315064f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=0.74
cc_2 VNB N_A_c_238_n 0.0361271f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=1.765
cc_3 VNB N_A_c_239_n 0.00241315f $X=-0.19 $Y=-0.245 $X2=0.71 $Y2=1.515
cc_4 VNB N_A_28_74#_c_267_n 0.0384485f $X=-0.19 $Y=-0.245 $X2=0.69 $Y2=1.515
cc_5 VNB N_A_28_74#_M1008_g 0.0254313f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_6 VNB N_A_28_74#_c_269_n 0.0277086f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_7 VNB N_A_28_74#_c_270_n 0.0240482f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_A_28_74#_c_271_n 0.00680342f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A_28_74#_c_272_n 0.00941963f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_28_74#_c_273_n 7.67056e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_28_74#_c_274_n 0.0309085f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_28_74#_c_275_n 0.00272939f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_28_74#_c_276_n 0.00935765f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_492_48#_M1014_g 0.034419f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_492_48#_c_373_n 0.0489586f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_492_48#_c_374_n 0.0307165f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_492_48#_M1025_g 0.0197088f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_492_48#_c_376_n 0.0531561f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_492_48#_M1027_g 0.0237855f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_492_48#_c_378_n 0.0123274f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_492_48#_c_379_n 0.00290227f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_492_48#_c_380_n 0.0143458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_492_48#_c_381_n 0.00159323f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_492_48#_c_382_n 0.00370531f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_492_48#_c_383_n 0.00146225f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_492_48#_c_384_n 0.00126249f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_492_48#_c_385_n 0.0140893f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_492_48#_c_386_n 0.00588023f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_492_48#_c_387_n 0.00271717f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_B_c_543_n 0.0160994f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=1.35
cc_31 VNB N_B_c_544_n 0.0861447f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=2.4
cc_32 VNB N_B_c_545_n 0.0123527f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_33 VNB N_B_M1031_g 0.0312285f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_B_c_547_n 0.0356568f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_B_c_548_n 0.00426041f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_B_c_549_n 0.0559851f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_B_c_550_n 0.00749069f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_B_c_551_n 0.0139891f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_B_c_552_n 0.0442797f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_B_c_553_n 0.018754f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB B 0.00807683f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_608_74#_c_685_n 0.0180887f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=2.4
cc_43 VNB N_A_608_74#_c_686_n 0.0234224f $X=-0.19 $Y=-0.245 $X2=0.65 $Y2=1.515
cc_44 VNB N_A_608_74#_M1018_g 0.00764536f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_A_608_74#_c_688_n 0.0278016f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_A_608_74#_c_689_n 0.00667824f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_608_74#_c_690_n 0.0184598f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_608_74#_c_691_n 0.00411066f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A_608_74#_c_692_n 0.00257604f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_A_608_74#_c_693_n 0.00423629f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_A_608_74#_c_694_n 0.00411475f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_A_608_74#_c_695_n 0.00202646f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_A_608_74#_c_696_n 0.00373666f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_A_608_74#_c_697_n 0.0121753f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_A_608_74#_c_698_n 0.0622779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_A_608_74#_c_699_n 0.00249927f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_A_608_74#_c_700_n 0.00357135f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_A_608_74#_c_701_n 0.0423682f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_A_430_418#_c_950_n 0.0185368f $X=-0.19 $Y=-0.245 $X2=0.69 $Y2=1.515
cc_60 VNB N_A_430_418#_c_951_n 0.0601382f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_A_430_418#_c_952_n 0.00809181f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_A_430_418#_c_953_n 0.0288231f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_A_430_418#_c_954_n 0.0196479f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_A_430_418#_c_955_n 0.0220679f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_A_430_418#_c_956_n 0.0143866f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_A_430_418#_c_957_n 0.0301313f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_A_430_418#_c_958_n 0.00399338f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_A_430_418#_c_959_n 0.00322214f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_CIN_c_1163_n 0.0186178f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_CIN_c_1164_n 0.0161662f $X=-0.19 $Y=-0.245 $X2=0.65 $Y2=1.515
cc_71 VNB CIN 0.00303624f $X=-0.19 $Y=-0.245 $X2=0.69 $Y2=1.515
cc_72 VNB N_CIN_c_1166_n 0.104245f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_A_1854_368#_c_1222_n 0.0202294f $X=-0.19 $Y=-0.245 $X2=0.65
+ $Y2=1.515
cc_74 VNB N_A_1854_368#_c_1223_n 0.00659559f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_A_1854_368#_c_1224_n 0.0060187f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_A_1854_368#_c_1225_n 0.0359566f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_A_1854_368#_c_1226_n 0.00288542f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_A_2004_136#_c_1317_n 0.0347631f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=2.4
cc_79 VNB N_A_2004_136#_c_1318_n 0.021195f $X=-0.19 $Y=-0.245 $X2=0.65 $Y2=1.515
cc_80 VNB N_A_2004_136#_c_1319_n 0.00405023f $X=-0.19 $Y=-0.245 $X2=0.69
+ $Y2=1.665
cc_81 VNB N_A_2004_136#_c_1320_n 0.00491697f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_82 VNB N_A_2004_136#_c_1321_n 0.0182706f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_83 VNB N_A_2004_136#_c_1322_n 0.00269518f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_84 VNB N_A_2004_136#_c_1323_n 0.00189369f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_85 VNB N_A_2004_136#_c_1324_n 0.00164386f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_86 VNB N_VPWR_c_1400_n 0.541827f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_87 VNB N_A_256_368#_c_1499_n 0.0123292f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_88 VNB N_A_256_368#_c_1500_n 0.00176057f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_89 VNB N_A_256_368#_c_1501_n 0.0143257f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_90 VNB N_A_256_368#_c_1502_n 0.00563003f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_91 VNB N_A_256_368#_c_1503_n 0.00496161f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_92 VNB N_A_256_368#_c_1504_n 0.00278665f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_93 VNB N_A_1197_368#_c_1593_n 0.00254826f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_94 VNB N_A_1197_368#_c_1594_n 0.00657764f $X=-0.19 $Y=-0.245 $X2=0.69
+ $Y2=1.665
cc_95 VNB N_A_1197_368#_c_1595_n 0.0044471f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_96 VNB N_COUT_c_1630_n 0.00726691f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_97 VNB N_COUT_c_1631_n 0.0103544f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_98 VNB N_A_1595_400#_c_1677_n 0.00303844f $X=-0.19 $Y=-0.245 $X2=0.69
+ $Y2=1.515
cc_99 VNB N_A_1595_400#_c_1678_n 0.0121901f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_100 VNB N_A_1595_400#_c_1679_n 0.00248754f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_101 VNB N_A_1967_384#_c_1706_n 2.80212e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_102 VNB N_A_1967_384#_c_1707_n 0.00677145f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_103 VNB SUM 0.0184457f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=2.4
cc_104 VNB SUM 0.03594f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_105 VNB N_VGND_c_1770_n 0.0107331f $X=-0.19 $Y=-0.245 $X2=0.69 $Y2=1.665
cc_106 VNB N_VGND_c_1771_n 0.0133606f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_107 VNB N_VGND_c_1772_n 0.0135101f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_108 VNB N_VGND_c_1773_n 0.0207581f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_109 VNB N_VGND_c_1774_n 0.0193106f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_110 VNB N_VGND_c_1775_n 0.106993f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_111 VNB N_VGND_c_1776_n 0.0730655f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_112 VNB N_VGND_c_1777_n 0.0695222f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_113 VNB N_VGND_c_1778_n 0.0195666f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_114 VNB N_VGND_c_1779_n 0.692691f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_115 VNB N_VGND_c_1780_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_116 VNB N_VGND_c_1781_n 0.00969062f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_117 VNB N_VGND_c_1782_n 0.00653982f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_118 VNB N_VGND_c_1783_n 0.0080786f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_119 VPB N_A_c_238_n 0.0377974f $X=-0.19 $Y=1.66 $X2=0.515 $Y2=1.765
cc_120 VPB N_A_c_239_n 0.00320363f $X=-0.19 $Y=1.66 $X2=0.71 $Y2=1.515
cc_121 VPB N_A_28_74#_c_267_n 0.0262877f $X=-0.19 $Y=1.66 $X2=0.69 $Y2=1.515
cc_122 VPB N_A_28_74#_c_270_n 0.0539701f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_123 VPB N_A_28_74#_c_279_n 0.00184963f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_124 VPB N_A_28_74#_c_280_n 0.0381768f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_125 VPB N_A_28_74#_c_281_n 0.00244277f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_126 VPB N_A_28_74#_c_282_n 0.00435773f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_127 VPB N_A_492_48#_c_388_n 0.0162835f $X=-0.19 $Y=1.66 $X2=0.71 $Y2=1.515
cc_128 VPB N_A_492_48#_c_389_n 0.0237245f $X=-0.19 $Y=1.66 $X2=0.69 $Y2=1.515
cc_129 VPB N_A_492_48#_c_373_n 0.023017f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_130 VPB N_A_492_48#_c_374_n 0.0410689f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_131 VPB N_A_492_48#_c_376_n 0.0245512f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_132 VPB N_A_492_48#_c_378_n 2.20132e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_133 VPB N_A_492_48#_c_394_n 0.00704552f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_134 VPB N_A_492_48#_c_384_n 0.00303878f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_135 VPB N_A_492_48#_c_385_n 0.0030902f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_136 VPB N_A_492_48#_c_397_n 0.0052784f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_137 VPB N_B_c_555_n 0.0137521f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_138 VPB N_B_c_556_n 0.08191f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_139 VPB N_B_c_557_n 0.0197011f $X=-0.19 $Y=1.66 $X2=0.65 $Y2=1.515
cc_140 VPB N_B_c_558_n 0.00698484f $X=-0.19 $Y=1.66 $X2=0.71 $Y2=1.515
cc_141 VPB N_B_c_559_n 0.0109377f $X=-0.19 $Y=1.66 $X2=0.71 $Y2=1.515
cc_142 VPB N_B_c_560_n 0.0160072f $X=-0.19 $Y=1.66 $X2=0.69 $Y2=1.515
cc_143 VPB N_B_c_561_n 0.0347272f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_144 VPB N_B_c_548_n 0.0767623f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_145 VPB N_B_c_563_n 0.0175183f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_146 VPB N_B_c_564_n 0.0089864f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_147 VPB N_B_c_552_n 0.00726359f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_148 VPB N_A_608_74#_c_685_n 0.0451694f $X=-0.19 $Y=1.66 $X2=0.515 $Y2=2.4
cc_149 VPB N_A_608_74#_c_689_n 0.00550662f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_150 VPB N_A_608_74#_c_704_n 0.0220558f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_151 VPB N_A_608_74#_c_705_n 5.58911e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_152 VPB N_A_608_74#_c_691_n 0.00260521f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_153 VPB N_A_608_74#_c_707_n 0.00489305f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_154 VPB N_A_608_74#_c_708_n 0.00126888f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_155 VPB N_A_608_74#_c_709_n 0.0104049f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_156 VPB N_A_608_74#_c_710_n 0.00159323f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_157 VPB N_A_608_74#_c_711_n 9.80449e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_158 VPB N_A_608_74#_c_712_n 0.00324116f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_159 VPB N_A_608_74#_c_713_n 0.00140424f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_160 VPB N_A_608_74#_c_714_n 0.033504f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_161 VPB N_A_608_74#_c_715_n 0.00611548f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_162 VPB N_A_608_74#_c_692_n 0.00411346f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_163 VPB N_A_608_74#_c_717_n 0.0159757f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_164 VPB N_A_608_74#_c_718_n 6.01039e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_165 VPB N_A_608_74#_c_693_n 0.00714486f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_166 VPB N_A_608_74#_c_720_n 0.00312651f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_167 VPB N_A_608_74#_c_699_n 9.06608e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_168 VPB N_A_608_74#_c_722_n 0.00122299f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_169 VPB N_A_430_418#_c_960_n 0.0366731f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_170 VPB N_A_430_418#_c_961_n 0.0187079f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_171 VPB N_A_430_418#_c_962_n 0.017637f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_172 VPB N_A_430_418#_c_953_n 0.0396387f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_173 VPB N_A_430_418#_c_955_n 0.00663468f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_174 VPB N_A_430_418#_c_956_n 0.0073459f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_175 VPB N_A_430_418#_c_966_n 0.00150798f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_176 VPB N_A_430_418#_c_967_n 0.00506007f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_177 VPB N_A_430_418#_c_968_n 0.0031884f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_178 VPB N_A_430_418#_c_969_n 0.0187719f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_179 VPB N_A_430_418#_c_970_n 7.2724e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_180 VPB N_A_430_418#_c_971_n 0.0115552f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_181 VPB N_A_430_418#_c_972_n 7.90628e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_182 VPB N_A_430_418#_c_973_n 0.0144569f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_183 VPB N_A_430_418#_c_974_n 0.00705926f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_184 VPB N_A_430_418#_c_957_n 0.00563137f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_185 VPB N_A_430_418#_c_958_n 0.00216373f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_186 VPB N_A_430_418#_c_959_n 0.00127727f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_187 VPB N_CIN_c_1167_n 0.0163015f $X=-0.19 $Y=1.66 $X2=0.5 $Y2=1.35
cc_188 VPB N_CIN_c_1168_n 0.0188223f $X=-0.19 $Y=1.66 $X2=0.515 $Y2=2.4
cc_189 VPB N_CIN_c_1166_n 0.0155732f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_190 VPB N_A_1854_368#_c_1227_n 0.0172624f $X=-0.19 $Y=1.66 $X2=0.69 $Y2=1.515
cc_191 VPB N_A_1854_368#_c_1228_n 0.0100535f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_192 VPB N_A_1854_368#_c_1229_n 0.00480016f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_193 VPB N_A_1854_368#_c_1230_n 0.0165534f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_194 VPB N_A_1854_368#_c_1231_n 0.00250967f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_195 VPB N_A_1854_368#_c_1232_n 0.00262687f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_196 VPB N_A_1854_368#_c_1223_n 0.00624422f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_197 VPB N_A_1854_368#_c_1234_n 0.0290493f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_198 VPB N_A_1854_368#_c_1235_n 0.00717098f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_199 VPB N_A_1854_368#_c_1225_n 0.0175713f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_200 VPB N_A_1854_368#_c_1226_n 4.25781e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_201 VPB N_A_2004_136#_c_1317_n 0.0371534f $X=-0.19 $Y=1.66 $X2=0.515 $Y2=2.4
cc_202 VPB N_A_2004_136#_c_1319_n 0.00181304f $X=-0.19 $Y=1.66 $X2=0.69
+ $Y2=1.665
cc_203 VPB N_A_2004_136#_c_1324_n 0.00205193f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_204 VPB N_VPWR_c_1401_n 0.00600159f $X=-0.19 $Y=1.66 $X2=0.69 $Y2=1.665
cc_205 VPB N_VPWR_c_1402_n 0.00859185f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_206 VPB N_VPWR_c_1403_n 0.00799841f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_207 VPB N_VPWR_c_1404_n 0.00598112f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_208 VPB N_VPWR_c_1405_n 0.0751118f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_209 VPB N_VPWR_c_1406_n 0.00324402f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_210 VPB N_VPWR_c_1407_n 0.0183065f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_211 VPB N_VPWR_c_1408_n 0.108695f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_212 VPB N_VPWR_c_1409_n 0.072584f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_213 VPB N_VPWR_c_1410_n 0.0180274f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_214 VPB N_VPWR_c_1400_n 0.150461f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_215 VPB N_VPWR_c_1412_n 0.00460249f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_216 VPB N_VPWR_c_1413_n 0.00671858f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_217 VPB N_VPWR_c_1414_n 0.00460249f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_218 VPB N_A_256_368#_c_1505_n 0.0101262f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_219 VPB N_A_256_368#_c_1506_n 0.0119515f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_220 VPB N_A_256_368#_c_1507_n 0.00378114f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_221 VPB N_A_256_368#_c_1508_n 0.00237322f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_222 VPB N_A_256_368#_c_1509_n 0.0109216f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_223 VPB N_A_256_368#_c_1501_n 0.0042336f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_224 VPB N_A_256_368#_c_1503_n 0.00555687f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_225 VPB N_A_1197_368#_c_1596_n 0.00292153f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_226 VPB N_A_1197_368#_c_1594_n 0.0023976f $X=-0.19 $Y=1.66 $X2=0.69 $Y2=1.665
cc_227 VPB N_COUT_c_1630_n 0.0062147f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_228 VPB N_A_1595_400#_c_1680_n 0.00267638f $X=-0.19 $Y=1.66 $X2=0.515 $Y2=2.4
cc_229 VPB N_A_1595_400#_c_1678_n 0.00307434f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_230 VPB N_A_1967_384#_c_1708_n 0.00262968f $X=-0.19 $Y=1.66 $X2=0.71
+ $Y2=1.515
cc_231 VPB N_A_1967_384#_c_1709_n 0.00925292f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_232 VPB N_A_1967_384#_c_1710_n 0.00649699f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_233 VPB N_A_1967_384#_c_1711_n 0.00360845f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_234 VPB N_A_1967_384#_c_1707_n 0.00399265f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_235 VPB SUM 0.0539684f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_236 N_A_M1017_g N_A_28_74#_c_267_n 8.11251e-19 $X=0.5 $Y=0.74 $X2=0 $Y2=0
cc_237 N_A_c_238_n N_A_28_74#_c_267_n 0.0305981f $X=0.515 $Y=1.765 $X2=0 $Y2=0
cc_238 N_A_c_239_n N_A_28_74#_c_267_n 6.29033e-19 $X=0.71 $Y=1.515 $X2=0 $Y2=0
cc_239 N_A_M1017_g N_A_28_74#_c_269_n 0.0108351f $X=0.5 $Y=0.74 $X2=0 $Y2=0
cc_240 N_A_M1017_g N_A_28_74#_c_270_n 0.0159847f $X=0.5 $Y=0.74 $X2=0 $Y2=0
cc_241 N_A_c_238_n N_A_28_74#_c_270_n 0.00788328f $X=0.515 $Y=1.765 $X2=0 $Y2=0
cc_242 N_A_c_239_n N_A_28_74#_c_270_n 0.0329871f $X=0.71 $Y=1.515 $X2=0 $Y2=0
cc_243 N_A_M1017_g N_A_28_74#_c_271_n 0.0160518f $X=0.5 $Y=0.74 $X2=0 $Y2=0
cc_244 N_A_c_238_n N_A_28_74#_c_271_n 0.0033642f $X=0.515 $Y=1.765 $X2=0 $Y2=0
cc_245 N_A_c_239_n N_A_28_74#_c_271_n 0.02209f $X=0.71 $Y=1.515 $X2=0 $Y2=0
cc_246 N_A_M1017_g N_A_28_74#_c_272_n 0.00257623f $X=0.5 $Y=0.74 $X2=0 $Y2=0
cc_247 N_A_c_238_n N_A_28_74#_c_272_n 0.00196095f $X=0.515 $Y=1.765 $X2=0 $Y2=0
cc_248 N_A_c_239_n N_A_28_74#_c_272_n 0.0225779f $X=0.71 $Y=1.515 $X2=0 $Y2=0
cc_249 N_A_c_238_n N_A_28_74#_c_279_n 0.00181871f $X=0.515 $Y=1.765 $X2=0 $Y2=0
cc_250 N_A_c_239_n N_A_28_74#_c_279_n 0.0115302f $X=0.71 $Y=1.515 $X2=0 $Y2=0
cc_251 N_A_M1017_g N_A_28_74#_c_273_n 0.00303494f $X=0.5 $Y=0.74 $X2=0 $Y2=0
cc_252 N_A_c_238_n N_A_28_74#_c_281_n 6.38314e-19 $X=0.515 $Y=1.765 $X2=0 $Y2=0
cc_253 N_A_M1017_g N_A_28_74#_c_276_n 0.00304554f $X=0.5 $Y=0.74 $X2=0 $Y2=0
cc_254 N_A_c_238_n N_VPWR_c_1401_n 0.0196325f $X=0.515 $Y=1.765 $X2=0 $Y2=0
cc_255 N_A_c_239_n N_VPWR_c_1401_n 0.0193147f $X=0.71 $Y=1.515 $X2=0 $Y2=0
cc_256 N_A_c_238_n N_VPWR_c_1407_n 0.00413917f $X=0.515 $Y=1.765 $X2=0 $Y2=0
cc_257 N_A_c_238_n N_VPWR_c_1400_n 0.00821254f $X=0.515 $Y=1.765 $X2=0 $Y2=0
cc_258 N_A_M1017_g N_VGND_c_1770_n 0.0141934f $X=0.5 $Y=0.74 $X2=0 $Y2=0
cc_259 N_A_M1017_g N_VGND_c_1774_n 0.00434272f $X=0.5 $Y=0.74 $X2=0 $Y2=0
cc_260 N_A_M1017_g N_VGND_c_1779_n 0.00828734f $X=0.5 $Y=0.74 $X2=0 $Y2=0
cc_261 N_A_28_74#_c_274_n N_A_492_48#_M1014_g 0.0136594f $X=2.585 $Y=0.34 $X2=0
+ $Y2=0
cc_262 N_A_28_74#_c_302_p N_A_492_48#_M1014_g 0.0106281f $X=2.75 $Y=0.55 $X2=0
+ $Y2=0
cc_263 N_A_28_74#_c_280_n N_A_492_48#_c_389_n 0.0121257f $X=3.685 $Y=2.99 $X2=0
+ $Y2=0
cc_264 N_A_28_74#_c_302_p N_A_492_48#_c_373_n 0.0028692f $X=2.75 $Y=0.55 $X2=0
+ $Y2=0
cc_265 N_A_28_74#_c_280_n N_A_492_48#_c_374_n 0.00347797f $X=3.685 $Y=2.99 $X2=0
+ $Y2=0
cc_266 N_A_28_74#_c_282_n N_A_492_48#_c_374_n 0.00764912f $X=3.85 $Y=2.43 $X2=0
+ $Y2=0
cc_267 N_A_28_74#_c_274_n N_B_c_543_n 9.18426e-19 $X=2.585 $Y=0.34 $X2=-0.19
+ $Y2=-0.245
cc_268 N_A_28_74#_c_280_n N_B_c_555_n 0.0112424f $X=3.685 $Y=2.99 $X2=0 $Y2=0
cc_269 N_A_28_74#_c_282_n N_B_c_555_n 0.00121631f $X=3.85 $Y=2.43 $X2=0 $Y2=0
cc_270 N_A_28_74#_c_280_n N_B_c_556_n 0.0166861f $X=3.685 $Y=2.99 $X2=0 $Y2=0
cc_271 N_A_28_74#_c_280_n N_B_c_557_n 0.00594174f $X=3.685 $Y=2.99 $X2=0 $Y2=0
cc_272 N_A_28_74#_c_282_n N_B_c_558_n 4.13106e-19 $X=3.85 $Y=2.43 $X2=0 $Y2=0
cc_273 N_A_28_74#_c_280_n N_B_c_559_n 0.00106333f $X=3.685 $Y=2.99 $X2=0 $Y2=0
cc_274 N_A_28_74#_c_282_n N_B_c_560_n 0.00175517f $X=3.85 $Y=2.43 $X2=0 $Y2=0
cc_275 N_A_28_74#_c_280_n N_A_608_74#_M1029_d 0.00266003f $X=3.685 $Y=2.99 $X2=0
+ $Y2=0
cc_276 N_A_28_74#_c_280_n N_A_608_74#_c_705_n 0.0228124f $X=3.685 $Y=2.99 $X2=0
+ $Y2=0
cc_277 N_A_28_74#_M1021_d N_A_608_74#_c_707_n 0.00589973f $X=3.65 $Y=1.895 $X2=0
+ $Y2=0
cc_278 N_A_28_74#_c_282_n N_A_608_74#_c_707_n 0.0137222f $X=3.85 $Y=2.43 $X2=0
+ $Y2=0
cc_279 N_A_28_74#_M1021_d N_A_608_74#_c_708_n 0.00738292f $X=3.65 $Y=1.895 $X2=0
+ $Y2=0
cc_280 N_A_28_74#_c_282_n N_A_608_74#_c_708_n 0.0493824f $X=3.85 $Y=2.43 $X2=0
+ $Y2=0
cc_281 N_A_28_74#_c_280_n N_A_608_74#_c_710_n 0.015927f $X=3.685 $Y=2.99 $X2=0
+ $Y2=0
cc_282 N_A_28_74#_c_274_n N_A_430_418#_M1014_s 0.00257204f $X=2.585 $Y=0.34
+ $X2=-0.19 $Y2=-0.245
cc_283 N_A_28_74#_c_280_n N_A_430_418#_M1011_s 0.00304846f $X=3.685 $Y=2.99
+ $X2=0 $Y2=0
cc_284 N_A_28_74#_M1008_g N_A_430_418#_c_955_n 0.00185792f $X=1.41 $Y=0.79 $X2=0
+ $Y2=0
cc_285 N_A_28_74#_c_274_n N_A_430_418#_c_955_n 0.016478f $X=2.585 $Y=0.34 $X2=0
+ $Y2=0
cc_286 N_A_28_74#_M1021_d N_A_430_418#_c_967_n 0.00981922f $X=3.65 $Y=1.895
+ $X2=0 $Y2=0
cc_287 N_A_28_74#_c_282_n N_A_430_418#_c_967_n 0.006835f $X=3.85 $Y=2.43 $X2=0
+ $Y2=0
cc_288 N_A_28_74#_c_279_n N_VPWR_M1005_d 0.0100571f $X=1.09 $Y=2.905 $X2=-0.19
+ $Y2=-0.245
cc_289 N_A_28_74#_c_267_n N_VPWR_c_1401_n 0.00308226f $X=1.205 $Y=1.765 $X2=0
+ $Y2=0
cc_290 N_A_28_74#_c_270_n N_VPWR_c_1401_n 0.067783f $X=0.29 $Y=1.985 $X2=0 $Y2=0
cc_291 N_A_28_74#_c_279_n N_VPWR_c_1401_n 0.068507f $X=1.09 $Y=2.905 $X2=0 $Y2=0
cc_292 N_A_28_74#_c_281_n N_VPWR_c_1401_n 0.0140789f $X=1.175 $Y=2.99 $X2=0
+ $Y2=0
cc_293 N_A_28_74#_c_270_n N_VPWR_c_1407_n 0.0112891f $X=0.29 $Y=1.985 $X2=0
+ $Y2=0
cc_294 N_A_28_74#_c_267_n N_VPWR_c_1408_n 7.43987e-19 $X=1.205 $Y=1.765 $X2=0
+ $Y2=0
cc_295 N_A_28_74#_c_280_n N_VPWR_c_1408_n 0.178139f $X=3.685 $Y=2.99 $X2=0 $Y2=0
cc_296 N_A_28_74#_c_281_n N_VPWR_c_1408_n 0.0121505f $X=1.175 $Y=2.99 $X2=0
+ $Y2=0
cc_297 N_A_28_74#_c_270_n N_VPWR_c_1400_n 0.00934413f $X=0.29 $Y=1.985 $X2=0
+ $Y2=0
cc_298 N_A_28_74#_c_280_n N_VPWR_c_1400_n 0.0998778f $X=3.685 $Y=2.99 $X2=0
+ $Y2=0
cc_299 N_A_28_74#_c_281_n N_VPWR_c_1400_n 0.00660392f $X=1.175 $Y=2.99 $X2=0
+ $Y2=0
cc_300 N_A_28_74#_c_280_n N_A_256_368#_M1011_d 0.00240242f $X=3.685 $Y=2.99
+ $X2=0 $Y2=0
cc_301 N_A_28_74#_c_280_n N_A_256_368#_c_1506_n 0.0501424f $X=3.685 $Y=2.99
+ $X2=0 $Y2=0
cc_302 N_A_28_74#_c_279_n N_A_256_368#_c_1507_n 0.013418f $X=1.09 $Y=2.905 $X2=0
+ $Y2=0
cc_303 N_A_28_74#_c_280_n N_A_256_368#_c_1507_n 0.0382734f $X=3.685 $Y=2.99
+ $X2=0 $Y2=0
cc_304 N_A_28_74#_c_280_n N_A_256_368#_c_1516_n 0.0182069f $X=3.685 $Y=2.99
+ $X2=0 $Y2=0
cc_305 N_A_28_74#_c_274_n N_A_256_368#_c_1517_n 0.0124901f $X=2.585 $Y=0.34
+ $X2=0 $Y2=0
cc_306 N_A_28_74#_c_267_n N_A_256_368#_c_1509_n 0.00930908f $X=1.205 $Y=1.765
+ $X2=0 $Y2=0
cc_307 N_A_28_74#_c_272_n N_A_256_368#_c_1509_n 0.00771297f $X=1.09 $Y=1.63
+ $X2=0 $Y2=0
cc_308 N_A_28_74#_c_279_n N_A_256_368#_c_1509_n 0.0568852f $X=1.09 $Y=2.905
+ $X2=0 $Y2=0
cc_309 N_A_28_74#_c_267_n N_A_256_368#_c_1501_n 0.00356111f $X=1.205 $Y=1.765
+ $X2=0 $Y2=0
cc_310 N_A_28_74#_M1008_g N_A_256_368#_c_1501_n 0.0141665f $X=1.41 $Y=0.79 $X2=0
+ $Y2=0
cc_311 N_A_28_74#_c_272_n N_A_256_368#_c_1501_n 0.0380023f $X=1.09 $Y=1.63 $X2=0
+ $Y2=0
cc_312 N_A_28_74#_c_279_n N_A_256_368#_c_1501_n 0.00677897f $X=1.09 $Y=2.905
+ $X2=0 $Y2=0
cc_313 N_A_28_74#_M1008_g N_A_256_368#_c_1502_n 0.00485468f $X=1.41 $Y=0.79
+ $X2=0 $Y2=0
cc_314 N_A_28_74#_c_274_n N_A_256_368#_c_1502_n 0.0224951f $X=2.585 $Y=0.34
+ $X2=0 $Y2=0
cc_315 N_A_28_74#_M1014_d N_A_256_368#_c_1504_n 0.00134007f $X=2.61 $Y=0.37
+ $X2=0 $Y2=0
cc_316 N_A_28_74#_c_302_p N_A_256_368#_c_1504_n 0.00182376f $X=2.75 $Y=0.55
+ $X2=0 $Y2=0
cc_317 N_A_28_74#_c_271_n N_VGND_M1017_d 0.00683277f $X=1.005 $Y=1.095 $X2=-0.19
+ $Y2=-0.245
cc_318 N_A_28_74#_c_272_n N_VGND_M1017_d 0.00669877f $X=1.09 $Y=1.63 $X2=-0.19
+ $Y2=-0.245
cc_319 N_A_28_74#_c_273_n N_VGND_M1017_d 0.0101547f $X=1.205 $Y=1.01 $X2=-0.19
+ $Y2=-0.245
cc_320 N_A_28_74#_M1008_g N_VGND_c_1770_n 0.00110513f $X=1.41 $Y=0.79 $X2=0
+ $Y2=0
cc_321 N_A_28_74#_c_269_n N_VGND_c_1770_n 0.0191765f $X=0.285 $Y=0.515 $X2=0
+ $Y2=0
cc_322 N_A_28_74#_c_271_n N_VGND_c_1770_n 0.0257907f $X=1.005 $Y=1.095 $X2=0
+ $Y2=0
cc_323 N_A_28_74#_c_273_n N_VGND_c_1770_n 0.0318061f $X=1.205 $Y=1.01 $X2=0
+ $Y2=0
cc_324 N_A_28_74#_c_275_n N_VGND_c_1770_n 0.0150382f $X=1.29 $Y=0.34 $X2=0 $Y2=0
cc_325 N_A_28_74#_c_269_n N_VGND_c_1774_n 0.0145639f $X=0.285 $Y=0.515 $X2=0
+ $Y2=0
cc_326 N_A_28_74#_M1008_g N_VGND_c_1775_n 7.64118e-19 $X=1.41 $Y=0.79 $X2=0
+ $Y2=0
cc_327 N_A_28_74#_c_274_n N_VGND_c_1775_n 0.100421f $X=2.585 $Y=0.34 $X2=0 $Y2=0
cc_328 N_A_28_74#_c_275_n N_VGND_c_1775_n 0.0121867f $X=1.29 $Y=0.34 $X2=0 $Y2=0
cc_329 N_A_28_74#_c_269_n N_VGND_c_1779_n 0.0119984f $X=0.285 $Y=0.515 $X2=0
+ $Y2=0
cc_330 N_A_28_74#_c_274_n N_VGND_c_1779_n 0.0576395f $X=2.585 $Y=0.34 $X2=0
+ $Y2=0
cc_331 N_A_28_74#_c_275_n N_VGND_c_1779_n 0.00660921f $X=1.29 $Y=0.34 $X2=0
+ $Y2=0
cc_332 N_A_492_48#_c_373_n N_B_c_543_n 0.00874716f $X=3.485 $Y=1.522 $X2=-0.19
+ $Y2=-0.245
cc_333 N_A_492_48#_M1025_g N_B_c_543_n 0.00681957f $X=3.645 $Y=0.915 $X2=-0.19
+ $Y2=-0.245
cc_334 N_A_492_48#_c_389_n N_B_c_555_n 0.0120822f $X=2.55 $Y=2.015 $X2=0 $Y2=0
cc_335 N_A_492_48#_c_373_n N_B_c_555_n 0.0080578f $X=3.485 $Y=1.522 $X2=0 $Y2=0
cc_336 N_A_492_48#_c_374_n N_B_c_555_n 0.0157531f $X=3.575 $Y=1.82 $X2=0 $Y2=0
cc_337 N_A_492_48#_M1025_g N_B_c_544_n 0.00897756f $X=3.645 $Y=0.915 $X2=0 $Y2=0
cc_338 N_A_492_48#_c_381_n N_B_c_544_n 0.00157877f $X=4.285 $Y=0.34 $X2=0 $Y2=0
cc_339 N_A_492_48#_M1014_g N_B_c_545_n 0.0215747f $X=2.535 $Y=0.69 $X2=0 $Y2=0
cc_340 N_A_492_48#_c_374_n N_B_c_556_n 0.00882199f $X=3.575 $Y=1.82 $X2=0 $Y2=0
cc_341 N_A_492_48#_c_389_n N_B_c_557_n 0.00204236f $X=2.55 $Y=2.015 $X2=0 $Y2=0
cc_342 N_A_492_48#_c_374_n N_B_c_558_n 7.79787e-19 $X=3.575 $Y=1.82 $X2=0 $Y2=0
cc_343 N_A_492_48#_c_374_n N_B_c_560_n 0.0164566f $X=3.575 $Y=1.82 $X2=0 $Y2=0
cc_344 N_A_492_48#_c_385_n N_B_c_560_n 0.00121094f $X=3.825 $Y=1.545 $X2=0 $Y2=0
cc_345 N_A_492_48#_M1025_g N_B_M1031_g 0.0128894f $X=3.645 $Y=0.915 $X2=0 $Y2=0
cc_346 N_A_492_48#_c_379_n N_B_M1031_g 0.0246091f $X=4.2 $Y=1.38 $X2=0 $Y2=0
cc_347 N_A_492_48#_c_380_n N_B_M1031_g 0.00900113f $X=4.965 $Y=0.34 $X2=0 $Y2=0
cc_348 N_A_492_48#_c_381_n N_B_M1031_g 0.00367885f $X=4.285 $Y=0.34 $X2=0 $Y2=0
cc_349 N_A_492_48#_c_380_n N_B_c_547_n 0.00469669f $X=4.965 $Y=0.34 $X2=0 $Y2=0
cc_350 N_A_492_48#_c_397_n N_B_c_548_n 0.00373656f $X=5.12 $Y=1.905 $X2=0 $Y2=0
cc_351 N_A_492_48#_c_379_n N_B_c_549_n 0.00137564f $X=4.2 $Y=1.38 $X2=0 $Y2=0
cc_352 N_A_492_48#_c_380_n N_B_c_549_n 0.0154235f $X=4.965 $Y=0.34 $X2=0 $Y2=0
cc_353 N_A_492_48#_c_382_n N_B_c_549_n 0.00863609f $X=5.13 $Y=0.585 $X2=0 $Y2=0
cc_354 N_A_492_48#_c_383_n N_B_c_549_n 0.00188605f $X=5.295 $Y=0.925 $X2=0 $Y2=0
cc_355 N_A_492_48#_c_376_n N_B_c_563_n 0.0287883f $X=5.91 $Y=1.765 $X2=0 $Y2=0
cc_356 N_A_492_48#_c_394_n N_B_c_563_n 0.013447f $X=5.63 $Y=1.905 $X2=0 $Y2=0
cc_357 N_A_492_48#_c_384_n N_B_c_563_n 0.00113245f $X=5.715 $Y=1.82 $X2=0 $Y2=0
cc_358 N_A_492_48#_c_397_n N_B_c_563_n 0.00667126f $X=5.12 $Y=1.905 $X2=0 $Y2=0
cc_359 N_A_492_48#_c_381_n N_B_c_550_n 4.71126e-19 $X=4.285 $Y=0.34 $X2=0 $Y2=0
cc_360 N_A_492_48#_c_376_n N_B_c_552_n 0.0225969f $X=5.91 $Y=1.765 $X2=0 $Y2=0
cc_361 N_A_492_48#_c_394_n N_B_c_552_n 7.05791e-19 $X=5.63 $Y=1.905 $X2=0 $Y2=0
cc_362 N_A_492_48#_c_383_n N_B_c_552_n 0.00127052f $X=5.295 $Y=0.925 $X2=0 $Y2=0
cc_363 N_A_492_48#_c_397_n N_B_c_552_n 0.00467581f $X=5.12 $Y=1.905 $X2=0 $Y2=0
cc_364 N_A_492_48#_c_386_n N_B_c_552_n 0.00578495f $X=5.84 $Y=1.42 $X2=0 $Y2=0
cc_365 N_A_492_48#_M1027_g N_B_c_553_n 0.0145618f $X=6.09 $Y=0.725 $X2=0 $Y2=0
cc_366 N_A_492_48#_c_380_n N_B_c_553_n 0.00354135f $X=4.965 $Y=0.34 $X2=0 $Y2=0
cc_367 N_A_492_48#_c_382_n N_B_c_553_n 0.0106025f $X=5.13 $Y=0.585 $X2=0 $Y2=0
cc_368 N_A_492_48#_c_440_p N_B_c_553_n 0.0143185f $X=5.63 $Y=0.925 $X2=0 $Y2=0
cc_369 N_A_492_48#_c_383_n N_B_c_553_n 6.11309e-19 $X=5.295 $Y=0.925 $X2=0 $Y2=0
cc_370 N_A_492_48#_c_387_n N_B_c_553_n 0.00578495f $X=5.8 $Y=1.255 $X2=0 $Y2=0
cc_371 N_A_492_48#_c_376_n B 2.88108e-19 $X=5.91 $Y=1.765 $X2=0 $Y2=0
cc_372 N_A_492_48#_c_383_n B 0.0211671f $X=5.295 $Y=0.925 $X2=0 $Y2=0
cc_373 N_A_492_48#_c_397_n B 0.0145403f $X=5.12 $Y=1.905 $X2=0 $Y2=0
cc_374 N_A_492_48#_c_387_n B 0.0163239f $X=5.8 $Y=1.255 $X2=0 $Y2=0
cc_375 N_A_492_48#_c_376_n N_A_608_74#_c_685_n 0.0316496f $X=5.91 $Y=1.765 $X2=0
+ $Y2=0
cc_376 N_A_492_48#_c_374_n N_A_608_74#_c_705_n 0.0103628f $X=3.575 $Y=1.82 $X2=0
+ $Y2=0
cc_377 N_A_492_48#_c_373_n N_A_608_74#_c_691_n 0.0161982f $X=3.485 $Y=1.522
+ $X2=0 $Y2=0
cc_378 N_A_492_48#_c_374_n N_A_608_74#_c_691_n 0.0159819f $X=3.575 $Y=1.82 $X2=0
+ $Y2=0
cc_379 N_A_492_48#_M1025_g N_A_608_74#_c_691_n 0.00392847f $X=3.645 $Y=0.915
+ $X2=0 $Y2=0
cc_380 N_A_492_48#_c_379_n N_A_608_74#_c_691_n 0.00601997f $X=4.2 $Y=1.38 $X2=0
+ $Y2=0
cc_381 N_A_492_48#_c_385_n N_A_608_74#_c_691_n 0.0242286f $X=3.825 $Y=1.545
+ $X2=0 $Y2=0
cc_382 N_A_492_48#_c_374_n N_A_608_74#_c_707_n 0.0180989f $X=3.575 $Y=1.82 $X2=0
+ $Y2=0
cc_383 N_A_492_48#_c_385_n N_A_608_74#_c_707_n 0.034138f $X=3.825 $Y=1.545 $X2=0
+ $Y2=0
cc_384 N_A_492_48#_c_374_n N_A_608_74#_c_708_n 0.00216189f $X=3.575 $Y=1.82
+ $X2=0 $Y2=0
cc_385 N_A_492_48#_M1007_s N_A_608_74#_c_709_n 6.70056e-19 $X=4.975 $Y=1.84
+ $X2=0 $Y2=0
cc_386 N_A_492_48#_M1007_s N_A_608_74#_c_741_n 0.00406933f $X=4.975 $Y=1.84
+ $X2=0 $Y2=0
cc_387 N_A_492_48#_M1007_s N_A_608_74#_c_742_n 0.00491282f $X=4.975 $Y=1.84
+ $X2=0 $Y2=0
cc_388 N_A_492_48#_c_376_n N_A_608_74#_c_742_n 0.0134577f $X=5.91 $Y=1.765 $X2=0
+ $Y2=0
cc_389 N_A_492_48#_c_394_n N_A_608_74#_c_742_n 0.0108f $X=5.63 $Y=1.905 $X2=0
+ $Y2=0
cc_390 N_A_492_48#_c_397_n N_A_608_74#_c_742_n 0.0131127f $X=5.12 $Y=1.905 $X2=0
+ $Y2=0
cc_391 N_A_492_48#_M1007_s N_A_608_74#_c_711_n 7.26895e-19 $X=4.975 $Y=1.84
+ $X2=0 $Y2=0
cc_392 N_A_492_48#_c_397_n N_A_608_74#_c_711_n 0.00722023f $X=5.12 $Y=1.905
+ $X2=0 $Y2=0
cc_393 N_A_492_48#_c_376_n N_A_608_74#_c_712_n 0.00650445f $X=5.91 $Y=1.765
+ $X2=0 $Y2=0
cc_394 N_A_492_48#_c_376_n N_A_608_74#_c_713_n 7.79828e-19 $X=5.91 $Y=1.765
+ $X2=0 $Y2=0
cc_395 N_A_492_48#_c_376_n N_A_608_74#_c_715_n 7.37926e-19 $X=5.91 $Y=1.765
+ $X2=0 $Y2=0
cc_396 N_A_492_48#_c_373_n N_A_608_74#_c_720_n 0.00670871f $X=3.485 $Y=1.522
+ $X2=0 $Y2=0
cc_397 N_A_492_48#_c_374_n N_A_608_74#_c_720_n 7.22214e-19 $X=3.575 $Y=1.82
+ $X2=0 $Y2=0
cc_398 N_A_492_48#_c_376_n N_A_608_74#_c_699_n 2.12915e-19 $X=5.91 $Y=1.765
+ $X2=0 $Y2=0
cc_399 N_A_492_48#_M1027_g N_A_430_418#_c_950_n 0.00791982f $X=6.09 $Y=0.725
+ $X2=0 $Y2=0
cc_400 N_A_492_48#_c_376_n N_A_430_418#_c_952_n 0.00791982f $X=5.91 $Y=1.765
+ $X2=0 $Y2=0
cc_401 N_A_492_48#_M1014_g N_A_430_418#_c_955_n 0.0259633f $X=2.535 $Y=0.69
+ $X2=0 $Y2=0
cc_402 N_A_492_48#_c_374_n N_A_430_418#_c_956_n 0.00157045f $X=3.575 $Y=1.82
+ $X2=0 $Y2=0
cc_403 N_A_492_48#_c_379_n N_A_430_418#_c_956_n 0.0516033f $X=4.2 $Y=1.38 $X2=0
+ $Y2=0
cc_404 N_A_492_48#_c_380_n N_A_430_418#_c_956_n 0.0141693f $X=4.965 $Y=0.34
+ $X2=0 $Y2=0
cc_405 N_A_492_48#_c_382_n N_A_430_418#_c_956_n 0.0102652f $X=5.13 $Y=0.585
+ $X2=0 $Y2=0
cc_406 N_A_492_48#_c_383_n N_A_430_418#_c_956_n 0.0109342f $X=5.295 $Y=0.925
+ $X2=0 $Y2=0
cc_407 N_A_492_48#_c_385_n N_A_430_418#_c_956_n 0.0204142f $X=3.825 $Y=1.545
+ $X2=0 $Y2=0
cc_408 N_A_492_48#_c_397_n N_A_430_418#_c_956_n 0.0216873f $X=5.12 $Y=1.905
+ $X2=0 $Y2=0
cc_409 N_A_492_48#_c_389_n N_A_430_418#_c_967_n 0.0117688f $X=2.55 $Y=2.015
+ $X2=0 $Y2=0
cc_410 N_A_492_48#_c_373_n N_A_430_418#_c_967_n 0.00623437f $X=3.485 $Y=1.522
+ $X2=0 $Y2=0
cc_411 N_A_492_48#_c_374_n N_A_430_418#_c_967_n 0.00615332f $X=3.575 $Y=1.82
+ $X2=0 $Y2=0
cc_412 N_A_492_48#_c_385_n N_A_430_418#_c_967_n 0.00415724f $X=3.825 $Y=1.545
+ $X2=0 $Y2=0
cc_413 N_A_492_48#_c_376_n N_A_430_418#_c_969_n 0.00454084f $X=5.91 $Y=1.765
+ $X2=0 $Y2=0
cc_414 N_A_492_48#_c_394_n N_A_430_418#_c_969_n 0.0277257f $X=5.63 $Y=1.905
+ $X2=0 $Y2=0
cc_415 N_A_492_48#_c_397_n N_A_430_418#_c_969_n 0.0200122f $X=5.12 $Y=1.905
+ $X2=0 $Y2=0
cc_416 N_A_492_48#_c_386_n N_A_430_418#_c_969_n 0.00557311f $X=5.84 $Y=1.42
+ $X2=0 $Y2=0
cc_417 N_A_492_48#_c_397_n N_A_430_418#_c_970_n 0.00250307f $X=5.12 $Y=1.905
+ $X2=0 $Y2=0
cc_418 N_A_492_48#_c_388_n N_A_430_418#_c_973_n 0.0031695f $X=2.55 $Y=1.925
+ $X2=0 $Y2=0
cc_419 N_A_492_48#_c_389_n N_A_430_418#_c_973_n 0.00537063f $X=2.55 $Y=2.015
+ $X2=0 $Y2=0
cc_420 N_A_492_48#_c_394_n N_VPWR_M1007_d 0.00441072f $X=5.63 $Y=1.905 $X2=0
+ $Y2=0
cc_421 N_A_492_48#_c_376_n N_VPWR_c_1402_n 0.00295065f $X=5.91 $Y=1.765 $X2=0
+ $Y2=0
cc_422 N_A_492_48#_c_376_n N_VPWR_c_1405_n 0.0049405f $X=5.91 $Y=1.765 $X2=0
+ $Y2=0
cc_423 N_A_492_48#_c_389_n N_VPWR_c_1408_n 9.29978e-19 $X=2.55 $Y=2.015 $X2=0
+ $Y2=0
cc_424 N_A_492_48#_c_376_n N_VPWR_c_1400_n 0.00508379f $X=5.91 $Y=1.765 $X2=0
+ $Y2=0
cc_425 N_A_492_48#_c_379_n N_A_256_368#_M1025_d 0.00657304f $X=4.2 $Y=1.38 $X2=0
+ $Y2=0
cc_426 N_A_492_48#_c_389_n N_A_256_368#_c_1505_n 0.00374685f $X=2.55 $Y=2.015
+ $X2=0 $Y2=0
cc_427 N_A_492_48#_c_389_n N_A_256_368#_c_1506_n 0.0115042f $X=2.55 $Y=2.015
+ $X2=0 $Y2=0
cc_428 N_A_492_48#_c_389_n N_A_256_368#_c_1508_n 5.56999e-19 $X=2.55 $Y=2.015
+ $X2=0 $Y2=0
cc_429 N_A_492_48#_c_373_n N_A_256_368#_c_1508_n 0.00430547f $X=3.485 $Y=1.522
+ $X2=0 $Y2=0
cc_430 N_A_492_48#_M1014_g N_A_256_368#_c_1534_n 6.2386e-19 $X=2.535 $Y=0.69
+ $X2=0 $Y2=0
cc_431 N_A_492_48#_M1025_g N_A_256_368#_c_1534_n 0.00147462f $X=3.645 $Y=0.915
+ $X2=0 $Y2=0
cc_432 N_A_492_48#_M1025_g N_A_256_368#_c_1499_n 0.00307819f $X=3.645 $Y=0.915
+ $X2=0 $Y2=0
cc_433 N_A_492_48#_c_381_n N_A_256_368#_c_1499_n 0.0159272f $X=4.285 $Y=0.34
+ $X2=0 $Y2=0
cc_434 N_A_492_48#_c_374_n N_A_256_368#_c_1500_n 0.00147467f $X=3.575 $Y=1.82
+ $X2=0 $Y2=0
cc_435 N_A_492_48#_M1025_g N_A_256_368#_c_1500_n 0.0123007f $X=3.645 $Y=0.915
+ $X2=0 $Y2=0
cc_436 N_A_492_48#_c_379_n N_A_256_368#_c_1500_n 0.052748f $X=4.2 $Y=1.38 $X2=0
+ $Y2=0
cc_437 N_A_492_48#_c_385_n N_A_256_368#_c_1500_n 0.0130785f $X=3.825 $Y=1.545
+ $X2=0 $Y2=0
cc_438 N_A_492_48#_M1014_g N_A_256_368#_c_1503_n 0.00534131f $X=2.535 $Y=0.69
+ $X2=0 $Y2=0
cc_439 N_A_492_48#_c_388_n N_A_256_368#_c_1503_n 0.00691306f $X=2.55 $Y=1.925
+ $X2=0 $Y2=0
cc_440 N_A_492_48#_c_373_n N_A_256_368#_c_1503_n 0.0221613f $X=3.485 $Y=1.522
+ $X2=0 $Y2=0
cc_441 N_A_492_48#_c_374_n N_A_256_368#_c_1503_n 0.00140042f $X=3.575 $Y=1.82
+ $X2=0 $Y2=0
cc_442 N_A_492_48#_M1014_g N_A_256_368#_c_1504_n 0.00141098f $X=2.535 $Y=0.69
+ $X2=0 $Y2=0
cc_443 N_A_492_48#_c_373_n N_A_256_368#_c_1504_n 0.00508507f $X=3.485 $Y=1.522
+ $X2=0 $Y2=0
cc_444 N_A_492_48#_M1027_g N_A_1197_368#_c_1593_n 0.0129141f $X=6.09 $Y=0.725
+ $X2=0 $Y2=0
cc_445 N_A_492_48#_c_440_p N_A_1197_368#_c_1593_n 0.00821874f $X=5.63 $Y=0.925
+ $X2=0 $Y2=0
cc_446 N_A_492_48#_c_376_n N_A_1197_368#_c_1596_n 0.0141571f $X=5.91 $Y=1.765
+ $X2=0 $Y2=0
cc_447 N_A_492_48#_c_394_n N_A_1197_368#_c_1596_n 0.00762374f $X=5.63 $Y=1.905
+ $X2=0 $Y2=0
cc_448 N_A_492_48#_c_376_n N_A_1197_368#_c_1594_n 0.0127319f $X=5.91 $Y=1.765
+ $X2=0 $Y2=0
cc_449 N_A_492_48#_M1027_g N_A_1197_368#_c_1594_n 0.00421254f $X=6.09 $Y=0.725
+ $X2=0 $Y2=0
cc_450 N_A_492_48#_c_384_n N_A_1197_368#_c_1594_n 0.0108481f $X=5.715 $Y=1.82
+ $X2=0 $Y2=0
cc_451 N_A_492_48#_c_386_n N_A_1197_368#_c_1594_n 0.0236229f $X=5.84 $Y=1.42
+ $X2=0 $Y2=0
cc_452 N_A_492_48#_M1027_g N_A_1197_368#_c_1595_n 0.00270236f $X=6.09 $Y=0.725
+ $X2=0 $Y2=0
cc_453 N_A_492_48#_c_387_n N_A_1197_368#_c_1595_n 0.0104428f $X=5.8 $Y=1.255
+ $X2=0 $Y2=0
cc_454 N_A_492_48#_c_376_n N_COUT_c_1631_n 2.07873e-19 $X=5.91 $Y=1.765 $X2=0
+ $Y2=0
cc_455 N_A_492_48#_c_440_p N_VGND_M1015_d 0.0125322f $X=5.63 $Y=0.925 $X2=0
+ $Y2=0
cc_456 N_A_492_48#_c_387_n N_VGND_M1015_d 0.00237231f $X=5.8 $Y=1.255 $X2=0
+ $Y2=0
cc_457 N_A_492_48#_c_376_n N_VGND_c_1771_n 0.00143519f $X=5.91 $Y=1.765 $X2=0
+ $Y2=0
cc_458 N_A_492_48#_M1027_g N_VGND_c_1771_n 0.00570238f $X=6.09 $Y=0.725 $X2=0
+ $Y2=0
cc_459 N_A_492_48#_c_380_n N_VGND_c_1771_n 0.0138907f $X=4.965 $Y=0.34 $X2=0
+ $Y2=0
cc_460 N_A_492_48#_c_440_p N_VGND_c_1771_n 0.0222657f $X=5.63 $Y=0.925 $X2=0
+ $Y2=0
cc_461 N_A_492_48#_c_386_n N_VGND_c_1771_n 0.00488384f $X=5.84 $Y=1.42 $X2=0
+ $Y2=0
cc_462 N_A_492_48#_M1014_g N_VGND_c_1775_n 0.00278247f $X=2.535 $Y=0.69 $X2=0
+ $Y2=0
cc_463 N_A_492_48#_c_380_n N_VGND_c_1775_n 0.0666882f $X=4.965 $Y=0.34 $X2=0
+ $Y2=0
cc_464 N_A_492_48#_c_381_n N_VGND_c_1775_n 0.0115566f $X=4.285 $Y=0.34 $X2=0
+ $Y2=0
cc_465 N_A_492_48#_M1027_g N_VGND_c_1776_n 0.00527282f $X=6.09 $Y=0.725 $X2=0
+ $Y2=0
cc_466 N_A_492_48#_M1014_g N_VGND_c_1779_n 0.00358523f $X=2.535 $Y=0.69 $X2=0
+ $Y2=0
cc_467 N_A_492_48#_M1027_g N_VGND_c_1779_n 0.00534666f $X=6.09 $Y=0.725 $X2=0
+ $Y2=0
cc_468 N_A_492_48#_c_380_n N_VGND_c_1779_n 0.0357004f $X=4.965 $Y=0.34 $X2=0
+ $Y2=0
cc_469 N_A_492_48#_c_381_n N_VGND_c_1779_n 0.00579705f $X=4.285 $Y=0.34 $X2=0
+ $Y2=0
cc_470 N_A_492_48#_c_440_p N_VGND_c_1779_n 0.00667209f $X=5.63 $Y=0.925 $X2=0
+ $Y2=0
cc_471 N_B_c_555_n N_A_608_74#_c_705_n 0.00613299f $X=3.04 $Y=3.005 $X2=0 $Y2=0
cc_472 N_B_c_543_n N_A_608_74#_c_691_n 0.00176537f $X=2.965 $Y=0.255 $X2=0 $Y2=0
cc_473 N_B_c_560_n N_A_608_74#_c_707_n 0.00574142f $X=4.29 $Y=2.81 $X2=0 $Y2=0
cc_474 N_B_c_558_n N_A_608_74#_c_708_n 0.00362613f $X=4.29 $Y=2.9 $X2=0 $Y2=0
cc_475 N_B_c_560_n N_A_608_74#_c_708_n 0.0187451f $X=4.29 $Y=2.81 $X2=0 $Y2=0
cc_476 N_B_c_548_n N_A_608_74#_c_708_n 7.27788e-19 $X=4.825 $Y=3.075 $X2=0 $Y2=0
cc_477 N_B_c_559_n N_A_608_74#_c_709_n 0.00948559f $X=4.29 $Y=3.075 $X2=0 $Y2=0
cc_478 N_B_c_561_n N_A_608_74#_c_709_n 0.004676f $X=4.75 $Y=3.15 $X2=0 $Y2=0
cc_479 N_B_c_548_n N_A_608_74#_c_709_n 0.0129047f $X=4.825 $Y=3.075 $X2=0 $Y2=0
cc_480 N_B_c_563_n N_A_608_74#_c_709_n 0.0015709f $X=5.345 $Y=1.765 $X2=0 $Y2=0
cc_481 N_B_c_556_n N_A_608_74#_c_710_n 0.00232404f $X=4.2 $Y=3.15 $X2=0 $Y2=0
cc_482 N_B_c_559_n N_A_608_74#_c_710_n 0.00391879f $X=4.29 $Y=3.075 $X2=0 $Y2=0
cc_483 N_B_c_564_n N_A_608_74#_c_710_n 6.42445e-19 $X=4.29 $Y=3.15 $X2=0 $Y2=0
cc_484 N_B_c_558_n N_A_608_74#_c_741_n 2.99669e-19 $X=4.29 $Y=2.9 $X2=0 $Y2=0
cc_485 N_B_c_560_n N_A_608_74#_c_741_n 2.67397e-19 $X=4.29 $Y=2.81 $X2=0 $Y2=0
cc_486 N_B_c_548_n N_A_608_74#_c_741_n 0.00819436f $X=4.825 $Y=3.075 $X2=0 $Y2=0
cc_487 N_B_c_563_n N_A_608_74#_c_741_n 0.00476127f $X=5.345 $Y=1.765 $X2=0 $Y2=0
cc_488 N_B_c_563_n N_A_608_74#_c_742_n 0.0136173f $X=5.345 $Y=1.765 $X2=0 $Y2=0
cc_489 N_B_c_548_n N_A_608_74#_c_711_n 0.00481538f $X=4.825 $Y=3.075 $X2=0 $Y2=0
cc_490 N_B_c_555_n N_A_608_74#_c_720_n 7.1167e-19 $X=3.04 $Y=3.005 $X2=0 $Y2=0
cc_491 N_B_c_560_n N_A_430_418#_c_956_n 0.00282109f $X=4.29 $Y=2.81 $X2=0 $Y2=0
cc_492 N_B_M1031_g N_A_430_418#_c_956_n 0.00362758f $X=4.305 $Y=0.915 $X2=0
+ $Y2=0
cc_493 N_B_c_549_n N_A_430_418#_c_956_n 0.0118737f $X=4.835 $Y=1.255 $X2=0 $Y2=0
cc_494 N_B_c_551_n N_A_430_418#_c_956_n 0.012449f $X=4.75 $Y=1.435 $X2=0 $Y2=0
cc_495 B N_A_430_418#_c_956_n 0.0313157f $X=4.955 $Y=1.21 $X2=0 $Y2=0
cc_496 N_B_c_560_n N_A_430_418#_c_966_n 0.00329463f $X=4.29 $Y=2.81 $X2=0 $Y2=0
cc_497 N_B_c_548_n N_A_430_418#_c_966_n 0.012449f $X=4.825 $Y=3.075 $X2=0 $Y2=0
cc_498 N_B_c_555_n N_A_430_418#_c_967_n 0.00890743f $X=3.04 $Y=3.005 $X2=0 $Y2=0
cc_499 N_B_c_560_n N_A_430_418#_c_967_n 0.00521341f $X=4.29 $Y=2.81 $X2=0 $Y2=0
cc_500 N_B_M1031_g N_A_430_418#_c_967_n 7.23332e-19 $X=4.305 $Y=0.915 $X2=0
+ $Y2=0
cc_501 N_B_c_548_n N_A_430_418#_c_969_n 0.013348f $X=4.825 $Y=3.075 $X2=0 $Y2=0
cc_502 N_B_c_563_n N_A_430_418#_c_969_n 0.00239266f $X=5.345 $Y=1.765 $X2=0
+ $Y2=0
cc_503 B N_A_430_418#_c_969_n 0.00418222f $X=4.955 $Y=1.21 $X2=0 $Y2=0
cc_504 N_B_c_548_n N_A_430_418#_c_970_n 0.00157474f $X=4.825 $Y=3.075 $X2=0
+ $Y2=0
cc_505 N_B_c_561_n N_VPWR_c_1402_n 0.00243239f $X=4.75 $Y=3.15 $X2=0 $Y2=0
cc_506 N_B_c_548_n N_VPWR_c_1402_n 3.07893e-19 $X=4.825 $Y=3.075 $X2=0 $Y2=0
cc_507 N_B_c_563_n N_VPWR_c_1402_n 0.00818159f $X=5.345 $Y=1.765 $X2=0 $Y2=0
cc_508 N_B_c_557_n N_VPWR_c_1408_n 0.0441946f $X=3.13 $Y=3.15 $X2=0 $Y2=0
cc_509 N_B_c_563_n N_VPWR_c_1408_n 0.00413917f $X=5.345 $Y=1.765 $X2=0 $Y2=0
cc_510 N_B_c_556_n N_VPWR_c_1400_n 0.0302019f $X=4.2 $Y=3.15 $X2=0 $Y2=0
cc_511 N_B_c_557_n N_VPWR_c_1400_n 0.00674634f $X=3.13 $Y=3.15 $X2=0 $Y2=0
cc_512 N_B_c_561_n N_VPWR_c_1400_n 0.0148287f $X=4.75 $Y=3.15 $X2=0 $Y2=0
cc_513 N_B_c_563_n N_VPWR_c_1400_n 0.00399275f $X=5.345 $Y=1.765 $X2=0 $Y2=0
cc_514 N_B_c_564_n N_VPWR_c_1400_n 0.00441518f $X=4.29 $Y=3.15 $X2=0 $Y2=0
cc_515 N_B_c_555_n N_A_256_368#_c_1508_n 0.00199825f $X=3.04 $Y=3.005 $X2=0
+ $Y2=0
cc_516 N_B_c_555_n N_A_256_368#_c_1516_n 0.00196378f $X=3.04 $Y=3.005 $X2=0
+ $Y2=0
cc_517 N_B_c_555_n N_A_256_368#_c_1550_n 0.00412674f $X=3.04 $Y=3.005 $X2=0
+ $Y2=0
cc_518 N_B_c_543_n N_A_256_368#_c_1534_n 0.0129263f $X=2.965 $Y=0.255 $X2=0
+ $Y2=0
cc_519 N_B_c_544_n N_A_256_368#_c_1499_n 0.015881f $X=4.23 $Y=0.18 $X2=0 $Y2=0
cc_520 N_B_M1031_g N_A_256_368#_c_1499_n 0.00101961f $X=4.305 $Y=0.915 $X2=0
+ $Y2=0
cc_521 N_B_c_543_n N_A_256_368#_c_1517_n 0.00591399f $X=2.965 $Y=0.255 $X2=0
+ $Y2=0
cc_522 N_B_c_544_n N_A_256_368#_c_1517_n 0.00217912f $X=4.23 $Y=0.18 $X2=0 $Y2=0
cc_523 N_B_c_545_n N_A_256_368#_c_1517_n 2.91242e-19 $X=3.04 $Y=0.18 $X2=0 $Y2=0
cc_524 N_B_c_543_n N_A_256_368#_c_1500_n 3.57076e-19 $X=2.965 $Y=0.255 $X2=0
+ $Y2=0
cc_525 N_B_M1031_g N_A_256_368#_c_1500_n 0.00221237f $X=4.305 $Y=0.915 $X2=0
+ $Y2=0
cc_526 N_B_c_543_n N_A_256_368#_c_1503_n 0.002458f $X=2.965 $Y=0.255 $X2=0 $Y2=0
cc_527 N_B_c_555_n N_A_256_368#_c_1503_n 0.0014973f $X=3.04 $Y=3.005 $X2=0 $Y2=0
cc_528 N_B_c_543_n N_A_256_368#_c_1504_n 0.0115084f $X=2.965 $Y=0.255 $X2=0
+ $Y2=0
cc_529 N_B_c_563_n N_A_1197_368#_c_1596_n 0.00135989f $X=5.345 $Y=1.765 $X2=0
+ $Y2=0
cc_530 N_B_c_547_n N_VGND_c_1771_n 0.00258065f $X=4.76 $Y=0.18 $X2=0 $Y2=0
cc_531 N_B_c_553_n N_VGND_c_1771_n 0.0033927f $X=5.345 $Y=1.255 $X2=0 $Y2=0
cc_532 N_B_c_545_n N_VGND_c_1775_n 0.047914f $X=3.04 $Y=0.18 $X2=0 $Y2=0
cc_533 N_B_c_553_n N_VGND_c_1775_n 0.00521619f $X=5.345 $Y=1.255 $X2=0 $Y2=0
cc_534 N_B_c_544_n N_VGND_c_1779_n 0.0332509f $X=4.23 $Y=0.18 $X2=0 $Y2=0
cc_535 N_B_c_545_n N_VGND_c_1779_n 0.0102556f $X=3.04 $Y=0.18 $X2=0 $Y2=0
cc_536 N_B_c_547_n N_VGND_c_1779_n 0.0151063f $X=4.76 $Y=0.18 $X2=0 $Y2=0
cc_537 N_B_c_550_n N_VGND_c_1779_n 0.00370842f $X=4.305 $Y=0.18 $X2=0 $Y2=0
cc_538 N_B_c_553_n N_VGND_c_1779_n 0.00499022f $X=5.345 $Y=1.255 $X2=0 $Y2=0
cc_539 N_A_608_74#_c_686_n N_A_430_418#_c_951_n 0.00103362f $X=8.085 $Y=1.155
+ $X2=0 $Y2=0
cc_540 N_A_608_74#_c_700_n N_A_430_418#_c_951_n 4.56844e-19 $X=7.91 $Y=1.32
+ $X2=0 $Y2=0
cc_541 N_A_608_74#_c_701_n N_A_430_418#_c_951_n 0.0211413f $X=8.085 $Y=1.32
+ $X2=0 $Y2=0
cc_542 N_A_608_74#_c_685_n N_A_430_418#_c_952_n 0.0182942f $X=6.495 $Y=1.925
+ $X2=0 $Y2=0
cc_543 N_A_608_74#_c_699_n N_A_430_418#_c_952_n 0.00114907f $X=6.605 $Y=1.675
+ $X2=0 $Y2=0
cc_544 N_A_608_74#_c_692_n N_A_430_418#_c_960_n 0.0101161f $X=7.87 $Y=2.905
+ $X2=0 $Y2=0
cc_545 N_A_608_74#_c_700_n N_A_430_418#_c_960_n 5.05061e-19 $X=7.91 $Y=1.32
+ $X2=0 $Y2=0
cc_546 N_A_608_74#_c_701_n N_A_430_418#_c_960_n 0.0132892f $X=8.085 $Y=1.32
+ $X2=0 $Y2=0
cc_547 N_A_608_74#_c_685_n N_A_430_418#_c_961_n 4.49838e-19 $X=6.495 $Y=1.925
+ $X2=0 $Y2=0
cc_548 N_A_608_74#_c_692_n N_A_430_418#_c_962_n 0.0322695f $X=7.87 $Y=2.905
+ $X2=0 $Y2=0
cc_549 N_A_608_74#_c_717_n N_A_430_418#_c_962_n 0.00230718f $X=8.545 $Y=2.99
+ $X2=0 $Y2=0
cc_550 N_A_608_74#_c_718_n N_A_430_418#_c_962_n 7.01078e-19 $X=8.63 $Y=2.905
+ $X2=0 $Y2=0
cc_551 N_A_608_74#_c_722_n N_A_430_418#_c_962_n 0.00448828f $X=7.87 $Y=2.99
+ $X2=0 $Y2=0
cc_552 N_A_608_74#_c_688_n N_A_430_418#_c_953_n 0.018548f $X=10.205 $Y=1.545
+ $X2=0 $Y2=0
cc_553 N_A_608_74#_c_704_n N_A_430_418#_c_953_n 0.0296667f $X=10.205 $Y=1.845
+ $X2=0 $Y2=0
cc_554 N_A_608_74#_c_688_n N_A_430_418#_c_954_n 5.77834e-19 $X=10.205 $Y=1.545
+ $X2=0 $Y2=0
cc_555 N_A_608_74#_c_698_n N_A_430_418#_c_954_n 0.00110913f $X=10.41 $Y=0.405
+ $X2=0 $Y2=0
cc_556 N_A_608_74#_c_707_n N_A_430_418#_c_966_n 0.0120951f $X=4.105 $Y=1.965
+ $X2=0 $Y2=0
cc_557 N_A_608_74#_M1029_d N_A_430_418#_c_967_n 0.00270048f $X=3.115 $Y=2.09
+ $X2=0 $Y2=0
cc_558 N_A_608_74#_c_705_n N_A_430_418#_c_967_n 0.0213703f $X=3.35 $Y=2.57 $X2=0
+ $Y2=0
cc_559 N_A_608_74#_c_707_n N_A_430_418#_c_967_n 0.0292954f $X=4.105 $Y=1.965
+ $X2=0 $Y2=0
cc_560 N_A_608_74#_c_708_n N_A_430_418#_c_967_n 0.0117692f $X=4.19 $Y=2.905
+ $X2=0 $Y2=0
cc_561 N_A_608_74#_c_720_n N_A_430_418#_c_967_n 0.012635f $X=3.35 $Y=2.04 $X2=0
+ $Y2=0
cc_562 N_A_608_74#_c_685_n N_A_430_418#_c_969_n 0.00555047f $X=6.495 $Y=1.925
+ $X2=0 $Y2=0
cc_563 N_A_608_74#_c_742_n N_A_430_418#_c_969_n 0.0206589f $X=6.15 $Y=2.475
+ $X2=0 $Y2=0
cc_564 N_A_608_74#_c_711_n N_A_430_418#_c_969_n 0.00420248f $X=5.045 $Y=2.475
+ $X2=0 $Y2=0
cc_565 N_A_608_74#_c_713_n N_A_430_418#_c_969_n 0.020978f $X=6.565 $Y=2.39 $X2=0
+ $Y2=0
cc_566 N_A_608_74#_c_801_p N_A_430_418#_c_969_n 0.0086273f $X=6.4 $Y=2.475 $X2=0
+ $Y2=0
cc_567 N_A_608_74#_c_699_n N_A_430_418#_c_969_n 0.00371687f $X=6.605 $Y=1.675
+ $X2=0 $Y2=0
cc_568 N_A_608_74#_c_707_n N_A_430_418#_c_970_n 0.0013519f $X=4.105 $Y=1.965
+ $X2=0 $Y2=0
cc_569 N_A_608_74#_c_708_n N_A_430_418#_c_970_n 0.00130949f $X=4.19 $Y=2.905
+ $X2=0 $Y2=0
cc_570 N_A_608_74#_c_688_n N_A_430_418#_c_971_n 0.00155821f $X=10.205 $Y=1.545
+ $X2=0 $Y2=0
cc_571 N_A_608_74#_c_704_n N_A_430_418#_c_971_n 0.00734195f $X=10.205 $Y=1.845
+ $X2=0 $Y2=0
cc_572 N_A_608_74#_c_692_n N_A_430_418#_c_971_n 0.0193609f $X=7.87 $Y=2.905
+ $X2=0 $Y2=0
cc_573 N_A_608_74#_c_718_n N_A_430_418#_c_971_n 0.0213523f $X=8.63 $Y=2.905
+ $X2=0 $Y2=0
cc_574 N_A_608_74#_c_693_n N_A_430_418#_c_971_n 0.024422f $X=9.215 $Y=1.74 $X2=0
+ $Y2=0
cc_575 N_A_608_74#_c_700_n N_A_430_418#_c_971_n 0.00375844f $X=7.91 $Y=1.32
+ $X2=0 $Y2=0
cc_576 N_A_608_74#_c_701_n N_A_430_418#_c_971_n 0.0021367f $X=8.085 $Y=1.32
+ $X2=0 $Y2=0
cc_577 N_A_608_74#_c_692_n N_A_430_418#_c_972_n 0.00257207f $X=7.87 $Y=2.905
+ $X2=0 $Y2=0
cc_578 N_A_608_74#_c_708_n N_A_430_418#_c_974_n 0.0489087f $X=4.19 $Y=2.905
+ $X2=0 $Y2=0
cc_579 N_A_608_74#_c_709_n N_A_430_418#_c_974_n 0.0200259f $X=4.875 $Y=2.99
+ $X2=0 $Y2=0
cc_580 N_A_608_74#_c_741_n N_A_430_418#_c_974_n 0.0129197f $X=4.96 $Y=2.905
+ $X2=0 $Y2=0
cc_581 N_A_608_74#_c_711_n N_A_430_418#_c_974_n 0.0140118f $X=5.045 $Y=2.475
+ $X2=0 $Y2=0
cc_582 N_A_608_74#_c_685_n N_A_430_418#_c_957_n 0.0070422f $X=6.495 $Y=1.925
+ $X2=0 $Y2=0
cc_583 N_A_608_74#_c_692_n N_A_430_418#_c_957_n 0.00150933f $X=7.87 $Y=2.905
+ $X2=0 $Y2=0
cc_584 N_A_608_74#_c_692_n N_A_430_418#_c_958_n 0.0358108f $X=7.87 $Y=2.905
+ $X2=0 $Y2=0
cc_585 N_A_608_74#_c_700_n N_A_430_418#_c_958_n 0.0226372f $X=7.91 $Y=1.32 $X2=0
+ $Y2=0
cc_586 N_A_608_74#_c_701_n N_A_430_418#_c_958_n 0.00183067f $X=8.085 $Y=1.32
+ $X2=0 $Y2=0
cc_587 N_A_608_74#_c_688_n N_A_430_418#_c_959_n 3.09256e-19 $X=10.205 $Y=1.545
+ $X2=0 $Y2=0
cc_588 N_A_608_74#_c_704_n N_A_430_418#_c_959_n 2.06554e-19 $X=10.205 $Y=1.845
+ $X2=0 $Y2=0
cc_589 N_A_608_74#_c_692_n N_CIN_c_1167_n 9.15402e-19 $X=7.87 $Y=2.905 $X2=-0.19
+ $Y2=-0.245
cc_590 N_A_608_74#_c_717_n N_CIN_c_1167_n 0.0108838f $X=8.545 $Y=2.99 $X2=-0.19
+ $Y2=-0.245
cc_591 N_A_608_74#_c_718_n N_CIN_c_1167_n 0.0251655f $X=8.63 $Y=2.905 $X2=-0.19
+ $Y2=-0.245
cc_592 N_A_608_74#_c_694_n N_CIN_c_1167_n 0.00172235f $X=8.715 $Y=1.74 $X2=-0.19
+ $Y2=-0.245
cc_593 N_A_608_74#_c_686_n N_CIN_c_1163_n 0.0155338f $X=8.085 $Y=1.155 $X2=0
+ $Y2=0
cc_594 N_A_608_74#_c_695_n N_CIN_c_1163_n 0.00433414f $X=9.3 $Y=1.655 $X2=0
+ $Y2=0
cc_595 N_A_608_74#_c_718_n N_CIN_c_1168_n 0.00393022f $X=8.63 $Y=2.905 $X2=0
+ $Y2=0
cc_596 N_A_608_74#_c_693_n N_CIN_c_1168_n 0.00525807f $X=9.215 $Y=1.74 $X2=0
+ $Y2=0
cc_597 N_A_608_74#_c_690_n N_CIN_c_1164_n 0.0078612f $X=10.02 $Y=0.405 $X2=0
+ $Y2=0
cc_598 N_A_608_74#_c_695_n N_CIN_c_1164_n 0.01354f $X=9.3 $Y=1.655 $X2=0 $Y2=0
cc_599 N_A_608_74#_c_697_n N_CIN_c_1164_n 0.0152526f $X=10.41 $Y=0.405 $X2=0
+ $Y2=0
cc_600 N_A_608_74#_c_693_n CIN 0.0231488f $X=9.215 $Y=1.74 $X2=0 $Y2=0
cc_601 N_A_608_74#_c_694_n CIN 7.37368e-19 $X=8.715 $Y=1.74 $X2=0 $Y2=0
cc_602 N_A_608_74#_c_695_n CIN 0.0231948f $X=9.3 $Y=1.655 $X2=0 $Y2=0
cc_603 N_A_608_74#_M1018_g N_CIN_c_1166_n 0.0078612f $X=9.945 $Y=1 $X2=0 $Y2=0
cc_604 N_A_608_74#_c_693_n N_CIN_c_1166_n 0.0179114f $X=9.215 $Y=1.74 $X2=0
+ $Y2=0
cc_605 N_A_608_74#_c_694_n N_CIN_c_1166_n 0.00753461f $X=8.715 $Y=1.74 $X2=0
+ $Y2=0
cc_606 N_A_608_74#_c_695_n N_CIN_c_1166_n 0.0186426f $X=9.3 $Y=1.655 $X2=0 $Y2=0
cc_607 N_A_608_74#_c_701_n N_CIN_c_1166_n 0.0172684f $X=8.085 $Y=1.32 $X2=0
+ $Y2=0
cc_608 N_A_608_74#_c_704_n N_A_1854_368#_c_1228_n 0.0046545f $X=10.205 $Y=1.845
+ $X2=0 $Y2=0
cc_609 N_A_608_74#_M1018_g N_A_1854_368#_c_1239_n 0.00465864f $X=9.945 $Y=1
+ $X2=0 $Y2=0
cc_610 N_A_608_74#_c_697_n N_A_1854_368#_c_1239_n 0.0227871f $X=10.41 $Y=0.405
+ $X2=0 $Y2=0
cc_611 N_A_608_74#_c_693_n N_A_1854_368#_c_1232_n 0.00843028f $X=9.215 $Y=1.74
+ $X2=0 $Y2=0
cc_612 N_A_608_74#_M1018_g N_A_1854_368#_c_1223_n 0.00235677f $X=9.945 $Y=1
+ $X2=0 $Y2=0
cc_613 N_A_608_74#_c_689_n N_A_1854_368#_c_1223_n 0.0053768f $X=10.205 $Y=1.755
+ $X2=0 $Y2=0
cc_614 N_A_608_74#_c_704_n N_A_1854_368#_c_1223_n 0.0016904f $X=10.205 $Y=1.845
+ $X2=0 $Y2=0
cc_615 N_A_608_74#_c_693_n N_A_1854_368#_c_1223_n 0.0143571f $X=9.215 $Y=1.74
+ $X2=0 $Y2=0
cc_616 N_A_608_74#_M1018_g N_A_1854_368#_c_1224_n 0.00322397f $X=9.945 $Y=1
+ $X2=0 $Y2=0
cc_617 N_A_608_74#_c_695_n N_A_1854_368#_c_1224_n 0.0245777f $X=9.3 $Y=1.655
+ $X2=0 $Y2=0
cc_618 N_A_608_74#_c_704_n N_A_1854_368#_c_1234_n 0.00512165f $X=10.205 $Y=1.845
+ $X2=0 $Y2=0
cc_619 N_A_608_74#_M1018_g N_A_2004_136#_c_1319_n 8.93644e-19 $X=9.945 $Y=1
+ $X2=0 $Y2=0
cc_620 N_A_608_74#_c_688_n N_A_2004_136#_c_1319_n 0.00572229f $X=10.205 $Y=1.545
+ $X2=0 $Y2=0
cc_621 N_A_608_74#_c_689_n N_A_2004_136#_c_1319_n 0.00614972f $X=10.205 $Y=1.755
+ $X2=0 $Y2=0
cc_622 N_A_608_74#_c_704_n N_A_2004_136#_c_1319_n 0.00789498f $X=10.205 $Y=1.845
+ $X2=0 $Y2=0
cc_623 N_A_608_74#_c_697_n N_A_2004_136#_c_1320_n 0.00627556f $X=10.41 $Y=0.405
+ $X2=0 $Y2=0
cc_624 N_A_608_74#_c_698_n N_A_2004_136#_c_1320_n 4.72354e-19 $X=10.41 $Y=0.405
+ $X2=0 $Y2=0
cc_625 N_A_608_74#_c_697_n N_A_2004_136#_c_1322_n 0.0151563f $X=10.41 $Y=0.405
+ $X2=0 $Y2=0
cc_626 N_A_608_74#_c_698_n N_A_2004_136#_c_1322_n 0.00132987f $X=10.41 $Y=0.405
+ $X2=0 $Y2=0
cc_627 N_A_608_74#_c_688_n N_A_2004_136#_c_1336_n 0.00910172f $X=10.205 $Y=1.545
+ $X2=0 $Y2=0
cc_628 N_A_608_74#_c_697_n N_A_2004_136#_c_1336_n 0.038646f $X=10.41 $Y=0.405
+ $X2=0 $Y2=0
cc_629 N_A_608_74#_c_698_n N_A_2004_136#_c_1336_n 0.011627f $X=10.41 $Y=0.405
+ $X2=0 $Y2=0
cc_630 N_A_608_74#_c_742_n N_VPWR_M1007_d 0.00812992f $X=6.15 $Y=2.475 $X2=0
+ $Y2=0
cc_631 N_A_608_74#_c_718_n N_VPWR_M1004_d 0.00953714f $X=8.63 $Y=2.905 $X2=0
+ $Y2=0
cc_632 N_A_608_74#_c_709_n N_VPWR_c_1402_n 0.00814477f $X=4.875 $Y=2.99 $X2=0
+ $Y2=0
cc_633 N_A_608_74#_c_741_n N_VPWR_c_1402_n 0.00728136f $X=4.96 $Y=2.905 $X2=0
+ $Y2=0
cc_634 N_A_608_74#_c_742_n N_VPWR_c_1402_n 0.0236929f $X=6.15 $Y=2.475 $X2=0
+ $Y2=0
cc_635 N_A_608_74#_c_712_n N_VPWR_c_1402_n 0.00817223f $X=6.4 $Y=2.905 $X2=0
+ $Y2=0
cc_636 N_A_608_74#_c_715_n N_VPWR_c_1402_n 0.00856798f $X=6.65 $Y=2.99 $X2=0
+ $Y2=0
cc_637 N_A_608_74#_c_717_n N_VPWR_c_1403_n 0.0142846f $X=8.545 $Y=2.99 $X2=0
+ $Y2=0
cc_638 N_A_608_74#_c_718_n N_VPWR_c_1403_n 0.0657339f $X=8.63 $Y=2.905 $X2=0
+ $Y2=0
cc_639 N_A_608_74#_c_693_n N_VPWR_c_1403_n 0.0110646f $X=9.215 $Y=1.74 $X2=0
+ $Y2=0
cc_640 N_A_608_74#_c_685_n N_VPWR_c_1405_n 7.25171e-19 $X=6.495 $Y=1.925 $X2=0
+ $Y2=0
cc_641 N_A_608_74#_c_714_n N_VPWR_c_1405_n 0.0730565f $X=7.785 $Y=2.99 $X2=0
+ $Y2=0
cc_642 N_A_608_74#_c_715_n N_VPWR_c_1405_n 0.0358565f $X=6.65 $Y=2.99 $X2=0
+ $Y2=0
cc_643 N_A_608_74#_c_717_n N_VPWR_c_1405_n 0.0501353f $X=8.545 $Y=2.99 $X2=0
+ $Y2=0
cc_644 N_A_608_74#_c_722_n N_VPWR_c_1405_n 0.0121143f $X=7.87 $Y=2.99 $X2=0
+ $Y2=0
cc_645 N_A_608_74#_c_709_n N_VPWR_c_1408_n 0.0500304f $X=4.875 $Y=2.99 $X2=0
+ $Y2=0
cc_646 N_A_608_74#_c_710_n N_VPWR_c_1408_n 0.0115566f $X=4.275 $Y=2.99 $X2=0
+ $Y2=0
cc_647 N_A_608_74#_c_709_n N_VPWR_c_1400_n 0.0264677f $X=4.875 $Y=2.99 $X2=0
+ $Y2=0
cc_648 N_A_608_74#_c_710_n N_VPWR_c_1400_n 0.00579705f $X=4.275 $Y=2.99 $X2=0
+ $Y2=0
cc_649 N_A_608_74#_c_742_n N_VPWR_c_1400_n 0.0271957f $X=6.15 $Y=2.475 $X2=0
+ $Y2=0
cc_650 N_A_608_74#_c_714_n N_VPWR_c_1400_n 0.0426655f $X=7.785 $Y=2.99 $X2=0
+ $Y2=0
cc_651 N_A_608_74#_c_715_n N_VPWR_c_1400_n 0.0194413f $X=6.65 $Y=2.99 $X2=0
+ $Y2=0
cc_652 N_A_608_74#_c_717_n N_VPWR_c_1400_n 0.0287839f $X=8.545 $Y=2.99 $X2=0
+ $Y2=0
cc_653 N_A_608_74#_c_722_n N_VPWR_c_1400_n 0.00659864f $X=7.87 $Y=2.99 $X2=0
+ $Y2=0
cc_654 N_A_608_74#_c_705_n N_A_256_368#_c_1508_n 0.033874f $X=3.35 $Y=2.57 $X2=0
+ $Y2=0
cc_655 N_A_608_74#_c_705_n N_A_256_368#_c_1516_n 0.0121155f $X=3.35 $Y=2.57
+ $X2=0 $Y2=0
cc_656 N_A_608_74#_M1006_d N_A_256_368#_c_1534_n 0.00562291f $X=3.04 $Y=0.37
+ $X2=0 $Y2=0
cc_657 N_A_608_74#_c_691_n N_A_256_368#_c_1534_n 0.0236057f $X=3.43 $Y=0.76
+ $X2=0 $Y2=0
cc_658 N_A_608_74#_M1006_d N_A_256_368#_c_1499_n 0.00455896f $X=3.04 $Y=0.37
+ $X2=0 $Y2=0
cc_659 N_A_608_74#_c_691_n N_A_256_368#_c_1499_n 0.0129709f $X=3.43 $Y=0.76
+ $X2=0 $Y2=0
cc_660 N_A_608_74#_c_691_n N_A_256_368#_c_1503_n 0.0322273f $X=3.43 $Y=0.76
+ $X2=0 $Y2=0
cc_661 N_A_608_74#_c_720_n N_A_256_368#_c_1503_n 0.0114639f $X=3.35 $Y=2.04
+ $X2=0 $Y2=0
cc_662 N_A_608_74#_M1006_d N_A_256_368#_c_1504_n 0.00105058f $X=3.04 $Y=0.37
+ $X2=0 $Y2=0
cc_663 N_A_608_74#_c_691_n N_A_256_368#_c_1504_n 0.0131266f $X=3.43 $Y=0.76
+ $X2=0 $Y2=0
cc_664 N_A_608_74#_c_742_n N_A_1197_368#_M1012_d 0.00308816f $X=6.15 $Y=2.475
+ $X2=0 $Y2=0
cc_665 N_A_608_74#_c_712_n N_A_1197_368#_M1012_d 0.00479816f $X=6.4 $Y=2.905
+ $X2=0 $Y2=0
cc_666 N_A_608_74#_c_801_p N_A_1197_368#_M1012_d 0.0032922f $X=6.4 $Y=2.475
+ $X2=0 $Y2=0
cc_667 N_A_608_74#_c_685_n N_A_1197_368#_c_1596_n 0.00224436f $X=6.495 $Y=1.925
+ $X2=0 $Y2=0
cc_668 N_A_608_74#_c_742_n N_A_1197_368#_c_1596_n 0.00877893f $X=6.15 $Y=2.475
+ $X2=0 $Y2=0
cc_669 N_A_608_74#_c_713_n N_A_1197_368#_c_1596_n 0.0258596f $X=6.565 $Y=2.39
+ $X2=0 $Y2=0
cc_670 N_A_608_74#_c_801_p N_A_1197_368#_c_1596_n 0.013336f $X=6.4 $Y=2.475
+ $X2=0 $Y2=0
cc_671 N_A_608_74#_c_685_n N_A_1197_368#_c_1594_n 0.0035823f $X=6.495 $Y=1.925
+ $X2=0 $Y2=0
cc_672 N_A_608_74#_c_699_n N_A_1197_368#_c_1594_n 0.0258596f $X=6.605 $Y=1.675
+ $X2=0 $Y2=0
cc_673 N_A_608_74#_c_685_n N_A_1197_368#_c_1595_n 0.00152634f $X=6.495 $Y=1.925
+ $X2=0 $Y2=0
cc_674 N_A_608_74#_c_712_n N_COUT_M1030_d 0.00874807f $X=6.4 $Y=2.905 $X2=0
+ $Y2=0
cc_675 N_A_608_74#_c_713_n N_COUT_M1030_d 0.00419945f $X=6.565 $Y=2.39 $X2=0
+ $Y2=0
cc_676 N_A_608_74#_c_801_p N_COUT_M1030_d 0.00188126f $X=6.4 $Y=2.475 $X2=0
+ $Y2=0
cc_677 N_A_608_74#_c_685_n N_COUT_c_1630_n 0.00767841f $X=6.495 $Y=1.925 $X2=0
+ $Y2=0
cc_678 N_A_608_74#_c_712_n N_COUT_c_1630_n 0.00916949f $X=6.4 $Y=2.905 $X2=0
+ $Y2=0
cc_679 N_A_608_74#_c_713_n N_COUT_c_1630_n 0.030697f $X=6.565 $Y=2.39 $X2=0
+ $Y2=0
cc_680 N_A_608_74#_c_714_n N_COUT_c_1630_n 0.0142433f $X=7.785 $Y=2.99 $X2=0
+ $Y2=0
cc_681 N_A_608_74#_c_801_p N_COUT_c_1630_n 0.0153274f $X=6.4 $Y=2.475 $X2=0
+ $Y2=0
cc_682 N_A_608_74#_c_699_n N_COUT_c_1630_n 0.0242846f $X=6.605 $Y=1.675 $X2=0
+ $Y2=0
cc_683 N_A_608_74#_c_714_n N_COUT_c_1643_n 0.029904f $X=7.785 $Y=2.99 $X2=0
+ $Y2=0
cc_684 N_A_608_74#_c_685_n N_COUT_c_1631_n 0.00145288f $X=6.495 $Y=1.925 $X2=0
+ $Y2=0
cc_685 N_A_608_74#_c_699_n N_COUT_c_1631_n 0.00663139f $X=6.605 $Y=1.675 $X2=0
+ $Y2=0
cc_686 N_A_608_74#_c_700_n N_COUT_c_1631_n 3.58087e-19 $X=7.91 $Y=1.32 $X2=0
+ $Y2=0
cc_687 N_A_608_74#_c_686_n COUT 0.00622306f $X=8.085 $Y=1.155 $X2=0 $Y2=0
cc_688 N_A_608_74#_c_700_n COUT 0.0215354f $X=7.91 $Y=1.32 $X2=0 $Y2=0
cc_689 N_A_608_74#_c_701_n COUT 0.00187528f $X=8.085 $Y=1.32 $X2=0 $Y2=0
cc_690 N_A_608_74#_c_692_n N_A_1595_400#_c_1680_n 0.0652283f $X=7.87 $Y=2.905
+ $X2=0 $Y2=0
cc_691 N_A_608_74#_c_718_n N_A_1595_400#_c_1680_n 0.0336618f $X=8.63 $Y=2.905
+ $X2=0 $Y2=0
cc_692 N_A_608_74#_c_701_n N_A_1595_400#_c_1680_n 0.00137994f $X=8.085 $Y=1.32
+ $X2=0 $Y2=0
cc_693 N_A_608_74#_c_717_n N_A_1595_400#_c_1685_n 0.018572f $X=8.545 $Y=2.99
+ $X2=0 $Y2=0
cc_694 N_A_608_74#_c_686_n N_A_1595_400#_c_1677_n 0.00457683f $X=8.085 $Y=1.155
+ $X2=0 $Y2=0
cc_695 N_A_608_74#_c_692_n N_A_1595_400#_c_1678_n 0.0188536f $X=7.87 $Y=2.905
+ $X2=0 $Y2=0
cc_696 N_A_608_74#_c_694_n N_A_1595_400#_c_1678_n 0.0135153f $X=8.715 $Y=1.74
+ $X2=0 $Y2=0
cc_697 N_A_608_74#_c_700_n N_A_1595_400#_c_1678_n 0.0245555f $X=7.91 $Y=1.32
+ $X2=0 $Y2=0
cc_698 N_A_608_74#_c_701_n N_A_1595_400#_c_1679_n 0.00457683f $X=8.085 $Y=1.32
+ $X2=0 $Y2=0
cc_699 N_A_608_74#_c_688_n N_A_1967_384#_c_1708_n 0.00641416f $X=10.205 $Y=1.545
+ $X2=0 $Y2=0
cc_700 N_A_608_74#_c_704_n N_A_1967_384#_c_1708_n 0.00681556f $X=10.205 $Y=1.845
+ $X2=0 $Y2=0
cc_701 N_A_608_74#_c_704_n N_A_1967_384#_c_1709_n 0.00948109f $X=10.205 $Y=1.845
+ $X2=0 $Y2=0
cc_702 N_A_608_74#_c_695_n N_VGND_M1019_d 0.0112075f $X=9.3 $Y=1.655 $X2=0 $Y2=0
cc_703 N_A_608_74#_c_693_n N_VGND_c_1772_n 3.03849e-19 $X=9.215 $Y=1.74 $X2=0
+ $Y2=0
cc_704 N_A_608_74#_c_695_n N_VGND_c_1772_n 0.0317803f $X=9.3 $Y=1.655 $X2=0
+ $Y2=0
cc_705 N_A_608_74#_c_696_n N_VGND_c_1772_n 0.0279244f $X=9.385 $Y=0.412 $X2=0
+ $Y2=0
cc_706 N_A_608_74#_c_686_n N_VGND_c_1776_n 0.00527342f $X=8.085 $Y=1.155 $X2=0
+ $Y2=0
cc_707 N_A_608_74#_c_690_n N_VGND_c_1777_n 0.0122133f $X=10.02 $Y=0.405 $X2=0
+ $Y2=0
cc_708 N_A_608_74#_c_696_n N_VGND_c_1777_n 0.0121867f $X=9.385 $Y=0.412 $X2=0
+ $Y2=0
cc_709 N_A_608_74#_c_697_n N_VGND_c_1777_n 0.077768f $X=10.41 $Y=0.405 $X2=0
+ $Y2=0
cc_710 N_A_608_74#_c_686_n N_VGND_c_1779_n 0.00534666f $X=8.085 $Y=1.155 $X2=0
+ $Y2=0
cc_711 N_A_608_74#_c_690_n N_VGND_c_1779_n 0.0035565f $X=10.02 $Y=0.405 $X2=0
+ $Y2=0
cc_712 N_A_608_74#_c_696_n N_VGND_c_1779_n 0.00660921f $X=9.385 $Y=0.412 $X2=0
+ $Y2=0
cc_713 N_A_608_74#_c_697_n N_VGND_c_1779_n 0.0421017f $X=10.41 $Y=0.405 $X2=0
+ $Y2=0
cc_714 N_A_608_74#_c_698_n N_VGND_c_1779_n 0.0122913f $X=10.41 $Y=0.405 $X2=0
+ $Y2=0
cc_715 N_A_430_418#_c_960_n N_CIN_c_1167_n 0.00333256f $X=7.81 $Y=1.8 $X2=-0.19
+ $Y2=-0.245
cc_716 N_A_430_418#_c_962_n N_CIN_c_1167_n 0.0216342f $X=7.9 $Y=1.925 $X2=-0.19
+ $Y2=-0.245
cc_717 N_A_430_418#_c_971_n N_CIN_c_1167_n 0.0120122f $X=10.655 $Y=2.035
+ $X2=-0.19 $Y2=-0.245
cc_718 N_A_430_418#_c_971_n N_CIN_c_1168_n 0.00684381f $X=10.655 $Y=2.035 $X2=0
+ $Y2=0
cc_719 N_A_430_418#_c_971_n CIN 5.45617e-19 $X=10.655 $Y=2.035 $X2=0 $Y2=0
cc_720 N_A_430_418#_c_960_n N_CIN_c_1166_n 9.38476e-19 $X=7.81 $Y=1.8 $X2=0
+ $Y2=0
cc_721 N_A_430_418#_c_971_n N_CIN_c_1166_n 0.00426106f $X=10.655 $Y=2.035 $X2=0
+ $Y2=0
cc_722 N_A_430_418#_c_971_n N_A_1854_368#_M1010_d 0.00400551f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_723 N_A_430_418#_c_1077_p N_A_1854_368#_M1028_d 0.00143427f $X=10.8 $Y=2.035
+ $X2=0 $Y2=0
cc_724 N_A_430_418#_c_959_n N_A_1854_368#_M1028_d 0.00551227f $X=10.85 $Y=1.595
+ $X2=0 $Y2=0
cc_725 N_A_430_418#_c_954_n N_A_1854_368#_c_1222_n 0.0113071f $X=10.89 $Y=1.43
+ $X2=0 $Y2=0
cc_726 N_A_430_418#_c_971_n N_A_1854_368#_c_1232_n 0.0362344f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_727 N_A_430_418#_c_971_n N_A_1854_368#_c_1223_n 0.0107117f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_728 N_A_430_418#_c_953_n N_A_1854_368#_c_1234_n 0.00512165f $X=10.655
+ $Y=1.845 $X2=0 $Y2=0
cc_729 N_A_430_418#_c_953_n N_A_1854_368#_c_1235_n 0.00623135f $X=10.655
+ $Y=1.845 $X2=0 $Y2=0
cc_730 N_A_430_418#_c_953_n N_A_1854_368#_c_1225_n 0.00771364f $X=10.655
+ $Y=1.845 $X2=0 $Y2=0
cc_731 N_A_430_418#_c_971_n N_A_2004_136#_M1024_d 0.00275654f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_732 N_A_430_418#_c_953_n N_A_2004_136#_c_1319_n 0.00623663f $X=10.655
+ $Y=1.845 $X2=0 $Y2=0
cc_733 N_A_430_418#_c_954_n N_A_2004_136#_c_1319_n 0.00405893f $X=10.89 $Y=1.43
+ $X2=0 $Y2=0
cc_734 N_A_430_418#_c_971_n N_A_2004_136#_c_1319_n 0.0227639f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_735 N_A_430_418#_c_1077_p N_A_2004_136#_c_1319_n 0.00233425f $X=10.8 $Y=2.035
+ $X2=0 $Y2=0
cc_736 N_A_430_418#_c_959_n N_A_2004_136#_c_1319_n 0.0530268f $X=10.85 $Y=1.595
+ $X2=0 $Y2=0
cc_737 N_A_430_418#_c_954_n N_A_2004_136#_c_1320_n 0.00797711f $X=10.89 $Y=1.43
+ $X2=0 $Y2=0
cc_738 N_A_430_418#_c_954_n N_A_2004_136#_c_1321_n 0.00232018f $X=10.89 $Y=1.43
+ $X2=0 $Y2=0
cc_739 N_A_430_418#_c_953_n N_A_2004_136#_c_1336_n 0.00642036f $X=10.655
+ $Y=1.845 $X2=0 $Y2=0
cc_740 N_A_430_418#_c_954_n N_A_2004_136#_c_1336_n 0.00967195f $X=10.89 $Y=1.43
+ $X2=0 $Y2=0
cc_741 N_A_430_418#_c_959_n N_A_2004_136#_c_1336_n 0.016795f $X=10.85 $Y=1.595
+ $X2=0 $Y2=0
cc_742 N_A_430_418#_c_969_n N_VPWR_M1007_d 0.00412872f $X=7.295 $Y=2.035 $X2=0
+ $Y2=0
cc_743 N_A_430_418#_c_971_n N_VPWR_M1004_d 0.0121108f $X=10.655 $Y=2.035 $X2=0
+ $Y2=0
cc_744 N_A_430_418#_c_971_n N_VPWR_c_1403_n 0.0137038f $X=10.655 $Y=2.035 $X2=0
+ $Y2=0
cc_745 N_A_430_418#_c_962_n N_VPWR_c_1405_n 7.43378e-19 $X=7.9 $Y=1.925 $X2=0
+ $Y2=0
cc_746 N_A_430_418#_c_967_n N_A_256_368#_M1011_d 3.14661e-19 $X=4.415 $Y=2.035
+ $X2=0 $Y2=0
cc_747 N_A_430_418#_M1011_s N_A_256_368#_c_1506_n 0.00682932f $X=2.15 $Y=2.09
+ $X2=0 $Y2=0
cc_748 N_A_430_418#_c_967_n N_A_256_368#_c_1506_n 0.0055145f $X=4.415 $Y=2.035
+ $X2=0 $Y2=0
cc_749 N_A_430_418#_c_968_n N_A_256_368#_c_1506_n 0.00227498f $X=2.305 $Y=2.035
+ $X2=0 $Y2=0
cc_750 N_A_430_418#_c_973_n N_A_256_368#_c_1506_n 0.02983f $X=2.16 $Y=2.035
+ $X2=0 $Y2=0
cc_751 N_A_430_418#_c_967_n N_A_256_368#_c_1508_n 0.0242931f $X=4.415 $Y=2.035
+ $X2=0 $Y2=0
cc_752 N_A_430_418#_c_968_n N_A_256_368#_c_1508_n 2.34713e-19 $X=2.305 $Y=2.035
+ $X2=0 $Y2=0
cc_753 N_A_430_418#_c_973_n N_A_256_368#_c_1508_n 0.0148549f $X=2.16 $Y=2.035
+ $X2=0 $Y2=0
cc_754 N_A_430_418#_c_968_n N_A_256_368#_c_1509_n 0.0074703f $X=2.305 $Y=2.035
+ $X2=0 $Y2=0
cc_755 N_A_430_418#_c_973_n N_A_256_368#_c_1509_n 0.0341781f $X=2.16 $Y=2.035
+ $X2=0 $Y2=0
cc_756 N_A_430_418#_c_955_n N_A_256_368#_c_1501_n 0.0436429f $X=2.32 $Y=0.78
+ $X2=0 $Y2=0
cc_757 N_A_430_418#_c_955_n N_A_256_368#_c_1502_n 0.0209605f $X=2.32 $Y=0.78
+ $X2=0 $Y2=0
cc_758 N_A_430_418#_c_955_n N_A_256_368#_c_1503_n 0.0334038f $X=2.32 $Y=0.78
+ $X2=0 $Y2=0
cc_759 N_A_430_418#_c_967_n N_A_256_368#_c_1503_n 0.00835823f $X=4.415 $Y=2.035
+ $X2=0 $Y2=0
cc_760 N_A_430_418#_c_968_n N_A_256_368#_c_1503_n 2.54236e-19 $X=2.305 $Y=2.035
+ $X2=0 $Y2=0
cc_761 N_A_430_418#_c_973_n N_A_256_368#_c_1503_n 0.00546571f $X=2.16 $Y=2.035
+ $X2=0 $Y2=0
cc_762 N_A_430_418#_c_955_n N_A_256_368#_c_1504_n 0.00554772f $X=2.32 $Y=0.78
+ $X2=0 $Y2=0
cc_763 N_A_430_418#_c_969_n N_A_1197_368#_M1012_d 0.00100298f $X=7.295 $Y=2.035
+ $X2=0 $Y2=0
cc_764 N_A_430_418#_c_950_n N_A_1197_368#_c_1593_n 0.00774505f $X=6.52 $Y=1.12
+ $X2=0 $Y2=0
cc_765 N_A_430_418#_c_969_n N_A_1197_368#_c_1596_n 0.026791f $X=7.295 $Y=2.035
+ $X2=0 $Y2=0
cc_766 N_A_430_418#_c_950_n N_A_1197_368#_c_1594_n 0.00183123f $X=6.52 $Y=1.12
+ $X2=0 $Y2=0
cc_767 N_A_430_418#_c_950_n N_A_1197_368#_c_1595_n 0.00242694f $X=6.52 $Y=1.12
+ $X2=0 $Y2=0
cc_768 N_A_430_418#_c_969_n N_COUT_M1030_d 0.0088082f $X=7.295 $Y=2.035 $X2=0
+ $Y2=0
cc_769 N_A_430_418#_c_971_n N_COUT_M1030_d 0.00678598f $X=10.655 $Y=2.035 $X2=0
+ $Y2=0
cc_770 N_A_430_418#_c_972_n N_COUT_M1030_d 0.00283248f $X=7.585 $Y=2.035 $X2=0
+ $Y2=0
cc_771 N_A_430_418#_c_958_n N_COUT_M1030_d 0.00550281f $X=7.37 $Y=1.335 $X2=0
+ $Y2=0
cc_772 N_A_430_418#_c_961_n N_COUT_c_1630_n 0.00450777f $X=7.535 $Y=1.8 $X2=0
+ $Y2=0
cc_773 N_A_430_418#_c_969_n N_COUT_c_1630_n 0.0274935f $X=7.295 $Y=2.035 $X2=0
+ $Y2=0
cc_774 N_A_430_418#_c_972_n N_COUT_c_1630_n 5.86129e-19 $X=7.585 $Y=2.035 $X2=0
+ $Y2=0
cc_775 N_A_430_418#_c_960_n N_COUT_c_1643_n 0.00166755f $X=7.81 $Y=1.8 $X2=0
+ $Y2=0
cc_776 N_A_430_418#_c_961_n N_COUT_c_1643_n 0.00242951f $X=7.535 $Y=1.8 $X2=0
+ $Y2=0
cc_777 N_A_430_418#_c_962_n N_COUT_c_1643_n 0.00236219f $X=7.9 $Y=1.925 $X2=0
+ $Y2=0
cc_778 N_A_430_418#_c_969_n N_COUT_c_1643_n 0.0081924f $X=7.295 $Y=2.035 $X2=0
+ $Y2=0
cc_779 N_A_430_418#_c_971_n N_COUT_c_1643_n 0.0013529f $X=10.655 $Y=2.035 $X2=0
+ $Y2=0
cc_780 N_A_430_418#_c_972_n N_COUT_c_1643_n 0.00361926f $X=7.585 $Y=2.035 $X2=0
+ $Y2=0
cc_781 N_A_430_418#_c_958_n N_COUT_c_1643_n 0.0201052f $X=7.37 $Y=1.335 $X2=0
+ $Y2=0
cc_782 N_A_430_418#_c_950_n N_COUT_c_1631_n 0.0135652f $X=6.52 $Y=1.12 $X2=0
+ $Y2=0
cc_783 N_A_430_418#_c_951_n N_COUT_c_1631_n 0.0279512f $X=7.205 $Y=1.195 $X2=0
+ $Y2=0
cc_784 N_A_430_418#_c_957_n N_COUT_c_1631_n 0.00450777f $X=7.37 $Y=1.335 $X2=0
+ $Y2=0
cc_785 N_A_430_418#_c_958_n N_COUT_c_1631_n 0.0728001f $X=7.37 $Y=1.335 $X2=0
+ $Y2=0
cc_786 N_A_430_418#_c_951_n COUT 0.0156322f $X=7.205 $Y=1.195 $X2=0 $Y2=0
cc_787 N_A_430_418#_c_958_n COUT 0.0251574f $X=7.37 $Y=1.335 $X2=0 $Y2=0
cc_788 N_A_430_418#_c_971_n N_A_1595_400#_M1026_d 0.00943568f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_789 N_A_430_418#_c_960_n N_A_1595_400#_c_1680_n 9.41618e-19 $X=7.81 $Y=1.8
+ $X2=0 $Y2=0
cc_790 N_A_430_418#_c_962_n N_A_1595_400#_c_1680_n 0.00595274f $X=7.9 $Y=1.925
+ $X2=0 $Y2=0
cc_791 N_A_430_418#_c_971_n N_A_1595_400#_c_1685_n 0.0317546f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_792 N_A_430_418#_c_960_n N_A_1595_400#_c_1678_n 8.6017e-19 $X=7.81 $Y=1.8
+ $X2=0 $Y2=0
cc_793 N_A_430_418#_c_971_n N_A_1967_384#_M1024_s 0.00576515f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_794 N_A_430_418#_c_971_n N_A_1967_384#_c_1708_n 0.0182448f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_795 N_A_430_418#_c_953_n N_A_1967_384#_c_1709_n 0.017922f $X=10.655 $Y=1.845
+ $X2=0 $Y2=0
cc_796 N_A_430_418#_c_971_n N_A_1967_384#_c_1709_n 0.0134585f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_797 N_A_430_418#_c_1077_p N_A_1967_384#_c_1709_n 0.0029808f $X=10.8 $Y=2.035
+ $X2=0 $Y2=0
cc_798 N_A_430_418#_c_959_n N_A_1967_384#_c_1709_n 0.0135704f $X=10.85 $Y=1.595
+ $X2=0 $Y2=0
cc_799 N_A_430_418#_c_954_n N_A_1967_384#_c_1706_n 0.00321553f $X=10.89 $Y=1.43
+ $X2=0 $Y2=0
cc_800 N_A_430_418#_c_954_n N_A_1967_384#_c_1723_n 0.00157686f $X=10.89 $Y=1.43
+ $X2=0 $Y2=0
cc_801 N_A_430_418#_c_953_n N_A_1967_384#_c_1710_n 0.00703602f $X=10.655
+ $Y=1.845 $X2=0 $Y2=0
cc_802 N_A_430_418#_c_1077_p N_A_1967_384#_c_1711_n 0.00153221f $X=10.8 $Y=2.035
+ $X2=0 $Y2=0
cc_803 N_A_430_418#_c_953_n N_A_1967_384#_c_1707_n 0.00439319f $X=10.655
+ $Y=1.845 $X2=0 $Y2=0
cc_804 N_A_430_418#_c_954_n N_A_1967_384#_c_1707_n 0.00357212f $X=10.89 $Y=1.43
+ $X2=0 $Y2=0
cc_805 N_A_430_418#_c_959_n N_A_1967_384#_c_1707_n 0.0530346f $X=10.85 $Y=1.595
+ $X2=0 $Y2=0
cc_806 N_A_430_418#_c_950_n N_VGND_c_1776_n 0.00527282f $X=6.52 $Y=1.12 $X2=0
+ $Y2=0
cc_807 N_A_430_418#_c_954_n N_VGND_c_1777_n 4.16716e-19 $X=10.89 $Y=1.43 $X2=0
+ $Y2=0
cc_808 N_A_430_418#_c_950_n N_VGND_c_1779_n 0.00534666f $X=6.52 $Y=1.12 $X2=0
+ $Y2=0
cc_809 N_CIN_c_1168_n N_A_1854_368#_c_1228_n 0.00706911f $X=9.195 $Y=1.765 $X2=0
+ $Y2=0
cc_810 N_CIN_c_1168_n N_A_1854_368#_c_1229_n 0.0046492f $X=9.195 $Y=1.765 $X2=0
+ $Y2=0
cc_811 N_CIN_c_1168_n N_A_1854_368#_c_1232_n 0.0021506f $X=9.195 $Y=1.765 $X2=0
+ $Y2=0
cc_812 N_CIN_c_1166_n N_A_1854_368#_c_1232_n 0.00489441f $X=9.195 $Y=1.46 $X2=0
+ $Y2=0
cc_813 N_CIN_c_1168_n N_A_1854_368#_c_1223_n 0.0036824f $X=9.195 $Y=1.765 $X2=0
+ $Y2=0
cc_814 N_CIN_c_1166_n N_A_1854_368#_c_1223_n 0.00232812f $X=9.195 $Y=1.46 $X2=0
+ $Y2=0
cc_815 N_CIN_c_1164_n N_A_1854_368#_c_1224_n 0.00110516f $X=9.47 $Y=1.395 $X2=0
+ $Y2=0
cc_816 N_CIN_c_1167_n N_VPWR_c_1403_n 0.00257417f $X=8.49 $Y=1.765 $X2=0 $Y2=0
cc_817 N_CIN_c_1168_n N_VPWR_c_1403_n 0.00789327f $X=9.195 $Y=1.765 $X2=0 $Y2=0
cc_818 N_CIN_c_1167_n N_VPWR_c_1405_n 7.44166e-19 $X=8.49 $Y=1.765 $X2=0 $Y2=0
cc_819 N_CIN_c_1168_n N_VPWR_c_1409_n 0.0044313f $X=9.195 $Y=1.765 $X2=0 $Y2=0
cc_820 N_CIN_c_1168_n N_VPWR_c_1400_n 0.00862964f $X=9.195 $Y=1.765 $X2=0 $Y2=0
cc_821 N_CIN_c_1163_n N_A_1595_400#_c_1677_n 0.00596212f $X=8.585 $Y=1.155 $X2=0
+ $Y2=0
cc_822 N_CIN_c_1167_n N_A_1595_400#_c_1678_n 0.00642478f $X=8.49 $Y=1.765 $X2=0
+ $Y2=0
cc_823 N_CIN_c_1163_n N_A_1595_400#_c_1678_n 0.00199024f $X=8.585 $Y=1.155 $X2=0
+ $Y2=0
cc_824 CIN N_A_1595_400#_c_1678_n 0.0151014f $X=8.795 $Y=1.21 $X2=0 $Y2=0
cc_825 N_CIN_c_1166_n N_A_1595_400#_c_1678_n 0.0130167f $X=9.195 $Y=1.46 $X2=0
+ $Y2=0
cc_826 N_CIN_c_1163_n N_A_1595_400#_c_1679_n 0.00584862f $X=8.585 $Y=1.155 $X2=0
+ $Y2=0
cc_827 N_CIN_c_1166_n N_A_1595_400#_c_1679_n 0.00575403f $X=9.195 $Y=1.46 $X2=0
+ $Y2=0
cc_828 N_CIN_c_1163_n N_VGND_c_1772_n 0.0163781f $X=8.585 $Y=1.155 $X2=0 $Y2=0
cc_829 N_CIN_c_1164_n N_VGND_c_1772_n 0.00135766f $X=9.47 $Y=1.395 $X2=0 $Y2=0
cc_830 CIN N_VGND_c_1772_n 0.0267264f $X=8.795 $Y=1.21 $X2=0 $Y2=0
cc_831 N_CIN_c_1166_n N_VGND_c_1772_n 0.0025546f $X=9.195 $Y=1.46 $X2=0 $Y2=0
cc_832 N_CIN_c_1163_n N_VGND_c_1776_n 0.00527282f $X=8.585 $Y=1.155 $X2=0 $Y2=0
cc_833 N_CIN_c_1164_n N_VGND_c_1777_n 5.88756e-19 $X=9.47 $Y=1.395 $X2=0 $Y2=0
cc_834 N_CIN_c_1163_n N_VGND_c_1779_n 0.00534666f $X=8.585 $Y=1.155 $X2=0 $Y2=0
cc_835 N_A_1854_368#_c_1227_n N_A_2004_136#_c_1317_n 0.0112607f $X=11.775
+ $Y=1.765 $X2=0 $Y2=0
cc_836 N_A_1854_368#_c_1230_n N_A_2004_136#_c_1317_n 6.31855e-19 $X=11.805
+ $Y=2.99 $X2=0 $Y2=0
cc_837 N_A_1854_368#_c_1231_n N_A_2004_136#_c_1317_n 0.00287306f $X=11.89
+ $Y=2.905 $X2=0 $Y2=0
cc_838 N_A_1854_368#_c_1225_n N_A_2004_136#_c_1317_n 0.0179413f $X=11.7 $Y=1.515
+ $X2=0 $Y2=0
cc_839 N_A_1854_368#_c_1226_n N_A_2004_136#_c_1317_n 0.00228376f $X=11.89
+ $Y=1.515 $X2=0 $Y2=0
cc_840 N_A_1854_368#_c_1223_n N_A_2004_136#_c_1319_n 0.0173801f $X=9.49 $Y=1.995
+ $X2=0 $Y2=0
cc_841 N_A_1854_368#_c_1224_n N_A_2004_136#_c_1319_n 0.00330702f $X=9.72 $Y=1.34
+ $X2=0 $Y2=0
cc_842 N_A_1854_368#_c_1222_n N_A_2004_136#_c_1320_n 0.0012124f $X=11.465
+ $Y=1.35 $X2=0 $Y2=0
cc_843 N_A_1854_368#_c_1222_n N_A_2004_136#_c_1321_n 0.00957183f $X=11.465
+ $Y=1.35 $X2=0 $Y2=0
cc_844 N_A_1854_368#_c_1222_n N_A_2004_136#_c_1323_n 0.0110418f $X=11.465
+ $Y=1.35 $X2=0 $Y2=0
cc_845 N_A_1854_368#_c_1225_n N_A_2004_136#_c_1360_n 0.00285464f $X=11.7
+ $Y=1.515 $X2=0 $Y2=0
cc_846 N_A_1854_368#_c_1226_n N_A_2004_136#_c_1360_n 0.0166605f $X=11.89
+ $Y=1.515 $X2=0 $Y2=0
cc_847 N_A_1854_368#_c_1225_n N_A_2004_136#_c_1362_n 0.00415388f $X=11.7
+ $Y=1.515 $X2=0 $Y2=0
cc_848 N_A_1854_368#_c_1226_n N_A_2004_136#_c_1362_n 0.0134553f $X=11.89
+ $Y=1.515 $X2=0 $Y2=0
cc_849 N_A_1854_368#_c_1222_n N_A_2004_136#_c_1324_n 0.00391168f $X=11.465
+ $Y=1.35 $X2=0 $Y2=0
cc_850 N_A_1854_368#_c_1225_n N_A_2004_136#_c_1324_n 3.25592e-19 $X=11.7
+ $Y=1.515 $X2=0 $Y2=0
cc_851 N_A_1854_368#_c_1226_n N_A_2004_136#_c_1324_n 0.0263839f $X=11.89
+ $Y=1.515 $X2=0 $Y2=0
cc_852 N_A_1854_368#_c_1231_n N_VPWR_M1013_d 0.0092342f $X=11.89 $Y=2.905 $X2=0
+ $Y2=0
cc_853 N_A_1854_368#_c_1229_n N_VPWR_c_1403_n 0.0119328f $X=9.725 $Y=2.99 $X2=0
+ $Y2=0
cc_854 N_A_1854_368#_c_1232_n N_VPWR_c_1403_n 0.0597126f $X=9.42 $Y=2.08 $X2=0
+ $Y2=0
cc_855 N_A_1854_368#_c_1227_n N_VPWR_c_1404_n 0.00332849f $X=11.775 $Y=1.765
+ $X2=0 $Y2=0
cc_856 N_A_1854_368#_c_1230_n N_VPWR_c_1404_n 0.0146661f $X=11.805 $Y=2.99 $X2=0
+ $Y2=0
cc_857 N_A_1854_368#_c_1231_n N_VPWR_c_1404_n 0.0789548f $X=11.89 $Y=2.905 $X2=0
+ $Y2=0
cc_858 N_A_1854_368#_c_1227_n N_VPWR_c_1409_n 7.43987e-19 $X=11.775 $Y=1.765
+ $X2=0 $Y2=0
cc_859 N_A_1854_368#_c_1229_n N_VPWR_c_1409_n 0.0336038f $X=9.725 $Y=2.99 $X2=0
+ $Y2=0
cc_860 N_A_1854_368#_c_1230_n N_VPWR_c_1409_n 0.0121867f $X=11.805 $Y=2.99 $X2=0
+ $Y2=0
cc_861 N_A_1854_368#_c_1234_n N_VPWR_c_1409_n 0.134995f $X=10.8 $Y=2.907 $X2=0
+ $Y2=0
cc_862 N_A_1854_368#_c_1229_n N_VPWR_c_1400_n 0.0181986f $X=9.725 $Y=2.99 $X2=0
+ $Y2=0
cc_863 N_A_1854_368#_c_1230_n N_VPWR_c_1400_n 0.00660921f $X=11.805 $Y=2.99
+ $X2=0 $Y2=0
cc_864 N_A_1854_368#_c_1234_n N_VPWR_c_1400_n 0.0783914f $X=10.8 $Y=2.907 $X2=0
+ $Y2=0
cc_865 N_A_1854_368#_c_1228_n N_A_1967_384#_c_1729_n 0.0284333f $X=9.42 $Y=2.815
+ $X2=0 $Y2=0
cc_866 N_A_1854_368#_c_1234_n N_A_1967_384#_c_1729_n 0.0130862f $X=10.8 $Y=2.907
+ $X2=0 $Y2=0
cc_867 N_A_1854_368#_c_1223_n N_A_1967_384#_c_1708_n 0.0382752f $X=9.49 $Y=1.995
+ $X2=0 $Y2=0
cc_868 N_A_1854_368#_M1028_d N_A_1967_384#_c_1709_n 0.0128589f $X=10.73 $Y=1.92
+ $X2=0 $Y2=0
cc_869 N_A_1854_368#_c_1230_n N_A_1967_384#_c_1709_n 0.0296055f $X=11.805
+ $Y=2.99 $X2=0 $Y2=0
cc_870 N_A_1854_368#_c_1231_n N_A_1967_384#_c_1709_n 0.0254201f $X=11.89
+ $Y=2.905 $X2=0 $Y2=0
cc_871 N_A_1854_368#_c_1234_n N_A_1967_384#_c_1709_n 0.0250603f $X=10.8 $Y=2.907
+ $X2=0 $Y2=0
cc_872 N_A_1854_368#_c_1235_n N_A_1967_384#_c_1709_n 0.0260578f $X=11.155
+ $Y=2.907 $X2=0 $Y2=0
cc_873 N_A_1854_368#_c_1222_n N_A_1967_384#_c_1706_n 0.00452331f $X=11.465
+ $Y=1.35 $X2=0 $Y2=0
cc_874 N_A_1854_368#_c_1222_n N_A_1967_384#_c_1723_n 0.00391079f $X=11.465
+ $Y=1.35 $X2=0 $Y2=0
cc_875 N_A_1854_368#_c_1227_n N_A_1967_384#_c_1711_n 0.00498109f $X=11.775
+ $Y=1.765 $X2=0 $Y2=0
cc_876 N_A_1854_368#_c_1231_n N_A_1967_384#_c_1711_n 0.0415787f $X=11.89
+ $Y=2.905 $X2=0 $Y2=0
cc_877 N_A_1854_368#_c_1225_n N_A_1967_384#_c_1711_n 0.00897356f $X=11.7
+ $Y=1.515 $X2=0 $Y2=0
cc_878 N_A_1854_368#_c_1226_n N_A_1967_384#_c_1711_n 0.00817548f $X=11.89
+ $Y=1.515 $X2=0 $Y2=0
cc_879 N_A_1854_368#_c_1222_n N_A_1967_384#_c_1707_n 0.00618787f $X=11.465
+ $Y=1.35 $X2=0 $Y2=0
cc_880 N_A_1854_368#_c_1227_n N_A_1967_384#_c_1707_n 0.00136495f $X=11.775
+ $Y=1.765 $X2=0 $Y2=0
cc_881 N_A_1854_368#_c_1231_n N_A_1967_384#_c_1707_n 0.00594434f $X=11.89
+ $Y=2.905 $X2=0 $Y2=0
cc_882 N_A_1854_368#_c_1225_n N_A_1967_384#_c_1707_n 8.45983e-19 $X=11.7
+ $Y=1.515 $X2=0 $Y2=0
cc_883 N_A_1854_368#_c_1226_n N_A_1967_384#_c_1707_n 0.0253231f $X=11.89
+ $Y=1.515 $X2=0 $Y2=0
cc_884 N_A_1854_368#_c_1231_n SUM 0.00526803f $X=11.89 $Y=2.905 $X2=0 $Y2=0
cc_885 N_A_1854_368#_c_1222_n N_VGND_c_1773_n 6.79189e-19 $X=11.465 $Y=1.35
+ $X2=0 $Y2=0
cc_886 N_A_1854_368#_c_1222_n N_VGND_c_1777_n 6.15596e-19 $X=11.465 $Y=1.35
+ $X2=0 $Y2=0
cc_887 N_A_2004_136#_c_1317_n N_VPWR_c_1404_n 0.0213474f $X=12.455 $Y=1.765
+ $X2=0 $Y2=0
cc_888 N_A_2004_136#_c_1324_n N_VPWR_c_1404_n 0.0190023f $X=12.285 $Y=1.515
+ $X2=0 $Y2=0
cc_889 N_A_2004_136#_c_1317_n N_VPWR_c_1410_n 0.00413917f $X=12.455 $Y=1.765
+ $X2=0 $Y2=0
cc_890 N_A_2004_136#_c_1317_n N_VPWR_c_1400_n 0.00821221f $X=12.455 $Y=1.765
+ $X2=0 $Y2=0
cc_891 N_A_2004_136#_c_1319_n N_A_1967_384#_c_1708_n 0.0197948f $X=10.43
+ $Y=2.065 $X2=0 $Y2=0
cc_892 N_A_2004_136#_M1024_d N_A_1967_384#_c_1709_n 0.00453512f $X=10.28 $Y=1.92
+ $X2=0 $Y2=0
cc_893 N_A_2004_136#_c_1319_n N_A_1967_384#_c_1709_n 0.0144706f $X=10.43
+ $Y=2.065 $X2=0 $Y2=0
cc_894 N_A_2004_136#_c_1320_n N_A_1967_384#_c_1706_n 0.00594961f $X=10.83
+ $Y=0.74 $X2=0 $Y2=0
cc_895 N_A_2004_136#_c_1321_n N_A_1967_384#_c_1706_n 0.0231392f $X=11.585
+ $Y=0.405 $X2=0 $Y2=0
cc_896 N_A_2004_136#_c_1336_n N_A_1967_384#_c_1706_n 0.0258345f $X=10.83 $Y=1
+ $X2=0 $Y2=0
cc_897 N_A_2004_136#_c_1336_n N_A_1967_384#_c_1723_n 0.0161207f $X=10.83 $Y=1
+ $X2=0 $Y2=0
cc_898 N_A_2004_136#_c_1336_n N_A_1967_384#_c_1707_n 4.55714e-19 $X=10.83 $Y=1
+ $X2=0 $Y2=0
cc_899 N_A_2004_136#_c_1318_n SUM 0.00782592f $X=12.465 $Y=1.35 $X2=0 $Y2=0
cc_900 N_A_2004_136#_c_1317_n SUM 0.018944f $X=12.455 $Y=1.765 $X2=0 $Y2=0
cc_901 N_A_2004_136#_c_1318_n SUM 0.00328088f $X=12.465 $Y=1.35 $X2=0 $Y2=0
cc_902 N_A_2004_136#_c_1324_n SUM 0.0357347f $X=12.285 $Y=1.515 $X2=0 $Y2=0
cc_903 N_A_2004_136#_c_1323_n N_VGND_M1001_d 0.00857919f $X=11.67 $Y=1.01 $X2=0
+ $Y2=0
cc_904 N_A_2004_136#_c_1360_n N_VGND_M1001_d 0.023077f $X=12.145 $Y=1.095 $X2=0
+ $Y2=0
cc_905 N_A_2004_136#_c_1362_n N_VGND_M1001_d 0.00277575f $X=11.755 $Y=1.095
+ $X2=0 $Y2=0
cc_906 N_A_2004_136#_c_1324_n N_VGND_M1001_d 0.00105494f $X=12.285 $Y=1.515
+ $X2=0 $Y2=0
cc_907 N_A_2004_136#_c_1317_n N_VGND_c_1773_n 8.18201e-19 $X=12.455 $Y=1.765
+ $X2=0 $Y2=0
cc_908 N_A_2004_136#_c_1318_n N_VGND_c_1773_n 0.0104405f $X=12.465 $Y=1.35 $X2=0
+ $Y2=0
cc_909 N_A_2004_136#_c_1321_n N_VGND_c_1773_n 0.0153023f $X=11.585 $Y=0.405
+ $X2=0 $Y2=0
cc_910 N_A_2004_136#_c_1323_n N_VGND_c_1773_n 0.02505f $X=11.67 $Y=1.01 $X2=0
+ $Y2=0
cc_911 N_A_2004_136#_c_1360_n N_VGND_c_1773_n 0.0307423f $X=12.145 $Y=1.095
+ $X2=0 $Y2=0
cc_912 N_A_2004_136#_c_1321_n N_VGND_c_1777_n 0.0392505f $X=11.585 $Y=0.405
+ $X2=0 $Y2=0
cc_913 N_A_2004_136#_c_1322_n N_VGND_c_1777_n 0.00832763f $X=10.915 $Y=0.405
+ $X2=0 $Y2=0
cc_914 N_A_2004_136#_c_1336_n N_VGND_c_1777_n 0.00259374f $X=10.83 $Y=1 $X2=0
+ $Y2=0
cc_915 N_A_2004_136#_c_1318_n N_VGND_c_1778_n 0.00466874f $X=12.465 $Y=1.35
+ $X2=0 $Y2=0
cc_916 N_A_2004_136#_c_1318_n N_VGND_c_1779_n 0.00505379f $X=12.465 $Y=1.35
+ $X2=0 $Y2=0
cc_917 N_A_2004_136#_c_1321_n N_VGND_c_1779_n 0.0305583f $X=11.585 $Y=0.405
+ $X2=0 $Y2=0
cc_918 N_A_2004_136#_c_1322_n N_VGND_c_1779_n 0.00629651f $X=10.915 $Y=0.405
+ $X2=0 $Y2=0
cc_919 N_A_2004_136#_c_1336_n N_VGND_c_1779_n 0.00575318f $X=10.83 $Y=1 $X2=0
+ $Y2=0
cc_920 N_VPWR_c_1404_n SUM 0.0742466f $X=12.23 $Y=2.015 $X2=0 $Y2=0
cc_921 N_VPWR_c_1410_n SUM 0.011066f $X=12.72 $Y=3.33 $X2=0 $Y2=0
cc_922 N_VPWR_c_1400_n SUM 0.00915947f $X=12.72 $Y=3.33 $X2=0 $Y2=0
cc_923 N_A_256_368#_c_1499_n N_VGND_c_1775_n 0.0504711f $X=3.695 $Y=0.34 $X2=0
+ $Y2=0
cc_924 N_A_256_368#_c_1517_n N_VGND_c_1775_n 0.0115381f $X=3.175 $Y=0.34 $X2=0
+ $Y2=0
cc_925 N_A_256_368#_c_1499_n N_VGND_c_1779_n 0.0260462f $X=3.695 $Y=0.34 $X2=0
+ $Y2=0
cc_926 N_A_256_368#_c_1517_n N_VGND_c_1779_n 0.00579326f $X=3.175 $Y=0.34 $X2=0
+ $Y2=0
cc_927 N_A_1197_368#_c_1594_n N_COUT_c_1630_n 0.00632803f $X=6.14 $Y=1.82 $X2=0
+ $Y2=0
cc_928 N_A_1197_368#_c_1593_n N_COUT_c_1631_n 0.0242367f $X=6.305 $Y=0.55 $X2=0
+ $Y2=0
cc_929 N_A_1197_368#_c_1594_n N_COUT_c_1631_n 0.0118325f $X=6.14 $Y=1.82 $X2=0
+ $Y2=0
cc_930 N_A_1197_368#_c_1593_n N_VGND_c_1771_n 0.0102236f $X=6.305 $Y=0.55 $X2=0
+ $Y2=0
cc_931 N_A_1197_368#_c_1593_n N_VGND_c_1776_n 0.0126924f $X=6.305 $Y=0.55 $X2=0
+ $Y2=0
cc_932 N_A_1197_368#_c_1593_n N_VGND_c_1779_n 0.0118128f $X=6.305 $Y=0.55 $X2=0
+ $Y2=0
cc_933 N_COUT_c_1631_n N_VGND_c_1776_n 0.013372f $X=6.805 $Y=0.56 $X2=0 $Y2=0
cc_934 COUT N_VGND_c_1776_n 0.029099f $X=7.835 $Y=0.47 $X2=0 $Y2=0
cc_935 N_COUT_c_1631_n N_VGND_c_1779_n 0.0149229f $X=6.805 $Y=0.56 $X2=0 $Y2=0
cc_936 COUT N_VGND_c_1779_n 0.0332939f $X=7.835 $Y=0.47 $X2=0 $Y2=0
cc_937 N_A_1595_400#_c_1677_n N_VGND_c_1772_n 0.02327f $X=8.37 $Y=0.55 $X2=0
+ $Y2=0
cc_938 N_A_1595_400#_c_1677_n N_VGND_c_1776_n 0.0127604f $X=8.37 $Y=0.55 $X2=0
+ $Y2=0
cc_939 N_A_1595_400#_c_1677_n N_VGND_c_1779_n 0.011834f $X=8.37 $Y=0.55 $X2=0
+ $Y2=0
cc_940 SUM N_VGND_c_1773_n 0.0164291f $X=12.635 $Y=0.47 $X2=0 $Y2=0
cc_941 SUM N_VGND_c_1778_n 0.010571f $X=12.635 $Y=0.47 $X2=0 $Y2=0
cc_942 SUM N_VGND_c_1779_n 0.0113586f $X=12.635 $Y=0.47 $X2=0 $Y2=0
