# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_hs__dlxtn_2
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_hs__dlxtn_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  7.200000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.208500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.300000 0.455000 1.780000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.638000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.260000 1.920000 6.635000 2.890000 ;
        RECT 6.320000 0.350000 6.585000 1.125000 ;
        RECT 6.415000 1.125000 6.585000 1.920000 ;
    END
  END Q
  PIN GATE_N
    ANTENNAGATEAREA  0.237000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.985000 1.450000 1.315000 1.780000 ;
    END
  END GATE_N
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 7.200000 0.085000 ;
        RECT 0.625000  0.085000 0.955000 0.410000 ;
        RECT 2.815000  0.085000 3.145000 1.055000 ;
        RECT 4.820000  0.085000 5.150000 0.975000 ;
        RECT 5.845000  0.085000 6.140000 1.125000 ;
        RECT 6.755000  0.085000 7.085000 1.130000 ;
      LAYER mcon ;
        RECT 0.155000 -0.085000 0.325000 0.085000 ;
        RECT 0.635000 -0.085000 0.805000 0.085000 ;
        RECT 1.115000 -0.085000 1.285000 0.085000 ;
        RECT 1.595000 -0.085000 1.765000 0.085000 ;
        RECT 2.075000 -0.085000 2.245000 0.085000 ;
        RECT 2.555000 -0.085000 2.725000 0.085000 ;
        RECT 3.035000 -0.085000 3.205000 0.085000 ;
        RECT 3.515000 -0.085000 3.685000 0.085000 ;
        RECT 3.995000 -0.085000 4.165000 0.085000 ;
        RECT 4.475000 -0.085000 4.645000 0.085000 ;
        RECT 4.955000 -0.085000 5.125000 0.085000 ;
        RECT 5.435000 -0.085000 5.605000 0.085000 ;
        RECT 5.915000 -0.085000 6.085000 0.085000 ;
        RECT 6.395000 -0.085000 6.565000 0.085000 ;
        RECT 6.875000 -0.085000 7.045000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.245000 7.200000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 3.245000 7.200000 3.415000 ;
        RECT 0.765000 2.290000 1.095000 3.245000 ;
        RECT 2.360000 2.780000 2.705000 3.245000 ;
        RECT 4.360000 2.625000 5.080000 3.245000 ;
        RECT 5.845000 1.820000 6.060000 3.245000 ;
        RECT 6.835000 1.820000 7.085000 3.245000 ;
      LAYER mcon ;
        RECT 0.155000 3.245000 0.325000 3.415000 ;
        RECT 0.635000 3.245000 0.805000 3.415000 ;
        RECT 1.115000 3.245000 1.285000 3.415000 ;
        RECT 1.595000 3.245000 1.765000 3.415000 ;
        RECT 2.075000 3.245000 2.245000 3.415000 ;
        RECT 2.555000 3.245000 2.725000 3.415000 ;
        RECT 3.035000 3.245000 3.205000 3.415000 ;
        RECT 3.515000 3.245000 3.685000 3.415000 ;
        RECT 3.995000 3.245000 4.165000 3.415000 ;
        RECT 4.475000 3.245000 4.645000 3.415000 ;
        RECT 4.955000 3.245000 5.125000 3.415000 ;
        RECT 5.435000 3.245000 5.605000 3.415000 ;
        RECT 5.915000 3.245000 6.085000 3.415000 ;
        RECT 6.395000 3.245000 6.565000 3.415000 ;
        RECT 6.875000 3.245000 7.045000 3.415000 ;
      LAYER met1 ;
        RECT 0.000000 3.085000 7.200000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.115000 0.580000 1.315000 0.750000 ;
      RECT 0.115000 0.750000 0.795000 1.130000 ;
      RECT 0.265000 1.950000 0.795000 2.120000 ;
      RECT 0.265000 2.120000 0.595000 2.980000 ;
      RECT 0.625000 1.130000 0.795000 1.950000 ;
      RECT 1.135000 0.920000 1.885000 1.170000 ;
      RECT 1.145000 0.255000 2.645000 0.425000 ;
      RECT 1.145000 0.425000 1.315000 0.580000 ;
      RECT 1.265000 2.100000 1.655000 2.440000 ;
      RECT 1.265000 2.440000 3.045000 2.610000 ;
      RECT 1.265000 2.610000 1.655000 2.980000 ;
      RECT 1.485000 0.760000 1.885000 0.920000 ;
      RECT 1.485000 1.170000 1.885000 1.770000 ;
      RECT 1.485000 1.770000 1.655000 2.100000 ;
      RECT 1.825000 1.940000 3.510000 1.970000 ;
      RECT 1.825000 1.970000 2.225000 2.270000 ;
      RECT 2.055000 0.595000 2.305000 1.800000 ;
      RECT 2.055000 1.800000 3.510000 1.940000 ;
      RECT 2.475000 0.425000 2.645000 1.300000 ;
      RECT 2.475000 1.300000 2.970000 1.630000 ;
      RECT 2.875000 2.610000 3.045000 2.905000 ;
      RECT 2.875000 2.905000 4.190000 3.075000 ;
      RECT 3.180000 1.470000 3.510000 1.800000 ;
      RECT 3.315000 0.255000 4.375000 0.585000 ;
      RECT 3.315000 0.585000 3.485000 1.470000 ;
      RECT 3.330000 2.140000 3.850000 2.735000 ;
      RECT 3.655000 0.805000 4.250000 1.055000 ;
      RECT 3.680000 1.055000 3.850000 2.140000 ;
      RECT 4.020000 1.485000 4.350000 1.815000 ;
      RECT 4.020000 1.815000 4.190000 2.905000 ;
      RECT 4.080000 1.055000 4.250000 1.145000 ;
      RECT 4.080000 1.145000 5.160000 1.295000 ;
      RECT 4.080000 1.295000 5.335000 1.315000 ;
      RECT 4.360000 2.025000 5.580000 2.355000 ;
      RECT 4.990000 1.315000 5.335000 1.625000 ;
      RECT 5.250000 1.795000 5.675000 1.965000 ;
      RECT 5.250000 1.965000 5.580000 2.025000 ;
      RECT 5.250000 2.355000 5.580000 2.955000 ;
      RECT 5.330000 0.355000 5.580000 0.955000 ;
      RECT 5.330000 0.955000 5.675000 1.125000 ;
      RECT 5.505000 1.125000 5.675000 1.295000 ;
      RECT 5.505000 1.295000 6.245000 1.625000 ;
      RECT 5.505000 1.625000 5.675000 1.795000 ;
  END
END sky130_fd_sc_hs__dlxtn_2
