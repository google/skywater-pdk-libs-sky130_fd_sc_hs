* File: sky130_fd_sc_hs__and3b_1.pxi.spice
* Created: Tue Sep  1 19:55:27 2020
* 
x_PM_SKY130_FD_SC_HS__AND3B_1%A_N N_A_N_M1008_g N_A_N_M1006_g N_A_N_c_69_n
+ N_A_N_c_70_n N_A_N_c_74_n N_A_N_c_75_n A_N A_N N_A_N_c_71_n N_A_N_c_72_n
+ PM_SKY130_FD_SC_HS__AND3B_1%A_N
x_PM_SKY130_FD_SC_HS__AND3B_1%A_114_74# N_A_114_74#_M1008_d N_A_114_74#_M1006_d
+ N_A_114_74#_c_99_n N_A_114_74#_c_100_n N_A_114_74#_c_101_n N_A_114_74#_M1004_g
+ N_A_114_74#_c_109_n N_A_114_74#_M1001_g N_A_114_74#_c_102_n
+ N_A_114_74#_c_103_n N_A_114_74#_c_110_n N_A_114_74#_c_104_n
+ N_A_114_74#_c_105_n N_A_114_74#_c_106_n N_A_114_74#_c_112_n
+ N_A_114_74#_c_107_n PM_SKY130_FD_SC_HS__AND3B_1%A_114_74#
x_PM_SKY130_FD_SC_HS__AND3B_1%B N_B_M1005_g N_B_c_168_n N_B_M1003_g B
+ N_B_c_170_n PM_SKY130_FD_SC_HS__AND3B_1%B
x_PM_SKY130_FD_SC_HS__AND3B_1%C N_C_M1009_g N_C_c_201_n N_C_M1000_g C
+ N_C_c_202_n PM_SKY130_FD_SC_HS__AND3B_1%C
x_PM_SKY130_FD_SC_HS__AND3B_1%A_266_94# N_A_266_94#_M1004_s N_A_266_94#_M1001_s
+ N_A_266_94#_M1003_d N_A_266_94#_c_228_n N_A_266_94#_M1007_g
+ N_A_266_94#_M1002_g N_A_266_94#_c_230_n N_A_266_94#_c_231_n
+ N_A_266_94#_c_232_n N_A_266_94#_c_250_n N_A_266_94#_c_233_n
+ N_A_266_94#_c_236_n N_A_266_94#_c_237_n PM_SKY130_FD_SC_HS__AND3B_1%A_266_94#
x_PM_SKY130_FD_SC_HS__AND3B_1%VPWR N_VPWR_M1006_s N_VPWR_M1001_d N_VPWR_M1000_d
+ N_VPWR_c_315_n N_VPWR_c_316_n N_VPWR_c_317_n N_VPWR_c_318_n N_VPWR_c_319_n
+ N_VPWR_c_320_n N_VPWR_c_321_n N_VPWR_c_322_n VPWR N_VPWR_c_323_n
+ N_VPWR_c_314_n PM_SKY130_FD_SC_HS__AND3B_1%VPWR
x_PM_SKY130_FD_SC_HS__AND3B_1%X N_X_M1002_d N_X_M1007_d N_X_c_359_n N_X_c_360_n
+ X X X X N_X_c_363_n N_X_c_361_n PM_SKY130_FD_SC_HS__AND3B_1%X
x_PM_SKY130_FD_SC_HS__AND3B_1%VGND N_VGND_M1008_s N_VGND_M1009_d N_VGND_c_382_n
+ N_VGND_c_383_n N_VGND_c_384_n VGND N_VGND_c_385_n N_VGND_c_386_n
+ N_VGND_c_387_n N_VGND_c_388_n PM_SKY130_FD_SC_HS__AND3B_1%VGND
cc_1 VNB N_A_N_M1008_g 0.0315936f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.645
cc_2 VNB N_A_N_c_69_n 0.0275245f $X=-0.19 $Y=-0.245 $X2=0.405 $Y2=1.615
cc_3 VNB N_A_N_c_70_n 0.0036645f $X=-0.19 $Y=-0.245 $X2=0.405 $Y2=1.78
cc_4 VNB N_A_N_c_71_n 0.0185743f $X=-0.19 $Y=-0.245 $X2=0.405 $Y2=1.275
cc_5 VNB N_A_N_c_72_n 0.0240162f $X=-0.19 $Y=-0.245 $X2=0.405 $Y2=1.275
cc_6 VNB N_A_114_74#_c_99_n 0.0344902f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=2.54
cc_7 VNB N_A_114_74#_c_100_n 0.0129028f $X=-0.19 $Y=-0.245 $X2=0.405 $Y2=1.615
cc_8 VNB N_A_114_74#_c_101_n 0.0161108f $X=-0.19 $Y=-0.245 $X2=0.405 $Y2=1.78
cc_9 VNB N_A_114_74#_c_102_n 0.010725f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_114_74#_c_103_n 0.00839405f $X=-0.19 $Y=-0.245 $X2=0.405 $Y2=1.275
cc_11 VNB N_A_114_74#_c_104_n 0.0205614f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_114_74#_c_105_n 0.00199474f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_114_74#_c_106_n 0.0493999f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_114_74#_c_107_n 9.31753e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_B_M1005_g 0.0236487f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.645
cc_16 VNB N_B_c_168_n 0.0258125f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.78
cc_17 VNB N_C_M1009_g 0.0263528f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.645
cc_18 VNB N_C_c_201_n 0.023975f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.78
cc_19 VNB N_C_c_202_n 0.00189186f $X=-0.19 $Y=-0.245 $X2=0.405 $Y2=1.615
cc_20 VNB N_A_266_94#_c_228_n 0.0358794f $X=-0.19 $Y=-0.245 $X2=0.405 $Y2=1.275
cc_21 VNB N_A_266_94#_M1002_g 0.0294556f $X=-0.19 $Y=-0.245 $X2=0.502 $Y2=2.045
cc_22 VNB N_A_266_94#_c_230_n 0.010932f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_266_94#_c_231_n 0.00257034f $X=-0.19 $Y=-0.245 $X2=0.405 $Y2=1.275
cc_24 VNB N_A_266_94#_c_232_n 0.0351178f $X=-0.19 $Y=-0.245 $X2=0.347 $Y2=1.295
cc_25 VNB N_A_266_94#_c_233_n 8.27411e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_VPWR_c_314_n 0.163682f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_X_c_359_n 0.0267746f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=2.54
cc_28 VNB N_X_c_360_n 0.0144258f $X=-0.19 $Y=-0.245 $X2=0.405 $Y2=1.78
cc_29 VNB N_X_c_361_n 0.0248166f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_382_n 0.0120272f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=2.045
cc_31 VNB N_VGND_c_383_n 0.0342445f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=2.54
cc_32 VNB N_VGND_c_384_n 0.0134281f $X=-0.19 $Y=-0.245 $X2=0.405 $Y2=1.78
cc_33 VNB N_VGND_c_385_n 0.0644827f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_34 VNB N_VGND_c_386_n 0.0191572f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_387_n 0.267554f $X=-0.19 $Y=-0.245 $X2=0.347 $Y2=1.295
cc_36 VNB N_VGND_c_388_n 0.0113485f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VPB N_A_N_c_70_n 0.0154589f $X=-0.19 $Y=1.66 $X2=0.405 $Y2=1.78
cc_38 VPB N_A_N_c_74_n 0.0135533f $X=-0.19 $Y=1.66 $X2=0.502 $Y2=1.94
cc_39 VPB N_A_N_c_75_n 0.0326515f $X=-0.19 $Y=1.66 $X2=0.502 $Y2=2.045
cc_40 VPB N_A_N_c_72_n 0.00817485f $X=-0.19 $Y=1.66 $X2=0.405 $Y2=1.275
cc_41 VPB N_A_114_74#_c_100_n 7.7196e-19 $X=-0.19 $Y=1.66 $X2=0.405 $Y2=1.615
cc_42 VPB N_A_114_74#_c_109_n 0.0255758f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.21
cc_43 VPB N_A_114_74#_c_110_n 0.024899f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_44 VPB N_A_114_74#_c_106_n 0.0122024f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_45 VPB N_A_114_74#_c_112_n 0.00906052f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_46 VPB N_A_114_74#_c_107_n 0.00814936f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_47 VPB N_B_c_168_n 0.0275208f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.78
cc_48 VPB N_B_c_170_n 0.00256745f $X=-0.19 $Y=1.66 $X2=0.405 $Y2=1.615
cc_49 VPB N_C_c_201_n 0.0273778f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.78
cc_50 VPB N_C_c_202_n 0.00583347f $X=-0.19 $Y=1.66 $X2=0.405 $Y2=1.615
cc_51 VPB N_A_266_94#_c_228_n 0.0295497f $X=-0.19 $Y=1.66 $X2=0.405 $Y2=1.275
cc_52 VPB N_A_266_94#_c_231_n 0.00419179f $X=-0.19 $Y=1.66 $X2=0.405 $Y2=1.275
cc_53 VPB N_A_266_94#_c_236_n 0.0142366f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_54 VPB N_A_266_94#_c_237_n 0.0040121f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_55 VPB N_VPWR_c_315_n 0.0120152f $X=-0.19 $Y=1.66 $X2=0.405 $Y2=1.275
cc_56 VPB N_VPWR_c_316_n 0.0462693f $X=-0.19 $Y=1.66 $X2=0.405 $Y2=1.615
cc_57 VPB N_VPWR_c_317_n 0.0336932f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.21
cc_58 VPB N_VPWR_c_318_n 0.0202787f $X=-0.19 $Y=1.66 $X2=0.405 $Y2=1.275
cc_59 VPB N_VPWR_c_319_n 0.0391783f $X=-0.19 $Y=1.66 $X2=0.347 $Y2=1.275
cc_60 VPB N_VPWR_c_320_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_61 VPB N_VPWR_c_321_n 0.0208961f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_62 VPB N_VPWR_c_322_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0.347 $Y2=1.665
cc_63 VPB N_VPWR_c_323_n 0.0201176f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_64 VPB N_VPWR_c_314_n 0.0881578f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_65 VPB X 0.0434696f $X=-0.19 $Y=1.66 $X2=0.347 $Y2=1.275
cc_66 VPB N_X_c_363_n 0.0159529f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_67 VPB N_X_c_361_n 0.00780005f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_68 N_A_N_M1008_g N_A_114_74#_c_103_n 0.00829387f $X=0.495 $Y=0.645 $X2=0
+ $Y2=0
cc_69 N_A_N_c_75_n N_A_114_74#_c_110_n 0.00406782f $X=0.502 $Y=2.045 $X2=0 $Y2=0
cc_70 N_A_N_M1008_g N_A_114_74#_c_104_n 0.00867488f $X=0.495 $Y=0.645 $X2=0
+ $Y2=0
cc_71 N_A_N_c_72_n N_A_114_74#_c_104_n 0.00725794f $X=0.405 $Y=1.275 $X2=0 $Y2=0
cc_72 N_A_N_c_71_n N_A_114_74#_c_105_n 0.00332712f $X=0.405 $Y=1.275 $X2=0 $Y2=0
cc_73 N_A_N_c_72_n N_A_114_74#_c_105_n 0.0397534f $X=0.405 $Y=1.275 $X2=0 $Y2=0
cc_74 N_A_N_M1008_g N_A_114_74#_c_106_n 0.0176124f $X=0.495 $Y=0.645 $X2=0 $Y2=0
cc_75 N_A_N_c_69_n N_A_114_74#_c_106_n 0.0176124f $X=0.405 $Y=1.615 $X2=0 $Y2=0
cc_76 N_A_N_c_72_n N_A_114_74#_c_106_n 7.04297e-19 $X=0.405 $Y=1.275 $X2=0 $Y2=0
cc_77 N_A_N_c_70_n N_A_114_74#_c_112_n 0.00332712f $X=0.405 $Y=1.78 $X2=0 $Y2=0
cc_78 N_A_N_c_75_n N_A_114_74#_c_112_n 0.00536561f $X=0.502 $Y=2.045 $X2=0 $Y2=0
cc_79 N_A_N_c_69_n N_A_114_74#_c_107_n 0.00332712f $X=0.405 $Y=1.615 $X2=0 $Y2=0
cc_80 N_A_N_c_70_n N_VPWR_c_316_n 0.00130639f $X=0.405 $Y=1.78 $X2=0 $Y2=0
cc_81 N_A_N_c_75_n N_VPWR_c_316_n 0.020185f $X=0.502 $Y=2.045 $X2=0 $Y2=0
cc_82 N_A_N_c_72_n N_VPWR_c_316_n 0.0181212f $X=0.405 $Y=1.275 $X2=0 $Y2=0
cc_83 N_A_N_c_75_n N_VPWR_c_319_n 0.00429299f $X=0.502 $Y=2.045 $X2=0 $Y2=0
cc_84 N_A_N_c_75_n N_VPWR_c_314_n 0.00852523f $X=0.502 $Y=2.045 $X2=0 $Y2=0
cc_85 N_A_N_M1008_g N_VGND_c_383_n 0.0180652f $X=0.495 $Y=0.645 $X2=0 $Y2=0
cc_86 N_A_N_c_71_n N_VGND_c_383_n 0.0014092f $X=0.405 $Y=1.275 $X2=0 $Y2=0
cc_87 N_A_N_c_72_n N_VGND_c_383_n 0.0287296f $X=0.405 $Y=1.275 $X2=0 $Y2=0
cc_88 N_A_N_M1008_g N_VGND_c_385_n 0.00383152f $X=0.495 $Y=0.645 $X2=0 $Y2=0
cc_89 N_A_N_M1008_g N_VGND_c_387_n 0.00762539f $X=0.495 $Y=0.645 $X2=0 $Y2=0
cc_90 N_A_114_74#_c_101_n N_B_M1005_g 0.0548083f $X=1.69 $Y=1.185 $X2=0 $Y2=0
cc_91 N_A_114_74#_c_102_n N_B_M1005_g 0.0101654f $X=1.61 $Y=1.185 $X2=0 $Y2=0
cc_92 N_A_114_74#_c_100_n N_B_c_168_n 0.0101654f $X=1.7 $Y=1.675 $X2=0 $Y2=0
cc_93 N_A_114_74#_c_109_n N_B_c_168_n 0.0243625f $X=1.7 $Y=1.765 $X2=0 $Y2=0
cc_94 N_A_114_74#_c_109_n N_B_c_170_n 8.62223e-19 $X=1.7 $Y=1.765 $X2=0 $Y2=0
cc_95 N_A_114_74#_c_102_n N_B_c_170_n 0.00101876f $X=1.61 $Y=1.185 $X2=0 $Y2=0
cc_96 N_A_114_74#_c_101_n N_A_266_94#_c_230_n 0.0112826f $X=1.69 $Y=1.185 $X2=0
+ $Y2=0
cc_97 N_A_114_74#_c_103_n N_A_266_94#_c_230_n 0.0159343f $X=0.78 $Y=0.645 $X2=0
+ $Y2=0
cc_98 N_A_114_74#_c_104_n N_A_266_94#_c_230_n 0.013901f $X=0.957 $Y=1.212 $X2=0
+ $Y2=0
cc_99 N_A_114_74#_c_99_n N_A_266_94#_c_231_n 0.00983996f $X=1.61 $Y=1.26 $X2=0
+ $Y2=0
cc_100 N_A_114_74#_c_100_n N_A_266_94#_c_231_n 0.00730149f $X=1.7 $Y=1.675 $X2=0
+ $Y2=0
cc_101 N_A_114_74#_c_109_n N_A_266_94#_c_231_n 0.0084038f $X=1.7 $Y=1.765 $X2=0
+ $Y2=0
cc_102 N_A_114_74#_c_102_n N_A_266_94#_c_231_n 0.00489741f $X=1.61 $Y=1.185
+ $X2=0 $Y2=0
cc_103 N_A_114_74#_c_105_n N_A_266_94#_c_231_n 0.0376823f $X=0.957 $Y=1.518
+ $X2=0 $Y2=0
cc_104 N_A_114_74#_c_106_n N_A_266_94#_c_231_n 0.00320796f $X=0.975 $Y=1.195
+ $X2=0 $Y2=0
cc_105 N_A_114_74#_c_112_n N_A_266_94#_c_231_n 0.0116419f $X=0.78 $Y=2.1 $X2=0
+ $Y2=0
cc_106 N_A_114_74#_c_101_n N_A_266_94#_c_232_n 0.00839128f $X=1.69 $Y=1.185
+ $X2=0 $Y2=0
cc_107 N_A_114_74#_c_102_n N_A_266_94#_c_232_n 0.00729494f $X=1.61 $Y=1.185
+ $X2=0 $Y2=0
cc_108 N_A_114_74#_c_109_n N_A_266_94#_c_250_n 0.0165054f $X=1.7 $Y=1.765 $X2=0
+ $Y2=0
cc_109 N_A_114_74#_c_99_n N_A_266_94#_c_233_n 0.00878777f $X=1.61 $Y=1.26 $X2=0
+ $Y2=0
cc_110 N_A_114_74#_c_101_n N_A_266_94#_c_233_n 0.00134888f $X=1.69 $Y=1.185
+ $X2=0 $Y2=0
cc_111 N_A_114_74#_c_102_n N_A_266_94#_c_233_n 2.23825e-19 $X=1.61 $Y=1.185
+ $X2=0 $Y2=0
cc_112 N_A_114_74#_c_104_n N_A_266_94#_c_233_n 0.013702f $X=0.957 $Y=1.212 $X2=0
+ $Y2=0
cc_113 N_A_114_74#_c_105_n N_A_266_94#_c_233_n 6.05e-19 $X=0.957 $Y=1.518 $X2=0
+ $Y2=0
cc_114 N_A_114_74#_c_106_n N_A_266_94#_c_233_n 6.14826e-19 $X=0.975 $Y=1.195
+ $X2=0 $Y2=0
cc_115 N_A_114_74#_c_109_n N_A_266_94#_c_236_n 0.01135f $X=1.7 $Y=1.765 $X2=0
+ $Y2=0
cc_116 N_A_114_74#_c_110_n N_A_266_94#_c_236_n 0.0284314f $X=0.78 $Y=2.265 $X2=0
+ $Y2=0
cc_117 N_A_114_74#_c_112_n N_A_266_94#_c_236_n 0.0084726f $X=0.78 $Y=2.1 $X2=0
+ $Y2=0
cc_118 N_A_114_74#_c_109_n N_A_266_94#_c_237_n 6.01988e-19 $X=1.7 $Y=1.765 $X2=0
+ $Y2=0
cc_119 N_A_114_74#_c_110_n N_VPWR_c_316_n 0.0346007f $X=0.78 $Y=2.265 $X2=0
+ $Y2=0
cc_120 N_A_114_74#_c_109_n N_VPWR_c_317_n 0.00570239f $X=1.7 $Y=1.765 $X2=0
+ $Y2=0
cc_121 N_A_114_74#_c_109_n N_VPWR_c_319_n 0.00393873f $X=1.7 $Y=1.765 $X2=0
+ $Y2=0
cc_122 N_A_114_74#_c_110_n N_VPWR_c_319_n 0.0146357f $X=0.78 $Y=2.265 $X2=0
+ $Y2=0
cc_123 N_A_114_74#_c_109_n N_VPWR_c_314_n 0.00462577f $X=1.7 $Y=1.765 $X2=0
+ $Y2=0
cc_124 N_A_114_74#_c_110_n N_VPWR_c_314_n 0.0121141f $X=0.78 $Y=2.265 $X2=0
+ $Y2=0
cc_125 N_A_114_74#_c_103_n N_VGND_c_383_n 0.0167375f $X=0.78 $Y=0.645 $X2=0
+ $Y2=0
cc_126 N_A_114_74#_c_104_n N_VGND_c_383_n 0.00701512f $X=0.957 $Y=1.212 $X2=0
+ $Y2=0
cc_127 N_A_114_74#_c_101_n N_VGND_c_385_n 0.00485498f $X=1.69 $Y=1.185 $X2=0
+ $Y2=0
cc_128 N_A_114_74#_c_103_n N_VGND_c_385_n 0.0145628f $X=0.78 $Y=0.645 $X2=0
+ $Y2=0
cc_129 N_A_114_74#_c_101_n N_VGND_c_387_n 0.00514438f $X=1.69 $Y=1.185 $X2=0
+ $Y2=0
cc_130 N_A_114_74#_c_103_n N_VGND_c_387_n 0.012086f $X=0.78 $Y=0.645 $X2=0 $Y2=0
cc_131 N_B_M1005_g N_C_M1009_g 0.0335091f $X=2.08 $Y=0.79 $X2=0 $Y2=0
cc_132 N_B_c_168_n N_C_c_201_n 0.0380832f $X=2.245 $Y=1.765 $X2=0 $Y2=0
cc_133 N_B_c_170_n N_C_c_201_n 4.88773e-19 $X=2.17 $Y=1.515 $X2=0 $Y2=0
cc_134 N_B_c_168_n N_C_c_202_n 0.00222599f $X=2.245 $Y=1.765 $X2=0 $Y2=0
cc_135 N_B_c_170_n N_C_c_202_n 0.0285913f $X=2.17 $Y=1.515 $X2=0 $Y2=0
cc_136 N_B_M1005_g N_A_266_94#_c_230_n 0.00297121f $X=2.08 $Y=0.79 $X2=0 $Y2=0
cc_137 N_B_M1005_g N_A_266_94#_c_231_n 0.00165534f $X=2.08 $Y=0.79 $X2=0 $Y2=0
cc_138 N_B_c_168_n N_A_266_94#_c_231_n 8.56404e-19 $X=2.245 $Y=1.765 $X2=0 $Y2=0
cc_139 N_B_c_170_n N_A_266_94#_c_231_n 0.0161999f $X=2.17 $Y=1.515 $X2=0 $Y2=0
cc_140 N_B_M1005_g N_A_266_94#_c_232_n 0.0152776f $X=2.08 $Y=0.79 $X2=0 $Y2=0
cc_141 N_B_c_168_n N_A_266_94#_c_232_n 0.00489479f $X=2.245 $Y=1.765 $X2=0 $Y2=0
cc_142 N_B_c_170_n N_A_266_94#_c_232_n 0.0245335f $X=2.17 $Y=1.515 $X2=0 $Y2=0
cc_143 N_B_c_168_n N_A_266_94#_c_250_n 0.0135176f $X=2.245 $Y=1.765 $X2=0 $Y2=0
cc_144 N_B_c_170_n N_A_266_94#_c_250_n 0.0210925f $X=2.17 $Y=1.515 $X2=0 $Y2=0
cc_145 N_B_c_168_n N_A_266_94#_c_236_n 5.36224e-19 $X=2.245 $Y=1.765 $X2=0 $Y2=0
cc_146 N_B_c_168_n N_A_266_94#_c_237_n 0.00807882f $X=2.245 $Y=1.765 $X2=0 $Y2=0
cc_147 N_B_c_170_n N_A_266_94#_c_237_n 0.00137314f $X=2.17 $Y=1.515 $X2=0 $Y2=0
cc_148 N_B_c_168_n N_VPWR_c_317_n 0.00360626f $X=2.245 $Y=1.765 $X2=0 $Y2=0
cc_149 N_B_c_168_n N_VPWR_c_321_n 0.00396914f $X=2.245 $Y=1.765 $X2=0 $Y2=0
cc_150 N_B_c_168_n N_VPWR_c_314_n 0.00462577f $X=2.245 $Y=1.765 $X2=0 $Y2=0
cc_151 N_B_M1005_g N_VGND_c_384_n 0.00268474f $X=2.08 $Y=0.79 $X2=0 $Y2=0
cc_152 N_B_M1005_g N_VGND_c_385_n 0.00507111f $X=2.08 $Y=0.79 $X2=0 $Y2=0
cc_153 N_B_M1005_g N_VGND_c_387_n 0.00514438f $X=2.08 $Y=0.79 $X2=0 $Y2=0
cc_154 N_C_M1009_g N_A_266_94#_c_228_n 0.00132954f $X=2.62 $Y=0.79 $X2=0 $Y2=0
cc_155 N_C_c_201_n N_A_266_94#_c_228_n 0.0426747f $X=2.7 $Y=1.765 $X2=0 $Y2=0
cc_156 N_C_c_202_n N_A_266_94#_c_228_n 0.00268644f $X=2.71 $Y=1.515 $X2=0 $Y2=0
cc_157 N_C_M1009_g N_A_266_94#_M1002_g 0.00939291f $X=2.62 $Y=0.79 $X2=0 $Y2=0
cc_158 N_C_M1009_g N_A_266_94#_c_232_n 0.0170163f $X=2.62 $Y=0.79 $X2=0 $Y2=0
cc_159 N_C_c_201_n N_A_266_94#_c_232_n 0.00691332f $X=2.7 $Y=1.765 $X2=0 $Y2=0
cc_160 N_C_c_202_n N_A_266_94#_c_232_n 0.0454831f $X=2.71 $Y=1.515 $X2=0 $Y2=0
cc_161 N_C_c_201_n N_A_266_94#_c_237_n 0.00918905f $X=2.7 $Y=1.765 $X2=0 $Y2=0
cc_162 N_C_c_202_n N_A_266_94#_c_237_n 0.00733542f $X=2.71 $Y=1.515 $X2=0 $Y2=0
cc_163 N_C_c_201_n N_VPWR_c_318_n 0.0105493f $X=2.7 $Y=1.765 $X2=0 $Y2=0
cc_164 N_C_c_202_n N_VPWR_c_318_n 0.00246882f $X=2.71 $Y=1.515 $X2=0 $Y2=0
cc_165 N_C_c_201_n N_VPWR_c_321_n 0.00393873f $X=2.7 $Y=1.765 $X2=0 $Y2=0
cc_166 N_C_c_201_n N_VPWR_c_314_n 0.00462577f $X=2.7 $Y=1.765 $X2=0 $Y2=0
cc_167 N_C_M1009_g N_X_c_359_n 6.21799e-19 $X=2.62 $Y=0.79 $X2=0 $Y2=0
cc_168 N_C_c_201_n N_X_c_363_n 7.37845e-19 $X=2.7 $Y=1.765 $X2=0 $Y2=0
cc_169 N_C_M1009_g N_VGND_c_384_n 0.0203753f $X=2.62 $Y=0.79 $X2=0 $Y2=0
cc_170 N_C_M1009_g N_VGND_c_385_n 0.00269285f $X=2.62 $Y=0.79 $X2=0 $Y2=0
cc_171 N_C_M1009_g N_VGND_c_387_n 0.00277796f $X=2.62 $Y=0.79 $X2=0 $Y2=0
cc_172 N_A_266_94#_c_250_n N_VPWR_M1001_d 0.0108794f $X=2.31 $Y=2.035 $X2=0
+ $Y2=0
cc_173 N_A_266_94#_c_250_n N_VPWR_c_317_n 0.0228618f $X=2.31 $Y=2.035 $X2=0
+ $Y2=0
cc_174 N_A_266_94#_c_236_n N_VPWR_c_317_n 0.0161747f $X=1.475 $Y=1.985 $X2=0
+ $Y2=0
cc_175 N_A_266_94#_c_237_n N_VPWR_c_317_n 0.0161747f $X=2.475 $Y=2.115 $X2=0
+ $Y2=0
cc_176 N_A_266_94#_c_228_n N_VPWR_c_318_n 0.0141373f $X=3.285 $Y=1.765 $X2=0
+ $Y2=0
cc_177 N_A_266_94#_c_232_n N_VPWR_c_318_n 0.00642764f $X=3.045 $Y=1.135 $X2=0
+ $Y2=0
cc_178 N_A_266_94#_c_237_n N_VPWR_c_318_n 0.0510966f $X=2.475 $Y=2.115 $X2=0
+ $Y2=0
cc_179 N_A_266_94#_c_236_n N_VPWR_c_319_n 0.0066794f $X=1.475 $Y=1.985 $X2=0
+ $Y2=0
cc_180 N_A_266_94#_c_237_n N_VPWR_c_321_n 0.00665021f $X=2.475 $Y=2.115 $X2=0
+ $Y2=0
cc_181 N_A_266_94#_c_228_n N_VPWR_c_323_n 0.00445602f $X=3.285 $Y=1.765 $X2=0
+ $Y2=0
cc_182 N_A_266_94#_c_228_n N_VPWR_c_314_n 0.00865368f $X=3.285 $Y=1.765 $X2=0
+ $Y2=0
cc_183 N_A_266_94#_c_236_n N_VPWR_c_314_n 0.00997343f $X=1.475 $Y=1.985 $X2=0
+ $Y2=0
cc_184 N_A_266_94#_c_237_n N_VPWR_c_314_n 0.0099564f $X=2.475 $Y=2.115 $X2=0
+ $Y2=0
cc_185 N_A_266_94#_M1002_g N_X_c_359_n 0.00888737f $X=3.335 $Y=0.74 $X2=0 $Y2=0
cc_186 N_A_266_94#_M1002_g N_X_c_360_n 0.00396511f $X=3.335 $Y=0.74 $X2=0 $Y2=0
cc_187 N_A_266_94#_c_232_n N_X_c_360_n 0.00630461f $X=3.045 $Y=1.135 $X2=0 $Y2=0
cc_188 N_A_266_94#_c_228_n X 0.0108779f $X=3.285 $Y=1.765 $X2=0 $Y2=0
cc_189 N_A_266_94#_c_228_n N_X_c_363_n 0.00477393f $X=3.285 $Y=1.765 $X2=0 $Y2=0
cc_190 N_A_266_94#_c_232_n N_X_c_363_n 0.00531127f $X=3.045 $Y=1.135 $X2=0 $Y2=0
cc_191 N_A_266_94#_c_228_n N_X_c_361_n 0.00699163f $X=3.285 $Y=1.765 $X2=0 $Y2=0
cc_192 N_A_266_94#_M1002_g N_X_c_361_n 0.00252147f $X=3.335 $Y=0.74 $X2=0 $Y2=0
cc_193 N_A_266_94#_c_232_n N_X_c_361_n 0.0306189f $X=3.045 $Y=1.135 $X2=0 $Y2=0
cc_194 N_A_266_94#_c_232_n N_VGND_M1009_d 0.00592064f $X=3.045 $Y=1.135 $X2=0
+ $Y2=0
cc_195 N_A_266_94#_c_228_n N_VGND_c_384_n 5.63838e-19 $X=3.285 $Y=1.765 $X2=0
+ $Y2=0
cc_196 N_A_266_94#_M1002_g N_VGND_c_384_n 0.00656426f $X=3.335 $Y=0.74 $X2=0
+ $Y2=0
cc_197 N_A_266_94#_c_232_n N_VGND_c_384_n 0.043095f $X=3.045 $Y=1.135 $X2=0
+ $Y2=0
cc_198 N_A_266_94#_c_230_n N_VGND_c_385_n 0.0103491f $X=1.475 $Y=0.615 $X2=0
+ $Y2=0
cc_199 N_A_266_94#_M1002_g N_VGND_c_386_n 0.00434272f $X=3.335 $Y=0.74 $X2=0
+ $Y2=0
cc_200 N_A_266_94#_M1002_g N_VGND_c_387_n 0.00828751f $X=3.335 $Y=0.74 $X2=0
+ $Y2=0
cc_201 N_A_266_94#_c_230_n N_VGND_c_387_n 0.0113354f $X=1.475 $Y=0.615 $X2=0
+ $Y2=0
cc_202 N_A_266_94#_c_232_n A_353_94# 0.0048076f $X=3.045 $Y=1.135 $X2=-0.19
+ $Y2=-0.245
cc_203 N_A_266_94#_c_232_n A_431_94# 0.0106289f $X=3.045 $Y=1.135 $X2=-0.19
+ $Y2=-0.245
cc_204 N_VPWR_c_323_n X 0.0181635f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_205 N_VPWR_c_314_n X 0.0150013f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_206 N_VPWR_c_318_n N_X_c_363_n 0.0407049f $X=3.01 $Y=2.115 $X2=0 $Y2=0
cc_207 N_X_c_359_n N_VGND_c_384_n 0.0211012f $X=3.55 $Y=0.515 $X2=0 $Y2=0
cc_208 N_X_c_359_n N_VGND_c_386_n 0.0163488f $X=3.55 $Y=0.515 $X2=0 $Y2=0
cc_209 N_X_c_359_n N_VGND_c_387_n 0.0134757f $X=3.55 $Y=0.515 $X2=0 $Y2=0
