* File: sky130_fd_sc_hs__and2_1.pxi.spice
* Created: Tue Sep  1 19:54:34 2020
* 
x_PM_SKY130_FD_SC_HS__AND2_1%A N_A_c_47_n N_A_M1003_g N_A_c_49_n N_A_c_54_n
+ N_A_M1004_g N_A_c_50_n A A N_A_c_52_n PM_SKY130_FD_SC_HS__AND2_1%A
x_PM_SKY130_FD_SC_HS__AND2_1%B N_B_M1001_g N_B_c_86_n N_B_c_87_n N_B_M1002_g B
+ N_B_c_84_n N_B_c_85_n PM_SKY130_FD_SC_HS__AND2_1%B
x_PM_SKY130_FD_SC_HS__AND2_1%A_56_136# N_A_56_136#_M1003_s N_A_56_136#_M1004_d
+ N_A_56_136#_c_132_n N_A_56_136#_M1000_g N_A_56_136#_c_133_n
+ N_A_56_136#_M1005_g N_A_56_136#_c_134_n N_A_56_136#_c_138_n
+ N_A_56_136#_c_139_n N_A_56_136#_c_140_n N_A_56_136#_c_141_n
+ N_A_56_136#_c_142_n N_A_56_136#_c_143_n N_A_56_136#_c_135_n
+ PM_SKY130_FD_SC_HS__AND2_1%A_56_136#
x_PM_SKY130_FD_SC_HS__AND2_1%VPWR N_VPWR_M1004_s N_VPWR_M1002_d N_VPWR_c_202_n
+ N_VPWR_c_203_n N_VPWR_c_204_n N_VPWR_c_205_n N_VPWR_c_206_n N_VPWR_c_207_n
+ VPWR N_VPWR_c_208_n N_VPWR_c_201_n PM_SKY130_FD_SC_HS__AND2_1%VPWR
x_PM_SKY130_FD_SC_HS__AND2_1%X N_X_M1005_d N_X_M1000_d N_X_c_231_n X X X
+ N_X_c_232_n X PM_SKY130_FD_SC_HS__AND2_1%X
x_PM_SKY130_FD_SC_HS__AND2_1%VGND N_VGND_M1001_d N_VGND_c_253_n N_VGND_c_254_n
+ N_VGND_c_255_n VGND N_VGND_c_256_n N_VGND_c_257_n
+ PM_SKY130_FD_SC_HS__AND2_1%VGND
cc_1 VNB N_A_c_47_n 0.02449f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=0.57
cc_2 VNB N_A_M1003_g 0.0120472f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1
cc_3 VNB N_A_c_49_n 0.00665438f $X=-0.19 $Y=-0.245 $X2=0.745 $Y2=1.955
cc_4 VNB N_A_c_50_n 0.0204235f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=1.545
cc_5 VNB A 0.0358286f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.47
cc_6 VNB N_A_c_52_n 0.0544958f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=0.405
cc_7 VNB B 0.00237204f $X=-0.19 $Y=-0.245 $X2=0.745 $Y2=2.045
cc_8 VNB N_B_c_84_n 0.0272161f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=1.395
cc_9 VNB N_B_c_85_n 0.0182698f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.47
cc_10 VNB N_A_56_136#_c_132_n 0.0289949f $X=-0.19 $Y=-0.245 $X2=0.745 $Y2=1.545
cc_11 VNB N_A_56_136#_c_133_n 0.0216407f $X=-0.19 $Y=-0.245 $X2=0.745 $Y2=2.54
cc_12 VNB N_A_56_136#_c_134_n 0.0335551f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.47
cc_13 VNB N_A_56_136#_c_135_n 0.00556882f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_VPWR_c_201_n 0.103974f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_X_c_231_n 0.0367857f $X=-0.19 $Y=-0.245 $X2=0.745 $Y2=2.54
cc_16 VNB N_X_c_232_n 0.02259f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_VGND_c_253_n 0.0186268f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1
cc_18 VNB N_VGND_c_254_n 0.037648f $X=-0.19 $Y=-0.245 $X2=0.745 $Y2=2.045
cc_19 VNB N_VGND_c_255_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0.745 $Y2=2.54
cc_20 VNB N_VGND_c_256_n 0.0224545f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=0.462
cc_21 VNB N_VGND_c_257_n 0.173493f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VPB N_A_c_49_n 0.0181314f $X=-0.19 $Y=1.66 $X2=0.745 $Y2=1.955
cc_23 VPB N_A_c_54_n 0.0272249f $X=-0.19 $Y=1.66 $X2=0.745 $Y2=2.045
cc_24 VPB N_B_c_86_n 0.0156915f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1
cc_25 VPB N_B_c_87_n 0.0225764f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1
cc_26 VPB B 0.00138105f $X=-0.19 $Y=1.66 $X2=0.745 $Y2=2.045
cc_27 VPB N_B_c_84_n 0.00562806f $X=-0.19 $Y=1.66 $X2=0.7 $Y2=1.395
cc_28 VPB N_A_56_136#_c_132_n 0.0328698f $X=-0.19 $Y=1.66 $X2=0.745 $Y2=1.545
cc_29 VPB N_A_56_136#_c_134_n 0.0101637f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=0.47
cc_30 VPB N_A_56_136#_c_138_n 0.00257779f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_31 VPB N_A_56_136#_c_139_n 0.0141715f $X=-0.19 $Y=1.66 $X2=0.67 $Y2=0.405
cc_32 VPB N_A_56_136#_c_140_n 0.00397788f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=0.462
cc_33 VPB N_A_56_136#_c_141_n 0.00402361f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_34 VPB N_A_56_136#_c_142_n 0.0018089f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_35 VPB N_A_56_136#_c_143_n 0.00948496f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_36 VPB N_A_56_136#_c_135_n 4.76351e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_37 VPB N_VPWR_c_202_n 0.0396256f $X=-0.19 $Y=1.66 $X2=0.745 $Y2=2.045
cc_38 VPB N_VPWR_c_203_n 0.00652655f $X=-0.19 $Y=1.66 $X2=0.7 $Y2=1.545
cc_39 VPB N_VPWR_c_204_n 0.013281f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_40 VPB N_VPWR_c_205_n 0.00623744f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_41 VPB N_VPWR_c_206_n 0.0195482f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=0.405
cc_42 VPB N_VPWR_c_207_n 0.00614127f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=0.405
cc_43 VPB N_VPWR_c_208_n 0.0205542f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_44 VPB N_VPWR_c_201_n 0.0661559f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_45 VPB X 0.0535235f $X=-0.19 $Y=1.66 $X2=0.7 $Y2=1.545
cc_46 VPB N_X_c_232_n 0.00905736f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_47 N_A_c_49_n N_B_c_86_n 0.00718885f $X=0.745 $Y=1.955 $X2=0 $Y2=0
cc_48 N_A_c_54_n N_B_c_87_n 0.0269971f $X=0.745 $Y=2.045 $X2=0 $Y2=0
cc_49 N_A_M1003_g B 0.00151136f $X=0.64 $Y=1 $X2=0 $Y2=0
cc_50 N_A_c_50_n B 0.00112834f $X=0.7 $Y=1.545 $X2=0 $Y2=0
cc_51 N_A_M1003_g N_B_c_84_n 0.00137655f $X=0.64 $Y=1 $X2=0 $Y2=0
cc_52 N_A_c_50_n N_B_c_84_n 0.0150816f $X=0.7 $Y=1.545 $X2=0 $Y2=0
cc_53 N_A_c_47_n N_B_c_85_n 0.00298419f $X=0.64 $Y=0.57 $X2=0 $Y2=0
cc_54 N_A_M1003_g N_B_c_85_n 0.0210976f $X=0.64 $Y=1 $X2=0 $Y2=0
cc_55 A N_B_c_85_n 0.00194518f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_56 N_A_M1003_g N_A_56_136#_c_134_n 0.014365f $X=0.64 $Y=1 $X2=0 $Y2=0
cc_57 N_A_c_49_n N_A_56_136#_c_134_n 0.0108936f $X=0.745 $Y=1.955 $X2=0 $Y2=0
cc_58 N_A_c_50_n N_A_56_136#_c_134_n 0.00648097f $X=0.7 $Y=1.545 $X2=0 $Y2=0
cc_59 A N_A_56_136#_c_134_n 0.0255901f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_60 N_A_c_52_n N_A_56_136#_c_134_n 0.00172729f $X=0.61 $Y=0.405 $X2=0 $Y2=0
cc_61 N_A_c_49_n N_A_56_136#_c_138_n 0.0129216f $X=0.745 $Y=1.955 $X2=0 $Y2=0
cc_62 N_A_c_54_n N_A_56_136#_c_138_n 0.0101329f $X=0.745 $Y=2.045 $X2=0 $Y2=0
cc_63 N_A_c_50_n N_A_56_136#_c_138_n 0.00232067f $X=0.7 $Y=1.545 $X2=0 $Y2=0
cc_64 N_A_c_54_n N_A_56_136#_c_140_n 0.00764413f $X=0.745 $Y=2.045 $X2=0 $Y2=0
cc_65 N_A_c_54_n N_VPWR_c_202_n 0.0151914f $X=0.745 $Y=2.045 $X2=0 $Y2=0
cc_66 N_A_c_54_n N_VPWR_c_206_n 0.00413917f $X=0.745 $Y=2.045 $X2=0 $Y2=0
cc_67 N_A_c_54_n N_VPWR_c_201_n 0.00818241f $X=0.745 $Y=2.045 $X2=0 $Y2=0
cc_68 N_A_c_47_n N_VGND_c_253_n 0.00157877f $X=0.64 $Y=0.57 $X2=0 $Y2=0
cc_69 A N_VGND_c_253_n 0.015731f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_70 A N_VGND_c_254_n 0.0478766f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_71 N_A_c_52_n N_VGND_c_254_n 0.0116176f $X=0.61 $Y=0.405 $X2=0 $Y2=0
cc_72 N_A_c_47_n N_VGND_c_257_n 0.00487856f $X=0.64 $Y=0.57 $X2=0 $Y2=0
cc_73 A N_VGND_c_257_n 0.0249126f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_74 N_A_c_52_n N_VGND_c_257_n 0.0101636f $X=0.61 $Y=0.405 $X2=0 $Y2=0
cc_75 N_B_c_86_n N_A_56_136#_c_132_n 0.0109781f $X=1.245 $Y=1.955 $X2=0 $Y2=0
cc_76 N_B_c_87_n N_A_56_136#_c_132_n 0.0164827f $X=1.245 $Y=2.045 $X2=0 $Y2=0
cc_77 B N_A_56_136#_c_132_n 3.66423e-19 $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_78 N_B_c_84_n N_A_56_136#_c_132_n 0.0174253f $X=1.24 $Y=1.515 $X2=0 $Y2=0
cc_79 B N_A_56_136#_c_133_n 0.00358991f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_80 N_B_c_85_n N_A_56_136#_c_133_n 0.0187211f $X=1.24 $Y=1.35 $X2=0 $Y2=0
cc_81 B N_A_56_136#_c_134_n 0.0171072f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_82 N_B_c_84_n N_A_56_136#_c_134_n 5.35461e-19 $X=1.24 $Y=1.515 $X2=0 $Y2=0
cc_83 N_B_c_85_n N_A_56_136#_c_134_n 0.00171729f $X=1.24 $Y=1.35 $X2=0 $Y2=0
cc_84 N_B_c_87_n N_A_56_136#_c_140_n 0.0160324f $X=1.245 $Y=2.045 $X2=0 $Y2=0
cc_85 N_B_c_86_n N_A_56_136#_c_141_n 0.00497599f $X=1.245 $Y=1.955 $X2=0 $Y2=0
cc_86 N_B_c_87_n N_A_56_136#_c_141_n 0.00830695f $X=1.245 $Y=2.045 $X2=0 $Y2=0
cc_87 B N_A_56_136#_c_141_n 0.0164847f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_88 N_B_c_84_n N_A_56_136#_c_141_n 4.86414e-19 $X=1.24 $Y=1.515 $X2=0 $Y2=0
cc_89 N_B_c_86_n N_A_56_136#_c_142_n 0.00334443f $X=1.245 $Y=1.955 $X2=0 $Y2=0
cc_90 N_B_c_86_n N_A_56_136#_c_143_n 0.00208396f $X=1.245 $Y=1.955 $X2=0 $Y2=0
cc_91 N_B_c_87_n N_A_56_136#_c_143_n 0.0010315f $X=1.245 $Y=2.045 $X2=0 $Y2=0
cc_92 B N_A_56_136#_c_143_n 0.00937184f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_93 N_B_c_84_n N_A_56_136#_c_143_n 6.23375e-19 $X=1.24 $Y=1.515 $X2=0 $Y2=0
cc_94 B N_A_56_136#_c_135_n 0.0258883f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_95 N_B_c_84_n N_A_56_136#_c_135_n 0.00201866f $X=1.24 $Y=1.515 $X2=0 $Y2=0
cc_96 N_B_c_87_n N_VPWR_c_202_n 7.15022e-19 $X=1.245 $Y=2.045 $X2=0 $Y2=0
cc_97 N_B_c_87_n N_VPWR_c_203_n 0.00984508f $X=1.245 $Y=2.045 $X2=0 $Y2=0
cc_98 N_B_c_87_n N_VPWR_c_206_n 0.00445347f $X=1.245 $Y=2.045 $X2=0 $Y2=0
cc_99 N_B_c_87_n N_VPWR_c_201_n 0.00858831f $X=1.245 $Y=2.045 $X2=0 $Y2=0
cc_100 N_B_c_85_n N_X_c_231_n 8.72408e-19 $X=1.24 $Y=1.35 $X2=0 $Y2=0
cc_101 B A_143_136# 8.67896e-19 $X=1.115 $Y=1.21 $X2=-0.19 $Y2=-0.245
cc_102 B N_VGND_M1001_d 0.00152312f $X=1.115 $Y=1.21 $X2=-0.19 $Y2=-0.245
cc_103 B N_VGND_c_253_n 0.00546541f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_104 N_B_c_84_n N_VGND_c_253_n 3.3155e-19 $X=1.24 $Y=1.515 $X2=0 $Y2=0
cc_105 N_B_c_85_n N_VGND_c_253_n 0.0043444f $X=1.24 $Y=1.35 $X2=0 $Y2=0
cc_106 N_B_c_85_n N_VGND_c_254_n 0.00428744f $X=1.24 $Y=1.35 $X2=0 $Y2=0
cc_107 N_B_c_85_n N_VGND_c_257_n 0.00476395f $X=1.24 $Y=1.35 $X2=0 $Y2=0
cc_108 N_A_56_136#_c_141_n N_VPWR_M1002_d 0.00754811f $X=1.58 $Y=1.935 $X2=0
+ $Y2=0
cc_109 N_A_56_136#_c_138_n N_VPWR_c_202_n 0.00498708f $X=0.855 $Y=1.935 $X2=0
+ $Y2=0
cc_110 N_A_56_136#_c_139_n N_VPWR_c_202_n 0.0219579f $X=0.59 $Y=1.935 $X2=0
+ $Y2=0
cc_111 N_A_56_136#_c_140_n N_VPWR_c_202_n 0.0320858f $X=1.02 $Y=2.265 $X2=0
+ $Y2=0
cc_112 N_A_56_136#_c_132_n N_VPWR_c_203_n 0.016211f $X=1.78 $Y=1.765 $X2=0 $Y2=0
cc_113 N_A_56_136#_c_140_n N_VPWR_c_203_n 0.0545031f $X=1.02 $Y=2.265 $X2=0
+ $Y2=0
cc_114 N_A_56_136#_c_141_n N_VPWR_c_203_n 0.0222798f $X=1.58 $Y=1.935 $X2=0
+ $Y2=0
cc_115 N_A_56_136#_c_140_n N_VPWR_c_206_n 0.0158666f $X=1.02 $Y=2.265 $X2=0
+ $Y2=0
cc_116 N_A_56_136#_c_132_n N_VPWR_c_208_n 0.00413917f $X=1.78 $Y=1.765 $X2=0
+ $Y2=0
cc_117 N_A_56_136#_c_132_n N_VPWR_c_201_n 0.00821544f $X=1.78 $Y=1.765 $X2=0
+ $Y2=0
cc_118 N_A_56_136#_c_140_n N_VPWR_c_201_n 0.012191f $X=1.02 $Y=2.265 $X2=0 $Y2=0
cc_119 N_A_56_136#_c_132_n N_X_c_231_n 0.00239376f $X=1.78 $Y=1.765 $X2=0 $Y2=0
cc_120 N_A_56_136#_c_133_n N_X_c_231_n 0.0106952f $X=1.79 $Y=1.35 $X2=0 $Y2=0
cc_121 N_A_56_136#_c_135_n N_X_c_231_n 0.00842104f $X=1.81 $Y=1.515 $X2=0 $Y2=0
cc_122 N_A_56_136#_c_132_n X 0.00958783f $X=1.78 $Y=1.765 $X2=0 $Y2=0
cc_123 N_A_56_136#_c_141_n X 0.0141946f $X=1.58 $Y=1.935 $X2=0 $Y2=0
cc_124 N_A_56_136#_c_135_n X 0.00445935f $X=1.81 $Y=1.515 $X2=0 $Y2=0
cc_125 N_A_56_136#_c_132_n N_X_c_232_n 0.00461053f $X=1.78 $Y=1.765 $X2=0 $Y2=0
cc_126 N_A_56_136#_c_133_n N_X_c_232_n 0.00348686f $X=1.79 $Y=1.35 $X2=0 $Y2=0
cc_127 N_A_56_136#_c_142_n N_X_c_232_n 0.00456343f $X=1.665 $Y=1.85 $X2=0 $Y2=0
cc_128 N_A_56_136#_c_135_n N_X_c_232_n 0.0251162f $X=1.81 $Y=1.515 $X2=0 $Y2=0
cc_129 N_A_56_136#_c_132_n N_VGND_c_253_n 4.5946e-19 $X=1.78 $Y=1.765 $X2=0
+ $Y2=0
cc_130 N_A_56_136#_c_133_n N_VGND_c_253_n 0.00769141f $X=1.79 $Y=1.35 $X2=0
+ $Y2=0
cc_131 N_A_56_136#_c_135_n N_VGND_c_253_n 0.00429544f $X=1.81 $Y=1.515 $X2=0
+ $Y2=0
cc_132 N_A_56_136#_c_133_n N_VGND_c_256_n 0.0046731f $X=1.79 $Y=1.35 $X2=0 $Y2=0
cc_133 N_A_56_136#_c_133_n N_VGND_c_257_n 0.00505379f $X=1.79 $Y=1.35 $X2=0
+ $Y2=0
cc_134 N_VPWR_c_203_n X 0.0549067f $X=1.555 $Y=2.355 $X2=0 $Y2=0
cc_135 N_VPWR_c_208_n X 0.017536f $X=2.16 $Y=3.33 $X2=0 $Y2=0
cc_136 N_VPWR_c_201_n X 0.0145148f $X=2.16 $Y=3.33 $X2=0 $Y2=0
cc_137 N_X_c_231_n N_VGND_c_253_n 0.0226294f $X=2.005 $Y=0.645 $X2=0 $Y2=0
cc_138 N_X_c_231_n N_VGND_c_256_n 0.0141483f $X=2.005 $Y=0.645 $X2=0 $Y2=0
cc_139 N_X_c_231_n N_VGND_c_257_n 0.0161522f $X=2.005 $Y=0.645 $X2=0 $Y2=0
