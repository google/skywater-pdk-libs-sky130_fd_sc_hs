* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hs__mux4_2 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
X0 a_909_74# S0 a_1152_392# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=150000u
X1 a_255_74# S0 a_333_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X2 VPWR a_1429_74# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X3 VGND a_1429_74# X VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X4 a_333_74# S0 a_618_392# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=150000u
X5 a_1152_392# A2 VPWR VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=150000u
X6 VGND A1 a_255_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X7 X a_1429_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X8 VGND A3 a_831_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X9 a_1429_74# a_1500_94# a_333_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X10 a_31_94# S0 VPWR VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=150000u
X11 a_1429_74# a_1500_94# a_909_74# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=150000u
X12 a_909_74# a_31_94# a_1047_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X13 a_1047_74# A2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X14 a_1500_94# S1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=150000u
X15 a_831_74# S0 a_909_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X16 VPWR A3 a_840_392# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=150000u
X17 a_1500_94# S1 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X18 a_333_74# a_31_94# a_507_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X19 a_507_74# A0 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X20 a_840_392# a_31_94# a_909_74# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=150000u
X21 a_618_392# A0 VPWR VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=150000u
X22 a_333_74# S1 a_1429_74# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=150000u
X23 a_31_94# S0 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X24 a_909_74# S1 a_1429_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X25 X a_1429_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X26 VPWR A1 a_264_392# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=150000u
X27 a_264_392# a_31_94# a_333_74# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=150000u
.ends
