* File: sky130_fd_sc_hs__nor2b_1.spice
* Created: Thu Aug 27 20:53:27 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hs__nor2b_1.pex.spice"
.subckt sky130_fd_sc_hs__nor2b_1  VNB VPB B_N A VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A	A
* B_N	B_N
* VPB	VPB
* VNB	VNB
MM1003 N_VGND_M1003_d N_B_N_M1003_g N_A_27_112#_M1003_s VNB NLOWVT L=0.15 W=0.55
+ AD=0.130955 AS=0.2805 PD=1.02326 PS=2.12 NRD=39.816 NRS=0 M=1 R=3.66667
+ SA=75000.4 SB=75001.4 A=0.0825 P=1.4 MULT=1
MM1005 N_Y_M1005_d N_A_M1005_g N_VGND_M1003_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.13135 AS=0.176195 PD=1.095 PS=1.37674 NRD=12.156 NRS=0 M=1 R=4.93333
+ SA=75000.8 SB=75000.8 A=0.111 P=1.78 MULT=1
MM1002 N_VGND_M1002_d N_A_27_112#_M1002_g N_Y_M1005_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.2627 AS=0.13135 PD=2.19 PS=1.095 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.3
+ SB=75000.3 A=0.111 P=1.78 MULT=1
MM1000 N_VPWR_M1000_d N_B_N_M1000_g N_A_27_112#_M1000_s VPB PSHORT L=0.15 W=0.84
+ AD=0.201 AS=0.2478 PD=1.35429 PS=2.27 NRD=39.8531 NRS=2.3443 M=1 R=5.6
+ SA=75000.2 SB=75001.3 A=0.126 P=1.98 MULT=1
MM1001 A_278_368# N_A_M1001_g N_VPWR_M1000_d VPB PSHORT L=0.15 W=1.12 AD=0.1512
+ AS=0.268 PD=1.39 PS=1.80571 NRD=14.0658 NRS=1.7533 M=1 R=7.46667 SA=75000.7
+ SB=75000.7 A=0.168 P=2.54 MULT=1
MM1004 N_Y_M1004_d N_A_27_112#_M1004_g A_278_368# VPB PSHORT L=0.15 W=1.12
+ AD=0.42 AS=0.1512 PD=2.99 PS=1.39 NRD=2.6201 NRS=14.0658 M=1 R=7.46667
+ SA=75001.1 SB=75000.3 A=0.168 P=2.54 MULT=1
DX6_noxref VNB VPB NWDIODE A=5.1708 P=9.28
*
.include "sky130_fd_sc_hs__nor2b_1.pxi.spice"
*
.ends
*
*
