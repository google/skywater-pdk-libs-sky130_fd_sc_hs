* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hs__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
M1000 VPWR a_81_264# X VPB pshort w=1.12e+06u l=150000u
+  ad=6.38e+11p pd=5.45e+06u as=3.08e+11p ps=2.79e+06u
M1001 a_364_392# B1 a_81_264# VPB pshort w=1e+06u l=150000u
+  ad=5.75e+11p pd=5.15e+06u as=2.75e+11p ps=2.55e+06u
M1002 a_364_392# A2 VPWR VPB pshort w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1003 VPWR A1 a_364_392# VPB pshort w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 VGND a_81_264# X VNB nlowvt w=740000u l=150000u
+  ad=4.541e+11p pd=4.09e+06u as=1.961e+11p ps=2.01e+06u
M1005 VGND A2 a_452_136# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=2.08e+11p ps=1.93e+06u
M1006 a_81_264# B1 VGND VNB nlowvt w=640000u l=150000u
+  ad=1.792e+11p pd=1.84e+06u as=0p ps=0u
M1007 a_452_136# A1 a_81_264# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
