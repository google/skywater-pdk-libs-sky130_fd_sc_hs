* File: sky130_fd_sc_hs__or2b_1.pxi.spice
* Created: Tue Sep  1 20:20:06 2020
* 
x_PM_SKY130_FD_SC_HS__OR2B_1%B_N N_B_N_c_59_n N_B_N_c_64_n N_B_N_c_65_n
+ N_B_N_M1005_g N_B_N_c_60_n N_B_N_c_61_n N_B_N_M1002_g B_N
+ PM_SKY130_FD_SC_HS__OR2B_1%B_N
x_PM_SKY130_FD_SC_HS__OR2B_1%A_27_112# N_A_27_112#_M1002_s N_A_27_112#_M1005_s
+ N_A_27_112#_M1000_g N_A_27_112#_c_100_n N_A_27_112#_M1004_g N_A_27_112#_c_94_n
+ N_A_27_112#_c_95_n N_A_27_112#_c_102_n N_A_27_112#_c_103_n N_A_27_112#_c_104_n
+ N_A_27_112#_c_117_n N_A_27_112#_c_96_n N_A_27_112#_c_97_n N_A_27_112#_c_98_n
+ N_A_27_112#_c_99_n PM_SKY130_FD_SC_HS__OR2B_1%A_27_112#
x_PM_SKY130_FD_SC_HS__OR2B_1%A N_A_M1001_g N_A_c_163_n N_A_M1006_g A N_A_c_164_n
+ PM_SKY130_FD_SC_HS__OR2B_1%A
x_PM_SKY130_FD_SC_HS__OR2B_1%A_264_368# N_A_264_368#_M1000_d
+ N_A_264_368#_M1004_s N_A_264_368#_c_194_n N_A_264_368#_M1003_g
+ N_A_264_368#_M1007_g N_A_264_368#_c_201_n N_A_264_368#_c_196_n
+ N_A_264_368#_c_197_n N_A_264_368#_c_198_n N_A_264_368#_c_203_n
+ N_A_264_368#_c_199_n PM_SKY130_FD_SC_HS__OR2B_1%A_264_368#
x_PM_SKY130_FD_SC_HS__OR2B_1%VPWR N_VPWR_M1005_d N_VPWR_M1006_d N_VPWR_c_263_n
+ N_VPWR_c_264_n N_VPWR_c_265_n N_VPWR_c_266_n VPWR N_VPWR_c_267_n
+ N_VPWR_c_268_n N_VPWR_c_262_n N_VPWR_c_270_n PM_SKY130_FD_SC_HS__OR2B_1%VPWR
x_PM_SKY130_FD_SC_HS__OR2B_1%X N_X_M1007_d N_X_M1003_d N_X_c_300_n N_X_c_301_n X
+ X X N_X_c_304_n N_X_c_302_n X PM_SKY130_FD_SC_HS__OR2B_1%X
x_PM_SKY130_FD_SC_HS__OR2B_1%VGND N_VGND_M1002_d N_VGND_M1001_d N_VGND_c_323_n
+ N_VGND_c_324_n N_VGND_c_325_n N_VGND_c_326_n VGND N_VGND_c_327_n
+ N_VGND_c_328_n N_VGND_c_329_n N_VGND_c_330_n PM_SKY130_FD_SC_HS__OR2B_1%VGND
cc_1 VNB N_B_N_c_59_n 0.0695094f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.7
cc_2 VNB N_B_N_c_60_n 0.02624f $X=-0.19 $Y=-0.245 $X2=0.805 $Y2=1.295
cc_3 VNB N_B_N_c_61_n 0.0243562f $X=-0.19 $Y=-0.245 $X2=0.88 $Y2=1.22
cc_4 VNB B_N 0.00771224f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_5 VNB N_A_27_112#_M1000_g 0.0236728f $X=-0.19 $Y=-0.245 $X2=0.88 $Y2=0.835
cc_6 VNB N_A_27_112#_c_94_n 0.0441328f $X=-0.19 $Y=-0.245 $X2=0.36 $Y2=1.385
cc_7 VNB N_A_27_112#_c_95_n 0.0137914f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.385
cc_8 VNB N_A_27_112#_c_96_n 0.00279704f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A_27_112#_c_97_n 0.00409161f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_27_112#_c_98_n 0.0155571f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_27_112#_c_99_n 0.0144242f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_M1001_g 0.0263428f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.045
cc_13 VNB N_A_c_163_n 0.0281461f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.54
cc_14 VNB N_A_c_164_n 0.00180753f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_264_368#_c_194_n 0.0364436f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=1.295
cc_16 VNB N_A_264_368#_M1007_g 0.0294109f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_264_368#_c_196_n 0.00325419f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.385
cc_18 VNB N_A_264_368#_c_197_n 0.00335286f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_264_368#_c_198_n 0.0202157f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_264_368#_c_199_n 0.00626634f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_VPWR_c_262_n 0.143779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_X_c_300_n 0.0272846f $X=-0.19 $Y=-0.245 $X2=0.88 $Y2=0.835
cc_23 VNB N_X_c_301_n 0.0154926f $X=-0.19 $Y=-0.245 $X2=0.36 $Y2=1.295
cc_24 VNB N_X_c_302_n 0.0248898f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_VGND_c_323_n 0.0346814f $X=-0.19 $Y=-0.245 $X2=0.88 $Y2=0.835
cc_26 VNB N_VGND_c_324_n 0.0188865f $X=-0.19 $Y=-0.245 $X2=0.36 $Y2=1.295
cc_27 VNB N_VGND_c_325_n 0.0216143f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.385
cc_28 VNB N_VGND_c_326_n 0.00798243f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.295
cc_29 VNB N_VGND_c_327_n 0.0310594f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.385
cc_30 VNB N_VGND_c_328_n 0.0206731f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_329_n 0.220663f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_330_n 0.0100982f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VPB N_B_N_c_59_n 0.00355203f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.7
cc_34 VPB N_B_N_c_64_n 0.0205008f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.955
cc_35 VPB N_B_N_c_65_n 0.0317089f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.045
cc_36 VPB N_A_27_112#_c_100_n 0.0179198f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.21
cc_37 VPB N_A_27_112#_c_95_n 0.00906645f $X=-0.19 $Y=1.66 $X2=0.29 $Y2=1.385
cc_38 VPB N_A_27_112#_c_102_n 0.0433096f $X=-0.19 $Y=1.66 $X2=0.29 $Y2=1.385
cc_39 VPB N_A_27_112#_c_103_n 0.00235784f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_40 VPB N_A_27_112#_c_104_n 0.00979329f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_41 VPB N_A_27_112#_c_97_n 0.0104101f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_42 VPB N_A_c_163_n 0.0280754f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.54
cc_43 VPB N_A_c_164_n 0.00483912f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_44 VPB N_A_264_368#_c_194_n 0.0296995f $X=-0.19 $Y=1.66 $X2=0.565 $Y2=1.295
cc_45 VPB N_A_264_368#_c_201_n 0.0175967f $X=-0.19 $Y=1.66 $X2=0.29 $Y2=1.385
cc_46 VPB N_A_264_368#_c_197_n 0.00138341f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_47 VPB N_A_264_368#_c_203_n 0.00692132f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_48 VPB N_VPWR_c_263_n 0.0269547f $X=-0.19 $Y=1.66 $X2=0.88 $Y2=0.835
cc_49 VPB N_VPWR_c_264_n 0.0142675f $X=-0.19 $Y=1.66 $X2=0.36 $Y2=1.295
cc_50 VPB N_VPWR_c_265_n 0.0395991f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_51 VPB N_VPWR_c_266_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_52 VPB N_VPWR_c_267_n 0.0191515f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_53 VPB N_VPWR_c_268_n 0.0227588f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_54 VPB N_VPWR_c_262_n 0.0906352f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_55 VPB N_VPWR_c_270_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_56 VPB X 0.046779f $X=-0.19 $Y=1.66 $X2=0.36 $Y2=1.385
cc_57 VPB N_X_c_304_n 0.0203147f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_58 VPB N_X_c_302_n 0.00790788f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_59 N_B_N_c_61_n N_A_27_112#_M1000_g 0.00726223f $X=0.88 $Y=1.22 $X2=0 $Y2=0
cc_60 N_B_N_c_59_n N_A_27_112#_c_94_n 0.00307942f $X=0.505 $Y=1.7 $X2=0 $Y2=0
cc_61 N_B_N_c_60_n N_A_27_112#_c_94_n 0.00389289f $X=0.805 $Y=1.295 $X2=0 $Y2=0
cc_62 N_B_N_c_64_n N_A_27_112#_c_102_n 0.00147973f $X=0.505 $Y=1.955 $X2=0 $Y2=0
cc_63 N_B_N_c_65_n N_A_27_112#_c_102_n 0.022519f $X=0.505 $Y=2.045 $X2=0 $Y2=0
cc_64 N_B_N_c_64_n N_A_27_112#_c_103_n 0.0166765f $X=0.505 $Y=1.955 $X2=0 $Y2=0
cc_65 N_B_N_c_60_n N_A_27_112#_c_103_n 0.0019038f $X=0.805 $Y=1.295 $X2=0 $Y2=0
cc_66 B_N N_A_27_112#_c_103_n 5.214e-19 $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_67 N_B_N_c_59_n N_A_27_112#_c_104_n 0.00222782f $X=0.505 $Y=1.7 $X2=0 $Y2=0
cc_68 N_B_N_c_64_n N_A_27_112#_c_104_n 0.00438675f $X=0.505 $Y=1.955 $X2=0 $Y2=0
cc_69 B_N N_A_27_112#_c_104_n 0.0230941f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_70 N_B_N_c_61_n N_A_27_112#_c_117_n 0.00400158f $X=0.88 $Y=1.22 $X2=0 $Y2=0
cc_71 N_B_N_c_60_n N_A_27_112#_c_96_n 0.00871279f $X=0.805 $Y=1.295 $X2=0 $Y2=0
cc_72 N_B_N_c_61_n N_A_27_112#_c_96_n 0.00795326f $X=0.88 $Y=1.22 $X2=0 $Y2=0
cc_73 B_N N_A_27_112#_c_96_n 0.0237254f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_74 N_B_N_c_59_n N_A_27_112#_c_97_n 0.00954145f $X=0.505 $Y=1.7 $X2=0 $Y2=0
cc_75 N_B_N_c_64_n N_A_27_112#_c_97_n 0.00138205f $X=0.505 $Y=1.955 $X2=0 $Y2=0
cc_76 N_B_N_c_60_n N_A_27_112#_c_97_n 0.00620548f $X=0.805 $Y=1.295 $X2=0 $Y2=0
cc_77 N_B_N_c_60_n N_A_27_112#_c_98_n 0.0101512f $X=0.805 $Y=1.295 $X2=0 $Y2=0
cc_78 N_B_N_c_59_n N_A_27_112#_c_99_n 0.0102304f $X=0.505 $Y=1.7 $X2=0 $Y2=0
cc_79 B_N N_A_27_112#_c_99_n 0.0271897f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_80 N_B_N_c_65_n N_VPWR_c_263_n 0.0220538f $X=0.505 $Y=2.045 $X2=0 $Y2=0
cc_81 N_B_N_c_65_n N_VPWR_c_267_n 0.00445602f $X=0.505 $Y=2.045 $X2=0 $Y2=0
cc_82 N_B_N_c_65_n N_VPWR_c_262_n 0.00865213f $X=0.505 $Y=2.045 $X2=0 $Y2=0
cc_83 N_B_N_c_61_n N_VGND_c_323_n 0.0059966f $X=0.88 $Y=1.22 $X2=0 $Y2=0
cc_84 N_B_N_c_61_n N_VGND_c_327_n 0.00434478f $X=0.88 $Y=1.22 $X2=0 $Y2=0
cc_85 N_B_N_c_61_n N_VGND_c_329_n 0.00487769f $X=0.88 $Y=1.22 $X2=0 $Y2=0
cc_86 N_A_27_112#_M1000_g N_A_M1001_g 0.014193f $X=1.665 $Y=0.835 $X2=0 $Y2=0
cc_87 N_A_27_112#_c_100_n N_A_c_163_n 0.0524311f $X=1.69 $Y=1.765 $X2=0 $Y2=0
cc_88 N_A_27_112#_c_95_n N_A_c_163_n 0.0290208f $X=1.59 $Y=1.3 $X2=0 $Y2=0
cc_89 N_A_27_112#_c_95_n N_A_c_164_n 4.28628e-19 $X=1.59 $Y=1.3 $X2=0 $Y2=0
cc_90 N_A_27_112#_c_100_n N_A_264_368#_c_201_n 0.0164217f $X=1.69 $Y=1.765 $X2=0
+ $Y2=0
cc_91 N_A_27_112#_M1000_g N_A_264_368#_c_196_n 0.00744356f $X=1.665 $Y=0.835
+ $X2=0 $Y2=0
cc_92 N_A_27_112#_M1000_g N_A_264_368#_c_197_n 0.00575302f $X=1.665 $Y=0.835
+ $X2=0 $Y2=0
cc_93 N_A_27_112#_c_100_n N_A_264_368#_c_197_n 0.0029102f $X=1.69 $Y=1.765 $X2=0
+ $Y2=0
cc_94 N_A_27_112#_c_95_n N_A_264_368#_c_197_n 0.0163386f $X=1.59 $Y=1.3 $X2=0
+ $Y2=0
cc_95 N_A_27_112#_c_98_n N_A_264_368#_c_197_n 0.0250314f $X=1.36 $Y=1.465 $X2=0
+ $Y2=0
cc_96 N_A_27_112#_c_100_n N_A_264_368#_c_203_n 0.013567f $X=1.69 $Y=1.765 $X2=0
+ $Y2=0
cc_97 N_A_27_112#_c_94_n N_A_264_368#_c_203_n 0.00775559f $X=1.59 $Y=1.465 $X2=0
+ $Y2=0
cc_98 N_A_27_112#_c_95_n N_A_264_368#_c_203_n 8.37984e-19 $X=1.59 $Y=1.3 $X2=0
+ $Y2=0
cc_99 N_A_27_112#_c_97_n N_A_264_368#_c_203_n 0.00447704f $X=0.83 $Y=1.465 $X2=0
+ $Y2=0
cc_100 N_A_27_112#_c_98_n N_A_264_368#_c_203_n 0.0155529f $X=1.36 $Y=1.465 $X2=0
+ $Y2=0
cc_101 N_A_27_112#_M1000_g N_A_264_368#_c_199_n 0.0056446f $X=1.665 $Y=0.835
+ $X2=0 $Y2=0
cc_102 N_A_27_112#_c_100_n N_VPWR_c_263_n 0.0040491f $X=1.69 $Y=1.765 $X2=0
+ $Y2=0
cc_103 N_A_27_112#_c_102_n N_VPWR_c_263_n 0.0346007f $X=0.28 $Y=2.265 $X2=0
+ $Y2=0
cc_104 N_A_27_112#_c_103_n N_VPWR_c_263_n 0.00371626f $X=0.66 $Y=1.845 $X2=0
+ $Y2=0
cc_105 N_A_27_112#_c_97_n N_VPWR_c_263_n 0.0157412f $X=0.83 $Y=1.465 $X2=0 $Y2=0
cc_106 N_A_27_112#_c_98_n N_VPWR_c_263_n 0.00497979f $X=1.36 $Y=1.465 $X2=0
+ $Y2=0
cc_107 N_A_27_112#_c_100_n N_VPWR_c_265_n 0.00481995f $X=1.69 $Y=1.765 $X2=0
+ $Y2=0
cc_108 N_A_27_112#_c_102_n N_VPWR_c_267_n 0.0145938f $X=0.28 $Y=2.265 $X2=0
+ $Y2=0
cc_109 N_A_27_112#_c_100_n N_VPWR_c_262_n 0.00508379f $X=1.69 $Y=1.765 $X2=0
+ $Y2=0
cc_110 N_A_27_112#_c_102_n N_VPWR_c_262_n 0.0120466f $X=0.28 $Y=2.265 $X2=0
+ $Y2=0
cc_111 N_A_27_112#_M1000_g N_VGND_c_323_n 0.00735506f $X=1.665 $Y=0.835 $X2=0
+ $Y2=0
cc_112 N_A_27_112#_c_94_n N_VGND_c_323_n 0.00766427f $X=1.59 $Y=1.465 $X2=0
+ $Y2=0
cc_113 N_A_27_112#_c_96_n N_VGND_c_323_n 0.00488088f $X=0.745 $Y=1.3 $X2=0 $Y2=0
cc_114 N_A_27_112#_c_98_n N_VGND_c_323_n 0.0449072f $X=1.36 $Y=1.465 $X2=0 $Y2=0
cc_115 N_A_27_112#_M1000_g N_VGND_c_325_n 0.00418801f $X=1.665 $Y=0.835 $X2=0
+ $Y2=0
cc_116 N_A_27_112#_c_117_n N_VGND_c_327_n 0.00243801f $X=0.745 $Y=1.01 $X2=0
+ $Y2=0
cc_117 N_A_27_112#_c_99_n N_VGND_c_327_n 0.00905393f $X=0.665 $Y=0.845 $X2=0
+ $Y2=0
cc_118 N_A_27_112#_M1000_g N_VGND_c_329_n 0.00487769f $X=1.665 $Y=0.835 $X2=0
+ $Y2=0
cc_119 N_A_27_112#_c_117_n N_VGND_c_329_n 0.00494557f $X=0.745 $Y=1.01 $X2=0
+ $Y2=0
cc_120 N_A_27_112#_c_99_n N_VGND_c_329_n 0.0154532f $X=0.665 $Y=0.845 $X2=0
+ $Y2=0
cc_121 N_A_M1001_g N_A_264_368#_c_194_n 0.00113203f $X=2.095 $Y=0.835 $X2=0
+ $Y2=0
cc_122 N_A_c_163_n N_A_264_368#_c_194_n 0.043529f $X=2.11 $Y=1.765 $X2=0 $Y2=0
cc_123 N_A_c_164_n N_A_264_368#_c_194_n 0.00292422f $X=2.2 $Y=1.515 $X2=0 $Y2=0
cc_124 N_A_M1001_g N_A_264_368#_M1007_g 0.0127273f $X=2.095 $Y=0.835 $X2=0 $Y2=0
cc_125 N_A_c_163_n N_A_264_368#_c_201_n 0.00259875f $X=2.11 $Y=1.765 $X2=0 $Y2=0
cc_126 N_A_M1001_g N_A_264_368#_c_196_n 0.0124806f $X=2.095 $Y=0.835 $X2=0 $Y2=0
cc_127 N_A_M1001_g N_A_264_368#_c_197_n 0.00428454f $X=2.095 $Y=0.835 $X2=0
+ $Y2=0
cc_128 N_A_c_163_n N_A_264_368#_c_197_n 9.01058e-19 $X=2.11 $Y=1.765 $X2=0 $Y2=0
cc_129 N_A_c_164_n N_A_264_368#_c_197_n 0.0322792f $X=2.2 $Y=1.515 $X2=0 $Y2=0
cc_130 N_A_M1001_g N_A_264_368#_c_198_n 0.013594f $X=2.095 $Y=0.835 $X2=0 $Y2=0
cc_131 N_A_c_163_n N_A_264_368#_c_198_n 0.00309794f $X=2.11 $Y=1.765 $X2=0 $Y2=0
cc_132 N_A_c_164_n N_A_264_368#_c_198_n 0.0466983f $X=2.2 $Y=1.515 $X2=0 $Y2=0
cc_133 N_A_c_163_n N_A_264_368#_c_203_n 0.00373365f $X=2.11 $Y=1.765 $X2=0 $Y2=0
cc_134 N_A_M1001_g N_A_264_368#_c_199_n 0.00300021f $X=2.095 $Y=0.835 $X2=0
+ $Y2=0
cc_135 N_A_c_164_n N_A_264_368#_c_199_n 7.33087e-19 $X=2.2 $Y=1.515 $X2=0 $Y2=0
cc_136 N_A_c_163_n N_VPWR_c_264_n 0.0177334f $X=2.11 $Y=1.765 $X2=0 $Y2=0
cc_137 N_A_c_164_n N_VPWR_c_264_n 0.00959142f $X=2.2 $Y=1.515 $X2=0 $Y2=0
cc_138 N_A_c_163_n N_VPWR_c_265_n 0.0049405f $X=2.11 $Y=1.765 $X2=0 $Y2=0
cc_139 N_A_c_163_n N_VPWR_c_262_n 0.00508379f $X=2.11 $Y=1.765 $X2=0 $Y2=0
cc_140 N_A_c_163_n N_X_c_304_n 7.65008e-19 $X=2.11 $Y=1.765 $X2=0 $Y2=0
cc_141 N_A_M1001_g N_VGND_c_324_n 0.00665253f $X=2.095 $Y=0.835 $X2=0 $Y2=0
cc_142 N_A_M1001_g N_VGND_c_325_n 0.0043356f $X=2.095 $Y=0.835 $X2=0 $Y2=0
cc_143 N_A_M1001_g N_VGND_c_329_n 0.00487769f $X=2.095 $Y=0.835 $X2=0 $Y2=0
cc_144 N_A_264_368#_c_201_n N_VPWR_c_263_n 0.0380372f $X=1.465 $Y=2.695 $X2=0
+ $Y2=0
cc_145 N_A_264_368#_c_194_n N_VPWR_c_264_n 0.0114591f $X=2.695 $Y=1.765 $X2=0
+ $Y2=0
cc_146 N_A_264_368#_c_201_n N_VPWR_c_264_n 0.0241168f $X=1.465 $Y=2.695 $X2=0
+ $Y2=0
cc_147 N_A_264_368#_c_198_n N_VPWR_c_264_n 0.0022447f $X=2.535 $Y=1.095 $X2=0
+ $Y2=0
cc_148 N_A_264_368#_c_203_n N_VPWR_c_264_n 0.00177012f $X=1.78 $Y=1.905 $X2=0
+ $Y2=0
cc_149 N_A_264_368#_c_201_n N_VPWR_c_265_n 0.0097982f $X=1.465 $Y=2.695 $X2=0
+ $Y2=0
cc_150 N_A_264_368#_c_194_n N_VPWR_c_268_n 0.00445602f $X=2.695 $Y=1.765 $X2=0
+ $Y2=0
cc_151 N_A_264_368#_c_194_n N_VPWR_c_262_n 0.00865635f $X=2.695 $Y=1.765 $X2=0
+ $Y2=0
cc_152 N_A_264_368#_c_201_n N_VPWR_c_262_n 0.0111907f $X=1.465 $Y=2.695 $X2=0
+ $Y2=0
cc_153 N_A_264_368#_c_203_n A_353_368# 0.00359365f $X=1.78 $Y=1.905 $X2=-0.19
+ $Y2=-0.245
cc_154 N_A_264_368#_M1007_g N_X_c_300_n 0.0113949f $X=2.825 $Y=0.74 $X2=0 $Y2=0
cc_155 N_A_264_368#_c_194_n N_X_c_301_n 2.77016e-19 $X=2.695 $Y=1.765 $X2=0
+ $Y2=0
cc_156 N_A_264_368#_M1007_g N_X_c_301_n 0.00556841f $X=2.825 $Y=0.74 $X2=0 $Y2=0
cc_157 N_A_264_368#_c_198_n N_X_c_301_n 0.0104368f $X=2.535 $Y=1.095 $X2=0 $Y2=0
cc_158 N_A_264_368#_c_194_n X 0.0103749f $X=2.695 $Y=1.765 $X2=0 $Y2=0
cc_159 N_A_264_368#_c_194_n N_X_c_304_n 0.00624725f $X=2.695 $Y=1.765 $X2=0
+ $Y2=0
cc_160 N_A_264_368#_c_198_n N_X_c_304_n 0.0138812f $X=2.535 $Y=1.095 $X2=0 $Y2=0
cc_161 N_A_264_368#_c_194_n N_X_c_302_n 0.00647696f $X=2.695 $Y=1.765 $X2=0
+ $Y2=0
cc_162 N_A_264_368#_M1007_g N_X_c_302_n 0.00246301f $X=2.825 $Y=0.74 $X2=0 $Y2=0
cc_163 N_A_264_368#_c_198_n N_X_c_302_n 0.0302873f $X=2.535 $Y=1.095 $X2=0 $Y2=0
cc_164 N_A_264_368#_c_198_n N_VGND_M1001_d 0.00843341f $X=2.535 $Y=1.095 $X2=0
+ $Y2=0
cc_165 N_A_264_368#_c_196_n N_VGND_c_323_n 0.0379888f $X=1.88 $Y=0.835 $X2=0
+ $Y2=0
cc_166 N_A_264_368#_c_199_n N_VGND_c_323_n 0.0102677f $X=1.87 $Y=1.095 $X2=0
+ $Y2=0
cc_167 N_A_264_368#_c_194_n N_VGND_c_324_n 3.08957e-19 $X=2.695 $Y=1.765 $X2=0
+ $Y2=0
cc_168 N_A_264_368#_M1007_g N_VGND_c_324_n 0.0110504f $X=2.825 $Y=0.74 $X2=0
+ $Y2=0
cc_169 N_A_264_368#_c_196_n N_VGND_c_324_n 0.0195637f $X=1.88 $Y=0.835 $X2=0
+ $Y2=0
cc_170 N_A_264_368#_c_198_n N_VGND_c_324_n 0.0347439f $X=2.535 $Y=1.095 $X2=0
+ $Y2=0
cc_171 N_A_264_368#_c_196_n N_VGND_c_325_n 0.00852231f $X=1.88 $Y=0.835 $X2=0
+ $Y2=0
cc_172 N_A_264_368#_M1007_g N_VGND_c_328_n 0.00434272f $X=2.825 $Y=0.74 $X2=0
+ $Y2=0
cc_173 N_A_264_368#_M1007_g N_VGND_c_329_n 0.00829406f $X=2.825 $Y=0.74 $X2=0
+ $Y2=0
cc_174 N_A_264_368#_c_196_n N_VGND_c_329_n 0.0112256f $X=1.88 $Y=0.835 $X2=0
+ $Y2=0
cc_175 N_VPWR_c_268_n X 0.0230718f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_176 N_VPWR_c_262_n X 0.0190639f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_177 N_VPWR_c_264_n N_X_c_304_n 0.0421814f $X=2.42 $Y=2.115 $X2=0 $Y2=0
cc_178 N_X_c_300_n N_VGND_c_324_n 0.0353629f $X=3.04 $Y=0.515 $X2=0 $Y2=0
cc_179 N_X_c_300_n N_VGND_c_328_n 0.0176874f $X=3.04 $Y=0.515 $X2=0 $Y2=0
cc_180 N_X_c_300_n N_VGND_c_329_n 0.0145837f $X=3.04 $Y=0.515 $X2=0 $Y2=0
