* File: sky130_fd_sc_hs__buf_8.pex.spice
* Created: Thu Aug 27 20:34:42 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HS__BUF_8%A 3 5 7 8 10 13 17 19 21 22 23 24 37 38
r67 38 39 1.2957 $w=3.72e-07 $l=1e-08 $layer=POLY_cond $X=1.4 $Y=1.557 $X2=1.41
+ $Y2=1.557
r68 36 38 17.4919 $w=3.72e-07 $l=1.35e-07 $layer=POLY_cond $X=1.265 $Y=1.557
+ $X2=1.4 $Y2=1.557
r69 36 37 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.265
+ $Y=1.515 $X2=1.265 $Y2=1.515
r70 34 36 38.2231 $w=3.72e-07 $l=2.95e-07 $layer=POLY_cond $X=0.97 $Y=1.557
+ $X2=1.265 $Y2=1.557
r71 33 34 1.2957 $w=3.72e-07 $l=1e-08 $layer=POLY_cond $X=0.96 $Y=1.557 $X2=0.97
+ $Y2=1.557
r72 31 33 48.5887 $w=3.72e-07 $l=3.75e-07 $layer=POLY_cond $X=0.585 $Y=1.557
+ $X2=0.96 $Y2=1.557
r73 31 32 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=0.585
+ $Y=1.515 $X2=0.585 $Y2=1.515
r74 29 31 9.71774 $w=3.72e-07 $l=7.5e-08 $layer=POLY_cond $X=0.51 $Y=1.557
+ $X2=0.585 $Y2=1.557
r75 28 29 1.94355 $w=3.72e-07 $l=1.5e-08 $layer=POLY_cond $X=0.495 $Y=1.557
+ $X2=0.51 $Y2=1.557
r76 24 37 1.74206 $w=4.28e-07 $l=6.5e-08 $layer=LI1_cond $X=1.2 $Y=1.565
+ $X2=1.265 $Y2=1.565
r77 23 24 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=0.72 $Y=1.565
+ $X2=1.2 $Y2=1.565
r78 23 32 3.61813 $w=4.28e-07 $l=1.35e-07 $layer=LI1_cond $X=0.72 $Y=1.565
+ $X2=0.585 $Y2=1.565
r79 22 32 9.24634 $w=4.28e-07 $l=3.45e-07 $layer=LI1_cond $X=0.24 $Y=1.565
+ $X2=0.585 $Y2=1.565
r80 19 39 24.0971 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=1.41 $Y=1.765
+ $X2=1.41 $Y2=1.557
r81 19 21 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.41 $Y=1.765
+ $X2=1.41 $Y2=2.4
r82 15 38 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.4 $Y=1.35 $X2=1.4
+ $Y2=1.557
r83 15 17 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.4 $Y=1.35 $X2=1.4
+ $Y2=0.74
r84 11 34 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.97 $Y=1.35
+ $X2=0.97 $Y2=1.557
r85 11 13 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=0.97 $Y=1.35
+ $X2=0.97 $Y2=0.74
r86 8 33 24.0971 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=0.96 $Y=1.765
+ $X2=0.96 $Y2=1.557
r87 8 10 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.96 $Y=1.765
+ $X2=0.96 $Y2=2.4
r88 5 29 24.0971 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=0.51 $Y=1.765
+ $X2=0.51 $Y2=1.557
r89 5 7 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.51 $Y=1.765
+ $X2=0.51 $Y2=2.4
r90 1 28 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.495 $Y=1.35
+ $X2=0.495 $Y2=1.557
r91 1 3 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=0.495 $Y=1.35
+ $X2=0.495 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HS__BUF_8%A_27_74# 1 2 3 4 15 17 19 22 24 26 29 31 33 36
+ 38 40 43 45 47 50 52 54 55 57 60 64 66 68 71 73 75 77 78 79 83 87 89 91 94 100
+ 106 107 108 127
c231 15 0 1.65559e-19 $X=1.83 $Y=0.74
r232 127 128 1.88281 $w=3.84e-07 $l=1.5e-08 $layer=POLY_cond $X=5.195 $Y=1.532
+ $X2=5.21 $Y2=1.532
r233 126 127 54.6016 $w=3.84e-07 $l=4.35e-07 $layer=POLY_cond $X=4.76 $Y=1.532
+ $X2=5.195 $Y2=1.532
r234 125 126 1.88281 $w=3.84e-07 $l=1.5e-08 $layer=POLY_cond $X=4.745 $Y=1.532
+ $X2=4.76 $Y2=1.532
r235 122 123 8.78646 $w=3.84e-07 $l=7e-08 $layer=POLY_cond $X=4.19 $Y=1.532
+ $X2=4.26 $Y2=1.532
r236 121 122 47.6979 $w=3.84e-07 $l=3.8e-07 $layer=POLY_cond $X=3.81 $Y=1.532
+ $X2=4.19 $Y2=1.532
r237 120 121 6.27604 $w=3.84e-07 $l=5e-08 $layer=POLY_cond $X=3.76 $Y=1.532
+ $X2=3.81 $Y2=1.532
r238 119 120 56.4844 $w=3.84e-07 $l=4.5e-07 $layer=POLY_cond $X=3.31 $Y=1.532
+ $X2=3.76 $Y2=1.532
r239 118 119 15.0625 $w=3.84e-07 $l=1.2e-07 $layer=POLY_cond $X=3.19 $Y=1.532
+ $X2=3.31 $Y2=1.532
r240 117 118 41.4219 $w=3.84e-07 $l=3.3e-07 $layer=POLY_cond $X=2.86 $Y=1.532
+ $X2=3.19 $Y2=1.532
r241 116 117 12.5521 $w=3.84e-07 $l=1e-07 $layer=POLY_cond $X=2.76 $Y=1.532
+ $X2=2.86 $Y2=1.532
r242 115 116 50.2083 $w=3.84e-07 $l=4e-07 $layer=POLY_cond $X=2.36 $Y=1.532
+ $X2=2.76 $Y2=1.532
r243 114 115 12.5521 $w=3.84e-07 $l=1e-07 $layer=POLY_cond $X=2.26 $Y=1.532
+ $X2=2.36 $Y2=1.532
r244 111 112 3.76562 $w=3.84e-07 $l=3e-08 $layer=POLY_cond $X=1.83 $Y=1.532
+ $X2=1.86 $Y2=1.532
r245 101 125 13.1797 $w=3.84e-07 $l=1.05e-07 $layer=POLY_cond $X=4.64 $Y=1.532
+ $X2=4.745 $Y2=1.532
r246 101 123 47.6979 $w=3.84e-07 $l=3.8e-07 $layer=POLY_cond $X=4.64 $Y=1.532
+ $X2=4.26 $Y2=1.532
r247 100 101 32.2844 $w=1.7e-07 $l=7.65e-07 $layer=licon1_POLY $count=4 $X=4.64
+ $Y=1.465 $X2=4.64 $Y2=1.465
r248 98 114 42.6771 $w=3.84e-07 $l=3.4e-07 $layer=POLY_cond $X=1.92 $Y=1.532
+ $X2=2.26 $Y2=1.532
r249 98 112 7.53125 $w=3.84e-07 $l=6e-08 $layer=POLY_cond $X=1.92 $Y=1.532
+ $X2=1.86 $Y2=1.532
r250 97 100 94.9892 $w=3.28e-07 $l=2.72e-06 $layer=LI1_cond $X=1.92 $Y=1.465
+ $X2=4.64 $Y2=1.465
r251 97 98 32.2844 $w=1.7e-07 $l=7.65e-07 $layer=licon1_POLY $count=4 $X=1.92
+ $Y=1.465 $X2=1.92 $Y2=1.465
r252 95 108 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=1.685 $Y=1.465
+ $X2=1.685 $Y2=1.095
r253 95 97 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=1.77 $Y=1.465
+ $X2=1.92 $Y2=1.465
r254 93 95 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=1.685 $Y=1.63
+ $X2=1.685 $Y2=1.465
r255 93 94 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=1.685 $Y=1.63
+ $X2=1.685 $Y2=1.95
r256 92 106 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.35 $Y=2.035
+ $X2=1.185 $Y2=2.035
r257 91 94 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.6 $Y=2.035
+ $X2=1.685 $Y2=1.95
r258 91 92 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=1.6 $Y=2.035
+ $X2=1.35 $Y2=2.035
r259 90 107 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.27 $Y=1.095
+ $X2=1.185 $Y2=1.095
r260 89 108 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.6 $Y=1.095
+ $X2=1.685 $Y2=1.095
r261 89 90 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=1.6 $Y=1.095
+ $X2=1.27 $Y2=1.095
r262 85 107 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.185 $Y=1.01
+ $X2=1.185 $Y2=1.095
r263 85 87 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=1.185 $Y=1.01
+ $X2=1.185 $Y2=0.515
r264 81 106 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.185 $Y=2.12
+ $X2=1.185 $Y2=2.035
r265 81 83 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=1.185 $Y=2.12
+ $X2=1.185 $Y2=2.815
r266 80 104 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.45 $Y=2.035
+ $X2=0.285 $Y2=2.035
r267 79 106 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.02 $Y=2.035
+ $X2=1.185 $Y2=2.035
r268 79 80 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=1.02 $Y=2.035
+ $X2=0.45 $Y2=2.035
r269 77 107 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.1 $Y=1.095
+ $X2=1.185 $Y2=1.095
r270 77 78 47.9519 $w=1.68e-07 $l=7.35e-07 $layer=LI1_cond $X=1.1 $Y=1.095
+ $X2=0.365 $Y2=1.095
r271 73 104 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.285 $Y=2.12
+ $X2=0.285 $Y2=2.035
r272 73 75 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=0.285 $Y=2.12
+ $X2=0.285 $Y2=2.815
r273 69 78 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.24 $Y=1.01
+ $X2=0.365 $Y2=1.095
r274 69 71 22.8184 $w=2.48e-07 $l=4.95e-07 $layer=LI1_cond $X=0.24 $Y=1.01
+ $X2=0.24 $Y2=0.515
r275 66 128 24.8669 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=5.21 $Y=1.765
+ $X2=5.21 $Y2=1.532
r276 66 68 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=5.21 $Y=1.765
+ $X2=5.21 $Y2=2.4
r277 62 127 24.8669 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=5.195 $Y=1.3
+ $X2=5.195 $Y2=1.532
r278 62 64 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=5.195 $Y=1.3
+ $X2=5.195 $Y2=0.74
r279 58 126 24.8669 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=4.76 $Y=1.3
+ $X2=4.76 $Y2=1.532
r280 58 60 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=4.76 $Y=1.3
+ $X2=4.76 $Y2=0.74
r281 55 125 24.8669 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=4.745 $Y=1.765
+ $X2=4.745 $Y2=1.532
r282 55 57 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=4.745 $Y=1.765
+ $X2=4.745 $Y2=2.4
r283 52 123 24.8669 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=4.26 $Y=1.765
+ $X2=4.26 $Y2=1.532
r284 52 54 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=4.26 $Y=1.765
+ $X2=4.26 $Y2=2.4
r285 48 122 24.8669 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=4.19 $Y=1.3
+ $X2=4.19 $Y2=1.532
r286 48 50 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=4.19 $Y=1.3
+ $X2=4.19 $Y2=0.74
r287 45 121 24.8669 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=3.81 $Y=1.765
+ $X2=3.81 $Y2=1.532
r288 45 47 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.81 $Y=1.765
+ $X2=3.81 $Y2=2.4
r289 41 120 24.8669 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=3.76 $Y=1.3
+ $X2=3.76 $Y2=1.532
r290 41 43 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=3.76 $Y=1.3
+ $X2=3.76 $Y2=0.74
r291 38 119 24.8669 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=3.31 $Y=1.765
+ $X2=3.31 $Y2=1.532
r292 38 40 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.31 $Y=1.765
+ $X2=3.31 $Y2=2.4
r293 34 118 24.8669 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=3.19 $Y=1.3
+ $X2=3.19 $Y2=1.532
r294 34 36 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=3.19 $Y=1.3
+ $X2=3.19 $Y2=0.74
r295 31 117 24.8669 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=2.86 $Y=1.765
+ $X2=2.86 $Y2=1.532
r296 31 33 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.86 $Y=1.765
+ $X2=2.86 $Y2=2.4
r297 27 116 24.8669 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=2.76 $Y=1.3
+ $X2=2.76 $Y2=1.532
r298 27 29 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=2.76 $Y=1.3
+ $X2=2.76 $Y2=0.74
r299 24 115 24.8669 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=2.36 $Y=1.765
+ $X2=2.36 $Y2=1.532
r300 24 26 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.36 $Y=1.765
+ $X2=2.36 $Y2=2.4
r301 20 114 24.8669 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=2.26 $Y=1.3
+ $X2=2.26 $Y2=1.532
r302 20 22 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=2.26 $Y=1.3
+ $X2=2.26 $Y2=0.74
r303 17 112 24.8669 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=1.86 $Y=1.765
+ $X2=1.86 $Y2=1.532
r304 17 19 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.86 $Y=1.765
+ $X2=1.86 $Y2=2.4
r305 13 111 24.8669 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=1.83 $Y=1.3
+ $X2=1.83 $Y2=1.532
r306 13 15 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=1.83 $Y=1.3
+ $X2=1.83 $Y2=0.74
r307 4 106 400 $w=1.7e-07 $l=3.4187e-07 $layer=licon1_PDIFF $count=1 $X=1.035
+ $Y=1.84 $X2=1.185 $Y2=2.115
r308 4 83 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=1.035
+ $Y=1.84 $X2=1.185 $Y2=2.815
r309 3 104 400 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_PDIFF $count=1 $X=0.14
+ $Y=1.84 $X2=0.285 $Y2=2.115
r310 3 75 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=0.14
+ $Y=1.84 $X2=0.285 $Y2=2.815
r311 2 87 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.045
+ $Y=0.37 $X2=1.185 $Y2=0.515
r312 1 71 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__BUF_8%VPWR 1 2 3 4 5 6 23 27 31 35 39 41 43 47 49 54
+ 59 64 69 75 78 81 84 87 91
r89 90 91 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r90 87 88 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r91 84 85 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r92 81 82 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r93 78 79 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r94 75 76 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r95 73 91 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=5.52 $Y2=3.33
r96 73 88 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=4.56 $Y2=3.33
r97 72 73 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r98 70 87 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.65 $Y=3.33
+ $X2=4.525 $Y2=3.33
r99 70 72 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=4.65 $Y=3.33
+ $X2=5.04 $Y2=3.33
r100 69 90 3.9577 $w=1.7e-07 $l=2.05e-07 $layer=LI1_cond $X=5.35 $Y=3.33
+ $X2=5.555 $Y2=3.33
r101 69 72 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=5.35 $Y=3.33
+ $X2=5.04 $Y2=3.33
r102 68 88 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=4.56 $Y2=3.33
r103 68 85 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=3.6 $Y2=3.33
r104 67 68 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r105 65 84 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.7 $Y=3.33
+ $X2=3.575 $Y2=3.33
r106 65 67 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=3.7 $Y=3.33
+ $X2=4.08 $Y2=3.33
r107 64 87 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.4 $Y=3.33
+ $X2=4.525 $Y2=3.33
r108 64 67 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=4.4 $Y=3.33 $X2=4.08
+ $Y2=3.33
r109 63 85 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=3.6 $Y2=3.33
r110 62 63 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r111 60 81 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.75 $Y=3.33
+ $X2=2.625 $Y2=3.33
r112 60 62 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=2.75 $Y=3.33
+ $X2=3.12 $Y2=3.33
r113 59 84 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.45 $Y=3.33
+ $X2=3.575 $Y2=3.33
r114 59 62 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=3.45 $Y=3.33
+ $X2=3.12 $Y2=3.33
r115 58 82 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r116 58 79 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.68 $Y2=3.33
r117 57 58 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r118 55 78 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.8 $Y=3.33
+ $X2=1.675 $Y2=3.33
r119 55 57 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=1.8 $Y=3.33
+ $X2=2.16 $Y2=3.33
r120 54 81 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.5 $Y=3.33
+ $X2=2.625 $Y2=3.33
r121 54 57 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=2.5 $Y=3.33
+ $X2=2.16 $Y2=3.33
r122 53 79 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=1.68 $Y2=3.33
r123 53 76 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r124 52 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r125 50 75 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.82 $Y=3.33
+ $X2=0.735 $Y2=3.33
r126 50 52 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=0.82 $Y=3.33
+ $X2=1.2 $Y2=3.33
r127 49 78 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.55 $Y=3.33
+ $X2=1.675 $Y2=3.33
r128 49 52 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=1.55 $Y=3.33
+ $X2=1.2 $Y2=3.33
r129 47 63 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.88 $Y=3.33
+ $X2=3.12 $Y2=3.33
r130 47 82 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.88 $Y=3.33
+ $X2=2.64 $Y2=3.33
r131 43 46 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=5.475 $Y=1.985
+ $X2=5.475 $Y2=2.815
r132 41 90 3.18546 $w=2.5e-07 $l=1.18427e-07 $layer=LI1_cond $X=5.475 $Y=3.245
+ $X2=5.555 $Y2=3.33
r133 41 46 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=5.475 $Y=3.245
+ $X2=5.475 $Y2=2.815
r134 37 87 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.525 $Y=3.245
+ $X2=4.525 $Y2=3.33
r135 37 39 43.3319 $w=2.48e-07 $l=9.4e-07 $layer=LI1_cond $X=4.525 $Y=3.245
+ $X2=4.525 $Y2=2.305
r136 33 84 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.575 $Y=3.245
+ $X2=3.575 $Y2=3.33
r137 33 35 43.3319 $w=2.48e-07 $l=9.4e-07 $layer=LI1_cond $X=3.575 $Y=3.245
+ $X2=3.575 $Y2=2.305
r138 29 81 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.625 $Y=3.245
+ $X2=2.625 $Y2=3.33
r139 29 31 43.3319 $w=2.48e-07 $l=9.4e-07 $layer=LI1_cond $X=2.625 $Y=3.245
+ $X2=2.625 $Y2=2.305
r140 25 78 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.675 $Y=3.245
+ $X2=1.675 $Y2=3.33
r141 25 27 36.4172 $w=2.48e-07 $l=7.9e-07 $layer=LI1_cond $X=1.675 $Y=3.245
+ $X2=1.675 $Y2=2.455
r142 21 75 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.735 $Y=3.245
+ $X2=0.735 $Y2=3.33
r143 21 23 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=0.735 $Y=3.245
+ $X2=0.735 $Y2=2.455
r144 6 46 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=5.285
+ $Y=1.84 $X2=5.435 $Y2=2.815
r145 6 43 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=5.285
+ $Y=1.84 $X2=5.435 $Y2=1.985
r146 5 39 300 $w=1.7e-07 $l=5.34766e-07 $layer=licon1_PDIFF $count=2 $X=4.335
+ $Y=1.84 $X2=4.485 $Y2=2.305
r147 4 35 300 $w=1.7e-07 $l=5.34766e-07 $layer=licon1_PDIFF $count=2 $X=3.385
+ $Y=1.84 $X2=3.535 $Y2=2.305
r148 3 31 300 $w=1.7e-07 $l=5.34766e-07 $layer=licon1_PDIFF $count=2 $X=2.435
+ $Y=1.84 $X2=2.585 $Y2=2.305
r149 2 27 300 $w=1.7e-07 $l=6.85912e-07 $layer=licon1_PDIFF $count=2 $X=1.485
+ $Y=1.84 $X2=1.635 $Y2=2.455
r150 1 23 300 $w=1.7e-07 $l=6.85912e-07 $layer=licon1_PDIFF $count=2 $X=0.585
+ $Y=1.84 $X2=0.735 $Y2=2.455
.ends

.subckt PM_SKY130_FD_SC_HS__BUF_8%X 1 2 3 4 5 6 7 8 27 31 35 36 37 38 41 45 49
+ 51 55 59 63 65 69 72 73 74 75 76 77 78 79 80 88
c155 36 0 1.65559e-19 $X=2.13 $Y=1.045
r156 85 88 0.516019 $w=3.33e-07 $l=1.5e-08 $layer=LI1_cond $X=4.987 $Y=1.97
+ $X2=4.987 $Y2=1.985
r157 79 80 12.7285 $w=3.33e-07 $l=3.7e-07 $layer=LI1_cond $X=4.987 $Y=2.405
+ $X2=4.987 $Y2=2.775
r158 78 85 3.67481 $w=2.52e-07 $l=8.5e-08 $layer=LI1_cond $X=4.987 $Y=1.885
+ $X2=4.987 $Y2=1.97
r159 78 79 12.3845 $w=3.33e-07 $l=3.6e-07 $layer=LI1_cond $X=4.987 $Y=2.045
+ $X2=4.987 $Y2=2.405
r160 78 88 2.06408 $w=3.33e-07 $l=6e-08 $layer=LI1_cond $X=4.987 $Y=2.045
+ $X2=4.987 $Y2=1.985
r161 72 78 3.67481 $w=2.52e-07 $l=1.15888e-07 $layer=LI1_cond $X=5.06 $Y=1.8
+ $X2=4.987 $Y2=1.885
r162 71 77 3.67481 $w=2.52e-07 $l=1.19499e-07 $layer=LI1_cond $X=5.06 $Y=1.13
+ $X2=4.977 $Y2=1.045
r163 71 72 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.06 $Y=1.13
+ $X2=5.06 $Y2=1.8
r164 67 77 3.67481 $w=2.52e-07 $l=8.5e-08 $layer=LI1_cond $X=4.977 $Y=0.96
+ $X2=4.977 $Y2=1.045
r165 67 69 15.3086 $w=3.33e-07 $l=4.45e-07 $layer=LI1_cond $X=4.977 $Y=0.96
+ $X2=4.977 $Y2=0.515
r166 66 76 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.2 $Y=1.885
+ $X2=4.035 $Y2=1.885
r167 65 78 2.79892 $w=1.7e-07 $l=1.67e-07 $layer=LI1_cond $X=4.82 $Y=1.885
+ $X2=4.987 $Y2=1.885
r168 65 66 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=4.82 $Y=1.885
+ $X2=4.2 $Y2=1.885
r169 64 75 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.14 $Y=1.045
+ $X2=3.975 $Y2=1.045
r170 63 77 2.79892 $w=1.7e-07 $l=1.67e-07 $layer=LI1_cond $X=4.81 $Y=1.045
+ $X2=4.977 $Y2=1.045
r171 63 64 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.81 $Y=1.045
+ $X2=4.14 $Y2=1.045
r172 59 61 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=4.035 $Y=1.985
+ $X2=4.035 $Y2=2.815
r173 57 76 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.035 $Y=1.97
+ $X2=4.035 $Y2=1.885
r174 57 59 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=4.035 $Y=1.97
+ $X2=4.035 $Y2=1.985
r175 53 75 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.975 $Y=0.96
+ $X2=3.975 $Y2=1.045
r176 53 55 15.5405 $w=3.28e-07 $l=4.45e-07 $layer=LI1_cond $X=3.975 $Y=0.96
+ $X2=3.975 $Y2=0.515
r177 52 74 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.25 $Y=1.885
+ $X2=3.085 $Y2=1.885
r178 51 76 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.87 $Y=1.885
+ $X2=4.035 $Y2=1.885
r179 51 52 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=3.87 $Y=1.885
+ $X2=3.25 $Y2=1.885
r180 50 73 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.14 $Y=1.045
+ $X2=2.975 $Y2=1.045
r181 49 75 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.81 $Y=1.045
+ $X2=3.975 $Y2=1.045
r182 49 50 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.81 $Y=1.045
+ $X2=3.14 $Y2=1.045
r183 45 47 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=3.085 $Y=1.985
+ $X2=3.085 $Y2=2.815
r184 43 74 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.085 $Y=1.97
+ $X2=3.085 $Y2=1.885
r185 43 45 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=3.085 $Y=1.97
+ $X2=3.085 $Y2=1.985
r186 39 73 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.975 $Y=0.96
+ $X2=2.975 $Y2=1.045
r187 39 41 15.5405 $w=3.28e-07 $l=4.45e-07 $layer=LI1_cond $X=2.975 $Y=0.96
+ $X2=2.975 $Y2=0.515
r188 37 74 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.92 $Y=1.885
+ $X2=3.085 $Y2=1.885
r189 37 38 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=2.92 $Y=1.885
+ $X2=2.3 $Y2=1.885
r190 35 73 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.81 $Y=1.045
+ $X2=2.975 $Y2=1.045
r191 35 36 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=2.81 $Y=1.045
+ $X2=2.13 $Y2=1.045
r192 31 33 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=2.135 $Y=1.985
+ $X2=2.135 $Y2=2.815
r193 29 38 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.135 $Y=1.97
+ $X2=2.3 $Y2=1.885
r194 29 31 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=2.135 $Y=1.97
+ $X2=2.135 $Y2=1.985
r195 25 36 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.045 $Y=0.96
+ $X2=2.13 $Y2=1.045
r196 25 27 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=2.045 $Y=0.96
+ $X2=2.045 $Y2=0.515
r197 8 80 400 $w=1.7e-07 $l=1.05428e-06 $layer=licon1_PDIFF $count=1 $X=4.82
+ $Y=1.84 $X2=4.985 $Y2=2.815
r198 8 88 400 $w=1.7e-07 $l=2.26164e-07 $layer=licon1_PDIFF $count=1 $X=4.82
+ $Y=1.84 $X2=4.985 $Y2=1.985
r199 7 61 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=3.885
+ $Y=1.84 $X2=4.035 $Y2=2.815
r200 7 59 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=3.885
+ $Y=1.84 $X2=4.035 $Y2=1.985
r201 6 47 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=2.935
+ $Y=1.84 $X2=3.085 $Y2=2.815
r202 6 45 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=2.935
+ $Y=1.84 $X2=3.085 $Y2=1.985
r203 5 33 400 $w=1.7e-07 $l=1.07034e-06 $layer=licon1_PDIFF $count=1 $X=1.935
+ $Y=1.84 $X2=2.135 $Y2=2.815
r204 5 31 400 $w=1.7e-07 $l=2.62678e-07 $layer=licon1_PDIFF $count=1 $X=1.935
+ $Y=1.84 $X2=2.135 $Y2=1.985
r205 4 69 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=4.835
+ $Y=0.37 $X2=4.975 $Y2=0.515
r206 3 55 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.835
+ $Y=0.37 $X2=3.975 $Y2=0.515
r207 2 41 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.835
+ $Y=0.37 $X2=2.975 $Y2=0.515
r208 1 27 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.905
+ $Y=0.37 $X2=2.045 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__BUF_8%VGND 1 2 3 4 5 6 21 25 29 33 37 39 41 44 45 47
+ 48 50 51 52 54 59 74 79 82 86
r92 85 86 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r93 82 83 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r94 79 80 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r95 77 86 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=5.52
+ $Y2=0
r96 76 77 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r97 74 85 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=5.315 $Y=0 $X2=5.537
+ $Y2=0
r98 74 76 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=5.315 $Y=0 $X2=5.04
+ $Y2=0
r99 73 77 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=5.04
+ $Y2=0
r100 72 73 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r101 70 73 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=4.08
+ $Y2=0
r102 69 70 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r103 67 83 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.68
+ $Y2=0
r104 66 67 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r105 64 82 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.78 $Y=0 $X2=1.615
+ $Y2=0
r106 64 66 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=1.78 $Y=0 $X2=2.16
+ $Y2=0
r107 63 83 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=1.68
+ $Y2=0
r108 63 80 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r109 62 63 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r110 60 79 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.875 $Y=0 $X2=0.71
+ $Y2=0
r111 60 62 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.875 $Y=0 $X2=1.2
+ $Y2=0
r112 59 82 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.45 $Y=0 $X2=1.615
+ $Y2=0
r113 59 62 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=1.45 $Y=0 $X2=1.2
+ $Y2=0
r114 57 80 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r115 56 57 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r116 54 79 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.545 $Y=0 $X2=0.71
+ $Y2=0
r117 54 56 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.545 $Y=0
+ $X2=0.24 $Y2=0
r118 52 70 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.88 $Y=0
+ $X2=3.12 $Y2=0
r119 52 67 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=2.88 $Y=0 $X2=2.16
+ $Y2=0
r120 50 72 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=4.31 $Y=0 $X2=4.08
+ $Y2=0
r121 50 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.31 $Y=0 $X2=4.475
+ $Y2=0
r122 49 76 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=4.64 $Y=0 $X2=5.04
+ $Y2=0
r123 49 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.64 $Y=0 $X2=4.475
+ $Y2=0
r124 47 69 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=3.31 $Y=0 $X2=3.12
+ $Y2=0
r125 47 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.31 $Y=0 $X2=3.475
+ $Y2=0
r126 46 72 28.7059 $w=1.68e-07 $l=4.4e-07 $layer=LI1_cond $X=3.64 $Y=0 $X2=4.08
+ $Y2=0
r127 46 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.64 $Y=0 $X2=3.475
+ $Y2=0
r128 44 66 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=2.31 $Y=0 $X2=2.16
+ $Y2=0
r129 44 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.31 $Y=0 $X2=2.475
+ $Y2=0
r130 43 69 31.3155 $w=1.68e-07 $l=4.8e-07 $layer=LI1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r131 43 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.64 $Y=0 $X2=2.475
+ $Y2=0
r132 39 85 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=5.48 $Y=0.085
+ $X2=5.537 $Y2=0
r133 39 41 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=5.48 $Y=0.085
+ $X2=5.48 $Y2=0.515
r134 35 51 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.475 $Y=0.085
+ $X2=4.475 $Y2=0
r135 35 37 18.8582 $w=3.28e-07 $l=5.4e-07 $layer=LI1_cond $X=4.475 $Y=0.085
+ $X2=4.475 $Y2=0.625
r136 31 48 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.475 $Y=0.085
+ $X2=3.475 $Y2=0
r137 31 33 18.8582 $w=3.28e-07 $l=5.4e-07 $layer=LI1_cond $X=3.475 $Y=0.085
+ $X2=3.475 $Y2=0.625
r138 27 45 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.475 $Y=0.085
+ $X2=2.475 $Y2=0
r139 27 29 18.8582 $w=3.28e-07 $l=5.4e-07 $layer=LI1_cond $X=2.475 $Y=0.085
+ $X2=2.475 $Y2=0.625
r140 23 82 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.615 $Y=0.085
+ $X2=1.615 $Y2=0
r141 23 25 20.6043 $w=3.28e-07 $l=5.9e-07 $layer=LI1_cond $X=1.615 $Y=0.085
+ $X2=1.615 $Y2=0.675
r142 19 79 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.71 $Y=0.085
+ $X2=0.71 $Y2=0
r143 19 21 20.6043 $w=3.28e-07 $l=5.9e-07 $layer=LI1_cond $X=0.71 $Y=0.085
+ $X2=0.71 $Y2=0.675
r144 6 41 91 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=2 $X=5.27
+ $Y=0.37 $X2=5.48 $Y2=0.515
r145 5 37 182 $w=1.7e-07 $l=3.44347e-07 $layer=licon1_NDIFF $count=1 $X=4.265
+ $Y=0.37 $X2=4.475 $Y2=0.625
r146 4 33 182 $w=1.7e-07 $l=3.44347e-07 $layer=licon1_NDIFF $count=1 $X=3.265
+ $Y=0.37 $X2=3.475 $Y2=0.625
r147 3 29 182 $w=1.7e-07 $l=3.17372e-07 $layer=licon1_NDIFF $count=1 $X=2.335
+ $Y=0.37 $X2=2.475 $Y2=0.625
r148 2 25 182 $w=1.7e-07 $l=3.68409e-07 $layer=licon1_NDIFF $count=1 $X=1.475
+ $Y=0.37 $X2=1.615 $Y2=0.675
r149 1 21 182 $w=1.7e-07 $l=3.68409e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.37 $X2=0.71 $Y2=0.675
.ends

