* File: sky130_fd_sc_hs__dlxtn_1.pxi.spice
* Created: Tue Sep  1 20:02:57 2020
* 
x_PM_SKY130_FD_SC_HS__DLXTN_1%D N_D_c_127_n N_D_M1005_g N_D_c_128_n N_D_c_132_n
+ N_D_M1001_g D N_D_c_130_n PM_SKY130_FD_SC_HS__DLXTN_1%D
x_PM_SKY130_FD_SC_HS__DLXTN_1%GATE_N N_GATE_N_c_155_n N_GATE_N_M1000_g
+ N_GATE_N_M1008_g GATE_N PM_SKY130_FD_SC_HS__DLXTN_1%GATE_N
x_PM_SKY130_FD_SC_HS__DLXTN_1%A_217_419# N_A_217_419#_M1008_d
+ N_A_217_419#_M1000_d N_A_217_419#_c_206_n N_A_217_419#_M1003_g
+ N_A_217_419#_c_194_n N_A_217_419#_M1004_g N_A_217_419#_c_195_n
+ N_A_217_419#_M1017_g N_A_217_419#_c_196_n N_A_217_419#_c_207_n
+ N_A_217_419#_c_208_n N_A_217_419#_M1010_g N_A_217_419#_c_197_n
+ N_A_217_419#_c_198_n N_A_217_419#_c_199_n N_A_217_419#_c_200_n
+ N_A_217_419#_c_209_n N_A_217_419#_c_237_p N_A_217_419#_c_210_n
+ N_A_217_419#_c_211_n N_A_217_419#_c_212_n N_A_217_419#_c_213_n
+ N_A_217_419#_c_214_n N_A_217_419#_c_201_n N_A_217_419#_c_202_n
+ N_A_217_419#_c_203_n N_A_217_419#_c_204_n N_A_217_419#_c_205_n
+ PM_SKY130_FD_SC_HS__DLXTN_1%A_217_419#
x_PM_SKY130_FD_SC_HS__DLXTN_1%A_27_115# N_A_27_115#_M1005_s N_A_27_115#_M1001_s
+ N_A_27_115#_c_350_n N_A_27_115#_c_351_n N_A_27_115#_c_362_n
+ N_A_27_115#_M1009_g N_A_27_115#_c_352_n N_A_27_115#_c_353_n
+ N_A_27_115#_M1016_g N_A_27_115#_c_363_n N_A_27_115#_c_354_n
+ N_A_27_115#_c_382_n N_A_27_115#_c_355_n N_A_27_115#_c_356_n
+ N_A_27_115#_c_357_n N_A_27_115#_c_358_n N_A_27_115#_c_359_n
+ N_A_27_115#_c_365_n N_A_27_115#_c_360_n PM_SKY130_FD_SC_HS__DLXTN_1%A_27_115#
x_PM_SKY130_FD_SC_HS__DLXTN_1%A_369_392# N_A_369_392#_M1004_s
+ N_A_369_392#_M1003_s N_A_369_392#_c_469_n N_A_369_392#_M1013_g
+ N_A_369_392#_M1007_g N_A_369_392#_c_470_n N_A_369_392#_c_479_n
+ N_A_369_392#_c_471_n N_A_369_392#_c_472_n N_A_369_392#_c_473_n
+ N_A_369_392#_c_480_n N_A_369_392#_c_474_n N_A_369_392#_c_475_n
+ N_A_369_392#_c_476_n PM_SKY130_FD_SC_HS__DLXTN_1%A_369_392#
x_PM_SKY130_FD_SC_HS__DLXTN_1%A_863_441# N_A_863_441#_M1014_d
+ N_A_863_441#_M1011_d N_A_863_441#_c_574_n N_A_863_441#_M1015_g
+ N_A_863_441#_M1012_g N_A_863_441#_c_576_n N_A_863_441#_M1006_g
+ N_A_863_441#_M1002_g N_A_863_441#_c_567_n N_A_863_441#_c_568_n
+ N_A_863_441#_c_578_n N_A_863_441#_c_579_n N_A_863_441#_c_569_n
+ N_A_863_441#_c_570_n N_A_863_441#_c_581_n N_A_863_441#_c_571_n
+ N_A_863_441#_c_572_n N_A_863_441#_c_573_n
+ PM_SKY130_FD_SC_HS__DLXTN_1%A_863_441#
x_PM_SKY130_FD_SC_HS__DLXTN_1%A_669_392# N_A_669_392#_M1017_d
+ N_A_669_392#_M1013_d N_A_669_392#_c_658_n N_A_669_392#_c_667_n
+ N_A_669_392#_M1011_g N_A_669_392#_M1014_g N_A_669_392#_c_660_n
+ N_A_669_392#_c_674_n N_A_669_392#_c_661_n N_A_669_392#_c_662_n
+ N_A_669_392#_c_663_n N_A_669_392#_c_664_n N_A_669_392#_c_668_n
+ N_A_669_392#_c_665_n PM_SKY130_FD_SC_HS__DLXTN_1%A_669_392#
x_PM_SKY130_FD_SC_HS__DLXTN_1%VPWR N_VPWR_M1001_d N_VPWR_M1003_d N_VPWR_M1015_d
+ N_VPWR_M1006_s N_VPWR_c_750_n N_VPWR_c_751_n N_VPWR_c_752_n N_VPWR_c_753_n
+ N_VPWR_c_754_n N_VPWR_c_755_n VPWR N_VPWR_c_756_n N_VPWR_c_757_n
+ N_VPWR_c_758_n N_VPWR_c_759_n N_VPWR_c_749_n N_VPWR_c_761_n N_VPWR_c_762_n
+ N_VPWR_c_763_n PM_SKY130_FD_SC_HS__DLXTN_1%VPWR
x_PM_SKY130_FD_SC_HS__DLXTN_1%Q N_Q_M1002_d N_Q_M1006_d Q Q Q Q Q Q Q
+ PM_SKY130_FD_SC_HS__DLXTN_1%Q
x_PM_SKY130_FD_SC_HS__DLXTN_1%VGND N_VGND_M1005_d N_VGND_M1004_d N_VGND_M1012_d
+ N_VGND_M1002_s N_VGND_c_843_n N_VGND_c_844_n N_VGND_c_845_n N_VGND_c_846_n
+ N_VGND_c_847_n N_VGND_c_848_n VGND N_VGND_c_849_n N_VGND_c_850_n
+ N_VGND_c_851_n N_VGND_c_852_n N_VGND_c_853_n N_VGND_c_854_n N_VGND_c_855_n
+ N_VGND_c_856_n PM_SKY130_FD_SC_HS__DLXTN_1%VGND
cc_1 VNB N_D_c_127_n 0.023907f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.235
cc_2 VNB N_D_c_128_n 0.00821356f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=1.93
cc_3 VNB D 0.00853519f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_4 VNB N_D_c_130_n 0.0608998f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.4
cc_5 VNB N_GATE_N_c_155_n 0.017563f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.235
cc_6 VNB N_GATE_N_M1008_g 0.0250566f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=2.02
cc_7 VNB GATE_N 0.00137191f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=2.515
cc_8 VNB N_A_217_419#_c_194_n 0.0183659f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A_217_419#_c_195_n 0.0142192f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.4
cc_10 VNB N_A_217_419#_c_196_n 0.01469f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_217_419#_c_197_n 0.0280101f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_217_419#_c_198_n 0.00799851f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_217_419#_c_199_n 0.00995015f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_217_419#_c_200_n 0.00246966f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_217_419#_c_201_n 0.0390372f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_217_419#_c_202_n 5.58375e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_217_419#_c_203_n 0.00370923f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_217_419#_c_204_n 0.0304702f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_217_419#_c_205_n 0.0696329f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_27_115#_c_350_n 0.044003f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=2.515
cc_21 VNB N_A_27_115#_c_351_n 0.00641988f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=2.515
cc_22 VNB N_A_27_115#_c_352_n 0.0183536f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.4
cc_23 VNB N_A_27_115#_c_353_n 0.0159209f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.4
cc_24 VNB N_A_27_115#_c_354_n 0.00843476f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_27_115#_c_355_n 0.0222777f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_27_115#_c_356_n 0.00508052f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_27_115#_c_357_n 0.0239123f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_27_115#_c_358_n 0.00292455f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_27_115#_c_359_n 0.00226844f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_27_115#_c_360_n 0.00713993f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_369_392#_c_469_n 0.0210812f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=2.515
cc_32 VNB N_A_369_392#_c_470_n 4.52811e-19 $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=1.4
cc_33 VNB N_A_369_392#_c_471_n 0.00214971f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_369_392#_c_472_n 0.00976848f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_369_392#_c_473_n 0.0388293f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_369_392#_c_474_n 0.00311606f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_369_392#_c_475_n 0.00784989f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_369_392#_c_476_n 0.0167827f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_863_441#_M1012_g 0.038971f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.4
cc_40 VNB N_A_863_441#_M1002_g 0.0292088f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.4
cc_41 VNB N_A_863_441#_c_567_n 0.0564819f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_863_441#_c_568_n 0.0191627f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_863_441#_c_569_n 0.0084573f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_863_441#_c_570_n 5.75951e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_A_863_441#_c_571_n 0.00882152f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_A_863_441#_c_572_n 0.0162964f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_863_441#_c_573_n 0.00301142f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_669_392#_c_658_n 0.00155105f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=2.515
cc_49 VNB N_A_669_392#_M1014_g 0.0256539f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.4
cc_50 VNB N_A_669_392#_c_660_n 0.00129139f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_A_669_392#_c_661_n 0.00184728f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_A_669_392#_c_662_n 0.00365233f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_A_669_392#_c_663_n 0.0103795f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_A_669_392#_c_664_n 0.0293462f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_A_669_392#_c_665_n 0.00398491f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_VPWR_c_749_n 0.283096f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB Q 0.054669f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=2.515
cc_58 VNB N_VGND_c_843_n 0.0163672f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=1.4
cc_59 VNB N_VGND_c_844_n 0.00970291f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.4
cc_60 VNB N_VGND_c_845_n 0.0197811f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_VGND_c_846_n 0.0213431f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_VGND_c_847_n 0.0442207f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_VGND_c_848_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_VGND_c_849_n 0.0195521f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_VGND_c_850_n 0.0440818f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_VGND_c_851_n 0.0211139f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_VGND_c_852_n 0.0195898f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_VGND_c_853_n 0.39755f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_VGND_c_854_n 0.00631593f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_VGND_c_855_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_VGND_c_856_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VPB N_D_c_128_n 0.0188286f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=1.93
cc_73 VPB N_D_c_132_n 0.0267653f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=2.02
cc_74 VPB N_GATE_N_c_155_n 0.0509986f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.235
cc_75 VPB GATE_N 0.00166466f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=2.515
cc_76 VPB N_A_217_419#_c_206_n 0.0184208f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=2.515
cc_77 VPB N_A_217_419#_c_207_n 0.0360483f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.4
cc_78 VPB N_A_217_419#_c_208_n 0.0219267f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_79 VPB N_A_217_419#_c_209_n 0.00645301f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_80 VPB N_A_217_419#_c_210_n 0.00765968f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_81 VPB N_A_217_419#_c_211_n 8.72539e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_82 VPB N_A_217_419#_c_212_n 0.00650481f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_83 VPB N_A_217_419#_c_213_n 0.0294051f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_84 VPB N_A_217_419#_c_214_n 0.00652782f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_85 VPB N_A_217_419#_c_202_n 0.0038176f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_86 VPB N_A_217_419#_c_203_n 0.00534526f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_87 VPB N_A_217_419#_c_204_n 0.0252147f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_88 VPB N_A_217_419#_c_205_n 0.0374181f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_89 VPB N_A_27_115#_c_351_n 0.0074381f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=2.515
cc_90 VPB N_A_27_115#_c_362_n 0.0214413f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.21
cc_91 VPB N_A_27_115#_c_363_n 0.0440992f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.4
cc_92 VPB N_A_27_115#_c_354_n 0.00160101f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_93 VPB N_A_27_115#_c_365_n 0.0143789f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_94 VPB N_A_369_392#_c_469_n 0.0351174f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=2.515
cc_95 VPB N_A_369_392#_c_470_n 2.66113e-19 $X=-0.19 $Y=1.66 $X2=0.51 $Y2=1.4
cc_96 VPB N_A_369_392#_c_479_n 0.0219988f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_97 VPB N_A_369_392#_c_480_n 0.00855098f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_98 VPB N_A_369_392#_c_474_n 0.00265032f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_99 VPB N_A_863_441#_c_574_n 0.0702192f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=2.515
cc_100 VPB N_A_863_441#_M1012_g 0.0226503f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.4
cc_101 VPB N_A_863_441#_c_576_n 0.0208633f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.4
cc_102 VPB N_A_863_441#_c_568_n 0.00918987f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_103 VPB N_A_863_441#_c_578_n 0.00200721f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_104 VPB N_A_863_441#_c_579_n 0.00961903f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_105 VPB N_A_863_441#_c_570_n 0.00573494f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_106 VPB N_A_863_441#_c_581_n 0.0115165f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_107 VPB N_A_669_392#_c_658_n 0.00866003f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=2.515
cc_108 VPB N_A_669_392#_c_667_n 0.0260701f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.21
cc_109 VPB N_A_669_392#_c_668_n 0.00299652f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_110 VPB N_A_669_392#_c_665_n 0.00380426f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_111 VPB N_VPWR_c_750_n 0.0159115f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=1.4
cc_112 VPB N_VPWR_c_751_n 0.014119f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.4
cc_113 VPB N_VPWR_c_752_n 0.012039f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_114 VPB N_VPWR_c_753_n 0.0214784f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_115 VPB N_VPWR_c_754_n 0.0210901f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_116 VPB N_VPWR_c_755_n 0.0047828f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_117 VPB N_VPWR_c_756_n 0.0194332f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_118 VPB N_VPWR_c_757_n 0.0384481f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_119 VPB N_VPWR_c_758_n 0.0426279f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_120 VPB N_VPWR_c_759_n 0.0200671f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_121 VPB N_VPWR_c_749_n 0.102585f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_122 VPB N_VPWR_c_761_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_123 VPB N_VPWR_c_762_n 0.00660399f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_124 VPB N_VPWR_c_763_n 0.0112431f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_125 VPB Q 0.0536572f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=2.515
cc_126 N_D_c_132_n N_GATE_N_c_155_n 0.0195844f $X=0.51 $Y=2.02 $X2=-0.19
+ $Y2=-0.245
cc_127 N_D_c_130_n N_GATE_N_c_155_n 0.0182426f $X=0.495 $Y=1.4 $X2=-0.19
+ $Y2=-0.245
cc_128 N_D_c_127_n N_GATE_N_M1008_g 0.0208145f $X=0.495 $Y=1.235 $X2=0 $Y2=0
cc_129 N_D_c_130_n N_GATE_N_M1008_g 0.00189512f $X=0.495 $Y=1.4 $X2=0 $Y2=0
cc_130 N_D_c_128_n N_A_27_115#_c_363_n 0.00105226f $X=0.51 $Y=1.93 $X2=0 $Y2=0
cc_131 N_D_c_132_n N_A_27_115#_c_363_n 0.018666f $X=0.51 $Y=2.02 $X2=0 $Y2=0
cc_132 N_D_c_127_n N_A_27_115#_c_354_n 0.0047087f $X=0.495 $Y=1.235 $X2=0 $Y2=0
cc_133 D N_A_27_115#_c_354_n 0.0288934f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_134 N_D_c_130_n N_A_27_115#_c_354_n 0.00608894f $X=0.495 $Y=1.4 $X2=0 $Y2=0
cc_135 N_D_c_127_n N_A_27_115#_c_355_n 0.0228518f $X=0.495 $Y=1.235 $X2=0 $Y2=0
cc_136 D N_A_27_115#_c_355_n 0.0247838f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_137 N_D_c_130_n N_A_27_115#_c_355_n 0.00186348f $X=0.495 $Y=1.4 $X2=0 $Y2=0
cc_138 N_D_c_127_n N_A_27_115#_c_356_n 7.68306e-19 $X=0.495 $Y=1.235 $X2=0 $Y2=0
cc_139 N_D_c_128_n N_A_27_115#_c_365_n 0.0218158f $X=0.51 $Y=1.93 $X2=0 $Y2=0
cc_140 D N_A_27_115#_c_365_n 0.0239444f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_141 N_D_c_130_n N_A_27_115#_c_365_n 0.00211484f $X=0.495 $Y=1.4 $X2=0 $Y2=0
cc_142 N_D_c_132_n N_VPWR_c_750_n 0.00797131f $X=0.51 $Y=2.02 $X2=0 $Y2=0
cc_143 N_D_c_132_n N_VPWR_c_756_n 0.00544739f $X=0.51 $Y=2.02 $X2=0 $Y2=0
cc_144 N_D_c_132_n N_VPWR_c_749_n 0.00537853f $X=0.51 $Y=2.02 $X2=0 $Y2=0
cc_145 N_D_c_127_n N_VGND_c_843_n 0.00130869f $X=0.495 $Y=1.235 $X2=0 $Y2=0
cc_146 N_D_c_127_n N_VGND_c_849_n 0.00341528f $X=0.495 $Y=1.235 $X2=0 $Y2=0
cc_147 N_D_c_127_n N_VGND_c_853_n 0.0048347f $X=0.495 $Y=1.235 $X2=0 $Y2=0
cc_148 N_GATE_N_c_155_n N_A_217_419#_c_198_n 0.00261996f $X=1.01 $Y=2.02 $X2=0
+ $Y2=0
cc_149 N_GATE_N_M1008_g N_A_217_419#_c_198_n 0.00581294f $X=1.085 $Y=0.94 $X2=0
+ $Y2=0
cc_150 GATE_N N_A_217_419#_c_198_n 0.014308f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_151 N_GATE_N_M1008_g N_A_217_419#_c_199_n 0.00371584f $X=1.085 $Y=0.94 $X2=0
+ $Y2=0
cc_152 N_GATE_N_c_155_n N_A_217_419#_c_200_n 0.0012472f $X=1.01 $Y=2.02 $X2=0
+ $Y2=0
cc_153 N_GATE_N_M1008_g N_A_217_419#_c_200_n 0.00359662f $X=1.085 $Y=0.94 $X2=0
+ $Y2=0
cc_154 GATE_N N_A_217_419#_c_200_n 0.0276849f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_155 N_GATE_N_c_155_n N_A_217_419#_c_213_n 0.0228562f $X=1.01 $Y=2.02 $X2=0
+ $Y2=0
cc_156 GATE_N N_A_217_419#_c_213_n 0.0103789f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_157 N_GATE_N_c_155_n N_A_217_419#_c_214_n 0.00673688f $X=1.01 $Y=2.02 $X2=0
+ $Y2=0
cc_158 N_GATE_N_M1008_g N_A_217_419#_c_201_n 0.0155068f $X=1.085 $Y=0.94 $X2=0
+ $Y2=0
cc_159 N_GATE_N_c_155_n N_A_217_419#_c_205_n 0.0122983f $X=1.01 $Y=2.02 $X2=0
+ $Y2=0
cc_160 GATE_N N_A_217_419#_c_205_n 8.12953e-19 $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_161 N_GATE_N_c_155_n N_A_27_115#_c_363_n 0.00107913f $X=1.01 $Y=2.02 $X2=0
+ $Y2=0
cc_162 N_GATE_N_c_155_n N_A_27_115#_c_354_n 0.00168379f $X=1.01 $Y=2.02 $X2=0
+ $Y2=0
cc_163 N_GATE_N_M1008_g N_A_27_115#_c_354_n 0.00608847f $X=1.085 $Y=0.94 $X2=0
+ $Y2=0
cc_164 GATE_N N_A_27_115#_c_354_n 0.0178278f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_165 N_GATE_N_c_155_n N_A_27_115#_c_382_n 0.00156749f $X=1.01 $Y=2.02 $X2=0
+ $Y2=0
cc_166 N_GATE_N_M1008_g N_A_27_115#_c_382_n 0.0140794f $X=1.085 $Y=0.94 $X2=0
+ $Y2=0
cc_167 GATE_N N_A_27_115#_c_382_n 0.00371492f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_168 N_GATE_N_M1008_g N_A_27_115#_c_355_n 0.00509262f $X=1.085 $Y=0.94 $X2=0
+ $Y2=0
cc_169 N_GATE_N_M1008_g N_A_27_115#_c_356_n 0.00773574f $X=1.085 $Y=0.94 $X2=0
+ $Y2=0
cc_170 N_GATE_N_c_155_n N_A_27_115#_c_365_n 0.00287212f $X=1.01 $Y=2.02 $X2=0
+ $Y2=0
cc_171 GATE_N N_A_27_115#_c_365_n 0.00791845f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_172 N_GATE_N_c_155_n N_VPWR_c_750_n 0.0197973f $X=1.01 $Y=2.02 $X2=0 $Y2=0
cc_173 N_GATE_N_c_155_n N_VPWR_c_757_n 0.00502391f $X=1.01 $Y=2.02 $X2=0 $Y2=0
cc_174 N_GATE_N_c_155_n N_VPWR_c_749_n 0.00487653f $X=1.01 $Y=2.02 $X2=0 $Y2=0
cc_175 N_GATE_N_M1008_g N_VGND_c_843_n 5.5317e-19 $X=1.085 $Y=0.94 $X2=0 $Y2=0
cc_176 N_GATE_N_M1008_g N_VGND_c_850_n 0.00318127f $X=1.085 $Y=0.94 $X2=0 $Y2=0
cc_177 N_GATE_N_M1008_g N_VGND_c_853_n 0.00438121f $X=1.085 $Y=0.94 $X2=0 $Y2=0
cc_178 N_A_217_419#_c_194_n N_A_27_115#_c_350_n 0.0028424f $X=2.355 $Y=1.185
+ $X2=0 $Y2=0
cc_179 N_A_217_419#_c_205_n N_A_27_115#_c_350_n 0.0150713f $X=2.215 $Y=1.535
+ $X2=0 $Y2=0
cc_180 N_A_217_419#_c_205_n N_A_27_115#_c_351_n 0.00879135f $X=2.215 $Y=1.535
+ $X2=0 $Y2=0
cc_181 N_A_217_419#_c_206_n N_A_27_115#_c_362_n 0.025151f $X=2.215 $Y=1.885
+ $X2=0 $Y2=0
cc_182 N_A_217_419#_c_209_n N_A_27_115#_c_362_n 0.0126958f $X=2.875 $Y=2.525
+ $X2=0 $Y2=0
cc_183 N_A_217_419#_c_237_p N_A_27_115#_c_362_n 0.00707689f $X=2.96 $Y=2.905
+ $X2=0 $Y2=0
cc_184 N_A_217_419#_c_211_n N_A_27_115#_c_362_n 0.00428477f $X=3.045 $Y=2.99
+ $X2=0 $Y2=0
cc_185 N_A_217_419#_c_197_n N_A_27_115#_c_352_n 0.0229755f $X=3.805 $Y=1.185
+ $X2=0 $Y2=0
cc_186 N_A_217_419#_c_194_n N_A_27_115#_c_353_n 0.00461218f $X=2.355 $Y=1.185
+ $X2=0 $Y2=0
cc_187 N_A_217_419#_c_195_n N_A_27_115#_c_353_n 0.0229755f $X=3.59 $Y=1.11 $X2=0
+ $Y2=0
cc_188 N_A_217_419#_c_198_n N_A_27_115#_c_354_n 0.0140297f $X=1.485 $Y=1.165
+ $X2=0 $Y2=0
cc_189 N_A_217_419#_M1008_d N_A_27_115#_c_382_n 0.00616067f $X=1.16 $Y=0.57
+ $X2=0 $Y2=0
cc_190 N_A_217_419#_c_198_n N_A_27_115#_c_382_n 0.00997713f $X=1.485 $Y=1.165
+ $X2=0 $Y2=0
cc_191 N_A_217_419#_c_199_n N_A_27_115#_c_382_n 0.00618319f $X=1.685 $Y=1.33
+ $X2=0 $Y2=0
cc_192 N_A_217_419#_c_201_n N_A_27_115#_c_382_n 2.54774e-19 $X=1.72 $Y=0.925
+ $X2=0 $Y2=0
cc_193 N_A_217_419#_c_198_n N_A_27_115#_c_355_n 4.39007e-19 $X=1.485 $Y=1.165
+ $X2=0 $Y2=0
cc_194 N_A_217_419#_M1008_d N_A_27_115#_c_356_n 0.00339584f $X=1.16 $Y=0.57
+ $X2=0 $Y2=0
cc_195 N_A_217_419#_c_194_n N_A_27_115#_c_357_n 0.0156819f $X=2.355 $Y=1.185
+ $X2=0 $Y2=0
cc_196 N_A_217_419#_c_198_n N_A_27_115#_c_357_n 0.00552911f $X=1.485 $Y=1.165
+ $X2=0 $Y2=0
cc_197 N_A_217_419#_c_199_n N_A_27_115#_c_357_n 0.0169889f $X=1.685 $Y=1.33
+ $X2=0 $Y2=0
cc_198 N_A_217_419#_c_201_n N_A_27_115#_c_357_n 0.00199179f $X=1.72 $Y=0.925
+ $X2=0 $Y2=0
cc_199 N_A_217_419#_c_194_n N_A_27_115#_c_359_n 0.00722178f $X=2.355 $Y=1.185
+ $X2=0 $Y2=0
cc_200 N_A_217_419#_c_205_n N_A_27_115#_c_360_n 0.00275434f $X=2.215 $Y=1.535
+ $X2=0 $Y2=0
cc_201 N_A_217_419#_c_209_n N_A_369_392#_M1003_s 0.00811065f $X=2.875 $Y=2.525
+ $X2=0 $Y2=0
cc_202 N_A_217_419#_c_207_n N_A_369_392#_c_469_n 0.00978818f $X=3.985 $Y=2.375
+ $X2=0 $Y2=0
cc_203 N_A_217_419#_c_208_n N_A_369_392#_c_469_n 0.0103911f $X=3.985 $Y=2.465
+ $X2=0 $Y2=0
cc_204 N_A_217_419#_c_209_n N_A_369_392#_c_469_n 0.00143509f $X=2.875 $Y=2.525
+ $X2=0 $Y2=0
cc_205 N_A_217_419#_c_237_p N_A_369_392#_c_469_n 0.00443826f $X=2.96 $Y=2.905
+ $X2=0 $Y2=0
cc_206 N_A_217_419#_c_210_n N_A_369_392#_c_469_n 0.0143782f $X=4.01 $Y=2.99
+ $X2=0 $Y2=0
cc_207 N_A_217_419#_c_212_n N_A_369_392#_c_469_n 0.00115231f $X=4.095 $Y=2.905
+ $X2=0 $Y2=0
cc_208 N_A_217_419#_c_204_n N_A_369_392#_c_469_n 0.0185905f $X=4.175 $Y=1.62
+ $X2=0 $Y2=0
cc_209 N_A_217_419#_c_194_n N_A_369_392#_c_470_n 0.0094035f $X=2.355 $Y=1.185
+ $X2=0 $Y2=0
cc_210 N_A_217_419#_c_199_n N_A_369_392#_c_470_n 0.044954f $X=1.685 $Y=1.33
+ $X2=0 $Y2=0
cc_211 N_A_217_419#_c_200_n N_A_369_392#_c_470_n 0.0295284f $X=1.685 $Y=1.57
+ $X2=0 $Y2=0
cc_212 N_A_217_419#_c_201_n N_A_369_392#_c_470_n 0.00156461f $X=1.72 $Y=0.925
+ $X2=0 $Y2=0
cc_213 N_A_217_419#_c_205_n N_A_369_392#_c_470_n 0.0291082f $X=2.215 $Y=1.535
+ $X2=0 $Y2=0
cc_214 N_A_217_419#_c_209_n N_A_369_392#_c_479_n 0.0207776f $X=2.875 $Y=2.525
+ $X2=0 $Y2=0
cc_215 N_A_217_419#_c_205_n N_A_369_392#_c_479_n 0.00409565f $X=2.215 $Y=1.535
+ $X2=0 $Y2=0
cc_216 N_A_217_419#_c_195_n N_A_369_392#_c_472_n 0.0201753f $X=3.59 $Y=1.11
+ $X2=0 $Y2=0
cc_217 N_A_217_419#_c_197_n N_A_369_392#_c_472_n 6.48245e-19 $X=3.805 $Y=1.185
+ $X2=0 $Y2=0
cc_218 N_A_217_419#_c_195_n N_A_369_392#_c_473_n 0.0103701f $X=3.59 $Y=1.11
+ $X2=0 $Y2=0
cc_219 N_A_217_419#_c_206_n N_A_369_392#_c_480_n 0.0142993f $X=2.215 $Y=1.885
+ $X2=0 $Y2=0
cc_220 N_A_217_419#_c_209_n N_A_369_392#_c_480_n 0.02864f $X=2.875 $Y=2.525
+ $X2=0 $Y2=0
cc_221 N_A_217_419#_c_214_n N_A_369_392#_c_480_n 0.0356523f $X=1.405 $Y=2.075
+ $X2=0 $Y2=0
cc_222 N_A_217_419#_c_202_n N_A_369_392#_c_480_n 0.0088212f $X=1.72 $Y=1.605
+ $X2=0 $Y2=0
cc_223 N_A_217_419#_c_205_n N_A_369_392#_c_480_n 0.0153271f $X=2.215 $Y=1.535
+ $X2=0 $Y2=0
cc_224 N_A_217_419#_c_204_n N_A_369_392#_c_474_n 3.42585e-19 $X=4.175 $Y=1.62
+ $X2=0 $Y2=0
cc_225 N_A_217_419#_c_195_n N_A_369_392#_c_475_n 0.00344145f $X=3.59 $Y=1.11
+ $X2=0 $Y2=0
cc_226 N_A_217_419#_c_196_n N_A_369_392#_c_475_n 0.00125106f $X=3.805 $Y=1.455
+ $X2=0 $Y2=0
cc_227 N_A_217_419#_c_195_n N_A_369_392#_c_476_n 0.0110573f $X=3.59 $Y=1.11
+ $X2=0 $Y2=0
cc_228 N_A_217_419#_c_197_n N_A_369_392#_c_476_n 0.00502885f $X=3.805 $Y=1.185
+ $X2=0 $Y2=0
cc_229 N_A_217_419#_c_203_n N_A_369_392#_c_476_n 6.07693e-19 $X=4.175 $Y=1.62
+ $X2=0 $Y2=0
cc_230 N_A_217_419#_c_204_n N_A_369_392#_c_476_n 0.00901901f $X=4.175 $Y=1.62
+ $X2=0 $Y2=0
cc_231 N_A_217_419#_c_207_n N_A_863_441#_c_574_n 0.0216769f $X=3.985 $Y=2.375
+ $X2=0 $Y2=0
cc_232 N_A_217_419#_c_208_n N_A_863_441#_c_574_n 0.0265789f $X=3.985 $Y=2.465
+ $X2=0 $Y2=0
cc_233 N_A_217_419#_c_210_n N_A_863_441#_c_574_n 0.00144847f $X=4.01 $Y=2.99
+ $X2=0 $Y2=0
cc_234 N_A_217_419#_c_212_n N_A_863_441#_c_574_n 0.00838792f $X=4.095 $Y=2.905
+ $X2=0 $Y2=0
cc_235 N_A_217_419#_c_204_n N_A_863_441#_c_574_n 6.7394e-19 $X=4.175 $Y=1.62
+ $X2=0 $Y2=0
cc_236 N_A_217_419#_c_207_n N_A_863_441#_M1012_g 0.00414193f $X=3.985 $Y=2.375
+ $X2=0 $Y2=0
cc_237 N_A_217_419#_c_197_n N_A_863_441#_M1012_g 0.00219948f $X=3.805 $Y=1.185
+ $X2=0 $Y2=0
cc_238 N_A_217_419#_c_212_n N_A_863_441#_M1012_g 0.00407454f $X=4.095 $Y=2.905
+ $X2=0 $Y2=0
cc_239 N_A_217_419#_c_203_n N_A_863_441#_M1012_g 0.0011566f $X=4.175 $Y=1.62
+ $X2=0 $Y2=0
cc_240 N_A_217_419#_c_204_n N_A_863_441#_M1012_g 0.0174593f $X=4.175 $Y=1.62
+ $X2=0 $Y2=0
cc_241 N_A_217_419#_c_207_n N_A_863_441#_c_578_n 3.34543e-19 $X=3.985 $Y=2.375
+ $X2=0 $Y2=0
cc_242 N_A_217_419#_c_212_n N_A_863_441#_c_578_n 0.0262118f $X=4.095 $Y=2.905
+ $X2=0 $Y2=0
cc_243 N_A_217_419#_c_210_n N_A_669_392#_M1013_d 0.0057923f $X=4.01 $Y=2.99
+ $X2=0 $Y2=0
cc_244 N_A_217_419#_c_197_n N_A_669_392#_c_660_n 0.00191766f $X=3.805 $Y=1.185
+ $X2=0 $Y2=0
cc_245 N_A_217_419#_c_203_n N_A_669_392#_c_660_n 0.0118013f $X=4.175 $Y=1.62
+ $X2=0 $Y2=0
cc_246 N_A_217_419#_c_204_n N_A_669_392#_c_660_n 0.00550226f $X=4.175 $Y=1.62
+ $X2=0 $Y2=0
cc_247 N_A_217_419#_c_195_n N_A_669_392#_c_674_n 0.00743237f $X=3.59 $Y=1.11
+ $X2=0 $Y2=0
cc_248 N_A_217_419#_c_197_n N_A_669_392#_c_674_n 2.03611e-19 $X=3.805 $Y=1.185
+ $X2=0 $Y2=0
cc_249 N_A_217_419#_c_197_n N_A_669_392#_c_661_n 6.85352e-19 $X=3.805 $Y=1.185
+ $X2=0 $Y2=0
cc_250 N_A_217_419#_c_196_n N_A_669_392#_c_662_n 0.001192f $X=3.805 $Y=1.455
+ $X2=0 $Y2=0
cc_251 N_A_217_419#_c_203_n N_A_669_392#_c_662_n 0.01518f $X=4.175 $Y=1.62 $X2=0
+ $Y2=0
cc_252 N_A_217_419#_c_204_n N_A_669_392#_c_662_n 0.00131112f $X=4.175 $Y=1.62
+ $X2=0 $Y2=0
cc_253 N_A_217_419#_c_208_n N_A_669_392#_c_668_n 0.00660021f $X=3.985 $Y=2.465
+ $X2=0 $Y2=0
cc_254 N_A_217_419#_c_209_n N_A_669_392#_c_668_n 0.00972995f $X=2.875 $Y=2.525
+ $X2=0 $Y2=0
cc_255 N_A_217_419#_c_237_p N_A_669_392#_c_668_n 0.00639531f $X=2.96 $Y=2.905
+ $X2=0 $Y2=0
cc_256 N_A_217_419#_c_210_n N_A_669_392#_c_668_n 0.0342344f $X=4.01 $Y=2.99
+ $X2=0 $Y2=0
cc_257 N_A_217_419#_c_212_n N_A_669_392#_c_668_n 0.0478039f $X=4.095 $Y=2.905
+ $X2=0 $Y2=0
cc_258 N_A_217_419#_c_195_n N_A_669_392#_c_665_n 6.1471e-19 $X=3.59 $Y=1.11
+ $X2=0 $Y2=0
cc_259 N_A_217_419#_c_196_n N_A_669_392#_c_665_n 0.00839087f $X=3.805 $Y=1.455
+ $X2=0 $Y2=0
cc_260 N_A_217_419#_c_207_n N_A_669_392#_c_665_n 0.00369358f $X=3.985 $Y=2.375
+ $X2=0 $Y2=0
cc_261 N_A_217_419#_c_197_n N_A_669_392#_c_665_n 0.0108592f $X=3.805 $Y=1.185
+ $X2=0 $Y2=0
cc_262 N_A_217_419#_c_203_n N_A_669_392#_c_665_n 0.0478039f $X=4.175 $Y=1.62
+ $X2=0 $Y2=0
cc_263 N_A_217_419#_c_204_n N_A_669_392#_c_665_n 0.0119327f $X=4.175 $Y=1.62
+ $X2=0 $Y2=0
cc_264 N_A_217_419#_c_209_n N_VPWR_M1003_d 0.0122282f $X=2.875 $Y=2.525 $X2=0
+ $Y2=0
cc_265 N_A_217_419#_c_213_n N_VPWR_c_750_n 0.0611759f $X=1.32 $Y=2.24 $X2=0
+ $Y2=0
cc_266 N_A_217_419#_c_206_n N_VPWR_c_751_n 0.00438753f $X=2.215 $Y=1.885 $X2=0
+ $Y2=0
cc_267 N_A_217_419#_c_209_n N_VPWR_c_751_n 0.0267961f $X=2.875 $Y=2.525 $X2=0
+ $Y2=0
cc_268 N_A_217_419#_c_237_p N_VPWR_c_751_n 0.00924851f $X=2.96 $Y=2.905 $X2=0
+ $Y2=0
cc_269 N_A_217_419#_c_211_n N_VPWR_c_751_n 0.0142284f $X=3.045 $Y=2.99 $X2=0
+ $Y2=0
cc_270 N_A_217_419#_c_208_n N_VPWR_c_752_n 5.74056e-19 $X=3.985 $Y=2.465 $X2=0
+ $Y2=0
cc_271 N_A_217_419#_c_210_n N_VPWR_c_752_n 0.00992039f $X=4.01 $Y=2.99 $X2=0
+ $Y2=0
cc_272 N_A_217_419#_c_212_n N_VPWR_c_752_n 0.0194917f $X=4.095 $Y=2.905 $X2=0
+ $Y2=0
cc_273 N_A_217_419#_c_206_n N_VPWR_c_757_n 0.00366846f $X=2.215 $Y=1.885 $X2=0
+ $Y2=0
cc_274 N_A_217_419#_c_209_n N_VPWR_c_757_n 0.00949357f $X=2.875 $Y=2.525 $X2=0
+ $Y2=0
cc_275 N_A_217_419#_c_213_n N_VPWR_c_757_n 0.0201915f $X=1.32 $Y=2.24 $X2=0
+ $Y2=0
cc_276 N_A_217_419#_c_208_n N_VPWR_c_758_n 0.00278223f $X=3.985 $Y=2.465 $X2=0
+ $Y2=0
cc_277 N_A_217_419#_c_209_n N_VPWR_c_758_n 0.00197454f $X=2.875 $Y=2.525 $X2=0
+ $Y2=0
cc_278 N_A_217_419#_c_210_n N_VPWR_c_758_n 0.0733589f $X=4.01 $Y=2.99 $X2=0
+ $Y2=0
cc_279 N_A_217_419#_c_211_n N_VPWR_c_758_n 0.0119496f $X=3.045 $Y=2.99 $X2=0
+ $Y2=0
cc_280 N_A_217_419#_c_206_n N_VPWR_c_749_n 0.0049649f $X=2.215 $Y=1.885 $X2=0
+ $Y2=0
cc_281 N_A_217_419#_c_208_n N_VPWR_c_749_n 0.00355603f $X=3.985 $Y=2.465 $X2=0
+ $Y2=0
cc_282 N_A_217_419#_c_209_n N_VPWR_c_749_n 0.0241361f $X=2.875 $Y=2.525 $X2=0
+ $Y2=0
cc_283 N_A_217_419#_c_210_n N_VPWR_c_749_n 0.0415125f $X=4.01 $Y=2.99 $X2=0
+ $Y2=0
cc_284 N_A_217_419#_c_211_n N_VPWR_c_749_n 0.00636858f $X=3.045 $Y=2.99 $X2=0
+ $Y2=0
cc_285 N_A_217_419#_c_213_n N_VPWR_c_749_n 0.0181131f $X=1.32 $Y=2.24 $X2=0
+ $Y2=0
cc_286 N_A_217_419#_c_209_n A_585_392# 0.00306281f $X=2.875 $Y=2.525 $X2=-0.19
+ $Y2=-0.245
cc_287 N_A_217_419#_c_237_p A_585_392# 0.00320536f $X=2.96 $Y=2.905 $X2=-0.19
+ $Y2=-0.245
cc_288 N_A_217_419#_c_210_n A_585_392# 0.00351031f $X=4.01 $Y=2.99 $X2=-0.19
+ $Y2=-0.245
cc_289 N_A_217_419#_c_210_n A_812_508# 5.9219e-19 $X=4.01 $Y=2.99 $X2=-0.19
+ $Y2=-0.245
cc_290 N_A_217_419#_c_212_n A_812_508# 0.00375576f $X=4.095 $Y=2.905 $X2=-0.19
+ $Y2=-0.245
cc_291 N_A_217_419#_c_194_n N_VGND_c_844_n 0.00196203f $X=2.355 $Y=1.185 $X2=0
+ $Y2=0
cc_292 N_A_217_419#_c_195_n N_VGND_c_844_n 3.86051e-19 $X=3.59 $Y=1.11 $X2=0
+ $Y2=0
cc_293 N_A_217_419#_c_195_n N_VGND_c_847_n 9.44495e-19 $X=3.59 $Y=1.11 $X2=0
+ $Y2=0
cc_294 N_A_217_419#_c_194_n N_VGND_c_850_n 0.00278271f $X=2.355 $Y=1.185 $X2=0
+ $Y2=0
cc_295 N_A_217_419#_c_194_n N_VGND_c_853_n 0.00363426f $X=2.355 $Y=1.185 $X2=0
+ $Y2=0
cc_296 N_A_27_115#_c_357_n N_A_369_392#_M1004_s 0.00441657f $X=2.475 $Y=0.34
+ $X2=-0.19 $Y2=-0.245
cc_297 N_A_27_115#_c_350_n N_A_369_392#_c_469_n 0.00535816f $X=2.85 $Y=1.555
+ $X2=0 $Y2=0
cc_298 N_A_27_115#_c_351_n N_A_369_392#_c_469_n 0.0183178f $X=2.85 $Y=1.795
+ $X2=0 $Y2=0
cc_299 N_A_27_115#_c_362_n N_A_369_392#_c_469_n 0.0556309f $X=2.85 $Y=1.885
+ $X2=0 $Y2=0
cc_300 N_A_27_115#_c_352_n N_A_369_392#_c_469_n 0.00637363f $X=3.125 $Y=1.185
+ $X2=0 $Y2=0
cc_301 N_A_27_115#_c_360_n N_A_369_392#_c_469_n 2.92453e-19 $X=2.805 $Y=1.39
+ $X2=0 $Y2=0
cc_302 N_A_27_115#_c_350_n N_A_369_392#_c_470_n 2.97794e-19 $X=2.85 $Y=1.555
+ $X2=0 $Y2=0
cc_303 N_A_27_115#_c_351_n N_A_369_392#_c_470_n 9.58777e-19 $X=2.85 $Y=1.795
+ $X2=0 $Y2=0
cc_304 N_A_27_115#_c_357_n N_A_369_392#_c_470_n 0.0144209f $X=2.475 $Y=0.34
+ $X2=0 $Y2=0
cc_305 N_A_27_115#_c_359_n N_A_369_392#_c_470_n 0.0269076f $X=2.56 $Y=1.225
+ $X2=0 $Y2=0
cc_306 N_A_27_115#_c_360_n N_A_369_392#_c_470_n 0.0264318f $X=2.805 $Y=1.39
+ $X2=0 $Y2=0
cc_307 N_A_27_115#_c_350_n N_A_369_392#_c_479_n 0.00340591f $X=2.85 $Y=1.555
+ $X2=0 $Y2=0
cc_308 N_A_27_115#_c_351_n N_A_369_392#_c_479_n 0.00538946f $X=2.85 $Y=1.795
+ $X2=0 $Y2=0
cc_309 N_A_27_115#_c_362_n N_A_369_392#_c_479_n 0.00857984f $X=2.85 $Y=1.885
+ $X2=0 $Y2=0
cc_310 N_A_27_115#_c_352_n N_A_369_392#_c_479_n 0.00407107f $X=3.125 $Y=1.185
+ $X2=0 $Y2=0
cc_311 N_A_27_115#_c_360_n N_A_369_392#_c_479_n 0.0372099f $X=2.805 $Y=1.39
+ $X2=0 $Y2=0
cc_312 N_A_27_115#_c_353_n N_A_369_392#_c_471_n 0.00172839f $X=3.2 $Y=1.11 $X2=0
+ $Y2=0
cc_313 N_A_27_115#_c_362_n N_A_369_392#_c_480_n 0.00182085f $X=2.85 $Y=1.885
+ $X2=0 $Y2=0
cc_314 N_A_27_115#_c_351_n N_A_369_392#_c_474_n 0.00122716f $X=2.85 $Y=1.795
+ $X2=0 $Y2=0
cc_315 N_A_27_115#_c_352_n N_A_369_392#_c_474_n 7.22068e-19 $X=3.125 $Y=1.185
+ $X2=0 $Y2=0
cc_316 N_A_27_115#_c_360_n N_A_369_392#_c_474_n 0.00550381f $X=2.805 $Y=1.39
+ $X2=0 $Y2=0
cc_317 N_A_27_115#_c_350_n N_A_369_392#_c_475_n 0.00126828f $X=2.85 $Y=1.555
+ $X2=0 $Y2=0
cc_318 N_A_27_115#_c_353_n N_A_369_392#_c_475_n 0.0045287f $X=3.2 $Y=1.11 $X2=0
+ $Y2=0
cc_319 N_A_27_115#_c_359_n N_A_369_392#_c_475_n 0.00474577f $X=2.56 $Y=1.225
+ $X2=0 $Y2=0
cc_320 N_A_27_115#_c_360_n N_A_369_392#_c_475_n 0.0111511f $X=2.805 $Y=1.39
+ $X2=0 $Y2=0
cc_321 N_A_27_115#_c_362_n N_A_669_392#_c_668_n 0.00205487f $X=2.85 $Y=1.885
+ $X2=0 $Y2=0
cc_322 N_A_27_115#_c_363_n N_VPWR_c_750_n 0.0346007f $X=0.285 $Y=2.24 $X2=0
+ $Y2=0
cc_323 N_A_27_115#_c_365_n N_VPWR_c_750_n 0.0129691f $X=0.69 $Y=1.82 $X2=0 $Y2=0
cc_324 N_A_27_115#_c_362_n N_VPWR_c_751_n 0.00522314f $X=2.85 $Y=1.885 $X2=0
+ $Y2=0
cc_325 N_A_27_115#_c_363_n N_VPWR_c_756_n 0.0132586f $X=0.285 $Y=2.24 $X2=0
+ $Y2=0
cc_326 N_A_27_115#_c_362_n N_VPWR_c_758_n 0.0031609f $X=2.85 $Y=1.885 $X2=0
+ $Y2=0
cc_327 N_A_27_115#_c_362_n N_VPWR_c_749_n 0.0041189f $X=2.85 $Y=1.885 $X2=0
+ $Y2=0
cc_328 N_A_27_115#_c_363_n N_VPWR_c_749_n 0.0119178f $X=0.285 $Y=2.24 $X2=0
+ $Y2=0
cc_329 N_A_27_115#_c_354_n N_VGND_M1005_d 0.00379202f $X=0.69 $Y=1.735 $X2=-0.19
+ $Y2=-0.245
cc_330 N_A_27_115#_c_382_n N_VGND_M1005_d 0.00840371f $X=1.145 $Y=0.745
+ $X2=-0.19 $Y2=-0.245
cc_331 N_A_27_115#_c_355_n N_VGND_M1005_d 0.00462497f $X=0.775 $Y=0.745
+ $X2=-0.19 $Y2=-0.245
cc_332 N_A_27_115#_c_357_n N_VGND_M1004_d 6.45227e-19 $X=2.475 $Y=0.34 $X2=0
+ $Y2=0
cc_333 N_A_27_115#_c_359_n N_VGND_M1004_d 0.0110386f $X=2.56 $Y=1.225 $X2=0
+ $Y2=0
cc_334 N_A_27_115#_c_382_n N_VGND_c_843_n 0.0137179f $X=1.145 $Y=0.745 $X2=0
+ $Y2=0
cc_335 N_A_27_115#_c_355_n N_VGND_c_843_n 0.0126353f $X=0.775 $Y=0.745 $X2=0
+ $Y2=0
cc_336 N_A_27_115#_c_356_n N_VGND_c_843_n 0.0045384f $X=1.23 $Y=0.66 $X2=0 $Y2=0
cc_337 N_A_27_115#_c_358_n N_VGND_c_843_n 0.0139003f $X=1.315 $Y=0.34 $X2=0
+ $Y2=0
cc_338 N_A_27_115#_c_350_n N_VGND_c_844_n 0.00944812f $X=2.85 $Y=1.555 $X2=0
+ $Y2=0
cc_339 N_A_27_115#_c_353_n N_VGND_c_844_n 0.0109791f $X=3.2 $Y=1.11 $X2=0 $Y2=0
cc_340 N_A_27_115#_c_357_n N_VGND_c_844_n 0.0148948f $X=2.475 $Y=0.34 $X2=0
+ $Y2=0
cc_341 N_A_27_115#_c_359_n N_VGND_c_844_n 0.0481399f $X=2.56 $Y=1.225 $X2=0
+ $Y2=0
cc_342 N_A_27_115#_c_360_n N_VGND_c_844_n 0.0129855f $X=2.805 $Y=1.39 $X2=0
+ $Y2=0
cc_343 N_A_27_115#_c_353_n N_VGND_c_847_n 0.00483734f $X=3.2 $Y=1.11 $X2=0 $Y2=0
cc_344 N_A_27_115#_c_355_n N_VGND_c_849_n 0.0102001f $X=0.775 $Y=0.745 $X2=0
+ $Y2=0
cc_345 N_A_27_115#_c_382_n N_VGND_c_850_n 0.00257035f $X=1.145 $Y=0.745 $X2=0
+ $Y2=0
cc_346 N_A_27_115#_c_357_n N_VGND_c_850_n 0.086417f $X=2.475 $Y=0.34 $X2=0 $Y2=0
cc_347 N_A_27_115#_c_358_n N_VGND_c_850_n 0.0120335f $X=1.315 $Y=0.34 $X2=0
+ $Y2=0
cc_348 N_A_27_115#_c_353_n N_VGND_c_853_n 0.00469725f $X=3.2 $Y=1.11 $X2=0 $Y2=0
cc_349 N_A_27_115#_c_382_n N_VGND_c_853_n 0.00597829f $X=1.145 $Y=0.745 $X2=0
+ $Y2=0
cc_350 N_A_27_115#_c_355_n N_VGND_c_853_n 0.0162516f $X=0.775 $Y=0.745 $X2=0
+ $Y2=0
cc_351 N_A_27_115#_c_357_n N_VGND_c_853_n 0.049532f $X=2.475 $Y=0.34 $X2=0 $Y2=0
cc_352 N_A_27_115#_c_358_n N_VGND_c_853_n 0.00658039f $X=1.315 $Y=0.34 $X2=0
+ $Y2=0
cc_353 N_A_369_392#_c_473_n N_A_863_441#_M1012_g 0.0360676f $X=4.19 $Y=0.42
+ $X2=0 $Y2=0
cc_354 N_A_369_392#_c_472_n N_A_669_392#_M1017_d 0.00212267f $X=4.19 $Y=0.42
+ $X2=-0.19 $Y2=-0.245
cc_355 N_A_369_392#_c_472_n N_A_669_392#_c_660_n 0.0290049f $X=4.19 $Y=0.42
+ $X2=0 $Y2=0
cc_356 N_A_369_392#_c_473_n N_A_669_392#_c_660_n 0.00378883f $X=4.19 $Y=0.42
+ $X2=0 $Y2=0
cc_357 N_A_369_392#_c_476_n N_A_669_392#_c_660_n 0.0155131f $X=4.19 $Y=0.585
+ $X2=0 $Y2=0
cc_358 N_A_369_392#_c_472_n N_A_669_392#_c_674_n 0.00839569f $X=4.19 $Y=0.42
+ $X2=0 $Y2=0
cc_359 N_A_369_392#_c_475_n N_A_669_392#_c_674_n 0.0112489f $X=3.34 $Y=1.47
+ $X2=0 $Y2=0
cc_360 N_A_369_392#_c_476_n N_A_669_392#_c_661_n 0.00195157f $X=4.19 $Y=0.585
+ $X2=0 $Y2=0
cc_361 N_A_369_392#_c_469_n N_A_669_392#_c_668_n 0.0238743f $X=3.27 $Y=1.885
+ $X2=0 $Y2=0
cc_362 N_A_369_392#_c_474_n N_A_669_392#_c_668_n 0.0127169f $X=3.345 $Y=1.635
+ $X2=0 $Y2=0
cc_363 N_A_369_392#_c_469_n N_A_669_392#_c_665_n 0.00535501f $X=3.27 $Y=1.885
+ $X2=0 $Y2=0
cc_364 N_A_369_392#_c_474_n N_A_669_392#_c_665_n 0.0322562f $X=3.345 $Y=1.635
+ $X2=0 $Y2=0
cc_365 N_A_369_392#_c_475_n N_A_669_392#_c_665_n 0.0287917f $X=3.34 $Y=1.47
+ $X2=0 $Y2=0
cc_366 N_A_369_392#_c_476_n N_A_669_392#_c_665_n 0.00100266f $X=4.19 $Y=0.585
+ $X2=0 $Y2=0
cc_367 N_A_369_392#_c_469_n N_VPWR_c_758_n 0.00278271f $X=3.27 $Y=1.885 $X2=0
+ $Y2=0
cc_368 N_A_369_392#_c_469_n N_VPWR_c_749_n 0.00355607f $X=3.27 $Y=1.885 $X2=0
+ $Y2=0
cc_369 N_A_369_392#_c_479_n N_VGND_c_844_n 0.00546692f $X=3.18 $Y=1.81 $X2=0
+ $Y2=0
cc_370 N_A_369_392#_c_471_n N_VGND_c_844_n 0.0189627f $X=3.485 $Y=0.42 $X2=0
+ $Y2=0
cc_371 N_A_369_392#_c_475_n N_VGND_c_844_n 0.0183504f $X=3.34 $Y=1.47 $X2=0
+ $Y2=0
cc_372 N_A_369_392#_c_472_n N_VGND_c_845_n 0.0120179f $X=4.19 $Y=0.42 $X2=0
+ $Y2=0
cc_373 N_A_369_392#_c_473_n N_VGND_c_845_n 0.00178328f $X=4.19 $Y=0.42 $X2=0
+ $Y2=0
cc_374 N_A_369_392#_c_471_n N_VGND_c_847_n 0.0121867f $X=3.485 $Y=0.42 $X2=0
+ $Y2=0
cc_375 N_A_369_392#_c_472_n N_VGND_c_847_n 0.0576446f $X=4.19 $Y=0.42 $X2=0
+ $Y2=0
cc_376 N_A_369_392#_c_473_n N_VGND_c_847_n 0.00783549f $X=4.19 $Y=0.42 $X2=0
+ $Y2=0
cc_377 N_A_369_392#_c_471_n N_VGND_c_853_n 0.00660921f $X=3.485 $Y=0.42 $X2=0
+ $Y2=0
cc_378 N_A_369_392#_c_472_n N_VGND_c_853_n 0.0330012f $X=4.19 $Y=0.42 $X2=0
+ $Y2=0
cc_379 N_A_369_392#_c_473_n N_VGND_c_853_n 0.011167f $X=4.19 $Y=0.42 $X2=0 $Y2=0
cc_380 N_A_369_392#_c_475_n A_655_79# 0.00191955f $X=3.34 $Y=1.47 $X2=-0.19
+ $Y2=-0.245
cc_381 N_A_863_441#_M1012_g N_A_669_392#_c_658_n 0.00996804f $X=4.67 $Y=0.905
+ $X2=0 $Y2=0
cc_382 N_A_863_441#_c_570_n N_A_669_392#_c_658_n 0.00851758f $X=5.57 $Y=1.94
+ $X2=0 $Y2=0
cc_383 N_A_863_441#_c_574_n N_A_669_392#_c_667_n 0.00587655f $X=4.405 $Y=2.465
+ $X2=0 $Y2=0
cc_384 N_A_863_441#_M1012_g N_A_669_392#_c_667_n 0.0146004f $X=4.67 $Y=0.905
+ $X2=0 $Y2=0
cc_385 N_A_863_441#_c_578_n N_A_669_392#_c_667_n 0.0184063f $X=5.265 $Y=2.19
+ $X2=0 $Y2=0
cc_386 N_A_863_441#_c_579_n N_A_669_392#_c_667_n 0.0127548f $X=5.43 $Y=2.815
+ $X2=0 $Y2=0
cc_387 N_A_863_441#_c_581_n N_A_669_392#_c_667_n 0.00330776f $X=5.43 $Y=2.105
+ $X2=0 $Y2=0
cc_388 N_A_863_441#_M1012_g N_A_669_392#_M1014_g 0.0110566f $X=4.67 $Y=0.905
+ $X2=0 $Y2=0
cc_389 N_A_863_441#_c_567_n N_A_669_392#_M1014_g 2.16706e-19 $X=6.125 $Y=1.465
+ $X2=0 $Y2=0
cc_390 N_A_863_441#_c_569_n N_A_669_392#_M1014_g 0.00592153f $X=5.445 $Y=0.62
+ $X2=0 $Y2=0
cc_391 N_A_863_441#_c_571_n N_A_669_392#_M1014_g 0.00271673f $X=5.467 $Y=1.135
+ $X2=0 $Y2=0
cc_392 N_A_863_441#_c_573_n N_A_669_392#_M1014_g 0.00399403f $X=5.685 $Y=1.3
+ $X2=0 $Y2=0
cc_393 N_A_863_441#_M1012_g N_A_669_392#_c_660_n 0.00822975f $X=4.67 $Y=0.905
+ $X2=0 $Y2=0
cc_394 N_A_863_441#_M1012_g N_A_669_392#_c_661_n 0.006717f $X=4.67 $Y=0.905
+ $X2=0 $Y2=0
cc_395 N_A_863_441#_c_574_n N_A_669_392#_c_662_n 0.00172761f $X=4.405 $Y=2.465
+ $X2=0 $Y2=0
cc_396 N_A_863_441#_M1012_g N_A_669_392#_c_662_n 0.00737738f $X=4.67 $Y=0.905
+ $X2=0 $Y2=0
cc_397 N_A_863_441#_c_578_n N_A_669_392#_c_662_n 0.00733394f $X=5.265 $Y=2.19
+ $X2=0 $Y2=0
cc_398 N_A_863_441#_M1012_g N_A_669_392#_c_663_n 0.00979471f $X=4.67 $Y=0.905
+ $X2=0 $Y2=0
cc_399 N_A_863_441#_c_567_n N_A_669_392#_c_663_n 3.52118e-19 $X=6.125 $Y=1.465
+ $X2=0 $Y2=0
cc_400 N_A_863_441#_c_578_n N_A_669_392#_c_663_n 0.0233661f $X=5.265 $Y=2.19
+ $X2=0 $Y2=0
cc_401 N_A_863_441#_c_581_n N_A_669_392#_c_663_n 0.0026587f $X=5.43 $Y=2.105
+ $X2=0 $Y2=0
cc_402 N_A_863_441#_c_571_n N_A_669_392#_c_663_n 0.00275913f $X=5.467 $Y=1.135
+ $X2=0 $Y2=0
cc_403 N_A_863_441#_c_572_n N_A_669_392#_c_663_n 0.02787f $X=5.72 $Y=1.465 $X2=0
+ $Y2=0
cc_404 N_A_863_441#_M1012_g N_A_669_392#_c_664_n 0.0180926f $X=4.67 $Y=0.905
+ $X2=0 $Y2=0
cc_405 N_A_863_441#_c_567_n N_A_669_392#_c_664_n 0.0179536f $X=6.125 $Y=1.465
+ $X2=0 $Y2=0
cc_406 N_A_863_441#_c_578_n N_A_669_392#_c_664_n 0.00239819f $X=5.265 $Y=2.19
+ $X2=0 $Y2=0
cc_407 N_A_863_441#_c_581_n N_A_669_392#_c_664_n 4.65026e-19 $X=5.43 $Y=2.105
+ $X2=0 $Y2=0
cc_408 N_A_863_441#_c_571_n N_A_669_392#_c_664_n 2.32562e-19 $X=5.467 $Y=1.135
+ $X2=0 $Y2=0
cc_409 N_A_863_441#_c_572_n N_A_669_392#_c_664_n 0.00115796f $X=5.72 $Y=1.465
+ $X2=0 $Y2=0
cc_410 N_A_863_441#_c_578_n N_VPWR_M1015_d 0.00690748f $X=5.265 $Y=2.19 $X2=0
+ $Y2=0
cc_411 N_A_863_441#_c_574_n N_VPWR_c_752_n 0.017332f $X=4.405 $Y=2.465 $X2=0
+ $Y2=0
cc_412 N_A_863_441#_c_578_n N_VPWR_c_752_n 0.0505306f $X=5.265 $Y=2.19 $X2=0
+ $Y2=0
cc_413 N_A_863_441#_c_579_n N_VPWR_c_752_n 0.0330734f $X=5.43 $Y=2.815 $X2=0
+ $Y2=0
cc_414 N_A_863_441#_c_576_n N_VPWR_c_753_n 0.0100009f $X=6.215 $Y=1.765 $X2=0
+ $Y2=0
cc_415 N_A_863_441#_c_567_n N_VPWR_c_753_n 0.00871615f $X=6.125 $Y=1.465 $X2=0
+ $Y2=0
cc_416 N_A_863_441#_c_579_n N_VPWR_c_753_n 0.0515947f $X=5.43 $Y=2.815 $X2=0
+ $Y2=0
cc_417 N_A_863_441#_c_570_n N_VPWR_c_753_n 0.00970239f $X=5.57 $Y=1.94 $X2=0
+ $Y2=0
cc_418 N_A_863_441#_c_581_n N_VPWR_c_753_n 0.0356788f $X=5.43 $Y=2.105 $X2=0
+ $Y2=0
cc_419 N_A_863_441#_c_572_n N_VPWR_c_753_n 0.00451871f $X=5.72 $Y=1.465 $X2=0
+ $Y2=0
cc_420 N_A_863_441#_c_579_n N_VPWR_c_754_n 0.0172711f $X=5.43 $Y=2.815 $X2=0
+ $Y2=0
cc_421 N_A_863_441#_c_574_n N_VPWR_c_758_n 0.00429299f $X=4.405 $Y=2.465 $X2=0
+ $Y2=0
cc_422 N_A_863_441#_c_576_n N_VPWR_c_759_n 0.00439937f $X=6.215 $Y=1.765 $X2=0
+ $Y2=0
cc_423 N_A_863_441#_c_574_n N_VPWR_c_749_n 0.00879947f $X=4.405 $Y=2.465 $X2=0
+ $Y2=0
cc_424 N_A_863_441#_c_576_n N_VPWR_c_749_n 0.00847542f $X=6.215 $Y=1.765 $X2=0
+ $Y2=0
cc_425 N_A_863_441#_c_579_n N_VPWR_c_749_n 0.0142626f $X=5.43 $Y=2.815 $X2=0
+ $Y2=0
cc_426 N_A_863_441#_c_576_n Q 0.0169287f $X=6.215 $Y=1.765 $X2=0 $Y2=0
cc_427 N_A_863_441#_M1002_g Q 0.0247184f $X=6.22 $Y=0.74 $X2=0 $Y2=0
cc_428 N_A_863_441#_c_568_n Q 0.0212435f $X=6.125 $Y=1.3 $X2=0 $Y2=0
cc_429 N_A_863_441#_c_570_n Q 0.00534926f $X=5.57 $Y=1.94 $X2=0 $Y2=0
cc_430 N_A_863_441#_c_571_n Q 0.00495431f $X=5.467 $Y=1.135 $X2=0 $Y2=0
cc_431 N_A_863_441#_c_572_n Q 0.0130363f $X=5.72 $Y=1.465 $X2=0 $Y2=0
cc_432 N_A_863_441#_M1012_g N_VGND_c_845_n 0.00853602f $X=4.67 $Y=0.905 $X2=0
+ $Y2=0
cc_433 N_A_863_441#_c_569_n N_VGND_c_845_n 0.026273f $X=5.445 $Y=0.62 $X2=0
+ $Y2=0
cc_434 N_A_863_441#_M1002_g N_VGND_c_846_n 0.00647412f $X=6.22 $Y=0.74 $X2=0
+ $Y2=0
cc_435 N_A_863_441#_c_567_n N_VGND_c_846_n 0.0094508f $X=6.125 $Y=1.465 $X2=0
+ $Y2=0
cc_436 N_A_863_441#_c_569_n N_VGND_c_846_n 0.0523445f $X=5.445 $Y=0.62 $X2=0
+ $Y2=0
cc_437 N_A_863_441#_c_572_n N_VGND_c_846_n 0.00364403f $X=5.72 $Y=1.465 $X2=0
+ $Y2=0
cc_438 N_A_863_441#_M1012_g N_VGND_c_847_n 0.00380268f $X=4.67 $Y=0.905 $X2=0
+ $Y2=0
cc_439 N_A_863_441#_c_569_n N_VGND_c_851_n 0.011607f $X=5.445 $Y=0.62 $X2=0
+ $Y2=0
cc_440 N_A_863_441#_M1002_g N_VGND_c_852_n 0.00434272f $X=6.22 $Y=0.74 $X2=0
+ $Y2=0
cc_441 N_A_863_441#_M1012_g N_VGND_c_853_n 0.0045051f $X=4.67 $Y=0.905 $X2=0
+ $Y2=0
cc_442 N_A_863_441#_M1002_g N_VGND_c_853_n 0.00828958f $X=6.22 $Y=0.74 $X2=0
+ $Y2=0
cc_443 N_A_863_441#_c_569_n N_VGND_c_853_n 0.0128499f $X=5.445 $Y=0.62 $X2=0
+ $Y2=0
cc_444 N_A_669_392#_c_667_n N_VPWR_c_752_n 0.00616536f $X=5.205 $Y=1.885 $X2=0
+ $Y2=0
cc_445 N_A_669_392#_c_667_n N_VPWR_c_753_n 0.00459327f $X=5.205 $Y=1.885 $X2=0
+ $Y2=0
cc_446 N_A_669_392#_c_667_n N_VPWR_c_754_n 0.00445602f $X=5.205 $Y=1.885 $X2=0
+ $Y2=0
cc_447 N_A_669_392#_c_667_n N_VPWR_c_749_n 0.00864807f $X=5.205 $Y=1.885 $X2=0
+ $Y2=0
cc_448 N_A_669_392#_M1014_g N_VGND_c_845_n 0.00509156f $X=5.23 $Y=0.795 $X2=0
+ $Y2=0
cc_449 N_A_669_392#_c_660_n N_VGND_c_845_n 0.0201918f $X=4.51 $Y=0.93 $X2=0
+ $Y2=0
cc_450 N_A_669_392#_c_661_n N_VGND_c_845_n 0.00578369f $X=4.595 $Y=1.305 $X2=0
+ $Y2=0
cc_451 N_A_669_392#_c_663_n N_VGND_c_845_n 0.0214678f $X=5.15 $Y=1.47 $X2=0
+ $Y2=0
cc_452 N_A_669_392#_c_664_n N_VGND_c_845_n 0.0026557f $X=5.15 $Y=1.47 $X2=0
+ $Y2=0
cc_453 N_A_669_392#_M1014_g N_VGND_c_846_n 0.00366693f $X=5.23 $Y=0.795 $X2=0
+ $Y2=0
cc_454 N_A_669_392#_M1014_g N_VGND_c_851_n 0.00482438f $X=5.23 $Y=0.795 $X2=0
+ $Y2=0
cc_455 N_A_669_392#_M1014_g N_VGND_c_853_n 0.00512916f $X=5.23 $Y=0.795 $X2=0
+ $Y2=0
cc_456 N_A_669_392#_c_660_n N_VGND_c_853_n 0.0132675f $X=4.51 $Y=0.93 $X2=0
+ $Y2=0
cc_457 N_A_669_392#_c_660_n A_871_139# 0.0065047f $X=4.51 $Y=0.93 $X2=-0.19
+ $Y2=-0.245
cc_458 N_A_669_392#_c_661_n A_871_139# 8.22496e-19 $X=4.595 $Y=1.305 $X2=-0.19
+ $Y2=-0.245
cc_459 N_VPWR_c_753_n Q 0.0794554f $X=5.99 $Y=1.985 $X2=0 $Y2=0
cc_460 N_VPWR_c_759_n Q 0.014802f $X=6.48 $Y=3.33 $X2=0 $Y2=0
cc_461 N_VPWR_c_749_n Q 0.0122072f $X=6.48 $Y=3.33 $X2=0 $Y2=0
cc_462 Q N_VGND_c_846_n 0.0294766f $X=6.395 $Y=0.47 $X2=0 $Y2=0
cc_463 Q N_VGND_c_852_n 0.014787f $X=6.395 $Y=0.47 $X2=0 $Y2=0
cc_464 Q N_VGND_c_853_n 0.012183f $X=6.395 $Y=0.47 $X2=0 $Y2=0
