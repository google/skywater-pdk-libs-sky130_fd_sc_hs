* File: sky130_fd_sc_hs__dlrbp_2.pex.spice
* Created: Thu Aug 27 20:41:18 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HS__DLRBP_2%D 3 5 7 8
c36 5 0 3.00127e-19 $X=0.505 $Y=1.885
r37 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.59
+ $Y=1.615 $X2=0.59 $Y2=1.615
r38 8 12 4.53993 $w=3.28e-07 $l=1.3e-07 $layer=LI1_cond $X=0.72 $Y=1.615
+ $X2=0.59 $Y2=1.615
r39 5 11 55.362 $w=3.01e-07 $l=3.07409e-07 $layer=POLY_cond $X=0.505 $Y=1.885
+ $X2=0.585 $Y2=1.615
r40 5 7 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=0.505 $Y=1.885
+ $X2=0.505 $Y2=2.38
r41 1 11 38.5481 $w=3.01e-07 $l=2.05122e-07 $layer=POLY_cond $X=0.495 $Y=1.45
+ $X2=0.585 $Y2=1.615
r42 1 3 315.351 $w=1.5e-07 $l=6.15e-07 $layer=POLY_cond $X=0.495 $Y=1.45
+ $X2=0.495 $Y2=0.835
.ends

.subckt PM_SKY130_FD_SC_HS__DLRBP_2%GATE 3 5 6 8 9 12 14
c40 14 0 2.61276e-20 $X=1.13 $Y=1.22
c41 9 0 1.09742e-19 $X=1.2 $Y=1.295
r42 12 15 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.13 $Y=1.385
+ $X2=1.13 $Y2=1.55
r43 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.13 $Y=1.385
+ $X2=1.13 $Y2=1.22
r44 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.13
+ $Y=1.385 $X2=1.13 $Y2=1.385
r45 9 13 3.3458 $w=3.08e-07 $l=9e-08 $layer=LI1_cond $X=1.13 $Y=1.295 $X2=1.13
+ $Y2=1.385
r46 6 8 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=1.125 $Y=1.885
+ $X2=1.125 $Y2=2.38
r47 5 6 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=1.125 $Y=1.795 $X2=1.125
+ $Y2=1.885
r48 5 15 95.2339 $w=1.8e-07 $l=2.45e-07 $layer=POLY_cond $X=1.125 $Y=1.795
+ $X2=1.125 $Y2=1.55
r49 3 14 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.075 $Y=0.74
+ $X2=1.075 $Y2=1.22
.ends

.subckt PM_SKY130_FD_SC_HS__DLRBP_2%A_230_74# 1 2 7 9 10 11 13 14 16 17 19 20 21
+ 25 30 31 33 35 36 39 46 49 51 57
c141 35 0 6.32864e-20 $X=3.73 $Y=0.345
c142 31 0 2.61276e-20 $X=2.81 $Y=0.665
c143 21 0 1.87347e-19 $X=3.265 $Y=1.765
c144 20 0 8.05161e-20 $X=3.715 $Y=1.765
c145 17 0 1.67788e-19 $X=3.175 $Y=1.885
r146 50 57 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=1.7 $Y=1.505 $X2=1.7
+ $Y2=1.415
r147 49 52 8.69073 $w=4.08e-07 $l=1.65e-07 $layer=LI1_cond $X=1.66 $Y=1.505
+ $X2=1.66 $Y2=1.67
r148 49 51 8.69073 $w=4.08e-07 $l=1.65e-07 $layer=LI1_cond $X=1.66 $Y=1.505
+ $X2=1.66 $Y2=1.34
r149 49 50 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.7
+ $Y=1.505 $X2=1.7 $Y2=1.505
r150 44 46 7.60612 $w=2.48e-07 $l=1.65e-07 $layer=LI1_cond $X=1.375 $Y=2.065
+ $X2=1.54 $Y2=2.065
r151 42 51 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=1.54 $Y=1.01
+ $X2=1.54 $Y2=1.34
r152 41 42 13.823 $w=4.98e-07 $l=3.45e-07 $layer=LI1_cond $X=1.375 $Y=0.665
+ $X2=1.375 $Y2=1.01
r153 39 41 3.58824 $w=4.98e-07 $l=1.5e-07 $layer=LI1_cond $X=1.375 $Y=0.515
+ $X2=1.375 $Y2=0.665
r154 36 63 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.73 $Y=0.345
+ $X2=3.73 $Y2=0.51
r155 35 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.73
+ $Y=0.345 $X2=3.73 $Y2=0.345
r156 33 55 18.4631 $w=1.68e-07 $l=2.83e-07 $layer=LI1_cond $X=2.895 $Y=0.382
+ $X2=2.895 $Y2=0.665
r157 33 35 33.8954 $w=2.53e-07 $l=7.5e-07 $layer=LI1_cond $X=2.98 $Y=0.382
+ $X2=3.73 $Y2=0.382
r158 32 41 7.15667 $w=1.7e-07 $l=2.5e-07 $layer=LI1_cond $X=1.625 $Y=0.665
+ $X2=1.375 $Y2=0.665
r159 31 55 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.81 $Y=0.665
+ $X2=2.895 $Y2=0.665
r160 31 32 77.3102 $w=1.68e-07 $l=1.185e-06 $layer=LI1_cond $X=2.81 $Y=0.665
+ $X2=1.625 $Y2=0.665
r161 30 46 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.54 $Y=1.94
+ $X2=1.54 $Y2=2.065
r162 30 52 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=1.54 $Y=1.94
+ $X2=1.54 $Y2=1.67
r163 25 63 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=3.79 $Y=0.83
+ $X2=3.79 $Y2=0.51
r164 23 25 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=3.79 $Y=1.69
+ $X2=3.79 $Y2=0.83
r165 20 23 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.715 $Y=1.765
+ $X2=3.79 $Y2=1.69
r166 20 21 230.745 $w=1.5e-07 $l=4.5e-07 $layer=POLY_cond $X=3.715 $Y=1.765
+ $X2=3.265 $Y2=1.765
r167 17 21 26.9307 $w=1.5e-07 $l=1.58745e-07 $layer=POLY_cond $X=3.175 $Y=1.885
+ $X2=3.265 $Y2=1.765
r168 17 19 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=3.175 $Y=1.885
+ $X2=3.175 $Y2=2.46
r169 14 16 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=2.185 $Y=1.885
+ $X2=2.185 $Y2=2.38
r170 11 26 53.0007 $w=1.77e-07 $l=1.94936e-07 $layer=POLY_cond $X=2.175 $Y=1.225
+ $X2=2.185 $Y2=1.415
r171 11 13 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=2.175 $Y=1.225
+ $X2=2.175 $Y2=0.78
r172 10 14 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=2.185 $Y=1.795
+ $X2=2.185 $Y2=1.885
r173 9 26 20.0833 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=2.185 $Y=1.49
+ $X2=2.185 $Y2=1.415
r174 9 10 118.556 $w=1.8e-07 $l=3.05e-07 $layer=POLY_cond $X=2.185 $Y=1.49
+ $X2=2.185 $Y2=1.795
r175 8 57 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.865 $Y=1.415
+ $X2=1.7 $Y2=1.415
r176 7 26 6.7465 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=2.095 $Y=1.415
+ $X2=2.185 $Y2=1.415
r177 7 8 117.936 $w=1.5e-07 $l=2.3e-07 $layer=POLY_cond $X=2.095 $Y=1.415
+ $X2=1.865 $Y2=1.415
r178 2 44 600 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=1.2
+ $Y=1.96 $X2=1.375 $Y2=2.105
r179 1 39 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.15
+ $Y=0.37 $X2=1.29 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__DLRBP_2%A_27_112# 1 2 7 9 12 14 20 21 22 25 28 30 31
c82 28 0 1.90385e-19 $X=0.265 $Y=1.13
c83 25 0 1.97327e-19 $X=2.65 $Y=1.635
c84 21 0 1.67788e-19 $X=2.485 $Y=2.445
r85 30 31 8.51103 $w=3.58e-07 $l=1.65e-07 $layer=LI1_cond $X=0.265 $Y=2.115
+ $X2=0.265 $Y2=1.95
r86 28 31 53.4973 $w=1.68e-07 $l=8.2e-07 $layer=LI1_cond $X=0.17 $Y=1.13
+ $X2=0.17 $Y2=1.95
r87 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.65
+ $Y=1.635 $X2=2.65 $Y2=1.635
r88 23 25 26.11 $w=3.18e-07 $l=7.25e-07 $layer=LI1_cond $X=2.645 $Y=2.36
+ $X2=2.645 $Y2=1.635
r89 21 23 7.68211 $w=1.7e-07 $l=1.9799e-07 $layer=LI1_cond $X=2.485 $Y=2.445
+ $X2=2.645 $Y2=2.36
r90 21 22 133.091 $w=1.68e-07 $l=2.04e-06 $layer=LI1_cond $X=2.485 $Y=2.445
+ $X2=0.445 $Y2=2.445
r91 20 22 8.02311 $w=1.7e-07 $l=2.18403e-07 $layer=LI1_cond $X=0.265 $Y=2.36
+ $X2=0.445 $Y2=2.445
r92 19 30 0.480185 $w=3.58e-07 $l=1.5e-08 $layer=LI1_cond $X=0.265 $Y=2.13
+ $X2=0.265 $Y2=2.115
r93 19 20 7.36283 $w=3.58e-07 $l=2.3e-07 $layer=LI1_cond $X=0.265 $Y=2.13
+ $X2=0.265 $Y2=2.36
r94 14 28 8.99121 $w=3.58e-07 $l=1.8e-07 $layer=LI1_cond $X=0.265 $Y=0.95
+ $X2=0.265 $Y2=1.13
r95 14 16 3.89722 $w=3.6e-07 $l=1.15e-07 $layer=LI1_cond $X=0.265 $Y=0.95
+ $X2=0.265 $Y2=0.835
r96 10 26 38.5615 $w=3.23e-07 $l=2.11069e-07 $layer=POLY_cond $X=2.77 $Y=1.47
+ $X2=2.665 $Y2=1.635
r97 10 12 384.574 $w=1.5e-07 $l=7.5e-07 $layer=POLY_cond $X=2.77 $Y=1.47
+ $X2=2.77 $Y2=0.72
r98 7 26 51.2457 $w=3.23e-07 $l=2.91548e-07 $layer=POLY_cond $X=2.755 $Y=1.885
+ $X2=2.665 $Y2=1.635
r99 7 9 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=2.755 $Y=1.885
+ $X2=2.755 $Y2=2.46
r100 2 30 300 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.96 $X2=0.28 $Y2=2.115
r101 1 16 182 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.56 $X2=0.28 $Y2=0.835
.ends

.subckt PM_SKY130_FD_SC_HS__DLRBP_2%A_363_82# 1 2 9 10 12 13 14 15 18 19 20 23
+ 32 34 38 41
c116 38 0 9.98003e-21 $X=3.22 $Y=1.315
c117 34 0 8.05161e-20 $X=3.18 $Y=1.215
r118 38 41 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.22 $Y=1.315
+ $X2=3.22 $Y2=1.15
r119 37 39 8.69073 $w=4.08e-07 $l=1.65e-07 $layer=LI1_cond $X=3.18 $Y=1.315
+ $X2=3.18 $Y2=1.48
r120 37 38 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.22
+ $Y=1.315 $X2=3.22 $Y2=1.315
r121 34 37 2.81084 $w=4.08e-07 $l=1e-07 $layer=LI1_cond $X=3.18 $Y=1.215
+ $X2=3.18 $Y2=1.315
r122 30 32 7.37564 $w=2.48e-07 $l=1.6e-07 $layer=LI1_cond $X=1.96 $Y=2.065
+ $X2=2.12 $Y2=2.065
r123 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.87
+ $Y=2.215 $X2=3.87 $Y2=2.215
r124 21 23 24.0965 $w=3.28e-07 $l=6.9e-07 $layer=LI1_cond $X=3.87 $Y=2.905
+ $X2=3.87 $Y2=2.215
r125 19 21 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.705 $Y=2.99
+ $X2=3.87 $Y2=2.905
r126 19 20 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=3.705 $Y=2.99
+ $X2=3.145 $Y2=2.99
r127 18 20 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.06 $Y=2.905
+ $X2=3.145 $Y2=2.99
r128 18 39 92.9679 $w=1.68e-07 $l=1.425e-06 $layer=LI1_cond $X=3.06 $Y=2.905
+ $X2=3.06 $Y2=1.48
r129 16 27 7.83486 $w=3.27e-07 $l=2.95212e-07 $layer=LI1_cond $X=2.205 $Y=1.215
+ $X2=2 $Y2=1.005
r130 15 34 5.92876 $w=1.7e-07 $l=2.05e-07 $layer=LI1_cond $X=2.975 $Y=1.215
+ $X2=3.18 $Y2=1.215
r131 15 16 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=2.975 $Y=1.215
+ $X2=2.205 $Y2=1.215
r132 14 32 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.12 $Y=1.94
+ $X2=2.12 $Y2=2.065
r133 13 16 5.97199 $w=3.27e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.12 $Y=1.3
+ $X2=2.205 $Y2=1.215
r134 13 14 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=2.12 $Y=1.3 $X2=2.12
+ $Y2=1.94
r135 10 24 50.1894 $w=3.66e-07 $l=3.02903e-07 $layer=POLY_cond $X=3.71 $Y=2.465
+ $X2=3.827 $Y2=2.215
r136 10 12 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=3.71 $Y=2.465
+ $X2=3.71 $Y2=2.75
r137 9 41 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=3.13 $Y=0.72
+ $X2=3.13 $Y2=1.15
r138 2 30 600 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=1.815
+ $Y=1.96 $X2=1.96 $Y2=2.105
r139 1 27 182 $w=1.7e-07 $l=6.63551e-07 $layer=licon1_NDIFF $count=1 $X=1.815
+ $Y=0.41 $X2=1.96 $Y2=1.005
.ends

.subckt PM_SKY130_FD_SC_HS__DLRBP_2%A_821_98# 1 2 7 9 11 12 14 17 19 21 24 26 28
+ 29 30 31 33 36 40 42 43 50 56 58 60 62 65 66 67
c159 67 0 1.03706e-19 $X=5.33 $Y=1.72
c160 58 0 1.02956e-19 $X=5.955 $Y=1.805
c161 43 0 1.27212e-20 $X=5.095 $Y=2.155
c162 31 0 1.30305e-19 $X=7.615 $Y=1.765
c163 24 0 1.93666e-19 $X=6.53 $Y=0.74
c164 7 0 6.32864e-20 $X=4.18 $Y=1.115
r165 77 78 6.59453 $w=4.02e-07 $l=5.5e-08 $layer=POLY_cond $X=6.1 $Y=1.532
+ $X2=6.155 $Y2=1.532
r166 70 71 5.27442 $w=4.68e-07 $l=1.65e-07 $layer=LI1_cond $X=5.33 $Y=2.155
+ $X2=5.33 $Y2=2.32
r167 69 70 4.32624 $w=4.68e-07 $l=1.7e-07 $layer=LI1_cond $X=5.33 $Y=1.985
+ $X2=5.33 $Y2=2.155
r168 66 69 4.58073 $w=4.68e-07 $l=1.8e-07 $layer=LI1_cond $X=5.33 $Y=1.805
+ $X2=5.33 $Y2=1.985
r169 66 67 7.30169 $w=4.68e-07 $l=8.5e-08 $layer=LI1_cond $X=5.33 $Y=1.805
+ $X2=5.33 $Y2=1.72
r170 65 67 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=5.18 $Y=1.13
+ $X2=5.18 $Y2=1.72
r171 63 80 8.99254 $w=4.02e-07 $l=7.5e-08 $layer=POLY_cond $X=6.53 $Y=1.532
+ $X2=6.605 $Y2=1.532
r172 63 78 44.9627 $w=4.02e-07 $l=3.75e-07 $layer=POLY_cond $X=6.53 $Y=1.532
+ $X2=6.155 $Y2=1.532
r173 62 63 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.53
+ $Y=1.465 $X2=6.53 $Y2=1.465
r174 60 74 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=6.04 $Y=1.465
+ $X2=6.04 $Y2=1.805
r175 60 62 14.1436 $w=3.28e-07 $l=4.05e-07 $layer=LI1_cond $X=6.125 $Y=1.465
+ $X2=6.53 $Y2=1.465
r176 59 66 6.76998 $w=1.7e-07 $l=2.35e-07 $layer=LI1_cond $X=5.565 $Y=1.805
+ $X2=5.33 $Y2=1.805
r177 58 74 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.955 $Y=1.805
+ $X2=6.04 $Y2=1.805
r178 58 59 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=5.955 $Y=1.805
+ $X2=5.565 $Y2=1.805
r179 56 71 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=5.4 $Y=2.4 $X2=5.4
+ $Y2=2.32
r180 48 65 11.1798 $w=4.73e-07 $l=2.37e-07 $layer=LI1_cond $X=5.027 $Y=0.893
+ $X2=5.027 $Y2=1.13
r181 48 50 9.51827 $w=4.73e-07 $l=3.78e-07 $layer=LI1_cond $X=5.027 $Y=0.893
+ $X2=5.027 $Y2=0.515
r182 45 46 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.41
+ $Y=2.155 $X2=4.41 $Y2=2.155
r183 43 70 2.80859 $w=3.3e-07 $l=2.35e-07 $layer=LI1_cond $X=5.095 $Y=2.155
+ $X2=5.33 $Y2=2.155
r184 43 45 23.9219 $w=3.28e-07 $l=6.85e-07 $layer=LI1_cond $X=5.095 $Y=2.155
+ $X2=4.41 $Y2=2.155
r185 38 40 71.7872 $w=1.5e-07 $l=1.4e-07 $layer=POLY_cond $X=4.18 $Y=1.19
+ $X2=4.32 $Y2=1.19
r186 34 42 37.0704 $w=1.5e-07 $l=2.36947e-07 $layer=POLY_cond $X=7.625 $Y=1.3
+ $X2=7.615 $Y2=1.532
r187 34 36 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=7.625 $Y=1.3
+ $X2=7.625 $Y2=0.79
r188 31 42 37.0704 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=7.615 $Y=1.765
+ $X2=7.615 $Y2=1.532
r189 31 33 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=7.615 $Y=1.765
+ $X2=7.615 $Y2=2.34
r190 30 80 12.4798 $w=4.02e-07 $l=1.1887e-07 $layer=POLY_cond $X=6.695 $Y=1.465
+ $X2=6.605 $Y2=1.532
r191 29 42 5.03009 $w=3.3e-07 $l=1.1887e-07 $layer=POLY_cond $X=7.525 $Y=1.465
+ $X2=7.615 $Y2=1.532
r192 29 30 145.135 $w=3.3e-07 $l=8.3e-07 $layer=POLY_cond $X=7.525 $Y=1.465
+ $X2=6.695 $Y2=1.465
r193 26 80 25.9839 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=6.605 $Y=1.765
+ $X2=6.605 $Y2=1.532
r194 26 28 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=6.605 $Y=1.765
+ $X2=6.605 $Y2=2.4
r195 22 63 25.9839 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=6.53 $Y=1.3
+ $X2=6.53 $Y2=1.532
r196 22 24 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=6.53 $Y=1.3
+ $X2=6.53 $Y2=0.74
r197 19 78 25.9839 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=6.155 $Y=1.765
+ $X2=6.155 $Y2=1.532
r198 19 21 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=6.155 $Y=1.765
+ $X2=6.155 $Y2=2.4
r199 15 77 25.9839 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=6.1 $Y=1.3 $X2=6.1
+ $Y2=1.532
r200 15 17 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=6.1 $Y=1.3 $X2=6.1
+ $Y2=0.74
r201 12 46 63.2868 $w=2.84e-07 $l=3.31738e-07 $layer=POLY_cond $X=4.365 $Y=2.465
+ $X2=4.41 $Y2=2.155
r202 12 14 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=4.365 $Y=2.465
+ $X2=4.365 $Y2=2.75
r203 11 46 38.6777 $w=2.84e-07 $l=2.05122e-07 $layer=POLY_cond $X=4.32 $Y=1.99
+ $X2=4.41 $Y2=2.155
r204 10 40 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.32 $Y=1.265
+ $X2=4.32 $Y2=1.19
r205 10 11 371.755 $w=1.5e-07 $l=7.25e-07 $layer=POLY_cond $X=4.32 $Y=1.265
+ $X2=4.32 $Y2=1.99
r206 7 38 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.18 $Y=1.115
+ $X2=4.18 $Y2=1.19
r207 7 9 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=4.18 $Y=1.115 $X2=4.18
+ $Y2=0.83
r208 2 69 600 $w=1.7e-07 $l=2.62678e-07 $layer=licon1_PDIFF $count=1 $X=5.2
+ $Y=1.84 $X2=5.4 $Y2=1.985
r209 2 56 300 $w=1.7e-07 $l=6.5238e-07 $layer=licon1_PDIFF $count=2 $X=5.2
+ $Y=1.84 $X2=5.4 $Y2=2.4
r210 1 50 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=4.81
+ $Y=0.37 $X2=4.955 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__DLRBP_2%A_641_80# 1 2 7 9 12 15 16 22 25 26 27 32
c83 7 0 2.50955e-19 $X=5.125 $Y=1.765
r84 32 35 7.92305 $w=3.18e-07 $l=2.2e-07 $layer=LI1_cond $X=4.765 $Y=1.515
+ $X2=4.765 $Y2=1.735
r85 32 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.77
+ $Y=1.515 $X2=4.77 $Y2=1.515
r86 28 30 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=3.4 $Y=1.735
+ $X2=3.655 $Y2=1.735
r87 27 30 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=3.74 $Y=1.735
+ $X2=3.655 $Y2=1.735
r88 26 35 4.44149 $w=1.7e-07 $l=1.6e-07 $layer=LI1_cond $X=4.605 $Y=1.735
+ $X2=4.765 $Y2=1.735
r89 26 27 56.4332 $w=1.68e-07 $l=8.65e-07 $layer=LI1_cond $X=4.605 $Y=1.735
+ $X2=3.74 $Y2=1.735
r90 25 30 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.655 $Y=1.65
+ $X2=3.655 $Y2=1.735
r91 24 25 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=3.655 $Y=0.96
+ $X2=3.655 $Y2=1.65
r92 20 28 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.4 $Y=1.82 $X2=3.4
+ $Y2=1.735
r93 20 22 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=3.4 $Y=1.82 $X2=3.4
+ $Y2=2.11
r94 16 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.57 $Y=0.875
+ $X2=3.655 $Y2=0.96
r95 16 18 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=3.57 $Y=0.875
+ $X2=3.46 $Y2=0.875
r96 15 33 46.3382 $w=3.3e-07 $l=2.65e-07 $layer=POLY_cond $X=5.035 $Y=1.515
+ $X2=4.77 $Y2=1.515
r97 10 15 44.1289 $w=1.9e-07 $l=1.79374e-07 $layer=POLY_cond $X=5.17 $Y=1.35
+ $X2=5.14 $Y2=1.515
r98 10 12 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=5.17 $Y=1.35
+ $X2=5.17 $Y2=0.74
r99 7 15 65.692 $w=1.9e-07 $l=2.57391e-07 $layer=POLY_cond $X=5.125 $Y=1.765
+ $X2=5.14 $Y2=1.515
r100 7 9 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=5.125 $Y=1.765
+ $X2=5.125 $Y2=2.4
r101 2 22 300 $w=1.7e-07 $l=2.12132e-07 $layer=licon1_PDIFF $count=2 $X=3.25
+ $Y=1.96 $X2=3.4 $Y2=2.11
r102 1 18 182 $w=1.7e-07 $l=5.88855e-07 $layer=licon1_NDIFF $count=1 $X=3.205
+ $Y=0.4 $X2=3.46 $Y2=0.875
.ends

.subckt PM_SKY130_FD_SC_HS__DLRBP_2%RESET_B 1 3 4 6 7 11
c34 11 0 1.47999e-19 $X=5.62 $Y=1.385
c35 4 0 1.27212e-20 $X=5.625 $Y=1.765
c36 1 0 2.71532e-19 $X=5.56 $Y=1.22
r37 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.62
+ $Y=1.385 $X2=5.62 $Y2=1.385
r38 7 11 3.11471 $w=3.68e-07 $l=1e-07 $layer=LI1_cond $X=5.52 $Y=1.365 $X2=5.62
+ $Y2=1.365
r39 4 10 77.2841 $w=2.7e-07 $l=3.82492e-07 $layer=POLY_cond $X=5.625 $Y=1.765
+ $X2=5.62 $Y2=1.385
r40 4 6 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=5.625 $Y=1.765
+ $X2=5.625 $Y2=2.4
r41 1 10 38.9026 $w=2.7e-07 $l=1.92678e-07 $layer=POLY_cond $X=5.56 $Y=1.22
+ $X2=5.62 $Y2=1.385
r42 1 3 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=5.56 $Y=1.22 $X2=5.56
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HS__DLRBP_2%A_1449_368# 1 2 7 9 12 14 16 19 23 26 29 35
+ 38 39 43
c70 38 0 1.93666e-19 $X=7.41 $Y=1.13
c71 7 0 1.00299e-19 $X=8.165 $Y=1.765
r72 43 44 1.23274 $w=3.91e-07 $l=1e-08 $layer=POLY_cond $X=8.615 $Y=1.532
+ $X2=8.625 $Y2=1.532
r73 42 43 51.7749 $w=3.91e-07 $l=4.2e-07 $layer=POLY_cond $X=8.195 $Y=1.532
+ $X2=8.615 $Y2=1.532
r74 41 42 3.69821 $w=3.91e-07 $l=3e-08 $layer=POLY_cond $X=8.165 $Y=1.532
+ $X2=8.195 $Y2=1.532
r75 36 41 10.4783 $w=3.91e-07 $l=8.5e-08 $layer=POLY_cond $X=8.08 $Y=1.532
+ $X2=8.165 $Y2=1.532
r76 35 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.08
+ $Y=1.465 $X2=8.08 $Y2=1.465
r77 33 39 1.11842 $w=3.3e-07 $l=1.55e-07 $layer=LI1_cond $X=7.555 $Y=1.465
+ $X2=7.4 $Y2=1.465
r78 33 35 18.3343 $w=3.28e-07 $l=5.25e-07 $layer=LI1_cond $X=7.555 $Y=1.465
+ $X2=8.08 $Y2=1.465
r79 29 31 26.3947 $w=3.08e-07 $l=7.1e-07 $layer=LI1_cond $X=7.4 $Y=1.985 $X2=7.4
+ $Y2=2.695
r80 27 39 5.44021 $w=3.1e-07 $l=1.65e-07 $layer=LI1_cond $X=7.4 $Y=1.63 $X2=7.4
+ $Y2=1.465
r81 27 29 13.1973 $w=3.08e-07 $l=3.55e-07 $layer=LI1_cond $X=7.4 $Y=1.63 $X2=7.4
+ $Y2=1.985
r82 26 39 5.44021 $w=3.1e-07 $l=1.65e-07 $layer=LI1_cond $X=7.4 $Y=1.3 $X2=7.4
+ $Y2=1.465
r83 26 38 6.31985 $w=3.08e-07 $l=1.7e-07 $layer=LI1_cond $X=7.4 $Y=1.3 $X2=7.4
+ $Y2=1.13
r84 21 38 5.81909 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=7.41 $Y=0.965
+ $X2=7.41 $Y2=1.13
r85 21 23 12.2229 $w=3.28e-07 $l=3.5e-07 $layer=LI1_cond $X=7.41 $Y=0.965
+ $X2=7.41 $Y2=0.615
r86 17 44 25.3065 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=8.625 $Y=1.3
+ $X2=8.625 $Y2=1.532
r87 17 19 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=8.625 $Y=1.3
+ $X2=8.625 $Y2=0.74
r88 14 43 25.3065 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=8.615 $Y=1.765
+ $X2=8.615 $Y2=1.532
r89 14 16 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=8.615 $Y=1.765
+ $X2=8.615 $Y2=2.4
r90 10 42 25.3065 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=8.195 $Y=1.3
+ $X2=8.195 $Y2=1.532
r91 10 12 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=8.195 $Y=1.3
+ $X2=8.195 $Y2=0.74
r92 7 41 25.3065 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=8.165 $Y=1.765
+ $X2=8.165 $Y2=1.532
r93 7 9 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=8.165 $Y=1.765
+ $X2=8.165 $Y2=2.4
r94 2 31 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=7.245
+ $Y=1.84 $X2=7.39 $Y2=2.695
r95 2 29 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=7.245
+ $Y=1.84 $X2=7.39 $Y2=1.985
r96 1 23 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=7.265
+ $Y=0.47 $X2=7.41 $Y2=0.615
.ends

.subckt PM_SKY130_FD_SC_HS__DLRBP_2%VPWR 1 2 3 4 5 6 7 26 30 34 40 44 48 50 55
+ 56 58 59 60 62 70 82 86 92 95 98 105 109
r110 108 109 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r111 105 106 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r112 98 101 9.62469 $w=6.38e-07 $l=5.15e-07 $layer=LI1_cond $X=4.745 $Y=2.815
+ $X2=4.745 $Y2=3.33
r113 95 96 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r114 92 93 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r115 90 109 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=3.33
+ $X2=8.88 $Y2=3.33
r116 90 106 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=3.33
+ $X2=7.92 $Y2=3.33
r117 89 90 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=3.33 $X2=8.4
+ $Y2=3.33
r118 87 105 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.055 $Y=3.33
+ $X2=7.89 $Y2=3.33
r119 87 89 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=8.055 $Y=3.33
+ $X2=8.4 $Y2=3.33
r120 86 108 4.01252 $w=1.7e-07 $l=1.82e-07 $layer=LI1_cond $X=8.755 $Y=3.33
+ $X2=8.937 $Y2=3.33
r121 86 89 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=8.755 $Y=3.33
+ $X2=8.4 $Y2=3.33
r122 85 106 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=7.92 $Y2=3.33
r123 84 85 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r124 82 105 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.725 $Y=3.33
+ $X2=7.89 $Y2=3.33
r125 82 84 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=7.725 $Y=3.33
+ $X2=7.44 $Y2=3.33
r126 81 85 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=7.44 $Y2=3.33
r127 80 81 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r128 78 81 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=6.48 $Y2=3.33
r129 77 78 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r130 75 101 8.73481 $w=1.7e-07 $l=3.2e-07 $layer=LI1_cond $X=5.065 $Y=3.33
+ $X2=4.745 $Y2=3.33
r131 75 77 29.6845 $w=1.68e-07 $l=4.55e-07 $layer=LI1_cond $X=5.065 $Y=3.33
+ $X2=5.52 $Y2=3.33
r132 74 96 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=2.64 $Y2=3.33
r133 73 74 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r134 71 95 9.23004 $w=1.7e-07 $l=1.83e-07 $layer=LI1_cond $X=2.695 $Y=3.33
+ $X2=2.512 $Y2=3.33
r135 71 73 90.3583 $w=1.68e-07 $l=1.385e-06 $layer=LI1_cond $X=2.695 $Y=3.33
+ $X2=4.08 $Y2=3.33
r136 70 101 8.73481 $w=1.7e-07 $l=3.2e-07 $layer=LI1_cond $X=4.425 $Y=3.33
+ $X2=4.745 $Y2=3.33
r137 70 73 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=4.425 $Y=3.33
+ $X2=4.08 $Y2=3.33
r138 69 96 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r139 68 69 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r140 66 69 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.16 $Y2=3.33
r141 66 93 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r142 65 68 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.2 $Y=3.33 $X2=2.16
+ $Y2=3.33
r143 65 66 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r144 63 92 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.98 $Y=3.33
+ $X2=0.815 $Y2=3.33
r145 63 65 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=0.98 $Y=3.33
+ $X2=1.2 $Y2=3.33
r146 62 95 9.23004 $w=1.7e-07 $l=1.82e-07 $layer=LI1_cond $X=2.33 $Y=3.33
+ $X2=2.512 $Y2=3.33
r147 62 68 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=2.33 $Y=3.33
+ $X2=2.16 $Y2=3.33
r148 60 78 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=5.52 $Y2=3.33
r149 60 74 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=4.08 $Y2=3.33
r150 60 101 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r151 58 80 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=6.665 $Y=3.33
+ $X2=6.48 $Y2=3.33
r152 58 59 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.665 $Y=3.33
+ $X2=6.83 $Y2=3.33
r153 57 84 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=6.995 $Y=3.33
+ $X2=7.44 $Y2=3.33
r154 57 59 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.995 $Y=3.33
+ $X2=6.83 $Y2=3.33
r155 55 77 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=5.735 $Y=3.33
+ $X2=5.52 $Y2=3.33
r156 55 56 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.735 $Y=3.33
+ $X2=5.9 $Y2=3.33
r157 54 80 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=6.065 $Y=3.33
+ $X2=6.48 $Y2=3.33
r158 54 56 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.065 $Y=3.33
+ $X2=5.9 $Y2=3.33
r159 50 53 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=8.88 $Y=1.985
+ $X2=8.88 $Y2=2.815
r160 48 108 3.13065 $w=2.5e-07 $l=1.09864e-07 $layer=LI1_cond $X=8.88 $Y=3.245
+ $X2=8.937 $Y2=3.33
r161 48 53 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=8.88 $Y=3.245
+ $X2=8.88 $Y2=2.815
r162 44 47 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=7.89 $Y=1.985
+ $X2=7.89 $Y2=2.695
r163 42 105 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.89 $Y=3.245
+ $X2=7.89 $Y2=3.33
r164 42 47 19.2074 $w=3.28e-07 $l=5.5e-07 $layer=LI1_cond $X=7.89 $Y=3.245
+ $X2=7.89 $Y2=2.695
r165 38 59 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.83 $Y=3.245
+ $X2=6.83 $Y2=3.33
r166 38 40 32.8272 $w=3.28e-07 $l=9.4e-07 $layer=LI1_cond $X=6.83 $Y=3.245
+ $X2=6.83 $Y2=2.305
r167 34 37 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=5.9 $Y=2.145
+ $X2=5.9 $Y2=2.825
r168 32 56 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.9 $Y=3.245 $X2=5.9
+ $Y2=3.33
r169 32 37 14.6675 $w=3.28e-07 $l=4.2e-07 $layer=LI1_cond $X=5.9 $Y=3.245
+ $X2=5.9 $Y2=2.825
r170 28 95 1.2012 $w=3.65e-07 $l=8.5e-08 $layer=LI1_cond $X=2.512 $Y=3.245
+ $X2=2.512 $Y2=3.33
r171 28 30 14.5239 $w=3.63e-07 $l=4.6e-07 $layer=LI1_cond $X=2.512 $Y=3.245
+ $X2=2.512 $Y2=2.785
r172 24 92 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.815 $Y=3.245
+ $X2=0.815 $Y2=3.33
r173 24 26 13.2706 $w=3.28e-07 $l=3.8e-07 $layer=LI1_cond $X=0.815 $Y=3.245
+ $X2=0.815 $Y2=2.865
r174 7 53 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=8.69
+ $Y=1.84 $X2=8.84 $Y2=2.815
r175 7 50 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=8.69
+ $Y=1.84 $X2=8.84 $Y2=1.985
r176 6 47 400 $w=1.7e-07 $l=9.4975e-07 $layer=licon1_PDIFF $count=1 $X=7.69
+ $Y=1.84 $X2=7.89 $Y2=2.695
r177 6 44 400 $w=1.7e-07 $l=2.62678e-07 $layer=licon1_PDIFF $count=1 $X=7.69
+ $Y=1.84 $X2=7.89 $Y2=1.985
r178 5 40 300 $w=1.7e-07 $l=5.34766e-07 $layer=licon1_PDIFF $count=2 $X=6.68
+ $Y=1.84 $X2=6.83 $Y2=2.305
r179 4 37 400 $w=1.7e-07 $l=1.08038e-06 $layer=licon1_PDIFF $count=1 $X=5.7
+ $Y=1.84 $X2=5.9 $Y2=2.825
r180 4 34 400 $w=1.7e-07 $l=3.9246e-07 $layer=licon1_PDIFF $count=1 $X=5.7
+ $Y=1.84 $X2=5.9 $Y2=2.145
r181 3 98 600 $w=1.7e-07 $l=4.20595e-07 $layer=licon1_PDIFF $count=1 $X=4.44
+ $Y=2.54 $X2=4.745 $Y2=2.815
r182 2 30 600 $w=1.7e-07 $l=9.4174e-07 $layer=licon1_PDIFF $count=1 $X=2.26
+ $Y=1.96 $X2=2.51 $Y2=2.785
r183 1 26 600 $w=1.7e-07 $l=1.01573e-06 $layer=licon1_PDIFF $count=1 $X=0.58
+ $Y=1.96 $X2=0.815 $Y2=2.865
.ends

.subckt PM_SKY130_FD_SC_HS__DLRBP_2%Q 1 2 9 13 17 18 19 20 23
c55 23 0 1.30305e-19 $X=6.96 $Y=1.295
c56 9 0 1.67826e-19 $X=6.315 $Y=0.515
r57 22 23 25.3036 $w=2.28e-07 $l=5.05e-07 $layer=LI1_cond $X=6.96 $Y=1.8
+ $X2=6.96 $Y2=1.295
r58 21 23 8.26753 $w=2.28e-07 $l=1.65e-07 $layer=LI1_cond $X=6.96 $Y=1.13
+ $X2=6.96 $Y2=1.295
r59 19 21 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=6.845 $Y=1.045
+ $X2=6.96 $Y2=1.13
r60 19 20 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=6.845 $Y=1.045
+ $X2=6.48 $Y2=1.045
r61 17 22 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=6.845 $Y=1.885
+ $X2=6.96 $Y2=1.8
r62 17 18 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=6.845 $Y=1.885
+ $X2=6.465 $Y2=1.885
r63 13 15 54.1497 $w=1.68e-07 $l=8.3e-07 $layer=LI1_cond $X=6.38 $Y=1.985
+ $X2=6.38 $Y2=2.815
r64 11 18 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.38 $Y=1.97
+ $X2=6.465 $Y2=1.885
r65 11 13 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=6.38 $Y=1.97
+ $X2=6.38 $Y2=1.985
r66 7 20 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=6.315 $Y=0.96
+ $X2=6.48 $Y2=1.045
r67 7 9 15.5405 $w=3.28e-07 $l=4.45e-07 $layer=LI1_cond $X=6.315 $Y=0.96
+ $X2=6.315 $Y2=0.515
r68 2 15 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=6.23
+ $Y=1.84 $X2=6.38 $Y2=2.815
r69 2 13 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=6.23
+ $Y=1.84 $X2=6.38 $Y2=1.985
r70 1 9 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=6.175
+ $Y=0.37 $X2=6.315 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__DLRBP_2%Q_N 1 2 9 13 14 19 25
c30 25 0 1.00299e-19 $X=8.405 $Y=1.82
r31 17 19 1.12043 $w=3.58e-07 $l=3.5e-08 $layer=LI1_cond $X=8.405 $Y=2 $X2=8.405
+ $Y2=2.035
r32 14 17 0.800308 $w=3.58e-07 $l=2.5e-08 $layer=LI1_cond $X=8.405 $Y=1.975
+ $X2=8.405 $Y2=2
r33 14 25 8.1909 $w=3.58e-07 $l=1.55e-07 $layer=LI1_cond $X=8.405 $Y=1.975
+ $X2=8.405 $Y2=1.82
r34 14 22 24.1693 $w=3.58e-07 $l=7.55e-07 $layer=LI1_cond $X=8.405 $Y=2.06
+ $X2=8.405 $Y2=2.815
r35 14 19 0.800308 $w=3.58e-07 $l=2.5e-08 $layer=LI1_cond $X=8.405 $Y=2.06
+ $X2=8.405 $Y2=2.035
r36 13 25 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=8.5 $Y=1.13 $X2=8.5
+ $Y2=1.82
r37 7 13 8.64139 $w=3.38e-07 $l=1.7e-07 $layer=LI1_cond $X=8.415 $Y=0.96
+ $X2=8.415 $Y2=1.13
r38 7 9 15.0834 $w=3.38e-07 $l=4.45e-07 $layer=LI1_cond $X=8.415 $Y=0.96
+ $X2=8.415 $Y2=0.515
r39 2 14 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=8.24
+ $Y=1.84 $X2=8.39 $Y2=1.985
r40 2 22 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=8.24
+ $Y=1.84 $X2=8.39 $Y2=2.815
r41 1 9 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=8.27
+ $Y=0.37 $X2=8.41 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__DLRBP_2%VGND 1 2 3 4 5 6 7 24 28 32 36 40 42 44 47
+ 54 55 57 58 60 61 62 64 91 95 101 104 108
r109 107 108 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=0
+ $X2=8.88 $Y2=0
r110 104 105 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=0
+ $X2=7.92 $Y2=0
r111 101 102 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0
+ $X2=0.72 $Y2=0
r112 99 108 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=0 $X2=8.88
+ $Y2=0
r113 99 105 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=0 $X2=7.92
+ $Y2=0
r114 98 99 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r115 96 104 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.075 $Y=0
+ $X2=7.91 $Y2=0
r116 96 98 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=8.075 $Y=0 $X2=8.4
+ $Y2=0
r117 95 107 4.01252 $w=1.7e-07 $l=1.82e-07 $layer=LI1_cond $X=8.755 $Y=0
+ $X2=8.937 $Y2=0
r118 95 98 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=8.755 $Y=0 $X2=8.4
+ $Y2=0
r119 94 105 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=0
+ $X2=7.92 $Y2=0
r120 93 94 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.44 $Y=0 $X2=7.44
+ $Y2=0
r121 91 104 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.745 $Y=0
+ $X2=7.91 $Y2=0
r122 91 93 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=7.745 $Y=0
+ $X2=7.44 $Y2=0
r123 90 94 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.48 $Y=0 $X2=7.44
+ $Y2=0
r124 89 90 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.48 $Y=0 $X2=6.48
+ $Y2=0
r125 87 90 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=6.48
+ $Y2=0
r126 86 87 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r127 83 86 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=4.56 $Y=0 $X2=5.52
+ $Y2=0
r128 80 81 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r129 78 81 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=2.64 $Y=0
+ $X2=4.08 $Y2=0
r130 77 80 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=2.64 $Y=0 $X2=4.08
+ $Y2=0
r131 77 78 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r132 75 78 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r133 74 75 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r134 72 75 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r135 72 102 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r136 71 74 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r137 71 72 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r138 69 101 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.955 $Y=0
+ $X2=0.79 $Y2=0
r139 69 71 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=0.955 $Y=0 $X2=1.2
+ $Y2=0
r140 67 102 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0
+ $X2=0.72 $Y2=0
r141 66 67 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r142 64 101 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.625 $Y=0
+ $X2=0.79 $Y2=0
r143 64 66 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=0.625 $Y=0
+ $X2=0.24 $Y2=0
r144 62 87 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=5.52
+ $Y2=0
r145 62 81 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=4.08
+ $Y2=0
r146 62 83 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r147 60 89 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=6.65 $Y=0 $X2=6.48
+ $Y2=0
r148 60 61 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.65 $Y=0 $X2=6.815
+ $Y2=0
r149 59 93 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=6.98 $Y=0 $X2=7.44
+ $Y2=0
r150 59 61 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.98 $Y=0 $X2=6.815
+ $Y2=0
r151 57 86 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=5.61 $Y=0 $X2=5.52
+ $Y2=0
r152 57 58 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.61 $Y=0 $X2=5.775
+ $Y2=0
r153 56 89 35.2299 $w=1.68e-07 $l=5.4e-07 $layer=LI1_cond $X=5.94 $Y=0 $X2=6.48
+ $Y2=0
r154 56 58 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.94 $Y=0 $X2=5.775
+ $Y2=0
r155 55 83 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.395 $Y=0 $X2=4.56
+ $Y2=0
r156 54 80 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=4.23 $Y=0 $X2=4.08
+ $Y2=0
r157 54 55 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.23 $Y=0 $X2=4.395
+ $Y2=0
r158 47 74 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=2.305 $Y=0
+ $X2=2.16 $Y2=0
r159 47 51 11.1804 $w=3.33e-07 $l=3.25e-07 $layer=LI1_cond $X=2.472 $Y=0
+ $X2=2.472 $Y2=0.325
r160 47 77 4.71304 $w=1.7e-07 $l=1.68e-07 $layer=LI1_cond $X=2.472 $Y=0 $X2=2.64
+ $Y2=0
r161 42 107 3.13065 $w=2.5e-07 $l=1.09864e-07 $layer=LI1_cond $X=8.88 $Y=0.085
+ $X2=8.937 $Y2=0
r162 42 44 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=8.88 $Y=0.085
+ $X2=8.88 $Y2=0.515
r163 38 104 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.91 $Y=0.085
+ $X2=7.91 $Y2=0
r164 38 40 18.5089 $w=3.28e-07 $l=5.3e-07 $layer=LI1_cond $X=7.91 $Y=0.085
+ $X2=7.91 $Y2=0.615
r165 34 61 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.815 $Y=0.085
+ $X2=6.815 $Y2=0
r166 34 36 18.3343 $w=3.28e-07 $l=5.25e-07 $layer=LI1_cond $X=6.815 $Y=0.085
+ $X2=6.815 $Y2=0.61
r167 30 58 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.775 $Y=0.085
+ $X2=5.775 $Y2=0
r168 30 32 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=5.775 $Y=0.085
+ $X2=5.775 $Y2=0.515
r169 26 55 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.395 $Y=0.085
+ $X2=4.395 $Y2=0
r170 26 28 26.0173 $w=3.28e-07 $l=7.45e-07 $layer=LI1_cond $X=4.395 $Y=0.085
+ $X2=4.395 $Y2=0.83
r171 22 101 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.79 $Y=0.085
+ $X2=0.79 $Y2=0
r172 22 24 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=0.79 $Y=0.085
+ $X2=0.79 $Y2=0.515
r173 7 44 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=8.7
+ $Y=0.37 $X2=8.84 $Y2=0.515
r174 6 40 91 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=2 $X=7.7
+ $Y=0.47 $X2=7.91 $Y2=0.615
r175 5 36 182 $w=1.7e-07 $l=3.28634e-07 $layer=licon1_NDIFF $count=1 $X=6.605
+ $Y=0.37 $X2=6.815 $Y2=0.61
r176 4 32 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=5.635
+ $Y=0.37 $X2=5.775 $Y2=0.515
r177 3 28 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=4.255
+ $Y=0.62 $X2=4.395 $Y2=0.83
r178 2 51 182 $w=1.7e-07 $l=2.59037e-07 $layer=licon1_NDIFF $count=1 $X=2.25
+ $Y=0.41 $X2=2.47 $Y2=0.325
r179 1 24 91 $w=1.7e-07 $l=2.41454e-07 $layer=licon1_NDIFF $count=2 $X=0.57
+ $Y=0.56 $X2=0.79 $Y2=0.515
.ends

