* NGSPICE file created from sky130_fd_sc_hs__dfxtp_1.ext - technology: sky130A

.subckt sky130_fd_sc_hs__dfxtp_1 CLK D VGND VNB VPB VPWR Q
M1000 Q a_1210_314# VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=3.304e+11p pd=2.83e+06u as=1.50923e+12p ps=1.272e+07u
M1001 a_454_503# D VPWR VPB pshort w=420000u l=150000u
+  ad=1.967e+11p pd=2.01e+06u as=0p ps=0u
M1002 a_1168_124# a_27_74# a_1011_424# VNB nlowvt w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=2.362e+11p ps=2.07e+06u
M1003 a_206_368# a_27_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.553e+11p pd=2.17e+06u as=1.27305e+12p ps=1.059e+07u
M1004 a_713_458# a_561_463# VGND VNB nlowvt w=550000u l=150000u
+  ad=2.18125e+11p pd=2.05e+06u as=0p ps=0u
M1005 VPWR a_1210_314# a_1118_508# VPB pshort w=420000u l=150000u
+  ad=0p pd=0u as=1.995e+11p ps=1.79e+06u
M1006 a_1011_424# a_206_368# a_713_458# VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_454_503# D VGND VNB nlowvt w=420000u l=150000u
+  ad=3.1125e+11p pd=2.43e+06u as=0p ps=0u
M1008 VPWR a_1011_424# a_1210_314# VPB pshort w=840000u l=150000u
+  ad=0p pd=0u as=2.478e+11p ps=2.27e+06u
M1009 VGND a_1011_424# a_1210_314# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=1.824e+11p ps=1.85e+06u
M1010 a_713_458# a_561_463# VPWR VPB pshort w=840000u l=150000u
+  ad=4.662e+11p pd=2.79e+06u as=0p ps=0u
M1011 a_1118_508# a_206_368# a_1011_424# VPB pshort w=420000u l=150000u
+  ad=0p pd=0u as=2.856e+11p ps=2.45e+06u
M1012 Q a_1210_314# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1013 VGND a_713_458# a_731_101# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=8.82e+10p ps=1.26e+06u
M1014 a_206_368# a_27_74# VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=3.304e+11p pd=2.83e+06u as=0p ps=0u
M1015 VPWR a_713_458# a_668_503# VPB pshort w=420000u l=150000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1016 VPWR CLK a_27_74# VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=3.304e+11p ps=2.83e+06u
M1017 a_731_101# a_206_368# a_561_463# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.575e+11p ps=1.73e+06u
M1018 a_1011_424# a_27_74# a_713_458# VPB pshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_561_463# a_27_74# a_454_503# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 VGND a_1210_314# a_1168_124# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 VGND CLK a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1022 a_668_503# a_27_74# a_561_463# VPB pshort w=420000u l=150000u
+  ad=0p pd=0u as=1.967e+11p ps=2.01e+06u
M1023 a_561_463# a_206_368# a_454_503# VPB pshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

