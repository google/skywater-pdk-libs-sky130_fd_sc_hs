* NGSPICE file created from sky130_fd_sc_hs__nand4b_4.ext - technology: sky130A

.subckt sky130_fd_sc_hs__nand4b_4 A_N B C D VGND VNB VPB VPWR Y
M1000 a_656_74# C a_1025_158# VNB nlowvt w=740000u l=150000u
+  ad=8.399e+11p pd=8.19e+06u as=1.0287e+12p ps=1.022e+07u
M1001 VGND D a_1025_158# VNB nlowvt w=740000u l=150000u
+  ad=6.9465e+11p pd=6.36e+06u as=0p ps=0u
M1002 Y B VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=2.2512e+12p pd=1.298e+07u as=5.0862e+12p ps=2.218e+07u
M1003 Y C VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_27_158# A_N VPWR VPB pshort w=840000u l=150000u
+  ad=2.52e+11p pd=2.28e+06u as=0p ps=0u
M1005 VPWR B Y VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VPWR A_N a_27_158# VPB pshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_225_74# B a_656_74# VNB nlowvt w=740000u l=150000u
+  ad=1.01295e+12p pd=1.022e+07u as=0p ps=0u
M1008 VPWR C Y VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_225_74# a_27_158# Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=4.144e+11p ps=4.08e+06u
M1010 a_1025_158# D VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_1025_158# C a_656_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_656_74# B a_225_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VPWR a_27_158# Y VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_225_74# a_27_158# Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 Y D VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_1025_158# C a_656_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_1025_158# D VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 VGND D a_1025_158# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 Y a_27_158# VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 VPWR D Y VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_225_74# B a_656_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_656_74# B a_225_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 VGND A_N a_27_158# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=1.962e+11p ps=2.05e+06u
M1024 Y a_27_158# a_225_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 Y a_27_158# a_225_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 a_656_74# C a_1025_158# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

