* File: sky130_fd_sc_hs__and2b_4.spice
* Created: Tue Sep  1 19:55:03 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hs__and2b_4.pex.spice"
.subckt sky130_fd_sc_hs__and2b_4  VNB VPB A_N B VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* B	B
* A_N	A_N
* VPB	VPB
* VNB	VNB
MM1011 N_VGND_M1011_d N_A_N_M1011_g N_A_27_392#_M1011_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.112 AS=0.1824 PD=0.99 PS=1.85 NRD=13.116 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75003.9 A=0.096 P=1.58 MULT=1
MM1007 N_A_233_74#_M1007_d N_B_M1007_g N_VGND_M1011_d VNB NLOWVT L=0.15 W=0.64
+ AD=0.112 AS=0.112 PD=0.99 PS=0.99 NRD=5.616 NRS=0 M=1 R=4.26667 SA=75000.7
+ SB=75003.4 A=0.096 P=1.58 MULT=1
MM1005 N_A_218_424#_M1005_d N_A_27_392#_M1005_g N_A_233_74#_M1007_d VNB NLOWVT
+ L=0.15 W=0.64 AD=0.0896 AS=0.112 PD=0.92 PS=0.99 NRD=0 NRS=7.488 M=1 R=4.26667
+ SA=75001.2 SB=75002.9 A=0.096 P=1.58 MULT=1
MM1015 N_A_218_424#_M1005_d N_A_27_392#_M1015_g N_A_233_74#_M1015_s VNB NLOWVT
+ L=0.15 W=0.64 AD=0.0896 AS=0.096 PD=0.92 PS=0.94 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75001.6 SB=75002.5 A=0.096 P=1.58 MULT=1
MM1017 N_A_233_74#_M1015_s N_B_M1017_g N_VGND_M1017_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.096 AS=0.111026 PD=0.94 PS=0.997101 NRD=3.744 NRS=9.372 M=1 R=4.26667
+ SA=75002.1 SB=75002 A=0.096 P=1.58 MULT=1
MM1000 N_VGND_M1017_s N_A_218_424#_M1000_g N_X_M1000_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.128374 AS=0.1073 PD=1.1529 PS=1.03 NRD=0.804 NRS=1.62 M=1 R=4.93333
+ SA=75002.3 SB=75001.5 A=0.111 P=1.78 MULT=1
MM1003 N_VGND_M1003_d N_A_218_424#_M1003_g N_X_M1000_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.11655 AS=0.1073 PD=1.055 PS=1.03 NRD=0 NRS=0 M=1 R=4.93333 SA=75002.7
+ SB=75001.1 A=0.111 P=1.78 MULT=1
MM1013 N_VGND_M1003_d N_A_218_424#_M1013_g N_X_M1013_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.11655 AS=0.1036 PD=1.055 PS=1.02 NRD=5.664 NRS=0 M=1 R=4.93333 SA=75003.2
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1014 N_VGND_M1014_d N_A_218_424#_M1014_g N_X_M1013_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.1036 PD=2.05 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75003.6
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1016 N_VPWR_M1016_d N_A_N_M1016_g N_A_27_392#_M1016_s VPB PSHORT L=0.15 W=1
+ AD=0.193261 AS=0.285 PD=1.48913 PS=2.57 NRD=1.9503 NRS=1.9503 M=1 R=6.66667
+ SA=75000.2 SB=75003.4 A=0.15 P=2.3 MULT=1
MM1001 N_A_218_424#_M1001_d N_A_27_392#_M1001_g N_VPWR_M1016_d VPB PSHORT L=0.15
+ W=0.84 AD=0.126 AS=0.162339 PD=1.14 PS=1.25087 NRD=2.3443 NRS=18.7544 M=1
+ R=5.6 SA=75000.7 SB=75003.5 A=0.126 P=1.98 MULT=1
MM1002 N_A_218_424#_M1001_d N_A_27_392#_M1002_g N_VPWR_M1002_s VPB PSHORT L=0.15
+ W=0.84 AD=0.126 AS=0.1554 PD=1.14 PS=1.21 NRD=2.3443 NRS=2.3443 M=1 R=5.6
+ SA=75001.2 SB=75003.1 A=0.126 P=1.98 MULT=1
MM1008 N_A_218_424#_M1008_d N_B_M1008_g N_VPWR_M1002_s VPB PSHORT L=0.15 W=0.84
+ AD=0.126 AS=0.1554 PD=1.14 PS=1.21 NRD=2.3443 NRS=18.7544 M=1 R=5.6 SA=75001.7
+ SB=75002.5 A=0.126 P=1.98 MULT=1
MM1010 N_A_218_424#_M1008_d N_B_M1010_g N_VPWR_M1010_s VPB PSHORT L=0.15 W=0.84
+ AD=0.126 AS=0.165 PD=1.14 PS=1.27714 NRD=2.3443 NRS=18.7544 M=1 R=5.6
+ SA=75002.1 SB=75002.1 A=0.126 P=1.98 MULT=1
MM1004 N_X_M1004_d N_A_218_424#_M1004_g N_VPWR_M1010_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.22 PD=1.42 PS=1.70286 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75002 SB=75001.6 A=0.168 P=2.54 MULT=1
MM1006 N_X_M1004_d N_A_218_424#_M1006_g N_VPWR_M1006_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75002.5 SB=75001.1 A=0.168 P=2.54 MULT=1
MM1009 N_X_M1009_d N_A_218_424#_M1009_g N_VPWR_M1006_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75002.9 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1012 N_X_M1009_d N_A_218_424#_M1012_g N_VPWR_M1012_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.3192 PD=1.42 PS=2.81 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75003.4 SB=75000.2 A=0.168 P=2.54 MULT=1
DX18_noxref VNB VPB NWDIODE A=9.6348 P=14.08
c_54 VNB 0 2.21145e-19 $X=0 $Y=0
c_108 VPB 0 1.47064e-19 $X=0 $Y=3.085
*
.include "sky130_fd_sc_hs__and2b_4.pxi.spice"
*
.ends
*
*
