* File: sky130_fd_sc_hs__dfrbp_1.pex.spice
* Created: Thu Aug 27 20:38:15 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HS__DFRBP_1%D 1 3 6 8 9 10 11 17 20 21
r31 20 22 45.79 $w=4.05e-07 $l=1.65e-07 $layer=POLY_cond $X=0.422 $Y=1.165
+ $X2=0.422 $Y2=1
r32 20 21 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=0.385
+ $Y=1.165 $X2=0.385 $Y2=1.165
r33 17 18 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=0.385
+ $Y=1.845 $X2=0.385 $Y2=1.845
r34 15 20 5.08091 $w=4.05e-07 $l=3.7e-08 $layer=POLY_cond $X=0.422 $Y=1.202
+ $X2=0.422 $Y2=1.165
r35 15 17 88.298 $w=4.05e-07 $l=6.43e-07 $layer=POLY_cond $X=0.422 $Y=1.202
+ $X2=0.422 $Y2=1.845
r36 11 18 5.5434 $w=3.93e-07 $l=1.9e-07 $layer=LI1_cond $X=0.322 $Y=2.035
+ $X2=0.322 $Y2=1.845
r37 10 18 5.25164 $w=3.93e-07 $l=1.8e-07 $layer=LI1_cond $X=0.322 $Y=1.665
+ $X2=0.322 $Y2=1.845
r38 9 10 10.795 $w=3.93e-07 $l=3.7e-07 $layer=LI1_cond $X=0.322 $Y=1.295
+ $X2=0.322 $Y2=1.665
r39 9 21 3.79285 $w=3.93e-07 $l=1.3e-07 $layer=LI1_cond $X=0.322 $Y=1.295
+ $X2=0.322 $Y2=1.165
r40 8 17 41.6085 $w=4.05e-07 $l=3.03e-07 $layer=POLY_cond $X=0.422 $Y=2.148
+ $X2=0.422 $Y2=1.845
r41 6 22 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=0.55 $Y=0.6 $X2=0.55
+ $Y2=1
r42 1 8 47.3046 $w=3.23e-07 $l=3.5609e-07 $layer=POLY_cond $X=0.505 $Y=2.465
+ $X2=0.422 $Y2=2.148
r43 1 3 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=0.505 $Y=2.465
+ $X2=0.505 $Y2=2.75
.ends

.subckt PM_SKY130_FD_SC_HS__DFRBP_1%RESET_B 3 6 8 9 11 14 16 17 19 22 24 26 27
+ 28 30 31 32 33 34 39 42 45 46 49 50 53 58
c191 50 0 7.11201e-21 $X=1.165 $Y=1.295
c192 49 0 1.15516e-19 $X=1.165 $Y=1.295
c193 39 0 6.85463e-20 $X=7.92 $Y=2.035
r194 57 58 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.135
+ $Y=2 $X2=8.135 $Y2=2
r195 53 55 41.4566 $w=4.65e-07 $l=1.65e-07 $layer=POLY_cond $X=1.097 $Y=1.975
+ $X2=1.097 $Y2=2.14
r196 53 54 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.165
+ $Y=1.975 $X2=1.165 $Y2=1.975
r197 50 54 29.0245 $w=2.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.165 $Y=1.295
+ $X2=1.165 $Y2=1.975
r198 49 51 47.3569 $w=4.65e-07 $l=1.65e-07 $layer=POLY_cond $X=1.097 $Y=1.295
+ $X2=1.097 $Y2=1.13
r199 49 50 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.165
+ $Y=1.295 $X2=1.165 $Y2=1.295
r200 45 46 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.395
+ $Y=1.99 $X2=5.395 $Y2=1.99
r201 42 54 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=2.035
+ $X2=1.2 $Y2=2.035
r202 40 58 7.50834 $w=3.28e-07 $l=2.15e-07 $layer=LI1_cond $X=7.92 $Y=2
+ $X2=8.135 $Y2=2
r203 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=2.035
+ $X2=7.92 $Y2=2.035
r204 36 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=2.035
+ $X2=5.52 $Y2=2.035
r205 34 36 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.665 $Y=2.035
+ $X2=5.52 $Y2=2.035
r206 33 39 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=7.775 $Y=2.035
+ $X2=7.92 $Y2=2.035
r207 33 34 2.61138 $w=1.4e-07 $l=2.11e-06 $layer=MET1_cond $X=7.775 $Y=2.035
+ $X2=5.665 $Y2=2.035
r208 32 42 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.345 $Y=2.035
+ $X2=1.2 $Y2=2.035
r209 31 36 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.375 $Y=2.035
+ $X2=5.52 $Y2=2.035
r210 31 32 4.98761 $w=1.4e-07 $l=4.03e-06 $layer=MET1_cond $X=5.375 $Y=2.035
+ $X2=1.345 $Y2=2.035
r211 29 45 65.573 $w=3.3e-07 $l=3.75e-07 $layer=POLY_cond $X=5.02 $Y=1.99
+ $X2=5.395 $Y2=1.99
r212 29 30 5.03009 $w=3.3e-07 $l=1.08995e-07 $layer=POLY_cond $X=5.02 $Y=1.99
+ $X2=4.93 $Y2=2.032
r213 27 28 49.7366 $w=2e-07 $l=1.5e-07 $layer=POLY_cond $X=4.89 $Y=1.085
+ $X2=4.89 $Y2=1.235
r214 24 57 57.6553 $w=2.91e-07 $l=3.01662e-07 $layer=POLY_cond $X=8.18 $Y=2.28
+ $X2=8.135 $Y2=2
r215 24 26 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=8.18 $Y=2.28
+ $X2=8.18 $Y2=2.565
r216 20 57 38.6072 $w=2.91e-07 $l=2.05122e-07 $layer=POLY_cond $X=8.045 $Y=1.835
+ $X2=8.135 $Y2=2
r217 20 22 643.521 $w=1.5e-07 $l=1.255e-06 $layer=POLY_cond $X=8.045 $Y=1.835
+ $X2=8.045 $Y2=0.58
r218 17 30 37.0704 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=4.93 $Y=2.24
+ $X2=4.93 $Y2=2.032
r219 17 19 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=4.93 $Y=2.24
+ $X2=4.93 $Y2=2.525
r220 16 30 37.0704 $w=1.5e-07 $l=2.14369e-07 $layer=POLY_cond $X=4.915 $Y=1.825
+ $X2=4.93 $Y2=2.032
r221 16 28 302.532 $w=1.5e-07 $l=5.9e-07 $layer=POLY_cond $X=4.915 $Y=1.825
+ $X2=4.915 $Y2=1.235
r222 14 27 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=4.865 $Y=0.8
+ $X2=4.865 $Y2=1.085
r223 9 11 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=0.955 $Y=2.465
+ $X2=0.955 $Y2=2.75
r224 8 9 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=0.955 $Y=2.375
+ $X2=0.955 $Y2=2.465
r225 8 55 91.3468 $w=1.8e-07 $l=2.35e-07 $layer=POLY_cond $X=0.955 $Y=2.375
+ $X2=0.955 $Y2=2.14
r226 6 53 8.0134 $w=4.65e-07 $l=6.7e-08 $layer=POLY_cond $X=1.097 $Y=1.908
+ $X2=1.097 $Y2=1.975
r227 5 49 8.0134 $w=4.65e-07 $l=6.7e-08 $layer=POLY_cond $X=1.097 $Y=1.362
+ $X2=1.097 $Y2=1.295
r228 5 6 65.3032 $w=4.65e-07 $l=5.46e-07 $layer=POLY_cond $X=1.097 $Y=1.362
+ $X2=1.097 $Y2=1.908
r229 3 51 271.766 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=0.94 $Y=0.6 $X2=0.94
+ $Y2=1.13
.ends

.subckt PM_SKY130_FD_SC_HS__DFRBP_1%CLK 1 3 6 8
c43 6 0 7.11201e-21 $X=1.97 $Y=0.74
c44 1 0 1.84834e-19 $X=1.965 $Y=1.725
r45 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.95
+ $Y=1.475 $X2=1.95 $Y2=1.475
r46 8 12 6.42105 $w=3.99e-07 $l=2.1e-07 $layer=LI1_cond $X=2.16 $Y=1.545
+ $X2=1.95 $Y2=1.545
r47 4 11 38.5562 $w=2.99e-07 $l=1.74714e-07 $layer=POLY_cond $X=1.97 $Y=1.31
+ $X2=1.95 $Y2=1.475
r48 4 6 292.277 $w=1.5e-07 $l=5.7e-07 $layer=POLY_cond $X=1.97 $Y=1.31 $X2=1.97
+ $Y2=0.74
r49 1 11 52.2586 $w=2.99e-07 $l=2.57391e-07 $layer=POLY_cond $X=1.965 $Y=1.725
+ $X2=1.95 $Y2=1.475
r50 1 3 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.965 $Y=1.725
+ $X2=1.965 $Y2=2.36
.ends

.subckt PM_SKY130_FD_SC_HS__DFRBP_1%A_498_360# 1 2 8 9 11 12 15 16 18 19 21 22
+ 23 24 26 29 32 33 35 37 41 42 43 45 46 47 50 52 53 55 61 66
c198 66 0 1.69357e-19 $X=3.385 $Y=1.65
c199 52 0 1.08581e-19 $X=6.735 $Y=1.865
c200 47 0 1.02732e-19 $X=6.255 $Y=1.065
c201 43 0 1.03779e-19 $X=4.52 $Y=0.665
c202 9 0 1.6736e-20 $X=3.455 $Y=2.24
r203 64 65 11.0397 $w=5.23e-07 $l=2.25e-07 $layer=LI1_cond $X=2.852 $Y=0.575
+ $X2=2.852 $Y2=0.8
r204 61 64 5.35387 $w=5.23e-07 $l=2.35e-07 $layer=LI1_cond $X=2.852 $Y=0.34
+ $X2=2.852 $Y2=0.575
r205 59 60 14.2883 $w=3.33e-07 $l=3.9e-07 $layer=LI1_cond $X=2.64 $Y=1.857
+ $X2=3.03 $Y2=1.857
r206 55 56 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.205
+ $Y=2.03 $X2=7.205 $Y2=2.03
r207 53 55 13.4452 $w=3.28e-07 $l=3.85e-07 $layer=LI1_cond $X=6.82 $Y=2.03
+ $X2=7.205 $Y2=2.03
r208 52 53 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=6.735 $Y=1.865
+ $X2=6.82 $Y2=2.03
r209 51 52 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=6.735 $Y=1.23
+ $X2=6.735 $Y2=1.865
r210 50 72 16.6118 $w=3.3e-07 $l=9.5e-08 $layer=POLY_cond $X=6.645 $Y=1.065
+ $X2=6.645 $Y2=1.16
r211 49 50 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.645
+ $Y=1.065 $X2=6.645 $Y2=1.065
r212 47 49 13.6198 $w=3.28e-07 $l=3.9e-07 $layer=LI1_cond $X=6.255 $Y=1.065
+ $X2=6.645 $Y2=1.065
r213 46 51 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=6.65 $Y=1.065
+ $X2=6.735 $Y2=1.23
r214 46 49 0.174613 $w=3.28e-07 $l=5e-09 $layer=LI1_cond $X=6.65 $Y=1.065
+ $X2=6.645 $Y2=1.065
r215 45 47 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=6.17 $Y=0.9
+ $X2=6.255 $Y2=1.065
r216 44 45 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=6.17 $Y=0.75
+ $X2=6.17 $Y2=0.9
r217 42 44 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.085 $Y=0.665
+ $X2=6.17 $Y2=0.75
r218 42 43 102.102 $w=1.68e-07 $l=1.565e-06 $layer=LI1_cond $X=6.085 $Y=0.665
+ $X2=4.52 $Y2=0.665
r219 41 43 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.435 $Y=0.58
+ $X2=4.52 $Y2=0.665
r220 40 41 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=4.435 $Y=0.425
+ $X2=4.435 $Y2=0.58
r221 38 69 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.385 $Y=1.74
+ $X2=3.385 $Y2=1.905
r222 38 66 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=3.385 $Y=1.74
+ $X2=3.385 $Y2=1.65
r223 37 38 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.385
+ $Y=1.74 $X2=3.385 $Y2=1.74
r224 35 60 3.11411 $w=3.33e-07 $l=1.53734e-07 $layer=LI1_cond $X=3.115 $Y=1.74
+ $X2=3.03 $Y2=1.857
r225 35 37 9.42908 $w=3.28e-07 $l=2.7e-07 $layer=LI1_cond $X=3.115 $Y=1.74
+ $X2=3.385 $Y2=1.74
r226 34 61 7.46409 $w=1.7e-07 $l=2.63e-07 $layer=LI1_cond $X=3.115 $Y=0.34
+ $X2=2.852 $Y2=0.34
r227 33 40 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.35 $Y=0.34
+ $X2=4.435 $Y2=0.425
r228 33 34 80.5722 $w=1.68e-07 $l=1.235e-06 $layer=LI1_cond $X=4.35 $Y=0.34
+ $X2=3.115 $Y2=0.34
r229 32 60 4.67747 $w=1.7e-07 $l=2.82e-07 $layer=LI1_cond $X=3.03 $Y=1.575
+ $X2=3.03 $Y2=1.857
r230 32 65 50.5615 $w=1.68e-07 $l=7.75e-07 $layer=LI1_cond $X=3.03 $Y=1.575
+ $X2=3.03 $Y2=0.8
r231 27 29 56.4043 $w=1.5e-07 $l=1.1e-07 $layer=POLY_cond $X=3.975 $Y=1.17
+ $X2=4.085 $Y2=1.17
r232 24 56 52.2586 $w=2.99e-07 $l=2.7157e-07 $layer=POLY_cond $X=7.25 $Y=2.28
+ $X2=7.205 $Y2=2.03
r233 24 26 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=7.25 $Y=2.28
+ $X2=7.25 $Y2=2.565
r234 22 72 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.48 $Y=1.16
+ $X2=6.645 $Y2=1.16
r235 22 23 184.596 $w=1.5e-07 $l=3.6e-07 $layer=POLY_cond $X=6.48 $Y=1.16
+ $X2=6.12 $Y2=1.16
r236 19 23 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=6.045 $Y=1.085
+ $X2=6.12 $Y2=1.16
r237 19 21 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=6.045 $Y=1.085
+ $X2=6.045 $Y2=0.69
r238 16 29 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.085 $Y=1.095
+ $X2=4.085 $Y2=1.17
r239 16 18 94.7933 $w=1.5e-07 $l=2.95e-07 $layer=POLY_cond $X=4.085 $Y=1.095
+ $X2=4.085 $Y2=0.8
r240 14 27 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.975 $Y=1.245
+ $X2=3.975 $Y2=1.17
r241 14 15 169.213 $w=1.5e-07 $l=3.3e-07 $layer=POLY_cond $X=3.975 $Y=1.245
+ $X2=3.975 $Y2=1.575
r242 13 66 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.55 $Y=1.65
+ $X2=3.385 $Y2=1.65
r243 12 15 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.9 $Y=1.65
+ $X2=3.975 $Y2=1.575
r244 12 13 179.468 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=3.9 $Y=1.65
+ $X2=3.55 $Y2=1.65
r245 9 11 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=3.455 $Y=2.24
+ $X2=3.455 $Y2=2.525
r246 8 9 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=3.455 $Y=2.15 $X2=3.455
+ $Y2=2.24
r247 8 69 95.2339 $w=1.8e-07 $l=2.45e-07 $layer=POLY_cond $X=3.455 $Y=2.15
+ $X2=3.455 $Y2=1.905
r248 2 59 600 $w=1.7e-07 $l=2.22711e-07 $layer=licon1_PDIFF $count=1 $X=2.49
+ $Y=1.8 $X2=2.64 $Y2=1.96
r249 1 64 182 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_NDIFF $count=1 $X=2.615
+ $Y=0.37 $X2=2.755 $Y2=0.575
.ends

.subckt PM_SKY130_FD_SC_HS__DFRBP_1%A_841_401# 1 2 7 9 12 14 19 20 22 23 24 25
+ 26 27 30
c113 23 0 1.58258e-20 $X=4.63 $Y=1.005
c114 12 0 1.63224e-19 $X=4.475 $Y=0.8
r115 30 32 32.7294 $w=2.48e-07 $l=7.1e-07 $layer=LI1_cond $X=6.355 $Y=1.88
+ $X2=6.355 $Y2=2.59
r116 28 30 14.2903 $w=2.48e-07 $l=3.1e-07 $layer=LI1_cond $X=6.355 $Y=1.57
+ $X2=6.355 $Y2=1.88
r117 26 28 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=6.23 $Y=1.485
+ $X2=6.355 $Y2=1.57
r118 26 27 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=6.23 $Y=1.485
+ $X2=5.915 $Y2=1.485
r119 25 27 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.83 $Y=1.4
+ $X2=5.915 $Y2=1.485
r120 24 35 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.83 $Y=1.09
+ $X2=5.83 $Y2=1.005
r121 24 25 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=5.83 $Y=1.09
+ $X2=5.83 $Y2=1.4
r122 22 35 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.745 $Y=1.005
+ $X2=5.83 $Y2=1.005
r123 22 23 72.7433 $w=1.68e-07 $l=1.115e-06 $layer=LI1_cond $X=5.745 $Y=1.005
+ $X2=4.63 $Y2=1.005
r124 19 20 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.465
+ $Y=1.65 $X2=4.465 $Y2=1.65
r125 17 23 7.36005 $w=1.7e-07 $l=1.77482e-07 $layer=LI1_cond $X=4.49 $Y=1.09
+ $X2=4.63 $Y2=1.005
r126 17 19 23.0489 $w=2.78e-07 $l=5.6e-07 $layer=LI1_cond $X=4.49 $Y=1.09
+ $X2=4.49 $Y2=1.65
r127 16 20 38.0424 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.465 $Y=1.485
+ $X2=4.465 $Y2=1.65
r128 14 20 62.0758 $w=3.3e-07 $l=3.55e-07 $layer=POLY_cond $X=4.465 $Y=2.005
+ $X2=4.465 $Y2=1.65
r129 12 16 351.245 $w=1.5e-07 $l=6.85e-07 $layer=POLY_cond $X=4.475 $Y=0.8
+ $X2=4.475 $Y2=1.485
r130 7 14 33.7113 $w=3.36e-07 $l=3.08504e-07 $layer=POLY_cond $X=4.295 $Y=2.24
+ $X2=4.465 $Y2=2.005
r131 7 9 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=4.295 $Y=2.24
+ $X2=4.295 $Y2=2.525
r132 2 32 400 $w=1.7e-07 $l=9.26971e-07 $layer=licon1_PDIFF $count=1 $X=6.165
+ $Y=1.735 $X2=6.315 $Y2=2.59
r133 2 30 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=6.165
+ $Y=1.735 $X2=6.315 $Y2=1.88
r134 1 35 182 $w=1.7e-07 $l=7.36834e-07 $layer=licon1_NDIFF $count=1 $X=5.53
+ $Y=0.37 $X2=5.75 $Y2=1.005
.ends

.subckt PM_SKY130_FD_SC_HS__DFRBP_1%A_706_463# 1 2 3 12 14 16 18 20 21 22 24 31
+ 33 36 37
c129 33 0 1.55214e-19 $X=4.975 $Y=1.45
c130 31 0 1.21504e-19 $X=4.095 $Y=0.812
c131 20 0 1.03565e-19 $X=4.095 $Y=2.415
c132 14 0 2.11313e-19 $X=6 $Y=1.54
r133 37 39 7.32792 $w=3.08e-07 $l=1.85e-07 $layer=LI1_cond $X=4.975 $Y=2.515
+ $X2=5.16 $Y2=2.515
r134 36 42 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=5.395 $Y=1.45
+ $X2=5.395 $Y2=1.54
r135 36 41 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.395 $Y=1.45
+ $X2=5.395 $Y2=1.285
r136 35 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.395
+ $Y=1.45 $X2=5.395 $Y2=1.45
r137 33 35 20.6613 $w=2.48e-07 $l=4.2e-07 $layer=LI1_cond $X=4.975 $Y=1.45
+ $X2=5.395 $Y2=1.45
r138 29 31 5.96091 $w=4.33e-07 $l=2.25e-07 $layer=LI1_cond $X=3.87 $Y=0.812
+ $X2=4.095 $Y2=0.812
r139 26 27 20.9215 $w=2.42e-07 $l=4.15e-07 $layer=LI1_cond $X=3.68 $Y=2.585
+ $X2=4.095 $Y2=2.585
r140 24 37 4.21588 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.975 $Y=2.35
+ $X2=4.975 $Y2=2.515
r141 23 33 2.94836 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.975 $Y=1.615
+ $X2=4.975 $Y2=1.45
r142 23 24 47.9519 $w=1.68e-07 $l=7.35e-07 $layer=LI1_cond $X=4.975 $Y=1.615
+ $X2=4.975 $Y2=2.35
r143 22 27 5.3796 $w=2.42e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.18 $Y=2.5
+ $X2=4.095 $Y2=2.585
r144 21 37 5.79756 $w=3.08e-07 $l=9.21954e-08 $layer=LI1_cond $X=4.89 $Y=2.5
+ $X2=4.975 $Y2=2.515
r145 21 22 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=4.89 $Y=2.5
+ $X2=4.18 $Y2=2.5
r146 20 27 2.80567 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=4.095 $Y=2.415
+ $X2=4.095 $Y2=2.585
r147 19 31 6.29128 $w=1.7e-07 $l=2.18e-07 $layer=LI1_cond $X=4.095 $Y=1.03
+ $X2=4.095 $Y2=0.812
r148 19 20 90.3583 $w=1.68e-07 $l=1.385e-06 $layer=LI1_cond $X=4.095 $Y=1.03
+ $X2=4.095 $Y2=2.415
r149 16 18 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=6.09 $Y=1.66
+ $X2=6.09 $Y2=2.235
r150 15 42 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.56 $Y=1.54
+ $X2=5.395 $Y2=1.54
r151 14 16 26.9307 $w=1.5e-07 $l=1.58745e-07 $layer=POLY_cond $X=6 $Y=1.54
+ $X2=6.09 $Y2=1.66
r152 14 15 225.617 $w=1.5e-07 $l=4.4e-07 $layer=POLY_cond $X=6 $Y=1.54 $X2=5.56
+ $Y2=1.54
r153 12 41 305.096 $w=1.5e-07 $l=5.95e-07 $layer=POLY_cond $X=5.455 $Y=0.69
+ $X2=5.455 $Y2=1.285
r154 3 39 600 $w=1.7e-07 $l=2.66458e-07 $layer=licon1_PDIFF $count=1 $X=5.005
+ $Y=2.315 $X2=5.16 $Y2=2.515
r155 2 26 600 $w=1.7e-07 $l=3.36749e-07 $layer=licon1_PDIFF $count=1 $X=3.53
+ $Y=2.315 $X2=3.68 $Y2=2.585
r156 1 29 182 $w=1.7e-07 $l=3.07571e-07 $layer=licon1_NDIFF $count=1 $X=3.66
+ $Y=0.59 $X2=3.87 $Y2=0.81
.ends

.subckt PM_SKY130_FD_SC_HS__DFRBP_1%A_319_360# 1 2 7 9 10 12 14 15 16 17 18 21
+ 23 24 25 27 28 30 31 35 36 37 40 42 45 48 49 53 56 60
c190 56 0 1.15516e-19 $X=1.695 $Y=1.055
c191 53 0 1.84834e-19 $X=2.61 $Y=1.385
c192 21 0 1.58258e-20 $X=3.585 $Y=0.8
c193 15 0 1.03565e-19 $X=3.51 $Y=1.26
c194 14 0 5.32615e-20 $X=2.935 $Y=3.075
r195 62 63 14.6951 $w=4.1e-07 $l=1.25e-07 $layer=POLY_cond $X=2.415 $Y=1.455
+ $X2=2.54 $Y2=1.455
r196 57 60 6.46067 $w=3.28e-07 $l=1.85e-07 $layer=LI1_cond $X=1.555 $Y=1.975
+ $X2=1.74 $Y2=1.975
r197 54 63 8.22927 $w=4.1e-07 $l=7e-08 $layer=POLY_cond $X=2.61 $Y=1.455
+ $X2=2.54 $Y2=1.455
r198 53 54 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.61
+ $Y=1.385 $X2=2.61 $Y2=1.385
r199 51 53 8.55602 $w=3.28e-07 $l=2.45e-07 $layer=LI1_cond $X=2.61 $Y=1.14
+ $X2=2.61 $Y2=1.385
r200 50 56 3.57226 $w=1.7e-07 $l=2.25e-07 $layer=LI1_cond $X=1.92 $Y=1.055
+ $X2=1.695 $Y2=1.055
r201 49 51 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.445 $Y=1.055
+ $X2=2.61 $Y2=1.14
r202 49 50 34.2513 $w=1.68e-07 $l=5.25e-07 $layer=LI1_cond $X=2.445 $Y=1.055
+ $X2=1.92 $Y2=1.055
r203 48 57 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.555 $Y=1.81
+ $X2=1.555 $Y2=1.975
r204 47 56 3.05675 $w=3.1e-07 $l=1.77482e-07 $layer=LI1_cond $X=1.555 $Y=1.14
+ $X2=1.695 $Y2=1.055
r205 47 48 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.555 $Y=1.14
+ $X2=1.555 $Y2=1.81
r206 43 56 3.05675 $w=3.1e-07 $l=8.5e-08 $layer=LI1_cond $X=1.695 $Y=0.97
+ $X2=1.695 $Y2=1.055
r207 43 45 12.0937 $w=4.48e-07 $l=4.55e-07 $layer=LI1_cond $X=1.695 $Y=0.97
+ $X2=1.695 $Y2=0.515
r208 38 40 458.926 $w=1.5e-07 $l=8.95e-07 $layer=POLY_cond $X=7.095 $Y=1.475
+ $X2=7.095 $Y2=0.58
r209 36 38 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=7.02 $Y=1.55
+ $X2=7.095 $Y2=1.475
r210 36 37 199.979 $w=1.5e-07 $l=3.9e-07 $layer=POLY_cond $X=7.02 $Y=1.55
+ $X2=6.63 $Y2=1.55
r211 33 35 294.84 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=6.54 $Y=2.81
+ $X2=6.54 $Y2=2.235
r212 32 37 26.9307 $w=1.5e-07 $l=1.48324e-07 $layer=POLY_cond $X=6.54 $Y=1.66
+ $X2=6.63 $Y2=1.55
r213 32 35 294.84 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=6.54 $Y=1.66
+ $X2=6.54 $Y2=2.235
r214 30 33 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=6.54 $Y=2.9 $X2=6.54
+ $Y2=2.81
r215 30 31 68.0242 $w=1.8e-07 $l=1.75e-07 $layer=POLY_cond $X=6.54 $Y=2.9
+ $X2=6.54 $Y2=3.075
r216 29 42 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=3.995 $Y=3.15
+ $X2=3.905 $Y2=3.15
r217 28 31 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=6.45 $Y=3.15
+ $X2=6.54 $Y2=3.075
r218 28 29 1258.84 $w=1.5e-07 $l=2.455e-06 $layer=POLY_cond $X=6.45 $Y=3.15
+ $X2=3.995 $Y2=3.15
r219 25 27 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=3.905 $Y=2.81
+ $X2=3.905 $Y2=2.525
r220 24 42 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=3.905 $Y=3.075
+ $X2=3.905 $Y2=3.15
r221 23 25 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=3.905 $Y=2.9
+ $X2=3.905 $Y2=2.81
r222 23 24 68.0242 $w=1.8e-07 $l=1.75e-07 $layer=POLY_cond $X=3.905 $Y=2.9
+ $X2=3.905 $Y2=3.075
r223 19 21 197.415 $w=1.5e-07 $l=3.85e-07 $layer=POLY_cond $X=3.585 $Y=1.185
+ $X2=3.585 $Y2=0.8
r224 17 42 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=3.815 $Y=3.15
+ $X2=3.905 $Y2=3.15
r225 17 18 412.777 $w=1.5e-07 $l=8.05e-07 $layer=POLY_cond $X=3.815 $Y=3.15
+ $X2=3.01 $Y2=3.15
r226 15 19 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.51 $Y=1.26
+ $X2=3.585 $Y2=1.185
r227 15 16 256.383 $w=1.5e-07 $l=5e-07 $layer=POLY_cond $X=3.51 $Y=1.26 $X2=3.01
+ $Y2=1.26
r228 14 18 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.935 $Y=3.075
+ $X2=3.01 $Y2=3.15
r229 13 16 29.2062 $w=4.1e-07 $l=2.29456e-07 $layer=POLY_cond $X=2.935 $Y=1.455
+ $X2=3.01 $Y2=1.26
r230 13 54 38.2073 $w=4.1e-07 $l=3.25e-07 $layer=POLY_cond $X=2.935 $Y=1.455
+ $X2=2.61 $Y2=1.455
r231 13 14 781.968 $w=1.5e-07 $l=1.525e-06 $layer=POLY_cond $X=2.935 $Y=1.55
+ $X2=2.935 $Y2=3.075
r232 10 63 26.4667 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=2.54 $Y=1.185
+ $X2=2.54 $Y2=1.455
r233 10 12 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=2.54 $Y=1.185
+ $X2=2.54 $Y2=0.74
r234 7 62 26.4667 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=2.415 $Y=1.725
+ $X2=2.415 $Y2=1.455
r235 7 9 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.415 $Y=1.725
+ $X2=2.415 $Y2=2.36
r236 2 60 600 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=1.595
+ $Y=1.8 $X2=1.74 $Y2=1.975
r237 1 45 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=1.61
+ $Y=0.37 $X2=1.755 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__DFRBP_1%A_1482_48# 1 2 7 9 11 12 14 15 18 21 24 25
+ 38 40 44
c95 38 0 6.85463e-20 $X=8.885 $Y=1.85
c96 15 0 1.98491e-19 $X=8.485 $Y=0.985
r97 36 38 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=8.555 $Y=1.85
+ $X2=8.885 $Y2=1.85
r98 29 44 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=7.595 $Y=1.065
+ $X2=7.67 $Y2=1.065
r99 29 41 19.2347 $w=3.3e-07 $l=1.1e-07 $layer=POLY_cond $X=7.595 $Y=1.065
+ $X2=7.485 $Y2=1.065
r100 28 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.595
+ $Y=1.065 $X2=7.595 $Y2=1.065
r101 25 28 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=7.595 $Y=0.985
+ $X2=7.595 $Y2=1.065
r102 24 38 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.885 $Y=1.765
+ $X2=8.885 $Y2=1.85
r103 23 40 2.90768 $w=3.27e-07 $l=1.95944e-07 $layer=LI1_cond $X=8.885 $Y=1.07
+ $X2=8.727 $Y2=0.985
r104 23 24 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=8.885 $Y=1.07
+ $X2=8.885 $Y2=1.765
r105 19 40 2.90768 $w=3.27e-07 $l=8.5e-08 $layer=LI1_cond $X=8.727 $Y=0.9
+ $X2=8.727 $Y2=0.985
r106 19 21 7.89165 $w=4.83e-07 $l=3.2e-07 $layer=LI1_cond $X=8.727 $Y=0.9
+ $X2=8.727 $Y2=0.58
r107 18 32 4.37637 $w=3.93e-07 $l=1.5e-07 $layer=LI1_cond $X=8.555 $Y=2.532
+ $X2=8.405 $Y2=2.532
r108 17 36 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.555 $Y=1.935
+ $X2=8.555 $Y2=1.85
r109 17 18 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=8.555 $Y=1.935
+ $X2=8.555 $Y2=2.335
r110 16 25 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.76 $Y=0.985
+ $X2=7.595 $Y2=0.985
r111 15 40 3.78066 $w=1.7e-07 $l=2.42e-07 $layer=LI1_cond $X=8.485 $Y=0.985
+ $X2=8.727 $Y2=0.985
r112 15 16 47.2995 $w=1.68e-07 $l=7.25e-07 $layer=LI1_cond $X=8.485 $Y=0.985
+ $X2=7.76 $Y2=0.985
r113 12 14 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=7.67 $Y=2.28
+ $X2=7.67 $Y2=2.565
r114 11 12 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=7.67 $Y=2.19 $X2=7.67
+ $Y2=2.28
r115 10 44 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=7.67 $Y=1.23
+ $X2=7.67 $Y2=1.065
r116 10 11 373.161 $w=1.8e-07 $l=9.6e-07 $layer=POLY_cond $X=7.67 $Y=1.23
+ $X2=7.67 $Y2=2.19
r117 7 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.485 $Y=0.9
+ $X2=7.485 $Y2=1.065
r118 7 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=7.485 $Y=0.9
+ $X2=7.485 $Y2=0.58
r119 2 32 600 $w=1.7e-07 $l=2.74955e-07 $layer=licon1_PDIFF $count=1 $X=8.255
+ $Y=2.355 $X2=8.405 $Y2=2.565
r120 1 21 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=8.51
+ $Y=0.37 $X2=8.65 $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_HS__DFRBP_1%A_1224_74# 1 2 9 12 13 15 16 17 18 20 23 25
+ 28 29 31 34 37 38 42 47 48 49 51 52 54 56
c164 51 0 1.04385e-19 $X=7.58 $Y=2.365
c165 29 0 1.79977e-19 $X=10.5 $Y=2.045
c166 17 0 1.98491e-19 $X=8.72 $Y=1.43
r167 57 64 23.6063 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=8.495 $Y=1.43
+ $X2=8.63 $Y2=1.43
r168 57 61 10.4917 $w=3.3e-07 $l=6e-08 $layer=POLY_cond $X=8.495 $Y=1.43
+ $X2=8.435 $Y2=1.43
r169 56 59 3.07318 $w=2.98e-07 $l=8e-08 $layer=LI1_cond $X=8.48 $Y=1.43 $X2=8.48
+ $Y2=1.51
r170 56 57 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.495
+ $Y=1.43 $X2=8.495 $Y2=1.43
r171 53 54 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.665 $Y=1.51
+ $X2=7.58 $Y2=1.51
r172 52 59 4.061 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=8.33 $Y=1.51 $X2=8.48
+ $Y2=1.51
r173 52 53 43.385 $w=1.68e-07 $l=6.65e-07 $layer=LI1_cond $X=8.33 $Y=1.51
+ $X2=7.665 $Y2=1.51
r174 50 54 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.58 $Y=1.595
+ $X2=7.58 $Y2=1.51
r175 50 51 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=7.58 $Y=1.595
+ $X2=7.58 $Y2=2.365
r176 48 54 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.495 $Y=1.51
+ $X2=7.58 $Y2=1.51
r177 48 49 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=7.495 $Y=1.51
+ $X2=7.16 $Y2=1.51
r178 47 49 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.075 $Y=1.425
+ $X2=7.16 $Y2=1.51
r179 46 47 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=7.075 $Y=0.73
+ $X2=7.075 $Y2=1.425
r180 42 51 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=7.495 $Y=2.53
+ $X2=7.58 $Y2=2.365
r181 42 44 21.1281 $w=3.28e-07 $l=6.05e-07 $layer=LI1_cond $X=7.495 $Y=2.53
+ $X2=6.89 $Y2=2.53
r182 38 46 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=6.99 $Y=0.565
+ $X2=7.075 $Y2=0.73
r183 38 40 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=6.99 $Y=0.565
+ $X2=6.695 $Y2=0.565
r184 32 37 34.7346 $w=1.65e-07 $l=1.72337e-07 $layer=POLY_cond $X=10.515
+ $Y=1.265 $X2=10.5 $Y2=1.43
r185 32 34 317.915 $w=1.5e-07 $l=6.2e-07 $layer=POLY_cond $X=10.515 $Y=1.265
+ $X2=10.515 $Y2=0.645
r186 29 31 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=10.5 $Y=2.045
+ $X2=10.5 $Y2=2.54
r187 28 29 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=10.5 $Y=1.955
+ $X2=10.5 $Y2=2.045
r188 27 37 34.7346 $w=1.65e-07 $l=1.65e-07 $layer=POLY_cond $X=10.5 $Y=1.595
+ $X2=10.5 $Y2=1.43
r189 27 28 139.935 $w=1.8e-07 $l=3.6e-07 $layer=POLY_cond $X=10.5 $Y=1.595
+ $X2=10.5 $Y2=1.955
r190 26 36 5.16599 $w=3.3e-07 $l=2.3e-07 $layer=POLY_cond $X=9.515 $Y=1.43
+ $X2=9.285 $Y2=1.43
r191 25 37 3.90195 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=10.41 $Y=1.43
+ $X2=10.5 $Y2=1.43
r192 25 26 156.501 $w=3.3e-07 $l=8.95e-07 $layer=POLY_cond $X=10.41 $Y=1.43
+ $X2=9.515 $Y2=1.43
r193 21 36 38.9663 $w=3.64e-07 $l=2.29783e-07 $layer=POLY_cond $X=9.44 $Y=1.265
+ $X2=9.285 $Y2=1.43
r194 21 23 269.202 $w=1.5e-07 $l=5.25e-07 $layer=POLY_cond $X=9.44 $Y=1.265
+ $X2=9.44 $Y2=0.74
r195 18 36 61.4773 $w=3.64e-07 $l=3.98905e-07 $layer=POLY_cond $X=9.145 $Y=1.765
+ $X2=9.285 $Y2=1.43
r196 18 20 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=9.145 $Y=1.765
+ $X2=9.145 $Y2=2.4
r197 17 64 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=8.72 $Y=1.43 $X2=8.63
+ $Y2=1.43
r198 16 36 5.16599 $w=3.3e-07 $l=2.3e-07 $layer=POLY_cond $X=9.055 $Y=1.43
+ $X2=9.285 $Y2=1.43
r199 16 17 58.5785 $w=3.3e-07 $l=3.35e-07 $layer=POLY_cond $X=9.055 $Y=1.43
+ $X2=8.72 $Y2=1.43
r200 13 15 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=8.63 $Y=2.28
+ $X2=8.63 $Y2=2.565
r201 12 13 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=8.63 $Y=2.19 $X2=8.63
+ $Y2=2.28
r202 11 64 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=8.63 $Y=1.595
+ $X2=8.63 $Y2=1.43
r203 11 12 231.282 $w=1.8e-07 $l=5.95e-07 $layer=POLY_cond $X=8.63 $Y=1.595
+ $X2=8.63 $Y2=2.19
r204 7 61 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.435 $Y=1.265
+ $X2=8.435 $Y2=1.43
r205 7 9 351.245 $w=1.5e-07 $l=6.85e-07 $layer=POLY_cond $X=8.435 $Y=1.265
+ $X2=8.435 $Y2=0.58
r206 2 44 600 $w=1.7e-07 $l=9.22307e-07 $layer=licon1_PDIFF $count=1 $X=6.615
+ $Y=1.735 $X2=6.89 $Y2=2.53
r207 1 40 182 $w=1.7e-07 $l=6.65395e-07 $layer=licon1_NDIFF $count=1 $X=6.12
+ $Y=0.37 $X2=6.695 $Y2=0.565
.ends

.subckt PM_SKY130_FD_SC_HS__DFRBP_1%A_2026_424# 1 2 9 11 13 16 20 24 27
r50 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.965
+ $Y=1.465 $X2=10.965 $Y2=1.465
r51 22 27 0.364692 $w=3.3e-07 $l=1.25e-07 $layer=LI1_cond $X=10.44 $Y=1.465
+ $X2=10.315 $Y2=1.465
r52 22 24 18.3343 $w=3.28e-07 $l=5.25e-07 $layer=LI1_cond $X=10.44 $Y=1.465
+ $X2=10.965 $Y2=1.465
r53 18 27 6.46576 $w=2.5e-07 $l=1.65e-07 $layer=LI1_cond $X=10.315 $Y=1.63
+ $X2=10.315 $Y2=1.465
r54 18 20 29.5025 $w=2.48e-07 $l=6.4e-07 $layer=LI1_cond $X=10.315 $Y=1.63
+ $X2=10.315 $Y2=2.27
r55 14 27 6.46576 $w=2.5e-07 $l=1.65e-07 $layer=LI1_cond $X=10.315 $Y=1.3
+ $X2=10.315 $Y2=1.465
r56 14 16 30.4245 $w=2.48e-07 $l=6.6e-07 $layer=LI1_cond $X=10.315 $Y=1.3
+ $X2=10.315 $Y2=0.64
r57 11 25 61.4066 $w=2.86e-07 $l=3.24037e-07 $layer=POLY_cond $X=11.015 $Y=1.765
+ $X2=10.965 $Y2=1.465
r58 11 13 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=11.015 $Y=1.765
+ $X2=11.015 $Y2=2.4
r59 7 25 38.6549 $w=2.86e-07 $l=1.88348e-07 $layer=POLY_cond $X=11.015 $Y=1.3
+ $X2=10.965 $Y2=1.465
r60 7 9 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=11.015 $Y=1.3
+ $X2=11.015 $Y2=0.74
r61 2 20 300 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=2 $X=10.13
+ $Y=2.12 $X2=10.275 $Y2=2.27
r62 1 16 182 $w=1.7e-07 $l=3.34739e-07 $layer=licon1_NDIFF $count=1 $X=10.155
+ $Y=0.37 $X2=10.3 $Y2=0.64
.ends

.subckt PM_SKY130_FD_SC_HS__DFRBP_1%VPWR 1 2 3 4 5 6 7 8 25 27 31 35 39 43 49 51
+ 55 59 63 65 70 75 83 88 93 103 104 110 113 116 119 122 125 128
r140 128 129 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.8 $Y=3.33
+ $X2=10.8 $Y2=3.33
r141 125 126 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r142 123 126 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=7.92 $Y=3.33
+ $X2=8.88 $Y2=3.33
r143 122 123 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r144 119 120 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r145 116 117 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r146 113 114 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r147 110 111 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r148 107 108 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r149 104 129 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.28 $Y=3.33
+ $X2=10.8 $Y2=3.33
r150 103 104 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.28 $Y=3.33
+ $X2=11.28 $Y2=3.33
r151 101 128 7.94884 $w=1.7e-07 $l=1.48e-07 $layer=LI1_cond $X=10.905 $Y=3.33
+ $X2=10.757 $Y2=3.33
r152 101 103 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=10.905 $Y=3.33
+ $X2=11.28 $Y2=3.33
r153 100 129 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.32 $Y=3.33
+ $X2=10.8 $Y2=3.33
r154 99 100 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=10.32 $Y=3.33
+ $X2=10.32 $Y2=3.33
r155 97 100 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=9.36 $Y=3.33
+ $X2=10.32 $Y2=3.33
r156 97 126 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.36 $Y=3.33
+ $X2=8.88 $Y2=3.33
r157 96 99 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=9.36 $Y=3.33
+ $X2=10.32 $Y2=3.33
r158 96 97 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=9.36 $Y=3.33
+ $X2=9.36 $Y2=3.33
r159 94 125 6.25164 $w=1.7e-07 $l=1.08e-07 $layer=LI1_cond $X=9.025 $Y=3.33
+ $X2=8.917 $Y2=3.33
r160 94 96 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=9.025 $Y=3.33
+ $X2=9.36 $Y2=3.33
r161 93 128 7.94884 $w=1.7e-07 $l=1.47e-07 $layer=LI1_cond $X=10.61 $Y=3.33
+ $X2=10.757 $Y2=3.33
r162 93 99 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=10.61 $Y=3.33
+ $X2=10.32 $Y2=3.33
r163 92 123 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=7.92 $Y2=3.33
r164 92 120 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=6 $Y2=3.33
r165 91 92 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r166 89 119 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.03 $Y=3.33
+ $X2=5.905 $Y2=3.33
r167 89 91 91.9893 $w=1.68e-07 $l=1.41e-06 $layer=LI1_cond $X=6.03 $Y=3.33
+ $X2=7.44 $Y2=3.33
r168 88 122 6.47928 $w=1.7e-07 $l=1.12e-07 $layer=LI1_cond $X=7.835 $Y=3.33
+ $X2=7.947 $Y2=3.33
r169 88 91 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=7.835 $Y=3.33
+ $X2=7.44 $Y2=3.33
r170 87 117 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=4.56 $Y2=3.33
r171 86 87 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r172 84 116 8.88104 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=4.785 $Y=3.33
+ $X2=4.612 $Y2=3.33
r173 84 86 47.9519 $w=1.68e-07 $l=7.35e-07 $layer=LI1_cond $X=4.785 $Y=3.33
+ $X2=5.52 $Y2=3.33
r174 83 119 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.78 $Y=3.33
+ $X2=5.905 $Y2=3.33
r175 83 86 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=5.78 $Y=3.33
+ $X2=5.52 $Y2=3.33
r176 82 117 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=4.56 $Y2=3.33
r177 81 82 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r178 79 82 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=4.08 $Y2=3.33
r179 79 114 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=2.16 $Y2=3.33
r180 78 81 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=2.64 $Y=3.33
+ $X2=4.08 $Y2=3.33
r181 78 79 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r182 76 113 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.355 $Y=3.33
+ $X2=2.19 $Y2=3.33
r183 76 78 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=2.355 $Y=3.33
+ $X2=2.64 $Y2=3.33
r184 75 116 8.88104 $w=1.7e-07 $l=1.72e-07 $layer=LI1_cond $X=4.44 $Y=3.33
+ $X2=4.612 $Y2=3.33
r185 75 81 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=4.44 $Y=3.33
+ $X2=4.08 $Y2=3.33
r186 74 114 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r187 74 111 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r188 73 74 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r189 71 110 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.345 $Y=3.33
+ $X2=1.22 $Y2=3.33
r190 71 73 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=1.345 $Y=3.33
+ $X2=1.68 $Y2=3.33
r191 70 113 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.025 $Y=3.33
+ $X2=2.19 $Y2=3.33
r192 70 73 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=2.025 $Y=3.33
+ $X2=1.68 $Y2=3.33
r193 69 111 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r194 69 108 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r195 68 69 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r196 66 107 4.00981 $w=1.7e-07 $l=1.83e-07 $layer=LI1_cond $X=0.365 $Y=3.33
+ $X2=0.182 $Y2=3.33
r197 66 68 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=0.365 $Y=3.33
+ $X2=0.72 $Y2=3.33
r198 65 110 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.095 $Y=3.33
+ $X2=1.22 $Y2=3.33
r199 65 68 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=1.095 $Y=3.33
+ $X2=0.72 $Y2=3.33
r200 63 120 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=5.76 $Y=3.33
+ $X2=6 $Y2=3.33
r201 63 87 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=5.76 $Y=3.33
+ $X2=5.52 $Y2=3.33
r202 59 62 16.2123 $w=2.93e-07 $l=4.15e-07 $layer=LI1_cond $X=10.757 $Y=1.985
+ $X2=10.757 $Y2=2.4
r203 57 128 0.543863 $w=2.95e-07 $l=8.5e-08 $layer=LI1_cond $X=10.757 $Y=3.245
+ $X2=10.757 $Y2=3.33
r204 57 62 33.0107 $w=2.93e-07 $l=8.45e-07 $layer=LI1_cond $X=10.757 $Y=3.245
+ $X2=10.757 $Y2=2.4
r205 53 125 0.512231 $w=2.15e-07 $l=8.5e-08 $layer=LI1_cond $X=8.917 $Y=3.245
+ $X2=8.917 $Y2=3.33
r206 53 55 52.262 $w=2.13e-07 $l=9.75e-07 $layer=LI1_cond $X=8.917 $Y=3.245
+ $X2=8.917 $Y2=2.27
r207 52 122 6.47928 $w=1.7e-07 $l=1.13e-07 $layer=LI1_cond $X=8.06 $Y=3.33
+ $X2=7.947 $Y2=3.33
r208 51 125 6.25164 $w=1.7e-07 $l=1.07e-07 $layer=LI1_cond $X=8.81 $Y=3.33
+ $X2=8.917 $Y2=3.33
r209 51 52 48.9305 $w=1.68e-07 $l=7.5e-07 $layer=LI1_cond $X=8.81 $Y=3.33
+ $X2=8.06 $Y2=3.33
r210 47 122 0.355529 $w=2.25e-07 $l=8.5e-08 $layer=LI1_cond $X=7.947 $Y=3.245
+ $X2=7.947 $Y2=3.33
r211 47 49 34.8294 $w=2.23e-07 $l=6.8e-07 $layer=LI1_cond $X=7.947 $Y=3.245
+ $X2=7.947 $Y2=2.565
r212 43 46 31.5769 $w=2.48e-07 $l=6.85e-07 $layer=LI1_cond $X=5.905 $Y=1.905
+ $X2=5.905 $Y2=2.59
r213 41 119 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.905 $Y=3.245
+ $X2=5.905 $Y2=3.33
r214 41 46 30.194 $w=2.48e-07 $l=6.55e-07 $layer=LI1_cond $X=5.905 $Y=3.245
+ $X2=5.905 $Y2=2.59
r215 37 116 1.03204 $w=3.45e-07 $l=8.5e-08 $layer=LI1_cond $X=4.612 $Y=3.245
+ $X2=4.612 $Y2=3.33
r216 37 39 13.5287 $w=3.43e-07 $l=4.05e-07 $layer=LI1_cond $X=4.612 $Y=3.245
+ $X2=4.612 $Y2=2.84
r217 33 113 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.19 $Y=3.245
+ $X2=2.19 $Y2=3.33
r218 33 35 17.112 $w=3.28e-07 $l=4.9e-07 $layer=LI1_cond $X=2.19 $Y=3.245
+ $X2=2.19 $Y2=2.755
r219 29 110 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.22 $Y=3.245
+ $X2=1.22 $Y2=3.33
r220 29 31 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=1.22 $Y=3.245
+ $X2=1.22 $Y2=2.815
r221 25 107 3.13335 $w=2.5e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.24 $Y=3.245
+ $X2=0.182 $Y2=3.33
r222 25 27 22.8184 $w=2.48e-07 $l=4.95e-07 $layer=LI1_cond $X=0.24 $Y=3.245
+ $X2=0.24 $Y2=2.75
r223 8 62 300 $w=1.7e-07 $l=3.60832e-07 $layer=licon1_PDIFF $count=2 $X=10.575
+ $Y=2.12 $X2=10.76 $Y2=2.4
r224 8 59 600 $w=1.7e-07 $l=2.74317e-07 $layer=licon1_PDIFF $count=1 $X=10.575
+ $Y=2.12 $X2=10.79 $Y2=1.985
r225 7 55 300 $w=1.7e-07 $l=2.53969e-07 $layer=licon1_PDIFF $count=2 $X=8.705
+ $Y=2.355 $X2=8.92 $Y2=2.27
r226 6 49 600 $w=1.7e-07 $l=2.84341e-07 $layer=licon1_PDIFF $count=1 $X=7.745
+ $Y=2.355 $X2=7.92 $Y2=2.565
r227 5 46 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=5.72
+ $Y=1.735 $X2=5.865 $Y2=2.59
r228 5 43 400 $w=1.7e-07 $l=2.31409e-07 $layer=licon1_PDIFF $count=1 $X=5.72
+ $Y=1.735 $X2=5.865 $Y2=1.905
r229 4 39 600 $w=1.7e-07 $l=6.33739e-07 $layer=licon1_PDIFF $count=1 $X=4.37
+ $Y=2.315 $X2=4.61 $Y2=2.84
r230 3 35 600 $w=1.7e-07 $l=1.02727e-06 $layer=licon1_PDIFF $count=1 $X=2.04
+ $Y=1.8 $X2=2.19 $Y2=2.755
r231 2 31 600 $w=1.7e-07 $l=3.4187e-07 $layer=licon1_PDIFF $count=1 $X=1.03
+ $Y=2.54 $X2=1.18 $Y2=2.815
r232 1 27 600 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.54 $X2=0.28 $Y2=2.75
.ends

.subckt PM_SKY130_FD_SC_HS__DFRBP_1%A_38_78# 1 2 3 4 13 16 17 21 23 26 28 32 35
+ 43
c107 26 0 5.32615e-20 $X=3.755 $Y=2.075
c108 23 0 1.69357e-19 $X=3.67 $Y=2.16
c109 17 0 1.6736e-20 $X=3.065 $Y=2.395
r110 37 39 4.53993 $w=3.28e-07 $l=1.3e-07 $layer=LI1_cond $X=3.23 $Y=2.395
+ $X2=3.23 $Y2=2.525
r111 35 37 8.20679 $w=3.28e-07 $l=2.35e-07 $layer=LI1_cond $X=3.23 $Y=2.16
+ $X2=3.23 $Y2=2.395
r112 32 34 14.9345 $w=2.9e-07 $l=3.55e-07 $layer=LI1_cond $X=0.73 $Y=2.395
+ $X2=0.73 $Y2=2.75
r113 28 30 5.06376 $w=3.28e-07 $l=1.45e-07 $layer=LI1_cond $X=0.335 $Y=0.6
+ $X2=0.335 $Y2=0.745
r114 25 43 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.755 $Y=1.37
+ $X2=3.755 $Y2=1.285
r115 25 26 45.9947 $w=1.68e-07 $l=7.05e-07 $layer=LI1_cond $X=3.755 $Y=1.37
+ $X2=3.755 $Y2=2.075
r116 24 35 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.395 $Y=2.16
+ $X2=3.23 $Y2=2.16
r117 23 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.67 $Y=2.16
+ $X2=3.755 $Y2=2.075
r118 23 24 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=3.67 $Y=2.16
+ $X2=3.395 $Y2=2.16
r119 19 43 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=3.41 $Y=1.285
+ $X2=3.755 $Y2=1.285
r120 19 21 17.9781 $w=2.48e-07 $l=3.9e-07 $layer=LI1_cond $X=3.41 $Y=1.2
+ $X2=3.41 $Y2=0.81
r121 18 32 3.86198 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.895 $Y=2.395
+ $X2=0.73 $Y2=2.395
r122 17 37 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.065 $Y=2.395
+ $X2=3.23 $Y2=2.395
r123 17 18 141.572 $w=1.68e-07 $l=2.17e-06 $layer=LI1_cond $X=3.065 $Y=2.395
+ $X2=0.895 $Y2=2.395
r124 16 32 5.64745 $w=2.9e-07 $l=1.05119e-07 $layer=LI1_cond $X=0.775 $Y=2.31
+ $X2=0.73 $Y2=2.395
r125 15 16 96.5562 $w=1.68e-07 $l=1.48e-06 $layer=LI1_cond $X=0.775 $Y=0.83
+ $X2=0.775 $Y2=2.31
r126 14 30 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.5 $Y=0.745
+ $X2=0.335 $Y2=0.745
r127 13 15 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.69 $Y=0.745
+ $X2=0.775 $Y2=0.83
r128 13 14 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=0.69 $Y=0.745
+ $X2=0.5 $Y2=0.745
r129 4 39 600 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_PDIFF $count=1 $X=3.085
+ $Y=2.315 $X2=3.23 $Y2=2.525
r130 3 34 600 $w=1.7e-07 $l=2.74955e-07 $layer=licon1_PDIFF $count=1 $X=0.58
+ $Y=2.54 $X2=0.73 $Y2=2.75
r131 2 21 182 $w=1.7e-07 $l=2.83373e-07 $layer=licon1_NDIFF $count=1 $X=3.225
+ $Y=0.59 $X2=3.37 $Y2=0.81
r132 1 28 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=0.19
+ $Y=0.39 $X2=0.335 $Y2=0.6
.ends

.subckt PM_SKY130_FD_SC_HS__DFRBP_1%Q_N 1 2 9 11 12 13 26
c24 12 0 1.79977e-19 $X=9.84 $Y=2.405
r25 26 27 5.27602 $w=6.88e-07 $l=1.75e-07 $layer=LI1_cond $X=9.605 $Y=1.985
+ $X2=9.605 $Y2=1.81
r26 13 23 0.693379 $w=6.88e-07 $l=4e-08 $layer=LI1_cond $X=9.605 $Y=2.775
+ $X2=9.605 $Y2=2.815
r27 12 13 6.41375 $w=6.88e-07 $l=3.7e-07 $layer=LI1_cond $X=9.605 $Y=2.405
+ $X2=9.605 $Y2=2.775
r28 12 17 4.33362 $w=6.88e-07 $l=2.5e-07 $layer=LI1_cond $X=9.605 $Y=2.405
+ $X2=9.605 $Y2=2.155
r29 11 17 2.08014 $w=6.88e-07 $l=1.2e-07 $layer=LI1_cond $X=9.605 $Y=2.035
+ $X2=9.605 $Y2=2.155
r30 11 26 0.866723 $w=6.88e-07 $l=5e-08 $layer=LI1_cond $X=9.605 $Y=2.035
+ $X2=9.605 $Y2=1.985
r31 9 27 38.267 $w=3.88e-07 $l=1.295e-06 $layer=LI1_cond $X=9.755 $Y=0.515
+ $X2=9.755 $Y2=1.81
r32 2 26 200 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=3 $X=9.22
+ $Y=1.84 $X2=9.37 $Y2=1.985
r33 2 23 200 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=3 $X=9.22
+ $Y=1.84 $X2=9.37 $Y2=2.815
r34 1 9 91 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=2 $X=9.515
+ $Y=0.37 $X2=9.725 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__DFRBP_1%Q 1 2 9 10 11 24 27 35
r22 33 35 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=11.35 $Y=1.13
+ $X2=11.35 $Y2=1.82
r23 25 27 1.12043 $w=3.58e-07 $l=3.5e-08 $layer=LI1_cond $X=11.255 $Y=2
+ $X2=11.255 $Y2=2.035
r24 17 24 0.622942 $w=3.68e-07 $l=2e-08 $layer=LI1_cond $X=11.25 $Y=0.945
+ $X2=11.25 $Y2=0.925
r25 11 25 0.800308 $w=3.58e-07 $l=2.5e-08 $layer=LI1_cond $X=11.255 $Y=1.975
+ $X2=11.255 $Y2=2
r26 11 35 8.1909 $w=3.58e-07 $l=1.55e-07 $layer=LI1_cond $X=11.255 $Y=1.975
+ $X2=11.255 $Y2=1.82
r27 11 30 24.1693 $w=3.58e-07 $l=7.55e-07 $layer=LI1_cond $X=11.255 $Y=2.06
+ $X2=11.255 $Y2=2.815
r28 11 27 0.800308 $w=3.58e-07 $l=2.5e-08 $layer=LI1_cond $X=11.255 $Y=2.06
+ $X2=11.255 $Y2=2.035
r29 10 33 8.16504 $w=3.68e-07 $l=1.53e-07 $layer=LI1_cond $X=11.25 $Y=0.977
+ $X2=11.25 $Y2=1.13
r30 10 17 0.996707 $w=3.68e-07 $l=3.2e-08 $layer=LI1_cond $X=11.25 $Y=0.977
+ $X2=11.25 $Y2=0.945
r31 10 24 1.02785 $w=3.68e-07 $l=3.3e-08 $layer=LI1_cond $X=11.25 $Y=0.892
+ $X2=11.25 $Y2=0.925
r32 9 10 11.7425 $w=3.68e-07 $l=3.77e-07 $layer=LI1_cond $X=11.25 $Y=0.515
+ $X2=11.25 $Y2=0.892
r33 2 11 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=11.09
+ $Y=1.84 $X2=11.24 $Y2=1.985
r34 2 30 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=11.09
+ $Y=1.84 $X2=11.24 $Y2=2.815
r35 1 9 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=11.09
+ $Y=0.37 $X2=11.23 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__DFRBP_1%VGND 1 2 3 4 5 6 21 23 27 31 35 39 43 45 50
+ 55 63 68 75 76 79 82 86 92 95 98
r113 98 99 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.8 $Y=0 $X2=10.8
+ $Y2=0
r114 95 96 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=9.36 $Y=0 $X2=9.36
+ $Y2=0
r115 92 93 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=7.92 $Y=0 $X2=7.92
+ $Y2=0
r116 86 89 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=5.16 $Y=0 $X2=5.16
+ $Y2=0.325
r117 86 87 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r118 82 83 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r119 80 83 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r120 79 80 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r121 76 99 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.28 $Y=0
+ $X2=10.8 $Y2=0
r122 75 76 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.28 $Y=0
+ $X2=11.28 $Y2=0
r123 73 98 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=10.895 $Y=0
+ $X2=10.77 $Y2=0
r124 73 75 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=10.895 $Y=0
+ $X2=11.28 $Y2=0
r125 72 99 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.32 $Y=0
+ $X2=10.8 $Y2=0
r126 72 96 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=10.32 $Y=0
+ $X2=9.36 $Y2=0
r127 71 72 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=10.32 $Y=0
+ $X2=10.32 $Y2=0
r128 69 95 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=9.39 $Y=0 $X2=9.265
+ $Y2=0
r129 69 71 60.6738 $w=1.68e-07 $l=9.3e-07 $layer=LI1_cond $X=9.39 $Y=0 $X2=10.32
+ $Y2=0
r130 68 98 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=10.645 $Y=0
+ $X2=10.77 $Y2=0
r131 68 71 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=10.645 $Y=0
+ $X2=10.32 $Y2=0
r132 67 96 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=0 $X2=9.36
+ $Y2=0
r133 67 93 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=8.88 $Y=0 $X2=7.92
+ $Y2=0
r134 66 67 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=8.88 $Y=0 $X2=8.88
+ $Y2=0
r135 64 92 10.7288 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=7.995 $Y=0 $X2=7.765
+ $Y2=0
r136 64 66 57.738 $w=1.68e-07 $l=8.85e-07 $layer=LI1_cond $X=7.995 $Y=0 $X2=8.88
+ $Y2=0
r137 63 95 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=9.14 $Y=0 $X2=9.265
+ $Y2=0
r138 63 66 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=9.14 $Y=0 $X2=8.88
+ $Y2=0
r139 62 93 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=0 $X2=7.92
+ $Y2=0
r140 61 62 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=7.44 $Y=0
+ $X2=7.44 $Y2=0
r141 59 87 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=5.04
+ $Y2=0
r142 58 61 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=5.52 $Y=0 $X2=7.44
+ $Y2=0
r143 58 59 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=5.52 $Y=0
+ $X2=5.52 $Y2=0
r144 56 86 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.325 $Y=0 $X2=5.16
+ $Y2=0
r145 56 58 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=5.325 $Y=0
+ $X2=5.52 $Y2=0
r146 55 92 10.7288 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=7.535 $Y=0 $X2=7.765
+ $Y2=0
r147 55 61 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=7.535 $Y=0 $X2=7.44
+ $Y2=0
r148 54 87 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=2.64 $Y=0 $X2=5.04
+ $Y2=0
r149 54 83 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=2.16
+ $Y2=0
r150 53 54 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r151 51 82 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.42 $Y=0 $X2=2.255
+ $Y2=0
r152 51 53 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=2.42 $Y=0 $X2=2.64
+ $Y2=0
r153 50 86 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.995 $Y=0 $X2=5.16
+ $Y2=0
r154 50 53 153.642 $w=1.68e-07 $l=2.355e-06 $layer=LI1_cond $X=4.995 $Y=0
+ $X2=2.64 $Y2=0
r155 48 80 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r156 47 48 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r157 45 79 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.03 $Y=0 $X2=1.155
+ $Y2=0
r158 45 47 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=1.03 $Y=0 $X2=0.72
+ $Y2=0
r159 43 62 0.468274 $w=4.9e-07 $l=1.68e-06 $layer=MET1_cond $X=5.76 $Y=0
+ $X2=7.44 $Y2=0
r160 43 59 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=5.76 $Y=0
+ $X2=5.52 $Y2=0
r161 39 41 20.744 $w=2.48e-07 $l=4.5e-07 $layer=LI1_cond $X=10.77 $Y=0.515
+ $X2=10.77 $Y2=0.965
r162 37 98 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=10.77 $Y=0.085
+ $X2=10.77 $Y2=0
r163 37 39 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=10.77 $Y=0.085
+ $X2=10.77 $Y2=0.515
r164 33 95 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=9.265 $Y=0.085
+ $X2=9.265 $Y2=0
r165 33 35 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=9.265 $Y=0.085
+ $X2=9.265 $Y2=0.515
r166 29 92 1.85547 $w=4.6e-07 $l=8.5e-08 $layer=LI1_cond $X=7.765 $Y=0.085
+ $X2=7.765 $Y2=0
r167 29 31 12.2208 $w=4.58e-07 $l=4.7e-07 $layer=LI1_cond $X=7.765 $Y=0.085
+ $X2=7.765 $Y2=0.555
r168 25 82 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.255 $Y=0.085
+ $X2=2.255 $Y2=0
r169 25 27 17.112 $w=3.28e-07 $l=4.9e-07 $layer=LI1_cond $X=2.255 $Y=0.085
+ $X2=2.255 $Y2=0.575
r170 24 79 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.28 $Y=0 $X2=1.155
+ $Y2=0
r171 23 82 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.09 $Y=0 $X2=2.255
+ $Y2=0
r172 23 24 52.8449 $w=1.68e-07 $l=8.1e-07 $layer=LI1_cond $X=2.09 $Y=0 $X2=1.28
+ $Y2=0
r173 19 79 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.155 $Y=0.085
+ $X2=1.155 $Y2=0
r174 19 21 23.7403 $w=2.48e-07 $l=5.15e-07 $layer=LI1_cond $X=1.155 $Y=0.085
+ $X2=1.155 $Y2=0.6
r175 6 41 182 $w=1.7e-07 $l=6.87768e-07 $layer=licon1_NDIFF $count=1 $X=10.59
+ $Y=0.37 $X2=10.79 $Y2=0.965
r176 6 39 182 $w=1.7e-07 $l=2.62678e-07 $layer=licon1_NDIFF $count=1 $X=10.59
+ $Y=0.37 $X2=10.79 $Y2=0.515
r177 5 35 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=9.08
+ $Y=0.37 $X2=9.225 $Y2=0.515
r178 4 31 182 $w=1.7e-07 $l=2.82754e-07 $layer=licon1_NDIFF $count=1 $X=7.56
+ $Y=0.37 $X2=7.765 $Y2=0.555
r179 3 89 182 $w=1.7e-07 $l=3.58504e-07 $layer=licon1_NDIFF $count=1 $X=4.94
+ $Y=0.59 $X2=5.16 $Y2=0.325
r180 2 27 182 $w=1.7e-07 $l=2.95212e-07 $layer=licon1_NDIFF $count=1 $X=2.045
+ $Y=0.37 $X2=2.255 $Y2=0.575
r181 1 21 182 $w=1.7e-07 $l=2.86182e-07 $layer=licon1_NDIFF $count=1 $X=1.015
+ $Y=0.39 $X2=1.195 $Y2=0.6
.ends

