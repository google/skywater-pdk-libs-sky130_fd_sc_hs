* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hs__o21ba_4 A1 A2 B1_N VGND VNB VPB VPWR X
M1000 a_193_48# a_27_368# VPWR VPB pshort w=840000u l=150000u
+  ad=5.52e+11p pd=4.88e+06u as=2.2288e+12p ps=1.517e+07u
M1001 VPWR a_27_368# a_193_48# VPB pshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1002 VGND a_193_48# X VNB nlowvt w=740000u l=150000u
+  ad=1.0914e+12p pd=1.012e+07u as=4.218e+11p ps=4.1e+06u
M1003 VGND A2 a_618_94# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=7.9445e+11p ps=7.84e+06u
M1004 a_892_392# A1 VPWR VPB pshort w=1e+06u l=150000u
+  ad=6e+11p pd=5.2e+06u as=0p ps=0u
M1005 VGND a_193_48# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_618_94# A1 VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_193_48# a_27_368# a_618_94# VNB nlowvt w=640000u l=150000u
+  ad=1.792e+11p pd=1.84e+06u as=0p ps=0u
M1008 a_193_48# A2 a_892_392# VPB pshort w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_618_94# A2 VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VGND A1 a_618_94# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 X a_193_48# VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=6.72e+11p pd=5.68e+06u as=0p ps=0u
M1012 VPWR a_193_48# X VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 X a_193_48# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 X a_193_48# VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_892_392# A2 a_193_48# VPB pshort w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VPWR B1_N a_27_368# VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=3.304e+11p ps=2.83e+06u
M1017 VPWR a_193_48# X VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 VPWR A1 a_892_392# VPB pshort w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_618_94# a_27_368# a_193_48# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 X a_193_48# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 VGND B1_N a_27_368# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
.ends
