* File: sky130_fd_sc_hs__or3b_2.spice
* Created: Tue Sep  1 20:20:50 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hs__or3b_2.pex.spice"
.subckt sky130_fd_sc_hs__or3b_2  VNB VPB C_N A B VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* B	B
* A	A
* C_N	C_N
* VPB	VPB
* VNB	VNB
MM1007 N_VGND_M1007_d N_C_N_M1007_g N_A_27_368#_M1007_s VNB NLOWVT L=0.15 W=0.55
+ AD=0.107506 AS=0.15675 PD=0.937984 PS=1.67 NRD=18.54 NRS=0 M=1 R=3.66667
+ SA=75000.2 SB=75002.9 A=0.0825 P=1.4 MULT=1
MM1006 N_X_M1006_d N_A_190_260#_M1006_g N_VGND_M1007_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.144644 PD=1.02 PS=1.26202 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.6
+ SB=75002.2 A=0.111 P=1.78 MULT=1
MM1011 N_X_M1006_d N_A_190_260#_M1011_g N_VGND_M1011_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.210739 PD=1.02 PS=1.41029 NRD=0 NRS=29.184 M=1 R=4.93333
+ SA=75001 SB=75001.8 A=0.111 P=1.78 MULT=1
MM1010 N_A_190_260#_M1010_d N_A_M1010_g N_VGND_M1011_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.112 AS=0.182261 PD=0.99 PS=1.21971 NRD=13.116 NRS=21.552 M=1 R=4.26667
+ SA=75001.8 SB=75001.3 A=0.096 P=1.58 MULT=1
MM1008 N_VGND_M1008_d N_B_M1008_g N_A_190_260#_M1010_d VNB NLOWVT L=0.15 W=0.64
+ AD=0.1344 AS=0.112 PD=1.06 PS=0.99 NRD=13.116 NRS=0 M=1 R=4.26667 SA=75002.3
+ SB=75000.8 A=0.096 P=1.58 MULT=1
MM1001 N_A_190_260#_M1001_d N_A_27_368#_M1001_g N_VGND_M1008_d VNB NLOWVT L=0.15
+ W=0.64 AD=0.1824 AS=0.1344 PD=1.85 PS=1.06 NRD=0 NRS=13.116 M=1 R=4.26667
+ SA=75002.9 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1009 N_VPWR_M1009_d N_C_N_M1009_g N_A_27_368#_M1009_s VPB PSHORT L=0.15 W=0.84
+ AD=0.174 AS=0.2478 PD=1.29 PS=2.27 NRD=35.6767 NRS=2.3443 M=1 R=5.6 SA=75000.2
+ SB=75002.9 A=0.126 P=1.98 MULT=1
MM1002 N_X_M1002_d N_A_190_260#_M1002_g N_VPWR_M1009_d VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.232 PD=1.42 PS=1.72 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.6 SB=75002.2 A=0.168 P=2.54 MULT=1
MM1003 N_X_M1002_d N_A_190_260#_M1003_g N_VPWR_M1003_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.336608 PD=1.42 PS=1.80151 NRD=1.7533 NRS=25.4918 M=1 R=7.46667
+ SA=75001.1 SB=75001.7 A=0.168 P=2.54 MULT=1
MM1005 A_458_368# N_A_M1005_g N_VPWR_M1003_s VPB PSHORT L=0.15 W=1 AD=0.135
+ AS=0.300542 PD=1.27 PS=1.60849 NRD=15.7403 NRS=30.5153 M=1 R=6.66667
+ SA=75001.8 SB=75001.2 A=0.15 P=2.3 MULT=1
MM1000 A_542_368# N_B_M1000_g A_458_368# VPB PSHORT L=0.15 W=1 AD=0.195 AS=0.135
+ PD=1.39 PS=1.27 NRD=27.5603 NRS=15.7403 M=1 R=6.66667 SA=75002.3 SB=75000.8
+ A=0.15 P=2.3 MULT=1
MM1004 N_A_190_260#_M1004_d N_A_27_368#_M1004_g A_542_368# VPB PSHORT L=0.15 W=1
+ AD=0.295 AS=0.195 PD=2.59 PS=1.39 NRD=1.9503 NRS=27.5603 M=1 R=6.66667
+ SA=75002.8 SB=75000.2 A=0.15 P=2.3 MULT=1
DX12_noxref VNB VPB NWDIODE A=7.8492 P=12.16
*
.include "sky130_fd_sc_hs__or3b_2.pxi.spice"
*
.ends
*
*
