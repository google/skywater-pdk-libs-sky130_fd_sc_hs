* File: sky130_fd_sc_hs__decap_4.pxi.spice
* Created: Tue Sep  1 19:59:09 2020
* 
x_PM_SKY130_FD_SC_HS__DECAP_4%VGND N_VGND_M1001_s N_VGND_M1000_g N_VGND_c_20_n
+ N_VGND_c_21_n N_VGND_c_22_n N_VGND_c_23_n N_VGND_c_24_n VGND N_VGND_c_25_n
+ N_VGND_c_26_n PM_SKY130_FD_SC_HS__DECAP_4%VGND
x_PM_SKY130_FD_SC_HS__DECAP_4%VPWR N_VPWR_M1000_s N_VPWR_M1001_g N_VPWR_c_45_n
+ N_VPWR_c_49_n N_VPWR_c_50_n N_VPWR_c_51_n N_VPWR_c_52_n N_VPWR_c_46_n
+ N_VPWR_c_47_n VPWR N_VPWR_c_48_n PM_SKY130_FD_SC_HS__DECAP_4%VPWR
cc_1 VNB N_VGND_c_20_n 0.0180938f $X=-0.19 $Y=-0.245 $X2=0.455 $Y2=0.085
cc_2 VNB N_VGND_c_21_n 0.0675204f $X=-0.19 $Y=-0.245 $X2=0.335 $Y2=0.64
cc_3 VNB N_VGND_c_22_n 0.042044f $X=-0.19 $Y=-0.245 $X2=0.575 $Y2=1.42
cc_4 VNB N_VGND_c_23_n 0.0127868f $X=-0.19 $Y=-0.245 $X2=1.615 $Y2=0.085
cc_5 VNB N_VGND_c_24_n 0.0274307f $X=-0.19 $Y=-0.245 $X2=1.615 $Y2=0.64
cc_6 VNB N_VGND_c_25_n 0.0221481f $X=-0.19 $Y=-0.245 $X2=1.45 $Y2=0
cc_7 VNB N_VGND_c_26_n 0.132293f $X=-0.19 $Y=-0.245 $X2=1.68 $Y2=0
cc_8 VNB N_VPWR_c_45_n 0.12629f $X=-0.19 $Y=-0.245 $X2=0.91 $Y2=1.83
cc_9 VNB N_VPWR_c_46_n 0.0216619f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_VPWR_c_47_n 0.0573234f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_VPWR_c_48_n 0.0840719f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VPB N_VGND_M1000_g 0.102919f $X=-0.19 $Y=1.66 $X2=0.91 $Y2=2.46
cc_13 VPB N_VGND_c_22_n 0.0193702f $X=-0.19 $Y=1.66 $X2=0.575 $Y2=1.42
cc_14 VPB N_VPWR_c_49_n 0.0113726f $X=-0.19 $Y=1.66 $X2=0.455 $Y2=0.64
cc_15 VPB N_VPWR_c_50_n 0.056103f $X=-0.19 $Y=1.66 $X2=0.455 $Y2=1.42
cc_16 VPB N_VPWR_c_51_n 0.0225322f $X=-0.19 $Y=1.66 $X2=1.615 $Y2=0.085
cc_17 VPB N_VPWR_c_52_n 0.0192666f $X=-0.19 $Y=1.66 $X2=1.615 $Y2=0.64
cc_18 VPB N_VPWR_c_46_n 0.0662839f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_19 VPB N_VPWR_c_48_n 0.0478118f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_20 N_VGND_c_21_n N_VPWR_c_45_n 0.0773177f $X=0.335 $Y=0.64 $X2=0 $Y2=0
cc_21 N_VGND_c_22_n N_VPWR_c_45_n 0.0173516f $X=0.575 $Y=1.42 $X2=0 $Y2=0
cc_22 N_VGND_c_24_n N_VPWR_c_45_n 0.0335332f $X=1.615 $Y=0.64 $X2=0 $Y2=0
cc_23 N_VGND_c_25_n N_VPWR_c_45_n 0.0220076f $X=1.45 $Y=0 $X2=0 $Y2=0
cc_24 N_VGND_c_26_n N_VPWR_c_45_n 0.0428939f $X=1.68 $Y=0 $X2=0 $Y2=0
cc_25 N_VGND_M1000_g N_VPWR_c_50_n 0.0605103f $X=0.91 $Y=2.46 $X2=0 $Y2=0
cc_26 N_VGND_c_21_n N_VPWR_c_50_n 0.0143348f $X=0.335 $Y=0.64 $X2=0 $Y2=0
cc_27 N_VGND_M1000_g N_VPWR_c_51_n 0.0221223f $X=0.91 $Y=2.46 $X2=0 $Y2=0
cc_28 N_VGND_M1000_g N_VPWR_c_46_n 0.108651f $X=0.91 $Y=2.46 $X2=0 $Y2=0
cc_29 N_VGND_c_21_n N_VPWR_c_46_n 0.0136195f $X=0.335 $Y=0.64 $X2=0 $Y2=0
cc_30 N_VGND_c_22_n N_VPWR_c_46_n 0.00969158f $X=0.575 $Y=1.42 $X2=0 $Y2=0
cc_31 N_VGND_c_24_n N_VPWR_c_46_n 0.0106491f $X=1.615 $Y=0.64 $X2=0 $Y2=0
cc_32 N_VGND_M1000_g N_VPWR_c_47_n 0.0139884f $X=0.91 $Y=2.46 $X2=0 $Y2=0
cc_33 N_VGND_c_21_n N_VPWR_c_47_n 0.00834649f $X=0.335 $Y=0.64 $X2=0 $Y2=0
cc_34 N_VGND_c_22_n N_VPWR_c_47_n 0.00887584f $X=0.575 $Y=1.42 $X2=0 $Y2=0
cc_35 N_VGND_M1000_g N_VPWR_c_48_n 0.0434015f $X=0.91 $Y=2.46 $X2=0 $Y2=0
