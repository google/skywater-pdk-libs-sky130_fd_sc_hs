* File: sky130_fd_sc_hs__a2111o_4.pxi.spice
* Created: Thu Aug 27 20:22:44 2020
* 
x_PM_SKY130_FD_SC_HS__A2111O_4%A_137_260# N_A_137_260#_M1017_d
+ N_A_137_260#_M1006_s N_A_137_260#_M1012_s N_A_137_260#_M1001_d
+ N_A_137_260#_M1010_d N_A_137_260#_c_176_n N_A_137_260#_M1008_g
+ N_A_137_260#_c_177_n N_A_137_260#_M1011_g N_A_137_260#_M1005_g
+ N_A_137_260#_c_178_n N_A_137_260#_M1013_g N_A_137_260#_M1016_g
+ N_A_137_260#_c_179_n N_A_137_260#_M1014_g N_A_137_260#_M1021_g
+ N_A_137_260#_M1025_g N_A_137_260#_c_162_n N_A_137_260#_c_163_n
+ N_A_137_260#_c_164_n N_A_137_260#_c_165_n N_A_137_260#_c_181_n
+ N_A_137_260#_c_166_n N_A_137_260#_c_167_n N_A_137_260#_c_168_n
+ N_A_137_260#_c_169_n N_A_137_260#_c_170_n N_A_137_260#_c_171_n
+ N_A_137_260#_c_172_n N_A_137_260#_c_173_n N_A_137_260#_c_182_n
+ N_A_137_260#_c_174_n N_A_137_260#_c_175_n
+ PM_SKY130_FD_SC_HS__A2111O_4%A_137_260#
x_PM_SKY130_FD_SC_HS__A2111O_4%D1 N_D1_M1017_g N_D1_c_341_n N_D1_c_347_n
+ N_D1_M1010_g N_D1_M1022_g N_D1_c_343_n N_D1_c_349_n N_D1_M1015_g D1
+ N_D1_c_344_n N_D1_c_345_n PM_SKY130_FD_SC_HS__A2111O_4%D1
x_PM_SKY130_FD_SC_HS__A2111O_4%C1 N_C1_M1006_g N_C1_c_413_n N_C1_M1018_g
+ N_C1_M1023_g N_C1_c_408_n N_C1_c_414_n N_C1_M1020_g N_C1_c_409_n N_C1_c_410_n
+ C1 C1 C1 N_C1_c_412_n PM_SKY130_FD_SC_HS__A2111O_4%C1
x_PM_SKY130_FD_SC_HS__A2111O_4%B1 N_B1_c_473_n N_B1_M1012_g N_B1_c_474_n
+ N_B1_c_475_n N_B1_c_476_n N_B1_M1026_g N_B1_c_479_n N_B1_M1000_g N_B1_c_480_n
+ N_B1_M1024_g B1 B1 N_B1_c_478_n PM_SKY130_FD_SC_HS__A2111O_4%B1
x_PM_SKY130_FD_SC_HS__A2111O_4%A1 N_A1_c_534_n N_A1_M1002_g N_A1_M1001_g
+ N_A1_c_535_n N_A1_M1003_g N_A1_M1019_g A1 A1 N_A1_c_533_n
+ PM_SKY130_FD_SC_HS__A2111O_4%A1
x_PM_SKY130_FD_SC_HS__A2111O_4%A2 N_A2_c_584_n N_A2_c_591_n N_A2_M1004_g
+ N_A2_M1009_g N_A2_c_586_n N_A2_c_593_n N_A2_M1007_g N_A2_M1027_g A2 A2
+ N_A2_c_589_n PM_SKY130_FD_SC_HS__A2111O_4%A2
x_PM_SKY130_FD_SC_HS__A2111O_4%VPWR N_VPWR_M1008_s N_VPWR_M1011_s N_VPWR_M1014_s
+ N_VPWR_M1002_d N_VPWR_M1004_d N_VPWR_c_634_n N_VPWR_c_635_n N_VPWR_c_636_n
+ N_VPWR_c_637_n N_VPWR_c_638_n N_VPWR_c_639_n N_VPWR_c_640_n N_VPWR_c_641_n
+ N_VPWR_c_642_n N_VPWR_c_643_n N_VPWR_c_644_n VPWR N_VPWR_c_645_n
+ N_VPWR_c_646_n N_VPWR_c_647_n N_VPWR_c_633_n N_VPWR_c_649_n N_VPWR_c_650_n
+ PM_SKY130_FD_SC_HS__A2111O_4%VPWR
x_PM_SKY130_FD_SC_HS__A2111O_4%X N_X_M1005_s N_X_M1021_s N_X_M1008_d N_X_M1013_d
+ N_X_c_734_n N_X_c_735_n N_X_c_741_n N_X_c_742_n N_X_c_743_n N_X_c_744_n
+ N_X_c_736_n N_X_c_737_n N_X_c_745_n N_X_c_738_n N_X_c_746_n N_X_c_739_n X X
+ PM_SKY130_FD_SC_HS__A2111O_4%X
x_PM_SKY130_FD_SC_HS__A2111O_4%A_549_392# N_A_549_392#_M1010_s
+ N_A_549_392#_M1015_s N_A_549_392#_M1020_s N_A_549_392#_c_812_n
+ N_A_549_392#_c_813_n N_A_549_392#_c_814_n N_A_549_392#_c_815_n
+ N_A_549_392#_c_816_n N_A_549_392#_c_817_n N_A_549_392#_c_818_n
+ PM_SKY130_FD_SC_HS__A2111O_4%A_549_392#
x_PM_SKY130_FD_SC_HS__A2111O_4%A_814_392# N_A_814_392#_M1018_d
+ N_A_814_392#_M1000_s N_A_814_392#_c_860_n N_A_814_392#_c_861_n
+ N_A_814_392#_c_862_n PM_SKY130_FD_SC_HS__A2111O_4%A_814_392#
x_PM_SKY130_FD_SC_HS__A2111O_4%A_1013_392# N_A_1013_392#_M1000_d
+ N_A_1013_392#_M1024_d N_A_1013_392#_M1003_s N_A_1013_392#_M1007_s
+ N_A_1013_392#_c_890_n N_A_1013_392#_c_891_n N_A_1013_392#_c_892_n
+ N_A_1013_392#_c_893_n N_A_1013_392#_c_928_n N_A_1013_392#_c_894_n
+ N_A_1013_392#_c_895_n N_A_1013_392#_c_896_n N_A_1013_392#_c_897_n
+ N_A_1013_392#_c_898_n N_A_1013_392#_c_899_n
+ PM_SKY130_FD_SC_HS__A2111O_4%A_1013_392#
x_PM_SKY130_FD_SC_HS__A2111O_4%VGND N_VGND_M1005_d N_VGND_M1016_d N_VGND_M1025_d
+ N_VGND_M1022_s N_VGND_M1023_d N_VGND_M1026_d N_VGND_M1009_s N_VGND_c_948_n
+ N_VGND_c_949_n N_VGND_c_950_n N_VGND_c_951_n N_VGND_c_952_n N_VGND_c_953_n
+ N_VGND_c_954_n N_VGND_c_955_n N_VGND_c_956_n N_VGND_c_957_n N_VGND_c_958_n
+ N_VGND_c_959_n N_VGND_c_960_n VGND N_VGND_c_961_n N_VGND_c_962_n
+ N_VGND_c_963_n N_VGND_c_964_n N_VGND_c_965_n N_VGND_c_966_n N_VGND_c_967_n
+ N_VGND_c_968_n N_VGND_c_969_n N_VGND_c_970_n PM_SKY130_FD_SC_HS__A2111O_4%VGND
x_PM_SKY130_FD_SC_HS__A2111O_4%A_1210_74# N_A_1210_74#_M1001_s
+ N_A_1210_74#_M1019_s N_A_1210_74#_M1027_d N_A_1210_74#_c_1062_n
+ N_A_1210_74#_c_1063_n N_A_1210_74#_c_1064_n N_A_1210_74#_c_1065_n
+ N_A_1210_74#_c_1066_n N_A_1210_74#_c_1067_n
+ PM_SKY130_FD_SC_HS__A2111O_4%A_1210_74#
cc_1 VNB N_A_137_260#_M1005_g 0.0246266f $X=-0.19 $Y=-0.245 $X2=1.285 $Y2=0.74
cc_2 VNB N_A_137_260#_M1016_g 0.0209331f $X=-0.19 $Y=-0.245 $X2=1.715 $Y2=0.74
cc_3 VNB N_A_137_260#_M1021_g 0.0209331f $X=-0.19 $Y=-0.245 $X2=2.145 $Y2=0.74
cc_4 VNB N_A_137_260#_M1025_g 0.021412f $X=-0.19 $Y=-0.245 $X2=2.575 $Y2=0.74
cc_5 VNB N_A_137_260#_c_162_n 0.0133831f $X=-0.19 $Y=-0.245 $X2=3.045 $Y2=1.465
cc_6 VNB N_A_137_260#_c_163_n 0.146983f $X=-0.19 $Y=-0.245 $X2=2.485 $Y2=1.465
cc_7 VNB N_A_137_260#_c_164_n 0.00206705f $X=-0.19 $Y=-0.245 $X2=3.265 $Y2=0.515
cc_8 VNB N_A_137_260#_c_165_n 0.00164495f $X=-0.19 $Y=-0.245 $X2=3.13 $Y2=1.3
cc_9 VNB N_A_137_260#_c_166_n 0.00791729f $X=-0.19 $Y=-0.245 $X2=4.05 $Y2=1.005
cc_10 VNB N_A_137_260#_c_167_n 0.00178908f $X=-0.19 $Y=-0.245 $X2=4.135
+ $Y2=0.515
cc_11 VNB N_A_137_260#_c_168_n 0.00917015f $X=-0.19 $Y=-0.245 $X2=4.92 $Y2=1.195
cc_12 VNB N_A_137_260#_c_169_n 0.003224f $X=-0.19 $Y=-0.245 $X2=5.005 $Y2=0.515
cc_13 VNB N_A_137_260#_c_170_n 0.0167045f $X=-0.19 $Y=-0.245 $X2=6.51 $Y2=1.195
cc_14 VNB N_A_137_260#_c_171_n 9.35553e-19 $X=-0.19 $Y=-0.245 $X2=6.605 $Y2=0.79
cc_15 VNB N_A_137_260#_c_172_n 0.00256255f $X=-0.19 $Y=-0.245 $X2=3.197
+ $Y2=1.005
cc_16 VNB N_A_137_260#_c_173_n 2.54259e-19 $X=-0.19 $Y=-0.245 $X2=3.13 $Y2=1.465
cc_17 VNB N_A_137_260#_c_174_n 0.00425475f $X=-0.19 $Y=-0.245 $X2=4.135
+ $Y2=1.005
cc_18 VNB N_A_137_260#_c_175_n 0.00159638f $X=-0.19 $Y=-0.245 $X2=5.005
+ $Y2=1.195
cc_19 VNB N_D1_M1017_g 0.0243515f $X=-0.19 $Y=-0.245 $X2=4.865 $Y2=0.37
cc_20 VNB N_D1_c_341_n 0.00424565f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_D1_M1022_g 0.0233084f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_D1_c_343_n 0.00307356f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_D1_c_344_n 0.00521187f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_D1_c_345_n 0.0395761f $X=-0.19 $Y=-0.245 $X2=1.675 $Y2=1.765
cc_25 VNB N_C1_M1006_g 0.0328076f $X=-0.19 $Y=-0.245 $X2=4.865 $Y2=0.37
cc_26 VNB N_C1_c_408_n 0.0162228f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_C1_c_409_n 0.0149068f $X=-0.19 $Y=-0.245 $X2=0.775 $Y2=1.765
cc_28 VNB N_C1_c_410_n 0.00789277f $X=-0.19 $Y=-0.245 $X2=0.775 $Y2=2.4
cc_29 VNB C1 0.00771653f $X=-0.19 $Y=-0.245 $X2=1.225 $Y2=2.4
cc_30 VNB N_C1_c_412_n 0.0348531f $X=-0.19 $Y=-0.245 $X2=1.675 $Y2=2.4
cc_31 VNB N_B1_c_473_n 0.0150917f $X=-0.19 $Y=-0.245 $X2=3.125 $Y2=0.37
cc_32 VNB N_B1_c_474_n 0.0151763f $X=-0.19 $Y=-0.245 $X2=6.465 $Y2=0.37
cc_33 VNB N_B1_c_475_n 0.00874277f $X=-0.19 $Y=-0.245 $X2=3.17 $Y2=1.96
cc_34 VNB N_B1_c_476_n 0.019199f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB B1 0.00301796f $X=-0.19 $Y=-0.245 $X2=0.775 $Y2=1.765
cc_36 VNB N_B1_c_478_n 0.0973357f $X=-0.19 $Y=-0.245 $X2=1.225 $Y2=2.4
cc_37 VNB N_A1_M1001_g 0.0384872f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A1_M1019_g 0.0324852f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB A1 0.00484998f $X=-0.19 $Y=-0.245 $X2=0.775 $Y2=1.765
cc_40 VNB N_A1_c_533_n 0.0272667f $X=-0.19 $Y=-0.245 $X2=1.285 $Y2=0.74
cc_41 VNB N_A2_c_584_n 0.00347224f $X=-0.19 $Y=-0.245 $X2=3.995 $Y2=0.37
cc_42 VNB N_A2_M1009_g 0.0233949f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A2_c_586_n 0.00418093f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A2_M1027_g 0.0324492f $X=-0.19 $Y=-0.245 $X2=0.775 $Y2=2.4
cc_45 VNB A2 0.0203442f $X=-0.19 $Y=-0.245 $X2=1.225 $Y2=2.4
cc_46 VNB N_A2_c_589_n 0.0436625f $X=-0.19 $Y=-0.245 $X2=1.715 $Y2=0.74
cc_47 VNB N_VPWR_c_633_n 0.342803f $X=-0.19 $Y=-0.245 $X2=6.51 $Y2=1.195
cc_48 VNB N_X_c_734_n 0.0153235f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_X_c_735_n 0.0316066f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_X_c_736_n 0.00206666f $X=-0.19 $Y=-0.245 $X2=1.675 $Y2=2.4
cc_51 VNB N_X_c_737_n 0.00423905f $X=-0.19 $Y=-0.245 $X2=1.715 $Y2=1.3
cc_52 VNB N_X_c_738_n 0.00206666f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_X_c_739_n 0.00178779f $X=-0.19 $Y=-0.245 $X2=3.045 $Y2=1.465
cc_54 VNB X 0.0359413f $X=-0.19 $Y=-0.245 $X2=1.035 $Y2=1.465
cc_55 VNB N_VGND_c_948_n 0.0254564f $X=-0.19 $Y=-0.245 $X2=1.285 $Y2=0.74
cc_56 VNB N_VGND_c_949_n 0.0065212f $X=-0.19 $Y=-0.245 $X2=1.675 $Y2=2.4
cc_57 VNB N_VGND_c_950_n 0.0172524f $X=-0.19 $Y=-0.245 $X2=1.715 $Y2=0.74
cc_58 VNB N_VGND_c_951_n 0.00424579f $X=-0.19 $Y=-0.245 $X2=2.125 $Y2=2.4
cc_59 VNB N_VGND_c_952_n 0.0182548f $X=-0.19 $Y=-0.245 $X2=2.145 $Y2=1.3
cc_60 VNB N_VGND_c_953_n 0.00266729f $X=-0.19 $Y=-0.245 $X2=2.575 $Y2=1.3
cc_61 VNB N_VGND_c_954_n 0.00250542f $X=-0.19 $Y=-0.245 $X2=3.045 $Y2=1.465
cc_62 VNB N_VGND_c_955_n 0.0158756f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_VGND_c_956_n 0.00396467f $X=-0.19 $Y=-0.245 $X2=3.197 $Y2=0.92
cc_64 VNB N_VGND_c_957_n 0.0309422f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_VGND_c_958_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=3.13 $Y2=1.09
cc_66 VNB N_VGND_c_959_n 0.0172524f $X=-0.19 $Y=-0.245 $X2=3.13 $Y2=1.3
cc_67 VNB N_VGND_c_960_n 0.00326991f $X=-0.19 $Y=-0.245 $X2=3.13 $Y2=1.63
cc_68 VNB N_VGND_c_961_n 0.0151736f $X=-0.19 $Y=-0.245 $X2=4.92 $Y2=1.195
cc_69 VNB N_VGND_c_962_n 0.0151736f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_VGND_c_963_n 0.0440384f $X=-0.19 $Y=-0.245 $X2=6.605 $Y2=0.79
cc_71 VNB N_VGND_c_964_n 0.0169136f $X=-0.19 $Y=-0.245 $X2=3.32 $Y2=2.115
cc_72 VNB N_VGND_c_965_n 0.481891f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_VGND_c_966_n 0.00461913f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_VGND_c_967_n 0.00622543f $X=-0.19 $Y=-0.245 $X2=1.035 $Y2=1.532
cc_75 VNB N_VGND_c_968_n 0.00622543f $X=-0.19 $Y=-0.245 $X2=1.675 $Y2=1.532
cc_76 VNB N_VGND_c_969_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=2.145 $Y2=1.532
cc_77 VNB N_VGND_c_970_n 0.00604233f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_A_1210_74#_c_1062_n 0.00750863f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VNB N_A_1210_74#_c_1063_n 0.00445625f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_A_1210_74#_c_1064_n 0.00514874f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_81 VNB N_A_1210_74#_c_1065_n 0.0137881f $X=-0.19 $Y=-0.245 $X2=1.225 $Y2=2.4
cc_82 VNB N_A_1210_74#_c_1066_n 0.00403069f $X=-0.19 $Y=-0.245 $X2=1.225 $Y2=2.4
cc_83 VNB N_A_1210_74#_c_1067_n 0.0237116f $X=-0.19 $Y=-0.245 $X2=1.285 $Y2=0.74
cc_84 VPB N_A_137_260#_c_176_n 0.0164045f $X=-0.19 $Y=1.66 $X2=0.775 $Y2=1.765
cc_85 VPB N_A_137_260#_c_177_n 0.0152454f $X=-0.19 $Y=1.66 $X2=1.225 $Y2=1.765
cc_86 VPB N_A_137_260#_c_178_n 0.015247f $X=-0.19 $Y=1.66 $X2=1.675 $Y2=1.765
cc_87 VPB N_A_137_260#_c_179_n 0.017577f $X=-0.19 $Y=1.66 $X2=2.125 $Y2=1.765
cc_88 VPB N_A_137_260#_c_163_n 0.0294594f $X=-0.19 $Y=1.66 $X2=2.485 $Y2=1.465
cc_89 VPB N_A_137_260#_c_181_n 0.00260106f $X=-0.19 $Y=1.66 $X2=3.13 $Y2=1.95
cc_90 VPB N_A_137_260#_c_182_n 0.00417182f $X=-0.19 $Y=1.66 $X2=3.32 $Y2=2.115
cc_91 VPB N_D1_c_341_n 0.0107116f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_92 VPB N_D1_c_347_n 0.0238409f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_93 VPB N_D1_c_343_n 0.0061435f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_94 VPB N_D1_c_349_n 0.0209442f $X=-0.19 $Y=1.66 $X2=0.775 $Y2=1.765
cc_95 VPB N_D1_c_344_n 0.00444206f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_96 VPB N_C1_c_413_n 0.0148234f $X=-0.19 $Y=1.66 $X2=3.17 $Y2=1.96
cc_97 VPB N_C1_c_414_n 0.0186803f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_98 VPB C1 0.00729324f $X=-0.19 $Y=1.66 $X2=1.225 $Y2=2.4
cc_99 VPB N_C1_c_412_n 0.0412126f $X=-0.19 $Y=1.66 $X2=1.675 $Y2=2.4
cc_100 VPB N_B1_c_479_n 0.0186946f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_101 VPB N_B1_c_480_n 0.014858f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_102 VPB B1 0.00430243f $X=-0.19 $Y=1.66 $X2=0.775 $Y2=1.765
cc_103 VPB N_B1_c_478_n 0.0360462f $X=-0.19 $Y=1.66 $X2=1.225 $Y2=2.4
cc_104 VPB N_A1_c_534_n 0.0152696f $X=-0.19 $Y=1.66 $X2=3.125 $Y2=0.37
cc_105 VPB N_A1_c_535_n 0.0152986f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_106 VPB A1 0.00274353f $X=-0.19 $Y=1.66 $X2=0.775 $Y2=1.765
cc_107 VPB N_A1_c_533_n 0.0319515f $X=-0.19 $Y=1.66 $X2=1.285 $Y2=0.74
cc_108 VPB N_A2_c_584_n 0.00681858f $X=-0.19 $Y=1.66 $X2=3.995 $Y2=0.37
cc_109 VPB N_A2_c_591_n 0.0209975f $X=-0.19 $Y=1.66 $X2=4.865 $Y2=0.37
cc_110 VPB N_A2_c_586_n 0.00847249f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_111 VPB N_A2_c_593_n 0.0291968f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_112 VPB A2 0.0104325f $X=-0.19 $Y=1.66 $X2=1.225 $Y2=2.4
cc_113 VPB N_VPWR_c_634_n 0.0434034f $X=-0.19 $Y=1.66 $X2=0.775 $Y2=2.4
cc_114 VPB N_VPWR_c_635_n 0.00799266f $X=-0.19 $Y=1.66 $X2=1.285 $Y2=1.3
cc_115 VPB N_VPWR_c_636_n 0.0229489f $X=-0.19 $Y=1.66 $X2=1.675 $Y2=1.765
cc_116 VPB N_VPWR_c_637_n 0.00329129f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_117 VPB N_VPWR_c_638_n 0.00504372f $X=-0.19 $Y=1.66 $X2=2.145 $Y2=1.3
cc_118 VPB N_VPWR_c_639_n 0.0143948f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_119 VPB N_VPWR_c_640_n 0.0047828f $X=-0.19 $Y=1.66 $X2=2.575 $Y2=1.3
cc_120 VPB N_VPWR_c_641_n 0.0206041f $X=-0.19 $Y=1.66 $X2=2.575 $Y2=0.74
cc_121 VPB N_VPWR_c_642_n 0.00324402f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_122 VPB N_VPWR_c_643_n 0.0206041f $X=-0.19 $Y=1.66 $X2=1.035 $Y2=1.465
cc_123 VPB N_VPWR_c_644_n 0.0047828f $X=-0.19 $Y=1.66 $X2=1.035 $Y2=1.465
cc_124 VPB N_VPWR_c_645_n 0.0909002f $X=-0.19 $Y=1.66 $X2=3.13 $Y2=1.95
cc_125 VPB N_VPWR_c_646_n 0.0164337f $X=-0.19 $Y=1.66 $X2=4.135 $Y2=0.515
cc_126 VPB N_VPWR_c_647_n 0.0197879f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_127 VPB N_VPWR_c_633_n 0.11901f $X=-0.19 $Y=1.66 $X2=6.51 $Y2=1.195
cc_128 VPB N_VPWR_c_649_n 0.00601644f $X=-0.19 $Y=1.66 $X2=6.64 $Y2=0.79
cc_129 VPB N_VPWR_c_650_n 0.00460249f $X=-0.19 $Y=1.66 $X2=3.197 $Y2=1.005
cc_130 VPB N_X_c_741_n 6.45555e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_131 VPB N_X_c_742_n 0.0199052f $X=-0.19 $Y=1.66 $X2=0.775 $Y2=1.765
cc_132 VPB N_X_c_743_n 0.00257348f $X=-0.19 $Y=1.66 $X2=1.225 $Y2=1.765
cc_133 VPB N_X_c_744_n 0.00363002f $X=-0.19 $Y=1.66 $X2=1.285 $Y2=0.74
cc_134 VPB N_X_c_745_n 0.00257348f $X=-0.19 $Y=1.66 $X2=2.125 $Y2=1.765
cc_135 VPB N_X_c_746_n 0.00188882f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_136 VPB X 0.00895317f $X=-0.19 $Y=1.66 $X2=1.035 $Y2=1.465
cc_137 VPB N_A_549_392#_c_812_n 0.00617724f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_138 VPB N_A_549_392#_c_813_n 0.00213603f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_139 VPB N_A_549_392#_c_814_n 0.00424137f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_140 VPB N_A_549_392#_c_815_n 0.00711978f $X=-0.19 $Y=1.66 $X2=0.775 $Y2=2.4
cc_141 VPB N_A_549_392#_c_816_n 0.00636f $X=-0.19 $Y=1.66 $X2=1.285 $Y2=1.3
cc_142 VPB N_A_549_392#_c_817_n 0.00587218f $X=-0.19 $Y=1.66 $X2=1.675 $Y2=1.765
cc_143 VPB N_A_549_392#_c_818_n 0.0021839f $X=-0.19 $Y=1.66 $X2=1.675 $Y2=2.4
cc_144 VPB N_A_814_392#_c_860_n 0.017897f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_145 VPB N_A_814_392#_c_861_n 0.00109997f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_146 VPB N_A_814_392#_c_862_n 0.00183558f $X=-0.19 $Y=1.66 $X2=0.775 $Y2=1.765
cc_147 VPB N_A_1013_392#_c_890_n 0.00585892f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_148 VPB N_A_1013_392#_c_891_n 0.00502224f $X=-0.19 $Y=1.66 $X2=0.775 $Y2=2.4
cc_149 VPB N_A_1013_392#_c_892_n 0.00398437f $X=-0.19 $Y=1.66 $X2=0.775 $Y2=2.4
cc_150 VPB N_A_1013_392#_c_893_n 0.00213609f $X=-0.19 $Y=1.66 $X2=1.225
+ $Y2=1.765
cc_151 VPB N_A_1013_392#_c_894_n 0.00319618f $X=-0.19 $Y=1.66 $X2=1.285 $Y2=0.74
cc_152 VPB N_A_1013_392#_c_895_n 0.00180921f $X=-0.19 $Y=1.66 $X2=1.675 $Y2=2.4
cc_153 VPB N_A_1013_392#_c_896_n 0.00424615f $X=-0.19 $Y=1.66 $X2=1.715 $Y2=1.3
cc_154 VPB N_A_1013_392#_c_897_n 0.0107381f $X=-0.19 $Y=1.66 $X2=1.715 $Y2=0.74
cc_155 VPB N_A_1013_392#_c_898_n 0.0360166f $X=-0.19 $Y=1.66 $X2=2.125 $Y2=1.765
cc_156 VPB N_A_1013_392#_c_899_n 0.00159638f $X=-0.19 $Y=1.66 $X2=2.145 $Y2=0.74
cc_157 N_A_137_260#_M1025_g N_D1_M1017_g 0.00920717f $X=2.575 $Y=0.74 $X2=0
+ $Y2=0
cc_158 N_A_137_260#_c_164_n N_D1_M1017_g 0.0088411f $X=3.265 $Y=0.515 $X2=0
+ $Y2=0
cc_159 N_A_137_260#_c_165_n N_D1_M1017_g 0.00468003f $X=3.13 $Y=1.3 $X2=0 $Y2=0
cc_160 N_A_137_260#_c_172_n N_D1_M1017_g 0.00383016f $X=3.197 $Y=1.005 $X2=0
+ $Y2=0
cc_161 N_A_137_260#_c_162_n N_D1_c_341_n 0.00190569f $X=3.045 $Y=1.465 $X2=0
+ $Y2=0
cc_162 N_A_137_260#_c_181_n N_D1_c_341_n 0.00875445f $X=3.13 $Y=1.95 $X2=0 $Y2=0
cc_163 N_A_137_260#_c_173_n N_D1_c_341_n 6.56895e-19 $X=3.13 $Y=1.465 $X2=0
+ $Y2=0
cc_164 N_A_137_260#_c_181_n N_D1_c_347_n 0.0060183f $X=3.13 $Y=1.95 $X2=0 $Y2=0
cc_165 N_A_137_260#_c_182_n N_D1_c_347_n 0.0154255f $X=3.32 $Y=2.115 $X2=0 $Y2=0
cc_166 N_A_137_260#_c_165_n N_D1_M1022_g 0.00341074f $X=3.13 $Y=1.3 $X2=0 $Y2=0
cc_167 N_A_137_260#_c_166_n N_D1_M1022_g 0.013218f $X=4.05 $Y=1.005 $X2=0 $Y2=0
cc_168 N_A_137_260#_c_181_n N_D1_c_343_n 0.00238825f $X=3.13 $Y=1.95 $X2=0 $Y2=0
cc_169 N_A_137_260#_c_181_n N_D1_c_349_n 0.0012221f $X=3.13 $Y=1.95 $X2=0 $Y2=0
cc_170 N_A_137_260#_c_182_n N_D1_c_349_n 0.00289319f $X=3.32 $Y=2.115 $X2=0
+ $Y2=0
cc_171 N_A_137_260#_c_165_n N_D1_c_344_n 0.00282261f $X=3.13 $Y=1.3 $X2=0 $Y2=0
cc_172 N_A_137_260#_c_181_n N_D1_c_344_n 0.0118515f $X=3.13 $Y=1.95 $X2=0 $Y2=0
cc_173 N_A_137_260#_c_166_n N_D1_c_344_n 0.0254454f $X=4.05 $Y=1.005 $X2=0 $Y2=0
cc_174 N_A_137_260#_c_173_n N_D1_c_344_n 0.0266866f $X=3.13 $Y=1.465 $X2=0 $Y2=0
cc_175 N_A_137_260#_c_182_n N_D1_c_344_n 0.00156971f $X=3.32 $Y=2.115 $X2=0
+ $Y2=0
cc_176 N_A_137_260#_c_174_n N_D1_c_344_n 9.88457e-19 $X=4.135 $Y=1.005 $X2=0
+ $Y2=0
cc_177 N_A_137_260#_c_162_n N_D1_c_345_n 0.00928659f $X=3.045 $Y=1.465 $X2=0
+ $Y2=0
cc_178 N_A_137_260#_c_163_n N_D1_c_345_n 0.0165426f $X=2.485 $Y=1.465 $X2=0
+ $Y2=0
cc_179 N_A_137_260#_c_165_n N_D1_c_345_n 0.00170063f $X=3.13 $Y=1.3 $X2=0 $Y2=0
cc_180 N_A_137_260#_c_166_n N_D1_c_345_n 5.5668e-19 $X=4.05 $Y=1.005 $X2=0 $Y2=0
cc_181 N_A_137_260#_c_172_n N_D1_c_345_n 0.00468078f $X=3.197 $Y=1.005 $X2=0
+ $Y2=0
cc_182 N_A_137_260#_c_173_n N_D1_c_345_n 0.00872384f $X=3.13 $Y=1.465 $X2=0
+ $Y2=0
cc_183 N_A_137_260#_c_182_n N_D1_c_345_n 0.00292383f $X=3.32 $Y=2.115 $X2=0
+ $Y2=0
cc_184 N_A_137_260#_c_166_n N_C1_M1006_g 0.016344f $X=4.05 $Y=1.005 $X2=0 $Y2=0
cc_185 N_A_137_260#_c_174_n N_C1_M1006_g 0.00443494f $X=4.135 $Y=1.005 $X2=0
+ $Y2=0
cc_186 N_A_137_260#_c_168_n N_C1_c_408_n 0.00385041f $X=4.92 $Y=1.195 $X2=0
+ $Y2=0
cc_187 N_A_137_260#_c_167_n N_C1_c_409_n 0.00126475f $X=4.135 $Y=0.515 $X2=0
+ $Y2=0
cc_188 N_A_137_260#_c_168_n N_C1_c_410_n 0.0102868f $X=4.92 $Y=1.195 $X2=0 $Y2=0
cc_189 N_A_137_260#_c_174_n N_C1_c_410_n 0.00150966f $X=4.135 $Y=1.005 $X2=0
+ $Y2=0
cc_190 N_A_137_260#_c_166_n C1 0.00353585f $X=4.05 $Y=1.005 $X2=0 $Y2=0
cc_191 N_A_137_260#_c_168_n C1 0.0532268f $X=4.92 $Y=1.195 $X2=0 $Y2=0
cc_192 N_A_137_260#_c_170_n C1 0.00511502f $X=6.51 $Y=1.195 $X2=0 $Y2=0
cc_193 N_A_137_260#_c_174_n C1 0.014169f $X=4.135 $Y=1.005 $X2=0 $Y2=0
cc_194 N_A_137_260#_c_175_n C1 0.0150362f $X=5.005 $Y=1.195 $X2=0 $Y2=0
cc_195 N_A_137_260#_c_168_n N_C1_c_412_n 0.00435093f $X=4.92 $Y=1.195 $X2=0
+ $Y2=0
cc_196 N_A_137_260#_c_174_n N_C1_c_412_n 0.00279548f $X=4.135 $Y=1.005 $X2=0
+ $Y2=0
cc_197 N_A_137_260#_c_169_n N_B1_c_473_n 0.00202516f $X=5.005 $Y=0.515 $X2=-0.19
+ $Y2=-0.245
cc_198 N_A_137_260#_c_168_n N_B1_c_474_n 0.00376958f $X=4.92 $Y=1.195 $X2=0
+ $Y2=0
cc_199 N_A_137_260#_c_169_n N_B1_c_474_n 0.00385868f $X=5.005 $Y=0.515 $X2=0
+ $Y2=0
cc_200 N_A_137_260#_c_170_n N_B1_c_474_n 0.00376958f $X=6.51 $Y=1.195 $X2=0
+ $Y2=0
cc_201 N_A_137_260#_c_175_n N_B1_c_474_n 0.00459246f $X=5.005 $Y=1.195 $X2=0
+ $Y2=0
cc_202 N_A_137_260#_c_168_n N_B1_c_475_n 0.0114299f $X=4.92 $Y=1.195 $X2=0 $Y2=0
cc_203 N_A_137_260#_c_169_n N_B1_c_476_n 0.00202516f $X=5.005 $Y=0.515 $X2=0
+ $Y2=0
cc_204 N_A_137_260#_c_170_n B1 0.0521988f $X=6.51 $Y=1.195 $X2=0 $Y2=0
cc_205 N_A_137_260#_c_170_n N_B1_c_478_n 0.0468085f $X=6.51 $Y=1.195 $X2=0 $Y2=0
cc_206 N_A_137_260#_c_170_n N_A1_M1001_g 0.0128558f $X=6.51 $Y=1.195 $X2=0 $Y2=0
cc_207 N_A_137_260#_c_171_n N_A1_M1001_g 0.00268505f $X=6.605 $Y=0.79 $X2=0
+ $Y2=0
cc_208 N_A_137_260#_c_170_n N_A1_M1019_g 0.00567167f $X=6.51 $Y=1.195 $X2=0
+ $Y2=0
cc_209 N_A_137_260#_c_171_n N_A1_M1019_g 0.00661126f $X=6.605 $Y=0.79 $X2=0
+ $Y2=0
cc_210 N_A_137_260#_c_170_n A1 0.0380613f $X=6.51 $Y=1.195 $X2=0 $Y2=0
cc_211 N_A_137_260#_c_170_n N_A1_c_533_n 0.0049516f $X=6.51 $Y=1.195 $X2=0 $Y2=0
cc_212 N_A_137_260#_c_170_n N_A2_M1009_g 7.22688e-19 $X=6.51 $Y=1.195 $X2=0
+ $Y2=0
cc_213 N_A_137_260#_c_170_n A2 6.93463e-19 $X=6.51 $Y=1.195 $X2=0 $Y2=0
cc_214 N_A_137_260#_c_176_n N_VPWR_c_634_n 0.00993564f $X=0.775 $Y=1.765 $X2=0
+ $Y2=0
cc_215 N_A_137_260#_c_177_n N_VPWR_c_635_n 0.00586501f $X=1.225 $Y=1.765 $X2=0
+ $Y2=0
cc_216 N_A_137_260#_c_178_n N_VPWR_c_635_n 0.00586501f $X=1.675 $Y=1.765 $X2=0
+ $Y2=0
cc_217 N_A_137_260#_c_179_n N_VPWR_c_636_n 0.0100892f $X=2.125 $Y=1.765 $X2=0
+ $Y2=0
cc_218 N_A_137_260#_c_162_n N_VPWR_c_636_n 0.0192372f $X=3.045 $Y=1.465 $X2=0
+ $Y2=0
cc_219 N_A_137_260#_c_163_n N_VPWR_c_636_n 0.00629085f $X=2.485 $Y=1.465 $X2=0
+ $Y2=0
cc_220 N_A_137_260#_c_181_n N_VPWR_c_636_n 0.00408142f $X=3.13 $Y=1.95 $X2=0
+ $Y2=0
cc_221 N_A_137_260#_c_182_n N_VPWR_c_636_n 0.00557626f $X=3.32 $Y=2.115 $X2=0
+ $Y2=0
cc_222 N_A_137_260#_c_176_n N_VPWR_c_641_n 0.00445602f $X=0.775 $Y=1.765 $X2=0
+ $Y2=0
cc_223 N_A_137_260#_c_177_n N_VPWR_c_641_n 0.00445602f $X=1.225 $Y=1.765 $X2=0
+ $Y2=0
cc_224 N_A_137_260#_c_178_n N_VPWR_c_643_n 0.00445602f $X=1.675 $Y=1.765 $X2=0
+ $Y2=0
cc_225 N_A_137_260#_c_179_n N_VPWR_c_643_n 0.00445602f $X=2.125 $Y=1.765 $X2=0
+ $Y2=0
cc_226 N_A_137_260#_c_176_n N_VPWR_c_633_n 0.00861697f $X=0.775 $Y=1.765 $X2=0
+ $Y2=0
cc_227 N_A_137_260#_c_177_n N_VPWR_c_633_n 0.00857589f $X=1.225 $Y=1.765 $X2=0
+ $Y2=0
cc_228 N_A_137_260#_c_178_n N_VPWR_c_633_n 0.00857589f $X=1.675 $Y=1.765 $X2=0
+ $Y2=0
cc_229 N_A_137_260#_c_179_n N_VPWR_c_633_n 0.00862391f $X=2.125 $Y=1.765 $X2=0
+ $Y2=0
cc_230 N_A_137_260#_M1005_g N_X_c_734_n 0.0145305f $X=1.285 $Y=0.74 $X2=0 $Y2=0
cc_231 N_A_137_260#_c_162_n N_X_c_734_n 0.040362f $X=3.045 $Y=1.465 $X2=0 $Y2=0
cc_232 N_A_137_260#_c_163_n N_X_c_734_n 0.013583f $X=2.485 $Y=1.465 $X2=0 $Y2=0
cc_233 N_A_137_260#_c_176_n N_X_c_741_n 0.0154002f $X=0.775 $Y=1.765 $X2=0 $Y2=0
cc_234 N_A_137_260#_c_163_n N_X_c_741_n 5.17675e-19 $X=2.485 $Y=1.465 $X2=0
+ $Y2=0
cc_235 N_A_137_260#_c_176_n N_X_c_743_n 0.017229f $X=0.775 $Y=1.765 $X2=0 $Y2=0
cc_236 N_A_137_260#_c_177_n N_X_c_743_n 0.0125029f $X=1.225 $Y=1.765 $X2=0 $Y2=0
cc_237 N_A_137_260#_c_178_n N_X_c_743_n 6.9119e-19 $X=1.675 $Y=1.765 $X2=0 $Y2=0
cc_238 N_A_137_260#_c_177_n N_X_c_744_n 0.0120074f $X=1.225 $Y=1.765 $X2=0 $Y2=0
cc_239 N_A_137_260#_c_178_n N_X_c_744_n 0.0129464f $X=1.675 $Y=1.765 $X2=0 $Y2=0
cc_240 N_A_137_260#_c_179_n N_X_c_744_n 0.00325815f $X=2.125 $Y=1.765 $X2=0
+ $Y2=0
cc_241 N_A_137_260#_c_162_n N_X_c_744_n 0.0694546f $X=3.045 $Y=1.465 $X2=0 $Y2=0
cc_242 N_A_137_260#_c_163_n N_X_c_744_n 0.0155728f $X=2.485 $Y=1.465 $X2=0 $Y2=0
cc_243 N_A_137_260#_M1005_g N_X_c_736_n 3.97481e-19 $X=1.285 $Y=0.74 $X2=0 $Y2=0
cc_244 N_A_137_260#_M1016_g N_X_c_736_n 0.00845522f $X=1.715 $Y=0.74 $X2=0 $Y2=0
cc_245 N_A_137_260#_M1021_g N_X_c_736_n 5.68006e-19 $X=2.145 $Y=0.74 $X2=0 $Y2=0
cc_246 N_A_137_260#_M1016_g N_X_c_737_n 0.0111034f $X=1.715 $Y=0.74 $X2=0 $Y2=0
cc_247 N_A_137_260#_M1021_g N_X_c_737_n 0.0120709f $X=2.145 $Y=0.74 $X2=0 $Y2=0
cc_248 N_A_137_260#_M1025_g N_X_c_737_n 2.99675e-19 $X=2.575 $Y=0.74 $X2=0 $Y2=0
cc_249 N_A_137_260#_c_162_n N_X_c_737_n 0.0598052f $X=3.045 $Y=1.465 $X2=0 $Y2=0
cc_250 N_A_137_260#_c_163_n N_X_c_737_n 0.00457162f $X=2.485 $Y=1.465 $X2=0
+ $Y2=0
cc_251 N_A_137_260#_c_165_n N_X_c_737_n 8.27816e-19 $X=3.13 $Y=1.3 $X2=0 $Y2=0
cc_252 N_A_137_260#_c_177_n N_X_c_745_n 6.9119e-19 $X=1.225 $Y=1.765 $X2=0 $Y2=0
cc_253 N_A_137_260#_c_178_n N_X_c_745_n 0.0125029f $X=1.675 $Y=1.765 $X2=0 $Y2=0
cc_254 N_A_137_260#_c_179_n N_X_c_745_n 0.0118573f $X=2.125 $Y=1.765 $X2=0 $Y2=0
cc_255 N_A_137_260#_M1016_g N_X_c_738_n 5.68006e-19 $X=1.715 $Y=0.74 $X2=0 $Y2=0
cc_256 N_A_137_260#_M1021_g N_X_c_738_n 0.00845522f $X=2.145 $Y=0.74 $X2=0 $Y2=0
cc_257 N_A_137_260#_M1025_g N_X_c_738_n 3.97481e-19 $X=2.575 $Y=0.74 $X2=0 $Y2=0
cc_258 N_A_137_260#_c_176_n N_X_c_746_n 0.00110979f $X=0.775 $Y=1.765 $X2=0
+ $Y2=0
cc_259 N_A_137_260#_c_177_n N_X_c_746_n 9.3899e-19 $X=1.225 $Y=1.765 $X2=0 $Y2=0
cc_260 N_A_137_260#_c_162_n N_X_c_746_n 0.0248105f $X=3.045 $Y=1.465 $X2=0 $Y2=0
cc_261 N_A_137_260#_c_163_n N_X_c_746_n 0.00733767f $X=2.485 $Y=1.465 $X2=0
+ $Y2=0
cc_262 N_A_137_260#_M1016_g N_X_c_739_n 9.7541e-19 $X=1.715 $Y=0.74 $X2=0 $Y2=0
cc_263 N_A_137_260#_c_162_n N_X_c_739_n 0.0209731f $X=3.045 $Y=1.465 $X2=0 $Y2=0
cc_264 N_A_137_260#_c_163_n N_X_c_739_n 0.00232957f $X=2.485 $Y=1.465 $X2=0
+ $Y2=0
cc_265 N_A_137_260#_c_176_n X 0.0015256f $X=0.775 $Y=1.765 $X2=0 $Y2=0
cc_266 N_A_137_260#_M1005_g X 0.00443048f $X=1.285 $Y=0.74 $X2=0 $Y2=0
cc_267 N_A_137_260#_c_162_n X 0.0234845f $X=3.045 $Y=1.465 $X2=0 $Y2=0
cc_268 N_A_137_260#_c_163_n X 0.0171147f $X=2.485 $Y=1.465 $X2=0 $Y2=0
cc_269 N_A_137_260#_c_162_n N_A_549_392#_c_812_n 0.00958133f $X=3.045 $Y=1.465
+ $X2=0 $Y2=0
cc_270 N_A_137_260#_c_182_n N_A_549_392#_c_812_n 0.0289859f $X=3.32 $Y=2.115
+ $X2=0 $Y2=0
cc_271 N_A_137_260#_M1010_d N_A_549_392#_c_813_n 0.00243452f $X=3.17 $Y=1.96
+ $X2=0 $Y2=0
cc_272 N_A_137_260#_c_182_n N_A_549_392#_c_813_n 0.0126885f $X=3.32 $Y=2.115
+ $X2=0 $Y2=0
cc_273 N_A_137_260#_c_182_n N_A_549_392#_c_815_n 0.0517083f $X=3.32 $Y=2.115
+ $X2=0 $Y2=0
cc_274 N_A_137_260#_c_170_n N_A_814_392#_c_860_n 0.00668474f $X=6.51 $Y=1.195
+ $X2=0 $Y2=0
cc_275 N_A_137_260#_c_170_n N_A_1013_392#_c_893_n 0.00193826f $X=6.51 $Y=1.195
+ $X2=0 $Y2=0
cc_276 N_A_137_260#_c_170_n N_A_1013_392#_c_894_n 0.00297895f $X=6.51 $Y=1.195
+ $X2=0 $Y2=0
cc_277 N_A_137_260#_c_166_n N_VGND_M1022_s 0.00187091f $X=4.05 $Y=1.005 $X2=0
+ $Y2=0
cc_278 N_A_137_260#_M1005_g N_VGND_c_948_n 0.0112604f $X=1.285 $Y=0.74 $X2=0
+ $Y2=0
cc_279 N_A_137_260#_M1016_g N_VGND_c_948_n 5.04273e-19 $X=1.715 $Y=0.74 $X2=0
+ $Y2=0
cc_280 N_A_137_260#_M1016_g N_VGND_c_949_n 0.0017512f $X=1.715 $Y=0.74 $X2=0
+ $Y2=0
cc_281 N_A_137_260#_M1021_g N_VGND_c_949_n 0.0017512f $X=2.145 $Y=0.74 $X2=0
+ $Y2=0
cc_282 N_A_137_260#_M1021_g N_VGND_c_950_n 0.00434272f $X=2.145 $Y=0.74 $X2=0
+ $Y2=0
cc_283 N_A_137_260#_M1025_g N_VGND_c_950_n 0.00383152f $X=2.575 $Y=0.74 $X2=0
+ $Y2=0
cc_284 N_A_137_260#_M1021_g N_VGND_c_951_n 5.77606e-19 $X=2.145 $Y=0.74 $X2=0
+ $Y2=0
cc_285 N_A_137_260#_M1025_g N_VGND_c_951_n 0.0112827f $X=2.575 $Y=0.74 $X2=0
+ $Y2=0
cc_286 N_A_137_260#_c_162_n N_VGND_c_951_n 0.0133944f $X=3.045 $Y=1.465 $X2=0
+ $Y2=0
cc_287 N_A_137_260#_c_164_n N_VGND_c_951_n 0.0430526f $X=3.265 $Y=0.515 $X2=0
+ $Y2=0
cc_288 N_A_137_260#_c_172_n N_VGND_c_951_n 0.0088844f $X=3.197 $Y=1.005 $X2=0
+ $Y2=0
cc_289 N_A_137_260#_c_164_n N_VGND_c_952_n 0.013284f $X=3.265 $Y=0.515 $X2=0
+ $Y2=0
cc_290 N_A_137_260#_c_164_n N_VGND_c_953_n 0.0151524f $X=3.265 $Y=0.515 $X2=0
+ $Y2=0
cc_291 N_A_137_260#_c_166_n N_VGND_c_953_n 0.0179755f $X=4.05 $Y=1.005 $X2=0
+ $Y2=0
cc_292 N_A_137_260#_c_167_n N_VGND_c_953_n 0.0150888f $X=4.135 $Y=0.515 $X2=0
+ $Y2=0
cc_293 N_A_137_260#_c_167_n N_VGND_c_954_n 0.0219298f $X=4.135 $Y=0.515 $X2=0
+ $Y2=0
cc_294 N_A_137_260#_c_168_n N_VGND_c_954_n 0.0223605f $X=4.92 $Y=1.195 $X2=0
+ $Y2=0
cc_295 N_A_137_260#_c_169_n N_VGND_c_954_n 0.0219298f $X=5.005 $Y=0.515 $X2=0
+ $Y2=0
cc_296 N_A_137_260#_c_169_n N_VGND_c_955_n 0.0218329f $X=5.005 $Y=0.515 $X2=0
+ $Y2=0
cc_297 N_A_137_260#_c_170_n N_VGND_c_955_n 0.0232912f $X=6.51 $Y=1.195 $X2=0
+ $Y2=0
cc_298 N_A_137_260#_M1005_g N_VGND_c_959_n 0.00383152f $X=1.285 $Y=0.74 $X2=0
+ $Y2=0
cc_299 N_A_137_260#_M1016_g N_VGND_c_959_n 0.00434272f $X=1.715 $Y=0.74 $X2=0
+ $Y2=0
cc_300 N_A_137_260#_c_167_n N_VGND_c_961_n 0.00749631f $X=4.135 $Y=0.515 $X2=0
+ $Y2=0
cc_301 N_A_137_260#_c_169_n N_VGND_c_962_n 0.00749631f $X=5.005 $Y=0.515 $X2=0
+ $Y2=0
cc_302 N_A_137_260#_M1005_g N_VGND_c_965_n 0.0075754f $X=1.285 $Y=0.74 $X2=0
+ $Y2=0
cc_303 N_A_137_260#_M1016_g N_VGND_c_965_n 0.00820284f $X=1.715 $Y=0.74 $X2=0
+ $Y2=0
cc_304 N_A_137_260#_M1021_g N_VGND_c_965_n 0.00820284f $X=2.145 $Y=0.74 $X2=0
+ $Y2=0
cc_305 N_A_137_260#_M1025_g N_VGND_c_965_n 0.0075754f $X=2.575 $Y=0.74 $X2=0
+ $Y2=0
cc_306 N_A_137_260#_c_164_n N_VGND_c_965_n 0.0108098f $X=3.265 $Y=0.515 $X2=0
+ $Y2=0
cc_307 N_A_137_260#_c_167_n N_VGND_c_965_n 0.0062048f $X=4.135 $Y=0.515 $X2=0
+ $Y2=0
cc_308 N_A_137_260#_c_169_n N_VGND_c_965_n 0.0062048f $X=5.005 $Y=0.515 $X2=0
+ $Y2=0
cc_309 N_A_137_260#_c_170_n N_A_1210_74#_c_1062_n 0.0243671f $X=6.51 $Y=1.195
+ $X2=0 $Y2=0
cc_310 N_A_137_260#_M1001_d N_A_1210_74#_c_1063_n 0.00176461f $X=6.465 $Y=0.37
+ $X2=0 $Y2=0
cc_311 N_A_137_260#_c_170_n N_A_1210_74#_c_1063_n 0.00338623f $X=6.51 $Y=1.195
+ $X2=0 $Y2=0
cc_312 N_A_137_260#_c_171_n N_A_1210_74#_c_1063_n 0.0143564f $X=6.605 $Y=0.79
+ $X2=0 $Y2=0
cc_313 N_A_137_260#_c_171_n N_A_1210_74#_c_1066_n 0.0094371f $X=6.605 $Y=0.79
+ $X2=0 $Y2=0
cc_314 N_D1_M1022_g N_C1_M1006_g 0.026984f $X=3.48 $Y=0.69 $X2=0 $Y2=0
cc_315 N_D1_c_344_n N_C1_M1006_g 0.00541691f $X=3.47 $Y=1.425 $X2=0 $Y2=0
cc_316 N_D1_c_345_n N_C1_M1006_g 0.0105371f $X=3.48 $Y=1.425 $X2=0 $Y2=0
cc_317 N_D1_c_349_n N_C1_c_413_n 0.00891721f $X=3.545 $Y=1.885 $X2=0 $Y2=0
cc_318 N_D1_c_344_n C1 0.0205928f $X=3.47 $Y=1.425 $X2=0 $Y2=0
cc_319 N_D1_c_345_n C1 3.19228e-19 $X=3.48 $Y=1.425 $X2=0 $Y2=0
cc_320 N_D1_c_343_n N_C1_c_412_n 0.0245077f $X=3.545 $Y=1.795 $X2=0 $Y2=0
cc_321 N_D1_c_344_n N_C1_c_412_n 0.00144306f $X=3.47 $Y=1.425 $X2=0 $Y2=0
cc_322 N_D1_c_347_n N_VPWR_c_636_n 0.0103599f $X=3.095 $Y=1.885 $X2=0 $Y2=0
cc_323 N_D1_c_347_n N_VPWR_c_645_n 0.00278257f $X=3.095 $Y=1.885 $X2=0 $Y2=0
cc_324 N_D1_c_349_n N_VPWR_c_645_n 0.00278257f $X=3.545 $Y=1.885 $X2=0 $Y2=0
cc_325 N_D1_c_347_n N_VPWR_c_633_n 0.00358623f $X=3.095 $Y=1.885 $X2=0 $Y2=0
cc_326 N_D1_c_349_n N_VPWR_c_633_n 0.00353905f $X=3.545 $Y=1.885 $X2=0 $Y2=0
cc_327 N_D1_c_347_n N_A_549_392#_c_812_n 0.0078738f $X=3.095 $Y=1.885 $X2=0
+ $Y2=0
cc_328 N_D1_c_349_n N_A_549_392#_c_812_n 5.7112e-19 $X=3.545 $Y=1.885 $X2=0
+ $Y2=0
cc_329 N_D1_c_347_n N_A_549_392#_c_813_n 0.0108414f $X=3.095 $Y=1.885 $X2=0
+ $Y2=0
cc_330 N_D1_c_349_n N_A_549_392#_c_813_n 0.0108414f $X=3.545 $Y=1.885 $X2=0
+ $Y2=0
cc_331 N_D1_c_347_n N_A_549_392#_c_814_n 0.00262934f $X=3.095 $Y=1.885 $X2=0
+ $Y2=0
cc_332 N_D1_c_347_n N_A_549_392#_c_815_n 6.80212e-19 $X=3.095 $Y=1.885 $X2=0
+ $Y2=0
cc_333 N_D1_c_349_n N_A_549_392#_c_815_n 0.0116699f $X=3.545 $Y=1.885 $X2=0
+ $Y2=0
cc_334 N_D1_c_344_n N_A_549_392#_c_815_n 0.00972896f $X=3.47 $Y=1.425 $X2=0
+ $Y2=0
cc_335 N_D1_c_349_n N_A_549_392#_c_818_n 0.00171731f $X=3.545 $Y=1.885 $X2=0
+ $Y2=0
cc_336 N_D1_M1017_g N_VGND_c_951_n 0.0034789f $X=3.05 $Y=0.69 $X2=0 $Y2=0
cc_337 N_D1_M1017_g N_VGND_c_952_n 0.00371957f $X=3.05 $Y=0.69 $X2=0 $Y2=0
cc_338 N_D1_M1022_g N_VGND_c_952_n 0.00383152f $X=3.48 $Y=0.69 $X2=0 $Y2=0
cc_339 N_D1_M1017_g N_VGND_c_953_n 4.71027e-19 $X=3.05 $Y=0.69 $X2=0 $Y2=0
cc_340 N_D1_M1022_g N_VGND_c_953_n 0.00870112f $X=3.48 $Y=0.69 $X2=0 $Y2=0
cc_341 N_D1_M1017_g N_VGND_c_965_n 0.00619993f $X=3.05 $Y=0.69 $X2=0 $Y2=0
cc_342 N_D1_M1022_g N_VGND_c_965_n 0.0075754f $X=3.48 $Y=0.69 $X2=0 $Y2=0
cc_343 N_C1_c_409_n N_B1_c_473_n 0.00859538f $X=4.36 $Y=1.085 $X2=-0.19
+ $Y2=-0.245
cc_344 N_C1_c_410_n N_B1_c_473_n 0.00368377f $X=4.36 $Y=1.235 $X2=-0.19
+ $Y2=-0.245
cc_345 N_C1_c_408_n N_B1_c_475_n 0.00368377f $X=4.37 $Y=1.45 $X2=0 $Y2=0
cc_346 C1 N_B1_c_475_n 0.00293335f $X=4.955 $Y=1.58 $X2=0 $Y2=0
cc_347 C1 B1 0.0219368f $X=4.955 $Y=1.58 $X2=0 $Y2=0
cc_348 C1 N_B1_c_478_n 0.00464261f $X=4.955 $Y=1.58 $X2=0 $Y2=0
cc_349 N_C1_c_412_n N_B1_c_478_n 0.00337788f $X=4.445 $Y=1.667 $X2=0 $Y2=0
cc_350 N_C1_c_413_n N_VPWR_c_645_n 0.00278257f $X=3.995 $Y=1.885 $X2=0 $Y2=0
cc_351 N_C1_c_414_n N_VPWR_c_645_n 0.00278257f $X=4.445 $Y=1.885 $X2=0 $Y2=0
cc_352 N_C1_c_413_n N_VPWR_c_633_n 0.00353905f $X=3.995 $Y=1.885 $X2=0 $Y2=0
cc_353 N_C1_c_414_n N_VPWR_c_633_n 0.00358623f $X=4.445 $Y=1.885 $X2=0 $Y2=0
cc_354 N_C1_c_413_n N_A_549_392#_c_815_n 0.0117317f $X=3.995 $Y=1.885 $X2=0
+ $Y2=0
cc_355 N_C1_c_414_n N_A_549_392#_c_815_n 6.7795e-19 $X=4.445 $Y=1.885 $X2=0
+ $Y2=0
cc_356 N_C1_c_412_n N_A_549_392#_c_815_n 0.003211f $X=4.445 $Y=1.667 $X2=0 $Y2=0
cc_357 N_C1_c_413_n N_A_549_392#_c_816_n 0.0108414f $X=3.995 $Y=1.885 $X2=0
+ $Y2=0
cc_358 N_C1_c_414_n N_A_549_392#_c_816_n 0.0134708f $X=4.445 $Y=1.885 $X2=0
+ $Y2=0
cc_359 N_C1_c_413_n N_A_549_392#_c_817_n 5.7112e-19 $X=3.995 $Y=1.885 $X2=0
+ $Y2=0
cc_360 N_C1_c_414_n N_A_549_392#_c_817_n 0.00766499f $X=4.445 $Y=1.885 $X2=0
+ $Y2=0
cc_361 N_C1_c_413_n N_A_549_392#_c_818_n 0.00171731f $X=3.995 $Y=1.885 $X2=0
+ $Y2=0
cc_362 N_C1_c_414_n N_A_814_392#_c_860_n 0.0146982f $X=4.445 $Y=1.885 $X2=0
+ $Y2=0
cc_363 C1 N_A_814_392#_c_860_n 0.0654719f $X=4.955 $Y=1.58 $X2=0 $Y2=0
cc_364 N_C1_c_412_n N_A_814_392#_c_860_n 0.00418405f $X=4.445 $Y=1.667 $X2=0
+ $Y2=0
cc_365 N_C1_c_413_n N_A_814_392#_c_861_n 0.00301095f $X=3.995 $Y=1.885 $X2=0
+ $Y2=0
cc_366 N_C1_c_414_n N_A_814_392#_c_861_n 0.00497407f $X=4.445 $Y=1.885 $X2=0
+ $Y2=0
cc_367 C1 N_A_814_392#_c_861_n 0.0143367f $X=4.955 $Y=1.58 $X2=0 $Y2=0
cc_368 N_C1_c_412_n N_A_814_392#_c_861_n 0.00435468f $X=4.445 $Y=1.667 $X2=0
+ $Y2=0
cc_369 N_C1_c_414_n N_A_1013_392#_c_892_n 5.73871e-19 $X=4.445 $Y=1.885 $X2=0
+ $Y2=0
cc_370 N_C1_M1006_g N_VGND_c_953_n 0.0084935f $X=3.92 $Y=0.69 $X2=0 $Y2=0
cc_371 N_C1_c_409_n N_VGND_c_953_n 4.44652e-19 $X=4.36 $Y=1.085 $X2=0 $Y2=0
cc_372 N_C1_M1006_g N_VGND_c_954_n 4.95643e-19 $X=3.92 $Y=0.69 $X2=0 $Y2=0
cc_373 N_C1_c_409_n N_VGND_c_954_n 0.010382f $X=4.36 $Y=1.085 $X2=0 $Y2=0
cc_374 N_C1_M1006_g N_VGND_c_961_n 0.00383152f $X=3.92 $Y=0.69 $X2=0 $Y2=0
cc_375 N_C1_c_409_n N_VGND_c_961_n 0.00383152f $X=4.36 $Y=1.085 $X2=0 $Y2=0
cc_376 N_C1_M1006_g N_VGND_c_965_n 0.0075754f $X=3.92 $Y=0.69 $X2=0 $Y2=0
cc_377 N_C1_c_409_n N_VGND_c_965_n 0.0075754f $X=4.36 $Y=1.085 $X2=0 $Y2=0
cc_378 N_B1_c_480_n N_A1_c_534_n 0.00827175f $X=5.865 $Y=1.885 $X2=-0.19
+ $Y2=-0.245
cc_379 N_B1_c_478_n N_A1_M1001_g 0.0128102f $X=5.57 $Y=1.615 $X2=0 $Y2=0
cc_380 B1 A1 0.0293403f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_381 N_B1_c_478_n A1 2.76139e-19 $X=5.57 $Y=1.615 $X2=0 $Y2=0
cc_382 B1 N_A1_c_533_n 0.00295361f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_383 N_B1_c_478_n N_A1_c_533_n 0.0188925f $X=5.57 $Y=1.615 $X2=0 $Y2=0
cc_384 N_B1_c_479_n N_VPWR_c_645_n 0.00278271f $X=5.415 $Y=1.885 $X2=0 $Y2=0
cc_385 N_B1_c_480_n N_VPWR_c_645_n 0.00278271f $X=5.865 $Y=1.885 $X2=0 $Y2=0
cc_386 N_B1_c_479_n N_VPWR_c_633_n 0.00358624f $X=5.415 $Y=1.885 $X2=0 $Y2=0
cc_387 N_B1_c_480_n N_VPWR_c_633_n 0.00353907f $X=5.865 $Y=1.885 $X2=0 $Y2=0
cc_388 N_B1_c_479_n N_A_549_392#_c_816_n 5.67935e-19 $X=5.415 $Y=1.885 $X2=0
+ $Y2=0
cc_389 N_B1_c_479_n N_A_814_392#_c_860_n 0.0149153f $X=5.415 $Y=1.885 $X2=0
+ $Y2=0
cc_390 B1 N_A_814_392#_c_860_n 0.00496499f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_391 N_B1_c_478_n N_A_814_392#_c_860_n 5.36244e-19 $X=5.57 $Y=1.615 $X2=0
+ $Y2=0
cc_392 N_B1_c_479_n N_A_814_392#_c_862_n 0.0140207f $X=5.415 $Y=1.885 $X2=0
+ $Y2=0
cc_393 N_B1_c_480_n N_A_814_392#_c_862_n 0.0101178f $X=5.865 $Y=1.885 $X2=0
+ $Y2=0
cc_394 B1 N_A_814_392#_c_862_n 0.0276944f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_395 N_B1_c_478_n N_A_814_392#_c_862_n 0.0082188f $X=5.57 $Y=1.615 $X2=0 $Y2=0
cc_396 N_B1_c_479_n N_A_1013_392#_c_891_n 0.0136535f $X=5.415 $Y=1.885 $X2=0
+ $Y2=0
cc_397 N_B1_c_480_n N_A_1013_392#_c_891_n 0.012504f $X=5.865 $Y=1.885 $X2=0
+ $Y2=0
cc_398 N_B1_c_480_n N_A_1013_392#_c_893_n 7.86054e-19 $X=5.865 $Y=1.885 $X2=0
+ $Y2=0
cc_399 B1 N_A_1013_392#_c_893_n 0.00973077f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_400 N_B1_c_473_n N_VGND_c_954_n 0.010382f $X=4.79 $Y=1.09 $X2=0 $Y2=0
cc_401 N_B1_c_476_n N_VGND_c_954_n 5.01309e-19 $X=5.22 $Y=1.09 $X2=0 $Y2=0
cc_402 N_B1_c_473_n N_VGND_c_955_n 5.01478e-19 $X=4.79 $Y=1.09 $X2=0 $Y2=0
cc_403 N_B1_c_476_n N_VGND_c_955_n 0.0114363f $X=5.22 $Y=1.09 $X2=0 $Y2=0
cc_404 N_B1_c_478_n N_VGND_c_955_n 0.00805342f $X=5.57 $Y=1.615 $X2=0 $Y2=0
cc_405 N_B1_c_473_n N_VGND_c_962_n 0.00383152f $X=4.79 $Y=1.09 $X2=0 $Y2=0
cc_406 N_B1_c_476_n N_VGND_c_962_n 0.00383152f $X=5.22 $Y=1.09 $X2=0 $Y2=0
cc_407 N_B1_c_473_n N_VGND_c_965_n 0.0075754f $X=4.79 $Y=1.09 $X2=0 $Y2=0
cc_408 N_B1_c_476_n N_VGND_c_965_n 0.0075754f $X=5.22 $Y=1.09 $X2=0 $Y2=0
cc_409 N_A1_c_533_n N_A2_c_584_n 0.0235898f $X=6.765 $Y=1.667 $X2=0 $Y2=0
cc_410 N_A1_c_535_n N_A2_c_591_n 0.00827302f $X=6.765 $Y=1.885 $X2=0 $Y2=0
cc_411 N_A1_M1019_g N_A2_M1009_g 0.0164018f $X=6.82 $Y=0.69 $X2=0 $Y2=0
cc_412 N_A1_M1019_g A2 9.03234e-19 $X=6.82 $Y=0.69 $X2=0 $Y2=0
cc_413 A1 A2 0.0291962f $X=6.875 $Y=1.58 $X2=0 $Y2=0
cc_414 N_A1_c_533_n A2 2.41572e-19 $X=6.765 $Y=1.667 $X2=0 $Y2=0
cc_415 N_A1_M1019_g N_A2_c_589_n 0.010226f $X=6.82 $Y=0.69 $X2=0 $Y2=0
cc_416 A1 N_A2_c_589_n 0.0027659f $X=6.875 $Y=1.58 $X2=0 $Y2=0
cc_417 N_A1_c_534_n N_VPWR_c_637_n 0.0106654f $X=6.315 $Y=1.885 $X2=0 $Y2=0
cc_418 N_A1_c_535_n N_VPWR_c_637_n 0.0113455f $X=6.765 $Y=1.885 $X2=0 $Y2=0
cc_419 N_A1_c_535_n N_VPWR_c_638_n 5.37805e-19 $X=6.765 $Y=1.885 $X2=0 $Y2=0
cc_420 N_A1_c_534_n N_VPWR_c_645_n 0.00413917f $X=6.315 $Y=1.885 $X2=0 $Y2=0
cc_421 N_A1_c_535_n N_VPWR_c_646_n 0.00413917f $X=6.765 $Y=1.885 $X2=0 $Y2=0
cc_422 N_A1_c_534_n N_VPWR_c_633_n 0.0081781f $X=6.315 $Y=1.885 $X2=0 $Y2=0
cc_423 N_A1_c_535_n N_VPWR_c_633_n 0.0081781f $X=6.765 $Y=1.885 $X2=0 $Y2=0
cc_424 N_A1_c_534_n N_A_1013_392#_c_891_n 0.00125031f $X=6.315 $Y=1.885 $X2=0
+ $Y2=0
cc_425 N_A1_c_534_n N_A_1013_392#_c_894_n 0.0133276f $X=6.315 $Y=1.885 $X2=0
+ $Y2=0
cc_426 N_A1_c_535_n N_A_1013_392#_c_894_n 0.0127476f $X=6.765 $Y=1.885 $X2=0
+ $Y2=0
cc_427 A1 N_A_1013_392#_c_894_n 0.0458106f $X=6.875 $Y=1.58 $X2=0 $Y2=0
cc_428 N_A1_c_533_n N_A_1013_392#_c_894_n 0.00873855f $X=6.765 $Y=1.667 $X2=0
+ $Y2=0
cc_429 N_A1_c_535_n N_A_1013_392#_c_895_n 0.00554978f $X=6.765 $Y=1.885 $X2=0
+ $Y2=0
cc_430 A1 N_A_1013_392#_c_899_n 0.0150385f $X=6.875 $Y=1.58 $X2=0 $Y2=0
cc_431 N_A1_M1019_g N_VGND_c_956_n 3.24085e-19 $X=6.82 $Y=0.69 $X2=0 $Y2=0
cc_432 N_A1_M1001_g N_VGND_c_963_n 0.00282582f $X=6.39 $Y=0.69 $X2=0 $Y2=0
cc_433 N_A1_M1019_g N_VGND_c_963_n 0.00282606f $X=6.82 $Y=0.69 $X2=0 $Y2=0
cc_434 N_A1_M1001_g N_VGND_c_965_n 0.00359239f $X=6.39 $Y=0.69 $X2=0 $Y2=0
cc_435 N_A1_M1019_g N_VGND_c_965_n 0.00354344f $X=6.82 $Y=0.69 $X2=0 $Y2=0
cc_436 N_A1_M1001_g N_A_1210_74#_c_1062_n 0.00667566f $X=6.39 $Y=0.69 $X2=0
+ $Y2=0
cc_437 N_A1_M1019_g N_A_1210_74#_c_1062_n 4.5114e-19 $X=6.82 $Y=0.69 $X2=0 $Y2=0
cc_438 N_A1_M1001_g N_A_1210_74#_c_1063_n 0.00828071f $X=6.39 $Y=0.69 $X2=0
+ $Y2=0
cc_439 N_A1_M1019_g N_A_1210_74#_c_1063_n 0.0119714f $X=6.82 $Y=0.69 $X2=0 $Y2=0
cc_440 N_A1_M1001_g N_A_1210_74#_c_1064_n 0.00224648f $X=6.39 $Y=0.69 $X2=0
+ $Y2=0
cc_441 N_A1_M1019_g N_A_1210_74#_c_1066_n 6.58764e-19 $X=6.82 $Y=0.69 $X2=0
+ $Y2=0
cc_442 A1 N_A_1210_74#_c_1066_n 0.006568f $X=6.875 $Y=1.58 $X2=0 $Y2=0
cc_443 N_A2_c_591_n N_VPWR_c_637_n 5.35985e-19 $X=7.215 $Y=1.885 $X2=0 $Y2=0
cc_444 N_A2_c_591_n N_VPWR_c_638_n 0.0106464f $X=7.215 $Y=1.885 $X2=0 $Y2=0
cc_445 N_A2_c_593_n N_VPWR_c_638_n 0.00526215f $X=7.665 $Y=1.885 $X2=0 $Y2=0
cc_446 N_A2_c_591_n N_VPWR_c_646_n 0.00413917f $X=7.215 $Y=1.885 $X2=0 $Y2=0
cc_447 N_A2_c_593_n N_VPWR_c_647_n 0.00445602f $X=7.665 $Y=1.885 $X2=0 $Y2=0
cc_448 N_A2_c_591_n N_VPWR_c_633_n 0.0081781f $X=7.215 $Y=1.885 $X2=0 $Y2=0
cc_449 N_A2_c_593_n N_VPWR_c_633_n 0.0086105f $X=7.665 $Y=1.885 $X2=0 $Y2=0
cc_450 N_A2_c_591_n N_A_1013_392#_c_895_n 0.00369429f $X=7.215 $Y=1.885 $X2=0
+ $Y2=0
cc_451 N_A2_c_591_n N_A_1013_392#_c_896_n 0.0171379f $X=7.215 $Y=1.885 $X2=0
+ $Y2=0
cc_452 N_A2_c_593_n N_A_1013_392#_c_896_n 0.0124546f $X=7.665 $Y=1.885 $X2=0
+ $Y2=0
cc_453 A2 N_A_1013_392#_c_896_n 0.0378485f $X=7.835 $Y=1.58 $X2=0 $Y2=0
cc_454 N_A2_c_589_n N_A_1013_392#_c_896_n 4.03951e-19 $X=7.68 $Y=1.425 $X2=0
+ $Y2=0
cc_455 N_A2_c_593_n N_A_1013_392#_c_897_n 0.00108926f $X=7.665 $Y=1.885 $X2=0
+ $Y2=0
cc_456 A2 N_A_1013_392#_c_897_n 0.0281455f $X=7.835 $Y=1.58 $X2=0 $Y2=0
cc_457 N_A2_c_591_n N_A_1013_392#_c_898_n 6.69308e-19 $X=7.215 $Y=1.885 $X2=0
+ $Y2=0
cc_458 N_A2_c_593_n N_A_1013_392#_c_898_n 0.0106911f $X=7.665 $Y=1.885 $X2=0
+ $Y2=0
cc_459 N_A2_M1009_g N_VGND_c_956_n 0.00825457f $X=7.25 $Y=0.69 $X2=0 $Y2=0
cc_460 N_A2_M1027_g N_VGND_c_956_n 0.0116536f $X=7.68 $Y=0.69 $X2=0 $Y2=0
cc_461 N_A2_M1009_g N_VGND_c_963_n 0.00383152f $X=7.25 $Y=0.69 $X2=0 $Y2=0
cc_462 N_A2_M1027_g N_VGND_c_964_n 0.00383152f $X=7.68 $Y=0.69 $X2=0 $Y2=0
cc_463 N_A2_M1009_g N_VGND_c_965_n 0.00757637f $X=7.25 $Y=0.69 $X2=0 $Y2=0
cc_464 N_A2_M1027_g N_VGND_c_965_n 0.00761145f $X=7.68 $Y=0.69 $X2=0 $Y2=0
cc_465 N_A2_M1009_g N_A_1210_74#_c_1063_n 7.00191e-19 $X=7.25 $Y=0.69 $X2=0
+ $Y2=0
cc_466 N_A2_M1009_g N_A_1210_74#_c_1065_n 0.0151262f $X=7.25 $Y=0.69 $X2=0 $Y2=0
cc_467 N_A2_M1027_g N_A_1210_74#_c_1065_n 0.0138099f $X=7.68 $Y=0.69 $X2=0 $Y2=0
cc_468 A2 N_A_1210_74#_c_1065_n 0.0639085f $X=7.835 $Y=1.58 $X2=0 $Y2=0
cc_469 N_A2_c_589_n N_A_1210_74#_c_1065_n 0.00442405f $X=7.68 $Y=1.425 $X2=0
+ $Y2=0
cc_470 N_A2_M1027_g N_A_1210_74#_c_1067_n 4.43891e-19 $X=7.68 $Y=0.69 $X2=0
+ $Y2=0
cc_471 N_VPWR_M1008_s N_X_c_742_n 0.00340242f $X=0.425 $Y=1.84 $X2=0 $Y2=0
cc_472 N_VPWR_c_634_n N_X_c_742_n 0.022498f $X=0.55 $Y=2.305 $X2=0 $Y2=0
cc_473 N_VPWR_c_634_n N_X_c_743_n 0.0563525f $X=0.55 $Y=2.305 $X2=0 $Y2=0
cc_474 N_VPWR_c_635_n N_X_c_743_n 0.0547423f $X=1.45 $Y=2.305 $X2=0 $Y2=0
cc_475 N_VPWR_c_641_n N_X_c_743_n 0.014552f $X=1.365 $Y=3.33 $X2=0 $Y2=0
cc_476 N_VPWR_c_633_n N_X_c_743_n 0.0119791f $X=7.92 $Y=3.33 $X2=0 $Y2=0
cc_477 N_VPWR_M1011_s N_X_c_744_n 0.00247267f $X=1.3 $Y=1.84 $X2=0 $Y2=0
cc_478 N_VPWR_c_635_n N_X_c_744_n 0.0136682f $X=1.45 $Y=2.305 $X2=0 $Y2=0
cc_479 N_VPWR_c_636_n N_X_c_744_n 0.0107081f $X=2.35 $Y=1.985 $X2=0 $Y2=0
cc_480 N_VPWR_c_635_n N_X_c_745_n 0.0547423f $X=1.45 $Y=2.305 $X2=0 $Y2=0
cc_481 N_VPWR_c_636_n N_X_c_745_n 0.0677182f $X=2.35 $Y=1.985 $X2=0 $Y2=0
cc_482 N_VPWR_c_643_n N_X_c_745_n 0.014552f $X=2.265 $Y=3.33 $X2=0 $Y2=0
cc_483 N_VPWR_c_633_n N_X_c_745_n 0.0119791f $X=7.92 $Y=3.33 $X2=0 $Y2=0
cc_484 N_VPWR_c_636_n N_A_549_392#_c_812_n 0.0463434f $X=2.35 $Y=1.985 $X2=0
+ $Y2=0
cc_485 N_VPWR_c_645_n N_A_549_392#_c_813_n 0.03588f $X=6.375 $Y=3.33 $X2=0 $Y2=0
cc_486 N_VPWR_c_633_n N_A_549_392#_c_813_n 0.0201952f $X=7.92 $Y=3.33 $X2=0
+ $Y2=0
cc_487 N_VPWR_c_636_n N_A_549_392#_c_814_n 0.0136296f $X=2.35 $Y=1.985 $X2=0
+ $Y2=0
cc_488 N_VPWR_c_645_n N_A_549_392#_c_814_n 0.0236039f $X=6.375 $Y=3.33 $X2=0
+ $Y2=0
cc_489 N_VPWR_c_633_n N_A_549_392#_c_814_n 0.012761f $X=7.92 $Y=3.33 $X2=0 $Y2=0
cc_490 N_VPWR_c_645_n N_A_549_392#_c_816_n 0.0594839f $X=6.375 $Y=3.33 $X2=0
+ $Y2=0
cc_491 N_VPWR_c_633_n N_A_549_392#_c_816_n 0.0329562f $X=7.92 $Y=3.33 $X2=0
+ $Y2=0
cc_492 N_VPWR_c_645_n N_A_549_392#_c_818_n 0.0235512f $X=6.375 $Y=3.33 $X2=0
+ $Y2=0
cc_493 N_VPWR_c_633_n N_A_549_392#_c_818_n 0.0126924f $X=7.92 $Y=3.33 $X2=0
+ $Y2=0
cc_494 N_VPWR_c_637_n N_A_1013_392#_c_891_n 0.0125885f $X=6.54 $Y=2.4 $X2=0
+ $Y2=0
cc_495 N_VPWR_c_645_n N_A_1013_392#_c_891_n 0.056348f $X=6.375 $Y=3.33 $X2=0
+ $Y2=0
cc_496 N_VPWR_c_633_n N_A_1013_392#_c_891_n 0.0315544f $X=7.92 $Y=3.33 $X2=0
+ $Y2=0
cc_497 N_VPWR_c_645_n N_A_1013_392#_c_892_n 0.0200723f $X=6.375 $Y=3.33 $X2=0
+ $Y2=0
cc_498 N_VPWR_c_633_n N_A_1013_392#_c_892_n 0.0108858f $X=7.92 $Y=3.33 $X2=0
+ $Y2=0
cc_499 N_VPWR_c_637_n N_A_1013_392#_c_928_n 0.040027f $X=6.54 $Y=2.4 $X2=0 $Y2=0
cc_500 N_VPWR_M1002_d N_A_1013_392#_c_894_n 0.00197722f $X=6.39 $Y=1.96 $X2=0
+ $Y2=0
cc_501 N_VPWR_c_637_n N_A_1013_392#_c_894_n 0.0171813f $X=6.54 $Y=2.4 $X2=0
+ $Y2=0
cc_502 N_VPWR_c_637_n N_A_1013_392#_c_895_n 0.0449718f $X=6.54 $Y=2.4 $X2=0
+ $Y2=0
cc_503 N_VPWR_c_638_n N_A_1013_392#_c_895_n 0.0440249f $X=7.44 $Y=2.455 $X2=0
+ $Y2=0
cc_504 N_VPWR_c_646_n N_A_1013_392#_c_895_n 0.00749631f $X=7.275 $Y=3.33 $X2=0
+ $Y2=0
cc_505 N_VPWR_c_633_n N_A_1013_392#_c_895_n 0.0062048f $X=7.92 $Y=3.33 $X2=0
+ $Y2=0
cc_506 N_VPWR_M1004_d N_A_1013_392#_c_896_n 0.00222494f $X=7.29 $Y=1.96 $X2=0
+ $Y2=0
cc_507 N_VPWR_c_638_n N_A_1013_392#_c_896_n 0.0154248f $X=7.44 $Y=2.455 $X2=0
+ $Y2=0
cc_508 N_VPWR_c_638_n N_A_1013_392#_c_898_n 0.0462948f $X=7.44 $Y=2.455 $X2=0
+ $Y2=0
cc_509 N_VPWR_c_647_n N_A_1013_392#_c_898_n 0.0145938f $X=7.92 $Y=3.33 $X2=0
+ $Y2=0
cc_510 N_VPWR_c_633_n N_A_1013_392#_c_898_n 0.0120466f $X=7.92 $Y=3.33 $X2=0
+ $Y2=0
cc_511 N_X_c_734_n N_VGND_M1005_d 0.00328964f $X=1.415 $Y=1.045 $X2=-0.19
+ $Y2=-0.245
cc_512 N_X_c_737_n N_VGND_M1016_d 0.00176461f $X=2.195 $Y=1.045 $X2=0 $Y2=0
cc_513 N_X_c_734_n N_VGND_c_948_n 0.0219406f $X=1.415 $Y=1.045 $X2=0 $Y2=0
cc_514 N_X_c_736_n N_VGND_c_948_n 0.0164981f $X=1.5 $Y=0.515 $X2=0 $Y2=0
cc_515 N_X_c_736_n N_VGND_c_949_n 0.0157999f $X=1.5 $Y=0.515 $X2=0 $Y2=0
cc_516 N_X_c_737_n N_VGND_c_949_n 0.0135055f $X=2.195 $Y=1.045 $X2=0 $Y2=0
cc_517 N_X_c_738_n N_VGND_c_949_n 0.0157999f $X=2.36 $Y=0.515 $X2=0 $Y2=0
cc_518 N_X_c_738_n N_VGND_c_950_n 0.0109942f $X=2.36 $Y=0.515 $X2=0 $Y2=0
cc_519 N_X_c_738_n N_VGND_c_951_n 0.0216805f $X=2.36 $Y=0.515 $X2=0 $Y2=0
cc_520 N_X_c_736_n N_VGND_c_959_n 0.0109942f $X=1.5 $Y=0.515 $X2=0 $Y2=0
cc_521 N_X_c_736_n N_VGND_c_965_n 0.00904371f $X=1.5 $Y=0.515 $X2=0 $Y2=0
cc_522 N_X_c_738_n N_VGND_c_965_n 0.00904371f $X=2.36 $Y=0.515 $X2=0 $Y2=0
cc_523 N_A_549_392#_c_816_n N_A_814_392#_M1018_d 0.00243452f $X=4.505 $Y=2.99
+ $X2=-0.19 $Y2=1.66
cc_524 N_A_549_392#_M1020_s N_A_814_392#_c_860_n 0.00315345f $X=4.52 $Y=1.96
+ $X2=0 $Y2=0
cc_525 N_A_549_392#_c_817_n N_A_814_392#_c_860_n 0.0220544f $X=4.67 $Y=2.455
+ $X2=0 $Y2=0
cc_526 N_A_549_392#_c_815_n N_A_814_392#_c_861_n 0.0524267f $X=3.77 $Y=2.115
+ $X2=0 $Y2=0
cc_527 N_A_549_392#_c_816_n N_A_814_392#_c_861_n 0.012787f $X=4.505 $Y=2.99
+ $X2=0 $Y2=0
cc_528 N_A_549_392#_c_817_n N_A_814_392#_c_861_n 0.0289859f $X=4.67 $Y=2.455
+ $X2=0 $Y2=0
cc_529 N_A_549_392#_c_817_n N_A_1013_392#_c_890_n 0.046699f $X=4.67 $Y=2.455
+ $X2=0 $Y2=0
cc_530 N_A_549_392#_c_816_n N_A_1013_392#_c_892_n 0.0147157f $X=4.505 $Y=2.99
+ $X2=0 $Y2=0
cc_531 N_A_814_392#_c_860_n N_A_1013_392#_M1000_d 0.00315345f $X=5.475 $Y=2.035
+ $X2=-0.19 $Y2=1.66
cc_532 N_A_814_392#_c_860_n N_A_1013_392#_c_890_n 0.0210301f $X=5.475 $Y=2.035
+ $X2=0 $Y2=0
cc_533 N_A_814_392#_M1000_s N_A_1013_392#_c_891_n 0.00197722f $X=5.49 $Y=1.96
+ $X2=0 $Y2=0
cc_534 N_A_814_392#_c_862_n N_A_1013_392#_c_891_n 0.0160777f $X=5.64 $Y=2.115
+ $X2=0 $Y2=0
cc_535 N_A_814_392#_c_862_n N_A_1013_392#_c_893_n 0.01311f $X=5.64 $Y=2.115
+ $X2=0 $Y2=0
cc_536 N_A_814_392#_c_862_n N_A_1013_392#_c_928_n 0.039994f $X=5.64 $Y=2.115
+ $X2=0 $Y2=0
cc_537 N_VGND_c_955_n N_A_1210_74#_c_1062_n 0.0219626f $X=5.435 $Y=0.515 $X2=0
+ $Y2=0
cc_538 N_VGND_c_956_n N_A_1210_74#_c_1063_n 0.00988046f $X=7.465 $Y=0.585 $X2=0
+ $Y2=0
cc_539 N_VGND_c_963_n N_A_1210_74#_c_1063_n 0.0425255f $X=7.3 $Y=0 $X2=0 $Y2=0
cc_540 N_VGND_c_965_n N_A_1210_74#_c_1063_n 0.0277484f $X=7.92 $Y=0 $X2=0 $Y2=0
cc_541 N_VGND_c_955_n N_A_1210_74#_c_1064_n 0.00816634f $X=5.435 $Y=0.515 $X2=0
+ $Y2=0
cc_542 N_VGND_c_963_n N_A_1210_74#_c_1064_n 0.019738f $X=7.3 $Y=0 $X2=0 $Y2=0
cc_543 N_VGND_c_965_n N_A_1210_74#_c_1064_n 0.012511f $X=7.92 $Y=0 $X2=0 $Y2=0
cc_544 N_VGND_M1009_s N_A_1210_74#_c_1065_n 0.00176461f $X=7.325 $Y=0.37 $X2=0
+ $Y2=0
cc_545 N_VGND_c_956_n N_A_1210_74#_c_1065_n 0.0170777f $X=7.465 $Y=0.585 $X2=0
+ $Y2=0
cc_546 N_VGND_c_956_n N_A_1210_74#_c_1067_n 0.0150645f $X=7.465 $Y=0.585 $X2=0
+ $Y2=0
cc_547 N_VGND_c_964_n N_A_1210_74#_c_1067_n 0.011066f $X=7.92 $Y=0 $X2=0 $Y2=0
cc_548 N_VGND_c_965_n N_A_1210_74#_c_1067_n 0.00915947f $X=7.92 $Y=0 $X2=0 $Y2=0
