# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_hs__a222o_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__a222o_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.800000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.925000 1.120000 3.255000 1.520000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.485000 1.120000 3.825000 1.545000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.220000 1.120000 2.755000 1.790000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.565000 1.180000 1.930000 1.760000 ;
    END
  END B2
  PIN C1
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.120000 0.550000 1.790000 ;
    END
  END C1
  PIN C2
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.060000 1.120000 1.390000 1.760000 ;
    END
  END C2
  PIN X
    ANTENNADIFFAREA  0.541300 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.355000 0.350000 4.710000 1.130000 ;
        RECT 4.355000 1.820000 4.710000 2.980000 ;
        RECT 4.540000 1.130000 4.710000 1.820000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 4.800000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 4.800000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.800000 0.085000 ;
      RECT 0.000000  3.245000 4.800000 3.415000 ;
      RECT 0.115000  1.960000 0.445000 2.905000 ;
      RECT 0.115000  2.905000 2.590000 3.075000 ;
      RECT 0.140000  0.350000 0.470000 0.780000 ;
      RECT 0.140000  0.780000 4.185000 0.950000 ;
      RECT 0.720000  0.950000 0.890000 1.930000 ;
      RECT 0.720000  1.930000 1.050000 2.735000 ;
      RECT 0.960000  0.085000 1.805000 0.600000 ;
      RECT 1.220000  1.930000 1.550000 2.905000 ;
      RECT 1.720000  1.930000 2.050000 1.960000 ;
      RECT 1.720000  1.960000 3.650000 2.130000 ;
      RECT 1.720000  2.130000 2.050000 2.735000 ;
      RECT 2.260000  2.300000 2.590000 2.905000 ;
      RECT 2.295000  0.330000 3.130000 0.780000 ;
      RECT 2.820000  2.300000 3.150000 3.245000 ;
      RECT 3.320000  1.895000 3.650000 1.960000 ;
      RECT 3.320000  2.130000 3.650000 2.935000 ;
      RECT 3.620000  0.085000 4.185000 0.610000 ;
      RECT 3.855000  1.895000 4.185000 3.245000 ;
      RECT 4.015000  0.950000 4.185000 1.300000 ;
      RECT 4.015000  1.300000 4.370000 1.630000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
  END
END sky130_fd_sc_hs__a222o_1
END LIBRARY
