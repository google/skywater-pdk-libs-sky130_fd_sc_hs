# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_hs__mux2i_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.840000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A0
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.525000 1.350000 2.865000 1.780000 ;
    END
  END A0
  PIN A1
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.395000 1.180000 3.725000 1.550000 ;
    END
  END A1
  PIN S
    ANTENNAGATEAREA  0.488000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.180000 0.550000 1.855000 ;
    END
  END S
  PIN Y
    ANTENNADIFFAREA  0.857700 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.495000 0.705000 3.225000 1.035000 ;
        RECT 3.035000 1.035000 3.225000 2.735000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 3.840000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 3.840000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.840000 0.085000 ;
      RECT 0.000000  3.245000 3.840000 3.415000 ;
      RECT 0.105000  2.100000 0.355000 3.245000 ;
      RECT 0.115000  0.085000 0.365000 0.905000 ;
      RECT 0.545000  0.405000 0.890000 0.905000 ;
      RECT 0.555000  2.100000 0.890000 2.980000 ;
      RECT 0.720000  0.905000 0.890000 1.350000 ;
      RECT 0.720000  1.350000 2.130000 1.520000 ;
      RECT 0.720000  1.520000 0.890000 2.100000 ;
      RECT 1.080000  1.820000 1.330000 1.950000 ;
      RECT 1.080000  1.950000 2.835000 2.120000 ;
      RECT 1.080000  2.120000 1.330000 2.980000 ;
      RECT 1.105000  0.350000 1.435000 1.010000 ;
      RECT 1.105000  1.010000 2.275000 1.180000 ;
      RECT 1.530000  2.290000 1.860000 3.245000 ;
      RECT 1.605000  0.085000 1.935000 0.840000 ;
      RECT 1.800000  1.520000 2.130000 1.680000 ;
      RECT 2.060000  2.290000 2.310000 2.905000 ;
      RECT 2.060000  2.905000 3.735000 3.075000 ;
      RECT 2.105000  0.350000 3.680000 0.520000 ;
      RECT 2.105000  0.520000 2.275000 1.010000 ;
      RECT 2.505000  2.120000 2.835000 2.735000 ;
      RECT 3.395000  0.520000 3.680000 1.010000 ;
      RECT 3.405000  1.820000 3.735000 2.905000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
  END
END sky130_fd_sc_hs__mux2i_1
END LIBRARY
