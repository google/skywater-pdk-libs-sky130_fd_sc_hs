* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hs__dfxtp_4 CLK D VGND VNB VPB VPWR Q
X0 a_27_74# CLK VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X1 a_651_503# a_696_458# VPWR VPB sky130_fd_pr__pfet_01v8 w=420000u l=150000u
X2 VGND a_1226_296# Q VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X3 VGND a_544_485# a_696_458# VNB sky130_fd_pr__nfet_01v8_lvt w=550000u l=150000u
X4 a_1034_424# a_27_74# a_1178_124# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X5 VGND a_1226_296# Q VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X6 a_1034_424# a_206_368# a_1141_508# VPB sky130_fd_pr__pfet_01v8 w=420000u l=150000u
X7 a_1226_296# a_1034_424# VPWR VPB sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X8 a_544_485# a_206_368# a_735_102# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X9 Q a_1226_296# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X10 a_1226_296# a_1034_424# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X11 Q a_1226_296# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X12 Q a_1226_296# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X13 Q a_1226_296# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X14 VGND a_27_74# a_206_368# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X15 a_437_503# a_206_368# a_544_485# VPB sky130_fd_pr__pfet_01v8 w=420000u l=150000u
X16 a_696_458# a_27_74# a_1034_424# VPB sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X17 VPWR a_27_74# a_206_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X18 VPWR a_1034_424# a_1226_296# VPB sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X19 VGND D a_437_503# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X20 a_735_102# a_696_458# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X21 a_1141_508# a_1226_296# VPWR VPB sky130_fd_pr__pfet_01v8 w=420000u l=150000u
X22 a_544_485# a_27_74# a_651_503# VPB sky130_fd_pr__pfet_01v8 w=420000u l=150000u
X23 VPWR a_1226_296# Q VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X24 a_696_458# a_206_368# a_1034_424# VNB sky130_fd_pr__nfet_01v8_lvt w=550000u l=150000u
X25 VPWR a_544_485# a_696_458# VPB sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X26 VPWR D a_437_503# VPB sky130_fd_pr__pfet_01v8 w=420000u l=150000u
X27 a_437_503# a_27_74# a_544_485# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X28 VPWR a_1226_296# Q VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X29 a_27_74# CLK VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X30 a_1178_124# a_1226_296# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
.ends
