* File: sky130_fd_sc_hs__or3b_4.pxi.spice
* Created: Tue Sep  1 20:20:57 2020
* 
x_PM_SKY130_FD_SC_HS__OR3B_4%C_N N_C_N_c_112_n N_C_N_c_113_n N_C_N_c_119_n
+ N_C_N_M1013_g N_C_N_M1017_g C_N N_C_N_c_115_n N_C_N_c_116_n N_C_N_c_117_n
+ PM_SKY130_FD_SC_HS__OR3B_4%C_N
x_PM_SKY130_FD_SC_HS__OR3B_4%A N_A_c_149_n N_A_M1000_g N_A_M1015_g N_A_c_150_n
+ N_A_c_158_n N_A_M1007_g N_A_c_151_n N_A_c_152_n N_A_c_165_n A N_A_c_154_n
+ N_A_c_155_n PM_SKY130_FD_SC_HS__OR3B_4%A
x_PM_SKY130_FD_SC_HS__OR3B_4%B N_B_c_242_n N_B_M1003_g N_B_c_243_n N_B_M1016_g
+ N_B_M1008_g B B B N_B_c_245_n B N_B_c_246_n PM_SKY130_FD_SC_HS__OR3B_4%B
x_PM_SKY130_FD_SC_HS__OR3B_4%A_27_392# N_A_27_392#_M1017_s N_A_27_392#_M1013_s
+ N_A_27_392#_c_306_n N_A_27_392#_c_307_n N_A_27_392#_c_321_n
+ N_A_27_392#_M1012_g N_A_27_392#_c_308_n N_A_27_392#_c_309_n
+ N_A_27_392#_c_323_n N_A_27_392#_M1014_g N_A_27_392#_c_310_n
+ N_A_27_392#_M1011_g N_A_27_392#_c_311_n N_A_27_392#_c_312_n
+ N_A_27_392#_c_313_n N_A_27_392#_c_314_n N_A_27_392#_c_315_n
+ N_A_27_392#_c_316_n N_A_27_392#_c_317_n N_A_27_392#_c_318_n
+ N_A_27_392#_c_319_n PM_SKY130_FD_SC_HS__OR3B_4%A_27_392#
x_PM_SKY130_FD_SC_HS__OR3B_4%A_409_392# N_A_409_392#_M1011_s
+ N_A_409_392#_M1008_d N_A_409_392#_M1012_d N_A_409_392#_M1002_g
+ N_A_409_392#_c_410_n N_A_409_392#_M1001_g N_A_409_392#_M1004_g
+ N_A_409_392#_c_411_n N_A_409_392#_M1005_g N_A_409_392#_c_412_n
+ N_A_409_392#_M1006_g N_A_409_392#_M1010_g N_A_409_392#_M1018_g
+ N_A_409_392#_c_413_n N_A_409_392#_M1009_g N_A_409_392#_c_403_n
+ N_A_409_392#_c_421_n N_A_409_392#_c_424_n N_A_409_392#_c_404_n
+ N_A_409_392#_c_405_n N_A_409_392#_c_428_n N_A_409_392#_c_406_n
+ N_A_409_392#_c_407_n N_A_409_392#_c_493_p N_A_409_392#_c_446_n
+ N_A_409_392#_c_436_n N_A_409_392#_c_408_n N_A_409_392#_c_409_n
+ PM_SKY130_FD_SC_HS__OR3B_4%A_409_392#
x_PM_SKY130_FD_SC_HS__OR3B_4%VPWR N_VPWR_M1013_d N_VPWR_M1007_s N_VPWR_M1005_s
+ N_VPWR_M1009_s N_VPWR_c_560_n N_VPWR_c_561_n N_VPWR_c_562_n N_VPWR_c_563_n
+ N_VPWR_c_564_n VPWR N_VPWR_c_565_n N_VPWR_c_566_n N_VPWR_c_567_n
+ N_VPWR_c_568_n N_VPWR_c_569_n N_VPWR_c_570_n N_VPWR_c_571_n N_VPWR_c_559_n
+ PM_SKY130_FD_SC_HS__OR3B_4%VPWR
x_PM_SKY130_FD_SC_HS__OR3B_4%A_217_392# N_A_217_392#_M1000_d
+ N_A_217_392#_M1016_s N_A_217_392#_c_633_n N_A_217_392#_c_631_n
+ N_A_217_392#_c_642_n N_A_217_392#_c_637_n N_A_217_392#_c_632_n
+ PM_SKY130_FD_SC_HS__OR3B_4%A_217_392#
x_PM_SKY130_FD_SC_HS__OR3B_4%A_307_392# N_A_307_392#_M1003_d
+ N_A_307_392#_M1014_s N_A_307_392#_c_669_n
+ PM_SKY130_FD_SC_HS__OR3B_4%A_307_392#
x_PM_SKY130_FD_SC_HS__OR3B_4%X N_X_M1002_d N_X_M1010_d N_X_M1001_d N_X_M1006_d
+ N_X_c_683_n N_X_c_690_n N_X_c_684_n N_X_c_685_n N_X_c_691_n N_X_c_692_n
+ N_X_c_693_n N_X_c_686_n N_X_c_687_n N_X_c_694_n N_X_c_695_n N_X_c_688_n X X
+ PM_SKY130_FD_SC_HS__OR3B_4%X
x_PM_SKY130_FD_SC_HS__OR3B_4%VGND N_VGND_M1017_d N_VGND_M1011_d N_VGND_M1015_d
+ N_VGND_M1004_s N_VGND_M1018_s N_VGND_c_766_n N_VGND_c_767_n N_VGND_c_768_n
+ N_VGND_c_769_n N_VGND_c_770_n N_VGND_c_771_n VGND N_VGND_c_772_n
+ N_VGND_c_773_n N_VGND_c_774_n N_VGND_c_775_n N_VGND_c_776_n N_VGND_c_777_n
+ N_VGND_c_778_n N_VGND_c_779_n N_VGND_c_780_n N_VGND_c_781_n
+ PM_SKY130_FD_SC_HS__OR3B_4%VGND
cc_1 VNB N_C_N_c_112_n 0.00611484f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=1.485
cc_2 VNB N_C_N_c_113_n 0.00993104f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=1.795
cc_3 VNB N_C_N_M1017_g 0.0140578f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=1
cc_4 VNB N_C_N_c_115_n 0.0423064f $X=-0.19 $Y=-0.245 $X2=0.44 $Y2=0.405
cc_5 VNB N_C_N_c_116_n 0.037815f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=0.405
cc_6 VNB N_C_N_c_117_n 0.0241483f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=0.405
cc_7 VNB N_A_c_149_n 0.0264634f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=1.485
cc_8 VNB N_A_c_150_n 0.00626383f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=1
cc_9 VNB N_A_c_151_n 0.00499407f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=0.405
cc_10 VNB N_A_c_152_n 0.0198957f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB A 0.0102241f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=0.405
cc_12 VNB N_A_c_154_n 0.0300625f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=0.447
cc_13 VNB N_A_c_155_n 0.0176886f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_B_c_242_n 0.0191765f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=1.485
cc_15 VNB N_B_c_243_n 0.0161262f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=2.46
cc_16 VNB N_B_M1008_g 0.0292928f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=1
cc_17 VNB N_B_c_245_n 0.00766314f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=0.447
cc_18 VNB N_B_c_246_n 0.00175805f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_27_392#_c_306_n 0.0161855f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=1
cc_20 VNB N_A_27_392#_c_307_n 0.0204404f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=1.395
cc_21 VNB N_A_27_392#_c_308_n 0.0123063f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=0.405
cc_22 VNB N_A_27_392#_c_309_n 0.0169405f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_27_392#_c_310_n 0.0182156f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=0.405
cc_24 VNB N_A_27_392#_c_311_n 0.00756635f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_27_392#_c_312_n 0.00533856f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_27_392#_c_313_n 0.00710076f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_27_392#_c_314_n 0.016362f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_27_392#_c_315_n 0.00704671f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_27_392#_c_316_n 0.00747682f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_27_392#_c_317_n 0.00262689f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_27_392#_c_318_n 0.0878232f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_27_392#_c_319_n 0.00931031f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_409_392#_M1002_g 0.0205516f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_409_392#_M1004_g 0.0212989f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=0.405
cc_35 VNB N_A_409_392#_M1010_g 0.0215504f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_409_392#_M1018_g 0.0232607f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_409_392#_c_403_n 0.00562827f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_409_392#_c_404_n 0.00131771f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_409_392#_c_405_n 0.00206397f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_409_392#_c_406_n 0.00130667f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_409_392#_c_407_n 2.89653e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_409_392#_c_408_n 0.00230657f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_409_392#_c_409_n 0.10325f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_VPWR_c_559_n 0.243291f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_X_c_683_n 0.00180052f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=0.405
cc_46 VNB N_X_c_684_n 0.00305083f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=0.447
cc_47 VNB N_X_c_685_n 0.00132324f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_X_c_686_n 0.00206666f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_X_c_687_n 0.00862347f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_X_c_688_n 0.00178779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB X 0.0263822f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_VGND_c_766_n 0.0157839f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=0.405
cc_53 VNB N_VGND_c_767_n 0.00577372f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_VGND_c_768_n 0.00499242f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=0.447
cc_55 VNB N_VGND_c_769_n 0.00425535f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_VGND_c_770_n 0.0120272f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_VGND_c_771_n 0.0258363f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_VGND_c_772_n 0.0256449f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_VGND_c_773_n 0.0318347f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_VGND_c_774_n 0.0169342f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_VGND_c_775_n 0.0159692f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_VGND_c_776_n 0.0188435f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_VGND_c_777_n 0.00894083f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_VGND_c_778_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_VGND_c_779_n 0.00632462f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_VGND_c_780_n 0.00461913f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_VGND_c_781_n 0.320408f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VPB N_C_N_c_113_n 0.00781167f $X=-0.19 $Y=1.66 $X2=0.5 $Y2=1.795
cc_69 VPB N_C_N_c_119_n 0.0257036f $X=-0.19 $Y=1.66 $X2=0.5 $Y2=1.885
cc_70 VPB N_A_c_149_n 0.0361617f $X=-0.19 $Y=1.66 $X2=0.5 $Y2=1.485
cc_71 VPB N_A_c_150_n 0.00771524f $X=-0.19 $Y=1.66 $X2=0.515 $Y2=1
cc_72 VPB N_A_c_158_n 0.0232443f $X=-0.19 $Y=1.66 $X2=0.515 $Y2=1
cc_73 VPB N_A_c_151_n 0.00237792f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=0.405
cc_74 VPB N_B_c_242_n 0.0348979f $X=-0.19 $Y=1.66 $X2=0.5 $Y2=1.485
cc_75 VPB N_B_c_243_n 0.0341358f $X=-0.19 $Y=1.66 $X2=0.5 $Y2=2.46
cc_76 VPB N_B_c_245_n 0.00935377f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=0.447
cc_77 VPB N_B_c_246_n 0.0011366f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_78 VPB N_A_27_392#_c_307_n 0.00578885f $X=-0.19 $Y=1.66 $X2=0.5 $Y2=1.395
cc_79 VPB N_A_27_392#_c_321_n 0.0224212f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=0.47
cc_80 VPB N_A_27_392#_c_309_n 0.00578885f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_81 VPB N_A_27_392#_c_323_n 0.0216821f $X=-0.19 $Y=1.66 $X2=0.515 $Y2=0.405
cc_82 VPB N_A_27_392#_c_314_n 0.0562726f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_83 VPB N_A_409_392#_c_410_n 0.015951f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=0.405
cc_84 VPB N_A_409_392#_c_411_n 0.0147332f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=0.405
cc_85 VPB N_A_409_392#_c_412_n 0.0152456f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_86 VPB N_A_409_392#_c_413_n 0.016407f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_87 VPB N_A_409_392#_c_407_n 0.00179663f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_88 VPB N_A_409_392#_c_409_n 0.0261127f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_89 VPB N_VPWR_c_560_n 0.016173f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=0.405
cc_90 VPB N_VPWR_c_561_n 0.00890487f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=0.405
cc_91 VPB N_VPWR_c_562_n 0.00507021f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_92 VPB N_VPWR_c_563_n 0.0103331f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=0.447
cc_93 VPB N_VPWR_c_564_n 0.0435928f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_94 VPB N_VPWR_c_565_n 0.0178682f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_95 VPB N_VPWR_c_566_n 0.0682215f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_96 VPB N_VPWR_c_567_n 0.0171897f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_97 VPB N_VPWR_c_568_n 0.0206041f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_98 VPB N_VPWR_c_569_n 0.00614127f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_99 VPB N_VPWR_c_570_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_100 VPB N_VPWR_c_571_n 0.00460249f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_101 VPB N_VPWR_c_559_n 0.0791685f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_102 VPB N_A_217_392#_c_631_n 0.00257348f $X=-0.19 $Y=1.66 $X2=0.44 $Y2=0.405
cc_103 VPB N_A_217_392#_c_632_n 0.00298292f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=0.405
cc_104 VPB N_A_307_392#_c_669_n 0.00814829f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=0.47
cc_105 VPB N_X_c_690_n 0.00181303f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=0.405
cc_106 VPB N_X_c_691_n 0.00217622f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_107 VPB N_X_c_692_n 0.00133248f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=0.447
cc_108 VPB N_X_c_693_n 0.00257348f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_109 VPB N_X_c_694_n 0.00809985f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_110 VPB N_X_c_695_n 0.00187476f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_111 VPB X 0.00685195f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_112 N_C_N_c_112_n N_A_c_149_n 0.0200572f $X=0.5 $Y=1.485 $X2=-0.19 $Y2=-0.245
cc_113 N_C_N_c_113_n N_A_c_149_n 0.00504292f $X=0.5 $Y=1.795 $X2=-0.19
+ $Y2=-0.245
cc_114 N_C_N_c_119_n N_A_c_149_n 0.0182393f $X=0.5 $Y=1.885 $X2=-0.19 $Y2=-0.245
cc_115 N_C_N_c_112_n N_A_c_151_n 0.00121813f $X=0.5 $Y=1.485 $X2=0 $Y2=0
cc_116 N_C_N_M1017_g N_A_c_151_n 0.00236605f $X=0.515 $Y=1 $X2=0 $Y2=0
cc_117 N_C_N_M1017_g N_A_c_165_n 0.00363967f $X=0.515 $Y=1 $X2=0 $Y2=0
cc_118 N_C_N_M1017_g N_A_27_392#_c_313_n 0.00756288f $X=0.515 $Y=1 $X2=0 $Y2=0
cc_119 N_C_N_c_112_n N_A_27_392#_c_314_n 0.0150652f $X=0.5 $Y=1.485 $X2=0 $Y2=0
cc_120 N_C_N_c_119_n N_A_27_392#_c_314_n 0.00653489f $X=0.5 $Y=1.885 $X2=0 $Y2=0
cc_121 N_C_N_M1017_g N_A_27_392#_c_314_n 0.00136405f $X=0.515 $Y=1 $X2=0 $Y2=0
cc_122 N_C_N_M1017_g N_A_27_392#_c_315_n 0.0131846f $X=0.515 $Y=1 $X2=0 $Y2=0
cc_123 N_C_N_c_116_n N_A_27_392#_c_315_n 9.73891e-19 $X=0.61 $Y=0.405 $X2=0
+ $Y2=0
cc_124 N_C_N_c_117_n N_A_27_392#_c_315_n 0.0210442f $X=0.61 $Y=0.405 $X2=0 $Y2=0
cc_125 N_C_N_M1017_g N_A_27_392#_c_316_n 0.00217394f $X=0.515 $Y=1 $X2=0 $Y2=0
cc_126 N_C_N_c_115_n N_A_27_392#_c_316_n 0.00202112f $X=0.44 $Y=0.405 $X2=0
+ $Y2=0
cc_127 N_C_N_c_117_n N_A_27_392#_c_316_n 0.0276654f $X=0.61 $Y=0.405 $X2=0 $Y2=0
cc_128 N_C_N_c_112_n N_A_27_392#_c_319_n 0.00155545f $X=0.5 $Y=1.485 $X2=0 $Y2=0
cc_129 N_C_N_M1017_g N_A_27_392#_c_319_n 0.00529261f $X=0.515 $Y=1 $X2=0 $Y2=0
cc_130 N_C_N_c_119_n N_VPWR_c_560_n 0.0194213f $X=0.5 $Y=1.885 $X2=0 $Y2=0
cc_131 N_C_N_c_119_n N_VPWR_c_565_n 0.00413917f $X=0.5 $Y=1.885 $X2=0 $Y2=0
cc_132 N_C_N_c_119_n N_VPWR_c_559_n 0.00821204f $X=0.5 $Y=1.885 $X2=0 $Y2=0
cc_133 N_C_N_M1017_g N_VGND_c_766_n 3.41717e-19 $X=0.515 $Y=1 $X2=0 $Y2=0
cc_134 N_C_N_c_116_n N_VGND_c_766_n 0.00302495f $X=0.61 $Y=0.405 $X2=0 $Y2=0
cc_135 N_C_N_c_117_n N_VGND_c_766_n 0.0332676f $X=0.61 $Y=0.405 $X2=0 $Y2=0
cc_136 N_C_N_c_115_n N_VGND_c_772_n 0.0116176f $X=0.44 $Y=0.405 $X2=0 $Y2=0
cc_137 N_C_N_c_117_n N_VGND_c_772_n 0.0435286f $X=0.61 $Y=0.405 $X2=0 $Y2=0
cc_138 N_C_N_c_115_n N_VGND_c_781_n 0.00740915f $X=0.44 $Y=0.405 $X2=0 $Y2=0
cc_139 N_C_N_c_116_n N_VGND_c_781_n 0.00763303f $X=0.61 $Y=0.405 $X2=0 $Y2=0
cc_140 N_C_N_c_117_n N_VGND_c_781_n 0.0225644f $X=0.61 $Y=0.405 $X2=0 $Y2=0
cc_141 N_A_c_149_n N_B_c_242_n 0.0340107f $X=1.01 $Y=1.885 $X2=-0.19 $Y2=-0.245
cc_142 N_A_c_151_n N_B_c_242_n 4.89617e-19 $X=0.965 $Y=1.595 $X2=-0.19
+ $Y2=-0.245
cc_143 N_A_c_152_n N_B_c_242_n 0.006956f $X=3.005 $Y=1.235 $X2=-0.19 $Y2=-0.245
cc_144 N_A_c_150_n N_B_c_243_n 0.0127442f $X=3.405 $Y=1.795 $X2=0 $Y2=0
cc_145 N_A_c_158_n N_B_c_243_n 0.0320046f $X=3.405 $Y=1.885 $X2=0 $Y2=0
cc_146 N_A_c_152_n N_B_c_243_n 0.00359328f $X=3.005 $Y=1.235 $X2=0 $Y2=0
cc_147 A N_B_c_243_n 0.00156846f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_148 N_A_c_154_n N_B_c_243_n 0.00503224f $X=3.45 $Y=1.385 $X2=0 $Y2=0
cc_149 N_A_c_152_n N_B_M1008_g 0.00776233f $X=3.005 $Y=1.235 $X2=0 $Y2=0
cc_150 A N_B_M1008_g 0.00564771f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_151 N_A_c_154_n N_B_M1008_g 0.0126306f $X=3.45 $Y=1.385 $X2=0 $Y2=0
cc_152 N_A_c_155_n N_B_M1008_g 0.0113667f $X=3.45 $Y=1.22 $X2=0 $Y2=0
cc_153 N_A_c_150_n N_B_c_245_n 0.00101641f $X=3.405 $Y=1.795 $X2=0 $Y2=0
cc_154 N_A_c_152_n N_B_c_245_n 0.0782005f $X=3.005 $Y=1.235 $X2=0 $Y2=0
cc_155 A N_B_c_245_n 0.00518511f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_156 N_A_c_149_n N_B_c_246_n 0.00119021f $X=1.01 $Y=1.885 $X2=0 $Y2=0
cc_157 N_A_c_151_n N_B_c_246_n 0.017898f $X=0.965 $Y=1.595 $X2=0 $Y2=0
cc_158 N_A_c_152_n N_B_c_246_n 0.0246172f $X=3.005 $Y=1.235 $X2=0 $Y2=0
cc_159 N_A_c_152_n N_A_27_392#_c_306_n 0.00745441f $X=3.005 $Y=1.235 $X2=0 $Y2=0
cc_160 N_A_c_152_n N_A_27_392#_c_308_n 0.00990197f $X=3.005 $Y=1.235 $X2=0 $Y2=0
cc_161 N_A_c_152_n N_A_27_392#_c_310_n 0.00345416f $X=3.005 $Y=1.235 $X2=0 $Y2=0
cc_162 N_A_c_152_n N_A_27_392#_c_311_n 0.00852274f $X=3.005 $Y=1.235 $X2=0 $Y2=0
cc_163 N_A_c_152_n N_A_27_392#_c_312_n 0.00707292f $X=3.005 $Y=1.235 $X2=0 $Y2=0
cc_164 A N_A_27_392#_c_312_n 3.00989e-19 $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_165 N_A_c_165_n N_A_27_392#_c_313_n 0.00835492f $X=1.13 $Y=1.235 $X2=0 $Y2=0
cc_166 N_A_c_151_n N_A_27_392#_c_314_n 0.0162724f $X=0.965 $Y=1.595 $X2=0 $Y2=0
cc_167 N_A_c_149_n N_A_27_392#_c_315_n 0.0012342f $X=1.01 $Y=1.885 $X2=0 $Y2=0
cc_168 N_A_c_152_n N_A_27_392#_c_315_n 0.0593467f $X=3.005 $Y=1.235 $X2=0 $Y2=0
cc_169 N_A_c_165_n N_A_27_392#_c_315_n 0.026613f $X=1.13 $Y=1.235 $X2=0 $Y2=0
cc_170 N_A_c_152_n N_A_27_392#_c_318_n 0.00179644f $X=3.005 $Y=1.235 $X2=0 $Y2=0
cc_171 N_A_c_151_n N_A_27_392#_c_319_n 9.34433e-19 $X=0.965 $Y=1.595 $X2=0 $Y2=0
cc_172 A N_A_409_392#_M1002_g 5.24353e-19 $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_173 N_A_c_154_n N_A_409_392#_M1002_g 0.020457f $X=3.45 $Y=1.385 $X2=0 $Y2=0
cc_174 N_A_c_155_n N_A_409_392#_M1002_g 0.0239844f $X=3.45 $Y=1.22 $X2=0 $Y2=0
cc_175 N_A_c_150_n N_A_409_392#_c_410_n 0.00371178f $X=3.405 $Y=1.795 $X2=0
+ $Y2=0
cc_176 N_A_c_158_n N_A_409_392#_c_410_n 0.0161754f $X=3.405 $Y=1.885 $X2=0 $Y2=0
cc_177 N_A_c_158_n N_A_409_392#_c_421_n 0.0169996f $X=3.405 $Y=1.885 $X2=0 $Y2=0
cc_178 A N_A_409_392#_c_421_n 0.0137967f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_179 N_A_c_154_n N_A_409_392#_c_421_n 0.00217592f $X=3.45 $Y=1.385 $X2=0 $Y2=0
cc_180 N_A_c_152_n N_A_409_392#_c_424_n 0.0382868f $X=3.005 $Y=1.235 $X2=0 $Y2=0
cc_181 A N_A_409_392#_c_424_n 0.00423902f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_182 N_A_c_152_n N_A_409_392#_c_404_n 0.0244317f $X=3.005 $Y=1.235 $X2=0 $Y2=0
cc_183 N_A_c_155_n N_A_409_392#_c_405_n 0.00691851f $X=3.45 $Y=1.22 $X2=0 $Y2=0
cc_184 A N_A_409_392#_c_428_n 0.0133644f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_185 N_A_c_154_n N_A_409_392#_c_428_n 0.00279603f $X=3.45 $Y=1.385 $X2=0 $Y2=0
cc_186 N_A_c_155_n N_A_409_392#_c_428_n 0.00882094f $X=3.45 $Y=1.22 $X2=0 $Y2=0
cc_187 A N_A_409_392#_c_406_n 0.012266f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_188 N_A_c_154_n N_A_409_392#_c_406_n 4.82359e-19 $X=3.45 $Y=1.385 $X2=0 $Y2=0
cc_189 N_A_c_155_n N_A_409_392#_c_406_n 0.00349115f $X=3.45 $Y=1.22 $X2=0 $Y2=0
cc_190 N_A_c_150_n N_A_409_392#_c_407_n 0.00341329f $X=3.405 $Y=1.795 $X2=0
+ $Y2=0
cc_191 N_A_c_158_n N_A_409_392#_c_407_n 0.00166763f $X=3.405 $Y=1.885 $X2=0
+ $Y2=0
cc_192 A N_A_409_392#_c_436_n 0.018439f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_193 N_A_c_155_n N_A_409_392#_c_436_n 7.15494e-19 $X=3.45 $Y=1.22 $X2=0 $Y2=0
cc_194 N_A_c_150_n N_A_409_392#_c_408_n 0.00100335f $X=3.405 $Y=1.795 $X2=0
+ $Y2=0
cc_195 A N_A_409_392#_c_408_n 0.0212197f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_196 N_A_c_154_n N_A_409_392#_c_408_n 0.00176166f $X=3.45 $Y=1.385 $X2=0 $Y2=0
cc_197 N_A_c_150_n N_A_409_392#_c_409_n 0.00715573f $X=3.405 $Y=1.795 $X2=0
+ $Y2=0
cc_198 N_A_c_149_n N_VPWR_c_560_n 0.00985716f $X=1.01 $Y=1.885 $X2=0 $Y2=0
cc_199 N_A_c_151_n N_VPWR_c_560_n 0.00745363f $X=0.965 $Y=1.595 $X2=0 $Y2=0
cc_200 N_A_c_158_n N_VPWR_c_561_n 0.0033662f $X=3.405 $Y=1.885 $X2=0 $Y2=0
cc_201 N_A_c_149_n N_VPWR_c_566_n 0.00445602f $X=1.01 $Y=1.885 $X2=0 $Y2=0
cc_202 N_A_c_158_n N_VPWR_c_566_n 0.00456932f $X=3.405 $Y=1.885 $X2=0 $Y2=0
cc_203 N_A_c_149_n N_VPWR_c_559_n 0.00857821f $X=1.01 $Y=1.885 $X2=0 $Y2=0
cc_204 N_A_c_158_n N_VPWR_c_559_n 0.00890787f $X=3.405 $Y=1.885 $X2=0 $Y2=0
cc_205 N_A_c_149_n N_A_217_392#_c_633_n 0.00401542f $X=1.01 $Y=1.885 $X2=0 $Y2=0
cc_206 N_A_c_151_n N_A_217_392#_c_633_n 0.0024991f $X=0.965 $Y=1.595 $X2=0 $Y2=0
cc_207 N_A_c_152_n N_A_217_392#_c_633_n 0.00581099f $X=3.005 $Y=1.235 $X2=0
+ $Y2=0
cc_208 N_A_c_149_n N_A_217_392#_c_631_n 0.0047544f $X=1.01 $Y=1.885 $X2=0 $Y2=0
cc_209 N_A_c_149_n N_A_217_392#_c_637_n 0.00167066f $X=1.01 $Y=1.885 $X2=0 $Y2=0
cc_210 N_A_c_158_n N_A_217_392#_c_632_n 0.00616038f $X=3.405 $Y=1.885 $X2=0
+ $Y2=0
cc_211 N_A_c_152_n N_VGND_M1017_d 0.00920587f $X=3.005 $Y=1.235 $X2=-0.19
+ $Y2=-0.245
cc_212 N_A_c_165_n N_VGND_M1017_d 0.00744673f $X=1.13 $Y=1.235 $X2=-0.19
+ $Y2=-0.245
cc_213 N_A_c_155_n N_VGND_c_767_n 4.30893e-19 $X=3.45 $Y=1.22 $X2=0 $Y2=0
cc_214 N_A_c_155_n N_VGND_c_768_n 0.00304076f $X=3.45 $Y=1.22 $X2=0 $Y2=0
cc_215 N_A_c_155_n N_VGND_c_774_n 0.00434272f $X=3.45 $Y=1.22 $X2=0 $Y2=0
cc_216 N_A_c_155_n N_VGND_c_781_n 0.00439488f $X=3.45 $Y=1.22 $X2=0 $Y2=0
cc_217 N_B_c_242_n N_A_27_392#_c_307_n 0.021193f $X=1.46 $Y=1.885 $X2=0 $Y2=0
cc_218 N_B_c_245_n N_A_27_392#_c_307_n 0.0122762f $X=2.91 $Y=1.635 $X2=0 $Y2=0
cc_219 N_B_c_246_n N_A_27_392#_c_307_n 4.00295e-19 $X=1.67 $Y=1.645 $X2=0 $Y2=0
cc_220 N_B_c_242_n N_A_27_392#_c_321_n 0.0381125f $X=1.46 $Y=1.885 $X2=0 $Y2=0
cc_221 N_B_c_245_n N_A_27_392#_c_321_n 0.00425914f $X=2.91 $Y=1.635 $X2=0 $Y2=0
cc_222 N_B_c_245_n N_A_27_392#_c_308_n 0.00218423f $X=2.91 $Y=1.635 $X2=0 $Y2=0
cc_223 N_B_c_243_n N_A_27_392#_c_309_n 0.0218359f $X=2.895 $Y=1.885 $X2=0 $Y2=0
cc_224 N_B_c_245_n N_A_27_392#_c_309_n 0.0122762f $X=2.91 $Y=1.635 $X2=0 $Y2=0
cc_225 N_B_c_243_n N_A_27_392#_c_323_n 0.0419538f $X=2.895 $Y=1.885 $X2=0 $Y2=0
cc_226 N_B_c_245_n N_A_27_392#_c_323_n 0.00237826f $X=2.91 $Y=1.635 $X2=0 $Y2=0
cc_227 N_B_M1008_g N_A_27_392#_c_310_n 0.0357543f $X=2.96 $Y=0.74 $X2=0 $Y2=0
cc_228 N_B_c_242_n N_A_27_392#_c_318_n 0.00168855f $X=1.46 $Y=1.885 $X2=0 $Y2=0
cc_229 N_B_M1008_g N_A_409_392#_c_403_n 6.67759e-19 $X=2.96 $Y=0.74 $X2=0 $Y2=0
cc_230 N_B_c_243_n N_A_409_392#_c_421_n 0.0146176f $X=2.895 $Y=1.885 $X2=0 $Y2=0
cc_231 N_B_M1008_g N_A_409_392#_c_424_n 0.00986262f $X=2.96 $Y=0.74 $X2=0 $Y2=0
cc_232 N_B_c_245_n N_A_409_392#_c_407_n 0.00482933f $X=2.91 $Y=1.635 $X2=0 $Y2=0
cc_233 N_B_c_242_n N_A_409_392#_c_446_n 6.62582e-19 $X=1.46 $Y=1.885 $X2=0 $Y2=0
cc_234 N_B_c_243_n N_A_409_392#_c_446_n 2.32791e-19 $X=2.895 $Y=1.885 $X2=0
+ $Y2=0
cc_235 N_B_c_245_n N_A_409_392#_c_446_n 0.066653f $X=2.91 $Y=1.635 $X2=0 $Y2=0
cc_236 N_B_c_245_n N_A_409_392#_c_408_n 0.00254086f $X=2.91 $Y=1.635 $X2=0 $Y2=0
cc_237 N_B_c_242_n N_VPWR_c_566_n 0.00445602f $X=1.46 $Y=1.885 $X2=0 $Y2=0
cc_238 N_B_c_243_n N_VPWR_c_566_n 0.00444483f $X=2.895 $Y=1.885 $X2=0 $Y2=0
cc_239 N_B_c_242_n N_VPWR_c_559_n 0.0044517f $X=1.46 $Y=1.885 $X2=0 $Y2=0
cc_240 N_B_c_243_n N_VPWR_c_559_n 0.00446127f $X=2.895 $Y=1.885 $X2=0 $Y2=0
cc_241 N_B_c_242_n N_A_217_392#_c_633_n 0.00745913f $X=1.46 $Y=1.885 $X2=0 $Y2=0
cc_242 N_B_c_246_n N_A_217_392#_c_633_n 0.00275075f $X=1.67 $Y=1.645 $X2=0 $Y2=0
cc_243 N_B_c_242_n N_A_217_392#_c_631_n 0.00627007f $X=1.46 $Y=1.885 $X2=0 $Y2=0
cc_244 N_B_c_242_n N_A_217_392#_c_642_n 0.0128702f $X=1.46 $Y=1.885 $X2=0 $Y2=0
cc_245 N_B_c_243_n N_A_217_392#_c_642_n 0.0123877f $X=2.895 $Y=1.885 $X2=0 $Y2=0
cc_246 N_B_c_246_n N_A_217_392#_c_642_n 0.016537f $X=1.67 $Y=1.645 $X2=0 $Y2=0
cc_247 N_B_c_242_n N_A_217_392#_c_637_n 2.24111e-19 $X=1.46 $Y=1.885 $X2=0 $Y2=0
cc_248 N_B_c_243_n N_A_217_392#_c_632_n 0.00253633f $X=2.895 $Y=1.885 $X2=0
+ $Y2=0
cc_249 N_B_c_242_n N_A_307_392#_c_669_n 0.00156215f $X=1.46 $Y=1.885 $X2=0 $Y2=0
cc_250 N_B_c_243_n N_A_307_392#_c_669_n 0.00323498f $X=2.895 $Y=1.885 $X2=0
+ $Y2=0
cc_251 N_B_M1008_g N_VGND_c_767_n 0.00740102f $X=2.96 $Y=0.74 $X2=0 $Y2=0
cc_252 N_B_M1008_g N_VGND_c_774_n 0.00383152f $X=2.96 $Y=0.74 $X2=0 $Y2=0
cc_253 N_B_M1008_g N_VGND_c_781_n 0.00377775f $X=2.96 $Y=0.74 $X2=0 $Y2=0
cc_254 N_A_27_392#_c_310_n N_A_409_392#_c_403_n 0.00669352f $X=2.46 $Y=1.185
+ $X2=0 $Y2=0
cc_255 N_A_27_392#_c_317_n N_A_409_392#_c_403_n 0.0363197f $X=1.745 $Y=0.475
+ $X2=0 $Y2=0
cc_256 N_A_27_392#_c_318_n N_A_409_392#_c_403_n 0.00458815f $X=1.745 $Y=0.475
+ $X2=0 $Y2=0
cc_257 N_A_27_392#_c_323_n N_A_409_392#_c_421_n 0.00813086f $X=2.445 $Y=1.885
+ $X2=0 $Y2=0
cc_258 N_A_27_392#_c_310_n N_A_409_392#_c_424_n 0.00877732f $X=2.46 $Y=1.185
+ $X2=0 $Y2=0
cc_259 N_A_27_392#_c_308_n N_A_409_392#_c_404_n 0.00125147f $X=2.355 $Y=1.26
+ $X2=0 $Y2=0
cc_260 N_A_27_392#_c_310_n N_A_409_392#_c_404_n 7.16501e-19 $X=2.46 $Y=1.185
+ $X2=0 $Y2=0
cc_261 N_A_27_392#_c_315_n N_A_409_392#_c_404_n 0.0151541f $X=1.58 $Y=0.895
+ $X2=0 $Y2=0
cc_262 N_A_27_392#_c_318_n N_A_409_392#_c_404_n 0.00180265f $X=1.745 $Y=0.475
+ $X2=0 $Y2=0
cc_263 N_A_27_392#_c_321_n N_A_409_392#_c_446_n 0.00449049f $X=1.97 $Y=1.885
+ $X2=0 $Y2=0
cc_264 N_A_27_392#_c_323_n N_A_409_392#_c_446_n 0.00149457f $X=2.445 $Y=1.885
+ $X2=0 $Y2=0
cc_265 N_A_27_392#_c_314_n N_VPWR_c_560_n 0.0697922f $X=0.275 $Y=2.105 $X2=0
+ $Y2=0
cc_266 N_A_27_392#_c_314_n N_VPWR_c_565_n 0.011066f $X=0.275 $Y=2.105 $X2=0
+ $Y2=0
cc_267 N_A_27_392#_c_321_n N_VPWR_c_566_n 0.00291649f $X=1.97 $Y=1.885 $X2=0
+ $Y2=0
cc_268 N_A_27_392#_c_323_n N_VPWR_c_566_n 0.00291649f $X=2.445 $Y=1.885 $X2=0
+ $Y2=0
cc_269 N_A_27_392#_c_321_n N_VPWR_c_559_n 0.00360347f $X=1.97 $Y=1.885 $X2=0
+ $Y2=0
cc_270 N_A_27_392#_c_323_n N_VPWR_c_559_n 0.00359835f $X=2.445 $Y=1.885 $X2=0
+ $Y2=0
cc_271 N_A_27_392#_c_314_n N_VPWR_c_559_n 0.00915947f $X=0.275 $Y=2.105 $X2=0
+ $Y2=0
cc_272 N_A_27_392#_c_321_n N_A_217_392#_c_633_n 0.00145661f $X=1.97 $Y=1.885
+ $X2=0 $Y2=0
cc_273 N_A_27_392#_c_321_n N_A_217_392#_c_631_n 6.39213e-19 $X=1.97 $Y=1.885
+ $X2=0 $Y2=0
cc_274 N_A_27_392#_c_321_n N_A_217_392#_c_642_n 0.0128326f $X=1.97 $Y=1.885
+ $X2=0 $Y2=0
cc_275 N_A_27_392#_c_323_n N_A_217_392#_c_642_n 0.011084f $X=2.445 $Y=1.885
+ $X2=0 $Y2=0
cc_276 N_A_27_392#_c_321_n N_A_307_392#_c_669_n 0.0114475f $X=1.97 $Y=1.885
+ $X2=0 $Y2=0
cc_277 N_A_27_392#_c_323_n N_A_307_392#_c_669_n 0.0114471f $X=2.445 $Y=1.885
+ $X2=0 $Y2=0
cc_278 N_A_27_392#_c_315_n N_VGND_M1017_d 0.0264369f $X=1.58 $Y=0.895 $X2=-0.19
+ $Y2=-0.245
cc_279 N_A_27_392#_c_315_n N_VGND_c_766_n 0.0368353f $X=1.58 $Y=0.895 $X2=0
+ $Y2=0
cc_280 N_A_27_392#_c_317_n N_VGND_c_766_n 0.0268466f $X=1.745 $Y=0.475 $X2=0
+ $Y2=0
cc_281 N_A_27_392#_c_318_n N_VGND_c_766_n 0.00807651f $X=1.745 $Y=0.475 $X2=0
+ $Y2=0
cc_282 N_A_27_392#_c_310_n N_VGND_c_767_n 0.00416056f $X=2.46 $Y=1.185 $X2=0
+ $Y2=0
cc_283 N_A_27_392#_c_317_n N_VGND_c_767_n 0.00110157f $X=1.745 $Y=0.475 $X2=0
+ $Y2=0
cc_284 N_A_27_392#_c_310_n N_VGND_c_773_n 0.00434272f $X=2.46 $Y=1.185 $X2=0
+ $Y2=0
cc_285 N_A_27_392#_c_317_n N_VGND_c_773_n 0.0163537f $X=1.745 $Y=0.475 $X2=0
+ $Y2=0
cc_286 N_A_27_392#_c_318_n N_VGND_c_773_n 0.00620834f $X=1.745 $Y=0.475 $X2=0
+ $Y2=0
cc_287 N_A_27_392#_c_310_n N_VGND_c_781_n 0.00444308f $X=2.46 $Y=1.185 $X2=0
+ $Y2=0
cc_288 N_A_27_392#_c_315_n N_VGND_c_781_n 0.014088f $X=1.58 $Y=0.895 $X2=0 $Y2=0
cc_289 N_A_27_392#_c_317_n N_VGND_c_781_n 0.0121533f $X=1.745 $Y=0.475 $X2=0
+ $Y2=0
cc_290 N_A_27_392#_c_318_n N_VGND_c_781_n 0.00425878f $X=1.745 $Y=0.475 $X2=0
+ $Y2=0
cc_291 N_A_409_392#_c_421_n N_VPWR_M1007_s 0.00751294f $X=3.715 $Y=2.055 $X2=0
+ $Y2=0
cc_292 N_A_409_392#_c_407_n N_VPWR_M1007_s 0.0015634f $X=3.8 $Y=1.97 $X2=0 $Y2=0
cc_293 N_A_409_392#_c_410_n N_VPWR_c_561_n 0.00196165f $X=3.915 $Y=1.765 $X2=0
+ $Y2=0
cc_294 N_A_409_392#_c_421_n N_VPWR_c_561_n 0.0205313f $X=3.715 $Y=2.055 $X2=0
+ $Y2=0
cc_295 N_A_409_392#_c_410_n N_VPWR_c_562_n 5.86327e-19 $X=3.915 $Y=1.765 $X2=0
+ $Y2=0
cc_296 N_A_409_392#_c_411_n N_VPWR_c_562_n 0.0133793f $X=4.365 $Y=1.765 $X2=0
+ $Y2=0
cc_297 N_A_409_392#_c_412_n N_VPWR_c_562_n 0.00630489f $X=4.815 $Y=1.765 $X2=0
+ $Y2=0
cc_298 N_A_409_392#_c_413_n N_VPWR_c_564_n 0.00993564f $X=5.265 $Y=1.765 $X2=0
+ $Y2=0
cc_299 N_A_409_392#_c_410_n N_VPWR_c_567_n 0.00461464f $X=3.915 $Y=1.765 $X2=0
+ $Y2=0
cc_300 N_A_409_392#_c_411_n N_VPWR_c_567_n 0.00413917f $X=4.365 $Y=1.765 $X2=0
+ $Y2=0
cc_301 N_A_409_392#_c_412_n N_VPWR_c_568_n 0.00445602f $X=4.815 $Y=1.765 $X2=0
+ $Y2=0
cc_302 N_A_409_392#_c_413_n N_VPWR_c_568_n 0.00445602f $X=5.265 $Y=1.765 $X2=0
+ $Y2=0
cc_303 N_A_409_392#_c_410_n N_VPWR_c_559_n 0.00908203f $X=3.915 $Y=1.765 $X2=0
+ $Y2=0
cc_304 N_A_409_392#_c_411_n N_VPWR_c_559_n 0.00817726f $X=4.365 $Y=1.765 $X2=0
+ $Y2=0
cc_305 N_A_409_392#_c_412_n N_VPWR_c_559_n 0.00857589f $X=4.815 $Y=1.765 $X2=0
+ $Y2=0
cc_306 N_A_409_392#_c_413_n N_VPWR_c_559_n 0.0086105f $X=5.265 $Y=1.765 $X2=0
+ $Y2=0
cc_307 N_A_409_392#_c_421_n N_A_217_392#_M1016_s 0.0069199f $X=3.715 $Y=2.055
+ $X2=0 $Y2=0
cc_308 N_A_409_392#_c_446_n N_A_217_392#_c_633_n 0.00577366f $X=2.385 $Y=2.08
+ $X2=0 $Y2=0
cc_309 N_A_409_392#_M1012_d N_A_217_392#_c_642_n 0.00445893f $X=2.045 $Y=1.96
+ $X2=0 $Y2=0
cc_310 N_A_409_392#_c_421_n N_A_217_392#_c_642_n 0.0268572f $X=3.715 $Y=2.055
+ $X2=0 $Y2=0
cc_311 N_A_409_392#_c_446_n N_A_217_392#_c_642_n 0.0176315f $X=2.385 $Y=2.08
+ $X2=0 $Y2=0
cc_312 N_A_409_392#_c_421_n N_A_217_392#_c_632_n 0.0203284f $X=3.715 $Y=2.055
+ $X2=0 $Y2=0
cc_313 N_A_409_392#_c_421_n N_A_307_392#_M1014_s 0.00415853f $X=3.715 $Y=2.055
+ $X2=0 $Y2=0
cc_314 N_A_409_392#_M1012_d N_A_307_392#_c_669_n 0.00228327f $X=2.045 $Y=1.96
+ $X2=0 $Y2=0
cc_315 N_A_409_392#_M1002_g N_X_c_683_n 0.00553314f $X=3.9 $Y=0.74 $X2=0 $Y2=0
cc_316 N_A_409_392#_M1004_g N_X_c_683_n 4.18509e-19 $X=4.355 $Y=0.74 $X2=0 $Y2=0
cc_317 N_A_409_392#_c_428_n N_X_c_683_n 0.0117533f $X=3.715 $Y=0.895 $X2=0 $Y2=0
cc_318 N_A_409_392#_c_410_n N_X_c_690_n 0.00637204f $X=3.915 $Y=1.765 $X2=0
+ $Y2=0
cc_319 N_A_409_392#_c_411_n N_X_c_690_n 0.00438646f $X=4.365 $Y=1.765 $X2=0
+ $Y2=0
cc_320 N_A_409_392#_c_421_n N_X_c_690_n 0.0133252f $X=3.715 $Y=2.055 $X2=0 $Y2=0
cc_321 N_A_409_392#_M1004_g N_X_c_684_n 0.0127369f $X=4.355 $Y=0.74 $X2=0 $Y2=0
cc_322 N_A_409_392#_M1010_g N_X_c_684_n 0.0113812f $X=4.835 $Y=0.74 $X2=0 $Y2=0
cc_323 N_A_409_392#_c_493_p N_X_c_684_n 0.048506f $X=5.01 $Y=1.465 $X2=0 $Y2=0
cc_324 N_A_409_392#_c_409_n N_X_c_684_n 0.00336308f $X=5.265 $Y=1.532 $X2=0
+ $Y2=0
cc_325 N_A_409_392#_M1002_g N_X_c_685_n 7.08499e-19 $X=3.9 $Y=0.74 $X2=0 $Y2=0
cc_326 N_A_409_392#_c_428_n N_X_c_685_n 0.00174806f $X=3.715 $Y=0.895 $X2=0
+ $Y2=0
cc_327 N_A_409_392#_c_406_n N_X_c_685_n 0.0118403f $X=3.8 $Y=1.3 $X2=0 $Y2=0
cc_328 N_A_409_392#_c_493_p N_X_c_685_n 0.0143376f $X=5.01 $Y=1.465 $X2=0 $Y2=0
cc_329 N_A_409_392#_c_409_n N_X_c_685_n 0.00291196f $X=5.265 $Y=1.532 $X2=0
+ $Y2=0
cc_330 N_A_409_392#_c_411_n N_X_c_691_n 0.0130724f $X=4.365 $Y=1.765 $X2=0 $Y2=0
cc_331 N_A_409_392#_c_412_n N_X_c_691_n 0.0119563f $X=4.815 $Y=1.765 $X2=0 $Y2=0
cc_332 N_A_409_392#_c_493_p N_X_c_691_n 0.0477127f $X=5.01 $Y=1.465 $X2=0 $Y2=0
cc_333 N_A_409_392#_c_409_n N_X_c_691_n 0.00923295f $X=5.265 $Y=1.532 $X2=0
+ $Y2=0
cc_334 N_A_409_392#_c_410_n N_X_c_692_n 8.18018e-19 $X=3.915 $Y=1.765 $X2=0
+ $Y2=0
cc_335 N_A_409_392#_c_407_n N_X_c_692_n 0.0134537f $X=3.8 $Y=1.97 $X2=0 $Y2=0
cc_336 N_A_409_392#_c_493_p N_X_c_692_n 0.0143367f $X=5.01 $Y=1.465 $X2=0 $Y2=0
cc_337 N_A_409_392#_c_409_n N_X_c_692_n 0.00413775f $X=5.265 $Y=1.532 $X2=0
+ $Y2=0
cc_338 N_A_409_392#_c_411_n N_X_c_693_n 7.68526e-19 $X=4.365 $Y=1.765 $X2=0
+ $Y2=0
cc_339 N_A_409_392#_c_412_n N_X_c_693_n 0.012705f $X=4.815 $Y=1.765 $X2=0 $Y2=0
cc_340 N_A_409_392#_c_413_n N_X_c_693_n 0.017229f $X=5.265 $Y=1.765 $X2=0 $Y2=0
cc_341 N_A_409_392#_M1004_g N_X_c_686_n 6.97985e-19 $X=4.355 $Y=0.74 $X2=0 $Y2=0
cc_342 N_A_409_392#_M1010_g N_X_c_686_n 0.00939045f $X=4.835 $Y=0.74 $X2=0 $Y2=0
cc_343 N_A_409_392#_M1018_g N_X_c_686_n 3.97481e-19 $X=5.265 $Y=0.74 $X2=0 $Y2=0
cc_344 N_A_409_392#_M1018_g N_X_c_687_n 0.0160624f $X=5.265 $Y=0.74 $X2=0 $Y2=0
cc_345 N_A_409_392#_c_493_p N_X_c_687_n 0.00296926f $X=5.01 $Y=1.465 $X2=0 $Y2=0
cc_346 N_A_409_392#_c_409_n N_X_c_687_n 4.34863e-19 $X=5.265 $Y=1.532 $X2=0
+ $Y2=0
cc_347 N_A_409_392#_c_413_n N_X_c_694_n 0.0152243f $X=5.265 $Y=1.765 $X2=0 $Y2=0
cc_348 N_A_409_392#_c_409_n N_X_c_694_n 5.17675e-19 $X=5.265 $Y=1.532 $X2=0
+ $Y2=0
cc_349 N_A_409_392#_c_412_n N_X_c_695_n 9.3899e-19 $X=4.815 $Y=1.765 $X2=0 $Y2=0
cc_350 N_A_409_392#_c_413_n N_X_c_695_n 0.00114764f $X=5.265 $Y=1.765 $X2=0
+ $Y2=0
cc_351 N_A_409_392#_c_493_p N_X_c_695_n 0.0252322f $X=5.01 $Y=1.465 $X2=0 $Y2=0
cc_352 N_A_409_392#_c_409_n N_X_c_695_n 0.00805362f $X=5.265 $Y=1.532 $X2=0
+ $Y2=0
cc_353 N_A_409_392#_M1010_g N_X_c_688_n 9.7541e-19 $X=4.835 $Y=0.74 $X2=0 $Y2=0
cc_354 N_A_409_392#_c_493_p N_X_c_688_n 0.0209731f $X=5.01 $Y=1.465 $X2=0 $Y2=0
cc_355 N_A_409_392#_c_409_n N_X_c_688_n 0.00232957f $X=5.265 $Y=1.532 $X2=0
+ $Y2=0
cc_356 N_A_409_392#_M1018_g X 0.0067245f $X=5.265 $Y=0.74 $X2=0 $Y2=0
cc_357 N_A_409_392#_c_413_n X 0.00135286f $X=5.265 $Y=1.765 $X2=0 $Y2=0
cc_358 N_A_409_392#_c_493_p X 0.0213231f $X=5.01 $Y=1.465 $X2=0 $Y2=0
cc_359 N_A_409_392#_c_409_n X 0.0159973f $X=5.265 $Y=1.532 $X2=0 $Y2=0
cc_360 N_A_409_392#_c_424_n N_VGND_M1011_d 0.00488266f $X=3.09 $Y=0.895 $X2=0
+ $Y2=0
cc_361 N_A_409_392#_c_428_n N_VGND_M1015_d 0.00765735f $X=3.715 $Y=0.895 $X2=0
+ $Y2=0
cc_362 N_A_409_392#_c_406_n N_VGND_M1015_d 0.00158921f $X=3.8 $Y=1.3 $X2=0 $Y2=0
cc_363 N_A_409_392#_c_403_n N_VGND_c_767_n 0.011672f $X=2.245 $Y=0.515 $X2=0
+ $Y2=0
cc_364 N_A_409_392#_c_424_n N_VGND_c_767_n 0.0204705f $X=3.09 $Y=0.895 $X2=0
+ $Y2=0
cc_365 N_A_409_392#_c_405_n N_VGND_c_767_n 0.011122f $X=3.175 $Y=0.515 $X2=0
+ $Y2=0
cc_366 N_A_409_392#_M1002_g N_VGND_c_768_n 0.00716586f $X=3.9 $Y=0.74 $X2=0
+ $Y2=0
cc_367 N_A_409_392#_M1004_g N_VGND_c_768_n 4.0977e-19 $X=4.355 $Y=0.74 $X2=0
+ $Y2=0
cc_368 N_A_409_392#_c_405_n N_VGND_c_768_n 0.00978394f $X=3.175 $Y=0.515 $X2=0
+ $Y2=0
cc_369 N_A_409_392#_c_428_n N_VGND_c_768_n 0.0183125f $X=3.715 $Y=0.895 $X2=0
+ $Y2=0
cc_370 N_A_409_392#_M1002_g N_VGND_c_769_n 4.55137e-19 $X=3.9 $Y=0.74 $X2=0
+ $Y2=0
cc_371 N_A_409_392#_M1004_g N_VGND_c_769_n 0.00898965f $X=4.355 $Y=0.74 $X2=0
+ $Y2=0
cc_372 N_A_409_392#_M1010_g N_VGND_c_769_n 0.00322767f $X=4.835 $Y=0.74 $X2=0
+ $Y2=0
cc_373 N_A_409_392#_M1010_g N_VGND_c_771_n 5.11007e-19 $X=4.835 $Y=0.74 $X2=0
+ $Y2=0
cc_374 N_A_409_392#_M1018_g N_VGND_c_771_n 0.0113385f $X=5.265 $Y=0.74 $X2=0
+ $Y2=0
cc_375 N_A_409_392#_c_403_n N_VGND_c_773_n 0.0144834f $X=2.245 $Y=0.515 $X2=0
+ $Y2=0
cc_376 N_A_409_392#_c_405_n N_VGND_c_774_n 0.0109336f $X=3.175 $Y=0.515 $X2=0
+ $Y2=0
cc_377 N_A_409_392#_M1002_g N_VGND_c_775_n 0.00383152f $X=3.9 $Y=0.74 $X2=0
+ $Y2=0
cc_378 N_A_409_392#_M1004_g N_VGND_c_775_n 0.00383152f $X=4.355 $Y=0.74 $X2=0
+ $Y2=0
cc_379 N_A_409_392#_M1010_g N_VGND_c_776_n 0.00434272f $X=4.835 $Y=0.74 $X2=0
+ $Y2=0
cc_380 N_A_409_392#_M1018_g N_VGND_c_776_n 0.00383152f $X=5.265 $Y=0.74 $X2=0
+ $Y2=0
cc_381 N_A_409_392#_M1002_g N_VGND_c_781_n 0.00649193f $X=3.9 $Y=0.74 $X2=0
+ $Y2=0
cc_382 N_A_409_392#_M1004_g N_VGND_c_781_n 0.00757785f $X=4.355 $Y=0.74 $X2=0
+ $Y2=0
cc_383 N_A_409_392#_M1010_g N_VGND_c_781_n 0.00821749f $X=4.835 $Y=0.74 $X2=0
+ $Y2=0
cc_384 N_A_409_392#_M1018_g N_VGND_c_781_n 0.0075754f $X=5.265 $Y=0.74 $X2=0
+ $Y2=0
cc_385 N_A_409_392#_c_403_n N_VGND_c_781_n 0.011967f $X=2.245 $Y=0.515 $X2=0
+ $Y2=0
cc_386 N_A_409_392#_c_424_n N_VGND_c_781_n 0.0117123f $X=3.09 $Y=0.895 $X2=0
+ $Y2=0
cc_387 N_A_409_392#_c_405_n N_VGND_c_781_n 0.00901999f $X=3.175 $Y=0.515 $X2=0
+ $Y2=0
cc_388 N_A_409_392#_c_428_n N_VGND_c_781_n 0.00763539f $X=3.715 $Y=0.895 $X2=0
+ $Y2=0
cc_389 N_VPWR_c_560_n N_A_217_392#_c_631_n 0.016852f $X=0.725 $Y=2.105 $X2=0
+ $Y2=0
cc_390 N_VPWR_c_566_n N_A_217_392#_c_631_n 0.014552f $X=3.505 $Y=3.33 $X2=0
+ $Y2=0
cc_391 N_VPWR_c_559_n N_A_217_392#_c_631_n 0.0119791f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_392 N_VPWR_c_559_n N_A_217_392#_c_642_n 0.01233f $X=5.52 $Y=3.33 $X2=0 $Y2=0
cc_393 N_VPWR_c_561_n N_A_217_392#_c_632_n 0.017638f $X=3.67 $Y=2.475 $X2=0
+ $Y2=0
cc_394 N_VPWR_c_566_n N_A_217_392#_c_632_n 0.0146079f $X=3.505 $Y=3.33 $X2=0
+ $Y2=0
cc_395 N_VPWR_c_559_n N_A_217_392#_c_632_n 0.0120887f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_396 N_VPWR_c_566_n N_A_307_392#_c_669_n 0.0515327f $X=3.505 $Y=3.33 $X2=0
+ $Y2=0
cc_397 N_VPWR_c_559_n N_A_307_392#_c_669_n 0.0435095f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_398 N_VPWR_c_561_n N_X_c_690_n 0.0207936f $X=3.67 $Y=2.475 $X2=0 $Y2=0
cc_399 N_VPWR_c_562_n N_X_c_690_n 0.0535896f $X=4.59 $Y=2.305 $X2=0 $Y2=0
cc_400 N_VPWR_c_567_n N_X_c_690_n 0.00749631f $X=4.425 $Y=3.33 $X2=0 $Y2=0
cc_401 N_VPWR_c_559_n N_X_c_690_n 0.0062048f $X=5.52 $Y=3.33 $X2=0 $Y2=0
cc_402 N_VPWR_M1005_s N_X_c_691_n 0.00222494f $X=4.44 $Y=1.84 $X2=0 $Y2=0
cc_403 N_VPWR_c_562_n N_X_c_691_n 0.0154248f $X=4.59 $Y=2.305 $X2=0 $Y2=0
cc_404 N_VPWR_c_562_n N_X_c_693_n 0.0563525f $X=4.59 $Y=2.305 $X2=0 $Y2=0
cc_405 N_VPWR_c_564_n N_X_c_693_n 0.0563525f $X=5.49 $Y=2.305 $X2=0 $Y2=0
cc_406 N_VPWR_c_568_n N_X_c_693_n 0.014552f $X=5.405 $Y=3.33 $X2=0 $Y2=0
cc_407 N_VPWR_c_559_n N_X_c_693_n 0.0119791f $X=5.52 $Y=3.33 $X2=0 $Y2=0
cc_408 N_VPWR_M1009_s N_X_c_694_n 0.00344613f $X=5.34 $Y=1.84 $X2=0 $Y2=0
cc_409 N_VPWR_c_564_n N_X_c_694_n 0.0206356f $X=5.49 $Y=2.305 $X2=0 $Y2=0
cc_410 N_A_217_392#_c_642_n N_A_307_392#_M1003_d 0.0070808f $X=3.005 $Y=2.445
+ $X2=-0.19 $Y2=1.66
cc_411 N_A_217_392#_c_642_n N_A_307_392#_M1014_s 0.00414445f $X=3.005 $Y=2.445
+ $X2=0 $Y2=0
cc_412 N_A_217_392#_c_631_n N_A_307_392#_c_669_n 0.0108142f $X=1.235 $Y=2.815
+ $X2=0 $Y2=0
cc_413 N_A_217_392#_c_642_n N_A_307_392#_c_669_n 0.0686384f $X=3.005 $Y=2.445
+ $X2=0 $Y2=0
cc_414 N_A_217_392#_c_632_n N_A_307_392#_c_669_n 0.0124625f $X=3.17 $Y=2.475
+ $X2=0 $Y2=0
cc_415 N_X_c_684_n N_VGND_M1004_s 0.00364486f $X=4.885 $Y=1.045 $X2=0 $Y2=0
cc_416 N_X_c_687_n N_VGND_M1018_s 0.00338075f $X=5.405 $Y=1.045 $X2=0 $Y2=0
cc_417 N_X_c_683_n N_VGND_c_768_n 0.0160427f $X=4.14 $Y=0.515 $X2=0 $Y2=0
cc_418 N_X_c_683_n N_VGND_c_769_n 0.0157999f $X=4.14 $Y=0.515 $X2=0 $Y2=0
cc_419 N_X_c_684_n N_VGND_c_769_n 0.015373f $X=4.885 $Y=1.045 $X2=0 $Y2=0
cc_420 N_X_c_686_n N_VGND_c_769_n 0.0259969f $X=5.05 $Y=0.515 $X2=0 $Y2=0
cc_421 N_X_c_686_n N_VGND_c_771_n 0.0164981f $X=5.05 $Y=0.515 $X2=0 $Y2=0
cc_422 N_X_c_687_n N_VGND_c_771_n 0.023173f $X=5.405 $Y=1.045 $X2=0 $Y2=0
cc_423 N_X_c_683_n N_VGND_c_775_n 0.00749631f $X=4.14 $Y=0.515 $X2=0 $Y2=0
cc_424 N_X_c_686_n N_VGND_c_776_n 0.0109942f $X=5.05 $Y=0.515 $X2=0 $Y2=0
cc_425 N_X_c_683_n N_VGND_c_781_n 0.0062048f $X=4.14 $Y=0.515 $X2=0 $Y2=0
cc_426 N_X_c_686_n N_VGND_c_781_n 0.00904371f $X=5.05 $Y=0.515 $X2=0 $Y2=0
