* File: sky130_fd_sc_hs__a2bb2o_4.pex.spice
* Created: Tue Sep  1 19:51:52 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HS__A2BB2O_4%A_162_48# 1 2 3 12 14 16 19 21 23 26 28 30
+ 33 35 37 38 43 46 47 48 50 51 52 53 54 57 61 63 67 71
c166 33 0 1.57686e-19 $X=2.175 $Y=0.74
r167 78 79 40.0639 $w=3.91e-07 $l=3.25e-07 $layer=POLY_cond $X=1.85 $Y=1.532
+ $X2=2.175 $Y2=1.532
r168 77 78 12.9437 $w=3.91e-07 $l=1.05e-07 $layer=POLY_cond $X=1.745 $Y=1.532
+ $X2=1.85 $Y2=1.532
r169 76 77 42.5294 $w=3.91e-07 $l=3.45e-07 $layer=POLY_cond $X=1.4 $Y=1.532
+ $X2=1.745 $Y2=1.532
r170 75 76 10.4783 $w=3.91e-07 $l=8.5e-08 $layer=POLY_cond $X=1.315 $Y=1.532
+ $X2=1.4 $Y2=1.532
r171 72 73 8.01279 $w=3.91e-07 $l=6.5e-08 $layer=POLY_cond $X=0.885 $Y=1.532
+ $X2=0.95 $Y2=1.532
r172 67 81 9.86189 $w=3.91e-07 $l=8e-08 $layer=POLY_cond $X=2.22 $Y=1.532
+ $X2=2.3 $Y2=1.532
r173 67 79 5.54731 $w=3.91e-07 $l=4.5e-08 $layer=POLY_cond $X=2.22 $Y=1.532
+ $X2=2.175 $Y2=1.532
r174 59 70 3.40825 $w=2.5e-07 $l=1.25e-07 $layer=LI1_cond $X=4.815 $Y=0.475
+ $X2=4.69 $Y2=0.475
r175 59 61 36.1867 $w=2.48e-07 $l=7.85e-07 $layer=LI1_cond $X=4.815 $Y=0.475
+ $X2=5.6 $Y2=0.475
r176 55 71 4.10697 $w=2.22e-07 $l=9.80051e-08 $layer=LI1_cond $X=4.662 $Y=1.18
+ $X2=4.69 $Y2=1.095
r177 55 57 52.6107 $w=1.93e-07 $l=9.25e-07 $layer=LI1_cond $X=4.662 $Y=1.18
+ $X2=4.662 $Y2=2.105
r178 54 71 4.10697 $w=2.22e-07 $l=8.5e-08 $layer=LI1_cond $X=4.69 $Y=1.01
+ $X2=4.69 $Y2=1.095
r179 53 70 3.40825 $w=2.5e-07 $l=1.25e-07 $layer=LI1_cond $X=4.69 $Y=0.6
+ $X2=4.69 $Y2=0.475
r180 53 54 18.9001 $w=2.48e-07 $l=4.1e-07 $layer=LI1_cond $X=4.69 $Y=0.6
+ $X2=4.69 $Y2=1.01
r181 51 71 2.32734 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.565 $Y=1.095
+ $X2=4.69 $Y2=1.095
r182 51 52 67.5241 $w=1.68e-07 $l=1.035e-06 $layer=LI1_cond $X=4.565 $Y=1.095
+ $X2=3.53 $Y2=1.095
r183 50 52 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.445 $Y=1.01
+ $X2=3.53 $Y2=1.095
r184 49 50 38.1658 $w=1.68e-07 $l=5.85e-07 $layer=LI1_cond $X=3.445 $Y=0.425
+ $X2=3.445 $Y2=1.01
r185 47 49 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.36 $Y=0.34
+ $X2=3.445 $Y2=0.425
r186 47 48 35.5561 $w=1.68e-07 $l=5.45e-07 $layer=LI1_cond $X=3.36 $Y=0.34
+ $X2=2.815 $Y2=0.34
r187 45 48 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.73 $Y=0.425
+ $X2=2.815 $Y2=0.34
r188 45 46 38.1658 $w=1.68e-07 $l=5.85e-07 $layer=LI1_cond $X=2.73 $Y=0.425
+ $X2=2.73 $Y2=1.01
r189 44 63 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.385 $Y=1.095
+ $X2=2.3 $Y2=1.095
r190 43 46 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.645 $Y=1.095
+ $X2=2.73 $Y2=1.01
r191 43 44 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=2.645 $Y=1.095
+ $X2=2.385 $Y2=1.095
r192 41 75 14.1765 $w=3.91e-07 $l=1.15e-07 $layer=POLY_cond $X=1.2 $Y=1.532
+ $X2=1.315 $Y2=1.532
r193 41 73 30.8184 $w=3.91e-07 $l=2.5e-07 $layer=POLY_cond $X=1.2 $Y=1.532
+ $X2=0.95 $Y2=1.532
r194 40 41 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.2
+ $Y=1.465 $X2=1.2 $Y2=1.465
r195 38 67 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.22
+ $Y=1.465 $X2=2.22 $Y2=1.465
r196 38 63 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=2.3 $Y=1.465 $X2=2.3
+ $Y2=1.095
r197 38 40 35.4464 $w=3.28e-07 $l=1.015e-06 $layer=LI1_cond $X=2.215 $Y=1.465
+ $X2=1.2 $Y2=1.465
r198 35 81 25.3065 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=2.3 $Y=1.765
+ $X2=2.3 $Y2=1.532
r199 35 37 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.3 $Y=1.765
+ $X2=2.3 $Y2=2.4
r200 31 79 25.3065 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=2.175 $Y=1.3
+ $X2=2.175 $Y2=1.532
r201 31 33 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=2.175 $Y=1.3
+ $X2=2.175 $Y2=0.74
r202 28 78 25.3065 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=1.85 $Y=1.765
+ $X2=1.85 $Y2=1.532
r203 28 30 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.85 $Y=1.765
+ $X2=1.85 $Y2=2.4
r204 24 77 25.3065 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=1.745 $Y=1.3
+ $X2=1.745 $Y2=1.532
r205 24 26 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=1.745 $Y=1.3
+ $X2=1.745 $Y2=0.74
r206 21 76 25.3065 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=1.4 $Y=1.765
+ $X2=1.4 $Y2=1.532
r207 21 23 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.4 $Y=1.765
+ $X2=1.4 $Y2=2.4
r208 17 75 25.3065 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=1.315 $Y=1.3
+ $X2=1.315 $Y2=1.532
r209 17 19 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=1.315 $Y=1.3
+ $X2=1.315 $Y2=0.74
r210 14 73 25.3065 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=0.95 $Y=1.765
+ $X2=0.95 $Y2=1.532
r211 14 16 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.95 $Y=1.765
+ $X2=0.95 $Y2=2.4
r212 10 72 25.3065 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=0.885 $Y=1.3
+ $X2=0.885 $Y2=1.532
r213 10 12 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=0.885 $Y=1.3
+ $X2=0.885 $Y2=0.74
r214 3 57 300 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=2 $X=4.525
+ $Y=1.96 $X2=4.675 $Y2=2.105
r215 2 61 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=5.46
+ $Y=0.37 $X2=5.6 $Y2=0.515
r216 1 70 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=4.51
+ $Y=0.37 $X2=4.65 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__A2BB2O_4%A1_N 1 3 6 8 12
r37 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.765
+ $Y=1.515 $X2=2.765 $Y2=1.515
r38 8 12 5.85988 $w=2.93e-07 $l=1.5e-07 $layer=LI1_cond $X=2.702 $Y=1.665
+ $X2=2.702 $Y2=1.515
r39 4 11 38.5562 $w=2.99e-07 $l=2.05122e-07 $layer=POLY_cond $X=2.855 $Y=1.35
+ $X2=2.765 $Y2=1.515
r40 4 6 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=2.855 $Y=1.35
+ $X2=2.855 $Y2=0.79
r41 1 11 52.2586 $w=2.99e-07 $l=2.85044e-07 $layer=POLY_cond $X=2.84 $Y=1.765
+ $X2=2.765 $Y2=1.515
r42 1 3 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.84 $Y=1.765
+ $X2=2.84 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_HS__A2BB2O_4%A2_N 1 3 6 8
r32 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.445
+ $Y=1.515 $X2=3.445 $Y2=1.515
r33 8 12 4.15415 $w=4.28e-07 $l=1.55e-07 $layer=LI1_cond $X=3.6 $Y=1.565
+ $X2=3.445 $Y2=1.565
r34 4 11 39.7867 $w=4.1e-07 $l=2.05122e-07 $layer=POLY_cond $X=3.285 $Y=1.35
+ $X2=3.375 $Y2=1.515
r35 4 6 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=3.285 $Y=1.35
+ $X2=3.285 $Y2=0.79
r36 1 11 49.7794 $w=4.1e-07 $l=3.14245e-07 $layer=POLY_cond $X=3.23 $Y=1.765
+ $X2=3.375 $Y2=1.515
r37 1 3 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.23 $Y=1.765
+ $X2=3.23 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_HS__A2BB2O_4%A_586_94# 1 2 7 11 13 15 16 18 20 21 23 27
+ 30 33 35 36 39 40 42
r89 43 46 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=3.105 $Y=2.035
+ $X2=3.455 $Y2=2.035
r90 40 49 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=3.985 $Y=1.635
+ $X2=3.985 $Y2=1.725
r91 39 40 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.985
+ $Y=1.635 $X2=3.985 $Y2=1.635
r92 37 39 12.3057 $w=2.93e-07 $l=3.15e-07 $layer=LI1_cond $X=4.002 $Y=1.95
+ $X2=4.002 $Y2=1.635
r93 36 46 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=3.62 $Y=2.035
+ $X2=3.455 $Y2=2.035
r94 35 37 7.47753 $w=1.7e-07 $l=1.84673e-07 $layer=LI1_cond $X=3.855 $Y=2.035
+ $X2=4.002 $Y2=1.95
r95 35 36 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=3.855 $Y=2.035
+ $X2=3.62 $Y2=2.035
r96 33 46 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=3.455 $Y=2.815
+ $X2=3.455 $Y2=2.12
r97 30 43 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.105 $Y=1.95
+ $X2=3.105 $Y2=2.035
r98 30 42 53.4973 $w=1.68e-07 $l=8.2e-07 $layer=LI1_cond $X=3.105 $Y=1.95
+ $X2=3.105 $Y2=1.13
r99 25 42 5.87448 $w=2.03e-07 $l=1.02e-07 $layer=LI1_cond $X=3.087 $Y=1.028
+ $X2=3.087 $Y2=1.13
r100 25 27 12.0647 $w=2.03e-07 $l=2.23e-07 $layer=LI1_cond $X=3.087 $Y=1.028
+ $X2=3.087 $Y2=0.805
r101 21 22 31.303 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=4.45 $Y=1.725
+ $X2=4.45 $Y2=1.65
r102 18 23 64.3434 $w=1.8e-07 $l=1.6e-07 $layer=POLY_cond $X=4.9 $Y=1.885
+ $X2=4.9 $Y2=1.725
r103 18 20 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=4.9 $Y=1.885
+ $X2=4.9 $Y2=2.46
r104 17 21 7.1379 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=4.54 $Y=1.725 $X2=4.45
+ $Y2=1.725
r105 16 23 7.1379 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=4.81 $Y=1.725 $X2=4.9
+ $Y2=1.725
r106 16 17 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=4.81 $Y=1.725
+ $X2=4.54 $Y2=1.725
r107 13 21 64.3434 $w=1.8e-07 $l=1.6e-07 $layer=POLY_cond $X=4.45 $Y=1.885
+ $X2=4.45 $Y2=1.725
r108 13 15 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=4.45 $Y=1.885
+ $X2=4.45 $Y2=2.46
r109 11 22 466.617 $w=1.5e-07 $l=9.1e-07 $layer=POLY_cond $X=4.435 $Y=0.74
+ $X2=4.435 $Y2=1.65
r110 8 49 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.15 $Y=1.725
+ $X2=3.985 $Y2=1.725
r111 7 21 7.1379 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=4.36 $Y=1.725 $X2=4.45
+ $Y2=1.725
r112 7 8 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=4.36 $Y=1.725
+ $X2=4.15 $Y2=1.725
r113 2 46 400 $w=1.7e-07 $l=3.4187e-07 $layer=licon1_PDIFF $count=1 $X=3.305
+ $Y=1.84 $X2=3.455 $Y2=2.115
r114 2 33 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=3.305
+ $Y=1.84 $X2=3.455 $Y2=2.815
r115 1 27 182 $w=1.7e-07 $l=3.98905e-07 $layer=licon1_NDIFF $count=1 $X=2.93
+ $Y=0.47 $X2=3.07 $Y2=0.805
.ends

.subckt PM_SKY130_FD_SC_HS__A2BB2O_4%B2 2 3 5 8 11 12 14 17 19 20 30
c53 17 0 1.56257e-19 $X=5.815 $Y=0.69
r54 29 30 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=5.8 $Y=1.425
+ $X2=5.815 $Y2=1.425
r55 27 29 40.2181 $w=3.3e-07 $l=2.3e-07 $layer=POLY_cond $X=5.57 $Y=1.425
+ $X2=5.8 $Y2=1.425
r56 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.57
+ $Y=1.425 $X2=5.57 $Y2=1.425
r57 25 27 32.3493 $w=3.3e-07 $l=1.85e-07 $layer=POLY_cond $X=5.385 $Y=1.425
+ $X2=5.57 $Y2=1.425
r58 23 25 6.12014 $w=3.3e-07 $l=3.5e-08 $layer=POLY_cond $X=5.35 $Y=1.425
+ $X2=5.385 $Y2=1.425
r59 20 28 9.89065 $w=5.18e-07 $l=4.3e-07 $layer=LI1_cond $X=6 $Y=1.52 $X2=5.57
+ $Y2=1.52
r60 19 28 1.15008 $w=5.18e-07 $l=5e-08 $layer=LI1_cond $X=5.52 $Y=1.52 $X2=5.57
+ $Y2=1.52
r61 15 30 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.815 $Y=1.26
+ $X2=5.815 $Y2=1.425
r62 15 17 292.277 $w=1.5e-07 $l=5.7e-07 $layer=POLY_cond $X=5.815 $Y=1.26
+ $X2=5.815 $Y2=0.69
r63 12 14 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=5.8 $Y=1.885
+ $X2=5.8 $Y2=2.46
r64 11 12 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=5.8 $Y=1.795 $X2=5.8
+ $Y2=1.885
r65 10 29 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=5.8 $Y=1.59 $X2=5.8
+ $Y2=1.425
r66 10 11 79.6855 $w=1.8e-07 $l=2.05e-07 $layer=POLY_cond $X=5.8 $Y=1.59 $X2=5.8
+ $Y2=1.795
r67 6 25 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.385 $Y=1.26
+ $X2=5.385 $Y2=1.425
r68 6 8 292.277 $w=1.5e-07 $l=5.7e-07 $layer=POLY_cond $X=5.385 $Y=1.26
+ $X2=5.385 $Y2=0.69
r69 3 5 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=5.35 $Y=1.885
+ $X2=5.35 $Y2=2.46
r70 2 3 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=5.35 $Y=1.795 $X2=5.35
+ $Y2=1.885
r71 1 23 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=5.35 $Y=1.59
+ $X2=5.35 $Y2=1.425
r72 1 2 79.6855 $w=1.8e-07 $l=2.05e-07 $layer=POLY_cond $X=5.35 $Y=1.59 $X2=5.35
+ $Y2=1.795
.ends

.subckt PM_SKY130_FD_SC_HS__A2BB2O_4%B1 2 5 7 9 11 12 14 17 19 20 30
c48 5 0 1.39795e-19 $X=6.245 $Y=0.69
r49 29 30 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=6.7 $Y=1.425
+ $X2=6.715 $Y2=1.425
r50 27 29 29.7264 $w=3.3e-07 $l=1.7e-07 $layer=POLY_cond $X=6.53 $Y=1.425
+ $X2=6.7 $Y2=1.425
r51 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.53
+ $Y=1.425 $X2=6.53 $Y2=1.425
r52 25 27 48.9612 $w=3.3e-07 $l=2.8e-07 $layer=POLY_cond $X=6.25 $Y=1.425
+ $X2=6.53 $Y2=1.425
r53 23 25 0.874306 $w=3.3e-07 $l=5e-09 $layer=POLY_cond $X=6.245 $Y=1.425
+ $X2=6.25 $Y2=1.425
r54 20 28 9.89065 $w=5.18e-07 $l=4.3e-07 $layer=LI1_cond $X=6.96 $Y=1.52
+ $X2=6.53 $Y2=1.52
r55 19 28 1.15008 $w=5.18e-07 $l=5e-08 $layer=LI1_cond $X=6.48 $Y=1.52 $X2=6.53
+ $Y2=1.52
r56 15 30 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.715 $Y=1.26
+ $X2=6.715 $Y2=1.425
r57 15 17 292.277 $w=1.5e-07 $l=5.7e-07 $layer=POLY_cond $X=6.715 $Y=1.26
+ $X2=6.715 $Y2=0.69
r58 12 14 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=6.7 $Y=1.885
+ $X2=6.7 $Y2=2.46
r59 11 12 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=6.7 $Y=1.795 $X2=6.7
+ $Y2=1.885
r60 10 29 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=6.7 $Y=1.59 $X2=6.7
+ $Y2=1.425
r61 10 11 79.6855 $w=1.8e-07 $l=2.05e-07 $layer=POLY_cond $X=6.7 $Y=1.59 $X2=6.7
+ $Y2=1.795
r62 7 9 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=6.25 $Y=1.885
+ $X2=6.25 $Y2=2.46
r63 3 23 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.245 $Y=1.26
+ $X2=6.245 $Y2=1.425
r64 3 5 292.277 $w=1.5e-07 $l=5.7e-07 $layer=POLY_cond $X=6.245 $Y=1.26
+ $X2=6.245 $Y2=0.69
r65 2 7 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=6.25 $Y=1.795 $X2=6.25
+ $Y2=1.885
r66 1 25 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=6.25 $Y=1.59
+ $X2=6.25 $Y2=1.425
r67 1 2 79.6855 $w=1.8e-07 $l=2.05e-07 $layer=POLY_cond $X=6.25 $Y=1.59 $X2=6.25
+ $Y2=1.795
.ends

.subckt PM_SKY130_FD_SC_HS__A2BB2O_4%VPWR 1 2 3 4 5 18 22 26 32 36 39 40 42 43
+ 44 46 55 59 72 73 76 79 82
r87 82 83 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r88 79 80 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r89 76 77 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r90 72 73 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r91 70 73 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6 $Y=3.33 $X2=6.96
+ $Y2=3.33
r92 70 83 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=3.33 $X2=5.52
+ $Y2=3.33
r93 69 70 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r94 67 82 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.66 $Y=3.33
+ $X2=5.535 $Y2=3.33
r95 67 69 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=5.66 $Y=3.33 $X2=6
+ $Y2=3.33
r96 66 83 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=5.52 $Y2=3.33
r97 65 66 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r98 63 80 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=2.64 $Y2=3.33
r99 62 65 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=3.12 $Y=3.33
+ $X2=5.04 $Y2=3.33
r100 62 63 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r101 60 79 9.31531 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=2.78 $Y=3.33
+ $X2=2.595 $Y2=3.33
r102 60 62 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=2.78 $Y=3.33
+ $X2=3.12 $Y2=3.33
r103 59 82 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.41 $Y=3.33
+ $X2=5.535 $Y2=3.33
r104 59 65 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=5.41 $Y=3.33
+ $X2=5.04 $Y2=3.33
r105 58 80 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r106 57 58 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r107 55 79 9.31531 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=2.41 $Y=3.33
+ $X2=2.595 $Y2=3.33
r108 55 57 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=2.41 $Y=3.33
+ $X2=2.16 $Y2=3.33
r109 54 58 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.16 $Y2=3.33
r110 54 77 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r111 53 54 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r112 51 76 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.81 $Y=3.33
+ $X2=0.685 $Y2=3.33
r113 51 53 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=0.81 $Y=3.33
+ $X2=1.2 $Y2=3.33
r114 49 77 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r115 48 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r116 46 76 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.56 $Y=3.33
+ $X2=0.685 $Y2=3.33
r117 46 48 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=0.56 $Y=3.33
+ $X2=0.24 $Y2=3.33
r118 44 66 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=5.04 $Y2=3.33
r119 44 63 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=3.12 $Y2=3.33
r120 42 69 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=6.39 $Y=3.33 $X2=6
+ $Y2=3.33
r121 42 43 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.39 $Y=3.33
+ $X2=6.475 $Y2=3.33
r122 41 72 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=6.56 $Y=3.33 $X2=6.96
+ $Y2=3.33
r123 41 43 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.56 $Y=3.33
+ $X2=6.475 $Y2=3.33
r124 39 53 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=1.54 $Y=3.33
+ $X2=1.2 $Y2=3.33
r125 39 40 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.54 $Y=3.33
+ $X2=1.625 $Y2=3.33
r126 38 57 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=1.71 $Y=3.33
+ $X2=2.16 $Y2=3.33
r127 38 40 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.71 $Y=3.33
+ $X2=1.625 $Y2=3.33
r128 34 43 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.475 $Y=3.245
+ $X2=6.475 $Y2=3.33
r129 34 36 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=6.475 $Y=3.245
+ $X2=6.475 $Y2=2.455
r130 30 82 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.535 $Y=3.245
+ $X2=5.535 $Y2=3.33
r131 30 32 36.4172 $w=2.48e-07 $l=7.9e-07 $layer=LI1_cond $X=5.535 $Y=3.245
+ $X2=5.535 $Y2=2.455
r132 26 29 21.803 $w=3.68e-07 $l=7e-07 $layer=LI1_cond $X=2.595 $Y=2.115
+ $X2=2.595 $Y2=2.815
r133 24 79 1.24149 $w=3.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.595 $Y=3.245
+ $X2=2.595 $Y2=3.33
r134 24 29 13.3933 $w=3.68e-07 $l=4.3e-07 $layer=LI1_cond $X=2.595 $Y=3.245
+ $X2=2.595 $Y2=2.815
r135 20 40 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.625 $Y=3.245
+ $X2=1.625 $Y2=3.33
r136 20 22 61.3262 $w=1.68e-07 $l=9.4e-07 $layer=LI1_cond $X=1.625 $Y=3.245
+ $X2=1.625 $Y2=2.305
r137 16 76 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.685 $Y=3.245
+ $X2=0.685 $Y2=3.33
r138 16 18 43.3319 $w=2.48e-07 $l=9.4e-07 $layer=LI1_cond $X=0.685 $Y=3.245
+ $X2=0.685 $Y2=2.305
r139 5 36 300 $w=1.7e-07 $l=5.65044e-07 $layer=licon1_PDIFF $count=2 $X=6.325
+ $Y=1.96 $X2=6.475 $Y2=2.455
r140 4 32 300 $w=1.7e-07 $l=5.65044e-07 $layer=licon1_PDIFF $count=2 $X=5.425
+ $Y=1.96 $X2=5.575 $Y2=2.455
r141 3 29 400 $w=1.7e-07 $l=1.07941e-06 $layer=licon1_PDIFF $count=1 $X=2.375
+ $Y=1.84 $X2=2.595 $Y2=2.815
r142 3 26 400 $w=1.7e-07 $l=3.68951e-07 $layer=licon1_PDIFF $count=1 $X=2.375
+ $Y=1.84 $X2=2.595 $Y2=2.115
r143 2 22 300 $w=1.7e-07 $l=5.34766e-07 $layer=licon1_PDIFF $count=2 $X=1.475
+ $Y=1.84 $X2=1.625 $Y2=2.305
r144 1 18 300 $w=1.7e-07 $l=5.23784e-07 $layer=licon1_PDIFF $count=2 $X=0.6
+ $Y=1.84 $X2=0.725 $Y2=2.305
.ends

.subckt PM_SKY130_FD_SC_HS__A2BB2O_4%X 1 2 3 4 13 14 17 21 25 27 31 35 39 40 42
c68 25 0 1.57686e-19 $X=1.795 $Y=1.045
r69 40 42 9.22205 $w=6.35e-07 $l=4.8e-07 $layer=LI1_cond $X=0.24 $Y=1.465
+ $X2=0.72 $Y2=1.465
r70 35 37 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=2.075 $Y=1.985
+ $X2=2.075 $Y2=2.815
r71 33 35 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=2.075 $Y=1.97
+ $X2=2.075 $Y2=1.985
r72 29 31 20.5135 $w=2.48e-07 $l=4.45e-07 $layer=LI1_cond $X=1.92 $Y=0.96
+ $X2=1.92 $Y2=0.515
r73 28 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.34 $Y=1.885
+ $X2=1.175 $Y2=1.885
r74 27 33 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.91 $Y=1.885
+ $X2=2.075 $Y2=1.97
r75 27 28 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=1.91 $Y=1.885
+ $X2=1.34 $Y2=1.885
r76 25 29 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.795 $Y=1.045
+ $X2=1.92 $Y2=0.96
r77 21 23 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=1.175 $Y=1.985
+ $X2=1.175 $Y2=2.815
r78 19 39 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.175 $Y=1.97
+ $X2=1.175 $Y2=1.885
r79 19 21 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=1.175 $Y=1.97
+ $X2=1.175 $Y2=1.985
r80 15 42 6.53228 $w=6.35e-07 $l=6.53242e-07 $layer=LI1_cond $X=1.06 $Y=0.96
+ $X2=0.72 $Y2=1.465
r81 15 17 20.5135 $w=2.48e-07 $l=4.45e-07 $layer=LI1_cond $X=1.06 $Y=0.96
+ $X2=1.06 $Y2=0.515
r82 14 15 9.82347 $w=6.35e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.185 $Y=1.045
+ $X2=1.06 $Y2=0.96
r83 14 25 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=1.185 $Y=1.045
+ $X2=1.795 $Y2=1.045
r84 13 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.01 $Y=1.885
+ $X2=1.175 $Y2=1.885
r85 13 14 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=1.01 $Y=1.885
+ $X2=0.835 $Y2=1.885
r86 4 37 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=1.925
+ $Y=1.84 $X2=2.075 $Y2=2.815
r87 4 35 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=1.925
+ $Y=1.84 $X2=2.075 $Y2=1.985
r88 3 23 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=1.025
+ $Y=1.84 $X2=1.175 $Y2=2.815
r89 3 21 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=1.025
+ $Y=1.84 $X2=1.175 $Y2=1.985
r90 2 31 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.82
+ $Y=0.37 $X2=1.96 $Y2=0.515
r91 1 17 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=0.96
+ $Y=0.37 $X2=1.1 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__A2BB2O_4%A_820_392# 1 2 3 4 15 17 18 19 22 23 27 29
+ 31 33 38
r65 31 40 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.925 $Y=2.12
+ $X2=6.925 $Y2=2.035
r66 31 33 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=6.925 $Y=2.12
+ $X2=6.925 $Y2=2.815
r67 30 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.19 $Y=2.035
+ $X2=6.025 $Y2=2.035
r68 29 40 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.76 $Y=2.035
+ $X2=6.925 $Y2=2.035
r69 29 30 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=6.76 $Y=2.035
+ $X2=6.19 $Y2=2.035
r70 25 38 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.025 $Y=2.12
+ $X2=6.025 $Y2=2.035
r71 25 27 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=6.025 $Y=2.12
+ $X2=6.025 $Y2=2.815
r72 24 36 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.21 $Y=2.035
+ $X2=5.085 $Y2=2.035
r73 23 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.86 $Y=2.035
+ $X2=6.025 $Y2=2.035
r74 23 24 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=5.86 $Y=2.035
+ $X2=5.21 $Y2=2.035
r75 20 22 4.14879 $w=2.48e-07 $l=9e-08 $layer=LI1_cond $X=5.085 $Y=2.905
+ $X2=5.085 $Y2=2.815
r76 19 36 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.085 $Y=2.12
+ $X2=5.085 $Y2=2.035
r77 19 22 32.0379 $w=2.48e-07 $l=6.95e-07 $layer=LI1_cond $X=5.085 $Y=2.12
+ $X2=5.085 $Y2=2.815
r78 17 20 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=4.96 $Y=2.99
+ $X2=5.085 $Y2=2.905
r79 17 18 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=4.96 $Y=2.99
+ $X2=4.39 $Y2=2.99
r80 13 18 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.225 $Y=2.905
+ $X2=4.39 $Y2=2.99
r81 13 15 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=4.225 $Y=2.905
+ $X2=4.225 $Y2=2.455
r82 4 40 400 $w=1.7e-07 $l=2.17428e-07 $layer=licon1_PDIFF $count=1 $X=6.775
+ $Y=1.96 $X2=6.925 $Y2=2.115
r83 4 33 400 $w=1.7e-07 $l=9.26971e-07 $layer=licon1_PDIFF $count=1 $X=6.775
+ $Y=1.96 $X2=6.925 $Y2=2.815
r84 3 38 400 $w=1.7e-07 $l=2.17428e-07 $layer=licon1_PDIFF $count=1 $X=5.875
+ $Y=1.96 $X2=6.025 $Y2=2.115
r85 3 27 400 $w=1.7e-07 $l=9.26971e-07 $layer=licon1_PDIFF $count=1 $X=5.875
+ $Y=1.96 $X2=6.025 $Y2=2.815
r86 2 36 400 $w=1.7e-07 $l=2.17428e-07 $layer=licon1_PDIFF $count=1 $X=4.975
+ $Y=1.96 $X2=5.125 $Y2=2.115
r87 2 22 400 $w=1.7e-07 $l=9.26971e-07 $layer=licon1_PDIFF $count=1 $X=4.975
+ $Y=1.96 $X2=5.125 $Y2=2.815
r88 1 15 300 $w=1.7e-07 $l=5.53986e-07 $layer=licon1_PDIFF $count=2 $X=4.1
+ $Y=1.96 $X2=4.225 $Y2=2.455
.ends

.subckt PM_SKY130_FD_SC_HS__A2BB2O_4%VGND 1 2 3 4 5 18 22 26 30 36 37 39 40 42
+ 43 45 46 49 50 51 63 78 79 82
r95 82 83 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r96 78 79 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=0 $X2=6.96
+ $Y2=0
r97 76 79 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=0 $X2=6.96
+ $Y2=0
r98 75 76 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6.48 $Y=0 $X2=6.48
+ $Y2=0
r99 73 76 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=4.56 $Y=0 $X2=6.48
+ $Y2=0
r100 73 83 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=4.08
+ $Y2=0
r101 72 75 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=4.56 $Y=0 $X2=6.48
+ $Y2=0
r102 72 73 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.56 $Y=0
+ $X2=4.56 $Y2=0
r103 70 82 13.5049 $w=1.7e-07 $l=3.43e-07 $layer=LI1_cond $X=4.385 $Y=0
+ $X2=4.042 $Y2=0
r104 70 72 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=4.385 $Y=0
+ $X2=4.56 $Y2=0
r105 65 68 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=2.64 $Y=0 $X2=3.6
+ $Y2=0
r106 65 66 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r107 63 82 13.5049 $w=1.7e-07 $l=3.42e-07 $layer=LI1_cond $X=3.7 $Y=0 $X2=4.042
+ $Y2=0
r108 63 68 6.52406 $w=1.68e-07 $l=1e-07 $layer=LI1_cond $X=3.7 $Y=0 $X2=3.6
+ $Y2=0
r109 62 66 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r110 61 62 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r111 59 62 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r112 58 59 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r113 55 59 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=1.2
+ $Y2=0
r114 54 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r115 51 83 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.08
+ $Y2=0
r116 51 66 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=2.64
+ $Y2=0
r117 51 68 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r118 49 75 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=6.495 $Y=0 $X2=6.48
+ $Y2=0
r119 49 50 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.495 $Y=0 $X2=6.58
+ $Y2=0
r120 48 78 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=6.665 $Y=0 $X2=6.96
+ $Y2=0
r121 48 50 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.665 $Y=0 $X2=6.58
+ $Y2=0
r122 45 46 9.62896 $w=3.68e-07 $l=2e-07 $layer=LI1_cond $X=6.48 $Y=0.55 $X2=6.48
+ $Y2=0.35
r123 42 61 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=2.225 $Y=0 $X2=2.16
+ $Y2=0
r124 42 43 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.225 $Y=0 $X2=2.35
+ $Y2=0
r125 41 65 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=2.475 $Y=0
+ $X2=2.64 $Y2=0
r126 41 43 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.475 $Y=0 $X2=2.35
+ $Y2=0
r127 39 58 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=1.365 $Y=0 $X2=1.2
+ $Y2=0
r128 39 40 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.365 $Y=0 $X2=1.49
+ $Y2=0
r129 38 61 35.5561 $w=1.68e-07 $l=5.45e-07 $layer=LI1_cond $X=1.615 $Y=0
+ $X2=2.16 $Y2=0
r130 38 40 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.615 $Y=0 $X2=1.49
+ $Y2=0
r131 36 54 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.505 $Y=0
+ $X2=0.24 $Y2=0
r132 36 37 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.505 $Y=0 $X2=0.63
+ $Y2=0
r133 35 58 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=0.755 $Y=0 $X2=1.2
+ $Y2=0
r134 35 37 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.755 $Y=0 $X2=0.63
+ $Y2=0
r135 33 50 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.58 $Y=0.085
+ $X2=6.58 $Y2=0
r136 33 46 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=6.58 $Y=0.085
+ $X2=6.58 $Y2=0.35
r137 28 82 2.81621 $w=6.85e-07 $l=8.5e-08 $layer=LI1_cond $X=4.042 $Y=0.085
+ $X2=4.042 $Y2=0
r138 28 30 10.302 $w=6.83e-07 $l=5.9e-07 $layer=LI1_cond $X=4.042 $Y=0.085
+ $X2=4.042 $Y2=0.675
r139 24 43 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.35 $Y=0.085
+ $X2=2.35 $Y2=0
r140 24 26 27.1977 $w=2.48e-07 $l=5.9e-07 $layer=LI1_cond $X=2.35 $Y=0.085
+ $X2=2.35 $Y2=0.675
r141 20 40 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.49 $Y=0.085
+ $X2=1.49 $Y2=0
r142 20 22 24.8928 $w=2.48e-07 $l=5.4e-07 $layer=LI1_cond $X=1.49 $Y=0.085
+ $X2=1.49 $Y2=0.625
r143 16 37 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.63 $Y=0.085
+ $X2=0.63 $Y2=0
r144 16 18 24.8928 $w=2.48e-07 $l=5.4e-07 $layer=LI1_cond $X=0.63 $Y=0.085
+ $X2=0.63 $Y2=0.625
r145 5 45 182 $w=1.7e-07 $l=2.47386e-07 $layer=licon1_NDIFF $count=1 $X=6.32
+ $Y=0.37 $X2=6.48 $Y2=0.55
r146 4 30 182 $w=1.7e-07 $l=9.57027e-07 $layer=licon1_NDIFF $count=1 $X=3.36
+ $Y=0.47 $X2=4.22 $Y2=0.675
r147 4 30 182 $w=1.7e-07 $l=5.17446e-07 $layer=licon1_NDIFF $count=1 $X=3.36
+ $Y=0.47 $X2=3.785 $Y2=0.675
r148 3 26 182 $w=1.7e-07 $l=3.68409e-07 $layer=licon1_NDIFF $count=1 $X=2.25
+ $Y=0.37 $X2=2.39 $Y2=0.675
r149 2 22 182 $w=1.7e-07 $l=3.17372e-07 $layer=licon1_NDIFF $count=1 $X=1.39
+ $Y=0.37 $X2=1.53 $Y2=0.625
r150 1 18 182 $w=1.7e-07 $l=3.11288e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.37 $X2=0.67 $Y2=0.625
.ends

.subckt PM_SKY130_FD_SC_HS__A2BB2O_4%A_1009_74# 1 2 3 10 16 18 22 25
c30 16 0 2.96052e-19 $X=6.03 $Y=0.515
r31 20 22 18.6696 $w=2.48e-07 $l=4.05e-07 $layer=LI1_cond $X=6.97 $Y=0.92
+ $X2=6.97 $Y2=0.515
r32 19 25 3.77418 $w=2.45e-07 $l=1.16619e-07 $layer=LI1_cond $X=6.115 $Y=1.005
+ $X2=6.03 $Y2=0.93
r33 18 20 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=6.845 $Y=1.005
+ $X2=6.97 $Y2=0.92
r34 18 19 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=6.845 $Y=1.005
+ $X2=6.115 $Y2=1.005
r35 14 25 2.68609 $w=1.7e-07 $l=1.6e-07 $layer=LI1_cond $X=6.03 $Y=0.77 $X2=6.03
+ $Y2=0.93
r36 14 16 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=6.03 $Y=0.77
+ $X2=6.03 $Y2=0.515
r37 10 25 3.77418 $w=2.45e-07 $l=8.5e-08 $layer=LI1_cond $X=5.945 $Y=0.93
+ $X2=6.03 $Y2=0.93
r38 10 12 27.9107 $w=3.18e-07 $l=7.75e-07 $layer=LI1_cond $X=5.945 $Y=0.93
+ $X2=5.17 $Y2=0.93
r39 3 22 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=6.79
+ $Y=0.37 $X2=6.93 $Y2=0.515
r40 2 25 182 $w=1.7e-07 $l=5.60647e-07 $layer=licon1_NDIFF $count=1 $X=5.89
+ $Y=0.37 $X2=6.03 $Y2=0.865
r41 2 16 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=5.89
+ $Y=0.37 $X2=6.03 $Y2=0.515
r42 1 12 182 $w=1.7e-07 $l=5.48954e-07 $layer=licon1_NDIFF $count=1 $X=5.045
+ $Y=0.37 $X2=5.17 $Y2=0.86
.ends

