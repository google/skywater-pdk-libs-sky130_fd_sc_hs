# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_hs__dlrtp_2
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_hs__dlrtp_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  7.200000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.208500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.450000 0.515000 1.780000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.567400 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.255000 0.350000 6.585000 0.960000 ;
        RECT 6.255000 0.960000 7.075000 1.130000 ;
        RECT 6.255000 2.060000 6.585000 2.980000 ;
        RECT 6.415000 1.800000 7.075000 1.970000 ;
        RECT 6.415000 1.970000 6.585000 2.060000 ;
        RECT 6.845000 1.130000 7.075000 1.800000 ;
    END
  END Q
  PIN RESET_B
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.435000 1.180000 5.840000 1.550000 ;
    END
  END RESET_B
  PIN GATE
    ANTENNAGATEAREA  0.237000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 1.025000 1.180000 1.285000 1.550000 ;
    END
  END GATE
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 7.200000 0.085000 ;
        RECT 0.650000  0.085000 0.980000 0.940000 ;
        RECT 2.305000  0.085000 2.635000 0.410000 ;
        RECT 4.285000  0.085000 4.615000 0.845000 ;
        RECT 5.755000  0.085000 6.085000 1.010000 ;
        RECT 6.755000  0.085000 7.085000 0.790000 ;
      LAYER mcon ;
        RECT 0.155000 -0.085000 0.325000 0.085000 ;
        RECT 0.635000 -0.085000 0.805000 0.085000 ;
        RECT 1.115000 -0.085000 1.285000 0.085000 ;
        RECT 1.595000 -0.085000 1.765000 0.085000 ;
        RECT 2.075000 -0.085000 2.245000 0.085000 ;
        RECT 2.555000 -0.085000 2.725000 0.085000 ;
        RECT 3.035000 -0.085000 3.205000 0.085000 ;
        RECT 3.515000 -0.085000 3.685000 0.085000 ;
        RECT 3.995000 -0.085000 4.165000 0.085000 ;
        RECT 4.475000 -0.085000 4.645000 0.085000 ;
        RECT 4.955000 -0.085000 5.125000 0.085000 ;
        RECT 5.435000 -0.085000 5.605000 0.085000 ;
        RECT 5.915000 -0.085000 6.085000 0.085000 ;
        RECT 6.395000 -0.085000 6.565000 0.085000 ;
        RECT 6.875000 -0.085000 7.045000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.245000 7.200000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 3.245000 7.200000 3.415000 ;
        RECT 0.650000 2.780000 0.980000 3.245000 ;
        RECT 2.280000 2.780000 2.610000 3.245000 ;
        RECT 4.450000 2.650000 5.085000 3.245000 ;
        RECT 5.755000 2.060000 6.085000 3.245000 ;
        RECT 6.755000 2.140000 7.085000 3.245000 ;
      LAYER mcon ;
        RECT 0.155000 3.245000 0.325000 3.415000 ;
        RECT 0.635000 3.245000 0.805000 3.415000 ;
        RECT 1.115000 3.245000 1.285000 3.415000 ;
        RECT 1.595000 3.245000 1.765000 3.415000 ;
        RECT 2.075000 3.245000 2.245000 3.415000 ;
        RECT 2.555000 3.245000 2.725000 3.415000 ;
        RECT 3.035000 3.245000 3.205000 3.415000 ;
        RECT 3.515000 3.245000 3.685000 3.415000 ;
        RECT 3.995000 3.245000 4.165000 3.415000 ;
        RECT 4.475000 3.245000 4.645000 3.415000 ;
        RECT 4.955000 3.245000 5.125000 3.415000 ;
        RECT 5.435000 3.245000 5.605000 3.415000 ;
        RECT 5.915000 3.245000 6.085000 3.415000 ;
        RECT 6.395000 3.245000 6.565000 3.415000 ;
        RECT 6.875000 3.245000 7.045000 3.415000 ;
      LAYER met1 ;
        RECT 0.000000 3.085000 7.200000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.115000 1.950000 0.855000 2.440000 ;
      RECT 0.115000 2.440000 2.680000 2.610000 ;
      RECT 0.115000 2.610000 0.445000 2.820000 ;
      RECT 0.140000 0.540000 0.470000 1.110000 ;
      RECT 0.140000 1.110000 0.855000 1.280000 ;
      RECT 0.685000 1.280000 0.855000 1.950000 ;
      RECT 1.150000 0.350000 1.625000 0.580000 ;
      RECT 1.150000 0.580000 2.975000 0.750000 ;
      RECT 1.150000 0.750000 1.625000 1.010000 ;
      RECT 1.185000 1.940000 1.625000 2.270000 ;
      RECT 1.455000 1.010000 1.625000 1.420000 ;
      RECT 1.455000 1.420000 1.890000 1.750000 ;
      RECT 1.455000 1.750000 1.625000 1.940000 ;
      RECT 1.795000 0.920000 2.230000 1.080000 ;
      RECT 1.795000 1.080000 3.315000 1.250000 ;
      RECT 1.825000 1.940000 2.230000 2.270000 ;
      RECT 2.060000 1.250000 2.230000 1.940000 ;
      RECT 2.510000 1.440000 2.840000 1.770000 ;
      RECT 2.510000 1.770000 2.680000 2.440000 ;
      RECT 2.805000 0.255000 4.090000 0.425000 ;
      RECT 2.805000 0.425000 2.975000 0.580000 ;
      RECT 2.890000 1.940000 3.220000 2.110000 ;
      RECT 2.890000 2.110000 3.060000 2.905000 ;
      RECT 2.890000 2.905000 4.060000 3.075000 ;
      RECT 3.050000 1.250000 3.315000 1.450000 ;
      RECT 3.050000 1.450000 3.220000 1.940000 ;
      RECT 3.205000 0.595000 3.715000 0.845000 ;
      RECT 3.230000 2.405000 3.560000 2.735000 ;
      RECT 3.390000 1.760000 4.925000 1.930000 ;
      RECT 3.390000 1.930000 3.560000 2.405000 ;
      RECT 3.485000 0.845000 3.655000 1.760000 ;
      RECT 3.730000 2.100000 4.060000 2.905000 ;
      RECT 3.825000 1.260000 4.090000 1.590000 ;
      RECT 3.920000 0.425000 4.090000 1.260000 ;
      RECT 4.300000 2.100000 5.585000 2.380000 ;
      RECT 4.660000 1.350000 4.925000 1.760000 ;
      RECT 4.845000 0.350000 5.265000 1.130000 ;
      RECT 5.095000 1.130000 5.265000 1.720000 ;
      RECT 5.095000 1.720000 6.220000 1.890000 ;
      RECT 5.095000 1.890000 5.585000 2.100000 ;
      RECT 5.255000 2.380000 5.585000 2.980000 ;
      RECT 6.050000 1.300000 6.675000 1.630000 ;
      RECT 6.050000 1.630000 6.220000 1.720000 ;
  END
END sky130_fd_sc_hs__dlrtp_2
