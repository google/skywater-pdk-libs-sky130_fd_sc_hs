* File: sky130_fd_sc_hs__o311ai_1.spice
* Created: Tue Sep  1 20:17:37 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hs__o311ai_1.pex.spice"
.subckt sky130_fd_sc_hs__o311ai_1  VNB VPB A1 A2 A3 B1 C1 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* C1	C1
* B1	B1
* A3	A3
* A2	A2
* A1	A1
* VPB	VPB
* VNB	VNB
MM1005 N_A_128_74#_M1005_d N_A1_M1005_g N_VGND_M1005_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.11285 AS=0.2627 PD=1.045 PS=2.19 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75000.3
+ SB=75002.4 A=0.111 P=1.78 MULT=1
MM1008 N_VGND_M1008_d N_A2_M1008_g N_A_128_74#_M1005_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.222 AS=0.11285 PD=1.34 PS=1.045 NRD=27.564 NRS=4.044 M=1 R=4.93333
+ SA=75000.7 SB=75001.9 A=0.111 P=1.78 MULT=1
MM1009 N_A_128_74#_M1009_d N_A3_M1009_g N_VGND_M1008_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.1295 AS=0.222 PD=1.09 PS=1.34 NRD=11.34 NRS=24.324 M=1 R=4.93333
+ SA=75001.5 SB=75001.2 A=0.111 P=1.78 MULT=1
MM1007 A_469_74# N_B1_M1007_g N_A_128_74#_M1009_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.1147 AS=0.1295 PD=1.05 PS=1.09 NRD=16.212 NRS=0 M=1 R=4.93333 SA=75002
+ SB=75000.7 A=0.111 P=1.78 MULT=1
MM1001 N_Y_M1001_d N_C1_M1001_g A_469_74# VNB NLOWVT L=0.15 W=0.74 AD=0.2109
+ AS=0.1147 PD=2.05 PS=1.05 NRD=0 NRS=16.212 M=1 R=4.93333 SA=75002.4 SB=75000.2
+ A=0.111 P=1.78 MULT=1
MM1006 A_138_368# N_A1_M1006_g N_VPWR_M1006_s VPB PSHORT L=0.15 W=1.12 AD=0.1512
+ AS=0.3304 PD=1.39 PS=2.83 NRD=14.0658 NRS=1.7533 M=1 R=7.46667 SA=75000.2
+ SB=75002.3 A=0.168 P=2.54 MULT=1
MM1003 A_222_368# N_A2_M1003_g A_138_368# VPB PSHORT L=0.15 W=1.12 AD=0.2352
+ AS=0.1512 PD=1.54 PS=1.39 NRD=27.2451 NRS=14.0658 M=1 R=7.46667 SA=75000.6
+ SB=75001.9 A=0.168 P=2.54 MULT=1
MM1000 N_Y_M1000_d N_A3_M1000_g A_222_368# VPB PSHORT L=0.15 W=1.12 AD=0.2352
+ AS=0.2352 PD=1.54 PS=1.54 NRD=22.852 NRS=27.2451 M=1 R=7.46667 SA=75001.2
+ SB=75001.4 A=0.168 P=2.54 MULT=1
MM1004 N_VPWR_M1004_d N_B1_M1004_g N_Y_M1000_d VPB PSHORT L=0.15 W=1.12
+ AD=0.2352 AS=0.2352 PD=1.54 PS=1.54 NRD=10.5395 NRS=1.7533 M=1 R=7.46667
+ SA=75001.8 SB=75000.8 A=0.168 P=2.54 MULT=1
MM1002 N_Y_M1002_d N_C1_M1002_g N_VPWR_M1004_d VPB PSHORT L=0.15 W=1.12
+ AD=0.3304 AS=0.2352 PD=2.83 PS=1.54 NRD=1.7533 NRS=14.0658 M=1 R=7.46667
+ SA=75002.3 SB=75000.2 A=0.168 P=2.54 MULT=1
DX10_noxref VNB VPB NWDIODE A=6.9564 P=11.2
*
.include "sky130_fd_sc_hs__o311ai_1.pxi.spice"
*
.ends
*
*
