* NGSPICE file created from sky130_fd_sc_hs__decap_8.ext - technology: sky130A

.subckt sky130_fd_sc_hs__decap_8 VGND VNB VPB VPWR
M1000 VPWR VGND VPWR VPB pshort w=1e+06u l=1e+06u
+  ad=8.35e+11p pd=7.67e+06u as=0p ps=0u
M1001 VGND VPWR VGND VNB nlowvt w=420000u l=1e+06u
+  ad=3.465e+11p pd=4.17e+06u as=0p ps=0u
M1002 VPWR VGND VPWR VPB pshort w=1e+06u l=1e+06u
+  ad=0p pd=0u as=0p ps=0u
M1003 VGND VPWR VGND VNB nlowvt w=420000u l=1e+06u
+  ad=0p pd=0u as=0p ps=0u
.ends

