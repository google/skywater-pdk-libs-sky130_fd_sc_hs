* File: sky130_fd_sc_hs__xnor2_2.pxi.spice
* Created: Tue Sep  1 20:25:16 2020
* 
x_PM_SKY130_FD_SC_HS__XNOR2_2%A N_A_c_91_n N_A_M1015_g N_A_c_92_n N_A_M1011_g
+ N_A_c_93_n N_A_M1008_g N_A_c_94_n N_A_M1004_g N_A_c_95_n N_A_M1009_g
+ N_A_M1005_g N_A_c_97_n N_A_c_108_n N_A_c_109_n A N_A_c_99_n N_A_c_100_n
+ N_A_c_101_n N_A_c_102_n N_A_c_103_n PM_SKY130_FD_SC_HS__XNOR2_2%A
x_PM_SKY130_FD_SC_HS__XNOR2_2%B N_B_M1010_g N_B_c_245_n N_B_M1003_g N_B_c_235_n
+ N_B_M1000_g N_B_c_246_n N_B_M1006_g N_B_c_236_n N_B_M1002_g N_B_c_247_n
+ N_B_M1007_g N_B_c_237_n N_B_c_238_n N_B_c_239_n N_B_c_251_n N_B_c_252_n
+ N_B_c_275_n N_B_c_253_n N_B_c_328_p N_B_c_240_n N_B_c_241_n N_B_c_242_n B
+ N_B_c_244_n PM_SKY130_FD_SC_HS__XNOR2_2%B
x_PM_SKY130_FD_SC_HS__XNOR2_2%A_133_368# N_A_133_368#_M1010_d
+ N_A_133_368#_M1015_d N_A_133_368#_c_392_n N_A_133_368#_M1012_g
+ N_A_133_368#_c_385_n N_A_133_368#_M1001_g N_A_133_368#_c_393_n
+ N_A_133_368#_M1013_g N_A_133_368#_c_386_n N_A_133_368#_M1014_g
+ N_A_133_368#_c_394_n N_A_133_368#_c_387_n N_A_133_368#_c_388_n
+ N_A_133_368#_c_389_n N_A_133_368#_c_390_n N_A_133_368#_c_391_n
+ PM_SKY130_FD_SC_HS__XNOR2_2%A_133_368#
x_PM_SKY130_FD_SC_HS__XNOR2_2%VPWR N_VPWR_M1015_s N_VPWR_M1003_d N_VPWR_M1013_s
+ N_VPWR_M1009_d N_VPWR_c_485_n N_VPWR_c_486_n N_VPWR_c_487_n N_VPWR_c_488_n
+ N_VPWR_c_489_n N_VPWR_c_490_n VPWR N_VPWR_c_491_n N_VPWR_c_492_n
+ N_VPWR_c_493_n N_VPWR_c_494_n N_VPWR_c_484_n PM_SKY130_FD_SC_HS__XNOR2_2%VPWR
x_PM_SKY130_FD_SC_HS__XNOR2_2%Y N_Y_M1001_d N_Y_M1012_d N_Y_M1006_d N_Y_c_551_n
+ N_Y_c_552_n N_Y_c_553_n N_Y_c_569_n N_Y_c_558_n N_Y_c_570_n N_Y_c_554_n
+ N_Y_c_572_n N_Y_c_555_n N_Y_c_556_n N_Y_c_573_n Y Y N_Y_c_574_n
+ PM_SKY130_FD_SC_HS__XNOR2_2%Y
x_PM_SKY130_FD_SC_HS__XNOR2_2%A_638_368# N_A_638_368#_M1008_s
+ N_A_638_368#_M1007_s N_A_638_368#_c_652_n N_A_638_368#_c_659_n
+ N_A_638_368#_c_653_n PM_SKY130_FD_SC_HS__XNOR2_2%A_638_368#
x_PM_SKY130_FD_SC_HS__XNOR2_2%VGND N_VGND_M1011_s N_VGND_M1004_d N_VGND_M1002_s
+ N_VGND_c_679_n N_VGND_c_680_n N_VGND_c_681_n N_VGND_c_682_n N_VGND_c_683_n
+ N_VGND_c_684_n VGND N_VGND_c_685_n N_VGND_c_686_n N_VGND_c_687_n
+ N_VGND_c_688_n PM_SKY130_FD_SC_HS__XNOR2_2%VGND
x_PM_SKY130_FD_SC_HS__XNOR2_2%A_340_107# N_A_340_107#_M1001_s
+ N_A_340_107#_M1014_s N_A_340_107#_M1000_d N_A_340_107#_M1005_s
+ N_A_340_107#_c_747_n N_A_340_107#_c_748_n N_A_340_107#_c_744_n
+ N_A_340_107#_c_745_n N_A_340_107#_c_754_n N_A_340_107#_c_758_n
+ N_A_340_107#_c_746_n PM_SKY130_FD_SC_HS__XNOR2_2%A_340_107#
cc_1 VNB N_A_c_91_n 0.0428131f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.765
cc_2 VNB N_A_c_92_n 0.017864f $X=-0.19 $Y=-0.245 $X2=0.68 $Y2=1.22
cc_3 VNB N_A_c_93_n 0.0396704f $X=-0.19 $Y=-0.245 $X2=3.115 $Y2=1.765
cc_4 VNB N_A_c_94_n 0.0186645f $X=-0.19 $Y=-0.245 $X2=3.135 $Y2=1.22
cc_5 VNB N_A_c_95_n 0.0276464f $X=-0.19 $Y=-0.245 $X2=4.695 $Y2=1.765
cc_6 VNB N_A_M1005_g 0.031366f $X=-0.19 $Y=-0.245 $X2=4.785 $Y2=0.74
cc_7 VNB N_A_c_97_n 0.00126095f $X=-0.19 $Y=-0.245 $X2=3.19 $Y2=1.72
cc_8 VNB A 0.00491569f $X=-0.19 $Y=-0.245 $X2=4.475 $Y2=1.58
cc_9 VNB N_A_c_99_n 0.0212635f $X=-0.19 $Y=-0.245 $X2=2.975 $Y2=1.295
cc_10 VNB N_A_c_100_n 0.00284076f $X=-0.19 $Y=-0.245 $X2=0.865 $Y2=1.295
cc_11 VNB N_A_c_101_n 0.00311998f $X=-0.19 $Y=-0.245 $X2=3.12 $Y2=1.295
cc_12 VNB N_A_c_102_n 0.00526995f $X=-0.19 $Y=-0.245 $X2=3.12 $Y2=1.295
cc_13 VNB N_A_c_103_n 0.00770753f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.385
cc_14 VNB N_B_M1010_g 0.0267022f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=2.34
cc_15 VNB N_B_c_235_n 0.0190023f $X=-0.19 $Y=-0.245 $X2=3.115 $Y2=2.4
cc_16 VNB N_B_c_236_n 0.0181813f $X=-0.19 $Y=-0.245 $X2=4.695 $Y2=2.4
cc_17 VNB N_B_c_237_n 0.0126266f $X=-0.19 $Y=-0.245 $X2=3.19 $Y2=1.72
cc_18 VNB N_B_c_238_n 0.00111425f $X=-0.19 $Y=-0.245 $X2=4.475 $Y2=1.58
cc_19 VNB N_B_c_239_n 0.0372654f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_B_c_240_n 0.0198025f $X=-0.19 $Y=-0.245 $X2=3.12 $Y2=1.295
cc_21 VNB N_B_c_241_n 7.72606e-19 $X=-0.19 $Y=-0.245 $X2=3.12 $Y2=1.295
cc_22 VNB N_B_c_242_n 0.0227111f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.385
cc_23 VNB B 0.00119299f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.385
cc_24 VNB N_B_c_244_n 0.0545105f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_133_368#_c_385_n 0.0206891f $X=-0.19 $Y=-0.245 $X2=3.135 $Y2=1.22
cc_26 VNB N_A_133_368#_c_386_n 0.0190849f $X=-0.19 $Y=-0.245 $X2=4.785 $Y2=1.35
cc_27 VNB N_A_133_368#_c_387_n 0.00311207f $X=-0.19 $Y=-0.245 $X2=4.475 $Y2=1.58
cc_28 VNB N_A_133_368#_c_388_n 0.00644617f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.295
cc_29 VNB N_A_133_368#_c_389_n 0.0075666f $X=-0.19 $Y=-0.245 $X2=3.12 $Y2=1.295
cc_30 VNB N_A_133_368#_c_390_n 0.00974138f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_133_368#_c_391_n 0.0705575f $X=-0.19 $Y=-0.245 $X2=3.19 $Y2=1.385
cc_32 VNB N_VPWR_c_484_n 0.223389f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_Y_c_551_n 0.0311889f $X=-0.19 $Y=-0.245 $X2=3.135 $Y2=0.74
cc_34 VNB N_Y_c_552_n 0.00487916f $X=-0.19 $Y=-0.245 $X2=3.135 $Y2=0.74
cc_35 VNB N_Y_c_553_n 0.00986386f $X=-0.19 $Y=-0.245 $X2=4.695 $Y2=1.765
cc_36 VNB N_Y_c_554_n 5.82374e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_Y_c_555_n 0.00409335f $X=-0.19 $Y=-0.245 $X2=3.355 $Y2=1.805
cc_38 VNB N_Y_c_556_n 0.0148451f $X=-0.19 $Y=-0.245 $X2=4.475 $Y2=1.58
cc_39 VNB N_VGND_c_679_n 0.0131748f $X=-0.19 $Y=-0.245 $X2=3.135 $Y2=1.22
cc_40 VNB N_VGND_c_680_n 0.0273582f $X=-0.19 $Y=-0.245 $X2=3.135 $Y2=0.74
cc_41 VNB N_VGND_c_681_n 0.00800128f $X=-0.19 $Y=-0.245 $X2=4.785 $Y2=1.35
cc_42 VNB N_VGND_c_682_n 0.00812389f $X=-0.19 $Y=-0.245 $X2=3.19 $Y2=1.55
cc_43 VNB N_VGND_c_683_n 0.0656586f $X=-0.19 $Y=-0.245 $X2=3.355 $Y2=1.805
cc_44 VNB N_VGND_c_684_n 0.0064126f $X=-0.19 $Y=-0.245 $X2=4.475 $Y2=1.58
cc_45 VNB N_VGND_c_685_n 0.0190098f $X=-0.19 $Y=-0.245 $X2=3.12 $Y2=1.295
cc_46 VNB N_VGND_c_686_n 0.0193317f $X=-0.19 $Y=-0.245 $X2=3.19 $Y2=1.385
cc_47 VNB N_VGND_c_687_n 0.291439f $X=-0.19 $Y=-0.245 $X2=3.19 $Y2=1.385
cc_48 VNB N_VGND_c_688_n 0.0066048f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A_340_107#_c_744_n 0.00274459f $X=-0.19 $Y=-0.245 $X2=4.445
+ $Y2=1.805
cc_50 VNB N_A_340_107#_c_745_n 0.0024006f $X=-0.19 $Y=-0.245 $X2=4.475 $Y2=1.58
cc_51 VNB N_A_340_107#_c_746_n 0.0136683f $X=-0.19 $Y=-0.245 $X2=3.12 $Y2=1.295
cc_52 VPB N_A_c_91_n 0.0237413f $X=-0.19 $Y=1.66 $X2=0.59 $Y2=1.765
cc_53 VPB N_A_c_93_n 0.0247506f $X=-0.19 $Y=1.66 $X2=3.115 $Y2=1.765
cc_54 VPB N_A_c_95_n 0.0278223f $X=-0.19 $Y=1.66 $X2=4.695 $Y2=1.765
cc_55 VPB N_A_c_97_n 6.82535e-19 $X=-0.19 $Y=1.66 $X2=3.19 $Y2=1.72
cc_56 VPB N_A_c_108_n 0.0175175f $X=-0.19 $Y=1.66 $X2=4.445 $Y2=1.805
cc_57 VPB N_A_c_109_n 9.57272e-19 $X=-0.19 $Y=1.66 $X2=3.355 $Y2=1.805
cc_58 VPB A 0.00150831f $X=-0.19 $Y=1.66 $X2=4.475 $Y2=1.58
cc_59 VPB N_B_c_245_n 0.016212f $X=-0.19 $Y=1.66 $X2=0.68 $Y2=0.74
cc_60 VPB N_B_c_246_n 0.015275f $X=-0.19 $Y=1.66 $X2=3.135 $Y2=0.74
cc_61 VPB N_B_c_247_n 0.0145086f $X=-0.19 $Y=1.66 $X2=4.785 $Y2=0.74
cc_62 VPB N_B_c_237_n 0.00676355f $X=-0.19 $Y=1.66 $X2=3.19 $Y2=1.72
cc_63 VPB N_B_c_238_n 6.80183e-19 $X=-0.19 $Y=1.66 $X2=4.475 $Y2=1.58
cc_64 VPB N_B_c_239_n 0.0165375f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_65 VPB N_B_c_251_n 0.00700242f $X=-0.19 $Y=1.66 $X2=0.865 $Y2=1.295
cc_66 VPB N_B_c_252_n 7.33567e-19 $X=-0.19 $Y=1.66 $X2=0.72 $Y2=1.295
cc_67 VPB N_B_c_253_n 0.0100484f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_68 VPB N_B_c_242_n 0.0168058f $X=-0.19 $Y=1.66 $X2=0.59 $Y2=1.385
cc_69 VPB N_B_c_244_n 0.0130587f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_70 VPB N_A_133_368#_c_392_n 0.0165606f $X=-0.19 $Y=1.66 $X2=3.115 $Y2=1.765
cc_71 VPB N_A_133_368#_c_393_n 0.0162233f $X=-0.19 $Y=1.66 $X2=4.695 $Y2=1.765
cc_72 VPB N_A_133_368#_c_394_n 0.00417671f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_73 VPB N_A_133_368#_c_387_n 0.00109243f $X=-0.19 $Y=1.66 $X2=4.475 $Y2=1.58
cc_74 VPB N_A_133_368#_c_391_n 0.0138569f $X=-0.19 $Y=1.66 $X2=3.19 $Y2=1.385
cc_75 VPB N_VPWR_c_485_n 0.0121909f $X=-0.19 $Y=1.66 $X2=4.695 $Y2=1.765
cc_76 VPB N_VPWR_c_486_n 0.0293161f $X=-0.19 $Y=1.66 $X2=4.695 $Y2=2.4
cc_77 VPB N_VPWR_c_487_n 0.020562f $X=-0.19 $Y=1.66 $X2=4.785 $Y2=0.74
cc_78 VPB N_VPWR_c_488_n 0.00863527f $X=-0.19 $Y=1.66 $X2=3.19 $Y2=1.72
cc_79 VPB N_VPWR_c_489_n 0.0131441f $X=-0.19 $Y=1.66 $X2=3.355 $Y2=1.805
cc_80 VPB N_VPWR_c_490_n 0.034301f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_81 VPB N_VPWR_c_491_n 0.0249485f $X=-0.19 $Y=1.66 $X2=0.72 $Y2=1.295
cc_82 VPB N_VPWR_c_492_n 0.0440036f $X=-0.19 $Y=1.66 $X2=3.12 $Y2=1.295
cc_83 VPB N_VPWR_c_493_n 0.0304202f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_84 VPB N_VPWR_c_494_n 0.00632133f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_85 VPB N_VPWR_c_484_n 0.0718057f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_86 VPB N_Y_c_551_n 0.0264068f $X=-0.19 $Y=1.66 $X2=3.135 $Y2=0.74
cc_87 VPB N_Y_c_558_n 0.00801979f $X=-0.19 $Y=1.66 $X2=4.695 $Y2=2.4
cc_88 VPB Y 0.00257348f $X=-0.19 $Y=1.66 $X2=3.12 $Y2=1.295
cc_89 VPB N_A_638_368#_c_652_n 0.00541183f $X=-0.19 $Y=1.66 $X2=3.115 $Y2=1.765
cc_90 VPB N_A_638_368#_c_653_n 0.00372668f $X=-0.19 $Y=1.66 $X2=4.695 $Y2=2.4
cc_91 N_A_c_92_n N_B_M1010_g 0.0342458f $X=0.68 $Y=1.22 $X2=0 $Y2=0
cc_92 N_A_c_99_n N_B_M1010_g 0.00113884f $X=2.975 $Y=1.295 $X2=0 $Y2=0
cc_93 N_A_c_100_n N_B_M1010_g 6.92697e-19 $X=0.865 $Y=1.295 $X2=0 $Y2=0
cc_94 N_A_c_103_n N_B_M1010_g 0.00207268f $X=0.59 $Y=1.385 $X2=0 $Y2=0
cc_95 N_A_c_91_n N_B_c_245_n 0.0315495f $X=0.59 $Y=1.765 $X2=0 $Y2=0
cc_96 N_A_c_94_n N_B_c_235_n 0.0238678f $X=3.135 $Y=1.22 $X2=0 $Y2=0
cc_97 N_A_c_102_n N_B_c_235_n 3.87669e-19 $X=3.12 $Y=1.295 $X2=0 $Y2=0
cc_98 N_A_c_93_n N_B_c_246_n 0.030742f $X=3.115 $Y=1.765 $X2=0 $Y2=0
cc_99 N_A_c_108_n N_B_c_246_n 0.00744475f $X=4.445 $Y=1.805 $X2=0 $Y2=0
cc_100 N_A_M1005_g N_B_c_236_n 0.0266017f $X=4.785 $Y=0.74 $X2=0 $Y2=0
cc_101 N_A_c_95_n N_B_c_247_n 0.0333918f $X=4.695 $Y=1.765 $X2=0 $Y2=0
cc_102 N_A_c_108_n N_B_c_247_n 0.00706013f $X=4.445 $Y=1.805 $X2=0 $Y2=0
cc_103 N_A_c_91_n N_B_c_237_n 0.0436281f $X=0.59 $Y=1.765 $X2=0 $Y2=0
cc_104 N_A_c_100_n N_B_c_237_n 7.45074e-19 $X=0.865 $Y=1.295 $X2=0 $Y2=0
cc_105 N_A_c_99_n N_B_c_238_n 0.0190018f $X=2.975 $Y=1.295 $X2=0 $Y2=0
cc_106 N_A_c_99_n N_B_c_239_n 0.0113639f $X=2.975 $Y=1.295 $X2=0 $Y2=0
cc_107 N_A_c_93_n N_B_c_251_n 7.99559e-19 $X=3.115 $Y=1.765 $X2=0 $Y2=0
cc_108 N_A_c_109_n N_B_c_251_n 0.0100113f $X=3.355 $Y=1.805 $X2=0 $Y2=0
cc_109 N_A_c_99_n N_B_c_251_n 0.0164056f $X=2.975 $Y=1.295 $X2=0 $Y2=0
cc_110 N_A_c_93_n N_B_c_275_n 0.0033756f $X=3.115 $Y=1.765 $X2=0 $Y2=0
cc_111 N_A_c_93_n N_B_c_253_n 0.0124823f $X=3.115 $Y=1.765 $X2=0 $Y2=0
cc_112 N_A_c_95_n N_B_c_253_n 0.0180765f $X=4.695 $Y=1.765 $X2=0 $Y2=0
cc_113 N_A_c_108_n N_B_c_253_n 0.0610814f $X=4.445 $Y=1.805 $X2=0 $Y2=0
cc_114 N_A_c_109_n N_B_c_253_n 0.0202855f $X=3.355 $Y=1.805 $X2=0 $Y2=0
cc_115 A N_B_c_253_n 0.0193337f $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_116 N_A_c_95_n N_B_c_240_n 0.00129526f $X=4.695 $Y=1.765 $X2=0 $Y2=0
cc_117 N_A_M1005_g N_B_c_240_n 0.01286f $X=4.785 $Y=0.74 $X2=0 $Y2=0
cc_118 N_A_c_108_n N_B_c_240_n 0.00627445f $X=4.445 $Y=1.805 $X2=0 $Y2=0
cc_119 A N_B_c_240_n 0.0314518f $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_120 N_A_c_95_n N_B_c_242_n 0.0093551f $X=4.695 $Y=1.765 $X2=0 $Y2=0
cc_121 N_A_M1005_g N_B_c_242_n 0.0132787f $X=4.785 $Y=0.74 $X2=0 $Y2=0
cc_122 A N_B_c_242_n 0.0348465f $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_123 N_A_c_93_n B 8.71298e-19 $X=3.115 $Y=1.765 $X2=0 $Y2=0
cc_124 N_A_c_95_n B 2.21532e-19 $X=4.695 $Y=1.765 $X2=0 $Y2=0
cc_125 N_A_M1005_g B 9.31443e-19 $X=4.785 $Y=0.74 $X2=0 $Y2=0
cc_126 N_A_c_108_n B 0.0251802f $X=4.445 $Y=1.805 $X2=0 $Y2=0
cc_127 A B 0.0148825f $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_128 N_A_c_102_n B 0.0105933f $X=3.12 $Y=1.295 $X2=0 $Y2=0
cc_129 N_A_c_93_n N_B_c_244_n 0.019199f $X=3.115 $Y=1.765 $X2=0 $Y2=0
cc_130 N_A_c_95_n N_B_c_244_n 0.0191121f $X=4.695 $Y=1.765 $X2=0 $Y2=0
cc_131 N_A_c_97_n N_B_c_244_n 0.00365567f $X=3.19 $Y=1.72 $X2=0 $Y2=0
cc_132 N_A_c_108_n N_B_c_244_n 0.015999f $X=4.445 $Y=1.805 $X2=0 $Y2=0
cc_133 A N_B_c_244_n 0.00553854f $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_134 N_A_c_102_n N_B_c_244_n 0.00162562f $X=3.12 $Y=1.295 $X2=0 $Y2=0
cc_135 N_A_c_93_n N_A_133_368#_c_393_n 0.027089f $X=3.115 $Y=1.765 $X2=0 $Y2=0
cc_136 N_A_c_109_n N_A_133_368#_c_393_n 2.67149e-19 $X=3.355 $Y=1.805 $X2=0
+ $Y2=0
cc_137 N_A_c_94_n N_A_133_368#_c_386_n 0.0132146f $X=3.135 $Y=1.22 $X2=0 $Y2=0
cc_138 N_A_c_101_n N_A_133_368#_c_386_n 6.76195e-19 $X=3.12 $Y=1.295 $X2=0 $Y2=0
cc_139 N_A_c_102_n N_A_133_368#_c_386_n 0.00119559f $X=3.12 $Y=1.295 $X2=0 $Y2=0
cc_140 N_A_c_91_n N_A_133_368#_c_394_n 0.00823039f $X=0.59 $Y=1.765 $X2=0 $Y2=0
cc_141 N_A_c_99_n N_A_133_368#_c_394_n 0.00510089f $X=2.975 $Y=1.295 $X2=0 $Y2=0
cc_142 N_A_c_100_n N_A_133_368#_c_394_n 0.00228802f $X=0.865 $Y=1.295 $X2=0
+ $Y2=0
cc_143 N_A_c_103_n N_A_133_368#_c_394_n 0.00948332f $X=0.59 $Y=1.385 $X2=0 $Y2=0
cc_144 N_A_c_91_n N_A_133_368#_c_387_n 0.00226182f $X=0.59 $Y=1.765 $X2=0 $Y2=0
cc_145 N_A_c_92_n N_A_133_368#_c_387_n 4.6081e-19 $X=0.68 $Y=1.22 $X2=0 $Y2=0
cc_146 N_A_c_99_n N_A_133_368#_c_387_n 0.0262593f $X=2.975 $Y=1.295 $X2=0 $Y2=0
cc_147 N_A_c_100_n N_A_133_368#_c_387_n 0.0026151f $X=0.865 $Y=1.295 $X2=0 $Y2=0
cc_148 N_A_c_103_n N_A_133_368#_c_387_n 0.0261005f $X=0.59 $Y=1.385 $X2=0 $Y2=0
cc_149 N_A_c_92_n N_A_133_368#_c_388_n 0.00147911f $X=0.68 $Y=1.22 $X2=0 $Y2=0
cc_150 N_A_c_99_n N_A_133_368#_c_388_n 0.0130897f $X=2.975 $Y=1.295 $X2=0 $Y2=0
cc_151 N_A_c_93_n N_A_133_368#_c_389_n 4.75044e-19 $X=3.115 $Y=1.765 $X2=0 $Y2=0
cc_152 N_A_c_99_n N_A_133_368#_c_389_n 0.0361112f $X=2.975 $Y=1.295 $X2=0 $Y2=0
cc_153 N_A_c_101_n N_A_133_368#_c_389_n 0.00234524f $X=3.12 $Y=1.295 $X2=0 $Y2=0
cc_154 N_A_c_102_n N_A_133_368#_c_389_n 0.0119148f $X=3.12 $Y=1.295 $X2=0 $Y2=0
cc_155 N_A_c_99_n N_A_133_368#_c_390_n 0.0150674f $X=2.975 $Y=1.295 $X2=0 $Y2=0
cc_156 N_A_c_93_n N_A_133_368#_c_391_n 0.0188805f $X=3.115 $Y=1.765 $X2=0 $Y2=0
cc_157 N_A_c_97_n N_A_133_368#_c_391_n 9.66247e-19 $X=3.19 $Y=1.72 $X2=0 $Y2=0
cc_158 N_A_c_99_n N_A_133_368#_c_391_n 0.0077648f $X=2.975 $Y=1.295 $X2=0 $Y2=0
cc_159 N_A_c_102_n N_A_133_368#_c_391_n 7.12902e-19 $X=3.12 $Y=1.295 $X2=0 $Y2=0
cc_160 N_A_c_91_n N_VPWR_c_486_n 0.0128232f $X=0.59 $Y=1.765 $X2=0 $Y2=0
cc_161 N_A_c_93_n N_VPWR_c_488_n 0.00422112f $X=3.115 $Y=1.765 $X2=0 $Y2=0
cc_162 N_A_c_95_n N_VPWR_c_490_n 0.01421f $X=4.695 $Y=1.765 $X2=0 $Y2=0
cc_163 N_A_c_91_n N_VPWR_c_491_n 0.0049405f $X=0.59 $Y=1.765 $X2=0 $Y2=0
cc_164 N_A_c_93_n N_VPWR_c_492_n 0.00339044f $X=3.115 $Y=1.765 $X2=0 $Y2=0
cc_165 N_A_c_95_n N_VPWR_c_492_n 0.0044313f $X=4.695 $Y=1.765 $X2=0 $Y2=0
cc_166 N_A_c_91_n N_VPWR_c_484_n 0.00508379f $X=0.59 $Y=1.765 $X2=0 $Y2=0
cc_167 N_A_c_93_n N_VPWR_c_484_n 0.00447202f $X=3.115 $Y=1.765 $X2=0 $Y2=0
cc_168 N_A_c_95_n N_VPWR_c_484_n 0.00856934f $X=4.695 $Y=1.765 $X2=0 $Y2=0
cc_169 N_A_c_108_n N_Y_M1006_d 0.00198204f $X=4.445 $Y=1.805 $X2=0 $Y2=0
cc_170 N_A_c_91_n N_Y_c_551_n 0.0225967f $X=0.59 $Y=1.765 $X2=0 $Y2=0
cc_171 N_A_c_92_n N_Y_c_551_n 0.00499812f $X=0.68 $Y=1.22 $X2=0 $Y2=0
cc_172 N_A_c_100_n N_Y_c_551_n 0.00117441f $X=0.865 $Y=1.295 $X2=0 $Y2=0
cc_173 N_A_c_103_n N_Y_c_551_n 0.0273196f $X=0.59 $Y=1.385 $X2=0 $Y2=0
cc_174 N_A_c_91_n N_Y_c_552_n 0.00101288f $X=0.59 $Y=1.765 $X2=0 $Y2=0
cc_175 N_A_c_92_n N_Y_c_552_n 0.0103528f $X=0.68 $Y=1.22 $X2=0 $Y2=0
cc_176 N_A_c_100_n N_Y_c_552_n 0.00665349f $X=0.865 $Y=1.295 $X2=0 $Y2=0
cc_177 N_A_c_103_n N_Y_c_552_n 0.0252708f $X=0.59 $Y=1.385 $X2=0 $Y2=0
cc_178 N_A_c_91_n N_Y_c_569_n 0.0179277f $X=0.59 $Y=1.765 $X2=0 $Y2=0
cc_179 N_A_c_92_n N_Y_c_570_n 0.0132561f $X=0.68 $Y=1.22 $X2=0 $Y2=0
cc_180 N_A_c_92_n N_Y_c_554_n 0.00474295f $X=0.68 $Y=1.22 $X2=0 $Y2=0
cc_181 N_A_c_93_n N_Y_c_572_n 0.0139502f $X=3.115 $Y=1.765 $X2=0 $Y2=0
cc_182 N_A_c_93_n N_Y_c_573_n 7.96419e-19 $X=3.115 $Y=1.765 $X2=0 $Y2=0
cc_183 N_A_c_93_n N_Y_c_574_n 0.001721f $X=3.115 $Y=1.765 $X2=0 $Y2=0
cc_184 N_A_c_108_n N_A_638_368#_M1008_s 0.00298271f $X=4.445 $Y=1.805 $X2=-0.19
+ $Y2=-0.245
cc_185 N_A_c_109_n N_A_638_368#_M1008_s 0.00118857f $X=3.355 $Y=1.805 $X2=-0.19
+ $Y2=-0.245
cc_186 N_A_c_108_n N_A_638_368#_M1007_s 0.00124676f $X=4.445 $Y=1.805 $X2=0
+ $Y2=0
cc_187 A N_A_638_368#_M1007_s 0.00129985f $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_188 N_A_c_95_n N_A_638_368#_c_652_n 0.00336833f $X=4.695 $Y=1.765 $X2=0 $Y2=0
cc_189 N_A_c_95_n N_A_638_368#_c_659_n 0.00520993f $X=4.695 $Y=1.765 $X2=0 $Y2=0
cc_190 N_A_c_93_n N_A_638_368#_c_653_n 0.00386526f $X=3.115 $Y=1.765 $X2=0 $Y2=0
cc_191 N_A_c_92_n N_VGND_c_680_n 0.00928014f $X=0.68 $Y=1.22 $X2=0 $Y2=0
cc_192 N_A_c_94_n N_VGND_c_681_n 0.00418692f $X=3.135 $Y=1.22 $X2=0 $Y2=0
cc_193 N_A_M1005_g N_VGND_c_682_n 0.00460763f $X=4.785 $Y=0.74 $X2=0 $Y2=0
cc_194 N_A_c_92_n N_VGND_c_683_n 0.00351461f $X=0.68 $Y=1.22 $X2=0 $Y2=0
cc_195 N_A_c_94_n N_VGND_c_683_n 0.00324657f $X=3.135 $Y=1.22 $X2=0 $Y2=0
cc_196 N_A_M1005_g N_VGND_c_686_n 0.00327532f $X=4.785 $Y=0.74 $X2=0 $Y2=0
cc_197 N_A_c_92_n N_VGND_c_687_n 0.00401739f $X=0.68 $Y=1.22 $X2=0 $Y2=0
cc_198 N_A_c_94_n N_VGND_c_687_n 0.00411282f $X=3.135 $Y=1.22 $X2=0 $Y2=0
cc_199 N_A_M1005_g N_VGND_c_687_n 0.00418429f $X=4.785 $Y=0.74 $X2=0 $Y2=0
cc_200 N_A_c_99_n N_A_340_107#_c_747_n 0.00521727f $X=2.975 $Y=1.295 $X2=0 $Y2=0
cc_201 N_A_M1005_g N_A_340_107#_c_748_n 0.00984289f $X=4.785 $Y=0.74 $X2=0 $Y2=0
cc_202 N_A_c_99_n N_A_340_107#_c_744_n 0.00314462f $X=2.975 $Y=1.295 $X2=0 $Y2=0
cc_203 N_A_c_94_n N_A_340_107#_c_745_n 0.0103404f $X=3.135 $Y=1.22 $X2=0 $Y2=0
cc_204 N_A_c_99_n N_A_340_107#_c_745_n 0.0107331f $X=2.975 $Y=1.295 $X2=0 $Y2=0
cc_205 N_A_c_101_n N_A_340_107#_c_745_n 0.00234562f $X=3.12 $Y=1.295 $X2=0 $Y2=0
cc_206 N_A_c_102_n N_A_340_107#_c_745_n 0.00358921f $X=3.12 $Y=1.295 $X2=0 $Y2=0
cc_207 N_A_c_93_n N_A_340_107#_c_754_n 6.51786e-19 $X=3.115 $Y=1.765 $X2=0 $Y2=0
cc_208 N_A_c_94_n N_A_340_107#_c_754_n 0.0104775f $X=3.135 $Y=1.22 $X2=0 $Y2=0
cc_209 N_A_c_101_n N_A_340_107#_c_754_n 0.00116104f $X=3.12 $Y=1.295 $X2=0 $Y2=0
cc_210 N_A_c_102_n N_A_340_107#_c_754_n 0.00891553f $X=3.12 $Y=1.295 $X2=0 $Y2=0
cc_211 N_A_c_94_n N_A_340_107#_c_758_n 7.68469e-19 $X=3.135 $Y=1.22 $X2=0 $Y2=0
cc_212 N_A_M1005_g N_A_340_107#_c_758_n 7.40195e-19 $X=4.785 $Y=0.74 $X2=0 $Y2=0
cc_213 N_A_M1005_g N_A_340_107#_c_746_n 0.00520058f $X=4.785 $Y=0.74 $X2=0 $Y2=0
cc_214 N_B_c_251_n N_A_133_368#_c_392_n 0.00885662f $X=2.605 $Y=1.805 $X2=0
+ $Y2=0
cc_215 N_B_c_251_n N_A_133_368#_c_393_n 0.00838209f $X=2.605 $Y=1.805 $X2=0
+ $Y2=0
cc_216 N_B_c_245_n N_A_133_368#_c_394_n 0.0117139f $X=1.085 $Y=1.765 $X2=0 $Y2=0
cc_217 N_B_c_237_n N_A_133_368#_c_394_n 4.8004e-19 $X=1.085 $Y=1.557 $X2=0 $Y2=0
cc_218 N_B_c_252_n N_A_133_368#_c_394_n 0.00404854f $X=1.675 $Y=1.805 $X2=0
+ $Y2=0
cc_219 N_B_M1010_g N_A_133_368#_c_387_n 0.00491928f $X=1.07 $Y=0.74 $X2=0 $Y2=0
cc_220 N_B_c_245_n N_A_133_368#_c_387_n 0.00172764f $X=1.085 $Y=1.765 $X2=0
+ $Y2=0
cc_221 N_B_c_237_n N_A_133_368#_c_387_n 0.0160919f $X=1.085 $Y=1.557 $X2=0 $Y2=0
cc_222 N_B_c_238_n N_A_133_368#_c_387_n 0.0263213f $X=1.51 $Y=1.515 $X2=0 $Y2=0
cc_223 N_B_c_252_n N_A_133_368#_c_387_n 0.00823729f $X=1.675 $Y=1.805 $X2=0
+ $Y2=0
cc_224 N_B_M1010_g N_A_133_368#_c_388_n 0.0171185f $X=1.07 $Y=0.74 $X2=0 $Y2=0
cc_225 N_B_c_238_n N_A_133_368#_c_388_n 0.00706196f $X=1.51 $Y=1.515 $X2=0 $Y2=0
cc_226 N_B_c_239_n N_A_133_368#_c_388_n 0.00720307f $X=1.51 $Y=1.515 $X2=0 $Y2=0
cc_227 N_B_c_238_n N_A_133_368#_c_389_n 0.0117923f $X=1.51 $Y=1.515 $X2=0 $Y2=0
cc_228 N_B_c_239_n N_A_133_368#_c_389_n 8.33861e-19 $X=1.51 $Y=1.515 $X2=0 $Y2=0
cc_229 N_B_c_251_n N_A_133_368#_c_389_n 0.0482043f $X=2.605 $Y=1.805 $X2=0 $Y2=0
cc_230 N_B_M1010_g N_A_133_368#_c_390_n 5.78457e-19 $X=1.07 $Y=0.74 $X2=0 $Y2=0
cc_231 N_B_c_238_n N_A_133_368#_c_390_n 0.0139809f $X=1.51 $Y=1.515 $X2=0 $Y2=0
cc_232 N_B_c_239_n N_A_133_368#_c_390_n 0.00157908f $X=1.51 $Y=1.515 $X2=0 $Y2=0
cc_233 N_B_c_251_n N_A_133_368#_c_390_n 0.00353018f $X=2.605 $Y=1.805 $X2=0
+ $Y2=0
cc_234 N_B_c_238_n N_A_133_368#_c_391_n 0.00241968f $X=1.51 $Y=1.515 $X2=0 $Y2=0
cc_235 N_B_c_239_n N_A_133_368#_c_391_n 0.018056f $X=1.51 $Y=1.515 $X2=0 $Y2=0
cc_236 N_B_c_251_n N_A_133_368#_c_391_n 0.0200172f $X=2.605 $Y=1.805 $X2=0 $Y2=0
cc_237 N_B_c_251_n N_VPWR_M1003_d 0.0041093f $X=2.605 $Y=1.805 $X2=0 $Y2=0
cc_238 N_B_c_252_n N_VPWR_M1003_d 0.00664633f $X=1.675 $Y=1.805 $X2=0 $Y2=0
cc_239 N_B_c_251_n N_VPWR_M1013_s 5.54636e-19 $X=2.605 $Y=1.805 $X2=0 $Y2=0
cc_240 N_B_c_275_n N_VPWR_M1013_s 0.00227421f $X=2.69 $Y=2.06 $X2=0 $Y2=0
cc_241 N_B_c_253_n N_VPWR_M1013_s 0.0107325f $X=5.025 $Y=2.145 $X2=0 $Y2=0
cc_242 N_B_c_328_p N_VPWR_M1013_s 0.00289755f $X=2.775 $Y=2.145 $X2=0 $Y2=0
cc_243 N_B_c_253_n N_VPWR_M1009_d 0.0112985f $X=5.025 $Y=2.145 $X2=0 $Y2=0
cc_244 N_B_c_242_n N_VPWR_M1009_d 0.00374217f $X=5.11 $Y=2.06 $X2=0 $Y2=0
cc_245 N_B_c_253_n N_VPWR_c_490_n 0.0259222f $X=5.025 $Y=2.145 $X2=0 $Y2=0
cc_246 N_B_c_245_n N_VPWR_c_491_n 0.0049405f $X=1.085 $Y=1.765 $X2=0 $Y2=0
cc_247 N_B_c_246_n N_VPWR_c_492_n 0.00278271f $X=3.745 $Y=1.765 $X2=0 $Y2=0
cc_248 N_B_c_247_n N_VPWR_c_492_n 0.00278271f $X=4.195 $Y=1.765 $X2=0 $Y2=0
cc_249 N_B_c_245_n N_VPWR_c_493_n 0.013982f $X=1.085 $Y=1.765 $X2=0 $Y2=0
cc_250 N_B_c_245_n N_VPWR_c_484_n 0.00508379f $X=1.085 $Y=1.765 $X2=0 $Y2=0
cc_251 N_B_c_246_n N_VPWR_c_484_n 0.0035438f $X=3.745 $Y=1.765 $X2=0 $Y2=0
cc_252 N_B_c_247_n N_VPWR_c_484_n 0.00354337f $X=4.195 $Y=1.765 $X2=0 $Y2=0
cc_253 N_B_c_251_n N_Y_M1012_d 0.00197722f $X=2.605 $Y=1.805 $X2=0 $Y2=0
cc_254 N_B_c_253_n N_Y_M1006_d 0.00385637f $X=5.025 $Y=2.145 $X2=0 $Y2=0
cc_255 N_B_M1010_g N_Y_c_552_n 0.00103342f $X=1.07 $Y=0.74 $X2=0 $Y2=0
cc_256 N_B_c_245_n N_Y_c_569_n 0.0141775f $X=1.085 $Y=1.765 $X2=0 $Y2=0
cc_257 N_B_c_239_n N_Y_c_569_n 0.00480167f $X=1.51 $Y=1.515 $X2=0 $Y2=0
cc_258 N_B_c_251_n N_Y_c_569_n 0.0111055f $X=2.605 $Y=1.805 $X2=0 $Y2=0
cc_259 N_B_c_252_n N_Y_c_569_n 0.0132626f $X=1.675 $Y=1.805 $X2=0 $Y2=0
cc_260 N_B_M1010_g N_Y_c_570_n 0.00535018f $X=1.07 $Y=0.74 $X2=0 $Y2=0
cc_261 N_B_c_246_n N_Y_c_572_n 0.0104878f $X=3.745 $Y=1.765 $X2=0 $Y2=0
cc_262 N_B_c_251_n N_Y_c_572_n 0.00373153f $X=2.605 $Y=1.805 $X2=0 $Y2=0
cc_263 N_B_c_253_n N_Y_c_572_n 0.0609726f $X=5.025 $Y=2.145 $X2=0 $Y2=0
cc_264 N_B_c_328_p N_Y_c_572_n 0.0117636f $X=2.775 $Y=2.145 $X2=0 $Y2=0
cc_265 N_B_M1010_g N_Y_c_556_n 0.0114851f $X=1.07 $Y=0.74 $X2=0 $Y2=0
cc_266 N_B_c_246_n N_Y_c_573_n 0.00449851f $X=3.745 $Y=1.765 $X2=0 $Y2=0
cc_267 N_B_c_247_n N_Y_c_573_n 0.00355574f $X=4.195 $Y=1.765 $X2=0 $Y2=0
cc_268 N_B_c_253_n N_Y_c_573_n 0.0162374f $X=5.025 $Y=2.145 $X2=0 $Y2=0
cc_269 N_B_c_251_n N_Y_c_574_n 0.0217519f $X=2.605 $Y=1.805 $X2=0 $Y2=0
cc_270 N_B_c_253_n N_A_638_368#_M1008_s 0.00876881f $X=5.025 $Y=2.145 $X2=-0.19
+ $Y2=-0.245
cc_271 N_B_c_253_n N_A_638_368#_M1007_s 0.0049608f $X=5.025 $Y=2.145 $X2=0 $Y2=0
cc_272 N_B_c_246_n N_A_638_368#_c_652_n 0.00963532f $X=3.745 $Y=1.765 $X2=0
+ $Y2=0
cc_273 N_B_c_247_n N_A_638_368#_c_652_n 0.0116689f $X=4.195 $Y=1.765 $X2=0 $Y2=0
cc_274 N_B_c_253_n N_A_638_368#_c_652_n 0.00292982f $X=5.025 $Y=2.145 $X2=0
+ $Y2=0
cc_275 N_B_c_253_n N_A_638_368#_c_659_n 0.0202127f $X=5.025 $Y=2.145 $X2=0 $Y2=0
cc_276 N_B_c_246_n N_A_638_368#_c_653_n 0.0052941f $X=3.745 $Y=1.765 $X2=0 $Y2=0
cc_277 N_B_c_240_n N_VGND_M1002_s 0.0041543f $X=5.025 $Y=1.095 $X2=0 $Y2=0
cc_278 N_B_c_235_n N_VGND_c_681_n 0.00455846f $X=3.73 $Y=1.22 $X2=0 $Y2=0
cc_279 N_B_c_236_n N_VGND_c_682_n 0.00460763f $X=4.18 $Y=1.22 $X2=0 $Y2=0
cc_280 N_B_M1010_g N_VGND_c_683_n 0.00278271f $X=1.07 $Y=0.74 $X2=0 $Y2=0
cc_281 N_B_c_235_n N_VGND_c_685_n 0.00326539f $X=3.73 $Y=1.22 $X2=0 $Y2=0
cc_282 N_B_c_236_n N_VGND_c_685_n 0.00329249f $X=4.18 $Y=1.22 $X2=0 $Y2=0
cc_283 N_B_M1010_g N_VGND_c_687_n 0.00358137f $X=1.07 $Y=0.74 $X2=0 $Y2=0
cc_284 N_B_c_235_n N_VGND_c_687_n 0.00416026f $X=3.73 $Y=1.22 $X2=0 $Y2=0
cc_285 N_B_c_236_n N_VGND_c_687_n 0.00421564f $X=4.18 $Y=1.22 $X2=0 $Y2=0
cc_286 N_B_c_241_n N_A_340_107#_M1000_d 0.00267476f $X=4.255 $Y=1.095 $X2=0
+ $Y2=0
cc_287 N_B_c_240_n N_A_340_107#_M1005_s 0.00246551f $X=5.025 $Y=1.095 $X2=0
+ $Y2=0
cc_288 N_B_c_236_n N_A_340_107#_c_748_n 0.0102985f $X=4.18 $Y=1.22 $X2=0 $Y2=0
cc_289 N_B_c_240_n N_A_340_107#_c_748_n 0.0332405f $X=5.025 $Y=1.095 $X2=0 $Y2=0
cc_290 N_B_M1010_g N_A_340_107#_c_744_n 6.43207e-19 $X=1.07 $Y=0.74 $X2=0 $Y2=0
cc_291 N_B_c_235_n N_A_340_107#_c_745_n 0.00164705f $X=3.73 $Y=1.22 $X2=0 $Y2=0
cc_292 N_B_c_235_n N_A_340_107#_c_754_n 0.0130102f $X=3.73 $Y=1.22 $X2=0 $Y2=0
cc_293 N_B_c_235_n N_A_340_107#_c_758_n 0.00555908f $X=3.73 $Y=1.22 $X2=0 $Y2=0
cc_294 N_B_c_236_n N_A_340_107#_c_758_n 0.00346836f $X=4.18 $Y=1.22 $X2=0 $Y2=0
cc_295 N_B_c_241_n N_A_340_107#_c_758_n 0.0214926f $X=4.255 $Y=1.095 $X2=0 $Y2=0
cc_296 N_B_c_244_n N_A_340_107#_c_758_n 0.00149766f $X=4.18 $Y=1.492 $X2=0 $Y2=0
cc_297 N_B_c_236_n N_A_340_107#_c_746_n 8.44873e-19 $X=4.18 $Y=1.22 $X2=0 $Y2=0
cc_298 N_B_c_240_n N_A_340_107#_c_746_n 0.022058f $X=5.025 $Y=1.095 $X2=0 $Y2=0
cc_299 N_A_133_368#_c_392_n N_VPWR_c_487_n 0.00377622f $X=2.045 $Y=1.765 $X2=0
+ $Y2=0
cc_300 N_A_133_368#_c_393_n N_VPWR_c_487_n 0.00335424f $X=2.495 $Y=1.765 $X2=0
+ $Y2=0
cc_301 N_A_133_368#_c_393_n N_VPWR_c_488_n 0.00555772f $X=2.495 $Y=1.765 $X2=0
+ $Y2=0
cc_302 N_A_133_368#_c_392_n N_VPWR_c_493_n 0.00625366f $X=2.045 $Y=1.765 $X2=0
+ $Y2=0
cc_303 N_A_133_368#_c_392_n N_VPWR_c_484_n 0.00415962f $X=2.045 $Y=1.765 $X2=0
+ $Y2=0
cc_304 N_A_133_368#_c_393_n N_VPWR_c_484_n 0.00436232f $X=2.495 $Y=1.765 $X2=0
+ $Y2=0
cc_305 N_A_133_368#_c_389_n N_Y_M1001_d 0.00456646f $X=2.42 $Y=1.385 $X2=-0.19
+ $Y2=-0.245
cc_306 N_A_133_368#_c_394_n N_Y_c_551_n 0.0131596f $X=1.005 $Y=1.985 $X2=0 $Y2=0
cc_307 N_A_133_368#_c_388_n N_Y_c_552_n 0.0143386f $X=1.285 $Y=0.8 $X2=0 $Y2=0
cc_308 N_A_133_368#_M1015_d N_Y_c_569_n 0.00710579f $X=0.665 $Y=1.84 $X2=0 $Y2=0
cc_309 N_A_133_368#_c_392_n N_Y_c_569_n 0.00941017f $X=2.045 $Y=1.765 $X2=0
+ $Y2=0
cc_310 N_A_133_368#_c_394_n N_Y_c_569_n 0.0300713f $X=1.005 $Y=1.985 $X2=0 $Y2=0
cc_311 N_A_133_368#_c_388_n N_Y_c_570_n 0.0154603f $X=1.285 $Y=0.8 $X2=0 $Y2=0
cc_312 N_A_133_368#_c_393_n N_Y_c_572_n 0.0125032f $X=2.495 $Y=1.765 $X2=0 $Y2=0
cc_313 N_A_133_368#_c_386_n N_Y_c_555_n 0.00431131f $X=2.705 $Y=1.22 $X2=0 $Y2=0
cc_314 N_A_133_368#_M1010_d N_Y_c_556_n 0.00245749f $X=1.145 $Y=0.37 $X2=0 $Y2=0
cc_315 N_A_133_368#_c_385_n N_Y_c_556_n 0.0123292f $X=2.06 $Y=1.22 $X2=0 $Y2=0
cc_316 N_A_133_368#_c_388_n N_Y_c_556_n 0.0236434f $X=1.285 $Y=0.8 $X2=0 $Y2=0
cc_317 N_A_133_368#_c_390_n N_Y_c_556_n 0.00734058f $X=1.915 $Y=1.28 $X2=0 $Y2=0
cc_318 N_A_133_368#_c_392_n Y 0.00974081f $X=2.045 $Y=1.765 $X2=0 $Y2=0
cc_319 N_A_133_368#_c_393_n Y 0.00641749f $X=2.495 $Y=1.765 $X2=0 $Y2=0
cc_320 N_A_133_368#_c_392_n N_Y_c_574_n 0.0192205f $X=2.045 $Y=1.765 $X2=0 $Y2=0
cc_321 N_A_133_368#_c_393_n N_Y_c_574_n 0.00609044f $X=2.495 $Y=1.765 $X2=0
+ $Y2=0
cc_322 N_A_133_368#_c_385_n N_VGND_c_683_n 0.00278271f $X=2.06 $Y=1.22 $X2=0
+ $Y2=0
cc_323 N_A_133_368#_c_386_n N_VGND_c_683_n 0.00324657f $X=2.705 $Y=1.22 $X2=0
+ $Y2=0
cc_324 N_A_133_368#_c_385_n N_VGND_c_687_n 0.00360197f $X=2.06 $Y=1.22 $X2=0
+ $Y2=0
cc_325 N_A_133_368#_c_386_n N_VGND_c_687_n 0.00412609f $X=2.705 $Y=1.22 $X2=0
+ $Y2=0
cc_326 N_A_133_368#_c_390_n N_A_340_107#_M1001_s 0.0020198f $X=1.915 $Y=1.28
+ $X2=-0.19 $Y2=-0.245
cc_327 N_A_133_368#_c_385_n N_A_340_107#_c_747_n 0.00868583f $X=2.06 $Y=1.22
+ $X2=0 $Y2=0
cc_328 N_A_133_368#_c_386_n N_A_340_107#_c_747_n 0.0106562f $X=2.705 $Y=1.22
+ $X2=0 $Y2=0
cc_329 N_A_133_368#_c_389_n N_A_340_107#_c_747_n 0.0285439f $X=2.42 $Y=1.385
+ $X2=0 $Y2=0
cc_330 N_A_133_368#_c_391_n N_A_340_107#_c_747_n 0.00135087f $X=2.495 $Y=1.492
+ $X2=0 $Y2=0
cc_331 N_A_133_368#_c_385_n N_A_340_107#_c_744_n 0.00263714f $X=2.06 $Y=1.22
+ $X2=0 $Y2=0
cc_332 N_A_133_368#_c_386_n N_A_340_107#_c_744_n 3.24573e-19 $X=2.705 $Y=1.22
+ $X2=0 $Y2=0
cc_333 N_A_133_368#_c_388_n N_A_340_107#_c_744_n 0.0147768f $X=1.285 $Y=0.8
+ $X2=0 $Y2=0
cc_334 N_A_133_368#_c_390_n N_A_340_107#_c_744_n 0.0285439f $X=1.915 $Y=1.28
+ $X2=0 $Y2=0
cc_335 N_A_133_368#_c_391_n N_A_340_107#_c_744_n 2.19227e-19 $X=2.495 $Y=1.492
+ $X2=0 $Y2=0
cc_336 N_A_133_368#_c_385_n N_A_340_107#_c_745_n 0.00164025f $X=2.06 $Y=1.22
+ $X2=0 $Y2=0
cc_337 N_A_133_368#_c_386_n N_A_340_107#_c_745_n 0.0106998f $X=2.705 $Y=1.22
+ $X2=0 $Y2=0
cc_338 N_VPWR_M1015_s N_Y_c_551_n 0.00907364f $X=0.135 $Y=1.84 $X2=0 $Y2=0
cc_339 N_VPWR_M1015_s N_Y_c_569_n 0.0106949f $X=0.135 $Y=1.84 $X2=0 $Y2=0
cc_340 N_VPWR_M1003_d N_Y_c_569_n 0.0230565f $X=1.16 $Y=1.84 $X2=0 $Y2=0
cc_341 N_VPWR_c_486_n N_Y_c_569_n 0.0150052f $X=0.28 $Y=2.825 $X2=0 $Y2=0
cc_342 N_VPWR_c_493_n N_Y_c_569_n 0.0511674f $X=1.79 $Y=2.825 $X2=0 $Y2=0
cc_343 N_VPWR_c_484_n N_Y_c_569_n 0.0342201f $X=5.04 $Y=3.33 $X2=0 $Y2=0
cc_344 N_VPWR_M1015_s N_Y_c_558_n 0.00242814f $X=0.135 $Y=1.84 $X2=0 $Y2=0
cc_345 N_VPWR_c_486_n N_Y_c_558_n 0.0122531f $X=0.28 $Y=2.825 $X2=0 $Y2=0
cc_346 N_VPWR_c_484_n N_Y_c_558_n 0.00170605f $X=5.04 $Y=3.33 $X2=0 $Y2=0
cc_347 N_VPWR_M1013_s N_Y_c_572_n 0.00874225f $X=2.57 $Y=1.84 $X2=0 $Y2=0
cc_348 N_VPWR_c_487_n N_Y_c_572_n 0.00224782f $X=2.64 $Y=3.33 $X2=0 $Y2=0
cc_349 N_VPWR_c_488_n N_Y_c_572_n 0.0258802f $X=2.805 $Y=2.905 $X2=0 $Y2=0
cc_350 N_VPWR_c_492_n N_Y_c_572_n 0.00304065f $X=4.805 $Y=3.33 $X2=0 $Y2=0
cc_351 N_VPWR_c_484_n N_Y_c_572_n 0.0137974f $X=5.04 $Y=3.33 $X2=0 $Y2=0
cc_352 N_VPWR_c_487_n Y 0.0170499f $X=2.64 $Y=3.33 $X2=0 $Y2=0
cc_353 N_VPWR_c_488_n Y 0.0163626f $X=2.805 $Y=2.905 $X2=0 $Y2=0
cc_354 N_VPWR_c_493_n Y 0.0265327f $X=1.79 $Y=2.825 $X2=0 $Y2=0
cc_355 N_VPWR_c_484_n Y 0.0139057f $X=5.04 $Y=3.33 $X2=0 $Y2=0
cc_356 N_VPWR_c_490_n N_A_638_368#_c_652_n 0.0119239f $X=4.97 $Y=2.485 $X2=0
+ $Y2=0
cc_357 N_VPWR_c_492_n N_A_638_368#_c_652_n 0.0681033f $X=4.805 $Y=3.33 $X2=0
+ $Y2=0
cc_358 N_VPWR_c_484_n N_A_638_368#_c_652_n 0.0378958f $X=5.04 $Y=3.33 $X2=0
+ $Y2=0
cc_359 N_VPWR_c_488_n N_A_638_368#_c_653_n 0.0185433f $X=2.805 $Y=2.905 $X2=0
+ $Y2=0
cc_360 N_VPWR_c_492_n N_A_638_368#_c_653_n 0.0229944f $X=4.805 $Y=3.33 $X2=0
+ $Y2=0
cc_361 N_VPWR_c_484_n N_A_638_368#_c_653_n 0.012911f $X=5.04 $Y=3.33 $X2=0 $Y2=0
cc_362 N_Y_c_572_n N_A_638_368#_M1008_s 0.00899578f $X=3.805 $Y=2.485 $X2=-0.19
+ $Y2=-0.245
cc_363 N_Y_M1006_d N_A_638_368#_c_652_n 0.00197722f $X=3.82 $Y=1.84 $X2=0 $Y2=0
cc_364 N_Y_c_572_n N_A_638_368#_c_652_n 0.0051463f $X=3.805 $Y=2.485 $X2=0 $Y2=0
cc_365 N_Y_c_573_n N_A_638_368#_c_652_n 0.015244f $X=3.97 $Y=2.485 $X2=0 $Y2=0
cc_366 N_Y_c_572_n N_A_638_368#_c_653_n 0.0251737f $X=3.805 $Y=2.485 $X2=0 $Y2=0
cc_367 N_Y_c_552_n N_VGND_M1011_s 0.00690923f $X=0.665 $Y=0.925 $X2=-0.19
+ $Y2=-0.245
cc_368 N_Y_c_552_n N_VGND_c_680_n 0.0192864f $X=0.665 $Y=0.925 $X2=0 $Y2=0
cc_369 N_Y_c_553_n N_VGND_c_680_n 0.0127101f $X=0.255 $Y=0.925 $X2=0 $Y2=0
cc_370 N_Y_c_570_n N_VGND_c_680_n 0.0183033f $X=0.75 $Y=0.84 $X2=0 $Y2=0
cc_371 N_Y_c_554_n N_VGND_c_680_n 0.0143324f $X=0.835 $Y=0.34 $X2=0 $Y2=0
cc_372 N_Y_c_554_n N_VGND_c_683_n 0.0118705f $X=0.835 $Y=0.34 $X2=0 $Y2=0
cc_373 N_Y_c_556_n N_VGND_c_683_n 0.111797f $X=2.19 $Y=0.377 $X2=0 $Y2=0
cc_374 N_Y_c_552_n N_VGND_c_687_n 0.00623186f $X=0.665 $Y=0.925 $X2=0 $Y2=0
cc_375 N_Y_c_553_n N_VGND_c_687_n 0.00172823f $X=0.255 $Y=0.925 $X2=0 $Y2=0
cc_376 N_Y_c_554_n N_VGND_c_687_n 0.0061974f $X=0.835 $Y=0.34 $X2=0 $Y2=0
cc_377 N_Y_c_556_n N_VGND_c_687_n 0.0641627f $X=2.19 $Y=0.377 $X2=0 $Y2=0
cc_378 N_Y_c_552_n A_151_74# 0.00170774f $X=0.665 $Y=0.925 $X2=-0.19 $Y2=-0.245
cc_379 N_Y_c_570_n A_151_74# 0.00411005f $X=0.75 $Y=0.84 $X2=-0.19 $Y2=-0.245
cc_380 N_Y_c_556_n A_151_74# 0.00389187f $X=2.19 $Y=0.377 $X2=-0.19 $Y2=-0.245
cc_381 N_Y_c_556_n N_A_340_107#_M1001_s 0.00226585f $X=2.19 $Y=0.377 $X2=-0.19
+ $Y2=-0.245
cc_382 N_Y_M1001_d N_A_340_107#_c_747_n 0.00860281f $X=2.135 $Y=0.37 $X2=0 $Y2=0
cc_383 N_Y_c_555_n N_A_340_107#_c_747_n 0.0271762f $X=2.38 $Y=0.415 $X2=0 $Y2=0
cc_384 N_Y_c_556_n N_A_340_107#_c_747_n 0.00570513f $X=2.19 $Y=0.377 $X2=0 $Y2=0
cc_385 N_Y_c_556_n N_A_340_107#_c_744_n 0.0191024f $X=2.19 $Y=0.377 $X2=0 $Y2=0
cc_386 N_Y_c_555_n N_A_340_107#_c_745_n 0.00621476f $X=2.38 $Y=0.415 $X2=0 $Y2=0
cc_387 N_VGND_c_683_n N_A_340_107#_c_747_n 0.00237563f $X=3.265 $Y=0 $X2=0 $Y2=0
cc_388 N_VGND_c_687_n N_A_340_107#_c_747_n 0.00549522f $X=5.04 $Y=0 $X2=0 $Y2=0
cc_389 N_VGND_M1002_s N_A_340_107#_c_748_n 0.00787506f $X=4.255 $Y=0.37 $X2=0
+ $Y2=0
cc_390 N_VGND_c_682_n N_A_340_107#_c_748_n 0.0262746f $X=4.48 $Y=0.335 $X2=0
+ $Y2=0
cc_391 N_VGND_c_685_n N_A_340_107#_c_748_n 0.00266206f $X=4.31 $Y=0 $X2=0 $Y2=0
cc_392 N_VGND_c_686_n N_A_340_107#_c_748_n 0.0023667f $X=5.04 $Y=0 $X2=0 $Y2=0
cc_393 N_VGND_c_687_n N_A_340_107#_c_748_n 0.0107342f $X=5.04 $Y=0 $X2=0 $Y2=0
cc_394 N_VGND_c_681_n N_A_340_107#_c_745_n 0.00613715f $X=3.43 $Y=0.335 $X2=0
+ $Y2=0
cc_395 N_VGND_c_683_n N_A_340_107#_c_745_n 0.0144609f $X=3.265 $Y=0 $X2=0 $Y2=0
cc_396 N_VGND_c_687_n N_A_340_107#_c_745_n 0.0118703f $X=5.04 $Y=0 $X2=0 $Y2=0
cc_397 N_VGND_M1004_d N_A_340_107#_c_754_n 0.0145608f $X=3.21 $Y=0.37 $X2=0
+ $Y2=0
cc_398 N_VGND_c_681_n N_A_340_107#_c_754_n 0.0255041f $X=3.43 $Y=0.335 $X2=0
+ $Y2=0
cc_399 N_VGND_c_683_n N_A_340_107#_c_754_n 0.0023667f $X=3.265 $Y=0 $X2=0 $Y2=0
cc_400 N_VGND_c_685_n N_A_340_107#_c_754_n 0.00236055f $X=4.31 $Y=0 $X2=0 $Y2=0
cc_401 N_VGND_c_687_n N_A_340_107#_c_754_n 0.0102361f $X=5.04 $Y=0 $X2=0 $Y2=0
cc_402 N_VGND_c_685_n N_A_340_107#_c_758_n 0.00723046f $X=4.31 $Y=0 $X2=0 $Y2=0
cc_403 N_VGND_c_687_n N_A_340_107#_c_758_n 0.0106441f $X=5.04 $Y=0 $X2=0 $Y2=0
cc_404 N_VGND_c_686_n N_A_340_107#_c_746_n 0.00789542f $X=5.04 $Y=0 $X2=0 $Y2=0
cc_405 N_VGND_c_687_n N_A_340_107#_c_746_n 0.0106304f $X=5.04 $Y=0 $X2=0 $Y2=0
