* File: sky130_fd_sc_hs__and3_4.pex.spice
* Created: Thu Aug 27 20:32:30 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HS__AND3_4%A_83_260# 1 2 3 4 13 15 18 22 24 26 29 31 33
+ 36 38 40 41 48 50 51 52 55 57 61 63 67 71 73 74 75 78 79 80 81
c177 73 0 1.40226e-19 $X=5.455 $Y=1.195
c178 48 0 1.82661e-19 $X=1.88 $Y=1.465
c179 36 0 1.59824e-19 $X=1.87 $Y=0.74
r180 88 89 45.2262 $w=3.89e-07 $l=3.65e-07 $layer=POLY_cond $X=1.505 $Y=1.532
+ $X2=1.87 $Y2=1.532
r181 87 88 8.05398 $w=3.89e-07 $l=6.5e-08 $layer=POLY_cond $X=1.44 $Y=1.532
+ $X2=1.505 $Y2=1.532
r182 84 85 1.85861 $w=3.89e-07 $l=1.5e-08 $layer=POLY_cond $X=0.94 $Y=1.532
+ $X2=0.955 $Y2=1.532
r183 83 84 53.2802 $w=3.89e-07 $l=4.3e-07 $layer=POLY_cond $X=0.51 $Y=1.532
+ $X2=0.94 $Y2=1.532
r184 82 83 0.619537 $w=3.89e-07 $l=5e-09 $layer=POLY_cond $X=0.505 $Y=1.532
+ $X2=0.51 $Y2=1.532
r185 77 78 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.54 $Y=1.28
+ $X2=5.54 $Y2=1.95
r186 76 81 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.145 $Y=2.035
+ $X2=4.98 $Y2=2.035
r187 75 78 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.455 $Y=2.035
+ $X2=5.54 $Y2=1.95
r188 75 76 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=5.455 $Y=2.035
+ $X2=5.145 $Y2=2.035
r189 73 77 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.455 $Y=1.195
+ $X2=5.54 $Y2=1.28
r190 73 74 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=5.455 $Y=1.195
+ $X2=5.14 $Y2=1.195
r191 69 81 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.98 $Y=2.12
+ $X2=4.98 $Y2=2.035
r192 69 71 5.06376 $w=3.28e-07 $l=1.45e-07 $layer=LI1_cond $X=4.98 $Y=2.12
+ $X2=4.98 $Y2=2.265
r193 65 74 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.975 $Y=1.11
+ $X2=5.14 $Y2=1.195
r194 65 67 12.2229 $w=3.28e-07 $l=3.5e-07 $layer=LI1_cond $X=4.975 $Y=1.11
+ $X2=4.975 $Y2=0.76
r195 64 80 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.145 $Y=2.035
+ $X2=3.98 $Y2=2.035
r196 63 81 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.815 $Y=2.035
+ $X2=4.98 $Y2=2.035
r197 63 64 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.815 $Y=2.035
+ $X2=4.145 $Y2=2.035
r198 59 80 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.98 $Y=2.12
+ $X2=3.98 $Y2=2.035
r199 59 61 5.06376 $w=3.28e-07 $l=1.45e-07 $layer=LI1_cond $X=3.98 $Y=2.12
+ $X2=3.98 $Y2=2.265
r200 58 79 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.895 $Y=2.035
+ $X2=2.73 $Y2=2.035
r201 57 80 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.815 $Y=2.035
+ $X2=3.98 $Y2=2.035
r202 57 58 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=3.815 $Y=2.035
+ $X2=2.895 $Y2=2.035
r203 53 79 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.73 $Y=2.12
+ $X2=2.73 $Y2=2.035
r204 53 55 5.06376 $w=3.28e-07 $l=1.45e-07 $layer=LI1_cond $X=2.73 $Y=2.12
+ $X2=2.73 $Y2=2.265
r205 51 79 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.565 $Y=2.035
+ $X2=2.73 $Y2=2.035
r206 51 52 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=2.565 $Y=2.035
+ $X2=2.235 $Y2=2.035
r207 50 52 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.15 $Y=1.95
+ $X2=2.235 $Y2=2.035
r208 49 50 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=2.15 $Y=1.63
+ $X2=2.15 $Y2=1.95
r209 48 91 9.29306 $w=3.89e-07 $l=7.5e-08 $layer=POLY_cond $X=1.88 $Y=1.532
+ $X2=1.955 $Y2=1.532
r210 48 89 1.23907 $w=3.89e-07 $l=1e-08 $layer=POLY_cond $X=1.88 $Y=1.532
+ $X2=1.87 $Y2=1.532
r211 47 48 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.88
+ $Y=1.465 $X2=1.88 $Y2=1.465
r212 44 87 29.7378 $w=3.89e-07 $l=2.4e-07 $layer=POLY_cond $X=1.2 $Y=1.532
+ $X2=1.44 $Y2=1.532
r213 44 85 30.3573 $w=3.89e-07 $l=2.45e-07 $layer=POLY_cond $X=1.2 $Y=1.532
+ $X2=0.955 $Y2=1.532
r214 43 47 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=1.2 $Y=1.465
+ $X2=1.88 $Y2=1.465
r215 43 44 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.2
+ $Y=1.465 $X2=1.2 $Y2=1.465
r216 41 49 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.065 $Y=1.465
+ $X2=2.15 $Y2=1.63
r217 41 47 6.46067 $w=3.28e-07 $l=1.85e-07 $layer=LI1_cond $X=2.065 $Y=1.465
+ $X2=1.88 $Y2=1.465
r218 38 91 25.1816 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=1.955 $Y=1.765
+ $X2=1.955 $Y2=1.532
r219 38 40 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.955 $Y=1.765
+ $X2=1.955 $Y2=2.4
r220 34 89 25.1816 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=1.87 $Y=1.3
+ $X2=1.87 $Y2=1.532
r221 34 36 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=1.87 $Y=1.3
+ $X2=1.87 $Y2=0.74
r222 31 88 25.1816 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=1.505 $Y=1.765
+ $X2=1.505 $Y2=1.532
r223 31 33 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.505 $Y=1.765
+ $X2=1.505 $Y2=2.4
r224 27 87 25.1816 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=1.44 $Y=1.3
+ $X2=1.44 $Y2=1.532
r225 27 29 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=1.44 $Y=1.3
+ $X2=1.44 $Y2=0.74
r226 24 85 25.1816 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=0.955 $Y=1.765
+ $X2=0.955 $Y2=1.532
r227 24 26 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.955 $Y=1.765
+ $X2=0.955 $Y2=2.4
r228 20 84 25.1816 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=0.94 $Y=1.3
+ $X2=0.94 $Y2=1.532
r229 20 22 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=0.94 $Y=1.3
+ $X2=0.94 $Y2=0.74
r230 16 83 25.1816 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=0.51 $Y=1.3
+ $X2=0.51 $Y2=1.532
r231 16 18 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=0.51 $Y=1.3
+ $X2=0.51 $Y2=0.74
r232 13 82 25.1816 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=0.505 $Y=1.765
+ $X2=0.505 $Y2=1.532
r233 13 15 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.505 $Y=1.765
+ $X2=0.505 $Y2=2.4
r234 4 71 300 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=2 $X=4.83
+ $Y=2.12 $X2=4.98 $Y2=2.265
r235 3 61 300 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=2 $X=3.83
+ $Y=2.12 $X2=3.98 $Y2=2.265
r236 2 55 300 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=2 $X=2.58
+ $Y=2.12 $X2=2.73 $Y2=2.265
r237 1 67 182 $w=1.7e-07 $l=4.83735e-07 $layer=licon1_NDIFF $count=1 $X=4.765
+ $Y=0.37 $X2=4.975 $Y2=0.76
.ends

.subckt PM_SKY130_FD_SC_HS__AND3_4%C 3 6 7 9 12 15 16 18 19 20 26
c66 20 0 1.82661e-19 $X=3.12 $Y=1.665
c67 12 0 1.44963e-19 $X=2.8 $Y=0.69
c68 6 0 4.56703e-20 $X=2.505 $Y=1.955
r69 28 29 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.03
+ $Y=1.615 $X2=3.03 $Y2=1.615
r70 26 28 11.8137 $w=3.06e-07 $l=7.5e-08 $layer=POLY_cond $X=2.955 $Y=1.615
+ $X2=3.03 $Y2=1.615
r71 25 26 24.415 $w=3.06e-07 $l=1.55e-07 $layer=POLY_cond $X=2.8 $Y=1.615
+ $X2=2.955 $Y2=1.615
r72 24 25 46.4673 $w=3.06e-07 $l=2.95e-07 $layer=POLY_cond $X=2.505 $Y=1.615
+ $X2=2.8 $Y2=1.615
r73 20 29 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=3.12 $Y=1.615 $X2=3.03
+ $Y2=1.615
r74 19 29 13.6198 $w=3.28e-07 $l=3.9e-07 $layer=LI1_cond $X=2.64 $Y=1.615
+ $X2=3.03 $Y2=1.615
r75 16 18 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=2.955 $Y=2.045
+ $X2=2.955 $Y2=2.54
r76 15 16 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=2.955 $Y=1.955
+ $X2=2.955 $Y2=2.045
r77 14 26 15.178 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=2.955 $Y=1.78
+ $X2=2.955 $Y2=1.615
r78 14 15 68.0242 $w=1.8e-07 $l=1.75e-07 $layer=POLY_cond $X=2.955 $Y=1.78
+ $X2=2.955 $Y2=1.955
r79 10 25 19.4347 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.8 $Y=1.45 $X2=2.8
+ $Y2=1.615
r80 10 12 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=2.8 $Y=1.45 $X2=2.8
+ $Y2=0.69
r81 7 9 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=2.505 $Y=2.045
+ $X2=2.505 $Y2=2.54
r82 6 7 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=2.505 $Y=1.955 $X2=2.505
+ $Y2=2.045
r83 5 24 15.178 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=2.505 $Y=1.78
+ $X2=2.505 $Y2=1.615
r84 5 6 68.0242 $w=1.8e-07 $l=1.75e-07 $layer=POLY_cond $X=2.505 $Y=1.78
+ $X2=2.505 $Y2=1.955
r85 1 24 21.2647 $w=3.06e-07 $l=2.22486e-07 $layer=POLY_cond $X=2.37 $Y=1.45
+ $X2=2.505 $Y2=1.615
r86 1 3 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=2.37 $Y=1.45 $X2=2.37
+ $Y2=0.69
.ends

.subckt PM_SKY130_FD_SC_HS__AND3_4%B 2 3 5 8 11 12 14 17 19 20 28 30
c63 11 0 7.64129e-20 $X=4.245 $Y=1.955
c64 2 0 7.64129e-20 $X=3.755 $Y=1.955
r65 29 30 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=4.245 $Y=1.49
+ $X2=4.26 $Y2=1.49
r66 27 29 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=4.17 $Y=1.49
+ $X2=4.245 $Y2=1.49
r67 27 28 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.17
+ $Y=1.49 $X2=4.17 $Y2=1.49
r68 25 27 66.4473 $w=3.3e-07 $l=3.8e-07 $layer=POLY_cond $X=3.79 $Y=1.49
+ $X2=4.17 $Y2=1.49
r69 23 25 6.12014 $w=3.3e-07 $l=3.5e-08 $layer=POLY_cond $X=3.755 $Y=1.49
+ $X2=3.79 $Y2=1.49
r70 20 28 2.36587 $w=4.53e-07 $l=9e-08 $layer=LI1_cond $X=4.08 $Y=1.552 $X2=4.17
+ $Y2=1.552
r71 19 20 12.618 $w=4.53e-07 $l=4.8e-07 $layer=LI1_cond $X=3.6 $Y=1.552 $X2=4.08
+ $Y2=1.552
r72 15 30 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.26 $Y=1.325
+ $X2=4.26 $Y2=1.49
r73 15 17 325.606 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=4.26 $Y=1.325
+ $X2=4.26 $Y2=0.69
r74 12 14 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=4.245 $Y=2.045
+ $X2=4.245 $Y2=2.54
r75 11 12 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=4.245 $Y=1.955
+ $X2=4.245 $Y2=2.045
r76 10 29 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=4.245 $Y=1.655
+ $X2=4.245 $Y2=1.49
r77 10 11 116.613 $w=1.8e-07 $l=3e-07 $layer=POLY_cond $X=4.245 $Y=1.655
+ $X2=4.245 $Y2=1.955
r78 6 25 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.79 $Y=1.325
+ $X2=3.79 $Y2=1.49
r79 6 8 325.606 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.79 $Y=1.325
+ $X2=3.79 $Y2=0.69
r80 3 5 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=3.755 $Y=2.045
+ $X2=3.755 $Y2=2.54
r81 2 3 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=3.755 $Y=1.955 $X2=3.755
+ $Y2=2.045
r82 1 23 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=3.755 $Y=1.655
+ $X2=3.755 $Y2=1.49
r83 1 2 116.613 $w=1.8e-07 $l=3e-07 $layer=POLY_cond $X=3.755 $Y=1.655 $X2=3.755
+ $Y2=1.955
.ends

.subckt PM_SKY130_FD_SC_HS__AND3_4%A 3 5 7 8 10 13 15 22
c55 22 0 1.40226e-19 $X=5.205 $Y=1.747
r56 22 23 0.424296 $w=5.68e-07 $l=5e-09 $layer=POLY_cond $X=5.205 $Y=1.747
+ $X2=5.21 $Y2=1.747
r57 20 22 7.21303 $w=5.68e-07 $l=8.5e-08 $layer=POLY_cond $X=5.12 $Y=1.747
+ $X2=5.205 $Y2=1.747
r58 18 20 30.9736 $w=5.68e-07 $l=3.65e-07 $layer=POLY_cond $X=4.755 $Y=1.747
+ $X2=5.12 $Y2=1.747
r59 17 18 5.51585 $w=5.68e-07 $l=6.5e-08 $layer=POLY_cond $X=4.69 $Y=1.747
+ $X2=4.755 $Y2=1.747
r60 15 20 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.12
+ $Y=1.615 $X2=5.12 $Y2=1.615
r61 11 23 34.6593 $w=1.5e-07 $l=2.97e-07 $layer=POLY_cond $X=5.21 $Y=1.45
+ $X2=5.21 $Y2=1.747
r62 11 13 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=5.21 $Y=1.45
+ $X2=5.21 $Y2=0.69
r63 8 22 34.6593 $w=1.5e-07 $l=2.98e-07 $layer=POLY_cond $X=5.205 $Y=2.045
+ $X2=5.205 $Y2=1.747
r64 8 10 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=5.205 $Y=2.045
+ $X2=5.205 $Y2=2.54
r65 5 18 34.6593 $w=1.5e-07 $l=2.98e-07 $layer=POLY_cond $X=4.755 $Y=2.045
+ $X2=4.755 $Y2=1.747
r66 5 7 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=4.755 $Y=2.045
+ $X2=4.755 $Y2=2.54
r67 1 17 34.6593 $w=1.5e-07 $l=2.97e-07 $layer=POLY_cond $X=4.69 $Y=1.45
+ $X2=4.69 $Y2=1.747
r68 1 3 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=4.69 $Y=1.45 $X2=4.69
+ $Y2=0.69
.ends

.subckt PM_SKY130_FD_SC_HS__AND3_4%VPWR 1 2 3 4 5 6 19 21 27 31 33 37 41 43 45
+ 47 49 54 59 64 73 76 79 82 86
r82 85 86 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r83 82 83 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r84 79 80 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r85 76 77 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r86 73 74 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r87 70 71 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r88 68 86 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=5.52 $Y2=3.33
r89 68 83 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=4.56 $Y2=3.33
r90 67 68 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r91 65 82 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.645 $Y=3.33
+ $X2=4.48 $Y2=3.33
r92 65 67 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=4.645 $Y=3.33
+ $X2=5.04 $Y2=3.33
r93 64 85 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=5.315 $Y=3.33
+ $X2=5.537 $Y2=3.33
r94 64 67 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=5.315 $Y=3.33
+ $X2=5.04 $Y2=3.33
r95 63 83 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=4.56 $Y2=3.33
r96 63 80 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=3.12 $Y2=3.33
r97 62 63 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r98 60 79 12.3201 $w=1.7e-07 $l=2.9e-07 $layer=LI1_cond $X=3.645 $Y=3.33
+ $X2=3.355 $Y2=3.33
r99 60 62 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=3.645 $Y=3.33
+ $X2=4.08 $Y2=3.33
r100 59 82 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.315 $Y=3.33
+ $X2=4.48 $Y2=3.33
r101 59 62 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=4.315 $Y=3.33
+ $X2=4.08 $Y2=3.33
r102 58 77 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r103 58 74 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r104 57 58 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r105 55 73 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.395 $Y=3.33
+ $X2=1.23 $Y2=3.33
r106 55 57 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=1.395 $Y=3.33
+ $X2=1.68 $Y2=3.33
r107 54 76 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.065 $Y=3.33
+ $X2=2.23 $Y2=3.33
r108 54 57 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=2.065 $Y=3.33
+ $X2=1.68 $Y2=3.33
r109 53 74 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r110 53 71 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r111 52 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r112 50 70 4.00981 $w=1.7e-07 $l=1.83e-07 $layer=LI1_cond $X=0.365 $Y=3.33
+ $X2=0.182 $Y2=3.33
r113 50 52 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=0.365 $Y=3.33
+ $X2=0.72 $Y2=3.33
r114 49 73 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.065 $Y=3.33
+ $X2=1.23 $Y2=3.33
r115 49 52 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.065 $Y=3.33
+ $X2=0.72 $Y2=3.33
r116 47 80 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.88 $Y=3.33
+ $X2=3.12 $Y2=3.33
r117 47 77 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=2.88 $Y=3.33
+ $X2=2.16 $Y2=3.33
r118 43 85 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=5.48 $Y=3.245
+ $X2=5.537 $Y2=3.33
r119 43 45 27.5888 $w=3.28e-07 $l=7.9e-07 $layer=LI1_cond $X=5.48 $Y=3.245
+ $X2=5.48 $Y2=2.455
r120 39 82 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.48 $Y=3.245
+ $X2=4.48 $Y2=3.33
r121 39 41 27.5888 $w=3.28e-07 $l=7.9e-07 $layer=LI1_cond $X=4.48 $Y=3.245
+ $X2=4.48 $Y2=2.455
r122 35 79 2.44113 $w=5.8e-07 $l=8.5e-08 $layer=LI1_cond $X=3.355 $Y=3.245
+ $X2=3.355 $Y2=3.33
r123 35 37 16.2914 $w=5.78e-07 $l=7.9e-07 $layer=LI1_cond $X=3.355 $Y=3.245
+ $X2=3.355 $Y2=2.455
r124 34 76 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.395 $Y=3.33
+ $X2=2.23 $Y2=3.33
r125 33 79 12.3201 $w=1.7e-07 $l=2.9e-07 $layer=LI1_cond $X=3.065 $Y=3.33
+ $X2=3.355 $Y2=3.33
r126 33 34 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.065 $Y=3.33
+ $X2=2.395 $Y2=3.33
r127 29 76 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.23 $Y=3.245
+ $X2=2.23 $Y2=3.33
r128 29 31 27.5888 $w=3.28e-07 $l=7.9e-07 $layer=LI1_cond $X=2.23 $Y=3.245
+ $X2=2.23 $Y2=2.455
r129 25 73 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.23 $Y=3.245
+ $X2=1.23 $Y2=3.33
r130 25 27 32.8272 $w=3.28e-07 $l=9.4e-07 $layer=LI1_cond $X=1.23 $Y=3.245
+ $X2=1.23 $Y2=2.305
r131 21 24 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=0.24 $Y=1.985
+ $X2=0.24 $Y2=2.815
r132 19 70 3.13335 $w=2.5e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.24 $Y=3.245
+ $X2=0.182 $Y2=3.33
r133 19 24 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=0.24 $Y=3.245
+ $X2=0.24 $Y2=2.815
r134 6 45 300 $w=1.7e-07 $l=4.2335e-07 $layer=licon1_PDIFF $count=2 $X=5.28
+ $Y=2.12 $X2=5.48 $Y2=2.455
r135 5 41 300 $w=1.7e-07 $l=4.07216e-07 $layer=licon1_PDIFF $count=2 $X=4.32
+ $Y=2.12 $X2=4.48 $Y2=2.455
r136 4 37 150 $w=1.7e-07 $l=6.40976e-07 $layer=licon1_PDIFF $count=4 $X=3.03
+ $Y=2.12 $X2=3.525 $Y2=2.455
r137 3 31 300 $w=1.7e-07 $l=7.07972e-07 $layer=licon1_PDIFF $count=2 $X=2.03
+ $Y=1.84 $X2=2.23 $Y2=2.455
r138 2 27 300 $w=1.7e-07 $l=5.5608e-07 $layer=licon1_PDIFF $count=2 $X=1.03
+ $Y=1.84 $X2=1.23 $Y2=2.305
r139 1 24 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.815
r140 1 21 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HS__AND3_4%X 1 2 3 4 13 15 19 23 27 28 29 30 31 32 33 50
+ 60
c69 15 0 4.56703e-20 $X=1.565 $Y=1.885
r70 57 60 0.516019 $w=3.33e-07 $l=1.5e-08 $layer=LI1_cond $X=0.727 $Y=1.97
+ $X2=0.727 $Y2=1.985
r71 43 50 1.22229 $w=3.28e-07 $l=3.5e-08 $layer=LI1_cond $X=0.725 $Y=0.96
+ $X2=0.725 $Y2=0.925
r72 32 33 12.7285 $w=3.33e-07 $l=3.7e-07 $layer=LI1_cond $X=0.727 $Y=2.405
+ $X2=0.727 $Y2=2.775
r73 31 52 3.10218 $w=3.05e-07 $l=9.88686e-08 $layer=LI1_cond $X=0.727 $Y=1.885
+ $X2=0.697 $Y2=1.8
r74 31 57 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.727 $Y=1.885
+ $X2=0.727 $Y2=1.97
r75 31 32 12.3845 $w=3.33e-07 $l=3.6e-07 $layer=LI1_cond $X=0.727 $Y=2.045
+ $X2=0.727 $Y2=2.405
r76 31 60 2.06408 $w=3.33e-07 $l=6e-08 $layer=LI1_cond $X=0.727 $Y=2.045
+ $X2=0.727 $Y2=1.985
r77 30 52 5.65745 $w=2.73e-07 $l=1.35e-07 $layer=LI1_cond $X=0.697 $Y=1.665
+ $X2=0.697 $Y2=1.8
r78 29 30 15.5056 $w=2.73e-07 $l=3.7e-07 $layer=LI1_cond $X=0.697 $Y=1.295
+ $X2=0.697 $Y2=1.665
r79 29 51 6.91466 $w=2.73e-07 $l=1.65e-07 $layer=LI1_cond $X=0.697 $Y=1.295
+ $X2=0.697 $Y2=1.13
r80 28 43 3.12539 $w=3.02e-07 $l=8.5e-08 $layer=LI1_cond $X=0.725 $Y=1.045
+ $X2=0.725 $Y2=0.96
r81 28 51 3.12539 $w=3.02e-07 $l=9.80051e-08 $layer=LI1_cond $X=0.725 $Y=1.045
+ $X2=0.697 $Y2=1.13
r82 28 50 0.873063 $w=3.28e-07 $l=2.5e-08 $layer=LI1_cond $X=0.725 $Y=0.9
+ $X2=0.725 $Y2=0.925
r83 27 28 13.4452 $w=3.28e-07 $l=3.85e-07 $layer=LI1_cond $X=0.725 $Y=0.515
+ $X2=0.725 $Y2=0.9
r84 23 25 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=1.73 $Y=1.985
+ $X2=1.73 $Y2=2.815
r85 21 23 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=1.73 $Y=1.97
+ $X2=1.73 $Y2=1.985
r86 17 19 20.5135 $w=2.48e-07 $l=4.45e-07 $layer=LI1_cond $X=1.615 $Y=0.96
+ $X2=1.615 $Y2=0.515
r87 16 31 3.51065 $w=1.7e-07 $l=1.68e-07 $layer=LI1_cond $X=0.895 $Y=1.885
+ $X2=0.727 $Y2=1.885
r88 15 21 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.565 $Y=1.885
+ $X2=1.73 $Y2=1.97
r89 15 16 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.565 $Y=1.885
+ $X2=0.895 $Y2=1.885
r90 14 28 3.47949 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.89 $Y=1.045
+ $X2=0.725 $Y2=1.045
r91 13 17 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.49 $Y=1.045
+ $X2=1.615 $Y2=0.96
r92 13 14 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=1.49 $Y=1.045 $X2=0.89
+ $Y2=1.045
r93 4 25 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=1.58
+ $Y=1.84 $X2=1.73 $Y2=2.815
r94 4 23 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=1.58
+ $Y=1.84 $X2=1.73 $Y2=1.985
r95 3 33 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=0.58
+ $Y=1.84 $X2=0.73 $Y2=2.815
r96 3 60 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=0.58
+ $Y=1.84 $X2=0.73 $Y2=1.985
r97 2 19 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.515
+ $Y=0.37 $X2=1.655 $Y2=0.515
r98 1 27 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=0.585
+ $Y=0.37 $X2=0.725 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__AND3_4%VGND 1 2 3 4 13 15 19 23 27 29 31 36 41 48 49
+ 55 58 61
r72 61 62 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r73 58 59 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r74 55 56 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r75 52 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r76 49 62 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=5.52 $Y=0 $X2=3.12
+ $Y2=0
r77 48 49 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r78 46 61 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.18 $Y=0 $X2=3.015
+ $Y2=0
r79 46 48 152.663 $w=1.68e-07 $l=2.34e-06 $layer=LI1_cond $X=3.18 $Y=0 $X2=5.52
+ $Y2=0
r80 45 59 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=2.16
+ $Y2=0
r81 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r82 42 58 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.25 $Y=0 $X2=2.085
+ $Y2=0
r83 42 44 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=2.25 $Y=0 $X2=2.64
+ $Y2=0
r84 41 61 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.85 $Y=0 $X2=3.015
+ $Y2=0
r85 41 44 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=2.85 $Y=0 $X2=2.64
+ $Y2=0
r86 40 59 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r87 40 56 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r88 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r89 37 55 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.32 $Y=0 $X2=1.195
+ $Y2=0
r90 37 39 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=1.32 $Y=0 $X2=1.68
+ $Y2=0
r91 36 58 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.92 $Y=0 $X2=2.085
+ $Y2=0
r92 36 39 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=1.92 $Y=0 $X2=1.68
+ $Y2=0
r93 35 56 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r94 35 53 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r95 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r96 32 52 3.99177 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.38 $Y=0 $X2=0.19
+ $Y2=0
r97 32 34 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=0.38 $Y=0 $X2=0.72
+ $Y2=0
r98 31 55 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.07 $Y=0 $X2=1.195
+ $Y2=0
r99 31 34 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=1.07 $Y=0 $X2=0.72
+ $Y2=0
r100 29 62 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.88 $Y=0
+ $X2=3.12 $Y2=0
r101 29 45 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.88 $Y=0
+ $X2=2.64 $Y2=0
r102 25 61 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.015 $Y=0.085
+ $X2=3.015 $Y2=0
r103 25 27 19.7312 $w=3.28e-07 $l=5.65e-07 $layer=LI1_cond $X=3.015 $Y=0.085
+ $X2=3.015 $Y2=0.65
r104 21 58 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.085 $Y=0.085
+ $X2=2.085 $Y2=0
r105 21 23 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=2.085 $Y=0.085
+ $X2=2.085 $Y2=0.515
r106 17 55 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.195 $Y=0.085
+ $X2=1.195 $Y2=0
r107 17 19 24.8928 $w=2.48e-07 $l=5.4e-07 $layer=LI1_cond $X=1.195 $Y=0.085
+ $X2=1.195 $Y2=0.625
r108 13 52 3.1514 $w=2.5e-07 $l=1.12916e-07 $layer=LI1_cond $X=0.255 $Y=0.085
+ $X2=0.19 $Y2=0
r109 13 15 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=0.255 $Y=0.085
+ $X2=0.255 $Y2=0.515
r110 4 27 182 $w=1.7e-07 $l=3.42929e-07 $layer=licon1_NDIFF $count=1 $X=2.875
+ $Y=0.37 $X2=3.015 $Y2=0.65
r111 3 23 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.945
+ $Y=0.37 $X2=2.085 $Y2=0.515
r112 2 19 182 $w=1.7e-07 $l=3.17372e-07 $layer=licon1_NDIFF $count=1 $X=1.015
+ $Y=0.37 $X2=1.155 $Y2=0.625
r113 1 15 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.15
+ $Y=0.37 $X2=0.295 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__AND3_4%A_489_74# 1 2 9 11 12 15
c31 9 0 3.04787e-19 $X=2.585 $Y=0.515
r32 13 15 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=4.005 $Y=0.985
+ $X2=4.005 $Y2=0.81
r33 11 13 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.92 $Y=1.07
+ $X2=4.005 $Y2=0.985
r34 11 12 81.5508 $w=1.68e-07 $l=1.25e-06 $layer=LI1_cond $X=3.92 $Y=1.07
+ $X2=2.67 $Y2=1.07
r35 7 12 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=2.545 $Y=0.985
+ $X2=2.67 $Y2=1.07
r36 7 9 21.6659 $w=2.48e-07 $l=4.7e-07 $layer=LI1_cond $X=2.545 $Y=0.985
+ $X2=2.545 $Y2=0.515
r37 2 15 182 $w=1.7e-07 $l=5.05173e-07 $layer=licon1_NDIFF $count=1 $X=3.865
+ $Y=0.37 $X2=4.005 $Y2=0.81
r38 1 9 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.445
+ $Y=0.37 $X2=2.585 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__AND3_4%A_686_74# 1 2 3 12 14 15 18 20 24 26
r45 22 24 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=5.475 $Y=0.425
+ $X2=5.475 $Y2=0.515
r46 21 26 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.64 $Y=0.34
+ $X2=4.475 $Y2=0.34
r47 20 22 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=5.31 $Y=0.34
+ $X2=5.475 $Y2=0.425
r48 20 21 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.31 $Y=0.34
+ $X2=4.64 $Y2=0.34
r49 16 26 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.475 $Y=0.425
+ $X2=4.475 $Y2=0.34
r50 16 18 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=4.475 $Y=0.425
+ $X2=4.475 $Y2=0.515
r51 14 26 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.31 $Y=0.34
+ $X2=4.475 $Y2=0.34
r52 14 15 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=4.31 $Y=0.34
+ $X2=3.74 $Y2=0.34
r53 10 15 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.575 $Y=0.425
+ $X2=3.74 $Y2=0.34
r54 10 12 7.85757 $w=3.28e-07 $l=2.25e-07 $layer=LI1_cond $X=3.575 $Y=0.425
+ $X2=3.575 $Y2=0.65
r55 3 24 91 $w=1.7e-07 $l=2.5229e-07 $layer=licon1_NDIFF $count=2 $X=5.285
+ $Y=0.37 $X2=5.475 $Y2=0.515
r56 2 18 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=4.335
+ $Y=0.37 $X2=4.475 $Y2=0.515
r57 1 12 182 $w=1.7e-07 $l=3.44964e-07 $layer=licon1_NDIFF $count=1 $X=3.43
+ $Y=0.37 $X2=3.575 $Y2=0.65
.ends

