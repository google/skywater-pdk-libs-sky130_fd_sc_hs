* File: sky130_fd_sc_hs__sedfxtp_1.spice
* Created: Tue Sep  1 20:24:33 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hs__sedfxtp_1.pex.spice"
.subckt sky130_fd_sc_hs__sedfxtp_1  VNB VPB D DE SCD SCE CLK VPWR Q VGND
* 
* VGND	VGND
* Q	Q
* VPWR	VPWR
* CLK	CLK
* SCE	SCE
* SCD	SCD
* DE	DE
* D	D
* VPB	VPB
* VNB	VNB
MM1017 A_143_74# N_D_M1017_g N_A_27_74#_M1017_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.0504 AS=0.1806 PD=0.66 PS=1.7 NRD=18.564 NRS=21.42 M=1 R=2.8 SA=75000.4
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1004 N_VGND_M1004_d N_DE_M1004_g A_143_74# VNB NLOWVT L=0.15 W=0.42 AD=0.1197
+ AS=0.0504 PD=1.41 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75000.7 SB=75000.2
+ A=0.063 P=1.14 MULT=1
MM1010 N_VGND_M1010_d N_DE_M1010_g N_A_159_404#_M1010_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.0588 AS=0.1197 PD=0.7 PS=1.41 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2 SB=75001.5
+ A=0.063 P=1.14 MULT=1
MM1012 A_505_111# N_A_159_404#_M1012_g N_VGND_M1010_d VNB NLOWVT L=0.15 W=0.42
+ AD=0.0504 AS=0.0588 PD=0.66 PS=0.7 NRD=18.564 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1038 N_A_27_74#_M1038_d N_A_547_301#_M1038_g A_505_111# VNB NLOWVT L=0.15
+ W=0.42 AD=0.0588 AS=0.0504 PD=0.7 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75001
+ SB=75000.7 A=0.063 P=1.14 MULT=1
MM1025 N_A_669_111#_M1025_d N_A_639_85#_M1025_g N_A_27_74#_M1038_d VNB NLOWVT
+ L=0.15 W=0.42 AD=0.1491 AS=0.0588 PD=1.55 PS=0.7 NRD=19.992 NRS=0 M=1 R=2.8
+ SA=75001.5 SB=75000.3 A=0.063 P=1.14 MULT=1
MM1041 N_VGND_M1041_d N_SCE_M1041_g N_A_639_85#_M1041_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.0588 AS=0.1176 PD=0.7 PS=1.4 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2 SB=75001
+ A=0.063 P=1.14 MULT=1
MM1031 A_1026_125# N_SCD_M1031_g N_VGND_M1041_d VNB NLOWVT L=0.15 W=0.42
+ AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1028 N_A_669_111#_M1028_d N_SCE_M1028_g A_1026_125# VNB NLOWVT L=0.15 W=0.42
+ AD=0.1176 AS=0.0441 PD=1.4 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75001
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1018 N_A_1295_74#_M1018_d N_CLK_M1018_g N_VGND_M1018_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.2072 AS=0.2109 PD=2.04 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1007 N_A_1492_74#_M1007_d N_A_1295_74#_M1007_g N_VGND_M1007_s VNB NLOWVT
+ L=0.15 W=0.74 AD=0.2072 AS=0.2109 PD=2.04 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1026 N_A_1688_97#_M1026_d N_A_1295_74#_M1026_g N_A_669_111#_M1026_s VNB NLOWVT
+ L=0.15 W=0.42 AD=0.1113 AS=0.1176 PD=0.95 PS=1.4 NRD=71.424 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75002.2 A=0.063 P=1.14 MULT=1
MM1032 A_1824_97# N_A_1492_74#_M1032_g N_A_1688_97#_M1026_d VNB NLOWVT L=0.15
+ W=0.42 AD=0.0903 AS=0.1113 PD=0.85 PS=0.95 NRD=45.708 NRS=0 M=1 R=2.8
+ SA=75000.9 SB=75001.5 A=0.063 P=1.14 MULT=1
MM1029 N_VGND_M1029_d N_A_1910_71#_M1029_g A_1824_97# VNB NLOWVT L=0.15 W=0.42
+ AD=0.135232 AS=0.0903 PD=0.986604 PS=0.85 NRD=22.848 NRS=45.708 M=1 R=2.8
+ SA=75001.5 SB=75001 A=0.063 P=1.14 MULT=1
MM1033 N_A_1910_71#_M1033_d N_A_1688_97#_M1033_g N_VGND_M1029_d VNB NLOWVT
+ L=0.15 W=0.64 AD=0.1824 AS=0.206068 PD=1.85 PS=1.5034 NRD=0 NRS=46.872 M=1
+ R=4.26667 SA=75001.6 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1022 A_2313_74# N_A_1910_71#_M1022_g N_VGND_M1022_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.0672 AS=0.1824 PD=0.85 PS=1.85 NRD=9.372 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75001.9 A=0.096 P=1.58 MULT=1
MM1024 N_A_2385_74#_M1024_d N_A_1492_74#_M1024_g A_2313_74# VNB NLOWVT L=0.15
+ W=0.64 AD=0.129147 AS=0.0672 PD=1.20755 PS=0.85 NRD=0 NRS=9.372 M=1 R=4.26667
+ SA=75000.6 SB=75001.5 A=0.096 P=1.58 MULT=1
MM1034 A_2487_74# N_A_1295_74#_M1034_g N_A_2385_74#_M1024_d VNB NLOWVT L=0.15
+ W=0.42 AD=0.0504 AS=0.0847528 PD=0.66 PS=0.792453 NRD=18.564 NRS=23.568 M=1
+ R=2.8 SA=75001.1 SB=75001.7 A=0.063 P=1.14 MULT=1
MM1035 N_VGND_M1035_d N_A_547_301#_M1035_g A_2487_74# VNB NLOWVT L=0.15 W=0.42
+ AD=0.20475 AS=0.0504 PD=1.395 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75001.5
+ SB=75001.3 A=0.063 P=1.14 MULT=1
MM1019 N_A_547_301#_M1019_d N_A_2385_74#_M1019_g N_VGND_M1035_d VNB NLOWVT
+ L=0.15 W=0.42 AD=0.1197 AS=0.20475 PD=1.41 PS=1.395 NRD=0 NRS=19.992 M=1 R=2.8
+ SA=75002.6 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1006 N_VGND_M1006_d N_A_2385_74#_M1006_g N_Q_M1006_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.2109 PD=2.05 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1037 A_114_464# N_D_M1037_g N_A_27_74#_M1037_s VPB PSHORT L=0.15 W=0.64
+ AD=0.0768 AS=0.1824 PD=0.88 PS=1.85 NRD=19.9955 NRS=3.0732 M=1 R=4.26667
+ SA=75000.2 SB=75000.6 A=0.096 P=1.58 MULT=1
MM1023 N_VPWR_M1023_d N_A_159_404#_M1023_g A_114_464# VPB PSHORT L=0.15 W=0.64
+ AD=0.1888 AS=0.0768 PD=1.87 PS=0.88 NRD=3.0732 NRS=19.9955 M=1 R=4.26667
+ SA=75000.6 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1036 N_VPWR_M1036_d N_DE_M1036_g N_A_159_404#_M1036_s VPB PSHORT L=0.15 W=0.64
+ AD=0.1696 AS=0.1888 PD=1.17 PS=1.87 NRD=73.8553 NRS=3.0732 M=1 R=4.26667
+ SA=75000.2 SB=75001.7 A=0.096 P=1.58 MULT=1
MM1013 A_554_463# N_DE_M1013_g N_VPWR_M1036_d VPB PSHORT L=0.15 W=0.64 AD=0.0768
+ AS=0.1696 PD=0.88 PS=1.17 NRD=19.9955 NRS=3.0732 M=1 R=4.26667 SA=75000.9
+ SB=75001 A=0.096 P=1.58 MULT=1
MM1000 N_A_27_74#_M1000_d N_A_547_301#_M1000_g A_554_463# VPB PSHORT L=0.15
+ W=0.64 AD=0.096 AS=0.0768 PD=0.94 PS=0.88 NRD=3.0732 NRS=19.9955 M=1 R=4.26667
+ SA=75001.3 SB=75000.6 A=0.096 P=1.58 MULT=1
MM1008 N_A_669_111#_M1008_d N_SCE_M1008_g N_A_27_74#_M1000_d VPB PSHORT L=0.15
+ W=0.64 AD=0.176 AS=0.096 PD=1.83 PS=0.94 NRD=3.0732 NRS=3.0732 M=1 R=4.26667
+ SA=75001.7 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1027 N_VPWR_M1027_d N_SCE_M1027_g N_A_639_85#_M1027_s VPB PSHORT L=0.15 W=0.64
+ AD=0.1696 AS=0.1792 PD=1.17 PS=1.84 NRD=73.8553 NRS=3.0732 M=1 R=4.26667
+ SA=75000.2 SB=75001.3 A=0.096 P=1.58 MULT=1
MM1016 A_1053_455# N_SCD_M1016_g N_VPWR_M1027_d VPB PSHORT L=0.15 W=0.64
+ AD=0.0768 AS=0.1696 PD=0.88 PS=1.17 NRD=19.9955 NRS=3.0732 M=1 R=4.26667
+ SA=75000.9 SB=75000.6 A=0.096 P=1.58 MULT=1
MM1002 N_A_669_111#_M1002_d N_A_639_85#_M1002_g A_1053_455# VPB PSHORT L=0.15
+ W=0.64 AD=0.176 AS=0.0768 PD=1.83 PS=0.88 NRD=3.0732 NRS=19.9955 M=1 R=4.26667
+ SA=75001.3 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1020 N_A_1295_74#_M1020_d N_CLK_M1020_g N_VPWR_M1020_s VPB PSHORT L=0.15
+ W=1.12 AD=0.308 AS=0.308 PD=2.79 PS=2.79 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75000.2 A=0.168 P=2.54 MULT=1
MM1030 N_A_1492_74#_M1030_d N_A_1295_74#_M1030_g N_VPWR_M1030_s VPB PSHORT
+ L=0.15 W=1.12 AD=0.308 AS=0.308 PD=2.79 PS=2.79 NRD=1.7533 NRS=1.7533 M=1
+ R=7.46667 SA=75000.2 SB=75000.2 A=0.168 P=2.54 MULT=1
MM1015 N_A_1688_97#_M1015_d N_A_1492_74#_M1015_g N_A_669_111#_M1015_s VPB PSHORT
+ L=0.15 W=0.42 AD=0.0735 AS=0.1176 PD=0.77 PS=1.4 NRD=28.1316 NRS=4.6886 M=1
+ R=2.8 SA=75000.2 SB=75001.5 A=0.063 P=1.14 MULT=1
MM1014 A_1890_508# N_A_1295_74#_M1014_g N_A_1688_97#_M1015_d VPB PSHORT L=0.15
+ W=0.42 AD=0.0588 AS=0.0735 PD=0.7 PS=0.77 NRD=39.8531 NRS=4.6886 M=1 R=2.8
+ SA=75000.7 SB=75001 A=0.063 P=1.14 MULT=1
MM1003 N_VPWR_M1003_d N_A_1910_71#_M1003_g A_1890_508# VPB PSHORT L=0.15 W=0.42
+ AD=0.0964833 AS=0.0588 PD=0.893333 PS=0.7 NRD=4.6886 NRS=39.8531 M=1 R=2.8
+ SA=75001.1 SB=75000.6 A=0.063 P=1.14 MULT=1
MM1039 N_A_1910_71#_M1039_d N_A_1688_97#_M1039_g N_VPWR_M1003_d VPB PSHORT
+ L=0.15 W=0.84 AD=0.231 AS=0.192967 PD=2.23 PS=1.78667 NRD=2.3443 NRS=19.9167
+ M=1 R=5.6 SA=75000.7 SB=75000.2 A=0.126 P=1.98 MULT=1
MM1009 A_2274_392# N_A_1910_71#_M1009_g N_VPWR_M1009_s VPB PSHORT L=0.15 W=1
+ AD=0.3925 AS=0.275 PD=1.785 PS=2.55 NRD=66.4678 NRS=1.9503 M=1 R=6.66667
+ SA=75000.2 SB=75001.8 A=0.15 P=2.3 MULT=1
MM1001 N_A_2385_74#_M1001_d N_A_1295_74#_M1001_g A_2274_392# VPB PSHORT L=0.15
+ W=1 AD=0.234366 AS=0.3925 PD=1.9507 PS=1.785 NRD=1.9503 NRS=66.4678 M=1
+ R=6.66667 SA=75001.1 SB=75000.9 A=0.15 P=2.3 MULT=1
MM1040 A_2568_508# N_A_1492_74#_M1040_g N_A_2385_74#_M1001_d VPB PSHORT L=0.15
+ W=0.42 AD=0.0567 AS=0.0984338 PD=0.69 PS=0.819296 NRD=37.5088 NRS=45.7237 M=1
+ R=2.8 SA=75001.7 SB=75001.3 A=0.063 P=1.14 MULT=1
MM1021 N_VPWR_M1021_d N_A_547_301#_M1021_g A_2568_508# VPB PSHORT L=0.15 W=0.42
+ AD=0.116292 AS=0.0567 PD=0.950943 PS=0.69 NRD=72.693 NRS=37.5088 M=1 R=2.8
+ SA=75002.1 SB=75000.9 A=0.063 P=1.14 MULT=1
MM1005 N_A_547_301#_M1005_d N_A_2385_74#_M1005_g N_VPWR_M1021_d VPB PSHORT
+ L=0.15 W=0.64 AD=0.176 AS=0.177208 PD=1.83 PS=1.44906 NRD=3.0732 NRS=38.4741
+ M=1 R=4.26667 SA=75001.9 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1011 N_VPWR_M1011_d N_A_2385_74#_M1011_g N_Q_M1011_s VPB PSHORT L=0.15 W=1.12
+ AD=0.3192 AS=0.308 PD=2.81 PS=2.79 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75000.2 A=0.168 P=2.54 MULT=1
DX42_noxref VNB VPB NWDIODE A=29.34 P=35.32
c_169 VNB 0 2.70131e-19 $X=0 $Y=0
c_328 VPB 0 8.71884e-20 $X=0 $Y=3.085
*
.include "sky130_fd_sc_hs__sedfxtp_1.pxi.spice"
*
.ends
*
*
