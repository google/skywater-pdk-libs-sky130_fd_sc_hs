# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_hs__nor3_1
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_hs__nor3_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  1.920000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105000 1.180000 0.360000 1.780000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.870000 1.300000 1.315000 1.780000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.485000 1.300000 1.815000 1.780000 ;
    END
  END C
  PIN Y
    ANTENNADIFFAREA  0.737300 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.530000 0.880000 1.805000 1.130000 ;
        RECT 0.530000 1.130000 0.700000 1.950000 ;
        RECT 0.530000 1.950000 1.815000 2.120000 ;
        RECT 0.605000 2.120000 1.815000 2.980000 ;
        RECT 0.615000 0.365000 0.805000 0.880000 ;
        RECT 1.475000 0.350000 1.805000 0.880000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 1.920000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 1.920000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 1.920000 0.085000 ;
      RECT 0.000000  3.245000 1.920000 3.415000 ;
      RECT 0.105000  1.950000 0.355000 2.325000 ;
      RECT 0.105000  2.325000 0.435000 3.245000 ;
      RECT 0.115000  0.085000 0.445000 0.710000 ;
      RECT 0.115000  0.710000 0.360000 1.010000 ;
      RECT 0.975000  0.085000 1.305000 0.710000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
  END
END sky130_fd_sc_hs__nor3_1
END LIBRARY
