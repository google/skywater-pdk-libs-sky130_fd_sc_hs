* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hs__a31o_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
X0 VPWR a_83_274# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X1 VGND a_83_274# X VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X2 VPWR A1 a_529_392# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=150000u
X3 X a_83_274# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X4 VPWR A3 a_529_392# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=150000u
X5 a_83_274# B1 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X6 a_529_392# B1 a_83_274# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=150000u
X7 a_83_274# A1 a_775_74# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X8 a_83_274# B1 a_529_392# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=150000u
X9 a_529_392# A2 VPWR VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=150000u
X10 a_529_392# A1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=150000u
X11 VGND a_83_274# X VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X12 VPWR a_83_274# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X13 a_1000_74# A2 a_775_74# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X14 X a_83_274# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X15 X a_83_274# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X16 VPWR A2 a_529_392# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=150000u
X17 a_1000_74# A3 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X18 X a_83_274# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X19 a_775_74# A2 a_1000_74# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X20 a_529_392# A3 VPWR VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=150000u
X21 VGND B1 a_83_274# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X22 a_775_74# A1 a_83_274# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X23 VGND A3 a_1000_74# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
.ends
