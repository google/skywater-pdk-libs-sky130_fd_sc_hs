* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hs__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
X0 VPWR A2 a_80_392# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=150000u
X1 a_431_392# D1 a_85_136# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=150000u
X2 VPWR a_85_136# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X3 a_80_392# A1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=150000u
X4 VGND B1 a_85_136# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X5 a_80_392# B1 a_353_392# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=150000u
X6 a_85_136# A1 a_168_136# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X7 VGND D1 a_85_136# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X8 a_85_136# C1 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X9 a_353_392# C1 a_431_392# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=150000u
X10 a_168_136# A2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X11 VGND a_85_136# X VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
.ends
