* File: sky130_fd_sc_hs__dfxtp_1.spice
* Created: Thu Aug 27 20:39:57 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hs__dfxtp_1.pex.spice"
.subckt sky130_fd_sc_hs__dfxtp_1  VNB VPB CLK D VPWR Q VGND
* 
* VGND	VGND
* Q	Q
* VPWR	VPWR
* D	D
* CLK	CLK
* VPB	VPB
* VNB	VNB
MM1021 N_VGND_M1021_d N_CLK_M1021_g N_A_27_74#_M1021_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1739 AS=0.2109 PD=1.21 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75000.9 A=0.111 P=1.78 MULT=1
MM1003 N_A_206_368#_M1003_d N_A_27_74#_M1003_g N_VGND_M1021_d VNB NLOWVT L=0.15
+ W=0.74 AD=0.2553 AS=0.1739 PD=2.17 PS=1.21 NRD=9.72 NRS=30.804 M=1 R=4.93333
+ SA=75000.8 SB=75000.3 A=0.111 P=1.78 MULT=1
MM1007 N_A_454_503#_M1007_d N_D_M1007_g N_VGND_M1007_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.155625 AS=0.23015 PD=1.215 PS=2.1 NRD=90.144 NRS=140.844 M=1 R=2.8
+ SA=75000.3 SB=75003 A=0.063 P=1.14 MULT=1
MM1019 N_A_561_463#_M1019_d N_A_27_74#_M1019_g N_A_454_503#_M1007_d VNB NLOWVT
+ L=0.15 W=0.42 AD=0.07875 AS=0.155625 PD=0.865 PS=1.215 NRD=1.428 NRS=90.144
+ M=1 R=2.8 SA=75000.9 SB=75002.4 A=0.063 P=1.14 MULT=1
MM1017 A_731_101# N_A_206_368#_M1017_g N_A_561_463#_M1019_d VNB NLOWVT L=0.15
+ W=0.42 AD=0.0441 AS=0.07875 PD=0.63 PS=0.865 NRD=14.28 NRS=11.424 M=1 R=2.8
+ SA=75001.1 SB=75002.5 A=0.063 P=1.14 MULT=1
MM1013 N_VGND_M1013_d N_A_713_458#_M1013_g A_731_101# VNB NLOWVT L=0.15 W=0.42
+ AD=0.142713 AS=0.0441 PD=1.07814 PS=0.63 NRD=81.36 NRS=14.28 M=1 R=2.8
+ SA=75001.4 SB=75002.2 A=0.063 P=1.14 MULT=1
MM1004 N_A_713_458#_M1004_d N_A_561_463#_M1004_g N_VGND_M1013_d VNB NLOWVT
+ L=0.15 W=0.55 AD=0.109062 AS=0.186887 PD=1.025 PS=1.41186 NRD=17.448
+ NRS=38.172 M=1 R=3.66667 SA=75001.7 SB=75001.2 A=0.0825 P=1.4 MULT=1
MM1006 N_A_1011_424#_M1006_d N_A_206_368#_M1006_g N_A_713_458#_M1004_d VNB
+ NLOWVT L=0.15 W=0.55 AD=0.133928 AS=0.109062 PD=1.17371 PS=1.025 NRD=21.816
+ NRS=0 M=1 R=3.66667 SA=75002.1 SB=75001 A=0.0825 P=1.4 MULT=1
MM1002 A_1168_124# N_A_27_74#_M1002_g N_A_1011_424#_M1006_d VNB NLOWVT L=0.15
+ W=0.42 AD=0.05565 AS=0.102272 PD=0.685 PS=0.896289 NRD=22.14 NRS=30 M=1 R=2.8
+ SA=75002.8 SB=75000.6 A=0.063 P=1.14 MULT=1
MM1020 N_VGND_M1020_d N_A_1210_314#_M1020_g A_1168_124# VNB NLOWVT L=0.15 W=0.42
+ AD=0.1197 AS=0.05565 PD=1.41 PS=0.685 NRD=0 NRS=22.14 M=1 R=2.8 SA=75003.3
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1009 N_VGND_M1009_d N_A_1011_424#_M1009_g N_A_1210_314#_M1009_s VNB NLOWVT
+ L=0.15 W=0.64 AD=0.113994 AS=0.1824 PD=1.00638 PS=1.85 NRD=5.616 NRS=0 M=1
+ R=4.26667 SA=75000.2 SB=75000.7 A=0.096 P=1.58 MULT=1
MM1012 N_Q_M1012_d N_A_1210_314#_M1012_g N_VGND_M1009_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.131806 PD=2.05 PS=1.16362 NRD=0 NRS=5.664 M=1 R=4.93333
+ SA=75000.6 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1016 N_VPWR_M1016_d N_CLK_M1016_g N_A_27_74#_M1016_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.3304 PD=1.42 PS=2.83 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1014 N_A_206_368#_M1014_d N_A_27_74#_M1014_g N_VPWR_M1016_d VPB PSHORT L=0.15
+ W=1.12 AD=0.3304 AS=0.168 PD=2.83 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.7 SB=75000.2 A=0.168 P=2.54 MULT=1
MM1001 N_A_454_503#_M1001_d N_D_M1001_g N_VPWR_M1001_s VPB PSHORT L=0.15 W=0.42
+ AD=0.09835 AS=0.2972 PD=1.005 PS=2.41 NRD=46.886 NRS=306.099 M=1 R=2.8
+ SA=75000.5 SB=75002.2 A=0.063 P=1.14 MULT=1
MM1023 N_A_561_463#_M1023_d N_A_206_368#_M1023_g N_A_454_503#_M1001_d VPB PSHORT
+ L=0.15 W=0.42 AD=0.09835 AS=0.09835 PD=1.005 PS=1.005 NRD=4.6886 NRS=4.6886
+ M=1 R=2.8 SA=75000.6 SB=75001.9 A=0.063 P=1.14 MULT=1
MM1022 A_668_503# N_A_27_74#_M1022_g N_A_561_463#_M1023_d VPB PSHORT L=0.15
+ W=0.42 AD=0.0504 AS=0.09835 PD=0.66 PS=1.005 NRD=30.4759 NRS=46.886 M=1 R=2.8
+ SA=75000.9 SB=75003 A=0.063 P=1.14 MULT=1
MM1015 N_VPWR_M1015_d N_A_713_458#_M1015_g A_668_503# VPB PSHORT L=0.15 W=0.42
+ AD=0.126575 AS=0.0504 PD=1.03 PS=0.66 NRD=115.541 NRS=30.4759 M=1 R=2.8
+ SA=75001.3 SB=75002.6 A=0.063 P=1.14 MULT=1
MM1010 N_A_713_458#_M1010_d N_A_561_463#_M1010_g N_VPWR_M1015_d VPB PSHORT
+ L=0.15 W=0.84 AD=0.2331 AS=0.25315 PD=1.395 PS=2.06 NRD=4.6886 NRS=57.7604 M=1
+ R=5.6 SA=75001 SB=75001.5 A=0.126 P=1.98 MULT=1
MM1018 N_A_1011_424#_M1018_d N_A_27_74#_M1018_g N_A_713_458#_M1010_d VPB PSHORT
+ L=0.15 W=0.84 AD=0.1904 AS=0.2331 PD=1.63333 PS=1.395 NRD=2.3443 NRS=59.7895
+ M=1 R=5.6 SA=75001.8 SB=75000.8 A=0.126 P=1.98 MULT=1
MM1011 A_1118_508# N_A_206_368#_M1011_g N_A_1011_424#_M1018_d VPB PSHORT L=0.15
+ W=0.42 AD=0.09975 AS=0.0952 PD=0.895 PS=0.816667 NRD=85.5965 NRS=46.886 M=1
+ R=2.8 SA=75003 SB=75000.8 A=0.063 P=1.14 MULT=1
MM1005 N_VPWR_M1005_d N_A_1210_314#_M1005_g A_1118_508# VPB PSHORT L=0.15 W=0.42
+ AD=0.1239 AS=0.09975 PD=1.43 PS=0.895 NRD=4.6886 NRS=85.5965 M=1 R=2.8
+ SA=75003.6 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1008 N_VPWR_M1008_d N_A_1011_424#_M1008_g N_A_1210_314#_M1008_s VPB PSHORT
+ L=0.15 W=0.84 AD=0.1596 AS=0.2478 PD=1.26429 PS=2.27 NRD=2.3443 NRS=2.3443 M=1
+ R=5.6 SA=75000.2 SB=75000.7 A=0.126 P=1.98 MULT=1
MM1000 N_Q_M1000_d N_A_1210_314#_M1000_g N_VPWR_M1008_d VPB PSHORT L=0.15 W=1.12
+ AD=0.3304 AS=0.2128 PD=2.83 PS=1.68571 NRD=1.7533 NRS=11.426 M=1 R=7.46667
+ SA=75000.6 SB=75000.2 A=0.168 P=2.54 MULT=1
DX24_noxref VNB VPB NWDIODE A=15.8844 P=20.8
*
.include "sky130_fd_sc_hs__dfxtp_1.pxi.spice"
*
.ends
*
*
