# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_hs__fa_1
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_hs__fa_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  8.640000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.984000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.885000 1.220000 1.215000 1.540000 ;
        RECT 1.045000 0.920000 4.710000 0.935000 ;
        RECT 1.045000 0.935000 5.980000 1.090000 ;
        RECT 1.045000 1.090000 1.215000 1.220000 ;
        RECT 3.300000 1.090000 3.630000 1.455000 ;
        RECT 4.380000 1.090000 5.980000 1.105000 ;
        RECT 4.380000 1.105000 4.710000 1.455000 ;
        RECT 5.810000 1.105000 5.980000 1.320000 ;
        RECT 5.810000 1.320000 6.210000 1.575000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.984000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.800000 1.320000 7.470000 1.780000 ;
    END
  END B
  PIN CIN
    ANTENNAGATEAREA  0.738000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.565000 1.260000 2.115000 1.575000 ;
        RECT 1.565000 1.575000 1.795000 1.780000 ;
        RECT 3.840000 1.260000 4.195000 1.780000 ;
        RECT 4.925000 1.275000 5.640000 1.575000 ;
        RECT 4.925000 1.575000 5.155000 1.780000 ;
      LAYER mcon ;
        RECT 1.595000 1.580000 1.765000 1.750000 ;
        RECT 3.995000 1.580000 4.165000 1.750000 ;
        RECT 4.955000 1.580000 5.125000 1.750000 ;
      LAYER met1 ;
        RECT 1.535000 1.550000 1.825000 1.595000 ;
        RECT 1.535000 1.595000 5.185000 1.735000 ;
        RECT 1.535000 1.735000 1.825000 1.780000 ;
        RECT 3.935000 1.550000 4.225000 1.595000 ;
        RECT 3.935000 1.735000 4.225000 1.780000 ;
        RECT 4.895000 1.550000 5.185000 1.595000 ;
        RECT 4.895000 1.735000 5.185000 1.780000 ;
    END
  END CIN
  PIN COUT
    ANTENNADIFFAREA  0.519000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.210000 0.350000 8.540000 1.130000 ;
        RECT 8.285000 1.130000 8.540000 2.980000 ;
    END
  END COUT
  PIN SUM
    ANTENNADIFFAREA  0.530100 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.350000 0.365000 1.130000 ;
        RECT 0.085000 1.130000 0.255000 1.820000 ;
        RECT 0.085000 1.820000 0.355000 2.980000 ;
    END
  END SUM
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 8.640000 0.085000 ;
        RECT 0.625000  0.085000 0.980000 0.410000 ;
        RECT 3.070000  0.085000 3.400000 0.410000 ;
        RECT 4.080000  0.085000 4.555000 0.710000 ;
        RECT 6.830000  0.085000 7.080000 0.470000 ;
        RECT 7.780000  0.085000 8.030000 0.770000 ;
      LAYER mcon ;
        RECT 0.155000 -0.085000 0.325000 0.085000 ;
        RECT 0.635000 -0.085000 0.805000 0.085000 ;
        RECT 1.115000 -0.085000 1.285000 0.085000 ;
        RECT 1.595000 -0.085000 1.765000 0.085000 ;
        RECT 2.075000 -0.085000 2.245000 0.085000 ;
        RECT 2.555000 -0.085000 2.725000 0.085000 ;
        RECT 3.035000 -0.085000 3.205000 0.085000 ;
        RECT 3.515000 -0.085000 3.685000 0.085000 ;
        RECT 3.995000 -0.085000 4.165000 0.085000 ;
        RECT 4.475000 -0.085000 4.645000 0.085000 ;
        RECT 4.955000 -0.085000 5.125000 0.085000 ;
        RECT 5.435000 -0.085000 5.605000 0.085000 ;
        RECT 5.915000 -0.085000 6.085000 0.085000 ;
        RECT 6.395000 -0.085000 6.565000 0.085000 ;
        RECT 6.875000 -0.085000 7.045000 0.085000 ;
        RECT 7.355000 -0.085000 7.525000 0.085000 ;
        RECT 7.835000 -0.085000 8.005000 0.085000 ;
        RECT 8.315000 -0.085000 8.485000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.245000 8.640000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 3.245000 8.640000 3.415000 ;
        RECT 0.555000 2.050000 0.885000 3.245000 ;
        RECT 3.080000 2.630000 3.410000 3.245000 ;
        RECT 4.105000 2.305000 4.435000 3.245000 ;
        RECT 6.120000 2.500000 6.825000 3.245000 ;
        RECT 7.755000 1.820000 8.085000 3.245000 ;
      LAYER mcon ;
        RECT 0.155000 3.245000 0.325000 3.415000 ;
        RECT 0.635000 3.245000 0.805000 3.415000 ;
        RECT 1.115000 3.245000 1.285000 3.415000 ;
        RECT 1.595000 3.245000 1.765000 3.415000 ;
        RECT 2.075000 3.245000 2.245000 3.415000 ;
        RECT 2.555000 3.245000 2.725000 3.415000 ;
        RECT 3.035000 3.245000 3.205000 3.415000 ;
        RECT 3.515000 3.245000 3.685000 3.415000 ;
        RECT 3.995000 3.245000 4.165000 3.415000 ;
        RECT 4.475000 3.245000 4.645000 3.415000 ;
        RECT 4.955000 3.245000 5.125000 3.415000 ;
        RECT 5.435000 3.245000 5.605000 3.415000 ;
        RECT 5.915000 3.245000 6.085000 3.415000 ;
        RECT 6.395000 3.245000 6.565000 3.415000 ;
        RECT 6.875000 3.245000 7.045000 3.415000 ;
        RECT 7.355000 3.245000 7.525000 3.415000 ;
        RECT 7.835000 3.245000 8.005000 3.415000 ;
        RECT 8.315000 3.245000 8.485000 3.415000 ;
      LAYER met1 ;
        RECT 0.000000 3.085000 8.640000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.425000 1.300000 0.705000 1.630000 ;
      RECT 0.535000 0.580000 2.270000 0.750000 ;
      RECT 0.535000 0.750000 0.705000 1.300000 ;
      RECT 0.535000 1.630000 0.705000 1.710000 ;
      RECT 0.535000 1.710000 1.225000 1.880000 ;
      RECT 1.055000 1.880000 1.225000 1.950000 ;
      RECT 1.055000 1.950000 2.410000 2.120000 ;
      RECT 1.940000 0.355000 2.270000 0.580000 ;
      RECT 2.080000 1.745000 2.410000 1.950000 ;
      RECT 2.080000 2.120000 2.410000 2.755000 ;
      RECT 2.325000 1.260000 2.750000 1.575000 ;
      RECT 2.480000 0.420000 2.890000 0.580000 ;
      RECT 2.480000 0.580000 3.910000 0.750000 ;
      RECT 2.580000 1.575000 2.750000 1.625000 ;
      RECT 2.580000 1.625000 3.200000 1.795000 ;
      RECT 2.610000 1.965000 2.860000 2.290000 ;
      RECT 2.610000 2.290000 3.930000 2.460000 ;
      RECT 2.610000 2.460000 2.860000 2.755000 ;
      RECT 3.030000 1.795000 3.200000 1.950000 ;
      RECT 3.030000 1.950000 5.495000 2.120000 ;
      RECT 3.580000 0.420000 3.910000 0.580000 ;
      RECT 3.600000 2.460000 3.930000 2.755000 ;
      RECT 5.045000 0.435000 5.375000 0.595000 ;
      RECT 5.045000 0.595000 6.320000 0.765000 ;
      RECT 5.070000 2.120000 5.495000 2.755000 ;
      RECT 5.325000 1.745000 6.550000 1.915000 ;
      RECT 5.325000 1.915000 5.495000 1.950000 ;
      RECT 5.555000 0.255000 6.660000 0.425000 ;
      RECT 5.665000 2.085000 7.320000 2.255000 ;
      RECT 5.665000 2.255000 5.950000 2.755000 ;
      RECT 6.150000 0.765000 6.320000 0.980000 ;
      RECT 6.150000 0.980000 8.040000 1.150000 ;
      RECT 6.380000 1.150000 6.550000 1.745000 ;
      RECT 6.490000 0.425000 6.660000 0.640000 ;
      RECT 6.490000 0.640000 7.590000 0.810000 ;
      RECT 6.990000 1.950000 7.320000 2.085000 ;
      RECT 7.000000 2.255000 7.320000 2.830000 ;
      RECT 7.260000 0.480000 7.590000 0.640000 ;
      RECT 7.710000 1.150000 8.040000 1.550000 ;
  END
END sky130_fd_sc_hs__fa_1
