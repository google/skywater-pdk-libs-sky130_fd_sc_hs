* File: sky130_fd_sc_hs__ha_2.pex.spice
* Created: Thu Aug 27 20:47:23 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HS__HA_2%B 5 9 10 12 13 15 16 17 20 27 28 30 31 32 33 34
c86 27 0 7.58277e-20 $X=0.385 $Y=1.465
c87 20 0 1.73571e-19 $X=1.955 $Y=1.615
r88 33 34 26.6182 $w=1.98e-07 $l=4.8e-07 $layer=LI1_cond $X=1.2 $Y=2.42 $X2=1.68
+ $Y2=2.42
r89 32 33 26.6182 $w=1.98e-07 $l=4.8e-07 $layer=LI1_cond $X=0.72 $Y=2.42 $X2=1.2
+ $Y2=2.42
r90 31 45 3.15876 $w=2e-07 $l=8.5e-08 $layer=LI1_cond $X=0.21 $Y=2.42 $X2=0.295
+ $Y2=2.42
r91 31 32 22.7364 $w=1.98e-07 $l=4.1e-07 $layer=LI1_cond $X=0.31 $Y=2.42
+ $X2=0.72 $Y2=2.42
r92 31 45 0.831818 $w=1.98e-07 $l=1.5e-08 $layer=LI1_cond $X=0.31 $Y=2.42
+ $X2=0.295 $Y2=2.42
r93 30 34 6.1 $w=1.98e-07 $l=1.1e-07 $layer=LI1_cond $X=1.79 $Y=2.42 $X2=1.68
+ $Y2=2.42
r94 28 43 45.3857 $w=3.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.395 $Y=1.465
+ $X2=0.395 $Y2=1.63
r95 28 42 46.4315 $w=3.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.395 $Y=1.465
+ $X2=0.395 $Y2=1.3
r96 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.385
+ $Y=1.465 $X2=0.385 $Y2=1.465
r97 24 31 26.9578 $w=3.08e-07 $l=6.9e-07 $layer=LI1_cond $X=0.21 $Y=1.63
+ $X2=0.21 $Y2=2.32
r98 23 27 6.11144 $w=3.28e-07 $l=1.75e-07 $layer=LI1_cond $X=0.21 $Y=1.465
+ $X2=0.385 $Y2=1.465
r99 23 24 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.21 $Y=1.465
+ $X2=0.21 $Y2=1.63
r100 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.955
+ $Y=1.615 $X2=1.955 $Y2=1.615
r101 18 30 7.36389 $w=2e-07 $l=2.09105e-07 $layer=LI1_cond $X=1.955 $Y=2.32
+ $X2=1.79 $Y2=2.42
r102 18 20 24.6204 $w=3.28e-07 $l=7.05e-07 $layer=LI1_cond $X=1.955 $Y=2.32
+ $X2=1.955 $Y2=1.615
r103 16 17 26.3127 $w=1.55e-07 $l=5.5e-08 $layer=POLY_cond $X=0.497 $Y=1.79
+ $X2=0.497 $Y2=1.845
r104 16 43 76.5459 $w=1.55e-07 $l=1.6e-07 $layer=POLY_cond $X=0.492 $Y=1.79
+ $X2=0.492 $Y2=1.63
r105 13 21 54.3118 $w=2.67e-07 $l=2.57391e-07 $layer=POLY_cond $X=1.88 $Y=1.865
+ $X2=1.895 $Y2=1.615
r106 13 15 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=1.88 $Y=1.865
+ $X2=1.88 $Y2=2.44
r107 10 21 86.8062 $w=2.67e-07 $l=4.994e-07 $layer=POLY_cond $X=1.745 $Y=1.185
+ $X2=1.895 $Y2=1.615
r108 10 12 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=1.745 $Y=1.185
+ $X2=1.745 $Y2=0.74
r109 9 17 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=0.505 $Y=2.42
+ $X2=0.505 $Y2=1.845
r110 5 42 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=0.495 $Y=0.74
+ $X2=0.495 $Y2=1.3
.ends

.subckt PM_SKY130_FD_SC_HS__HA_2%A 3 5 7 10 12 14 15 22
c55 22 0 2.15518e-19 $X=1.315 $Y=1.632
r56 22 23 20.258 $w=3.45e-07 $l=1.45e-07 $layer=POLY_cond $X=1.315 $Y=1.632
+ $X2=1.46 $Y2=1.632
r57 20 22 12.5739 $w=3.45e-07 $l=9e-08 $layer=POLY_cond $X=1.225 $Y=1.632
+ $X2=1.315 $Y2=1.632
r58 18 20 37.7217 $w=3.45e-07 $l=2.7e-07 $layer=POLY_cond $X=0.955 $Y=1.632
+ $X2=1.225 $Y2=1.632
r59 17 18 9.77971 $w=3.45e-07 $l=7e-08 $layer=POLY_cond $X=0.885 $Y=1.632
+ $X2=0.955 $Y2=1.632
r60 15 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.225
+ $Y=1.595 $X2=1.225 $Y2=1.595
r61 12 23 22.2839 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=1.46 $Y=1.865
+ $X2=1.46 $Y2=1.632
r62 12 14 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=1.46 $Y=1.865
+ $X2=1.46 $Y2=2.44
r63 8 22 22.2839 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=1.315 $Y=1.4
+ $X2=1.315 $Y2=1.632
r64 8 10 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.315 $Y=1.4
+ $X2=1.315 $Y2=0.74
r65 5 18 22.2839 $w=1.5e-07 $l=2.13e-07 $layer=POLY_cond $X=0.955 $Y=1.845
+ $X2=0.955 $Y2=1.632
r66 5 7 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=0.955 $Y=1.845
+ $X2=0.955 $Y2=2.42
r67 1 17 22.2839 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=0.885 $Y=1.4
+ $X2=0.885 $Y2=1.632
r68 1 3 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.885 $Y=1.4 $X2=0.885
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HS__HA_2%A_27_74# 1 2 11 17 18 20 23 25 27 30 32 33 36
+ 38 39 41 42 45 48 49 51 52 54 56 59 62 64 72
c161 56 0 1.3969e-19 $X=0.73 $Y=2.065
c162 49 0 1.73571e-19 $X=2.87 $Y=1.445
c163 25 0 3.7278e-20 $X=5.255 $Y=1.765
r164 71 72 1.28191 $w=3.76e-07 $l=1e-08 $layer=POLY_cond $X=5.255 $Y=1.532
+ $X2=5.265 $Y2=1.532
r165 70 71 53.8404 $w=3.76e-07 $l=4.2e-07 $layer=POLY_cond $X=4.835 $Y=1.532
+ $X2=5.255 $Y2=1.532
r166 69 70 3.84574 $w=3.76e-07 $l=3e-08 $layer=POLY_cond $X=4.805 $Y=1.532
+ $X2=4.835 $Y2=1.532
r167 65 72 16.0239 $w=3.76e-07 $l=1.25e-07 $layer=POLY_cond $X=5.39 $Y=1.532
+ $X2=5.265 $Y2=1.532
r168 64 67 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=5.39 $Y=1.465
+ $X2=5.39 $Y2=1.63
r169 64 65 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.39
+ $Y=1.465 $X2=5.39 $Y2=1.465
r170 59 61 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=0.805 $Y=1.045
+ $X2=0.805 $Y2=1.195
r171 54 67 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=5.47 $Y=2.34
+ $X2=5.47 $Y2=1.63
r172 51 54 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.385 $Y=2.425
+ $X2=5.47 $Y2=2.34
r173 51 52 190.829 $w=1.68e-07 $l=2.925e-06 $layer=LI1_cond $X=5.385 $Y=2.425
+ $X2=2.46 $Y2=2.425
r174 48 49 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.87
+ $Y=1.445 $X2=2.87 $Y2=1.445
r175 46 62 3.70735 $w=2.5e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.46 $Y=1.445
+ $X2=2.375 $Y2=1.36
r176 46 48 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=2.46 $Y=1.445
+ $X2=2.87 $Y2=1.445
r177 45 52 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.375 $Y=2.34
+ $X2=2.46 $Y2=2.425
r178 44 62 2.76166 $w=1.7e-07 $l=2.5e-07 $layer=LI1_cond $X=2.375 $Y=1.61
+ $X2=2.375 $Y2=1.36
r179 44 45 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=2.375 $Y=1.61
+ $X2=2.375 $Y2=2.34
r180 43 61 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.89 $Y=1.195
+ $X2=0.805 $Y2=1.195
r181 42 62 3.70735 $w=2.5e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.29 $Y=1.195
+ $X2=2.375 $Y2=1.36
r182 42 43 91.3369 $w=1.68e-07 $l=1.4e-06 $layer=LI1_cond $X=2.29 $Y=1.195
+ $X2=0.89 $Y2=1.195
r183 41 56 0.716491 $w=1.7e-07 $l=1.16619e-07 $layer=LI1_cond $X=0.805 $Y=1.98
+ $X2=0.73 $Y2=2.065
r184 40 61 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=0.805 $Y=1.28
+ $X2=0.805 $Y2=1.195
r185 40 41 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=0.805 $Y=1.28
+ $X2=0.805 $Y2=1.98
r186 38 59 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.72 $Y=1.045
+ $X2=0.805 $Y2=1.045
r187 38 39 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=0.72 $Y=1.045
+ $X2=0.445 $Y2=1.045
r188 34 39 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.28 $Y=0.96
+ $X2=0.445 $Y2=1.045
r189 34 36 15.5405 $w=3.28e-07 $l=4.45e-07 $layer=LI1_cond $X=0.28 $Y=0.96
+ $X2=0.28 $Y2=0.515
r190 32 33 32.6715 $w=1.65e-07 $l=7.5e-08 $layer=POLY_cond $X=3.012 $Y=1.79
+ $X2=3.012 $Y2=1.865
r191 28 72 24.356 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=5.265 $Y=1.3
+ $X2=5.265 $Y2=1.532
r192 28 30 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=5.265 $Y=1.3
+ $X2=5.265 $Y2=0.74
r193 25 71 24.356 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=5.255 $Y=1.765
+ $X2=5.255 $Y2=1.532
r194 25 27 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=5.255 $Y=1.765
+ $X2=5.255 $Y2=2.4
r195 21 70 24.356 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=4.835 $Y=1.3
+ $X2=4.835 $Y2=1.532
r196 21 23 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=4.835 $Y=1.3
+ $X2=4.835 $Y2=0.74
r197 18 69 24.356 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=4.805 $Y=1.765
+ $X2=4.805 $Y2=1.532
r198 18 20 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=4.805 $Y=1.765
+ $X2=4.805 $Y2=2.4
r199 17 33 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=3.02 $Y=2.44
+ $X2=3.02 $Y2=1.865
r200 13 49 37.0704 $w=1.5e-07 $l=1.81659e-07 $layer=POLY_cond $X=3.005 $Y=1.61
+ $X2=2.97 $Y2=1.445
r201 13 32 92.2979 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=3.005 $Y=1.61
+ $X2=3.005 $Y2=1.79
r202 9 49 37.0704 $w=1.5e-07 $l=1.81659e-07 $layer=POLY_cond $X=2.935 $Y=1.28
+ $X2=2.97 $Y2=1.445
r203 9 11 276.894 $w=1.5e-07 $l=5.4e-07 $layer=POLY_cond $X=2.935 $Y=1.28
+ $X2=2.935 $Y2=0.74
r204 2 56 600 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=0.58
+ $Y=1.92 $X2=0.73 $Y2=2.065
r205 1 36 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__HA_2%A_391_388# 1 2 7 9 10 12 13 15 16 18 19 25 27
+ 28 30 33 36 41 47
c87 16 0 1.1278e-19 $X=4.405 $Y=1.22
r88 47 48 5.52752 $w=4.36e-07 $l=5e-08 $layer=POLY_cond $X=4.355 $Y=1.492
+ $X2=4.405 $Y2=1.492
r89 44 45 2.21101 $w=4.36e-07 $l=2e-08 $layer=POLY_cond $X=3.905 $Y=1.492
+ $X2=3.925 $Y2=1.492
r90 41 44 12.9125 $w=4.36e-07 $l=1.45186e-07 $layer=POLY_cond $X=3.815 $Y=1.385
+ $X2=3.905 $Y2=1.492
r91 40 41 57.7042 $w=3.3e-07 $l=3.3e-07 $layer=POLY_cond $X=3.485 $Y=1.385
+ $X2=3.815 $Y2=1.385
r92 39 40 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=3.485
+ $Y=1.385 $X2=3.485 $Y2=1.385
r93 36 39 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=3.405 $Y=1.025
+ $X2=3.405 $Y2=1.385
r94 34 47 21.0046 $w=4.36e-07 $l=1.9e-07 $layer=POLY_cond $X=4.165 $Y=1.492
+ $X2=4.355 $Y2=1.492
r95 34 45 26.5321 $w=4.36e-07 $l=2.4e-07 $layer=POLY_cond $X=4.165 $Y=1.492
+ $X2=3.925 $Y2=1.492
r96 33 39 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=4.165 $Y=1.385
+ $X2=3.49 $Y2=1.385
r97 33 34 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=4.165
+ $Y=1.385 $X2=4.165 $Y2=1.385
r98 29 39 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=3.405 $Y=1.55
+ $X2=3.405 $Y2=1.385
r99 29 30 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=3.405 $Y=1.55
+ $X2=3.405 $Y2=1.92
r100 27 36 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.32 $Y=1.025
+ $X2=3.405 $Y2=1.025
r101 27 28 33.5989 $w=1.68e-07 $l=5.15e-07 $layer=LI1_cond $X=3.32 $Y=1.025
+ $X2=2.805 $Y2=1.025
r102 23 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.72 $Y=0.94
+ $X2=2.805 $Y2=1.025
r103 23 25 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=2.72 $Y=0.94 $X2=2.72
+ $Y2=0.85
r104 19 30 7.14316 $w=2.5e-07 $l=1.62019e-07 $layer=LI1_cond $X=3.32 $Y=2.045
+ $X2=3.405 $Y2=1.92
r105 19 21 24.2013 $w=2.48e-07 $l=5.25e-07 $layer=LI1_cond $X=3.32 $Y=2.045
+ $X2=2.795 $Y2=2.045
r106 16 48 27.9822 $w=1.5e-07 $l=2.72e-07 $layer=POLY_cond $X=4.405 $Y=1.22
+ $X2=4.405 $Y2=1.492
r107 16 18 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=4.405 $Y=1.22
+ $X2=4.405 $Y2=0.74
r108 13 47 27.9822 $w=1.5e-07 $l=2.73e-07 $layer=POLY_cond $X=4.355 $Y=1.765
+ $X2=4.355 $Y2=1.492
r109 13 15 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=4.355 $Y=1.765
+ $X2=4.355 $Y2=2.4
r110 10 45 27.9822 $w=1.5e-07 $l=2.72e-07 $layer=POLY_cond $X=3.925 $Y=1.22
+ $X2=3.925 $Y2=1.492
r111 10 12 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=3.925 $Y=1.22
+ $X2=3.925 $Y2=0.74
r112 7 44 27.9822 $w=1.5e-07 $l=2.73e-07 $layer=POLY_cond $X=3.905 $Y=1.765
+ $X2=3.905 $Y2=1.492
r113 7 9 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.905 $Y=1.765
+ $X2=3.905 $Y2=2.4
r114 2 21 600 $w=1.7e-07 $l=9.09615e-07 $layer=licon1_PDIFF $count=1 $X=1.955
+ $Y=1.94 $X2=2.795 $Y2=2.085
r115 1 25 182 $w=1.7e-07 $l=2.98831e-07 $layer=licon1_NDIFF $count=1 $X=2.575
+ $Y=0.615 $X2=2.72 $Y2=0.85
.ends

.subckt PM_SKY130_FD_SC_HS__HA_2%VPWR 1 2 3 4 5 16 18 22 26 28 30 32 34 44 49 58
+ 63 71 73 77
c67 4 0 1.85225e-19 $X=4.43 $Y=1.84
r68 76 77 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r69 73 74 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r70 70 71 11.0283 $w=7.33e-07 $l=1.65e-07 $layer=LI1_cond $X=3.68 $Y=3.047
+ $X2=3.845 $Y2=3.047
r71 67 70 1.30185 $w=7.33e-07 $l=8e-08 $layer=LI1_cond $X=3.6 $Y=3.047 $X2=3.68
+ $Y2=3.047
r72 67 68 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r73 65 67 5.77698 $w=7.33e-07 $l=3.55e-07 $layer=LI1_cond $X=3.245 $Y=3.047
+ $X2=3.6 $Y2=3.047
r74 62 68 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=3.6 $Y2=3.33
r75 61 65 2.03415 $w=7.33e-07 $l=1.25e-07 $layer=LI1_cond $X=3.12 $Y=3.047
+ $X2=3.245 $Y2=3.047
r76 61 63 8.99415 $w=7.33e-07 $l=4e-08 $layer=LI1_cond $X=3.12 $Y=3.047 $X2=3.08
+ $Y2=3.047
r77 61 62 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r78 58 59 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r79 55 56 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r80 53 77 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=5.52 $Y2=3.33
r81 53 74 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=4.56 $Y2=3.33
r82 52 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r83 50 73 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.745 $Y=3.33
+ $X2=4.58 $Y2=3.33
r84 50 52 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=4.745 $Y=3.33
+ $X2=5.04 $Y2=3.33
r85 49 76 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=5.315 $Y=3.33
+ $X2=5.537 $Y2=3.33
r86 49 52 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=5.315 $Y=3.33
+ $X2=5.04 $Y2=3.33
r87 48 74 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=4.56 $Y2=3.33
r88 48 68 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=3.6 $Y2=3.33
r89 47 71 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=4.08 $Y=3.33
+ $X2=3.845 $Y2=3.33
r90 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r91 44 73 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.415 $Y=3.33
+ $X2=4.58 $Y2=3.33
r92 44 47 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=4.415 $Y=3.33
+ $X2=4.08 $Y2=3.33
r93 43 59 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r94 42 63 91.3369 $w=1.68e-07 $l=1.4e-06 $layer=LI1_cond $X=1.68 $Y=3.33
+ $X2=3.08 $Y2=3.33
r95 42 43 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r96 40 58 9.56655 $w=1.7e-07 $l=1.93e-07 $layer=LI1_cond $X=1.4 $Y=3.33
+ $X2=1.207 $Y2=3.33
r97 40 42 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=1.4 $Y=3.33 $X2=1.68
+ $Y2=3.33
r98 38 59 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r99 38 56 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r100 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r101 35 55 4.73185 $w=1.7e-07 $l=2.23e-07 $layer=LI1_cond $X=0.445 $Y=3.33
+ $X2=0.222 $Y2=3.33
r102 35 37 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=0.445 $Y=3.33
+ $X2=0.72 $Y2=3.33
r103 34 58 9.56655 $w=1.7e-07 $l=1.92e-07 $layer=LI1_cond $X=1.015 $Y=3.33
+ $X2=1.207 $Y2=3.33
r104 34 37 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=1.015 $Y=3.33
+ $X2=0.72 $Y2=3.33
r105 32 62 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.88 $Y=3.33
+ $X2=3.12 $Y2=3.33
r106 32 43 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=2.88 $Y=3.33
+ $X2=1.68 $Y2=3.33
r107 28 76 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=5.48 $Y=3.245
+ $X2=5.537 $Y2=3.33
r108 28 30 15.8897 $w=3.28e-07 $l=4.55e-07 $layer=LI1_cond $X=5.48 $Y=3.245
+ $X2=5.48 $Y2=2.79
r109 24 73 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.58 $Y=3.245
+ $X2=4.58 $Y2=3.33
r110 24 26 15.8897 $w=3.28e-07 $l=4.55e-07 $layer=LI1_cond $X=4.58 $Y=3.245
+ $X2=4.58 $Y2=2.79
r111 20 58 1.35792 $w=3.85e-07 $l=8.5e-08 $layer=LI1_cond $X=1.207 $Y=3.245
+ $X2=1.207 $Y2=3.33
r112 20 22 14.0688 $w=3.83e-07 $l=4.7e-07 $layer=LI1_cond $X=1.207 $Y=3.245
+ $X2=1.207 $Y2=2.775
r113 16 55 3.03433 $w=3.3e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.28 $Y=3.245
+ $X2=0.222 $Y2=3.33
r114 16 18 16.4136 $w=3.28e-07 $l=4.7e-07 $layer=LI1_cond $X=0.28 $Y=3.245
+ $X2=0.28 $Y2=2.775
r115 5 30 600 $w=1.7e-07 $l=1.02225e-06 $layer=licon1_PDIFF $count=1 $X=5.33
+ $Y=1.84 $X2=5.48 $Y2=2.79
r116 4 26 600 $w=1.7e-07 $l=1.02225e-06 $layer=licon1_PDIFF $count=1 $X=4.43
+ $Y=1.84 $X2=4.58 $Y2=2.79
r117 3 70 600 $w=1.7e-07 $l=1.13027e-06 $layer=licon1_PDIFF $count=1 $X=3.095
+ $Y=1.94 $X2=3.68 $Y2=2.815
r118 3 65 600 $w=1.7e-07 $l=9.47035e-07 $layer=licon1_PDIFF $count=1 $X=3.095
+ $Y=1.94 $X2=3.245 $Y2=2.815
r119 2 22 600 $w=1.7e-07 $l=9.3843e-07 $layer=licon1_PDIFF $count=1 $X=1.03
+ $Y=1.92 $X2=1.205 $Y2=2.775
r120 1 18 600 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.92 $X2=0.28 $Y2=2.775
.ends

.subckt PM_SKY130_FD_SC_HS__HA_2%SUM 1 2 7 12 13 14 18
c32 18 0 1.85225e-19 $X=4.505 $Y=1.995
r33 14 18 2.59474 $w=3.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.59 $Y=1.995
+ $X2=4.505 $Y2=1.995
r34 14 18 0.493904 $w=3.48e-07 $l=1.5e-08 $layer=LI1_cond $X=4.49 $Y=1.995
+ $X2=4.505 $Y2=1.995
r35 13 14 13.5 $w=3.48e-07 $l=4.1e-07 $layer=LI1_cond $X=4.08 $Y=1.995 $X2=4.49
+ $Y2=1.995
r36 12 14 5.34211 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=4.59 $Y=1.82
+ $X2=4.59 $Y2=1.995
r37 11 12 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=4.59 $Y=1.05
+ $X2=4.59 $Y2=1.82
r38 7 11 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.505 $Y=0.965
+ $X2=4.59 $Y2=1.05
r39 7 9 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=4.505 $Y=0.965
+ $X2=4.165 $Y2=0.965
r40 2 13 600 $w=1.7e-07 $l=2.17428e-07 $layer=licon1_PDIFF $count=1 $X=3.98
+ $Y=1.84 $X2=4.13 $Y2=1.995
r41 1 9 182 $w=1.7e-07 $l=6.72458e-07 $layer=licon1_NDIFF $count=1 $X=4 $Y=0.37
+ $X2=4.165 $Y2=0.965
.ends

.subckt PM_SKY130_FD_SC_HS__HA_2%COUT 1 2 10 11 13 14 25
c31 14 0 1.1278e-19 $X=4.955 $Y=0.84
c32 11 0 3.7278e-20 $X=5.03 $Y=1.82
r33 18 25 1.3969 $w=3.28e-07 $l=4e-08 $layer=LI1_cond $X=5.05 $Y=0.965 $X2=5.05
+ $Y2=0.925
r34 14 27 7.69388 $w=3.28e-07 $l=1.43e-07 $layer=LI1_cond $X=5.05 $Y=0.987
+ $X2=5.05 $Y2=1.13
r35 14 18 0.768295 $w=3.28e-07 $l=2.2e-08 $layer=LI1_cond $X=5.05 $Y=0.987
+ $X2=5.05 $Y2=0.965
r36 14 25 0.803218 $w=3.28e-07 $l=2.3e-08 $layer=LI1_cond $X=5.05 $Y=0.902
+ $X2=5.05 $Y2=0.925
r37 13 14 13.515 $w=3.28e-07 $l=3.87e-07 $layer=LI1_cond $X=5.05 $Y=0.515
+ $X2=5.05 $Y2=0.902
r38 11 27 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=4.97 $Y=1.82 $X2=4.97
+ $Y2=1.13
r39 10 11 8.8114 $w=3.28e-07 $l=1.75e-07 $layer=LI1_cond $X=5.03 $Y=1.995
+ $X2=5.03 $Y2=1.82
r40 2 10 600 $w=1.7e-07 $l=2.17428e-07 $layer=licon1_PDIFF $count=1 $X=4.88
+ $Y=1.84 $X2=5.03 $Y2=1.995
r41 1 13 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=4.91
+ $Y=0.37 $X2=5.05 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__HA_2%VGND 1 2 3 4 5 18 22 26 30 32 34 37 38 40 41 42
+ 51 55 60 66 69 73
r73 72 73 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r74 69 70 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r75 66 67 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r76 64 73 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=5.52
+ $Y2=0
r77 64 70 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=4.56
+ $Y2=0
r78 63 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r79 61 69 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.705 $Y=0 $X2=4.58
+ $Y2=0
r80 61 63 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=4.705 $Y=0 $X2=5.04
+ $Y2=0
r81 60 72 4.01252 $w=1.7e-07 $l=1.82e-07 $layer=LI1_cond $X=5.395 $Y=0 $X2=5.577
+ $Y2=0
r82 60 63 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=5.395 $Y=0 $X2=5.04
+ $Y2=0
r83 59 70 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=4.56
+ $Y2=0
r84 59 67 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=3.6
+ $Y2=0
r85 58 59 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r86 56 66 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.875 $Y=0 $X2=3.71
+ $Y2=0
r87 56 58 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=3.875 $Y=0 $X2=4.08
+ $Y2=0
r88 55 69 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.455 $Y=0 $X2=4.58
+ $Y2=0
r89 55 58 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=4.455 $Y=0 $X2=4.08
+ $Y2=0
r90 53 54 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r91 51 66 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.545 $Y=0 $X2=3.71
+ $Y2=0
r92 51 53 90.3583 $w=1.68e-07 $l=1.385e-06 $layer=LI1_cond $X=3.545 $Y=0
+ $X2=2.16 $Y2=0
r93 50 54 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r94 49 50 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r95 46 50 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r96 45 46 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r97 42 67 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=2.88 $Y=0 $X2=3.6
+ $Y2=0
r98 42 54 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=2.88 $Y=0 $X2=2.16
+ $Y2=0
r99 40 49 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=1.795 $Y=0 $X2=1.68
+ $Y2=0
r100 40 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.795 $Y=0 $X2=1.96
+ $Y2=0
r101 39 53 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=2.125 $Y=0 $X2=2.16
+ $Y2=0
r102 39 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.125 $Y=0 $X2=1.96
+ $Y2=0
r103 37 45 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=0.935 $Y=0
+ $X2=0.72 $Y2=0
r104 37 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.935 $Y=0 $X2=1.1
+ $Y2=0
r105 36 49 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=1.265 $Y=0
+ $X2=1.68 $Y2=0
r106 36 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.265 $Y=0 $X2=1.1
+ $Y2=0
r107 32 72 3.13065 $w=2.5e-07 $l=1.09864e-07 $layer=LI1_cond $X=5.52 $Y=0.085
+ $X2=5.577 $Y2=0
r108 32 34 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=5.52 $Y=0.085
+ $X2=5.52 $Y2=0.515
r109 28 69 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.58 $Y=0.085
+ $X2=4.58 $Y2=0
r110 28 30 20.5135 $w=2.48e-07 $l=4.45e-07 $layer=LI1_cond $X=4.58 $Y=0.085
+ $X2=4.58 $Y2=0.53
r111 24 66 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.71 $Y=0.085
+ $X2=3.71 $Y2=0
r112 24 26 15.5405 $w=3.28e-07 $l=4.45e-07 $layer=LI1_cond $X=3.71 $Y=0.085
+ $X2=3.71 $Y2=0.53
r113 20 41 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.96 $Y=0.085
+ $X2=1.96 $Y2=0
r114 20 22 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=1.96 $Y=0.085
+ $X2=1.96 $Y2=0.515
r115 16 38 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.1 $Y=0.085 $X2=1.1
+ $Y2=0
r116 16 18 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=1.1 $Y=0.085
+ $X2=1.1 $Y2=0.515
r117 5 34 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=5.34
+ $Y=0.37 $X2=5.48 $Y2=0.515
r118 4 30 182 $w=1.7e-07 $l=2.19089e-07 $layer=licon1_NDIFF $count=1 $X=4.48
+ $Y=0.37 $X2=4.62 $Y2=0.53
r119 3 26 182 $w=1.7e-07 $l=2.20907e-07 $layer=licon1_NDIFF $count=1 $X=3.565
+ $Y=0.37 $X2=3.71 $Y2=0.53
r120 2 22 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=1.82
+ $Y=0.37 $X2=1.96 $Y2=0.515
r121 1 18 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=0.96
+ $Y=0.37 $X2=1.1 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__HA_2%A_278_74# 1 2 7 12 13 14 17
r38 15 17 6.11144 $w=3.28e-07 $l=1.75e-07 $layer=LI1_cond $X=3.15 $Y=0.425
+ $X2=3.15 $Y2=0.6
r39 13 15 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.985 $Y=0.34
+ $X2=3.15 $Y2=0.425
r40 13 14 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=2.985 $Y=0.34
+ $X2=2.465 $Y2=0.34
r41 11 14 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.38 $Y=0.425
+ $X2=2.465 $Y2=0.34
r42 11 12 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=2.38 $Y=0.425
+ $X2=2.38 $Y2=0.77
r43 7 12 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.295 $Y=0.855
+ $X2=2.38 $Y2=0.77
r44 7 9 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=2.295 $Y=0.855
+ $X2=1.53 $Y2=0.855
r45 2 17 182 $w=1.7e-07 $l=2.91719e-07 $layer=licon1_NDIFF $count=1 $X=3.01
+ $Y=0.37 $X2=3.15 $Y2=0.6
r46 1 9 182 $w=1.7e-07 $l=5.50568e-07 $layer=licon1_NDIFF $count=1 $X=1.39
+ $Y=0.37 $X2=1.53 $Y2=0.855
.ends

