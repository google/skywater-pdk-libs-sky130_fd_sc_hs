* File: sky130_fd_sc_hs__o41a_4.spice
* Created: Tue Sep  1 20:19:23 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hs__o41a_4.pex.spice"
.subckt sky130_fd_sc_hs__o41a_4  VNB VPB B1 A4 A3 A1 A2 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A2	A2
* A1	A1
* A3	A3
* A4	A4
* B1	B1
* VPB	VPB
* VNB	VNB
MM1009 N_X_M1009_d N_A_110_48#_M1009_g N_VGND_M1009_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.2627 PD=1.02 PS=2.19 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75000.3
+ SB=75001.6 A=0.111 P=1.78 MULT=1
MM1013 N_X_M1009_d N_A_110_48#_M1013_g N_VGND_M1013_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1295 PD=1.02 PS=1.09 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.7
+ SB=75001.1 A=0.111 P=1.78 MULT=1
MM1015 N_X_M1015_d N_A_110_48#_M1015_g N_VGND_M1013_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1295 PD=1.02 PS=1.09 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75001.2
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1023 N_X_M1015_d N_A_110_48#_M1023_g N_VGND_M1023_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.2109 PD=1.02 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.6
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1005 N_A_523_124#_M1005_d N_B1_M1005_g N_A_110_48#_M1005_s VNB NLOWVT L=0.15
+ W=0.64 AD=0.1824 AS=0.0896 PD=1.85 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75004.5 A=0.096 P=1.58 MULT=1
MM1012 N_A_523_124#_M1012_d N_B1_M1012_g N_A_110_48#_M1005_s VNB NLOWVT L=0.15
+ W=0.64 AD=0.1184 AS=0.0896 PD=1.01 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.6 SB=75004 A=0.096 P=1.58 MULT=1
MM1003 N_A_523_124#_M1012_d N_A3_M1003_g N_VGND_M1003_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.1184 AS=0.19135 PD=1.01 PS=1.26 NRD=16.872 NRS=60 M=1 R=4.26667
+ SA=75001.2 SB=75003.5 A=0.096 P=1.58 MULT=1
MM1000 N_A_523_124#_M1000_d N_A4_M1000_g N_VGND_M1003_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.0896 AS=0.19135 PD=0.92 PS=1.26 NRD=0 NRS=0 M=1 R=4.26667 SA=75001.9
+ SB=75002.9 A=0.096 P=1.58 MULT=1
MM1027 N_A_523_124#_M1000_d N_A4_M1027_g N_VGND_M1027_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.0896 AS=0.0896 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667 SA=75002.3
+ SB=75002.4 A=0.096 P=1.58 MULT=1
MM1014 N_A_523_124#_M1014_d N_A3_M1014_g N_VGND_M1027_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.0928 AS=0.0896 PD=0.93 PS=0.92 NRD=0.936 NRS=0 M=1 R=4.26667 SA=75002.7
+ SB=75002 A=0.096 P=1.58 MULT=1
MM1008 N_A_523_124#_M1014_d N_A2_M1008_g N_VGND_M1008_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.0928 AS=0.0896 PD=0.93 PS=0.92 NRD=0.936 NRS=0 M=1 R=4.26667 SA=75003.2
+ SB=75001.6 A=0.096 P=1.58 MULT=1
MM1010 N_A_523_124#_M1010_d N_A1_M1010_g N_VGND_M1008_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.0896 AS=0.0896 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667 SA=75003.6
+ SB=75001.1 A=0.096 P=1.58 MULT=1
MM1011 N_A_523_124#_M1010_d N_A1_M1011_g N_VGND_M1011_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.0896 AS=0.113125 PD=0.92 PS=1.005 NRD=0 NRS=0 M=1 R=4.26667 SA=75004
+ SB=75000.7 A=0.096 P=1.58 MULT=1
MM1017 N_A_523_124#_M1017_d N_A2_M1017_g N_VGND_M1011_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.1824 AS=0.113125 PD=1.85 PS=1.005 NRD=0 NRS=13.116 M=1 R=4.26667
+ SA=75004.5 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1019 N_X_M1019_d N_A_110_48#_M1019_g N_VPWR_M1019_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.3304 PD=1.42 PS=2.83 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75002.3 A=0.168 P=2.54 MULT=1
MM1022 N_X_M1019_d N_A_110_48#_M1022_g N_VPWR_M1022_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.7 SB=75001.9 A=0.168 P=2.54 MULT=1
MM1024 N_X_M1024_d N_A_110_48#_M1024_g N_VPWR_M1022_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.1 SB=75001.4 A=0.168 P=2.54 MULT=1
MM1025 N_X_M1024_d N_A_110_48#_M1025_g N_VPWR_M1025_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.228743 PD=1.42 PS=1.72 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.6 SB=75001 A=0.168 P=2.54 MULT=1
MM1016 N_A_110_48#_M1016_d N_B1_M1016_g N_VPWR_M1025_s VPB PSHORT L=0.15 W=0.84
+ AD=0.126 AS=0.171557 PD=1.14 PS=1.29 NRD=2.3443 NRS=22.261 M=1 R=5.6
+ SA=75002.1 SB=75000.7 A=0.126 P=1.98 MULT=1
MM1020 N_A_110_48#_M1016_d N_B1_M1020_g N_VPWR_M1020_s VPB PSHORT L=0.15 W=0.84
+ AD=0.126 AS=0.2478 PD=1.14 PS=2.27 NRD=2.3443 NRS=2.3443 M=1 R=5.6 SA=75002.6
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1001 N_A_851_368#_M1001_d N_A3_M1001_g N_A_762_368#_M1001_s VPB PSHORT L=0.15
+ W=1.12 AD=0.168 AS=0.3304 PD=1.42 PS=2.83 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75003.5 A=0.168 P=2.54 MULT=1
MM1004 N_A_110_48#_M1004_d N_A4_M1004_g N_A_851_368#_M1001_d VPB PSHORT L=0.15
+ W=1.12 AD=0.1736 AS=0.168 PD=1.43 PS=1.42 NRD=2.6201 NRS=1.7533 M=1 R=7.46667
+ SA=75000.7 SB=75003.1 A=0.168 P=2.54 MULT=1
MM1026 N_A_110_48#_M1004_d N_A4_M1026_g N_A_851_368#_M1026_s VPB PSHORT L=0.15
+ W=1.12 AD=0.1736 AS=0.168 PD=1.43 PS=1.42 NRD=2.6201 NRS=1.7533 M=1 R=7.46667
+ SA=75001.1 SB=75002.6 A=0.168 P=2.54 MULT=1
MM1002 N_A_851_368#_M1026_s N_A3_M1002_g N_A_762_368#_M1002_s VPB PSHORT L=0.15
+ W=1.12 AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.6 SB=75002.2 A=0.168 P=2.54 MULT=1
MM1006 N_A_1213_368#_M1006_d N_A2_M1006_g N_A_762_368#_M1002_s VPB PSHORT L=0.15
+ W=1.12 AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75002 SB=75001.7 A=0.168 P=2.54 MULT=1
MM1007 N_VPWR_M1007_d N_A1_M1007_g N_A_1213_368#_M1006_d VPB PSHORT L=0.15
+ W=1.12 AD=0.1904 AS=0.168 PD=1.46 PS=1.42 NRD=5.2599 NRS=1.7533 M=1 R=7.46667
+ SA=75002.5 SB=75001.3 A=0.168 P=2.54 MULT=1
MM1021 N_VPWR_M1007_d N_A1_M1021_g N_A_1213_368#_M1021_s VPB PSHORT L=0.15
+ W=1.12 AD=0.1904 AS=0.196 PD=1.46 PS=1.47 NRD=5.2599 NRS=10.5395 M=1 R=7.46667
+ SA=75003 SB=75000.8 A=0.168 P=2.54 MULT=1
MM1018 N_A_1213_368#_M1021_s N_A2_M1018_g N_A_762_368#_M1018_s VPB PSHORT L=0.15
+ W=1.12 AD=0.196 AS=0.3864 PD=1.47 PS=2.93 NRD=1.7533 NRS=10.5395 M=1 R=7.46667
+ SA=75003.5 SB=75000.3 A=0.168 P=2.54 MULT=1
DX28_noxref VNB VPB NWDIODE A=15.8844 P=20.8
*
.include "sky130_fd_sc_hs__o41a_4.pxi.spice"
*
.ends
*
*
