# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_hs__einvn_8
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_hs__einvn_8 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  9.120000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  2.232000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.995000 1.350000 8.995000 1.780000 ;
    END
  END A
  PIN TE_B
    ANTENNAGATEAREA  1.623000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105000 1.180000 0.435000 1.630000 ;
    END
  END TE_B
  PIN Z
    ANTENNADIFFAREA  2.332400 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.925000 1.550000 5.725000 1.780000 ;
        RECT 5.455000 0.770000 6.645000 1.010000 ;
        RECT 5.455000 1.010000 8.505000 1.130000 ;
        RECT 5.455000 1.130000 5.725000 1.550000 ;
        RECT 5.555000 1.780000 5.725000 1.950000 ;
        RECT 5.555000 1.950000 8.555000 2.120000 ;
        RECT 5.555000 2.120000 5.725000 2.735000 ;
        RECT 6.315000 1.130000 8.505000 1.180000 ;
        RECT 6.425000 2.120000 6.755000 2.735000 ;
        RECT 7.325000 0.615000 7.495000 1.010000 ;
        RECT 7.325000 2.120000 7.655000 2.735000 ;
        RECT 8.175000 0.615000 8.505000 1.010000 ;
        RECT 8.225000 2.120000 8.555000 2.735000 ;
    END
  END Z
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 9.120000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 9.120000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 9.120000 0.085000 ;
      RECT 0.000000  3.245000 9.120000 3.415000 ;
      RECT 0.115000  1.820000 0.445000 3.245000 ;
      RECT 0.175000  0.085000 0.505000 0.990000 ;
      RECT 0.615000  1.130000 1.355000 1.335000 ;
      RECT 0.615000  1.335000 0.945000 2.980000 ;
      RECT 0.685000  0.325000 1.355000 1.130000 ;
      RECT 1.175000  1.665000 4.495000 1.835000 ;
      RECT 1.175000  1.835000 1.425000 2.980000 ;
      RECT 1.525000  0.350000 1.695000 1.300000 ;
      RECT 1.525000  1.300000 5.275000 1.380000 ;
      RECT 1.525000  1.380000 4.415000 1.470000 ;
      RECT 1.625000  2.005000 1.955000 3.245000 ;
      RECT 1.875000  0.085000 2.125000 1.130000 ;
      RECT 2.125000  1.835000 2.375000 2.980000 ;
      RECT 2.305000  0.350000 2.555000 1.300000 ;
      RECT 2.575000  2.005000 2.905000 3.245000 ;
      RECT 2.735000  0.085000 3.065000 1.130000 ;
      RECT 3.075000  1.835000 3.325000 2.980000 ;
      RECT 3.235000  0.350000 3.485000 1.300000 ;
      RECT 3.525000  2.005000 3.855000 3.245000 ;
      RECT 3.665000  0.085000 3.995000 1.130000 ;
      RECT 4.025000  1.835000 4.495000 1.950000 ;
      RECT 4.025000  1.950000 5.355000 2.120000 ;
      RECT 4.025000  2.120000 4.355000 2.980000 ;
      RECT 4.165000  0.350000 4.415000 1.210000 ;
      RECT 4.165000  1.210000 5.275000 1.300000 ;
      RECT 4.525000  2.290000 4.855000 3.245000 ;
      RECT 4.595000  0.085000 4.925000 1.040000 ;
      RECT 5.025000  2.120000 5.355000 2.905000 ;
      RECT 5.025000  2.905000 9.005000 3.075000 ;
      RECT 5.105000  0.255000 9.005000 0.425000 ;
      RECT 5.105000  0.425000 7.145000 0.600000 ;
      RECT 5.105000  0.600000 5.275000 1.210000 ;
      RECT 5.925000  2.290000 6.255000 2.905000 ;
      RECT 6.815000  0.600000 7.145000 0.825000 ;
      RECT 6.955000  2.290000 7.125000 2.905000 ;
      RECT 7.675000  0.425000 8.005000 0.825000 ;
      RECT 7.855000  2.290000 8.025000 2.905000 ;
      RECT 8.675000  0.425000 9.005000 1.130000 ;
      RECT 8.755000  1.950000 9.005000 2.905000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
      RECT 7.835000 -0.085000 8.005000 0.085000 ;
      RECT 7.835000  3.245000 8.005000 3.415000 ;
      RECT 8.315000 -0.085000 8.485000 0.085000 ;
      RECT 8.315000  3.245000 8.485000 3.415000 ;
      RECT 8.795000 -0.085000 8.965000 0.085000 ;
      RECT 8.795000  3.245000 8.965000 3.415000 ;
  END
END sky130_fd_sc_hs__einvn_8
