* File: sky130_fd_sc_hs__dfrtn_1.pex.spice
* Created: Thu Aug 27 20:38:30 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HS__DFRTN_1%D 2 3 4 5 7 10 14 16 21 22 23 28 29
r37 28 29 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.27
+ $Y=1.125 $X2=0.27 $Y2=1.125
r38 22 23 16.0907 $w=2.63e-07 $l=3.7e-07 $layer=LI1_cond $X=0.237 $Y=1.665
+ $X2=0.237 $Y2=2.035
r39 21 22 16.0907 $w=2.63e-07 $l=3.7e-07 $layer=LI1_cond $X=0.237 $Y=1.295
+ $X2=0.237 $Y2=1.665
r40 21 29 7.39303 $w=2.63e-07 $l=1.7e-07 $layer=LI1_cond $X=0.237 $Y=1.295
+ $X2=0.237 $Y2=1.125
r41 15 28 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=0.27 $Y=1.465
+ $X2=0.27 $Y2=1.125
r42 15 16 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.27 $Y=1.465
+ $X2=0.27 $Y2=1.63
r43 14 28 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=0.27 $Y=1.11
+ $X2=0.27 $Y2=1.125
r44 13 14 43.5886 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=0.352 $Y=0.96
+ $X2=0.352 $Y2=1.11
r45 10 13 194.851 $w=1.5e-07 $l=3.8e-07 $layer=POLY_cond $X=0.525 $Y=0.58
+ $X2=0.525 $Y2=0.96
r46 5 7 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=0.5 $Y=2.465 $X2=0.5
+ $Y2=2.75
r47 4 5 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=0.5 $Y=2.375 $X2=0.5
+ $Y2=2.465
r48 3 17 71.7872 $w=1.5e-07 $l=1.4e-07 $layer=POLY_cond $X=0.5 $Y=1.995 $X2=0.36
+ $Y2=1.995
r49 3 4 118.556 $w=1.8e-07 $l=3.05e-07 $layer=POLY_cond $X=0.5 $Y=2.07 $X2=0.5
+ $Y2=2.375
r50 2 17 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.36 $Y=1.92 $X2=0.36
+ $Y2=1.995
r51 2 16 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=0.36 $Y=1.92 $X2=0.36
+ $Y2=1.63
.ends

.subckt PM_SKY130_FD_SC_HS__DFRTN_1%RESET_B 3 6 7 9 12 15 16 18 21 24 25 27 28
+ 29 30 31 36 37 39 42 47 48 52 59
c201 42 0 1.59754e-19 $X=0.975 $Y=1.515
c202 7 0 1.83104e-19 $X=0.95 $Y=2.465
r203 52 55 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=8.545 $Y=1.63
+ $X2=8.545 $Y2=1.795
r204 52 54 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=8.545 $Y=1.63
+ $X2=8.545 $Y2=1.465
r205 47 50 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.985 $Y=1.635
+ $X2=4.985 $Y2=1.8
r206 47 49 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.985 $Y=1.635
+ $X2=4.985 $Y2=1.47
r207 47 48 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.985
+ $Y=1.635 $X2=4.985 $Y2=1.635
r208 43 59 6.03022 $w=4.28e-07 $l=2.25e-07 $layer=LI1_cond $X=0.975 $Y=1.565
+ $X2=1.2 $Y2=1.565
r209 42 45 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.975 $Y=1.515
+ $X2=0.975 $Y2=1.68
r210 42 44 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.975 $Y=1.515
+ $X2=0.975 $Y2=1.35
r211 42 43 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.975
+ $Y=1.515 $X2=0.975 $Y2=1.515
r212 39 59 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=1.665
+ $X2=1.2 $Y2=1.665
r213 37 52 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.545
+ $Y=1.63 $X2=8.545 $Y2=1.63
r214 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=1.665
+ $X2=8.4 $Y2=1.665
r215 33 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=1.665
+ $X2=5.04 $Y2=1.665
r216 31 33 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.185 $Y=1.665
+ $X2=5.04 $Y2=1.665
r217 30 36 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=8.255 $Y=1.665
+ $X2=8.4 $Y2=1.665
r218 30 31 3.7995 $w=1.4e-07 $l=3.07e-06 $layer=MET1_cond $X=8.255 $Y=1.665
+ $X2=5.185 $Y2=1.665
r219 29 39 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.345 $Y=1.665
+ $X2=1.2 $Y2=1.665
r220 28 33 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.895 $Y=1.665
+ $X2=5.04 $Y2=1.665
r221 28 29 4.39356 $w=1.4e-07 $l=3.55e-06 $layer=MET1_cond $X=4.895 $Y=1.665
+ $X2=1.345 $Y2=1.665
r222 25 27 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=8.62 $Y=2.465
+ $X2=8.62 $Y2=2.75
r223 24 25 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=8.62 $Y=2.375
+ $X2=8.62 $Y2=2.465
r224 24 55 225.452 $w=1.8e-07 $l=5.8e-07 $layer=POLY_cond $X=8.62 $Y=2.375
+ $X2=8.62 $Y2=1.795
r225 21 54 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=8.605 $Y=0.805
+ $X2=8.605 $Y2=1.465
r226 16 18 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=4.91 $Y=2.465
+ $X2=4.91 $Y2=2.75
r227 15 16 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=4.91 $Y=2.375
+ $X2=4.91 $Y2=2.465
r228 15 50 223.508 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.91 $Y=2.375
+ $X2=4.91 $Y2=1.8
r229 12 49 320.479 $w=1.5e-07 $l=6.25e-07 $layer=POLY_cond $X=4.895 $Y=0.845
+ $X2=4.895 $Y2=1.47
r230 7 9 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=0.95 $Y=2.465 $X2=0.95
+ $Y2=2.75
r231 6 7 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=0.95 $Y=2.375 $X2=0.95
+ $Y2=2.465
r232 6 45 270.153 $w=1.8e-07 $l=6.95e-07 $layer=POLY_cond $X=0.95 $Y=2.375
+ $X2=0.95 $Y2=1.68
r233 3 44 394.83 $w=1.5e-07 $l=7.7e-07 $layer=POLY_cond $X=0.915 $Y=0.58
+ $X2=0.915 $Y2=1.35
.ends

.subckt PM_SKY130_FD_SC_HS__DFRTN_1%CLK_N 1 3 4 6 7
c36 7 0 1.59754e-19 $X=1.68 $Y=1.295
r37 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.54
+ $Y=1.385 $X2=1.54 $Y2=1.385
r38 7 11 4.3606 $w=3.68e-07 $l=1.4e-07 $layer=LI1_cond $X=1.68 $Y=1.365 $X2=1.54
+ $Y2=1.365
r39 4 10 75.0274 $w=2.85e-07 $l=4.14439e-07 $layer=POLY_cond $X=1.455 $Y=1.765
+ $X2=1.527 $Y2=1.385
r40 4 6 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.455 $Y=1.765
+ $X2=1.455 $Y2=2.4
r41 1 10 38.666 $w=2.85e-07 $l=2.09893e-07 $layer=POLY_cond $X=1.425 $Y=1.22
+ $X2=1.527 $Y2=1.385
r42 1 3 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.425 $Y=1.22 $X2=1.425
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HS__DFRTN_1%A_507_368# 1 2 9 11 12 15 16 18 20 21 23 25
+ 26 28 30 32 33 37 38 43 44 47 48 49 51 52 53 55 57 58 60 61 64 70 71 72 79
c199 79 0 1.01786e-19 $X=7.42 $Y=1.29
c200 60 0 2.79847e-19 $X=7.255 $Y=1.29
c201 58 0 2.84298e-19 $X=7.08 $Y=1.29
c202 57 0 2.21313e-20 $X=6.535 $Y=1.21
c203 38 0 1.21692e-19 $X=3.55 $Y=1.94
c204 37 0 5.2417e-20 $X=3.55 $Y=1.94
c205 25 0 1.07929e-19 $X=6.9 $Y=1.29
c206 15 0 1.32597e-19 $X=4.01 $Y=2.375
c207 12 0 1.09116e-19 $X=3.92 $Y=2.015
r208 70 71 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.54
+ $Y=0.36 $X2=3.54 $Y2=0.36
r209 64 66 8.2628 $w=2.63e-07 $l=1.9e-07 $layer=LI1_cond $X=2.807 $Y=1.14
+ $X2=2.807 $Y2=1.33
r210 61 79 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=7.255 $Y=1.29
+ $X2=7.42 $Y2=1.29
r211 60 61 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=7.255
+ $Y=1.29 $X2=7.255 $Y2=1.29
r212 58 72 14.2244 $w=3.28e-07 $l=3.3e-07 $layer=LI1_cond $X=7.08 $Y=1.29
+ $X2=6.75 $Y2=1.29
r213 58 60 6.11144 $w=3.28e-07 $l=1.75e-07 $layer=LI1_cond $X=7.08 $Y=1.29
+ $X2=7.255 $Y2=1.29
r214 57 72 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=6.535 $Y=1.21
+ $X2=6.75 $Y2=1.21
r215 55 57 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.45 $Y=1.125
+ $X2=6.535 $Y2=1.21
r216 54 55 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=6.45 $Y=0.425
+ $X2=6.45 $Y2=1.125
r217 52 54 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.365 $Y=0.34
+ $X2=6.45 $Y2=0.425
r218 52 53 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=6.365 $Y=0.34
+ $X2=5.695 $Y2=0.34
r219 50 53 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.61 $Y=0.425
+ $X2=5.695 $Y2=0.34
r220 50 51 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=5.61 $Y=0.425
+ $X2=5.61 $Y2=0.79
r221 48 51 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.525 $Y=0.875
+ $X2=5.61 $Y2=0.79
r222 48 49 69.1551 $w=1.68e-07 $l=1.06e-06 $layer=LI1_cond $X=5.525 $Y=0.875
+ $X2=4.465 $Y2=0.875
r223 47 49 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.38 $Y=0.79
+ $X2=4.465 $Y2=0.875
r224 46 47 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=4.38 $Y=0.465
+ $X2=4.38 $Y2=0.79
r225 45 70 4.3182 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=3.705 $Y=0.36
+ $X2=3.62 $Y2=0.36
r226 44 46 6.91519 $w=2.1e-07 $l=1.41244e-07 $layer=LI1_cond $X=4.295 $Y=0.36
+ $X2=4.38 $Y2=0.465
r227 44 45 31.1602 $w=2.08e-07 $l=5.9e-07 $layer=LI1_cond $X=4.295 $Y=0.36
+ $X2=3.705 $Y2=0.36
r228 42 70 2.11342 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=3.62 $Y=0.465
+ $X2=3.62 $Y2=0.36
r229 42 43 50.8877 $w=1.68e-07 $l=7.8e-07 $layer=LI1_cond $X=3.62 $Y=0.465
+ $X2=3.62 $Y2=1.245
r230 38 76 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=3.55 $Y=1.94
+ $X2=3.55 $Y2=2.015
r231 37 38 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.55
+ $Y=1.94 $X2=3.55 $Y2=1.94
r232 35 68 3.13371 $w=3.3e-07 $l=1.4265e-07 $layer=LI1_cond $X=2.94 $Y=1.94
+ $X2=2.807 $Y2=1.96
r233 35 37 21.3027 $w=3.28e-07 $l=6.1e-07 $layer=LI1_cond $X=2.94 $Y=1.94
+ $X2=3.55 $Y2=1.94
r234 34 66 3.33486 $w=1.7e-07 $l=1.33e-07 $layer=LI1_cond $X=2.94 $Y=1.33
+ $X2=2.807 $Y2=1.33
r235 33 43 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.535 $Y=1.33
+ $X2=3.62 $Y2=1.245
r236 33 34 38.8182 $w=1.68e-07 $l=5.95e-07 $layer=LI1_cond $X=3.535 $Y=1.33
+ $X2=2.94 $Y2=1.33
r237 32 68 3.78913 $w=2.65e-07 $l=1.85e-07 $layer=LI1_cond $X=2.807 $Y=1.775
+ $X2=2.807 $Y2=1.96
r238 31 66 3.69652 $w=2.63e-07 $l=8.5e-08 $layer=LI1_cond $X=2.807 $Y=1.415
+ $X2=2.807 $Y2=1.33
r239 31 32 15.6558 $w=2.63e-07 $l=3.6e-07 $layer=LI1_cond $X=2.807 $Y=1.415
+ $X2=2.807 $Y2=1.775
r240 28 30 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=7.675 $Y=1.125
+ $X2=7.675 $Y2=0.805
r241 26 28 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=7.6 $Y=1.2
+ $X2=7.675 $Y2=1.125
r242 26 79 92.2979 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=7.6 $Y=1.2 $X2=7.42
+ $Y2=1.2
r243 25 61 62.0758 $w=3.3e-07 $l=3.55e-07 $layer=POLY_cond $X=6.9 $Y=1.29
+ $X2=7.255 $Y2=1.29
r244 21 23 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=6.81 $Y=1.885
+ $X2=6.81 $Y2=2.46
r245 20 21 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=6.81 $Y=1.795
+ $X2=6.81 $Y2=1.885
r246 19 25 18.0464 $w=4.25e-07 $l=2.05122e-07 $layer=POLY_cond $X=6.81 $Y=1.455
+ $X2=6.9 $Y2=1.29
r247 19 20 132.161 $w=1.8e-07 $l=3.4e-07 $layer=POLY_cond $X=6.81 $Y=1.455
+ $X2=6.81 $Y2=1.795
r248 16 18 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=4.01 $Y=2.465
+ $X2=4.01 $Y2=2.75
r249 15 16 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=4.01 $Y=2.375
+ $X2=4.01 $Y2=2.465
r250 14 15 104.952 $w=1.8e-07 $l=2.7e-07 $layer=POLY_cond $X=4.01 $Y=2.105
+ $X2=4.01 $Y2=2.375
r251 13 76 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=3.715 $Y=2.015
+ $X2=3.55 $Y2=2.015
r252 12 14 31.7871 $w=1.52e-07 $l=1.27279e-07 $layer=POLY_cond $X=3.92 $Y=2.015
+ $X2=4.01 $Y2=2.105
r253 12 13 79.6855 $w=1.8e-07 $l=2.05e-07 $layer=POLY_cond $X=3.92 $Y=2.015
+ $X2=3.715 $Y2=2.015
r254 9 71 19.9604 $w=1.5e-07 $l=1.95653e-07 $layer=POLY_cond $X=3.495 $Y=0.525
+ $X2=3.562 $Y2=0.36
r255 9 11 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=3.495 $Y=0.525
+ $X2=3.495 $Y2=0.845
r256 2 68 600 $w=1.7e-07 $l=2.91719e-07 $layer=licon1_PDIFF $count=1 $X=2.535
+ $Y=1.84 $X2=2.765 $Y2=1.98
r257 1 64 182 $w=1.7e-07 $l=7.37564e-07 $layer=licon1_NDIFF $count=1 $X=2.55
+ $Y=0.5 $X2=2.76 $Y2=1.14
.ends

.subckt PM_SKY130_FD_SC_HS__DFRTN_1%A_856_304# 1 2 8 9 11 14 18 19 22 28 31 32
+ 33 35 37 38
c99 37 0 2.21313e-20 $X=6.11 $Y=2.135
c100 35 0 2.66816e-19 $X=6.03 $Y=1.215
c101 31 0 2.7349e-20 $X=4.445 $Y=1.685
c102 8 0 5.2417e-20 $X=4.4 $Y=2.375
r103 37 39 0.373936 $w=8.33e-07 $l=5e-09 $layer=LI1_cond $X=6.282 $Y=2.135
+ $X2=6.282 $Y2=2.14
r104 37 38 11.6472 $w=8.33e-07 $l=1.65e-07 $layer=LI1_cond $X=6.282 $Y=2.135
+ $X2=6.282 $Y2=1.97
r105 32 42 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.445 $Y=1.685
+ $X2=4.445 $Y2=1.85
r106 32 41 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.445 $Y=1.685
+ $X2=4.445 $Y2=1.52
r107 31 33 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=4.445 $Y=1.685
+ $X2=4.445 $Y2=1.52
r108 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.445
+ $Y=1.685 $X2=4.445 $Y2=1.685
r109 28 39 11.3712 $w=7.08e-07 $l=6.75e-07 $layer=LI1_cond $X=6.345 $Y=2.815
+ $X2=6.345 $Y2=2.14
r110 24 35 3.70735 $w=2.5e-07 $l=1.18427e-07 $layer=LI1_cond $X=5.95 $Y=1.3
+ $X2=6.03 $Y2=1.215
r111 24 38 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.95 $Y=1.3
+ $X2=5.95 $Y2=1.97
r112 20 35 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.03 $Y=1.13
+ $X2=6.03 $Y2=1.215
r113 20 22 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=6.03 $Y=1.13
+ $X2=6.03 $Y2=0.76
r114 18 35 2.76166 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.865 $Y=1.215
+ $X2=6.03 $Y2=1.215
r115 18 19 81.877 $w=1.68e-07 $l=1.255e-06 $layer=LI1_cond $X=5.865 $Y=1.215
+ $X2=4.61 $Y2=1.215
r116 16 19 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.525 $Y=1.3
+ $X2=4.61 $Y2=1.215
r117 16 33 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=4.525 $Y=1.3
+ $X2=4.525 $Y2=1.52
r118 14 41 346.117 $w=1.5e-07 $l=6.75e-07 $layer=POLY_cond $X=4.535 $Y=0.845
+ $X2=4.535 $Y2=1.52
r119 9 11 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=4.4 $Y=2.465 $X2=4.4
+ $Y2=2.75
r120 8 9 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=4.4 $Y=2.375 $X2=4.4
+ $Y2=2.465
r121 8 42 204.073 $w=1.8e-07 $l=5.25e-07 $layer=POLY_cond $X=4.4 $Y=2.375
+ $X2=4.4 $Y2=1.85
r122 2 37 200 $w=1.7e-07 $l=2.40312e-07 $layer=licon1_PDIFF $count=3 $X=5.955
+ $Y=1.96 $X2=6.11 $Y2=2.135
r123 2 28 200 $w=1.7e-07 $l=9.29274e-07 $layer=licon1_PDIFF $count=3 $X=5.955
+ $Y=1.96 $X2=6.11 $Y2=2.815
r124 1 22 91 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=2 $X=5.89
+ $Y=0.595 $X2=6.03 $Y2=0.76
.ends

.subckt PM_SKY130_FD_SC_HS__DFRTN_1%A_714_127# 1 2 3 12 14 16 18 21 24 26 27 31
+ 33 35 41 43 44
c119 41 0 1.09116e-19 $X=3.97 $Y=2.75
r120 39 41 4.81032 $w=4.58e-07 $l=1.85e-07 $layer=LI1_cond $X=3.785 $Y=2.75
+ $X2=3.97 $Y2=2.75
r121 35 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.53
+ $Y=1.635 $X2=5.53 $Y2=1.635
r122 33 35 13.4452 $w=3.28e-07 $l=3.85e-07 $layer=LI1_cond $X=5.53 $Y=2.02
+ $X2=5.53 $Y2=1.635
r123 29 33 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=5.135 $Y=2.105
+ $X2=5.53 $Y2=2.105
r124 29 31 19.5566 $w=3.28e-07 $l=5.6e-07 $layer=LI1_cond $X=5.135 $Y=2.19
+ $X2=5.135 $Y2=2.75
r125 28 44 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.055 $Y=2.105
+ $X2=3.97 $Y2=2.105
r126 27 29 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=4.97 $Y=2.105
+ $X2=5.135 $Y2=2.105
r127 27 28 59.6952 $w=1.68e-07 $l=9.15e-07 $layer=LI1_cond $X=4.97 $Y=2.105
+ $X2=4.055 $Y2=2.105
r128 26 41 6.6364 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=3.97 $Y=2.52 $X2=3.97
+ $Y2=2.75
r129 25 44 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.97 $Y=2.19
+ $X2=3.97 $Y2=2.105
r130 25 26 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=3.97 $Y=2.19
+ $X2=3.97 $Y2=2.52
r131 24 44 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.97 $Y=2.02
+ $X2=3.97 $Y2=2.105
r132 24 43 61.6524 $w=1.68e-07 $l=9.45e-07 $layer=LI1_cond $X=3.97 $Y=2.02
+ $X2=3.97 $Y2=1.075
r133 19 43 6.71194 $w=2.48e-07 $l=1.25e-07 $layer=LI1_cond $X=4 $Y=0.95 $X2=4
+ $Y2=1.075
r134 19 21 4.37928 $w=2.48e-07 $l=9.5e-08 $layer=LI1_cond $X=4 $Y=0.95 $X2=4
+ $Y2=0.855
r135 18 36 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=5.74 $Y=1.635
+ $X2=5.53 $Y2=1.635
r136 14 18 59.8433 $w=2.19e-07 $l=2.62202e-07 $layer=POLY_cond $X=5.88 $Y=1.885
+ $X2=5.855 $Y2=1.635
r137 14 16 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=5.88 $Y=1.885
+ $X2=5.88 $Y2=2.46
r138 10 18 41.1355 $w=2.19e-07 $l=1.83916e-07 $layer=POLY_cond $X=5.815 $Y=1.47
+ $X2=5.855 $Y2=1.635
r139 10 12 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=5.815 $Y=1.47
+ $X2=5.815 $Y2=0.965
r140 3 31 600 $w=1.7e-07 $l=2.74955e-07 $layer=licon1_PDIFF $count=1 $X=4.985
+ $Y=2.54 $X2=5.135 $Y2=2.75
r141 2 39 600 $w=1.7e-07 $l=2.74955e-07 $layer=licon1_PDIFF $count=1 $X=3.635
+ $Y=2.54 $X2=3.785 $Y2=2.75
r142 1 21 182 $w=1.7e-07 $l=4.8775e-07 $layer=licon1_NDIFF $count=1 $X=3.57
+ $Y=0.635 $X2=3.96 $Y2=0.855
.ends

.subckt PM_SKY130_FD_SC_HS__DFRTN_1%A_300_74# 1 2 7 9 10 12 13 16 17 19 20 21 23
+ 27 28 29 33 34 36 37 38 39 41 42 49 51 55 56 59 62 63
c206 56 0 1.21652e-19 $X=7.475 $Y=1.86
c207 17 0 2.7349e-20 $X=3.81 $Y=1.47
r208 63 72 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.345 $Y=1.635
+ $X2=6.345 $Y2=1.47
r209 62 65 3.0228 $w=3.03e-07 $l=8e-08 $layer=LI1_cond $X=6.357 $Y=1.635
+ $X2=6.357 $Y2=1.715
r210 62 63 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.345
+ $Y=1.635 $X2=6.345 $Y2=1.635
r211 59 60 9.78865 $w=5.11e-07 $l=4.1e-07 $layer=LI1_cond $X=1.64 $Y=0.68
+ $X2=2.05 $Y2=0.68
r212 55 56 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=7.475
+ $Y=1.86 $X2=7.475 $Y2=1.86
r213 53 55 2.76586 $w=2.48e-07 $l=6e-08 $layer=LI1_cond $X=7.435 $Y=1.8
+ $X2=7.435 $Y2=1.86
r214 52 65 4.15824 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=6.51 $Y=1.715
+ $X2=6.357 $Y2=1.715
r215 51 53 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=7.31 $Y=1.715
+ $X2=7.435 $Y2=1.8
r216 51 52 52.1925 $w=1.68e-07 $l=8e-07 $layer=LI1_cond $X=7.31 $Y=1.715
+ $X2=6.51 $Y2=1.715
r217 49 50 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.08
+ $Y=1.515 $X2=2.08 $Y2=1.515
r218 47 49 15.2824 $w=2.28e-07 $l=3.05e-07 $layer=LI1_cond $X=2.05 $Y=1.82
+ $X2=2.05 $Y2=1.515
r219 46 60 5.43104 $w=2.3e-07 $l=3.3e-07 $layer=LI1_cond $X=2.05 $Y=1.01
+ $X2=2.05 $Y2=0.68
r220 46 49 25.3036 $w=2.28e-07 $l=5.05e-07 $layer=LI1_cond $X=2.05 $Y=1.01
+ $X2=2.05 $Y2=1.515
r221 42 47 7.07951 $w=3.25e-07 $l=2.11835e-07 $layer=LI1_cond $X=1.935 $Y=1.982
+ $X2=2.05 $Y2=1.82
r222 42 44 9.04224 $w=3.23e-07 $l=2.55e-07 $layer=LI1_cond $X=1.935 $Y=1.982
+ $X2=1.68 $Y2=1.982
r223 41 56 40.6942 $w=4.1e-07 $l=3e-07 $layer=POLY_cond $X=7.515 $Y=2.16
+ $X2=7.515 $Y2=1.86
r224 37 50 50.7098 $w=3.3e-07 $l=2.9e-07 $layer=POLY_cond $X=2.37 $Y=1.515
+ $X2=2.08 $Y2=1.515
r225 37 38 6.91837 $w=3.3e-07 $l=1.08995e-07 $layer=POLY_cond $X=2.37 $Y=1.515
+ $X2=2.46 $Y2=1.557
r226 34 41 44.6839 $w=3.29e-07 $l=3.70473e-07 $layer=POLY_cond $X=7.66 $Y=2.465
+ $X2=7.515 $Y2=2.16
r227 34 36 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=7.66 $Y=2.465
+ $X2=7.66 $Y2=2.75
r228 33 72 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=6.255 $Y=0.965
+ $X2=6.255 $Y2=1.47
r229 30 33 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=6.255 $Y=0.255
+ $X2=6.255 $Y2=0.965
r230 28 30 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=6.18 $Y=0.18
+ $X2=6.255 $Y2=0.255
r231 28 29 989.638 $w=1.5e-07 $l=1.93e-06 $layer=POLY_cond $X=6.18 $Y=0.18
+ $X2=4.25 $Y2=0.18
r232 25 40 13.7767 $w=1.5e-07 $l=1.5e-07 $layer=POLY_cond $X=4.175 $Y=1.13
+ $X2=4.175 $Y2=1.28
r233 25 27 146.138 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=4.175 $Y=1.13
+ $X2=4.175 $Y2=0.845
r234 24 29 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.175 $Y=0.255
+ $X2=4.25 $Y2=0.18
r235 24 27 302.532 $w=1.5e-07 $l=5.9e-07 $layer=POLY_cond $X=4.175 $Y=0.255
+ $X2=4.175 $Y2=0.845
r236 21 23 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=3.56 $Y=2.465
+ $X2=3.56 $Y2=2.75
r237 19 21 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.485 $Y=2.39
+ $X2=3.56 $Y2=2.465
r238 19 20 174.34 $w=1.5e-07 $l=3.4e-07 $layer=POLY_cond $X=3.485 $Y=2.39
+ $X2=3.145 $Y2=2.39
r239 18 39 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.145 $Y=1.47
+ $X2=3.07 $Y2=1.47
r240 17 40 80.0453 $w=2.4e-07 $l=4.50083e-07 $layer=POLY_cond $X=3.81 $Y=1.47
+ $X2=4.175 $Y2=1.28
r241 17 18 340.989 $w=1.5e-07 $l=6.65e-07 $layer=POLY_cond $X=3.81 $Y=1.47
+ $X2=3.145 $Y2=1.47
r242 16 20 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.07 $Y=2.315
+ $X2=3.145 $Y2=2.39
r243 15 39 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.07 $Y=1.545
+ $X2=3.07 $Y2=1.47
r244 15 16 394.83 $w=1.5e-07 $l=7.7e-07 $layer=POLY_cond $X=3.07 $Y=1.545
+ $X2=3.07 $Y2=2.315
r245 14 38 6.91837 $w=1.5e-07 $l=1.26214e-07 $layer=POLY_cond $X=2.55 $Y=1.47
+ $X2=2.46 $Y2=1.557
r246 13 39 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.995 $Y=1.47
+ $X2=3.07 $Y2=1.47
r247 13 14 228.181 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=2.995 $Y=1.47
+ $X2=2.55 $Y2=1.47
r248 10 38 18.1359 $w=1.5e-07 $l=2.14369e-07 $layer=POLY_cond $X=2.475 $Y=1.35
+ $X2=2.46 $Y2=1.557
r249 10 12 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=2.475 $Y=1.35
+ $X2=2.475 $Y2=0.87
r250 7 38 18.1359 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=2.46 $Y=1.765
+ $X2=2.46 $Y2=1.557
r251 7 9 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.46 $Y=1.765
+ $X2=2.46 $Y2=2.4
r252 2 44 600 $w=1.7e-07 $l=2.43721e-07 $layer=licon1_PDIFF $count=1 $X=1.53
+ $Y=1.84 $X2=1.68 $Y2=2.02
r253 1 59 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.5
+ $Y=0.37 $X2=1.64 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__DFRTN_1%A_1598_93# 1 2 9 11 13 14 21 23 26 27 31
c89 9 0 1.58195e-19 $X=8.065 $Y=0.805
r90 29 31 8.03677 $w=3.78e-07 $l=2.65e-07 $layer=LI1_cond $X=9.21 $Y=0.765
+ $X2=9.475 $Y2=0.765
r91 25 31 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=9.475 $Y=0.955
+ $X2=9.475 $Y2=0.765
r92 25 26 65.8931 $w=1.68e-07 $l=1.01e-06 $layer=LI1_cond $X=9.475 $Y=0.955
+ $X2=9.475 $Y2=1.965
r93 24 27 6.08426 $w=2.7e-07 $l=2.29619e-07 $layer=LI1_cond $X=9.05 $Y=2.05
+ $X2=8.865 $Y2=2.15
r94 23 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.39 $Y=2.05
+ $X2=9.475 $Y2=1.965
r95 23 24 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=9.39 $Y=2.05
+ $X2=9.05 $Y2=2.05
r96 19 27 0.630948 $w=3.3e-07 $l=1.94743e-07 $layer=LI1_cond $X=8.845 $Y=2.335
+ $X2=8.865 $Y2=2.15
r97 19 21 14.4928 $w=3.28e-07 $l=4.15e-07 $layer=LI1_cond $X=8.845 $Y=2.335
+ $X2=8.845 $Y2=2.75
r98 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.155
+ $Y=2.17 $X2=8.155 $Y2=2.17
r99 14 27 6.08426 $w=2.7e-07 $l=1.85e-07 $layer=LI1_cond $X=8.68 $Y=2.15
+ $X2=8.865 $Y2=2.15
r100 14 16 16.3522 $w=3.68e-07 $l=5.25e-07 $layer=LI1_cond $X=8.68 $Y=2.15
+ $X2=8.155 $Y2=2.15
r101 11 17 60.4771 $w=2.87e-07 $l=3.30379e-07 $layer=POLY_cond $X=8.08 $Y=2.465
+ $X2=8.155 $Y2=2.17
r102 11 13 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=8.08 $Y=2.465
+ $X2=8.08 $Y2=2.75
r103 7 17 38.6443 $w=2.87e-07 $l=2.05122e-07 $layer=POLY_cond $X=8.065 $Y=2.005
+ $X2=8.155 $Y2=2.17
r104 7 9 615.319 $w=1.5e-07 $l=1.2e-06 $layer=POLY_cond $X=8.065 $Y=2.005
+ $X2=8.065 $Y2=0.805
r105 2 21 600 $w=1.7e-07 $l=2.74955e-07 $layer=licon1_PDIFF $count=1 $X=8.695
+ $Y=2.54 $X2=8.845 $Y2=2.75
r106 1 29 182 $w=1.7e-07 $l=2.29565e-07 $layer=licon1_NDIFF $count=1 $X=9.07
+ $Y=0.595 $X2=9.21 $Y2=0.765
.ends

.subckt PM_SKY130_FD_SC_HS__DFRTN_1%A_1266_119# 1 2 7 9 10 11 12 14 15 17 19 21
+ 22 24 26 29 33 38 40 41 46 48 50 51
c138 48 0 2.64234e-19 $X=7.815 $Y=1.21
r139 50 51 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=9.085
+ $Y=1.29 $X2=9.085 $Y2=1.29
r140 46 47 20.5133 $w=2.26e-07 $l=3.8e-07 $layer=LI1_cond $X=7.435 $Y=2.7
+ $X2=7.815 $Y2=2.7
r141 42 48 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.9 $Y=1.21
+ $X2=7.815 $Y2=1.21
r142 41 50 4.79851 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=8.92 $Y=1.21
+ $X2=9.07 $Y2=1.21
r143 41 42 66.5455 $w=1.68e-07 $l=1.02e-06 $layer=LI1_cond $X=8.92 $Y=1.21
+ $X2=7.9 $Y2=1.21
r144 40 47 2.4068 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.815 $Y=2.535
+ $X2=7.815 $Y2=2.7
r145 39 48 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.815 $Y=1.295
+ $X2=7.815 $Y2=1.21
r146 39 40 80.8984 $w=1.68e-07 $l=1.24e-06 $layer=LI1_cond $X=7.815 $Y=1.295
+ $X2=7.815 $Y2=2.535
r147 38 48 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.815 $Y=1.125
+ $X2=7.815 $Y2=1.21
r148 37 38 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=7.815 $Y=0.955
+ $X2=7.815 $Y2=1.125
r149 33 46 1.22073 $w=3.3e-07 $l=1.75152e-07 $layer=LI1_cond $X=7.435 $Y=2.7
+ $X2=7.435 $Y2=2.7
r150 33 35 13.969 $w=3.28e-07 $l=4e-07 $layer=LI1_cond $X=7.435 $Y=2.7 $X2=7.035
+ $Y2=2.7
r151 29 37 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=7.73 $Y=0.79
+ $X2=7.815 $Y2=0.955
r152 29 31 9.42908 $w=3.28e-07 $l=2.7e-07 $layer=LI1_cond $X=7.73 $Y=0.79
+ $X2=7.46 $Y2=0.79
r153 27 51 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=9.085 $Y=1.63
+ $X2=9.085 $Y2=1.29
r154 27 28 50.3824 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=9.085 $Y=1.63
+ $X2=9.085 $Y2=1.97
r155 25 51 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=9.085 $Y=1.275
+ $X2=9.085 $Y2=1.29
r156 25 26 13.5877 $w=2.4e-07 $l=7.5e-08 $layer=POLY_cond $X=9.085 $Y=1.275
+ $X2=9.085 $Y2=1.2
r157 22 24 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=10.04 $Y=2.045
+ $X2=10.04 $Y2=2.54
r158 19 21 122.107 $w=1.5e-07 $l=3.8e-07 $layer=POLY_cond $X=10.03 $Y=1.125
+ $X2=10.03 $Y2=0.745
r159 18 28 18.414 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.25 $Y=1.97
+ $X2=9.085 $Y2=1.97
r160 17 22 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=9.965 $Y=1.97
+ $X2=10.04 $Y2=2.045
r161 17 18 366.628 $w=1.5e-07 $l=7.15e-07 $layer=POLY_cond $X=9.965 $Y=1.97
+ $X2=9.25 $Y2=1.97
r162 16 26 12.1617 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.25 $Y=1.2
+ $X2=9.085 $Y2=1.2
r163 15 19 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=9.955 $Y=1.2
+ $X2=10.03 $Y2=1.125
r164 15 16 361.5 $w=1.5e-07 $l=7.05e-07 $layer=POLY_cond $X=9.955 $Y=1.2
+ $X2=9.25 $Y2=1.2
r165 12 14 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=9.07 $Y=2.465
+ $X2=9.07 $Y2=2.75
r166 11 12 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=9.07 $Y=2.375
+ $X2=9.07 $Y2=2.465
r167 10 28 19.4594 $w=2.93e-07 $l=8.21584e-08 $layer=POLY_cond $X=9.07 $Y=2.045
+ $X2=9.085 $Y2=1.97
r168 10 11 128.274 $w=1.8e-07 $l=3.3e-07 $layer=POLY_cond $X=9.07 $Y=2.045
+ $X2=9.07 $Y2=2.375
r169 7 26 13.5877 $w=2.4e-07 $l=1.21861e-07 $layer=POLY_cond $X=8.995 $Y=1.125
+ $X2=9.085 $Y2=1.2
r170 7 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=8.995 $Y=1.125
+ $X2=8.995 $Y2=0.805
r171 2 46 600 $w=1.7e-07 $l=9.77036e-07 $layer=licon1_PDIFF $count=1 $X=6.885
+ $Y=1.96 $X2=7.435 $Y2=2.7
r172 2 35 600 $w=1.7e-07 $l=8.11542e-07 $layer=licon1_PDIFF $count=1 $X=6.885
+ $Y=1.96 $X2=7.035 $Y2=2.7
r173 1 31 91 $w=1.7e-07 $l=1.22362e-06 $layer=licon1_NDIFF $count=2 $X=6.33
+ $Y=0.595 $X2=7.46 $Y2=0.79
.ends

.subckt PM_SKY130_FD_SC_HS__DFRTN_1%A_1934_94# 1 2 7 9 10 12 13 15 19 24 27 31
r60 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.48
+ $Y=1.485 $X2=10.48 $Y2=1.485
r61 25 31 0.364692 $w=3.3e-07 $l=1.25e-07 $layer=LI1_cond $X=9.98 $Y=1.485
+ $X2=9.855 $Y2=1.485
r62 25 27 17.4613 $w=3.28e-07 $l=5e-07 $layer=LI1_cond $X=9.98 $Y=1.485
+ $X2=10.48 $Y2=1.485
r63 24 30 1.61342 $w=2.48e-07 $l=3.5e-08 $layer=LI1_cond $X=9.855 $Y=2.27
+ $X2=9.855 $Y2=2.305
r64 21 31 6.46576 $w=2.5e-07 $l=1.65e-07 $layer=LI1_cond $X=9.855 $Y=1.65
+ $X2=9.855 $Y2=1.485
r65 21 24 28.5806 $w=2.48e-07 $l=6.2e-07 $layer=LI1_cond $X=9.855 $Y=1.65
+ $X2=9.855 $Y2=2.27
r66 17 31 6.46576 $w=2.5e-07 $l=1.65e-07 $layer=LI1_cond $X=9.855 $Y=1.32
+ $X2=9.855 $Y2=1.485
r67 17 19 26.5062 $w=2.48e-07 $l=5.75e-07 $layer=LI1_cond $X=9.855 $Y=1.32
+ $X2=9.855 $Y2=0.745
r68 13 30 6.46688 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=9.815 $Y=2.47
+ $X2=9.815 $Y2=2.305
r69 13 15 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=9.815 $Y=2.47
+ $X2=9.815 $Y2=2.815
r70 10 28 57.6553 $w=2.91e-07 $l=3.10805e-07 $layer=POLY_cond $X=10.545 $Y=1.765
+ $X2=10.48 $Y2=1.485
r71 10 12 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=10.545 $Y=1.765
+ $X2=10.545 $Y2=2.4
r72 7 28 38.6072 $w=2.91e-07 $l=1.92678e-07 $layer=POLY_cond $X=10.54 $Y=1.32
+ $X2=10.48 $Y2=1.485
r73 7 9 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=10.54 $Y=1.32 $X2=10.54
+ $Y2=0.84
r74 2 24 600 $w=1.7e-07 $l=2.03101e-07 $layer=licon1_PDIFF $count=1 $X=9.69
+ $Y=2.12 $X2=9.815 $Y2=2.27
r75 2 15 600 $w=1.7e-07 $l=7.54917e-07 $layer=licon1_PDIFF $count=1 $X=9.69
+ $Y=2.12 $X2=9.815 $Y2=2.815
r76 1 19 182 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_NDIFF $count=1 $X=9.67
+ $Y=0.47 $X2=9.815 $Y2=0.745
.ends

.subckt PM_SKY130_FD_SC_HS__DFRTN_1%VPWR 1 2 3 4 5 6 7 8 25 27 31 35 39 41 45 49
+ 53 57 60 61 63 64 65 67 72 77 92 101 102 108 111 114 117 120
r134 120 121 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.36 $Y=3.33
+ $X2=9.36 $Y2=3.33
r135 114 115 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r136 111 112 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r137 108 109 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r138 105 106 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r139 101 102 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.8 $Y=3.33
+ $X2=10.8 $Y2=3.33
r140 99 102 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=9.84 $Y=3.33
+ $X2=10.8 $Y2=3.33
r141 99 121 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.84 $Y=3.33
+ $X2=9.36 $Y2=3.33
r142 98 99 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.84 $Y=3.33
+ $X2=9.84 $Y2=3.33
r143 96 120 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=9.46 $Y=3.33
+ $X2=9.335 $Y2=3.33
r144 96 98 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=9.46 $Y=3.33
+ $X2=9.84 $Y2=3.33
r145 95 121 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=3.33
+ $X2=9.36 $Y2=3.33
r146 94 95 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r147 92 120 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=9.21 $Y=3.33
+ $X2=9.335 $Y2=3.33
r148 92 94 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=9.21 $Y=3.33
+ $X2=8.88 $Y2=3.33
r149 91 95 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=7.92 $Y=3.33
+ $X2=8.88 $Y2=3.33
r150 90 91 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r151 88 91 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=6 $Y=3.33
+ $X2=7.92 $Y2=3.33
r152 87 90 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=6 $Y=3.33 $X2=7.92
+ $Y2=3.33
r153 87 88 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r154 85 117 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.82 $Y=3.33
+ $X2=5.655 $Y2=3.33
r155 85 87 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=5.82 $Y=3.33 $X2=6
+ $Y2=3.33
r156 84 115 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=4.56 $Y2=3.33
r157 83 84 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r158 81 84 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=4.08 $Y2=3.33
r159 81 112 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=2.16 $Y2=3.33
r160 80 83 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=2.64 $Y=3.33
+ $X2=4.08 $Y2=3.33
r161 80 81 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r162 78 111 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.4 $Y=3.33
+ $X2=2.235 $Y2=3.33
r163 78 80 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=2.4 $Y=3.33
+ $X2=2.64 $Y2=3.33
r164 77 114 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.46 $Y=3.33
+ $X2=4.625 $Y2=3.33
r165 77 83 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=4.46 $Y=3.33
+ $X2=4.08 $Y2=3.33
r166 76 112 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r167 76 109 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r168 75 76 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r169 73 108 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.39 $Y=3.33
+ $X2=1.225 $Y2=3.33
r170 73 75 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=1.39 $Y=3.33
+ $X2=1.68 $Y2=3.33
r171 72 111 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.07 $Y=3.33
+ $X2=2.235 $Y2=3.33
r172 72 75 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=2.07 $Y=3.33
+ $X2=1.68 $Y2=3.33
r173 71 109 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r174 71 106 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r175 70 71 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r176 68 105 4.746 $w=1.7e-07 $l=2.2e-07 $layer=LI1_cond $X=0.44 $Y=3.33 $X2=0.22
+ $Y2=3.33
r177 68 70 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=0.44 $Y=3.33
+ $X2=0.72 $Y2=3.33
r178 67 108 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.06 $Y=3.33
+ $X2=1.225 $Y2=3.33
r179 67 70 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=1.06 $Y=3.33
+ $X2=0.72 $Y2=3.33
r180 65 88 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=3.33 $X2=6
+ $Y2=3.33
r181 65 115 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=4.56 $Y2=3.33
r182 65 117 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r183 63 98 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=10.15 $Y=3.33
+ $X2=9.84 $Y2=3.33
r184 63 64 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=10.15 $Y=3.33
+ $X2=10.275 $Y2=3.33
r185 62 101 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=10.4 $Y=3.33
+ $X2=10.8 $Y2=3.33
r186 62 64 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=10.4 $Y=3.33
+ $X2=10.275 $Y2=3.33
r187 60 90 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=8.14 $Y=3.33
+ $X2=7.92 $Y2=3.33
r188 60 61 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.14 $Y=3.33
+ $X2=8.305 $Y2=3.33
r189 59 94 26.7487 $w=1.68e-07 $l=4.1e-07 $layer=LI1_cond $X=8.47 $Y=3.33
+ $X2=8.88 $Y2=3.33
r190 59 61 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.47 $Y=3.33
+ $X2=8.305 $Y2=3.33
r191 55 64 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=10.275 $Y=3.245
+ $X2=10.275 $Y2=3.33
r192 55 57 45.1758 $w=2.48e-07 $l=9.8e-07 $layer=LI1_cond $X=10.275 $Y=3.245
+ $X2=10.275 $Y2=2.265
r193 51 120 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=9.335 $Y=3.245
+ $X2=9.335 $Y2=3.33
r194 51 53 22.8184 $w=2.48e-07 $l=4.95e-07 $layer=LI1_cond $X=9.335 $Y=3.245
+ $X2=9.335 $Y2=2.75
r195 47 61 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.305 $Y=3.245
+ $X2=8.305 $Y2=3.33
r196 47 49 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=8.305 $Y=3.245
+ $X2=8.305 $Y2=2.75
r197 43 117 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.655 $Y=3.245
+ $X2=5.655 $Y2=3.33
r198 43 45 27.938 $w=3.28e-07 $l=8e-07 $layer=LI1_cond $X=5.655 $Y=3.245
+ $X2=5.655 $Y2=2.445
r199 42 114 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.79 $Y=3.33
+ $X2=4.625 $Y2=3.33
r200 41 117 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.49 $Y=3.33
+ $X2=5.655 $Y2=3.33
r201 41 42 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=5.49 $Y=3.33 $X2=4.79
+ $Y2=3.33
r202 37 114 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.625 $Y=3.245
+ $X2=4.625 $Y2=3.33
r203 37 39 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=4.625 $Y=3.245
+ $X2=4.625 $Y2=2.75
r204 33 111 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.235 $Y=3.245
+ $X2=2.235 $Y2=3.33
r205 33 35 14.8421 $w=3.28e-07 $l=4.25e-07 $layer=LI1_cond $X=2.235 $Y=3.245
+ $X2=2.235 $Y2=2.82
r206 29 108 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.225 $Y=3.245
+ $X2=1.225 $Y2=3.33
r207 29 31 16.4136 $w=3.28e-07 $l=4.7e-07 $layer=LI1_cond $X=1.225 $Y=3.245
+ $X2=1.225 $Y2=2.775
r208 25 105 3.02018 $w=3.3e-07 $l=1.09087e-07 $layer=LI1_cond $X=0.275 $Y=3.245
+ $X2=0.22 $Y2=3.33
r209 25 27 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=0.275 $Y=3.245
+ $X2=0.275 $Y2=2.75
r210 8 57 300 $w=1.7e-07 $l=2.62678e-07 $layer=licon1_PDIFF $count=2 $X=10.115
+ $Y=2.12 $X2=10.315 $Y2=2.265
r211 7 53 600 $w=1.7e-07 $l=2.74955e-07 $layer=licon1_PDIFF $count=1 $X=9.145
+ $Y=2.54 $X2=9.295 $Y2=2.75
r212 6 49 600 $w=1.7e-07 $l=2.74955e-07 $layer=licon1_PDIFF $count=1 $X=8.155
+ $Y=2.54 $X2=8.305 $Y2=2.75
r213 5 45 300 $w=1.7e-07 $l=5.43921e-07 $layer=licon1_PDIFF $count=2 $X=5.53
+ $Y=1.96 $X2=5.655 $Y2=2.445
r214 4 39 600 $w=1.7e-07 $l=2.74955e-07 $layer=licon1_PDIFF $count=1 $X=4.475
+ $Y=2.54 $X2=4.625 $Y2=2.75
r215 3 35 600 $w=1.7e-07 $l=1.05e-06 $layer=licon1_PDIFF $count=1 $X=2.09
+ $Y=1.84 $X2=2.235 $Y2=2.82
r216 2 31 600 $w=1.7e-07 $l=3.19726e-07 $layer=licon1_PDIFF $count=1 $X=1.025
+ $Y=2.54 $X2=1.225 $Y2=2.775
r217 1 27 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.54 $X2=0.275 $Y2=2.75
.ends

.subckt PM_SKY130_FD_SC_HS__DFRTN_1%A_33_74# 1 2 3 4 14 17 19 20 22 23 24 25 29
+ 34 38 39
c116 25 0 2.54289e-19 $X=3.17 $Y=2.4
c117 20 0 1.83104e-19 $X=1.23 $Y=2.4
c118 14 0 1.52323e-19 $X=0.625 $Y=2.18
r119 39 42 6.22319 $w=2.48e-07 $l=1.35e-07 $layer=LI1_cond $X=3.24 $Y=0.72
+ $X2=3.24 $Y2=0.855
r120 32 34 8.25044 $w=4.38e-07 $l=3.15e-07 $layer=LI1_cond $X=0.31 $Y=0.57
+ $X2=0.625 $Y2=0.57
r121 27 29 12.2159 $w=2.48e-07 $l=2.65e-07 $layer=LI1_cond $X=3.295 $Y=2.485
+ $X2=3.295 $Y2=2.75
r122 26 38 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.505 $Y=2.4
+ $X2=2.42 $Y2=2.4
r123 25 27 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=3.17 $Y=2.4
+ $X2=3.295 $Y2=2.485
r124 25 26 43.385 $w=1.68e-07 $l=6.65e-07 $layer=LI1_cond $X=3.17 $Y=2.4
+ $X2=2.505 $Y2=2.4
r125 23 39 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.115 $Y=0.72
+ $X2=3.24 $Y2=0.72
r126 23 24 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=3.115 $Y=0.72
+ $X2=2.505 $Y2=0.72
r127 22 38 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.42 $Y=2.315
+ $X2=2.42 $Y2=2.4
r128 21 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.42 $Y=0.805
+ $X2=2.505 $Y2=0.72
r129 21 22 98.5134 $w=1.68e-07 $l=1.51e-06 $layer=LI1_cond $X=2.42 $Y=0.805
+ $X2=2.42 $Y2=2.315
r130 19 38 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.335 $Y=2.4
+ $X2=2.42 $Y2=2.4
r131 19 20 72.0909 $w=1.68e-07 $l=1.105e-06 $layer=LI1_cond $X=2.335 $Y=2.4
+ $X2=1.23 $Y2=2.4
r132 15 20 28.304 $w=2.03e-07 $l=4.9784e-07 $layer=LI1_cond $X=0.765 $Y=2.332
+ $X2=1.23 $Y2=2.4
r133 15 36 8.41379 $w=2.03e-07 $l=1.4e-07 $layer=LI1_cond $X=0.765 $Y=2.332
+ $X2=0.625 $Y2=2.332
r134 15 17 18.4391 $w=2.48e-07 $l=4e-07 $layer=LI1_cond $X=0.765 $Y=2.35
+ $X2=0.765 $Y2=2.75
r135 14 36 1.77774 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=0.625 $Y=2.18
+ $X2=0.625 $Y2=2.332
r136 13 34 6.36164 $w=1.7e-07 $l=2.2e-07 $layer=LI1_cond $X=0.625 $Y=0.79
+ $X2=0.625 $Y2=0.57
r137 13 14 90.6845 $w=1.68e-07 $l=1.39e-06 $layer=LI1_cond $X=0.625 $Y=0.79
+ $X2=0.625 $Y2=2.18
r138 4 29 600 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_PDIFF $count=1 $X=3.19
+ $Y=2.54 $X2=3.335 $Y2=2.75
r139 3 17 600 $w=1.7e-07 $l=2.74955e-07 $layer=licon1_PDIFF $count=1 $X=0.575
+ $Y=2.54 $X2=0.725 $Y2=2.75
r140 2 42 182 $w=1.7e-07 $l=2.755e-07 $layer=licon1_NDIFF $count=1 $X=3.155
+ $Y=0.635 $X2=3.28 $Y2=0.855
r141 1 32 182 $w=1.7e-07 $l=2.62678e-07 $layer=licon1_NDIFF $count=1 $X=0.165
+ $Y=0.37 $X2=0.31 $Y2=0.57
.ends

.subckt PM_SKY130_FD_SC_HS__DFRTN_1%Q 1 2 9 13 14 15 16 23 32
r26 21 23 1.31708 $w=3.48e-07 $l=4e-08 $layer=LI1_cond $X=10.78 $Y=1.995
+ $X2=10.78 $Y2=2.035
r27 15 16 12.183 $w=3.48e-07 $l=3.7e-07 $layer=LI1_cond $X=10.78 $Y=2.405
+ $X2=10.78 $Y2=2.775
r28 14 21 0.75732 $w=3.48e-07 $l=2.3e-08 $layer=LI1_cond $X=10.78 $Y=1.972
+ $X2=10.78 $Y2=1.995
r29 14 32 8.06043 $w=3.48e-07 $l=1.52e-07 $layer=LI1_cond $X=10.78 $Y=1.972
+ $X2=10.78 $Y2=1.82
r30 14 15 11.4586 $w=3.48e-07 $l=3.48e-07 $layer=LI1_cond $X=10.78 $Y=2.057
+ $X2=10.78 $Y2=2.405
r31 14 23 0.724393 $w=3.48e-07 $l=2.2e-08 $layer=LI1_cond $X=10.78 $Y=2.057
+ $X2=10.78 $Y2=2.035
r32 13 32 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=10.87 $Y=1.15
+ $X2=10.87 $Y2=1.82
r33 7 13 9.06106 $w=3.63e-07 $l=1.82e-07 $layer=LI1_cond $X=10.772 $Y=0.968
+ $X2=10.772 $Y2=1.15
r34 7 9 11.4613 $w=3.63e-07 $l=3.63e-07 $layer=LI1_cond $X=10.772 $Y=0.968
+ $X2=10.772 $Y2=0.605
r35 2 14 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=10.62
+ $Y=1.84 $X2=10.77 $Y2=1.985
r36 2 16 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=10.62
+ $Y=1.84 $X2=10.77 $Y2=2.815
r37 1 9 91 $w=1.7e-07 $l=1.96214e-07 $layer=licon1_NDIFF $count=2 $X=10.615
+ $Y=0.47 $X2=10.755 $Y2=0.605
.ends

.subckt PM_SKY130_FD_SC_HS__DFRTN_1%VGND 1 2 3 4 5 18 22 26 30 34 36 38 43 48 53
+ 61 71 72 75 78 81 84 87
r110 87 88 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.32 $Y=0
+ $X2=10.32 $Y2=0
r111 84 85 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r112 81 82 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r113 78 79 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r114 75 76 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r115 72 88 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.8 $Y=0
+ $X2=10.32 $Y2=0
r116 71 72 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.8 $Y=0 $X2=10.8
+ $Y2=0
r117 69 87 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=10.41 $Y=0
+ $X2=10.285 $Y2=0
r118 69 71 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=10.41 $Y=0 $X2=10.8
+ $Y2=0
r119 68 88 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.84 $Y=0
+ $X2=10.32 $Y2=0
r120 67 68 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=9.84 $Y=0 $X2=9.84
+ $Y2=0
r121 65 68 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=8.88 $Y=0 $X2=9.84
+ $Y2=0
r122 65 85 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=0 $X2=8.4
+ $Y2=0
r123 64 67 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=8.88 $Y=0 $X2=9.84
+ $Y2=0
r124 64 65 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=8.88 $Y=0 $X2=8.88
+ $Y2=0
r125 62 84 10.4332 $w=1.7e-07 $l=2.2e-07 $layer=LI1_cond $X=8.555 $Y=0 $X2=8.335
+ $Y2=0
r126 62 64 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=8.555 $Y=0
+ $X2=8.88 $Y2=0
r127 61 87 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=10.16 $Y=0
+ $X2=10.285 $Y2=0
r128 61 67 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=10.16 $Y=0 $X2=9.84
+ $Y2=0
r129 60 85 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=0 $X2=8.4
+ $Y2=0
r130 59 60 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=7.92 $Y=0 $X2=7.92
+ $Y2=0
r131 56 59 156.578 $w=1.68e-07 $l=2.4e-06 $layer=LI1_cond $X=5.52 $Y=0 $X2=7.92
+ $Y2=0
r132 54 81 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.355 $Y=0 $X2=5.19
+ $Y2=0
r133 54 56 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=5.355 $Y=0
+ $X2=5.52 $Y2=0
r134 53 84 10.4332 $w=1.7e-07 $l=2.2e-07 $layer=LI1_cond $X=8.115 $Y=0 $X2=8.335
+ $Y2=0
r135 53 59 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=8.115 $Y=0
+ $X2=7.92 $Y2=0
r136 52 82 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=2.64 $Y=0 $X2=5.04
+ $Y2=0
r137 52 79 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=2.16
+ $Y2=0
r138 51 52 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r139 49 78 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.35 $Y=0 $X2=2.185
+ $Y2=0
r140 49 51 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=2.35 $Y=0 $X2=2.64
+ $Y2=0
r141 48 81 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.025 $Y=0 $X2=5.19
+ $Y2=0
r142 48 51 155.599 $w=1.68e-07 $l=2.385e-06 $layer=LI1_cond $X=5.025 $Y=0
+ $X2=2.64 $Y2=0
r143 47 79 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r144 47 76 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r145 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r146 44 75 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.295 $Y=0 $X2=1.17
+ $Y2=0
r147 44 46 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=1.295 $Y=0
+ $X2=1.68 $Y2=0
r148 43 78 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.02 $Y=0 $X2=2.185
+ $Y2=0
r149 43 46 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=2.02 $Y=0 $X2=1.68
+ $Y2=0
r150 41 76 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r151 40 41 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r152 38 75 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.045 $Y=0 $X2=1.17
+ $Y2=0
r153 38 40 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=1.045 $Y=0
+ $X2=0.72 $Y2=0
r154 36 60 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=5.52 $Y=0 $X2=7.92
+ $Y2=0
r155 36 82 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=5.04
+ $Y2=0
r156 36 56 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r157 32 87 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=10.285 $Y=0.085
+ $X2=10.285 $Y2=0
r158 32 34 23.9708 $w=2.48e-07 $l=5.2e-07 $layer=LI1_cond $X=10.285 $Y=0.085
+ $X2=10.285 $Y2=0.605
r159 28 84 1.73497 $w=4.4e-07 $l=8.5e-08 $layer=LI1_cond $X=8.335 $Y=0.085
+ $X2=8.335 $Y2=0
r160 28 30 17.1557 $w=4.38e-07 $l=6.55e-07 $layer=LI1_cond $X=8.335 $Y=0.085
+ $X2=8.335 $Y2=0.74
r161 24 81 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.19 $Y=0.085
+ $X2=5.19 $Y2=0
r162 24 26 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=5.19 $Y=0.085
+ $X2=5.19 $Y2=0.535
r163 20 78 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.185 $Y=0.085
+ $X2=2.185 $Y2=0
r164 20 22 7.50834 $w=3.28e-07 $l=2.15e-07 $layer=LI1_cond $X=2.185 $Y=0.085
+ $X2=2.185 $Y2=0.3
r165 16 75 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.17 $Y=0.085
+ $X2=1.17 $Y2=0
r166 16 18 22.8184 $w=2.48e-07 $l=4.95e-07 $layer=LI1_cond $X=1.17 $Y=0.085
+ $X2=1.17 $Y2=0.58
r167 5 34 91 $w=1.7e-07 $l=2.79464e-07 $layer=licon1_NDIFF $count=2 $X=10.105
+ $Y=0.47 $X2=10.325 $Y2=0.605
r168 4 30 182 $w=1.7e-07 $l=2.57488e-07 $layer=licon1_NDIFF $count=1 $X=8.14
+ $Y=0.595 $X2=8.335 $Y2=0.74
r169 3 26 182 $w=1.7e-07 $l=2.6533e-07 $layer=licon1_NDIFF $count=1 $X=4.97
+ $Y=0.635 $X2=5.19 $Y2=0.535
r170 2 22 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=2.045
+ $Y=0.155 $X2=2.185 $Y2=0.3
r171 1 18 182 $w=1.7e-07 $l=3.07571e-07 $layer=licon1_NDIFF $count=1 $X=0.99
+ $Y=0.37 $X2=1.21 $Y2=0.58
.ends

