* NGSPICE file created from sky130_fd_sc_hs__a221o_4.ext - technology: sky130A

.subckt sky130_fd_sc_hs__a221o_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
M1000 VPWR a_154_135# X VPB pshort w=1.12e+06u l=150000u
+  ad=2.157e+12p pd=1.483e+07u as=6.72e+11p ps=5.68e+06u
M1001 a_157_376# A1 VPWR VPB pshort w=1e+06u l=150000u
+  ad=1.36e+12p pd=1.072e+07u as=0p ps=0u
M1002 X a_154_135# VGND VNB nlowvt w=740000u l=150000u
+  ad=4.144e+11p pd=4.08e+06u as=1.62282e+12p ps=1.315e+07u
M1003 a_154_135# C1 a_1102_392# VPB pshort w=1e+06u l=150000u
+  ad=3e+11p pd=2.6e+06u as=1.44e+12p ps=1.088e+07u
M1004 VPWR A1 a_157_376# VPB pshort w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_154_135# A1 a_71_135# VNB nlowvt w=640000u l=150000u
+  ad=5.376e+11p pd=5.52e+06u as=5.184e+11p ps=5.46e+06u
M1006 a_1102_392# C1 a_154_135# VPB pshort w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_71_135# A1 a_154_135# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_157_376# B2 a_1102_392# VPB pshort w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_1102_392# B2 a_157_376# VPB pshort w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_157_376# B1 a_1102_392# VPB pshort w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_154_135# B1 a_1346_123# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=5.632e+11p ps=5.6e+06u
M1012 VGND a_154_135# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_157_376# A2 VPWR VPB pshort w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_1346_123# B2 VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VPWR A2 a_157_376# VPB pshort w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VGND B2 a_1346_123# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 X a_154_135# VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_1346_123# B1 a_154_135# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VPWR a_154_135# X VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 VGND a_154_135# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_1102_392# B1 a_157_376# VPB pshort w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_71_135# A2 VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 X a_154_135# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 a_154_135# C1 VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 X a_154_135# VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 VGND C1 a_154_135# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 VGND A2 a_71_135# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

