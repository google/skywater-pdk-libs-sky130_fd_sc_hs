* NGSPICE file created from sky130_fd_sc_hs__a21bo_2.ext - technology: sky130A

.subckt sky130_fd_sc_hs__a21bo_2 A1 A2 B1_N VGND VNB VPB VPWR X
M1000 VGND a_187_244# X VNB nlowvt w=740000u l=150000u
+  ad=9.689e+11p pd=7.11e+06u as=2.072e+11p ps=2.04e+06u
M1001 a_187_244# a_32_368# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.072e+11p pd=2.04e+06u as=0p ps=0u
M1002 VPWR B1_N a_32_368# VPB pshort w=840000u l=150000u
+  ad=9.916e+11p pd=8.36e+06u as=2.31e+11p ps=2.23e+06u
M1003 X a_187_244# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 VGND A2 a_587_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.368e+11p ps=2.12e+06u
M1005 a_504_392# a_32_368# a_187_244# VPB pshort w=1e+06u l=150000u
+  ad=5.75e+11p pd=5.15e+06u as=2.75e+11p ps=2.55e+06u
M1006 VPWR A1 a_504_392# VPB pshort w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 X a_187_244# VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=3.36e+11p pd=2.84e+06u as=0p ps=0u
M1008 a_504_392# A2 VPWR VPB pshort w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VGND B1_N a_32_368# VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=1.4575e+11p ps=1.63e+06u
M1010 a_587_74# A1 a_187_244# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VPWR a_187_244# X VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

