* File: sky130_fd_sc_hs__o22ai_4.pex.spice
* Created: Thu Aug 27 21:00:43 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HS__O22AI_4%A1 3 5 7 8 10 13 17 19 21 22 24 27 29 36 45
+ 48 49 58 62 66
c126 29 0 8.50911e-20 $X=1.38 $Y=1.485
c127 22 0 2.61514e-19 $X=3.76 $Y=1.765
c128 17 0 3.15663e-20 $X=1.425 $Y=0.74
c129 13 0 7.73112e-20 $X=0.995 $Y=0.74
c130 8 0 8.10185e-20 $X=0.96 $Y=1.765
c131 5 0 1.60269e-20 $X=0.51 $Y=1.765
r132 58 59 4.39323 $w=3.84e-07 $l=3.5e-08 $layer=POLY_cond $X=1.425 $Y=1.542
+ $X2=1.46 $Y2=1.542
r133 55 56 4.39323 $w=3.84e-07 $l=3.5e-08 $layer=POLY_cond $X=0.96 $Y=1.542
+ $X2=0.995 $Y2=1.542
r134 52 53 1.88281 $w=3.84e-07 $l=1.5e-08 $layer=POLY_cond $X=0.495 $Y=1.542
+ $X2=0.51 $Y2=1.542
r135 49 66 7.44484 $w=4.28e-07 $l=1.15e-07 $layer=LI1_cond $X=3.12 $Y=1.935
+ $X2=3.235 $Y2=1.935
r136 48 49 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=2.64 $Y=1.935
+ $X2=3.12 $Y2=1.935
r137 48 62 7.44484 $w=4.28e-07 $l=1.15e-07 $layer=LI1_cond $X=2.64 $Y=1.935
+ $X2=2.525 $Y2=1.935
r138 45 47 13.2509 $w=2.67e-07 $l=2.9e-07 $layer=LI1_cond $X=3.805 $Y=1.515
+ $X2=3.805 $Y2=1.805
r139 45 46 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.805
+ $Y=1.515 $X2=3.805 $Y2=1.515
r140 41 58 5.02083 $w=3.84e-07 $l=4e-08 $layer=POLY_cond $X=1.385 $Y=1.542
+ $X2=1.425 $Y2=1.542
r141 41 56 48.9531 $w=3.84e-07 $l=3.9e-07 $layer=POLY_cond $X=1.385 $Y=1.542
+ $X2=0.995 $Y2=1.542
r142 36 47 3.37873 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.64 $Y=1.805
+ $X2=3.805 $Y2=1.805
r143 36 66 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=3.64 $Y=1.805
+ $X2=3.235 $Y2=1.805
r144 35 42 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.55 $Y=1.805
+ $X2=1.465 $Y2=1.805
r145 35 62 63.6096 $w=1.68e-07 $l=9.75e-07 $layer=LI1_cond $X=1.55 $Y=1.805
+ $X2=2.525 $Y2=1.805
r146 32 55 32.0078 $w=3.84e-07 $l=2.55e-07 $layer=POLY_cond $X=0.705 $Y=1.542
+ $X2=0.96 $Y2=1.542
r147 32 53 24.4766 $w=3.84e-07 $l=1.95e-07 $layer=POLY_cond $X=0.705 $Y=1.542
+ $X2=0.51 $Y2=1.542
r148 31 32 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=0.705
+ $Y=1.485 $X2=0.705 $Y2=1.485
r149 29 42 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=1.465 $Y=1.485
+ $X2=1.465 $Y2=1.805
r150 29 41 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.385
+ $Y=1.485 $X2=1.385 $Y2=1.485
r151 29 31 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=1.38 $Y=1.485
+ $X2=0.705 $Y2=1.485
r152 25 46 38.5562 $w=2.99e-07 $l=1.88348e-07 $layer=POLY_cond $X=3.855 $Y=1.35
+ $X2=3.805 $Y2=1.515
r153 25 27 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=3.855 $Y=1.35
+ $X2=3.855 $Y2=0.74
r154 22 46 52.2586 $w=2.99e-07 $l=2.7157e-07 $layer=POLY_cond $X=3.76 $Y=1.765
+ $X2=3.805 $Y2=1.515
r155 22 24 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.76 $Y=1.765
+ $X2=3.76 $Y2=2.4
r156 19 59 24.8669 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=1.46 $Y=1.765
+ $X2=1.46 $Y2=1.542
r157 19 21 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.46 $Y=1.765
+ $X2=1.46 $Y2=2.4
r158 15 58 24.8669 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=1.425 $Y=1.32
+ $X2=1.425 $Y2=1.542
r159 15 17 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=1.425 $Y=1.32
+ $X2=1.425 $Y2=0.74
r160 11 56 24.8669 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=0.995 $Y=1.32
+ $X2=0.995 $Y2=1.542
r161 11 13 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=0.995 $Y=1.32
+ $X2=0.995 $Y2=0.74
r162 8 55 24.8669 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=0.96 $Y=1.765
+ $X2=0.96 $Y2=1.542
r163 8 10 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.96 $Y=1.765
+ $X2=0.96 $Y2=2.4
r164 5 53 24.8669 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=0.51 $Y=1.765
+ $X2=0.51 $Y2=1.542
r165 5 7 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.51 $Y=1.765
+ $X2=0.51 $Y2=2.4
r166 1 52 24.8669 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=0.495 $Y=1.32
+ $X2=0.495 $Y2=1.542
r167 1 3 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=0.495 $Y=1.32
+ $X2=0.495 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HS__O22AI_4%A2 1 3 4 6 7 9 10 12 13 15 16 18 19 21 22 24
+ 25 26 27 46
c88 27 0 1.98342e-19 $X=3.12 $Y=1.295
c89 10 0 4.72982e-20 $X=2.41 $Y=1.765
c90 1 0 8.50911e-20 $X=1.91 $Y=1.765
r91 46 47 1.71734 $w=4.21e-07 $l=1.5e-08 $layer=POLY_cond $X=3.31 $Y=1.492
+ $X2=3.325 $Y2=1.492
r92 44 46 27.4774 $w=4.21e-07 $l=2.4e-07 $layer=POLY_cond $X=3.07 $Y=1.492
+ $X2=3.31 $Y2=1.492
r93 44 45 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.07
+ $Y=1.385 $X2=3.07 $Y2=1.385
r94 42 44 24.0428 $w=4.21e-07 $l=2.1e-07 $layer=POLY_cond $X=2.86 $Y=1.492
+ $X2=3.07 $Y2=1.492
r95 41 42 0.572447 $w=4.21e-07 $l=5e-09 $layer=POLY_cond $X=2.855 $Y=1.492
+ $X2=2.86 $Y2=1.492
r96 40 45 10.59 $w=3.68e-07 $l=3.4e-07 $layer=LI1_cond $X=2.73 $Y=1.365 $X2=3.07
+ $Y2=1.365
r97 39 41 14.3112 $w=4.21e-07 $l=1.25e-07 $layer=POLY_cond $X=2.73 $Y=1.492
+ $X2=2.855 $Y2=1.492
r98 39 40 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.73
+ $Y=1.385 $X2=2.73 $Y2=1.385
r99 37 39 36.6366 $w=4.21e-07 $l=3.2e-07 $layer=POLY_cond $X=2.41 $Y=1.492
+ $X2=2.73 $Y2=1.492
r100 36 37 6.29691 $w=4.21e-07 $l=5.5e-08 $layer=POLY_cond $X=2.355 $Y=1.492
+ $X2=2.41 $Y2=1.492
r101 34 36 34.9192 $w=4.21e-07 $l=3.05e-07 $layer=POLY_cond $X=2.05 $Y=1.492
+ $X2=2.355 $Y2=1.492
r102 34 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.05
+ $Y=1.385 $X2=2.05 $Y2=1.385
r103 32 34 14.3112 $w=4.21e-07 $l=1.25e-07 $layer=POLY_cond $X=1.925 $Y=1.492
+ $X2=2.05 $Y2=1.492
r104 31 32 1.71734 $w=4.21e-07 $l=1.5e-08 $layer=POLY_cond $X=1.91 $Y=1.492
+ $X2=1.925 $Y2=1.492
r105 27 45 1.55736 $w=3.68e-07 $l=5e-08 $layer=LI1_cond $X=3.12 $Y=1.365
+ $X2=3.07 $Y2=1.365
r106 26 40 2.80324 $w=3.68e-07 $l=9e-08 $layer=LI1_cond $X=2.64 $Y=1.365
+ $X2=2.73 $Y2=1.365
r107 25 26 14.9506 $w=3.68e-07 $l=4.8e-07 $layer=LI1_cond $X=2.16 $Y=1.365
+ $X2=2.64 $Y2=1.365
r108 25 35 3.42618 $w=3.68e-07 $l=1.1e-07 $layer=LI1_cond $X=2.16 $Y=1.365
+ $X2=2.05 $Y2=1.365
r109 22 47 27.1176 $w=1.5e-07 $l=2.72e-07 $layer=POLY_cond $X=3.325 $Y=1.22
+ $X2=3.325 $Y2=1.492
r110 22 24 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=3.325 $Y=1.22
+ $X2=3.325 $Y2=0.74
r111 19 46 27.1176 $w=1.5e-07 $l=2.73e-07 $layer=POLY_cond $X=3.31 $Y=1.765
+ $X2=3.31 $Y2=1.492
r112 19 21 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.31 $Y=1.765
+ $X2=3.31 $Y2=2.4
r113 16 42 27.1176 $w=1.5e-07 $l=2.73e-07 $layer=POLY_cond $X=2.86 $Y=1.765
+ $X2=2.86 $Y2=1.492
r114 16 18 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.86 $Y=1.765
+ $X2=2.86 $Y2=2.4
r115 13 41 27.1176 $w=1.5e-07 $l=2.72e-07 $layer=POLY_cond $X=2.855 $Y=1.22
+ $X2=2.855 $Y2=1.492
r116 13 15 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=2.855 $Y=1.22
+ $X2=2.855 $Y2=0.74
r117 10 37 27.1176 $w=1.5e-07 $l=2.73e-07 $layer=POLY_cond $X=2.41 $Y=1.765
+ $X2=2.41 $Y2=1.492
r118 10 12 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.41 $Y=1.765
+ $X2=2.41 $Y2=2.4
r119 7 36 27.1176 $w=1.5e-07 $l=2.72e-07 $layer=POLY_cond $X=2.355 $Y=1.22
+ $X2=2.355 $Y2=1.492
r120 7 9 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=2.355 $Y=1.22
+ $X2=2.355 $Y2=0.74
r121 4 32 27.1176 $w=1.5e-07 $l=2.72e-07 $layer=POLY_cond $X=1.925 $Y=1.22
+ $X2=1.925 $Y2=1.492
r122 4 6 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.925 $Y=1.22
+ $X2=1.925 $Y2=0.74
r123 1 31 27.1176 $w=1.5e-07 $l=2.73e-07 $layer=POLY_cond $X=1.91 $Y=1.765
+ $X2=1.91 $Y2=1.492
r124 1 3 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.91 $Y=1.765
+ $X2=1.91 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_HS__O22AI_4%B1 3 5 7 8 10 13 15 17 20 22 24 25 27 28 36
+ 38 44 52 55
c121 13 0 7.5396e-20 $X=4.785 $Y=0.74
r122 52 53 1.82116 $w=3.97e-07 $l=1.5e-08 $layer=POLY_cond $X=5.21 $Y=1.532
+ $X2=5.225 $Y2=1.532
r123 49 50 3.03526 $w=3.97e-07 $l=2.5e-08 $layer=POLY_cond $X=4.76 $Y=1.532
+ $X2=4.785 $Y2=1.532
r124 46 47 1.82116 $w=3.97e-07 $l=1.5e-08 $layer=POLY_cond $X=4.295 $Y=1.532
+ $X2=4.31 $Y2=1.532
r125 44 55 6.01275 $w=2.28e-07 $l=1.2e-07 $layer=LI1_cond $X=5.52 $Y=1.295
+ $X2=5.52 $Y2=1.175
r126 41 42 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.565
+ $Y=1.385 $X2=7.565 $Y2=1.385
r127 38 41 7.33373 $w=3.28e-07 $l=2.1e-07 $layer=LI1_cond $X=7.565 $Y=1.175
+ $X2=7.565 $Y2=1.385
r128 37 55 2.50919 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=5.635 $Y=1.175
+ $X2=5.52 $Y2=1.175
r129 36 38 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.4 $Y=1.175
+ $X2=7.565 $Y2=1.175
r130 36 37 115.15 $w=1.68e-07 $l=1.765e-06 $layer=LI1_cond $X=7.4 $Y=1.175
+ $X2=5.635 $Y2=1.175
r131 35 52 9.10579 $w=3.97e-07 $l=7.5e-08 $layer=POLY_cond $X=5.135 $Y=1.532
+ $X2=5.21 $Y2=1.532
r132 35 50 42.4937 $w=3.97e-07 $l=3.5e-07 $layer=POLY_cond $X=5.135 $Y=1.532
+ $X2=4.785 $Y2=1.532
r133 34 35 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=5.135
+ $Y=1.465 $X2=5.135 $Y2=1.465
r134 31 49 37.0302 $w=3.97e-07 $l=3.05e-07 $layer=POLY_cond $X=4.455 $Y=1.532
+ $X2=4.76 $Y2=1.532
r135 31 47 17.6045 $w=3.97e-07 $l=1.45e-07 $layer=POLY_cond $X=4.455 $Y=1.532
+ $X2=4.31 $Y2=1.532
r136 30 34 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=4.455 $Y=1.465
+ $X2=5.135 $Y2=1.465
r137 30 31 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=4.455
+ $Y=1.465 $X2=4.455 $Y2=1.465
r138 28 44 8.51806 $w=2.28e-07 $l=1.7e-07 $layer=LI1_cond $X=5.52 $Y=1.465
+ $X2=5.52 $Y2=1.295
r139 28 34 9.42908 $w=3.28e-07 $l=2.7e-07 $layer=LI1_cond $X=5.405 $Y=1.465
+ $X2=5.135 $Y2=1.465
r140 25 42 38.9026 $w=2.7e-07 $l=1.74714e-07 $layer=POLY_cond $X=7.585 $Y=1.22
+ $X2=7.565 $Y2=1.385
r141 25 27 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=7.585 $Y=1.22
+ $X2=7.585 $Y2=0.74
r142 22 42 77.2841 $w=2.7e-07 $l=3.82492e-07 $layer=POLY_cond $X=7.56 $Y=1.765
+ $X2=7.565 $Y2=1.385
r143 22 24 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=7.56 $Y=1.765
+ $X2=7.56 $Y2=2.4
r144 18 53 25.678 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=5.225 $Y=1.3
+ $X2=5.225 $Y2=1.532
r145 18 20 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=5.225 $Y=1.3
+ $X2=5.225 $Y2=0.74
r146 15 52 25.678 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=5.21 $Y=1.765
+ $X2=5.21 $Y2=1.532
r147 15 17 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=5.21 $Y=1.765
+ $X2=5.21 $Y2=2.4
r148 11 50 25.678 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=4.785 $Y=1.3
+ $X2=4.785 $Y2=1.532
r149 11 13 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=4.785 $Y=1.3
+ $X2=4.785 $Y2=0.74
r150 8 49 25.678 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=4.76 $Y=1.765
+ $X2=4.76 $Y2=1.532
r151 8 10 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=4.76 $Y=1.765
+ $X2=4.76 $Y2=2.4
r152 5 47 25.678 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=4.31 $Y=1.765
+ $X2=4.31 $Y2=1.532
r153 5 7 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=4.31 $Y=1.765
+ $X2=4.31 $Y2=2.4
r154 1 46 25.678 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=4.295 $Y=1.3
+ $X2=4.295 $Y2=1.532
r155 1 3 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=4.295 $Y=1.3
+ $X2=4.295 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HS__O22AI_4%B2 3 5 7 10 12 14 17 19 21 22 24 27 34 35 47
+ 48 50 56
c87 22 0 6.40318e-20 $X=7.07 $Y=1.765
c88 5 0 1.73237e-19 $X=5.71 $Y=1.765
r89 48 49 1.96467 $w=3.68e-07 $l=1.5e-08 $layer=POLY_cond $X=7.07 $Y=1.557
+ $X2=7.085 $Y2=1.557
r90 46 48 10.4783 $w=3.68e-07 $l=8e-08 $layer=POLY_cond $X=6.99 $Y=1.557
+ $X2=7.07 $Y2=1.557
r91 46 47 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.99
+ $Y=1.515 $X2=6.99 $Y2=1.515
r92 44 46 49.7717 $w=3.68e-07 $l=3.8e-07 $layer=POLY_cond $X=6.61 $Y=1.557
+ $X2=6.99 $Y2=1.557
r93 43 44 3.27446 $w=3.68e-07 $l=2.5e-08 $layer=POLY_cond $X=6.585 $Y=1.557
+ $X2=6.61 $Y2=1.557
r94 40 41 9.82337 $w=3.68e-07 $l=7.5e-08 $layer=POLY_cond $X=6.085 $Y=1.557
+ $X2=6.16 $Y2=1.557
r95 39 40 49.1168 $w=3.68e-07 $l=3.75e-07 $layer=POLY_cond $X=5.71 $Y=1.557
+ $X2=6.085 $Y2=1.557
r96 38 39 7.2038 $w=3.68e-07 $l=5.5e-08 $layer=POLY_cond $X=5.655 $Y=1.557
+ $X2=5.71 $Y2=1.557
r97 35 47 0.987808 $w=3.48e-07 $l=3e-08 $layer=LI1_cond $X=6.96 $Y=1.605
+ $X2=6.99 $Y2=1.605
r98 35 50 8.0671 $w=3.48e-07 $l=2.45e-07 $layer=LI1_cond $X=6.96 $Y=1.605
+ $X2=6.715 $Y2=1.605
r99 34 50 7.73783 $w=3.48e-07 $l=2.35e-07 $layer=LI1_cond $X=6.48 $Y=1.605
+ $X2=6.715 $Y2=1.605
r100 34 56 4.74445 $w=3.48e-07 $l=1.15e-07 $layer=LI1_cond $X=6.48 $Y=1.605
+ $X2=6.365 $Y2=1.605
r101 32 43 36.019 $w=3.68e-07 $l=2.75e-07 $layer=POLY_cond $X=6.31 $Y=1.557
+ $X2=6.585 $Y2=1.557
r102 32 41 19.6467 $w=3.68e-07 $l=1.5e-07 $layer=POLY_cond $X=6.31 $Y=1.557
+ $X2=6.16 $Y2=1.557
r103 31 56 2.53537 $w=2.48e-07 $l=5.5e-08 $layer=LI1_cond $X=6.31 $Y=1.555
+ $X2=6.365 $Y2=1.555
r104 31 32 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.31
+ $Y=1.515 $X2=6.31 $Y2=1.515
r105 25 49 23.8357 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=7.085 $Y=1.35
+ $X2=7.085 $Y2=1.557
r106 25 27 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=7.085 $Y=1.35
+ $X2=7.085 $Y2=0.74
r107 22 48 23.8357 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=7.07 $Y=1.765
+ $X2=7.07 $Y2=1.557
r108 22 24 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=7.07 $Y=1.765
+ $X2=7.07 $Y2=2.4
r109 19 44 23.8357 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=6.61 $Y=1.765
+ $X2=6.61 $Y2=1.557
r110 19 21 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=6.61 $Y=1.765
+ $X2=6.61 $Y2=2.4
r111 15 43 23.8357 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=6.585 $Y=1.35
+ $X2=6.585 $Y2=1.557
r112 15 17 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=6.585 $Y=1.35
+ $X2=6.585 $Y2=0.74
r113 12 41 23.8357 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=6.16 $Y=1.765
+ $X2=6.16 $Y2=1.557
r114 12 14 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=6.16 $Y=1.765
+ $X2=6.16 $Y2=2.4
r115 8 40 23.8357 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=6.085 $Y=1.35
+ $X2=6.085 $Y2=1.557
r116 8 10 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=6.085 $Y=1.35
+ $X2=6.085 $Y2=0.74
r117 5 39 23.8357 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=5.71 $Y=1.765
+ $X2=5.71 $Y2=1.557
r118 5 7 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=5.71 $Y=1.765
+ $X2=5.71 $Y2=2.4
r119 1 38 23.8357 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=5.655 $Y=1.35
+ $X2=5.655 $Y2=1.557
r120 1 3 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=5.655 $Y=1.35
+ $X2=5.655 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HS__O22AI_4%VPWR 1 2 3 4 5 16 18 24 28 32 34 36 38 40 45
+ 53 58 70 73 76 80
c97 32 0 1.73237e-19 $X=4.985 $Y=2.755
r98 79 80 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r99 76 77 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r100 70 71 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r101 67 68 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r102 65 80 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=7.92 $Y2=3.33
r103 64 65 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r104 62 65 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=7.44 $Y2=3.33
r105 62 77 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=5.04 $Y2=3.33
r106 61 64 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=5.52 $Y=3.33
+ $X2=7.44 $Y2=3.33
r107 61 62 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r108 59 76 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.15 $Y=3.33
+ $X2=5.025 $Y2=3.33
r109 59 61 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=5.15 $Y=3.33
+ $X2=5.52 $Y2=3.33
r110 58 79 4.64076 $w=1.7e-07 $l=2.45e-07 $layer=LI1_cond $X=7.67 $Y=3.33
+ $X2=7.915 $Y2=3.33
r111 58 64 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=7.67 $Y=3.33
+ $X2=7.44 $Y2=3.33
r112 57 77 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=5.04 $Y2=3.33
r113 56 57 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r114 54 73 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.2 $Y=3.33
+ $X2=4.035 $Y2=3.33
r115 54 56 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=4.2 $Y=3.33
+ $X2=4.56 $Y2=3.33
r116 53 76 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.9 $Y=3.33
+ $X2=5.025 $Y2=3.33
r117 53 56 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=4.9 $Y=3.33
+ $X2=4.56 $Y2=3.33
r118 51 52 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r119 49 52 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=3.6 $Y2=3.33
r120 49 71 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r121 48 51 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=1.68 $Y=3.33
+ $X2=3.6 $Y2=3.33
r122 48 49 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r123 46 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.35 $Y=3.33
+ $X2=1.185 $Y2=3.33
r124 46 48 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=1.35 $Y=3.33
+ $X2=1.68 $Y2=3.33
r125 45 73 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.87 $Y=3.33
+ $X2=4.035 $Y2=3.33
r126 45 51 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=3.87 $Y=3.33 $X2=3.6
+ $Y2=3.33
r127 44 71 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r128 44 68 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r129 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r130 41 67 4.0045 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=0.37 $Y=3.33
+ $X2=0.185 $Y2=3.33
r131 41 43 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=0.37 $Y=3.33
+ $X2=0.72 $Y2=3.33
r132 40 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.02 $Y=3.33
+ $X2=1.185 $Y2=3.33
r133 40 43 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=1.02 $Y=3.33 $X2=0.72
+ $Y2=3.33
r134 38 57 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=4.56 $Y2=3.33
r135 38 52 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=3.6 $Y2=3.33
r136 38 73 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r137 34 79 3.12541 $w=3.3e-07 $l=1.18427e-07 $layer=LI1_cond $X=7.835 $Y=3.245
+ $X2=7.915 $Y2=3.33
r138 34 36 27.5888 $w=3.28e-07 $l=7.9e-07 $layer=LI1_cond $X=7.835 $Y=3.245
+ $X2=7.835 $Y2=2.455
r139 30 76 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.025 $Y=3.245
+ $X2=5.025 $Y2=3.33
r140 30 32 22.5879 $w=2.48e-07 $l=4.9e-07 $layer=LI1_cond $X=5.025 $Y=3.245
+ $X2=5.025 $Y2=2.755
r141 26 73 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.035 $Y=3.245
+ $X2=4.035 $Y2=3.33
r142 26 28 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=4.035 $Y=3.245
+ $X2=4.035 $Y2=2.78
r143 22 70 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.185 $Y=3.245
+ $X2=1.185 $Y2=3.33
r144 22 24 26.5411 $w=3.28e-07 $l=7.6e-07 $layer=LI1_cond $X=1.185 $Y=3.245
+ $X2=1.185 $Y2=2.485
r145 18 21 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=0.245 $Y=1.985
+ $X2=0.245 $Y2=2.815
r146 16 67 3.13866 $w=2.5e-07 $l=1.11018e-07 $layer=LI1_cond $X=0.245 $Y=3.245
+ $X2=0.185 $Y2=3.33
r147 16 21 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=0.245 $Y=3.245
+ $X2=0.245 $Y2=2.815
r148 5 36 300 $w=1.7e-07 $l=7.07972e-07 $layer=licon1_PDIFF $count=2 $X=7.635
+ $Y=1.84 $X2=7.835 $Y2=2.455
r149 4 32 600 $w=1.7e-07 $l=9.87155e-07 $layer=licon1_PDIFF $count=1 $X=4.835
+ $Y=1.84 $X2=4.985 $Y2=2.755
r150 3 28 600 $w=1.7e-07 $l=1.03518e-06 $layer=licon1_PDIFF $count=1 $X=3.835
+ $Y=1.84 $X2=4.035 $Y2=2.78
r151 2 24 300 $w=1.7e-07 $l=7.16083e-07 $layer=licon1_PDIFF $count=2 $X=1.035
+ $Y=1.84 $X2=1.185 $Y2=2.485
r152 1 21 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=0.14
+ $Y=1.84 $X2=0.285 $Y2=2.815
r153 1 18 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.14
+ $Y=1.84 $X2=0.285 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HS__O22AI_4%A_117_368# 1 2 3 4 15 17 19 20 21 25 28
c51 21 0 8.10185e-20 $X=1.85 $Y=2.82
c52 19 0 4.72982e-20 $X=1.685 $Y=2.23
c53 17 0 1.60269e-20 $X=1.52 $Y=2.145
r54 30 31 3.26614 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=0.735 $Y=2.145
+ $X2=0.735 $Y2=2.23
r55 28 30 5.5876 $w=3.28e-07 $l=1.6e-07 $layer=LI1_cond $X=0.735 $Y=1.985
+ $X2=0.735 $Y2=2.145
r56 23 25 32.4125 $w=3.18e-07 $l=9e-07 $layer=LI1_cond $X=2.635 $Y=2.82
+ $X2=3.535 $Y2=2.82
r57 21 23 28.2709 $w=3.18e-07 $l=7.85e-07 $layer=LI1_cond $X=1.85 $Y=2.82
+ $X2=2.635 $Y2=2.82
r58 20 21 6.81859 $w=3.2e-07 $l=2.31571e-07 $layer=LI1_cond $X=1.685 $Y=2.66
+ $X2=1.85 $Y2=2.82
r59 19 33 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.685 $Y=2.23
+ $X2=1.685 $Y2=2.145
r60 19 20 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=1.685 $Y=2.23
+ $X2=1.685 $Y2=2.66
r61 18 30 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.9 $Y=2.145
+ $X2=0.735 $Y2=2.145
r62 17 33 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.52 $Y=2.145
+ $X2=1.685 $Y2=2.145
r63 17 18 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=1.52 $Y=2.145
+ $X2=0.9 $Y2=2.145
r64 15 31 6.99698 $w=2.78e-07 $l=1.7e-07 $layer=LI1_cond $X=0.71 $Y=2.4 $X2=0.71
+ $Y2=2.23
r65 4 25 600 $w=1.7e-07 $l=1.01223e-06 $layer=licon1_PDIFF $count=1 $X=3.385
+ $Y=1.84 $X2=3.535 $Y2=2.78
r66 3 23 600 $w=1.7e-07 $l=1.01223e-06 $layer=licon1_PDIFF $count=1 $X=2.485
+ $Y=1.84 $X2=2.635 $Y2=2.78
r67 2 33 300 $w=1.7e-07 $l=4.53845e-07 $layer=licon1_PDIFF $count=2 $X=1.535
+ $Y=1.84 $X2=1.685 $Y2=2.225
r68 1 28 600 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=1.84 $X2=0.735 $Y2=1.985
r69 1 15 300 $w=1.7e-07 $l=6.30555e-07 $layer=licon1_PDIFF $count=2 $X=0.585
+ $Y=1.84 $X2=0.735 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_HS__O22AI_4%Y 1 2 3 4 5 6 7 8 25 30 31 32 39 45 47 50 52
+ 57 60 61 63 66 67 68 69 73 80 82
c142 63 0 6.40318e-20 $X=6.835 $Y=2.115
r143 73 80 2.27456 $w=3.78e-07 $l=7.5e-08 $layer=LI1_cond $X=4.965 $Y=0.94
+ $X2=5.04 $Y2=0.94
r144 69 82 6.90319 $w=3.78e-07 $l=1.1e-07 $layer=LI1_cond $X=5.045 $Y=0.94
+ $X2=5.155 $Y2=0.94
r145 69 80 0.151637 $w=3.78e-07 $l=5e-09 $layer=LI1_cond $X=5.045 $Y=0.94
+ $X2=5.04 $Y2=0.94
r146 69 73 0.151637 $w=3.78e-07 $l=5e-09 $layer=LI1_cond $X=4.96 $Y=0.94
+ $X2=4.965 $Y2=0.94
r147 68 69 12.131 $w=3.78e-07 $l=4e-07 $layer=LI1_cond $X=4.56 $Y=0.94 $X2=4.96
+ $Y2=0.94
r148 65 67 8.46017 $w=3.23e-07 $l=1.65e-07 $layer=LI1_cond $X=7.37 $Y=0.757
+ $X2=7.535 $Y2=0.757
r149 65 66 8.46017 $w=3.23e-07 $l=1.65e-07 $layer=LI1_cond $X=7.37 $Y=0.757
+ $X2=7.205 $Y2=0.757
r150 61 66 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=6.535 $Y=0.835
+ $X2=7.205 $Y2=0.835
r151 59 61 8.46017 $w=3.23e-07 $l=1.65e-07 $layer=LI1_cond $X=6.37 $Y=0.757
+ $X2=6.535 $Y2=0.757
r152 59 60 8.46017 $w=3.23e-07 $l=1.65e-07 $layer=LI1_cond $X=6.37 $Y=0.757
+ $X2=6.205 $Y2=0.757
r153 52 54 4.53993 $w=3.28e-07 $l=1.3e-07 $layer=LI1_cond $X=2.185 $Y=2.275
+ $X2=2.185 $Y2=2.405
r154 49 50 67.1979 $w=1.68e-07 $l=1.03e-06 $layer=LI1_cond $X=7.985 $Y=0.92
+ $X2=7.985 $Y2=1.95
r155 47 49 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.9 $Y=0.835
+ $X2=7.985 $Y2=0.92
r156 47 67 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=7.9 $Y=0.835
+ $X2=7.535 $Y2=0.835
r157 46 63 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7 $Y=2.035
+ $X2=6.835 $Y2=2.035
r158 45 50 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.9 $Y=2.035
+ $X2=7.985 $Y2=1.95
r159 45 46 58.7166 $w=1.68e-07 $l=9e-07 $layer=LI1_cond $X=7.9 $Y=2.035 $X2=7
+ $Y2=2.035
r160 40 57 8.61065 $w=1.7e-07 $l=1.88348e-07 $layer=LI1_cond $X=6.1 $Y=2.035
+ $X2=5.935 $Y2=1.985
r161 39 63 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.67 $Y=2.035
+ $X2=6.835 $Y2=2.035
r162 39 40 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=6.67 $Y=2.035
+ $X2=6.1 $Y2=2.035
r163 36 60 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=5.44 $Y=0.835
+ $X2=6.205 $Y2=0.835
r164 36 82 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=5.44 $Y=0.835
+ $X2=5.155 $Y2=0.835
r165 31 57 8.61065 $w=1.7e-07 $l=1.88348e-07 $layer=LI1_cond $X=5.77 $Y=1.935
+ $X2=5.935 $Y2=1.985
r166 31 32 105.69 $w=1.68e-07 $l=1.62e-06 $layer=LI1_cond $X=5.77 $Y=1.935
+ $X2=4.15 $Y2=1.935
r167 29 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.065 $Y=2.02
+ $X2=4.15 $Y2=1.935
r168 29 30 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=4.065 $Y=2.02
+ $X2=4.065 $Y2=2.32
r169 26 54 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.35 $Y=2.405
+ $X2=2.185 $Y2=2.405
r170 26 28 47.9519 $w=1.68e-07 $l=7.35e-07 $layer=LI1_cond $X=2.35 $Y=2.405
+ $X2=3.085 $Y2=2.405
r171 25 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.98 $Y=2.405
+ $X2=4.065 $Y2=2.32
r172 25 28 58.3904 $w=1.68e-07 $l=8.95e-07 $layer=LI1_cond $X=3.98 $Y=2.405
+ $X2=3.085 $Y2=2.405
r173 8 63 300 $w=1.7e-07 $l=3.4187e-07 $layer=licon1_PDIFF $count=2 $X=6.685
+ $Y=1.84 $X2=6.835 $Y2=2.115
r174 7 57 300 $w=1.7e-07 $l=2.38485e-07 $layer=licon1_PDIFF $count=2 $X=5.785
+ $Y=1.84 $X2=5.935 $Y2=2.015
r175 6 28 600 $w=1.7e-07 $l=6.3559e-07 $layer=licon1_PDIFF $count=1 $X=2.935
+ $Y=1.84 $X2=3.085 $Y2=2.405
r176 5 52 600 $w=1.7e-07 $l=5.25571e-07 $layer=licon1_PDIFF $count=1 $X=1.985
+ $Y=1.84 $X2=2.185 $Y2=2.275
r177 4 65 182 $w=1.7e-07 $l=4.37579e-07 $layer=licon1_NDIFF $count=1 $X=7.16
+ $Y=0.37 $X2=7.37 $Y2=0.715
r178 3 59 182 $w=1.7e-07 $l=4.37579e-07 $layer=licon1_NDIFF $count=1 $X=6.16
+ $Y=0.37 $X2=6.37 $Y2=0.715
r179 2 36 182 $w=1.7e-07 $l=5.30401e-07 $layer=licon1_NDIFF $count=1 $X=5.3
+ $Y=0.37 $X2=5.44 $Y2=0.835
r180 1 68 182 $w=1.7e-07 $l=6.62495e-07 $layer=licon1_NDIFF $count=1 $X=4.37
+ $Y=0.37 $X2=4.57 $Y2=0.94
.ends

.subckt PM_SKY130_FD_SC_HS__O22AI_4%A_877_368# 1 2 3 4 15 17 18 19 20 23 25 29
+ 32 35
c54 32 0 6.31714e-20 $X=4.535 $Y=2.355
r55 27 29 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=7.335 $Y=2.905
+ $X2=7.335 $Y2=2.455
r56 26 35 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.47 $Y=2.99
+ $X2=6.385 $Y2=2.99
r57 25 27 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=7.17 $Y=2.99
+ $X2=7.335 $Y2=2.905
r58 25 26 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=7.17 $Y=2.99 $X2=6.47
+ $Y2=2.99
r59 21 35 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.385 $Y=2.905
+ $X2=6.385 $Y2=2.99
r60 21 23 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=6.385 $Y=2.905
+ $X2=6.385 $Y2=2.455
r61 19 35 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.3 $Y=2.99 $X2=6.385
+ $Y2=2.99
r62 19 20 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=6.3 $Y=2.99 $X2=5.57
+ $Y2=2.99
r63 18 20 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=5.445 $Y=2.905
+ $X2=5.57 $Y2=2.99
r64 17 34 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.445 $Y=2.36
+ $X2=5.445 $Y2=2.275
r65 17 18 25.1233 $w=2.48e-07 $l=5.45e-07 $layer=LI1_cond $X=5.445 $Y=2.36
+ $X2=5.445 $Y2=2.905
r66 16 32 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.7 $Y=2.275
+ $X2=4.535 $Y2=2.275
r67 15 34 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.32 $Y=2.275
+ $X2=5.445 $Y2=2.275
r68 15 16 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=5.32 $Y=2.275
+ $X2=4.7 $Y2=2.275
r69 4 29 300 $w=1.7e-07 $l=7.03616e-07 $layer=licon1_PDIFF $count=2 $X=7.145
+ $Y=1.84 $X2=7.335 $Y2=2.455
r70 3 23 300 $w=1.7e-07 $l=6.85912e-07 $layer=licon1_PDIFF $count=2 $X=6.235
+ $Y=1.84 $X2=6.385 $Y2=2.455
r71 2 34 300 $w=1.7e-07 $l=6.06815e-07 $layer=licon1_PDIFF $count=2 $X=5.285
+ $Y=1.84 $X2=5.485 $Y2=2.355
r72 1 32 300 $w=1.7e-07 $l=5.85214e-07 $layer=licon1_PDIFF $count=2 $X=4.385
+ $Y=1.84 $X2=4.535 $Y2=2.355
.ends

.subckt PM_SKY130_FD_SC_HS__O22AI_4%A_27_74# 1 2 3 4 5 6 7 8 9 30 32 33 36 38 42
+ 44 48 50 52 53 54 64 68 70 73 76 77 79 80
c126 64 0 7.73112e-20 $X=1.25 $Y=0.925
c127 50 0 7.5396e-20 $X=3.905 $Y=0.925
c128 32 0 3.15663e-20 $X=1.125 $Y=1.065
r129 79 80 8.46017 $w=3.23e-07 $l=1.65e-07 $layer=LI1_cond $X=7.88 $Y=0.417
+ $X2=7.715 $Y2=0.417
r130 77 80 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=7.035 $Y=0.34
+ $X2=7.715 $Y2=0.34
r131 75 77 8.46017 $w=3.23e-07 $l=1.65e-07 $layer=LI1_cond $X=6.87 $Y=0.417
+ $X2=7.035 $Y2=0.417
r132 75 76 8.46017 $w=3.23e-07 $l=1.65e-07 $layer=LI1_cond $X=6.87 $Y=0.417
+ $X2=6.705 $Y2=0.417
r133 73 76 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=6.035 $Y=0.34
+ $X2=6.705 $Y2=0.34
r134 64 65 6.45368 $w=2.48e-07 $l=1.4e-07 $layer=LI1_cond $X=1.25 $Y=0.925
+ $X2=1.25 $Y2=1.065
r135 57 59 30.6727 $w=3.23e-07 $l=8.65e-07 $layer=LI1_cond $X=5.005 $Y=0.417
+ $X2=5.87 $Y2=0.417
r136 55 72 3.42929 $w=3.25e-07 $l=1.65e-07 $layer=LI1_cond $X=4.235 $Y=0.417
+ $X2=4.07 $Y2=0.417
r137 55 57 27.304 $w=3.23e-07 $l=7.7e-07 $layer=LI1_cond $X=4.235 $Y=0.417
+ $X2=5.005 $Y2=0.417
r138 54 73 8.35379 $w=3.23e-07 $l=1.62e-07 $layer=LI1_cond $X=5.873 $Y=0.417
+ $X2=6.035 $Y2=0.417
r139 54 59 0.106379 $w=3.23e-07 $l=3e-09 $layer=LI1_cond $X=5.873 $Y=0.417
+ $X2=5.87 $Y2=0.417
r140 52 72 3.38772 $w=3.3e-07 $l=1.63e-07 $layer=LI1_cond $X=4.07 $Y=0.58
+ $X2=4.07 $Y2=0.417
r141 52 53 9.07985 $w=3.28e-07 $l=2.6e-07 $layer=LI1_cond $X=4.07 $Y=0.58
+ $X2=4.07 $Y2=0.84
r142 51 70 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.235 $Y=0.925
+ $X2=3.11 $Y2=0.925
r143 50 53 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.905 $Y=0.925
+ $X2=4.07 $Y2=0.84
r144 50 51 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.905 $Y=0.925
+ $X2=3.235 $Y2=0.925
r145 46 70 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.11 $Y=0.84
+ $X2=3.11 $Y2=0.925
r146 46 48 14.9818 $w=2.48e-07 $l=3.25e-07 $layer=LI1_cond $X=3.11 $Y=0.84
+ $X2=3.11 $Y2=0.515
r147 45 68 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.305 $Y=0.925
+ $X2=2.18 $Y2=0.925
r148 44 70 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.985 $Y=0.925
+ $X2=3.11 $Y2=0.925
r149 44 45 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=2.985 $Y=0.925
+ $X2=2.305 $Y2=0.925
r150 40 68 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.18 $Y=0.84
+ $X2=2.18 $Y2=0.925
r151 40 42 14.9818 $w=2.48e-07 $l=3.25e-07 $layer=LI1_cond $X=2.18 $Y=0.84
+ $X2=2.18 $Y2=0.515
r152 39 64 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.375 $Y=0.925
+ $X2=1.25 $Y2=0.925
r153 38 68 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.055 $Y=0.925
+ $X2=2.18 $Y2=0.925
r154 38 39 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=2.055 $Y=0.925
+ $X2=1.375 $Y2=0.925
r155 34 64 3.91831 $w=2.48e-07 $l=8.5e-08 $layer=LI1_cond $X=1.25 $Y=0.84
+ $X2=1.25 $Y2=0.925
r156 34 36 14.9818 $w=2.48e-07 $l=3.25e-07 $layer=LI1_cond $X=1.25 $Y=0.84
+ $X2=1.25 $Y2=0.515
r157 32 65 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.125 $Y=1.065
+ $X2=1.25 $Y2=1.065
r158 32 33 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.125 $Y=1.065
+ $X2=0.445 $Y2=1.065
r159 28 33 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.28 $Y=0.98
+ $X2=0.445 $Y2=1.065
r160 28 30 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=0.28 $Y=0.98
+ $X2=0.28 $Y2=0.515
r161 9 79 182 $w=1.7e-07 $l=2.41454e-07 $layer=licon1_NDIFF $count=1 $X=7.66
+ $Y=0.37 $X2=7.88 $Y2=0.415
r162 8 75 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=6.66
+ $Y=0.37 $X2=6.87 $Y2=0.495
r163 7 59 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=5.73
+ $Y=0.37 $X2=5.87 $Y2=0.495
r164 6 57 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=4.86
+ $Y=0.37 $X2=5.005 $Y2=0.495
r165 5 72 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.93
+ $Y=0.37 $X2=4.07 $Y2=0.515
r166 4 70 182 $w=1.7e-07 $l=6.21068e-07 $layer=licon1_NDIFF $count=1 $X=2.93
+ $Y=0.37 $X2=3.07 $Y2=0.925
r167 4 48 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=2.93
+ $Y=0.37 $X2=3.07 $Y2=0.515
r168 3 68 182 $w=1.7e-07 $l=6.21068e-07 $layer=licon1_NDIFF $count=1 $X=2
+ $Y=0.37 $X2=2.14 $Y2=0.925
r169 3 42 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=2
+ $Y=0.37 $X2=2.14 $Y2=0.515
r170 2 36 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.07
+ $Y=0.37 $X2=1.21 $Y2=0.515
r171 1 30 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__O22AI_4%VGND 1 2 3 4 15 19 23 27 29 31 36 41 46 56
+ 57 60 63 66 69
r90 69 70 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r91 66 67 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r92 63 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r93 60 61 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r94 56 57 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=7.92 $Y=0
+ $X2=7.92 $Y2=0
r95 53 56 250.524 $w=1.68e-07 $l=3.84e-06 $layer=LI1_cond $X=4.08 $Y=0 $X2=7.92
+ $Y2=0
r96 51 69 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.735 $Y=0 $X2=3.57
+ $Y2=0
r97 51 53 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=3.735 $Y=0 $X2=4.08
+ $Y2=0
r98 50 70 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=3.6
+ $Y2=0
r99 50 67 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=2.64
+ $Y2=0
r100 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r101 47 66 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.805 $Y=0 $X2=2.64
+ $Y2=0
r102 47 49 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=2.805 $Y=0
+ $X2=3.12 $Y2=0
r103 46 69 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.405 $Y=0 $X2=3.57
+ $Y2=0
r104 46 49 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=3.405 $Y=0
+ $X2=3.12 $Y2=0
r105 45 67 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r106 45 64 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.68
+ $Y2=0
r107 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r108 42 63 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.875 $Y=0 $X2=1.71
+ $Y2=0
r109 42 44 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=1.875 $Y=0
+ $X2=2.16 $Y2=0
r110 41 66 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.475 $Y=0 $X2=2.64
+ $Y2=0
r111 41 44 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=2.475 $Y=0
+ $X2=2.16 $Y2=0
r112 40 64 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=1.68
+ $Y2=0
r113 40 61 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r114 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r115 37 60 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.945 $Y=0 $X2=0.78
+ $Y2=0
r116 37 39 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.945 $Y=0 $X2=1.2
+ $Y2=0
r117 36 63 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.545 $Y=0 $X2=1.71
+ $Y2=0
r118 36 39 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.545 $Y=0 $X2=1.2
+ $Y2=0
r119 34 61 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r120 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r121 31 60 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.615 $Y=0 $X2=0.78
+ $Y2=0
r122 31 33 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=0.615 $Y=0
+ $X2=0.24 $Y2=0
r123 29 57 1.07034 $w=4.9e-07 $l=3.84e-06 $layer=MET1_cond $X=4.08 $Y=0 $X2=7.92
+ $Y2=0
r124 29 70 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=3.6
+ $Y2=0
r125 29 53 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=4.08 $Y=0
+ $X2=4.08 $Y2=0
r126 25 69 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.57 $Y=0.085
+ $X2=3.57 $Y2=0
r127 25 27 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=3.57 $Y=0.085
+ $X2=3.57 $Y2=0.55
r128 21 66 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.64 $Y=0.085
+ $X2=2.64 $Y2=0
r129 21 23 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=2.64 $Y=0.085
+ $X2=2.64 $Y2=0.55
r130 17 63 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.71 $Y=0.085
+ $X2=1.71 $Y2=0
r131 17 19 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=1.71 $Y=0.085
+ $X2=1.71 $Y2=0.55
r132 13 60 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.78 $Y=0.085
+ $X2=0.78 $Y2=0
r133 13 15 18.6835 $w=3.28e-07 $l=5.35e-07 $layer=LI1_cond $X=0.78 $Y=0.085
+ $X2=0.78 $Y2=0.62
r134 4 27 182 $w=1.7e-07 $l=2.50998e-07 $layer=licon1_NDIFF $count=1 $X=3.4
+ $Y=0.37 $X2=3.57 $Y2=0.55
r135 3 23 182 $w=1.7e-07 $l=2.86182e-07 $layer=licon1_NDIFF $count=1 $X=2.43
+ $Y=0.37 $X2=2.64 $Y2=0.55
r136 2 19 182 $w=1.7e-07 $l=2.86182e-07 $layer=licon1_NDIFF $count=1 $X=1.5
+ $Y=0.37 $X2=1.71 $Y2=0.55
r137 1 15 182 $w=1.7e-07 $l=3.39116e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.37 $X2=0.78 $Y2=0.62
.ends

