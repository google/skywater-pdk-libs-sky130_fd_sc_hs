* File: sky130_fd_sc_hs__nor2b_4.spice
* Created: Tue Sep  1 20:11:20 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hs__nor2b_4.pex.spice"
.subckt sky130_fd_sc_hs__nor2b_4  VNB VPB A B_N VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* B_N	B_N
* A	A
* VPB	VPB
* VNB	VNB
MM1004 N_Y_M1004_d N_A_353_323#_M1004_g N_VGND_M1004_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.3223 PD=1.02 PS=2.57 NRD=0 NRS=61.704 M=1 R=4.93333 SA=75000.3
+ SB=75003 A=0.111 P=1.78 MULT=1
MM1009 N_Y_M1004_d N_A_353_323#_M1009_g N_VGND_M1009_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.4097 PD=1.02 PS=1.84 NRD=0 NRS=80.856 M=1 R=4.93333 SA=75000.7
+ SB=75002.6 A=0.111 P=1.78 MULT=1
MM1001 N_Y_M1001_d N_A_M1001_g N_VGND_M1009_s VNB NLOWVT L=0.15 W=0.74 AD=0.1036
+ AS=0.4097 PD=1.02 PS=1.84 NRD=0 NRS=80.856 M=1 R=4.93333 SA=75001.8 SB=75001.5
+ A=0.111 P=1.78 MULT=1
MM1005 N_Y_M1001_d N_A_M1005_g N_VGND_M1005_s VNB NLOWVT L=0.15 W=0.74 AD=0.1036
+ AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75002.2 SB=75001.1
+ A=0.111 P=1.78 MULT=1
MM1000 N_A_353_323#_M1000_d N_B_N_M1000_g N_VGND_M1005_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.518 AS=0.1036 PD=2.88 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75002.6
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1006 N_VPWR_M1006_d N_A_M1006_g N_A_116_368#_M1006_s VPB PSHORT L=0.15 W=1.12
+ AD=0.3304 AS=0.168 PD=2.83 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75004.2 A=0.168 P=2.54 MULT=1
MM1007 N_VPWR_M1007_d N_A_M1007_g N_A_116_368#_M1006_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.7 SB=75003.8 A=0.168 P=2.54 MULT=1
MM1008 N_VPWR_M1007_d N_A_M1008_g N_A_116_368#_M1008_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.1 SB=75003.3 A=0.168 P=2.54 MULT=1
MM1010 N_Y_M1010_d N_A_353_323#_M1010_g N_A_116_368#_M1008_s VPB PSHORT L=0.15
+ W=1.12 AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.6 SB=75002.9 A=0.168 P=2.54 MULT=1
MM1011 N_Y_M1010_d N_A_353_323#_M1011_g N_A_116_368#_M1011_s VPB PSHORT L=0.15
+ W=1.12 AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75002 SB=75002.4 A=0.168 P=2.54 MULT=1
MM1012 N_Y_M1012_d N_A_353_323#_M1012_g N_A_116_368#_M1011_s VPB PSHORT L=0.15
+ W=1.12 AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75002.5 SB=75002 A=0.168 P=2.54 MULT=1
MM1013 N_Y_M1012_d N_A_353_323#_M1013_g N_A_116_368#_M1013_s VPB PSHORT L=0.15
+ W=1.12 AD=0.168 AS=0.196 PD=1.42 PS=1.47 NRD=1.7533 NRS=10.5395 M=1 R=7.46667
+ SA=75002.9 SB=75001.5 A=0.168 P=2.54 MULT=1
MM1014 N_VPWR_M1014_d N_A_M1014_g N_A_116_368#_M1013_s VPB PSHORT L=0.15 W=1.12
+ AD=0.264 AS=0.196 PD=1.77714 PS=1.47 NRD=10.5395 NRS=1.7533 M=1 R=7.46667
+ SA=75003.4 SB=75001 A=0.168 P=2.54 MULT=1
MM1002 N_A_353_323#_M1002_d N_B_N_M1002_g N_VPWR_M1014_d VPB PSHORT L=0.15
+ W=0.84 AD=0.126 AS=0.198 PD=1.14 PS=1.33286 NRD=2.3443 NRS=22.655 M=1 R=5.6
+ SA=75004 SB=75000.7 A=0.126 P=1.98 MULT=1
MM1003 N_A_353_323#_M1002_d N_B_N_M1003_g N_VPWR_M1003_s VPB PSHORT L=0.15
+ W=0.84 AD=0.126 AS=0.2478 PD=1.14 PS=2.27 NRD=2.3443 NRS=2.3443 M=1 R=5.6
+ SA=75004.5 SB=75000.2 A=0.126 P=1.98 MULT=1
DX15_noxref VNB VPB NWDIODE A=10.5276 P=15.04
*
.include "sky130_fd_sc_hs__nor2b_4.pxi.spice"
*
.ends
*
*
