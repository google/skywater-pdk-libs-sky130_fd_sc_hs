* File: sky130_fd_sc_hs__a31oi_2.pex.spice
* Created: Tue Sep  1 19:53:13 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HS__A31OI_2%A3 1 3 4 6 7 9 10 12 13 15 21 27
c78 27 0 7.8613e-20 $X=0.27 $Y=1.175
c79 15 0 1.24498e-19 $X=1.95 $Y=1.175
c80 7 0 2.26479e-19 $X=1.925 $Y=1.22
r81 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.27
+ $Y=1.385 $X2=0.27 $Y2=1.385
r82 21 25 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=0.27 $Y=1.295 $X2=0.27
+ $Y2=1.385
r83 21 27 4.1907 $w=3.28e-07 $l=1.2e-07 $layer=LI1_cond $X=0.27 $Y=1.295
+ $X2=0.27 $Y2=1.175
r84 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.95
+ $Y=1.385 $X2=1.95 $Y2=1.385
r85 15 18 7.33373 $w=3.28e-07 $l=2.1e-07 $layer=LI1_cond $X=1.95 $Y=1.175
+ $X2=1.95 $Y2=1.385
r86 14 27 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.435 $Y=1.175
+ $X2=0.27 $Y2=1.175
r87 13 15 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.785 $Y=1.175
+ $X2=1.95 $Y2=1.175
r88 13 14 88.0749 $w=1.68e-07 $l=1.35e-06 $layer=LI1_cond $X=1.785 $Y=1.175
+ $X2=0.435 $Y2=1.175
r89 10 19 77.2841 $w=2.7e-07 $l=3.82492e-07 $layer=POLY_cond $X=1.955 $Y=1.765
+ $X2=1.95 $Y2=1.385
r90 10 12 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.955 $Y=1.765
+ $X2=1.955 $Y2=2.4
r91 7 19 38.9026 $w=2.7e-07 $l=1.77059e-07 $layer=POLY_cond $X=1.925 $Y=1.22
+ $X2=1.95 $Y2=1.385
r92 7 9 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.925 $Y=1.22 $X2=1.925
+ $Y2=0.74
r93 4 24 67.2473 $w=3.67e-07 $l=4.50888e-07 $layer=POLY_cond $X=0.505 $Y=1.765
+ $X2=0.35 $Y2=1.385
r94 4 6 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.505 $Y=1.765
+ $X2=0.505 $Y2=2.4
r95 1 24 39.0103 $w=3.67e-07 $l=2.26164e-07 $layer=POLY_cond $X=0.495 $Y=1.22
+ $X2=0.35 $Y2=1.385
r96 1 3 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=0.495 $Y=1.22 $X2=0.495
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HS__A31OI_2%A2 3 5 7 10 12 14 15 16 23 24
c55 24 0 7.8613e-20 $X=1.425 $Y=1.557
c56 5 0 1.71574e-19 $X=0.965 $Y=1.765
r57 24 25 3.94005 $w=3.67e-07 $l=3e-08 $layer=POLY_cond $X=1.425 $Y=1.557
+ $X2=1.455 $Y2=1.557
r58 22 24 5.91008 $w=3.67e-07 $l=4.5e-08 $layer=POLY_cond $X=1.38 $Y=1.557
+ $X2=1.425 $Y2=1.557
r59 22 23 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.38
+ $Y=1.515 $X2=1.38 $Y2=1.515
r60 20 22 54.5041 $w=3.67e-07 $l=4.15e-07 $layer=POLY_cond $X=0.965 $Y=1.557
+ $X2=1.38 $Y2=1.557
r61 19 20 5.25341 $w=3.67e-07 $l=4e-08 $layer=POLY_cond $X=0.925 $Y=1.557
+ $X2=0.965 $Y2=1.557
r62 16 23 5.92685 $w=3.48e-07 $l=1.8e-07 $layer=LI1_cond $X=1.2 $Y=1.605
+ $X2=1.38 $Y2=1.605
r63 15 16 15.8049 $w=3.48e-07 $l=4.8e-07 $layer=LI1_cond $X=0.72 $Y=1.605
+ $X2=1.2 $Y2=1.605
r64 12 25 23.77 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=1.455 $Y=1.765
+ $X2=1.455 $Y2=1.557
r65 12 14 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.455 $Y=1.765
+ $X2=1.455 $Y2=2.4
r66 8 24 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.425 $Y=1.35
+ $X2=1.425 $Y2=1.557
r67 8 10 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.425 $Y=1.35
+ $X2=1.425 $Y2=0.74
r68 5 20 23.77 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=0.965 $Y=1.765
+ $X2=0.965 $Y2=1.557
r69 5 7 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.965 $Y=1.765
+ $X2=0.965 $Y2=2.4
r70 1 19 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.925 $Y=1.35
+ $X2=0.925 $Y2=1.557
r71 1 3 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=0.925 $Y=1.35
+ $X2=0.925 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HS__A31OI_2%B1 1 3 4 6 7 9 10 15
c46 10 0 1.92056e-19 $X=2.64 $Y=1.295
r47 15 17 3.79101 $w=4.45e-07 $l=3.5e-08 $layer=POLY_cond $X=2.83 $Y=1.492
+ $X2=2.865 $Y2=1.492
r48 15 16 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.83
+ $Y=1.385 $X2=2.83 $Y2=1.385
r49 13 15 36.2854 $w=4.45e-07 $l=3.35e-07 $layer=POLY_cond $X=2.495 $Y=1.492
+ $X2=2.83 $Y2=1.492
r50 12 13 8.66517 $w=4.45e-07 $l=8e-08 $layer=POLY_cond $X=2.415 $Y=1.492
+ $X2=2.495 $Y2=1.492
r51 10 16 1.60667 $w=6.68e-07 $l=9e-08 $layer=LI1_cond $X=2.66 $Y=1.295 $X2=2.66
+ $Y2=1.385
r52 7 17 28.4889 $w=1.5e-07 $l=2.73e-07 $layer=POLY_cond $X=2.865 $Y=1.765
+ $X2=2.865 $Y2=1.492
r53 7 9 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.865 $Y=1.765
+ $X2=2.865 $Y2=2.4
r54 4 13 28.4889 $w=1.5e-07 $l=2.72e-07 $layer=POLY_cond $X=2.495 $Y=1.22
+ $X2=2.495 $Y2=1.492
r55 4 6 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=2.495 $Y=1.22 $X2=2.495
+ $Y2=0.74
r56 1 12 28.4889 $w=1.5e-07 $l=2.73e-07 $layer=POLY_cond $X=2.415 $Y=1.765
+ $X2=2.415 $Y2=1.492
r57 1 3 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.415 $Y=1.765
+ $X2=2.415 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_HS__A31OI_2%A1 3 5 7 10 12 14 15 22
c52 22 0 5.16637e-20 $X=3.755 $Y=1.557
r53 22 23 7.94506 $w=3.64e-07 $l=6e-08 $layer=POLY_cond $X=3.755 $Y=1.557
+ $X2=3.815 $Y2=1.557
r54 20 22 1.98626 $w=3.64e-07 $l=1.5e-08 $layer=POLY_cond $X=3.74 $Y=1.557
+ $X2=3.755 $Y2=1.557
r55 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.74
+ $Y=1.515 $X2=3.74 $Y2=1.515
r56 18 20 49.6566 $w=3.64e-07 $l=3.75e-07 $layer=POLY_cond $X=3.365 $Y=1.557
+ $X2=3.74 $Y2=1.557
r57 17 18 7.28297 $w=3.64e-07 $l=5.5e-08 $layer=POLY_cond $X=3.31 $Y=1.557
+ $X2=3.365 $Y2=1.557
r58 15 21 11.1952 $w=3.48e-07 $l=3.4e-07 $layer=LI1_cond $X=4.08 $Y=1.605
+ $X2=3.74 $Y2=1.605
r59 12 23 23.572 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=3.815 $Y=1.765
+ $X2=3.815 $Y2=1.557
r60 12 14 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.815 $Y=1.765
+ $X2=3.815 $Y2=2.4
r61 8 22 23.572 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.755 $Y=1.35
+ $X2=3.755 $Y2=1.557
r62 8 10 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=3.755 $Y=1.35
+ $X2=3.755 $Y2=0.74
r63 5 18 23.572 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=3.365 $Y=1.765
+ $X2=3.365 $Y2=1.557
r64 5 7 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.365 $Y=1.765
+ $X2=3.365 $Y2=2.4
r65 1 17 23.572 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.31 $Y=1.35 $X2=3.31
+ $Y2=1.557
r66 1 3 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=3.31 $Y=1.35 $X2=3.31
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HS__A31OI_2%A_27_368# 1 2 3 4 5 16 18 20 24 26 28 31 32
+ 33 34 38 40 42 47
c68 24 0 1.71574e-19 $X=1.23 $Y=2.815
r69 40 53 3.15431 $w=2.8e-07 $l=1.51987e-07 $layer=LI1_cond $X=4.065 $Y=2.23
+ $X2=4.04 $Y2=2.09
r70 40 42 9.67229 $w=2.78e-07 $l=2.35e-07 $layer=LI1_cond $X=4.065 $Y=2.23
+ $X2=4.065 $Y2=2.465
r71 39 51 4.57959 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=3.255 $Y=2.145
+ $X2=3.115 $Y2=2.145
r72 38 53 4.20574 $w=1.7e-07 $l=1.90526e-07 $layer=LI1_cond $X=3.875 $Y=2.145
+ $X2=4.04 $Y2=2.09
r73 38 39 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=3.875 $Y=2.145
+ $X2=3.255 $Y2=2.145
r74 35 37 17.2866 $w=2.78e-07 $l=4.2e-07 $layer=LI1_cond $X=3.115 $Y=2.905
+ $X2=3.115 $Y2=2.485
r75 34 51 2.78046 $w=2.8e-07 $l=8.5e-08 $layer=LI1_cond $X=3.115 $Y=2.23
+ $X2=3.115 $Y2=2.145
r76 34 37 10.4955 $w=2.78e-07 $l=2.55e-07 $layer=LI1_cond $X=3.115 $Y=2.23
+ $X2=3.115 $Y2=2.485
r77 32 35 7.36005 $w=1.7e-07 $l=1.77482e-07 $layer=LI1_cond $X=2.975 $Y=2.99
+ $X2=3.115 $Y2=2.905
r78 32 33 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=2.975 $Y=2.99
+ $X2=2.275 $Y2=2.99
r79 29 33 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=2.145 $Y=2.905
+ $X2=2.275 $Y2=2.99
r80 29 31 4.87572 $w=2.58e-07 $l=1.1e-07 $layer=LI1_cond $X=2.145 $Y=2.905
+ $X2=2.145 $Y2=2.795
r81 28 49 2.85134 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=2.145 $Y=2.12
+ $X2=2.145 $Y2=2.035
r82 28 31 29.9192 $w=2.58e-07 $l=6.75e-07 $layer=LI1_cond $X=2.145 $Y=2.12
+ $X2=2.145 $Y2=2.795
r83 27 47 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.395 $Y=2.035
+ $X2=1.23 $Y2=2.035
r84 26 49 4.36088 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.015 $Y=2.035
+ $X2=2.145 $Y2=2.035
r85 26 27 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=2.015 $Y=2.035
+ $X2=1.395 $Y2=2.035
r86 22 47 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.23 $Y=2.12 $X2=1.23
+ $Y2=2.035
r87 22 24 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=1.23 $Y=2.12
+ $X2=1.23 $Y2=2.815
r88 21 45 3.99177 $w=1.7e-07 $l=1.5411e-07 $layer=LI1_cond $X=0.365 $Y=2.035
+ $X2=0.24 $Y2=1.97
r89 20 47 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.065 $Y=2.035
+ $X2=1.23 $Y2=2.035
r90 20 21 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=1.065 $Y=2.035
+ $X2=0.365 $Y2=2.035
r91 16 45 3.1514 $w=2.5e-07 $l=1.5e-07 $layer=LI1_cond $X=0.24 $Y=2.12 $X2=0.24
+ $Y2=1.97
r92 16 18 12.9074 $w=2.48e-07 $l=2.8e-07 $layer=LI1_cond $X=0.24 $Y=2.12
+ $X2=0.24 $Y2=2.4
r93 5 53 600 $w=1.7e-07 $l=3.4187e-07 $layer=licon1_PDIFF $count=1 $X=3.89
+ $Y=1.84 $X2=4.04 $Y2=2.115
r94 5 42 300 $w=1.7e-07 $l=6.95971e-07 $layer=licon1_PDIFF $count=2 $X=3.89
+ $Y=1.84 $X2=4.04 $Y2=2.465
r95 4 51 600 $w=1.7e-07 $l=3.9246e-07 $layer=licon1_PDIFF $count=1 $X=2.94
+ $Y=1.84 $X2=3.14 $Y2=2.145
r96 4 37 300 $w=1.7e-07 $l=7.38258e-07 $layer=licon1_PDIFF $count=2 $X=2.94
+ $Y=1.84 $X2=3.14 $Y2=2.485
r97 3 49 400 $w=1.7e-07 $l=3.43875e-07 $layer=licon1_PDIFF $count=1 $X=2.03
+ $Y=1.84 $X2=2.185 $Y2=2.115
r98 3 31 400 $w=1.7e-07 $l=1.02959e-06 $layer=licon1_PDIFF $count=1 $X=2.03
+ $Y=1.84 $X2=2.185 $Y2=2.795
r99 2 47 400 $w=1.7e-07 $l=2.79285e-07 $layer=licon1_PDIFF $count=1 $X=1.04
+ $Y=1.84 $X2=1.23 $Y2=2.04
r100 2 24 400 $w=1.7e-07 $l=1.06577e-06 $layer=licon1_PDIFF $count=1 $X=1.04
+ $Y=1.84 $X2=1.23 $Y2=2.815
r101 1 45 600 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=1.985
r102 1 18 300 $w=1.7e-07 $l=6.28331e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_HS__A31OI_2%VPWR 1 2 3 12 16 20 22 24 29 34 44 45 48 51
+ 54
r58 54 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r59 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r60 48 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r61 45 55 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=3.6 $Y2=3.33
r62 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r63 42 54 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.755 $Y=3.33
+ $X2=3.59 $Y2=3.33
r64 42 44 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=3.755 $Y=3.33
+ $X2=4.08 $Y2=3.33
r65 41 55 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=3.6 $Y2=3.33
r66 40 41 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r67 37 40 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=2.16 $Y=3.33 $X2=3.12
+ $Y2=3.33
r68 35 51 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.845 $Y=3.33
+ $X2=1.72 $Y2=3.33
r69 35 37 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=1.845 $Y=3.33
+ $X2=2.16 $Y2=3.33
r70 34 54 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.425 $Y=3.33
+ $X2=3.59 $Y2=3.33
r71 34 40 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=3.425 $Y=3.33
+ $X2=3.12 $Y2=3.33
r72 33 52 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=1.68 $Y2=3.33
r73 33 49 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r74 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r75 30 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.895 $Y=3.33
+ $X2=0.73 $Y2=3.33
r76 30 32 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.895 $Y=3.33
+ $X2=1.2 $Y2=3.33
r77 29 51 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.595 $Y=3.33
+ $X2=1.72 $Y2=3.33
r78 29 32 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=1.595 $Y=3.33
+ $X2=1.2 $Y2=3.33
r79 27 49 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r80 26 27 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r81 24 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.565 $Y=3.33
+ $X2=0.73 $Y2=3.33
r82 24 26 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.565 $Y=3.33
+ $X2=0.24 $Y2=3.33
r83 22 41 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=3.12 $Y2=3.33
r84 22 52 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.68 $Y2=3.33
r85 22 37 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r86 18 54 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.59 $Y=3.245
+ $X2=3.59 $Y2=3.33
r87 18 20 26.1919 $w=3.28e-07 $l=7.5e-07 $layer=LI1_cond $X=3.59 $Y=3.245
+ $X2=3.59 $Y2=2.495
r88 14 51 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.72 $Y=3.245
+ $X2=1.72 $Y2=3.33
r89 14 16 36.4172 $w=2.48e-07 $l=7.9e-07 $layer=LI1_cond $X=1.72 $Y=3.245
+ $X2=1.72 $Y2=2.455
r90 10 48 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.73 $Y=3.245
+ $X2=0.73 $Y2=3.33
r91 10 12 29.1603 $w=3.28e-07 $l=8.35e-07 $layer=LI1_cond $X=0.73 $Y=3.245
+ $X2=0.73 $Y2=2.41
r92 3 20 300 $w=1.7e-07 $l=7.26137e-07 $layer=licon1_PDIFF $count=2 $X=3.44
+ $Y=1.84 $X2=3.59 $Y2=2.495
r93 2 16 300 $w=1.7e-07 $l=6.85912e-07 $layer=licon1_PDIFF $count=2 $X=1.53
+ $Y=1.84 $X2=1.68 $Y2=2.455
r94 1 12 300 $w=1.7e-07 $l=6.40625e-07 $layer=licon1_PDIFF $count=2 $X=0.58
+ $Y=1.84 $X2=0.73 $Y2=2.41
.ends

.subckt PM_SKY130_FD_SC_HS__A31OI_2%Y 1 2 3 12 16 20 21 23 24 26 27 28 31 32
r65 31 32 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=4.04 $Y=0.515
+ $X2=4.04 $Y2=0.925
r66 30 32 5.76222 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=4.04 $Y=1.09
+ $X2=4.04 $Y2=0.925
r67 29 31 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=4.04 $Y=0.425 $X2=4.04
+ $Y2=0.515
r68 26 30 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.875 $Y=1.175
+ $X2=4.04 $Y2=1.09
r69 26 27 35.2299 $w=1.68e-07 $l=5.4e-07 $layer=LI1_cond $X=3.875 $Y=1.175
+ $X2=3.335 $Y2=1.175
r70 24 29 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.875 $Y=0.34
+ $X2=4.04 $Y2=0.425
r71 24 28 40.123 $w=1.68e-07 $l=6.15e-07 $layer=LI1_cond $X=3.875 $Y=0.34
+ $X2=3.26 $Y2=0.34
r72 22 27 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.25 $Y=1.26
+ $X2=3.335 $Y2=1.175
r73 22 23 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=3.25 $Y=1.26
+ $X2=3.25 $Y2=1.72
r74 20 23 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.165 $Y=1.805
+ $X2=3.25 $Y2=1.72
r75 20 21 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=3.165 $Y=1.805
+ $X2=2.805 $Y2=1.805
r76 16 28 8.35379 $w=3.23e-07 $l=1.62e-07 $layer=LI1_cond $X=3.098 $Y=0.417
+ $X2=3.26 $Y2=0.417
r77 16 18 0.106379 $w=3.23e-07 $l=3e-09 $layer=LI1_cond $X=3.098 $Y=0.417
+ $X2=3.095 $Y2=0.417
r78 12 14 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=2.64 $Y=1.965
+ $X2=2.64 $Y2=2.645
r79 10 21 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.64 $Y=1.89
+ $X2=2.805 $Y2=1.805
r80 10 12 2.61919 $w=3.28e-07 $l=7.5e-08 $layer=LI1_cond $X=2.64 $Y=1.89
+ $X2=2.64 $Y2=1.965
r81 3 14 400 $w=1.7e-07 $l=8.76798e-07 $layer=licon1_PDIFF $count=1 $X=2.49
+ $Y=1.84 $X2=2.64 $Y2=2.645
r82 3 12 400 $w=1.7e-07 $l=2.03101e-07 $layer=licon1_PDIFF $count=1 $X=2.49
+ $Y=1.84 $X2=2.64 $Y2=1.965
r83 2 31 91 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=2 $X=3.83
+ $Y=0.37 $X2=4.04 $Y2=0.515
r84 1 18 91 $w=1.7e-07 $l=5.84166e-07 $layer=licon1_NDIFF $count=2 $X=2.57
+ $Y=0.37 $X2=3.095 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_HS__A31OI_2%VGND 1 2 7 9 13 15 17 30 31 37
r46 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r47 30 31 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r48 28 31 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=2.64 $Y=0 $X2=4.08
+ $Y2=0
r49 27 30 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=2.64 $Y=0 $X2=4.08
+ $Y2=0
r50 27 28 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r51 25 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.375 $Y=0 $X2=2.21
+ $Y2=0
r52 25 27 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=2.375 $Y=0 $X2=2.64
+ $Y2=0
r53 23 24 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r54 21 24 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r55 21 35 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r56 20 23 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r57 20 21 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r58 18 34 4.00981 $w=1.7e-07 $l=1.83e-07 $layer=LI1_cond $X=0.365 $Y=0 $X2=0.182
+ $Y2=0
r59 18 20 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=0.365 $Y=0 $X2=0.72
+ $Y2=0
r60 17 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.045 $Y=0 $X2=2.21
+ $Y2=0
r61 17 23 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=2.045 $Y=0 $X2=1.68
+ $Y2=0
r62 15 28 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r63 15 24 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.68
+ $Y2=0
r64 15 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r65 11 37 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.21 $Y=0.085
+ $X2=2.21 $Y2=0
r66 11 13 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=2.21 $Y=0.085
+ $X2=2.21 $Y2=0.495
r67 7 34 3.13335 $w=2.5e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.24 $Y=0.085
+ $X2=0.182 $Y2=0
r68 7 9 29.5025 $w=2.48e-07 $l=6.4e-07 $layer=LI1_cond $X=0.24 $Y=0.085 $X2=0.24
+ $Y2=0.725
r69 2 13 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=2 $Y=0.37
+ $X2=2.21 $Y2=0.495
r70 1 9 182 $w=1.7e-07 $l=4.21307e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.725
.ends

.subckt PM_SKY130_FD_SC_HS__A31OI_2%A_114_74# 1 2 9 11 12 13
c29 11 0 8.60869e-20 $X=1.545 $Y=0.34
c30 2 0 1.24498e-19 $X=1.5 $Y=0.37
r31 13 16 5.41299 $w=3.28e-07 $l=1.55e-07 $layer=LI1_cond $X=1.71 $Y=0.34
+ $X2=1.71 $Y2=0.495
r32 11 13 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.545 $Y=0.34
+ $X2=1.71 $Y2=0.34
r33 11 12 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.545 $Y=0.34
+ $X2=0.875 $Y2=0.34
r34 7 12 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.71 $Y=0.425
+ $X2=0.875 $Y2=0.34
r35 7 9 2.44458 $w=3.28e-07 $l=7e-08 $layer=LI1_cond $X=0.71 $Y=0.425 $X2=0.71
+ $Y2=0.495
r36 2 16 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=1.5
+ $Y=0.37 $X2=1.71 $Y2=0.495
r37 1 9 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=0.57
+ $Y=0.37 $X2=0.71 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_HS__A31OI_2%A_200_74# 1 2 12 14 15
r31 14 15 6.2579 $w=2.48e-07 $l=1.1e-07 $layer=LI1_cond $X=3.54 $Y=0.795
+ $X2=3.43 $Y2=0.795
r32 12 15 134.07 $w=1.68e-07 $l=2.055e-06 $layer=LI1_cond $X=1.375 $Y=0.835
+ $X2=3.43 $Y2=0.835
r33 10 12 8.46017 $w=3.23e-07 $l=1.65e-07 $layer=LI1_cond $X=1.21 $Y=0.757
+ $X2=1.375 $Y2=0.757
r34 2 14 182 $w=1.7e-07 $l=5.36936e-07 $layer=licon1_NDIFF $count=1 $X=3.385
+ $Y=0.37 $X2=3.54 $Y2=0.835
r35 1 10 182 $w=1.7e-07 $l=5.19495e-07 $layer=licon1_NDIFF $count=1 $X=1 $Y=0.37
+ $X2=1.21 $Y2=0.795
.ends

