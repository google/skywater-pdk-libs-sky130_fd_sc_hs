* File: sky130_fd_sc_hs__ha_1.pxi.spice
* Created: Tue Sep  1 20:06:29 2020
* 
x_PM_SKY130_FD_SC_HS__HA_1%A_83_260# N_A_83_260#_M1009_s N_A_83_260#_M1007_d
+ N_A_83_260#_M1012_g N_A_83_260#_c_89_n N_A_83_260#_M1006_g N_A_83_260#_c_90_n
+ N_A_83_260#_c_91_n N_A_83_260#_c_92_n N_A_83_260#_c_100_p N_A_83_260#_c_126_p
+ N_A_83_260#_c_93_n N_A_83_260#_c_96_n PM_SKY130_FD_SC_HS__HA_1%A_83_260#
x_PM_SKY130_FD_SC_HS__HA_1%A_239_294# N_A_239_294#_M1001_s N_A_239_294#_M1002_d
+ N_A_239_294#_c_147_n N_A_239_294#_M1007_g N_A_239_294#_M1009_g
+ N_A_239_294#_c_149_n N_A_239_294#_M1000_g N_A_239_294#_c_150_n
+ N_A_239_294#_M1003_g N_A_239_294#_c_151_n N_A_239_294#_c_158_n
+ N_A_239_294#_c_178_n N_A_239_294#_c_152_n N_A_239_294#_c_159_n
+ N_A_239_294#_c_160_n N_A_239_294#_c_153_n N_A_239_294#_c_154_n
+ N_A_239_294#_c_162_n PM_SKY130_FD_SC_HS__HA_1%A_239_294#
x_PM_SKY130_FD_SC_HS__HA_1%B N_B_c_259_n N_B_M1005_g N_B_M1010_g N_B_c_267_n
+ N_B_c_268_n N_B_M1002_g N_B_M1001_g N_B_c_262_n B N_B_c_264_n N_B_c_265_n
+ PM_SKY130_FD_SC_HS__HA_1%B
x_PM_SKY130_FD_SC_HS__HA_1%A N_A_M1013_g N_A_c_325_n N_A_c_326_n N_A_c_332_n
+ N_A_M1008_g N_A_c_327_n N_A_c_333_n N_A_M1004_g N_A_c_334_n N_A_M1011_g A
+ N_A_c_329_n N_A_c_330_n PM_SKY130_FD_SC_HS__HA_1%A
x_PM_SKY130_FD_SC_HS__HA_1%SUM N_SUM_M1012_s N_SUM_M1006_s SUM SUM SUM SUM SUM
+ SUM SUM SUM SUM PM_SKY130_FD_SC_HS__HA_1%SUM
x_PM_SKY130_FD_SC_HS__HA_1%VPWR N_VPWR_M1006_d N_VPWR_M1008_d N_VPWR_M1004_d
+ N_VPWR_c_419_n N_VPWR_c_420_n N_VPWR_c_421_n N_VPWR_c_422_n N_VPWR_c_423_n
+ VPWR N_VPWR_c_424_n N_VPWR_c_425_n N_VPWR_c_426_n N_VPWR_c_418_n
+ N_VPWR_c_428_n N_VPWR_c_429_n PM_SKY130_FD_SC_HS__HA_1%VPWR
x_PM_SKY130_FD_SC_HS__HA_1%COUT N_COUT_M1003_d N_COUT_M1000_d N_COUT_c_480_n
+ N_COUT_c_481_n COUT COUT COUT N_COUT_c_482_n PM_SKY130_FD_SC_HS__HA_1%COUT
x_PM_SKY130_FD_SC_HS__HA_1%VGND N_VGND_M1012_d N_VGND_M1010_d N_VGND_M1011_d
+ N_VGND_c_504_n N_VGND_c_505_n N_VGND_c_506_n N_VGND_c_507_n N_VGND_c_508_n
+ VGND N_VGND_c_509_n N_VGND_c_510_n N_VGND_c_511_n N_VGND_c_512_n
+ N_VGND_c_513_n N_VGND_c_514_n PM_SKY130_FD_SC_HS__HA_1%VGND
x_PM_SKY130_FD_SC_HS__HA_1%A_305_130# N_A_305_130#_M1009_d N_A_305_130#_M1013_d
+ N_A_305_130#_c_559_n N_A_305_130#_c_560_n N_A_305_130#_c_561_n
+ N_A_305_130#_c_562_n PM_SKY130_FD_SC_HS__HA_1%A_305_130#
cc_1 VNB N_A_83_260#_M1012_g 0.027038f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_2 VNB N_A_83_260#_c_89_n 0.04702f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.765
cc_3 VNB N_A_83_260#_c_90_n 0.01342f $X=-0.19 $Y=-0.245 $X2=0.77 $Y2=1.63
cc_4 VNB N_A_83_260#_c_91_n 4.54332e-19 $X=-0.19 $Y=-0.245 $X2=0.77 $Y2=2.31
cc_5 VNB N_A_83_260#_c_92_n 0.0148545f $X=-0.19 $Y=-0.245 $X2=1.07 $Y2=1.215
cc_6 VNB N_A_83_260#_c_93_n 0.0112018f $X=-0.19 $Y=-0.245 $X2=1.235 $Y2=1.105
cc_7 VNB N_A_239_294#_c_147_n 0.0194828f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.3
cc_8 VNB N_A_239_294#_M1009_g 0.0239995f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_9 VNB N_A_239_294#_c_149_n 0.0284825f $X=-0.19 $Y=-0.245 $X2=0.77 $Y2=1.63
cc_10 VNB N_A_239_294#_c_150_n 0.0216579f $X=-0.19 $Y=-0.245 $X2=0.855 $Y2=1.215
cc_11 VNB N_A_239_294#_c_151_n 0.00167715f $X=-0.19 $Y=-0.245 $X2=0.69 $Y2=1.465
cc_12 VNB N_A_239_294#_c_152_n 0.00810984f $X=-0.19 $Y=-0.245 $X2=1.575
+ $Y2=2.395
cc_13 VNB N_A_239_294#_c_153_n 0.00508564f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_239_294#_c_154_n 0.00648904f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_B_c_259_n 0.0224338f $X=-0.19 $Y=-0.245 $X2=1.09 $Y2=0.93
cc_16 VNB N_B_M1010_g 0.0215777f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_B_M1001_g 0.0251318f $X=-0.19 $Y=-0.245 $X2=0.77 $Y2=2.31
cc_18 VNB N_B_c_262_n 0.00305816f $X=-0.19 $Y=-0.245 $X2=0.69 $Y2=1.465
cc_19 VNB B 0.00105506f $X=-0.19 $Y=-0.245 $X2=1.235 $Y2=1.105
cc_20 VNB N_B_c_264_n 0.0341314f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_B_c_265_n 0.0124882f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_M1013_g 0.0132214f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_c_325_n 0.00793984f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_c_326_n 0.0144568f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_c_327_n 0.0792528f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_M1011_g 0.0417945f $X=-0.19 $Y=-0.245 $X2=1.41 $Y2=2.395
cc_27 VNB N_A_c_329_n 0.0734688f $X=-0.19 $Y=-0.245 $X2=0.69 $Y2=1.465
cc_28 VNB N_A_c_330_n 0.00343837f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB SUM 0.0259999f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.3
cc_30 VNB SUM 0.00884344f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_31 VNB SUM 0.0260472f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_32 VNB N_VPWR_c_418_n 0.203486f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_COUT_c_480_n 0.0250027f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_34 VNB N_COUT_c_481_n 0.00842165f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_35 VNB N_COUT_c_482_n 0.0224443f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_504_n 0.0224413f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_37 VNB N_VGND_c_505_n 0.0219598f $X=-0.19 $Y=-0.245 $X2=1.07 $Y2=1.215
cc_38 VNB N_VGND_c_506_n 0.00977234f $X=-0.19 $Y=-0.245 $X2=0.69 $Y2=1.215
cc_39 VNB N_VGND_c_507_n 0.042621f $X=-0.19 $Y=-0.245 $X2=0.69 $Y2=1.465
cc_40 VNB N_VGND_c_508_n 0.00513431f $X=-0.19 $Y=-0.245 $X2=1.235 $Y2=1.105
cc_41 VNB N_VGND_c_509_n 0.0194697f $X=-0.19 $Y=-0.245 $X2=1.235 $Y2=1.215
cc_42 VNB N_VGND_c_510_n 0.0327532f $X=-0.19 $Y=-0.245 $X2=1.575 $Y2=2.555
cc_43 VNB N_VGND_c_511_n 0.0206833f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_512_n 0.294725f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_VGND_c_513_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_VGND_c_514_n 0.00672884f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_305_130#_c_559_n 0.00261785f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_48 VNB N_A_305_130#_c_560_n 0.00125648f $X=-0.19 $Y=-0.245 $X2=0.505
+ $Y2=1.765
cc_49 VNB N_A_305_130#_c_561_n 0.00296164f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_50 VNB N_A_305_130#_c_562_n 0.00837552f $X=-0.19 $Y=-0.245 $X2=0.77 $Y2=1.63
cc_51 VPB N_A_83_260#_c_89_n 0.0290015f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.765
cc_52 VPB N_A_83_260#_c_91_n 0.00409439f $X=-0.19 $Y=1.66 $X2=0.77 $Y2=2.31
cc_53 VPB N_A_83_260#_c_96_n 3.75654e-19 $X=-0.19 $Y=1.66 $X2=1.575 $Y2=2.395
cc_54 VPB N_A_239_294#_c_147_n 0.0385744f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.3
cc_55 VPB N_A_239_294#_c_149_n 0.0337705f $X=-0.19 $Y=1.66 $X2=0.77 $Y2=1.63
cc_56 VPB N_A_239_294#_c_151_n 0.00333531f $X=-0.19 $Y=1.66 $X2=0.69 $Y2=1.465
cc_57 VPB N_A_239_294#_c_158_n 0.00436551f $X=-0.19 $Y=1.66 $X2=1.235 $Y2=1.105
cc_58 VPB N_A_239_294#_c_159_n 0.00243101f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_59 VPB N_A_239_294#_c_160_n 0.00391423f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_60 VPB N_A_239_294#_c_154_n 0.00347087f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_61 VPB N_A_239_294#_c_162_n 0.00145462f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_62 VPB N_B_c_259_n 0.0295763f $X=-0.19 $Y=1.66 $X2=1.09 $Y2=0.93
cc_63 VPB N_B_c_267_n 0.0106065f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.74
cc_64 VPB N_B_c_268_n 0.0225647f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_65 VPB N_B_c_264_n 0.0117015f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_66 VPB N_B_c_265_n 0.00647563f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_67 VPB N_A_c_326_n 6.97741e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_68 VPB N_A_c_332_n 0.0254321f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.3
cc_69 VPB N_A_c_333_n 0.0164489f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.4
cc_70 VPB N_A_c_334_n 0.0157028f $X=-0.19 $Y=1.66 $X2=1.07 $Y2=1.215
cc_71 VPB N_A_M1011_g 0.011206f $X=-0.19 $Y=1.66 $X2=1.41 $Y2=2.395
cc_72 VPB SUM 0.00764839f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.74
cc_73 VPB SUM 0.0494776f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.765
cc_74 VPB N_VPWR_c_419_n 0.0154148f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.4
cc_75 VPB N_VPWR_c_420_n 0.00667644f $X=-0.19 $Y=1.66 $X2=1.07 $Y2=1.215
cc_76 VPB N_VPWR_c_421_n 0.010309f $X=-0.19 $Y=1.66 $X2=0.69 $Y2=1.215
cc_77 VPB N_VPWR_c_422_n 0.0173363f $X=-0.19 $Y=1.66 $X2=0.69 $Y2=1.465
cc_78 VPB N_VPWR_c_423_n 0.00632158f $X=-0.19 $Y=1.66 $X2=1.235 $Y2=1.105
cc_79 VPB N_VPWR_c_424_n 0.0191515f $X=-0.19 $Y=1.66 $X2=1.235 $Y2=1.215
cc_80 VPB N_VPWR_c_425_n 0.0387125f $X=-0.19 $Y=1.66 $X2=1.575 $Y2=2.555
cc_81 VPB N_VPWR_c_426_n 0.0199976f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_82 VPB N_VPWR_c_418_n 0.082349f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_83 VPB N_VPWR_c_428_n 0.0113226f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_84 VPB N_VPWR_c_429_n 0.013174f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_85 VPB COUT 0.0504915f $X=-0.19 $Y=1.66 $X2=0.77 $Y2=1.63
cc_86 VPB N_COUT_c_482_n 0.00919412f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_87 N_A_83_260#_c_89_n N_A_239_294#_c_147_n 0.019895f $X=0.505 $Y=1.765 $X2=0
+ $Y2=0
cc_88 N_A_83_260#_c_90_n N_A_239_294#_c_147_n 6.56648e-19 $X=0.77 $Y=1.63 $X2=0
+ $Y2=0
cc_89 N_A_83_260#_c_91_n N_A_239_294#_c_147_n 0.00571062f $X=0.77 $Y=2.31 $X2=0
+ $Y2=0
cc_90 N_A_83_260#_c_100_p N_A_239_294#_c_147_n 0.0110652f $X=1.41 $Y=2.395 $X2=0
+ $Y2=0
cc_91 N_A_83_260#_c_93_n N_A_239_294#_c_147_n 0.00133607f $X=1.235 $Y=1.105
+ $X2=0 $Y2=0
cc_92 N_A_83_260#_c_96_n N_A_239_294#_c_147_n 0.0115268f $X=1.575 $Y=2.395 $X2=0
+ $Y2=0
cc_93 N_A_83_260#_c_89_n N_A_239_294#_M1009_g 0.00305941f $X=0.505 $Y=1.765
+ $X2=0 $Y2=0
cc_94 N_A_83_260#_c_90_n N_A_239_294#_M1009_g 8.95785e-19 $X=0.77 $Y=1.63 $X2=0
+ $Y2=0
cc_95 N_A_83_260#_c_93_n N_A_239_294#_M1009_g 0.00554476f $X=1.235 $Y=1.105
+ $X2=0 $Y2=0
cc_96 N_A_83_260#_c_89_n N_A_239_294#_c_151_n 2.02974e-19 $X=0.505 $Y=1.765
+ $X2=0 $Y2=0
cc_97 N_A_83_260#_c_90_n N_A_239_294#_c_151_n 0.00690853f $X=0.77 $Y=1.63 $X2=0
+ $Y2=0
cc_98 N_A_83_260#_c_91_n N_A_239_294#_c_151_n 0.0158825f $X=0.77 $Y=2.31 $X2=0
+ $Y2=0
cc_99 N_A_83_260#_c_93_n N_A_239_294#_c_151_n 0.0172163f $X=1.235 $Y=1.105 $X2=0
+ $Y2=0
cc_100 N_A_83_260#_M1007_d N_A_239_294#_c_158_n 0.00717012f $X=1.425 $Y=1.96
+ $X2=0 $Y2=0
cc_101 N_A_83_260#_c_96_n N_A_239_294#_c_158_n 0.0156509f $X=1.575 $Y=2.395
+ $X2=0 $Y2=0
cc_102 N_A_83_260#_M1007_d N_A_239_294#_c_178_n 4.64572e-19 $X=1.425 $Y=1.96
+ $X2=0 $Y2=0
cc_103 N_A_83_260#_c_91_n N_A_239_294#_c_178_n 0.00829137f $X=0.77 $Y=2.31 $X2=0
+ $Y2=0
cc_104 N_A_83_260#_c_100_p N_A_239_294#_c_178_n 0.0120951f $X=1.41 $Y=2.395
+ $X2=0 $Y2=0
cc_105 N_A_83_260#_c_96_n N_A_239_294#_c_178_n 0.00489071f $X=1.575 $Y=2.395
+ $X2=0 $Y2=0
cc_106 N_A_83_260#_M1012_g SUM 0.0128374f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_107 N_A_83_260#_c_93_n SUM 0.00647958f $X=1.235 $Y=1.105 $X2=0 $Y2=0
cc_108 N_A_83_260#_M1012_g SUM 0.00515125f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_109 N_A_83_260#_c_89_n SUM 2.30445e-19 $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_110 N_A_83_260#_M1012_g SUM 0.00409755f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_111 N_A_83_260#_c_89_n SUM 0.0137115f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_112 N_A_83_260#_c_90_n SUM 0.0344043f $X=0.77 $Y=1.63 $X2=0 $Y2=0
cc_113 N_A_83_260#_c_91_n SUM 0.0092039f $X=0.77 $Y=2.31 $X2=0 $Y2=0
cc_114 N_A_83_260#_c_89_n SUM 0.0217542f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_115 N_A_83_260#_c_91_n SUM 0.0277247f $X=0.77 $Y=2.31 $X2=0 $Y2=0
cc_116 N_A_83_260#_c_126_p SUM 0.0107657f $X=0.855 $Y=2.395 $X2=0 $Y2=0
cc_117 N_A_83_260#_c_91_n N_VPWR_M1006_d 0.0133604f $X=0.77 $Y=2.31 $X2=-0.19
+ $Y2=-0.245
cc_118 N_A_83_260#_c_100_p N_VPWR_M1006_d 0.0193014f $X=1.41 $Y=2.395 $X2=-0.19
+ $Y2=-0.245
cc_119 N_A_83_260#_c_126_p N_VPWR_M1006_d 0.00510195f $X=0.855 $Y=2.395
+ $X2=-0.19 $Y2=-0.245
cc_120 N_A_83_260#_c_89_n N_VPWR_c_419_n 0.00866457f $X=0.505 $Y=1.765 $X2=0
+ $Y2=0
cc_121 N_A_83_260#_c_100_p N_VPWR_c_419_n 0.0277606f $X=1.41 $Y=2.395 $X2=0
+ $Y2=0
cc_122 N_A_83_260#_c_126_p N_VPWR_c_419_n 0.0148861f $X=0.855 $Y=2.395 $X2=0
+ $Y2=0
cc_123 N_A_83_260#_c_96_n N_VPWR_c_419_n 0.0105551f $X=1.575 $Y=2.395 $X2=0
+ $Y2=0
cc_124 N_A_83_260#_c_89_n N_VPWR_c_424_n 0.00445602f $X=0.505 $Y=1.765 $X2=0
+ $Y2=0
cc_125 N_A_83_260#_c_96_n N_VPWR_c_425_n 0.00707049f $X=1.575 $Y=2.395 $X2=0
+ $Y2=0
cc_126 N_A_83_260#_c_89_n N_VPWR_c_418_n 0.00865213f $X=0.505 $Y=1.765 $X2=0
+ $Y2=0
cc_127 N_A_83_260#_c_100_p N_VPWR_c_418_n 0.00770325f $X=1.41 $Y=2.395 $X2=0
+ $Y2=0
cc_128 N_A_83_260#_c_126_p N_VPWR_c_418_n 6.0606e-19 $X=0.855 $Y=2.395 $X2=0
+ $Y2=0
cc_129 N_A_83_260#_c_96_n N_VPWR_c_418_n 0.0105792f $X=1.575 $Y=2.395 $X2=0
+ $Y2=0
cc_130 N_A_83_260#_M1012_g N_VGND_c_504_n 0.0065091f $X=0.495 $Y=0.74 $X2=0
+ $Y2=0
cc_131 N_A_83_260#_c_89_n N_VGND_c_504_n 0.00129532f $X=0.505 $Y=1.765 $X2=0
+ $Y2=0
cc_132 N_A_83_260#_c_90_n N_VGND_c_504_n 0.0117358f $X=0.77 $Y=1.63 $X2=0 $Y2=0
cc_133 N_A_83_260#_c_92_n N_VGND_c_504_n 9.77913e-19 $X=1.07 $Y=1.215 $X2=0
+ $Y2=0
cc_134 N_A_83_260#_M1012_g N_VGND_c_509_n 0.00434272f $X=0.495 $Y=0.74 $X2=0
+ $Y2=0
cc_135 N_A_83_260#_M1012_g N_VGND_c_512_n 0.00828941f $X=0.495 $Y=0.74 $X2=0
+ $Y2=0
cc_136 N_A_83_260#_c_93_n N_A_305_130#_c_561_n 0.00652315f $X=1.235 $Y=1.105
+ $X2=0 $Y2=0
cc_137 N_A_239_294#_c_147_n N_B_c_259_n 0.0480285f $X=1.35 $Y=1.885 $X2=-0.19
+ $Y2=-0.245
cc_138 N_A_239_294#_c_151_n N_B_c_259_n 0.00415077f $X=1.36 $Y=1.635 $X2=-0.19
+ $Y2=-0.245
cc_139 N_A_239_294#_c_158_n N_B_c_259_n 0.0193896f $X=3.36 $Y=2.055 $X2=-0.19
+ $Y2=-0.245
cc_140 N_A_239_294#_M1009_g N_B_M1010_g 0.0147051f $X=1.45 $Y=0.97 $X2=0 $Y2=0
cc_141 N_A_239_294#_c_158_n N_B_c_268_n 0.0179661f $X=3.36 $Y=2.055 $X2=0 $Y2=0
cc_142 N_A_239_294#_c_159_n N_B_c_268_n 9.00673e-19 $X=3.475 $Y=2.265 $X2=0
+ $Y2=0
cc_143 N_A_239_294#_c_152_n N_B_M1001_g 0.0087538f $X=3.185 $Y=0.74 $X2=0 $Y2=0
cc_144 N_A_239_294#_c_153_n N_B_M1001_g 0.0260005f $X=3.64 $Y=1.515 $X2=0 $Y2=0
cc_145 N_A_239_294#_c_147_n N_B_c_262_n 0.00120624f $X=1.35 $Y=1.885 $X2=0 $Y2=0
cc_146 N_A_239_294#_c_151_n N_B_c_262_n 0.0195858f $X=1.36 $Y=1.635 $X2=0 $Y2=0
cc_147 N_A_239_294#_c_158_n N_B_c_262_n 0.10735f $X=3.36 $Y=2.055 $X2=0 $Y2=0
cc_148 N_A_239_294#_c_160_n B 0.00947173f $X=3.555 $Y=1.97 $X2=0 $Y2=0
cc_149 N_A_239_294#_c_153_n B 0.0374191f $X=3.64 $Y=1.515 $X2=0 $Y2=0
cc_150 N_A_239_294#_c_158_n N_B_c_264_n 0.00493107f $X=3.36 $Y=2.055 $X2=0 $Y2=0
cc_151 N_A_239_294#_c_160_n N_B_c_264_n 0.00466205f $X=3.555 $Y=1.97 $X2=0 $Y2=0
cc_152 N_A_239_294#_c_153_n N_B_c_264_n 0.0122493f $X=3.64 $Y=1.515 $X2=0 $Y2=0
cc_153 N_A_239_294#_c_162_n N_B_c_264_n 0.00439489f $X=3.5 $Y=2.055 $X2=0 $Y2=0
cc_154 N_A_239_294#_c_152_n N_A_M1013_g 0.00519877f $X=3.185 $Y=0.74 $X2=0 $Y2=0
cc_155 N_A_239_294#_c_158_n N_A_c_332_n 0.0166792f $X=3.36 $Y=2.055 $X2=0 $Y2=0
cc_156 N_A_239_294#_c_152_n N_A_c_327_n 0.00622038f $X=3.185 $Y=0.74 $X2=0 $Y2=0
cc_157 N_A_239_294#_c_149_n N_A_c_333_n 0.0217546f $X=4.25 $Y=1.765 $X2=0 $Y2=0
cc_158 N_A_239_294#_c_159_n N_A_c_333_n 0.0100476f $X=3.475 $Y=2.265 $X2=0 $Y2=0
cc_159 N_A_239_294#_c_162_n N_A_c_333_n 0.00235472f $X=3.5 $Y=2.055 $X2=0 $Y2=0
cc_160 N_A_239_294#_c_149_n N_A_c_334_n 9.94165e-19 $X=4.25 $Y=1.765 $X2=0 $Y2=0
cc_161 N_A_239_294#_c_160_n N_A_c_334_n 0.00389188f $X=3.555 $Y=1.97 $X2=0 $Y2=0
cc_162 N_A_239_294#_c_154_n N_A_c_334_n 0.00195502f $X=4.21 $Y=1.515 $X2=0 $Y2=0
cc_163 N_A_239_294#_c_162_n N_A_c_334_n 0.00285756f $X=3.5 $Y=2.055 $X2=0 $Y2=0
cc_164 N_A_239_294#_c_149_n N_A_M1011_g 0.0333546f $X=4.25 $Y=1.765 $X2=0 $Y2=0
cc_165 N_A_239_294#_c_150_n N_A_M1011_g 0.0192035f $X=4.26 $Y=1.35 $X2=0 $Y2=0
cc_166 N_A_239_294#_c_152_n N_A_M1011_g 0.00138729f $X=3.185 $Y=0.74 $X2=0 $Y2=0
cc_167 N_A_239_294#_c_160_n N_A_M1011_g 0.00437042f $X=3.555 $Y=1.97 $X2=0 $Y2=0
cc_168 N_A_239_294#_c_153_n N_A_M1011_g 0.00328653f $X=3.64 $Y=1.515 $X2=0 $Y2=0
cc_169 N_A_239_294#_c_154_n N_A_M1011_g 0.0232629f $X=4.21 $Y=1.515 $X2=0 $Y2=0
cc_170 N_A_239_294#_c_152_n N_A_c_330_n 0.00617654f $X=3.185 $Y=0.74 $X2=0 $Y2=0
cc_171 N_A_239_294#_c_178_n N_VPWR_M1006_d 0.00259449f $X=1.525 $Y=2.055
+ $X2=-0.19 $Y2=-0.245
cc_172 N_A_239_294#_c_158_n N_VPWR_M1008_d 0.00918987f $X=3.36 $Y=2.055 $X2=0
+ $Y2=0
cc_173 N_A_239_294#_c_147_n N_VPWR_c_419_n 0.00637936f $X=1.35 $Y=1.885 $X2=0
+ $Y2=0
cc_174 N_A_239_294#_c_158_n N_VPWR_c_420_n 0.0476908f $X=3.36 $Y=2.055 $X2=0
+ $Y2=0
cc_175 N_A_239_294#_c_159_n N_VPWR_c_420_n 0.0290034f $X=3.475 $Y=2.265 $X2=0
+ $Y2=0
cc_176 N_A_239_294#_c_149_n N_VPWR_c_421_n 0.010284f $X=4.25 $Y=1.765 $X2=0
+ $Y2=0
cc_177 N_A_239_294#_c_159_n N_VPWR_c_421_n 0.0314893f $X=3.475 $Y=2.265 $X2=0
+ $Y2=0
cc_178 N_A_239_294#_c_154_n N_VPWR_c_421_n 0.0140709f $X=4.21 $Y=1.515 $X2=0
+ $Y2=0
cc_179 N_A_239_294#_c_162_n N_VPWR_c_421_n 0.00247877f $X=3.5 $Y=2.055 $X2=0
+ $Y2=0
cc_180 N_A_239_294#_c_159_n N_VPWR_c_422_n 0.0123628f $X=3.475 $Y=2.265 $X2=0
+ $Y2=0
cc_181 N_A_239_294#_c_147_n N_VPWR_c_425_n 0.00458182f $X=1.35 $Y=1.885 $X2=0
+ $Y2=0
cc_182 N_A_239_294#_c_149_n N_VPWR_c_426_n 0.00445602f $X=4.25 $Y=1.765 $X2=0
+ $Y2=0
cc_183 N_A_239_294#_c_147_n N_VPWR_c_418_n 0.0049649f $X=1.35 $Y=1.885 $X2=0
+ $Y2=0
cc_184 N_A_239_294#_c_149_n N_VPWR_c_418_n 0.00861459f $X=4.25 $Y=1.765 $X2=0
+ $Y2=0
cc_185 N_A_239_294#_c_159_n N_VPWR_c_418_n 0.0101999f $X=3.475 $Y=2.265 $X2=0
+ $Y2=0
cc_186 N_A_239_294#_c_158_n A_386_392# 0.0152207f $X=3.36 $Y=2.055 $X2=-0.19
+ $Y2=-0.245
cc_187 N_A_239_294#_c_150_n N_COUT_c_480_n 0.0058436f $X=4.26 $Y=1.35 $X2=0
+ $Y2=0
cc_188 N_A_239_294#_c_150_n N_COUT_c_481_n 0.00239802f $X=4.26 $Y=1.35 $X2=0
+ $Y2=0
cc_189 N_A_239_294#_c_154_n N_COUT_c_481_n 0.00338703f $X=4.21 $Y=1.515 $X2=0
+ $Y2=0
cc_190 N_A_239_294#_c_149_n COUT 0.014428f $X=4.25 $Y=1.765 $X2=0 $Y2=0
cc_191 N_A_239_294#_c_160_n COUT 0.00278963f $X=3.555 $Y=1.97 $X2=0 $Y2=0
cc_192 N_A_239_294#_c_154_n COUT 0.00296045f $X=4.21 $Y=1.515 $X2=0 $Y2=0
cc_193 N_A_239_294#_c_162_n COUT 0.00330848f $X=3.5 $Y=2.055 $X2=0 $Y2=0
cc_194 N_A_239_294#_c_149_n N_COUT_c_482_n 0.00629291f $X=4.25 $Y=1.765 $X2=0
+ $Y2=0
cc_195 N_A_239_294#_c_150_n N_COUT_c_482_n 0.00391901f $X=4.26 $Y=1.35 $X2=0
+ $Y2=0
cc_196 N_A_239_294#_c_154_n N_COUT_c_482_n 0.0262124f $X=4.21 $Y=1.515 $X2=0
+ $Y2=0
cc_197 N_A_239_294#_M1009_g N_VGND_c_504_n 0.0069746f $X=1.45 $Y=0.97 $X2=0
+ $Y2=0
cc_198 N_A_239_294#_M1009_g N_VGND_c_505_n 6.34279e-19 $X=1.45 $Y=0.97 $X2=0
+ $Y2=0
cc_199 N_A_239_294#_c_149_n N_VGND_c_506_n 0.00215627f $X=4.25 $Y=1.765 $X2=0
+ $Y2=0
cc_200 N_A_239_294#_c_150_n N_VGND_c_506_n 0.00685808f $X=4.26 $Y=1.35 $X2=0
+ $Y2=0
cc_201 N_A_239_294#_c_152_n N_VGND_c_506_n 0.0170465f $X=3.185 $Y=0.74 $X2=0
+ $Y2=0
cc_202 N_A_239_294#_c_154_n N_VGND_c_506_n 0.0247894f $X=4.21 $Y=1.515 $X2=0
+ $Y2=0
cc_203 N_A_239_294#_c_152_n N_VGND_c_507_n 0.00749462f $X=3.185 $Y=0.74 $X2=0
+ $Y2=0
cc_204 N_A_239_294#_M1009_g N_VGND_c_510_n 0.00402388f $X=1.45 $Y=0.97 $X2=0
+ $Y2=0
cc_205 N_A_239_294#_c_150_n N_VGND_c_511_n 0.00470409f $X=4.26 $Y=1.35 $X2=0
+ $Y2=0
cc_206 N_A_239_294#_M1009_g N_VGND_c_512_n 0.00462577f $X=1.45 $Y=0.97 $X2=0
+ $Y2=0
cc_207 N_A_239_294#_c_150_n N_VGND_c_512_n 0.00506877f $X=4.26 $Y=1.35 $X2=0
+ $Y2=0
cc_208 N_A_239_294#_c_152_n N_VGND_c_512_n 0.00907254f $X=3.185 $Y=0.74 $X2=0
+ $Y2=0
cc_209 N_A_239_294#_M1009_g N_A_305_130#_c_559_n 4.5765e-19 $X=1.45 $Y=0.97
+ $X2=0 $Y2=0
cc_210 N_A_239_294#_c_158_n N_A_305_130#_c_561_n 0.00487746f $X=3.36 $Y=2.055
+ $X2=0 $Y2=0
cc_211 N_A_239_294#_c_152_n N_A_305_130#_c_562_n 0.0164838f $X=3.185 $Y=0.74
+ $X2=0 $Y2=0
cc_212 N_A_239_294#_c_153_n N_A_305_130#_c_562_n 0.0120732f $X=3.64 $Y=1.515
+ $X2=0 $Y2=0
cc_213 N_A_239_294#_c_153_n A_695_119# 0.00433061f $X=3.64 $Y=1.515 $X2=-0.19
+ $Y2=-0.245
cc_214 N_B_c_259_n N_A_c_325_n 0.0177686f $X=1.855 $Y=1.885 $X2=0 $Y2=0
cc_215 N_B_c_262_n N_A_c_325_n 5.18945e-19 $X=2.095 $Y=1.635 $X2=0 $Y2=0
cc_216 B N_A_c_325_n 4.44378e-19 $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_217 N_B_c_264_n N_A_c_325_n 0.00747088f $X=3.25 $Y=1.635 $X2=0 $Y2=0
cc_218 N_B_c_265_n N_A_c_326_n 0.0134311f $X=2.97 $Y=1.635 $X2=0 $Y2=0
cc_219 N_B_c_259_n N_A_c_332_n 0.037895f $X=1.855 $Y=1.885 $X2=0 $Y2=0
cc_220 N_B_c_267_n N_A_c_332_n 0.00484081f $X=3.25 $Y=1.955 $X2=0 $Y2=0
cc_221 N_B_c_268_n N_A_c_332_n 0.00403015f $X=3.25 $Y=2.045 $X2=0 $Y2=0
cc_222 N_B_c_265_n N_A_c_332_n 0.00237826f $X=2.97 $Y=1.635 $X2=0 $Y2=0
cc_223 N_B_M1001_g N_A_c_327_n 0.0103003f $X=3.4 $Y=0.915 $X2=0 $Y2=0
cc_224 N_B_c_268_n N_A_c_333_n 0.0138118f $X=3.25 $Y=2.045 $X2=0 $Y2=0
cc_225 N_B_c_267_n N_A_c_334_n 0.00825442f $X=3.25 $Y=1.955 $X2=0 $Y2=0
cc_226 N_B_M1001_g N_A_M1011_g 0.0684309f $X=3.4 $Y=0.915 $X2=0 $Y2=0
cc_227 N_B_c_264_n N_A_M1011_g 0.00683016f $X=3.25 $Y=1.635 $X2=0 $Y2=0
cc_228 N_B_M1010_g N_A_c_329_n 0.0227537f $X=1.88 $Y=0.97 $X2=0 $Y2=0
cc_229 N_B_M1001_g N_A_c_329_n 0.00289061f $X=3.4 $Y=0.915 $X2=0 $Y2=0
cc_230 N_B_M1001_g N_A_c_330_n 7.51436e-19 $X=3.4 $Y=0.915 $X2=0 $Y2=0
cc_231 N_B_c_259_n N_VPWR_c_419_n 0.00439808f $X=1.855 $Y=1.885 $X2=0 $Y2=0
cc_232 N_B_c_259_n N_VPWR_c_420_n 0.00348125f $X=1.855 $Y=1.885 $X2=0 $Y2=0
cc_233 N_B_c_268_n N_VPWR_c_420_n 0.0120472f $X=3.25 $Y=2.045 $X2=0 $Y2=0
cc_234 N_B_c_268_n N_VPWR_c_422_n 0.00413917f $X=3.25 $Y=2.045 $X2=0 $Y2=0
cc_235 N_B_c_259_n N_VPWR_c_425_n 0.00461464f $X=1.855 $Y=1.885 $X2=0 $Y2=0
cc_236 N_B_c_259_n N_VPWR_c_418_n 0.00915569f $X=1.855 $Y=1.885 $X2=0 $Y2=0
cc_237 N_B_c_268_n N_VPWR_c_418_n 0.0081781f $X=3.25 $Y=2.045 $X2=0 $Y2=0
cc_238 N_B_M1010_g N_VGND_c_505_n 0.00800137f $X=1.88 $Y=0.97 $X2=0 $Y2=0
cc_239 N_B_M1001_g N_VGND_c_506_n 0.00201272f $X=3.4 $Y=0.915 $X2=0 $Y2=0
cc_240 N_B_M1010_g N_VGND_c_510_n 0.00334468f $X=1.88 $Y=0.97 $X2=0 $Y2=0
cc_241 N_B_M1010_g N_VGND_c_512_n 0.00388565f $X=1.88 $Y=0.97 $X2=0 $Y2=0
cc_242 N_B_M1001_g N_VGND_c_512_n 9.39239e-19 $X=3.4 $Y=0.915 $X2=0 $Y2=0
cc_243 N_B_c_259_n N_A_305_130#_c_560_n 0.00415048f $X=1.855 $Y=1.885 $X2=0
+ $Y2=0
cc_244 N_B_M1010_g N_A_305_130#_c_560_n 0.0125952f $X=1.88 $Y=0.97 $X2=0 $Y2=0
cc_245 N_B_c_262_n N_A_305_130#_c_560_n 0.0242269f $X=2.095 $Y=1.635 $X2=0 $Y2=0
cc_246 N_B_c_265_n N_A_305_130#_c_560_n 0.0187108f $X=2.97 $Y=1.635 $X2=0 $Y2=0
cc_247 N_B_M1010_g N_A_305_130#_c_562_n 0.00106355f $X=1.88 $Y=0.97 $X2=0 $Y2=0
cc_248 N_B_M1001_g N_A_305_130#_c_562_n 0.00329625f $X=3.4 $Y=0.915 $X2=0 $Y2=0
cc_249 N_B_c_265_n N_A_305_130#_c_562_n 0.0249273f $X=2.97 $Y=1.635 $X2=0 $Y2=0
cc_250 N_A_c_332_n N_VPWR_c_420_n 0.0203642f $X=2.425 $Y=1.885 $X2=0 $Y2=0
cc_251 N_A_c_333_n N_VPWR_c_420_n 5.8387e-19 $X=3.7 $Y=2.045 $X2=0 $Y2=0
cc_252 N_A_c_333_n N_VPWR_c_421_n 0.00711687f $X=3.7 $Y=2.045 $X2=0 $Y2=0
cc_253 N_A_c_334_n N_VPWR_c_421_n 8.24724e-19 $X=3.76 $Y=1.86 $X2=0 $Y2=0
cc_254 N_A_c_333_n N_VPWR_c_422_n 0.00445602f $X=3.7 $Y=2.045 $X2=0 $Y2=0
cc_255 N_A_c_332_n N_VPWR_c_425_n 0.00413917f $X=2.425 $Y=1.885 $X2=0 $Y2=0
cc_256 N_A_c_332_n N_VPWR_c_418_n 0.00818781f $X=2.425 $Y=1.885 $X2=0 $Y2=0
cc_257 N_A_c_333_n N_VPWR_c_418_n 0.00857909f $X=3.7 $Y=2.045 $X2=0 $Y2=0
cc_258 N_A_M1011_g N_COUT_c_480_n 2.20852e-19 $X=3.76 $Y=0.915 $X2=0 $Y2=0
cc_259 N_A_c_333_n COUT 3.44411e-19 $X=3.7 $Y=2.045 $X2=0 $Y2=0
cc_260 N_A_M1011_g COUT 5.22968e-19 $X=3.76 $Y=0.915 $X2=0 $Y2=0
cc_261 N_A_c_329_n N_VGND_c_505_n 0.0167899f $X=2.557 $Y=0.18 $X2=0 $Y2=0
cc_262 N_A_c_330_n N_VGND_c_505_n 0.032955f $X=2.615 $Y=0.42 $X2=0 $Y2=0
cc_263 N_A_c_327_n N_VGND_c_506_n 0.00763335f $X=3.685 $Y=0.18 $X2=0 $Y2=0
cc_264 N_A_M1011_g N_VGND_c_506_n 0.0253391f $X=3.76 $Y=0.915 $X2=0 $Y2=0
cc_265 N_A_c_329_n N_VGND_c_507_n 0.0458086f $X=2.557 $Y=0.18 $X2=0 $Y2=0
cc_266 N_A_c_330_n N_VGND_c_507_n 0.0215843f $X=2.615 $Y=0.42 $X2=0 $Y2=0
cc_267 N_A_c_327_n N_VGND_c_512_n 0.0456613f $X=3.685 $Y=0.18 $X2=0 $Y2=0
cc_268 N_A_c_329_n N_VGND_c_512_n 0.017183f $X=2.557 $Y=0.18 $X2=0 $Y2=0
cc_269 N_A_c_330_n N_VGND_c_512_n 0.0110944f $X=2.615 $Y=0.42 $X2=0 $Y2=0
cc_270 N_A_M1013_g N_A_305_130#_c_560_n 0.0124342f $X=2.41 $Y=1.015 $X2=0 $Y2=0
cc_271 N_A_c_330_n N_A_305_130#_c_560_n 2.92673e-19 $X=2.615 $Y=0.42 $X2=0 $Y2=0
cc_272 N_A_M1013_g N_A_305_130#_c_562_n 0.0098681f $X=2.41 $Y=1.015 $X2=0 $Y2=0
cc_273 N_A_c_325_n N_A_305_130#_c_562_n 9.07186e-19 $X=2.425 $Y=1.5 $X2=0 $Y2=0
cc_274 N_A_c_329_n N_A_305_130#_c_562_n 0.00166975f $X=2.557 $Y=0.18 $X2=0 $Y2=0
cc_275 N_A_c_330_n N_A_305_130#_c_562_n 0.0244297f $X=2.615 $Y=0.42 $X2=0 $Y2=0
cc_276 SUM N_VPWR_c_419_n 0.0132454f $X=0.155 $Y=1.95 $X2=0 $Y2=0
cc_277 SUM N_VPWR_c_424_n 0.0145938f $X=0.155 $Y=1.95 $X2=0 $Y2=0
cc_278 SUM N_VPWR_c_418_n 0.0120466f $X=0.155 $Y=1.95 $X2=0 $Y2=0
cc_279 SUM N_VGND_c_504_n 0.0166774f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_280 SUM N_VGND_c_509_n 0.0145639f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_281 SUM N_VGND_c_512_n 0.0119984f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_282 N_VPWR_c_421_n COUT 0.0348613f $X=3.975 $Y=2.265 $X2=0 $Y2=0
cc_283 N_VPWR_c_426_n COUT 0.0179404f $X=4.56 $Y=3.33 $X2=0 $Y2=0
cc_284 N_VPWR_c_418_n COUT 0.0148166f $X=4.56 $Y=3.33 $X2=0 $Y2=0
cc_285 N_COUT_c_480_n N_VGND_c_506_n 0.0280471f $X=4.475 $Y=0.64 $X2=0 $Y2=0
cc_286 N_COUT_c_480_n N_VGND_c_511_n 0.0118732f $X=4.475 $Y=0.64 $X2=0 $Y2=0
cc_287 N_COUT_c_480_n N_VGND_c_512_n 0.0137068f $X=4.475 $Y=0.64 $X2=0 $Y2=0
cc_288 N_VGND_c_505_n N_A_305_130#_c_559_n 0.0126212f $X=2.105 $Y=0.795 $X2=0
+ $Y2=0
cc_289 N_VGND_c_510_n N_A_305_130#_c_559_n 0.00343395f $X=1.93 $Y=0 $X2=0 $Y2=0
cc_290 N_VGND_c_512_n N_A_305_130#_c_559_n 0.00511344f $X=4.56 $Y=0 $X2=0 $Y2=0
cc_291 N_VGND_M1010_d N_A_305_130#_c_560_n 0.00540456f $X=1.955 $Y=0.65 $X2=0
+ $Y2=0
cc_292 N_VGND_c_505_n N_A_305_130#_c_560_n 0.0234275f $X=2.105 $Y=0.795 $X2=0
+ $Y2=0
cc_293 N_VGND_c_512_n N_A_305_130#_c_562_n 8.74981e-19 $X=4.56 $Y=0 $X2=0 $Y2=0
