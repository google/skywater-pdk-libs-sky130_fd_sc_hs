* File: sky130_fd_sc_hs__decap_8.spice
* Created: Thu Aug 27 20:37:42 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hs__decap_8.pex.spice"
.subckt sky130_fd_sc_hs__decap_8  VNB VPB VGND VPWR
* 
* VPWR	VPWR
* VGND	VGND
* VPB	VPB
* VNB	VNB
MM1001 N_VGND_M1001_s N_VPWR_M1001_g N_VGND_M1001_s VNB NLOWVT L=1 W=0.42
+ AD=0.05775 AS=0.1113 PD=0.695 PS=1.37 NRD=0 NRS=0 M=1 R=0.42 SA=500000
+ SB=500001 A=0.42 P=2.84 MULT=1
MM1003 N_VGND_M1001_s N_VPWR_M1003_g N_VGND_M1001_s VNB NLOWVT L=1 W=0.42
+ AD=0.1197 AS=0.05775 PD=1.41 PS=0.695 NRD=0 NRS=0 M=1 R=0.42 SA=500001
+ SB=500000 A=0.42 P=2.84 MULT=1
MM1000 N_VPWR_M1000_s N_VGND_M1000_g N_VPWR_M1000_s VPB PSHORT L=1 W=1 AD=0.1375
+ AS=0.275 PD=1.275 PS=2.55 NRD=0 NRS=1.9503 M=1 R=1 SA=500000 SB=500001 A=1 P=4
+ MULT=1
MM1002 N_VPWR_M1000_s N_VGND_M1002_g N_VPWR_M1000_s VPB PSHORT L=1 W=1 AD=0.285
+ AS=0.1375 PD=2.57 PS=1.275 NRD=0 NRS=0 M=1 R=1 SA=500001 SB=500000 A=1 P=4
+ MULT=1
DX4_noxref VNB VPB NWDIODE A=7.8492 P=12.16
*
.include "sky130_fd_sc_hs__decap_8.pxi.spice"
*
.ends
*
*
