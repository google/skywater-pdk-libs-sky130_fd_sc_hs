* File: sky130_fd_sc_hs__o311a_4.spice
* Created: Thu Aug 27 21:01:56 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hs__o311a_4.pex.spice"
.subckt sky130_fd_sc_hs__o311a_4  VNB VPB B1 C1 A3 A2 A1 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A1	A1
* A2	A2
* A3	A3
* C1	C1
* B1	B1
* VPB	VPB
* VNB	VNB
MM1000 N_X_M1000_d N_A_83_244#_M1000_g N_VGND_M1000_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.2627 PD=1.02 PS=2.19 NRD=0 NRS=5.664 M=1 R=4.93333 SA=75000.3
+ SB=75001.8 A=0.111 P=1.78 MULT=1
MM1008 N_X_M1000_d N_A_83_244#_M1008_g N_VGND_M1008_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.20165 PD=1.02 PS=1.285 NRD=0 NRS=21.072 M=1 R=4.93333
+ SA=75000.7 SB=75001.4 A=0.111 P=1.78 MULT=1
MM1009 N_X_M1009_d N_A_83_244#_M1009_g N_VGND_M1008_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1295 AS=0.20165 PD=1.09 PS=1.285 NRD=0 NRS=21.888 M=1 R=4.93333
+ SA=75001.4 SB=75000.7 A=0.111 P=1.78 MULT=1
MM1025 N_X_M1009_d N_A_83_244#_M1025_g N_VGND_M1025_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1295 AS=0.2109 PD=1.09 PS=2.05 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75001.9
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1003 N_A_651_78#_M1003_d N_B1_M1003_g N_A_564_78#_M1003_s VNB NLOWVT L=0.15
+ W=0.64 AD=0.2544 AS=0.178025 PD=1.435 PS=1.85 NRD=13.116 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75005.2 A=0.096 P=1.58 MULT=1
MM1012 N_A_83_244#_M1012_d N_C1_M1012_g N_A_651_78#_M1003_d VNB NLOWVT L=0.15
+ W=0.64 AD=0.171975 AS=0.2544 PD=1.295 PS=1.435 NRD=40.068 NRS=0 M=1 R=4.26667
+ SA=75001.1 SB=75004.2 A=0.096 P=1.58 MULT=1
MM1022 N_A_83_244#_M1012_d N_C1_M1022_g N_A_651_78#_M1022_s VNB NLOWVT L=0.15
+ W=0.64 AD=0.171975 AS=0.0896 PD=1.295 PS=0.92 NRD=40.068 NRS=0 M=1 R=4.26667
+ SA=75001.7 SB=75003.6 A=0.096 P=1.58 MULT=1
MM1026 N_A_651_78#_M1022_s N_B1_M1026_g N_A_564_78#_M1026_s VNB NLOWVT L=0.15
+ W=0.64 AD=0.0896 AS=0.1216 PD=0.92 PS=1.02 NRD=0 NRS=13.116 M=1 R=4.26667
+ SA=75002.2 SB=75003.2 A=0.096 P=1.58 MULT=1
MM1018 N_A_564_78#_M1026_s N_A3_M1018_g N_VGND_M1018_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.1216 AS=0.1232 PD=1.02 PS=1.025 NRD=5.616 NRS=7.488 M=1 R=4.26667
+ SA=75002.7 SB=75002.7 A=0.096 P=1.58 MULT=1
MM1023 N_A_564_78#_M1023_d N_A3_M1023_g N_VGND_M1018_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.0912 AS=0.1232 PD=0.925 PS=1.025 NRD=0.936 NRS=12.18 M=1 R=4.26667
+ SA=75003.2 SB=75002.1 A=0.096 P=1.58 MULT=1
MM1010 N_A_564_78#_M1023_d N_A2_M1010_g N_VGND_M1010_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.0912 AS=0.12 PD=0.925 PS=1.015 NRD=0 NRS=13.116 M=1 R=4.26667 SA=75003.7
+ SB=75001.7 A=0.096 P=1.58 MULT=1
MM1001 N_A_564_78#_M1001_d N_A1_M1001_g N_VGND_M1010_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.1216 AS=0.12 PD=1.02 PS=1.015 NRD=8.436 NRS=4.68 M=1 R=4.26667 SA=75004.2
+ SB=75001.2 A=0.096 P=1.58 MULT=1
MM1027 N_A_564_78#_M1001_d N_A1_M1027_g N_VGND_M1027_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.1216 AS=0.0944 PD=1.02 PS=0.935 NRD=10.308 NRS=2.808 M=1 R=4.26667
+ SA=75004.7 SB=75000.7 A=0.096 P=1.58 MULT=1
MM1019 N_A_564_78#_M1019_d N_A2_M1019_g N_VGND_M1027_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.1824 AS=0.0944 PD=1.85 PS=0.935 NRD=0 NRS=0 M=1 R=4.26667 SA=75005.2
+ SB=75000.2 A=0.096 P=1.58 MULT=1
MM1013 N_VPWR_M1013_d N_A_83_244#_M1013_g N_X_M1013_s VPB PSHORT L=0.15 W=1.12
+ AD=0.3304 AS=0.168 PD=2.83 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75004 A=0.168 P=2.54 MULT=1
MM1014 N_VPWR_M1014_d N_A_83_244#_M1014_g N_X_M1013_s VPB PSHORT L=0.15 W=1.12
+ AD=0.196 AS=0.168 PD=1.47 PS=1.42 NRD=10.5395 NRS=1.7533 M=1 R=7.46667
+ SA=75000.7 SB=75003.5 A=0.168 P=2.54 MULT=1
MM1016 N_VPWR_M1014_d N_A_83_244#_M1016_g N_X_M1016_s VPB PSHORT L=0.15 W=1.12
+ AD=0.196 AS=0.2716 PD=1.47 PS=1.605 NRD=1.7533 NRS=10.5395 M=1 R=7.46667
+ SA=75001.2 SB=75003 A=0.168 P=2.54 MULT=1
MM1024 N_VPWR_M1024_d N_A_83_244#_M1024_g N_X_M1016_s VPB PSHORT L=0.15 W=1.12
+ AD=0.204347 AS=0.2716 PD=1.55849 PS=1.605 NRD=1.7533 NRS=25.4918 M=1 R=7.46667
+ SA=75001.8 SB=75002.4 A=0.168 P=2.54 MULT=1
MM1002 N_VPWR_M1024_d N_B1_M1002_g N_A_83_244#_M1002_s VPB PSHORT L=0.15 W=1
+ AD=0.182453 AS=0.21 PD=1.39151 PS=1.42 NRD=12.7853 NRS=1.9503 M=1 R=6.66667
+ SA=75002.3 SB=75002.2 A=0.15 P=2.3 MULT=1
MM1004 N_A_83_244#_M1002_s N_C1_M1004_g N_VPWR_M1004_s VPB PSHORT L=0.15 W=1
+ AD=0.21 AS=0.3575 PD=1.42 PS=1.715 NRD=25.5903 NRS=1.9503 M=1 R=6.66667
+ SA=75002.9 SB=75001.6 A=0.15 P=2.3 MULT=1
MM1005 N_A_83_244#_M1005_d N_C1_M1005_g N_VPWR_M1004_s VPB PSHORT L=0.15 W=1
+ AD=0.175 AS=0.3575 PD=1.35 PS=1.715 NRD=1.9503 NRS=1.9503 M=1 R=6.66667
+ SA=75003.7 SB=75000.7 A=0.15 P=2.3 MULT=1
MM1006 N_VPWR_M1006_d N_B1_M1006_g N_A_83_244#_M1005_d VPB PSHORT L=0.15 W=1
+ AD=0.295 AS=0.175 PD=2.59 PS=1.35 NRD=1.9503 NRS=11.8003 M=1 R=6.66667
+ SA=75004.2 SB=75000.2 A=0.15 P=2.3 MULT=1
MM1011 N_A_83_244#_M1011_d N_A3_M1011_g N_A_1034_392#_M1011_s VPB PSHORT L=0.15
+ W=1 AD=0.16 AS=0.445 PD=1.32 PS=2.89 NRD=3.9203 NRS=16.7253 M=1 R=6.66667
+ SA=75000.4 SB=75002.7 A=0.15 P=2.3 MULT=1
MM1015 N_A_83_244#_M1011_d N_A3_M1015_g N_A_1034_392#_M1015_s VPB PSHORT L=0.15
+ W=1 AD=0.16 AS=0.1525 PD=1.32 PS=1.305 NRD=3.9203 NRS=1.9503 M=1 R=6.66667
+ SA=75000.8 SB=75002.2 A=0.15 P=2.3 MULT=1
MM1007 N_A_1338_392#_M1007_d N_A2_M1007_g N_A_1034_392#_M1015_s VPB PSHORT
+ L=0.15 W=1 AD=0.21 AS=0.1525 PD=1.42 PS=1.305 NRD=17.73 NRS=2.9353 M=1
+ R=6.66667 SA=75001.3 SB=75001.7 A=0.15 P=2.3 MULT=1
MM1017 N_VPWR_M1017_d N_A1_M1017_g N_A_1338_392#_M1007_d VPB PSHORT L=0.15 W=1
+ AD=0.15 AS=0.21 PD=1.3 PS=1.42 NRD=1.9503 NRS=9.8303 M=1 R=6.66667 SA=75001.9
+ SB=75001.2 A=0.15 P=2.3 MULT=1
MM1020 N_VPWR_M1017_d N_A1_M1020_g N_A_1338_392#_M1020_s VPB PSHORT L=0.15 W=1
+ AD=0.15 AS=0.16 PD=1.3 PS=1.32 NRD=1.9503 NRS=1.9503 M=1 R=6.66667 SA=75002.3
+ SB=75000.7 A=0.15 P=2.3 MULT=1
MM1021 N_A_1338_392#_M1020_s N_A2_M1021_g N_A_1034_392#_M1021_s VPB PSHORT
+ L=0.15 W=1 AD=0.16 AS=0.325 PD=1.32 PS=2.65 NRD=5.8903 NRS=7.8603 M=1
+ R=6.66667 SA=75002.8 SB=75000.2 A=0.15 P=2.3 MULT=1
DX28_noxref VNB VPB NWDIODE A=16.7772 P=21.76
*
.include "sky130_fd_sc_hs__o311a_4.pxi.spice"
*
.ends
*
*
