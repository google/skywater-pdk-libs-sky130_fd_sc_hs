* NGSPICE file created from sky130_fd_sc_hs__a2bb2o_1.ext - technology: sky130A

.subckt sky130_fd_sc_hs__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
M1000 a_530_392# B1 VPWR VPB pshort w=1e+06u l=150000u
+  ad=5.75e+11p pd=5.15e+06u as=7.28e+11p ps=5.63e+06u
M1001 a_93_264# a_257_126# VGND VNB nlowvt w=640000u l=150000u
+  ad=1.792e+11p pd=1.84e+06u as=8.3095e+11p ps=6.71e+06u
M1002 VPWR a_93_264# X VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=3.08e+11p ps=2.79e+06u
M1003 a_258_392# A1_N VPWR VPB pshort w=1e+06u l=150000u
+  ad=2.4e+11p pd=2.48e+06u as=0p ps=0u
M1004 a_605_126# B2 a_93_264# VNB nlowvt w=640000u l=150000u
+  ad=2.496e+11p pd=2.06e+06u as=0p ps=0u
M1005 a_530_392# a_257_126# a_93_264# VPB pshort w=1e+06u l=150000u
+  ad=0p pd=0u as=2.75e+11p ps=2.55e+06u
M1006 a_257_126# A1_N VGND VNB nlowvt w=550000u l=150000u
+  ad=1.54e+11p pd=1.66e+06u as=0p ps=0u
M1007 VGND A2_N a_257_126# VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VGND a_93_264# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=1.961e+11p ps=2.01e+06u
M1009 VPWR B2 a_530_392# VPB pshort w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VGND B1 a_605_126# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_257_126# A2_N a_258_392# VPB pshort w=1e+06u l=150000u
+  ad=2.75e+11p pd=2.55e+06u as=0p ps=0u
.ends

