* File: sky130_fd_sc_hs__a32oi_1.spice
* Created: Thu Aug 27 20:30:18 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hs__a32oi_1.pex.spice"
.subckt sky130_fd_sc_hs__a32oi_1  VNB VPB B2 B1 A1 A2 A3 Y VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* Y	Y
* A3	A3
* A2	A2
* A1	A1
* B1	B1
* B2	B2
* VPB	VPB
* VNB	VNB
MM1002 A_119_74# N_B2_M1002_g N_VGND_M1002_s VNB NLOWVT L=0.15 W=0.74 AD=0.0888
+ AS=0.2294 PD=0.98 PS=2.1 NRD=10.536 NRS=4.044 M=1 R=4.93333 SA=75000.2
+ SB=75002.5 A=0.111 P=1.78 MULT=1
MM1000 N_Y_M1000_d N_B1_M1000_g A_119_74# VNB NLOWVT L=0.15 W=0.74 AD=0.3034
+ AS=0.0888 PD=1.56 PS=0.98 NRD=0 NRS=10.536 M=1 R=4.93333 SA=75000.6 SB=75002.1
+ A=0.111 P=1.78 MULT=1
MM1006 A_391_74# N_A1_M1006_g N_Y_M1000_d VNB NLOWVT L=0.15 W=0.74 AD=0.0888
+ AS=0.3034 PD=0.98 PS=1.56 NRD=10.536 NRS=0 M=1 R=4.93333 SA=75001.6 SB=75001.2
+ A=0.111 P=1.78 MULT=1
MM1009 A_469_74# N_A2_M1009_g A_391_74# VNB NLOWVT L=0.15 W=0.74 AD=0.1554
+ AS=0.0888 PD=1.16 PS=0.98 NRD=25.128 NRS=10.536 M=1 R=4.93333 SA=75002
+ SB=75000.8 A=0.111 P=1.78 MULT=1
MM1001 N_VGND_M1001_d N_A3_M1001_g A_469_74# VNB NLOWVT L=0.15 W=0.74 AD=0.2109
+ AS=0.1554 PD=2.05 PS=1.16 NRD=0 NRS=25.128 M=1 R=4.93333 SA=75002.6 SB=75000.2
+ A=0.111 P=1.78 MULT=1
MM1004 N_Y_M1004_d N_B2_M1004_g N_A_27_368#_M1004_s VPB PSHORT L=0.15 W=1.12
+ AD=0.196 AS=0.3304 PD=1.47 PS=2.83 NRD=10.5395 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75002.6 A=0.168 P=2.54 MULT=1
MM1003 N_A_27_368#_M1003_d N_B1_M1003_g N_Y_M1004_d VPB PSHORT L=0.15 W=1.12
+ AD=0.2576 AS=0.196 PD=1.58 PS=1.47 NRD=10.5395 NRS=1.7533 M=1 R=7.46667
+ SA=75000.7 SB=75002.1 A=0.168 P=2.54 MULT=1
MM1008 N_VPWR_M1008_d N_A1_M1008_g N_A_27_368#_M1003_d VPB PSHORT L=0.15 W=1.12
+ AD=0.3584 AS=0.2576 PD=1.76 PS=1.58 NRD=1.7533 NRS=21.0987 M=1 R=7.46667
+ SA=75001.3 SB=75001.5 A=0.168 P=2.54 MULT=1
MM1005 N_A_27_368#_M1005_d N_A2_M1005_g N_VPWR_M1008_d VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.3584 PD=1.42 PS=1.76 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75002.1 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1007 N_VPWR_M1007_d N_A3_M1007_g N_A_27_368#_M1005_d VPB PSHORT L=0.15 W=1.12
+ AD=0.3304 AS=0.168 PD=2.83 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75002.6 SB=75000.2 A=0.168 P=2.54 MULT=1
DX10_noxref VNB VPB NWDIODE A=6.9564 P=11.2
c_351 A_119_74# 0 1.22712e-19 $X=0.595 $Y=0.37
*
.include "sky130_fd_sc_hs__a32oi_1.pxi.spice"
*
.ends
*
*
