* File: sky130_fd_sc_hs__or4b_2.pxi.spice
* Created: Thu Aug 27 21:07:12 2020
* 
x_PM_SKY130_FD_SC_HS__OR4B_2%D_N N_D_N_c_80_n N_D_N_M1006_g N_D_N_M1010_g D_N
+ N_D_N_c_82_n PM_SKY130_FD_SC_HS__OR4B_2%D_N
x_PM_SKY130_FD_SC_HS__OR4B_2%A_190_48# N_A_190_48#_M1004_d N_A_190_48#_M1002_d
+ N_A_190_48#_M1008_d N_A_190_48#_M1005_g N_A_190_48#_c_107_n
+ N_A_190_48#_c_123_n N_A_190_48#_M1000_g N_A_190_48#_c_108_n
+ N_A_190_48#_M1013_g N_A_190_48#_c_110_n N_A_190_48#_M1001_g
+ N_A_190_48#_c_111_n N_A_190_48#_c_112_n N_A_190_48#_c_113_n
+ N_A_190_48#_c_190_p N_A_190_48#_c_114_n N_A_190_48#_c_115_n
+ N_A_190_48#_c_116_n N_A_190_48#_c_125_n N_A_190_48#_c_117_n
+ N_A_190_48#_c_118_n N_A_190_48#_c_119_n N_A_190_48#_c_120_n
+ N_A_190_48#_c_126_n N_A_190_48#_c_121_n PM_SKY130_FD_SC_HS__OR4B_2%A_190_48#
x_PM_SKY130_FD_SC_HS__OR4B_2%A N_A_M1004_g N_A_c_228_n N_A_M1007_g A A
+ N_A_c_229_n PM_SKY130_FD_SC_HS__OR4B_2%A
x_PM_SKY130_FD_SC_HS__OR4B_2%B N_B_c_266_n N_B_M1012_g N_B_M1009_g B B
+ PM_SKY130_FD_SC_HS__OR4B_2%B
x_PM_SKY130_FD_SC_HS__OR4B_2%C N_C_c_300_n N_C_M1003_g N_C_M1002_g C C C
+ PM_SKY130_FD_SC_HS__OR4B_2%C
x_PM_SKY130_FD_SC_HS__OR4B_2%A_27_368# N_A_27_368#_M1010_s N_A_27_368#_M1006_s
+ N_A_27_368#_c_330_n N_A_27_368#_M1008_g N_A_27_368#_M1011_g
+ N_A_27_368#_c_332_n N_A_27_368#_c_333_n N_A_27_368#_c_334_n
+ N_A_27_368#_c_335_n N_A_27_368#_c_365_n N_A_27_368#_c_339_n
+ N_A_27_368#_c_377_n N_A_27_368#_c_368_n N_A_27_368#_c_398_p
+ N_A_27_368#_c_340_n N_A_27_368#_c_336_n PM_SKY130_FD_SC_HS__OR4B_2%A_27_368#
x_PM_SKY130_FD_SC_HS__OR4B_2%VPWR N_VPWR_M1006_d N_VPWR_M1001_s N_VPWR_c_427_n
+ VPWR N_VPWR_c_428_n N_VPWR_c_429_n N_VPWR_c_426_n N_VPWR_c_431_n
+ N_VPWR_c_432_n PM_SKY130_FD_SC_HS__OR4B_2%VPWR
x_PM_SKY130_FD_SC_HS__OR4B_2%X N_X_M1005_d N_X_M1000_d N_X_c_471_n N_X_c_472_n X
+ N_X_c_473_n PM_SKY130_FD_SC_HS__OR4B_2%X
x_PM_SKY130_FD_SC_HS__OR4B_2%VGND N_VGND_M1010_d N_VGND_M1013_s N_VGND_M1009_d
+ N_VGND_M1011_d N_VGND_c_517_n N_VGND_c_518_n N_VGND_c_519_n N_VGND_c_520_n
+ N_VGND_c_521_n VGND N_VGND_c_522_n N_VGND_c_523_n N_VGND_c_524_n
+ N_VGND_c_525_n N_VGND_c_526_n N_VGND_c_527_n N_VGND_c_528_n
+ PM_SKY130_FD_SC_HS__OR4B_2%VGND
cc_1 VNB N_D_N_c_80_n 0.0339337f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.765
cc_2 VNB N_D_N_M1010_g 0.0335586f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=0.835
cc_3 VNB N_D_N_c_82_n 0.0147527f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.515
cc_4 VNB N_A_190_48#_M1005_g 0.0217322f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.515
cc_5 VNB N_A_190_48#_c_107_n 0.0110629f $X=-0.19 $Y=-0.245 $X2=0.337 $Y2=1.665
cc_6 VNB N_A_190_48#_c_108_n 0.0134199f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_7 VNB N_A_190_48#_M1013_g 0.0229022f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_A_190_48#_c_110_n 0.0328645f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A_190_48#_c_111_n 0.00626877f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_190_48#_c_112_n 0.00305584f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_190_48#_c_113_n 0.00740858f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_190_48#_c_114_n 0.00379109f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_190_48#_c_115_n 0.00326291f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_190_48#_c_116_n 0.0126446f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_190_48#_c_117_n 0.00293951f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_190_48#_c_118_n 0.00951601f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_190_48#_c_119_n 0.0103969f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_190_48#_c_120_n 0.00809499f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_190_48#_c_121_n 0.0186681f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_M1004_g 0.0266404f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.26
cc_21 VNB N_A_c_228_n 0.0268397f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=0.835
cc_22 VNB N_A_c_229_n 0.00183238f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_B_c_266_n 0.0180474f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.765
cc_24 VNB N_B_M1009_g 0.0350429f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=0.835
cc_25 VNB B 0.00220385f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_26 VNB N_C_c_300_n 0.0168465f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.765
cc_27 VNB N_C_M1002_g 0.0343028f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=0.835
cc_28 VNB C 0.00367115f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_29 VNB N_A_27_368#_c_330_n 0.020756f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_27_368#_M1011_g 0.0311486f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.515
cc_31 VNB N_A_27_368#_c_332_n 0.0214174f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_27_368#_c_333_n 0.00531827f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_27_368#_c_334_n 0.00942464f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_27_368#_c_335_n 0.0086419f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_27_368#_c_336_n 0.00386761f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_VPWR_c_426_n 0.183584f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_X_c_471_n 0.00240191f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_X_c_472_n 0.00434772f $X=-0.19 $Y=-0.245 $X2=0.337 $Y2=1.515
cc_39 VNB N_X_c_473_n 0.00226257f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_517_n 0.0157056f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_518_n 0.0117064f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_519_n 0.0147881f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_520_n 0.0122168f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_521_n 0.0366542f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_VGND_c_522_n 0.0190549f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_VGND_c_523_n 0.0197882f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_VGND_c_524_n 0.0191517f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_VGND_c_525_n 0.0255552f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_VGND_c_526_n 0.0080786f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_VGND_c_527_n 0.0100021f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_VGND_c_528_n 0.265964f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VPB N_D_N_c_80_n 0.0352417f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.765
cc_53 VPB N_D_N_c_82_n 0.00743971f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.515
cc_54 VPB N_A_190_48#_c_107_n 7.52477e-19 $X=-0.19 $Y=1.66 $X2=0.337 $Y2=1.665
cc_55 VPB N_A_190_48#_c_123_n 0.0226643f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_56 VPB N_A_190_48#_c_110_n 0.0238332f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_57 VPB N_A_190_48#_c_125_n 0.0377253f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_58 VPB N_A_190_48#_c_126_n 0.0104317f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_59 VPB N_A_190_48#_c_121_n 0.0133271f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_60 VPB N_A_c_228_n 0.0340501f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=0.835
cc_61 VPB N_A_c_229_n 0.00366723f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_62 VPB N_B_c_266_n 0.0342672f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.765
cc_63 VPB B 0.00208534f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_64 VPB N_C_c_300_n 0.0346567f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.765
cc_65 VPB C 0.0029668f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_66 VPB N_A_27_368#_c_330_n 0.043269f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_67 VPB N_A_27_368#_c_335_n 0.00325164f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_68 VPB N_A_27_368#_c_339_n 0.0351409f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_69 VPB N_A_27_368#_c_340_n 0.00132971f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_70 VPB N_A_27_368#_c_336_n 0.00178662f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_71 VPB N_VPWR_c_427_n 0.0164215f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.515
cc_72 VPB N_VPWR_c_428_n 0.0177898f $X=-0.19 $Y=1.66 $X2=0.337 $Y2=1.665
cc_73 VPB N_VPWR_c_429_n 0.0603644f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_74 VPB N_VPWR_c_426_n 0.0720666f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_75 VPB N_VPWR_c_431_n 0.0274851f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_76 VPB N_VPWR_c_432_n 0.0159477f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_77 VPB X 0.00215253f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_78 VPB N_X_c_473_n 0.00105626f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_79 N_D_N_M1010_g N_A_190_48#_M1005_g 0.0151226f $X=0.51 $Y=0.835 $X2=0 $Y2=0
cc_80 N_D_N_c_80_n N_A_190_48#_c_107_n 0.0151226f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_81 N_D_N_c_80_n N_A_190_48#_c_123_n 0.0247093f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_82 N_D_N_M1010_g N_A_27_368#_c_332_n 0.00872945f $X=0.51 $Y=0.835 $X2=0 $Y2=0
cc_83 N_D_N_M1010_g N_A_27_368#_c_333_n 0.0120646f $X=0.51 $Y=0.835 $X2=0 $Y2=0
cc_84 N_D_N_c_82_n N_A_27_368#_c_333_n 0.00649299f $X=0.385 $Y=1.515 $X2=0 $Y2=0
cc_85 N_D_N_c_80_n N_A_27_368#_c_334_n 0.0016835f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_86 N_D_N_M1010_g N_A_27_368#_c_334_n 0.00377477f $X=0.51 $Y=0.835 $X2=0 $Y2=0
cc_87 N_D_N_c_82_n N_A_27_368#_c_334_n 0.0286137f $X=0.385 $Y=1.515 $X2=0 $Y2=0
cc_88 N_D_N_c_80_n N_A_27_368#_c_335_n 0.0039228f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_89 N_D_N_M1010_g N_A_27_368#_c_335_n 0.00700193f $X=0.51 $Y=0.835 $X2=0 $Y2=0
cc_90 N_D_N_c_82_n N_A_27_368#_c_335_n 0.0329136f $X=0.385 $Y=1.515 $X2=0 $Y2=0
cc_91 N_D_N_c_80_n N_A_27_368#_c_339_n 0.0274905f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_92 N_D_N_c_82_n N_A_27_368#_c_339_n 0.0339846f $X=0.385 $Y=1.515 $X2=0 $Y2=0
cc_93 N_D_N_c_80_n N_VPWR_c_427_n 0.00343137f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_94 N_D_N_c_80_n N_VPWR_c_426_n 0.00462577f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_95 N_D_N_c_80_n N_VPWR_c_431_n 0.00393265f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_96 N_D_N_M1010_g N_X_c_471_n 6.35749e-19 $X=0.51 $Y=0.835 $X2=0 $Y2=0
cc_97 N_D_N_M1010_g N_VGND_c_517_n 0.00459404f $X=0.51 $Y=0.835 $X2=0 $Y2=0
cc_98 N_D_N_M1010_g N_VGND_c_525_n 0.0043356f $X=0.51 $Y=0.835 $X2=0 $Y2=0
cc_99 N_D_N_M1010_g N_VGND_c_528_n 0.00487769f $X=0.51 $Y=0.835 $X2=0 $Y2=0
cc_100 N_A_190_48#_M1013_g N_A_M1004_g 0.0160656f $X=1.455 $Y=0.74 $X2=0 $Y2=0
cc_101 N_A_190_48#_c_110_n N_A_M1004_g 0.00252021f $X=1.49 $Y=1.765 $X2=0 $Y2=0
cc_102 N_A_190_48#_c_112_n N_A_M1004_g 0.00351998f $X=1.66 $Y=1.3 $X2=0 $Y2=0
cc_103 N_A_190_48#_c_113_n N_A_M1004_g 0.0156668f $X=2.175 $Y=1.045 $X2=0 $Y2=0
cc_104 N_A_190_48#_c_114_n N_A_M1004_g 0.00321875f $X=2.34 $Y=0.615 $X2=0 $Y2=0
cc_105 N_A_190_48#_c_117_n N_A_M1004_g 0.00107033f $X=1.66 $Y=1.465 $X2=0 $Y2=0
cc_106 N_A_190_48#_c_110_n N_A_c_228_n 0.0466218f $X=1.49 $Y=1.765 $X2=0 $Y2=0
cc_107 N_A_190_48#_c_113_n N_A_c_228_n 5.20343e-19 $X=2.175 $Y=1.045 $X2=0 $Y2=0
cc_108 N_A_190_48#_c_117_n N_A_c_228_n 0.00161664f $X=1.66 $Y=1.465 $X2=0 $Y2=0
cc_109 N_A_190_48#_c_118_n N_A_c_228_n 7.46984e-19 $X=2.34 $Y=1.045 $X2=0 $Y2=0
cc_110 N_A_190_48#_c_110_n N_A_c_229_n 0.00634756f $X=1.49 $Y=1.765 $X2=0 $Y2=0
cc_111 N_A_190_48#_c_113_n N_A_c_229_n 0.0144509f $X=2.175 $Y=1.045 $X2=0 $Y2=0
cc_112 N_A_190_48#_c_117_n N_A_c_229_n 0.0197025f $X=1.66 $Y=1.465 $X2=0 $Y2=0
cc_113 N_A_190_48#_c_118_n N_A_c_229_n 0.00726462f $X=2.34 $Y=1.045 $X2=0 $Y2=0
cc_114 N_A_190_48#_c_119_n N_B_c_266_n 9.60875e-19 $X=3.375 $Y=1.115 $X2=-0.19
+ $Y2=-0.245
cc_115 N_A_190_48#_c_114_n N_B_M1009_g 0.00321875f $X=2.34 $Y=0.615 $X2=0 $Y2=0
cc_116 N_A_190_48#_c_119_n N_B_M1009_g 0.016738f $X=3.375 $Y=1.115 $X2=0 $Y2=0
cc_117 N_A_190_48#_c_118_n B 0.00100747f $X=2.34 $Y=1.045 $X2=0 $Y2=0
cc_118 N_A_190_48#_c_119_n B 0.0140616f $X=3.375 $Y=1.115 $X2=0 $Y2=0
cc_119 N_A_190_48#_c_119_n N_C_c_300_n 0.00108395f $X=3.375 $Y=1.115 $X2=-0.19
+ $Y2=-0.245
cc_120 N_A_190_48#_c_119_n N_C_M1002_g 0.0148482f $X=3.375 $Y=1.115 $X2=0 $Y2=0
cc_121 N_A_190_48#_c_120_n N_C_M1002_g 0.00468012f $X=3.705 $Y=1.115 $X2=0 $Y2=0
cc_122 N_A_190_48#_c_119_n C 0.0160291f $X=3.375 $Y=1.115 $X2=0 $Y2=0
cc_123 N_A_190_48#_c_116_n N_A_27_368#_c_330_n 0.00145734f $X=4.065 $Y=1.185
+ $X2=0 $Y2=0
cc_124 N_A_190_48#_c_120_n N_A_27_368#_c_330_n 0.00303118f $X=3.705 $Y=1.115
+ $X2=0 $Y2=0
cc_125 N_A_190_48#_c_126_n N_A_27_368#_c_330_n 0.0240966f $X=4.03 $Y=2.105 $X2=0
+ $Y2=0
cc_126 N_A_190_48#_c_121_n N_A_27_368#_c_330_n 0.00536146f $X=4.05 $Y=1.94 $X2=0
+ $Y2=0
cc_127 N_A_190_48#_c_115_n N_A_27_368#_M1011_g 0.00700031f $X=3.54 $Y=0.615
+ $X2=0 $Y2=0
cc_128 N_A_190_48#_c_116_n N_A_27_368#_M1011_g 0.0127639f $X=4.065 $Y=1.185
+ $X2=0 $Y2=0
cc_129 N_A_190_48#_c_120_n N_A_27_368#_M1011_g 0.0092772f $X=3.705 $Y=1.115
+ $X2=0 $Y2=0
cc_130 N_A_190_48#_c_121_n N_A_27_368#_M1011_g 0.00539566f $X=4.05 $Y=1.94 $X2=0
+ $Y2=0
cc_131 N_A_190_48#_M1005_g N_A_27_368#_c_332_n 5.93853e-19 $X=1.025 $Y=0.74
+ $X2=0 $Y2=0
cc_132 N_A_190_48#_M1005_g N_A_27_368#_c_333_n 0.0015418f $X=1.025 $Y=0.74 $X2=0
+ $Y2=0
cc_133 N_A_190_48#_M1005_g N_A_27_368#_c_335_n 0.00506278f $X=1.025 $Y=0.74
+ $X2=0 $Y2=0
cc_134 N_A_190_48#_c_123_n N_A_27_368#_c_335_n 0.00146864f $X=1.04 $Y=1.765
+ $X2=0 $Y2=0
cc_135 N_A_190_48#_c_123_n N_A_27_368#_c_365_n 0.0153188f $X=1.04 $Y=1.765 $X2=0
+ $Y2=0
cc_136 N_A_190_48#_c_110_n N_A_27_368#_c_365_n 0.0200438f $X=1.49 $Y=1.765 $X2=0
+ $Y2=0
cc_137 N_A_190_48#_c_123_n N_A_27_368#_c_339_n 0.00787275f $X=1.04 $Y=1.765
+ $X2=0 $Y2=0
cc_138 N_A_190_48#_c_125_n N_A_27_368#_c_368_n 0.0141265f $X=4.03 $Y=2.815 $X2=0
+ $Y2=0
cc_139 N_A_190_48#_c_126_n N_A_27_368#_c_340_n 0.0559689f $X=4.03 $Y=2.105 $X2=0
+ $Y2=0
cc_140 N_A_190_48#_c_121_n N_A_27_368#_c_340_n 0.00677891f $X=4.05 $Y=1.94 $X2=0
+ $Y2=0
cc_141 N_A_190_48#_c_120_n N_A_27_368#_c_336_n 0.0280161f $X=3.705 $Y=1.115
+ $X2=0 $Y2=0
cc_142 N_A_190_48#_c_126_n N_A_27_368#_c_336_n 0.00244567f $X=4.03 $Y=2.105
+ $X2=0 $Y2=0
cc_143 N_A_190_48#_c_121_n N_A_27_368#_c_336_n 0.0249903f $X=4.05 $Y=1.94 $X2=0
+ $Y2=0
cc_144 N_A_190_48#_c_123_n N_VPWR_c_427_n 0.0106424f $X=1.04 $Y=1.765 $X2=0
+ $Y2=0
cc_145 N_A_190_48#_c_110_n N_VPWR_c_427_n 0.00139697f $X=1.49 $Y=1.765 $X2=0
+ $Y2=0
cc_146 N_A_190_48#_c_123_n N_VPWR_c_428_n 0.00413917f $X=1.04 $Y=1.765 $X2=0
+ $Y2=0
cc_147 N_A_190_48#_c_110_n N_VPWR_c_428_n 0.00415318f $X=1.49 $Y=1.765 $X2=0
+ $Y2=0
cc_148 N_A_190_48#_c_125_n N_VPWR_c_429_n 0.0164205f $X=4.03 $Y=2.815 $X2=0
+ $Y2=0
cc_149 N_A_190_48#_c_123_n N_VPWR_c_426_n 0.00414505f $X=1.04 $Y=1.765 $X2=0
+ $Y2=0
cc_150 N_A_190_48#_c_110_n N_VPWR_c_426_n 0.00414505f $X=1.49 $Y=1.765 $X2=0
+ $Y2=0
cc_151 N_A_190_48#_c_125_n N_VPWR_c_426_n 0.0135915f $X=4.03 $Y=2.815 $X2=0
+ $Y2=0
cc_152 N_A_190_48#_c_123_n N_VPWR_c_432_n 0.00106133f $X=1.04 $Y=1.765 $X2=0
+ $Y2=0
cc_153 N_A_190_48#_c_110_n N_VPWR_c_432_n 0.0134772f $X=1.49 $Y=1.765 $X2=0
+ $Y2=0
cc_154 N_A_190_48#_M1005_g N_X_c_471_n 0.00922867f $X=1.025 $Y=0.74 $X2=0 $Y2=0
cc_155 N_A_190_48#_M1013_g N_X_c_471_n 0.00930665f $X=1.455 $Y=0.74 $X2=0 $Y2=0
cc_156 N_A_190_48#_M1005_g N_X_c_472_n 0.0026107f $X=1.025 $Y=0.74 $X2=0 $Y2=0
cc_157 N_A_190_48#_c_108_n N_X_c_472_n 0.00246648f $X=1.38 $Y=1.375 $X2=0 $Y2=0
cc_158 N_A_190_48#_M1013_g N_X_c_472_n 0.00294637f $X=1.455 $Y=0.74 $X2=0 $Y2=0
cc_159 N_A_190_48#_c_190_p N_X_c_472_n 0.00733863f $X=1.745 $Y=1.045 $X2=0 $Y2=0
cc_160 N_A_190_48#_c_123_n X 0.0050636f $X=1.04 $Y=1.765 $X2=0 $Y2=0
cc_161 N_A_190_48#_c_108_n X 0.00501807f $X=1.38 $Y=1.375 $X2=0 $Y2=0
cc_162 N_A_190_48#_c_110_n X 0.00775563f $X=1.49 $Y=1.765 $X2=0 $Y2=0
cc_163 N_A_190_48#_c_117_n X 0.00206229f $X=1.66 $Y=1.465 $X2=0 $Y2=0
cc_164 N_A_190_48#_M1005_g N_X_c_473_n 0.00330399f $X=1.025 $Y=0.74 $X2=0 $Y2=0
cc_165 N_A_190_48#_c_107_n N_X_c_473_n 0.00437136f $X=1.04 $Y=1.675 $X2=0 $Y2=0
cc_166 N_A_190_48#_c_123_n N_X_c_473_n 0.00336883f $X=1.04 $Y=1.765 $X2=0 $Y2=0
cc_167 N_A_190_48#_c_108_n N_X_c_473_n 0.00668903f $X=1.38 $Y=1.375 $X2=0 $Y2=0
cc_168 N_A_190_48#_M1013_g N_X_c_473_n 9.29964e-19 $X=1.455 $Y=0.74 $X2=0 $Y2=0
cc_169 N_A_190_48#_c_110_n N_X_c_473_n 0.00400434f $X=1.49 $Y=1.765 $X2=0 $Y2=0
cc_170 N_A_190_48#_c_111_n N_X_c_473_n 0.00212694f $X=1.04 $Y=1.375 $X2=0 $Y2=0
cc_171 N_A_190_48#_c_112_n N_X_c_473_n 0.00551929f $X=1.66 $Y=1.3 $X2=0 $Y2=0
cc_172 N_A_190_48#_c_117_n N_X_c_473_n 0.0242992f $X=1.66 $Y=1.465 $X2=0 $Y2=0
cc_173 N_A_190_48#_c_113_n N_VGND_M1013_s 0.00218122f $X=2.175 $Y=1.045 $X2=0
+ $Y2=0
cc_174 N_A_190_48#_c_190_p N_VGND_M1013_s 0.00305443f $X=1.745 $Y=1.045 $X2=0
+ $Y2=0
cc_175 N_A_190_48#_c_119_n N_VGND_M1009_d 0.00526182f $X=3.375 $Y=1.115 $X2=0
+ $Y2=0
cc_176 N_A_190_48#_c_116_n N_VGND_M1011_d 0.00330281f $X=4.065 $Y=1.185 $X2=0
+ $Y2=0
cc_177 N_A_190_48#_M1005_g N_VGND_c_517_n 0.00709895f $X=1.025 $Y=0.74 $X2=0
+ $Y2=0
cc_178 N_A_190_48#_M1013_g N_VGND_c_518_n 0.00743057f $X=1.455 $Y=0.74 $X2=0
+ $Y2=0
cc_179 N_A_190_48#_c_110_n N_VGND_c_518_n 5.79784e-19 $X=1.49 $Y=1.765 $X2=0
+ $Y2=0
cc_180 N_A_190_48#_c_113_n N_VGND_c_518_n 0.0147668f $X=2.175 $Y=1.045 $X2=0
+ $Y2=0
cc_181 N_A_190_48#_c_190_p N_VGND_c_518_n 0.0129834f $X=1.745 $Y=1.045 $X2=0
+ $Y2=0
cc_182 N_A_190_48#_c_114_n N_VGND_c_518_n 0.0130314f $X=2.34 $Y=0.615 $X2=0
+ $Y2=0
cc_183 N_A_190_48#_c_114_n N_VGND_c_519_n 0.0134386f $X=2.34 $Y=0.615 $X2=0
+ $Y2=0
cc_184 N_A_190_48#_c_115_n N_VGND_c_519_n 0.00163718f $X=3.54 $Y=0.615 $X2=0
+ $Y2=0
cc_185 N_A_190_48#_c_119_n N_VGND_c_519_n 0.0314461f $X=3.375 $Y=1.115 $X2=0
+ $Y2=0
cc_186 N_A_190_48#_c_115_n N_VGND_c_521_n 0.0188012f $X=3.54 $Y=0.615 $X2=0
+ $Y2=0
cc_187 N_A_190_48#_c_116_n N_VGND_c_521_n 0.027045f $X=4.065 $Y=1.185 $X2=0
+ $Y2=0
cc_188 N_A_190_48#_M1005_g N_VGND_c_522_n 0.00417277f $X=1.025 $Y=0.74 $X2=0
+ $Y2=0
cc_189 N_A_190_48#_M1013_g N_VGND_c_522_n 0.00434272f $X=1.455 $Y=0.74 $X2=0
+ $Y2=0
cc_190 N_A_190_48#_c_114_n N_VGND_c_523_n 0.010412f $X=2.34 $Y=0.615 $X2=0 $Y2=0
cc_191 N_A_190_48#_c_115_n N_VGND_c_524_n 0.010139f $X=3.54 $Y=0.615 $X2=0 $Y2=0
cc_192 N_A_190_48#_M1005_g N_VGND_c_528_n 0.00770365f $X=1.025 $Y=0.74 $X2=0
+ $Y2=0
cc_193 N_A_190_48#_M1013_g N_VGND_c_528_n 0.00825059f $X=1.455 $Y=0.74 $X2=0
+ $Y2=0
cc_194 N_A_190_48#_c_114_n N_VGND_c_528_n 0.0113592f $X=2.34 $Y=0.615 $X2=0
+ $Y2=0
cc_195 N_A_190_48#_c_115_n N_VGND_c_528_n 0.0112086f $X=3.54 $Y=0.615 $X2=0
+ $Y2=0
cc_196 N_A_c_228_n N_B_c_266_n 0.0780322f $X=2.185 $Y=1.885 $X2=-0.19 $Y2=-0.245
cc_197 N_A_c_229_n N_B_c_266_n 0.00162913f $X=2.11 $Y=1.515 $X2=-0.19 $Y2=-0.245
cc_198 N_A_M1004_g N_B_M1009_g 0.0230804f $X=2.045 $Y=0.79 $X2=0 $Y2=0
cc_199 N_A_c_228_n N_B_M1009_g 0.00559311f $X=2.185 $Y=1.885 $X2=0 $Y2=0
cc_200 N_A_c_229_n N_B_M1009_g 7.46398e-19 $X=2.11 $Y=1.515 $X2=0 $Y2=0
cc_201 N_A_c_228_n B 0.00199525f $X=2.185 $Y=1.885 $X2=0 $Y2=0
cc_202 N_A_c_229_n B 0.0319684f $X=2.11 $Y=1.515 $X2=0 $Y2=0
cc_203 N_A_c_228_n N_A_27_368#_c_365_n 0.0126655f $X=2.185 $Y=1.885 $X2=0 $Y2=0
cc_204 N_A_c_229_n N_A_27_368#_c_365_n 0.0201317f $X=2.11 $Y=1.515 $X2=0 $Y2=0
cc_205 N_A_c_229_n N_VPWR_M1001_s 0.00403572f $X=2.11 $Y=1.515 $X2=0 $Y2=0
cc_206 N_A_c_228_n N_VPWR_c_429_n 0.00415318f $X=2.185 $Y=1.885 $X2=0 $Y2=0
cc_207 N_A_c_228_n N_VPWR_c_426_n 0.00414311f $X=2.185 $Y=1.885 $X2=0 $Y2=0
cc_208 N_A_c_228_n N_VPWR_c_432_n 0.0126617f $X=2.185 $Y=1.885 $X2=0 $Y2=0
cc_209 N_A_M1004_g N_X_c_471_n 8.75421e-19 $X=2.045 $Y=0.79 $X2=0 $Y2=0
cc_210 N_A_c_228_n X 2.76067e-19 $X=2.185 $Y=1.885 $X2=0 $Y2=0
cc_211 N_A_c_229_n X 0.0111406f $X=2.11 $Y=1.515 $X2=0 $Y2=0
cc_212 N_A_M1004_g N_VGND_c_518_n 0.00862467f $X=2.045 $Y=0.79 $X2=0 $Y2=0
cc_213 N_A_M1004_g N_VGND_c_519_n 5.59444e-19 $X=2.045 $Y=0.79 $X2=0 $Y2=0
cc_214 N_A_M1004_g N_VGND_c_523_n 0.00421418f $X=2.045 $Y=0.79 $X2=0 $Y2=0
cc_215 N_A_M1004_g N_VGND_c_528_n 0.00432128f $X=2.045 $Y=0.79 $X2=0 $Y2=0
cc_216 N_B_c_266_n N_C_c_300_n 0.0642377f $X=2.605 $Y=1.885 $X2=-0.19 $Y2=-0.245
cc_217 B N_C_c_300_n 0.00163768f $X=2.555 $Y=1.58 $X2=-0.19 $Y2=-0.245
cc_218 N_B_M1009_g N_C_M1002_g 0.0250853f $X=2.635 $Y=0.79 $X2=0 $Y2=0
cc_219 N_B_c_266_n C 0.00247798f $X=2.605 $Y=1.885 $X2=0 $Y2=0
cc_220 B C 0.0434889f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_221 N_B_c_266_n N_A_27_368#_c_365_n 0.00242272f $X=2.605 $Y=1.885 $X2=0 $Y2=0
cc_222 N_B_c_266_n N_A_27_368#_c_377_n 0.00429727f $X=2.605 $Y=1.885 $X2=0 $Y2=0
cc_223 N_B_c_266_n N_A_27_368#_c_368_n 0.0124461f $X=2.605 $Y=1.885 $X2=0 $Y2=0
cc_224 B N_A_27_368#_c_368_n 0.0070622f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_225 N_B_c_266_n N_VPWR_c_429_n 0.00307159f $X=2.605 $Y=1.885 $X2=0 $Y2=0
cc_226 N_B_c_266_n N_VPWR_c_426_n 0.00378101f $X=2.605 $Y=1.885 $X2=0 $Y2=0
cc_227 N_B_c_266_n N_VPWR_c_432_n 0.00120756f $X=2.605 $Y=1.885 $X2=0 $Y2=0
cc_228 B A_536_392# 0.00324694f $X=2.555 $Y=1.58 $X2=-0.19 $Y2=-0.245
cc_229 N_B_M1009_g N_VGND_c_518_n 5.60991e-19 $X=2.635 $Y=0.79 $X2=0 $Y2=0
cc_230 N_B_M1009_g N_VGND_c_519_n 0.0142125f $X=2.635 $Y=0.79 $X2=0 $Y2=0
cc_231 N_B_M1009_g N_VGND_c_523_n 0.00421418f $X=2.635 $Y=0.79 $X2=0 $Y2=0
cc_232 N_B_M1009_g N_VGND_c_528_n 0.00432128f $X=2.635 $Y=0.79 $X2=0 $Y2=0
cc_233 N_C_c_300_n N_A_27_368#_c_330_n 0.0385279f $X=3.115 $Y=1.885 $X2=0 $Y2=0
cc_234 N_C_M1002_g N_A_27_368#_c_330_n 0.0223905f $X=3.28 $Y=0.79 $X2=0 $Y2=0
cc_235 C N_A_27_368#_c_330_n 0.00281736f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_236 N_C_M1002_g N_A_27_368#_M1011_g 0.0173114f $X=3.28 $Y=0.79 $X2=0 $Y2=0
cc_237 N_C_c_300_n N_A_27_368#_c_368_n 0.0116346f $X=3.115 $Y=1.885 $X2=0 $Y2=0
cc_238 C N_A_27_368#_c_368_n 0.0195203f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_239 N_C_c_300_n N_A_27_368#_c_340_n 9.4827e-19 $X=3.115 $Y=1.885 $X2=0 $Y2=0
cc_240 C N_A_27_368#_c_340_n 0.037626f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_241 N_C_M1002_g N_A_27_368#_c_336_n 0.00238017f $X=3.28 $Y=0.79 $X2=0 $Y2=0
cc_242 C N_A_27_368#_c_336_n 0.0240984f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_243 N_C_c_300_n N_VPWR_c_429_n 0.00307159f $X=3.115 $Y=1.885 $X2=0 $Y2=0
cc_244 N_C_c_300_n N_VPWR_c_426_n 0.00379127f $X=3.115 $Y=1.885 $X2=0 $Y2=0
cc_245 C A_638_392# 0.00605657f $X=3.035 $Y=1.58 $X2=-0.19 $Y2=-0.245
cc_246 N_C_M1002_g N_VGND_c_519_n 0.00481242f $X=3.28 $Y=0.79 $X2=0 $Y2=0
cc_247 N_C_M1002_g N_VGND_c_524_n 0.00505936f $X=3.28 $Y=0.79 $X2=0 $Y2=0
cc_248 N_C_M1002_g N_VGND_c_528_n 0.00514438f $X=3.28 $Y=0.79 $X2=0 $Y2=0
cc_249 N_A_27_368#_c_335_n N_VPWR_M1006_d 0.00286058f $X=0.805 $Y=1.95 $X2=-0.19
+ $Y2=-0.245
cc_250 N_A_27_368#_c_365_n N_VPWR_M1006_d 8.26908e-19 $X=2.295 $Y=2.405
+ $X2=-0.19 $Y2=-0.245
cc_251 N_A_27_368#_c_339_n N_VPWR_M1006_d 0.0122292f $X=0.89 $Y=2.405 $X2=-0.19
+ $Y2=-0.245
cc_252 N_A_27_368#_c_365_n N_VPWR_M1001_s 0.0182031f $X=2.295 $Y=2.405 $X2=0
+ $Y2=0
cc_253 N_A_27_368#_c_365_n N_VPWR_c_427_n 0.00239871f $X=2.295 $Y=2.405 $X2=0
+ $Y2=0
cc_254 N_A_27_368#_c_339_n N_VPWR_c_427_n 0.023618f $X=0.89 $Y=2.405 $X2=0 $Y2=0
cc_255 N_A_27_368#_c_330_n N_VPWR_c_429_n 0.00343069f $X=3.655 $Y=1.885 $X2=0
+ $Y2=0
cc_256 N_A_27_368#_c_368_n N_VPWR_c_429_n 0.0290018f $X=3.525 $Y=2.775 $X2=0
+ $Y2=0
cc_257 N_A_27_368#_c_398_p N_VPWR_c_429_n 0.00455517f $X=2.465 $Y=2.775 $X2=0
+ $Y2=0
cc_258 N_A_27_368#_c_330_n N_VPWR_c_426_n 0.00506439f $X=3.655 $Y=1.885 $X2=0
+ $Y2=0
cc_259 N_A_27_368#_c_365_n N_VPWR_c_426_n 0.0251488f $X=2.295 $Y=2.405 $X2=0
+ $Y2=0
cc_260 N_A_27_368#_c_339_n N_VPWR_c_426_n 0.0183179f $X=0.89 $Y=2.405 $X2=0
+ $Y2=0
cc_261 N_A_27_368#_c_368_n N_VPWR_c_426_n 0.0380899f $X=3.525 $Y=2.775 $X2=0
+ $Y2=0
cc_262 N_A_27_368#_c_398_p N_VPWR_c_426_n 0.00575379f $X=2.465 $Y=2.775 $X2=0
+ $Y2=0
cc_263 N_A_27_368#_c_339_n N_VPWR_c_431_n 0.00671799f $X=0.89 $Y=2.405 $X2=0
+ $Y2=0
cc_264 N_A_27_368#_c_365_n N_VPWR_c_432_n 0.0272735f $X=2.295 $Y=2.405 $X2=0
+ $Y2=0
cc_265 N_A_27_368#_c_365_n N_X_M1000_d 0.00571673f $X=2.295 $Y=2.405 $X2=0 $Y2=0
cc_266 N_A_27_368#_c_332_n N_X_c_471_n 0.00448258f $X=0.295 $Y=0.835 $X2=0 $Y2=0
cc_267 N_A_27_368#_c_333_n N_X_c_472_n 0.0143703f $X=0.72 $Y=1.095 $X2=0 $Y2=0
cc_268 N_A_27_368#_c_365_n X 0.0195872f $X=2.295 $Y=2.405 $X2=0 $Y2=0
cc_269 N_A_27_368#_c_339_n X 0.016649f $X=0.89 $Y=2.405 $X2=0 $Y2=0
cc_270 N_A_27_368#_c_335_n N_X_c_473_n 0.0556308f $X=0.805 $Y=1.95 $X2=0 $Y2=0
cc_271 N_A_27_368#_c_365_n A_452_392# 0.0090591f $X=2.295 $Y=2.405 $X2=-0.19
+ $Y2=-0.245
cc_272 N_A_27_368#_c_377_n A_452_392# 0.00230601f $X=2.38 $Y=2.69 $X2=-0.19
+ $Y2=-0.245
cc_273 N_A_27_368#_c_368_n A_452_392# 3.64674e-19 $X=3.525 $Y=2.775 $X2=-0.19
+ $Y2=-0.245
cc_274 N_A_27_368#_c_398_p A_452_392# 0.00245088f $X=2.465 $Y=2.775 $X2=-0.19
+ $Y2=-0.245
cc_275 N_A_27_368#_c_368_n A_536_392# 0.0113255f $X=3.525 $Y=2.775 $X2=-0.19
+ $Y2=-0.245
cc_276 N_A_27_368#_c_368_n A_638_392# 0.0117123f $X=3.525 $Y=2.775 $X2=-0.19
+ $Y2=-0.245
cc_277 N_A_27_368#_c_333_n N_VGND_M1010_d 0.0041785f $X=0.72 $Y=1.095 $X2=-0.19
+ $Y2=-0.245
cc_278 N_A_27_368#_c_332_n N_VGND_c_517_n 0.0114804f $X=0.295 $Y=0.835 $X2=0
+ $Y2=0
cc_279 N_A_27_368#_c_333_n N_VGND_c_517_n 0.0215468f $X=0.72 $Y=1.095 $X2=0
+ $Y2=0
cc_280 N_A_27_368#_M1011_g N_VGND_c_521_n 0.0126413f $X=3.755 $Y=0.79 $X2=0
+ $Y2=0
cc_281 N_A_27_368#_M1011_g N_VGND_c_524_n 0.00485498f $X=3.755 $Y=0.79 $X2=0
+ $Y2=0
cc_282 N_A_27_368#_c_332_n N_VGND_c_525_n 0.00811255f $X=0.295 $Y=0.835 $X2=0
+ $Y2=0
cc_283 N_A_27_368#_M1011_g N_VGND_c_528_n 0.00514438f $X=3.755 $Y=0.79 $X2=0
+ $Y2=0
cc_284 N_A_27_368#_c_332_n N_VGND_c_528_n 0.0106114f $X=0.295 $Y=0.835 $X2=0
+ $Y2=0
cc_285 N_X_c_471_n N_VGND_c_517_n 0.0373918f $X=1.24 $Y=0.515 $X2=0 $Y2=0
cc_286 N_X_c_471_n N_VGND_c_518_n 0.0170646f $X=1.24 $Y=0.515 $X2=0 $Y2=0
cc_287 N_X_c_471_n N_VGND_c_522_n 0.0151167f $X=1.24 $Y=0.515 $X2=0 $Y2=0
cc_288 N_X_c_471_n N_VGND_c_528_n 0.0123643f $X=1.24 $Y=0.515 $X2=0 $Y2=0
