* File: sky130_fd_sc_hs__or3_2.pex.spice
* Created: Thu Aug 27 21:05:55 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HS__OR3_2%C 3 5 6 8 9 10 14 15 16
c38 16 0 4.32539e-20 $X=0.592 $Y=1.12
r39 14 16 46.3655 $w=3.45e-07 $l=1.65e-07 $layer=POLY_cond $X=0.592 $Y=1.285
+ $X2=0.592 $Y2=1.12
r40 14 15 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.6
+ $Y=1.285 $X2=0.6 $Y2=1.285
r41 9 10 10.6601 $w=3.98e-07 $l=3.7e-07 $layer=LI1_cond $X=0.635 $Y=1.295
+ $X2=0.635 $Y2=1.665
r42 9 15 0.288111 $w=3.98e-07 $l=1e-08 $layer=LI1_cond $X=0.635 $Y=1.295
+ $X2=0.635 $Y2=1.285
r43 6 8 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=0.675 $Y=1.885
+ $X2=0.675 $Y2=2.46
r44 5 6 44.9979 $w=2.86e-07 $l=3.05696e-07 $layer=POLY_cond $X=0.592 $Y=1.618
+ $X2=0.675 $Y2=1.885
r45 4 14 1.17081 $w=3.45e-07 $l=7e-09 $layer=POLY_cond $X=0.592 $Y=1.292
+ $X2=0.592 $Y2=1.285
r46 4 5 54.5263 $w=3.45e-07 $l=3.26e-07 $layer=POLY_cond $X=0.592 $Y=1.292
+ $X2=0.592 $Y2=1.618
r47 3 16 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=0.495 $Y=0.69
+ $X2=0.495 $Y2=1.12
.ends

.subckt PM_SKY130_FD_SC_HS__OR3_2%B 1 3 6 8 9 10 11 12 17 18
c47 1 0 1.74045e-19 $X=1.095 $Y=1.885
r48 17 18 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.17
+ $Y=1.295 $X2=1.17 $Y2=1.295
r49 11 12 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.17 $Y=2.405
+ $X2=1.17 $Y2=2.775
r50 10 11 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.17 $Y=2.035
+ $X2=1.17 $Y2=2.405
r51 10 18 25.8427 $w=3.28e-07 $l=7.4e-07 $layer=LI1_cond $X=1.17 $Y=2.035
+ $X2=1.17 $Y2=1.295
r52 9 17 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.17 $Y=1.635
+ $X2=1.17 $Y2=1.295
r53 8 17 38.6168 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.17 $Y=1.13
+ $X2=1.17 $Y2=1.295
r54 6 8 141.387 $w=1.5e-07 $l=4.4e-07 $layer=POLY_cond $X=1.15 $Y=0.69 $X2=1.15
+ $Y2=1.13
r55 1 9 43.19 $w=2.79e-07 $l=2.85044e-07 $layer=POLY_cond $X=1.095 $Y=1.885
+ $X2=1.17 $Y2=1.635
r56 1 3 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=1.095 $Y=1.885
+ $X2=1.095 $Y2=2.46
.ends

.subckt PM_SKY130_FD_SC_HS__OR3_2%A 3 6 7 9 10 13
r43 13 16 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.74 $Y=1.385
+ $X2=1.74 $Y2=1.55
r44 13 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.74 $Y=1.385
+ $X2=1.74 $Y2=1.22
r45 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.74
+ $Y=1.385 $X2=1.74 $Y2=1.385
r46 10 14 3.05058 $w=3.38e-07 $l=9e-08 $layer=LI1_cond $X=1.735 $Y=1.295
+ $X2=1.735 $Y2=1.385
r47 7 9 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=1.665 $Y=1.885
+ $X2=1.665 $Y2=2.46
r48 6 7 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=1.665 $Y=1.795 $X2=1.665
+ $Y2=1.885
r49 6 16 95.2339 $w=1.8e-07 $l=2.45e-07 $layer=POLY_cond $X=1.665 $Y=1.795
+ $X2=1.665 $Y2=1.55
r50 3 15 271.766 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=1.65 $Y=0.69 $X2=1.65
+ $Y2=1.22
.ends

.subckt PM_SKY130_FD_SC_HS__OR3_2%A_27_74# 1 2 3 10 12 15 17 19 22 26 29 32 34
+ 36 39 42 43 45 48 52 54 58
c107 54 0 4.32539e-20 $X=1.365 $Y=0.87
c108 52 0 1.74045e-19 $X=0.45 $Y=2.125
r109 58 59 8.8094 $w=3.83e-07 $l=7e-08 $layer=POLY_cond $X=2.725 $Y=1.532
+ $X2=2.795 $Y2=1.532
r110 55 56 11.3264 $w=3.83e-07 $l=9e-08 $layer=POLY_cond $X=2.275 $Y=1.532
+ $X2=2.365 $Y2=1.532
r111 49 52 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=0.18 $Y=2.045
+ $X2=0.45 $Y2=2.045
r112 46 58 9.43864 $w=3.83e-07 $l=7.5e-08 $layer=POLY_cond $X=2.65 $Y=1.532
+ $X2=2.725 $Y2=1.532
r113 46 56 35.8668 $w=3.83e-07 $l=2.85e-07 $layer=POLY_cond $X=2.65 $Y=1.532
+ $X2=2.365 $Y2=1.532
r114 45 46 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.65
+ $Y=1.465 $X2=2.65 $Y2=1.465
r115 43 45 14.1436 $w=3.28e-07 $l=4.05e-07 $layer=LI1_cond $X=2.245 $Y=1.465
+ $X2=2.65 $Y2=1.465
r116 42 43 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.16 $Y=1.3
+ $X2=2.245 $Y2=1.465
r117 41 42 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=2.16 $Y=0.96
+ $X2=2.16 $Y2=1.3
r118 40 54 8.61065 $w=1.7e-07 $l=1.67481e-07 $layer=LI1_cond $X=1.53 $Y=0.875
+ $X2=1.365 $Y2=0.87
r119 39 41 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.075 $Y=0.875
+ $X2=2.16 $Y2=0.96
r120 39 40 35.5561 $w=1.68e-07 $l=5.45e-07 $layer=LI1_cond $X=2.075 $Y=0.875
+ $X2=1.53 $Y2=0.875
r121 36 54 0.89609 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=1.365 $Y=0.78
+ $X2=1.365 $Y2=0.87
r122 36 38 4.62121 $w=3.3e-07 $l=1.25e-07 $layer=LI1_cond $X=1.365 $Y=0.78
+ $X2=1.365 $Y2=0.655
r123 35 48 2.90867 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=0.445 $Y=0.865
+ $X2=0.27 $Y2=0.865
r124 34 54 8.61065 $w=1.7e-07 $l=1.67481e-07 $layer=LI1_cond $X=1.2 $Y=0.865
+ $X2=1.365 $Y2=0.87
r125 34 35 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=1.2 $Y=0.865
+ $X2=0.445 $Y2=0.865
r126 32 52 23.9219 $w=3.28e-07 $l=6.85e-07 $layer=LI1_cond $X=0.45 $Y=2.815
+ $X2=0.45 $Y2=2.13
r127 29 49 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.18 $Y=1.96
+ $X2=0.18 $Y2=2.045
r128 28 48 3.58051 $w=2.6e-07 $l=1.25499e-07 $layer=LI1_cond $X=0.18 $Y=0.95
+ $X2=0.27 $Y2=0.865
r129 28 29 65.8931 $w=1.68e-07 $l=1.01e-06 $layer=LI1_cond $X=0.18 $Y=0.95
+ $X2=0.18 $Y2=1.96
r130 24 48 3.58051 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=0.27 $Y=0.78
+ $X2=0.27 $Y2=0.865
r131 24 26 4.2805 $w=3.48e-07 $l=1.3e-07 $layer=LI1_cond $X=0.27 $Y=0.78
+ $X2=0.27 $Y2=0.65
r132 20 59 24.8035 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=2.795 $Y=1.3
+ $X2=2.795 $Y2=1.532
r133 20 22 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=2.795 $Y=1.3
+ $X2=2.795 $Y2=0.74
r134 17 58 24.8035 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=2.725 $Y=1.765
+ $X2=2.725 $Y2=1.532
r135 17 19 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.725 $Y=1.765
+ $X2=2.725 $Y2=2.4
r136 13 56 24.8035 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=2.365 $Y=1.3
+ $X2=2.365 $Y2=1.532
r137 13 15 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=2.365 $Y=1.3
+ $X2=2.365 $Y2=0.74
r138 10 55 24.8035 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=2.275 $Y=1.765
+ $X2=2.275 $Y2=1.532
r139 10 12 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.275 $Y=1.765
+ $X2=2.275 $Y2=2.4
r140 3 52 400 $w=1.7e-07 $l=2.26164e-07 $layer=licon1_PDIFF $count=1 $X=0.305
+ $Y=1.96 $X2=0.45 $Y2=2.125
r141 3 32 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=0.305
+ $Y=1.96 $X2=0.45 $Y2=2.815
r142 2 38 182 $w=1.7e-07 $l=3.4803e-07 $layer=licon1_NDIFF $count=1 $X=1.225
+ $Y=0.37 $X2=1.365 $Y2=0.655
r143 1 26 182 $w=1.7e-07 $l=3.44964e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.65
.ends

.subckt PM_SKY130_FD_SC_HS__OR3_2%VPWR 1 2 9 13 15 18 19 20 29 35
r36 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r37 32 35 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r38 31 32 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r39 29 34 4.58274 $w=1.7e-07 $l=2.62e-07 $layer=LI1_cond $X=2.835 $Y=3.33
+ $X2=3.097 $Y2=3.33
r40 29 31 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=2.835 $Y=3.33
+ $X2=2.64 $Y2=3.33
r41 23 27 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=0.24 $Y=3.33
+ $X2=1.68 $Y2=3.33
r42 23 24 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r43 20 32 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.64 $Y2=3.33
r44 20 24 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=0.24 $Y2=3.33
r45 20 27 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r46 18 27 2.93583 $w=1.68e-07 $l=4.5e-08 $layer=LI1_cond $X=1.725 $Y=3.33
+ $X2=1.68 $Y2=3.33
r47 18 19 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.725 $Y=3.33
+ $X2=1.89 $Y2=3.33
r48 17 31 38.1658 $w=1.68e-07 $l=5.85e-07 $layer=LI1_cond $X=2.055 $Y=3.33
+ $X2=2.64 $Y2=3.33
r49 17 19 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.055 $Y=3.33
+ $X2=1.89 $Y2=3.33
r50 13 34 3.18343 $w=3.3e-07 $l=1.32868e-07 $layer=LI1_cond $X=3 $Y=3.245
+ $X2=3.097 $Y2=3.33
r51 13 15 35.621 $w=3.28e-07 $l=1.02e-06 $layer=LI1_cond $X=3 $Y=3.245 $X2=3
+ $Y2=2.225
r52 9 12 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=1.89 $Y=2.105 $X2=1.89
+ $Y2=2.815
r53 7 19 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.89 $Y=3.245 $X2=1.89
+ $Y2=3.33
r54 7 12 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=1.89 $Y=3.245
+ $X2=1.89 $Y2=2.815
r55 2 15 300 $w=1.7e-07 $l=4.74579e-07 $layer=licon1_PDIFF $count=2 $X=2.8
+ $Y=1.84 $X2=3 $Y2=2.225
r56 1 12 400 $w=1.7e-07 $l=9.26971e-07 $layer=licon1_PDIFF $count=1 $X=1.74
+ $Y=1.96 $X2=1.89 $Y2=2.815
r57 1 9 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=1.74
+ $Y=1.96 $X2=1.89 $Y2=2.105
.ends

.subckt PM_SKY130_FD_SC_HS__OR3_2%X 1 2 9 15 17 18 19 20 23 24
r46 23 24 18.5393 $w=2.28e-07 $l=3.7e-07 $layer=LI1_cond $X=3.12 $Y=1.295
+ $X2=3.12 $Y2=1.665
r47 22 24 6.76434 $w=2.28e-07 $l=1.35e-07 $layer=LI1_cond $X=3.12 $Y=1.8
+ $X2=3.12 $Y2=1.665
r48 21 23 8.26753 $w=2.28e-07 $l=1.65e-07 $layer=LI1_cond $X=3.12 $Y=1.13
+ $X2=3.12 $Y2=1.295
r49 19 21 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=3.005 $Y=1.045
+ $X2=3.12 $Y2=1.13
r50 19 20 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=3.005 $Y=1.045
+ $X2=2.745 $Y2=1.045
r51 17 22 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=3.005 $Y=1.885
+ $X2=3.12 $Y2=1.8
r52 17 18 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=3.005 $Y=1.885
+ $X2=2.665 $Y2=1.885
r53 13 20 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.58 $Y=0.96
+ $X2=2.745 $Y2=1.045
r54 13 15 15.5405 $w=3.28e-07 $l=4.45e-07 $layer=LI1_cond $X=2.58 $Y=0.96
+ $X2=2.58 $Y2=0.515
r55 9 11 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=2.5 $Y=1.985 $X2=2.5
+ $Y2=2.815
r56 7 18 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.5 $Y=1.97
+ $X2=2.665 $Y2=1.885
r57 7 9 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=2.5 $Y=1.97 $X2=2.5
+ $Y2=1.985
r58 2 11 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=2.35
+ $Y=1.84 $X2=2.5 $Y2=2.815
r59 2 9 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=2.35
+ $Y=1.84 $X2=2.5 $Y2=1.985
r60 1 15 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.44
+ $Y=0.37 $X2=2.58 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__OR3_2%VGND 1 2 3 12 14 16 18 20 25 30 36 47
r42 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r43 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r44 34 47 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r45 34 41 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=2.16
+ $Y2=0
r46 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r47 31 33 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=2.245 $Y=0 $X2=2.64
+ $Y2=0
r48 30 46 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=2.915 $Y=0 $X2=3.137
+ $Y2=0
r49 30 33 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=2.915 $Y=0 $X2=2.64
+ $Y2=0
r50 26 36 10.0494 $w=1.7e-07 $l=2.08e-07 $layer=LI1_cond $X=1.03 $Y=0 $X2=0.822
+ $Y2=0
r51 26 28 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=1.03 $Y=0 $X2=1.68
+ $Y2=0
r52 25 43 11.3024 $w=5.43e-07 $l=5.15e-07 $layer=LI1_cond $X=1.972 $Y=0
+ $X2=1.972 $Y2=0.515
r53 25 31 7.70116 $w=1.7e-07 $l=2.73e-07 $layer=LI1_cond $X=1.972 $Y=0 $X2=2.245
+ $Y2=0
r54 25 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r55 25 28 1.30481 $w=1.68e-07 $l=2e-08 $layer=LI1_cond $X=1.7 $Y=0 $X2=1.68
+ $Y2=0
r56 23 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r57 22 23 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r58 20 36 10.0494 $w=1.7e-07 $l=2.07e-07 $layer=LI1_cond $X=0.615 $Y=0 $X2=0.822
+ $Y2=0
r59 20 22 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=0.615 $Y=0 $X2=0.24
+ $Y2=0
r60 18 41 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r61 18 37 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=0.72
+ $Y2=0
r62 18 28 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r63 14 46 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=3.08 $Y=0.085
+ $X2=3.137 $Y2=0
r64 14 16 16.9374 $w=3.28e-07 $l=4.85e-07 $layer=LI1_cond $X=3.08 $Y=0.085
+ $X2=3.08 $Y2=0.57
r65 10 36 1.57254 $w=4.15e-07 $l=8.5e-08 $layer=LI1_cond $X=0.822 $Y=0.085
+ $X2=0.822 $Y2=0
r66 10 12 11.941 $w=4.13e-07 $l=4.3e-07 $layer=LI1_cond $X=0.822 $Y=0.085
+ $X2=0.822 $Y2=0.515
r67 3 16 182 $w=1.7e-07 $l=2.93428e-07 $layer=licon1_NDIFF $count=1 $X=2.87
+ $Y=0.37 $X2=3.08 $Y2=0.57
r68 2 43 182 $w=1.7e-07 $l=3.09112e-07 $layer=licon1_NDIFF $count=1 $X=1.725
+ $Y=0.37 $X2=1.97 $Y2=0.515
r69 1 12 182 $w=1.7e-07 $l=3.14245e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.37 $X2=0.82 $Y2=0.515
.ends

