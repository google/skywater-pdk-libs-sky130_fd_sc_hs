* File: sky130_fd_sc_hs__xor2_4.spice
* Created: Thu Aug 27 21:13:09 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hs__xor2_4.pex.spice"
.subckt sky130_fd_sc_hs__xor2_4  VNB VPB A B VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* B	B
* A	A
* VPB	VPB
* VNB	VNB
MM1001 N_A_160_98#_M1001_d N_A_M1001_g N_VGND_M1001_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.3811 PD=1.02 PS=2.51 NRD=0 NRS=40.536 M=1 R=4.93333 SA=75000.4
+ SB=75003.2 A=0.111 P=1.78 MULT=1
MM1022 N_A_160_98#_M1001_d N_A_M1022_g N_VGND_M1022_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.20775 PD=1.02 PS=1.49 NRD=0 NRS=36.6 M=1 R=4.93333 SA=75000.9
+ SB=75002.8 A=0.111 P=1.78 MULT=1
MM1023 N_A_160_98#_M1023_d N_B_M1023_g N_VGND_M1022_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1443 AS=0.20775 PD=1.13 PS=1.49 NRD=8.916 NRS=36.6 M=1 R=4.93333
+ SA=75001.5 SB=75002.2 A=0.111 P=1.78 MULT=1
MM1028 N_A_160_98#_M1023_d N_B_M1028_g N_VGND_M1028_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1443 AS=0.20775 PD=1.13 PS=1.49 NRD=8.916 NRS=36.6 M=1 R=4.93333 SA=75002
+ SB=75001.7 A=0.111 P=1.78 MULT=1
MM1011 N_VGND_M1028_s N_A_160_98#_M1011_g N_X_M1011_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.20775 AS=0.20905 PD=1.49 PS=1.305 NRD=36.6 NRS=46.212 M=1 R=4.93333
+ SA=75002.6 SB=75001.1 A=0.111 P=1.78 MULT=1
MM1029 N_VGND_M1029_d N_A_160_98#_M1029_g N_X_M1011_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.44175 AS=0.20905 PD=2.96 PS=1.305 NRD=87.876 NRS=0 M=1 R=4.93333
+ SA=75003.3 SB=75000.4 A=0.111 P=1.78 MULT=1
MM1012 N_VGND_M1012_d N_A_M1012_g N_A_877_74#_M1012_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1889 AS=0.2109 PD=1.36 PS=2.05 NRD=32.472 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75003.6 A=0.111 P=1.78 MULT=1
MM1014 N_VGND_M1012_d N_A_M1014_g N_A_877_74#_M1014_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1889 AS=0.1036 PD=1.36 PS=1.02 NRD=32.472 NRS=0 M=1 R=4.93333 SA=75000.8
+ SB=75003 A=0.111 P=1.78 MULT=1
MM1025 N_VGND_M1025_d N_A_M1025_g N_A_877_74#_M1014_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1889 AS=0.1036 PD=1.36 PS=1.02 NRD=32.472 NRS=0 M=1 R=4.93333 SA=75001.2
+ SB=75002.6 A=0.111 P=1.78 MULT=1
MM1026 N_VGND_M1025_d N_A_M1026_g N_A_877_74#_M1026_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1889 AS=0.1036 PD=1.36 PS=1.02 NRD=32.472 NRS=0 M=1 R=4.93333 SA=75001.8
+ SB=75002 A=0.111 P=1.78 MULT=1
MM1006 N_X_M1006_d N_B_M1006_g N_A_877_74#_M1026_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75002.2
+ SB=75001.6 A=0.111 P=1.78 MULT=1
MM1009 N_X_M1006_d N_B_M1009_g N_A_877_74#_M1009_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1295 PD=1.02 PS=1.09 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75002.7
+ SB=75001.1 A=0.111 P=1.78 MULT=1
MM1021 N_X_M1021_d N_B_M1021_g N_A_877_74#_M1009_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1295 PD=1.02 PS=1.09 NRD=0 NRS=0 M=1 R=4.93333 SA=75003.2
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1024 N_X_M1021_d N_B_M1024_g N_A_877_74#_M1024_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.2109 PD=1.02 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333 SA=75003.6
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1013 N_A_36_392#_M1013_d N_A_M1013_g N_VPWR_M1013_s VPB PSHORT L=0.15 W=1
+ AD=0.295 AS=0.175 PD=2.59 PS=1.35 NRD=1.9503 NRS=1.9503 M=1 R=6.66667
+ SA=75000.2 SB=75001.6 A=0.15 P=2.3 MULT=1
MM1018 N_A_36_392#_M1018_d N_A_M1018_g N_VPWR_M1013_s VPB PSHORT L=0.15 W=1
+ AD=0.15 AS=0.175 PD=1.3 PS=1.35 NRD=1.9503 NRS=11.8003 M=1 R=6.66667
+ SA=75000.7 SB=75001.1 A=0.15 P=2.3 MULT=1
MM1017 N_A_160_98#_M1017_d N_B_M1017_g N_A_36_392#_M1018_d VPB PSHORT L=0.15 W=1
+ AD=0.15 AS=0.15 PD=1.3 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=6.66667 SA=75001.2
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1020 N_A_160_98#_M1017_d N_B_M1020_g N_A_36_392#_M1020_s VPB PSHORT L=0.15 W=1
+ AD=0.15 AS=0.275 PD=1.3 PS=2.55 NRD=1.9503 NRS=1.9503 M=1 R=6.66667 SA=75001.6
+ SB=75000.2 A=0.15 P=2.3 MULT=1
MM1000 N_A_514_368#_M1000_d N_A_160_98#_M1000_g N_X_M1000_s VPB PSHORT L=0.15
+ W=1.12 AD=0.3136 AS=0.168 PD=2.8 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75005.4 A=0.168 P=2.54 MULT=1
MM1002 N_A_514_368#_M1002_d N_A_160_98#_M1002_g N_X_M1000_s VPB PSHORT L=0.15
+ W=1.12 AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.7 SB=75005 A=0.168 P=2.54 MULT=1
MM1003 N_A_514_368#_M1002_d N_A_160_98#_M1003_g N_X_M1003_s VPB PSHORT L=0.15
+ W=1.12 AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.1 SB=75004.5 A=0.168 P=2.54 MULT=1
MM1027 N_A_514_368#_M1027_d N_A_160_98#_M1027_g N_X_M1003_s VPB PSHORT L=0.15
+ W=1.12 AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.6 SB=75004.1 A=0.168 P=2.54 MULT=1
MM1004 N_A_514_368#_M1027_d N_A_M1004_g N_VPWR_M1004_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.27695 PD=1.42 PS=1.795 NRD=1.7533 NRS=33.8052 M=1 R=7.46667
+ SA=75002 SB=75003.6 A=0.168 P=2.54 MULT=1
MM1005 N_A_514_368#_M1005_d N_A_M1005_g N_VPWR_M1004_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.27695 PD=1.42 PS=1.795 NRD=1.7533 NRS=33.8052 M=1 R=7.46667
+ SA=75002.6 SB=75003 A=0.168 P=2.54 MULT=1
MM1010 N_A_514_368#_M1005_d N_A_M1010_g N_VPWR_M1010_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.270175 PD=1.42 PS=1.785 NRD=1.7533 NRS=32.7414 M=1 R=7.46667
+ SA=75003 SB=75002.6 A=0.168 P=2.54 MULT=1
MM1015 N_A_514_368#_M1015_d N_A_M1015_g N_VPWR_M1010_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.270175 PD=1.42 PS=1.785 NRD=1.7533 NRS=32.7414 M=1 R=7.46667
+ SA=75003.6 SB=75002 A=0.168 P=2.54 MULT=1
MM1007 N_VPWR_M1007_d N_B_M1007_g N_A_514_368#_M1015_d VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75004.1 SB=75001.6 A=0.168 P=2.54 MULT=1
MM1008 N_VPWR_M1007_d N_B_M1008_g N_A_514_368#_M1008_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75004.5 SB=75001.1 A=0.168 P=2.54 MULT=1
MM1016 N_VPWR_M1016_d N_B_M1016_g N_A_514_368#_M1008_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667 SA=75005
+ SB=75000.7 A=0.168 P=2.54 MULT=1
MM1019 N_VPWR_M1016_d N_B_M1019_g N_A_514_368#_M1019_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.3192 PD=1.42 PS=2.81 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75005.4 SB=75000.2 A=0.168 P=2.54 MULT=1
DX30_noxref VNB VPB NWDIODE A=16.7772 P=21.76
*
.include "sky130_fd_sc_hs__xor2_4.pxi.spice"
*
.ends
*
*
