* File: sky130_fd_sc_hs__nor2_2.pxi.spice
* Created: Tue Sep  1 20:10:50 2020
* 
x_PM_SKY130_FD_SC_HS__NOR2_2%B N_B_M1004_g N_B_M1003_g N_B_c_40_n N_B_c_45_n
+ N_B_M1005_g N_B_c_41_n N_B_c_42_n N_B_c_47_n B PM_SKY130_FD_SC_HS__NOR2_2%B
x_PM_SKY130_FD_SC_HS__NOR2_2%A N_A_c_80_n N_A_M1002_g N_A_c_81_n N_A_c_82_n
+ N_A_c_88_n N_A_M1000_g N_A_c_89_n N_A_M1001_g A A A N_A_c_85_n N_A_c_86_n
+ N_A_c_87_n PM_SKY130_FD_SC_HS__NOR2_2%A
x_PM_SKY130_FD_SC_HS__NOR2_2%A_35_368# N_A_35_368#_M1004_s N_A_35_368#_M1005_s
+ N_A_35_368#_M1001_s N_A_35_368#_c_126_n N_A_35_368#_c_127_n
+ N_A_35_368#_c_128_n N_A_35_368#_c_137_n N_A_35_368#_c_129_n
+ N_A_35_368#_c_130_n N_A_35_368#_c_131_n PM_SKY130_FD_SC_HS__NOR2_2%A_35_368#
x_PM_SKY130_FD_SC_HS__NOR2_2%Y N_Y_M1003_d N_Y_M1004_d N_Y_c_167_n Y Y Y
+ PM_SKY130_FD_SC_HS__NOR2_2%Y
x_PM_SKY130_FD_SC_HS__NOR2_2%VPWR N_VPWR_M1000_d N_VPWR_c_191_n N_VPWR_c_192_n
+ N_VPWR_c_193_n VPWR N_VPWR_c_194_n N_VPWR_c_190_n
+ PM_SKY130_FD_SC_HS__NOR2_2%VPWR
x_PM_SKY130_FD_SC_HS__NOR2_2%VGND N_VGND_M1003_s N_VGND_M1002_d N_VGND_c_217_n
+ N_VGND_c_218_n N_VGND_c_219_n VGND N_VGND_c_220_n N_VGND_c_221_n
+ N_VGND_c_222_n N_VGND_c_223_n PM_SKY130_FD_SC_HS__NOR2_2%VGND
cc_1 VNB N_B_c_40_n 0.0140756f $X=-0.19 $Y=-0.245 $X2=0.92 $Y2=1.69
cc_2 VNB N_B_c_41_n 0.0736776f $X=-0.19 $Y=-0.245 $X2=0.455 $Y2=1.385
cc_3 VNB N_B_c_42_n 0.0196224f $X=-0.19 $Y=-0.245 $X2=0.547 $Y2=1.22
cc_4 VNB B 0.0105321f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_5 VNB N_A_c_80_n 0.0173873f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=1.765
cc_6 VNB N_A_c_81_n 0.0177118f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=1.22
cc_7 VNB N_A_c_82_n 0.00722892f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=0.74
cc_8 VNB A 0.0193805f $X=-0.19 $Y=-0.245 $X2=0.455 $Y2=1.385
cc_9 VNB A 0.0201373f $X=-0.19 $Y=-0.245 $X2=0.547 $Y2=1.22
cc_10 VNB N_A_c_85_n 0.0955767f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=1.385
cc_11 VNB N_A_c_86_n 0.0910742f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=1.385
cc_12 VNB N_A_c_87_n 0.0251329f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_Y_c_167_n 0.00598888f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=1.765
cc_14 VNB N_VPWR_c_190_n 0.103974f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_VGND_c_217_n 0.0122168f $X=-0.19 $Y=-0.245 $X2=0.92 $Y2=1.69
cc_16 VNB N_VGND_c_218_n 0.0370023f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=1.765
cc_17 VNB N_VGND_c_219_n 0.0207786f $X=-0.19 $Y=-0.245 $X2=0.455 $Y2=1.385
cc_18 VNB N_VGND_c_220_n 0.0186948f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_19 VNB N_VGND_c_221_n 0.0282826f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_VGND_c_222_n 0.174237f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_VGND_c_223_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VPB N_B_c_40_n 0.0111346f $X=-0.19 $Y=1.66 $X2=0.92 $Y2=1.69
cc_23 VPB N_B_c_45_n 0.0145537f $X=-0.19 $Y=1.66 $X2=0.995 $Y2=1.765
cc_24 VPB N_B_c_41_n 0.00859226f $X=-0.19 $Y=1.66 $X2=0.455 $Y2=1.385
cc_25 VPB N_B_c_47_n 0.0181066f $X=-0.19 $Y=1.66 $X2=0.547 $Y2=1.765
cc_26 VPB N_A_c_88_n 0.0147219f $X=-0.19 $Y=1.66 $X2=0.565 $Y2=0.74
cc_27 VPB N_A_c_89_n 0.0196299f $X=-0.19 $Y=1.66 $X2=0.995 $Y2=1.765
cc_28 VPB N_A_c_86_n 0.016078f $X=-0.19 $Y=1.66 $X2=0.28 $Y2=1.385
cc_29 VPB N_A_35_368#_c_126_n 0.0419699f $X=-0.19 $Y=1.66 $X2=0.547 $Y2=1.385
cc_30 VPB N_A_35_368#_c_127_n 0.00523584f $X=-0.19 $Y=1.66 $X2=0.547 $Y2=1.765
cc_31 VPB N_A_35_368#_c_128_n 0.00935849f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.21
cc_32 VPB N_A_35_368#_c_129_n 0.0140223f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_33 VPB N_A_35_368#_c_130_n 0.00254452f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_34 VPB N_A_35_368#_c_131_n 0.042041f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_35 VPB N_VPWR_c_191_n 0.00571271f $X=-0.19 $Y=1.66 $X2=0.565 $Y2=0.74
cc_36 VPB N_VPWR_c_192_n 0.0387879f $X=-0.19 $Y=1.66 $X2=0.995 $Y2=1.765
cc_37 VPB N_VPWR_c_193_n 0.00460249f $X=-0.19 $Y=1.66 $X2=0.995 $Y2=2.4
cc_38 VPB N_VPWR_c_194_n 0.0201062f $X=-0.19 $Y=1.66 $X2=0.28 $Y2=1.385
cc_39 VPB N_VPWR_c_190_n 0.0608378f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_40 N_B_c_42_n N_A_c_80_n 0.00920383f $X=0.547 $Y=1.22 $X2=-0.19 $Y2=-0.245
cc_41 N_B_c_40_n N_A_c_82_n 0.0100444f $X=0.92 $Y=1.69 $X2=0 $Y2=0
cc_42 N_B_c_41_n N_A_c_82_n 0.00920383f $X=0.455 $Y=1.385 $X2=0 $Y2=0
cc_43 N_B_c_45_n N_A_c_88_n 0.00918371f $X=0.995 $Y=1.765 $X2=0 $Y2=0
cc_44 N_B_c_40_n N_A_c_86_n 0.00816756f $X=0.92 $Y=1.69 $X2=0 $Y2=0
cc_45 N_B_c_41_n N_A_c_86_n 0.00301946f $X=0.455 $Y=1.385 $X2=0 $Y2=0
cc_46 N_B_c_41_n N_A_35_368#_c_126_n 0.00185549f $X=0.455 $Y=1.385 $X2=0 $Y2=0
cc_47 N_B_c_47_n N_A_35_368#_c_126_n 0.00807154f $X=0.547 $Y=1.765 $X2=0 $Y2=0
cc_48 B N_A_35_368#_c_126_n 0.0149782f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_49 N_B_c_45_n N_A_35_368#_c_127_n 0.0121982f $X=0.995 $Y=1.765 $X2=0 $Y2=0
cc_50 N_B_c_47_n N_A_35_368#_c_127_n 0.013579f $X=0.547 $Y=1.765 $X2=0 $Y2=0
cc_51 N_B_c_45_n N_A_35_368#_c_137_n 0.00588035f $X=0.995 $Y=1.765 $X2=0 $Y2=0
cc_52 N_B_c_45_n N_A_35_368#_c_130_n 9.96784e-19 $X=0.995 $Y=1.765 $X2=0 $Y2=0
cc_53 N_B_c_40_n N_Y_c_167_n 0.0167438f $X=0.92 $Y=1.69 $X2=0 $Y2=0
cc_54 N_B_c_45_n N_Y_c_167_n 0.00129998f $X=0.995 $Y=1.765 $X2=0 $Y2=0
cc_55 N_B_c_41_n N_Y_c_167_n 0.0209871f $X=0.455 $Y=1.385 $X2=0 $Y2=0
cc_56 N_B_c_42_n N_Y_c_167_n 0.01725f $X=0.547 $Y=1.22 $X2=0 $Y2=0
cc_57 N_B_c_47_n N_Y_c_167_n 0.00286674f $X=0.547 $Y=1.765 $X2=0 $Y2=0
cc_58 B N_Y_c_167_n 0.0278923f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_59 N_B_c_45_n Y 0.00203343f $X=0.995 $Y=1.765 $X2=0 $Y2=0
cc_60 N_B_c_47_n Y 0.00253587f $X=0.547 $Y=1.765 $X2=0 $Y2=0
cc_61 N_B_c_45_n Y 0.010703f $X=0.995 $Y=1.765 $X2=0 $Y2=0
cc_62 N_B_c_47_n Y 0.010622f $X=0.547 $Y=1.765 $X2=0 $Y2=0
cc_63 N_B_c_45_n N_VPWR_c_192_n 0.00278271f $X=0.995 $Y=1.765 $X2=0 $Y2=0
cc_64 N_B_c_47_n N_VPWR_c_192_n 0.00278271f $X=0.547 $Y=1.765 $X2=0 $Y2=0
cc_65 N_B_c_45_n N_VPWR_c_190_n 0.00353907f $X=0.995 $Y=1.765 $X2=0 $Y2=0
cc_66 N_B_c_47_n N_VPWR_c_190_n 0.00357443f $X=0.547 $Y=1.765 $X2=0 $Y2=0
cc_67 N_B_c_41_n N_VGND_c_218_n 0.0022982f $X=0.455 $Y=1.385 $X2=0 $Y2=0
cc_68 N_B_c_42_n N_VGND_c_218_n 0.0161039f $X=0.547 $Y=1.22 $X2=0 $Y2=0
cc_69 B N_VGND_c_218_n 0.0283463f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_70 N_B_c_42_n N_VGND_c_220_n 0.00434272f $X=0.547 $Y=1.22 $X2=0 $Y2=0
cc_71 N_B_c_42_n N_VGND_c_222_n 0.00824032f $X=0.547 $Y=1.22 $X2=0 $Y2=0
cc_72 N_A_c_88_n N_A_35_368#_c_127_n 0.00125031f $X=1.445 $Y=1.765 $X2=0 $Y2=0
cc_73 N_A_c_88_n N_A_35_368#_c_137_n 0.00413798f $X=1.445 $Y=1.765 $X2=0 $Y2=0
cc_74 N_A_c_81_n N_A_35_368#_c_129_n 8.34335e-19 $X=1.355 $Y=1.26 $X2=0 $Y2=0
cc_75 N_A_c_88_n N_A_35_368#_c_129_n 0.0164228f $X=1.445 $Y=1.765 $X2=0 $Y2=0
cc_76 N_A_c_89_n N_A_35_368#_c_129_n 0.0137005f $X=1.895 $Y=1.765 $X2=0 $Y2=0
cc_77 A N_A_35_368#_c_129_n 0.0351284f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_78 N_A_c_86_n N_A_35_368#_c_129_n 0.0139189f $X=1.97 $Y=1.44 $X2=0 $Y2=0
cc_79 N_A_c_81_n N_A_35_368#_c_130_n 0.00332308f $X=1.355 $Y=1.26 $X2=0 $Y2=0
cc_80 N_A_c_88_n N_A_35_368#_c_131_n 7.87297e-19 $X=1.445 $Y=1.765 $X2=0 $Y2=0
cc_81 N_A_c_89_n N_A_35_368#_c_131_n 0.0134887f $X=1.895 $Y=1.765 $X2=0 $Y2=0
cc_82 N_A_c_80_n N_Y_c_167_n 0.0126271f $X=0.995 $Y=1.185 $X2=0 $Y2=0
cc_83 N_A_c_82_n N_Y_c_167_n 0.00958281f $X=1.07 $Y=1.26 $X2=0 $Y2=0
cc_84 N_A_c_86_n N_Y_c_167_n 0.00698924f $X=1.97 $Y=1.44 $X2=0 $Y2=0
cc_85 N_A_c_88_n N_VPWR_c_191_n 0.0131585f $X=1.445 $Y=1.765 $X2=0 $Y2=0
cc_86 N_A_c_89_n N_VPWR_c_191_n 0.00650058f $X=1.895 $Y=1.765 $X2=0 $Y2=0
cc_87 N_A_c_88_n N_VPWR_c_192_n 0.00413917f $X=1.445 $Y=1.765 $X2=0 $Y2=0
cc_88 N_A_c_89_n N_VPWR_c_194_n 0.00445602f $X=1.895 $Y=1.765 $X2=0 $Y2=0
cc_89 N_A_c_88_n N_VPWR_c_190_n 0.0081781f $X=1.445 $Y=1.765 $X2=0 $Y2=0
cc_90 N_A_c_89_n N_VPWR_c_190_n 0.00861084f $X=1.895 $Y=1.765 $X2=0 $Y2=0
cc_91 N_A_c_80_n N_VGND_c_219_n 0.0184907f $X=0.995 $Y=1.185 $X2=0 $Y2=0
cc_92 N_A_c_81_n N_VGND_c_219_n 0.00953674f $X=1.355 $Y=1.26 $X2=0 $Y2=0
cc_93 A N_VGND_c_219_n 0.0211138f $X=2.075 $Y=0.84 $X2=0 $Y2=0
cc_94 N_A_c_85_n N_VGND_c_219_n 0.0118488f $X=1.97 $Y=0.42 $X2=0 $Y2=0
cc_95 N_A_c_87_n N_VGND_c_219_n 0.0193455f $X=2.04 $Y=0.675 $X2=0 $Y2=0
cc_96 N_A_c_80_n N_VGND_c_220_n 0.00434272f $X=0.995 $Y=1.185 $X2=0 $Y2=0
cc_97 N_A_c_85_n N_VGND_c_221_n 0.00214182f $X=1.97 $Y=0.42 $X2=0 $Y2=0
cc_98 N_A_c_87_n N_VGND_c_221_n 0.0270748f $X=2.04 $Y=0.675 $X2=0 $Y2=0
cc_99 N_A_c_80_n N_VGND_c_222_n 0.00825157f $X=0.995 $Y=1.185 $X2=0 $Y2=0
cc_100 N_A_c_87_n N_VGND_c_222_n 0.0175158f $X=2.04 $Y=0.675 $X2=0 $Y2=0
cc_101 N_A_35_368#_c_127_n N_Y_M1004_d 0.00197722f $X=1.135 $Y=2.99 $X2=0 $Y2=0
cc_102 N_A_35_368#_c_130_n N_Y_c_167_n 0.012982f $X=1.305 $Y=1.86 $X2=0 $Y2=0
cc_103 N_A_35_368#_c_126_n Y 0.0614863f $X=0.32 $Y=1.985 $X2=0 $Y2=0
cc_104 N_A_35_368#_c_137_n Y 0.0535858f $X=1.22 $Y=1.985 $X2=0 $Y2=0
cc_105 N_A_35_368#_c_127_n Y 0.0167902f $X=1.135 $Y=2.99 $X2=0 $Y2=0
cc_106 N_A_35_368#_c_129_n N_VPWR_M1000_d 0.00222494f $X=1.955 $Y=1.86 $X2=-0.19
+ $Y2=1.66
cc_107 N_A_35_368#_c_127_n N_VPWR_c_191_n 0.0123543f $X=1.135 $Y=2.99 $X2=0
+ $Y2=0
cc_108 N_A_35_368#_c_137_n N_VPWR_c_191_n 0.0503418f $X=1.22 $Y=1.985 $X2=0
+ $Y2=0
cc_109 N_A_35_368#_c_129_n N_VPWR_c_191_n 0.0154248f $X=1.955 $Y=1.86 $X2=0
+ $Y2=0
cc_110 N_A_35_368#_c_131_n N_VPWR_c_191_n 0.0580287f $X=2.12 $Y=1.985 $X2=0
+ $Y2=0
cc_111 N_A_35_368#_c_127_n N_VPWR_c_192_n 0.0582805f $X=1.135 $Y=2.99 $X2=0
+ $Y2=0
cc_112 N_A_35_368#_c_128_n N_VPWR_c_192_n 0.0179217f $X=0.405 $Y=2.99 $X2=0
+ $Y2=0
cc_113 N_A_35_368#_c_131_n N_VPWR_c_194_n 0.0145938f $X=2.12 $Y=1.985 $X2=0
+ $Y2=0
cc_114 N_A_35_368#_c_127_n N_VPWR_c_190_n 0.0326824f $X=1.135 $Y=2.99 $X2=0
+ $Y2=0
cc_115 N_A_35_368#_c_128_n N_VPWR_c_190_n 0.00971942f $X=0.405 $Y=2.99 $X2=0
+ $Y2=0
cc_116 N_A_35_368#_c_131_n N_VPWR_c_190_n 0.0120466f $X=2.12 $Y=1.985 $X2=0
+ $Y2=0
cc_117 N_A_35_368#_c_129_n N_VGND_c_219_n 0.00427368f $X=1.955 $Y=1.86 $X2=0
+ $Y2=0
cc_118 N_A_35_368#_c_130_n N_VGND_c_219_n 0.00618439f $X=1.305 $Y=1.86 $X2=0
+ $Y2=0
cc_119 N_Y_c_167_n N_VGND_c_218_n 0.0255553f $X=0.78 $Y=0.515 $X2=0 $Y2=0
cc_120 N_Y_c_167_n N_VGND_c_219_n 0.0308485f $X=0.78 $Y=0.515 $X2=0 $Y2=0
cc_121 N_Y_c_167_n N_VGND_c_220_n 0.0144922f $X=0.78 $Y=0.515 $X2=0 $Y2=0
cc_122 N_Y_c_167_n N_VGND_c_222_n 0.0118826f $X=0.78 $Y=0.515 $X2=0 $Y2=0
