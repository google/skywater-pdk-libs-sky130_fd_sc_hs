* File: sky130_fd_sc_hs__dfstp_2.spice
* Created: Thu Aug 27 20:39:26 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hs__dfstp_2.pex.spice"
.subckt sky130_fd_sc_hs__dfstp_2  VNB VPB D CLK SET_B VPWR Q VGND
* 
* VGND	VGND
* Q	Q
* VPWR	VPWR
* SET_B	SET_B
* CLK	CLK
* D	D
* VPB	VPB
* VNB	VNB
MM1030 N_VGND_M1030_d N_D_M1030_g N_A_27_74#_M1030_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.1197 AS=0.1197 PD=1.41 PS=1.41 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1031 N_VGND_M1031_d N_CLK_M1031_g N_A_225_74#_M1031_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.2109 PD=1.02 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1018 N_A_398_74#_M1018_d N_A_225_74#_M1018_g N_VGND_M1031_d VNB NLOWVT L=0.15
+ W=0.74 AD=0.2109 AS=0.1036 PD=2.05 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.6 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1020 N_A_612_74#_M1020_d N_A_225_74#_M1020_g N_A_27_74#_M1020_s VNB NLOWVT
+ L=0.15 W=0.42 AD=0.14595 AS=0.18665 PD=1.115 PS=1.8 NRD=71.424 NRS=24.276 M=1
+ R=2.8 SA=75000.3 SB=75001.4 A=0.063 P=1.14 MULT=1
MM1015 A_781_74# N_A_398_74#_M1015_g N_A_612_74#_M1020_d VNB NLOWVT L=0.15
+ W=0.42 AD=0.0504 AS=0.14595 PD=0.66 PS=1.115 NRD=18.564 NRS=47.136 M=1 R=2.8
+ SA=75001.1 SB=75000.6 A=0.063 P=1.14 MULT=1
MM1022 N_VGND_M1022_d N_A_767_384#_M1022_g A_781_74# VNB NLOWVT L=0.15 W=0.42
+ AD=0.1197 AS=0.0504 PD=1.41 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75001.5
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1006 A_1057_118# N_A_612_74#_M1006_g N_A_767_384#_M1006_s VNB NLOWVT L=0.15
+ W=0.42 AD=0.0504 AS=0.1197 PD=0.66 PS=1.41 NRD=18.564 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75004.5 A=0.063 P=1.14 MULT=1
MM1021 N_VGND_M1021_d N_SET_B_M1021_g A_1057_118# VNB NLOWVT L=0.15 W=0.42
+ AD=0.120611 AS=0.0504 PD=0.954906 PS=0.66 NRD=38.568 NRS=18.564 M=1 R=2.8
+ SA=75000.6 SB=75004.1 A=0.063 P=1.14 MULT=1
MM1002 A_1278_74# N_A_612_74#_M1002_g N_VGND_M1021_d VNB NLOWVT L=0.15 W=0.64
+ AD=0.0768 AS=0.183789 PD=0.88 PS=1.45509 NRD=12.18 NRS=28.584 M=1 R=4.26667
+ SA=75000.9 SB=75002.4 A=0.096 P=1.58 MULT=1
MM1003 N_A_1356_74#_M1003_d N_A_398_74#_M1003_g A_1278_74# VNB NLOWVT L=0.15
+ W=0.64 AD=0.163804 AS=0.0768 PD=1.39472 PS=0.88 NRD=21.552 NRS=12.18 M=1
+ R=4.26667 SA=75001.3 SB=75002 A=0.096 P=1.58 MULT=1
MM1011 A_1489_118# N_A_225_74#_M1011_g N_A_1356_74#_M1003_d VNB NLOWVT L=0.15
+ W=0.42 AD=0.08085 AS=0.107496 PD=0.805 PS=0.915283 NRD=39.276 NRS=34.284 M=1
+ R=2.8 SA=75002.4 SB=75002.3 A=0.063 P=1.14 MULT=1
MM1028 A_1596_118# N_A_1566_92#_M1028_g A_1489_118# VNB NLOWVT L=0.15 W=0.42
+ AD=0.0882 AS=0.08085 PD=0.84 PS=0.805 NRD=44.28 NRS=39.276 M=1 R=2.8
+ SA=75002.9 SB=75001.8 A=0.063 P=1.14 MULT=1
MM1007 N_VGND_M1007_d N_SET_B_M1007_g A_1596_118# VNB NLOWVT L=0.15 W=0.42
+ AD=0.17955 AS=0.0882 PD=1.275 PS=0.84 NRD=0 NRS=44.28 M=1 R=2.8 SA=75003.5
+ SB=75001.2 A=0.063 P=1.14 MULT=1
MM1026 N_A_1566_92#_M1026_d N_A_1356_74#_M1026_g N_VGND_M1007_d VNB NLOWVT
+ L=0.15 W=0.42 AD=0.1197 AS=0.17955 PD=1.41 PS=1.275 NRD=0 NRS=19.992 M=1 R=2.8
+ SA=75004.5 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1016 N_VGND_M1016_d N_A_1356_74#_M1016_g N_A_2022_94#_M1016_s VNB NLOWVT
+ L=0.15 W=0.64 AD=0.144093 AS=0.1824 PD=1.08522 PS=1.85 NRD=15.468 NRS=0 M=1
+ R=4.26667 SA=75000.2 SB=75001.2 A=0.096 P=1.58 MULT=1
MM1008 N_VGND_M1016_d N_A_2022_94#_M1008_g N_Q_M1008_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.166607 AS=0.1036 PD=1.25478 PS=1.02 NRD=11.34 NRS=0 M=1 R=4.93333
+ SA=75000.7 SB=75000.7 A=0.111 P=1.78 MULT=1
MM1023 N_VGND_M1023_d N_A_2022_94#_M1023_g N_Q_M1008_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.2294 AS=0.1036 PD=2.1 PS=1.02 NRD=4.044 NRS=0 M=1 R=4.93333 SA=75001.2
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1000 N_VPWR_M1000_d N_D_M1000_g N_A_27_74#_M1000_s VPB PSHORT L=0.15 W=0.42
+ AD=0.1239 AS=0.1239 PD=1.43 PS=1.43 NRD=4.6886 NRS=4.6886 M=1 R=2.8 SA=75000.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1024 N_VPWR_M1024_d N_CLK_M1024_g N_A_225_74#_M1024_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.3304 PD=1.42 PS=2.83 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1029 N_A_398_74#_M1029_d N_A_225_74#_M1029_g N_VPWR_M1024_d VPB PSHORT L=0.15
+ W=1.12 AD=0.3304 AS=0.168 PD=2.83 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.7 SB=75000.2 A=0.168 P=2.54 MULT=1
MM1004 N_A_612_74#_M1004_d N_A_398_74#_M1004_g N_A_27_74#_M1004_s VPB PSHORT
+ L=0.15 W=0.42 AD=0.0735 AS=0.1239 PD=0.77 PS=1.43 NRD=28.1316 NRS=4.6886 M=1
+ R=2.8 SA=75000.2 SB=75004.6 A=0.063 P=1.14 MULT=1
MM1001 A_716_456# N_A_225_74#_M1001_g N_A_612_74#_M1004_d VPB PSHORT L=0.15
+ W=0.42 AD=0.0567 AS=0.0735 PD=0.69 PS=0.77 NRD=37.5088 NRS=4.6886 M=1 R=2.8
+ SA=75000.7 SB=75004.1 A=0.063 P=1.14 MULT=1
MM1017 N_VPWR_M1017_d N_A_767_384#_M1017_g A_716_456# VPB PSHORT L=0.15 W=0.42
+ AD=0.246825 AS=0.0567 PD=1.575 PS=0.69 NRD=86.7588 NRS=37.5088 M=1 R=2.8
+ SA=75001.1 SB=75003.7 A=0.063 P=1.14 MULT=1
MM1019 N_A_767_384#_M1019_d N_A_612_74#_M1019_g N_VPWR_M1017_d VPB PSHORT L=0.15
+ W=0.42 AD=0.063 AS=0.246825 PD=0.72 PS=1.575 NRD=0 NRS=249.835 M=1 R=2.8
+ SA=75002.3 SB=75002.6 A=0.063 P=1.14 MULT=1
MM1027 N_VPWR_M1027_d N_SET_B_M1027_g N_A_767_384#_M1019_d VPB PSHORT L=0.15
+ W=0.42 AD=0.14476 AS=0.063 PD=1.11211 PS=0.72 NRD=135.851 NRS=4.6886 M=1 R=2.8
+ SA=75002.7 SB=75002.1 A=0.063 P=1.14 MULT=1
MM1025 A_1266_341# N_A_612_74#_M1025_g N_VPWR_M1027_d VPB PSHORT L=0.15 W=1
+ AD=0.199812 AS=0.344665 PD=1.61 PS=2.64789 NRD=28.5256 NRS=57.0512 M=1
+ R=6.66667 SA=75001.6 SB=75000.9 A=0.15 P=2.3 MULT=1
MM1012 N_A_1356_74#_M1012_d N_A_225_74#_M1012_g A_1266_341# VPB PSHORT L=0.15
+ W=1 AD=0.303873 AS=0.199812 PD=2.28169 PS=1.61 NRD=22.9702 NRS=28.5256 M=1
+ R=6.66667 SA=75001.9 SB=75000.9 A=0.15 P=2.3 MULT=1
MM1032 A_1521_508# N_A_398_74#_M1032_g N_A_1356_74#_M1012_d VPB PSHORT L=0.15
+ W=0.42 AD=0.0567 AS=0.127627 PD=0.69 PS=0.95831 NRD=37.5088 NRS=80.9079 M=1
+ R=2.8 SA=75002.4 SB=75001.2 A=0.063 P=1.14 MULT=1
MM1009 N_VPWR_M1009_d N_A_1566_92#_M1009_g A_1521_508# VPB PSHORT L=0.15 W=0.42
+ AD=0.0819 AS=0.0567 PD=0.81 PS=0.69 NRD=46.886 NRS=37.5088 M=1 R=2.8
+ SA=75002.8 SB=75000.8 A=0.063 P=1.14 MULT=1
MM1014 N_A_1356_74#_M1014_d N_SET_B_M1014_g N_VPWR_M1009_d VPB PSHORT L=0.15
+ W=0.42 AD=0.1239 AS=0.0819 PD=1.43 PS=0.81 NRD=4.6886 NRS=4.6886 M=1 R=2.8
+ SA=75003.4 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1033 N_A_1566_92#_M1033_d N_A_1356_74#_M1033_g N_VPWR_M1033_s VPB PSHORT
+ L=0.15 W=0.42 AD=0.1239 AS=0.1239 PD=1.43 PS=1.43 NRD=4.6886 NRS=4.6886 M=1
+ R=2.8 SA=75000.2 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1013 N_VPWR_M1013_d N_A_1356_74#_M1013_g N_A_2022_94#_M1013_s VPB PSHORT
+ L=0.15 W=1 AD=0.198302 AS=0.295 PD=1.41981 PS=2.59 NRD=19.1878 NRS=1.9503 M=1
+ R=6.66667 SA=75000.2 SB=75001.2 A=0.15 P=2.3 MULT=1
MM1005 N_Q_M1005_d N_A_2022_94#_M1005_g N_VPWR_M1013_d VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.222098 PD=1.42 PS=1.59019 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.7 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1010 N_Q_M1005_d N_A_2022_94#_M1010_g N_VPWR_M1010_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.3304 PD=1.42 PS=2.83 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.1 SB=75000.2 A=0.168 P=2.54 MULT=1
DX34_noxref VNB VPB NWDIODE A=23.4057 P=28.75
c_1646 A_716_456# 0 1.50276e-19 $X=3.58 $Y=2.28
*
.include "sky130_fd_sc_hs__dfstp_2.pxi.spice"
*
.ends
*
*
