* NGSPICE file created from sky130_fd_sc_hs__a31o_2.ext - technology: sky130A

.subckt sky130_fd_sc_hs__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
M1000 VGND B1 a_97_296# VNB nlowvt w=740000u l=150000u
+  ad=9.435e+11p pd=6.99e+06u as=3.108e+11p ps=2.32e+06u
M1001 a_97_296# B1 a_362_368# VPB pshort w=1e+06u l=150000u
+  ad=3.05e+11p pd=2.61e+06u as=6.5e+11p ps=5.3e+06u
M1002 a_371_74# A3 VGND VNB nlowvt w=740000u l=150000u
+  ad=1.776e+11p pd=1.96e+06u as=0p ps=0u
M1003 a_362_368# A1 VPWR VPB pshort w=1e+06u l=150000u
+  ad=0p pd=0u as=1.4332e+12p ps=9.17e+06u
M1004 a_449_74# A2 a_371_74# VNB nlowvt w=740000u l=150000u
+  ad=3.108e+11p pd=2.32e+06u as=0p ps=0u
M1005 VGND a_97_296# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.072e+11p ps=2.04e+06u
M1006 X a_97_296# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_97_296# A1 a_449_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 X a_97_296# VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=3.36e+11p pd=2.84e+06u as=0p ps=0u
M1009 VPWR a_97_296# X VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_362_368# A3 VPWR VPB pshort w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VPWR A2 a_362_368# VPB pshort w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

