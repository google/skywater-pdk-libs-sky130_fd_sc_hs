* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hs__sdfrtp_1 CLK D RESET_B SCD SCE VGND VNB VPB VPWR Q
M1000 a_1319_118# a_1034_368# a_1233_118# VNB nlowvt w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=1.176e+11p ps=1.4e+06u
M1001 a_1367_92# a_1233_118# VPWR VPB pshort w=1e+06u l=150000u
+  ad=3e+11p pd=2.6e+06u as=2.23208e+12p ps=1.888e+07u
M1002 VPWR a_1367_92# a_1343_461# VPB pshort w=420000u l=150000u
+  ad=0p pd=0u as=1.134e+11p ps=1.38e+06u
M1003 a_1034_368# a_855_368# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=1.4802e+12p ps=1.325e+07u
M1004 a_1745_74# a_855_368# a_1367_92# VPB pshort w=1e+06u l=150000u
+  ad=4.42975e+11p pd=3.64e+06u as=0p ps=0u
M1005 VGND a_1997_272# a_1972_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=8.82e+10p ps=1.26e+06u
M1006 VPWR SCD a_538_464# VPB pshort w=640000u l=150000u
+  ad=0p pd=0u as=1.728e+11p ps=1.82e+06u
M1007 a_1972_74# a_855_368# a_1745_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=4.687e+11p ps=3.25e+06u
M1008 VGND CLK a_855_368# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1009 a_1233_118# a_855_368# a_300_464# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=3.822e+11p ps=3.5e+06u
M1010 a_1745_74# a_1034_368# a_1367_92# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=1.792e+11p ps=1.84e+06u
M1011 Q a_2399_424# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1012 a_312_81# a_27_88# a_225_81# VNB nlowvt w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=3.15e+11p ps=3.18e+06u
M1013 a_300_464# D a_312_81# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 VPWR a_1997_272# a_1993_508# VPB pshort w=420000u l=150000u
+  ad=0p pd=0u as=1.134e+11p ps=1.38e+06u
M1015 a_1997_272# RESET_B VPWR VPB pshort w=420000u l=150000u
+  ad=1.26e+11p pd=1.44e+06u as=0p ps=0u
M1016 VGND RESET_B a_225_81# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_2399_424# a_1745_74# VPWR VPB pshort w=840000u l=150000u
+  ad=2.478e+11p pd=2.27e+06u as=0p ps=0u
M1018 VPWR a_1745_74# a_1997_272# VPB pshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VGND RESET_B a_1397_118# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1020 a_216_464# SCE VPWR VPB pshort w=640000u l=150000u
+  ad=1.728e+11p pd=1.82e+06u as=0p ps=0u
M1021 a_225_81# SCD a_545_81# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1022 VPWR CLK a_855_368# VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=3.304e+11p ps=2.83e+06u
M1023 VPWR SCE a_27_88# VPB pshort w=640000u l=150000u
+  ad=0p pd=0u as=1.888e+11p ps=1.87e+06u
M1024 a_538_464# a_27_88# a_300_464# VPB pshort w=640000u l=150000u
+  ad=0p pd=0u as=9.783e+11p ps=6.66e+06u
M1025 a_1993_508# a_1034_368# a_1745_74# VPB pshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 a_1233_118# a_1034_368# a_300_464# VPB pshort w=420000u l=150000u
+  ad=2.765e+11p pd=3.02e+06u as=0p ps=0u
M1027 a_1397_118# a_1367_92# a_1319_118# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1028 a_1997_272# a_1745_74# a_2135_74# VNB nlowvt w=420000u l=150000u
+  ad=1.197e+11p pd=1.41e+06u as=8.82e+10p ps=1.26e+06u
M1029 a_1034_368# a_855_368# VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=3.304e+11p pd=2.83e+06u as=0p ps=0u
M1030 a_545_81# SCE a_300_464# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1031 a_2399_424# a_1745_74# VGND VNB nlowvt w=550000u l=150000u
+  ad=1.5675e+11p pd=1.67e+06u as=0p ps=0u
M1032 a_1343_461# a_855_368# a_1233_118# VPB pshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1033 a_1367_92# a_1233_118# VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1034 a_1233_118# RESET_B VPWR VPB pshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1035 Q a_2399_424# VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=3.304e+11p pd=2.83e+06u as=0p ps=0u
M1036 a_300_464# D a_216_464# VPB pshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1037 VGND SCE a_27_88# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.197e+11p ps=1.41e+06u
M1038 a_2135_74# RESET_B VGND VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1039 a_300_464# RESET_B VPWR VPB pshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
