* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hs__o21a_4 A1 A2 B1 VGND VNB VPB VPWR X
M1000 VPWR a_216_387# X VPB pshort w=1.12e+06u l=150000u
+  ad=2.0608e+12p pd=1.474e+07u as=6.72e+11p ps=5.68e+06u
M1001 VGND a_216_387# X VNB nlowvt w=740000u l=150000u
+  ad=1.1573e+12p pd=1.034e+07u as=4.144e+11p ps=4.08e+06u
M1002 X a_216_387# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1003 VPWR B1 a_216_387# VPB pshort w=840000u l=150000u
+  ad=0p pd=0u as=6.192e+11p ps=5.04e+06u
M1004 a_216_387# B1 VPWR VPB pshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_27_125# A2 VGND VNB nlowvt w=640000u l=150000u
+  ad=7.744e+11p pd=7.54e+06u as=0p ps=0u
M1006 VGND A2 a_27_125# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 X a_216_387# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VGND a_216_387# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_27_125# B1 a_216_387# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=1.792e+11p ps=1.84e+06u
M1010 VGND A1 a_27_125# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 X a_216_387# VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_27_125# A1 VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 X a_216_387# VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_216_387# B1 a_27_125# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_216_387# A2 a_116_387# VPB pshort w=1e+06u l=150000u
+  ad=0p pd=0u as=7e+11p ps=5.4e+06u
M1016 VPWR a_216_387# X VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 VPWR A1 a_116_387# VPB pshort w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_116_387# A2 a_216_387# VPB pshort w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_116_387# A1 VPWR VPB pshort w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
