* File: sky130_fd_sc_hs__or3b_1.spice
* Created: Thu Aug 27 21:06:13 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hs__or3b_1.pex.spice"
.subckt sky130_fd_sc_hs__or3b_1  VNB VPB C_N B A VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A	A
* B	B
* C_N	C_N
* VPB	VPB
* VNB	VNB
MM1008 N_A_124_424#_M1008_d N_C_N_M1008_g N_VGND_M1008_s VNB NLOWVT L=0.15
+ W=0.55 AD=0.1595 AS=0.1925 PD=1.68 PS=1.8 NRD=1.08 NRS=14.172 M=1 R=3.66667
+ SA=75000.3 SB=75000.2 A=0.0825 P=1.4 MULT=1
MM1004 N_VGND_M1004_d N_A_124_424#_M1004_g N_A_239_74#_M1004_s VNB NLOWVT L=0.15
+ W=0.55 AD=0.1155 AS=0.15675 PD=0.97 PS=1.67 NRD=15.264 NRS=0 M=1 R=3.66667
+ SA=75000.2 SB=75002 A=0.0825 P=1.4 MULT=1
MM1000 N_A_239_74#_M1000_d N_B_M1000_g N_VGND_M1004_d VNB NLOWVT L=0.15 W=0.55
+ AD=0.086625 AS=0.1155 PD=0.865 PS=0.97 NRD=0 NRS=15.264 M=1 R=3.66667
+ SA=75000.8 SB=75001.4 A=0.0825 P=1.4 MULT=1
MM1003 N_VGND_M1003_d N_A_M1003_g N_A_239_74#_M1000_d VNB NLOWVT L=0.15 W=0.55
+ AD=0.162122 AS=0.086625 PD=1.1469 PS=0.865 NRD=31.632 NRS=7.632 M=1 R=3.66667
+ SA=75001.2 SB=75001 A=0.0825 P=1.4 MULT=1
MM1006 N_X_M1006_d N_A_239_74#_M1006_g N_VGND_M1003_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.218128 PD=2.05 PS=1.5431 NRD=0 NRS=29.184 M=1 R=4.93333
+ SA=75001.5 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1001 N_A_124_424#_M1001_d N_C_N_M1001_g N_VPWR_M1001_s VPB PSHORT L=0.15
+ W=0.84 AD=0.2562 AS=0.2814 PD=2.29 PS=2.35 NRD=4.6886 NRS=11.7215 M=1 R=5.6
+ SA=75000.3 SB=75000.2 A=0.126 P=1.98 MULT=1
MM1002 A_368_391# N_A_124_424#_M1002_g N_A_239_74#_M1002_s VPB PSHORT L=0.15 W=1
+ AD=0.135 AS=0.295 PD=1.27 PS=2.59 NRD=15.7403 NRS=1.9503 M=1 R=6.66667
+ SA=75000.2 SB=75001.6 A=0.15 P=2.3 MULT=1
MM1007 A_452_391# N_B_M1007_g A_368_391# VPB PSHORT L=0.15 W=1 AD=0.135 AS=0.135
+ PD=1.27 PS=1.27 NRD=15.7403 NRS=15.7403 M=1 R=6.66667 SA=75000.6 SB=75001.2
+ A=0.15 P=2.3 MULT=1
MM1009 N_VPWR_M1009_d N_A_M1009_g A_452_391# VPB PSHORT L=0.15 W=1 AD=0.224717
+ AS=0.135 PD=1.46698 PS=1.27 NRD=18.715 NRS=15.7403 M=1 R=6.66667 SA=75001.1
+ SB=75000.8 A=0.15 P=2.3 MULT=1
MM1005 N_X_M1005_d N_A_239_74#_M1005_g N_VPWR_M1009_d VPB PSHORT L=0.15 W=1.12
+ AD=0.3304 AS=0.251683 PD=2.83 PS=1.64302 NRD=1.7533 NRS=10.5395 M=1 R=7.46667
+ SA=75001.5 SB=75000.2 A=0.168 P=2.54 MULT=1
DX10_noxref VNB VPB NWDIODE A=7.8492 P=12.16
*
.include "sky130_fd_sc_hs__or3b_1.pxi.spice"
*
.ends
*
*
