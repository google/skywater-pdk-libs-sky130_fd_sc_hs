* File: sky130_fd_sc_hs__dlxtn_2.spice
* Created: Tue Sep  1 20:03:03 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hs__dlxtn_2.pex.spice"
.subckt sky130_fd_sc_hs__dlxtn_2  VNB VPB D GATE_N VPWR Q VGND
* 
* VGND	VGND
* Q	Q
* VPWR	VPWR
* GATE_N	GATE_N
* D	D
* VPB	VPB
* VNB	VNB
MM1017 N_VGND_M1017_d N_D_M1017_g N_A_27_120#_M1017_s VNB NLOWVT L=0.15 W=0.55
+ AD=0.161184 AS=0.15675 PD=1.20233 PS=1.67 NRD=51.936 NRS=0 M=1 R=3.66667
+ SA=75000.2 SB=75000.8 A=0.0825 P=1.4 MULT=1
MM1003 N_A_232_82#_M1003_d N_GATE_N_M1003_g N_VGND_M1017_d VNB NLOWVT L=0.15
+ W=0.74 AD=0.2109 AS=0.216866 PD=2.05 PS=1.61767 NRD=0 NRS=38.604 M=1 R=4.93333
+ SA=75000.7 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1009 N_VGND_M1009_d N_A_232_82#_M1009_g N_A_369_392#_M1009_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.25707 AS=0.2109 PD=1.55507 PS=2.05 NRD=66.48 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75002 A=0.111 P=1.78 MULT=1
MM1002 A_658_79# N_A_27_120#_M1002_g N_VGND_M1009_d VNB NLOWVT L=0.15 W=0.64
+ AD=0.0768 AS=0.22233 PD=0.88 PS=1.34493 NRD=12.18 NRS=3.744 M=1 R=4.26667
+ SA=75001.1 SB=75001.4 A=0.096 P=1.58 MULT=1
MM1001 N_A_669_392#_M1001_d N_A_232_82#_M1001_g A_658_79# VNB NLOWVT L=0.15
+ W=0.64 AD=0.169238 AS=0.0768 PD=1.52755 PS=0.88 NRD=24.372 NRS=12.18 M=1
+ R=4.26667 SA=75001.5 SB=75001 A=0.096 P=1.58 MULT=1
MM1015 A_875_139# N_A_369_392#_M1015_g N_A_669_392#_M1001_d VNB NLOWVT L=0.15
+ W=0.42 AD=0.0504 AS=0.111062 PD=0.66 PS=1.00245 NRD=18.564 NRS=38.568 M=1
+ R=2.8 SA=75001.8 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1005 N_VGND_M1005_d N_A_842_405#_M1005_g A_875_139# VNB NLOWVT L=0.15 W=0.42
+ AD=0.0877655 AS=0.0504 PD=0.796552 PS=0.66 NRD=22.848 NRS=18.564 M=1 R=2.8
+ SA=75002.2 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1014 N_A_842_405#_M1014_d N_A_669_392#_M1014_g N_VGND_M1005_d VNB NLOWVT
+ L=0.15 W=0.74 AD=0.2109 AS=0.154634 PD=2.05 PS=1.40345 NRD=0 NRS=0 M=1
+ R=4.93333 SA=75001.6 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1000 N_Q_M1000_d N_A_842_405#_M1000_g N_VGND_M1000_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1258 AS=0.2109 PD=1.08 PS=2.05 NRD=0.804 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75000.7 A=0.111 P=1.78 MULT=1
MM1012 N_Q_M1000_d N_A_842_405#_M1012_g N_VGND_M1012_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1258 AS=0.2294 PD=1.08 PS=2.1 NRD=8.916 NRS=4.044 M=1 R=4.93333
+ SA=75000.7 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1008 N_VPWR_M1008_d N_D_M1008_g N_A_27_120#_M1008_s VPB PSHORT L=0.15 W=0.84
+ AD=0.168 AS=0.2478 PD=1.24 PS=2.27 NRD=14.0658 NRS=2.3443 M=1 R=5.6 SA=75000.2
+ SB=75000.8 A=0.126 P=1.98 MULT=1
MM1004 N_A_232_82#_M1004_d N_GATE_N_M1004_g N_VPWR_M1008_d VPB PSHORT L=0.15
+ W=0.84 AD=0.2478 AS=0.168 PD=2.27 PS=1.24 NRD=2.3443 NRS=14.0658 M=1 R=5.6
+ SA=75000.8 SB=75000.2 A=0.126 P=1.98 MULT=1
MM1006 N_VPWR_M1006_d N_A_232_82#_M1006_g N_A_369_392#_M1006_s VPB PSHORT L=0.15
+ W=0.84 AD=0.23294 AS=0.2478 PD=1.47457 PS=2.27 NRD=52.1262 NRS=2.3443 M=1
+ R=5.6 SA=75000.2 SB=75002 A=0.126 P=1.98 MULT=1
MM1016 A_585_392# N_A_27_120#_M1016_g N_VPWR_M1006_d VPB PSHORT L=0.15 W=1
+ AD=0.135 AS=0.27731 PD=1.27 PS=1.75543 NRD=15.7403 NRS=21.6503 M=1 R=6.66667
+ SA=75000.8 SB=75001.5 A=0.15 P=2.3 MULT=1
MM1018 N_A_669_392#_M1018_d N_A_369_392#_M1018_g A_585_392# VPB PSHORT L=0.15
+ W=1 AD=0.285335 AS=0.135 PD=2.05634 PS=1.27 NRD=8.8453 NRS=15.7403 M=1
+ R=6.66667 SA=75001.2 SB=75001.1 A=0.15 P=2.3 MULT=1
MM1010 A_791_503# N_A_232_82#_M1010_g N_A_669_392#_M1018_d VPB PSHORT L=0.15
+ W=0.42 AD=0.0567 AS=0.11984 PD=0.69 PS=0.863662 NRD=37.5088 NRS=63.3158 M=1
+ R=2.8 SA=75001.7 SB=75001.5 A=0.063 P=1.14 MULT=1
MM1013 N_VPWR_M1013_d N_A_842_405#_M1013_g A_791_503# VPB PSHORT L=0.15 W=0.42
+ AD=0.135355 AS=0.0567 PD=1.01455 PS=0.69 NRD=4.6886 NRS=37.5088 M=1 R=2.8
+ SA=75002.1 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1019 N_A_842_405#_M1019_d N_A_669_392#_M1019_g N_VPWR_M1013_d VPB PSHORT
+ L=0.15 W=1.12 AD=0.3304 AS=0.360945 PD=2.83 PS=2.70545 NRD=1.7533 NRS=2.6201
+ M=1 R=7.46667 SA=75001.3 SB=75000.2 A=0.168 P=2.54 MULT=1
MM1007 N_Q_M1007_d N_A_842_405#_M1007_g N_VPWR_M1007_s VPB PSHORT L=0.15 W=1.12
+ AD=0.1932 AS=0.3304 PD=1.465 PS=2.83 NRD=5.2599 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1011 N_Q_M1007_d N_A_842_405#_M1011_g N_VPWR_M1011_s VPB PSHORT L=0.15 W=1.12
+ AD=0.1932 AS=0.3304 PD=1.465 PS=2.83 NRD=6.1464 NRS=1.7533 M=1 R=7.46667
+ SA=75000.7 SB=75000.2 A=0.168 P=2.54 MULT=1
DX20_noxref VNB VPB NWDIODE A=14.1255 P=18.93
c_75 VNB 0 1.98766e-19 $X=0 $Y=0
c_972 A_658_79# 0 3.15497e-20 $X=3.29 $Y=0.395
*
.include "sky130_fd_sc_hs__dlxtn_2.pxi.spice"
*
.ends
*
*
