* File: sky130_fd_sc_hs__dfbbn_1.pex.spice
* Created: Tue Sep  1 19:59:21 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HS__DFBBN_1%CLK_N 3 5 7 8 12
c31 5 0 1.54433e-19 $X=0.495 $Y=1.765
r32 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.33
+ $Y=1.465 $X2=0.33 $Y2=1.465
r33 8 12 6.22942 $w=3.68e-07 $l=2e-07 $layer=LI1_cond $X=0.31 $Y=1.665 $X2=0.31
+ $Y2=1.465
r34 5 11 57.3754 $w=3.5e-07 $l=3.54965e-07 $layer=POLY_cond $X=0.495 $Y=1.765
+ $X2=0.375 $Y2=1.465
r35 5 7 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.495 $Y=1.765
+ $X2=0.495 $Y2=2.4
r36 1 11 38.7839 $w=3.5e-07 $l=2.16852e-07 $layer=POLY_cond $X=0.495 $Y=1.3
+ $X2=0.375 $Y2=1.465
r37 1 3 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=0.495 $Y=1.3 $X2=0.495
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HS__DFBBN_1%D 3 6 7 9 10 11 18
r43 16 18 13.9889 $w=3.3e-07 $l=8e-08 $layer=POLY_cond $X=2.01 $Y=1.345 $X2=2.09
+ $Y2=1.345
r44 14 16 16.6118 $w=3.3e-07 $l=9.5e-08 $layer=POLY_cond $X=1.915 $Y=1.345
+ $X2=2.01 $Y2=1.345
r45 10 11 19.2074 $w=3.28e-07 $l=5.5e-07 $layer=LI1_cond $X=2.09 $Y=1.345
+ $X2=2.64 $Y2=1.345
r46 10 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.09
+ $Y=1.345 $X2=2.09 $Y2=1.345
r47 7 9 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=2.01 $Y=2.44 $X2=2.01
+ $Y2=2.725
r48 6 7 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=2.01 $Y=2.35 $X2=2.01
+ $Y2=2.44
r49 5 16 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=2.01 $Y=1.51
+ $X2=2.01 $Y2=1.345
r50 5 6 326.516 $w=1.8e-07 $l=8.4e-07 $layer=POLY_cond $X=2.01 $Y=1.51 $X2=2.01
+ $Y2=2.35
r51 1 14 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.915 $Y=1.18
+ $X2=1.915 $Y2=1.345
r52 1 3 192.287 $w=1.5e-07 $l=3.75e-07 $layer=POLY_cond $X=1.915 $Y=1.18
+ $X2=1.915 $Y2=0.805
.ends

.subckt PM_SKY130_FD_SC_HS__DFBBN_1%A_474_405# 1 2 3 12 14 16 19 21 23 25 26 27
+ 29 30 31 32 36 38 42 49 55 60
c170 14 0 1.49698e-19 $X=2.61 $Y=2.44
r171 46 49 6.46067 $w=3.28e-07 $l=1.85e-07 $layer=LI1_cond $X=2.535 $Y=2.19
+ $X2=2.72 $Y2=2.19
r172 46 47 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.535
+ $Y=2.19 $X2=2.535 $Y2=2.19
r173 42 43 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.285
+ $Y=1.795 $X2=6.285 $Y2=1.795
r174 40 42 18.3343 $w=3.28e-07 $l=5.25e-07 $layer=LI1_cond $X=6.285 $Y=2.32
+ $X2=6.285 $Y2=1.795
r175 39 60 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.82 $Y=2.405
+ $X2=5.695 $Y2=2.405
r176 38 40 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=6.12 $Y=2.405
+ $X2=6.285 $Y2=2.32
r177 38 39 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=6.12 $Y=2.405
+ $X2=5.82 $Y2=2.405
r178 34 60 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.695 $Y=2.49
+ $X2=5.695 $Y2=2.405
r179 34 36 14.9818 $w=2.48e-07 $l=3.25e-07 $layer=LI1_cond $X=5.695 $Y=2.49
+ $X2=5.695 $Y2=2.815
r180 32 60 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.57 $Y=2.405
+ $X2=5.695 $Y2=2.405
r181 32 55 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=5.57 $Y=2.405
+ $X2=4.815 $Y2=2.405
r182 31 55 5.18835 $w=1.83e-07 $l=8.5e-08 $layer=LI1_cond $X=4.73 $Y=2.397
+ $X2=4.815 $Y2=2.397
r183 31 52 21.8821 $w=1.83e-07 $l=3.65e-07 $layer=LI1_cond $X=4.73 $Y=2.397
+ $X2=4.365 $Y2=2.397
r184 30 58 8.61582 $w=3.54e-07 $l=3.44601e-07 $layer=LI1_cond $X=4.73 $Y=1.165
+ $X2=4.98 $Y2=0.94
r185 30 31 74.3743 $w=1.68e-07 $l=1.14e-06 $layer=LI1_cond $X=4.73 $Y=1.165
+ $X2=4.73 $Y2=2.305
r186 29 52 14.4928 $w=3.28e-07 $l=4.15e-07 $layer=LI1_cond $X=4.365 $Y=2.905
+ $X2=4.365 $Y2=2.49
r187 26 29 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.2 $Y=2.99
+ $X2=4.365 $Y2=2.905
r188 26 27 91.0107 $w=1.68e-07 $l=1.395e-06 $layer=LI1_cond $X=4.2 $Y=2.99
+ $X2=2.805 $Y2=2.99
r189 25 27 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.72 $Y=2.905
+ $X2=2.805 $Y2=2.99
r190 24 49 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.72 $Y=2.355
+ $X2=2.72 $Y2=2.19
r191 24 25 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=2.72 $Y=2.355
+ $X2=2.72 $Y2=2.905
r192 21 43 50.756 $w=3.39e-07 $l=2.95804e-07 $layer=POLY_cond $X=6.41 $Y=2.045
+ $X2=6.31 $Y2=1.795
r193 21 23 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=6.41 $Y=2.045
+ $X2=6.41 $Y2=2.54
r194 17 43 38.6704 $w=3.39e-07 $l=2.14942e-07 $layer=POLY_cond $X=6.195 $Y=1.63
+ $X2=6.31 $Y2=1.795
r195 17 19 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=6.195 $Y=1.63
+ $X2=6.195 $Y2=0.87
r196 14 47 52.2586 $w=2.99e-07 $l=2.85044e-07 $layer=POLY_cond $X=2.61 $Y=2.44
+ $X2=2.535 $Y2=2.19
r197 14 16 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=2.61 $Y=2.44
+ $X2=2.61 $Y2=2.725
r198 10 47 38.5562 $w=2.99e-07 $l=1.67481e-07 $layer=POLY_cond $X=2.54 $Y=2.025
+ $X2=2.535 $Y2=2.19
r199 10 12 625.574 $w=1.5e-07 $l=1.22e-06 $layer=POLY_cond $X=2.54 $Y=2.025
+ $X2=2.54 $Y2=0.805
r200 3 60 600 $w=1.7e-07 $l=3.52101e-07 $layer=licon1_PDIFF $count=1 $X=5.505
+ $Y=2.12 $X2=5.655 $Y2=2.405
r201 3 36 600 $w=1.7e-07 $l=7.66339e-07 $layer=licon1_PDIFF $count=1 $X=5.505
+ $Y=2.12 $X2=5.655 $Y2=2.815
r202 2 52 300 $w=1.7e-07 $l=3.28634e-07 $layer=licon1_PDIFF $count=2 $X=4.235
+ $Y=2.12 $X2=4.365 $Y2=2.39
r203 1 58 182 $w=1.7e-07 $l=3.756e-07 $layer=licon1_NDIFF $count=1 $X=4.77
+ $Y=0.595 $X2=4.98 $Y2=0.88
.ends

.subckt PM_SKY130_FD_SC_HS__DFBBN_1%A_200_74# 1 2 7 9 12 13 15 16 18 22 25 29 30
+ 32 33 34 36 39 42 44 49 53 54 55 56 57 58 64 69 70 71 76
c221 76 0 1.02788e-19 $X=7.98 $Y=1.395
c222 70 0 5.14108e-20 $X=3.35 $Y=1.29
c223 58 0 7.83046e-20 $X=3.265 $Y=1.295
c224 57 0 7.98666e-20 $X=6.815 $Y=1.295
c225 56 0 1.63798e-20 $X=3.107 $Y=1.77
c226 53 0 1.54433e-19 $X=1.17 $Y=1.985
c227 36 0 9.67413e-20 $X=3.107 $Y=1.685
c228 34 0 1.55193e-19 $X=2.125 $Y=1.77
c229 16 0 1.47104e-19 $X=7.98 $Y=1.23
c230 13 0 1.06589e-20 $X=6.8 $Y=2.045
r231 69 71 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.35 $Y=1.29
+ $X2=3.35 $Y2=1.125
r232 69 70 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.35
+ $Y=1.29 $X2=3.35 $Y2=1.29
r233 64 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=1.295
+ $X2=6.96 $Y2=1.295
r234 61 70 8.03218 $w=3.28e-07 $l=2.3e-07 $layer=LI1_cond $X=3.12 $Y=1.29
+ $X2=3.35 $Y2=1.29
r235 61 78 0.453993 $w=3.28e-07 $l=1.3e-08 $layer=LI1_cond $X=3.12 $Y=1.29
+ $X2=3.107 $Y2=1.29
r236 60 61 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=1.295
+ $X2=3.12 $Y2=1.295
r237 58 60 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.265 $Y=1.295
+ $X2=3.12 $Y2=1.295
r238 57 64 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.815 $Y=1.295
+ $X2=6.96 $Y2=1.295
r239 57 58 4.39356 $w=1.4e-07 $l=3.55e-06 $layer=MET1_cond $X=6.815 $Y=1.295
+ $X2=3.265 $Y2=1.295
r240 54 55 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.33 $Y=1.82
+ $X2=1.33 $Y2=1.13
r241 53 54 8.69073 $w=4.08e-07 $l=1.65e-07 $layer=LI1_cond $X=1.21 $Y=1.985
+ $X2=1.21 $Y2=1.82
r242 50 76 35.8466 $w=3.3e-07 $l=2.05e-07 $layer=POLY_cond $X=7.775 $Y=1.395
+ $X2=7.98 $Y2=1.395
r243 49 50 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.775
+ $Y=1.395 $X2=7.775 $Y2=1.395
r244 47 65 3.34605 $w=3.8e-07 $l=1.83e-07 $layer=LI1_cond $X=7.075 $Y=1.37
+ $X2=6.892 $Y2=1.37
r245 47 49 21.2292 $w=3.78e-07 $l=7e-07 $layer=LI1_cond $X=7.075 $Y=1.37
+ $X2=7.775 $Y2=1.37
r246 44 45 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.875
+ $Y=1.765 $X2=6.875 $Y2=1.765
r247 42 65 3.47404 $w=3.65e-07 $l=1.9e-07 $layer=LI1_cond $X=6.892 $Y=1.56
+ $X2=6.892 $Y2=1.37
r248 42 44 6.47263 $w=3.63e-07 $l=2.05e-07 $layer=LI1_cond $X=6.892 $Y=1.56
+ $X2=6.892 $Y2=1.765
r249 39 40 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.075
+ $Y=2.19 $X2=3.075 $Y2=2.19
r250 37 56 3.52026 $w=2.65e-07 $l=8.5e-08 $layer=LI1_cond $X=3.107 $Y=1.855
+ $X2=3.107 $Y2=1.77
r251 37 39 14.5686 $w=2.63e-07 $l=3.35e-07 $layer=LI1_cond $X=3.107 $Y=1.855
+ $X2=3.107 $Y2=2.19
r252 36 56 3.52026 $w=2.65e-07 $l=8.5e-08 $layer=LI1_cond $X=3.107 $Y=1.685
+ $X2=3.107 $Y2=1.77
r253 35 78 2.04284 $w=2.65e-07 $l=1.65e-07 $layer=LI1_cond $X=3.107 $Y=1.455
+ $X2=3.107 $Y2=1.29
r254 35 36 10.0023 $w=2.63e-07 $l=2.3e-07 $layer=LI1_cond $X=3.107 $Y=1.455
+ $X2=3.107 $Y2=1.685
r255 33 56 2.98021 $w=1.7e-07 $l=1.32e-07 $layer=LI1_cond $X=2.975 $Y=1.77
+ $X2=3.107 $Y2=1.77
r256 33 34 55.4545 $w=1.68e-07 $l=8.5e-07 $layer=LI1_cond $X=2.975 $Y=1.77
+ $X2=2.125 $Y2=1.77
r257 31 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.04 $Y=1.855
+ $X2=2.125 $Y2=1.77
r258 31 32 68.5027 $w=1.68e-07 $l=1.05e-06 $layer=LI1_cond $X=2.04 $Y=1.855
+ $X2=2.04 $Y2=2.905
r259 29 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.955 $Y=2.99
+ $X2=2.04 $Y2=2.905
r260 29 30 35.2299 $w=1.68e-07 $l=5.4e-07 $layer=LI1_cond $X=1.955 $Y=2.99
+ $X2=1.415 $Y2=2.99
r261 23 55 8.99121 $w=3.58e-07 $l=1.8e-07 $layer=LI1_cond $X=1.235 $Y=0.95
+ $X2=1.235 $Y2=1.13
r262 23 25 13.9254 $w=3.58e-07 $l=4.35e-07 $layer=LI1_cond $X=1.235 $Y=0.95
+ $X2=1.235 $Y2=0.515
r263 20 30 8.45803 $w=1.7e-07 $l=2.43824e-07 $layer=LI1_cond $X=1.21 $Y=2.905
+ $X2=1.415 $Y2=2.99
r264 20 22 2.52975 $w=4.08e-07 $l=9e-08 $layer=LI1_cond $X=1.21 $Y=2.905
+ $X2=1.21 $Y2=2.815
r265 19 53 1.12433 $w=4.08e-07 $l=4e-08 $layer=LI1_cond $X=1.21 $Y=2.025
+ $X2=1.21 $Y2=1.985
r266 19 22 22.2056 $w=4.08e-07 $l=7.9e-07 $layer=LI1_cond $X=1.21 $Y=2.025
+ $X2=1.21 $Y2=2.815
r267 16 76 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.98 $Y=1.23
+ $X2=7.98 $Y2=1.395
r268 16 18 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=7.98 $Y=1.23
+ $X2=7.98 $Y2=0.91
r269 13 45 57.6553 $w=2.91e-07 $l=3.15278e-07 $layer=POLY_cond $X=6.8 $Y=2.045
+ $X2=6.875 $Y2=1.765
r270 13 15 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=6.8 $Y=2.045
+ $X2=6.8 $Y2=2.54
r271 12 71 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=3.33 $Y=0.805
+ $X2=3.33 $Y2=1.125
r272 7 40 52.2586 $w=2.99e-07 $l=2.7157e-07 $layer=POLY_cond $X=3.03 $Y=2.44
+ $X2=3.075 $Y2=2.19
r273 7 9 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=3.03 $Y=2.44 $X2=3.03
+ $Y2=2.725
r274 2 53 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=1.02
+ $Y=1.84 $X2=1.17 $Y2=1.985
r275 2 22 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=1.02
+ $Y=1.84 $X2=1.17 $Y2=2.815
r276 1 25 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1 $Y=0.37
+ $X2=1.14 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__DFBBN_1%A_595_119# 1 2 7 10 11 13 16 18 19 23 26 28
+ 30 35 39
c108 39 0 6.77906e-20 $X=3.975 $Y=1.47
c109 35 0 7.83046e-20 $X=3.72 $Y=1.595
c110 30 0 7.98666e-20 $X=3.115 $Y=0.775
c111 19 0 1.49698e-19 $X=3.41 $Y=2.65
c112 10 0 1.21772e-19 $X=4.59 $Y=1.955
r113 38 39 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=3.975 $Y=1.56
+ $X2=3.975 $Y2=1.47
r114 37 38 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.975
+ $Y=1.56 $X2=3.975 $Y2=1.56
r115 35 37 9.48476 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=3.72 $Y=1.595
+ $X2=3.975 $Y2=1.595
r116 30 32 3.31764 $w=3.28e-07 $l=9.5e-08 $layer=LI1_cond $X=3.115 $Y=0.775
+ $X2=3.115 $Y2=0.87
r117 28 35 4.5877 $w=1.7e-07 $l=2e-07 $layer=LI1_cond $X=3.72 $Y=1.395 $X2=3.72
+ $Y2=1.595
r118 27 28 28.7059 $w=1.68e-07 $l=4.4e-07 $layer=LI1_cond $X=3.72 $Y=0.955
+ $X2=3.72 $Y2=1.395
r119 25 35 8.3689 $w=3.28e-07 $l=3.09233e-07 $layer=LI1_cond $X=3.495 $Y=1.795
+ $X2=3.72 $Y2=1.595
r120 25 26 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=3.495 $Y=1.795
+ $X2=3.495 $Y2=2.565
r121 24 32 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.28 $Y=0.87
+ $X2=3.115 $Y2=0.87
r122 23 27 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.635 $Y=0.87
+ $X2=3.72 $Y2=0.955
r123 23 24 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=3.635 $Y=0.87
+ $X2=3.28 $Y2=0.87
r124 19 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.41 $Y=2.65
+ $X2=3.495 $Y2=2.565
r125 19 21 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=3.41 $Y=2.65
+ $X2=3.285 $Y2=2.65
r126 14 18 18.8402 $w=1.65e-07 $l=1.00623e-07 $layer=POLY_cond $X=4.695 $Y=1.395
+ $X2=4.635 $Y2=1.47
r127 14 16 269.202 $w=1.5e-07 $l=5.25e-07 $layer=POLY_cond $X=4.695 $Y=1.395
+ $X2=4.695 $Y2=0.87
r128 11 13 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=4.59 $Y=2.045
+ $X2=4.59 $Y2=2.54
r129 10 11 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=4.59 $Y=1.955
+ $X2=4.59 $Y2=2.045
r130 9 18 18.8402 $w=1.65e-07 $l=9.48683e-08 $layer=POLY_cond $X=4.59 $Y=1.545
+ $X2=4.635 $Y2=1.47
r131 9 10 159.371 $w=1.8e-07 $l=4.1e-07 $layer=POLY_cond $X=4.59 $Y=1.545
+ $X2=4.59 $Y2=1.955
r132 8 39 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.14 $Y=1.47
+ $X2=3.975 $Y2=1.47
r133 7 18 6.66866 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=4.5 $Y=1.47
+ $X2=4.635 $Y2=1.47
r134 7 8 184.596 $w=1.5e-07 $l=3.6e-07 $layer=POLY_cond $X=4.5 $Y=1.47 $X2=4.14
+ $Y2=1.47
r135 2 21 600 $w=1.7e-07 $l=2.38118e-07 $layer=licon1_PDIFF $count=1 $X=3.105
+ $Y=2.515 $X2=3.285 $Y2=2.65
r136 1 30 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=2.975
+ $Y=0.595 $X2=3.115 $Y2=0.775
.ends

.subckt PM_SKY130_FD_SC_HS__DFBBN_1%A_978_357# 1 2 7 9 12 16 18 19 21 22 25 26
+ 27 29 30 31 34 35 37 40 43 45 47 49 55 56 59
c179 55 0 1.32454e-19 $X=9.465 $Y=1.02
c180 49 0 1.21772e-19 $X=5.125 $Y=1.42
c181 47 0 1.48898e-19 $X=10.685 $Y=2.035
c182 35 0 5.09967e-20 $X=9.465 $Y=1.395
c183 34 0 3.62021e-19 $X=9.465 $Y=1.395
c184 31 0 1.47104e-19 $X=8.545 $Y=1.02
c185 22 0 7.44062e-20 $X=6.315 $Y=1.42
r186 52 53 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.145
+ $Y=1.5 $X2=5.145 $Y2=1.5
r187 49 52 3.29269 $w=2.78e-07 $l=8e-08 $layer=LI1_cond $X=5.125 $Y=1.42
+ $X2=5.125 $Y2=1.5
r188 45 47 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=10.515 $Y=2.035
+ $X2=10.685 $Y2=2.035
r189 41 56 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.515 $Y=1.02
+ $X2=10.43 $Y2=1.02
r190 41 43 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=10.515 $Y=1.02
+ $X2=10.725 $Y2=1.02
r191 40 45 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=10.43 $Y=1.95
+ $X2=10.515 $Y2=2.035
r192 39 56 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.43 $Y=1.105
+ $X2=10.43 $Y2=1.02
r193 39 40 55.1283 $w=1.68e-07 $l=8.45e-07 $layer=LI1_cond $X=10.43 $Y=1.105
+ $X2=10.43 $Y2=1.95
r194 38 55 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.63 $Y=1.02
+ $X2=9.465 $Y2=1.02
r195 37 56 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.345 $Y=1.02
+ $X2=10.43 $Y2=1.02
r196 37 38 46.6471 $w=1.68e-07 $l=7.15e-07 $layer=LI1_cond $X=10.345 $Y=1.02
+ $X2=9.63 $Y2=1.02
r197 35 60 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=9.465 $Y=1.395
+ $X2=9.465 $Y2=1.56
r198 35 59 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=9.465 $Y=1.395
+ $X2=9.465 $Y2=1.23
r199 34 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.465
+ $Y=1.395 $X2=9.465 $Y2=1.395
r200 32 55 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.465 $Y=1.105
+ $X2=9.465 $Y2=1.02
r201 32 34 10.1275 $w=3.28e-07 $l=2.9e-07 $layer=LI1_cond $X=9.465 $Y=1.105
+ $X2=9.465 $Y2=1.395
r202 30 55 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.3 $Y=1.02
+ $X2=9.465 $Y2=1.02
r203 30 31 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=9.3 $Y=1.02
+ $X2=8.545 $Y2=1.02
r204 29 31 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.46 $Y=0.935
+ $X2=8.545 $Y2=1.02
r205 28 29 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=8.46 $Y=0.51
+ $X2=8.46 $Y2=0.935
r206 26 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.375 $Y=0.425
+ $X2=8.46 $Y2=0.51
r207 26 27 123.305 $w=1.68e-07 $l=1.89e-06 $layer=LI1_cond $X=8.375 $Y=0.425
+ $X2=6.485 $Y2=0.425
r208 24 27 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.4 $Y=0.51
+ $X2=6.485 $Y2=0.425
r209 24 25 53.8235 $w=1.68e-07 $l=8.25e-07 $layer=LI1_cond $X=6.4 $Y=0.51
+ $X2=6.4 $Y2=1.335
r210 23 49 3.65648 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=5.265 $Y=1.42
+ $X2=5.125 $Y2=1.42
r211 22 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.315 $Y=1.42
+ $X2=6.4 $Y2=1.335
r212 22 23 68.5027 $w=1.68e-07 $l=1.05e-06 $layer=LI1_cond $X=6.315 $Y=1.42
+ $X2=5.265 $Y2=1.42
r213 19 21 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=9.51 $Y=1.885
+ $X2=9.51 $Y2=2.46
r214 18 19 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=9.51 $Y=1.795
+ $X2=9.51 $Y2=1.885
r215 18 60 91.3468 $w=1.8e-07 $l=2.35e-07 $layer=POLY_cond $X=9.51 $Y=1.795
+ $X2=9.51 $Y2=1.56
r216 16 59 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=9.445 $Y=0.75
+ $X2=9.445 $Y2=1.23
r217 10 53 39.2307 $w=2.57e-07 $l=2.07123e-07 $layer=POLY_cond $X=5.195 $Y=1.335
+ $X2=5.1 $Y2=1.5
r218 10 12 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=5.195 $Y=1.335
+ $X2=5.195 $Y2=0.87
r219 7 53 110.499 $w=2.57e-07 $l=6.02017e-07 $layer=POLY_cond $X=4.98 $Y=2.045
+ $X2=5.1 $Y2=1.5
r220 7 9 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=4.98 $Y=2.045
+ $X2=4.98 $Y2=2.54
r221 2 47 600 $w=1.7e-07 $l=2.51744e-07 $layer=licon1_PDIFF $count=1 $X=10.555
+ $Y=1.84 $X2=10.685 $Y2=2.035
r222 1 43 182 $w=1.7e-07 $l=3.33729e-07 $layer=licon1_NDIFF $count=1 $X=10.595
+ $Y=0.745 $X2=10.725 $Y2=1.02
.ends

.subckt PM_SKY130_FD_SC_HS__DFBBN_1%SET_B 1 3 6 8 9 10 12 15 17 18 23 27 30
c130 18 0 1.56839e-19 $X=5.665 $Y=2.035
c131 17 0 1.03371e-20 $X=8.735 $Y=2.035
c132 15 0 5.31324e-20 $X=9.015 $Y=0.75
c133 10 0 5.15029e-20 $X=8.89 $Y=1.885
r134 30 34 21.652 $w=3.28e-07 $l=6.2e-07 $layer=LI1_cond $X=8.895 $Y=1.415
+ $X2=8.895 $Y2=2.035
r135 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.895
+ $Y=1.415 $X2=8.895 $Y2=1.415
r136 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.685
+ $Y=1.795 $X2=5.685 $Y2=1.795
r137 23 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=2.035
+ $X2=8.88 $Y2=2.035
r138 21 27 8.8997 $w=3.29e-07 $l=2.94754e-07 $layer=LI1_cond $X=5.52 $Y=2.035
+ $X2=5.642 $Y2=1.795
r139 20 21 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=2.035
+ $X2=5.52 $Y2=2.035
r140 18 20 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.665 $Y=2.035
+ $X2=5.52 $Y2=2.035
r141 17 23 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=8.735 $Y=2.035
+ $X2=8.88 $Y2=2.035
r142 17 18 3.7995 $w=1.4e-07 $l=3.07e-06 $layer=MET1_cond $X=8.735 $Y=2.035
+ $X2=5.665 $Y2=2.035
r143 13 29 38.7084 $w=3.43e-07 $l=2.11069e-07 $layer=POLY_cond $X=9.015 $Y=1.25
+ $X2=8.91 $Y2=1.415
r144 13 15 256.383 $w=1.5e-07 $l=5e-07 $layer=POLY_cond $X=9.015 $Y=1.25
+ $X2=9.015 $Y2=0.75
r145 10 12 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=8.89 $Y=1.885
+ $X2=8.89 $Y2=2.46
r146 9 10 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=8.89 $Y=1.795 $X2=8.89
+ $Y2=1.885
r147 8 29 34.0194 $w=3.43e-07 $l=1.74714e-07 $layer=POLY_cond $X=8.89 $Y=1.58
+ $X2=8.91 $Y2=1.415
r148 8 9 83.5726 $w=1.8e-07 $l=2.15e-07 $layer=POLY_cond $X=8.89 $Y=1.58
+ $X2=8.89 $Y2=1.795
r149 4 26 39.3407 $w=3.87e-07 $l=2.09105e-07 $layer=POLY_cond $X=5.695 $Y=1.63
+ $X2=5.595 $Y2=1.795
r150 4 6 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=5.695 $Y=1.63
+ $X2=5.695 $Y2=0.87
r151 1 26 49.9272 $w=3.87e-07 $l=3.22102e-07 $layer=POLY_cond $X=5.43 $Y=2.045
+ $X2=5.595 $Y2=1.795
r152 1 3 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=5.43 $Y=2.045
+ $X2=5.43 $Y2=2.54
.ends

.subckt PM_SKY130_FD_SC_HS__DFBBN_1%A_27_74# 1 2 10 11 13 14 15 19 20 22 23 26
+ 27 28 30 34 35 36 39 40 41 43 44 45 46 47 49 53 55 56 57 60 62 68
c185 41 0 3.08859e-20 $X=7.34 $Y=2.465
c186 40 0 1.51042e-19 $X=7.34 $Y=2.375
c187 36 0 7.44062e-20 $X=6.745 $Y=1.27
c188 35 0 1.71071e-19 $X=7.25 $Y=1.27
c189 19 0 6.36774e-20 $X=2.9 $Y=0.805
r190 68 69 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.96
+ $Y=1.465 $X2=0.96 $Y2=1.465
r191 65 68 7.33373 $w=3.28e-07 $l=2.1e-07 $layer=LI1_cond $X=0.75 $Y=1.465
+ $X2=0.96 $Y2=1.465
r192 61 65 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.75 $Y=1.63
+ $X2=0.75 $Y2=1.465
r193 61 62 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=0.75 $Y=1.63
+ $X2=0.75 $Y2=1.95
r194 60 65 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.75 $Y=1.3
+ $X2=0.75 $Y2=1.465
r195 59 60 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=0.75 $Y=1.13
+ $X2=0.75 $Y2=1.3
r196 58 64 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.435 $Y=2.035
+ $X2=0.27 $Y2=2.035
r197 57 62 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.665 $Y=2.035
+ $X2=0.75 $Y2=1.95
r198 57 58 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=0.665 $Y=2.035
+ $X2=0.435 $Y2=2.035
r199 55 59 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.665 $Y=1.045
+ $X2=0.75 $Y2=1.13
r200 55 56 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=0.665 $Y=1.045
+ $X2=0.365 $Y2=1.045
r201 51 56 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.24 $Y=0.96
+ $X2=0.365 $Y2=1.045
r202 51 53 20.5135 $w=2.48e-07 $l=4.45e-07 $layer=LI1_cond $X=0.24 $Y=0.96
+ $X2=0.24 $Y2=0.515
r203 47 64 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.27 $Y=2.12 $X2=0.27
+ $Y2=2.035
r204 47 49 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=0.27 $Y=2.12
+ $X2=0.27 $Y2=2.815
r205 41 43 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=7.34 $Y=2.465
+ $X2=7.34 $Y2=2.75
r206 40 41 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=7.34 $Y=2.375
+ $X2=7.34 $Y2=2.465
r207 39 46 37.1337 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=7.34 $Y=1.89 $X2=7.34
+ $Y2=1.8
r208 39 40 188.524 $w=1.8e-07 $l=4.85e-07 $layer=POLY_cond $X=7.34 $Y=1.89
+ $X2=7.34 $Y2=2.375
r209 37 46 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=7.325 $Y=1.345
+ $X2=7.325 $Y2=1.8
r210 35 37 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=7.25 $Y=1.27
+ $X2=7.325 $Y2=1.345
r211 35 36 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=7.25 $Y=1.27
+ $X2=6.745 $Y2=1.27
r212 32 36 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=6.67 $Y=1.195
+ $X2=6.745 $Y2=1.27
r213 32 34 179.468 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=6.67 $Y=1.195
+ $X2=6.67 $Y2=0.845
r214 31 34 302.532 $w=1.5e-07 $l=5.9e-07 $layer=POLY_cond $X=6.67 $Y=0.255
+ $X2=6.67 $Y2=0.845
r215 28 30 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=3.54 $Y=2.44
+ $X2=3.54 $Y2=2.725
r216 27 28 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=3.54 $Y=2.35 $X2=3.54
+ $Y2=2.44
r217 26 45 37.1337 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=3.54 $Y=2.055
+ $X2=3.54 $Y2=1.965
r218 26 27 114.669 $w=1.8e-07 $l=2.95e-07 $layer=POLY_cond $X=3.54 $Y=2.055
+ $X2=3.54 $Y2=2.35
r219 24 45 76.9149 $w=1.5e-07 $l=1.5e-07 $layer=POLY_cond $X=3.525 $Y=1.815
+ $X2=3.525 $Y2=1.965
r220 22 24 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.45 $Y=1.74
+ $X2=3.525 $Y2=1.815
r221 22 23 243.564 $w=1.5e-07 $l=4.75e-07 $layer=POLY_cond $X=3.45 $Y=1.74
+ $X2=2.975 $Y2=1.74
r222 21 44 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.975 $Y=0.18
+ $X2=2.9 $Y2=0.18
r223 20 31 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=6.595 $Y=0.18
+ $X2=6.67 $Y2=0.255
r224 20 21 1856.21 $w=1.5e-07 $l=3.62e-06 $layer=POLY_cond $X=6.595 $Y=0.18
+ $X2=2.975 $Y2=0.18
r225 17 23 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.9 $Y=1.665
+ $X2=2.975 $Y2=1.74
r226 17 19 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=2.9 $Y=1.665
+ $X2=2.9 $Y2=0.805
r227 16 44 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.9 $Y=0.255
+ $X2=2.9 $Y2=0.18
r228 16 19 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=2.9 $Y=0.255
+ $X2=2.9 $Y2=0.805
r229 14 44 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.825 $Y=0.18
+ $X2=2.9 $Y2=0.18
r230 14 15 935.798 $w=1.5e-07 $l=1.825e-06 $layer=POLY_cond $X=2.825 $Y=0.18
+ $X2=1 $Y2=0.18
r231 11 69 61.4066 $w=2.86e-07 $l=3.07409e-07 $layer=POLY_cond $X=0.945 $Y=1.765
+ $X2=0.96 $Y2=1.465
r232 11 13 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.945 $Y=1.765
+ $X2=0.945 $Y2=2.4
r233 8 69 38.6549 $w=2.86e-07 $l=1.81659e-07 $layer=POLY_cond $X=0.925 $Y=1.3
+ $X2=0.96 $Y2=1.465
r234 8 10 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=0.925 $Y=1.3
+ $X2=0.925 $Y2=0.74
r235 7 15 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.925 $Y=0.255
+ $X2=1 $Y2=0.18
r236 7 10 248.691 $w=1.5e-07 $l=4.85e-07 $layer=POLY_cond $X=0.925 $Y=0.255
+ $X2=0.925 $Y2=0.74
r237 2 64 400 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.27 $Y2=2.115
r238 2 49 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.27 $Y2=2.815
r239 1 53 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__DFBBN_1%A_1534_446# 1 2 3 10 12 15 17 19 22 24 25 27
+ 29 30 32 33 35 38 40 43 47 48 51 52 54 58 59 60 65 68 69 73 75
c211 65 0 5.76555e-20 $X=11.3 $Y=2.29
c212 54 0 5.31324e-20 $X=11.215 $Y=0.68
c213 47 0 1.02788e-19 $X=8.055 $Y=2.215
c214 25 0 6.25621e-20 $X=11.585 $Y=1.477
c215 17 0 2.31979e-19 $X=11.435 $Y=1.765
c216 1 0 1.81011e-19 $X=9.52 $Y=0.38
r217 81 82 8.60714 $w=3.92e-07 $l=7e-08 $layer=POLY_cond $X=11.435 $Y=1.542
+ $X2=11.505 $Y2=1.542
r218 74 81 1.84439 $w=3.92e-07 $l=1.5e-08 $layer=POLY_cond $X=11.42 $Y=1.542
+ $X2=11.435 $Y2=1.542
r219 73 76 8.53881 $w=3.68e-07 $l=1.65e-07 $layer=LI1_cond $X=11.4 $Y=1.485
+ $X2=11.4 $Y2=1.65
r220 73 75 8.53881 $w=3.68e-07 $l=1.65e-07 $layer=LI1_cond $X=11.4 $Y=1.485
+ $X2=11.4 $Y2=1.32
r221 73 74 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=11.42
+ $Y=1.485 $X2=11.42 $Y2=1.485
r222 67 69 8.48848 $w=3.48e-07 $l=1.65e-07 $layer=LI1_cond $X=8.665 $Y=2.805
+ $X2=8.83 $Y2=2.805
r223 67 68 8.48848 $w=3.48e-07 $l=1.65e-07 $layer=LI1_cond $X=8.665 $Y=2.805
+ $X2=8.5 $Y2=2.805
r224 65 76 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=11.3 $Y=2.29
+ $X2=11.3 $Y2=1.65
r225 62 75 36.2086 $w=1.68e-07 $l=5.55e-07 $layer=LI1_cond $X=11.3 $Y=0.765
+ $X2=11.3 $Y2=1.32
r226 61 71 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.32 $Y=2.375
+ $X2=10.155 $Y2=2.375
r227 60 65 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=11.215 $Y=2.375
+ $X2=11.3 $Y2=2.29
r228 60 61 58.3904 $w=1.68e-07 $l=8.95e-07 $layer=LI1_cond $X=11.215 $Y=2.375
+ $X2=10.32 $Y2=2.375
r229 58 71 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=10.155 $Y=2.46
+ $X2=10.155 $Y2=2.375
r230 58 59 5.93683 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=10.155 $Y=2.46
+ $X2=10.155 $Y2=2.63
r231 54 62 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=11.215 $Y=0.68
+ $X2=11.3 $Y2=0.765
r232 54 56 100.144 $w=1.68e-07 $l=1.535e-06 $layer=LI1_cond $X=11.215 $Y=0.68
+ $X2=9.68 $Y2=0.68
r233 52 59 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=9.99 $Y=2.715
+ $X2=10.155 $Y2=2.63
r234 52 69 75.6791 $w=1.68e-07 $l=1.16e-06 $layer=LI1_cond $X=9.99 $Y=2.715
+ $X2=8.83 $Y2=2.715
r235 51 68 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=8.22 $Y=2.715
+ $X2=8.5 $Y2=2.715
r236 48 79 50.9497 $w=2.98e-07 $l=3.15e-07 $layer=POLY_cond $X=8.055 $Y=2.257
+ $X2=8.37 $Y2=2.257
r237 48 77 47.7148 $w=2.98e-07 $l=2.95e-07 $layer=POLY_cond $X=8.055 $Y=2.257
+ $X2=7.76 $Y2=2.257
r238 47 48 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.055
+ $Y=2.215 $X2=8.055 $Y2=2.215
r239 45 51 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=8.055 $Y=2.63
+ $X2=8.22 $Y2=2.715
r240 45 47 14.4928 $w=3.28e-07 $l=4.15e-07 $layer=LI1_cond $X=8.055 $Y=2.63
+ $X2=8.055 $Y2=2.215
r241 41 43 117.936 $w=1.5e-07 $l=2.3e-07 $layer=POLY_cond $X=12.19 $Y=1.9
+ $X2=12.42 $Y2=1.9
r242 36 38 141.011 $w=1.5e-07 $l=2.75e-07 $layer=POLY_cond $X=12.19 $Y=0.94
+ $X2=12.465 $Y2=0.94
r243 33 38 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=12.465 $Y=0.865
+ $X2=12.465 $Y2=0.94
r244 33 35 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=12.465 $Y=0.865
+ $X2=12.465 $Y2=0.58
r245 30 43 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=12.42 $Y=1.975
+ $X2=12.42 $Y2=1.9
r246 30 32 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=12.42 $Y=1.975
+ $X2=12.42 $Y2=2.47
r247 29 41 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=12.19 $Y=1.825
+ $X2=12.19 $Y2=1.9
r248 28 40 35.9208 $w=1.5e-07 $l=1.58e-07 $layer=POLY_cond $X=12.19 $Y=1.635
+ $X2=12.19 $Y2=1.477
r249 28 29 97.4255 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=12.19 $Y=1.635
+ $X2=12.19 $Y2=1.825
r250 27 40 35.9208 $w=1.5e-07 $l=1.57e-07 $layer=POLY_cond $X=12.19 $Y=1.32
+ $X2=12.19 $Y2=1.477
r251 26 36 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=12.19 $Y=1.015
+ $X2=12.19 $Y2=0.94
r252 26 27 156.394 $w=1.5e-07 $l=3.05e-07 $layer=POLY_cond $X=12.19 $Y=1.015
+ $X2=12.19 $Y2=1.32
r253 25 82 11.8363 $w=3.92e-07 $l=1.07703e-07 $layer=POLY_cond $X=11.585
+ $Y=1.477 $X2=11.505 $Y2=1.542
r254 24 40 4.4846 $w=3.15e-07 $l=7.5e-08 $layer=POLY_cond $X=12.115 $Y=1.477
+ $X2=12.19 $Y2=1.477
r255 24 25 97.0896 $w=3.15e-07 $l=5.3e-07 $layer=POLY_cond $X=12.115 $Y=1.477
+ $X2=11.585 $Y2=1.477
r256 20 82 25.3688 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=11.505 $Y=1.32
+ $X2=11.505 $Y2=1.542
r257 20 22 269.202 $w=1.5e-07 $l=5.25e-07 $layer=POLY_cond $X=11.505 $Y=1.32
+ $X2=11.505 $Y2=0.795
r258 17 81 25.3688 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=11.435 $Y=1.765
+ $X2=11.435 $Y2=1.542
r259 17 19 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=11.435 $Y=1.765
+ $X2=11.435 $Y2=2.4
r260 13 79 18.8112 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=8.37 $Y=2.05
+ $X2=8.37 $Y2=2.257
r261 13 15 584.553 $w=1.5e-07 $l=1.14e-06 $layer=POLY_cond $X=8.37 $Y=2.05
+ $X2=8.37 $Y2=0.91
r262 10 77 18.8112 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=7.76 $Y=2.465
+ $X2=7.76 $Y2=2.257
r263 10 12 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=7.76 $Y=2.465
+ $X2=7.76 $Y2=2.75
r264 3 71 300 $w=1.7e-07 $l=5.65044e-07 $layer=licon1_PDIFF $count=2 $X=10.005
+ $Y=1.96 $X2=10.155 $Y2=2.455
r265 2 67 600 $w=1.7e-07 $l=9.14631e-07 $layer=licon1_PDIFF $count=1 $X=8.52
+ $Y=1.96 $X2=8.665 $Y2=2.805
r266 1 56 182 $w=1.7e-07 $l=3.71484e-07 $layer=licon1_NDIFF $count=1 $X=9.52
+ $Y=0.38 $X2=9.68 $Y2=0.68
.ends

.subckt PM_SKY130_FD_SC_HS__DFBBN_1%A_1349_114# 1 2 9 11 13 14 22 26 27 29 30 33
+ 34 35 37 38 39 42 46 47 48
c150 46 0 3.08859e-20 $X=7.025 $Y=2.265
c151 30 0 5.15029e-20 $X=8.39 $Y=1.815
c152 29 0 1.39048e-19 $X=8.12 $Y=1.73
c153 27 0 1.72728e-19 $X=7.415 $Y=1.815
c154 14 0 1.06589e-20 $X=8.035 $Y=0.845
r155 46 47 9.86413 $w=5.53e-07 $l=1.65e-07 $layer=LI1_cond $X=7.137 $Y=2.265
+ $X2=7.137 $Y2=2.1
r156 42 43 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.005
+ $Y=1.585 $X2=10.005 $Y2=1.585
r157 40 42 12.7467 $w=3.28e-07 $l=3.65e-07 $layer=LI1_cond $X=10.005 $Y=1.95
+ $X2=10.005 $Y2=1.585
r158 38 40 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=9.84 $Y=2.035
+ $X2=10.005 $Y2=1.95
r159 38 39 28.7059 $w=1.68e-07 $l=4.4e-07 $layer=LI1_cond $X=9.84 $Y=2.035
+ $X2=9.4 $Y2=2.035
r160 36 39 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.315 $Y=2.12
+ $X2=9.4 $Y2=2.035
r161 36 37 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=9.315 $Y=2.12
+ $X2=9.315 $Y2=2.29
r162 34 37 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.23 $Y=2.375
+ $X2=9.315 $Y2=2.29
r163 34 35 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=9.23 $Y=2.375
+ $X2=8.56 $Y2=2.375
r164 33 35 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.475 $Y=2.29
+ $X2=8.56 $Y2=2.375
r165 32 33 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=8.475 $Y=1.9
+ $X2=8.475 $Y2=2.29
r166 31 48 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.205 $Y=1.815
+ $X2=8.12 $Y2=1.815
r167 30 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.39 $Y=1.815
+ $X2=8.475 $Y2=1.9
r168 30 31 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=8.39 $Y=1.815
+ $X2=8.205 $Y2=1.815
r169 29 48 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.12 $Y=1.73
+ $X2=8.12 $Y2=1.815
r170 28 29 46.9733 $w=1.68e-07 $l=7.2e-07 $layer=LI1_cond $X=8.12 $Y=1.01
+ $X2=8.12 $Y2=1.73
r171 26 48 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.035 $Y=1.815
+ $X2=8.12 $Y2=1.815
r172 26 27 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=8.035 $Y=1.815
+ $X2=7.415 $Y2=1.815
r173 24 27 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.33 $Y=1.9
+ $X2=7.415 $Y2=1.815
r174 24 47 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=7.33 $Y=1.9 $X2=7.33
+ $Y2=2.1
r175 20 46 2.41371 $w=5.53e-07 $l=1.12e-07 $layer=LI1_cond $X=7.137 $Y=2.377
+ $X2=7.137 $Y2=2.265
r176 20 22 9.43932 $w=5.53e-07 $l=4.38e-07 $layer=LI1_cond $X=7.137 $Y=2.377
+ $X2=7.137 $Y2=2.815
r177 16 19 27.938 $w=3.28e-07 $l=8e-07 $layer=LI1_cond $X=6.885 $Y=0.845
+ $X2=7.685 $Y2=0.845
r178 14 28 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=8.035 $Y=0.845
+ $X2=8.12 $Y2=1.01
r179 14 19 12.2229 $w=3.28e-07 $l=3.5e-07 $layer=LI1_cond $X=8.035 $Y=0.845
+ $X2=7.685 $Y2=0.845
r180 11 43 61.4066 $w=2.86e-07 $l=3.3541e-07 $layer=POLY_cond $X=9.93 $Y=1.885
+ $X2=10.005 $Y2=1.585
r181 11 13 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=9.93 $Y=1.885
+ $X2=9.93 $Y2=2.46
r182 7 43 38.6549 $w=2.86e-07 $l=2.05122e-07 $layer=POLY_cond $X=9.915 $Y=1.42
+ $X2=10.005 $Y2=1.585
r183 7 9 343.553 $w=1.5e-07 $l=6.7e-07 $layer=POLY_cond $X=9.915 $Y=1.42
+ $X2=9.915 $Y2=0.75
r184 2 46 600 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=6.875
+ $Y=2.12 $X2=7.025 $Y2=2.265
r185 2 22 600 $w=1.7e-07 $l=7.66339e-07 $layer=licon1_PDIFF $count=1 $X=6.875
+ $Y=2.12 $X2=7.025 $Y2=2.815
r186 1 19 121.333 $w=1.7e-07 $l=1.06869e-06 $layer=licon1_NDIFF $count=1
+ $X=6.745 $Y=0.57 $X2=7.685 $Y2=0.845
r187 1 16 121.333 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1
+ $X=6.745 $Y=0.57 $X2=6.885 $Y2=0.845
.ends

.subckt PM_SKY130_FD_SC_HS__DFBBN_1%RESET_B 1 3 6 8 12
c32 12 0 4.16644e-20 $X=10.85 $Y=1.515
c33 6 0 1.78363e-19 $X=10.94 $Y=0.955
r34 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.85
+ $Y=1.515 $X2=10.85 $Y2=1.515
r35 8 12 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=10.85 $Y=1.665
+ $X2=10.85 $Y2=1.515
r36 4 11 38.5562 $w=2.99e-07 $l=2.05122e-07 $layer=POLY_cond $X=10.94 $Y=1.35
+ $X2=10.85 $Y2=1.515
r37 4 6 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=10.94 $Y=1.35
+ $X2=10.94 $Y2=0.955
r38 1 11 52.2586 $w=2.99e-07 $l=2.78388e-07 $layer=POLY_cond $X=10.91 $Y=1.765
+ $X2=10.85 $Y2=1.515
r39 1 3 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=10.91 $Y=1.765
+ $X2=10.91 $Y2=2.16
.ends

.subckt PM_SKY130_FD_SC_HS__DFBBN_1%A_2412_410# 1 2 7 9 12 15 19 23 27 30
c57 15 0 1.18517e-19 $X=12.855 $Y=1.42
r58 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=12.67
+ $Y=1.42 $X2=12.67 $Y2=1.42
r59 25 30 0.364692 $w=3.3e-07 $l=1.25e-07 $layer=LI1_cond $X=12.36 $Y=1.42
+ $X2=12.235 $Y2=1.42
r60 25 27 10.826 $w=3.28e-07 $l=3.1e-07 $layer=LI1_cond $X=12.36 $Y=1.42
+ $X2=12.67 $Y2=1.42
r61 21 30 6.46576 $w=2.5e-07 $l=1.65e-07 $layer=LI1_cond $X=12.235 $Y=1.585
+ $X2=12.235 $Y2=1.42
r62 21 23 28.1196 $w=2.48e-07 $l=6.1e-07 $layer=LI1_cond $X=12.235 $Y=1.585
+ $X2=12.235 $Y2=2.195
r63 17 30 6.46576 $w=2.5e-07 $l=1.65e-07 $layer=LI1_cond $X=12.235 $Y=1.255
+ $X2=12.235 $Y2=1.42
r64 17 19 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=12.235 $Y=1.255
+ $X2=12.235 $Y2=0.58
r65 15 28 32.3493 $w=3.3e-07 $l=1.85e-07 $layer=POLY_cond $X=12.855 $Y=1.42
+ $X2=12.67 $Y2=1.42
r66 15 16 66.2869 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=12.945 $Y=1.42
+ $X2=12.945 $Y2=1.255
r67 12 16 264.074 $w=1.5e-07 $l=5.15e-07 $layer=POLY_cond $X=12.96 $Y=0.74
+ $X2=12.96 $Y2=1.255
r68 7 15 136.255 $w=1.8e-07 $l=3.45e-07 $layer=POLY_cond $X=12.945 $Y=1.765
+ $X2=12.945 $Y2=1.42
r69 7 9 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=12.945 $Y=1.765
+ $X2=12.945 $Y2=2.4
r70 2 23 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=12.06
+ $Y=2.05 $X2=12.195 $Y2=2.195
r71 1 19 182 $w=1.7e-07 $l=2.67208e-07 $layer=licon1_NDIFF $count=1 $X=12.12
+ $Y=0.37 $X2=12.25 $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_HS__DFBBN_1%VPWR 1 2 3 4 5 6 7 8 27 31 35 39 43 47 52 53
+ 55 56 57 59 71 79 83 88 93 100 101 104 107 110 117 124 127
r160 127 128 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.72 $Y=3.33
+ $X2=12.72 $Y2=3.33
r161 124 125 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.28 $Y=3.33
+ $X2=11.28 $Y2=3.33
r162 120 121 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.36 $Y=3.33
+ $X2=9.36 $Y2=3.33
r163 117 120 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=9.2 $Y=3.055
+ $X2=9.2 $Y2=3.33
r164 107 108 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r165 104 105 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r166 101 128 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=13.2 $Y=3.33
+ $X2=12.72 $Y2=3.33
r167 100 101 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.2 $Y=3.33
+ $X2=13.2 $Y2=3.33
r168 98 127 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=12.805 $Y=3.33
+ $X2=12.68 $Y2=3.33
r169 98 100 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=12.805 $Y=3.33
+ $X2=13.2 $Y2=3.33
r170 97 128 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.24 $Y=3.33
+ $X2=12.72 $Y2=3.33
r171 97 125 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=12.24 $Y=3.33
+ $X2=11.28 $Y2=3.33
r172 96 97 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=12.24 $Y=3.33
+ $X2=12.24 $Y2=3.33
r173 94 124 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.375 $Y=3.33
+ $X2=11.21 $Y2=3.33
r174 94 96 56.4332 $w=1.68e-07 $l=8.65e-07 $layer=LI1_cond $X=11.375 $Y=3.33
+ $X2=12.24 $Y2=3.33
r175 93 127 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=12.555 $Y=3.33
+ $X2=12.68 $Y2=3.33
r176 93 96 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=12.555 $Y=3.33
+ $X2=12.24 $Y2=3.33
r177 92 125 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.8 $Y=3.33
+ $X2=11.28 $Y2=3.33
r178 92 121 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=10.8 $Y=3.33
+ $X2=9.36 $Y2=3.33
r179 91 92 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.8 $Y=3.33
+ $X2=10.8 $Y2=3.33
r180 89 120 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.365 $Y=3.33
+ $X2=9.2 $Y2=3.33
r181 89 91 93.6203 $w=1.68e-07 $l=1.435e-06 $layer=LI1_cond $X=9.365 $Y=3.33
+ $X2=10.8 $Y2=3.33
r182 88 124 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.045 $Y=3.33
+ $X2=11.21 $Y2=3.33
r183 88 91 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=11.045 $Y=3.33
+ $X2=10.8 $Y2=3.33
r184 87 121 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=3.33
+ $X2=9.36 $Y2=3.33
r185 87 114 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=8.88 $Y=3.33
+ $X2=7.92 $Y2=3.33
r186 86 87 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r187 84 86 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=8.27 $Y=3.33
+ $X2=8.88 $Y2=3.33
r188 83 120 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.035 $Y=3.33
+ $X2=9.2 $Y2=3.33
r189 83 86 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=9.035 $Y=3.33
+ $X2=8.88 $Y2=3.33
r190 81 82 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r191 79 84 5.2253 $w=1.7e-07 $l=1.83e-07 $layer=LI1_cond $X=8.087 $Y=3.33
+ $X2=8.27 $Y2=3.33
r192 79 114 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r193 79 110 8.68279 $w=3.63e-07 $l=2.75e-07 $layer=LI1_cond $X=8.087 $Y=3.33
+ $X2=8.087 $Y2=3.055
r194 79 81 92.9679 $w=1.68e-07 $l=1.425e-06 $layer=LI1_cond $X=7.905 $Y=3.33
+ $X2=6.48 $Y2=3.33
r195 78 82 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=3.33 $X2=6.48
+ $Y2=3.33
r196 78 108 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6 $Y=3.33
+ $X2=5.04 $Y2=3.33
r197 77 78 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r198 75 107 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.37 $Y=3.33
+ $X2=5.205 $Y2=3.33
r199 75 77 41.1016 $w=1.68e-07 $l=6.3e-07 $layer=LI1_cond $X=5.37 $Y=3.33 $X2=6
+ $Y2=3.33
r200 74 108 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=5.04 $Y2=3.33
r201 73 74 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r202 71 107 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.04 $Y=3.33
+ $X2=5.205 $Y2=3.33
r203 71 73 156.578 $w=1.68e-07 $l=2.4e-06 $layer=LI1_cond $X=5.04 $Y=3.33
+ $X2=2.64 $Y2=3.33
r204 70 74 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r205 69 70 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r206 67 70 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.16 $Y2=3.33
r207 67 105 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r208 66 69 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.2 $Y=3.33 $X2=2.16
+ $Y2=3.33
r209 66 67 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r210 64 104 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.805 $Y=3.33
+ $X2=0.72 $Y2=3.33
r211 64 66 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=0.805 $Y=3.33
+ $X2=1.2 $Y2=3.33
r212 62 105 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r213 61 62 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r214 59 104 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.635 $Y=3.33
+ $X2=0.72 $Y2=3.33
r215 59 61 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=0.635 $Y=3.33
+ $X2=0.24 $Y2=3.33
r216 57 114 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=6.72 $Y=3.33
+ $X2=7.92 $Y2=3.33
r217 57 82 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=6.72 $Y=3.33
+ $X2=6.48 $Y2=3.33
r218 55 77 1.30481 $w=1.68e-07 $l=2e-08 $layer=LI1_cond $X=6.02 $Y=3.33 $X2=6
+ $Y2=3.33
r219 55 56 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.02 $Y=3.33
+ $X2=6.185 $Y2=3.33
r220 54 81 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=6.35 $Y=3.33
+ $X2=6.48 $Y2=3.33
r221 54 56 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.35 $Y=3.33
+ $X2=6.185 $Y2=3.33
r222 52 69 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=2.295 $Y=3.33
+ $X2=2.16 $Y2=3.33
r223 52 53 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.295 $Y=3.33
+ $X2=2.38 $Y2=3.33
r224 51 73 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=2.465 $Y=3.33
+ $X2=2.64 $Y2=3.33
r225 51 53 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.465 $Y=3.33
+ $X2=2.38 $Y2=3.33
r226 47 50 19.1306 $w=2.48e-07 $l=4.15e-07 $layer=LI1_cond $X=12.68 $Y=1.985
+ $X2=12.68 $Y2=2.4
r227 45 127 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=12.68 $Y=3.245
+ $X2=12.68 $Y2=3.33
r228 45 50 38.9526 $w=2.48e-07 $l=8.45e-07 $layer=LI1_cond $X=12.68 $Y=3.245
+ $X2=12.68 $Y2=2.4
r229 41 124 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=11.21 $Y=3.245
+ $X2=11.21 $Y2=3.33
r230 41 43 15.3659 $w=3.28e-07 $l=4.4e-07 $layer=LI1_cond $X=11.21 $Y=3.245
+ $X2=11.21 $Y2=2.805
r231 37 56 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.185 $Y=3.245
+ $X2=6.185 $Y2=3.33
r232 37 39 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=6.185 $Y=3.245
+ $X2=6.185 $Y2=2.78
r233 33 107 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.205 $Y=3.245
+ $X2=5.205 $Y2=3.33
r234 33 35 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=5.205 $Y=3.245
+ $X2=5.205 $Y2=2.78
r235 29 53 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.38 $Y=3.245
+ $X2=2.38 $Y2=3.33
r236 29 31 32.9465 $w=1.68e-07 $l=5.05e-07 $layer=LI1_cond $X=2.38 $Y=3.245
+ $X2=2.38 $Y2=2.74
r237 25 104 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.72 $Y=3.245
+ $X2=0.72 $Y2=3.33
r238 25 27 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=0.72 $Y=3.245
+ $X2=0.72 $Y2=2.455
r239 8 50 300 $w=1.7e-07 $l=4.48609e-07 $layer=licon1_PDIFF $count=2 $X=12.495
+ $Y=2.05 $X2=12.72 $Y2=2.4
r240 8 47 600 $w=1.7e-07 $l=2.55441e-07 $layer=licon1_PDIFF $count=1 $X=12.495
+ $Y=2.05 $X2=12.72 $Y2=1.985
r241 7 43 600 $w=1.7e-07 $l=1.07161e-06 $layer=licon1_PDIFF $count=1 $X=10.985
+ $Y=1.84 $X2=11.21 $Y2=2.805
r242 6 117 600 $w=1.7e-07 $l=1.20679e-06 $layer=licon1_PDIFF $count=1 $X=8.965
+ $Y=1.96 $X2=9.2 $Y2=3.055
r243 5 110 600 $w=1.7e-07 $l=6.27674e-07 $layer=licon1_PDIFF $count=1 $X=7.835
+ $Y=2.54 $X2=8.085 $Y2=3.055
r244 4 39 600 $w=1.7e-07 $l=7.2208e-07 $layer=licon1_PDIFF $count=1 $X=6.055
+ $Y=2.12 $X2=6.185 $Y2=2.78
r245 3 35 600 $w=1.7e-07 $l=7.31163e-07 $layer=licon1_PDIFF $count=1 $X=5.055
+ $Y=2.12 $X2=5.205 $Y2=2.78
r246 2 31 600 $w=1.7e-07 $l=3.91663e-07 $layer=licon1_PDIFF $count=1 $X=2.085
+ $Y=2.515 $X2=2.38 $Y2=2.74
r247 1 27 300 $w=1.7e-07 $l=6.85912e-07 $layer=licon1_PDIFF $count=2 $X=0.57
+ $Y=1.84 $X2=0.72 $Y2=2.455
.ends

.subckt PM_SKY130_FD_SC_HS__DFBBN_1%A_311_119# 1 2 3 4 15 18 20 21 22 27 30 31
+ 32 34 36 41 42 44 47
r122 45 47 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=4.06 $Y=1.08
+ $X2=4.39 $Y2=1.08
r123 41 42 9.43135 $w=1.98e-07 $l=1.65e-07 $layer=LI1_cond $X=1.685 $Y=2.57
+ $X2=1.685 $Y2=2.405
r124 39 42 91.0107 $w=1.68e-07 $l=1.395e-06 $layer=LI1_cond $X=1.67 $Y=1.01
+ $X2=1.67 $Y2=2.405
r125 38 39 5.26419 $w=2.78e-07 $l=8.5e-08 $layer=LI1_cond $X=1.725 $Y=0.925
+ $X2=1.725 $Y2=1.01
r126 36 38 5.55642 $w=2.78e-07 $l=1.35e-07 $layer=LI1_cond $X=1.725 $Y=0.79
+ $X2=1.725 $Y2=0.925
r127 33 47 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.39 $Y=1.165
+ $X2=4.39 $Y2=1.08
r128 33 34 52.1925 $w=1.68e-07 $l=8e-07 $layer=LI1_cond $X=4.39 $Y=1.165
+ $X2=4.39 $Y2=1.965
r129 31 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.305 $Y=2.05
+ $X2=4.39 $Y2=1.965
r130 31 32 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=4.305 $Y=2.05
+ $X2=4 $Y2=2.05
r131 30 45 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.06 $Y=0.995
+ $X2=4.06 $Y2=1.08
r132 29 30 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=4.06 $Y=0.615
+ $X2=4.06 $Y2=0.995
r133 25 32 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=3.875 $Y=2.135
+ $X2=4 $Y2=2.05
r134 25 27 20.0525 $w=2.48e-07 $l=4.35e-07 $layer=LI1_cond $X=3.875 $Y=2.135
+ $X2=3.875 $Y2=2.57
r135 22 44 8.99121 $w=3.58e-07 $l=1.8e-07 $layer=LI1_cond $X=3.64 $Y=0.435
+ $X2=3.46 $Y2=0.435
r136 22 24 4.1616 $w=3.58e-07 $l=1.3e-07 $layer=LI1_cond $X=3.64 $Y=0.435
+ $X2=3.77 $Y2=0.435
r137 21 29 8.02311 $w=3.6e-07 $l=2.18403e-07 $layer=LI1_cond $X=3.975 $Y=0.435
+ $X2=4.06 $Y2=0.615
r138 21 24 6.56252 $w=3.58e-07 $l=2.05e-07 $layer=LI1_cond $X=3.975 $Y=0.435
+ $X2=3.77 $Y2=0.435
r139 20 44 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=2.75 $Y=0.34
+ $X2=3.46 $Y2=0.34
r140 17 20 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.665 $Y=0.425
+ $X2=2.75 $Y2=0.34
r141 17 18 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=2.665 $Y=0.425
+ $X2=2.665 $Y2=0.84
r142 16 38 3.65648 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=1.865 $Y=0.925
+ $X2=1.725 $Y2=0.925
r143 15 18 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.58 $Y=0.925
+ $X2=2.665 $Y2=0.84
r144 15 16 46.6471 $w=1.68e-07 $l=7.15e-07 $layer=LI1_cond $X=2.58 $Y=0.925
+ $X2=1.865 $Y2=0.925
r145 4 27 600 $w=1.7e-07 $l=2.45967e-07 $layer=licon1_PDIFF $count=1 $X=3.615
+ $Y=2.515 $X2=3.835 $Y2=2.57
r146 3 41 600 $w=1.7e-07 $l=1.99687e-07 $layer=licon1_PDIFF $count=1 $X=1.57
+ $Y=2.425 $X2=1.7 $Y2=2.57
r147 2 24 182 $w=1.7e-07 $l=3.96169e-07 $layer=licon1_NDIFF $count=1 $X=3.405
+ $Y=0.595 $X2=3.77 $Y2=0.53
r148 1 36 182 $w=1.7e-07 $l=2.57488e-07 $layer=licon1_NDIFF $count=1 $X=1.555
+ $Y=0.595 $X2=1.7 $Y2=0.79
.ends

.subckt PM_SKY130_FD_SC_HS__DFBBN_1%Q_N 1 2 9 13 14 15 16 23 33
c37 33 0 1.59934e-19 $X=11.75 $Y=1.82
c38 14 0 6.25621e-20 $X=11.675 $Y=1.95
c39 9 0 1.78363e-19 $X=11.72 $Y=0.57
r40 21 35 0.329269 $w=3.48e-07 $l=1e-08 $layer=LI1_cond $X=11.75 $Y=1.995
+ $X2=11.75 $Y2=1.985
r41 21 23 1.31708 $w=3.48e-07 $l=4e-08 $layer=LI1_cond $X=11.75 $Y=1.995
+ $X2=11.75 $Y2=2.035
r42 16 30 1.31708 $w=3.48e-07 $l=4e-08 $layer=LI1_cond $X=11.75 $Y=2.775
+ $X2=11.75 $Y2=2.815
r43 15 16 12.183 $w=3.48e-07 $l=3.7e-07 $layer=LI1_cond $X=11.75 $Y=2.405
+ $X2=11.75 $Y2=2.775
r44 14 35 0.42805 $w=3.48e-07 $l=1.3e-08 $layer=LI1_cond $X=11.75 $Y=1.972
+ $X2=11.75 $Y2=1.985
r45 14 33 8.06043 $w=3.48e-07 $l=1.52e-07 $layer=LI1_cond $X=11.75 $Y=1.972
+ $X2=11.75 $Y2=1.82
r46 14 15 11.4586 $w=3.48e-07 $l=3.48e-07 $layer=LI1_cond $X=11.75 $Y=2.057
+ $X2=11.75 $Y2=2.405
r47 14 23 0.724393 $w=3.48e-07 $l=2.2e-08 $layer=LI1_cond $X=11.75 $Y=2.057
+ $X2=11.75 $Y2=2.035
r48 13 33 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=11.84 $Y=1.15
+ $X2=11.84 $Y2=1.82
r49 7 13 9.16175 $w=3.68e-07 $l=1.85e-07 $layer=LI1_cond $X=11.74 $Y=0.965
+ $X2=11.74 $Y2=1.15
r50 7 9 12.3031 $w=3.68e-07 $l=3.95e-07 $layer=LI1_cond $X=11.74 $Y=0.965
+ $X2=11.74 $Y2=0.57
r51 2 35 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=11.51
+ $Y=1.84 $X2=11.66 $Y2=1.985
r52 2 30 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=11.51
+ $Y=1.84 $X2=11.66 $Y2=2.815
r53 1 9 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=11.58
+ $Y=0.425 $X2=11.72 $Y2=0.57
.ends

.subckt PM_SKY130_FD_SC_HS__DFBBN_1%Q 1 2 7 8 9 10 11 12 13
r15 12 13 12.7285 $w=3.33e-07 $l=3.7e-07 $layer=LI1_cond $X=13.172 $Y=2.405
+ $X2=13.172 $Y2=2.775
r16 11 12 14.4485 $w=3.33e-07 $l=4.2e-07 $layer=LI1_cond $X=13.172 $Y=1.985
+ $X2=13.172 $Y2=2.405
r17 10 11 11.0084 $w=3.33e-07 $l=3.2e-07 $layer=LI1_cond $X=13.172 $Y=1.665
+ $X2=13.172 $Y2=1.985
r18 9 10 12.7285 $w=3.33e-07 $l=3.7e-07 $layer=LI1_cond $X=13.172 $Y=1.295
+ $X2=13.172 $Y2=1.665
r19 8 9 12.7285 $w=3.33e-07 $l=3.7e-07 $layer=LI1_cond $X=13.172 $Y=0.925
+ $X2=13.172 $Y2=1.295
r20 7 8 14.1045 $w=3.33e-07 $l=4.1e-07 $layer=LI1_cond $X=13.172 $Y=0.515
+ $X2=13.172 $Y2=0.925
r21 2 13 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=13.02
+ $Y=1.84 $X2=13.17 $Y2=2.815
r22 2 11 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=13.02
+ $Y=1.84 $X2=13.17 $Y2=1.985
r23 1 7 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=13.035
+ $Y=0.37 $X2=13.175 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__DFBBN_1%VGND 1 2 3 4 5 6 21 25 29 33 37 41 43 45 50
+ 55 63 71 76 83 84 87 90 93 96 99 102
r130 102 103 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.72 $Y=0
+ $X2=12.72 $Y2=0
r131 99 100 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.28 $Y=0
+ $X2=11.28 $Y2=0
r132 96 97 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=8.88 $Y=0
+ $X2=8.88 $Y2=0
r133 93 94 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=0 $X2=6 $Y2=0
r134 90 91 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r135 87 88 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r136 84 103 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=13.2 $Y=0
+ $X2=12.72 $Y2=0
r137 83 84 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.2 $Y=0 $X2=13.2
+ $Y2=0
r138 81 102 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=12.83 $Y=0
+ $X2=12.705 $Y2=0
r139 81 83 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=12.83 $Y=0 $X2=13.2
+ $Y2=0
r140 80 103 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.24 $Y=0
+ $X2=12.72 $Y2=0
r141 80 100 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=12.24 $Y=0
+ $X2=11.28 $Y2=0
r142 79 80 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=12.24 $Y=0
+ $X2=12.24 $Y2=0
r143 77 99 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.385 $Y=0
+ $X2=11.22 $Y2=0
r144 77 79 55.7807 $w=1.68e-07 $l=8.55e-07 $layer=LI1_cond $X=11.385 $Y=0
+ $X2=12.24 $Y2=0
r145 76 102 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=12.58 $Y=0
+ $X2=12.705 $Y2=0
r146 76 79 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=12.58 $Y=0
+ $X2=12.24 $Y2=0
r147 75 100 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.8 $Y=0
+ $X2=11.28 $Y2=0
r148 75 97 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=10.8 $Y=0
+ $X2=8.88 $Y2=0
r149 74 75 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=10.8 $Y=0
+ $X2=10.8 $Y2=0
r150 72 96 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.885 $Y=0 $X2=8.8
+ $Y2=0
r151 72 74 124.936 $w=1.68e-07 $l=1.915e-06 $layer=LI1_cond $X=8.885 $Y=0
+ $X2=10.8 $Y2=0
r152 71 99 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.055 $Y=0
+ $X2=11.22 $Y2=0
r153 71 74 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=11.055 $Y=0
+ $X2=10.8 $Y2=0
r154 70 97 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=0 $X2=8.88
+ $Y2=0
r155 69 70 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r156 67 94 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=0 $X2=6
+ $Y2=0
r157 66 69 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=6.48 $Y=0 $X2=8.4
+ $Y2=0
r158 66 67 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6.48 $Y=0
+ $X2=6.48 $Y2=0
r159 64 93 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.145 $Y=0 $X2=5.98
+ $Y2=0
r160 64 66 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=6.145 $Y=0
+ $X2=6.48 $Y2=0
r161 63 96 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.715 $Y=0 $X2=8.8
+ $Y2=0
r162 63 69 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=8.715 $Y=0 $X2=8.4
+ $Y2=0
r163 62 94 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=6
+ $Y2=0
r164 61 62 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=5.52 $Y=0
+ $X2=5.52 $Y2=0
r165 59 62 0.802756 $w=4.9e-07 $l=2.88e-06 $layer=MET1_cond $X=2.64 $Y=0
+ $X2=5.52 $Y2=0
r166 59 91 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=2.16
+ $Y2=0
r167 58 61 187.893 $w=1.68e-07 $l=2.88e-06 $layer=LI1_cond $X=2.64 $Y=0 $X2=5.52
+ $Y2=0
r168 58 59 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=2.64 $Y=0
+ $X2=2.64 $Y2=0
r169 56 90 9.23004 $w=1.7e-07 $l=1.83e-07 $layer=LI1_cond $X=2.41 $Y=0 $X2=2.227
+ $Y2=0
r170 56 58 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=2.41 $Y=0 $X2=2.64
+ $Y2=0
r171 55 93 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.815 $Y=0 $X2=5.98
+ $Y2=0
r172 55 61 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=5.815 $Y=0 $X2=5.52
+ $Y2=0
r173 54 91 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r174 54 88 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=0.72
+ $Y2=0
r175 53 54 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r176 51 87 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.875 $Y=0 $X2=0.71
+ $Y2=0
r177 51 53 52.5187 $w=1.68e-07 $l=8.05e-07 $layer=LI1_cond $X=0.875 $Y=0
+ $X2=1.68 $Y2=0
r178 50 90 9.23004 $w=1.7e-07 $l=1.82e-07 $layer=LI1_cond $X=2.045 $Y=0
+ $X2=2.227 $Y2=0
r179 50 53 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=2.045 $Y=0
+ $X2=1.68 $Y2=0
r180 48 88 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r181 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r182 45 87 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.545 $Y=0 $X2=0.71
+ $Y2=0
r183 45 47 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.545 $Y=0
+ $X2=0.24 $Y2=0
r184 43 70 0.468274 $w=4.9e-07 $l=1.68e-06 $layer=MET1_cond $X=6.72 $Y=0 $X2=8.4
+ $Y2=0
r185 43 67 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=6.72 $Y=0
+ $X2=6.48 $Y2=0
r186 39 102 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=12.705 $Y=0.085
+ $X2=12.705 $Y2=0
r187 39 41 22.8184 $w=2.48e-07 $l=4.95e-07 $layer=LI1_cond $X=12.705 $Y=0.085
+ $X2=12.705 $Y2=0.58
r188 35 99 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=11.22 $Y=0.085
+ $X2=11.22 $Y2=0
r189 35 37 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=11.22 $Y=0.085
+ $X2=11.22 $Y2=0.34
r190 31 96 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.8 $Y=0.085 $X2=8.8
+ $Y2=0
r191 31 33 30.9893 $w=1.68e-07 $l=4.75e-07 $layer=LI1_cond $X=8.8 $Y=0.085
+ $X2=8.8 $Y2=0.56
r192 27 93 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.98 $Y=0.085
+ $X2=5.98 $Y2=0
r193 27 29 27.4142 $w=3.28e-07 $l=7.85e-07 $layer=LI1_cond $X=5.98 $Y=0.085
+ $X2=5.98 $Y2=0.87
r194 23 90 1.2012 $w=3.65e-07 $l=8.5e-08 $layer=LI1_cond $X=2.227 $Y=0.085
+ $X2=2.227 $Y2=0
r195 23 25 13.261 $w=3.63e-07 $l=4.2e-07 $layer=LI1_cond $X=2.227 $Y=0.085
+ $X2=2.227 $Y2=0.505
r196 19 87 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.71 $Y=0.085
+ $X2=0.71 $Y2=0
r197 19 21 18.8582 $w=3.28e-07 $l=5.4e-07 $layer=LI1_cond $X=0.71 $Y=0.085
+ $X2=0.71 $Y2=0.625
r198 6 41 182 $w=1.7e-07 $l=2.95212e-07 $layer=licon1_NDIFF $count=1 $X=12.54
+ $Y=0.37 $X2=12.745 $Y2=0.58
r199 5 37 182 $w=1.7e-07 $l=4.97041e-07 $layer=licon1_NDIFF $count=1 $X=11.015
+ $Y=0.745 $X2=11.22 $Y2=0.34
r200 4 33 182 $w=1.7e-07 $l=4.19196e-07 $layer=licon1_NDIFF $count=1 $X=8.445
+ $Y=0.7 $X2=8.8 $Y2=0.56
r201 3 29 182 $w=1.7e-07 $l=3.65205e-07 $layer=licon1_NDIFF $count=1 $X=5.77
+ $Y=0.595 $X2=5.98 $Y2=0.87
r202 2 25 182 $w=1.7e-07 $l=2.7636e-07 $layer=licon1_NDIFF $count=1 $X=1.99
+ $Y=0.595 $X2=2.225 $Y2=0.505
r203 1 21 182 $w=1.7e-07 $l=3.17372e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.37 $X2=0.71 $Y2=0.625
.ends

.subckt PM_SKY130_FD_SC_HS__DFBBN_1%A_867_119# 1 2 9 11 12 15
r29 13 15 15.5405 $w=3.28e-07 $l=4.45e-07 $layer=LI1_cond $X=5.48 $Y=0.425
+ $X2=5.48 $Y2=0.87
r30 11 13 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=5.315 $Y=0.34
+ $X2=5.48 $Y2=0.425
r31 11 12 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.315 $Y=0.34
+ $X2=4.645 $Y2=0.34
r32 7 12 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.48 $Y=0.425
+ $X2=4.645 $Y2=0.34
r33 7 9 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=4.48 $Y=0.425
+ $X2=4.48 $Y2=0.74
r34 2 15 182 $w=1.7e-07 $l=3.65205e-07 $layer=licon1_NDIFF $count=1 $X=5.27
+ $Y=0.595 $X2=5.48 $Y2=0.87
r35 1 9 182 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=1 $X=4.335
+ $Y=0.595 $X2=4.48 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HS__DFBBN_1%A_1818_76# 1 2 9 11 13
c20 9 0 5.09967e-20 $X=9.23 $Y=0.56
c21 1 0 3.13464e-19 $X=9.09 $Y=0.38
r22 11 13 57.4118 $w=1.68e-07 $l=8.8e-07 $layer=LI1_cond $X=9.315 $Y=0.34
+ $X2=10.195 $Y2=0.34
r23 7 11 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=9.19 $Y=0.425
+ $X2=9.315 $Y2=0.34
r24 7 9 6.22319 $w=2.48e-07 $l=1.35e-07 $layer=LI1_cond $X=9.19 $Y=0.425
+ $X2=9.19 $Y2=0.56
r25 2 13 182 $w=1.7e-07 $l=2.24109e-07 $layer=licon1_NDIFF $count=1 $X=9.99
+ $Y=0.38 $X2=10.195 $Y2=0.34
r26 1 9 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=9.09 $Y=0.38
+ $X2=9.23 $Y2=0.56
.ends

