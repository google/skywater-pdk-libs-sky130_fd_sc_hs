* File: sky130_fd_sc_hs__inv_8.spice
* Created: Tue Sep  1 20:07:11 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hs__inv_8.pex.spice"
.subckt sky130_fd_sc_hs__inv_8  VNB VPB A VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A	A
* VPB	VPB
* VNB	VNB
MM1000 N_VGND_M1000_d N_A_M1000_g N_Y_M1000_s VNB NLOWVT L=0.15 W=0.74 AD=0.2109
+ AS=0.1036 PD=2.05 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2 SB=75003.4
+ A=0.111 P=1.78 MULT=1
MM1001 N_VGND_M1001_d N_A_M1001_g N_Y_M1000_s VNB NLOWVT L=0.15 W=0.74 AD=0.1036
+ AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.6 SB=75003
+ A=0.111 P=1.78 MULT=1
MM1004 N_VGND_M1001_d N_A_M1004_g N_Y_M1004_s VNB NLOWVT L=0.15 W=0.74 AD=0.1036
+ AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.1 SB=75002.6
+ A=0.111 P=1.78 MULT=1
MM1007 N_VGND_M1007_d N_A_M1007_g N_Y_M1004_s VNB NLOWVT L=0.15 W=0.74 AD=0.1295
+ AS=0.1036 PD=1.09 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.5 SB=75002.1
+ A=0.111 P=1.78 MULT=1
MM1012 N_VGND_M1007_d N_A_M1012_g N_Y_M1012_s VNB NLOWVT L=0.15 W=0.74 AD=0.1295
+ AS=0.1036 PD=1.09 PS=1.02 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75002 SB=75001.6
+ A=0.111 P=1.78 MULT=1
MM1013 N_VGND_M1013_d N_A_M1013_g N_Y_M1012_s VNB NLOWVT L=0.15 W=0.74 AD=0.1554
+ AS=0.1036 PD=1.16 PS=1.02 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75002.4 SB=75001.2
+ A=0.111 P=1.78 MULT=1
MM1014 N_VGND_M1013_d N_A_M1014_g N_Y_M1014_s VNB NLOWVT L=0.15 W=0.74 AD=0.1554
+ AS=0.1036 PD=1.16 PS=1.02 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75003 SB=75000.6
+ A=0.111 P=1.78 MULT=1
MM1015 N_VGND_M1015_d N_A_M1015_g N_Y_M1014_s VNB NLOWVT L=0.15 W=0.74 AD=0.2146
+ AS=0.1036 PD=2.06 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75003.4 SB=75000.2
+ A=0.111 P=1.78 MULT=1
MM1002 N_VPWR_M1002_d N_A_M1002_g N_Y_M1002_s VPB PSHORT L=0.15 W=1.12 AD=0.3304
+ AS=0.168 PD=2.83 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667 SA=75000.2
+ SB=75003.5 A=0.168 P=2.54 MULT=1
MM1003 N_VPWR_M1003_d N_A_M1003_g N_Y_M1002_s VPB PSHORT L=0.15 W=1.12 AD=0.196
+ AS=0.168 PD=1.47 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667 SA=75000.7
+ SB=75003.1 A=0.168 P=2.54 MULT=1
MM1005 N_VPWR_M1003_d N_A_M1005_g N_Y_M1005_s VPB PSHORT L=0.15 W=1.12 AD=0.196
+ AS=0.168 PD=1.47 PS=1.42 NRD=10.5395 NRS=1.7533 M=1 R=7.46667 SA=75001.2
+ SB=75002.6 A=0.168 P=2.54 MULT=1
MM1006 N_VPWR_M1006_d N_A_M1006_g N_Y_M1005_s VPB PSHORT L=0.15 W=1.12 AD=0.168
+ AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667 SA=75001.6
+ SB=75002.1 A=0.168 P=2.54 MULT=1
MM1008 N_VPWR_M1006_d N_A_M1008_g N_Y_M1008_s VPB PSHORT L=0.15 W=1.12 AD=0.168
+ AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667 SA=75002.1
+ SB=75001.7 A=0.168 P=2.54 MULT=1
MM1009 N_VPWR_M1009_d N_A_M1009_g N_Y_M1008_s VPB PSHORT L=0.15 W=1.12 AD=0.196
+ AS=0.168 PD=1.47 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667 SA=75002.5
+ SB=75001.2 A=0.168 P=2.54 MULT=1
MM1010 N_VPWR_M1009_d N_A_M1010_g N_Y_M1010_s VPB PSHORT L=0.15 W=1.12 AD=0.196
+ AS=0.168 PD=1.47 PS=1.42 NRD=10.5395 NRS=1.7533 M=1 R=7.46667 SA=75003
+ SB=75000.7 A=0.168 P=2.54 MULT=1
MM1011 N_VPWR_M1011_d N_A_M1011_g N_Y_M1010_s VPB PSHORT L=0.15 W=1.12 AD=0.3864
+ AS=0.168 PD=2.93 PS=1.42 NRD=10.5395 NRS=1.7533 M=1 R=7.46667 SA=75003.5
+ SB=75000.3 A=0.168 P=2.54 MULT=1
DX16_noxref VNB VPB NWDIODE A=8.742 P=13.12
*
.include "sky130_fd_sc_hs__inv_8.pxi.spice"
*
.ends
*
*
