* File: sky130_fd_sc_hs__fahcin_1.spice
* Created: Thu Aug 27 20:46:36 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hs__fahcin_1.pex.spice"
.subckt sky130_fd_sc_hs__fahcin_1  VNB VPB A B CIN VPWR COUT SUM VGND
* 
* VGND	VGND
* SUM	SUM
* COUT	COUT
* VPWR	VPWR
* CIN	CIN
* B	B
* A	A
* VPB	VPB
* VNB	VNB
MM1017 N_VGND_M1017_d N_A_M1017_g N_A_28_74#_M1017_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.279859 AS=0.2109 PD=1.6087 PS=2.05 NRD=11.34 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75001 A=0.111 P=1.78 MULT=1
MM1008 N_A_256_368#_M1008_d N_A_28_74#_M1008_g N_VGND_M1017_d VNB NLOWVT L=0.15
+ W=0.64 AD=0.1824 AS=0.242041 PD=1.85 PS=1.3913 NRD=0 NRS=76.872 M=1 R=4.26667
+ SA=75001.1 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1014 N_A_28_74#_M1014_d N_A_492_48#_M1014_g N_A_430_418#_M1014_s VNB NLOWVT
+ L=0.15 W=0.64 AD=0.0896 AS=0.1696 PD=0.92 PS=1.81 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75001.5 A=0.096 P=1.58 MULT=1
MM1006 N_A_608_74#_M1006_d N_B_M1006_g N_A_28_74#_M1014_d VNB NLOWVT L=0.15
+ W=0.64 AD=0.170162 AS=0.0896 PD=1.395 PS=0.92 NRD=46.872 NRS=0 M=1 R=4.26667
+ SA=75000.6 SB=75001.1 A=0.096 P=1.58 MULT=1
MM1025 N_A_256_368#_M1025_d N_A_492_48#_M1025_g N_A_608_74#_M1006_d VNB NLOWVT
+ L=0.15 W=0.64 AD=0.1632 AS=0.170162 PD=1.15 PS=1.395 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.9 SB=75000.9 A=0.096 P=1.58 MULT=1
MM1031 N_A_430_418#_M1031_d N_B_M1031_g N_A_256_368#_M1025_d VNB NLOWVT L=0.15
+ W=0.64 AD=0.1952 AS=0.1632 PD=1.89 PS=1.15 NRD=3.744 NRS=43.116 M=1 R=4.26667
+ SA=75001.6 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1015 N_VGND_M1015_d N_B_M1015_g N_A_492_48#_M1015_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.212455 AS=0.222 PD=1.41565 PS=2.08 NRD=22.692 NRS=2.424 M=1 R=4.93333
+ SA=75000.2 SB=75005 A=0.111 P=1.78 MULT=1
MM1027 N_A_1197_368#_M1027_d N_A_492_48#_M1027_g N_VGND_M1015_d VNB NLOWVT
+ L=0.15 W=0.64 AD=0.0896 AS=0.183745 PD=0.92 PS=1.22435 NRD=0 NRS=29.988 M=1
+ R=4.26667 SA=75001 SB=75005.1 A=0.096 P=1.58 MULT=1
MM1002 N_COUT_M1002_d N_A_430_418#_M1002_g N_A_1197_368#_M1027_d VNB NLOWVT
+ L=0.15 W=0.64 AD=0.4528 AS=0.0896 PD=2.055 PS=0.92 NRD=13.116 NRS=0 M=1
+ R=4.26667 SA=75001.4 SB=75004.6 A=0.096 P=1.58 MULT=1
MM1023 N_A_1595_400#_M1023_d N_A_608_74#_M1023_g N_COUT_M1002_d VNB NLOWVT
+ L=0.15 W=0.64 AD=0.112 AS=0.4528 PD=0.99 PS=2.055 NRD=13.116 NRS=0 M=1
+ R=4.26667 SA=75002.9 SB=75003.1 A=0.096 P=1.58 MULT=1
MM1019 N_VGND_M1019_d N_CIN_M1019_g N_A_1595_400#_M1023_d VNB NLOWVT L=0.15
+ W=0.64 AD=0.220012 AS=0.112 PD=1.53043 PS=0.99 NRD=14.052 NRS=0 M=1 R=4.26667
+ SA=75003.4 SB=75002.6 A=0.096 P=1.58 MULT=1
MM1003 N_A_1854_368#_M1003_d N_CIN_M1003_g N_VGND_M1019_d VNB NLOWVT L=0.15
+ W=0.74 AD=0.124942 AS=0.254388 PD=1.14217 PS=1.76957 NRD=5.664 NRS=62.016 M=1
+ R=4.93333 SA=75002.8 SB=75002.6 A=0.111 P=1.78 MULT=1
MM1018 N_A_2004_136#_M1018_d N_A_608_74#_M1018_g N_A_1854_368#_M1003_d VNB
+ NLOWVT L=0.15 W=0.64 AD=0.2544 AS=0.108058 PD=1.435 PS=0.987826 NRD=14.052
+ NRS=1.872 M=1 R=4.26667 SA=75003 SB=75002.5 A=0.096 P=1.58 MULT=1
MM1009 N_A_1967_384#_M1009_d N_A_430_418#_M1009_g N_A_2004_136#_M1018_d VNB
+ NLOWVT L=0.15 W=0.64 AD=0.1404 AS=0.2544 PD=1.145 PS=1.435 NRD=27.648 NRS=0
+ M=1 R=4.26667 SA=75004 SB=75001.6 A=0.096 P=1.58 MULT=1
MM1001 N_VGND_M1001_d N_A_1854_368#_M1001_g N_A_1967_384#_M1009_d VNB NLOWVT
+ L=0.15 W=0.64 AD=0.276638 AS=0.1404 PD=1.47478 PS=1.145 NRD=78.744 NRS=0 M=1
+ R=4.26667 SA=75004.3 SB=75001.2 A=0.096 P=1.58 MULT=1
MM1020 N_SUM_M1020_d N_A_2004_136#_M1020_g N_VGND_M1001_d VNB NLOWVT L=0.15
+ W=0.74 AD=0.2109 AS=0.319862 PD=2.05 PS=1.70522 NRD=0 NRS=25.128 M=1 R=4.93333
+ SA=75004.6 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1005 N_VPWR_M1005_d N_A_M1005_g N_A_28_74#_M1005_s VPB PSHORT L=0.15 W=1.12
+ AD=0.303985 AS=0.3304 PD=1.75396 PS=2.83 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75000.8 A=0.168 P=2.54 MULT=1
MM1000 N_A_256_368#_M1000_d N_A_28_74#_M1000_g N_VPWR_M1005_d VPB PSHORT L=0.15
+ W=1 AD=0.295 AS=0.271415 PD=2.59 PS=1.56604 NRD=1.9503 NRS=49.5652 M=1
+ R=6.66667 SA=75000.9 SB=75000.2 A=0.15 P=2.3 MULT=1
MM1011 N_A_256_368#_M1011_d N_A_492_48#_M1011_g N_A_430_418#_M1011_s VPB PSHORT
+ L=0.15 W=0.84 AD=0.1428 AS=0.273 PD=1.18 PS=2.33 NRD=11.7215 NRS=3.5066 M=1
+ R=5.6 SA=75000.2 SB=75001.7 A=0.126 P=1.98 MULT=1
MM1029 N_A_608_74#_M1029_d N_B_M1029_g N_A_256_368#_M1011_d VPB PSHORT L=0.15
+ W=0.84 AD=0.178762 AS=0.1428 PD=1.42 PS=1.18 NRD=58.6272 NRS=0 M=1 R=5.6
+ SA=75000.7 SB=75001.2 A=0.126 P=1.98 MULT=1
MM1021 N_A_28_74#_M1021_d N_A_492_48#_M1021_g N_A_608_74#_M1029_d VPB PSHORT
+ L=0.15 W=0.84 AD=0.2373 AS=0.178762 PD=1.405 PS=1.42 NRD=14.0658 NRS=2.3443
+ M=1 R=5.6 SA=75001 SB=75001 A=0.126 P=1.98 MULT=1
MM1016 N_A_430_418#_M1016_d N_B_M1016_g N_A_28_74#_M1021_d VPB PSHORT L=0.15
+ W=0.84 AD=0.2604 AS=0.2373 PD=2.3 PS=1.405 NRD=5.8509 NRS=52.7566 M=1 R=5.6
+ SA=75001.7 SB=75000.2 A=0.126 P=1.98 MULT=1
MM1007 N_VPWR_M1007_d N_B_M1007_g N_A_492_48#_M1007_s VPB PSHORT L=0.15 W=1.12
+ AD=0.239849 AS=0.3304 PD=1.62189 PS=2.83 NRD=4.3931 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75003.2 A=0.168 P=2.54 MULT=1
MM1012 N_A_1197_368#_M1012_d N_A_492_48#_M1012_g N_VPWR_M1007_d VPB PSHORT
+ L=0.15 W=1 AD=0.224239 AS=0.214151 PD=1.55978 PS=1.44811 NRD=1.9503
+ NRS=22.6353 M=1 R=6.66667 SA=75000.8 SB=75003 A=0.15 P=2.3 MULT=1
MM1030 N_COUT_M1030_d N_A_608_74#_M1030_g N_A_1197_368#_M1012_d VPB PSHORT
+ L=0.15 W=0.84 AD=0.5271 AS=0.188361 PD=2.095 PS=1.31022 NRD=49.2303
+ NRS=35.1645 M=1 R=5.6 SA=75001.4 SB=75002.9 A=0.126 P=1.98 MULT=1
MM1026 N_A_1595_400#_M1026_d N_A_430_418#_M1026_g N_COUT_M1030_d VPB PSHORT
+ L=0.15 W=0.84 AD=0.194296 AS=0.5271 PD=1.31478 PS=2.095 NRD=22.852 NRS=43.3794
+ M=1 R=5.6 SA=75002.8 SB=75001.5 A=0.126 P=1.98 MULT=1
MM1004 N_VPWR_M1004_d N_CIN_M1004_g N_A_1595_400#_M1026_d VPB PSHORT L=0.15 W=1
+ AD=0.278491 AS=0.231304 PD=1.58019 PS=1.56522 NRD=52.6975 NRS=12.7853 M=1
+ R=6.66667 SA=75002.9 SB=75000.9 A=0.15 P=2.3 MULT=1
MM1010 N_A_1854_368#_M1010_d N_CIN_M1010_g N_VPWR_M1004_d VPB PSHORT L=0.15
+ W=1.12 AD=0.3304 AS=0.311909 PD=2.83 PS=1.76981 NRD=1.7533 NRS=1.7533 M=1
+ R=7.46667 SA=75003.2 SB=75000.2 A=0.168 P=2.54 MULT=1
MM1024 N_A_2004_136#_M1024_d N_A_608_74#_M1024_g N_A_1967_384#_M1024_s VPB
+ PSHORT L=0.15 W=0.84 AD=0.126 AS=0.2478 PD=1.14 PS=2.27 NRD=2.3443 NRS=2.3443
+ M=1 R=5.6 SA=75000.2 SB=75000.8 A=0.126 P=1.98 MULT=1
MM1028 N_A_1854_368#_M1028_d N_A_430_418#_M1028_g N_A_2004_136#_M1024_d VPB
+ PSHORT L=0.15 W=0.84 AD=0.43155 AS=0.126 PD=3.07 PS=1.14 NRD=107.582
+ NRS=2.3443 M=1 R=5.6 SA=75000.7 SB=75000.3 A=0.126 P=1.98 MULT=1
MM1013 N_VPWR_M1013_d N_A_1854_368#_M1013_g N_A_1967_384#_M1013_s VPB PSHORT
+ L=0.15 W=1 AD=0.266698 AS=0.295 PD=1.5566 PS=2.59 NRD=47.5952 NRS=1.9503 M=1
+ R=6.66667 SA=75000.2 SB=75000.9 A=0.15 P=2.3 MULT=1
MM1022 N_SUM_M1022_d N_A_2004_136#_M1022_g N_VPWR_M1013_d VPB PSHORT L=0.15
+ W=1.12 AD=0.3304 AS=0.298702 PD=2.83 PS=1.7434 NRD=1.7533 NRS=1.7533 M=1
+ R=7.46667 SA=75000.8 SB=75000.2 A=0.168 P=2.54 MULT=1
DX32_noxref VNB VPB NWDIODE A=24.8124 P=30.4
c_119 VNB 0 2.57866e-19 $X=0 $Y=0
*
.include "sky130_fd_sc_hs__fahcin_1.pxi.spice"
*
.ends
*
*
