* File: sky130_fd_sc_hs__dfrtp_1.pxi.spice
* Created: Tue Sep  1 19:59:57 2020
* 
x_PM_SKY130_FD_SC_HS__DFRTP_1%D N_D_c_236_n N_D_c_241_n N_D_c_242_n N_D_M1013_g
+ N_D_M1025_g D D D N_D_c_238_n N_D_c_239_n N_D_c_244_n
+ PM_SKY130_FD_SC_HS__DFRTP_1%D
x_PM_SKY130_FD_SC_HS__DFRTP_1%RESET_B N_RESET_B_M1016_g N_RESET_B_c_269_n
+ N_RESET_B_c_277_n N_RESET_B_c_278_n N_RESET_B_M1014_g N_RESET_B_c_270_n
+ N_RESET_B_M1010_g N_RESET_B_c_279_n N_RESET_B_M1029_g N_RESET_B_c_271_n
+ N_RESET_B_M1002_g N_RESET_B_c_282_n N_RESET_B_M1000_g N_RESET_B_c_273_n
+ N_RESET_B_c_283_n N_RESET_B_c_284_n N_RESET_B_c_285_n N_RESET_B_c_286_n
+ N_RESET_B_c_287_n N_RESET_B_c_288_n RESET_B N_RESET_B_c_274_n
+ N_RESET_B_c_275_n N_RESET_B_c_290_n N_RESET_B_c_291_n N_RESET_B_c_292_n
+ PM_SKY130_FD_SC_HS__DFRTP_1%RESET_B
x_PM_SKY130_FD_SC_HS__DFRTP_1%CLK N_CLK_M1003_g N_CLK_c_470_n N_CLK_M1005_g CLK
+ PM_SKY130_FD_SC_HS__DFRTP_1%CLK
x_PM_SKY130_FD_SC_HS__DFRTP_1%A_490_366# N_A_490_366#_M1030_d
+ N_A_490_366#_M1008_d N_A_490_366#_c_531_n N_A_490_366#_c_532_n
+ N_A_490_366#_M1012_g N_A_490_366#_c_512_n N_A_490_366#_c_513_n
+ N_A_490_366#_M1001_g N_A_490_366#_c_515_n N_A_490_366#_M1026_g
+ N_A_490_366#_c_516_n N_A_490_366#_c_517_n N_A_490_366#_c_535_n
+ N_A_490_366#_M1023_g N_A_490_366#_c_536_n N_A_490_366#_c_518_n
+ N_A_490_366#_c_519_n N_A_490_366#_c_537_n N_A_490_366#_c_520_n
+ N_A_490_366#_c_521_n N_A_490_366#_c_554_p N_A_490_366#_c_522_n
+ N_A_490_366#_c_523_n N_A_490_366#_c_524_n N_A_490_366#_c_525_n
+ N_A_490_366#_c_526_n N_A_490_366#_c_527_n N_A_490_366#_c_528_n
+ N_A_490_366#_c_529_n N_A_490_366#_c_530_n
+ PM_SKY130_FD_SC_HS__DFRTP_1%A_490_366#
x_PM_SKY130_FD_SC_HS__DFRTP_1%A_830_359# N_A_830_359#_M1031_d
+ N_A_830_359#_M1017_d N_A_830_359#_c_717_n N_A_830_359#_M1007_g
+ N_A_830_359#_M1018_g N_A_830_359#_c_714_n N_A_830_359#_c_732_n
+ N_A_830_359#_c_748_n N_A_830_359#_c_720_n N_A_830_359#_c_715_n
+ N_A_830_359#_c_716_n PM_SKY130_FD_SC_HS__DFRTP_1%A_830_359#
x_PM_SKY130_FD_SC_HS__DFRTP_1%A_695_457# N_A_695_457#_M1004_d
+ N_A_695_457#_M1012_d N_A_695_457#_M1029_d N_A_695_457#_M1031_g
+ N_A_695_457#_c_806_n N_A_695_457#_M1017_g N_A_695_457#_c_800_n
+ N_A_695_457#_c_816_n N_A_695_457#_c_808_n N_A_695_457#_c_801_n
+ N_A_695_457#_c_802_n N_A_695_457#_c_803_n N_A_695_457#_c_804_n
+ N_A_695_457#_c_811_n N_A_695_457#_c_805_n N_A_695_457#_c_840_n
+ PM_SKY130_FD_SC_HS__DFRTP_1%A_695_457#
x_PM_SKY130_FD_SC_HS__DFRTP_1%A_306_74# N_A_306_74#_M1003_s N_A_306_74#_M1005_s
+ N_A_306_74#_c_939_n N_A_306_74#_M1008_g N_A_306_74#_c_926_n
+ N_A_306_74#_M1030_g N_A_306_74#_c_927_n N_A_306_74#_c_928_n
+ N_A_306_74#_c_929_n N_A_306_74#_c_942_n N_A_306_74#_c_943_n
+ N_A_306_74#_c_930_n N_A_306_74#_M1004_g N_A_306_74#_c_944_n
+ N_A_306_74#_c_945_n N_A_306_74#_c_946_n N_A_306_74#_M1015_g
+ N_A_306_74#_c_947_n N_A_306_74#_M1022_g N_A_306_74#_c_931_n
+ N_A_306_74#_c_932_n N_A_306_74#_M1020_g N_A_306_74#_c_951_n
+ N_A_306_74#_c_952_n N_A_306_74#_c_934_n N_A_306_74#_c_935_n
+ N_A_306_74#_c_936_n N_A_306_74#_c_937_n N_A_306_74#_c_938_n
+ N_A_306_74#_c_954_n PM_SKY130_FD_SC_HS__DFRTP_1%A_306_74#
x_PM_SKY130_FD_SC_HS__DFRTP_1%A_1518_203# N_A_1518_203#_M1021_d
+ N_A_1518_203#_M1000_d N_A_1518_203#_c_1124_n N_A_1518_203#_c_1125_n
+ N_A_1518_203#_c_1126_n N_A_1518_203#_M1011_g N_A_1518_203#_M1019_g
+ N_A_1518_203#_c_1117_n N_A_1518_203#_c_1118_n N_A_1518_203#_c_1119_n
+ N_A_1518_203#_c_1128_n N_A_1518_203#_c_1129_n N_A_1518_203#_c_1120_n
+ N_A_1518_203#_c_1121_n N_A_1518_203#_c_1122_n N_A_1518_203#_c_1131_n
+ N_A_1518_203#_c_1132_n N_A_1518_203#_c_1123_n
+ PM_SKY130_FD_SC_HS__DFRTP_1%A_1518_203#
x_PM_SKY130_FD_SC_HS__DFRTP_1%A_1266_74# N_A_1266_74#_M1026_d
+ N_A_1266_74#_M1022_d N_A_1266_74#_M1021_g N_A_1266_74#_c_1249_n
+ N_A_1266_74#_c_1250_n N_A_1266_74#_M1006_g N_A_1266_74#_c_1236_n
+ N_A_1266_74#_c_1237_n N_A_1266_74#_c_1238_n N_A_1266_74#_c_1253_n
+ N_A_1266_74#_c_1254_n N_A_1266_74#_M1028_g N_A_1266_74#_c_1239_n
+ N_A_1266_74#_c_1240_n N_A_1266_74#_c_1241_n N_A_1266_74#_M1027_g
+ N_A_1266_74#_c_1242_n N_A_1266_74#_c_1283_n N_A_1266_74#_c_1243_n
+ N_A_1266_74#_c_1256_n N_A_1266_74#_c_1244_n N_A_1266_74#_c_1269_n
+ N_A_1266_74#_c_1379_p N_A_1266_74#_c_1257_n N_A_1266_74#_c_1245_n
+ N_A_1266_74#_c_1246_n N_A_1266_74#_c_1247_n N_A_1266_74#_c_1248_n
+ PM_SKY130_FD_SC_HS__DFRTP_1%A_1266_74#
x_PM_SKY130_FD_SC_HS__DFRTP_1%A_1864_409# N_A_1864_409#_M1027_d
+ N_A_1864_409#_M1028_d N_A_1864_409#_c_1401_n N_A_1864_409#_M1024_g
+ N_A_1864_409#_M1009_g N_A_1864_409#_c_1397_n N_A_1864_409#_c_1398_n
+ N_A_1864_409#_c_1404_n N_A_1864_409#_c_1399_n N_A_1864_409#_c_1400_n
+ PM_SKY130_FD_SC_HS__DFRTP_1%A_1864_409#
x_PM_SKY130_FD_SC_HS__DFRTP_1%VPWR N_VPWR_M1013_s N_VPWR_M1014_d N_VPWR_M1005_d
+ N_VPWR_M1007_d N_VPWR_M1017_s N_VPWR_M1011_d N_VPWR_M1006_d N_VPWR_M1024_d
+ N_VPWR_c_1451_n N_VPWR_c_1452_n N_VPWR_c_1453_n N_VPWR_c_1454_n
+ N_VPWR_c_1455_n N_VPWR_c_1456_n N_VPWR_c_1457_n N_VPWR_c_1458_n
+ N_VPWR_c_1459_n N_VPWR_c_1460_n N_VPWR_c_1461_n N_VPWR_c_1462_n VPWR
+ N_VPWR_c_1463_n N_VPWR_c_1464_n N_VPWR_c_1465_n N_VPWR_c_1466_n
+ N_VPWR_c_1467_n N_VPWR_c_1468_n N_VPWR_c_1469_n N_VPWR_c_1470_n
+ N_VPWR_c_1471_n N_VPWR_c_1472_n N_VPWR_c_1473_n N_VPWR_c_1450_n
+ PM_SKY130_FD_SC_HS__DFRTP_1%VPWR
x_PM_SKY130_FD_SC_HS__DFRTP_1%A_30_78# N_A_30_78#_M1025_s N_A_30_78#_M1004_s
+ N_A_30_78#_M1013_d N_A_30_78#_M1012_s N_A_30_78#_c_1590_n N_A_30_78#_c_1591_n
+ N_A_30_78#_c_1597_n N_A_30_78#_c_1592_n N_A_30_78#_c_1598_n
+ N_A_30_78#_c_1593_n N_A_30_78#_c_1594_n N_A_30_78#_c_1600_n
+ N_A_30_78#_c_1601_n N_A_30_78#_c_1602_n N_A_30_78#_c_1603_n
+ N_A_30_78#_c_1595_n PM_SKY130_FD_SC_HS__DFRTP_1%A_30_78#
x_PM_SKY130_FD_SC_HS__DFRTP_1%Q N_Q_M1009_s N_Q_M1024_s N_Q_c_1715_n
+ N_Q_c_1716_n Q Q Q N_Q_c_1717_n PM_SKY130_FD_SC_HS__DFRTP_1%Q
x_PM_SKY130_FD_SC_HS__DFRTP_1%VGND N_VGND_M1016_d N_VGND_M1003_d N_VGND_M1010_d
+ N_VGND_M1019_d N_VGND_M1027_s N_VGND_M1009_d N_VGND_c_1745_n N_VGND_c_1746_n
+ N_VGND_c_1747_n N_VGND_c_1748_n N_VGND_c_1749_n N_VGND_c_1750_n
+ N_VGND_c_1751_n N_VGND_c_1752_n VGND N_VGND_c_1753_n N_VGND_c_1754_n
+ N_VGND_c_1755_n N_VGND_c_1756_n N_VGND_c_1757_n N_VGND_c_1758_n
+ N_VGND_c_1759_n N_VGND_c_1760_n N_VGND_c_1761_n
+ PM_SKY130_FD_SC_HS__DFRTP_1%VGND
cc_1 VNB N_D_c_236_n 0.0406028f $X=-0.19 $Y=-0.245 $X2=0.402 $Y2=1.828
cc_2 VNB N_D_M1025_g 0.0286471f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=0.6
cc_3 VNB N_D_c_238_n 0.0216279f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.165
cc_4 VNB N_D_c_239_n 0.0281582f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.165
cc_5 VNB N_RESET_B_M1016_g 0.0285646f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.01
cc_6 VNB N_RESET_B_c_269_n 0.0250069f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.75
cc_7 VNB N_RESET_B_c_270_n 0.0155478f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_8 VNB N_RESET_B_c_271_n 0.0176719f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.165
cc_9 VNB N_RESET_B_M1002_g 0.0510668f $X=-0.19 $Y=-0.245 $X2=0.402 $Y2=1.845
cc_10 VNB N_RESET_B_c_273_n 0.0134203f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_RESET_B_c_274_n 0.0343812f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_RESET_B_c_275_n 0.00330649f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_CLK_M1003_g 0.0258498f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.01
cc_14 VNB N_CLK_c_470_n 0.0323697f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.465
cc_15 VNB CLK 0.00636154f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=1
cc_16 VNB N_A_490_366#_c_512_n 0.0101009f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_17 VNB N_A_490_366#_c_513_n 0.0206887f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.95
cc_18 VNB N_A_490_366#_M1001_g 0.0240392f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_490_366#_c_515_n 0.0192767f $X=-0.19 $Y=-0.245 $X2=0.402 $Y2=1.165
cc_20 VNB N_A_490_366#_c_516_n 0.0205614f $X=-0.19 $Y=-0.245 $X2=0.402 $Y2=1
cc_21 VNB N_A_490_366#_c_517_n 0.0110312f $X=-0.19 $Y=-0.245 $X2=0.402 $Y2=1.845
cc_22 VNB N_A_490_366#_c_518_n 0.0105327f $X=-0.19 $Y=-0.245 $X2=0.32 $Y2=1.845
cc_23 VNB N_A_490_366#_c_519_n 0.0380469f $X=-0.19 $Y=-0.245 $X2=0.32 $Y2=2.035
cc_24 VNB N_A_490_366#_c_520_n 0.00138276f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_490_366#_c_521_n 0.00360885f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_490_366#_c_522_n 0.0169659f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_490_366#_c_523_n 9.76919e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_490_366#_c_524_n 0.00385029f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_490_366#_c_525_n 0.0019226f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_490_366#_c_526_n 0.0145565f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_490_366#_c_527_n 0.0120426f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_490_366#_c_528_n 0.0313598f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_490_366#_c_529_n 0.00797767f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_490_366#_c_530_n 0.00958036f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_830_359#_M1018_g 0.0352959f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_36 VNB N_A_830_359#_c_714_n 0.00330276f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_830_359#_c_715_n 0.00275035f $X=-0.19 $Y=-0.245 $X2=0.32 $Y2=1.295
cc_38 VNB N_A_830_359#_c_716_n 0.00947395f $X=-0.19 $Y=-0.245 $X2=0.32 $Y2=1.845
cc_39 VNB N_A_695_457#_M1031_g 0.0226589f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_40 VNB N_A_695_457#_c_800_n 0.00571098f $X=-0.19 $Y=-0.245 $X2=0.402
+ $Y2=1.165
cc_41 VNB N_A_695_457#_c_801_n 0.0011075f $X=-0.19 $Y=-0.245 $X2=0.402 $Y2=1.845
cc_42 VNB N_A_695_457#_c_802_n 0.00289685f $X=-0.19 $Y=-0.245 $X2=0.385
+ $Y2=1.845
cc_43 VNB N_A_695_457#_c_803_n 0.00804496f $X=-0.19 $Y=-0.245 $X2=0.402 $Y2=2.01
cc_44 VNB N_A_695_457#_c_804_n 0.0411633f $X=-0.19 $Y=-0.245 $X2=0.32 $Y2=1.165
cc_45 VNB N_A_695_457#_c_805_n 0.00300764f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_A_306_74#_c_926_n 0.0196868f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=0.6
cc_47 VNB N_A_306_74#_c_927_n 0.00468316f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.95
cc_48 VNB N_A_306_74#_c_928_n 0.0362722f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A_306_74#_c_929_n 0.0569372f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_A_306_74#_c_930_n 0.0179002f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.165
cc_51 VNB N_A_306_74#_c_931_n 0.0226279f $X=-0.19 $Y=-0.245 $X2=0.32 $Y2=2.035
cc_52 VNB N_A_306_74#_c_932_n 0.0014655f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_A_306_74#_M1020_g 0.0517191f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_A_306_74#_c_934_n 0.00994826f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_A_306_74#_c_935_n 0.00952551f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_A_306_74#_c_936_n 0.0033915f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_A_306_74#_c_937_n 0.00172158f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_A_306_74#_c_938_n 0.00486147f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_A_1518_203#_M1019_g 0.0207732f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_A_1518_203#_c_1117_n 0.0156636f $X=-0.19 $Y=-0.245 $X2=0.402
+ $Y2=1.165
cc_61 VNB N_A_1518_203#_c_1118_n 0.0155514f $X=-0.19 $Y=-0.245 $X2=0.385
+ $Y2=1.165
cc_62 VNB N_A_1518_203#_c_1119_n 0.0105463f $X=-0.19 $Y=-0.245 $X2=0.402
+ $Y2=2.01
cc_63 VNB N_A_1518_203#_c_1120_n 0.0023345f $X=-0.19 $Y=-0.245 $X2=0.32
+ $Y2=1.665
cc_64 VNB N_A_1518_203#_c_1121_n 0.00392193f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_A_1518_203#_c_1122_n 0.0310153f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_A_1518_203#_c_1123_n 0.0124417f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_A_1266_74#_M1021_g 0.04091f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=0.6
cc_68 VNB N_A_1266_74#_c_1236_n 0.0182931f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_A_1266_74#_c_1237_n 0.016718f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_A_1266_74#_c_1238_n 0.0126324f $X=-0.19 $Y=-0.245 $X2=0.385
+ $Y2=1.165
cc_71 VNB N_A_1266_74#_c_1239_n 0.0232568f $X=-0.19 $Y=-0.245 $X2=0.402 $Y2=2.01
cc_72 VNB N_A_1266_74#_c_1240_n 0.0100399f $X=-0.19 $Y=-0.245 $X2=0.32 $Y2=1.165
cc_73 VNB N_A_1266_74#_c_1241_n 0.0210614f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_A_1266_74#_c_1242_n 0.0123873f $X=-0.19 $Y=-0.245 $X2=0.32 $Y2=1.665
cc_75 VNB N_A_1266_74#_c_1243_n 0.00445288f $X=-0.19 $Y=-0.245 $X2=0.32
+ $Y2=1.845
cc_76 VNB N_A_1266_74#_c_1244_n 0.00403288f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_A_1266_74#_c_1245_n 0.00637997f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_A_1266_74#_c_1246_n 0.00599516f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VNB N_A_1266_74#_c_1247_n 0.00266453f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_A_1266_74#_c_1248_n 0.00109446f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_81 VNB N_A_1864_409#_M1009_g 0.0383367f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_82 VNB N_A_1864_409#_c_1397_n 0.0564146f $X=-0.19 $Y=-0.245 $X2=0.155
+ $Y2=1.95
cc_83 VNB N_A_1864_409#_c_1398_n 0.0212559f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_84 VNB N_A_1864_409#_c_1399_n 0.014962f $X=-0.19 $Y=-0.245 $X2=0.402
+ $Y2=1.845
cc_85 VNB N_A_1864_409#_c_1400_n 0.00445066f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_86 VNB N_VPWR_c_1450_n 0.462217f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_87 VNB N_A_30_78#_c_1590_n 0.003401f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_88 VNB N_A_30_78#_c_1591_n 0.00542054f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_89 VNB N_A_30_78#_c_1592_n 0.00295332f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.845
cc_90 VNB N_A_30_78#_c_1593_n 0.00365277f $X=-0.19 $Y=-0.245 $X2=0.32 $Y2=1.295
cc_91 VNB N_A_30_78#_c_1594_n 0.0223919f $X=-0.19 $Y=-0.245 $X2=0.32 $Y2=1.665
cc_92 VNB N_A_30_78#_c_1595_n 0.00700512f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_93 VNB N_Q_c_1715_n 0.00811762f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=0.6
cc_94 VNB N_Q_c_1716_n 0.00208381f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_95 VNB N_Q_c_1717_n 0.00535471f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_96 VNB N_VGND_c_1745_n 0.0162008f $X=-0.19 $Y=-0.245 $X2=0.402 $Y2=1
cc_97 VNB N_VGND_c_1746_n 0.00641543f $X=-0.19 $Y=-0.245 $X2=0.402 $Y2=2.01
cc_98 VNB N_VGND_c_1747_n 0.0111809f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_99 VNB N_VGND_c_1748_n 0.0145996f $X=-0.19 $Y=-0.245 $X2=0.32 $Y2=2.035
cc_100 VNB N_VGND_c_1749_n 0.010678f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_101 VNB N_VGND_c_1750_n 0.0505973f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_102 VNB N_VGND_c_1751_n 0.0307721f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_103 VNB N_VGND_c_1752_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_104 VNB N_VGND_c_1753_n 0.0201745f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_105 VNB N_VGND_c_1754_n 0.0818466f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_106 VNB N_VGND_c_1755_n 0.0580863f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_107 VNB N_VGND_c_1756_n 0.0325483f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_108 VNB N_VGND_c_1757_n 0.0345892f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_109 VNB N_VGND_c_1758_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_110 VNB N_VGND_c_1759_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_111 VNB N_VGND_c_1760_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_112 VNB N_VGND_c_1761_n 0.628803f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_113 VPB N_D_c_236_n 0.0142152f $X=-0.19 $Y=1.66 $X2=0.402 $Y2=1.828
cc_114 VPB N_D_c_241_n 0.0278711f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=2.375
cc_115 VPB N_D_c_242_n 0.0266297f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=2.465
cc_116 VPB N_D_c_239_n 0.0243342f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.165
cc_117 VPB N_D_c_244_n 0.0207718f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.845
cc_118 VPB N_RESET_B_c_269_n 0.0211247f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=2.75
cc_119 VPB N_RESET_B_c_277_n 0.0182428f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=1
cc_120 VPB N_RESET_B_c_278_n 0.0236024f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=0.6
cc_121 VPB N_RESET_B_c_279_n 0.0169736f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_122 VPB N_RESET_B_c_271_n 0.0111344f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.165
cc_123 VPB N_RESET_B_M1002_g 0.0151047f $X=-0.19 $Y=1.66 $X2=0.402 $Y2=1.845
cc_124 VPB N_RESET_B_c_282_n 0.0572287f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.845
cc_125 VPB N_RESET_B_c_283_n 0.01931f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_126 VPB N_RESET_B_c_284_n 0.00380287f $X=-0.19 $Y=1.66 $X2=0.32 $Y2=1.845
cc_127 VPB N_RESET_B_c_285_n 0.0198788f $X=-0.19 $Y=1.66 $X2=0.32 $Y2=2.035
cc_128 VPB N_RESET_B_c_286_n 0.00169127f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_129 VPB N_RESET_B_c_287_n 0.00495528f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_130 VPB N_RESET_B_c_288_n 0.00335799f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_131 VPB N_RESET_B_c_275_n 9.70225e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_132 VPB N_RESET_B_c_290_n 0.0304851f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_133 VPB N_RESET_B_c_291_n 0.0539371f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_134 VPB N_RESET_B_c_292_n 0.00620787f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_135 VPB N_CLK_c_470_n 0.0235518f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=2.465
cc_136 VPB CLK 0.00483282f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=1
cc_137 VPB N_A_490_366#_c_531_n 0.0143302f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=1
cc_138 VPB N_A_490_366#_c_532_n 0.0198055f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=0.6
cc_139 VPB N_A_490_366#_c_512_n 0.0099424f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.21
cc_140 VPB N_A_490_366#_c_513_n 0.00567537f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.95
cc_141 VPB N_A_490_366#_c_535_n 0.0624804f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.845
cc_142 VPB N_A_490_366#_c_536_n 0.00298582f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_143 VPB N_A_490_366#_c_537_n 0.00718131f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_144 VPB N_A_490_366#_c_520_n 9.36995e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_145 VPB N_A_490_366#_c_524_n 0.00559228f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_146 VPB N_A_490_366#_c_530_n 0.0192067f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_147 VPB N_A_830_359#_c_717_n 0.0637903f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=2.75
cc_148 VPB N_A_830_359#_M1018_g 0.00868606f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.21
cc_149 VPB N_A_830_359#_c_714_n 0.00245885f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_150 VPB N_A_830_359#_c_720_n 0.00215186f $X=-0.19 $Y=1.66 $X2=0.402 $Y2=2.01
cc_151 VPB N_A_830_359#_c_716_n 0.00382281f $X=-0.19 $Y=1.66 $X2=0.32 $Y2=1.845
cc_152 VPB N_A_695_457#_c_806_n 0.0172536f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.95
cc_153 VPB N_A_695_457#_c_800_n 0.00914592f $X=-0.19 $Y=1.66 $X2=0.402 $Y2=1.165
cc_154 VPB N_A_695_457#_c_808_n 0.00288458f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.165
cc_155 VPB N_A_695_457#_c_801_n 0.00577088f $X=-0.19 $Y=1.66 $X2=0.402 $Y2=1.845
cc_156 VPB N_A_695_457#_c_804_n 0.0241647f $X=-0.19 $Y=1.66 $X2=0.32 $Y2=1.165
cc_157 VPB N_A_695_457#_c_811_n 0.00256103f $X=-0.19 $Y=1.66 $X2=0.32 $Y2=1.665
cc_158 VPB N_A_306_74#_c_939_n 0.0145665f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=2.75
cc_159 VPB N_A_306_74#_c_927_n 0.0780956f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.95
cc_160 VPB N_A_306_74#_c_929_n 0.00705161f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_161 VPB N_A_306_74#_c_942_n 0.0560324f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_162 VPB N_A_306_74#_c_943_n 0.0125195f $X=-0.19 $Y=1.66 $X2=0.402 $Y2=1.165
cc_163 VPB N_A_306_74#_c_944_n 0.00711287f $X=-0.19 $Y=1.66 $X2=0.402 $Y2=1.845
cc_164 VPB N_A_306_74#_c_945_n 0.0192293f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.845
cc_165 VPB N_A_306_74#_c_946_n 0.0145254f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.845
cc_166 VPB N_A_306_74#_c_947_n 0.178904f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_167 VPB N_A_306_74#_M1022_g 0.0110598f $X=-0.19 $Y=1.66 $X2=0.32 $Y2=1.845
cc_168 VPB N_A_306_74#_c_931_n 0.0299618f $X=-0.19 $Y=1.66 $X2=0.32 $Y2=2.035
cc_169 VPB N_A_306_74#_c_932_n 0.012343f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_170 VPB N_A_306_74#_c_951_n 0.0089867f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_171 VPB N_A_306_74#_c_952_n 0.0254973f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_172 VPB N_A_306_74#_c_935_n 0.00363871f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_173 VPB N_A_306_74#_c_954_n 0.0069841f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_174 VPB N_A_1518_203#_c_1124_n 0.0069195f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=0.6
cc_175 VPB N_A_1518_203#_c_1125_n 0.0240163f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=0.6
cc_176 VPB N_A_1518_203#_c_1126_n 0.0216466f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_177 VPB N_A_1518_203#_c_1117_n 0.0041544f $X=-0.19 $Y=1.66 $X2=0.402
+ $Y2=1.165
cc_178 VPB N_A_1518_203#_c_1128_n 0.00705277f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_179 VPB N_A_1518_203#_c_1129_n 0.00198797f $X=-0.19 $Y=1.66 $X2=0.32
+ $Y2=1.295
cc_180 VPB N_A_1518_203#_c_1120_n 0.00168296f $X=-0.19 $Y=1.66 $X2=0.32
+ $Y2=1.665
cc_181 VPB N_A_1518_203#_c_1131_n 0.00942442f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_182 VPB N_A_1518_203#_c_1132_n 0.00312494f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_183 VPB N_A_1266_74#_c_1249_n 0.0330758f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.21
cc_184 VPB N_A_1266_74#_c_1250_n 0.0210347f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_185 VPB N_A_1266_74#_c_1236_n 0.00533618f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_186 VPB N_A_1266_74#_c_1237_n 0.003846f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_187 VPB N_A_1266_74#_c_1253_n 0.0108549f $X=-0.19 $Y=1.66 $X2=0.402 $Y2=1
cc_188 VPB N_A_1266_74#_c_1254_n 0.022831f $X=-0.19 $Y=1.66 $X2=0.402 $Y2=1.845
cc_189 VPB N_A_1266_74#_c_1242_n 9.60226e-19 $X=-0.19 $Y=1.66 $X2=0.32 $Y2=1.665
cc_190 VPB N_A_1266_74#_c_1256_n 0.00279628f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_191 VPB N_A_1266_74#_c_1257_n 0.00553847f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_192 VPB N_A_1266_74#_c_1245_n 0.00921317f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_193 VPB N_A_1266_74#_c_1247_n 2.00274e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_194 VPB N_A_1266_74#_c_1248_n 9.16426e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_195 VPB N_A_1864_409#_c_1401_n 0.0221503f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=2.75
cc_196 VPB N_A_1864_409#_c_1397_n 0.0304841f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.95
cc_197 VPB N_A_1864_409#_c_1398_n 0.00967318f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_198 VPB N_A_1864_409#_c_1404_n 0.00988755f $X=-0.19 $Y=1.66 $X2=0.402
+ $Y2=1.165
cc_199 VPB N_A_1864_409#_c_1400_n 0.00279207f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_200 VPB N_VPWR_c_1451_n 0.0103331f $X=-0.19 $Y=1.66 $X2=0.402 $Y2=2.01
cc_201 VPB N_VPWR_c_1452_n 0.0321941f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_202 VPB N_VPWR_c_1453_n 0.0127001f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_203 VPB N_VPWR_c_1454_n 0.00364482f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_204 VPB N_VPWR_c_1455_n 0.0150197f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_205 VPB N_VPWR_c_1456_n 0.0203282f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_206 VPB N_VPWR_c_1457_n 0.0249158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_207 VPB N_VPWR_c_1458_n 0.019026f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_208 VPB N_VPWR_c_1459_n 0.0204007f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_209 VPB N_VPWR_c_1460_n 0.0144553f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_210 VPB N_VPWR_c_1461_n 0.0120152f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_211 VPB N_VPWR_c_1462_n 0.0660664f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_212 VPB N_VPWR_c_1463_n 0.0205885f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_213 VPB N_VPWR_c_1464_n 0.0205285f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_214 VPB N_VPWR_c_1465_n 0.0598701f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_215 VPB N_VPWR_c_1466_n 0.0543442f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_216 VPB N_VPWR_c_1467_n 0.0380491f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_217 VPB N_VPWR_c_1468_n 0.0047828f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_218 VPB N_VPWR_c_1469_n 0.00613849f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_219 VPB N_VPWR_c_1470_n 0.00436844f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_220 VPB N_VPWR_c_1471_n 0.00436868f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_221 VPB N_VPWR_c_1472_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_222 VPB N_VPWR_c_1473_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_223 VPB N_VPWR_c_1450_n 0.115612f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_224 VPB N_A_30_78#_c_1591_n 0.00572962f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_225 VPB N_A_30_78#_c_1597_n 0.00384561f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.165
cc_226 VPB N_A_30_78#_c_1598_n 0.00755855f $X=-0.19 $Y=1.66 $X2=0.402 $Y2=2.01
cc_227 VPB N_A_30_78#_c_1593_n 0.00556354f $X=-0.19 $Y=1.66 $X2=0.32 $Y2=1.295
cc_228 VPB N_A_30_78#_c_1600_n 0.00883443f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_229 VPB N_A_30_78#_c_1601_n 0.0112127f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_230 VPB N_A_30_78#_c_1602_n 0.00239385f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_231 VPB N_A_30_78#_c_1603_n 0.00923877f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_232 VPB Q 0.0106664f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.95
cc_233 VPB Q 0.0225117f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_234 VPB N_Q_c_1717_n 0.00313086f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_235 N_D_M1025_g N_RESET_B_M1016_g 0.0243394f $X=0.51 $Y=0.6 $X2=0 $Y2=0
cc_236 N_D_c_239_n N_RESET_B_M1016_g 9.94104e-19 $X=0.385 $Y=1.165 $X2=0 $Y2=0
cc_237 N_D_c_236_n N_RESET_B_c_269_n 0.0243394f $X=0.402 $Y=1.828 $X2=0 $Y2=0
cc_238 N_D_c_241_n N_RESET_B_c_277_n 0.00650355f $X=0.495 $Y=2.375 $X2=0 $Y2=0
cc_239 N_D_c_242_n N_RESET_B_c_278_n 0.0156828f $X=0.495 $Y=2.465 $X2=0 $Y2=0
cc_240 N_D_c_238_n N_RESET_B_c_274_n 0.0243394f $X=0.385 $Y=1.165 $X2=0 $Y2=0
cc_241 N_D_c_244_n N_RESET_B_c_290_n 0.0243394f $X=0.385 $Y=1.845 $X2=0 $Y2=0
cc_242 N_D_c_242_n N_VPWR_c_1452_n 0.00729224f $X=0.495 $Y=2.465 $X2=0 $Y2=0
cc_243 N_D_c_239_n N_VPWR_c_1452_n 0.0129077f $X=0.385 $Y=1.165 $X2=0 $Y2=0
cc_244 N_D_c_244_n N_VPWR_c_1452_n 7.18884e-19 $X=0.385 $Y=1.845 $X2=0 $Y2=0
cc_245 N_D_c_242_n N_VPWR_c_1463_n 0.00444469f $X=0.495 $Y=2.465 $X2=0 $Y2=0
cc_246 N_D_c_242_n N_VPWR_c_1450_n 0.00895293f $X=0.495 $Y=2.465 $X2=0 $Y2=0
cc_247 N_D_M1025_g N_A_30_78#_c_1590_n 0.0108589f $X=0.51 $Y=0.6 $X2=0 $Y2=0
cc_248 N_D_c_239_n N_A_30_78#_c_1590_n 0.00411346f $X=0.385 $Y=1.165 $X2=0 $Y2=0
cc_249 N_D_M1025_g N_A_30_78#_c_1591_n 0.0145237f $X=0.51 $Y=0.6 $X2=0 $Y2=0
cc_250 N_D_c_239_n N_A_30_78#_c_1591_n 0.0884076f $X=0.385 $Y=1.165 $X2=0 $Y2=0
cc_251 N_D_M1025_g N_A_30_78#_c_1594_n 0.00806237f $X=0.51 $Y=0.6 $X2=0 $Y2=0
cc_252 N_D_c_238_n N_A_30_78#_c_1594_n 0.00161806f $X=0.385 $Y=1.165 $X2=0 $Y2=0
cc_253 N_D_c_239_n N_A_30_78#_c_1594_n 0.0286676f $X=0.385 $Y=1.165 $X2=0 $Y2=0
cc_254 N_D_c_241_n N_A_30_78#_c_1600_n 0.00464415f $X=0.495 $Y=2.375 $X2=0 $Y2=0
cc_255 N_D_c_242_n N_A_30_78#_c_1600_n 0.00887442f $X=0.495 $Y=2.465 $X2=0 $Y2=0
cc_256 N_D_M1025_g N_VGND_c_1751_n 0.00429844f $X=0.51 $Y=0.6 $X2=0 $Y2=0
cc_257 N_D_M1025_g N_VGND_c_1761_n 0.00539454f $X=0.51 $Y=0.6 $X2=0 $Y2=0
cc_258 N_RESET_B_c_274_n N_CLK_M1003_g 0.00301935f $X=1.155 $Y=1.295 $X2=0 $Y2=0
cc_259 N_RESET_B_c_269_n N_CLK_c_470_n 0.00635814f $X=1.072 $Y=1.893 $X2=0 $Y2=0
cc_260 N_RESET_B_c_283_n N_CLK_c_470_n 0.00427837f $X=4.895 $Y=2.035 $X2=0 $Y2=0
cc_261 N_RESET_B_c_274_n N_CLK_c_470_n 0.00730469f $X=1.155 $Y=1.295 $X2=0 $Y2=0
cc_262 N_RESET_B_c_283_n CLK 0.0140372f $X=4.895 $Y=2.035 $X2=0 $Y2=0
cc_263 N_RESET_B_c_283_n N_A_490_366#_M1008_d 0.00124406f $X=4.895 $Y=2.035
+ $X2=0 $Y2=0
cc_264 N_RESET_B_c_283_n N_A_490_366#_c_531_n 0.00357409f $X=4.895 $Y=2.035
+ $X2=0 $Y2=0
cc_265 N_RESET_B_c_283_n N_A_490_366#_c_512_n 0.0042766f $X=4.895 $Y=2.035 $X2=0
+ $Y2=0
cc_266 N_RESET_B_c_285_n N_A_490_366#_c_535_n 0.00268688f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_267 N_RESET_B_c_283_n N_A_490_366#_c_536_n 0.019565f $X=4.895 $Y=2.035 $X2=0
+ $Y2=0
cc_268 N_RESET_B_c_283_n N_A_490_366#_c_537_n 0.00843104f $X=4.895 $Y=2.035
+ $X2=0 $Y2=0
cc_269 N_RESET_B_c_283_n N_A_490_366#_c_520_n 0.0103491f $X=4.895 $Y=2.035 $X2=0
+ $Y2=0
cc_270 N_RESET_B_c_270_n N_A_490_366#_c_521_n 0.0109286f $X=4.785 $Y=1.185 $X2=0
+ $Y2=0
cc_271 N_RESET_B_c_285_n N_A_490_366#_c_524_n 0.0220527f $X=7.775 $Y=2.035 $X2=0
+ $Y2=0
cc_272 N_RESET_B_c_283_n N_A_490_366#_c_530_n 0.00382987f $X=4.895 $Y=2.035
+ $X2=0 $Y2=0
cc_273 N_RESET_B_c_285_n N_A_830_359#_M1017_d 0.00144653f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_274 N_RESET_B_c_279_n N_A_830_359#_c_717_n 0.0139713f $X=4.86 $Y=2.21 $X2=0
+ $Y2=0
cc_275 N_RESET_B_c_283_n N_A_830_359#_c_717_n 0.0113341f $X=4.895 $Y=2.035 $X2=0
+ $Y2=0
cc_276 N_RESET_B_c_291_n N_A_830_359#_c_717_n 0.0191507f $X=4.875 $Y=2.002 $X2=0
+ $Y2=0
cc_277 N_RESET_B_c_270_n N_A_830_359#_M1018_g 0.041724f $X=4.785 $Y=1.185 $X2=0
+ $Y2=0
cc_278 N_RESET_B_c_271_n N_A_830_359#_M1018_g 0.0138167f $X=4.875 $Y=1.795 $X2=0
+ $Y2=0
cc_279 N_RESET_B_c_270_n N_A_830_359#_c_714_n 0.00105936f $X=4.785 $Y=1.185
+ $X2=0 $Y2=0
cc_280 N_RESET_B_c_271_n N_A_830_359#_c_714_n 2.9783e-19 $X=4.875 $Y=1.795 $X2=0
+ $Y2=0
cc_281 N_RESET_B_c_283_n N_A_830_359#_c_714_n 0.0170583f $X=4.895 $Y=2.035 $X2=0
+ $Y2=0
cc_282 N_RESET_B_c_291_n N_A_830_359#_c_714_n 3.3918e-19 $X=4.875 $Y=2.002 $X2=0
+ $Y2=0
cc_283 N_RESET_B_c_270_n N_A_830_359#_c_732_n 0.0111445f $X=4.785 $Y=1.185 $X2=0
+ $Y2=0
cc_284 N_RESET_B_c_273_n N_A_830_359#_c_732_n 0.00240316f $X=4.875 $Y=1.26 $X2=0
+ $Y2=0
cc_285 N_RESET_B_c_285_n N_A_830_359#_c_720_n 0.0389295f $X=7.775 $Y=2.035 $X2=0
+ $Y2=0
cc_286 N_RESET_B_c_270_n N_A_695_457#_M1031_g 0.0148805f $X=4.785 $Y=1.185 $X2=0
+ $Y2=0
cc_287 N_RESET_B_c_273_n N_A_695_457#_M1031_g 0.00219471f $X=4.875 $Y=1.26 $X2=0
+ $Y2=0
cc_288 N_RESET_B_c_285_n N_A_695_457#_c_806_n 0.0113891f $X=7.775 $Y=2.035 $X2=0
+ $Y2=0
cc_289 N_RESET_B_c_283_n N_A_695_457#_c_800_n 0.0186344f $X=4.895 $Y=2.035 $X2=0
+ $Y2=0
cc_290 N_RESET_B_c_283_n N_A_695_457#_c_816_n 0.0138374f $X=4.895 $Y=2.035 $X2=0
+ $Y2=0
cc_291 N_RESET_B_c_283_n N_A_695_457#_c_808_n 0.008098f $X=4.895 $Y=2.035 $X2=0
+ $Y2=0
cc_292 N_RESET_B_c_279_n N_A_695_457#_c_801_n 0.00234023f $X=4.86 $Y=2.21 $X2=0
+ $Y2=0
cc_293 N_RESET_B_c_271_n N_A_695_457#_c_801_n 0.0056545f $X=4.875 $Y=1.795 $X2=0
+ $Y2=0
cc_294 N_RESET_B_c_283_n N_A_695_457#_c_801_n 0.0207498f $X=4.895 $Y=2.035 $X2=0
+ $Y2=0
cc_295 N_RESET_B_c_286_n N_A_695_457#_c_801_n 0.00237384f $X=5.185 $Y=2.035
+ $X2=0 $Y2=0
cc_296 N_RESET_B_c_287_n N_A_695_457#_c_801_n 0.0234789f $X=5.04 $Y=2.035 $X2=0
+ $Y2=0
cc_297 N_RESET_B_c_291_n N_A_695_457#_c_801_n 0.0103538f $X=4.875 $Y=2.002 $X2=0
+ $Y2=0
cc_298 N_RESET_B_c_273_n N_A_695_457#_c_802_n 0.00393752f $X=4.875 $Y=1.26 $X2=0
+ $Y2=0
cc_299 N_RESET_B_c_271_n N_A_695_457#_c_803_n 0.0121734f $X=4.875 $Y=1.795 $X2=0
+ $Y2=0
cc_300 N_RESET_B_c_273_n N_A_695_457#_c_803_n 0.00449896f $X=4.875 $Y=1.26 $X2=0
+ $Y2=0
cc_301 N_RESET_B_c_283_n N_A_695_457#_c_803_n 0.00353489f $X=4.895 $Y=2.035
+ $X2=0 $Y2=0
cc_302 N_RESET_B_c_285_n N_A_695_457#_c_803_n 0.0084128f $X=7.775 $Y=2.035 $X2=0
+ $Y2=0
cc_303 N_RESET_B_c_286_n N_A_695_457#_c_803_n 0.00351517f $X=5.185 $Y=2.035
+ $X2=0 $Y2=0
cc_304 N_RESET_B_c_287_n N_A_695_457#_c_803_n 0.01951f $X=5.04 $Y=2.035 $X2=0
+ $Y2=0
cc_305 N_RESET_B_c_291_n N_A_695_457#_c_803_n 0.00785354f $X=4.875 $Y=2.002
+ $X2=0 $Y2=0
cc_306 N_RESET_B_c_273_n N_A_695_457#_c_804_n 0.0103083f $X=4.875 $Y=1.26 $X2=0
+ $Y2=0
cc_307 N_RESET_B_c_285_n N_A_695_457#_c_804_n 0.00409962f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_308 N_RESET_B_c_279_n N_A_695_457#_c_811_n 0.00887731f $X=4.86 $Y=2.21 $X2=0
+ $Y2=0
cc_309 N_RESET_B_c_283_n N_A_695_457#_c_811_n 0.0041068f $X=4.895 $Y=2.035 $X2=0
+ $Y2=0
cc_310 N_RESET_B_c_285_n N_A_695_457#_c_811_n 4.57663e-19 $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_311 N_RESET_B_c_286_n N_A_695_457#_c_811_n 0.00893467f $X=5.185 $Y=2.035
+ $X2=0 $Y2=0
cc_312 N_RESET_B_c_287_n N_A_695_457#_c_811_n 0.0191542f $X=5.04 $Y=2.035 $X2=0
+ $Y2=0
cc_313 N_RESET_B_c_291_n N_A_695_457#_c_811_n 0.00191227f $X=4.875 $Y=2.002
+ $X2=0 $Y2=0
cc_314 N_RESET_B_c_279_n N_A_695_457#_c_840_n 0.00379552f $X=4.86 $Y=2.21 $X2=0
+ $Y2=0
cc_315 N_RESET_B_c_283_n N_A_306_74#_c_939_n 0.00909591f $X=4.895 $Y=2.035 $X2=0
+ $Y2=0
cc_316 N_RESET_B_c_283_n N_A_306_74#_c_927_n 0.00509095f $X=4.895 $Y=2.035 $X2=0
+ $Y2=0
cc_317 N_RESET_B_c_283_n N_A_306_74#_c_929_n 7.8631e-19 $X=4.895 $Y=2.035 $X2=0
+ $Y2=0
cc_318 N_RESET_B_c_283_n N_A_306_74#_c_946_n 0.00260456f $X=4.895 $Y=2.035 $X2=0
+ $Y2=0
cc_319 N_RESET_B_c_279_n N_A_306_74#_c_947_n 0.00852675f $X=4.86 $Y=2.21 $X2=0
+ $Y2=0
cc_320 N_RESET_B_c_285_n N_A_306_74#_M1022_g 0.00898574f $X=7.775 $Y=2.035 $X2=0
+ $Y2=0
cc_321 N_RESET_B_c_285_n N_A_306_74#_c_931_n 0.00802201f $X=7.775 $Y=2.035 $X2=0
+ $Y2=0
cc_322 N_RESET_B_c_285_n N_A_306_74#_c_932_n 3.42215e-19 $X=7.775 $Y=2.035 $X2=0
+ $Y2=0
cc_323 N_RESET_B_M1016_g N_A_306_74#_c_934_n 0.00308278f $X=0.9 $Y=0.6 $X2=0
+ $Y2=0
cc_324 N_RESET_B_c_283_n N_A_306_74#_c_935_n 8.85602e-19 $X=4.895 $Y=2.035 $X2=0
+ $Y2=0
cc_325 N_RESET_B_c_274_n N_A_306_74#_c_935_n 0.00644445f $X=1.155 $Y=1.295 $X2=0
+ $Y2=0
cc_326 N_RESET_B_c_275_n N_A_306_74#_c_935_n 0.049377f $X=1.155 $Y=1.295 $X2=0
+ $Y2=0
cc_327 N_RESET_B_c_283_n N_A_306_74#_c_937_n 0.00333482f $X=4.895 $Y=2.035 $X2=0
+ $Y2=0
cc_328 N_RESET_B_M1016_g N_A_306_74#_c_938_n 0.00279264f $X=0.9 $Y=0.6 $X2=0
+ $Y2=0
cc_329 N_RESET_B_c_275_n N_A_306_74#_c_938_n 8.29766e-19 $X=1.155 $Y=1.295 $X2=0
+ $Y2=0
cc_330 N_RESET_B_c_269_n N_A_306_74#_c_954_n 0.00298572f $X=1.072 $Y=1.893 $X2=0
+ $Y2=0
cc_331 N_RESET_B_c_283_n N_A_306_74#_c_954_n 0.0250468f $X=4.895 $Y=2.035 $X2=0
+ $Y2=0
cc_332 N_RESET_B_c_284_n N_A_306_74#_c_954_n 0.00246785f $X=1.345 $Y=2.035 $X2=0
+ $Y2=0
cc_333 N_RESET_B_c_275_n N_A_306_74#_c_954_n 0.0236266f $X=1.155 $Y=1.295 $X2=0
+ $Y2=0
cc_334 N_RESET_B_M1002_g N_A_1518_203#_c_1124_n 0.00652196f $X=8.205 $Y=0.615
+ $X2=0 $Y2=0
cc_335 N_RESET_B_c_282_n N_A_1518_203#_c_1125_n 0.022618f $X=8.26 $Y=2.39 $X2=0
+ $Y2=0
cc_336 N_RESET_B_c_285_n N_A_1518_203#_c_1125_n 0.00706641f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_337 N_RESET_B_c_288_n N_A_1518_203#_c_1125_n 0.00231702f $X=7.92 $Y=2.035
+ $X2=0 $Y2=0
cc_338 N_RESET_B_c_292_n N_A_1518_203#_c_1125_n 0.00228452f $X=8.18 $Y=2.09
+ $X2=0 $Y2=0
cc_339 N_RESET_B_c_282_n N_A_1518_203#_c_1126_n 0.012219f $X=8.26 $Y=2.39 $X2=0
+ $Y2=0
cc_340 N_RESET_B_M1002_g N_A_1518_203#_M1019_g 0.0166359f $X=8.205 $Y=0.615
+ $X2=0 $Y2=0
cc_341 N_RESET_B_M1002_g N_A_1518_203#_c_1117_n 0.0133984f $X=8.205 $Y=0.615
+ $X2=0 $Y2=0
cc_342 N_RESET_B_M1002_g N_A_1518_203#_c_1118_n 0.0149634f $X=8.205 $Y=0.615
+ $X2=0 $Y2=0
cc_343 N_RESET_B_M1002_g N_A_1518_203#_c_1119_n 0.00216035f $X=8.205 $Y=0.615
+ $X2=0 $Y2=0
cc_344 N_RESET_B_M1002_g N_A_1518_203#_c_1129_n 0.00169886f $X=8.205 $Y=0.615
+ $X2=0 $Y2=0
cc_345 N_RESET_B_c_282_n N_A_1518_203#_c_1129_n 6.9451e-19 $X=8.26 $Y=2.39 $X2=0
+ $Y2=0
cc_346 N_RESET_B_c_288_n N_A_1518_203#_c_1129_n 4.76192e-19 $X=7.92 $Y=2.035
+ $X2=0 $Y2=0
cc_347 N_RESET_B_c_292_n N_A_1518_203#_c_1129_n 0.00873148f $X=8.18 $Y=2.09
+ $X2=0 $Y2=0
cc_348 N_RESET_B_M1002_g N_A_1518_203#_c_1121_n 0.00118187f $X=8.205 $Y=0.615
+ $X2=0 $Y2=0
cc_349 N_RESET_B_c_285_n N_A_1518_203#_c_1121_n 3.17521e-19 $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_350 N_RESET_B_M1002_g N_A_1518_203#_c_1122_n 0.021263f $X=8.205 $Y=0.615
+ $X2=0 $Y2=0
cc_351 N_RESET_B_c_282_n N_A_1518_203#_c_1131_n 0.00637785f $X=8.26 $Y=2.39
+ $X2=0 $Y2=0
cc_352 N_RESET_B_c_292_n N_A_1518_203#_c_1131_n 0.00174345f $X=8.18 $Y=2.09
+ $X2=0 $Y2=0
cc_353 N_RESET_B_c_282_n N_A_1518_203#_c_1132_n 0.00534913f $X=8.26 $Y=2.39
+ $X2=0 $Y2=0
cc_354 N_RESET_B_c_288_n N_A_1518_203#_c_1132_n 5.01506e-19 $X=7.92 $Y=2.035
+ $X2=0 $Y2=0
cc_355 N_RESET_B_c_292_n N_A_1518_203#_c_1132_n 0.0175397f $X=8.18 $Y=2.09 $X2=0
+ $Y2=0
cc_356 N_RESET_B_c_285_n N_A_1266_74#_M1022_d 0.00283611f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_357 N_RESET_B_M1002_g N_A_1266_74#_M1021_g 0.0757442f $X=8.205 $Y=0.615 $X2=0
+ $Y2=0
cc_358 N_RESET_B_M1002_g N_A_1266_74#_c_1249_n 0.00953304f $X=8.205 $Y=0.615
+ $X2=0 $Y2=0
cc_359 N_RESET_B_c_282_n N_A_1266_74#_c_1249_n 0.0206573f $X=8.26 $Y=2.39 $X2=0
+ $Y2=0
cc_360 N_RESET_B_c_292_n N_A_1266_74#_c_1249_n 3.48207e-19 $X=8.18 $Y=2.09 $X2=0
+ $Y2=0
cc_361 N_RESET_B_c_282_n N_A_1266_74#_c_1250_n 0.00915627f $X=8.26 $Y=2.39 $X2=0
+ $Y2=0
cc_362 N_RESET_B_M1002_g N_A_1266_74#_c_1237_n 0.00996674f $X=8.205 $Y=0.615
+ $X2=0 $Y2=0
cc_363 N_RESET_B_c_285_n N_A_1266_74#_c_1256_n 0.0174694f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_364 N_RESET_B_c_285_n N_A_1266_74#_c_1269_n 0.0206747f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_365 N_RESET_B_M1002_g N_A_1266_74#_c_1257_n 0.00109662f $X=8.205 $Y=0.615
+ $X2=0 $Y2=0
cc_366 N_RESET_B_c_282_n N_A_1266_74#_c_1257_n 0.00116333f $X=8.26 $Y=2.39 $X2=0
+ $Y2=0
cc_367 N_RESET_B_c_285_n N_A_1266_74#_c_1257_n 0.0211228f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_368 N_RESET_B_c_288_n N_A_1266_74#_c_1257_n 0.00228452f $X=7.92 $Y=2.035
+ $X2=0 $Y2=0
cc_369 N_RESET_B_c_292_n N_A_1266_74#_c_1257_n 0.0236542f $X=8.18 $Y=2.09 $X2=0
+ $Y2=0
cc_370 N_RESET_B_M1002_g N_A_1266_74#_c_1245_n 0.011972f $X=8.205 $Y=0.615 $X2=0
+ $Y2=0
cc_371 N_RESET_B_c_282_n N_A_1266_74#_c_1245_n 0.00135016f $X=8.26 $Y=2.39 $X2=0
+ $Y2=0
cc_372 N_RESET_B_c_285_n N_A_1266_74#_c_1245_n 0.00476106f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_373 N_RESET_B_c_288_n N_A_1266_74#_c_1245_n 0.00823149f $X=7.92 $Y=2.035
+ $X2=0 $Y2=0
cc_374 N_RESET_B_c_292_n N_A_1266_74#_c_1245_n 0.02904f $X=8.18 $Y=2.09 $X2=0
+ $Y2=0
cc_375 N_RESET_B_c_285_n N_A_1266_74#_c_1247_n 0.00599756f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_376 N_RESET_B_M1002_g N_A_1266_74#_c_1248_n 0.00110907f $X=8.205 $Y=0.615
+ $X2=0 $Y2=0
cc_377 N_RESET_B_c_283_n N_VPWR_M1005_d 0.00544297f $X=4.895 $Y=2.035 $X2=0
+ $Y2=0
cc_378 N_RESET_B_c_278_n N_VPWR_c_1453_n 0.00589882f $X=0.945 $Y=2.465 $X2=0
+ $Y2=0
cc_379 N_RESET_B_c_279_n N_VPWR_c_1455_n 0.00274139f $X=4.86 $Y=2.21 $X2=0 $Y2=0
cc_380 N_RESET_B_c_279_n N_VPWR_c_1457_n 0.0078214f $X=4.86 $Y=2.21 $X2=0 $Y2=0
cc_381 N_RESET_B_c_271_n N_VPWR_c_1457_n 0.00126145f $X=4.875 $Y=1.795 $X2=0
+ $Y2=0
cc_382 N_RESET_B_c_285_n N_VPWR_c_1457_n 0.0317336f $X=7.775 $Y=2.035 $X2=0
+ $Y2=0
cc_383 N_RESET_B_c_286_n N_VPWR_c_1457_n 5.51604e-19 $X=5.185 $Y=2.035 $X2=0
+ $Y2=0
cc_384 N_RESET_B_c_287_n N_VPWR_c_1457_n 0.023147f $X=5.04 $Y=2.035 $X2=0 $Y2=0
cc_385 N_RESET_B_c_291_n N_VPWR_c_1457_n 0.00289108f $X=4.875 $Y=2.002 $X2=0
+ $Y2=0
cc_386 N_RESET_B_c_282_n N_VPWR_c_1458_n 0.00888753f $X=8.26 $Y=2.39 $X2=0 $Y2=0
cc_387 N_RESET_B_c_288_n N_VPWR_c_1458_n 0.00171912f $X=7.92 $Y=2.035 $X2=0
+ $Y2=0
cc_388 N_RESET_B_c_292_n N_VPWR_c_1458_n 0.0244512f $X=8.18 $Y=2.09 $X2=0 $Y2=0
cc_389 N_RESET_B_c_282_n N_VPWR_c_1459_n 0.00510653f $X=8.26 $Y=2.39 $X2=0 $Y2=0
cc_390 N_RESET_B_c_278_n N_VPWR_c_1463_n 0.00444469f $X=0.945 $Y=2.465 $X2=0
+ $Y2=0
cc_391 N_RESET_B_c_278_n N_VPWR_c_1450_n 0.0046079f $X=0.945 $Y=2.465 $X2=0
+ $Y2=0
cc_392 N_RESET_B_c_279_n N_VPWR_c_1450_n 9.49986e-19 $X=4.86 $Y=2.21 $X2=0 $Y2=0
cc_393 N_RESET_B_c_282_n N_VPWR_c_1450_n 0.0052212f $X=8.26 $Y=2.39 $X2=0 $Y2=0
cc_394 N_RESET_B_M1016_g N_A_30_78#_c_1590_n 0.00429043f $X=0.9 $Y=0.6 $X2=0
+ $Y2=0
cc_395 N_RESET_B_M1016_g N_A_30_78#_c_1591_n 0.00821385f $X=0.9 $Y=0.6 $X2=0
+ $Y2=0
cc_396 N_RESET_B_c_269_n N_A_30_78#_c_1591_n 0.0115982f $X=1.072 $Y=1.893 $X2=0
+ $Y2=0
cc_397 N_RESET_B_c_277_n N_A_30_78#_c_1591_n 0.00433638f $X=0.945 $Y=2.375 $X2=0
+ $Y2=0
cc_398 N_RESET_B_c_284_n N_A_30_78#_c_1591_n 0.00186952f $X=1.345 $Y=2.035 $X2=0
+ $Y2=0
cc_399 N_RESET_B_c_274_n N_A_30_78#_c_1591_n 0.00558005f $X=1.155 $Y=1.295 $X2=0
+ $Y2=0
cc_400 N_RESET_B_c_275_n N_A_30_78#_c_1591_n 0.069302f $X=1.155 $Y=1.295 $X2=0
+ $Y2=0
cc_401 N_RESET_B_c_290_n N_A_30_78#_c_1591_n 0.00619346f $X=1.155 $Y=1.975 $X2=0
+ $Y2=0
cc_402 N_RESET_B_c_283_n N_A_30_78#_c_1597_n 0.0311901f $X=4.895 $Y=2.035 $X2=0
+ $Y2=0
cc_403 N_RESET_B_c_283_n N_A_30_78#_c_1598_n 0.018683f $X=4.895 $Y=2.035 $X2=0
+ $Y2=0
cc_404 N_RESET_B_c_283_n N_A_30_78#_c_1593_n 0.00949005f $X=4.895 $Y=2.035 $X2=0
+ $Y2=0
cc_405 N_RESET_B_M1016_g N_A_30_78#_c_1594_n 9.29579e-19 $X=0.9 $Y=0.6 $X2=0
+ $Y2=0
cc_406 N_RESET_B_c_277_n N_A_30_78#_c_1600_n 0.00222596f $X=0.945 $Y=2.375 $X2=0
+ $Y2=0
cc_407 N_RESET_B_c_278_n N_A_30_78#_c_1600_n 0.0129415f $X=0.945 $Y=2.465 $X2=0
+ $Y2=0
cc_408 N_RESET_B_c_277_n N_A_30_78#_c_1601_n 0.0087036f $X=0.945 $Y=2.375 $X2=0
+ $Y2=0
cc_409 N_RESET_B_c_278_n N_A_30_78#_c_1601_n 0.00725597f $X=0.945 $Y=2.465 $X2=0
+ $Y2=0
cc_410 N_RESET_B_c_283_n N_A_30_78#_c_1601_n 0.00637217f $X=4.895 $Y=2.035 $X2=0
+ $Y2=0
cc_411 N_RESET_B_c_284_n N_A_30_78#_c_1601_n 0.00929883f $X=1.345 $Y=2.035 $X2=0
+ $Y2=0
cc_412 N_RESET_B_c_275_n N_A_30_78#_c_1601_n 0.0168504f $X=1.155 $Y=1.295 $X2=0
+ $Y2=0
cc_413 N_RESET_B_c_290_n N_A_30_78#_c_1601_n 0.00294352f $X=1.155 $Y=1.975 $X2=0
+ $Y2=0
cc_414 N_RESET_B_c_278_n N_A_30_78#_c_1602_n 5.09312e-19 $X=0.945 $Y=2.465 $X2=0
+ $Y2=0
cc_415 N_RESET_B_c_283_n N_A_30_78#_c_1603_n 0.0162799f $X=4.895 $Y=2.035 $X2=0
+ $Y2=0
cc_416 N_RESET_B_c_283_n N_A_30_78#_c_1595_n 0.00385939f $X=4.895 $Y=2.035 $X2=0
+ $Y2=0
cc_417 N_RESET_B_M1016_g N_VGND_c_1745_n 0.00603227f $X=0.9 $Y=0.6 $X2=0 $Y2=0
cc_418 N_RESET_B_c_274_n N_VGND_c_1745_n 0.00181416f $X=1.155 $Y=1.295 $X2=0
+ $Y2=0
cc_419 N_RESET_B_c_275_n N_VGND_c_1745_n 0.0144384f $X=1.155 $Y=1.295 $X2=0
+ $Y2=0
cc_420 N_RESET_B_M1002_g N_VGND_c_1747_n 0.0058325f $X=8.205 $Y=0.615 $X2=0
+ $Y2=0
cc_421 N_RESET_B_M1016_g N_VGND_c_1751_n 0.0053757f $X=0.9 $Y=0.6 $X2=0 $Y2=0
cc_422 N_RESET_B_c_270_n N_VGND_c_1754_n 0.00293358f $X=4.785 $Y=1.185 $X2=0
+ $Y2=0
cc_423 N_RESET_B_M1002_g N_VGND_c_1756_n 0.00552345f $X=8.205 $Y=0.615 $X2=0
+ $Y2=0
cc_424 N_RESET_B_M1016_g N_VGND_c_1761_n 0.00539454f $X=0.9 $Y=0.6 $X2=0 $Y2=0
cc_425 N_RESET_B_c_270_n N_VGND_c_1761_n 0.00451834f $X=4.785 $Y=1.185 $X2=0
+ $Y2=0
cc_426 N_RESET_B_M1002_g N_VGND_c_1761_n 0.00534666f $X=8.205 $Y=0.615 $X2=0
+ $Y2=0
cc_427 CLK N_A_490_366#_c_518_n 2.80033e-19 $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_428 CLK N_A_490_366#_c_537_n 0.0091781f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_429 N_CLK_c_470_n N_A_306_74#_c_939_n 0.0412532f $X=1.925 $Y=1.755 $X2=0
+ $Y2=0
cc_430 CLK N_A_306_74#_c_939_n 2.22405e-19 $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_431 N_CLK_M1003_g N_A_306_74#_c_926_n 0.023755f $X=1.89 $Y=0.74 $X2=0 $Y2=0
cc_432 N_CLK_M1003_g N_A_306_74#_c_929_n 0.00456314f $X=1.89 $Y=0.74 $X2=0 $Y2=0
cc_433 N_CLK_c_470_n N_A_306_74#_c_929_n 0.0252834f $X=1.925 $Y=1.755 $X2=0
+ $Y2=0
cc_434 CLK N_A_306_74#_c_929_n 0.00493727f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_435 N_CLK_M1003_g N_A_306_74#_c_934_n 0.00981385f $X=1.89 $Y=0.74 $X2=0 $Y2=0
cc_436 N_CLK_M1003_g N_A_306_74#_c_935_n 0.00375487f $X=1.89 $Y=0.74 $X2=0 $Y2=0
cc_437 N_CLK_c_470_n N_A_306_74#_c_935_n 0.00491363f $X=1.925 $Y=1.755 $X2=0
+ $Y2=0
cc_438 CLK N_A_306_74#_c_935_n 0.0314125f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_439 N_CLK_M1003_g N_A_306_74#_c_936_n 0.0114775f $X=1.89 $Y=0.74 $X2=0 $Y2=0
cc_440 N_CLK_c_470_n N_A_306_74#_c_936_n 7.71603e-19 $X=1.925 $Y=1.755 $X2=0
+ $Y2=0
cc_441 CLK N_A_306_74#_c_936_n 0.0336979f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_442 N_CLK_M1003_g N_A_306_74#_c_937_n 7.72463e-19 $X=1.89 $Y=0.74 $X2=0 $Y2=0
cc_443 CLK N_A_306_74#_c_937_n 0.0192888f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_444 N_CLK_M1003_g N_A_306_74#_c_938_n 0.00130048f $X=1.89 $Y=0.74 $X2=0 $Y2=0
cc_445 N_CLK_c_470_n N_A_306_74#_c_938_n 0.00166711f $X=1.925 $Y=1.755 $X2=0
+ $Y2=0
cc_446 CLK N_A_306_74#_c_938_n 0.00370093f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_447 N_CLK_c_470_n N_A_306_74#_c_954_n 0.00839664f $X=1.925 $Y=1.755 $X2=0
+ $Y2=0
cc_448 CLK N_A_306_74#_c_954_n 0.00517175f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_449 N_CLK_c_470_n N_VPWR_c_1453_n 0.00714164f $X=1.925 $Y=1.755 $X2=0 $Y2=0
cc_450 N_CLK_c_470_n N_VPWR_c_1454_n 0.0105821f $X=1.925 $Y=1.755 $X2=0 $Y2=0
cc_451 N_CLK_c_470_n N_VPWR_c_1464_n 0.00512473f $X=1.925 $Y=1.755 $X2=0 $Y2=0
cc_452 N_CLK_c_470_n N_VPWR_c_1450_n 0.00492022f $X=1.925 $Y=1.755 $X2=0 $Y2=0
cc_453 N_CLK_c_470_n N_A_30_78#_c_1597_n 0.0141336f $X=1.925 $Y=1.755 $X2=0
+ $Y2=0
cc_454 CLK N_A_30_78#_c_1597_n 0.00297855f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_455 N_CLK_c_470_n N_A_30_78#_c_1602_n 0.00118571f $X=1.925 $Y=1.755 $X2=0
+ $Y2=0
cc_456 N_CLK_M1003_g N_VGND_c_1745_n 0.00342433f $X=1.89 $Y=0.74 $X2=0 $Y2=0
cc_457 N_CLK_M1003_g N_VGND_c_1746_n 0.00550183f $X=1.89 $Y=0.74 $X2=0 $Y2=0
cc_458 N_CLK_M1003_g N_VGND_c_1753_n 0.00434272f $X=1.89 $Y=0.74 $X2=0 $Y2=0
cc_459 N_CLK_M1003_g N_VGND_c_1761_n 0.00825771f $X=1.89 $Y=0.74 $X2=0 $Y2=0
cc_460 N_A_490_366#_c_521_n N_A_830_359#_M1031_d 0.00330812f $X=5.48 $Y=0.65
+ $X2=-0.19 $Y2=-0.245
cc_461 N_A_490_366#_c_554_p N_A_830_359#_M1031_d 0.00218198f $X=5.565 $Y=0.565
+ $X2=-0.19 $Y2=-0.245
cc_462 N_A_490_366#_c_522_n N_A_830_359#_M1031_d 0.00764003f $X=7.25 $Y=0.34
+ $X2=-0.19 $Y2=-0.245
cc_463 N_A_490_366#_c_531_n N_A_830_359#_c_717_n 0.00346941f $X=3.4 $Y=2.12
+ $X2=0 $Y2=0
cc_464 N_A_490_366#_c_530_n N_A_830_359#_c_717_n 9.8574e-19 $X=3.33 $Y=1.635
+ $X2=0 $Y2=0
cc_465 N_A_490_366#_c_513_n N_A_830_359#_M1018_g 0.00466149f $X=4.005 $Y=1.405
+ $X2=0 $Y2=0
cc_466 N_A_490_366#_M1001_g N_A_830_359#_M1018_g 0.0529943f $X=4.005 $Y=0.9
+ $X2=0 $Y2=0
cc_467 N_A_490_366#_c_521_n N_A_830_359#_M1018_g 0.00367082f $X=5.48 $Y=0.65
+ $X2=0 $Y2=0
cc_468 N_A_490_366#_c_527_n N_A_830_359#_M1018_g 0.00687536f $X=4.35 $Y=0.415
+ $X2=0 $Y2=0
cc_469 N_A_490_366#_c_513_n N_A_830_359#_c_714_n 3.67416e-19 $X=4.005 $Y=1.405
+ $X2=0 $Y2=0
cc_470 N_A_490_366#_M1001_g N_A_830_359#_c_714_n 0.00134011f $X=4.005 $Y=0.9
+ $X2=0 $Y2=0
cc_471 N_A_490_366#_c_521_n N_A_830_359#_c_732_n 0.0658997f $X=5.48 $Y=0.65
+ $X2=0 $Y2=0
cc_472 N_A_490_366#_c_522_n N_A_830_359#_c_732_n 0.00571426f $X=7.25 $Y=0.34
+ $X2=0 $Y2=0
cc_473 N_A_490_366#_c_521_n N_A_830_359#_c_748_n 7.61753e-19 $X=5.48 $Y=0.65
+ $X2=0 $Y2=0
cc_474 N_A_490_366#_c_527_n N_A_830_359#_c_748_n 0.00928432f $X=4.35 $Y=0.415
+ $X2=0 $Y2=0
cc_475 N_A_490_366#_c_517_n N_A_830_359#_c_720_n 0.00388841f $X=6.33 $Y=1.27
+ $X2=0 $Y2=0
cc_476 N_A_490_366#_c_515_n N_A_830_359#_c_715_n 0.00184952f $X=6.255 $Y=1.195
+ $X2=0 $Y2=0
cc_477 N_A_490_366#_c_521_n N_A_830_359#_c_715_n 0.00596144f $X=5.48 $Y=0.65
+ $X2=0 $Y2=0
cc_478 N_A_490_366#_c_522_n N_A_830_359#_c_715_n 0.0168368f $X=7.25 $Y=0.34
+ $X2=0 $Y2=0
cc_479 N_A_490_366#_c_517_n N_A_830_359#_c_716_n 0.00184952f $X=6.33 $Y=1.27
+ $X2=0 $Y2=0
cc_480 N_A_490_366#_c_515_n N_A_695_457#_M1031_g 0.00895705f $X=6.255 $Y=1.195
+ $X2=0 $Y2=0
cc_481 N_A_490_366#_c_521_n N_A_695_457#_M1031_g 0.0118282f $X=5.48 $Y=0.65
+ $X2=0 $Y2=0
cc_482 N_A_490_366#_c_554_p N_A_695_457#_M1031_g 0.00736306f $X=5.565 $Y=0.565
+ $X2=0 $Y2=0
cc_483 N_A_490_366#_c_523_n N_A_695_457#_M1031_g 0.00665672f $X=5.65 $Y=0.34
+ $X2=0 $Y2=0
cc_484 N_A_490_366#_c_531_n N_A_695_457#_c_800_n 3.96425e-19 $X=3.4 $Y=2.12
+ $X2=0 $Y2=0
cc_485 N_A_490_366#_c_513_n N_A_695_457#_c_800_n 0.0113903f $X=4.005 $Y=1.405
+ $X2=0 $Y2=0
cc_486 N_A_490_366#_M1001_g N_A_695_457#_c_800_n 0.00880363f $X=4.005 $Y=0.9
+ $X2=0 $Y2=0
cc_487 N_A_490_366#_c_532_n N_A_695_457#_c_808_n 0.00398891f $X=3.4 $Y=2.21
+ $X2=0 $Y2=0
cc_488 N_A_490_366#_c_512_n N_A_695_457#_c_808_n 0.00109304f $X=3.79 $Y=1.635
+ $X2=0 $Y2=0
cc_489 N_A_490_366#_c_517_n N_A_695_457#_c_804_n 0.00170129f $X=6.33 $Y=1.27
+ $X2=0 $Y2=0
cc_490 N_A_490_366#_c_512_n N_A_695_457#_c_805_n 9.27017e-19 $X=3.79 $Y=1.635
+ $X2=0 $Y2=0
cc_491 N_A_490_366#_c_513_n N_A_695_457#_c_805_n 0.00364191f $X=4.005 $Y=1.405
+ $X2=0 $Y2=0
cc_492 N_A_490_366#_M1001_g N_A_695_457#_c_805_n 0.00809644f $X=4.005 $Y=0.9
+ $X2=0 $Y2=0
cc_493 N_A_490_366#_c_519_n N_A_695_457#_c_805_n 0.0352685f $X=4.265 $Y=0.415
+ $X2=0 $Y2=0
cc_494 N_A_490_366#_c_527_n N_A_695_457#_c_805_n 0.00147443f $X=4.35 $Y=0.415
+ $X2=0 $Y2=0
cc_495 N_A_490_366#_c_537_n N_A_306_74#_c_939_n 0.0022767f $X=3.035 $Y=1.725
+ $X2=0 $Y2=0
cc_496 N_A_490_366#_c_518_n N_A_306_74#_c_926_n 0.00552525f $X=2.95 $Y=1.56
+ $X2=0 $Y2=0
cc_497 N_A_490_366#_c_526_n N_A_306_74#_c_926_n 0.009246f $X=2.772 $Y=0.415
+ $X2=0 $Y2=0
cc_498 N_A_490_366#_c_531_n N_A_306_74#_c_927_n 0.0107254f $X=3.4 $Y=2.12 $X2=0
+ $Y2=0
cc_499 N_A_490_366#_c_532_n N_A_306_74#_c_927_n 0.0124685f $X=3.4 $Y=2.21 $X2=0
+ $Y2=0
cc_500 N_A_490_366#_c_536_n N_A_306_74#_c_927_n 0.00516557f $X=2.6 $Y=1.99 $X2=0
+ $Y2=0
cc_501 N_A_490_366#_c_518_n N_A_306_74#_c_927_n 3.10799e-19 $X=2.95 $Y=1.56
+ $X2=0 $Y2=0
cc_502 N_A_490_366#_c_537_n N_A_306_74#_c_927_n 0.0168163f $X=3.035 $Y=1.725
+ $X2=0 $Y2=0
cc_503 N_A_490_366#_c_530_n N_A_306_74#_c_927_n 0.021379f $X=3.33 $Y=1.635 $X2=0
+ $Y2=0
cc_504 N_A_490_366#_c_518_n N_A_306_74#_c_928_n 0.00679735f $X=2.95 $Y=1.56
+ $X2=0 $Y2=0
cc_505 N_A_490_366#_c_520_n N_A_306_74#_c_928_n 0.00510949f $X=3.33 $Y=1.725
+ $X2=0 $Y2=0
cc_506 N_A_490_366#_c_530_n N_A_306_74#_c_928_n 0.0263533f $X=3.33 $Y=1.635
+ $X2=0 $Y2=0
cc_507 N_A_490_366#_c_518_n N_A_306_74#_c_929_n 0.0117273f $X=2.95 $Y=1.56 $X2=0
+ $Y2=0
cc_508 N_A_490_366#_c_537_n N_A_306_74#_c_929_n 0.00288476f $X=3.035 $Y=1.725
+ $X2=0 $Y2=0
cc_509 N_A_490_366#_c_526_n N_A_306_74#_c_929_n 0.00673784f $X=2.772 $Y=0.415
+ $X2=0 $Y2=0
cc_510 N_A_490_366#_c_532_n N_A_306_74#_c_942_n 0.00899632f $X=3.4 $Y=2.21 $X2=0
+ $Y2=0
cc_511 N_A_490_366#_M1001_g N_A_306_74#_c_930_n 0.0189665f $X=4.005 $Y=0.9 $X2=0
+ $Y2=0
cc_512 N_A_490_366#_c_519_n N_A_306_74#_c_930_n 0.00661564f $X=4.265 $Y=0.415
+ $X2=0 $Y2=0
cc_513 N_A_490_366#_c_526_n N_A_306_74#_c_930_n 0.00461825f $X=2.772 $Y=0.415
+ $X2=0 $Y2=0
cc_514 N_A_490_366#_c_532_n N_A_306_74#_c_944_n 0.00278823f $X=3.4 $Y=2.21 $X2=0
+ $Y2=0
cc_515 N_A_490_366#_c_532_n N_A_306_74#_c_946_n 0.00991521f $X=3.4 $Y=2.21 $X2=0
+ $Y2=0
cc_516 N_A_490_366#_c_512_n N_A_306_74#_c_946_n 0.00449188f $X=3.79 $Y=1.635
+ $X2=0 $Y2=0
cc_517 N_A_490_366#_c_535_n N_A_306_74#_M1022_g 0.00735807f $X=7.265 $Y=2.39
+ $X2=0 $Y2=0
cc_518 N_A_490_366#_c_516_n N_A_306_74#_c_931_n 0.0196234f $X=6.69 $Y=1.27 $X2=0
+ $Y2=0
cc_519 N_A_490_366#_c_535_n N_A_306_74#_c_931_n 0.0220783f $X=7.265 $Y=2.39
+ $X2=0 $Y2=0
cc_520 N_A_490_366#_c_524_n N_A_306_74#_c_931_n 0.0164562f $X=7.13 $Y=2.14 $X2=0
+ $Y2=0
cc_521 N_A_490_366#_c_529_n N_A_306_74#_c_931_n 0.00266664f $X=7.335 $Y=1.18
+ $X2=0 $Y2=0
cc_522 N_A_490_366#_c_517_n N_A_306_74#_c_932_n 0.0196234f $X=6.33 $Y=1.27 $X2=0
+ $Y2=0
cc_523 N_A_490_366#_c_522_n N_A_306_74#_M1020_g 0.0088085f $X=7.25 $Y=0.34 $X2=0
+ $Y2=0
cc_524 N_A_490_366#_c_524_n N_A_306_74#_M1020_g 0.00923892f $X=7.13 $Y=2.14
+ $X2=0 $Y2=0
cc_525 N_A_490_366#_c_525_n N_A_306_74#_M1020_g 0.0233298f $X=7.335 $Y=1.015
+ $X2=0 $Y2=0
cc_526 N_A_490_366#_c_528_n N_A_306_74#_M1020_g 0.0213806f $X=6.855 $Y=1.18
+ $X2=0 $Y2=0
cc_527 N_A_490_366#_c_529_n N_A_306_74#_M1020_g 0.011895f $X=7.335 $Y=1.18 $X2=0
+ $Y2=0
cc_528 N_A_490_366#_c_535_n N_A_306_74#_c_952_n 0.00118457f $X=7.265 $Y=2.39
+ $X2=0 $Y2=0
cc_529 N_A_490_366#_M1030_d N_A_306_74#_c_936_n 0.00358564f $X=2.465 $Y=0.37
+ $X2=0 $Y2=0
cc_530 N_A_490_366#_c_518_n N_A_306_74#_c_936_n 0.01411f $X=2.95 $Y=1.56 $X2=0
+ $Y2=0
cc_531 N_A_490_366#_c_526_n N_A_306_74#_c_936_n 0.0150014f $X=2.772 $Y=0.415
+ $X2=0 $Y2=0
cc_532 N_A_490_366#_c_518_n N_A_306_74#_c_937_n 0.0290616f $X=2.95 $Y=1.56 $X2=0
+ $Y2=0
cc_533 N_A_490_366#_c_537_n N_A_306_74#_c_937_n 0.014588f $X=3.035 $Y=1.725
+ $X2=0 $Y2=0
cc_534 N_A_490_366#_c_536_n N_A_306_74#_c_954_n 0.00440098f $X=2.6 $Y=1.99 $X2=0
+ $Y2=0
cc_535 N_A_490_366#_c_537_n N_A_306_74#_c_954_n 0.00231522f $X=3.035 $Y=1.725
+ $X2=0 $Y2=0
cc_536 N_A_490_366#_c_535_n N_A_1518_203#_c_1125_n 0.0222944f $X=7.265 $Y=2.39
+ $X2=0 $Y2=0
cc_537 N_A_490_366#_c_524_n N_A_1518_203#_c_1125_n 3.6309e-19 $X=7.13 $Y=2.14
+ $X2=0 $Y2=0
cc_538 N_A_490_366#_c_535_n N_A_1518_203#_c_1126_n 0.029186f $X=7.265 $Y=2.39
+ $X2=0 $Y2=0
cc_539 N_A_490_366#_c_522_n N_A_1518_203#_M1019_g 0.00107872f $X=7.25 $Y=0.34
+ $X2=0 $Y2=0
cc_540 N_A_490_366#_c_525_n N_A_1518_203#_M1019_g 0.0045389f $X=7.335 $Y=1.015
+ $X2=0 $Y2=0
cc_541 N_A_490_366#_c_524_n N_A_1518_203#_c_1117_n 0.00240511f $X=7.13 $Y=2.14
+ $X2=0 $Y2=0
cc_542 N_A_490_366#_c_529_n N_A_1518_203#_c_1121_n 0.0276613f $X=7.335 $Y=1.18
+ $X2=0 $Y2=0
cc_543 N_A_490_366#_c_529_n N_A_1518_203#_c_1122_n 0.00201148f $X=7.335 $Y=1.18
+ $X2=0 $Y2=0
cc_544 N_A_490_366#_c_522_n N_A_1266_74#_M1026_d 0.00949775f $X=7.25 $Y=0.34
+ $X2=-0.19 $Y2=-0.245
cc_545 N_A_490_366#_c_515_n N_A_1266_74#_c_1283_n 0.0033591f $X=6.255 $Y=1.195
+ $X2=0 $Y2=0
cc_546 N_A_490_366#_c_521_n N_A_1266_74#_c_1283_n 0.00205017f $X=5.48 $Y=0.65
+ $X2=0 $Y2=0
cc_547 N_A_490_366#_c_522_n N_A_1266_74#_c_1283_n 0.00851496f $X=7.25 $Y=0.34
+ $X2=0 $Y2=0
cc_548 N_A_490_366#_c_515_n N_A_1266_74#_c_1243_n 0.00750067f $X=6.255 $Y=1.195
+ $X2=0 $Y2=0
cc_549 N_A_490_366#_c_516_n N_A_1266_74#_c_1243_n 0.00921579f $X=6.69 $Y=1.27
+ $X2=0 $Y2=0
cc_550 N_A_490_366#_c_517_n N_A_1266_74#_c_1243_n 0.00149703f $X=6.33 $Y=1.27
+ $X2=0 $Y2=0
cc_551 N_A_490_366#_c_524_n N_A_1266_74#_c_1243_n 0.00662434f $X=7.13 $Y=2.14
+ $X2=0 $Y2=0
cc_552 N_A_490_366#_c_528_n N_A_1266_74#_c_1243_n 6.18001e-19 $X=6.855 $Y=1.18
+ $X2=0 $Y2=0
cc_553 N_A_490_366#_c_529_n N_A_1266_74#_c_1243_n 0.0224751f $X=7.335 $Y=1.18
+ $X2=0 $Y2=0
cc_554 N_A_490_366#_c_535_n N_A_1266_74#_c_1256_n 0.00556629f $X=7.265 $Y=2.39
+ $X2=0 $Y2=0
cc_555 N_A_490_366#_c_524_n N_A_1266_74#_c_1256_n 0.0279379f $X=7.13 $Y=2.14
+ $X2=0 $Y2=0
cc_556 N_A_490_366#_c_516_n N_A_1266_74#_c_1244_n 0.00430336f $X=6.69 $Y=1.27
+ $X2=0 $Y2=0
cc_557 N_A_490_366#_c_522_n N_A_1266_74#_c_1244_n 0.0414158f $X=7.25 $Y=0.34
+ $X2=0 $Y2=0
cc_558 N_A_490_366#_c_525_n N_A_1266_74#_c_1244_n 0.0196081f $X=7.335 $Y=1.015
+ $X2=0 $Y2=0
cc_559 N_A_490_366#_c_528_n N_A_1266_74#_c_1244_n 0.00746605f $X=6.855 $Y=1.18
+ $X2=0 $Y2=0
cc_560 N_A_490_366#_c_529_n N_A_1266_74#_c_1244_n 0.030444f $X=7.335 $Y=1.18
+ $X2=0 $Y2=0
cc_561 N_A_490_366#_c_535_n N_A_1266_74#_c_1269_n 0.0145082f $X=7.265 $Y=2.39
+ $X2=0 $Y2=0
cc_562 N_A_490_366#_c_524_n N_A_1266_74#_c_1269_n 0.0232672f $X=7.13 $Y=2.14
+ $X2=0 $Y2=0
cc_563 N_A_490_366#_c_535_n N_A_1266_74#_c_1257_n 0.00566122f $X=7.265 $Y=2.39
+ $X2=0 $Y2=0
cc_564 N_A_490_366#_c_524_n N_A_1266_74#_c_1257_n 0.0462528f $X=7.13 $Y=2.14
+ $X2=0 $Y2=0
cc_565 N_A_490_366#_c_524_n N_A_1266_74#_c_1246_n 0.0142973f $X=7.13 $Y=2.14
+ $X2=0 $Y2=0
cc_566 N_A_490_366#_c_516_n N_A_1266_74#_c_1247_n 0.0016242f $X=6.69 $Y=1.27
+ $X2=0 $Y2=0
cc_567 N_A_490_366#_c_524_n N_A_1266_74#_c_1247_n 0.00830682f $X=7.13 $Y=2.14
+ $X2=0 $Y2=0
cc_568 N_A_490_366#_c_535_n N_VPWR_c_1466_n 0.00391396f $X=7.265 $Y=2.39 $X2=0
+ $Y2=0
cc_569 N_A_490_366#_c_532_n N_VPWR_c_1450_n 9.49986e-19 $X=3.4 $Y=2.21 $X2=0
+ $Y2=0
cc_570 N_A_490_366#_c_535_n N_VPWR_c_1450_n 0.0052212f $X=7.265 $Y=2.39 $X2=0
+ $Y2=0
cc_571 N_A_490_366#_M1008_d N_A_30_78#_c_1597_n 0.00662255f $X=2.45 $Y=1.83
+ $X2=0 $Y2=0
cc_572 N_A_490_366#_c_536_n N_A_30_78#_c_1597_n 0.0181445f $X=2.6 $Y=1.99 $X2=0
+ $Y2=0
cc_573 N_A_490_366#_c_537_n N_A_30_78#_c_1597_n 0.00414618f $X=3.035 $Y=1.725
+ $X2=0 $Y2=0
cc_574 N_A_490_366#_M1001_g N_A_30_78#_c_1592_n 2.75531e-19 $X=4.005 $Y=0.9
+ $X2=0 $Y2=0
cc_575 N_A_490_366#_c_519_n N_A_30_78#_c_1592_n 0.0194639f $X=4.265 $Y=0.415
+ $X2=0 $Y2=0
cc_576 N_A_490_366#_c_526_n N_A_30_78#_c_1592_n 0.0427756f $X=2.772 $Y=0.415
+ $X2=0 $Y2=0
cc_577 N_A_490_366#_c_531_n N_A_30_78#_c_1598_n 0.00448462f $X=3.4 $Y=2.12 $X2=0
+ $Y2=0
cc_578 N_A_490_366#_c_532_n N_A_30_78#_c_1598_n 0.0101252f $X=3.4 $Y=2.21 $X2=0
+ $Y2=0
cc_579 N_A_490_366#_c_512_n N_A_30_78#_c_1598_n 0.00156196f $X=3.79 $Y=1.635
+ $X2=0 $Y2=0
cc_580 N_A_490_366#_c_520_n N_A_30_78#_c_1598_n 0.0097192f $X=3.33 $Y=1.725
+ $X2=0 $Y2=0
cc_581 N_A_490_366#_c_530_n N_A_30_78#_c_1598_n 0.00122679f $X=3.33 $Y=1.635
+ $X2=0 $Y2=0
cc_582 N_A_490_366#_c_531_n N_A_30_78#_c_1593_n 0.00412111f $X=3.4 $Y=2.12 $X2=0
+ $Y2=0
cc_583 N_A_490_366#_c_512_n N_A_30_78#_c_1593_n 0.0131241f $X=3.79 $Y=1.635
+ $X2=0 $Y2=0
cc_584 N_A_490_366#_c_513_n N_A_30_78#_c_1593_n 0.00396133f $X=4.005 $Y=1.405
+ $X2=0 $Y2=0
cc_585 N_A_490_366#_c_518_n N_A_30_78#_c_1593_n 0.00565419f $X=2.95 $Y=1.56
+ $X2=0 $Y2=0
cc_586 N_A_490_366#_c_520_n N_A_30_78#_c_1593_n 0.0254409f $X=3.33 $Y=1.725
+ $X2=0 $Y2=0
cc_587 N_A_490_366#_c_530_n N_A_30_78#_c_1593_n 0.00325156f $X=3.33 $Y=1.635
+ $X2=0 $Y2=0
cc_588 N_A_490_366#_c_531_n N_A_30_78#_c_1603_n 3.7627e-19 $X=3.4 $Y=2.12 $X2=0
+ $Y2=0
cc_589 N_A_490_366#_c_532_n N_A_30_78#_c_1603_n 0.00332132f $X=3.4 $Y=2.21 $X2=0
+ $Y2=0
cc_590 N_A_490_366#_c_536_n N_A_30_78#_c_1603_n 0.00626245f $X=2.6 $Y=1.99 $X2=0
+ $Y2=0
cc_591 N_A_490_366#_c_537_n N_A_30_78#_c_1603_n 0.00177774f $X=3.035 $Y=1.725
+ $X2=0 $Y2=0
cc_592 N_A_490_366#_c_520_n N_A_30_78#_c_1603_n 0.0153036f $X=3.33 $Y=1.725
+ $X2=0 $Y2=0
cc_593 N_A_490_366#_c_530_n N_A_30_78#_c_1603_n 0.00209501f $X=3.33 $Y=1.635
+ $X2=0 $Y2=0
cc_594 N_A_490_366#_c_512_n N_A_30_78#_c_1595_n 8.36337e-19 $X=3.79 $Y=1.635
+ $X2=0 $Y2=0
cc_595 N_A_490_366#_M1001_g N_A_30_78#_c_1595_n 8.19151e-19 $X=4.005 $Y=0.9
+ $X2=0 $Y2=0
cc_596 N_A_490_366#_c_518_n N_A_30_78#_c_1595_n 0.0128908f $X=2.95 $Y=1.56 $X2=0
+ $Y2=0
cc_597 N_A_490_366#_c_520_n N_A_30_78#_c_1595_n 0.0153589f $X=3.33 $Y=1.725
+ $X2=0 $Y2=0
cc_598 N_A_490_366#_c_530_n N_A_30_78#_c_1595_n 0.00300406f $X=3.33 $Y=1.635
+ $X2=0 $Y2=0
cc_599 N_A_490_366#_c_521_n N_VGND_M1010_d 0.00922416f $X=5.48 $Y=0.65 $X2=0
+ $Y2=0
cc_600 N_A_490_366#_c_526_n N_VGND_c_1746_n 0.019376f $X=2.772 $Y=0.415 $X2=0
+ $Y2=0
cc_601 N_A_490_366#_c_522_n N_VGND_c_1747_n 0.00831292f $X=7.25 $Y=0.34 $X2=0
+ $Y2=0
cc_602 N_A_490_366#_c_525_n N_VGND_c_1747_n 0.00983536f $X=7.335 $Y=1.015 $X2=0
+ $Y2=0
cc_603 N_A_490_366#_c_519_n N_VGND_c_1754_n 0.0538921f $X=4.265 $Y=0.415 $X2=0
+ $Y2=0
cc_604 N_A_490_366#_c_521_n N_VGND_c_1754_n 0.0390983f $X=5.48 $Y=0.65 $X2=0
+ $Y2=0
cc_605 N_A_490_366#_c_523_n N_VGND_c_1754_n 0.0107916f $X=5.65 $Y=0.34 $X2=0
+ $Y2=0
cc_606 N_A_490_366#_c_526_n N_VGND_c_1754_n 0.0249143f $X=2.772 $Y=0.415 $X2=0
+ $Y2=0
cc_607 N_A_490_366#_c_527_n N_VGND_c_1754_n 0.0104006f $X=4.35 $Y=0.415 $X2=0
+ $Y2=0
cc_608 N_A_490_366#_c_515_n N_VGND_c_1755_n 0.00278271f $X=6.255 $Y=1.195 $X2=0
+ $Y2=0
cc_609 N_A_490_366#_c_521_n N_VGND_c_1755_n 0.00286598f $X=5.48 $Y=0.65 $X2=0
+ $Y2=0
cc_610 N_A_490_366#_c_522_n N_VGND_c_1755_n 0.114761f $X=7.25 $Y=0.34 $X2=0
+ $Y2=0
cc_611 N_A_490_366#_c_523_n N_VGND_c_1755_n 0.0117553f $X=5.65 $Y=0.34 $X2=0
+ $Y2=0
cc_612 N_A_490_366#_c_515_n N_VGND_c_1761_n 0.00361111f $X=6.255 $Y=1.195 $X2=0
+ $Y2=0
cc_613 N_A_490_366#_c_519_n N_VGND_c_1761_n 0.044091f $X=4.265 $Y=0.415 $X2=0
+ $Y2=0
cc_614 N_A_490_366#_c_521_n N_VGND_c_1761_n 0.0209417f $X=5.48 $Y=0.65 $X2=0
+ $Y2=0
cc_615 N_A_490_366#_c_522_n N_VGND_c_1761_n 0.0660751f $X=7.25 $Y=0.34 $X2=0
+ $Y2=0
cc_616 N_A_490_366#_c_523_n N_VGND_c_1761_n 0.00639038f $X=5.65 $Y=0.34 $X2=0
+ $Y2=0
cc_617 N_A_490_366#_c_526_n N_VGND_c_1761_n 0.0193906f $X=2.772 $Y=0.415 $X2=0
+ $Y2=0
cc_618 N_A_490_366#_c_527_n N_VGND_c_1761_n 0.00617686f $X=4.35 $Y=0.415 $X2=0
+ $Y2=0
cc_619 N_A_490_366#_c_521_n A_894_138# 0.00134267f $X=5.48 $Y=0.65 $X2=-0.19
+ $Y2=-0.245
cc_620 N_A_830_359#_c_732_n N_A_695_457#_M1031_g 0.0122404f $X=5.82 $Y=0.99
+ $X2=0 $Y2=0
cc_621 N_A_830_359#_c_715_n N_A_695_457#_M1031_g 0.00563857f $X=5.985 $Y=0.855
+ $X2=0 $Y2=0
cc_622 N_A_830_359#_c_716_n N_A_695_457#_M1031_g 0.0019205f $X=6.145 $Y=1.865
+ $X2=0 $Y2=0
cc_623 N_A_830_359#_c_716_n N_A_695_457#_c_806_n 0.00373472f $X=6.145 $Y=1.865
+ $X2=0 $Y2=0
cc_624 N_A_830_359#_c_717_n N_A_695_457#_c_800_n 0.00706419f $X=4.24 $Y=2.21
+ $X2=0 $Y2=0
cc_625 N_A_830_359#_M1018_g N_A_695_457#_c_800_n 0.00220779f $X=4.395 $Y=0.9
+ $X2=0 $Y2=0
cc_626 N_A_830_359#_c_714_n N_A_695_457#_c_800_n 0.0748432f $X=4.355 $Y=1.96
+ $X2=0 $Y2=0
cc_627 N_A_830_359#_c_717_n N_A_695_457#_c_816_n 0.0157202f $X=4.24 $Y=2.21
+ $X2=0 $Y2=0
cc_628 N_A_830_359#_c_714_n N_A_695_457#_c_816_n 0.00719989f $X=4.355 $Y=1.96
+ $X2=0 $Y2=0
cc_629 N_A_830_359#_c_717_n N_A_695_457#_c_808_n 7.54883e-19 $X=4.24 $Y=2.21
+ $X2=0 $Y2=0
cc_630 N_A_830_359#_c_717_n N_A_695_457#_c_801_n 0.00376557f $X=4.24 $Y=2.21
+ $X2=0 $Y2=0
cc_631 N_A_830_359#_M1018_g N_A_695_457#_c_801_n 0.00139327f $X=4.395 $Y=0.9
+ $X2=0 $Y2=0
cc_632 N_A_830_359#_c_714_n N_A_695_457#_c_801_n 0.0386689f $X=4.355 $Y=1.96
+ $X2=0 $Y2=0
cc_633 N_A_830_359#_M1018_g N_A_695_457#_c_802_n 0.00230788f $X=4.395 $Y=0.9
+ $X2=0 $Y2=0
cc_634 N_A_830_359#_c_714_n N_A_695_457#_c_802_n 0.026724f $X=4.355 $Y=1.96
+ $X2=0 $Y2=0
cc_635 N_A_830_359#_c_732_n N_A_695_457#_c_802_n 0.0115313f $X=5.82 $Y=0.99
+ $X2=0 $Y2=0
cc_636 N_A_830_359#_c_732_n N_A_695_457#_c_803_n 0.0585986f $X=5.82 $Y=0.99
+ $X2=0 $Y2=0
cc_637 N_A_830_359#_c_716_n N_A_695_457#_c_803_n 0.0159069f $X=6.145 $Y=1.865
+ $X2=0 $Y2=0
cc_638 N_A_830_359#_c_732_n N_A_695_457#_c_804_n 0.00636706f $X=5.82 $Y=0.99
+ $X2=0 $Y2=0
cc_639 N_A_830_359#_c_715_n N_A_695_457#_c_804_n 0.00593666f $X=5.985 $Y=0.855
+ $X2=0 $Y2=0
cc_640 N_A_830_359#_c_716_n N_A_695_457#_c_804_n 0.00831051f $X=6.145 $Y=1.865
+ $X2=0 $Y2=0
cc_641 N_A_830_359#_c_717_n N_A_695_457#_c_840_n 8.29006e-19 $X=4.24 $Y=2.21
+ $X2=0 $Y2=0
cc_642 N_A_830_359#_c_717_n N_A_306_74#_c_944_n 0.00323347f $X=4.24 $Y=2.21
+ $X2=0 $Y2=0
cc_643 N_A_830_359#_c_717_n N_A_306_74#_c_946_n 0.0314576f $X=4.24 $Y=2.21 $X2=0
+ $Y2=0
cc_644 N_A_830_359#_c_717_n N_A_306_74#_c_947_n 0.00852675f $X=4.24 $Y=2.21
+ $X2=0 $Y2=0
cc_645 N_A_830_359#_c_720_n N_A_306_74#_c_947_n 0.00611621f $X=6.145 $Y=2.03
+ $X2=0 $Y2=0
cc_646 N_A_830_359#_c_720_n N_A_306_74#_M1022_g 0.00116389f $X=6.145 $Y=2.03
+ $X2=0 $Y2=0
cc_647 N_A_830_359#_c_716_n N_A_306_74#_M1022_g 4.46008e-19 $X=6.145 $Y=1.865
+ $X2=0 $Y2=0
cc_648 N_A_830_359#_c_720_n N_A_306_74#_c_932_n 6.78448e-19 $X=6.145 $Y=2.03
+ $X2=0 $Y2=0
cc_649 N_A_830_359#_c_716_n N_A_306_74#_c_932_n 0.00196898f $X=6.145 $Y=1.865
+ $X2=0 $Y2=0
cc_650 N_A_830_359#_c_715_n N_A_1266_74#_c_1243_n 0.03852f $X=5.985 $Y=0.855
+ $X2=0 $Y2=0
cc_651 N_A_830_359#_c_720_n N_A_1266_74#_c_1256_n 0.0206296f $X=6.145 $Y=2.03
+ $X2=0 $Y2=0
cc_652 N_A_830_359#_c_716_n N_A_1266_74#_c_1256_n 0.00813918f $X=6.145 $Y=1.865
+ $X2=0 $Y2=0
cc_653 N_A_830_359#_c_716_n N_A_1266_74#_c_1247_n 0.0129729f $X=6.145 $Y=1.865
+ $X2=0 $Y2=0
cc_654 N_A_830_359#_c_717_n N_VPWR_c_1455_n 0.00274139f $X=4.24 $Y=2.21 $X2=0
+ $Y2=0
cc_655 N_A_830_359#_c_732_n N_VPWR_c_1457_n 0.00363609f $X=5.82 $Y=0.99 $X2=0
+ $Y2=0
cc_656 N_A_830_359#_c_720_n N_VPWR_c_1457_n 0.0405057f $X=6.145 $Y=2.03 $X2=0
+ $Y2=0
cc_657 N_A_830_359#_c_720_n N_VPWR_c_1466_n 0.00670512f $X=6.145 $Y=2.03 $X2=0
+ $Y2=0
cc_658 N_A_830_359#_c_717_n N_VPWR_c_1450_n 9.49986e-19 $X=4.24 $Y=2.21 $X2=0
+ $Y2=0
cc_659 N_A_830_359#_c_720_n N_VPWR_c_1450_n 0.00907985f $X=6.145 $Y=2.03 $X2=0
+ $Y2=0
cc_660 N_A_830_359#_c_732_n N_VGND_M1010_d 0.00954133f $X=5.82 $Y=0.99 $X2=0
+ $Y2=0
cc_661 N_A_830_359#_M1018_g N_VGND_c_1754_n 0.00110217f $X=4.395 $Y=0.9 $X2=0
+ $Y2=0
cc_662 N_A_830_359#_M1018_g N_VGND_c_1761_n 0.0010844f $X=4.395 $Y=0.9 $X2=0
+ $Y2=0
cc_663 N_A_830_359#_c_732_n A_894_138# 0.00510431f $X=5.82 $Y=0.99 $X2=-0.19
+ $Y2=-0.245
cc_664 N_A_695_457#_c_800_n N_A_306_74#_c_928_n 2.82786e-19 $X=4.01 $Y=2.4 $X2=0
+ $Y2=0
cc_665 N_A_695_457#_c_808_n N_A_306_74#_c_942_n 0.00372484f $X=4.095 $Y=2.485
+ $X2=0 $Y2=0
cc_666 N_A_695_457#_c_800_n N_A_306_74#_c_930_n 9.66665e-19 $X=4.01 $Y=2.4 $X2=0
+ $Y2=0
cc_667 N_A_695_457#_c_805_n N_A_306_74#_c_930_n 0.00203896f $X=4.01 $Y=0.86
+ $X2=0 $Y2=0
cc_668 N_A_695_457#_c_808_n N_A_306_74#_c_944_n 4.95605e-19 $X=4.095 $Y=2.485
+ $X2=0 $Y2=0
cc_669 N_A_695_457#_c_800_n N_A_306_74#_c_946_n 0.00175753f $X=4.01 $Y=2.4 $X2=0
+ $Y2=0
cc_670 N_A_695_457#_c_808_n N_A_306_74#_c_946_n 0.0120351f $X=4.095 $Y=2.485
+ $X2=0 $Y2=0
cc_671 N_A_695_457#_c_806_n N_A_306_74#_c_947_n 0.0104018f $X=5.88 $Y=1.66 $X2=0
+ $Y2=0
cc_672 N_A_695_457#_c_816_n N_A_306_74#_c_947_n 0.00293629f $X=4.615 $Y=2.485
+ $X2=0 $Y2=0
cc_673 N_A_695_457#_c_808_n N_A_306_74#_c_947_n 0.00246339f $X=4.095 $Y=2.485
+ $X2=0 $Y2=0
cc_674 N_A_695_457#_c_811_n N_A_306_74#_c_947_n 0.00523168f $X=5.085 $Y=2.485
+ $X2=0 $Y2=0
cc_675 N_A_695_457#_c_840_n N_A_306_74#_c_947_n 0.001324f $X=4.7 $Y=2.445 $X2=0
+ $Y2=0
cc_676 N_A_695_457#_c_806_n N_A_306_74#_M1022_g 0.00888826f $X=5.88 $Y=1.66
+ $X2=0 $Y2=0
cc_677 N_A_695_457#_c_806_n N_A_306_74#_c_932_n 0.00427682f $X=5.88 $Y=1.66
+ $X2=0 $Y2=0
cc_678 N_A_695_457#_c_804_n N_A_306_74#_c_932_n 0.00245186f $X=5.485 $Y=1.41
+ $X2=0 $Y2=0
cc_679 N_A_695_457#_c_816_n N_VPWR_M1007_d 0.00582643f $X=4.615 $Y=2.485 $X2=0
+ $Y2=0
cc_680 N_A_695_457#_c_801_n N_VPWR_M1007_d 4.45955e-19 $X=4.7 $Y=2.32 $X2=0
+ $Y2=0
cc_681 N_A_695_457#_c_840_n N_VPWR_M1007_d 0.00220216f $X=4.7 $Y=2.445 $X2=0
+ $Y2=0
cc_682 N_A_695_457#_c_816_n N_VPWR_c_1455_n 0.0180683f $X=4.615 $Y=2.485 $X2=0
+ $Y2=0
cc_683 N_A_695_457#_c_840_n N_VPWR_c_1455_n 0.00862169f $X=4.7 $Y=2.445 $X2=0
+ $Y2=0
cc_684 N_A_695_457#_c_811_n N_VPWR_c_1456_n 0.00589153f $X=5.085 $Y=2.485 $X2=0
+ $Y2=0
cc_685 N_A_695_457#_c_840_n N_VPWR_c_1456_n 5.93009e-19 $X=4.7 $Y=2.445 $X2=0
+ $Y2=0
cc_686 N_A_695_457#_c_806_n N_VPWR_c_1457_n 0.0131452f $X=5.88 $Y=1.66 $X2=0
+ $Y2=0
cc_687 N_A_695_457#_c_803_n N_VPWR_c_1457_n 0.0133374f $X=5.485 $Y=1.41 $X2=0
+ $Y2=0
cc_688 N_A_695_457#_c_804_n N_VPWR_c_1457_n 0.00741213f $X=5.485 $Y=1.41 $X2=0
+ $Y2=0
cc_689 N_A_695_457#_c_811_n N_VPWR_c_1457_n 0.0177113f $X=5.085 $Y=2.485 $X2=0
+ $Y2=0
cc_690 N_A_695_457#_c_816_n N_VPWR_c_1465_n 0.00300657f $X=4.615 $Y=2.485 $X2=0
+ $Y2=0
cc_691 N_A_695_457#_c_808_n N_VPWR_c_1465_n 0.0104385f $X=4.095 $Y=2.485 $X2=0
+ $Y2=0
cc_692 N_A_695_457#_c_806_n N_VPWR_c_1450_n 9.14192e-19 $X=5.88 $Y=1.66 $X2=0
+ $Y2=0
cc_693 N_A_695_457#_c_816_n N_VPWR_c_1450_n 0.00708968f $X=4.615 $Y=2.485 $X2=0
+ $Y2=0
cc_694 N_A_695_457#_c_808_n N_VPWR_c_1450_n 0.0154047f $X=4.095 $Y=2.485 $X2=0
+ $Y2=0
cc_695 N_A_695_457#_c_811_n N_VPWR_c_1450_n 0.0102762f $X=5.085 $Y=2.485 $X2=0
+ $Y2=0
cc_696 N_A_695_457#_c_840_n N_VPWR_c_1450_n 0.0021032f $X=4.7 $Y=2.445 $X2=0
+ $Y2=0
cc_697 N_A_695_457#_c_800_n N_A_30_78#_c_1592_n 0.00468745f $X=4.01 $Y=2.4 $X2=0
+ $Y2=0
cc_698 N_A_695_457#_c_805_n N_A_30_78#_c_1592_n 0.014451f $X=4.01 $Y=0.86 $X2=0
+ $Y2=0
cc_699 N_A_695_457#_c_800_n N_A_30_78#_c_1598_n 0.0135316f $X=4.01 $Y=2.4 $X2=0
+ $Y2=0
cc_700 N_A_695_457#_c_808_n N_A_30_78#_c_1598_n 0.0195289f $X=4.095 $Y=2.485
+ $X2=0 $Y2=0
cc_701 N_A_695_457#_c_800_n N_A_30_78#_c_1593_n 0.0482482f $X=4.01 $Y=2.4 $X2=0
+ $Y2=0
cc_702 N_A_695_457#_c_800_n N_A_30_78#_c_1603_n 0.00318453f $X=4.01 $Y=2.4 $X2=0
+ $Y2=0
cc_703 N_A_695_457#_c_808_n N_A_30_78#_c_1603_n 0.0225697f $X=4.095 $Y=2.485
+ $X2=0 $Y2=0
cc_704 N_A_695_457#_c_800_n N_A_30_78#_c_1595_n 0.0139397f $X=4.01 $Y=2.4 $X2=0
+ $Y2=0
cc_705 N_A_695_457#_c_805_n N_A_30_78#_c_1595_n 0.00972762f $X=4.01 $Y=0.86
+ $X2=0 $Y2=0
cc_706 N_A_695_457#_c_800_n A_785_457# 0.00135518f $X=4.01 $Y=2.4 $X2=-0.19
+ $Y2=-0.245
cc_707 N_A_695_457#_c_816_n A_785_457# 3.73291e-19 $X=4.615 $Y=2.485 $X2=-0.19
+ $Y2=-0.245
cc_708 N_A_695_457#_c_808_n A_785_457# 0.00191536f $X=4.095 $Y=2.485 $X2=-0.19
+ $Y2=-0.245
cc_709 N_A_695_457#_M1031_g N_VGND_c_1754_n 0.00366947f $X=5.44 $Y=0.74 $X2=0
+ $Y2=0
cc_710 N_A_695_457#_M1031_g N_VGND_c_1755_n 0.00309023f $X=5.44 $Y=0.74 $X2=0
+ $Y2=0
cc_711 N_A_695_457#_M1031_g N_VGND_c_1761_n 0.00393738f $X=5.44 $Y=0.74 $X2=0
+ $Y2=0
cc_712 N_A_306_74#_M1020_g N_A_1518_203#_M1019_g 0.0368892f $X=7.305 $Y=0.615
+ $X2=0 $Y2=0
cc_713 N_A_306_74#_M1020_g N_A_1518_203#_c_1117_n 0.0235039f $X=7.305 $Y=0.615
+ $X2=0 $Y2=0
cc_714 N_A_306_74#_M1020_g N_A_1518_203#_c_1121_n 3.81559e-19 $X=7.305 $Y=0.615
+ $X2=0 $Y2=0
cc_715 N_A_306_74#_M1020_g N_A_1518_203#_c_1122_n 0.0205557f $X=7.305 $Y=0.615
+ $X2=0 $Y2=0
cc_716 N_A_306_74#_c_932_n N_A_1266_74#_c_1243_n 2.4837e-19 $X=6.475 $Y=1.66
+ $X2=0 $Y2=0
cc_717 N_A_306_74#_M1022_g N_A_1266_74#_c_1256_n 0.00801796f $X=6.385 $Y=2.385
+ $X2=0 $Y2=0
cc_718 N_A_306_74#_c_931_n N_A_1266_74#_c_1256_n 0.00695524f $X=7.23 $Y=1.66
+ $X2=0 $Y2=0
cc_719 N_A_306_74#_c_932_n N_A_1266_74#_c_1256_n 0.00199946f $X=6.475 $Y=1.66
+ $X2=0 $Y2=0
cc_720 N_A_306_74#_M1020_g N_A_1266_74#_c_1244_n 0.00507341f $X=7.305 $Y=0.615
+ $X2=0 $Y2=0
cc_721 N_A_306_74#_c_931_n N_A_1266_74#_c_1257_n 3.51038e-19 $X=7.23 $Y=1.66
+ $X2=0 $Y2=0
cc_722 N_A_306_74#_M1020_g N_A_1266_74#_c_1246_n 0.00127921f $X=7.305 $Y=0.615
+ $X2=0 $Y2=0
cc_723 N_A_306_74#_c_931_n N_A_1266_74#_c_1247_n 0.00490084f $X=7.23 $Y=1.66
+ $X2=0 $Y2=0
cc_724 N_A_306_74#_c_932_n N_A_1266_74#_c_1247_n 0.00528124f $X=6.475 $Y=1.66
+ $X2=0 $Y2=0
cc_725 N_A_306_74#_M1020_g N_A_1266_74#_c_1247_n 2.86702e-19 $X=7.305 $Y=0.615
+ $X2=0 $Y2=0
cc_726 N_A_306_74#_c_939_n N_VPWR_c_1454_n 0.00953832f $X=2.375 $Y=1.755 $X2=0
+ $Y2=0
cc_727 N_A_306_74#_c_927_n N_VPWR_c_1454_n 0.00194465f $X=2.88 $Y=3.075 $X2=0
+ $Y2=0
cc_728 N_A_306_74#_c_943_n N_VPWR_c_1454_n 0.00263858f $X=2.955 $Y=3.15 $X2=0
+ $Y2=0
cc_729 N_A_306_74#_c_944_n N_VPWR_c_1455_n 0.00685937f $X=3.85 $Y=2.87 $X2=0
+ $Y2=0
cc_730 N_A_306_74#_c_947_n N_VPWR_c_1455_n 0.0250293f $X=6.295 $Y=3.15 $X2=0
+ $Y2=0
cc_731 N_A_306_74#_c_947_n N_VPWR_c_1456_n 0.0218819f $X=6.295 $Y=3.15 $X2=0
+ $Y2=0
cc_732 N_A_306_74#_c_947_n N_VPWR_c_1457_n 0.0259878f $X=6.295 $Y=3.15 $X2=0
+ $Y2=0
cc_733 N_A_306_74#_M1022_g N_VPWR_c_1457_n 0.00308789f $X=6.385 $Y=2.385 $X2=0
+ $Y2=0
cc_734 N_A_306_74#_c_952_n N_VPWR_c_1457_n 0.00312383f $X=6.385 $Y=3.15 $X2=0
+ $Y2=0
cc_735 N_A_306_74#_c_939_n N_VPWR_c_1465_n 0.00512473f $X=2.375 $Y=1.755 $X2=0
+ $Y2=0
cc_736 N_A_306_74#_c_943_n N_VPWR_c_1465_n 0.0455433f $X=2.955 $Y=3.15 $X2=0
+ $Y2=0
cc_737 N_A_306_74#_c_947_n N_VPWR_c_1466_n 0.0203278f $X=6.295 $Y=3.15 $X2=0
+ $Y2=0
cc_738 N_A_306_74#_c_939_n N_VPWR_c_1450_n 0.00492022f $X=2.375 $Y=1.755 $X2=0
+ $Y2=0
cc_739 N_A_306_74#_c_942_n N_VPWR_c_1450_n 0.0243846f $X=3.76 $Y=3.15 $X2=0
+ $Y2=0
cc_740 N_A_306_74#_c_943_n N_VPWR_c_1450_n 0.00710688f $X=2.955 $Y=3.15 $X2=0
+ $Y2=0
cc_741 N_A_306_74#_c_947_n N_VPWR_c_1450_n 0.0536469f $X=6.295 $Y=3.15 $X2=0
+ $Y2=0
cc_742 N_A_306_74#_c_951_n N_VPWR_c_1450_n 0.00541294f $X=3.85 $Y=3.15 $X2=0
+ $Y2=0
cc_743 N_A_306_74#_c_952_n N_VPWR_c_1450_n 0.0128115f $X=6.385 $Y=3.15 $X2=0
+ $Y2=0
cc_744 N_A_306_74#_c_934_n N_A_30_78#_c_1591_n 0.00411959f $X=1.675 $Y=0.515
+ $X2=0 $Y2=0
cc_745 N_A_306_74#_c_938_n N_A_30_78#_c_1591_n 0.00499191f $X=1.647 $Y=1.055
+ $X2=0 $Y2=0
cc_746 N_A_306_74#_M1005_s N_A_30_78#_c_1597_n 0.00354211f $X=1.57 $Y=1.83 $X2=0
+ $Y2=0
cc_747 N_A_306_74#_c_939_n N_A_30_78#_c_1597_n 0.01258f $X=2.375 $Y=1.755 $X2=0
+ $Y2=0
cc_748 N_A_306_74#_c_927_n N_A_30_78#_c_1597_n 0.012732f $X=2.88 $Y=3.075 $X2=0
+ $Y2=0
cc_749 N_A_306_74#_c_954_n N_A_30_78#_c_1597_n 0.00796796f $X=1.7 $Y=1.975 $X2=0
+ $Y2=0
cc_750 N_A_306_74#_c_928_n N_A_30_78#_c_1592_n 0.00482311f $X=3.43 $Y=1.275
+ $X2=0 $Y2=0
cc_751 N_A_306_74#_c_930_n N_A_30_78#_c_1592_n 0.00917108f $X=3.505 $Y=1.2 $X2=0
+ $Y2=0
cc_752 N_A_306_74#_c_946_n N_A_30_78#_c_1598_n 6.36667e-19 $X=3.85 $Y=2.78 $X2=0
+ $Y2=0
cc_753 N_A_306_74#_c_929_n N_A_30_78#_c_1593_n 5.58713e-19 $X=2.955 $Y=1.275
+ $X2=0 $Y2=0
cc_754 N_A_306_74#_c_954_n N_A_30_78#_c_1601_n 0.0157663f $X=1.7 $Y=1.975 $X2=0
+ $Y2=0
cc_755 N_A_306_74#_M1005_s N_A_30_78#_c_1602_n 0.00464207f $X=1.57 $Y=1.83 $X2=0
+ $Y2=0
cc_756 N_A_306_74#_c_927_n N_A_30_78#_c_1603_n 0.0117672f $X=2.88 $Y=3.075 $X2=0
+ $Y2=0
cc_757 N_A_306_74#_c_942_n N_A_30_78#_c_1603_n 0.00422515f $X=3.76 $Y=3.15 $X2=0
+ $Y2=0
cc_758 N_A_306_74#_c_928_n N_A_30_78#_c_1595_n 0.0147846f $X=3.43 $Y=1.275 $X2=0
+ $Y2=0
cc_759 N_A_306_74#_c_936_n N_VGND_M1003_d 0.00250873f $X=2.445 $Y=1.055 $X2=0
+ $Y2=0
cc_760 N_A_306_74#_c_934_n N_VGND_c_1745_n 0.0388154f $X=1.675 $Y=0.515 $X2=0
+ $Y2=0
cc_761 N_A_306_74#_c_926_n N_VGND_c_1746_n 0.0116945f $X=2.39 $Y=1.2 $X2=0 $Y2=0
cc_762 N_A_306_74#_c_934_n N_VGND_c_1746_n 0.0180786f $X=1.675 $Y=0.515 $X2=0
+ $Y2=0
cc_763 N_A_306_74#_c_936_n N_VGND_c_1746_n 0.0210288f $X=2.445 $Y=1.055 $X2=0
+ $Y2=0
cc_764 N_A_306_74#_M1020_g N_VGND_c_1747_n 5.78056e-19 $X=7.305 $Y=0.615 $X2=0
+ $Y2=0
cc_765 N_A_306_74#_c_934_n N_VGND_c_1753_n 0.0170181f $X=1.675 $Y=0.515 $X2=0
+ $Y2=0
cc_766 N_A_306_74#_c_926_n N_VGND_c_1754_n 0.00383152f $X=2.39 $Y=1.2 $X2=0
+ $Y2=0
cc_767 N_A_306_74#_M1020_g N_VGND_c_1755_n 9.33926e-19 $X=7.305 $Y=0.615 $X2=0
+ $Y2=0
cc_768 N_A_306_74#_c_926_n N_VGND_c_1761_n 0.00762539f $X=2.39 $Y=1.2 $X2=0
+ $Y2=0
cc_769 N_A_306_74#_c_934_n N_VGND_c_1761_n 0.0140297f $X=1.675 $Y=0.515 $X2=0
+ $Y2=0
cc_770 N_A_1518_203#_c_1118_n N_A_1266_74#_M1021_g 0.0107164f $X=8.615 $Y=1.1
+ $X2=0 $Y2=0
cc_771 N_A_1518_203#_c_1119_n N_A_1266_74#_M1021_g 0.0159617f $X=8.78 $Y=0.615
+ $X2=0 $Y2=0
cc_772 N_A_1518_203#_c_1120_n N_A_1266_74#_M1021_g 0.00301146f $X=9.105 $Y=1.855
+ $X2=0 $Y2=0
cc_773 N_A_1518_203#_c_1123_n N_A_1266_74#_M1021_g 0.00389282f $X=9.105 $Y=1.1
+ $X2=0 $Y2=0
cc_774 N_A_1518_203#_c_1128_n N_A_1266_74#_c_1249_n 0.0107968f $X=9.02 $Y=1.94
+ $X2=0 $Y2=0
cc_775 N_A_1518_203#_c_1129_n N_A_1266_74#_c_1249_n 0.00310966f $X=8.685 $Y=1.94
+ $X2=0 $Y2=0
cc_776 N_A_1518_203#_c_1120_n N_A_1266_74#_c_1249_n 0.00343619f $X=9.105
+ $Y=1.855 $X2=0 $Y2=0
cc_777 N_A_1518_203#_c_1132_n N_A_1266_74#_c_1249_n 0.00678514f $X=8.502
+ $Y=2.445 $X2=0 $Y2=0
cc_778 N_A_1518_203#_c_1131_n N_A_1266_74#_c_1250_n 0.006945f $X=8.485 $Y=2.675
+ $X2=0 $Y2=0
cc_779 N_A_1518_203#_c_1132_n N_A_1266_74#_c_1250_n 0.00313845f $X=8.502
+ $Y=2.445 $X2=0 $Y2=0
cc_780 N_A_1518_203#_c_1128_n N_A_1266_74#_c_1236_n 0.00354772f $X=9.02 $Y=1.94
+ $X2=0 $Y2=0
cc_781 N_A_1518_203#_c_1120_n N_A_1266_74#_c_1236_n 0.0103302f $X=9.105 $Y=1.855
+ $X2=0 $Y2=0
cc_782 N_A_1518_203#_c_1123_n N_A_1266_74#_c_1236_n 0.00508985f $X=9.105 $Y=1.1
+ $X2=0 $Y2=0
cc_783 N_A_1518_203#_c_1129_n N_A_1266_74#_c_1237_n 7.74206e-19 $X=8.685 $Y=1.94
+ $X2=0 $Y2=0
cc_784 N_A_1518_203#_c_1123_n N_A_1266_74#_c_1237_n 8.2291e-19 $X=9.105 $Y=1.1
+ $X2=0 $Y2=0
cc_785 N_A_1518_203#_c_1120_n N_A_1266_74#_c_1238_n 0.00511666f $X=9.105
+ $Y=1.855 $X2=0 $Y2=0
cc_786 N_A_1518_203#_c_1123_n N_A_1266_74#_c_1238_n 0.00147647f $X=9.105 $Y=1.1
+ $X2=0 $Y2=0
cc_787 N_A_1518_203#_c_1128_n N_A_1266_74#_c_1253_n 6.47767e-19 $X=9.02 $Y=1.94
+ $X2=0 $Y2=0
cc_788 N_A_1518_203#_c_1120_n N_A_1266_74#_c_1253_n 0.00358035f $X=9.105
+ $Y=1.855 $X2=0 $Y2=0
cc_789 N_A_1518_203#_c_1128_n N_A_1266_74#_c_1254_n 0.00455214f $X=9.02 $Y=1.94
+ $X2=0 $Y2=0
cc_790 N_A_1518_203#_c_1132_n N_A_1266_74#_c_1254_n 9.14342e-19 $X=8.502
+ $Y=2.445 $X2=0 $Y2=0
cc_791 N_A_1518_203#_c_1119_n N_A_1266_74#_c_1240_n 2.88416e-19 $X=8.78 $Y=0.615
+ $X2=0 $Y2=0
cc_792 N_A_1518_203#_c_1123_n N_A_1266_74#_c_1240_n 0.00670166f $X=9.105 $Y=1.1
+ $X2=0 $Y2=0
cc_793 N_A_1518_203#_c_1119_n N_A_1266_74#_c_1241_n 0.00317724f $X=8.78 $Y=0.615
+ $X2=0 $Y2=0
cc_794 N_A_1518_203#_c_1120_n N_A_1266_74#_c_1242_n 0.00419613f $X=9.105
+ $Y=1.855 $X2=0 $Y2=0
cc_795 N_A_1518_203#_c_1126_n N_A_1266_74#_c_1269_n 0.00757243f $X=7.685 $Y=2.39
+ $X2=0 $Y2=0
cc_796 N_A_1518_203#_c_1124_n N_A_1266_74#_c_1257_n 0.00331106f $X=7.685
+ $Y=1.835 $X2=0 $Y2=0
cc_797 N_A_1518_203#_c_1125_n N_A_1266_74#_c_1257_n 0.0103166f $X=7.685 $Y=2.3
+ $X2=0 $Y2=0
cc_798 N_A_1518_203#_c_1126_n N_A_1266_74#_c_1257_n 0.0046186f $X=7.685 $Y=2.39
+ $X2=0 $Y2=0
cc_799 N_A_1518_203#_c_1117_n N_A_1266_74#_c_1257_n 0.0015543f $X=7.685 $Y=1.745
+ $X2=0 $Y2=0
cc_800 N_A_1518_203#_c_1124_n N_A_1266_74#_c_1245_n 8.26265e-19 $X=7.685
+ $Y=1.835 $X2=0 $Y2=0
cc_801 N_A_1518_203#_c_1117_n N_A_1266_74#_c_1245_n 0.00762694f $X=7.685
+ $Y=1.745 $X2=0 $Y2=0
cc_802 N_A_1518_203#_c_1118_n N_A_1266_74#_c_1245_n 0.0272699f $X=8.615 $Y=1.1
+ $X2=0 $Y2=0
cc_803 N_A_1518_203#_c_1129_n N_A_1266_74#_c_1245_n 4.22281e-19 $X=8.685 $Y=1.94
+ $X2=0 $Y2=0
cc_804 N_A_1518_203#_c_1121_n N_A_1266_74#_c_1245_n 0.0204811f $X=7.755 $Y=1.1
+ $X2=0 $Y2=0
cc_805 N_A_1518_203#_c_1122_n N_A_1266_74#_c_1245_n 0.00111936f $X=7.755 $Y=1.18
+ $X2=0 $Y2=0
cc_806 N_A_1518_203#_c_1117_n N_A_1266_74#_c_1246_n 0.00211774f $X=7.685
+ $Y=1.745 $X2=0 $Y2=0
cc_807 N_A_1518_203#_c_1121_n N_A_1266_74#_c_1246_n 0.0034757f $X=7.755 $Y=1.1
+ $X2=0 $Y2=0
cc_808 N_A_1518_203#_c_1118_n N_A_1266_74#_c_1248_n 0.0242574f $X=8.615 $Y=1.1
+ $X2=0 $Y2=0
cc_809 N_A_1518_203#_c_1128_n N_A_1266_74#_c_1248_n 0.0118853f $X=9.02 $Y=1.94
+ $X2=0 $Y2=0
cc_810 N_A_1518_203#_c_1129_n N_A_1266_74#_c_1248_n 0.0136054f $X=8.685 $Y=1.94
+ $X2=0 $Y2=0
cc_811 N_A_1518_203#_c_1120_n N_A_1266_74#_c_1248_n 0.0235661f $X=9.105 $Y=1.855
+ $X2=0 $Y2=0
cc_812 N_A_1518_203#_c_1120_n N_A_1864_409#_c_1397_n 2.38456e-19 $X=9.105
+ $Y=1.855 $X2=0 $Y2=0
cc_813 N_A_1518_203#_c_1128_n N_A_1864_409#_c_1404_n 0.0121572f $X=9.02 $Y=1.94
+ $X2=0 $Y2=0
cc_814 N_A_1518_203#_c_1120_n N_A_1864_409#_c_1404_n 0.00900265f $X=9.105
+ $Y=1.855 $X2=0 $Y2=0
cc_815 N_A_1518_203#_c_1119_n N_A_1864_409#_c_1399_n 0.00478045f $X=8.78
+ $Y=0.615 $X2=0 $Y2=0
cc_816 N_A_1518_203#_c_1120_n N_A_1864_409#_c_1399_n 0.0077671f $X=9.105
+ $Y=1.855 $X2=0 $Y2=0
cc_817 N_A_1518_203#_c_1123_n N_A_1864_409#_c_1399_n 0.00665068f $X=9.105 $Y=1.1
+ $X2=0 $Y2=0
cc_818 N_A_1518_203#_c_1120_n N_A_1864_409#_c_1400_n 0.0234089f $X=9.105
+ $Y=1.855 $X2=0 $Y2=0
cc_819 N_A_1518_203#_c_1126_n N_VPWR_c_1458_n 0.00654507f $X=7.685 $Y=2.39 $X2=0
+ $Y2=0
cc_820 N_A_1518_203#_c_1131_n N_VPWR_c_1458_n 0.0178695f $X=8.485 $Y=2.675 $X2=0
+ $Y2=0
cc_821 N_A_1518_203#_c_1131_n N_VPWR_c_1459_n 0.0120785f $X=8.485 $Y=2.675 $X2=0
+ $Y2=0
cc_822 N_A_1518_203#_c_1128_n N_VPWR_c_1460_n 0.0259196f $X=9.02 $Y=1.94 $X2=0
+ $Y2=0
cc_823 N_A_1518_203#_c_1132_n N_VPWR_c_1460_n 0.0548082f $X=8.502 $Y=2.445 $X2=0
+ $Y2=0
cc_824 N_A_1518_203#_c_1126_n N_VPWR_c_1466_n 0.00501877f $X=7.685 $Y=2.39 $X2=0
+ $Y2=0
cc_825 N_A_1518_203#_c_1126_n N_VPWR_c_1450_n 0.0052212f $X=7.685 $Y=2.39 $X2=0
+ $Y2=0
cc_826 N_A_1518_203#_c_1131_n N_VPWR_c_1450_n 0.0126247f $X=8.485 $Y=2.675 $X2=0
+ $Y2=0
cc_827 N_A_1518_203#_M1019_g N_VGND_c_1747_n 0.0107187f $X=7.695 $Y=0.615 $X2=0
+ $Y2=0
cc_828 N_A_1518_203#_c_1118_n N_VGND_c_1747_n 0.0130069f $X=8.615 $Y=1.1 $X2=0
+ $Y2=0
cc_829 N_A_1518_203#_c_1119_n N_VGND_c_1747_n 0.00738736f $X=8.78 $Y=0.615 $X2=0
+ $Y2=0
cc_830 N_A_1518_203#_c_1121_n N_VGND_c_1747_n 0.0145528f $X=7.755 $Y=1.1 $X2=0
+ $Y2=0
cc_831 N_A_1518_203#_c_1122_n N_VGND_c_1747_n 0.0011793f $X=7.755 $Y=1.18 $X2=0
+ $Y2=0
cc_832 N_A_1518_203#_c_1119_n N_VGND_c_1748_n 0.0303742f $X=8.78 $Y=0.615 $X2=0
+ $Y2=0
cc_833 N_A_1518_203#_c_1123_n N_VGND_c_1748_n 0.00112954f $X=9.105 $Y=1.1 $X2=0
+ $Y2=0
cc_834 N_A_1518_203#_M1019_g N_VGND_c_1755_n 0.0045897f $X=7.695 $Y=0.615 $X2=0
+ $Y2=0
cc_835 N_A_1518_203#_c_1119_n N_VGND_c_1756_n 0.0126905f $X=8.78 $Y=0.615 $X2=0
+ $Y2=0
cc_836 N_A_1518_203#_M1019_g N_VGND_c_1761_n 0.0044912f $X=7.695 $Y=0.615 $X2=0
+ $Y2=0
cc_837 N_A_1518_203#_c_1119_n N_VGND_c_1761_n 0.0118012f $X=8.78 $Y=0.615 $X2=0
+ $Y2=0
cc_838 N_A_1266_74#_c_1239_n N_A_1864_409#_c_1397_n 0.00139534f $X=9.48 $Y=1.07
+ $X2=0 $Y2=0
cc_839 N_A_1266_74#_c_1242_n N_A_1864_409#_c_1397_n 0.0154815f $X=9.245 $Y=1.52
+ $X2=0 $Y2=0
cc_840 N_A_1266_74#_c_1253_n N_A_1864_409#_c_1404_n 0.00590965f $X=9.245 $Y=1.88
+ $X2=0 $Y2=0
cc_841 N_A_1266_74#_c_1254_n N_A_1864_409#_c_1404_n 0.0105256f $X=9.245 $Y=1.97
+ $X2=0 $Y2=0
cc_842 N_A_1266_74#_c_1238_n N_A_1864_409#_c_1399_n 0.00400367f $X=9.23 $Y=1.355
+ $X2=0 $Y2=0
cc_843 N_A_1266_74#_c_1239_n N_A_1864_409#_c_1399_n 0.00708838f $X=9.48 $Y=1.07
+ $X2=0 $Y2=0
cc_844 N_A_1266_74#_c_1241_n N_A_1864_409#_c_1399_n 0.0140899f $X=9.555 $Y=0.995
+ $X2=0 $Y2=0
cc_845 N_A_1266_74#_c_1242_n N_A_1864_409#_c_1399_n 7.91947e-19 $X=9.245 $Y=1.52
+ $X2=0 $Y2=0
cc_846 N_A_1266_74#_c_1239_n N_A_1864_409#_c_1400_n 0.0079216f $X=9.48 $Y=1.07
+ $X2=0 $Y2=0
cc_847 N_A_1266_74#_c_1242_n N_A_1864_409#_c_1400_n 0.00324958f $X=9.245 $Y=1.52
+ $X2=0 $Y2=0
cc_848 N_A_1266_74#_c_1257_n N_VPWR_c_1458_n 0.00177331f $X=7.55 $Y=2.475 $X2=0
+ $Y2=0
cc_849 N_A_1266_74#_c_1250_n N_VPWR_c_1459_n 0.00477303f $X=8.71 $Y=2.39 $X2=0
+ $Y2=0
cc_850 N_A_1266_74#_c_1249_n N_VPWR_c_1460_n 0.001714f $X=8.71 $Y=2.3 $X2=0
+ $Y2=0
cc_851 N_A_1266_74#_c_1250_n N_VPWR_c_1460_n 0.00744434f $X=8.71 $Y=2.39 $X2=0
+ $Y2=0
cc_852 N_A_1266_74#_c_1236_n N_VPWR_c_1460_n 3.97376e-19 $X=9.155 $Y=1.52 $X2=0
+ $Y2=0
cc_853 N_A_1266_74#_c_1254_n N_VPWR_c_1460_n 0.0126982f $X=9.245 $Y=1.97 $X2=0
+ $Y2=0
cc_854 N_A_1266_74#_c_1269_n N_VPWR_c_1466_n 0.0213832f $X=7.465 $Y=2.64 $X2=0
+ $Y2=0
cc_855 N_A_1266_74#_c_1379_p N_VPWR_c_1466_n 0.00379401f $X=6.65 $Y=2.64 $X2=0
+ $Y2=0
cc_856 N_A_1266_74#_c_1254_n N_VPWR_c_1467_n 0.00470366f $X=9.245 $Y=1.97 $X2=0
+ $Y2=0
cc_857 N_A_1266_74#_c_1250_n N_VPWR_c_1450_n 0.0052212f $X=8.71 $Y=2.39 $X2=0
+ $Y2=0
cc_858 N_A_1266_74#_c_1254_n N_VPWR_c_1450_n 0.00473388f $X=9.245 $Y=1.97 $X2=0
+ $Y2=0
cc_859 N_A_1266_74#_c_1269_n N_VPWR_c_1450_n 0.0313462f $X=7.465 $Y=2.64 $X2=0
+ $Y2=0
cc_860 N_A_1266_74#_c_1379_p N_VPWR_c_1450_n 0.00557315f $X=6.65 $Y=2.64 $X2=0
+ $Y2=0
cc_861 N_A_1266_74#_c_1269_n A_1468_493# 0.00358233f $X=7.465 $Y=2.64 $X2=-0.19
+ $Y2=-0.245
cc_862 N_A_1266_74#_c_1241_n N_Q_c_1715_n 0.00112501f $X=9.555 $Y=0.995 $X2=0
+ $Y2=0
cc_863 N_A_1266_74#_c_1239_n N_Q_c_1716_n 0.00112501f $X=9.48 $Y=1.07 $X2=0
+ $Y2=0
cc_864 N_A_1266_74#_c_1254_n Q 0.00322019f $X=9.245 $Y=1.97 $X2=0 $Y2=0
cc_865 N_A_1266_74#_M1021_g N_VGND_c_1748_n 0.00359522f $X=8.565 $Y=0.615 $X2=0
+ $Y2=0
cc_866 N_A_1266_74#_c_1240_n N_VGND_c_1748_n 0.0104251f $X=9.305 $Y=1.07 $X2=0
+ $Y2=0
cc_867 N_A_1266_74#_c_1241_n N_VGND_c_1748_n 0.0065091f $X=9.555 $Y=0.995 $X2=0
+ $Y2=0
cc_868 N_A_1266_74#_M1021_g N_VGND_c_1756_n 0.00527282f $X=8.565 $Y=0.615 $X2=0
+ $Y2=0
cc_869 N_A_1266_74#_c_1241_n N_VGND_c_1757_n 0.00434272f $X=9.555 $Y=0.995 $X2=0
+ $Y2=0
cc_870 N_A_1266_74#_M1021_g N_VGND_c_1761_n 0.00534666f $X=8.565 $Y=0.615 $X2=0
+ $Y2=0
cc_871 N_A_1266_74#_c_1241_n N_VGND_c_1761_n 0.00830282f $X=9.555 $Y=0.995 $X2=0
+ $Y2=0
cc_872 N_A_1864_409#_c_1404_n N_VPWR_c_1460_n 0.0462745f $X=9.47 $Y=2.19 $X2=0
+ $Y2=0
cc_873 N_A_1864_409#_c_1401_n N_VPWR_c_1462_n 0.0203918f $X=10.53 $Y=1.765 $X2=0
+ $Y2=0
cc_874 N_A_1864_409#_c_1398_n N_VPWR_c_1462_n 8.22785e-19 $X=10.53 $Y=1.575
+ $X2=0 $Y2=0
cc_875 N_A_1864_409#_c_1401_n N_VPWR_c_1467_n 0.00429299f $X=10.53 $Y=1.765
+ $X2=0 $Y2=0
cc_876 N_A_1864_409#_c_1404_n N_VPWR_c_1467_n 0.00575213f $X=9.47 $Y=2.19 $X2=0
+ $Y2=0
cc_877 N_A_1864_409#_c_1401_n N_VPWR_c_1450_n 0.00852523f $X=10.53 $Y=1.765
+ $X2=0 $Y2=0
cc_878 N_A_1864_409#_c_1404_n N_VPWR_c_1450_n 0.00591657f $X=9.47 $Y=2.19 $X2=0
+ $Y2=0
cc_879 N_A_1864_409#_M1009_g N_Q_c_1715_n 0.00853833f $X=10.545 $Y=0.74 $X2=0
+ $Y2=0
cc_880 N_A_1864_409#_c_1399_n N_Q_c_1715_n 0.0694074f $X=9.77 $Y=0.645 $X2=0
+ $Y2=0
cc_881 N_A_1864_409#_M1009_g N_Q_c_1716_n 0.00343176f $X=10.545 $Y=0.74 $X2=0
+ $Y2=0
cc_882 N_A_1864_409#_c_1397_n N_Q_c_1716_n 0.00187014f $X=10.44 $Y=1.55 $X2=0
+ $Y2=0
cc_883 N_A_1864_409#_c_1397_n Q 0.0150903f $X=10.44 $Y=1.55 $X2=0 $Y2=0
cc_884 N_A_1864_409#_c_1404_n Q 0.0848083f $X=9.47 $Y=2.19 $X2=0 $Y2=0
cc_885 N_A_1864_409#_c_1400_n Q 0.017588f $X=9.77 $Y=1.55 $X2=0 $Y2=0
cc_886 N_A_1864_409#_c_1401_n N_Q_c_1717_n 0.00351033f $X=10.53 $Y=1.765 $X2=0
+ $Y2=0
cc_887 N_A_1864_409#_M1009_g N_Q_c_1717_n 0.0104864f $X=10.545 $Y=0.74 $X2=0
+ $Y2=0
cc_888 N_A_1864_409#_c_1397_n N_Q_c_1717_n 0.0395686f $X=10.44 $Y=1.55 $X2=0
+ $Y2=0
cc_889 N_A_1864_409#_c_1398_n N_Q_c_1717_n 0.00217631f $X=10.53 $Y=1.575 $X2=0
+ $Y2=0
cc_890 N_A_1864_409#_c_1404_n N_Q_c_1717_n 0.00535008f $X=9.47 $Y=2.19 $X2=0
+ $Y2=0
cc_891 N_A_1864_409#_c_1400_n N_Q_c_1717_n 0.0198451f $X=9.77 $Y=1.55 $X2=0
+ $Y2=0
cc_892 N_A_1864_409#_c_1399_n N_VGND_c_1748_n 0.0184694f $X=9.77 $Y=0.645 $X2=0
+ $Y2=0
cc_893 N_A_1864_409#_c_1400_n N_VGND_c_1748_n 0.00144181f $X=9.77 $Y=1.55 $X2=0
+ $Y2=0
cc_894 N_A_1864_409#_M1009_g N_VGND_c_1750_n 0.00647412f $X=10.545 $Y=0.74 $X2=0
+ $Y2=0
cc_895 N_A_1864_409#_M1009_g N_VGND_c_1757_n 0.00434272f $X=10.545 $Y=0.74 $X2=0
+ $Y2=0
cc_896 N_A_1864_409#_c_1399_n N_VGND_c_1757_n 0.0145639f $X=9.77 $Y=0.645 $X2=0
+ $Y2=0
cc_897 N_A_1864_409#_M1009_g N_VGND_c_1761_n 0.00828941f $X=10.545 $Y=0.74 $X2=0
+ $Y2=0
cc_898 N_A_1864_409#_c_1399_n N_VGND_c_1761_n 0.0119984f $X=9.77 $Y=0.645 $X2=0
+ $Y2=0
cc_899 N_VPWR_M1005_d N_A_30_78#_c_1597_n 0.00501542f $X=2 $Y=1.83 $X2=0 $Y2=0
cc_900 N_VPWR_c_1454_n N_A_30_78#_c_1597_n 0.0162734f $X=2.15 $Y=2.785 $X2=0
+ $Y2=0
cc_901 N_VPWR_c_1450_n N_A_30_78#_c_1597_n 0.0237846f $X=10.8 $Y=3.33 $X2=0
+ $Y2=0
cc_902 N_VPWR_c_1452_n N_A_30_78#_c_1600_n 0.0310355f $X=0.27 $Y=2.75 $X2=0
+ $Y2=0
cc_903 N_VPWR_c_1453_n N_A_30_78#_c_1600_n 0.0222518f $X=1.17 $Y=2.815 $X2=0
+ $Y2=0
cc_904 N_VPWR_c_1463_n N_A_30_78#_c_1600_n 0.0144752f $X=1.085 $Y=3.33 $X2=0
+ $Y2=0
cc_905 N_VPWR_c_1450_n N_A_30_78#_c_1600_n 0.0119811f $X=10.8 $Y=3.33 $X2=0
+ $Y2=0
cc_906 N_VPWR_c_1453_n N_A_30_78#_c_1601_n 0.0193435f $X=1.17 $Y=2.815 $X2=0
+ $Y2=0
cc_907 N_VPWR_c_1450_n N_A_30_78#_c_1601_n 0.0125344f $X=10.8 $Y=3.33 $X2=0
+ $Y2=0
cc_908 N_VPWR_c_1450_n N_A_30_78#_c_1602_n 0.0165252f $X=10.8 $Y=3.33 $X2=0
+ $Y2=0
cc_909 N_VPWR_c_1465_n N_A_30_78#_c_1603_n 0.0053349f $X=4.385 $Y=3.33 $X2=0
+ $Y2=0
cc_910 N_VPWR_c_1450_n N_A_30_78#_c_1603_n 0.00670625f $X=10.8 $Y=3.33 $X2=0
+ $Y2=0
cc_911 N_VPWR_c_1460_n Q 0.00265735f $X=9.02 $Y=2.36 $X2=0 $Y2=0
cc_912 N_VPWR_c_1467_n Q 0.0311454f $X=10.595 $Y=3.33 $X2=0 $Y2=0
cc_913 N_VPWR_c_1450_n Q 0.0257795f $X=10.8 $Y=3.33 $X2=0 $Y2=0
cc_914 N_VPWR_c_1462_n N_Q_c_1717_n 0.045174f $X=10.76 $Y=1.985 $X2=0 $Y2=0
cc_915 N_A_30_78#_c_1590_n A_117_78# 0.00231141f $X=0.685 $Y=0.745 $X2=-0.19
+ $Y2=-0.245
cc_916 N_A_30_78#_c_1590_n N_VGND_c_1745_n 0.00719261f $X=0.685 $Y=0.745 $X2=0
+ $Y2=0
cc_917 N_A_30_78#_c_1594_n N_VGND_c_1745_n 0.00436551f $X=0.295 $Y=0.6 $X2=0
+ $Y2=0
cc_918 N_A_30_78#_c_1590_n N_VGND_c_1751_n 0.00570266f $X=0.685 $Y=0.745 $X2=0
+ $Y2=0
cc_919 N_A_30_78#_c_1594_n N_VGND_c_1751_n 0.0131067f $X=0.295 $Y=0.6 $X2=0
+ $Y2=0
cc_920 N_A_30_78#_c_1590_n N_VGND_c_1761_n 0.0111915f $X=0.685 $Y=0.745 $X2=0
+ $Y2=0
cc_921 N_A_30_78#_c_1594_n N_VGND_c_1761_n 0.0117869f $X=0.295 $Y=0.6 $X2=0
+ $Y2=0
cc_922 N_Q_c_1715_n N_VGND_c_1750_n 0.0293763f $X=10.33 $Y=0.515 $X2=0 $Y2=0
cc_923 N_Q_c_1715_n N_VGND_c_1757_n 0.0145639f $X=10.33 $Y=0.515 $X2=0 $Y2=0
cc_924 N_Q_c_1715_n N_VGND_c_1761_n 0.0119984f $X=10.33 $Y=0.515 $X2=0 $Y2=0
