* File: sky130_fd_sc_hs__a32oi_2.spice
* Created: Thu Aug 27 20:30:26 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hs__a32oi_2.pex.spice"
.subckt sky130_fd_sc_hs__a32oi_2  VNB VPB B2 B1 A1 A2 A3 Y VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* Y	Y
* A3	A3
* A2	A2
* A1	A1
* B1	B1
* B2	B2
* VPB	VPB
* VNB	VNB
MM1015 N_A_27_74#_M1015_d N_B2_M1015_g N_VGND_M1015_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.1221 PD=2.05 PS=1.07 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75001.6 A=0.111 P=1.78 MULT=1
MM1018 N_A_27_74#_M1018_d N_B2_M1018_g N_VGND_M1015_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1221 PD=1.02 PS=1.07 NRD=0 NRS=8.1 M=1 R=4.93333 SA=75000.7
+ SB=75001.1 A=0.111 P=1.78 MULT=1
MM1003 N_Y_M1003_d N_B1_M1003_g N_A_27_74#_M1018_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.1
+ SB=75000.7 A=0.111 P=1.78 MULT=1
MM1014 N_Y_M1003_d N_B1_M1014_g N_A_27_74#_M1014_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.2627 PD=1.02 PS=2.19 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75001.6
+ SB=75000.3 A=0.111 P=1.78 MULT=1
MM1012 N_Y_M1012_d N_A1_M1012_g N_A_507_74#_M1012_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.2109 PD=1.02 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75001.6 A=0.111 P=1.78 MULT=1
MM1019 N_Y_M1012_d N_A1_M1019_g N_A_507_74#_M1019_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.11285 PD=1.02 PS=1.045 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.6
+ SB=75001.2 A=0.111 P=1.78 MULT=1
MM1016 N_A_507_74#_M1019_s N_A2_M1016_g N_A_771_74#_M1016_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.11285 AS=0.14615 PD=1.045 PS=1.135 NRD=4.044 NRS=7.296 M=1
+ R=4.93333 SA=75001.1 SB=75000.8 A=0.111 P=1.78 MULT=1
MM1017 N_A_507_74#_M1017_d N_A2_M1017_g N_A_771_74#_M1016_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.2109 AS=0.14615 PD=2.05 PS=1.135 NRD=0 NRS=11.34 M=1 R=4.93333
+ SA=75001.6 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1002 N_A_771_74#_M1002_d N_A3_M1002_g N_VGND_M1002_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.2109 PD=1.02 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1013 N_A_771_74#_M1002_d N_A3_M1013_g N_VGND_M1013_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.2109 PD=1.02 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.6
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1004 N_Y_M1004_d N_B2_M1004_g N_A_27_368#_M1004_s VPB PSHORT L=0.15 W=1.12
+ AD=0.1932 AS=0.336 PD=1.465 PS=2.84 NRD=9.6727 NRS=2.6201 M=1 R=7.46667
+ SA=75000.2 SB=75005.2 A=0.168 P=2.54 MULT=1
MM1010 N_Y_M1004_d N_B2_M1010_g N_A_27_368#_M1010_s VPB PSHORT L=0.15 W=1.12
+ AD=0.1932 AS=0.196 PD=1.465 PS=1.47 NRD=1.7533 NRS=10.5395 M=1 R=7.46667
+ SA=75000.7 SB=75004.7 A=0.168 P=2.54 MULT=1
MM1007 N_A_27_368#_M1010_s N_B1_M1007_g N_Y_M1007_s VPB PSHORT L=0.15 W=1.12
+ AD=0.196 AS=0.196 PD=1.47 PS=1.47 NRD=1.7533 NRS=10.5395 M=1 R=7.46667
+ SA=75001.2 SB=75004.2 A=0.168 P=2.54 MULT=1
MM1011 N_A_27_368#_M1011_d N_B1_M1011_g N_Y_M1007_s VPB PSHORT L=0.15 W=1.12
+ AD=0.196 AS=0.196 PD=1.47 PS=1.47 NRD=10.5395 NRS=1.7533 M=1 R=7.46667
+ SA=75001.7 SB=75003.7 A=0.168 P=2.54 MULT=1
MM1000 N_A_27_368#_M1011_d N_A1_M1000_g N_VPWR_M1000_s VPB PSHORT L=0.15 W=1.12
+ AD=0.196 AS=0.3864 PD=1.47 PS=1.81 NRD=1.7533 NRS=2.6201 M=1 R=7.46667
+ SA=75002.2 SB=75003.2 A=0.168 P=2.54 MULT=1
MM1006 N_A_27_368#_M1006_d N_A1_M1006_g N_VPWR_M1000_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.3864 PD=1.42 PS=1.81 NRD=1.7533 NRS=2.6201 M=1 R=7.46667
+ SA=75003.1 SB=75002.4 A=0.168 P=2.54 MULT=1
MM1001 N_VPWR_M1001_d N_A2_M1001_g N_A_27_368#_M1006_d VPB PSHORT L=0.15 W=1.12
+ AD=0.2044 AS=0.168 PD=1.485 PS=1.42 NRD=11.426 NRS=1.7533 M=1 R=7.46667
+ SA=75003.5 SB=75001.9 A=0.168 P=2.54 MULT=1
MM1008 N_VPWR_M1001_d N_A2_M1008_g N_A_27_368#_M1008_s VPB PSHORT L=0.15 W=1.12
+ AD=0.2044 AS=0.266 PD=1.485 PS=1.595 NRD=3.5066 NRS=17.8679 M=1 R=7.46667
+ SA=75004 SB=75001.4 A=0.168 P=2.54 MULT=1
MM1005 N_VPWR_M1005_d N_A3_M1005_g N_A_27_368#_M1008_s VPB PSHORT L=0.15 W=1.12
+ AD=0.224 AS=0.266 PD=1.52 PS=1.595 NRD=10.5395 NRS=16.4101 M=1 R=7.46667
+ SA=75004.6 SB=75000.8 A=0.168 P=2.54 MULT=1
MM1009 N_VPWR_M1005_d N_A3_M1009_g N_A_27_368#_M1009_s VPB PSHORT L=0.15 W=1.12
+ AD=0.224 AS=0.3304 PD=1.52 PS=2.83 NRD=10.5395 NRS=1.7533 M=1 R=7.46667
+ SA=75005.2 SB=75000.2 A=0.168 P=2.54 MULT=1
DX20_noxref VNB VPB NWDIODE A=12.3132 P=16.96
*
.include "sky130_fd_sc_hs__a32oi_2.pxi.spice"
*
.ends
*
*
