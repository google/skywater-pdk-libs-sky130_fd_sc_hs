* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hs__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
X0 X a_83_260# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X1 a_83_260# B2 a_693_384# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=150000u
X2 a_83_260# a_233_384# a_588_74# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X3 VPWR A1_N a_233_384# VPB sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X4 a_693_384# B1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=150000u
X5 a_233_384# A2_N VPWR VPB sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X6 VPWR a_233_384# a_83_260# VPB sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X7 a_588_74# B2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X8 a_253_94# A2_N a_233_384# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X9 X a_83_260# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X10 VGND A1_N a_253_94# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X11 VGND B1 a_588_74# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
.ends
