* File: sky130_fd_sc_hs__nor3b_1.spice
* Created: Tue Sep  1 20:11:44 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hs__nor3b_1.pex.spice"
.subckt sky130_fd_sc_hs__nor3b_1  VNB VPB C_N A B VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* B	B
* A	A
* C_N	C_N
* VPB	VPB
* VNB	VNB
MM1005 N_VGND_M1005_d N_C_N_M1005_g N_A_27_112#_M1005_s VNB NLOWVT L=0.15 W=0.55
+ AD=0.116971 AS=0.2695 PD=0.963566 PS=2.08 NRD=18 NRS=0 M=1 R=3.66667
+ SA=75000.4 SB=75001.8 A=0.0825 P=1.4 MULT=1
MM1007 N_Y_M1007_d N_A_M1007_g N_VGND_M1005_d VNB NLOWVT L=0.15 W=0.74 AD=0.1184
+ AS=0.157379 PD=1.06 PS=1.29643 NRD=6.48 NRS=4.86 M=1 R=4.93333 SA=75000.8
+ SB=75001.2 A=0.111 P=1.78 MULT=1
MM1006 N_VGND_M1006_d N_B_M1006_g N_Y_M1007_d VNB NLOWVT L=0.15 W=0.74 AD=0.1554
+ AS=0.1184 PD=1.16 PS=1.06 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75001.2 SB=75000.8
+ A=0.111 P=1.78 MULT=1
MM1000 N_Y_M1000_d N_A_27_112#_M1000_g N_VGND_M1006_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.1554 PD=2.05 PS=1.16 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75001.8
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1001 N_VPWR_M1001_d N_C_N_M1001_g N_A_27_112#_M1001_s VPB PSHORT L=0.15 W=0.84
+ AD=0.1866 AS=0.2478 PD=1.32 PS=2.27 NRD=30.4759 NRS=2.3443 M=1 R=5.6
+ SA=75000.2 SB=75001.8 A=0.126 P=1.98 MULT=1
MM1002 A_260_368# N_A_M1002_g N_VPWR_M1001_d VPB PSHORT L=0.15 W=1.12 AD=0.1512
+ AS=0.2488 PD=1.39 PS=1.76 NRD=14.0658 NRS=1.7533 M=1 R=7.46667 SA=75000.6
+ SB=75001.2 A=0.168 P=2.54 MULT=1
MM1004 A_344_368# N_B_M1004_g A_260_368# VPB PSHORT L=0.15 W=1.12 AD=0.2352
+ AS=0.1512 PD=1.54 PS=1.39 NRD=27.2451 NRS=14.0658 M=1 R=7.46667 SA=75001.1
+ SB=75000.8 A=0.168 P=2.54 MULT=1
MM1003 N_Y_M1003_d N_A_27_112#_M1003_g A_344_368# VPB PSHORT L=0.15 W=1.12
+ AD=0.3304 AS=0.2352 PD=2.83 PS=1.54 NRD=1.7533 NRS=27.2451 M=1 R=7.46667
+ SA=75001.6 SB=75000.2 A=0.168 P=2.54 MULT=1
DX8_noxref VNB VPB NWDIODE A=6.0636 P=10.24
*
.include "sky130_fd_sc_hs__nor3b_1.pxi.spice"
*
.ends
*
*
