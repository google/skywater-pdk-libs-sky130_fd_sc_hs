* File: sky130_fd_sc_hs__a31oi_1.spice
* Created: Tue Sep  1 19:53:07 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hs__a31oi_1.pex.spice"
.subckt sky130_fd_sc_hs__a31oi_1  VNB VPB A3 A2 A1 B1 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* B1	B1
* A1	A1
* A2	A2
* A3	A3
* VPB	VPB
* VNB	VNB
MM1007 A_145_74# N_A3_M1007_g N_VGND_M1007_s VNB NLOWVT L=0.15 W=0.74 AD=0.0888
+ AS=0.3182 PD=0.98 PS=2.34 NRD=10.536 NRS=23.508 M=1 R=4.93333 SA=75000.4
+ SB=75001.7 A=0.111 P=1.78 MULT=1
MM1005 A_223_74# N_A2_M1005_g A_145_74# VNB NLOWVT L=0.15 W=0.74 AD=0.1554
+ AS=0.0888 PD=1.16 PS=0.98 NRD=25.128 NRS=10.536 M=1 R=4.93333 SA=75000.7
+ SB=75001.4 A=0.111 P=1.78 MULT=1
MM1001 N_Y_M1001_d N_A1_M1001_g A_223_74# VNB NLOWVT L=0.15 W=0.74 AD=0.1554
+ AS=0.1554 PD=1.16 PS=1.16 NRD=11.34 NRS=25.128 M=1 R=4.93333 SA=75001.3
+ SB=75000.8 A=0.111 P=1.78 MULT=1
MM1006 N_VGND_M1006_d N_B1_M1006_g N_Y_M1001_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.1554 PD=2.05 PS=1.16 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75001.9
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1000 N_A_136_368#_M1000_d N_A3_M1000_g N_VPWR_M1000_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.4312 PD=1.42 PS=3.01 NRD=1.7533 NRS=17.5724 M=1 R=7.46667
+ SA=75000.3 SB=75001.8 A=0.168 P=2.54 MULT=1
MM1002 N_VPWR_M1002_d N_A2_M1002_g N_A_136_368#_M1000_d VPB PSHORT L=0.15 W=1.12
+ AD=0.2744 AS=0.168 PD=1.61 PS=1.42 NRD=17.5724 NRS=1.7533 M=1 R=7.46667
+ SA=75000.8 SB=75001.4 A=0.168 P=2.54 MULT=1
MM1004 N_A_136_368#_M1004_d N_A1_M1004_g N_VPWR_M1002_d VPB PSHORT L=0.15 W=1.12
+ AD=0.196 AS=0.2744 PD=1.47 PS=1.61 NRD=1.7533 NRS=19.3454 M=1 R=7.46667
+ SA=75001.4 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1003 N_Y_M1003_d N_B1_M1003_g N_A_136_368#_M1004_d VPB PSHORT L=0.15 W=1.12
+ AD=0.3304 AS=0.196 PD=2.83 PS=1.47 NRD=1.7533 NRS=10.5395 M=1 R=7.46667
+ SA=75001.9 SB=75000.2 A=0.168 P=2.54 MULT=1
DX8_noxref VNB VPB NWDIODE A=6.0636 P=10.24
*
.include "sky130_fd_sc_hs__a31oi_1.pxi.spice"
*
.ends
*
*
