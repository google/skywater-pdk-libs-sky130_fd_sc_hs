* File: sky130_fd_sc_hs__dlclkp_2.pxi.spice
* Created: Thu Aug 27 20:40:37 2020
* 
x_PM_SKY130_FD_SC_HS__DLCLKP_2%A_83_244# N_A_83_244#_M1013_d N_A_83_244#_M1004_d
+ N_A_83_244#_c_139_n N_A_83_244#_M1020_g N_A_83_244#_c_140_n
+ N_A_83_244#_M1012_g N_A_83_244#_c_141_n N_A_83_244#_c_142_n
+ N_A_83_244#_c_147_n N_A_83_244#_c_206_p N_A_83_244#_c_143_n
+ N_A_83_244#_c_164_p N_A_83_244#_c_194_p N_A_83_244#_c_163_p
+ N_A_83_244#_c_181_p N_A_83_244#_c_165_p N_A_83_244#_c_144_n
+ PM_SKY130_FD_SC_HS__DLCLKP_2%A_83_244#
x_PM_SKY130_FD_SC_HS__DLCLKP_2%GATE N_GATE_c_224_n N_GATE_M1000_g N_GATE_M1014_g
+ GATE PM_SKY130_FD_SC_HS__DLCLKP_2%GATE
x_PM_SKY130_FD_SC_HS__DLCLKP_2%A_315_48# N_A_315_48#_M1015_s N_A_315_48#_M1002_s
+ N_A_315_48#_c_259_n N_A_315_48#_M1013_g N_A_315_48#_c_273_n
+ N_A_315_48#_M1007_g N_A_315_48#_c_260_n N_A_315_48#_M1016_g
+ N_A_315_48#_M1011_g N_A_315_48#_c_262_n N_A_315_48#_c_263_n
+ N_A_315_48#_c_264_n N_A_315_48#_c_277_n N_A_315_48#_c_278_n
+ N_A_315_48#_c_279_n N_A_315_48#_c_265_n N_A_315_48#_c_266_n
+ N_A_315_48#_c_267_n N_A_315_48#_c_280_n N_A_315_48#_c_281_n
+ N_A_315_48#_c_268_n N_A_315_48#_c_269_n N_A_315_48#_c_270_n
+ N_A_315_48#_c_271_n N_A_315_48#_c_284_n N_A_315_48#_c_285_n
+ N_A_315_48#_c_272_n PM_SKY130_FD_SC_HS__DLCLKP_2%A_315_48#
x_PM_SKY130_FD_SC_HS__DLCLKP_2%A_315_338# N_A_315_338#_M1011_d
+ N_A_315_338#_M1016_d N_A_315_338#_c_415_n N_A_315_338#_M1004_g
+ N_A_315_338#_c_405_n N_A_315_338#_c_406_n N_A_315_338#_M1006_g
+ N_A_315_338#_c_408_n N_A_315_338#_c_409_n N_A_315_338#_c_410_n
+ N_A_315_338#_c_411_n N_A_315_338#_c_420_n N_A_315_338#_c_412_n
+ N_A_315_338#_c_413_n N_A_315_338#_c_414_n
+ PM_SKY130_FD_SC_HS__DLCLKP_2%A_315_338#
x_PM_SKY130_FD_SC_HS__DLCLKP_2%CLK N_CLK_c_507_n N_CLK_c_508_n N_CLK_M1002_g
+ N_CLK_c_503_n N_CLK_M1015_g N_CLK_c_509_n N_CLK_M1017_g N_CLK_c_504_n
+ N_CLK_M1019_g CLK N_CLK_c_506_n PM_SKY130_FD_SC_HS__DLCLKP_2%CLK
x_PM_SKY130_FD_SC_HS__DLCLKP_2%A_27_74# N_A_27_74#_M1020_s N_A_27_74#_M1012_s
+ N_A_27_74#_M1010_g N_A_27_74#_c_566_n N_A_27_74#_c_567_n N_A_27_74#_c_568_n
+ N_A_27_74#_M1021_g N_A_27_74#_c_554_n N_A_27_74#_M1018_g N_A_27_74#_c_556_n
+ N_A_27_74#_c_570_n N_A_27_74#_M1009_g N_A_27_74#_c_557_n N_A_27_74#_c_558_n
+ N_A_27_74#_c_571_n N_A_27_74#_c_577_n N_A_27_74#_c_581_n N_A_27_74#_c_559_n
+ N_A_27_74#_c_560_n N_A_27_74#_c_561_n N_A_27_74#_c_572_n N_A_27_74#_c_562_n
+ N_A_27_74#_c_563_n N_A_27_74#_c_564_n PM_SKY130_FD_SC_HS__DLCLKP_2%A_27_74#
x_PM_SKY130_FD_SC_HS__DLCLKP_2%A_1041_387# N_A_1041_387#_M1018_d
+ N_A_1041_387#_M1017_d N_A_1041_387#_c_685_n N_A_1041_387#_c_686_n
+ N_A_1041_387#_c_687_n N_A_1041_387#_M1003_g N_A_1041_387#_M1001_g
+ N_A_1041_387#_c_689_n N_A_1041_387#_c_690_n N_A_1041_387#_M1005_g
+ N_A_1041_387#_c_691_n N_A_1041_387#_M1008_g N_A_1041_387#_c_698_n
+ N_A_1041_387#_c_692_n N_A_1041_387#_c_711_n N_A_1041_387#_c_693_n
+ N_A_1041_387#_c_694_n N_A_1041_387#_c_695_n
+ PM_SKY130_FD_SC_HS__DLCLKP_2%A_1041_387#
x_PM_SKY130_FD_SC_HS__DLCLKP_2%VPWR N_VPWR_M1012_d N_VPWR_M1021_d N_VPWR_M1002_d
+ N_VPWR_M1009_d N_VPWR_M1005_s N_VPWR_c_750_n N_VPWR_c_751_n N_VPWR_c_752_n
+ N_VPWR_c_753_n N_VPWR_c_754_n N_VPWR_c_755_n N_VPWR_c_756_n N_VPWR_c_757_n
+ VPWR N_VPWR_c_758_n N_VPWR_c_759_n N_VPWR_c_760_n N_VPWR_c_761_n
+ N_VPWR_c_762_n N_VPWR_c_763_n N_VPWR_c_749_n PM_SKY130_FD_SC_HS__DLCLKP_2%VPWR
x_PM_SKY130_FD_SC_HS__DLCLKP_2%GCLK N_GCLK_M1001_d N_GCLK_M1003_d GCLK GCLK GCLK
+ GCLK GCLK GCLK GCLK PM_SKY130_FD_SC_HS__DLCLKP_2%GCLK
x_PM_SKY130_FD_SC_HS__DLCLKP_2%VGND N_VGND_M1020_d N_VGND_M1010_d N_VGND_M1015_d
+ N_VGND_M1001_s N_VGND_M1008_s N_VGND_c_849_n N_VGND_c_867_n N_VGND_c_850_n
+ N_VGND_c_851_n N_VGND_c_852_n N_VGND_c_853_n N_VGND_c_854_n N_VGND_c_855_n
+ N_VGND_c_856_n VGND N_VGND_c_857_n N_VGND_c_858_n N_VGND_c_859_n
+ N_VGND_c_860_n N_VGND_c_861_n N_VGND_c_862_n N_VGND_c_863_n N_VGND_c_864_n
+ PM_SKY130_FD_SC_HS__DLCLKP_2%VGND
cc_1 VNB N_A_83_244#_c_139_n 0.0220218f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.22
cc_2 VNB N_A_83_244#_c_140_n 0.0431823f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.765
cc_3 VNB N_A_83_244#_c_141_n 0.00153124f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=1.95
cc_4 VNB N_A_83_244#_c_142_n 0.0152926f $X=-0.19 $Y=-0.245 $X2=1.39 $Y2=1.195
cc_5 VNB N_A_83_244#_c_143_n 0.00177418f $X=-0.19 $Y=-0.245 $X2=1.475 $Y2=1.11
cc_6 VNB N_A_83_244#_c_144_n 0.00400117f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.195
cc_7 VNB N_GATE_c_224_n 0.0282691f $X=-0.19 $Y=-0.245 $X2=1.725 $Y2=0.37
cc_8 VNB N_GATE_M1014_g 0.0359138f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB GATE 0.00166024f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_10 VNB N_A_315_48#_c_259_n 0.0194382f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.22
cc_11 VNB N_A_315_48#_c_260_n 0.0100498f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=1.55
cc_12 VNB N_A_315_48#_M1011_g 0.0270544f $X=-0.19 $Y=-0.245 $X2=0.785 $Y2=2.035
cc_13 VNB N_A_315_48#_c_262_n 0.0179051f $X=-0.19 $Y=-0.245 $X2=1.475 $Y2=1.11
cc_14 VNB N_A_315_48#_c_263_n 0.0220269f $X=-0.19 $Y=-0.245 $X2=1.985 $Y2=0.785
cc_15 VNB N_A_315_48#_c_264_n 0.00427785f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_315_48#_c_265_n 0.00821628f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=1.385
cc_17 VNB N_A_315_48#_c_266_n 0.00450361f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_315_48#_c_267_n 0.0444201f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_315_48#_c_268_n 0.00306113f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_315_48#_c_269_n 0.00809643f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_315_48#_c_270_n 0.00466113f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_315_48#_c_271_n 0.00191868f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_315_48#_c_272_n 0.0209823f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_315_338#_c_405_n 0.0186275f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.765
cc_25 VNB N_A_315_338#_c_406_n 0.00664977f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_26 VNB N_A_315_338#_M1006_g 0.0386613f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=1.95
cc_27 VNB N_A_315_338#_c_408_n 0.00235348f $X=-0.19 $Y=-0.245 $X2=0.785
+ $Y2=2.035
cc_28 VNB N_A_315_338#_c_409_n 0.0235511f $X=-0.19 $Y=-0.245 $X2=1.475 $Y2=0.95
cc_29 VNB N_A_315_338#_c_410_n 0.0217428f $X=-0.19 $Y=-0.245 $X2=1.62 $Y2=2.12
cc_30 VNB N_A_315_338#_c_411_n 0.00831277f $X=-0.19 $Y=-0.245 $X2=1.62 $Y2=2.55
cc_31 VNB N_A_315_338#_c_412_n 0.00764425f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.195
cc_32 VNB N_A_315_338#_c_413_n 0.00361802f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.385
cc_33 VNB N_A_315_338#_c_414_n 0.00241587f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=1.385
cc_34 VNB N_CLK_c_503_n 0.0193105f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_CLK_c_504_n 0.0143329f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_36 VNB CLK 0.00198218f $X=-0.19 $Y=-0.245 $X2=1.39 $Y2=1.195
cc_37 VNB N_CLK_c_506_n 0.0376276f $X=-0.19 $Y=-0.245 $X2=1.62 $Y2=2.55
cc_38 VNB N_A_27_74#_M1010_g 0.0450427f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.765
cc_39 VNB N_A_27_74#_c_554_n 0.181798f $X=-0.19 $Y=-0.245 $X2=0.785 $Y2=1.195
cc_40 VNB N_A_27_74#_M1018_g 0.0314802f $X=-0.19 $Y=-0.245 $X2=1.62 $Y2=2.12
cc_41 VNB N_A_27_74#_c_556_n 0.0139968f $X=-0.19 $Y=-0.245 $X2=1.56 $Y2=0.785
cc_42 VNB N_A_27_74#_c_557_n 0.0134447f $X=-0.19 $Y=-0.245 $X2=2.24 $Y2=2.715
cc_43 VNB N_A_27_74#_c_558_n 0.0184195f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_27_74#_c_559_n 0.0311942f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_A_27_74#_c_560_n 0.00181663f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_A_27_74#_c_561_n 0.00717518f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_27_74#_c_562_n 0.0319566f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_27_74#_c_563_n 0.00198487f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A_27_74#_c_564_n 0.0598204f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_A_1041_387#_c_685_n 0.0235679f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.22
cc_51 VNB N_A_1041_387#_c_686_n 0.0213858f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_52 VNB N_A_1041_387#_c_687_n 0.00939179f $X=-0.19 $Y=-0.245 $X2=0.495
+ $Y2=0.74
cc_53 VNB N_A_1041_387#_M1001_g 0.01958f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=1.95
cc_54 VNB N_A_1041_387#_c_689_n 0.0165324f $X=-0.19 $Y=-0.245 $X2=0.785
+ $Y2=1.195
cc_55 VNB N_A_1041_387#_c_690_n 0.0267295f $X=-0.19 $Y=-0.245 $X2=0.785
+ $Y2=2.035
cc_56 VNB N_A_1041_387#_c_691_n 0.018904f $X=-0.19 $Y=-0.245 $X2=1.62 $Y2=2.12
cc_57 VNB N_A_1041_387#_c_692_n 0.0128974f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=1.385
cc_58 VNB N_A_1041_387#_c_693_n 0.0011398f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_A_1041_387#_c_694_n 0.0152157f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_A_1041_387#_c_695_n 0.04777f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_VPWR_c_749_n 0.322901f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB GCLK 0.00279061f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.22
cc_63 VNB N_VGND_c_849_n 0.00624343f $X=-0.19 $Y=-0.245 $X2=0.785 $Y2=2.035
cc_64 VNB N_VGND_c_850_n 0.0138044f $X=-0.19 $Y=-0.245 $X2=1.985 $Y2=0.785
cc_65 VNB N_VGND_c_851_n 0.0127026f $X=-0.19 $Y=-0.245 $X2=2.24 $Y2=2.715
cc_66 VNB N_VGND_c_852_n 0.0322141f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_VGND_c_853_n 0.010678f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=1.385
cc_68 VNB N_VGND_c_854_n 0.0517326f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.55
cc_69 VNB N_VGND_c_855_n 0.0562641f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_VGND_c_856_n 0.0025968f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_VGND_c_857_n 0.0172347f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_VGND_c_858_n 0.0335133f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_VGND_c_859_n 0.0357493f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_VGND_c_860_n 0.0194281f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_VGND_c_861_n 0.00622845f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_VGND_c_862_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_VGND_c_863_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_VGND_c_864_n 0.41597f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VPB N_A_83_244#_c_140_n 0.0303696f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.765
cc_80 VPB N_A_83_244#_c_141_n 0.00350692f $X=-0.19 $Y=1.66 $X2=0.7 $Y2=1.95
cc_81 VPB N_A_83_244#_c_147_n 0.00768499f $X=-0.19 $Y=1.66 $X2=1.535 $Y2=2.035
cc_82 VPB N_GATE_c_224_n 0.0342485f $X=-0.19 $Y=1.66 $X2=1.725 $Y2=0.37
cc_83 VPB GATE 0.00138199f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.74
cc_84 VPB N_A_315_48#_c_273_n 0.0559614f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.765
cc_85 VPB N_A_315_48#_c_260_n 0.0371568f $X=-0.19 $Y=1.66 $X2=0.7 $Y2=1.55
cc_86 VPB N_A_315_48#_c_263_n 0.0160353f $X=-0.19 $Y=1.66 $X2=1.985 $Y2=0.785
cc_87 VPB N_A_315_48#_c_264_n 0.00830448f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_88 VPB N_A_315_48#_c_277_n 7.40136e-19 $X=-0.19 $Y=1.66 $X2=2.24 $Y2=2.715
cc_89 VPB N_A_315_48#_c_278_n 0.0204424f $X=-0.19 $Y=1.66 $X2=2.24 $Y2=2.715
cc_90 VPB N_A_315_48#_c_279_n 0.00281294f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_91 VPB N_A_315_48#_c_280_n 0.0038784f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_92 VPB N_A_315_48#_c_281_n 0.00348569f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_93 VPB N_A_315_48#_c_268_n 0.00593009f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_94 VPB N_A_315_48#_c_269_n 0.00924015f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_95 VPB N_A_315_48#_c_284_n 0.0181262f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_96 VPB N_A_315_48#_c_285_n 0.00337784f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_97 VPB N_A_315_48#_c_272_n 0.0161977f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_98 VPB N_A_315_338#_c_415_n 0.0176083f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.22
cc_99 VPB N_A_315_338#_c_405_n 0.0182164f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.765
cc_100 VPB N_A_315_338#_c_406_n 0.00571473f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.4
cc_101 VPB N_A_315_338#_c_408_n 0.00229055f $X=-0.19 $Y=1.66 $X2=0.785 $Y2=2.035
cc_102 VPB N_A_315_338#_c_409_n 0.00699468f $X=-0.19 $Y=1.66 $X2=1.475 $Y2=0.95
cc_103 VPB N_A_315_338#_c_420_n 0.0130417f $X=-0.19 $Y=1.66 $X2=1.705 $Y2=2.715
cc_104 VPB N_A_315_338#_c_414_n 0.0037762f $X=-0.19 $Y=1.66 $X2=0.6 $Y2=1.385
cc_105 VPB N_CLK_c_507_n 0.00861795f $X=-0.19 $Y=1.66 $X2=1.74 $Y2=1.96
cc_106 VPB N_CLK_c_508_n 0.0261208f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_107 VPB N_CLK_c_509_n 0.0154607f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.74
cc_108 VPB CLK 0.00387263f $X=-0.19 $Y=1.66 $X2=1.39 $Y2=1.195
cc_109 VPB N_CLK_c_506_n 0.0177503f $X=-0.19 $Y=1.66 $X2=1.62 $Y2=2.55
cc_110 VPB N_A_27_74#_M1010_g 0.0249593f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.765
cc_111 VPB N_A_27_74#_c_566_n 0.00552919f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.4
cc_112 VPB N_A_27_74#_c_567_n 0.0100286f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.4
cc_113 VPB N_A_27_74#_c_568_n 0.0236416f $X=-0.19 $Y=1.66 $X2=0.7 $Y2=1.55
cc_114 VPB N_A_27_74#_c_556_n 0.00113446f $X=-0.19 $Y=1.66 $X2=1.56 $Y2=0.785
cc_115 VPB N_A_27_74#_c_570_n 0.0256225f $X=-0.19 $Y=1.66 $X2=1.985 $Y2=0.785
cc_116 VPB N_A_27_74#_c_571_n 0.0413071f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_117 VPB N_A_27_74#_c_572_n 0.0131772f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_118 VPB N_A_27_74#_c_562_n 0.00751948f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_119 VPB N_A_1041_387#_c_687_n 0.0281292f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.74
cc_120 VPB N_A_1041_387#_c_690_n 0.0270667f $X=-0.19 $Y=1.66 $X2=0.785 $Y2=2.035
cc_121 VPB N_A_1041_387#_c_698_n 0.00301826f $X=-0.19 $Y=1.66 $X2=2.24 $Y2=2.715
cc_122 VPB N_A_1041_387#_c_693_n 0.00164874f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_123 VPB N_VPWR_c_750_n 0.0106565f $X=-0.19 $Y=1.66 $X2=1.475 $Y2=1.11
cc_124 VPB N_VPWR_c_751_n 0.00880467f $X=-0.19 $Y=1.66 $X2=1.985 $Y2=0.785
cc_125 VPB N_VPWR_c_752_n 0.0124551f $X=-0.19 $Y=1.66 $X2=2.24 $Y2=2.715
cc_126 VPB N_VPWR_c_753_n 0.0174362f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_127 VPB N_VPWR_c_754_n 0.0106521f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=1.55
cc_128 VPB N_VPWR_c_755_n 0.058526f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_129 VPB N_VPWR_c_756_n 0.0340382f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_130 VPB N_VPWR_c_757_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_131 VPB N_VPWR_c_758_n 0.05371f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_132 VPB N_VPWR_c_759_n 0.0191831f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_133 VPB N_VPWR_c_760_n 0.019013f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_134 VPB N_VPWR_c_761_n 0.0286985f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_135 VPB N_VPWR_c_762_n 0.0101806f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_136 VPB N_VPWR_c_763_n 0.0173816f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_137 VPB N_VPWR_c_749_n 0.116558f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_138 VPB GCLK 0.00343907f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.22
cc_139 N_A_83_244#_c_140_n N_GATE_c_224_n 0.0278162f $X=0.505 $Y=1.765 $X2=-0.19
+ $Y2=-0.245
cc_140 N_A_83_244#_c_141_n N_GATE_c_224_n 0.00310124f $X=0.7 $Y=1.95 $X2=-0.19
+ $Y2=-0.245
cc_141 N_A_83_244#_c_142_n N_GATE_c_224_n 0.00125994f $X=1.39 $Y=1.195 $X2=-0.19
+ $Y2=-0.245
cc_142 N_A_83_244#_c_147_n N_GATE_c_224_n 0.0179878f $X=1.535 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_143 N_A_83_244#_c_144_n N_GATE_c_224_n 0.00235935f $X=0.61 $Y=1.195 $X2=-0.19
+ $Y2=-0.245
cc_144 N_A_83_244#_c_139_n N_GATE_M1014_g 0.012465f $X=0.495 $Y=1.22 $X2=0 $Y2=0
cc_145 N_A_83_244#_c_140_n N_GATE_M1014_g 0.00568186f $X=0.505 $Y=1.765 $X2=0
+ $Y2=0
cc_146 N_A_83_244#_c_142_n N_GATE_M1014_g 0.0140883f $X=1.39 $Y=1.195 $X2=0
+ $Y2=0
cc_147 N_A_83_244#_c_143_n N_GATE_M1014_g 0.00251346f $X=1.475 $Y=1.11 $X2=0
+ $Y2=0
cc_148 N_A_83_244#_c_144_n N_GATE_M1014_g 0.00341679f $X=0.61 $Y=1.195 $X2=0
+ $Y2=0
cc_149 N_A_83_244#_c_142_n GATE 0.0242156f $X=1.39 $Y=1.195 $X2=0 $Y2=0
cc_150 N_A_83_244#_c_147_n GATE 0.0242115f $X=1.535 $Y=2.035 $X2=0 $Y2=0
cc_151 N_A_83_244#_c_144_n GATE 0.020776f $X=0.61 $Y=1.195 $X2=0 $Y2=0
cc_152 N_A_83_244#_c_142_n N_A_315_48#_c_259_n 0.00182637f $X=1.39 $Y=1.195
+ $X2=0 $Y2=0
cc_153 N_A_83_244#_c_143_n N_A_315_48#_c_259_n 0.00265217f $X=1.475 $Y=1.11
+ $X2=0 $Y2=0
cc_154 N_A_83_244#_c_163_p N_A_315_48#_c_259_n 0.0220272f $X=1.985 $Y=0.785
+ $X2=0 $Y2=0
cc_155 N_A_83_244#_c_164_p N_A_315_48#_c_273_n 0.00101661f $X=1.62 $Y=2.55 $X2=0
+ $Y2=0
cc_156 N_A_83_244#_c_165_p N_A_315_48#_c_273_n 0.00945707f $X=2.24 $Y=2.715
+ $X2=0 $Y2=0
cc_157 N_A_83_244#_M1004_d N_A_315_48#_c_264_n 9.27736e-19 $X=1.74 $Y=1.96 $X2=0
+ $Y2=0
cc_158 N_A_83_244#_c_147_n N_A_315_48#_c_264_n 0.00783655f $X=1.535 $Y=2.035
+ $X2=0 $Y2=0
cc_159 N_A_83_244#_M1004_d N_A_315_48#_c_277_n 0.00454028f $X=1.74 $Y=1.96 $X2=0
+ $Y2=0
cc_160 N_A_83_244#_c_147_n N_A_315_48#_c_277_n 0.00611828f $X=1.535 $Y=2.035
+ $X2=0 $Y2=0
cc_161 N_A_83_244#_c_164_p N_A_315_48#_c_277_n 0.00785901f $X=1.62 $Y=2.55 $X2=0
+ $Y2=0
cc_162 N_A_83_244#_c_165_p N_A_315_48#_c_277_n 0.00892168f $X=2.24 $Y=2.715
+ $X2=0 $Y2=0
cc_163 N_A_83_244#_c_142_n N_A_315_48#_c_266_n 0.0134482f $X=1.39 $Y=1.195 $X2=0
+ $Y2=0
cc_164 N_A_83_244#_c_163_p N_A_315_48#_c_266_n 0.0231063f $X=1.985 $Y=0.785
+ $X2=0 $Y2=0
cc_165 N_A_83_244#_c_147_n N_A_315_48#_c_267_n 5.1943e-19 $X=1.535 $Y=2.035
+ $X2=0 $Y2=0
cc_166 N_A_83_244#_c_163_p N_A_315_48#_c_267_n 0.00218947f $X=1.985 $Y=0.785
+ $X2=0 $Y2=0
cc_167 N_A_83_244#_c_165_p N_A_315_48#_c_280_n 0.00866848f $X=2.24 $Y=2.715
+ $X2=0 $Y2=0
cc_168 N_A_83_244#_c_164_p N_A_315_48#_c_281_n 0.00456122f $X=1.62 $Y=2.55 $X2=0
+ $Y2=0
cc_169 N_A_83_244#_c_165_p N_A_315_48#_c_281_n 0.0116105f $X=2.24 $Y=2.715 $X2=0
+ $Y2=0
cc_170 N_A_83_244#_c_147_n N_A_315_338#_c_415_n 0.00700798f $X=1.535 $Y=2.035
+ $X2=0 $Y2=0
cc_171 N_A_83_244#_c_164_p N_A_315_338#_c_415_n 0.0122485f $X=1.62 $Y=2.55 $X2=0
+ $Y2=0
cc_172 N_A_83_244#_c_181_p N_A_315_338#_c_415_n 0.00671935f $X=1.705 $Y=2.715
+ $X2=0 $Y2=0
cc_173 N_A_83_244#_c_165_p N_A_315_338#_c_415_n 0.00307308f $X=2.24 $Y=2.715
+ $X2=0 $Y2=0
cc_174 N_A_83_244#_c_147_n N_A_315_338#_c_406_n 7.08935e-19 $X=1.535 $Y=2.035
+ $X2=0 $Y2=0
cc_175 N_A_83_244#_c_163_p N_A_315_338#_M1006_g 0.00839955f $X=1.985 $Y=0.785
+ $X2=0 $Y2=0
cc_176 N_A_83_244#_c_165_p N_A_27_74#_c_568_n 0.00112965f $X=2.24 $Y=2.715 $X2=0
+ $Y2=0
cc_177 N_A_83_244#_c_139_n N_A_27_74#_c_558_n 0.00197738f $X=0.495 $Y=1.22 $X2=0
+ $Y2=0
cc_178 N_A_83_244#_c_140_n N_A_27_74#_c_571_n 0.018212f $X=0.505 $Y=1.765 $X2=0
+ $Y2=0
cc_179 N_A_83_244#_c_139_n N_A_27_74#_c_577_n 0.0132268f $X=0.495 $Y=1.22 $X2=0
+ $Y2=0
cc_180 N_A_83_244#_c_140_n N_A_27_74#_c_577_n 9.35735e-19 $X=0.505 $Y=1.765
+ $X2=0 $Y2=0
cc_181 N_A_83_244#_c_142_n N_A_27_74#_c_577_n 0.0308414f $X=1.39 $Y=1.195 $X2=0
+ $Y2=0
cc_182 N_A_83_244#_c_144_n N_A_27_74#_c_577_n 0.0250509f $X=0.61 $Y=1.195 $X2=0
+ $Y2=0
cc_183 N_A_83_244#_c_139_n N_A_27_74#_c_581_n 0.00234284f $X=0.495 $Y=1.22 $X2=0
+ $Y2=0
cc_184 N_A_83_244#_M1013_d N_A_27_74#_c_559_n 0.00224052f $X=1.725 $Y=0.37 $X2=0
+ $Y2=0
cc_185 N_A_83_244#_c_194_p N_A_27_74#_c_559_n 0.00850309f $X=1.56 $Y=0.785 $X2=0
+ $Y2=0
cc_186 N_A_83_244#_c_163_p N_A_27_74#_c_559_n 0.0387841f $X=1.985 $Y=0.785 $X2=0
+ $Y2=0
cc_187 N_A_83_244#_c_139_n N_A_27_74#_c_560_n 3.77494e-19 $X=0.495 $Y=1.22 $X2=0
+ $Y2=0
cc_188 N_A_83_244#_c_140_n N_A_27_74#_c_572_n 0.00341081f $X=0.505 $Y=1.765
+ $X2=0 $Y2=0
cc_189 N_A_83_244#_c_141_n N_A_27_74#_c_572_n 0.00563688f $X=0.7 $Y=1.95 $X2=0
+ $Y2=0
cc_190 N_A_83_244#_c_144_n N_A_27_74#_c_572_n 4.51339e-19 $X=0.61 $Y=1.195 $X2=0
+ $Y2=0
cc_191 N_A_83_244#_c_139_n N_A_27_74#_c_562_n 0.00629621f $X=0.495 $Y=1.22 $X2=0
+ $Y2=0
cc_192 N_A_83_244#_c_140_n N_A_27_74#_c_562_n 0.0125629f $X=0.505 $Y=1.765 $X2=0
+ $Y2=0
cc_193 N_A_83_244#_c_141_n N_A_27_74#_c_562_n 0.00999482f $X=0.7 $Y=1.95 $X2=0
+ $Y2=0
cc_194 N_A_83_244#_c_144_n N_A_27_74#_c_562_n 0.0331796f $X=0.61 $Y=1.195 $X2=0
+ $Y2=0
cc_195 N_A_83_244#_c_141_n N_VPWR_M1012_d 0.00239213f $X=0.7 $Y=1.95 $X2=-0.19
+ $Y2=-0.245
cc_196 N_A_83_244#_c_147_n N_VPWR_M1012_d 0.00754708f $X=1.535 $Y=2.035
+ $X2=-0.19 $Y2=-0.245
cc_197 N_A_83_244#_c_206_p N_VPWR_M1012_d 0.00468752f $X=0.785 $Y=2.035
+ $X2=-0.19 $Y2=-0.245
cc_198 N_A_83_244#_c_140_n N_VPWR_c_750_n 0.0109702f $X=0.505 $Y=1.765 $X2=0
+ $Y2=0
cc_199 N_A_83_244#_c_147_n N_VPWR_c_750_n 0.0234761f $X=1.535 $Y=2.035 $X2=0
+ $Y2=0
cc_200 N_A_83_244#_c_206_p N_VPWR_c_750_n 0.00888093f $X=0.785 $Y=2.035 $X2=0
+ $Y2=0
cc_201 N_A_83_244#_c_165_p N_VPWR_c_751_n 0.00732265f $X=2.24 $Y=2.715 $X2=0
+ $Y2=0
cc_202 N_A_83_244#_c_181_p N_VPWR_c_758_n 0.00425285f $X=1.705 $Y=2.715 $X2=0
+ $Y2=0
cc_203 N_A_83_244#_c_165_p N_VPWR_c_758_n 0.0188311f $X=2.24 $Y=2.715 $X2=0
+ $Y2=0
cc_204 N_A_83_244#_c_140_n N_VPWR_c_761_n 0.00445602f $X=0.505 $Y=1.765 $X2=0
+ $Y2=0
cc_205 N_A_83_244#_c_140_n N_VPWR_c_749_n 0.00863959f $X=0.505 $Y=1.765 $X2=0
+ $Y2=0
cc_206 N_A_83_244#_c_181_p N_VPWR_c_749_n 0.00531278f $X=1.705 $Y=2.715 $X2=0
+ $Y2=0
cc_207 N_A_83_244#_c_165_p N_VPWR_c_749_n 0.02329f $X=2.24 $Y=2.715 $X2=0 $Y2=0
cc_208 N_A_83_244#_c_147_n A_264_392# 0.00595227f $X=1.535 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_209 N_A_83_244#_c_144_n N_VGND_M1020_d 0.00236742f $X=0.61 $Y=1.195 $X2=-0.19
+ $Y2=-0.245
cc_210 N_A_83_244#_c_139_n N_VGND_c_849_n 0.0103149f $X=0.495 $Y=1.22 $X2=0
+ $Y2=0
cc_211 N_A_83_244#_c_163_p N_VGND_c_867_n 0.00553878f $X=1.985 $Y=0.785 $X2=0
+ $Y2=0
cc_212 N_A_83_244#_c_139_n N_VGND_c_857_n 0.00383152f $X=0.495 $Y=1.22 $X2=0
+ $Y2=0
cc_213 N_A_83_244#_c_139_n N_VGND_c_864_n 0.00372928f $X=0.495 $Y=1.22 $X2=0
+ $Y2=0
cc_214 N_A_83_244#_c_194_p A_267_74# 0.00141515f $X=1.56 $Y=0.785 $X2=-0.19
+ $Y2=-0.245
cc_215 N_GATE_M1014_g N_A_315_48#_c_259_n 0.0626206f $X=1.26 $Y=0.69 $X2=0 $Y2=0
cc_216 N_GATE_c_224_n N_A_315_48#_c_264_n 0.00449067f $X=1.245 $Y=1.885 $X2=0
+ $Y2=0
cc_217 GATE N_A_315_48#_c_264_n 0.0100164f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_218 N_GATE_M1014_g N_A_315_48#_c_266_n 9.06551e-19 $X=1.26 $Y=0.69 $X2=0
+ $Y2=0
cc_219 N_GATE_c_224_n N_A_315_338#_c_415_n 0.0539653f $X=1.245 $Y=1.885 $X2=0
+ $Y2=0
cc_220 N_GATE_c_224_n N_A_315_338#_c_406_n 0.0116062f $X=1.245 $Y=1.885 $X2=0
+ $Y2=0
cc_221 GATE N_A_315_338#_c_406_n 4.43419e-19 $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_222 N_GATE_M1014_g N_A_27_74#_c_577_n 0.00567107f $X=1.26 $Y=0.69 $X2=0 $Y2=0
cc_223 N_GATE_M1014_g N_A_27_74#_c_581_n 0.00933344f $X=1.26 $Y=0.69 $X2=0 $Y2=0
cc_224 N_GATE_M1014_g N_A_27_74#_c_559_n 0.00912427f $X=1.26 $Y=0.69 $X2=0 $Y2=0
cc_225 N_GATE_M1014_g N_A_27_74#_c_560_n 0.00289683f $X=1.26 $Y=0.69 $X2=0 $Y2=0
cc_226 N_GATE_c_224_n N_VPWR_c_750_n 0.0148788f $X=1.245 $Y=1.885 $X2=0 $Y2=0
cc_227 N_GATE_c_224_n N_VPWR_c_758_n 0.00461464f $X=1.245 $Y=1.885 $X2=0 $Y2=0
cc_228 N_GATE_c_224_n N_VPWR_c_749_n 0.00911543f $X=1.245 $Y=1.885 $X2=0 $Y2=0
cc_229 N_GATE_M1014_g N_VGND_c_849_n 0.00139764f $X=1.26 $Y=0.69 $X2=0 $Y2=0
cc_230 N_GATE_M1014_g N_VGND_c_855_n 0.00278237f $X=1.26 $Y=0.69 $X2=0 $Y2=0
cc_231 N_GATE_M1014_g N_VGND_c_864_n 0.00355577f $X=1.26 $Y=0.69 $X2=0 $Y2=0
cc_232 N_A_315_48#_c_273_n N_A_315_338#_c_415_n 0.0132581f $X=2.465 $Y=2.465
+ $X2=0 $Y2=0
cc_233 N_A_315_48#_c_264_n N_A_315_338#_c_415_n 0.00428065f $X=1.96 $Y=2.05
+ $X2=0 $Y2=0
cc_234 N_A_315_48#_c_277_n N_A_315_338#_c_415_n 0.00152992f $X=2.045 $Y=2.135
+ $X2=0 $Y2=0
cc_235 N_A_315_48#_c_281_n N_A_315_338#_c_415_n 5.8937e-19 $X=2.555 $Y=2.215
+ $X2=0 $Y2=0
cc_236 N_A_315_48#_c_273_n N_A_315_338#_c_405_n 0.021418f $X=2.465 $Y=2.465
+ $X2=0 $Y2=0
cc_237 N_A_315_48#_c_264_n N_A_315_338#_c_405_n 0.0127355f $X=1.96 $Y=2.05 $X2=0
+ $Y2=0
cc_238 N_A_315_48#_c_280_n N_A_315_338#_c_405_n 0.00586957f $X=2.225 $Y=2.215
+ $X2=0 $Y2=0
cc_239 N_A_315_48#_c_281_n N_A_315_338#_c_405_n 2.04762e-19 $X=2.555 $Y=2.215
+ $X2=0 $Y2=0
cc_240 N_A_315_48#_c_264_n N_A_315_338#_c_406_n 0.00166063f $X=1.96 $Y=2.05
+ $X2=0 $Y2=0
cc_241 N_A_315_48#_c_266_n N_A_315_338#_c_406_n 9.44863e-19 $X=1.88 $Y=1.285
+ $X2=0 $Y2=0
cc_242 N_A_315_48#_c_267_n N_A_315_338#_c_406_n 0.0274533f $X=1.88 $Y=1.285
+ $X2=0 $Y2=0
cc_243 N_A_315_48#_c_259_n N_A_315_338#_M1006_g 0.0124539f $X=1.65 $Y=1.12 $X2=0
+ $Y2=0
cc_244 N_A_315_48#_c_264_n N_A_315_338#_M1006_g 3.45059e-19 $X=1.96 $Y=2.05
+ $X2=0 $Y2=0
cc_245 N_A_315_48#_c_266_n N_A_315_338#_M1006_g 8.72535e-19 $X=1.88 $Y=1.285
+ $X2=0 $Y2=0
cc_246 N_A_315_48#_c_267_n N_A_315_338#_M1006_g 0.015433f $X=1.88 $Y=1.285 $X2=0
+ $Y2=0
cc_247 N_A_315_48#_c_273_n N_A_315_338#_c_408_n 0.00112784f $X=2.465 $Y=2.465
+ $X2=0 $Y2=0
cc_248 N_A_315_48#_c_266_n N_A_315_338#_c_408_n 0.0290018f $X=1.88 $Y=1.285
+ $X2=0 $Y2=0
cc_249 N_A_315_48#_c_267_n N_A_315_338#_c_408_n 4.40082e-19 $X=1.88 $Y=1.285
+ $X2=0 $Y2=0
cc_250 N_A_315_48#_c_281_n N_A_315_338#_c_408_n 0.0219306f $X=2.555 $Y=2.215
+ $X2=0 $Y2=0
cc_251 N_A_315_48#_c_268_n N_A_315_338#_c_408_n 0.00787853f $X=3.32 $Y=1.72
+ $X2=0 $Y2=0
cc_252 N_A_315_48#_c_264_n N_A_315_338#_c_409_n 0.0039305f $X=1.96 $Y=2.05 $X2=0
+ $Y2=0
cc_253 N_A_315_48#_c_281_n N_A_315_338#_c_409_n 3.75836e-19 $X=2.555 $Y=2.215
+ $X2=0 $Y2=0
cc_254 N_A_315_48#_M1011_g N_A_315_338#_c_410_n 0.0110475f $X=3.655 $Y=0.995
+ $X2=0 $Y2=0
cc_255 N_A_315_48#_c_263_n N_A_315_338#_c_410_n 0.00616339f $X=3.505 $Y=1.72
+ $X2=0 $Y2=0
cc_256 N_A_315_48#_c_278_n N_A_315_338#_c_410_n 0.0154262f $X=3.155 $Y=2.135
+ $X2=0 $Y2=0
cc_257 N_A_315_48#_c_268_n N_A_315_338#_c_410_n 0.0254905f $X=3.32 $Y=1.72 $X2=0
+ $Y2=0
cc_258 N_A_315_48#_c_266_n N_A_315_338#_c_411_n 0.0121988f $X=1.88 $Y=1.285
+ $X2=0 $Y2=0
cc_259 N_A_315_48#_c_267_n N_A_315_338#_c_411_n 0.00125415f $X=1.88 $Y=1.285
+ $X2=0 $Y2=0
cc_260 N_A_315_48#_c_260_n N_A_315_338#_c_420_n 0.018309f $X=3.595 $Y=2.045
+ $X2=0 $Y2=0
cc_261 N_A_315_48#_c_262_n N_A_315_338#_c_420_n 0.00514999f $X=3.995 $Y=1.63
+ $X2=0 $Y2=0
cc_262 N_A_315_48#_c_284_n N_A_315_338#_c_420_n 0.0585246f $X=4.38 $Y=2.24 $X2=0
+ $Y2=0
cc_263 N_A_315_48#_M1011_g N_A_315_338#_c_412_n 0.0152461f $X=3.655 $Y=0.995
+ $X2=0 $Y2=0
cc_264 N_A_315_48#_c_265_n N_A_315_338#_c_412_n 0.0502697f $X=4.43 $Y=0.74 $X2=0
+ $Y2=0
cc_265 N_A_315_48#_M1011_g N_A_315_338#_c_413_n 0.0041661f $X=3.655 $Y=0.995
+ $X2=0 $Y2=0
cc_266 N_A_315_48#_c_262_n N_A_315_338#_c_413_n 0.0070159f $X=3.995 $Y=1.63
+ $X2=0 $Y2=0
cc_267 N_A_315_48#_c_269_n N_A_315_338#_c_413_n 0.00330505f $X=4.16 $Y=1.72
+ $X2=0 $Y2=0
cc_268 N_A_315_48#_c_271_n N_A_315_338#_c_413_n 0.0147462f $X=4.402 $Y=1.275
+ $X2=0 $Y2=0
cc_269 N_A_315_48#_c_272_n N_A_315_338#_c_413_n 3.08675e-19 $X=4.16 $Y=1.63
+ $X2=0 $Y2=0
cc_270 N_A_315_48#_c_260_n N_A_315_338#_c_414_n 0.013422f $X=3.595 $Y=2.045
+ $X2=0 $Y2=0
cc_271 N_A_315_48#_M1011_g N_A_315_338#_c_414_n 0.0108872f $X=3.655 $Y=0.995
+ $X2=0 $Y2=0
cc_272 N_A_315_48#_c_262_n N_A_315_338#_c_414_n 0.00784757f $X=3.995 $Y=1.63
+ $X2=0 $Y2=0
cc_273 N_A_315_48#_c_278_n N_A_315_338#_c_414_n 0.00866805f $X=3.155 $Y=2.135
+ $X2=0 $Y2=0
cc_274 N_A_315_48#_c_279_n N_A_315_338#_c_414_n 0.0073632f $X=3.24 $Y=2.05 $X2=0
+ $Y2=0
cc_275 N_A_315_48#_c_268_n N_A_315_338#_c_414_n 0.024238f $X=3.32 $Y=1.72 $X2=0
+ $Y2=0
cc_276 N_A_315_48#_c_269_n N_A_315_338#_c_414_n 0.0245357f $X=4.16 $Y=1.72 $X2=0
+ $Y2=0
cc_277 N_A_315_48#_c_270_n N_A_315_338#_c_414_n 0.00511456f $X=4.187 $Y=1.555
+ $X2=0 $Y2=0
cc_278 N_A_315_48#_c_285_n N_A_315_338#_c_414_n 0.00716634f $X=4.377 $Y=2.075
+ $X2=0 $Y2=0
cc_279 N_A_315_48#_c_272_n N_A_315_338#_c_414_n 0.00124916f $X=4.16 $Y=1.63
+ $X2=0 $Y2=0
cc_280 N_A_315_48#_c_269_n N_CLK_c_507_n 0.00389336f $X=4.16 $Y=1.72 $X2=0 $Y2=0
cc_281 N_A_315_48#_c_284_n N_CLK_c_508_n 0.00466733f $X=4.38 $Y=2.24 $X2=0 $Y2=0
cc_282 N_A_315_48#_c_285_n N_CLK_c_508_n 0.00404765f $X=4.377 $Y=2.075 $X2=0
+ $Y2=0
cc_283 N_A_315_48#_c_265_n N_CLK_c_503_n 0.00589627f $X=4.43 $Y=0.74 $X2=0 $Y2=0
cc_284 N_A_315_48#_c_270_n N_CLK_c_503_n 0.00400418f $X=4.187 $Y=1.555 $X2=0
+ $Y2=0
cc_285 N_A_315_48#_c_271_n N_CLK_c_503_n 0.00229573f $X=4.402 $Y=1.275 $X2=0
+ $Y2=0
cc_286 N_A_315_48#_c_270_n CLK 0.0276167f $X=4.187 $Y=1.555 $X2=0 $Y2=0
cc_287 N_A_315_48#_c_271_n CLK 0.00263579f $X=4.402 $Y=1.275 $X2=0 $Y2=0
cc_288 N_A_315_48#_c_272_n CLK 2.40403e-19 $X=4.16 $Y=1.63 $X2=0 $Y2=0
cc_289 N_A_315_48#_c_270_n N_CLK_c_506_n 0.00389336f $X=4.187 $Y=1.555 $X2=0
+ $Y2=0
cc_290 N_A_315_48#_c_272_n N_CLK_c_506_n 0.0210768f $X=4.16 $Y=1.63 $X2=0 $Y2=0
cc_291 N_A_315_48#_c_273_n N_A_27_74#_M1010_g 0.0225424f $X=2.465 $Y=2.465 $X2=0
+ $Y2=0
cc_292 N_A_315_48#_c_260_n N_A_27_74#_M1010_g 0.003095f $X=3.595 $Y=2.045 $X2=0
+ $Y2=0
cc_293 N_A_315_48#_M1011_g N_A_27_74#_M1010_g 0.0113463f $X=3.655 $Y=0.995 $X2=0
+ $Y2=0
cc_294 N_A_315_48#_c_263_n N_A_27_74#_M1010_g 0.0214198f $X=3.505 $Y=1.72 $X2=0
+ $Y2=0
cc_295 N_A_315_48#_c_278_n N_A_27_74#_M1010_g 0.00730665f $X=3.155 $Y=2.135
+ $X2=0 $Y2=0
cc_296 N_A_315_48#_c_279_n N_A_27_74#_M1010_g 0.0036304f $X=3.24 $Y=2.05 $X2=0
+ $Y2=0
cc_297 N_A_315_48#_c_268_n N_A_27_74#_M1010_g 0.00140735f $X=3.32 $Y=1.72 $X2=0
+ $Y2=0
cc_298 N_A_315_48#_c_260_n N_A_27_74#_c_566_n 0.00711088f $X=3.595 $Y=2.045
+ $X2=0 $Y2=0
cc_299 N_A_315_48#_c_278_n N_A_27_74#_c_566_n 0.00434335f $X=3.155 $Y=2.135
+ $X2=0 $Y2=0
cc_300 N_A_315_48#_c_278_n N_A_27_74#_c_567_n 0.00724123f $X=3.155 $Y=2.135
+ $X2=0 $Y2=0
cc_301 N_A_315_48#_c_281_n N_A_27_74#_c_567_n 0.00104714f $X=2.555 $Y=2.215
+ $X2=0 $Y2=0
cc_302 N_A_315_48#_c_273_n N_A_27_74#_c_568_n 0.0289004f $X=2.465 $Y=2.465 $X2=0
+ $Y2=0
cc_303 N_A_315_48#_c_260_n N_A_27_74#_c_568_n 0.0101963f $X=3.595 $Y=2.045 $X2=0
+ $Y2=0
cc_304 N_A_315_48#_M1011_g N_A_27_74#_c_554_n 0.00895007f $X=3.655 $Y=0.995
+ $X2=0 $Y2=0
cc_305 N_A_315_48#_c_265_n N_A_27_74#_c_554_n 0.00735365f $X=4.43 $Y=0.74 $X2=0
+ $Y2=0
cc_306 N_A_315_48#_c_259_n N_A_27_74#_c_581_n 0.00111122f $X=1.65 $Y=1.12 $X2=0
+ $Y2=0
cc_307 N_A_315_48#_c_259_n N_A_27_74#_c_559_n 0.0110834f $X=1.65 $Y=1.12 $X2=0
+ $Y2=0
cc_308 N_A_315_48#_M1011_g N_A_27_74#_c_564_n 0.00187881f $X=3.655 $Y=0.995
+ $X2=0 $Y2=0
cc_309 N_A_315_48#_c_278_n N_VPWR_M1021_d 0.00276374f $X=3.155 $Y=2.135 $X2=0
+ $Y2=0
cc_310 N_A_315_48#_c_273_n N_VPWR_c_751_n 0.00168108f $X=2.465 $Y=2.465 $X2=0
+ $Y2=0
cc_311 N_A_315_48#_c_260_n N_VPWR_c_751_n 0.00634677f $X=3.595 $Y=2.045 $X2=0
+ $Y2=0
cc_312 N_A_315_48#_c_278_n N_VPWR_c_751_n 0.0152878f $X=3.155 $Y=2.135 $X2=0
+ $Y2=0
cc_313 N_A_315_48#_c_284_n N_VPWR_c_752_n 0.00316551f $X=4.38 $Y=2.24 $X2=0
+ $Y2=0
cc_314 N_A_315_48#_c_260_n N_VPWR_c_756_n 0.00445602f $X=3.595 $Y=2.045 $X2=0
+ $Y2=0
cc_315 N_A_315_48#_c_284_n N_VPWR_c_756_n 0.0135015f $X=4.38 $Y=2.24 $X2=0 $Y2=0
cc_316 N_A_315_48#_c_273_n N_VPWR_c_758_n 0.00445785f $X=2.465 $Y=2.465 $X2=0
+ $Y2=0
cc_317 N_A_315_48#_c_273_n N_VPWR_c_749_n 0.00893057f $X=2.465 $Y=2.465 $X2=0
+ $Y2=0
cc_318 N_A_315_48#_c_260_n N_VPWR_c_749_n 0.00863669f $X=3.595 $Y=2.045 $X2=0
+ $Y2=0
cc_319 N_A_315_48#_c_284_n N_VPWR_c_749_n 0.0121118f $X=4.38 $Y=2.24 $X2=0 $Y2=0
cc_320 N_A_315_48#_M1011_g N_VGND_c_850_n 0.00302736f $X=3.655 $Y=0.995 $X2=0
+ $Y2=0
cc_321 N_A_315_48#_c_265_n N_VGND_c_850_n 9.16406e-19 $X=4.43 $Y=0.74 $X2=0
+ $Y2=0
cc_322 N_A_315_48#_c_265_n N_VGND_c_851_n 0.0276447f $X=4.43 $Y=0.74 $X2=0 $Y2=0
cc_323 N_A_315_48#_c_259_n N_VGND_c_855_n 0.00278271f $X=1.65 $Y=1.12 $X2=0
+ $Y2=0
cc_324 N_A_315_48#_c_265_n N_VGND_c_858_n 0.00877136f $X=4.43 $Y=0.74 $X2=0
+ $Y2=0
cc_325 N_A_315_48#_c_259_n N_VGND_c_864_n 0.00358137f $X=1.65 $Y=1.12 $X2=0
+ $Y2=0
cc_326 N_A_315_48#_M1011_g N_VGND_c_864_n 9.49986e-19 $X=3.655 $Y=0.995 $X2=0
+ $Y2=0
cc_327 N_A_315_48#_c_265_n N_VGND_c_864_n 0.0106073f $X=4.43 $Y=0.74 $X2=0 $Y2=0
cc_328 N_A_315_338#_c_420_n N_CLK_c_508_n 0.00199604f $X=3.82 $Y=2.265 $X2=0
+ $Y2=0
cc_329 N_A_315_338#_c_413_n N_CLK_c_503_n 4.074e-19 $X=3.845 $Y=1.3 $X2=0 $Y2=0
cc_330 N_A_315_338#_c_408_n N_A_27_74#_M1010_g 0.00424756f $X=2.42 $Y=1.675
+ $X2=0 $Y2=0
cc_331 N_A_315_338#_c_409_n N_A_27_74#_M1010_g 0.0210112f $X=2.42 $Y=1.675 $X2=0
+ $Y2=0
cc_332 N_A_315_338#_c_410_n N_A_27_74#_M1010_g 0.0166946f $X=3.655 $Y=1.3 $X2=0
+ $Y2=0
cc_333 N_A_315_338#_c_420_n N_A_27_74#_c_567_n 5.25341e-19 $X=3.82 $Y=2.265
+ $X2=0 $Y2=0
cc_334 N_A_315_338#_c_420_n N_A_27_74#_c_568_n 0.00147927f $X=3.82 $Y=2.265
+ $X2=0 $Y2=0
cc_335 N_A_315_338#_c_412_n N_A_27_74#_c_554_n 0.00610504f $X=3.87 $Y=0.77 $X2=0
+ $Y2=0
cc_336 N_A_315_338#_M1006_g N_A_27_74#_c_559_n 0.00721522f $X=2.395 $Y=0.8 $X2=0
+ $Y2=0
cc_337 N_A_315_338#_M1006_g N_A_27_74#_c_563_n 7.06434e-19 $X=2.395 $Y=0.8 $X2=0
+ $Y2=0
cc_338 N_A_315_338#_c_410_n N_A_27_74#_c_563_n 0.00214479f $X=3.655 $Y=1.3 $X2=0
+ $Y2=0
cc_339 N_A_315_338#_M1006_g N_A_27_74#_c_564_n 0.04087f $X=2.395 $Y=0.8 $X2=0
+ $Y2=0
cc_340 N_A_315_338#_c_420_n N_VPWR_c_751_n 0.0132339f $X=3.82 $Y=2.265 $X2=0
+ $Y2=0
cc_341 N_A_315_338#_c_420_n N_VPWR_c_756_n 0.0145938f $X=3.82 $Y=2.265 $X2=0
+ $Y2=0
cc_342 N_A_315_338#_c_415_n N_VPWR_c_758_n 0.0030458f $X=1.665 $Y=1.885 $X2=0
+ $Y2=0
cc_343 N_A_315_338#_c_415_n N_VPWR_c_749_n 0.00376093f $X=1.665 $Y=1.885 $X2=0
+ $Y2=0
cc_344 N_A_315_338#_c_420_n N_VPWR_c_749_n 0.0120466f $X=3.82 $Y=2.265 $X2=0
+ $Y2=0
cc_345 N_A_315_338#_c_410_n N_VGND_M1010_d 0.00281417f $X=3.655 $Y=1.3 $X2=0
+ $Y2=0
cc_346 N_A_315_338#_M1006_g N_VGND_c_867_n 8.6539e-19 $X=2.395 $Y=0.8 $X2=0
+ $Y2=0
cc_347 N_A_315_338#_c_410_n N_VGND_c_867_n 0.0253449f $X=3.655 $Y=1.3 $X2=0
+ $Y2=0
cc_348 N_A_315_338#_c_410_n N_VGND_c_850_n 0.0126838f $X=3.655 $Y=1.3 $X2=0
+ $Y2=0
cc_349 N_A_315_338#_c_412_n N_VGND_c_850_n 0.00635827f $X=3.87 $Y=0.77 $X2=0
+ $Y2=0
cc_350 N_A_315_338#_c_412_n N_VGND_c_858_n 0.00701036f $X=3.87 $Y=0.77 $X2=0
+ $Y2=0
cc_351 N_A_315_338#_c_412_n N_VGND_c_864_n 0.00885159f $X=3.87 $Y=0.77 $X2=0
+ $Y2=0
cc_352 N_CLK_c_503_n N_A_27_74#_c_554_n 0.0103003f $X=4.645 $Y=1.445 $X2=0 $Y2=0
cc_353 N_CLK_c_504_n N_A_27_74#_c_554_n 0.0103107f $X=5.145 $Y=1.445 $X2=0 $Y2=0
cc_354 N_CLK_c_504_n N_A_27_74#_M1018_g 0.0322821f $X=5.145 $Y=1.445 $X2=0 $Y2=0
cc_355 CLK N_A_27_74#_c_556_n 2.24258e-19 $X=4.955 $Y=1.58 $X2=0 $Y2=0
cc_356 N_CLK_c_506_n N_A_27_74#_c_556_n 0.0123722f $X=5.13 $Y=1.652 $X2=0 $Y2=0
cc_357 N_CLK_c_509_n N_A_27_74#_c_570_n 0.00694438f $X=5.13 $Y=1.86 $X2=0 $Y2=0
cc_358 N_CLK_c_506_n N_A_27_74#_c_557_n 0.0322821f $X=5.13 $Y=1.652 $X2=0 $Y2=0
cc_359 N_CLK_c_504_n N_A_1041_387#_c_692_n 9.93468e-19 $X=5.145 $Y=1.445 $X2=0
+ $Y2=0
cc_360 N_CLK_c_509_n N_A_1041_387#_c_693_n 0.00179242f $X=5.13 $Y=1.86 $X2=0
+ $Y2=0
cc_361 CLK N_A_1041_387#_c_693_n 0.0134897f $X=4.955 $Y=1.58 $X2=0 $Y2=0
cc_362 N_CLK_c_506_n N_A_1041_387#_c_693_n 0.00223607f $X=5.13 $Y=1.652 $X2=0
+ $Y2=0
cc_363 N_CLK_c_504_n N_A_1041_387#_c_694_n 0.00396135f $X=5.145 $Y=1.445 $X2=0
+ $Y2=0
cc_364 CLK N_A_1041_387#_c_694_n 0.0145166f $X=4.955 $Y=1.58 $X2=0 $Y2=0
cc_365 N_CLK_c_506_n N_A_1041_387#_c_694_n 6.25973e-19 $X=5.13 $Y=1.652 $X2=0
+ $Y2=0
cc_366 N_CLK_c_508_n N_VPWR_c_752_n 0.00450659f $X=4.625 $Y=2.02 $X2=0 $Y2=0
cc_367 N_CLK_c_509_n N_VPWR_c_752_n 0.0043597f $X=5.13 $Y=1.86 $X2=0 $Y2=0
cc_368 CLK N_VPWR_c_752_n 0.017905f $X=4.955 $Y=1.58 $X2=0 $Y2=0
cc_369 N_CLK_c_506_n N_VPWR_c_752_n 0.00220066f $X=5.13 $Y=1.652 $X2=0 $Y2=0
cc_370 N_CLK_c_508_n N_VPWR_c_756_n 0.00559701f $X=4.625 $Y=2.02 $X2=0 $Y2=0
cc_371 N_CLK_c_509_n N_VPWR_c_759_n 0.00559701f $X=5.13 $Y=1.86 $X2=0 $Y2=0
cc_372 N_CLK_c_508_n N_VPWR_c_749_n 0.00537853f $X=4.625 $Y=2.02 $X2=0 $Y2=0
cc_373 N_CLK_c_509_n N_VPWR_c_749_n 0.00537853f $X=5.13 $Y=1.86 $X2=0 $Y2=0
cc_374 N_CLK_c_503_n N_VGND_c_851_n 0.00683202f $X=4.645 $Y=1.445 $X2=0 $Y2=0
cc_375 N_CLK_c_504_n N_VGND_c_851_n 0.0140738f $X=5.145 $Y=1.445 $X2=0 $Y2=0
cc_376 CLK N_VGND_c_851_n 0.023955f $X=4.955 $Y=1.58 $X2=0 $Y2=0
cc_377 N_CLK_c_506_n N_VGND_c_851_n 0.00396026f $X=5.13 $Y=1.652 $X2=0 $Y2=0
cc_378 N_CLK_c_503_n N_VGND_c_864_n 9.39239e-19 $X=4.645 $Y=1.445 $X2=0 $Y2=0
cc_379 N_CLK_c_504_n N_VGND_c_864_n 7.88961e-19 $X=5.145 $Y=1.445 $X2=0 $Y2=0
cc_380 N_A_27_74#_c_557_n N_A_1041_387#_c_686_n 0.00908904f $X=5.562 $Y=1.56
+ $X2=0 $Y2=0
cc_381 N_A_27_74#_c_570_n N_A_1041_387#_c_698_n 0.00967397f $X=5.605 $Y=1.86
+ $X2=0 $Y2=0
cc_382 N_A_27_74#_M1018_g N_A_1041_387#_c_692_n 0.00687676f $X=5.505 $Y=0.965
+ $X2=0 $Y2=0
cc_383 N_A_27_74#_c_557_n N_A_1041_387#_c_692_n 2.72517e-19 $X=5.562 $Y=1.56
+ $X2=0 $Y2=0
cc_384 N_A_27_74#_c_570_n N_A_1041_387#_c_711_n 0.00189113f $X=5.605 $Y=1.86
+ $X2=0 $Y2=0
cc_385 N_A_27_74#_c_556_n N_A_1041_387#_c_693_n 0.00800492f $X=5.605 $Y=1.77
+ $X2=0 $Y2=0
cc_386 N_A_27_74#_c_570_n N_A_1041_387#_c_693_n 0.00901125f $X=5.605 $Y=1.86
+ $X2=0 $Y2=0
cc_387 N_A_27_74#_c_557_n N_A_1041_387#_c_693_n 7.73634e-19 $X=5.562 $Y=1.56
+ $X2=0 $Y2=0
cc_388 N_A_27_74#_M1018_g N_A_1041_387#_c_694_n 0.0162742f $X=5.505 $Y=0.965
+ $X2=0 $Y2=0
cc_389 N_A_27_74#_c_556_n N_A_1041_387#_c_694_n 0.0088198f $X=5.605 $Y=1.77
+ $X2=0 $Y2=0
cc_390 N_A_27_74#_c_557_n N_A_1041_387#_c_694_n 0.00971201f $X=5.562 $Y=1.56
+ $X2=0 $Y2=0
cc_391 N_A_27_74#_M1018_g N_A_1041_387#_c_695_n 0.00849677f $X=5.505 $Y=0.965
+ $X2=0 $Y2=0
cc_392 N_A_27_74#_c_571_n N_VPWR_c_750_n 0.0418595f $X=0.28 $Y=2.815 $X2=0 $Y2=0
cc_393 N_A_27_74#_c_568_n N_VPWR_c_751_n 0.0163301f $X=2.885 $Y=2.465 $X2=0
+ $Y2=0
cc_394 N_A_27_74#_c_570_n N_VPWR_c_753_n 0.00560846f $X=5.605 $Y=1.86 $X2=0
+ $Y2=0
cc_395 N_A_27_74#_c_568_n N_VPWR_c_758_n 0.00413917f $X=2.885 $Y=2.465 $X2=0
+ $Y2=0
cc_396 N_A_27_74#_c_570_n N_VPWR_c_759_n 0.00528708f $X=5.605 $Y=1.86 $X2=0
+ $Y2=0
cc_397 N_A_27_74#_c_571_n N_VPWR_c_761_n 0.0154862f $X=0.28 $Y=2.815 $X2=0 $Y2=0
cc_398 N_A_27_74#_c_568_n N_VPWR_c_749_n 0.0085536f $X=2.885 $Y=2.465 $X2=0
+ $Y2=0
cc_399 N_A_27_74#_c_570_n N_VPWR_c_749_n 0.00537853f $X=5.605 $Y=1.86 $X2=0
+ $Y2=0
cc_400 N_A_27_74#_c_571_n N_VPWR_c_749_n 0.0127853f $X=0.28 $Y=2.815 $X2=0 $Y2=0
cc_401 N_A_27_74#_c_577_n N_VGND_M1020_d 0.0131464f $X=1.05 $Y=0.855 $X2=-0.19
+ $Y2=-0.245
cc_402 N_A_27_74#_c_581_n N_VGND_M1020_d 0.00419505f $X=1.135 $Y=0.77 $X2=-0.19
+ $Y2=-0.245
cc_403 N_A_27_74#_c_560_n N_VGND_M1020_d 5.38677e-19 $X=1.22 $Y=0.34 $X2=-0.19
+ $Y2=-0.245
cc_404 N_A_27_74#_c_558_n N_VGND_c_849_n 0.00971749f $X=0.28 $Y=0.645 $X2=0
+ $Y2=0
cc_405 N_A_27_74#_c_577_n N_VGND_c_849_n 0.0216654f $X=1.05 $Y=0.855 $X2=0 $Y2=0
cc_406 N_A_27_74#_c_581_n N_VGND_c_849_n 0.0133532f $X=1.135 $Y=0.77 $X2=0 $Y2=0
cc_407 N_A_27_74#_c_560_n N_VGND_c_849_n 0.0148722f $X=1.22 $Y=0.34 $X2=0 $Y2=0
cc_408 N_A_27_74#_M1010_g N_VGND_c_867_n 0.00566712f $X=2.87 $Y=0.905 $X2=0
+ $Y2=0
cc_409 N_A_27_74#_c_554_n N_VGND_c_867_n 0.00146902f $X=5.43 $Y=0.18 $X2=0 $Y2=0
cc_410 N_A_27_74#_c_563_n N_VGND_c_867_n 0.0154871f $X=2.995 $Y=0.34 $X2=0 $Y2=0
cc_411 N_A_27_74#_c_564_n N_VGND_c_867_n 0.00140632f $X=2.977 $Y=0.18 $X2=0
+ $Y2=0
cc_412 N_A_27_74#_M1010_g N_VGND_c_850_n 0.0028708f $X=2.87 $Y=0.905 $X2=0 $Y2=0
cc_413 N_A_27_74#_c_554_n N_VGND_c_850_n 0.0183632f $X=5.43 $Y=0.18 $X2=0 $Y2=0
cc_414 N_A_27_74#_c_563_n N_VGND_c_850_n 0.0240076f $X=2.995 $Y=0.34 $X2=0 $Y2=0
cc_415 N_A_27_74#_c_564_n N_VGND_c_850_n 0.00620031f $X=2.977 $Y=0.18 $X2=0
+ $Y2=0
cc_416 N_A_27_74#_c_554_n N_VGND_c_851_n 0.0256157f $X=5.43 $Y=0.18 $X2=0 $Y2=0
cc_417 N_A_27_74#_M1018_g N_VGND_c_851_n 0.00840262f $X=5.505 $Y=0.965 $X2=0
+ $Y2=0
cc_418 N_A_27_74#_c_559_n N_VGND_c_855_n 0.102814f $X=2.83 $Y=0.34 $X2=0 $Y2=0
cc_419 N_A_27_74#_c_560_n N_VGND_c_855_n 0.0120704f $X=1.22 $Y=0.34 $X2=0 $Y2=0
cc_420 N_A_27_74#_c_563_n N_VGND_c_855_n 0.0212434f $X=2.995 $Y=0.34 $X2=0 $Y2=0
cc_421 N_A_27_74#_c_564_n N_VGND_c_855_n 0.01344f $X=2.977 $Y=0.18 $X2=0 $Y2=0
cc_422 N_A_27_74#_c_558_n N_VGND_c_857_n 0.011913f $X=0.28 $Y=0.645 $X2=0 $Y2=0
cc_423 N_A_27_74#_c_554_n N_VGND_c_858_n 0.0354459f $X=5.43 $Y=0.18 $X2=0 $Y2=0
cc_424 N_A_27_74#_c_554_n N_VGND_c_859_n 0.017704f $X=5.43 $Y=0.18 $X2=0 $Y2=0
cc_425 N_A_27_74#_c_554_n N_VGND_c_864_n 0.0725918f $X=5.43 $Y=0.18 $X2=0 $Y2=0
cc_426 N_A_27_74#_c_558_n N_VGND_c_864_n 0.00988061f $X=0.28 $Y=0.645 $X2=0
+ $Y2=0
cc_427 N_A_27_74#_c_577_n N_VGND_c_864_n 0.0131405f $X=1.05 $Y=0.855 $X2=0 $Y2=0
cc_428 N_A_27_74#_c_559_n N_VGND_c_864_n 0.0591639f $X=2.83 $Y=0.34 $X2=0 $Y2=0
cc_429 N_A_27_74#_c_560_n N_VGND_c_864_n 0.00645034f $X=1.22 $Y=0.34 $X2=0 $Y2=0
cc_430 N_A_27_74#_c_563_n N_VGND_c_864_n 0.0110272f $X=2.995 $Y=0.34 $X2=0 $Y2=0
cc_431 N_A_27_74#_c_564_n N_VGND_c_864_n 0.0111058f $X=2.977 $Y=0.18 $X2=0 $Y2=0
cc_432 N_A_27_74#_c_559_n A_267_74# 0.00142017f $X=2.83 $Y=0.34 $X2=-0.19
+ $Y2=-0.245
cc_433 N_A_1041_387#_c_698_n N_VPWR_c_752_n 0.00158629f $X=5.38 $Y=2.81 $X2=0
+ $Y2=0
cc_434 N_A_1041_387#_c_686_n N_VPWR_c_753_n 0.0194855f $X=6.305 $Y=1.49 $X2=0
+ $Y2=0
cc_435 N_A_1041_387#_c_687_n N_VPWR_c_753_n 0.0057847f $X=6.725 $Y=1.765 $X2=0
+ $Y2=0
cc_436 N_A_1041_387#_c_711_n N_VPWR_c_753_n 0.0388118f $X=5.38 $Y=2.095 $X2=0
+ $Y2=0
cc_437 N_A_1041_387#_c_694_n N_VPWR_c_753_n 0.0302304f $X=6.14 $Y=1.105 $X2=0
+ $Y2=0
cc_438 N_A_1041_387#_c_690_n N_VPWR_c_755_n 0.00972643f $X=7.175 $Y=1.765 $X2=0
+ $Y2=0
cc_439 N_A_1041_387#_c_698_n N_VPWR_c_759_n 0.0138236f $X=5.38 $Y=2.81 $X2=0
+ $Y2=0
cc_440 N_A_1041_387#_c_687_n N_VPWR_c_760_n 0.00461464f $X=6.725 $Y=1.765 $X2=0
+ $Y2=0
cc_441 N_A_1041_387#_c_690_n N_VPWR_c_760_n 0.00422942f $X=7.175 $Y=1.765 $X2=0
+ $Y2=0
cc_442 N_A_1041_387#_c_687_n N_VPWR_c_749_n 0.00912633f $X=6.725 $Y=1.765 $X2=0
+ $Y2=0
cc_443 N_A_1041_387#_c_690_n N_VPWR_c_749_n 0.0078771f $X=7.175 $Y=1.765 $X2=0
+ $Y2=0
cc_444 N_A_1041_387#_c_698_n N_VPWR_c_749_n 0.0124505f $X=5.38 $Y=2.81 $X2=0
+ $Y2=0
cc_445 N_A_1041_387#_c_687_n GCLK 0.0182089f $X=6.725 $Y=1.765 $X2=0 $Y2=0
cc_446 N_A_1041_387#_M1001_g GCLK 0.0216129f $X=6.755 $Y=0.83 $X2=0 $Y2=0
cc_447 N_A_1041_387#_c_689_n GCLK 0.0144436f $X=7.085 $Y=1.49 $X2=0 $Y2=0
cc_448 N_A_1041_387#_c_690_n GCLK 0.0413205f $X=7.175 $Y=1.765 $X2=0 $Y2=0
cc_449 N_A_1041_387#_c_691_n GCLK 0.0149078f $X=7.185 $Y=1.31 $X2=0 $Y2=0
cc_450 N_A_1041_387#_c_694_n GCLK 0.0220232f $X=6.14 $Y=1.105 $X2=0 $Y2=0
cc_451 N_A_1041_387#_c_695_n GCLK 4.46319e-19 $X=6.14 $Y=1.105 $X2=0 $Y2=0
cc_452 N_A_1041_387#_c_692_n N_VGND_c_851_n 0.0122119f $X=5.72 $Y=0.74 $X2=0
+ $Y2=0
cc_453 N_A_1041_387#_c_685_n N_VGND_c_852_n 0.00536837f $X=6.635 $Y=1.49 $X2=0
+ $Y2=0
cc_454 N_A_1041_387#_M1001_g N_VGND_c_852_n 0.011131f $X=6.755 $Y=0.83 $X2=0
+ $Y2=0
cc_455 N_A_1041_387#_c_692_n N_VGND_c_852_n 0.00869348f $X=5.72 $Y=0.74 $X2=0
+ $Y2=0
cc_456 N_A_1041_387#_c_691_n N_VGND_c_854_n 0.00650727f $X=7.185 $Y=1.31 $X2=0
+ $Y2=0
cc_457 N_A_1041_387#_c_692_n N_VGND_c_859_n 0.00717288f $X=5.72 $Y=0.74 $X2=0
+ $Y2=0
cc_458 N_A_1041_387#_M1001_g N_VGND_c_860_n 0.00491683f $X=6.755 $Y=0.83 $X2=0
+ $Y2=0
cc_459 N_A_1041_387#_c_691_n N_VGND_c_860_n 0.00491683f $X=7.185 $Y=1.31 $X2=0
+ $Y2=0
cc_460 N_A_1041_387#_M1001_g N_VGND_c_864_n 0.00517496f $X=6.755 $Y=0.83 $X2=0
+ $Y2=0
cc_461 N_A_1041_387#_c_691_n N_VGND_c_864_n 0.00517496f $X=7.185 $Y=1.31 $X2=0
+ $Y2=0
cc_462 N_A_1041_387#_c_692_n N_VGND_c_864_n 0.0100033f $X=5.72 $Y=0.74 $X2=0
+ $Y2=0
cc_463 N_VPWR_c_753_n GCLK 0.00167254f $X=5.835 $Y=2.115 $X2=0 $Y2=0
cc_464 N_VPWR_c_755_n GCLK 0.0844051f $X=7.4 $Y=1.985 $X2=0 $Y2=0
cc_465 N_VPWR_c_760_n GCLK 0.014534f $X=7.315 $Y=3.33 $X2=0 $Y2=0
cc_466 N_VPWR_c_749_n GCLK 0.0119501f $X=7.44 $Y=3.33 $X2=0 $Y2=0
cc_467 N_VPWR_c_755_n N_VGND_c_854_n 0.0096123f $X=7.4 $Y=1.985 $X2=0 $Y2=0
cc_468 GCLK N_VGND_c_852_n 0.0131729f $X=6.875 $Y=0.47 $X2=0 $Y2=0
cc_469 GCLK N_VGND_c_854_n 0.0294122f $X=6.875 $Y=0.47 $X2=0 $Y2=0
cc_470 GCLK N_VGND_c_860_n 0.0105983f $X=6.875 $Y=0.47 $X2=0 $Y2=0
cc_471 GCLK N_VGND_c_864_n 0.0113894f $X=6.875 $Y=0.47 $X2=0 $Y2=0
