* File: sky130_fd_sc_hs__a22o_1.pxi.spice
* Created: Thu Aug 27 20:26:51 2020
* 
x_PM_SKY130_FD_SC_HS__A22O_1%A2 N_A2_c_57_n N_A2_c_58_n N_A2_c_63_n N_A2_M1009_g
+ N_A2_M1002_g A2 N_A2_c_61_n PM_SKY130_FD_SC_HS__A22O_1%A2
x_PM_SKY130_FD_SC_HS__A22O_1%B2 N_B2_c_88_n N_B2_M1003_g N_B2_M1004_g B2 B2
+ N_B2_c_90_n PM_SKY130_FD_SC_HS__A22O_1%B2
x_PM_SKY130_FD_SC_HS__A22O_1%B1 N_B1_M1000_g N_B1_c_123_n N_B1_c_124_n
+ N_B1_M1006_g N_B1_c_125_n N_B1_c_126_n B1 PM_SKY130_FD_SC_HS__A22O_1%B1
x_PM_SKY130_FD_SC_HS__A22O_1%A1 N_A1_c_159_n N_A1_M1005_g N_A1_c_160_n
+ N_A1_M1001_g A1 N_A1_c_161_n PM_SKY130_FD_SC_HS__A22O_1%A1
x_PM_SKY130_FD_SC_HS__A22O_1%A_222_392# N_A_222_392#_M1000_d
+ N_A_222_392#_M1003_d N_A_222_392#_c_194_n N_A_222_392#_M1007_g
+ N_A_222_392#_M1008_g N_A_222_392#_c_204_n N_A_222_392#_c_196_n
+ N_A_222_392#_c_197_n N_A_222_392#_c_201_n N_A_222_392#_c_198_n
+ PM_SKY130_FD_SC_HS__A22O_1%A_222_392#
x_PM_SKY130_FD_SC_HS__A22O_1%VPWR N_VPWR_M1009_s N_VPWR_M1001_d N_VPWR_c_252_n
+ N_VPWR_c_253_n N_VPWR_c_254_n VPWR N_VPWR_c_255_n N_VPWR_c_256_n
+ N_VPWR_c_251_n N_VPWR_c_258_n PM_SKY130_FD_SC_HS__A22O_1%VPWR
x_PM_SKY130_FD_SC_HS__A22O_1%A_132_392# N_A_132_392#_M1009_d
+ N_A_132_392#_M1006_d N_A_132_392#_c_288_n N_A_132_392#_c_286_n
+ N_A_132_392#_c_287_n N_A_132_392#_c_295_n
+ PM_SKY130_FD_SC_HS__A22O_1%A_132_392#
x_PM_SKY130_FD_SC_HS__A22O_1%X N_X_M1008_d N_X_M1007_d X X X X X X X
+ PM_SKY130_FD_SC_HS__A22O_1%X
x_PM_SKY130_FD_SC_HS__A22O_1%A_52_123# N_A_52_123#_M1002_s N_A_52_123#_M1005_d
+ N_A_52_123#_c_321_n N_A_52_123#_c_322_n N_A_52_123#_c_323_n
+ N_A_52_123#_c_324_n N_A_52_123#_c_325_n PM_SKY130_FD_SC_HS__A22O_1%A_52_123#
x_PM_SKY130_FD_SC_HS__A22O_1%VGND N_VGND_M1002_d N_VGND_M1008_s N_VGND_c_364_n
+ N_VGND_c_365_n N_VGND_c_366_n N_VGND_c_367_n VGND N_VGND_c_368_n
+ N_VGND_c_369_n N_VGND_c_370_n N_VGND_c_371_n PM_SKY130_FD_SC_HS__A22O_1%VGND
cc_1 VNB N_A2_c_57_n 0.00865851f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.42
cc_2 VNB N_A2_c_58_n 0.015328f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.795
cc_3 VNB N_A2_M1002_g 0.0113873f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=0.935
cc_4 VNB A2 0.0232559f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.47
cc_5 VNB N_A2_c_61_n 0.0570677f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=0.34
cc_6 VNB N_B2_c_88_n 0.0149141f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.42
cc_7 VNB N_B2_M1004_g 0.0316329f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=0.505
cc_8 VNB N_B2_c_90_n 0.0183584f $X=-0.19 $Y=-0.245 $X2=0.395 $Y2=0.34
cc_9 VNB N_B1_c_123_n 0.0120262f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=2.46
cc_10 VNB N_B1_c_124_n 0.0152531f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=0.505
cc_11 VNB N_B1_c_125_n 0.0137133f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=0.935
cc_12 VNB N_B1_c_126_n 0.0133794f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.33
cc_13 VNB B1 0.00283269f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.47
cc_14 VNB N_A1_c_159_n 0.0163683f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.42
cc_15 VNB N_A1_c_160_n 0.0588577f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=2.46
cc_16 VNB N_A1_c_161_n 0.00166777f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.47
cc_17 VNB N_A_222_392#_c_194_n 0.0487841f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=1.33
cc_18 VNB N_A_222_392#_M1008_g 0.0295424f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_222_392#_c_196_n 0.0190281f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_222_392#_c_197_n 0.00233602f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_222_392#_c_198_n 0.00179529f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_VPWR_c_251_n 0.143779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB X 0.0565573f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=1.33
cc_24 VNB N_A_52_123#_c_321_n 0.00794929f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=1.33
cc_25 VNB N_A_52_123#_c_322_n 5.74149e-19 $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.33
cc_26 VNB N_A_52_123#_c_323_n 0.00120814f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.47
cc_27 VNB N_A_52_123#_c_324_n 0.00843668f $X=-0.19 $Y=-0.245 $X2=0.395 $Y2=0.34
cc_28 VNB N_A_52_123#_c_325_n 0.0209393f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_364_n 0.0106411f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=0.935
cc_30 VNB N_VGND_c_365_n 0.0161981f $X=-0.19 $Y=-0.245 $X2=0.395 $Y2=0.34
cc_31 VNB N_VGND_c_366_n 0.021055f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_367_n 0.00413177f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=0.34
cc_33 VNB N_VGND_c_368_n 0.0408693f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_369_n 0.0191515f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_370_n 0.221318f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_371_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VPB N_A2_c_58_n 0.00776182f $X=-0.19 $Y=1.66 $X2=0.585 $Y2=1.795
cc_38 VPB N_A2_c_63_n 0.0266633f $X=-0.19 $Y=1.66 $X2=0.585 $Y2=1.885
cc_39 VPB N_B2_c_88_n 0.0341619f $X=-0.19 $Y=1.66 $X2=0.585 $Y2=1.42
cc_40 VPB N_B2_c_90_n 0.0163607f $X=-0.19 $Y=1.66 $X2=0.395 $Y2=0.34
cc_41 VPB N_B1_c_124_n 0.0332355f $X=-0.19 $Y=1.66 $X2=0.6 $Y2=0.505
cc_42 VPB B1 0.00222003f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=0.47
cc_43 VPB N_A1_c_160_n 0.0372369f $X=-0.19 $Y=1.66 $X2=0.585 $Y2=2.46
cc_44 VPB N_A1_c_161_n 0.00217948f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=0.47
cc_45 VPB N_A_222_392#_c_194_n 0.0274486f $X=-0.19 $Y=1.66 $X2=0.6 $Y2=1.33
cc_46 VPB N_A_222_392#_c_197_n 0.00156669f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_47 VPB N_VPWR_c_252_n 0.013204f $X=-0.19 $Y=1.66 $X2=0.6 $Y2=1.33
cc_48 VPB N_VPWR_c_253_n 0.0494415f $X=-0.19 $Y=1.66 $X2=0.6 $Y2=0.935
cc_49 VPB N_VPWR_c_254_n 0.00854384f $X=-0.19 $Y=1.66 $X2=0.395 $Y2=0.34
cc_50 VPB N_VPWR_c_255_n 0.0414615f $X=-0.19 $Y=1.66 $X2=0.342 $Y2=0.34
cc_51 VPB N_VPWR_c_256_n 0.0196299f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_52 VPB N_VPWR_c_251_n 0.0648288f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_53 VPB N_VPWR_c_258_n 0.0105616f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_54 VPB N_A_132_392#_c_286_n 0.0057356f $X=-0.19 $Y=1.66 $X2=0.395 $Y2=0.34
cc_55 VPB N_A_132_392#_c_287_n 0.00171072f $X=-0.19 $Y=1.66 $X2=0.395 $Y2=0.34
cc_56 VPB X 0.0604865f $X=-0.19 $Y=1.66 $X2=0.6 $Y2=1.33
cc_57 N_A2_c_58_n N_B2_c_88_n 0.0213265f $X=0.585 $Y=1.795 $X2=-0.19 $Y2=-0.245
cc_58 N_A2_c_63_n N_B2_c_88_n 0.0135242f $X=0.585 $Y=1.885 $X2=-0.19 $Y2=-0.245
cc_59 N_A2_c_61_n N_B2_M1004_g 0.0292353f $X=0.6 $Y=0.34 $X2=0 $Y2=0
cc_60 N_A2_c_58_n N_B2_c_90_n 0.0175612f $X=0.585 $Y=1.795 $X2=0 $Y2=0
cc_61 N_A2_c_63_n N_B2_c_90_n 0.00747944f $X=0.585 $Y=1.885 $X2=0 $Y2=0
cc_62 N_A2_c_63_n N_VPWR_c_253_n 0.00655454f $X=0.585 $Y=1.885 $X2=0 $Y2=0
cc_63 N_A2_c_63_n N_VPWR_c_255_n 0.0044313f $X=0.585 $Y=1.885 $X2=0 $Y2=0
cc_64 N_A2_c_63_n N_VPWR_c_251_n 0.00857176f $X=0.585 $Y=1.885 $X2=0 $Y2=0
cc_65 N_A2_c_63_n N_A_132_392#_c_288_n 0.0102221f $X=0.585 $Y=1.885 $X2=0 $Y2=0
cc_66 N_A2_c_63_n N_A_132_392#_c_287_n 0.00332677f $X=0.585 $Y=1.885 $X2=0 $Y2=0
cc_67 A2 N_A_52_123#_M1002_s 0.00167987f $X=0.155 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_68 N_A2_M1002_g N_A_52_123#_c_321_n 0.011742f $X=0.6 $Y=0.935 $X2=0 $Y2=0
cc_69 A2 N_A_52_123#_c_321_n 2.3751e-19 $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_70 N_A2_M1002_g N_A_52_123#_c_322_n 5.89712e-19 $X=0.6 $Y=0.935 $X2=0 $Y2=0
cc_71 N_A2_c_57_n N_A_52_123#_c_325_n 9.3169e-19 $X=0.585 $Y=1.42 $X2=0 $Y2=0
cc_72 N_A2_M1002_g N_A_52_123#_c_325_n 0.00748439f $X=0.6 $Y=0.935 $X2=0 $Y2=0
cc_73 A2 N_A_52_123#_c_325_n 0.0179561f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_74 N_A2_c_61_n N_A_52_123#_c_325_n 0.00159699f $X=0.6 $Y=0.34 $X2=0 $Y2=0
cc_75 A2 N_VGND_c_364_n 0.0257619f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_76 N_A2_c_61_n N_VGND_c_364_n 0.00658794f $X=0.6 $Y=0.34 $X2=0 $Y2=0
cc_77 A2 N_VGND_c_366_n 0.0285096f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_78 N_A2_c_61_n N_VGND_c_366_n 0.010364f $X=0.6 $Y=0.34 $X2=0 $Y2=0
cc_79 A2 N_VGND_c_370_n 0.0151033f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_80 N_A2_c_61_n N_VGND_c_370_n 0.0170069f $X=0.6 $Y=0.34 $X2=0 $Y2=0
cc_81 N_B2_M1004_g N_B1_c_123_n 0.0103623f $X=1.075 $Y=0.715 $X2=0 $Y2=0
cc_82 N_B2_c_88_n N_B1_c_124_n 0.0419214f $X=1.035 $Y=1.885 $X2=0 $Y2=0
cc_83 N_B2_c_90_n N_B1_c_124_n 4.10923e-19 $X=1.05 $Y=1.635 $X2=0 $Y2=0
cc_84 N_B2_M1004_g N_B1_c_125_n 0.0600955f $X=1.075 $Y=0.715 $X2=0 $Y2=0
cc_85 N_B2_c_88_n B1 4.14342e-19 $X=1.035 $Y=1.885 $X2=0 $Y2=0
cc_86 N_B2_c_90_n B1 0.0223685f $X=1.05 $Y=1.635 $X2=0 $Y2=0
cc_87 N_B2_c_88_n N_A_222_392#_c_201_n 0.0107492f $X=1.035 $Y=1.885 $X2=0 $Y2=0
cc_88 N_B2_c_90_n N_A_222_392#_c_201_n 0.00726805f $X=1.05 $Y=1.635 $X2=0 $Y2=0
cc_89 N_B2_M1004_g N_A_222_392#_c_198_n 3.18622e-19 $X=1.075 $Y=0.715 $X2=0
+ $Y2=0
cc_90 N_B2_c_90_n N_VPWR_c_253_n 0.0215684f $X=1.05 $Y=1.635 $X2=0 $Y2=0
cc_91 N_B2_c_88_n N_VPWR_c_255_n 0.00278271f $X=1.035 $Y=1.885 $X2=0 $Y2=0
cc_92 N_B2_c_88_n N_VPWR_c_251_n 0.00354253f $X=1.035 $Y=1.885 $X2=0 $Y2=0
cc_93 N_B2_c_88_n N_A_132_392#_c_288_n 2.09661e-19 $X=1.035 $Y=1.885 $X2=0 $Y2=0
cc_94 N_B2_c_90_n N_A_132_392#_c_288_n 0.0187042f $X=1.05 $Y=1.635 $X2=0 $Y2=0
cc_95 N_B2_c_88_n N_A_132_392#_c_286_n 0.0129118f $X=1.035 $Y=1.885 $X2=0 $Y2=0
cc_96 N_B2_c_88_n N_A_52_123#_c_321_n 0.00426646f $X=1.035 $Y=1.885 $X2=0 $Y2=0
cc_97 N_B2_M1004_g N_A_52_123#_c_321_n 0.0125893f $X=1.075 $Y=0.715 $X2=0 $Y2=0
cc_98 N_B2_c_90_n N_A_52_123#_c_321_n 0.0506736f $X=1.05 $Y=1.635 $X2=0 $Y2=0
cc_99 N_B2_M1004_g N_A_52_123#_c_322_n 0.00951806f $X=1.075 $Y=0.715 $X2=0 $Y2=0
cc_100 N_B2_M1004_g N_A_52_123#_c_323_n 0.00535541f $X=1.075 $Y=0.715 $X2=0
+ $Y2=0
cc_101 N_B2_M1004_g N_A_52_123#_c_325_n 6.05736e-19 $X=1.075 $Y=0.715 $X2=0
+ $Y2=0
cc_102 N_B2_c_90_n N_A_52_123#_c_325_n 0.0278161f $X=1.05 $Y=1.635 $X2=0 $Y2=0
cc_103 N_B2_M1004_g N_VGND_c_364_n 0.00384771f $X=1.075 $Y=0.715 $X2=0 $Y2=0
cc_104 N_B2_M1004_g N_VGND_c_368_n 0.00522295f $X=1.075 $Y=0.715 $X2=0 $Y2=0
cc_105 N_B2_M1004_g N_VGND_c_370_n 0.00537853f $X=1.075 $Y=0.715 $X2=0 $Y2=0
cc_106 N_B1_c_125_n N_A1_c_159_n 0.0232104f $X=1.467 $Y=1.11 $X2=-0.19
+ $Y2=-0.245
cc_107 N_B1_c_123_n N_A1_c_160_n 0.00726285f $X=1.5 $Y=1.47 $X2=0 $Y2=0
cc_108 N_B1_c_124_n N_A1_c_160_n 0.0479932f $X=1.515 $Y=1.885 $X2=0 $Y2=0
cc_109 N_B1_c_126_n N_A1_c_160_n 0.00974511f $X=1.467 $Y=1.26 $X2=0 $Y2=0
cc_110 B1 N_A1_c_160_n 0.00230326f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_111 N_B1_c_123_n N_A1_c_161_n 6.90997e-19 $X=1.5 $Y=1.47 $X2=0 $Y2=0
cc_112 N_B1_c_124_n N_A1_c_161_n 3.55575e-19 $X=1.515 $Y=1.885 $X2=0 $Y2=0
cc_113 B1 N_A1_c_161_n 0.024799f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_114 N_B1_c_124_n N_A_222_392#_c_204_n 0.0167844f $X=1.515 $Y=1.885 $X2=0
+ $Y2=0
cc_115 B1 N_A_222_392#_c_204_n 0.0244721f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_116 N_B1_c_124_n N_A_222_392#_c_198_n 0.00388761f $X=1.515 $Y=1.885 $X2=0
+ $Y2=0
cc_117 N_B1_c_125_n N_A_222_392#_c_198_n 0.00452641f $X=1.467 $Y=1.11 $X2=0
+ $Y2=0
cc_118 N_B1_c_126_n N_A_222_392#_c_198_n 0.00482129f $X=1.467 $Y=1.26 $X2=0
+ $Y2=0
cc_119 B1 N_A_222_392#_c_198_n 0.0164626f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_120 N_B1_c_124_n N_VPWR_c_255_n 0.00278271f $X=1.515 $Y=1.885 $X2=0 $Y2=0
cc_121 N_B1_c_124_n N_VPWR_c_251_n 0.00355001f $X=1.515 $Y=1.885 $X2=0 $Y2=0
cc_122 N_B1_c_124_n N_A_132_392#_c_286_n 0.0145199f $X=1.515 $Y=1.885 $X2=0
+ $Y2=0
cc_123 N_B1_c_123_n N_A_52_123#_c_321_n 0.00113592f $X=1.5 $Y=1.47 $X2=0 $Y2=0
cc_124 N_B1_c_126_n N_A_52_123#_c_321_n 0.00280224f $X=1.467 $Y=1.26 $X2=0 $Y2=0
cc_125 N_B1_c_125_n N_A_52_123#_c_322_n 0.00585891f $X=1.467 $Y=1.11 $X2=0 $Y2=0
cc_126 N_B1_c_125_n N_A_52_123#_c_324_n 0.016242f $X=1.467 $Y=1.11 $X2=0 $Y2=0
cc_127 N_B1_c_125_n N_VGND_c_368_n 0.00399513f $X=1.467 $Y=1.11 $X2=0 $Y2=0
cc_128 N_B1_c_125_n N_VGND_c_370_n 0.00537853f $X=1.467 $Y=1.11 $X2=0 $Y2=0
cc_129 N_A1_c_160_n N_A_222_392#_c_194_n 0.0362092f $X=2.055 $Y=1.885 $X2=0
+ $Y2=0
cc_130 N_A1_c_161_n N_A_222_392#_c_194_n 0.00134044f $X=2.13 $Y=1.515 $X2=0
+ $Y2=0
cc_131 N_A1_c_160_n N_A_222_392#_M1008_g 0.00183582f $X=2.055 $Y=1.885 $X2=0
+ $Y2=0
cc_132 N_A1_c_160_n N_A_222_392#_c_204_n 0.0171902f $X=2.055 $Y=1.885 $X2=0
+ $Y2=0
cc_133 N_A1_c_161_n N_A_222_392#_c_204_n 0.0206885f $X=2.13 $Y=1.515 $X2=0 $Y2=0
cc_134 N_A1_c_159_n N_A_222_392#_c_196_n 0.00648271f $X=1.865 $Y=1.11 $X2=0
+ $Y2=0
cc_135 N_A1_c_160_n N_A_222_392#_c_196_n 0.0153045f $X=2.055 $Y=1.885 $X2=0
+ $Y2=0
cc_136 N_A1_c_161_n N_A_222_392#_c_196_n 0.0247243f $X=2.13 $Y=1.515 $X2=0 $Y2=0
cc_137 N_A1_c_160_n N_A_222_392#_c_197_n 0.00812537f $X=2.055 $Y=1.885 $X2=0
+ $Y2=0
cc_138 N_A1_c_161_n N_A_222_392#_c_197_n 0.0277121f $X=2.13 $Y=1.515 $X2=0 $Y2=0
cc_139 N_A1_c_159_n N_A_222_392#_c_198_n 0.0110654f $X=1.865 $Y=1.11 $X2=0 $Y2=0
cc_140 N_A1_c_160_n N_A_222_392#_c_198_n 0.00186216f $X=2.055 $Y=1.885 $X2=0
+ $Y2=0
cc_141 N_A1_c_160_n N_VPWR_c_254_n 0.00391322f $X=2.055 $Y=1.885 $X2=0 $Y2=0
cc_142 N_A1_c_160_n N_VPWR_c_255_n 0.0044313f $X=2.055 $Y=1.885 $X2=0 $Y2=0
cc_143 N_A1_c_160_n N_VPWR_c_251_n 0.00855581f $X=2.055 $Y=1.885 $X2=0 $Y2=0
cc_144 N_A1_c_160_n N_A_132_392#_c_286_n 0.00350048f $X=2.055 $Y=1.885 $X2=0
+ $Y2=0
cc_145 N_A1_c_160_n N_A_132_392#_c_295_n 0.00610669f $X=2.055 $Y=1.885 $X2=0
+ $Y2=0
cc_146 N_A1_c_159_n N_A_52_123#_c_324_n 0.01135f $X=1.865 $Y=1.11 $X2=0 $Y2=0
cc_147 N_A1_c_160_n N_A_52_123#_c_324_n 7.37405e-19 $X=2.055 $Y=1.885 $X2=0
+ $Y2=0
cc_148 N_A1_c_159_n N_VGND_c_365_n 0.00705117f $X=1.865 $Y=1.11 $X2=0 $Y2=0
cc_149 N_A1_c_159_n N_VGND_c_368_n 0.00399513f $X=1.865 $Y=1.11 $X2=0 $Y2=0
cc_150 N_A1_c_159_n N_VGND_c_370_n 0.00537853f $X=1.865 $Y=1.11 $X2=0 $Y2=0
cc_151 N_A_222_392#_c_204_n N_VPWR_M1001_d 0.0160249f $X=2.505 $Y=2.055 $X2=0
+ $Y2=0
cc_152 N_A_222_392#_c_197_n N_VPWR_M1001_d 0.00193534f $X=2.67 $Y=1.465 $X2=0
+ $Y2=0
cc_153 N_A_222_392#_c_194_n N_VPWR_c_254_n 0.021624f $X=2.785 $Y=1.765 $X2=0
+ $Y2=0
cc_154 N_A_222_392#_c_204_n N_VPWR_c_254_n 0.0402772f $X=2.505 $Y=2.055 $X2=0
+ $Y2=0
cc_155 N_A_222_392#_c_194_n N_VPWR_c_256_n 0.00413917f $X=2.785 $Y=1.765 $X2=0
+ $Y2=0
cc_156 N_A_222_392#_c_194_n N_VPWR_c_251_n 0.00821431f $X=2.785 $Y=1.765 $X2=0
+ $Y2=0
cc_157 N_A_222_392#_c_204_n N_A_132_392#_M1006_d 0.00941364f $X=2.505 $Y=2.055
+ $X2=0 $Y2=0
cc_158 N_A_222_392#_c_201_n N_A_132_392#_c_288_n 0.0519649f $X=1.26 $Y=2.135
+ $X2=0 $Y2=0
cc_159 N_A_222_392#_M1003_d N_A_132_392#_c_286_n 0.00229612f $X=1.11 $Y=1.96
+ $X2=0 $Y2=0
cc_160 N_A_222_392#_c_201_n N_A_132_392#_c_286_n 0.0174007f $X=1.26 $Y=2.135
+ $X2=0 $Y2=0
cc_161 N_A_222_392#_c_204_n N_A_132_392#_c_295_n 0.0234793f $X=2.505 $Y=2.055
+ $X2=0 $Y2=0
cc_162 N_A_222_392#_c_194_n X 0.0242695f $X=2.785 $Y=1.765 $X2=0 $Y2=0
cc_163 N_A_222_392#_M1008_g X 0.0214406f $X=2.875 $Y=0.74 $X2=0 $Y2=0
cc_164 N_A_222_392#_c_204_n X 0.0140085f $X=2.505 $Y=2.055 $X2=0 $Y2=0
cc_165 N_A_222_392#_c_196_n X 0.00962585f $X=2.505 $Y=1.095 $X2=0 $Y2=0
cc_166 N_A_222_392#_c_197_n X 0.0603011f $X=2.67 $Y=1.465 $X2=0 $Y2=0
cc_167 N_A_222_392#_c_196_n N_A_52_123#_M1005_d 0.00358528f $X=2.505 $Y=1.095
+ $X2=0 $Y2=0
cc_168 N_A_222_392#_c_201_n N_A_52_123#_c_321_n 0.00236654f $X=1.26 $Y=2.135
+ $X2=0 $Y2=0
cc_169 N_A_222_392#_c_198_n N_A_52_123#_c_321_n 0.00373163f $X=1.65 $Y=0.885
+ $X2=0 $Y2=0
cc_170 N_A_222_392#_c_198_n N_A_52_123#_c_322_n 0.0218843f $X=1.65 $Y=0.885
+ $X2=0 $Y2=0
cc_171 N_A_222_392#_M1000_d N_A_52_123#_c_324_n 0.00177578f $X=1.51 $Y=0.395
+ $X2=0 $Y2=0
cc_172 N_A_222_392#_c_196_n N_A_52_123#_c_324_n 0.014733f $X=2.505 $Y=1.095
+ $X2=0 $Y2=0
cc_173 N_A_222_392#_c_198_n N_A_52_123#_c_324_n 0.0162725f $X=1.65 $Y=0.885
+ $X2=0 $Y2=0
cc_174 N_A_222_392#_c_196_n N_VGND_M1008_s 0.00345306f $X=2.505 $Y=1.095 $X2=0
+ $Y2=0
cc_175 N_A_222_392#_c_194_n N_VGND_c_365_n 9.99993e-19 $X=2.785 $Y=1.765 $X2=0
+ $Y2=0
cc_176 N_A_222_392#_M1008_g N_VGND_c_365_n 0.00698798f $X=2.875 $Y=0.74 $X2=0
+ $Y2=0
cc_177 N_A_222_392#_c_196_n N_VGND_c_365_n 0.0222869f $X=2.505 $Y=1.095 $X2=0
+ $Y2=0
cc_178 N_A_222_392#_M1008_g N_VGND_c_369_n 0.00434272f $X=2.875 $Y=0.74 $X2=0
+ $Y2=0
cc_179 N_A_222_392#_M1008_g N_VGND_c_370_n 0.00828906f $X=2.875 $Y=0.74 $X2=0
+ $Y2=0
cc_180 N_VPWR_c_253_n N_A_132_392#_c_288_n 0.0613781f $X=0.36 $Y=2.135 $X2=0
+ $Y2=0
cc_181 N_VPWR_c_254_n N_A_132_392#_c_286_n 0.01232f $X=2.56 $Y=2.43 $X2=0 $Y2=0
cc_182 N_VPWR_c_255_n N_A_132_392#_c_286_n 0.0727832f $X=2.165 $Y=3.33 $X2=0
+ $Y2=0
cc_183 N_VPWR_c_251_n N_A_132_392#_c_286_n 0.0404277f $X=3.12 $Y=3.33 $X2=0
+ $Y2=0
cc_184 N_VPWR_c_253_n N_A_132_392#_c_287_n 0.012272f $X=0.36 $Y=2.135 $X2=0
+ $Y2=0
cc_185 N_VPWR_c_255_n N_A_132_392#_c_287_n 0.017869f $X=2.165 $Y=3.33 $X2=0
+ $Y2=0
cc_186 N_VPWR_c_251_n N_A_132_392#_c_287_n 0.00965079f $X=3.12 $Y=3.33 $X2=0
+ $Y2=0
cc_187 N_VPWR_c_254_n X 0.0477818f $X=2.56 $Y=2.43 $X2=0 $Y2=0
cc_188 N_VPWR_c_256_n X 0.0146357f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_189 N_VPWR_c_251_n X 0.0121141f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_190 X N_VGND_c_365_n 0.0182902f $X=3.035 $Y=0.47 $X2=0 $Y2=0
cc_191 X N_VGND_c_369_n 0.0145639f $X=3.035 $Y=0.47 $X2=0 $Y2=0
cc_192 X N_VGND_c_370_n 0.0119984f $X=3.035 $Y=0.47 $X2=0 $Y2=0
cc_193 N_A_52_123#_c_321_n N_VGND_M1002_d 0.00205163f $X=1.115 $Y=1.215
+ $X2=-0.19 $Y2=-0.245
cc_194 N_A_52_123#_c_321_n N_VGND_c_364_n 0.0172284f $X=1.115 $Y=1.215 $X2=0
+ $Y2=0
cc_195 N_A_52_123#_c_323_n N_VGND_c_364_n 0.011275f $X=1.285 $Y=0.5 $X2=0 $Y2=0
cc_196 N_A_52_123#_c_324_n N_VGND_c_365_n 0.0164198f $X=2.08 $Y=0.54 $X2=0 $Y2=0
cc_197 N_A_52_123#_c_323_n N_VGND_c_368_n 0.00679203f $X=1.285 $Y=0.5 $X2=0
+ $Y2=0
cc_198 N_A_52_123#_c_324_n N_VGND_c_368_n 0.0353785f $X=2.08 $Y=0.54 $X2=0 $Y2=0
cc_199 N_A_52_123#_c_323_n N_VGND_c_370_n 0.00615299f $X=1.285 $Y=0.5 $X2=0
+ $Y2=0
cc_200 N_A_52_123#_c_324_n N_VGND_c_370_n 0.033495f $X=2.08 $Y=0.54 $X2=0 $Y2=0
cc_201 N_A_52_123#_c_322_n A_230_79# 0.00395173f $X=1.2 $Y=1.13 $X2=-0.19
+ $Y2=-0.245
cc_202 N_A_52_123#_c_324_n A_230_79# 6.79616e-19 $X=2.08 $Y=0.54 $X2=-0.19
+ $Y2=-0.245
