* File: sky130_fd_sc_hs__edfxtp_1.spice
* Created: Tue Sep  1 20:04:27 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hs__edfxtp_1.pex.spice"
.subckt sky130_fd_sc_hs__edfxtp_1  VNB VPB D DE CLK VPWR Q VGND
* 
* VGND	VGND
* Q	Q
* VPWR	VPWR
* CLK	CLK
* DE	DE
* D	D
* VPB	VPB
* VNB	VNB
MM1013 A_131_74# N_D_M1013_g N_A_27_508#_M1013_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.0504 AS=0.1197 PD=0.66 PS=1.41 NRD=18.564 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1009 N_VGND_M1009_d N_DE_M1009_g A_131_74# VNB NLOWVT L=0.15 W=0.42 AD=0.1176
+ AS=0.0504 PD=1.4 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75000.6 SB=75000.2
+ A=0.063 P=1.14 MULT=1
MM1014 N_VGND_M1014_d N_DE_M1014_g N_A_159_446#_M1014_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.0588 AS=0.1176 PD=0.7 PS=1.4 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2 SB=75001
+ A=0.063 P=1.14 MULT=1
MM1023 A_491_87# N_A_159_446#_M1023_g N_VGND_M1014_d VNB NLOWVT L=0.15 W=0.42
+ AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1025 N_A_27_508#_M1025_d N_A_533_61#_M1025_g A_491_87# VNB NLOWVT L=0.15
+ W=0.42 AD=0.1197 AS=0.0441 PD=1.41 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75001
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1017 N_A_763_74#_M1017_d N_CLK_M1017_g N_VGND_M1017_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.2035 AS=0.2109 PD=2.03 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1033 N_A_958_74#_M1033_d N_A_763_74#_M1033_g N_VGND_M1033_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.2109 AS=0.2072 PD=2.05 PS=2.04 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1028 N_A_1156_90#_M1028_d N_A_763_74#_M1028_g N_A_27_508#_M1028_s VNB NLOWVT
+ L=0.15 W=0.42 AD=0.17115 AS=0.1197 PD=1.235 PS=1.41 NRD=134.28 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75002.3 A=0.063 P=1.14 MULT=1
MM1031 A_1349_90# N_A_958_74#_M1031_g N_A_1156_90#_M1028_d VNB NLOWVT L=0.15
+ W=0.42 AD=0.063 AS=0.17115 PD=0.72 PS=1.235 NRD=27.132 NRS=18.564 M=1 R=2.8
+ SA=75001.2 SB=75001.3 A=0.063 P=1.14 MULT=1
MM1001 N_VGND_M1001_d N_A_1409_64#_M1001_g A_1349_90# VNB NLOWVT L=0.15 W=0.42
+ AD=0.109992 AS=0.063 PD=0.92717 PS=0.72 NRD=0 NRS=27.132 M=1 R=2.8 SA=75001.6
+ SB=75000.9 A=0.063 P=1.14 MULT=1
MM1008 N_A_1409_64#_M1008_d N_A_1156_90#_M1008_g N_VGND_M1001_d VNB NLOWVT
+ L=0.15 W=0.64 AD=0.1824 AS=0.167608 PD=1.85 PS=1.41283 NRD=0 NRS=46.872 M=1
+ R=4.26667 SA=75001.6 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1018 A_1797_74# N_A_1409_64#_M1018_g N_VGND_M1018_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1258 AS=0.2109 PD=1.08 PS=2.05 NRD=18.648 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75001.8 A=0.111 P=1.78 MULT=1
MM1032 N_A_1895_74#_M1032_d N_A_958_74#_M1032_g A_1797_74# VNB NLOWVT L=0.15
+ W=0.74 AD=0.154634 AS=0.1258 PD=1.40345 PS=1.08 NRD=0 NRS=18.648 M=1 R=4.93333
+ SA=75000.7 SB=75001.3 A=0.111 P=1.78 MULT=1
MM1011 A_1997_74# N_A_763_74#_M1011_g N_A_1895_74#_M1032_d VNB NLOWVT L=0.15
+ W=0.42 AD=0.0504 AS=0.0877655 PD=0.66 PS=0.796552 NRD=18.564 NRS=22.848 M=1
+ R=2.8 SA=75001.2 SB=75001.7 A=0.063 P=1.14 MULT=1
MM1005 N_VGND_M1005_d N_A_533_61#_M1005_g A_1997_74# VNB NLOWVT L=0.15 W=0.42
+ AD=0.20055 AS=0.0504 PD=1.375 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75001.6
+ SB=75001.3 A=0.063 P=1.14 MULT=1
MM1007 N_A_533_61#_M1007_d N_A_1895_74#_M1007_g N_VGND_M1005_d VNB NLOWVT L=0.15
+ W=0.42 AD=0.1197 AS=0.20055 PD=1.41 PS=1.375 NRD=0 NRS=0 M=1 R=2.8 SA=75002.7
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1022 N_VGND_M1022_d N_A_1895_74#_M1022_g N_Q_M1022_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.2627 AS=0.2109 PD=2.19 PS=2.05 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75000.3 A=0.111 P=1.78 MULT=1
MM1020 A_114_508# N_D_M1020_g N_A_27_508#_M1020_s VPB PSHORT L=0.15 W=0.42
+ AD=0.0504 AS=0.1197 PD=0.66 PS=1.41 NRD=30.4759 NRS=4.6886 M=1 R=2.8
+ SA=75000.2 SB=75000.6 A=0.063 P=1.14 MULT=1
MM1003 N_VPWR_M1003_d N_A_159_446#_M1003_g A_114_508# VPB PSHORT L=0.15 W=0.42
+ AD=0.1239 AS=0.0504 PD=1.43 PS=0.66 NRD=4.6886 NRS=30.4759 M=1 R=2.8
+ SA=75000.6 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1012 N_VPWR_M1012_d N_DE_M1012_g N_A_159_446#_M1012_s VPB PSHORT L=0.15 W=0.64
+ AD=0.1696 AS=0.1888 PD=1.41283 PS=1.87 NRD=73.8553 NRS=3.0732 M=1 R=4.26667
+ SA=75000.2 SB=75000.9 A=0.096 P=1.58 MULT=1
MM1026 A_554_436# N_DE_M1026_g N_VPWR_M1012_d VPB PSHORT L=0.15 W=0.42 AD=0.0504
+ AS=0.1113 PD=0.66 PS=0.92717 NRD=30.4759 NRS=4.6886 M=1 R=2.8 SA=75000.9
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1016 N_A_27_508#_M1016_d N_A_533_61#_M1016_g A_554_436# VPB PSHORT L=0.15
+ W=0.42 AD=0.1155 AS=0.0504 PD=1.39 PS=0.66 NRD=4.6886 NRS=30.4759 M=1 R=2.8
+ SA=75001.3 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1002 N_A_763_74#_M1002_d N_CLK_M1002_g N_VPWR_M1002_s VPB PSHORT L=0.15 W=1.12
+ AD=0.308 AS=0.3136 PD=2.79 PS=2.8 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75000.2 A=0.168 P=2.54 MULT=1
MM1019 N_A_958_74#_M1019_d N_A_763_74#_M1019_g N_VPWR_M1019_s VPB PSHORT L=0.15
+ W=1.12 AD=0.308 AS=0.308 PD=2.79 PS=2.79 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75000.2 A=0.168 P=2.54 MULT=1
MM1000 N_A_1156_90#_M1000_d N_A_958_74#_M1000_g N_A_27_508#_M1000_s VPB PSHORT
+ L=0.15 W=0.42 AD=0.063 AS=0.1176 PD=0.72 PS=1.4 NRD=4.6886 NRS=4.6886 M=1
+ R=2.8 SA=75000.2 SB=75001.6 A=0.063 P=1.14 MULT=1
MM1004 A_1382_508# N_A_763_74#_M1004_g N_A_1156_90#_M1000_d VPB PSHORT L=0.15
+ W=0.42 AD=0.07455 AS=0.063 PD=0.775 PS=0.72 NRD=57.4452 NRS=4.6886 M=1 R=2.8
+ SA=75000.7 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1030 N_VPWR_M1030_d N_A_1409_64#_M1030_g A_1382_508# VPB PSHORT L=0.15 W=0.42
+ AD=0.0979417 AS=0.07455 PD=0.886667 PS=0.775 NRD=9.3772 NRS=57.4452 M=1 R=2.8
+ SA=75001.2 SB=75000.6 A=0.063 P=1.14 MULT=1
MM1015 N_A_1409_64#_M1015_d N_A_1156_90#_M1015_g N_VPWR_M1030_d VPB PSHORT
+ L=0.15 W=0.84 AD=0.2478 AS=0.195883 PD=2.27 PS=1.77333 NRD=2.3443 NRS=23.443
+ M=1 R=5.6 SA=75000.8 SB=75000.2 A=0.126 P=1.98 MULT=1
MM1029 A_1794_392# N_A_1409_64#_M1029_g N_VPWR_M1029_s VPB PSHORT L=0.15 W=1
+ AD=0.3925 AS=0.295 PD=1.785 PS=2.59 NRD=66.4678 NRS=1.9503 M=1 R=6.66667
+ SA=75000.2 SB=75001.8 A=0.15 P=2.3 MULT=1
MM1021 N_A_1895_74#_M1021_d N_A_763_74#_M1021_g A_1794_392# VPB PSHORT L=0.15
+ W=1 AD=0.234366 AS=0.3925 PD=1.9507 PS=1.785 NRD=1.9503 NRS=66.4678 M=1
+ R=6.66667 SA=75001.2 SB=75000.9 A=0.15 P=2.3 MULT=1
MM1006 A_2088_502# N_A_958_74#_M1006_g N_A_1895_74#_M1021_d VPB PSHORT L=0.15
+ W=0.42 AD=0.0567 AS=0.0984338 PD=0.69 PS=0.819296 NRD=37.5088 NRS=45.7237 M=1
+ R=2.8 SA=75001.7 SB=75001.3 A=0.063 P=1.14 MULT=1
MM1024 N_VPWR_M1024_d N_A_533_61#_M1024_g A_2088_502# VPB PSHORT L=0.15 W=0.42
+ AD=0.116292 AS=0.0567 PD=0.950943 PS=0.69 NRD=65.6601 NRS=37.5088 M=1 R=2.8
+ SA=75002.1 SB=75000.9 A=0.063 P=1.14 MULT=1
MM1027 N_A_533_61#_M1027_d N_A_1895_74#_M1027_g N_VPWR_M1024_d VPB PSHORT L=0.15
+ W=0.64 AD=0.176 AS=0.177208 PD=1.83 PS=1.44906 NRD=3.0732 NRS=43.0839 M=1
+ R=4.26667 SA=75001.9 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1010 N_VPWR_M1010_d N_A_1895_74#_M1010_g N_Q_M1010_s VPB PSHORT L=0.15 W=1.12
+ AD=0.3192 AS=0.308 PD=2.81 PS=2.79 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75000.2 A=0.168 P=2.54 MULT=1
DX34_noxref VNB VPB NWDIODE A=24.8976 P=30.56
c_143 VNB 0 4.56061e-19 $X=0 $Y=0
*
.include "sky130_fd_sc_hs__edfxtp_1.pxi.spice"
*
.ends
*
*
