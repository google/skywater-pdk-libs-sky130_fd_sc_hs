* File: sky130_fd_sc_hs__a41oi_4.pex.spice
* Created: Tue Sep  1 19:54:28 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HS__A41OI_4%B1 3 5 7 10 12 14 15 17 18 19 20 22 23 24 25
+ 38
c78 20 0 4.79772e-20 $X=1.955 $Y=1.765
c79 19 0 1.97368e-19 $X=1.595 $Y=1.64
r80 37 39 29.8915 $w=3.87e-07 $l=2.4e-07 $layer=POLY_cond $X=1.265 $Y=1.557
+ $X2=1.505 $Y2=1.557
r81 37 38 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.265
+ $Y=1.515 $X2=1.265 $Y2=1.515
r82 35 37 32.3824 $w=3.87e-07 $l=2.6e-07 $layer=POLY_cond $X=1.005 $Y=1.557
+ $X2=1.265 $Y2=1.557
r83 34 35 1.24548 $w=3.87e-07 $l=1e-08 $layer=POLY_cond $X=0.995 $Y=1.557
+ $X2=1.005 $Y2=1.557
r84 32 34 51.0646 $w=3.87e-07 $l=4.1e-07 $layer=POLY_cond $X=0.585 $Y=1.557
+ $X2=0.995 $Y2=1.557
r85 32 33 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=0.585
+ $Y=1.515 $X2=0.585 $Y2=1.515
r86 30 32 9.34109 $w=3.87e-07 $l=7.5e-08 $layer=POLY_cond $X=0.51 $Y=1.557
+ $X2=0.585 $Y2=1.557
r87 29 30 1.86822 $w=3.87e-07 $l=1.5e-08 $layer=POLY_cond $X=0.495 $Y=1.557
+ $X2=0.51 $Y2=1.557
r88 25 38 1.74206 $w=4.28e-07 $l=6.5e-08 $layer=LI1_cond $X=1.2 $Y=1.565
+ $X2=1.265 $Y2=1.565
r89 24 25 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=0.72 $Y=1.565
+ $X2=1.2 $Y2=1.565
r90 24 33 3.61813 $w=4.28e-07 $l=1.35e-07 $layer=LI1_cond $X=0.72 $Y=1.565
+ $X2=0.585 $Y2=1.565
r91 23 33 9.24634 $w=4.28e-07 $l=3.45e-07 $layer=LI1_cond $X=0.24 $Y=1.565
+ $X2=0.585 $Y2=1.565
r92 20 22 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.955 $Y=1.765
+ $X2=1.955 $Y2=2.4
r93 19 39 29.9996 $w=3.87e-07 $l=1.2478e-07 $layer=POLY_cond $X=1.595 $Y=1.64
+ $X2=1.505 $Y2=1.557
r94 18 20 26.9307 $w=1.5e-07 $l=1.63936e-07 $layer=POLY_cond $X=1.865 $Y=1.64
+ $X2=1.955 $Y2=1.765
r95 18 19 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=1.865 $Y=1.64
+ $X2=1.595 $Y2=1.64
r96 15 39 25.0561 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=1.505 $Y=1.765
+ $X2=1.505 $Y2=1.557
r97 15 17 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.505 $Y=1.765
+ $X2=1.505 $Y2=2.4
r98 12 35 25.0561 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=1.005 $Y=1.765
+ $X2=1.005 $Y2=1.557
r99 12 14 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.005 $Y=1.765
+ $X2=1.005 $Y2=2.4
r100 8 34 25.0561 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.995 $Y=1.35
+ $X2=0.995 $Y2=1.557
r101 8 10 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=0.995 $Y=1.35
+ $X2=0.995 $Y2=0.74
r102 5 30 25.0561 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=0.51 $Y=1.765
+ $X2=0.51 $Y2=1.557
r103 5 7 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.51 $Y=1.765
+ $X2=0.51 $Y2=2.4
r104 1 29 25.0561 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.495 $Y=1.35
+ $X2=0.495 $Y2=1.557
r105 1 3 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=0.495 $Y=1.35
+ $X2=0.495 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HS__A41OI_4%A1 1 3 4 5 6 8 9 11 12 14 15 17 18 20 21 23
+ 24 26 27 28 39 42
c108 39 0 4.79772e-20 $X=3.13 $Y=1.515
c109 18 0 1.42322e-19 $X=3.405 $Y=1.765
c110 5 0 3.74663e-19 $X=2.06 $Y=1.28
r111 41 42 27.3753 $w=4.93e-07 $l=2.8e-07 $layer=POLY_cond $X=3.405 $Y=1.485
+ $X2=3.685 $Y2=1.485
r112 40 41 14.6653 $w=4.93e-07 $l=1.5e-07 $layer=POLY_cond $X=3.255 $Y=1.485
+ $X2=3.405 $Y2=1.485
r113 38 40 12.2211 $w=4.93e-07 $l=1.25e-07 $layer=POLY_cond $X=3.13 $Y=1.485
+ $X2=3.255 $Y2=1.485
r114 38 39 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=3.13
+ $Y=1.515 $X2=3.13 $Y2=1.515
r115 36 38 17.1095 $w=4.93e-07 $l=1.75e-07 $layer=POLY_cond $X=2.955 $Y=1.485
+ $X2=3.13 $Y2=1.485
r116 35 36 45.9513 $w=4.93e-07 $l=4.7e-07 $layer=POLY_cond $X=2.485 $Y=1.485
+ $X2=2.955 $Y2=1.485
r117 33 35 3.42191 $w=4.93e-07 $l=3.5e-08 $layer=POLY_cond $X=2.45 $Y=1.485
+ $X2=2.485 $Y2=1.485
r118 33 34 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=2.45
+ $Y=1.515 $X2=2.45 $Y2=1.515
r119 31 33 4.39959 $w=4.93e-07 $l=4.5e-08 $layer=POLY_cond $X=2.405 $Y=1.485
+ $X2=2.45 $Y2=1.485
r120 28 39 0.26801 $w=4.28e-07 $l=1e-08 $layer=LI1_cond $X=3.12 $Y=1.565
+ $X2=3.13 $Y2=1.565
r121 27 28 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=2.64 $Y=1.565
+ $X2=3.12 $Y2=1.565
r122 27 34 5.09219 $w=4.28e-07 $l=1.9e-07 $layer=LI1_cond $X=2.64 $Y=1.565
+ $X2=2.45 $Y2=1.565
r123 24 42 21.998 $w=4.93e-07 $l=3.76032e-07 $layer=POLY_cond $X=3.91 $Y=1.765
+ $X2=3.685 $Y2=1.485
r124 24 26 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.91 $Y=1.765
+ $X2=3.91 $Y2=2.4
r125 21 42 31.0522 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=3.685 $Y=1.205
+ $X2=3.685 $Y2=1.485
r126 21 23 149.42 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=3.685 $Y=1.205
+ $X2=3.685 $Y2=0.74
r127 18 41 31.0522 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=3.405 $Y=1.765
+ $X2=3.405 $Y2=1.485
r128 18 20 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.405 $Y=1.765
+ $X2=3.405 $Y2=2.4
r129 15 40 31.0522 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=3.255 $Y=1.205
+ $X2=3.255 $Y2=1.485
r130 15 17 149.42 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=3.255 $Y=1.205
+ $X2=3.255 $Y2=0.74
r131 12 36 31.0522 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=2.955 $Y=1.765
+ $X2=2.955 $Y2=1.485
r132 12 14 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.955 $Y=1.765
+ $X2=2.955 $Y2=2.4
r133 9 35 31.0522 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=2.485 $Y=1.205
+ $X2=2.485 $Y2=1.485
r134 9 11 149.42 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=2.485 $Y=1.205
+ $X2=2.485 $Y2=0.74
r135 6 31 31.0522 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=2.405 $Y=1.765
+ $X2=2.405 $Y2=1.485
r136 6 8 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.405 $Y=1.765
+ $X2=2.405 $Y2=2.4
r137 4 31 37.346 $w=4.93e-07 $l=2.58118e-07 $layer=POLY_cond $X=2.285 $Y=1.28
+ $X2=2.405 $Y2=1.485
r138 4 5 115.372 $w=1.5e-07 $l=2.25e-07 $layer=POLY_cond $X=2.285 $Y=1.28
+ $X2=2.06 $Y2=1.28
r139 1 5 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.985 $Y=1.205
+ $X2=2.06 $Y2=1.28
r140 1 3 149.42 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=1.985 $Y=1.205
+ $X2=1.985 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HS__A41OI_4%A2 1 3 4 6 7 9 10 12 13 15 16 18 19 21 22 24
+ 27 30 31 44 46 53
c91 53 0 1.1015e-19 $X=4.675 $Y=1.55
c92 46 0 1.45948e-19 $X=4.445 $Y=1.55
c93 44 0 2.95129e-19 $X=5.545 $Y=1.485
c94 16 0 5.93691e-20 $X=5.32 $Y=1.765
c95 1 0 1.63532e-19 $X=4.185 $Y=1.205
r96 41 42 23.6954 $w=4.17e-07 $l=2.05e-07 $layer=POLY_cond $X=5.115 $Y=1.485
+ $X2=5.32 $Y2=1.485
r97 40 41 28.3189 $w=4.17e-07 $l=2.45e-07 $layer=POLY_cond $X=4.87 $Y=1.485
+ $X2=5.115 $Y2=1.485
r98 39 40 21.3837 $w=4.17e-07 $l=1.85e-07 $layer=POLY_cond $X=4.685 $Y=1.485
+ $X2=4.87 $Y2=1.485
r99 38 46 0.260017 $w=4.58e-07 $l=1e-08 $layer=LI1_cond $X=4.435 $Y=1.55
+ $X2=4.445 $Y2=1.55
r100 37 39 28.8969 $w=4.17e-07 $l=2.5e-07 $layer=POLY_cond $X=4.435 $Y=1.485
+ $X2=4.685 $Y2=1.485
r101 37 38 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.435
+ $Y=1.485 $X2=4.435 $Y2=1.485
r102 35 37 8.66906 $w=4.17e-07 $l=7.5e-08 $layer=POLY_cond $X=4.36 $Y=1.485
+ $X2=4.435 $Y2=1.485
r103 31 53 3.96409 $w=4.58e-07 $l=1.15e-07 $layer=LI1_cond $X=4.56 $Y=1.55
+ $X2=4.675 $Y2=1.55
r104 31 46 2.9902 $w=4.58e-07 $l=1.15e-07 $layer=LI1_cond $X=4.56 $Y=1.55
+ $X2=4.445 $Y2=1.55
r105 30 38 9.23061 $w=4.58e-07 $l=3.55e-07 $layer=LI1_cond $X=4.08 $Y=1.55
+ $X2=4.435 $Y2=1.55
r106 28 44 10.4029 $w=4.17e-07 $l=9e-08 $layer=POLY_cond $X=5.455 $Y=1.485
+ $X2=5.545 $Y2=1.485
r107 28 42 15.6043 $w=4.17e-07 $l=1.35e-07 $layer=POLY_cond $X=5.455 $Y=1.485
+ $X2=5.32 $Y2=1.485
r108 27 53 27.2396 $w=3.28e-07 $l=7.8e-07 $layer=LI1_cond $X=5.455 $Y=1.485
+ $X2=4.675 $Y2=1.485
r109 27 28 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.455
+ $Y=1.485 $X2=5.455 $Y2=1.485
r110 22 44 31.7866 $w=4.17e-07 $l=3.94208e-07 $layer=POLY_cond $X=5.82 $Y=1.765
+ $X2=5.545 $Y2=1.485
r111 22 24 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=5.82 $Y=1.765
+ $X2=5.82 $Y2=2.4
r112 19 44 26.8826 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=5.545 $Y=1.205
+ $X2=5.545 $Y2=1.485
r113 19 21 149.42 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=5.545 $Y=1.205
+ $X2=5.545 $Y2=0.74
r114 16 42 26.8826 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=5.32 $Y=1.765
+ $X2=5.32 $Y2=1.485
r115 16 18 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=5.32 $Y=1.765
+ $X2=5.32 $Y2=2.4
r116 13 41 26.8826 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=5.115 $Y=1.205
+ $X2=5.115 $Y2=1.485
r117 13 15 149.42 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=5.115 $Y=1.205
+ $X2=5.115 $Y2=0.74
r118 10 40 26.8826 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=4.87 $Y=1.765
+ $X2=4.87 $Y2=1.485
r119 10 12 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=4.87 $Y=1.765
+ $X2=4.87 $Y2=2.4
r120 7 39 26.8826 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=4.685 $Y=1.205
+ $X2=4.685 $Y2=1.485
r121 7 9 149.42 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=4.685 $Y=1.205
+ $X2=4.685 $Y2=0.74
r122 4 35 26.8826 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=4.36 $Y=1.765
+ $X2=4.36 $Y2=1.485
r123 4 6 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=4.36 $Y=1.765
+ $X2=4.36 $Y2=2.4
r124 1 35 20.2278 $w=4.17e-07 $l=3.56931e-07 $layer=POLY_cond $X=4.185 $Y=1.205
+ $X2=4.36 $Y2=1.485
r125 1 3 149.42 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=4.185 $Y=1.205
+ $X2=4.185 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HS__A41OI_4%A3 1 3 6 8 10 13 15 17 20 22 24 27 29 30 31
+ 32 33 51
c87 33 0 1.87135e-19 $X=7.92 $Y=1.665
c88 22 0 9.95466e-21 $X=7.72 $Y=1.765
c89 13 0 1.85629e-19 $X=6.965 $Y=0.74
r90 51 52 13.8658 $w=3.65e-07 $l=1.05e-07 $layer=POLY_cond $X=7.72 $Y=1.557
+ $X2=7.825 $Y2=1.557
r91 49 51 1.98082 $w=3.65e-07 $l=1.5e-08 $layer=POLY_cond $X=7.705 $Y=1.557
+ $X2=7.72 $Y2=1.557
r92 49 50 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=7.705
+ $Y=1.515 $X2=7.705 $Y2=1.515
r93 47 49 40.937 $w=3.65e-07 $l=3.1e-07 $layer=POLY_cond $X=7.395 $Y=1.557
+ $X2=7.705 $Y2=1.557
r94 46 47 23.1096 $w=3.65e-07 $l=1.75e-07 $layer=POLY_cond $X=7.22 $Y=1.557
+ $X2=7.395 $Y2=1.557
r95 45 46 33.674 $w=3.65e-07 $l=2.55e-07 $layer=POLY_cond $X=6.965 $Y=1.557
+ $X2=7.22 $Y2=1.557
r96 44 45 25.7507 $w=3.65e-07 $l=1.95e-07 $layer=POLY_cond $X=6.77 $Y=1.557
+ $X2=6.965 $Y2=1.557
r97 43 44 31.0329 $w=3.65e-07 $l=2.35e-07 $layer=POLY_cond $X=6.535 $Y=1.557
+ $X2=6.77 $Y2=1.557
r98 41 43 25.0904 $w=3.65e-07 $l=1.9e-07 $layer=POLY_cond $X=6.345 $Y=1.557
+ $X2=6.535 $Y2=1.557
r99 41 42 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=6.345
+ $Y=1.515 $X2=6.345 $Y2=1.515
r100 39 41 9.90411 $w=3.65e-07 $l=7.5e-08 $layer=POLY_cond $X=6.27 $Y=1.557
+ $X2=6.345 $Y2=1.557
r101 33 50 5.76222 $w=4.28e-07 $l=2.15e-07 $layer=LI1_cond $X=7.92 $Y=1.565
+ $X2=7.705 $Y2=1.565
r102 32 50 7.10226 $w=4.28e-07 $l=2.65e-07 $layer=LI1_cond $X=7.44 $Y=1.565
+ $X2=7.705 $Y2=1.565
r103 31 32 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=6.96 $Y=1.565
+ $X2=7.44 $Y2=1.565
r104 30 31 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=6.48 $Y=1.565
+ $X2=6.96 $Y2=1.565
r105 30 42 3.61813 $w=4.28e-07 $l=1.35e-07 $layer=LI1_cond $X=6.48 $Y=1.565
+ $X2=6.345 $Y2=1.565
r106 29 42 9.24634 $w=4.28e-07 $l=3.45e-07 $layer=LI1_cond $X=6 $Y=1.565
+ $X2=6.345 $Y2=1.565
r107 25 52 23.6381 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=7.825 $Y=1.35
+ $X2=7.825 $Y2=1.557
r108 25 27 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=7.825 $Y=1.35
+ $X2=7.825 $Y2=0.74
r109 22 51 23.6381 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=7.72 $Y=1.765
+ $X2=7.72 $Y2=1.557
r110 22 24 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=7.72 $Y=1.765
+ $X2=7.72 $Y2=2.4
r111 18 47 23.6381 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=7.395 $Y=1.35
+ $X2=7.395 $Y2=1.557
r112 18 20 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=7.395 $Y=1.35
+ $X2=7.395 $Y2=0.74
r113 15 46 23.6381 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=7.22 $Y=1.765
+ $X2=7.22 $Y2=1.557
r114 15 17 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=7.22 $Y=1.765
+ $X2=7.22 $Y2=2.4
r115 11 45 23.6381 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=6.965 $Y=1.35
+ $X2=6.965 $Y2=1.557
r116 11 13 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=6.965 $Y=1.35
+ $X2=6.965 $Y2=0.74
r117 8 44 23.6381 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=6.77 $Y=1.765
+ $X2=6.77 $Y2=1.557
r118 8 10 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=6.77 $Y=1.765
+ $X2=6.77 $Y2=2.4
r119 4 43 23.6381 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=6.535 $Y=1.35
+ $X2=6.535 $Y2=1.557
r120 4 6 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=6.535 $Y=1.35
+ $X2=6.535 $Y2=0.74
r121 1 39 23.6381 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=6.27 $Y=1.765
+ $X2=6.27 $Y2=1.557
r122 1 3 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=6.27 $Y=1.765
+ $X2=6.27 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_HS__A41OI_4%A4 1 3 6 8 10 13 17 19 21 22 24 27 29 30 31
+ 32 49
c78 32 0 9.95466e-21 $X=9.84 $Y=1.665
c79 6 0 2.04552e-19 $X=8.255 $Y=0.74
c80 1 0 1.27766e-19 $X=8.22 $Y=1.765
r81 49 50 1.95405 $w=3.7e-07 $l=1.5e-08 $layer=POLY_cond $X=9.57 $Y=1.557
+ $X2=9.585 $Y2=1.557
r82 47 49 13.027 $w=3.7e-07 $l=1e-07 $layer=POLY_cond $X=9.47 $Y=1.557 $X2=9.57
+ $Y2=1.557
r83 47 48 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=9.47
+ $Y=1.515 $X2=9.47 $Y2=1.515
r84 45 47 45.5946 $w=3.7e-07 $l=3.5e-07 $layer=POLY_cond $X=9.12 $Y=1.557
+ $X2=9.47 $Y2=1.557
r85 44 45 0.651351 $w=3.7e-07 $l=5e-09 $layer=POLY_cond $X=9.115 $Y=1.557
+ $X2=9.12 $Y2=1.557
r86 43 44 56.0162 $w=3.7e-07 $l=4.3e-07 $layer=POLY_cond $X=8.685 $Y=1.557
+ $X2=9.115 $Y2=1.557
r87 42 43 1.95405 $w=3.7e-07 $l=1.5e-08 $layer=POLY_cond $X=8.67 $Y=1.557
+ $X2=8.685 $Y2=1.557
r88 40 42 28.6595 $w=3.7e-07 $l=2.2e-07 $layer=POLY_cond $X=8.45 $Y=1.557
+ $X2=8.67 $Y2=1.557
r89 40 41 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=8.45
+ $Y=1.515 $X2=8.45 $Y2=1.515
r90 38 40 25.4027 $w=3.7e-07 $l=1.95e-07 $layer=POLY_cond $X=8.255 $Y=1.557
+ $X2=8.45 $Y2=1.557
r91 37 38 4.55946 $w=3.7e-07 $l=3.5e-08 $layer=POLY_cond $X=8.22 $Y=1.557
+ $X2=8.255 $Y2=1.557
r92 32 48 9.91637 $w=4.28e-07 $l=3.7e-07 $layer=LI1_cond $X=9.84 $Y=1.565
+ $X2=9.47 $Y2=1.565
r93 31 48 2.94811 $w=4.28e-07 $l=1.1e-07 $layer=LI1_cond $X=9.36 $Y=1.565
+ $X2=9.47 $Y2=1.565
r94 30 31 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=8.88 $Y=1.565
+ $X2=9.36 $Y2=1.565
r95 30 41 11.5244 $w=4.28e-07 $l=4.3e-07 $layer=LI1_cond $X=8.88 $Y=1.565
+ $X2=8.45 $Y2=1.565
r96 29 41 1.34005 $w=4.28e-07 $l=5e-08 $layer=LI1_cond $X=8.4 $Y=1.565 $X2=8.45
+ $Y2=1.565
r97 25 50 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=9.585 $Y=1.35
+ $X2=9.585 $Y2=1.557
r98 25 27 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=9.585 $Y=1.35
+ $X2=9.585 $Y2=0.74
r99 22 49 23.9667 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=9.57 $Y=1.765
+ $X2=9.57 $Y2=1.557
r100 22 24 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=9.57 $Y=1.765
+ $X2=9.57 $Y2=2.4
r101 19 45 23.9667 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=9.12 $Y=1.765
+ $X2=9.12 $Y2=1.557
r102 19 21 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=9.12 $Y=1.765
+ $X2=9.12 $Y2=2.4
r103 15 44 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=9.115 $Y=1.35
+ $X2=9.115 $Y2=1.557
r104 15 17 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=9.115 $Y=1.35
+ $X2=9.115 $Y2=0.74
r105 11 43 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=8.685 $Y=1.35
+ $X2=8.685 $Y2=1.557
r106 11 13 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=8.685 $Y=1.35
+ $X2=8.685 $Y2=0.74
r107 8 42 23.9667 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=8.67 $Y=1.765
+ $X2=8.67 $Y2=1.557
r108 8 10 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=8.67 $Y=1.765
+ $X2=8.67 $Y2=2.4
r109 4 38 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=8.255 $Y=1.35
+ $X2=8.255 $Y2=1.557
r110 4 6 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=8.255 $Y=1.35
+ $X2=8.255 $Y2=0.74
r111 1 37 23.9667 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=8.22 $Y=1.765
+ $X2=8.22 $Y2=1.557
r112 1 3 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=8.22 $Y=1.765
+ $X2=8.22 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_HS__A41OI_4%A_27_368# 1 2 3 4 5 6 7 8 9 10 11 36 40 41
+ 44 46 48 49 50 54 56 57 60 62 66 68 72 74 78 80 84 86 90 92 94 96 98 102 105
+ 107 109 111 113 115
c197 56 0 1.32152e-19 $X=4.135 $Y=2.12
c198 54 0 1.35778e-19 $X=3.97 $Y=2.375
r199 94 117 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.795 $Y=2.12
+ $X2=9.795 $Y2=2.035
r200 94 96 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=9.795 $Y=2.12
+ $X2=9.795 $Y2=2.815
r201 93 115 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.06 $Y=2.035
+ $X2=8.895 $Y2=2.035
r202 92 117 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.63 $Y=2.035
+ $X2=9.795 $Y2=2.035
r203 92 93 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=9.63 $Y=2.035
+ $X2=9.06 $Y2=2.035
r204 88 115 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.895 $Y=2.12
+ $X2=8.895 $Y2=2.035
r205 88 90 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=8.895 $Y=2.12
+ $X2=8.895 $Y2=2.815
r206 87 113 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.11 $Y=2.035
+ $X2=7.945 $Y2=2.035
r207 86 115 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.73 $Y=2.035
+ $X2=8.895 $Y2=2.035
r208 86 87 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=8.73 $Y=2.035
+ $X2=8.11 $Y2=2.035
r209 82 113 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.945 $Y=2.12
+ $X2=7.945 $Y2=2.035
r210 82 84 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=7.945 $Y=2.12
+ $X2=7.945 $Y2=2.425
r211 81 111 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.16 $Y=2.035
+ $X2=6.995 $Y2=2.035
r212 80 113 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.78 $Y=2.035
+ $X2=7.945 $Y2=2.035
r213 80 81 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=7.78 $Y=2.035
+ $X2=7.16 $Y2=2.035
r214 76 111 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.995 $Y=2.12
+ $X2=6.995 $Y2=2.035
r215 76 78 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=6.995 $Y=2.12
+ $X2=6.995 $Y2=2.815
r216 75 109 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.21 $Y=2.035
+ $X2=6.045 $Y2=2.035
r217 74 111 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.83 $Y=2.035
+ $X2=6.995 $Y2=2.035
r218 74 75 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=6.83 $Y=2.035
+ $X2=6.21 $Y2=2.035
r219 70 109 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.045 $Y=2.12
+ $X2=6.045 $Y2=2.035
r220 70 72 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=6.045 $Y=2.12
+ $X2=6.045 $Y2=2.815
r221 69 107 8.61065 $w=1.7e-07 $l=1.94808e-07 $layer=LI1_cond $X=5.26 $Y=2.035
+ $X2=5.095 $Y2=1.97
r222 68 109 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.88 $Y=2.035
+ $X2=6.045 $Y2=2.035
r223 68 69 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=5.88 $Y=2.035
+ $X2=5.26 $Y2=2.035
r224 64 107 0.89609 $w=3.3e-07 $l=1.5e-07 $layer=LI1_cond $X=5.095 $Y=2.12
+ $X2=5.095 $Y2=1.97
r225 64 66 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=5.095 $Y=2.12
+ $X2=5.095 $Y2=2.815
r226 63 104 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.3 $Y=2.035
+ $X2=4.135 $Y2=2.035
r227 62 107 8.61065 $w=1.7e-07 $l=1.94808e-07 $layer=LI1_cond $X=4.93 $Y=2.035
+ $X2=5.095 $Y2=1.97
r228 62 63 41.1016 $w=1.68e-07 $l=6.3e-07 $layer=LI1_cond $X=4.93 $Y=2.035
+ $X2=4.3 $Y2=2.035
r229 58 105 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.135 $Y=2.46
+ $X2=4.135 $Y2=2.375
r230 58 60 12.3975 $w=3.28e-07 $l=3.55e-07 $layer=LI1_cond $X=4.135 $Y=2.46
+ $X2=4.135 $Y2=2.815
r231 57 105 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.135 $Y=2.29
+ $X2=4.135 $Y2=2.375
r232 56 104 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.135 $Y=2.12
+ $X2=4.135 $Y2=2.035
r233 56 57 5.93683 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=4.135 $Y=2.12
+ $X2=4.135 $Y2=2.29
r234 55 102 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.345 $Y=2.375
+ $X2=3.18 $Y2=2.375
r235 54 105 3.80956 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.97 $Y=2.375
+ $X2=4.135 $Y2=2.375
r236 54 55 40.7754 $w=1.68e-07 $l=6.25e-07 $layer=LI1_cond $X=3.97 $Y=2.375
+ $X2=3.345 $Y2=2.375
r237 51 100 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.345 $Y=2.375
+ $X2=2.18 $Y2=2.375
r238 50 102 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.015 $Y=2.375
+ $X2=3.18 $Y2=2.375
r239 50 51 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.015 $Y=2.375
+ $X2=2.345 $Y2=2.375
r240 48 100 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.18 $Y=2.46
+ $X2=2.18 $Y2=2.375
r241 48 49 15.5405 $w=3.28e-07 $l=4.45e-07 $layer=LI1_cond $X=2.18 $Y=2.46
+ $X2=2.18 $Y2=2.905
r242 47 98 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.445 $Y=2.99
+ $X2=1.28 $Y2=2.99
r243 46 49 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.015 $Y=2.99
+ $X2=2.18 $Y2=2.905
r244 46 47 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=2.015 $Y=2.99
+ $X2=1.445 $Y2=2.99
r245 42 98 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.28 $Y=2.905
+ $X2=1.28 $Y2=2.99
r246 42 44 17.4613 $w=3.28e-07 $l=5e-07 $layer=LI1_cond $X=1.28 $Y=2.905
+ $X2=1.28 $Y2=2.405
r247 40 98 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.115 $Y=2.99
+ $X2=1.28 $Y2=2.99
r248 40 41 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.115 $Y=2.99
+ $X2=0.445 $Y2=2.99
r249 36 39 27.2396 $w=3.28e-07 $l=7.8e-07 $layer=LI1_cond $X=0.28 $Y=2.035
+ $X2=0.28 $Y2=2.815
r250 34 41 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.28 $Y=2.905
+ $X2=0.445 $Y2=2.99
r251 34 39 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=0.28 $Y=2.905
+ $X2=0.28 $Y2=2.815
r252 11 117 400 $w=1.7e-07 $l=2.59374e-07 $layer=licon1_PDIFF $count=1 $X=9.645
+ $Y=1.84 $X2=9.795 $Y2=2.035
r253 11 96 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=9.645
+ $Y=1.84 $X2=9.795 $Y2=2.815
r254 10 115 400 $w=1.7e-07 $l=2.59374e-07 $layer=licon1_PDIFF $count=1 $X=8.745
+ $Y=1.84 $X2=8.895 $Y2=2.035
r255 10 90 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=8.745
+ $Y=1.84 $X2=8.895 $Y2=2.815
r256 9 113 600 $w=1.7e-07 $l=2.59374e-07 $layer=licon1_PDIFF $count=1 $X=7.795
+ $Y=1.84 $X2=7.945 $Y2=2.035
r257 9 84 300 $w=1.7e-07 $l=6.55725e-07 $layer=licon1_PDIFF $count=2 $X=7.795
+ $Y=1.84 $X2=7.945 $Y2=2.425
r258 8 111 400 $w=1.7e-07 $l=2.59374e-07 $layer=licon1_PDIFF $count=1 $X=6.845
+ $Y=1.84 $X2=6.995 $Y2=2.035
r259 8 78 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=6.845
+ $Y=1.84 $X2=6.995 $Y2=2.815
r260 7 109 400 $w=1.7e-07 $l=2.59374e-07 $layer=licon1_PDIFF $count=1 $X=5.895
+ $Y=1.84 $X2=6.045 $Y2=2.035
r261 7 72 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=5.895
+ $Y=1.84 $X2=6.045 $Y2=2.815
r262 6 107 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=4.945
+ $Y=1.84 $X2=5.095 $Y2=1.985
r263 6 66 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=4.945
+ $Y=1.84 $X2=5.095 $Y2=2.815
r264 5 104 400 $w=1.7e-07 $l=2.59374e-07 $layer=licon1_PDIFF $count=1 $X=3.985
+ $Y=1.84 $X2=4.135 $Y2=2.035
r265 5 60 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=3.985
+ $Y=1.84 $X2=4.135 $Y2=2.815
r266 4 102 300 $w=1.7e-07 $l=6.05372e-07 $layer=licon1_PDIFF $count=2 $X=3.03
+ $Y=1.84 $X2=3.18 $Y2=2.375
r267 3 100 300 $w=1.7e-07 $l=6.05372e-07 $layer=licon1_PDIFF $count=2 $X=2.03
+ $Y=1.84 $X2=2.18 $Y2=2.375
r268 2 44 300 $w=1.7e-07 $l=6.57438e-07 $layer=licon1_PDIFF $count=2 $X=1.08
+ $Y=1.84 $X2=1.28 $Y2=2.405
r269 1 39 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.815
r270 1 36 400 $w=1.7e-07 $l=2.57488e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.035
.ends

.subckt PM_SKY130_FD_SC_HS__A41OI_4%Y 1 2 3 4 5 18 22 23 28 31 32 34 36 41 44 46
+ 51 55 61 63
c110 61 0 1.73187e-19 $X=3.59 $Y=1.55
c111 55 0 1.21942e-19 $X=3.515 $Y=1.58
c112 51 0 1.63532e-19 $X=3.47 $Y=0.785
c113 46 0 1.77296e-19 $X=2.105 $Y=1.97
r114 58 63 0.460977 $w=2.48e-07 $l=1e-08 $layer=LI1_cond $X=3.59 $Y=1.675
+ $X2=3.59 $Y2=1.665
r115 55 63 1.75171 $w=2.48e-07 $l=3.8e-08 $layer=LI1_cond $X=3.59 $Y=1.627
+ $X2=3.59 $Y2=1.665
r116 55 61 4.73668 $w=2.48e-07 $l=7.7e-08 $layer=LI1_cond $X=3.59 $Y=1.627
+ $X2=3.59 $Y2=1.55
r117 55 58 1.70562 $w=2.48e-07 $l=3.7e-08 $layer=LI1_cond $X=3.59 $Y=1.712
+ $X2=3.59 $Y2=1.675
r118 54 55 10.9713 $w=2.48e-07 $l=2.38e-07 $layer=LI1_cond $X=3.59 $Y=1.95
+ $X2=3.59 $Y2=1.712
r119 53 61 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=3.55 $Y=1 $X2=3.55
+ $Y2=1.55
r120 51 53 10.2083 $w=3.28e-07 $l=2.15e-07 $layer=LI1_cond $X=3.47 $Y=0.785
+ $X2=3.47 $Y2=1
r121 45 46 7.71634 $w=2.98e-07 $l=1.45e-07 $layer=LI1_cond $X=1.96 $Y=1.97
+ $X2=2.105 $Y2=1.97
r122 43 45 8.8354 $w=2.98e-07 $l=2.3e-07 $layer=LI1_cond $X=1.73 $Y=1.97
+ $X2=1.96 $Y2=1.97
r123 43 44 5.41145 $w=2.98e-07 $l=8.5e-08 $layer=LI1_cond $X=1.73 $Y=1.97
+ $X2=1.645 $Y2=1.97
r124 36 54 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=3.465 $Y=2.035
+ $X2=3.59 $Y2=1.95
r125 36 46 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=3.465 $Y=2.035
+ $X2=2.105 $Y2=2.035
r126 32 34 8.73063 $w=3.28e-07 $l=2.5e-07 $layer=LI1_cond $X=2.27 $Y=1.01
+ $X2=2.27 $Y2=0.76
r127 31 45 0.922372 $w=2.9e-07 $l=1.5e-07 $layer=LI1_cond $X=1.96 $Y=1.82
+ $X2=1.96 $Y2=1.97
r128 30 32 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=1.96 $Y=1.095
+ $X2=2.27 $Y2=1.095
r129 30 31 25.4332 $w=2.88e-07 $l=6.4e-07 $layer=LI1_cond $X=1.96 $Y=1.18
+ $X2=1.96 $Y2=1.82
r130 26 43 4.061 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=1.73 $Y=2.12 $X2=1.73
+ $Y2=1.97
r131 26 28 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=1.73 $Y=2.12
+ $X2=1.73 $Y2=2.57
r132 25 41 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.945 $Y=2.035
+ $X2=0.78 $Y2=2.035
r133 25 44 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=0.945 $Y=2.035
+ $X2=1.645 $Y2=2.035
r134 22 30 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=1.815 $Y=1.095
+ $X2=1.96 $Y2=1.095
r135 22 23 61.3262 $w=1.68e-07 $l=9.4e-07 $layer=LI1_cond $X=1.815 $Y=1.095
+ $X2=0.875 $Y2=1.095
r136 16 23 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.71 $Y=1.01
+ $X2=0.875 $Y2=1.095
r137 16 18 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=0.71 $Y=1.01
+ $X2=0.71 $Y2=0.515
r138 5 43 600 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=1.58
+ $Y=1.84 $X2=1.73 $Y2=1.985
r139 5 28 600 $w=1.7e-07 $l=8.01499e-07 $layer=licon1_PDIFF $count=1 $X=1.58
+ $Y=1.84 $X2=1.73 $Y2=2.57
r140 4 41 300 $w=1.7e-07 $l=3.17884e-07 $layer=licon1_PDIFF $count=2 $X=0.585
+ $Y=1.84 $X2=0.78 $Y2=2.075
r141 3 51 182 $w=1.7e-07 $l=4.79922e-07 $layer=licon1_NDIFF $count=1 $X=3.33
+ $Y=0.37 $X2=3.47 $Y2=0.785
r142 2 34 182 $w=1.7e-07 $l=4.83735e-07 $layer=licon1_NDIFF $count=1 $X=2.06
+ $Y=0.37 $X2=2.27 $Y2=0.76
r143 1 18 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=0.57
+ $Y=0.37 $X2=0.71 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__A41OI_4%VPWR 1 2 3 4 5 6 7 8 27 29 33 35 39 41 45 47
+ 51 53 57 61 65 68 69 70 72 80 90 91 94 97 100 103 106 109 112
r144 112 113 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=3.33
+ $X2=8.4 $Y2=3.33
r145 109 110 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r146 107 110 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=7.44 $Y2=3.33
r147 106 107 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r148 104 107 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=6.48 $Y2=3.33
r149 103 104 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r150 100 101 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r151 98 101 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.56 $Y2=3.33
r152 97 98 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r153 95 98 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.6 $Y2=3.33
r154 94 95 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r155 90 91 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.84 $Y=3.33
+ $X2=9.84 $Y2=3.33
r156 88 91 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=8.88 $Y=3.33
+ $X2=9.84 $Y2=3.33
r157 88 113 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=3.33
+ $X2=8.4 $Y2=3.33
r158 87 88 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r159 85 112 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.53 $Y=3.33
+ $X2=8.405 $Y2=3.33
r160 85 87 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=8.53 $Y=3.33
+ $X2=8.88 $Y2=3.33
r161 84 113 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=3.33
+ $X2=8.4 $Y2=3.33
r162 84 110 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=3.33
+ $X2=7.44 $Y2=3.33
r163 83 84 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r164 81 109 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.61 $Y=3.33
+ $X2=7.485 $Y2=3.33
r165 81 83 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=7.61 $Y=3.33
+ $X2=7.92 $Y2=3.33
r166 80 112 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.28 $Y=3.33
+ $X2=8.405 $Y2=3.33
r167 80 83 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=8.28 $Y=3.33
+ $X2=7.92 $Y2=3.33
r168 79 95 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r169 78 79 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r170 75 79 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=2.16 $Y2=3.33
r171 74 78 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=0.24 $Y=3.33
+ $X2=2.16 $Y2=3.33
r172 74 75 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r173 72 94 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.515 $Y=3.33
+ $X2=2.68 $Y2=3.33
r174 72 78 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=2.515 $Y=3.33
+ $X2=2.16 $Y2=3.33
r175 70 104 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=5.52 $Y2=3.33
r176 70 101 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=4.56 $Y2=3.33
r177 68 87 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=9.26 $Y=3.33
+ $X2=8.88 $Y2=3.33
r178 68 69 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.26 $Y=3.33
+ $X2=9.345 $Y2=3.33
r179 67 90 26.7487 $w=1.68e-07 $l=4.1e-07 $layer=LI1_cond $X=9.43 $Y=3.33
+ $X2=9.84 $Y2=3.33
r180 67 69 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.43 $Y=3.33
+ $X2=9.345 $Y2=3.33
r181 63 69 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.345 $Y=3.245
+ $X2=9.345 $Y2=3.33
r182 63 65 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=9.345 $Y=3.245
+ $X2=9.345 $Y2=2.455
r183 59 112 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=8.405 $Y=3.245
+ $X2=8.405 $Y2=3.33
r184 59 61 36.4172 $w=2.48e-07 $l=7.9e-07 $layer=LI1_cond $X=8.405 $Y=3.245
+ $X2=8.405 $Y2=2.455
r185 55 109 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=7.485 $Y=3.245
+ $X2=7.485 $Y2=3.33
r186 55 57 36.4172 $w=2.48e-07 $l=7.9e-07 $layer=LI1_cond $X=7.485 $Y=3.245
+ $X2=7.485 $Y2=2.455
r187 54 106 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.66 $Y=3.33
+ $X2=6.535 $Y2=3.33
r188 53 109 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.36 $Y=3.33
+ $X2=7.485 $Y2=3.33
r189 53 54 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=7.36 $Y=3.33 $X2=6.66
+ $Y2=3.33
r190 49 106 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.535 $Y=3.245
+ $X2=6.535 $Y2=3.33
r191 49 51 36.4172 $w=2.48e-07 $l=7.9e-07 $layer=LI1_cond $X=6.535 $Y=3.245
+ $X2=6.535 $Y2=2.455
r192 48 103 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.71 $Y=3.33
+ $X2=5.585 $Y2=3.33
r193 47 106 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.41 $Y=3.33
+ $X2=6.535 $Y2=3.33
r194 47 48 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=6.41 $Y=3.33 $X2=5.71
+ $Y2=3.33
r195 43 103 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.585 $Y=3.245
+ $X2=5.585 $Y2=3.33
r196 43 45 36.4172 $w=2.48e-07 $l=7.9e-07 $layer=LI1_cond $X=5.585 $Y=3.245
+ $X2=5.585 $Y2=2.455
r197 42 100 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.75 $Y=3.33
+ $X2=4.625 $Y2=3.33
r198 41 103 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.46 $Y=3.33
+ $X2=5.585 $Y2=3.33
r199 41 42 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=5.46 $Y=3.33
+ $X2=4.75 $Y2=3.33
r200 37 100 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.625 $Y=3.245
+ $X2=4.625 $Y2=3.33
r201 37 39 36.4172 $w=2.48e-07 $l=7.9e-07 $layer=LI1_cond $X=4.625 $Y=3.245
+ $X2=4.625 $Y2=2.455
r202 36 97 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.795 $Y=3.33
+ $X2=3.67 $Y2=3.33
r203 35 100 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.5 $Y=3.33
+ $X2=4.625 $Y2=3.33
r204 35 36 45.9947 $w=1.68e-07 $l=7.05e-07 $layer=LI1_cond $X=4.5 $Y=3.33
+ $X2=3.795 $Y2=3.33
r205 31 97 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.67 $Y=3.245
+ $X2=3.67 $Y2=3.33
r206 31 33 20.744 $w=2.48e-07 $l=4.5e-07 $layer=LI1_cond $X=3.67 $Y=3.245
+ $X2=3.67 $Y2=2.795
r207 30 94 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.845 $Y=3.33
+ $X2=2.68 $Y2=3.33
r208 29 97 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.545 $Y=3.33
+ $X2=3.67 $Y2=3.33
r209 29 30 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=3.545 $Y=3.33
+ $X2=2.845 $Y2=3.33
r210 25 94 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.68 $Y=3.245
+ $X2=2.68 $Y2=3.33
r211 25 27 17.8105 $w=3.28e-07 $l=5.1e-07 $layer=LI1_cond $X=2.68 $Y=3.245
+ $X2=2.68 $Y2=2.735
r212 8 65 300 $w=1.7e-07 $l=6.85912e-07 $layer=licon1_PDIFF $count=2 $X=9.195
+ $Y=1.84 $X2=9.345 $Y2=2.455
r213 7 61 300 $w=1.7e-07 $l=6.85912e-07 $layer=licon1_PDIFF $count=2 $X=8.295
+ $Y=1.84 $X2=8.445 $Y2=2.455
r214 6 57 300 $w=1.7e-07 $l=6.85912e-07 $layer=licon1_PDIFF $count=2 $X=7.295
+ $Y=1.84 $X2=7.445 $Y2=2.455
r215 5 51 300 $w=1.7e-07 $l=6.85912e-07 $layer=licon1_PDIFF $count=2 $X=6.345
+ $Y=1.84 $X2=6.495 $Y2=2.455
r216 4 45 300 $w=1.7e-07 $l=6.85912e-07 $layer=licon1_PDIFF $count=2 $X=5.395
+ $Y=1.84 $X2=5.545 $Y2=2.455
r217 3 39 300 $w=1.7e-07 $l=6.85912e-07 $layer=licon1_PDIFF $count=2 $X=4.435
+ $Y=1.84 $X2=4.585 $Y2=2.455
r218 2 33 600 $w=1.7e-07 $l=1.02727e-06 $layer=licon1_PDIFF $count=1 $X=3.48
+ $Y=1.84 $X2=3.63 $Y2=2.795
r219 1 27 600 $w=1.7e-07 $l=9.89962e-07 $layer=licon1_PDIFF $count=1 $X=2.48
+ $Y=1.84 $X2=2.68 $Y2=2.735
.ends

.subckt PM_SKY130_FD_SC_HS__A41OI_4%VGND 1 2 3 4 13 15 19 23 27 29 31 36 44 51
+ 52 58 61 64
r99 64 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.36 $Y=0 $X2=9.36
+ $Y2=0
r100 61 62 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r101 58 59 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r102 55 56 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r103 52 65 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.84 $Y=0 $X2=9.36
+ $Y2=0
r104 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.84 $Y=0 $X2=9.84
+ $Y2=0
r105 49 64 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.495 $Y=0 $X2=9.33
+ $Y2=0
r106 49 51 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=9.495 $Y=0 $X2=9.84
+ $Y2=0
r107 48 65 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=0 $X2=9.36
+ $Y2=0
r108 48 62 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=0 $X2=8.4
+ $Y2=0
r109 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=0 $X2=8.88
+ $Y2=0
r110 45 61 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.635 $Y=0 $X2=8.47
+ $Y2=0
r111 45 47 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=8.635 $Y=0 $X2=8.88
+ $Y2=0
r112 44 64 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.165 $Y=0 $X2=9.33
+ $Y2=0
r113 44 47 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=9.165 $Y=0
+ $X2=8.88 $Y2=0
r114 43 62 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=0 $X2=8.4
+ $Y2=0
r115 42 43 1.32857 $w=1.7e-07 $l=1.19e-06 $layer=mcon $count=7 $X=7.92 $Y=0
+ $X2=7.92 $Y2=0
r116 40 59 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r117 39 42 407.102 $w=1.68e-07 $l=6.24e-06 $layer=LI1_cond $X=1.68 $Y=0 $X2=7.92
+ $Y2=0
r118 39 40 1.32857 $w=1.7e-07 $l=1.19e-06 $layer=mcon $count=7 $X=1.68 $Y=0
+ $X2=1.68 $Y2=0
r119 37 58 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.375 $Y=0 $X2=1.21
+ $Y2=0
r120 37 39 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.375 $Y=0
+ $X2=1.68 $Y2=0
r121 36 61 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.305 $Y=0 $X2=8.47
+ $Y2=0
r122 36 42 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=8.305 $Y=0
+ $X2=7.92 $Y2=0
r123 35 59 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r124 35 56 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r125 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r126 32 55 4.00981 $w=1.7e-07 $l=1.83e-07 $layer=LI1_cond $X=0.365 $Y=0
+ $X2=0.182 $Y2=0
r127 32 34 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=0.365 $Y=0
+ $X2=0.72 $Y2=0
r128 31 58 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.045 $Y=0 $X2=1.21
+ $Y2=0
r129 31 34 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=1.045 $Y=0
+ $X2=0.72 $Y2=0
r130 29 43 0.802756 $w=4.9e-07 $l=2.88e-06 $layer=MET1_cond $X=5.04 $Y=0
+ $X2=7.92 $Y2=0
r131 29 40 0.936549 $w=4.9e-07 $l=3.36e-06 $layer=MET1_cond $X=5.04 $Y=0
+ $X2=1.68 $Y2=0
r132 25 64 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.33 $Y=0.085
+ $X2=9.33 $Y2=0
r133 25 27 20.6043 $w=3.28e-07 $l=5.9e-07 $layer=LI1_cond $X=9.33 $Y=0.085
+ $X2=9.33 $Y2=0.675
r134 21 61 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.47 $Y=0.085
+ $X2=8.47 $Y2=0
r135 21 23 20.6043 $w=3.28e-07 $l=5.9e-07 $layer=LI1_cond $X=8.47 $Y=0.085
+ $X2=8.47 $Y2=0.675
r136 17 58 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.21 $Y=0.085
+ $X2=1.21 $Y2=0
r137 17 19 20.6043 $w=3.28e-07 $l=5.9e-07 $layer=LI1_cond $X=1.21 $Y=0.085
+ $X2=1.21 $Y2=0.675
r138 13 55 3.13335 $w=2.5e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.24 $Y=0.085
+ $X2=0.182 $Y2=0
r139 13 15 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=0.24 $Y=0.085
+ $X2=0.24 $Y2=0.515
r140 4 27 182 $w=1.7e-07 $l=3.68409e-07 $layer=licon1_NDIFF $count=1 $X=9.19
+ $Y=0.37 $X2=9.33 $Y2=0.675
r141 3 23 182 $w=1.7e-07 $l=3.68409e-07 $layer=licon1_NDIFF $count=1 $X=8.33
+ $Y=0.37 $X2=8.47 $Y2=0.675
r142 2 19 182 $w=1.7e-07 $l=3.68409e-07 $layer=licon1_NDIFF $count=1 $X=1.07
+ $Y=0.37 $X2=1.21 $Y2=0.675
r143 1 15 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__A41OI_4%A_325_74# 1 2 3 4 5 18 20 21 24 26 34 36 38
r63 32 34 27.1535 $w=3.63e-07 $l=8.6e-07 $layer=LI1_cond $X=4.9 $Y=0.437
+ $X2=5.76 $Y2=0.437
r64 30 38 6.12952 $w=2.67e-07 $l=1.65e-07 $layer=LI1_cond $X=4.135 $Y=0.437
+ $X2=3.97 $Y2=0.437
r65 30 32 24.1539 $w=3.63e-07 $l=7.65e-07 $layer=LI1_cond $X=4.135 $Y=0.437
+ $X2=4.9 $Y2=0.437
r66 27 36 11.6921 $w=1.7e-07 $l=2.65e-07 $layer=LI1_cond $X=3.135 $Y=0.34
+ $X2=2.87 $Y2=0.34
r67 26 38 6.12952 $w=2.67e-07 $l=2.07918e-07 $layer=LI1_cond $X=3.805 $Y=0.34
+ $X2=3.97 $Y2=0.437
r68 26 27 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.805 $Y=0.34
+ $X2=3.135 $Y2=0.34
r69 22 36 2.222 $w=5.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.87 $Y=0.425 $X2=2.87
+ $Y2=0.34
r70 22 24 2.03108 $w=5.28e-07 $l=9e-08 $layer=LI1_cond $X=2.87 $Y=0.425 $X2=2.87
+ $Y2=0.515
r71 20 36 11.6921 $w=1.7e-07 $l=2.65e-07 $layer=LI1_cond $X=2.605 $Y=0.34
+ $X2=2.87 $Y2=0.34
r72 20 21 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.605 $Y=0.34
+ $X2=1.935 $Y2=0.34
r73 16 21 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.77 $Y=0.425
+ $X2=1.935 $Y2=0.34
r74 16 18 8.03218 $w=3.28e-07 $l=2.3e-07 $layer=LI1_cond $X=1.77 $Y=0.425
+ $X2=1.77 $Y2=0.655
r75 5 34 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=5.62
+ $Y=0.37 $X2=5.76 $Y2=0.515
r76 4 32 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=4.76
+ $Y=0.37 $X2=4.9 $Y2=0.515
r77 3 38 91 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=2 $X=3.76
+ $Y=0.37 $X2=3.97 $Y2=0.515
r78 2 24 45.5 $w=1.7e-07 $l=5.47723e-07 $layer=licon1_NDIFF $count=4 $X=2.56
+ $Y=0.37 $X2=3.04 $Y2=0.515
r79 1 18 182 $w=1.7e-07 $l=3.50071e-07 $layer=licon1_NDIFF $count=1 $X=1.625
+ $Y=0.37 $X2=1.77 $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_HS__A41OI_4%A_852_74# 1 2 3 4 22 23
c31 22 0 1.35727e-19 $X=7.61 $Y=0.95
r32 22 23 5.33064 $w=3.58e-07 $l=1.65e-07 $layer=LI1_cond $X=7.61 $Y=0.95
+ $X2=7.445 $Y2=0.95
r33 20 23 23.5573 $w=3.38e-07 $l=6.95e-07 $layer=LI1_cond $X=6.75 $Y=0.96
+ $X2=7.445 $Y2=0.96
r34 18 20 48.1314 $w=3.38e-07 $l=1.42e-06 $layer=LI1_cond $X=5.33 $Y=0.96
+ $X2=6.75 $Y2=0.96
r35 15 18 29.15 $w=3.38e-07 $l=8.6e-07 $layer=LI1_cond $X=4.47 $Y=0.96 $X2=5.33
+ $Y2=0.96
r36 4 22 182 $w=1.7e-07 $l=6.4622e-07 $layer=licon1_NDIFF $count=1 $X=7.47
+ $Y=0.37 $X2=7.61 $Y2=0.95
r37 3 20 182 $w=1.7e-07 $l=6.56277e-07 $layer=licon1_NDIFF $count=1 $X=6.61
+ $Y=0.37 $X2=6.75 $Y2=0.96
r38 2 18 182 $w=1.7e-07 $l=6.4622e-07 $layer=licon1_NDIFF $count=1 $X=5.19
+ $Y=0.37 $X2=5.33 $Y2=0.95
r39 1 15 182 $w=1.7e-07 $l=6.76905e-07 $layer=licon1_NDIFF $count=1 $X=4.26
+ $Y=0.37 $X2=4.47 $Y2=0.95
.ends

.subckt PM_SKY130_FD_SC_HS__A41OI_4%A_1235_74# 1 2 3 4 5 16 20 24 25 28 30 34 39
+ 42
c55 39 0 9.28144e-20 $X=6.485 $Y=0.485
c56 20 0 1.6164e-19 $X=8.04 $Y=0.6
r57 37 39 7.12439 $w=2.68e-07 $l=1.65e-07 $layer=LI1_cond $X=6.32 $Y=0.485
+ $X2=6.485 $Y2=0.485
r58 32 34 22.8184 $w=2.48e-07 $l=4.95e-07 $layer=LI1_cond $X=9.84 $Y=1.01
+ $X2=9.84 $Y2=0.515
r59 31 42 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.985 $Y=1.095
+ $X2=8.9 $Y2=1.095
r60 30 32 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=9.715 $Y=1.095
+ $X2=9.84 $Y2=1.01
r61 30 31 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=9.715 $Y=1.095
+ $X2=8.985 $Y2=1.095
r62 26 42 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.9 $Y=1.01 $X2=8.9
+ $Y2=1.095
r63 26 28 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=8.9 $Y=1.01 $X2=8.9
+ $Y2=0.515
r64 24 42 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.815 $Y=1.095
+ $X2=8.9 $Y2=1.095
r65 24 25 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=8.815 $Y=1.095
+ $X2=8.125 $Y2=1.095
r66 21 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.04 $Y=1.01
+ $X2=8.125 $Y2=1.095
r67 21 23 2.93583 $w=1.68e-07 $l=4.5e-08 $layer=LI1_cond $X=8.04 $Y=1.01
+ $X2=8.04 $Y2=0.965
r68 20 41 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.04 $Y=0.6 $X2=8.04
+ $Y2=0.475
r69 20 23 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=8.04 $Y=0.6
+ $X2=8.04 $Y2=0.965
r70 19 39 32.0379 $w=2.48e-07 $l=6.95e-07 $layer=LI1_cond $X=7.18 $Y=0.475
+ $X2=6.485 $Y2=0.475
r71 16 41 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=7.955 $Y=0.475
+ $X2=8.04 $Y2=0.475
r72 16 19 35.7257 $w=2.48e-07 $l=7.75e-07 $layer=LI1_cond $X=7.955 $Y=0.475
+ $X2=7.18 $Y2=0.475
r73 5 34 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=9.66
+ $Y=0.37 $X2=9.8 $Y2=0.515
r74 4 28 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=8.76
+ $Y=0.37 $X2=8.9 $Y2=0.515
r75 3 41 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=7.9
+ $Y=0.37 $X2=8.04 $Y2=0.515
r76 3 23 182 $w=1.7e-07 $l=6.61306e-07 $layer=licon1_NDIFF $count=1 $X=7.9
+ $Y=0.37 $X2=8.04 $Y2=0.965
r77 2 19 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=7.04
+ $Y=0.37 $X2=7.18 $Y2=0.515
r78 1 37 182 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_NDIFF $count=1 $X=6.175
+ $Y=0.37 $X2=6.32 $Y2=0.525
.ends

