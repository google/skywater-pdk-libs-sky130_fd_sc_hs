* File: sky130_fd_sc_hs__or4bb_4.pxi.spice
* Created: Tue Sep  1 20:21:53 2020
* 
x_PM_SKY130_FD_SC_HS__OR4BB_4%D_N N_D_N_M1004_g N_D_N_c_139_n N_D_N_M1013_g D_N
+ N_D_N_c_140_n PM_SKY130_FD_SC_HS__OR4BB_4%D_N
x_PM_SKY130_FD_SC_HS__OR4BB_4%A_193_277# N_A_193_277#_M1011_d
+ N_A_193_277#_M1007_d N_A_193_277#_M1020_d N_A_193_277#_c_189_n
+ N_A_193_277#_M1008_g N_A_193_277#_c_173_n N_A_193_277#_M1000_g
+ N_A_193_277#_c_174_n N_A_193_277#_M1009_g N_A_193_277#_c_190_n
+ N_A_193_277#_M1010_g N_A_193_277#_c_175_n N_A_193_277#_c_176_n
+ N_A_193_277#_c_177_n N_A_193_277#_M1014_g N_A_193_277#_c_178_n
+ N_A_193_277#_M1012_g N_A_193_277#_c_179_n N_A_193_277#_c_180_n
+ N_A_193_277#_M1023_g N_A_193_277#_c_181_n N_A_193_277#_M1018_g
+ N_A_193_277#_c_182_n N_A_193_277#_c_183_n N_A_193_277#_c_195_n
+ N_A_193_277#_c_289_p N_A_193_277#_c_213_p N_A_193_277#_c_196_n
+ N_A_193_277#_c_197_n N_A_193_277#_c_184_n N_A_193_277#_c_185_n
+ N_A_193_277#_c_186_n N_A_193_277#_c_187_n N_A_193_277#_c_188_n
+ PM_SKY130_FD_SC_HS__OR4BB_4%A_193_277#
x_PM_SKY130_FD_SC_HS__OR4BB_4%C_N N_C_N_c_354_n N_C_N_M1006_g N_C_N_M1005_g C_N
+ N_C_N_c_356_n PM_SKY130_FD_SC_HS__OR4BB_4%C_N
x_PM_SKY130_FD_SC_HS__OR4BB_4%A_27_94# N_A_27_94#_M1004_s N_A_27_94#_M1013_s
+ N_A_27_94#_c_391_n N_A_27_94#_c_401_n N_A_27_94#_M1020_g N_A_27_94#_c_392_n
+ N_A_27_94#_M1011_g N_A_27_94#_c_393_n N_A_27_94#_c_403_n N_A_27_94#_M1022_g
+ N_A_27_94#_c_394_n N_A_27_94#_c_404_n N_A_27_94#_c_413_n N_A_27_94#_c_405_n
+ N_A_27_94#_c_395_n N_A_27_94#_c_396_n N_A_27_94#_c_515_p N_A_27_94#_c_407_n
+ N_A_27_94#_c_408_n N_A_27_94#_c_460_n N_A_27_94#_c_397_n N_A_27_94#_c_409_n
+ N_A_27_94#_c_398_n N_A_27_94#_c_399_n PM_SKY130_FD_SC_HS__OR4BB_4%A_27_94#
x_PM_SKY130_FD_SC_HS__OR4BB_4%A_678_368# N_A_678_368#_M1005_d
+ N_A_678_368#_M1006_d N_A_678_368#_c_536_n N_A_678_368#_c_550_n
+ N_A_678_368#_M1001_g N_A_678_368#_c_537_n N_A_678_368#_c_552_n
+ N_A_678_368#_M1002_g N_A_678_368#_c_538_n N_A_678_368#_M1021_g
+ N_A_678_368#_c_553_n N_A_678_368#_c_540_n N_A_678_368#_c_541_n
+ N_A_678_368#_c_542_n N_A_678_368#_c_543_n N_A_678_368#_c_544_n
+ N_A_678_368#_c_545_n N_A_678_368#_c_546_n N_A_678_368#_c_547_n
+ N_A_678_368#_c_548_n PM_SKY130_FD_SC_HS__OR4BB_4%A_678_368#
x_PM_SKY130_FD_SC_HS__OR4BB_4%B N_B_c_640_n N_B_M1015_g N_B_M1007_g N_B_c_641_n
+ N_B_M1016_g B B N_B_c_639_n PM_SKY130_FD_SC_HS__OR4BB_4%B
x_PM_SKY130_FD_SC_HS__OR4BB_4%A N_A_c_692_n N_A_M1003_g N_A_c_693_n N_A_c_698_n
+ N_A_M1017_g N_A_c_694_n N_A_c_700_n N_A_M1019_g A A N_A_c_696_n
+ PM_SKY130_FD_SC_HS__OR4BB_4%A
x_PM_SKY130_FD_SC_HS__OR4BB_4%VPWR N_VPWR_M1013_d N_VPWR_M1010_s N_VPWR_M1023_s
+ N_VPWR_M1017_s N_VPWR_c_739_n N_VPWR_c_740_n N_VPWR_c_741_n N_VPWR_c_742_n
+ VPWR N_VPWR_c_743_n N_VPWR_c_744_n N_VPWR_c_745_n N_VPWR_c_746_n
+ N_VPWR_c_738_n N_VPWR_c_748_n N_VPWR_c_749_n N_VPWR_c_750_n N_VPWR_c_751_n
+ PM_SKY130_FD_SC_HS__OR4BB_4%VPWR
x_PM_SKY130_FD_SC_HS__OR4BB_4%X N_X_M1000_s N_X_M1012_s N_X_M1008_d N_X_M1014_d
+ N_X_c_827_n N_X_c_831_n N_X_c_821_n N_X_c_836_n X X X N_X_c_826_n N_X_c_847_n
+ X PM_SKY130_FD_SC_HS__OR4BB_4%X
x_PM_SKY130_FD_SC_HS__OR4BB_4%A_791_392# N_A_791_392#_M1020_s
+ N_A_791_392#_M1022_s N_A_791_392#_M1002_s N_A_791_392#_c_875_n
+ N_A_791_392#_c_876_n N_A_791_392#_c_877_n N_A_791_392#_c_878_n
+ PM_SKY130_FD_SC_HS__OR4BB_4%A_791_392#
x_PM_SKY130_FD_SC_HS__OR4BB_4%A_1060_392# N_A_1060_392#_M1001_d
+ N_A_1060_392#_M1015_d N_A_1060_392#_c_916_n N_A_1060_392#_c_911_n
+ N_A_1060_392#_c_909_n N_A_1060_392#_c_910_n
+ PM_SKY130_FD_SC_HS__OR4BB_4%A_1060_392#
x_PM_SKY130_FD_SC_HS__OR4BB_4%A_1273_392# N_A_1273_392#_M1015_s
+ N_A_1273_392#_M1016_s N_A_1273_392#_M1019_d N_A_1273_392#_c_939_n
+ N_A_1273_392#_c_940_n N_A_1273_392#_c_941_n N_A_1273_392#_c_942_n
+ N_A_1273_392#_c_954_n N_A_1273_392#_c_943_n N_A_1273_392#_c_944_n
+ N_A_1273_392#_c_945_n PM_SKY130_FD_SC_HS__OR4BB_4%A_1273_392#
x_PM_SKY130_FD_SC_HS__OR4BB_4%VGND N_VGND_M1004_d N_VGND_M1009_d N_VGND_M1018_d
+ N_VGND_M1011_s N_VGND_M1021_d N_VGND_M1003_d N_VGND_c_992_n N_VGND_c_993_n
+ N_VGND_c_994_n N_VGND_c_995_n N_VGND_c_996_n N_VGND_c_997_n VGND
+ N_VGND_c_998_n N_VGND_c_999_n N_VGND_c_1000_n N_VGND_c_1001_n N_VGND_c_1002_n
+ N_VGND_c_1003_n N_VGND_c_1004_n N_VGND_c_1005_n N_VGND_c_1006_n
+ N_VGND_c_1007_n N_VGND_c_1008_n N_VGND_c_1009_n
+ PM_SKY130_FD_SC_HS__OR4BB_4%VGND
cc_1 VNB N_D_N_M1004_g 0.0311889f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.79
cc_2 VNB N_D_N_c_139_n 0.0272782f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.765
cc_3 VNB N_D_N_c_140_n 0.00610691f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.515
cc_4 VNB N_A_193_277#_c_173_n 0.0188063f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.515
cc_5 VNB N_A_193_277#_c_174_n 0.0186392f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_6 VNB N_A_193_277#_c_175_n 0.0244654f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_7 VNB N_A_193_277#_c_176_n 0.0447675f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_A_193_277#_c_177_n 0.0134803f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A_193_277#_c_178_n 0.0224215f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_193_277#_c_179_n 0.0377119f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_193_277#_c_180_n 0.0276005f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_193_277#_c_181_n 0.0225662f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_193_277#_c_182_n 0.00710369f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_193_277#_c_183_n 0.00201567f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_193_277#_c_184_n 0.00563574f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_193_277#_c_185_n 0.0122806f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_193_277#_c_186_n 0.00284323f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_193_277#_c_187_n 0.0106936f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_193_277#_c_188_n 0.0100439f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_C_N_c_354_n 0.0365396f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.35
cc_21 VNB N_C_N_M1005_g 0.0285893f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.34
cc_22 VNB N_C_N_c_356_n 0.00501603f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.515
cc_23 VNB N_A_27_94#_c_391_n 0.010657f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_24 VNB N_A_27_94#_c_392_n 0.111068f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.515
cc_25 VNB N_A_27_94#_c_393_n 0.00918813f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_27_94#_c_394_n 0.0231612f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_27_94#_c_395_n 0.00342592f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_27_94#_c_396_n 0.00823713f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_27_94#_c_397_n 0.0137595f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_27_94#_c_398_n 0.0250566f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_27_94#_c_399_n 0.00304223f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_678_368#_c_536_n 0.00393626f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_33 VNB N_A_678_368#_c_537_n 0.00419329f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.515
cc_34 VNB N_A_678_368#_c_538_n 0.0416302f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_678_368#_M1021_g 0.0256758f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_678_368#_c_540_n 0.0148767f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_678_368#_c_541_n 0.0011454f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_678_368#_c_542_n 0.00641518f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_678_368#_c_543_n 0.00178187f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_678_368#_c_544_n 0.00112108f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_678_368#_c_545_n 0.00565779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_678_368#_c_546_n 0.00832903f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_678_368#_c_547_n 0.00159323f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_678_368#_c_548_n 0.053577f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_B_M1007_g 0.0354061f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.34
cc_46 VNB B 0.00503944f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.515
cc_47 VNB N_B_c_639_n 0.0363457f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_c_692_n 0.0228205f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.35
cc_49 VNB N_A_c_693_n 0.00621485f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.765
cc_50 VNB N_A_c_694_n 0.0093909f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.515
cc_51 VNB A 0.0298057f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.665
cc_52 VNB N_A_c_696_n 0.0917685f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_VPWR_c_738_n 0.362705f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_X_c_821_n 0.00240191f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_VGND_c_992_n 0.018935f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_VGND_c_993_n 0.0192538f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_VGND_c_994_n 0.010143f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_VGND_c_995_n 0.0469473f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_VGND_c_996_n 0.00981447f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_VGND_c_997_n 0.0395568f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_VGND_c_998_n 0.0194159f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_VGND_c_999_n 0.0259476f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_VGND_c_1000_n 0.024583f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_VGND_c_1001_n 0.0126445f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_VGND_c_1002_n 0.476723f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_VGND_c_1003_n 0.00577043f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_VGND_c_1004_n 0.014232f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_VGND_c_1005_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_VGND_c_1006_n 0.0202358f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_VGND_c_1007_n 0.0240707f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_VGND_c_1008_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_VGND_c_1009_n 0.0126977f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VPB N_D_N_c_139_n 0.0311716f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.765
cc_74 VPB N_D_N_c_140_n 0.00510901f $X=-0.19 $Y=1.66 $X2=0.59 $Y2=1.515
cc_75 VPB N_A_193_277#_c_189_n 0.0169301f $X=-0.19 $Y=1.66 $X2=0.585 $Y2=1.515
cc_76 VPB N_A_193_277#_c_190_n 0.0154322f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_77 VPB N_A_193_277#_c_176_n 0.0128195f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_78 VPB N_A_193_277#_c_177_n 0.0242072f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_79 VPB N_A_193_277#_c_180_n 0.0258773f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_80 VPB N_A_193_277#_c_183_n 0.0032578f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_81 VPB N_A_193_277#_c_195_n 0.0128867f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_82 VPB N_A_193_277#_c_196_n 0.0275319f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_83 VPB N_A_193_277#_c_197_n 0.00227691f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_84 VPB N_A_193_277#_c_184_n 0.00225952f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_85 VPB N_C_N_c_354_n 0.0351089f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.35
cc_86 VPB N_C_N_c_356_n 0.00389748f $X=-0.19 $Y=1.66 $X2=0.59 $Y2=1.515
cc_87 VPB N_A_27_94#_c_391_n 0.0078368f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_88 VPB N_A_27_94#_c_401_n 0.0247617f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_89 VPB N_A_27_94#_c_393_n 0.00703503f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_90 VPB N_A_27_94#_c_403_n 0.0196279f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_91 VPB N_A_27_94#_c_404_n 0.0101859f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_92 VPB N_A_27_94#_c_405_n 0.022783f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_93 VPB N_A_27_94#_c_395_n 7.52822e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_94 VPB N_A_27_94#_c_407_n 0.00718545f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_95 VPB N_A_27_94#_c_408_n 0.00129137f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_96 VPB N_A_27_94#_c_409_n 0.00710642f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_97 VPB N_A_27_94#_c_398_n 0.0127995f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_98 VPB N_A_678_368#_c_536_n 0.00729098f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_99 VPB N_A_678_368#_c_550_n 0.0199305f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_100 VPB N_A_678_368#_c_537_n 0.00818147f $X=-0.19 $Y=1.66 $X2=0.63 $Y2=1.515
cc_101 VPB N_A_678_368#_c_552_n 0.0248602f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_102 VPB N_A_678_368#_c_553_n 0.0103092f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_103 VPB N_A_678_368#_c_541_n 0.00718291f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_104 VPB N_B_c_640_n 0.0178631f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.35
cc_105 VPB N_B_c_641_n 0.0148373f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_106 VPB B 0.00455295f $X=-0.19 $Y=1.66 $X2=0.59 $Y2=1.515
cc_107 VPB N_B_c_639_n 0.0363742f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_108 VPB N_A_c_693_n 0.00762212f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.765
cc_109 VPB N_A_c_698_n 0.0214597f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.34
cc_110 VPB N_A_c_694_n 0.0115448f $X=-0.19 $Y=1.66 $X2=0.585 $Y2=1.515
cc_111 VPB N_A_c_700_n 0.0285871f $X=-0.19 $Y=1.66 $X2=0.59 $Y2=1.515
cc_112 VPB N_VPWR_c_739_n 0.0105338f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_113 VPB N_VPWR_c_740_n 0.00366295f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_114 VPB N_VPWR_c_741_n 0.0110932f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_115 VPB N_VPWR_c_742_n 0.00610411f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_116 VPB N_VPWR_c_743_n 0.0177589f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_117 VPB N_VPWR_c_744_n 0.0266691f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_118 VPB N_VPWR_c_745_n 0.114116f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_119 VPB N_VPWR_c_746_n 0.0177898f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_120 VPB N_VPWR_c_738_n 0.12312f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_121 VPB N_VPWR_c_748_n 0.0270295f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_122 VPB N_VPWR_c_749_n 0.00778858f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_123 VPB N_VPWR_c_750_n 0.00614151f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_124 VPB N_VPWR_c_751_n 0.00613757f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_125 VPB N_A_791_392#_c_875_n 0.00677025f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_126 VPB N_A_791_392#_c_876_n 0.00428226f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_127 VPB N_A_791_392#_c_877_n 0.0114725f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_128 VPB N_A_791_392#_c_878_n 0.00217178f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_129 VPB N_A_1060_392#_c_909_n 0.00256834f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_130 VPB N_A_1060_392#_c_910_n 0.0136866f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_131 VPB N_A_1273_392#_c_939_n 0.00430123f $X=-0.19 $Y=1.66 $X2=0.59 $Y2=1.515
cc_132 VPB N_A_1273_392#_c_940_n 0.00431993f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_133 VPB N_A_1273_392#_c_941_n 0.0042859f $X=-0.19 $Y=1.66 $X2=0.63 $Y2=1.665
cc_134 VPB N_A_1273_392#_c_942_n 0.0103852f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_135 VPB N_A_1273_392#_c_943_n 0.00391181f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_136 VPB N_A_1273_392#_c_944_n 0.0154052f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_137 VPB N_A_1273_392#_c_945_n 0.0305744f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_138 N_D_N_c_139_n N_A_193_277#_c_189_n 0.0294858f $X=0.505 $Y=1.765 $X2=0
+ $Y2=0
cc_139 N_D_N_M1004_g N_A_193_277#_c_173_n 0.0217683f $X=0.495 $Y=0.79 $X2=0
+ $Y2=0
cc_140 N_D_N_c_139_n N_A_193_277#_c_176_n 0.0230184f $X=0.505 $Y=1.765 $X2=0
+ $Y2=0
cc_141 N_D_N_c_140_n N_A_193_277#_c_176_n 0.0033148f $X=0.59 $Y=1.515 $X2=0
+ $Y2=0
cc_142 N_D_N_M1004_g N_A_27_94#_c_394_n 0.00583778f $X=0.495 $Y=0.79 $X2=0 $Y2=0
cc_143 N_D_N_c_139_n N_A_27_94#_c_404_n 0.00664588f $X=0.505 $Y=1.765 $X2=0
+ $Y2=0
cc_144 N_D_N_c_139_n N_A_27_94#_c_413_n 0.0111908f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_145 N_D_N_c_140_n N_A_27_94#_c_413_n 0.0107011f $X=0.59 $Y=1.515 $X2=0 $Y2=0
cc_146 N_D_N_c_139_n N_A_27_94#_c_405_n 0.00780197f $X=0.505 $Y=1.765 $X2=0
+ $Y2=0
cc_147 N_D_N_M1004_g N_A_27_94#_c_397_n 0.00284854f $X=0.495 $Y=0.79 $X2=0 $Y2=0
cc_148 N_D_N_c_139_n N_A_27_94#_c_397_n 2.14231e-19 $X=0.505 $Y=1.765 $X2=0
+ $Y2=0
cc_149 N_D_N_c_140_n N_A_27_94#_c_397_n 0.00119546f $X=0.59 $Y=1.515 $X2=0 $Y2=0
cc_150 N_D_N_c_139_n N_A_27_94#_c_409_n 0.00362985f $X=0.505 $Y=1.765 $X2=0
+ $Y2=0
cc_151 N_D_N_c_140_n N_A_27_94#_c_409_n 0.00127779f $X=0.59 $Y=1.515 $X2=0 $Y2=0
cc_152 N_D_N_M1004_g N_A_27_94#_c_398_n 0.00583479f $X=0.495 $Y=0.79 $X2=0 $Y2=0
cc_153 N_D_N_c_139_n N_A_27_94#_c_398_n 0.013423f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_154 N_D_N_c_140_n N_A_27_94#_c_398_n 0.0329253f $X=0.59 $Y=1.515 $X2=0 $Y2=0
cc_155 N_D_N_c_139_n N_VPWR_c_739_n 0.00432031f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_156 N_D_N_c_139_n N_VPWR_c_738_n 0.00508379f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_157 N_D_N_c_139_n N_VPWR_c_748_n 0.00481134f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_158 N_D_N_M1004_g N_X_c_821_n 4.0795e-19 $X=0.495 $Y=0.79 $X2=0 $Y2=0
cc_159 N_D_N_M1004_g X 8.14457e-19 $X=0.495 $Y=0.79 $X2=0 $Y2=0
cc_160 N_D_N_c_139_n X 0.00151491f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_161 N_D_N_c_140_n X 0.0261069f $X=0.59 $Y=1.515 $X2=0 $Y2=0
cc_162 N_D_N_c_139_n N_X_c_826_n 5.4667e-19 $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_163 N_D_N_M1004_g N_VGND_c_992_n 0.0074594f $X=0.495 $Y=0.79 $X2=0 $Y2=0
cc_164 N_D_N_c_139_n N_VGND_c_992_n 0.00106565f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_165 N_D_N_c_140_n N_VGND_c_992_n 0.0158407f $X=0.59 $Y=1.515 $X2=0 $Y2=0
cc_166 N_D_N_M1004_g N_VGND_c_998_n 0.00485498f $X=0.495 $Y=0.79 $X2=0 $Y2=0
cc_167 N_D_N_M1004_g N_VGND_c_1002_n 0.00514438f $X=0.495 $Y=0.79 $X2=0 $Y2=0
cc_168 N_A_193_277#_c_180_n N_C_N_c_354_n 0.0442062f $X=2.78 $Y=1.765 $X2=-0.19
+ $Y2=-0.245
cc_169 N_A_193_277#_c_182_n N_C_N_c_354_n 0.00182565f $X=3.035 $Y=1.4 $X2=-0.19
+ $Y2=-0.245
cc_170 N_A_193_277#_c_183_n N_C_N_c_354_n 0.00638266f $X=3.12 $Y=2.29 $X2=-0.19
+ $Y2=-0.245
cc_171 N_A_193_277#_c_195_n N_C_N_c_354_n 0.0206868f $X=4.385 $Y=2.375 $X2=-0.19
+ $Y2=-0.245
cc_172 N_A_193_277#_c_181_n N_C_N_M1005_g 0.0274612f $X=2.895 $Y=1.235 $X2=0
+ $Y2=0
cc_173 N_A_193_277#_c_182_n N_C_N_M1005_g 0.00269182f $X=3.035 $Y=1.4 $X2=0
+ $Y2=0
cc_174 N_A_193_277#_c_182_n N_C_N_c_356_n 0.0160535f $X=3.035 $Y=1.4 $X2=0 $Y2=0
cc_175 N_A_193_277#_c_183_n N_C_N_c_356_n 0.0180008f $X=3.12 $Y=2.29 $X2=0 $Y2=0
cc_176 N_A_193_277#_c_197_n N_A_27_94#_c_391_n 0.00137329f $X=4.715 $Y=1.845
+ $X2=0 $Y2=0
cc_177 N_A_193_277#_c_195_n N_A_27_94#_c_401_n 0.0151987f $X=4.385 $Y=2.375
+ $X2=0 $Y2=0
cc_178 N_A_193_277#_c_213_p N_A_27_94#_c_401_n 0.0107909f $X=4.55 $Y=2.2 $X2=0
+ $Y2=0
cc_179 N_A_193_277#_c_197_n N_A_27_94#_c_401_n 0.0040125f $X=4.715 $Y=1.845
+ $X2=0 $Y2=0
cc_180 N_A_193_277#_c_197_n N_A_27_94#_c_392_n 5.27313e-19 $X=4.715 $Y=1.845
+ $X2=0 $Y2=0
cc_181 N_A_193_277#_c_187_n N_A_27_94#_c_392_n 0.0155743f $X=5.975 $Y=0.805
+ $X2=0 $Y2=0
cc_182 N_A_193_277#_c_196_n N_A_27_94#_c_393_n 0.00287682f $X=5.975 $Y=1.845
+ $X2=0 $Y2=0
cc_183 N_A_193_277#_c_197_n N_A_27_94#_c_393_n 9.24928e-19 $X=4.715 $Y=1.845
+ $X2=0 $Y2=0
cc_184 N_A_193_277#_c_195_n N_A_27_94#_c_403_n 0.00416368f $X=4.385 $Y=2.375
+ $X2=0 $Y2=0
cc_185 N_A_193_277#_c_213_p N_A_27_94#_c_403_n 0.00740763f $X=4.55 $Y=2.2 $X2=0
+ $Y2=0
cc_186 N_A_193_277#_c_196_n N_A_27_94#_c_403_n 0.0095072f $X=5.975 $Y=1.845
+ $X2=0 $Y2=0
cc_187 N_A_193_277#_c_197_n N_A_27_94#_c_403_n 0.00226144f $X=4.715 $Y=1.845
+ $X2=0 $Y2=0
cc_188 N_A_193_277#_c_189_n N_A_27_94#_c_413_n 0.0154267f $X=1.055 $Y=1.765
+ $X2=0 $Y2=0
cc_189 N_A_193_277#_c_190_n N_A_27_94#_c_413_n 0.0122666f $X=1.505 $Y=1.765
+ $X2=0 $Y2=0
cc_190 N_A_193_277#_c_177_n N_A_27_94#_c_413_n 0.0134306f $X=2.05 $Y=1.765 $X2=0
+ $Y2=0
cc_191 N_A_193_277#_c_180_n N_A_27_94#_c_413_n 0.0102436f $X=2.78 $Y=1.765 $X2=0
+ $Y2=0
cc_192 N_A_193_277#_c_189_n N_A_27_94#_c_405_n 5.08122e-19 $X=1.055 $Y=1.765
+ $X2=0 $Y2=0
cc_193 N_A_193_277#_c_174_n N_A_27_94#_c_395_n 0.00126052f $X=1.5 $Y=1.235 $X2=0
+ $Y2=0
cc_194 N_A_193_277#_c_175_n N_A_27_94#_c_395_n 0.0204722f $X=1.96 $Y=1.4 $X2=0
+ $Y2=0
cc_195 N_A_193_277#_c_176_n N_A_27_94#_c_395_n 0.00127741f $X=1.595 $Y=1.4 $X2=0
+ $Y2=0
cc_196 N_A_193_277#_c_177_n N_A_27_94#_c_395_n 0.00313425f $X=2.05 $Y=1.765
+ $X2=0 $Y2=0
cc_197 N_A_193_277#_c_178_n N_A_27_94#_c_395_n 0.00299548f $X=2.09 $Y=1.235
+ $X2=0 $Y2=0
cc_198 N_A_193_277#_c_182_n N_A_27_94#_c_395_n 0.0211767f $X=3.035 $Y=1.4 $X2=0
+ $Y2=0
cc_199 N_A_193_277#_c_175_n N_A_27_94#_c_396_n 0.00396956f $X=1.96 $Y=1.4 $X2=0
+ $Y2=0
cc_200 N_A_193_277#_c_178_n N_A_27_94#_c_396_n 0.0124511f $X=2.09 $Y=1.235 $X2=0
+ $Y2=0
cc_201 N_A_193_277#_c_179_n N_A_27_94#_c_396_n 0.0114432f $X=2.69 $Y=1.4 $X2=0
+ $Y2=0
cc_202 N_A_193_277#_c_181_n N_A_27_94#_c_396_n 0.0161776f $X=2.895 $Y=1.235
+ $X2=0 $Y2=0
cc_203 N_A_193_277#_c_182_n N_A_27_94#_c_396_n 0.0837177f $X=3.035 $Y=1.4 $X2=0
+ $Y2=0
cc_204 N_A_193_277#_c_175_n N_A_27_94#_c_407_n 0.00221754f $X=1.96 $Y=1.4 $X2=0
+ $Y2=0
cc_205 N_A_193_277#_c_177_n N_A_27_94#_c_407_n 0.0129876f $X=2.05 $Y=1.765 $X2=0
+ $Y2=0
cc_206 N_A_193_277#_c_179_n N_A_27_94#_c_407_n 0.0086439f $X=2.69 $Y=1.4 $X2=0
+ $Y2=0
cc_207 N_A_193_277#_c_180_n N_A_27_94#_c_407_n 0.00956705f $X=2.78 $Y=1.765
+ $X2=0 $Y2=0
cc_208 N_A_193_277#_c_182_n N_A_27_94#_c_407_n 0.0671678f $X=3.035 $Y=1.4 $X2=0
+ $Y2=0
cc_209 N_A_193_277#_c_183_n N_A_27_94#_c_407_n 0.0121409f $X=3.12 $Y=2.29 $X2=0
+ $Y2=0
cc_210 N_A_193_277#_c_190_n N_A_27_94#_c_408_n 9.6103e-19 $X=1.505 $Y=1.765
+ $X2=0 $Y2=0
cc_211 N_A_193_277#_c_176_n N_A_27_94#_c_408_n 5.4975e-19 $X=1.595 $Y=1.4 $X2=0
+ $Y2=0
cc_212 N_A_193_277#_c_180_n N_A_27_94#_c_460_n 0.0141965f $X=2.78 $Y=1.765 $X2=0
+ $Y2=0
cc_213 N_A_193_277#_c_189_n N_A_27_94#_c_409_n 0.00159154f $X=1.055 $Y=1.765
+ $X2=0 $Y2=0
cc_214 N_A_193_277#_c_195_n N_A_678_368#_M1006_d 0.0124752f $X=4.385 $Y=2.375
+ $X2=0 $Y2=0
cc_215 N_A_193_277#_c_196_n N_A_678_368#_c_536_n 0.00383754f $X=5.975 $Y=1.845
+ $X2=0 $Y2=0
cc_216 N_A_193_277#_c_195_n N_A_678_368#_c_550_n 5.09572e-19 $X=4.385 $Y=2.375
+ $X2=0 $Y2=0
cc_217 N_A_193_277#_c_213_p N_A_678_368#_c_550_n 0.00137514f $X=4.55 $Y=2.2
+ $X2=0 $Y2=0
cc_218 N_A_193_277#_c_196_n N_A_678_368#_c_550_n 0.0125799f $X=5.975 $Y=1.845
+ $X2=0 $Y2=0
cc_219 N_A_193_277#_c_196_n N_A_678_368#_c_537_n 0.00426441f $X=5.975 $Y=1.845
+ $X2=0 $Y2=0
cc_220 N_A_193_277#_c_196_n N_A_678_368#_c_552_n 0.00919154f $X=5.975 $Y=1.845
+ $X2=0 $Y2=0
cc_221 N_A_193_277#_c_196_n N_A_678_368#_c_538_n 0.00304271f $X=5.975 $Y=1.845
+ $X2=0 $Y2=0
cc_222 N_A_193_277#_c_184_n N_A_678_368#_c_538_n 0.0141645f $X=6.06 $Y=1.76
+ $X2=0 $Y2=0
cc_223 N_A_193_277#_c_188_n N_A_678_368#_c_538_n 0.0145968f $X=6.28 $Y=0.805
+ $X2=0 $Y2=0
cc_224 N_A_193_277#_c_185_n N_A_678_368#_M1021_g 0.0139922f $X=7.025 $Y=1.175
+ $X2=0 $Y2=0
cc_225 N_A_193_277#_c_186_n N_A_678_368#_M1021_g 8.77017e-19 $X=7.19 $Y=0.515
+ $X2=0 $Y2=0
cc_226 N_A_193_277#_c_188_n N_A_678_368#_M1021_g 0.0155215f $X=6.28 $Y=0.805
+ $X2=0 $Y2=0
cc_227 N_A_193_277#_c_195_n N_A_678_368#_c_553_n 0.047293f $X=4.385 $Y=2.375
+ $X2=0 $Y2=0
cc_228 N_A_193_277#_c_213_p N_A_678_368#_c_553_n 0.00845113f $X=4.55 $Y=2.2
+ $X2=0 $Y2=0
cc_229 N_A_193_277#_c_213_p N_A_678_368#_c_541_n 8.70168e-19 $X=4.55 $Y=2.2
+ $X2=0 $Y2=0
cc_230 N_A_193_277#_c_197_n N_A_678_368#_c_541_n 0.00819458f $X=4.715 $Y=1.845
+ $X2=0 $Y2=0
cc_231 N_A_193_277#_c_197_n N_A_678_368#_c_542_n 0.00479296f $X=4.715 $Y=1.845
+ $X2=0 $Y2=0
cc_232 N_A_193_277#_c_196_n N_A_678_368#_c_545_n 0.0811325f $X=5.975 $Y=1.845
+ $X2=0 $Y2=0
cc_233 N_A_193_277#_c_197_n N_A_678_368#_c_545_n 0.00856509f $X=4.715 $Y=1.845
+ $X2=0 $Y2=0
cc_234 N_A_193_277#_c_184_n N_A_678_368#_c_545_n 0.0256549f $X=6.06 $Y=1.76
+ $X2=0 $Y2=0
cc_235 N_A_193_277#_c_187_n N_A_678_368#_c_545_n 0.0823028f $X=5.975 $Y=0.805
+ $X2=0 $Y2=0
cc_236 N_A_193_277#_c_197_n N_A_678_368#_c_547_n 0.0159627f $X=4.715 $Y=1.845
+ $X2=0 $Y2=0
cc_237 N_A_193_277#_c_196_n N_A_678_368#_c_548_n 0.00313888f $X=5.975 $Y=1.845
+ $X2=0 $Y2=0
cc_238 N_A_193_277#_c_184_n N_A_678_368#_c_548_n 0.0107278f $X=6.06 $Y=1.76
+ $X2=0 $Y2=0
cc_239 N_A_193_277#_c_187_n N_A_678_368#_c_548_n 0.0222475f $X=5.975 $Y=0.805
+ $X2=0 $Y2=0
cc_240 N_A_193_277#_c_196_n N_B_c_640_n 0.00127717f $X=5.975 $Y=1.845 $X2=-0.19
+ $Y2=-0.245
cc_241 N_A_193_277#_c_185_n N_B_M1007_g 0.0150592f $X=7.025 $Y=1.175 $X2=0 $Y2=0
cc_242 N_A_193_277#_c_186_n N_B_M1007_g 0.0119556f $X=7.19 $Y=0.515 $X2=0 $Y2=0
cc_243 N_A_193_277#_c_188_n N_B_M1007_g 8.32625e-19 $X=6.28 $Y=0.805 $X2=0 $Y2=0
cc_244 N_A_193_277#_c_196_n B 0.00148823f $X=5.975 $Y=1.845 $X2=0 $Y2=0
cc_245 N_A_193_277#_c_184_n B 0.0218154f $X=6.06 $Y=1.76 $X2=0 $Y2=0
cc_246 N_A_193_277#_c_185_n B 0.0499003f $X=7.025 $Y=1.175 $X2=0 $Y2=0
cc_247 N_A_193_277#_c_196_n N_B_c_639_n 0.00322327f $X=5.975 $Y=1.845 $X2=0
+ $Y2=0
cc_248 N_A_193_277#_c_184_n N_B_c_639_n 0.00115822f $X=6.06 $Y=1.76 $X2=0 $Y2=0
cc_249 N_A_193_277#_c_185_n N_B_c_639_n 0.0161532f $X=7.025 $Y=1.175 $X2=0 $Y2=0
cc_250 N_A_193_277#_c_185_n N_A_c_692_n 0.00345375f $X=7.025 $Y=1.175 $X2=-0.19
+ $Y2=-0.245
cc_251 N_A_193_277#_c_186_n N_A_c_692_n 0.00866944f $X=7.19 $Y=0.515 $X2=-0.19
+ $Y2=-0.245
cc_252 N_A_193_277#_c_185_n A 0.00700079f $X=7.025 $Y=1.175 $X2=0 $Y2=0
cc_253 N_A_193_277#_c_183_n N_VPWR_M1023_s 0.006159f $X=3.12 $Y=2.29 $X2=0 $Y2=0
cc_254 N_A_193_277#_c_289_p N_VPWR_M1023_s 0.00417055f $X=3.205 $Y=2.375 $X2=0
+ $Y2=0
cc_255 N_A_193_277#_c_189_n N_VPWR_c_739_n 0.00935875f $X=1.055 $Y=1.765 $X2=0
+ $Y2=0
cc_256 N_A_193_277#_c_190_n N_VPWR_c_739_n 0.00106439f $X=1.505 $Y=1.765 $X2=0
+ $Y2=0
cc_257 N_A_193_277#_c_189_n N_VPWR_c_740_n 0.00106313f $X=1.055 $Y=1.765 $X2=0
+ $Y2=0
cc_258 N_A_193_277#_c_190_n N_VPWR_c_740_n 0.00878039f $X=1.505 $Y=1.765 $X2=0
+ $Y2=0
cc_259 N_A_193_277#_c_177_n N_VPWR_c_740_n 0.0217711f $X=2.05 $Y=1.765 $X2=0
+ $Y2=0
cc_260 N_A_193_277#_c_180_n N_VPWR_c_741_n 0.0182443f $X=2.78 $Y=1.765 $X2=0
+ $Y2=0
cc_261 N_A_193_277#_c_289_p N_VPWR_c_741_n 0.00853854f $X=3.205 $Y=2.375 $X2=0
+ $Y2=0
cc_262 N_A_193_277#_c_189_n N_VPWR_c_743_n 0.00413917f $X=1.055 $Y=1.765 $X2=0
+ $Y2=0
cc_263 N_A_193_277#_c_190_n N_VPWR_c_743_n 0.00413917f $X=1.505 $Y=1.765 $X2=0
+ $Y2=0
cc_264 N_A_193_277#_c_177_n N_VPWR_c_744_n 0.00413917f $X=2.05 $Y=1.765 $X2=0
+ $Y2=0
cc_265 N_A_193_277#_c_180_n N_VPWR_c_744_n 0.00413917f $X=2.78 $Y=1.765 $X2=0
+ $Y2=0
cc_266 N_A_193_277#_c_189_n N_VPWR_c_738_n 0.00398641f $X=1.055 $Y=1.765 $X2=0
+ $Y2=0
cc_267 N_A_193_277#_c_190_n N_VPWR_c_738_n 0.00398641f $X=1.505 $Y=1.765 $X2=0
+ $Y2=0
cc_268 N_A_193_277#_c_177_n N_VPWR_c_738_n 0.00400736f $X=2.05 $Y=1.765 $X2=0
+ $Y2=0
cc_269 N_A_193_277#_c_180_n N_VPWR_c_738_n 0.00400509f $X=2.78 $Y=1.765 $X2=0
+ $Y2=0
cc_270 N_A_193_277#_c_190_n N_X_c_827_n 0.0121284f $X=1.505 $Y=1.765 $X2=0 $Y2=0
cc_271 N_A_193_277#_c_175_n N_X_c_827_n 4.83617e-19 $X=1.96 $Y=1.4 $X2=0 $Y2=0
cc_272 N_A_193_277#_c_177_n N_X_c_827_n 0.00905247f $X=2.05 $Y=1.765 $X2=0 $Y2=0
cc_273 N_A_193_277#_c_180_n N_X_c_827_n 7.96173e-19 $X=2.78 $Y=1.765 $X2=0 $Y2=0
cc_274 N_A_193_277#_c_174_n N_X_c_831_n 7.13739e-19 $X=1.5 $Y=1.235 $X2=0 $Y2=0
cc_275 N_A_193_277#_c_178_n N_X_c_831_n 0.00456788f $X=2.09 $Y=1.235 $X2=0 $Y2=0
cc_276 N_A_193_277#_c_173_n N_X_c_821_n 0.00539925f $X=1.07 $Y=1.235 $X2=0 $Y2=0
cc_277 N_A_193_277#_c_174_n N_X_c_821_n 0.00599814f $X=1.5 $Y=1.235 $X2=0 $Y2=0
cc_278 N_A_193_277#_c_178_n N_X_c_821_n 0.00163425f $X=2.09 $Y=1.235 $X2=0 $Y2=0
cc_279 N_A_193_277#_c_174_n N_X_c_836_n 0.0137427f $X=1.5 $Y=1.235 $X2=0 $Y2=0
cc_280 N_A_193_277#_c_175_n N_X_c_836_n 6.21176e-19 $X=1.96 $Y=1.4 $X2=0 $Y2=0
cc_281 N_A_193_277#_c_178_n N_X_c_836_n 0.00890041f $X=2.09 $Y=1.235 $X2=0 $Y2=0
cc_282 N_A_193_277#_c_189_n X 0.0069092f $X=1.055 $Y=1.765 $X2=0 $Y2=0
cc_283 N_A_193_277#_c_173_n X 0.00366835f $X=1.07 $Y=1.235 $X2=0 $Y2=0
cc_284 N_A_193_277#_c_174_n X 0.0012083f $X=1.5 $Y=1.235 $X2=0 $Y2=0
cc_285 N_A_193_277#_c_190_n X 0.00540334f $X=1.505 $Y=1.765 $X2=0 $Y2=0
cc_286 N_A_193_277#_c_176_n X 0.0352056f $X=1.595 $Y=1.4 $X2=0 $Y2=0
cc_287 N_A_193_277#_c_177_n X 9.2319e-19 $X=2.05 $Y=1.765 $X2=0 $Y2=0
cc_288 N_A_193_277#_c_189_n N_X_c_826_n 0.00430681f $X=1.055 $Y=1.765 $X2=0
+ $Y2=0
cc_289 N_A_193_277#_c_190_n N_X_c_826_n 6.43337e-19 $X=1.505 $Y=1.765 $X2=0
+ $Y2=0
cc_290 N_A_193_277#_c_173_n N_X_c_847_n 0.00627859f $X=1.07 $Y=1.235 $X2=0 $Y2=0
cc_291 N_A_193_277#_c_174_n N_X_c_847_n 0.00719601f $X=1.5 $Y=1.235 $X2=0 $Y2=0
cc_292 N_A_193_277#_c_195_n N_A_791_392#_M1020_s 0.00993401f $X=4.385 $Y=2.375
+ $X2=-0.19 $Y2=-0.245
cc_293 N_A_193_277#_M1020_d N_A_791_392#_c_877_n 0.00202164f $X=4.4 $Y=1.96
+ $X2=0 $Y2=0
cc_294 N_A_193_277#_c_195_n N_A_791_392#_c_877_n 0.0478336f $X=4.385 $Y=2.375
+ $X2=0 $Y2=0
cc_295 N_A_193_277#_c_196_n N_A_1060_392#_c_911_n 0.0234894f $X=5.975 $Y=1.845
+ $X2=0 $Y2=0
cc_296 N_A_193_277#_c_196_n N_A_1060_392#_c_910_n 0.0340408f $X=5.975 $Y=1.845
+ $X2=0 $Y2=0
cc_297 N_A_193_277#_c_185_n N_VGND_M1021_d 0.0059537f $X=7.025 $Y=1.175 $X2=0
+ $Y2=0
cc_298 N_A_193_277#_c_173_n N_VGND_c_992_n 0.0115201f $X=1.07 $Y=1.235 $X2=0
+ $Y2=0
cc_299 N_A_193_277#_c_173_n N_VGND_c_993_n 0.00434272f $X=1.07 $Y=1.235 $X2=0
+ $Y2=0
cc_300 N_A_193_277#_c_174_n N_VGND_c_993_n 0.00316493f $X=1.5 $Y=1.235 $X2=0
+ $Y2=0
cc_301 N_A_193_277#_c_181_n N_VGND_c_994_n 0.0144484f $X=2.895 $Y=1.235 $X2=0
+ $Y2=0
cc_302 N_A_193_277#_c_187_n N_VGND_c_995_n 0.0662709f $X=5.975 $Y=0.805 $X2=0
+ $Y2=0
cc_303 N_A_193_277#_c_185_n N_VGND_c_996_n 0.0257907f $X=7.025 $Y=1.175 $X2=0
+ $Y2=0
cc_304 N_A_193_277#_c_186_n N_VGND_c_996_n 0.0334599f $X=7.19 $Y=0.515 $X2=0
+ $Y2=0
cc_305 N_A_193_277#_c_188_n N_VGND_c_996_n 0.0247207f $X=6.28 $Y=0.805 $X2=0
+ $Y2=0
cc_306 N_A_193_277#_c_186_n N_VGND_c_997_n 0.0350086f $X=7.19 $Y=0.515 $X2=0
+ $Y2=0
cc_307 N_A_193_277#_c_178_n N_VGND_c_999_n 0.0031692f $X=2.09 $Y=1.235 $X2=0
+ $Y2=0
cc_308 N_A_193_277#_c_181_n N_VGND_c_999_n 0.00383152f $X=2.895 $Y=1.235 $X2=0
+ $Y2=0
cc_309 N_A_193_277#_c_186_n N_VGND_c_1000_n 0.0145639f $X=7.19 $Y=0.515 $X2=0
+ $Y2=0
cc_310 N_A_193_277#_c_173_n N_VGND_c_1002_n 0.00825843f $X=1.07 $Y=1.235 $X2=0
+ $Y2=0
cc_311 N_A_193_277#_c_174_n N_VGND_c_1002_n 0.00393209f $X=1.5 $Y=1.235 $X2=0
+ $Y2=0
cc_312 N_A_193_277#_c_178_n N_VGND_c_1002_n 0.00398424f $X=2.09 $Y=1.235 $X2=0
+ $Y2=0
cc_313 N_A_193_277#_c_181_n N_VGND_c_1002_n 0.00760226f $X=2.895 $Y=1.235 $X2=0
+ $Y2=0
cc_314 N_A_193_277#_c_186_n N_VGND_c_1002_n 0.0119984f $X=7.19 $Y=0.515 $X2=0
+ $Y2=0
cc_315 N_A_193_277#_c_187_n N_VGND_c_1002_n 0.0549344f $X=5.975 $Y=0.805 $X2=0
+ $Y2=0
cc_316 N_A_193_277#_c_174_n N_VGND_c_1004_n 0.00360677f $X=1.5 $Y=1.235 $X2=0
+ $Y2=0
cc_317 N_A_193_277#_c_178_n N_VGND_c_1004_n 0.00397703f $X=2.09 $Y=1.235 $X2=0
+ $Y2=0
cc_318 N_A_193_277#_c_187_n N_VGND_c_1007_n 0.00313546f $X=5.975 $Y=0.805 $X2=0
+ $Y2=0
cc_319 N_C_N_c_354_n N_A_27_94#_c_391_n 0.00350303f $X=3.315 $Y=1.765 $X2=0
+ $Y2=0
cc_320 N_C_N_c_356_n N_A_27_94#_c_391_n 4.91898e-19 $X=3.54 $Y=1.515 $X2=0 $Y2=0
cc_321 N_C_N_c_354_n N_A_27_94#_c_392_n 0.00672943f $X=3.315 $Y=1.765 $X2=0
+ $Y2=0
cc_322 N_C_N_M1005_g N_A_27_94#_c_392_n 0.012031f $X=3.405 $Y=0.79 $X2=0 $Y2=0
cc_323 N_C_N_c_356_n N_A_27_94#_c_392_n 0.00173987f $X=3.54 $Y=1.515 $X2=0 $Y2=0
cc_324 N_C_N_c_354_n N_A_27_94#_c_396_n 0.00431721f $X=3.315 $Y=1.765 $X2=0
+ $Y2=0
cc_325 N_C_N_M1005_g N_A_27_94#_c_396_n 0.0170424f $X=3.405 $Y=0.79 $X2=0 $Y2=0
cc_326 N_C_N_c_356_n N_A_27_94#_c_396_n 0.0167123f $X=3.54 $Y=1.515 $X2=0 $Y2=0
cc_327 N_C_N_M1005_g N_A_27_94#_c_399_n 9.86457e-19 $X=3.405 $Y=0.79 $X2=0 $Y2=0
cc_328 N_C_N_c_354_n N_A_678_368#_c_553_n 0.00352482f $X=3.315 $Y=1.765 $X2=0
+ $Y2=0
cc_329 N_C_N_c_356_n N_A_678_368#_c_553_n 0.0248792f $X=3.54 $Y=1.515 $X2=0
+ $Y2=0
cc_330 N_C_N_c_354_n N_A_678_368#_c_541_n 0.00349763f $X=3.315 $Y=1.765 $X2=0
+ $Y2=0
cc_331 N_C_N_c_356_n N_A_678_368#_c_541_n 0.0150609f $X=3.54 $Y=1.515 $X2=0
+ $Y2=0
cc_332 N_C_N_c_354_n N_A_678_368#_c_543_n 7.37734e-19 $X=3.315 $Y=1.765 $X2=0
+ $Y2=0
cc_333 N_C_N_c_356_n N_A_678_368#_c_543_n 0.0150668f $X=3.54 $Y=1.515 $X2=0
+ $Y2=0
cc_334 N_C_N_M1005_g N_A_678_368#_c_546_n 0.00414295f $X=3.405 $Y=0.79 $X2=0
+ $Y2=0
cc_335 N_C_N_c_354_n N_VPWR_c_741_n 0.00669475f $X=3.315 $Y=1.765 $X2=0 $Y2=0
cc_336 N_C_N_c_354_n N_VPWR_c_745_n 0.0049405f $X=3.315 $Y=1.765 $X2=0 $Y2=0
cc_337 N_C_N_c_354_n N_VPWR_c_738_n 0.00508379f $X=3.315 $Y=1.765 $X2=0 $Y2=0
cc_338 N_C_N_c_354_n N_A_791_392#_c_877_n 0.00942085f $X=3.315 $Y=1.765 $X2=0
+ $Y2=0
cc_339 N_C_N_M1005_g N_VGND_c_994_n 0.00474761f $X=3.405 $Y=0.79 $X2=0 $Y2=0
cc_340 N_C_N_M1005_g N_VGND_c_1002_n 0.00514438f $X=3.405 $Y=0.79 $X2=0 $Y2=0
cc_341 N_C_N_M1005_g N_VGND_c_1006_n 0.00484614f $X=3.405 $Y=0.79 $X2=0 $Y2=0
cc_342 N_C_N_M1005_g N_VGND_c_1007_n 0.00188628f $X=3.405 $Y=0.79 $X2=0 $Y2=0
cc_343 N_A_27_94#_c_396_n N_A_678_368#_M1005_d 0.00515716f $X=3.945 $Y=1.005
+ $X2=-0.19 $Y2=-0.245
cc_344 N_A_27_94#_c_393_n N_A_678_368#_c_536_n 0.0102597f $X=4.775 $Y=1.795
+ $X2=0 $Y2=0
cc_345 N_A_27_94#_c_403_n N_A_678_368#_c_550_n 0.0448752f $X=4.775 $Y=1.885
+ $X2=0 $Y2=0
cc_346 N_A_27_94#_c_401_n N_A_678_368#_c_553_n 0.00368671f $X=4.325 $Y=1.885
+ $X2=0 $Y2=0
cc_347 N_A_27_94#_c_392_n N_A_678_368#_c_540_n 0.00410571f $X=4.735 $Y=1.185
+ $X2=0 $Y2=0
cc_348 N_A_27_94#_c_399_n N_A_678_368#_c_540_n 0.0247729f $X=4.11 $Y=1.005 $X2=0
+ $Y2=0
cc_349 N_A_27_94#_c_391_n N_A_678_368#_c_541_n 0.00747141f $X=4.325 $Y=1.795
+ $X2=0 $Y2=0
cc_350 N_A_27_94#_c_401_n N_A_678_368#_c_541_n 0.00129524f $X=4.325 $Y=1.885
+ $X2=0 $Y2=0
cc_351 N_A_27_94#_c_391_n N_A_678_368#_c_542_n 0.0121978f $X=4.325 $Y=1.795
+ $X2=0 $Y2=0
cc_352 N_A_27_94#_c_392_n N_A_678_368#_c_542_n 0.0120826f $X=4.735 $Y=1.185
+ $X2=0 $Y2=0
cc_353 N_A_27_94#_c_399_n N_A_678_368#_c_542_n 0.0156872f $X=4.11 $Y=1.005 $X2=0
+ $Y2=0
cc_354 N_A_27_94#_c_392_n N_A_678_368#_c_543_n 0.00488271f $X=4.735 $Y=1.185
+ $X2=0 $Y2=0
cc_355 N_A_27_94#_c_396_n N_A_678_368#_c_543_n 0.0032032f $X=3.945 $Y=1.005
+ $X2=0 $Y2=0
cc_356 N_A_27_94#_c_399_n N_A_678_368#_c_543_n 0.00876668f $X=4.11 $Y=1.005
+ $X2=0 $Y2=0
cc_357 N_A_27_94#_c_392_n N_A_678_368#_c_544_n 0.0164876f $X=4.735 $Y=1.185
+ $X2=0 $Y2=0
cc_358 N_A_27_94#_c_399_n N_A_678_368#_c_544_n 0.0243077f $X=4.11 $Y=1.005 $X2=0
+ $Y2=0
cc_359 N_A_27_94#_c_392_n N_A_678_368#_c_545_n 0.0161378f $X=4.735 $Y=1.185
+ $X2=0 $Y2=0
cc_360 N_A_27_94#_c_393_n N_A_678_368#_c_545_n 0.00723871f $X=4.775 $Y=1.795
+ $X2=0 $Y2=0
cc_361 N_A_27_94#_c_396_n N_A_678_368#_c_546_n 0.0326607f $X=3.945 $Y=1.005
+ $X2=0 $Y2=0
cc_362 N_A_27_94#_c_392_n N_A_678_368#_c_547_n 0.0126745f $X=4.735 $Y=1.185
+ $X2=0 $Y2=0
cc_363 N_A_27_94#_c_392_n N_A_678_368#_c_548_n 0.0102597f $X=4.735 $Y=1.185
+ $X2=0 $Y2=0
cc_364 N_A_27_94#_c_413_n N_VPWR_M1013_d 0.0108196f $X=2.695 $Y=2.475 $X2=-0.19
+ $Y2=-0.245
cc_365 N_A_27_94#_c_413_n N_VPWR_M1010_s 0.00624799f $X=2.695 $Y=2.475 $X2=0
+ $Y2=0
cc_366 N_A_27_94#_c_407_n N_VPWR_M1010_s 0.00135333f $X=2.695 $Y=1.795 $X2=0
+ $Y2=0
cc_367 N_A_27_94#_c_408_n N_VPWR_M1010_s 0.00195263f $X=1.79 $Y=1.795 $X2=0
+ $Y2=0
cc_368 N_A_27_94#_c_413_n N_VPWR_c_739_n 0.0225065f $X=2.695 $Y=2.475 $X2=0
+ $Y2=0
cc_369 N_A_27_94#_c_405_n N_VPWR_c_739_n 0.0088922f $X=0.445 $Y=2.475 $X2=0
+ $Y2=0
cc_370 N_A_27_94#_c_413_n N_VPWR_c_740_n 0.0242551f $X=2.695 $Y=2.475 $X2=0
+ $Y2=0
cc_371 N_A_27_94#_c_413_n N_VPWR_c_741_n 0.00110619f $X=2.695 $Y=2.475 $X2=0
+ $Y2=0
cc_372 N_A_27_94#_c_401_n N_VPWR_c_745_n 0.00291649f $X=4.325 $Y=1.885 $X2=0
+ $Y2=0
cc_373 N_A_27_94#_c_403_n N_VPWR_c_745_n 0.00290311f $X=4.775 $Y=1.885 $X2=0
+ $Y2=0
cc_374 N_A_27_94#_c_401_n N_VPWR_c_738_n 0.00364317f $X=4.325 $Y=1.885 $X2=0
+ $Y2=0
cc_375 N_A_27_94#_c_403_n N_VPWR_c_738_n 0.0035903f $X=4.775 $Y=1.885 $X2=0
+ $Y2=0
cc_376 N_A_27_94#_c_413_n N_VPWR_c_738_n 0.0589664f $X=2.695 $Y=2.475 $X2=0
+ $Y2=0
cc_377 N_A_27_94#_c_405_n N_VPWR_c_738_n 0.0122756f $X=0.445 $Y=2.475 $X2=0
+ $Y2=0
cc_378 N_A_27_94#_c_405_n N_VPWR_c_748_n 0.0107406f $X=0.445 $Y=2.475 $X2=0
+ $Y2=0
cc_379 N_A_27_94#_c_396_n N_X_M1012_s 0.0130244f $X=3.945 $Y=1.005 $X2=0 $Y2=0
cc_380 N_A_27_94#_c_413_n N_X_M1008_d 0.00549025f $X=2.695 $Y=2.475 $X2=0 $Y2=0
cc_381 N_A_27_94#_c_413_n N_X_M1014_d 0.016577f $X=2.695 $Y=2.475 $X2=0 $Y2=0
cc_382 N_A_27_94#_c_407_n N_X_M1014_d 0.00613992f $X=2.695 $Y=1.795 $X2=0 $Y2=0
cc_383 N_A_27_94#_c_413_n N_X_c_827_n 0.0642339f $X=2.695 $Y=2.475 $X2=0 $Y2=0
cc_384 N_A_27_94#_c_407_n N_X_c_827_n 0.0443071f $X=2.695 $Y=1.795 $X2=0 $Y2=0
cc_385 N_A_27_94#_c_408_n N_X_c_827_n 0.0124479f $X=1.79 $Y=1.795 $X2=0 $Y2=0
cc_386 N_A_27_94#_c_396_n N_X_c_836_n 0.0636566f $X=3.945 $Y=1.005 $X2=0 $Y2=0
cc_387 N_A_27_94#_c_515_p N_X_c_836_n 0.0128546f $X=1.79 $Y=1.005 $X2=0 $Y2=0
cc_388 N_A_27_94#_c_408_n X 0.0124843f $X=1.79 $Y=1.795 $X2=0 $Y2=0
cc_389 N_A_27_94#_c_409_n X 0.00251271f $X=0.28 $Y=2.115 $X2=0 $Y2=0
cc_390 N_A_27_94#_c_413_n N_X_c_826_n 0.0199998f $X=2.695 $Y=2.475 $X2=0 $Y2=0
cc_391 N_A_27_94#_c_409_n N_X_c_826_n 0.00450247f $X=0.28 $Y=2.115 $X2=0 $Y2=0
cc_392 N_A_27_94#_c_395_n N_X_c_847_n 0.0447261f $X=1.705 $Y=1.71 $X2=0 $Y2=0
cc_393 N_A_27_94#_c_401_n N_A_791_392#_c_877_n 0.0132453f $X=4.325 $Y=1.885
+ $X2=0 $Y2=0
cc_394 N_A_27_94#_c_403_n N_A_791_392#_c_877_n 0.0160557f $X=4.775 $Y=1.885
+ $X2=0 $Y2=0
cc_395 N_A_27_94#_c_401_n N_A_791_392#_c_878_n 4.4235e-19 $X=4.325 $Y=1.885
+ $X2=0 $Y2=0
cc_396 N_A_27_94#_c_403_n N_A_791_392#_c_878_n 0.00445357f $X=4.775 $Y=1.885
+ $X2=0 $Y2=0
cc_397 N_A_27_94#_c_395_n N_VGND_M1009_d 2.29386e-19 $X=1.705 $Y=1.71 $X2=0
+ $Y2=0
cc_398 N_A_27_94#_c_396_n N_VGND_M1009_d 0.00453009f $X=3.945 $Y=1.005 $X2=0
+ $Y2=0
cc_399 N_A_27_94#_c_515_p N_VGND_M1009_d 0.00287212f $X=1.79 $Y=1.005 $X2=0
+ $Y2=0
cc_400 N_A_27_94#_c_396_n N_VGND_M1018_d 0.00586681f $X=3.945 $Y=1.005 $X2=0
+ $Y2=0
cc_401 N_A_27_94#_c_394_n N_VGND_c_992_n 0.0273776f $X=0.28 $Y=0.615 $X2=0 $Y2=0
cc_402 N_A_27_94#_c_396_n N_VGND_c_994_n 0.0218424f $X=3.945 $Y=1.005 $X2=0
+ $Y2=0
cc_403 N_A_27_94#_c_392_n N_VGND_c_995_n 0.00433162f $X=4.735 $Y=1.185 $X2=0
+ $Y2=0
cc_404 N_A_27_94#_c_394_n N_VGND_c_998_n 0.0113014f $X=0.28 $Y=0.615 $X2=0 $Y2=0
cc_405 N_A_27_94#_c_392_n N_VGND_c_1002_n 0.00826608f $X=4.735 $Y=1.185 $X2=0
+ $Y2=0
cc_406 N_A_27_94#_c_394_n N_VGND_c_1002_n 0.0123744f $X=0.28 $Y=0.615 $X2=0
+ $Y2=0
cc_407 N_A_27_94#_c_392_n N_VGND_c_1007_n 0.00617278f $X=4.735 $Y=1.185 $X2=0
+ $Y2=0
cc_408 N_A_678_368#_M1021_g N_B_M1007_g 0.0220507f $X=6.33 $Y=0.74 $X2=0 $Y2=0
cc_409 N_A_678_368#_c_537_n B 6.83796e-19 $X=5.725 $Y=1.795 $X2=0 $Y2=0
cc_410 N_A_678_368#_c_538_n B 0.00126201f $X=6.255 $Y=1.335 $X2=0 $Y2=0
cc_411 N_A_678_368#_c_550_n N_VPWR_c_745_n 0.00278271f $X=5.225 $Y=1.885 $X2=0
+ $Y2=0
cc_412 N_A_678_368#_c_552_n N_VPWR_c_745_n 0.00278271f $X=5.725 $Y=1.885 $X2=0
+ $Y2=0
cc_413 N_A_678_368#_c_550_n N_VPWR_c_738_n 0.00354368f $X=5.225 $Y=1.885 $X2=0
+ $Y2=0
cc_414 N_A_678_368#_c_552_n N_VPWR_c_738_n 0.00359085f $X=5.725 $Y=1.885 $X2=0
+ $Y2=0
cc_415 N_A_678_368#_c_553_n N_A_791_392#_M1020_s 0.00383711f $X=3.885 $Y=2.035
+ $X2=-0.19 $Y2=-0.245
cc_416 N_A_678_368#_c_550_n N_A_791_392#_c_875_n 0.0111147f $X=5.225 $Y=1.885
+ $X2=0 $Y2=0
cc_417 N_A_678_368#_c_552_n N_A_791_392#_c_875_n 0.0129254f $X=5.725 $Y=1.885
+ $X2=0 $Y2=0
cc_418 N_A_678_368#_c_552_n N_A_791_392#_c_876_n 0.00659721f $X=5.725 $Y=1.885
+ $X2=0 $Y2=0
cc_419 N_A_678_368#_c_550_n N_A_791_392#_c_878_n 0.00682172f $X=5.225 $Y=1.885
+ $X2=0 $Y2=0
cc_420 N_A_678_368#_c_552_n N_A_791_392#_c_878_n 5.29259e-19 $X=5.725 $Y=1.885
+ $X2=0 $Y2=0
cc_421 N_A_678_368#_c_552_n N_A_1060_392#_c_911_n 0.0118723f $X=5.725 $Y=1.885
+ $X2=0 $Y2=0
cc_422 N_A_678_368#_c_552_n N_A_1060_392#_c_910_n 0.0117671f $X=5.725 $Y=1.885
+ $X2=0 $Y2=0
cc_423 N_A_678_368#_c_538_n N_A_1060_392#_c_910_n 0.00549121f $X=6.255 $Y=1.335
+ $X2=0 $Y2=0
cc_424 N_A_678_368#_c_552_n N_A_1273_392#_c_941_n 7.0304e-19 $X=5.725 $Y=1.885
+ $X2=0 $Y2=0
cc_425 N_A_678_368#_c_540_n N_VGND_M1011_s 0.00433267f $X=4.445 $Y=0.665 $X2=0
+ $Y2=0
cc_426 N_A_678_368#_c_544_n N_VGND_M1011_s 0.0101248f $X=4.53 $Y=1.26 $X2=0
+ $Y2=0
cc_427 N_A_678_368#_c_546_n N_VGND_c_994_n 0.0121688f $X=3.785 $Y=0.6 $X2=0
+ $Y2=0
cc_428 N_A_678_368#_M1021_g N_VGND_c_995_n 0.00433162f $X=6.33 $Y=0.74 $X2=0
+ $Y2=0
cc_429 N_A_678_368#_M1021_g N_VGND_c_996_n 0.0073183f $X=6.33 $Y=0.74 $X2=0
+ $Y2=0
cc_430 N_A_678_368#_M1021_g N_VGND_c_1002_n 0.00823168f $X=6.33 $Y=0.74 $X2=0
+ $Y2=0
cc_431 N_A_678_368#_c_540_n N_VGND_c_1002_n 0.0102144f $X=4.445 $Y=0.665 $X2=0
+ $Y2=0
cc_432 N_A_678_368#_c_546_n N_VGND_c_1002_n 0.0110483f $X=3.785 $Y=0.6 $X2=0
+ $Y2=0
cc_433 N_A_678_368#_c_540_n N_VGND_c_1006_n 0.00471384f $X=4.445 $Y=0.665 $X2=0
+ $Y2=0
cc_434 N_A_678_368#_c_546_n N_VGND_c_1006_n 0.0097989f $X=3.785 $Y=0.6 $X2=0
+ $Y2=0
cc_435 N_A_678_368#_c_540_n N_VGND_c_1007_n 0.0454526f $X=4.445 $Y=0.665 $X2=0
+ $Y2=0
cc_436 N_B_M1007_g N_A_c_692_n 0.0190243f $X=6.975 $Y=0.74 $X2=-0.19 $Y2=-0.245
cc_437 B N_A_c_693_n 9.85347e-19 $X=6.875 $Y=1.58 $X2=0 $Y2=0
cc_438 N_B_c_639_n N_A_c_693_n 0.0182767f $X=6.975 $Y=1.667 $X2=0 $Y2=0
cc_439 N_B_c_641_n N_A_c_698_n 0.00887032f $X=7.185 $Y=1.885 $X2=0 $Y2=0
cc_440 N_B_M1007_g A 0.00107976f $X=6.975 $Y=0.74 $X2=0 $Y2=0
cc_441 B A 0.00375953f $X=6.875 $Y=1.58 $X2=0 $Y2=0
cc_442 N_B_c_639_n A 4.5002e-19 $X=6.975 $Y=1.667 $X2=0 $Y2=0
cc_443 B N_A_c_696_n 3.12382e-19 $X=6.875 $Y=1.58 $X2=0 $Y2=0
cc_444 N_B_c_639_n N_A_c_696_n 0.00604191f $X=6.975 $Y=1.667 $X2=0 $Y2=0
cc_445 N_B_c_640_n N_VPWR_c_745_n 0.00278257f $X=6.735 $Y=1.885 $X2=0 $Y2=0
cc_446 N_B_c_641_n N_VPWR_c_745_n 0.00278257f $X=7.185 $Y=1.885 $X2=0 $Y2=0
cc_447 N_B_c_640_n N_VPWR_c_738_n 0.00358623f $X=6.735 $Y=1.885 $X2=0 $Y2=0
cc_448 N_B_c_641_n N_VPWR_c_738_n 0.00353905f $X=7.185 $Y=1.885 $X2=0 $Y2=0
cc_449 N_B_c_640_n N_A_791_392#_c_875_n 7.11409e-19 $X=6.735 $Y=1.885 $X2=0
+ $Y2=0
cc_450 N_B_c_640_n N_A_791_392#_c_876_n 9.78316e-19 $X=6.735 $Y=1.885 $X2=0
+ $Y2=0
cc_451 N_B_c_640_n N_A_1060_392#_c_916_n 0.00452035f $X=6.735 $Y=1.885 $X2=0
+ $Y2=0
cc_452 N_B_c_641_n N_A_1060_392#_c_916_n 0.0017515f $X=7.185 $Y=1.885 $X2=0
+ $Y2=0
cc_453 N_B_c_640_n N_A_1060_392#_c_909_n 0.0171646f $X=6.735 $Y=1.885 $X2=0
+ $Y2=0
cc_454 N_B_c_641_n N_A_1060_392#_c_909_n 0.00136805f $X=7.185 $Y=1.885 $X2=0
+ $Y2=0
cc_455 B N_A_1060_392#_c_909_n 0.0367818f $X=6.875 $Y=1.58 $X2=0 $Y2=0
cc_456 N_B_c_639_n N_A_1060_392#_c_909_n 0.00639846f $X=6.975 $Y=1.667 $X2=0
+ $Y2=0
cc_457 B N_A_1060_392#_c_910_n 0.0104107f $X=6.875 $Y=1.58 $X2=0 $Y2=0
cc_458 N_B_c_640_n N_A_1273_392#_c_939_n 0.00826735f $X=6.735 $Y=1.885 $X2=0
+ $Y2=0
cc_459 N_B_c_641_n N_A_1273_392#_c_939_n 5.25524e-19 $X=7.185 $Y=1.885 $X2=0
+ $Y2=0
cc_460 N_B_c_640_n N_A_1273_392#_c_940_n 0.00868057f $X=6.735 $Y=1.885 $X2=0
+ $Y2=0
cc_461 N_B_c_641_n N_A_1273_392#_c_940_n 0.0125587f $X=7.185 $Y=1.885 $X2=0
+ $Y2=0
cc_462 N_B_c_640_n N_A_1273_392#_c_941_n 0.00376944f $X=6.735 $Y=1.885 $X2=0
+ $Y2=0
cc_463 N_B_c_641_n N_A_1273_392#_c_942_n 0.00378482f $X=7.185 $Y=1.885 $X2=0
+ $Y2=0
cc_464 N_B_c_639_n N_A_1273_392#_c_942_n 7.69601e-19 $X=6.975 $Y=1.667 $X2=0
+ $Y2=0
cc_465 N_B_c_640_n N_A_1273_392#_c_954_n 5.79764e-19 $X=6.735 $Y=1.885 $X2=0
+ $Y2=0
cc_466 N_B_c_641_n N_A_1273_392#_c_954_n 0.00796422f $X=7.185 $Y=1.885 $X2=0
+ $Y2=0
cc_467 N_B_M1007_g N_VGND_c_996_n 0.00863466f $X=6.975 $Y=0.74 $X2=0 $Y2=0
cc_468 N_B_M1007_g N_VGND_c_997_n 7.12736e-19 $X=6.975 $Y=0.74 $X2=0 $Y2=0
cc_469 N_B_M1007_g N_VGND_c_1000_n 0.00434272f $X=6.975 $Y=0.74 $X2=0 $Y2=0
cc_470 N_B_M1007_g N_VGND_c_1002_n 0.00824595f $X=6.975 $Y=0.74 $X2=0 $Y2=0
cc_471 N_A_c_698_n N_VPWR_c_742_n 0.00432608f $X=7.635 $Y=1.885 $X2=0 $Y2=0
cc_472 N_A_c_700_n N_VPWR_c_742_n 0.0120535f $X=8.135 $Y=1.885 $X2=0 $Y2=0
cc_473 N_A_c_698_n N_VPWR_c_745_n 0.0044313f $X=7.635 $Y=1.885 $X2=0 $Y2=0
cc_474 N_A_c_700_n N_VPWR_c_746_n 0.00413917f $X=8.135 $Y=1.885 $X2=0 $Y2=0
cc_475 N_A_c_698_n N_VPWR_c_738_n 0.00853234f $X=7.635 $Y=1.885 $X2=0 $Y2=0
cc_476 N_A_c_700_n N_VPWR_c_738_n 0.00821221f $X=8.135 $Y=1.885 $X2=0 $Y2=0
cc_477 N_A_c_698_n N_A_1273_392#_c_940_n 0.00312124f $X=7.635 $Y=1.885 $X2=0
+ $Y2=0
cc_478 N_A_c_698_n N_A_1273_392#_c_942_n 0.00135864f $X=7.635 $Y=1.885 $X2=0
+ $Y2=0
cc_479 A N_A_1273_392#_c_942_n 0.00217576f $X=8.315 $Y=1.21 $X2=0 $Y2=0
cc_480 N_A_c_696_n N_A_1273_392#_c_942_n 8.44698e-19 $X=8.37 $Y=1.385 $X2=0
+ $Y2=0
cc_481 N_A_c_698_n N_A_1273_392#_c_954_n 0.00798141f $X=7.635 $Y=1.885 $X2=0
+ $Y2=0
cc_482 N_A_c_700_n N_A_1273_392#_c_954_n 2.70506e-19 $X=8.135 $Y=1.885 $X2=0
+ $Y2=0
cc_483 N_A_c_698_n N_A_1273_392#_c_943_n 0.0175539f $X=7.635 $Y=1.885 $X2=0
+ $Y2=0
cc_484 N_A_c_700_n N_A_1273_392#_c_943_n 0.0170908f $X=8.135 $Y=1.885 $X2=0
+ $Y2=0
cc_485 A N_A_1273_392#_c_943_n 0.0247357f $X=8.315 $Y=1.21 $X2=0 $Y2=0
cc_486 N_A_c_696_n N_A_1273_392#_c_943_n 0.00270933f $X=8.37 $Y=1.385 $X2=0
+ $Y2=0
cc_487 N_A_c_700_n N_A_1273_392#_c_944_n 0.00245361f $X=8.135 $Y=1.885 $X2=0
+ $Y2=0
cc_488 A N_A_1273_392#_c_944_n 0.0148879f $X=8.315 $Y=1.21 $X2=0 $Y2=0
cc_489 N_A_c_696_n N_A_1273_392#_c_944_n 0.00607805f $X=8.37 $Y=1.385 $X2=0
+ $Y2=0
cc_490 N_A_c_700_n N_A_1273_392#_c_945_n 6.79657e-19 $X=8.135 $Y=1.885 $X2=0
+ $Y2=0
cc_491 N_A_c_692_n N_VGND_c_997_n 0.0147238f $X=7.59 $Y=1.22 $X2=0 $Y2=0
cc_492 A N_VGND_c_997_n 0.0503712f $X=8.315 $Y=1.21 $X2=0 $Y2=0
cc_493 N_A_c_696_n N_VGND_c_997_n 0.00433572f $X=8.37 $Y=1.385 $X2=0 $Y2=0
cc_494 N_A_c_692_n N_VGND_c_1000_n 0.00383152f $X=7.59 $Y=1.22 $X2=0 $Y2=0
cc_495 N_A_c_692_n N_VGND_c_1002_n 0.00759105f $X=7.59 $Y=1.22 $X2=0 $Y2=0
cc_496 N_VPWR_M1010_s N_X_c_827_n 0.00607354f $X=1.58 $Y=1.84 $X2=0 $Y2=0
cc_497 N_VPWR_c_745_n N_A_791_392#_c_875_n 0.0178297f $X=7.745 $Y=3.33 $X2=0
+ $Y2=0
cc_498 N_VPWR_c_738_n N_A_791_392#_c_875_n 0.00970209f $X=8.4 $Y=3.33 $X2=0
+ $Y2=0
cc_499 N_VPWR_c_745_n N_A_791_392#_c_877_n 0.0373432f $X=7.745 $Y=3.33 $X2=0
+ $Y2=0
cc_500 N_VPWR_c_738_n N_A_791_392#_c_877_n 0.0311309f $X=8.4 $Y=3.33 $X2=0 $Y2=0
cc_501 N_VPWR_c_745_n N_A_791_392#_c_878_n 0.066876f $X=7.745 $Y=3.33 $X2=0
+ $Y2=0
cc_502 N_VPWR_c_738_n N_A_791_392#_c_878_n 0.0375607f $X=8.4 $Y=3.33 $X2=0 $Y2=0
cc_503 N_VPWR_c_742_n N_A_1273_392#_c_940_n 0.0119239f $X=7.91 $Y=2.495 $X2=0
+ $Y2=0
cc_504 N_VPWR_c_745_n N_A_1273_392#_c_940_n 0.0594312f $X=7.745 $Y=3.33 $X2=0
+ $Y2=0
cc_505 N_VPWR_c_738_n N_A_1273_392#_c_940_n 0.0328875f $X=8.4 $Y=3.33 $X2=0
+ $Y2=0
cc_506 N_VPWR_c_745_n N_A_1273_392#_c_941_n 0.0234827f $X=7.745 $Y=3.33 $X2=0
+ $Y2=0
cc_507 N_VPWR_c_738_n N_A_1273_392#_c_941_n 0.0127381f $X=8.4 $Y=3.33 $X2=0
+ $Y2=0
cc_508 N_VPWR_M1017_s N_A_1273_392#_c_943_n 0.00255032f $X=7.71 $Y=1.96 $X2=0
+ $Y2=0
cc_509 N_VPWR_c_742_n N_A_1273_392#_c_943_n 0.0209821f $X=7.91 $Y=2.495 $X2=0
+ $Y2=0
cc_510 N_VPWR_c_742_n N_A_1273_392#_c_945_n 0.0224125f $X=7.91 $Y=2.495 $X2=0
+ $Y2=0
cc_511 N_VPWR_c_746_n N_A_1273_392#_c_945_n 0.0126901f $X=8.4 $Y=3.33 $X2=0
+ $Y2=0
cc_512 N_VPWR_c_738_n N_A_1273_392#_c_945_n 0.010143f $X=8.4 $Y=3.33 $X2=0 $Y2=0
cc_513 N_X_c_836_n N_VGND_M1009_d 0.00717704f $X=2.14 $Y=0.585 $X2=0 $Y2=0
cc_514 N_X_c_821_n N_VGND_c_992_n 0.0520689f $X=1.285 $Y=0.515 $X2=0 $Y2=0
cc_515 N_X_c_821_n N_VGND_c_993_n 0.0144922f $X=1.285 $Y=0.515 $X2=0 $Y2=0
cc_516 N_X_c_836_n N_VGND_c_993_n 0.0029521f $X=2.14 $Y=0.585 $X2=0 $Y2=0
cc_517 N_X_c_831_n N_VGND_c_999_n 0.0192751f $X=2.305 $Y=0.585 $X2=0 $Y2=0
cc_518 N_X_c_836_n N_VGND_c_999_n 0.00294479f $X=2.14 $Y=0.585 $X2=0 $Y2=0
cc_519 N_X_c_831_n N_VGND_c_1002_n 0.0216949f $X=2.305 $Y=0.585 $X2=0 $Y2=0
cc_520 N_X_c_821_n N_VGND_c_1002_n 0.0118826f $X=1.285 $Y=0.515 $X2=0 $Y2=0
cc_521 N_X_c_836_n N_VGND_c_1002_n 0.0111994f $X=2.14 $Y=0.585 $X2=0 $Y2=0
cc_522 N_X_c_821_n N_VGND_c_1004_n 0.0029097f $X=1.285 $Y=0.515 $X2=0 $Y2=0
cc_523 N_X_c_836_n N_VGND_c_1004_n 0.0243979f $X=2.14 $Y=0.585 $X2=0 $Y2=0
cc_524 N_A_791_392#_c_875_n N_A_1060_392#_M1001_d 0.00250873f $X=5.865 $Y=2.99
+ $X2=-0.19 $Y2=1.66
cc_525 N_A_791_392#_c_875_n N_A_1060_392#_c_911_n 0.0188235f $X=5.865 $Y=2.99
+ $X2=0 $Y2=0
cc_526 N_A_791_392#_c_876_n N_A_1060_392#_c_911_n 0.0197801f $X=5.95 $Y=2.605
+ $X2=0 $Y2=0
cc_527 N_A_791_392#_M1002_s N_A_1060_392#_c_910_n 0.006022f $X=5.8 $Y=1.96 $X2=0
+ $Y2=0
cc_528 N_A_791_392#_c_875_n N_A_1060_392#_c_910_n 0.00325039f $X=5.865 $Y=2.99
+ $X2=0 $Y2=0
cc_529 N_A_791_392#_c_876_n N_A_1060_392#_c_910_n 0.0201229f $X=5.95 $Y=2.605
+ $X2=0 $Y2=0
cc_530 N_A_791_392#_c_876_n N_A_1273_392#_c_939_n 0.0306384f $X=5.95 $Y=2.605
+ $X2=0 $Y2=0
cc_531 N_A_791_392#_c_875_n N_A_1273_392#_c_941_n 0.0128665f $X=5.865 $Y=2.99
+ $X2=0 $Y2=0
cc_532 N_A_1060_392#_c_909_n N_A_1273_392#_M1015_s 0.00634569f $X=6.96 $Y=2.115
+ $X2=-0.19 $Y2=1.66
cc_533 N_A_1060_392#_c_910_n N_A_1273_392#_M1015_s 0.00623141f $X=6.575 $Y=2.11
+ $X2=-0.19 $Y2=1.66
cc_534 N_A_1060_392#_c_916_n N_A_1273_392#_c_939_n 0.0192154f $X=6.96 $Y=2.57
+ $X2=0 $Y2=0
cc_535 N_A_1060_392#_c_910_n N_A_1273_392#_c_939_n 0.0219832f $X=6.575 $Y=2.11
+ $X2=0 $Y2=0
cc_536 N_A_1060_392#_M1015_d N_A_1273_392#_c_940_n 0.00227576f $X=6.81 $Y=1.96
+ $X2=0 $Y2=0
cc_537 N_A_1060_392#_c_916_n N_A_1273_392#_c_940_n 0.012422f $X=6.96 $Y=2.57
+ $X2=0 $Y2=0
cc_538 N_A_1060_392#_c_909_n N_A_1273_392#_c_940_n 0.00347484f $X=6.96 $Y=2.115
+ $X2=0 $Y2=0
cc_539 N_A_1060_392#_c_909_n N_A_1273_392#_c_942_n 0.0219546f $X=6.96 $Y=2.115
+ $X2=0 $Y2=0
cc_540 N_A_1060_392#_c_916_n N_A_1273_392#_c_954_n 0.0302886f $X=6.96 $Y=2.57
+ $X2=0 $Y2=0
cc_541 N_A_1060_392#_c_909_n N_A_1273_392#_c_954_n 0.0020791f $X=6.96 $Y=2.115
+ $X2=0 $Y2=0
