# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_hs__dlrtn_2
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_hs__dlrtn_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  8.160000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.208500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.435000 1.450000 0.835000 1.780000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.543200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.845000 1.820000 7.535000 2.980000 ;
        RECT 7.205000 0.350000 7.535000 1.470000 ;
        RECT 7.365000 1.470000 7.535000 1.820000 ;
    END
  END Q
  PIN RESET_B
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.885000 1.180000 6.305000 1.550000 ;
    END
  END RESET_B
  PIN GATE_N
    ANTENNAGATEAREA  0.237000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 1.005000 1.450000 1.335000 1.780000 ;
    END
  END GATE_N
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 8.160000 0.085000 ;
        RECT 0.625000  0.085000 0.955000 0.410000 ;
        RECT 2.380000  0.085000 3.280000 0.410000 ;
        RECT 4.750000  0.085000 5.080000 0.680000 ;
        RECT 6.130000  0.085000 7.035000 1.010000 ;
        RECT 7.705000  0.085000 8.035000 1.130000 ;
      LAYER mcon ;
        RECT 0.155000 -0.085000 0.325000 0.085000 ;
        RECT 0.635000 -0.085000 0.805000 0.085000 ;
        RECT 1.115000 -0.085000 1.285000 0.085000 ;
        RECT 1.595000 -0.085000 1.765000 0.085000 ;
        RECT 2.075000 -0.085000 2.245000 0.085000 ;
        RECT 2.555000 -0.085000 2.725000 0.085000 ;
        RECT 3.035000 -0.085000 3.205000 0.085000 ;
        RECT 3.515000 -0.085000 3.685000 0.085000 ;
        RECT 3.995000 -0.085000 4.165000 0.085000 ;
        RECT 4.475000 -0.085000 4.645000 0.085000 ;
        RECT 4.955000 -0.085000 5.125000 0.085000 ;
        RECT 5.435000 -0.085000 5.605000 0.085000 ;
        RECT 5.915000 -0.085000 6.085000 0.085000 ;
        RECT 6.395000 -0.085000 6.565000 0.085000 ;
        RECT 6.875000 -0.085000 7.045000 0.085000 ;
        RECT 7.355000 -0.085000 7.525000 0.085000 ;
        RECT 7.835000 -0.085000 8.005000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.245000 8.160000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 3.245000 8.160000 3.415000 ;
        RECT 0.785000 1.950000 1.115000 3.245000 ;
        RECT 2.380000 2.860000 2.710000 3.245000 ;
        RECT 4.715000 2.630000 5.545000 3.245000 ;
        RECT 6.320000 2.060000 6.650000 3.245000 ;
        RECT 7.705000 1.820000 8.045000 3.245000 ;
      LAYER mcon ;
        RECT 0.155000 3.245000 0.325000 3.415000 ;
        RECT 0.635000 3.245000 0.805000 3.415000 ;
        RECT 1.115000 3.245000 1.285000 3.415000 ;
        RECT 1.595000 3.245000 1.765000 3.415000 ;
        RECT 2.075000 3.245000 2.245000 3.415000 ;
        RECT 2.555000 3.245000 2.725000 3.415000 ;
        RECT 3.035000 3.245000 3.205000 3.415000 ;
        RECT 3.515000 3.245000 3.685000 3.415000 ;
        RECT 3.995000 3.245000 4.165000 3.415000 ;
        RECT 4.475000 3.245000 4.645000 3.415000 ;
        RECT 4.955000 3.245000 5.125000 3.415000 ;
        RECT 5.435000 3.245000 5.605000 3.415000 ;
        RECT 5.915000 3.245000 6.085000 3.415000 ;
        RECT 6.395000 3.245000 6.565000 3.415000 ;
        RECT 6.875000 3.245000 7.045000 3.415000 ;
        RECT 7.355000 3.245000 7.525000 3.415000 ;
        RECT 7.835000 3.245000 8.005000 3.415000 ;
      LAYER met1 ;
        RECT 0.000000 3.085000 8.160000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.095000 0.580000 2.945000 0.750000 ;
      RECT 0.095000 0.750000 0.445000 1.250000 ;
      RECT 0.095000 1.250000 0.265000 1.950000 ;
      RECT 0.095000 1.950000 0.615000 2.830000 ;
      RECT 1.135000 0.920000 1.675000 1.250000 ;
      RECT 1.285000 1.950000 1.675000 2.520000 ;
      RECT 1.285000 2.520000 4.325000 2.690000 ;
      RECT 1.285000 2.690000 1.675000 2.830000 ;
      RECT 1.505000 1.250000 1.675000 1.340000 ;
      RECT 1.505000 1.340000 1.905000 1.670000 ;
      RECT 1.505000 1.670000 1.675000 1.950000 ;
      RECT 1.845000 0.920000 2.245000 1.170000 ;
      RECT 1.845000 1.840000 3.485000 2.010000 ;
      RECT 1.845000 2.010000 2.245000 2.350000 ;
      RECT 2.075000 1.170000 2.245000 1.840000 ;
      RECT 2.615000 0.750000 2.945000 1.590000 ;
      RECT 3.155000 1.190000 4.415000 1.520000 ;
      RECT 3.155000 1.520000 3.485000 1.840000 ;
      RECT 3.335000 2.180000 3.825000 2.350000 ;
      RECT 3.655000 1.690000 5.375000 1.860000 ;
      RECT 3.655000 1.860000 3.825000 2.180000 ;
      RECT 3.895000 0.350000 4.225000 0.850000 ;
      RECT 3.895000 0.850000 5.140000 1.020000 ;
      RECT 3.995000 2.030000 4.325000 2.520000 ;
      RECT 4.565000 2.030000 6.045000 2.360000 ;
      RECT 4.970000 1.020000 5.140000 1.350000 ;
      RECT 4.970000 1.350000 5.375000 1.690000 ;
      RECT 5.310000 0.350000 5.715000 1.130000 ;
      RECT 5.545000 1.130000 5.715000 1.720000 ;
      RECT 5.545000 1.720000 6.675000 1.890000 ;
      RECT 5.545000 1.890000 6.045000 2.030000 ;
      RECT 5.715000 2.360000 6.045000 2.980000 ;
      RECT 6.505000 1.320000 6.845000 1.650000 ;
      RECT 6.505000 1.650000 6.675000 1.720000 ;
  END
END sky130_fd_sc_hs__dlrtn_2
