# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_hs__nor4bb_1
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_hs__nor4bb_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.800000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.075000 1.350000 1.405000 2.150000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.915000 1.350000 2.275000 1.780000 ;
    END
  END B
  PIN C_N
    ANTENNAGATEAREA  0.208500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105000 1.180000 0.435000 1.550000 ;
    END
  END C_N
  PIN D_N
    ANTENNAGATEAREA  0.208500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.965000 1.450000 4.345000 1.780000 ;
    END
  END D_N
  PIN Y
    ANTENNADIFFAREA  0.848400 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.445000 0.350000 1.775000 0.880000 ;
        RECT 1.445000 0.880000 3.235000 1.050000 ;
        RECT 1.445000 1.050000 1.775000 1.130000 ;
        RECT 1.575000 1.130000 1.745000 2.060000 ;
        RECT 1.575000 2.060000 3.455000 2.390000 ;
        RECT 2.860000 0.350000 3.235000 0.880000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 4.800000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 4.800000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.800000 0.085000 ;
      RECT 0.000000  3.245000 4.800000 3.415000 ;
      RECT 0.115000  0.680000 0.775000 1.010000 ;
      RECT 0.115000  1.820000 0.775000 2.560000 ;
      RECT 0.115000  2.560000 3.795000 2.730000 ;
      RECT 0.605000  1.010000 0.775000 1.820000 ;
      RECT 0.650000  2.900000 1.345000 3.245000 ;
      RECT 0.945000  0.085000 1.275000 1.130000 ;
      RECT 1.945000  0.085000 2.690000 0.680000 ;
      RECT 2.485000  1.350000 2.815000 1.720000 ;
      RECT 2.485000  1.720000 3.795000 1.890000 ;
      RECT 3.070000  1.220000 4.685000 1.260000 ;
      RECT 3.070000  1.260000 3.740000 1.550000 ;
      RECT 3.405000  0.085000 4.175000 0.920000 ;
      RECT 3.570000  1.090000 4.685000 1.220000 ;
      RECT 3.625000  1.890000 3.795000 2.560000 ;
      RECT 3.965000  2.100000 4.185000 3.245000 ;
      RECT 4.355000  0.540000 4.685000 1.090000 ;
      RECT 4.355000  2.100000 4.685000 2.980000 ;
      RECT 4.515000  1.260000 4.685000 2.100000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
  END
END sky130_fd_sc_hs__nor4bb_1
END LIBRARY
