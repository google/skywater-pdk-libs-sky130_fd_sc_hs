* File: sky130_fd_sc_hs__a211o_4.pex.spice
* Created: Thu Aug 27 20:23:33 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HS__A211O_4%A_105_280# 1 2 3 4 13 15 16 18 20 23 25 27
+ 28 30 31 33 34 36 37 39 40 42 45 48 49 51 53 57 59 61 63 65 69 75
c170 75 0 1.0197e-19 $X=5.89 $Y=1.105
c171 61 0 1.45535e-19 $X=5.725 $Y=1.195
c172 57 0 1.44395e-19 $X=3.195 $Y=0.615
c173 45 0 6.27654e-20 $X=2.13 $Y=1.385
r174 83 84 14.9641 $w=3.06e-07 $l=9.5e-08 $layer=POLY_cond $X=1.965 $Y=1.492
+ $X2=2.06 $Y2=1.492
r175 82 83 52.768 $w=3.06e-07 $l=3.35e-07 $layer=POLY_cond $X=1.63 $Y=1.492
+ $X2=1.965 $Y2=1.492
r176 81 82 18.1144 $w=3.06e-07 $l=1.15e-07 $layer=POLY_cond $X=1.515 $Y=1.492
+ $X2=1.63 $Y2=1.492
r177 75 77 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=5.89 $Y=1.105
+ $X2=5.89 $Y2=1.195
r178 65 66 12.4848 $w=2.38e-07 $l=2.6e-07 $layer=LI1_cond $X=3.16 $Y=0.955
+ $X2=3.16 $Y2=1.215
r179 62 72 3.76007 $w=1.7e-07 $l=1.43e-07 $layer=LI1_cond $X=4.245 $Y=1.195
+ $X2=4.102 $Y2=1.195
r180 61 77 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.725 $Y=1.195
+ $X2=5.89 $Y2=1.195
r181 61 62 96.5562 $w=1.68e-07 $l=1.48e-06 $layer=LI1_cond $X=5.725 $Y=1.195
+ $X2=4.245 $Y2=1.195
r182 60 65 2.75731 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=3.28 $Y=0.955
+ $X2=3.16 $Y2=0.955
r183 59 72 9.70478 $w=2.83e-07 $l=2.4e-07 $layer=LI1_cond $X=4.102 $Y=0.955
+ $X2=4.102 $Y2=1.195
r184 59 69 2.4262 $w=2.83e-07 $l=6e-08 $layer=LI1_cond $X=4.102 $Y=0.955
+ $X2=4.102 $Y2=0.895
r185 59 60 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=3.96 $Y=0.955
+ $X2=3.28 $Y2=0.955
r186 55 65 4.08157 $w=2.38e-07 $l=8.5e-08 $layer=LI1_cond $X=3.16 $Y=0.87
+ $X2=3.16 $Y2=0.955
r187 55 57 12.2447 $w=2.38e-07 $l=2.55e-07 $layer=LI1_cond $X=3.16 $Y=0.87
+ $X2=3.16 $Y2=0.615
r188 51 53 68.1765 $w=1.68e-07 $l=1.045e-06 $layer=LI1_cond $X=2.615 $Y=2.145
+ $X2=3.66 $Y2=2.145
r189 50 63 3.19717 $w=2.95e-07 $l=1.62019e-07 $layer=LI1_cond $X=2.615 $Y=1.215
+ $X2=2.53 $Y2=1.34
r190 49 66 2.75731 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=3.04 $Y=1.215
+ $X2=3.16 $Y2=1.215
r191 49 50 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=3.04 $Y=1.215
+ $X2=2.615 $Y2=1.215
r192 48 51 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.53 $Y=2.06
+ $X2=2.615 $Y2=2.145
r193 47 63 3.3845 $w=1.7e-07 $l=2.1e-07 $layer=LI1_cond $X=2.53 $Y=1.55 $X2=2.53
+ $Y2=1.34
r194 47 48 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=2.53 $Y=1.55
+ $X2=2.53 $Y2=2.06
r195 45 84 11.0261 $w=3.06e-07 $l=7e-08 $layer=POLY_cond $X=2.13 $Y=1.492
+ $X2=2.06 $Y2=1.492
r196 44 45 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.13
+ $Y=1.385 $X2=2.13 $Y2=1.385
r197 42 63 3.19717 $w=2.95e-07 $l=8.5e-08 $layer=LI1_cond $X=2.445 $Y=1.34
+ $X2=2.53 $Y2=1.34
r198 42 44 8.64332 $w=4.18e-07 $l=3.15e-07 $layer=LI1_cond $X=2.445 $Y=1.34
+ $X2=2.13 $Y2=1.34
r199 37 45 56.7059 $w=3.06e-07 $l=4.76991e-07 $layer=POLY_cond $X=2.49 $Y=1.22
+ $X2=2.13 $Y2=1.492
r200 37 39 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=2.49 $Y=1.22
+ $X2=2.49 $Y2=0.74
r201 34 84 19.4347 $w=1.5e-07 $l=2.72e-07 $layer=POLY_cond $X=2.06 $Y=1.22
+ $X2=2.06 $Y2=1.492
r202 34 36 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=2.06 $Y=1.22
+ $X2=2.06 $Y2=0.74
r203 31 83 19.4347 $w=1.5e-07 $l=2.73e-07 $layer=POLY_cond $X=1.965 $Y=1.765
+ $X2=1.965 $Y2=1.492
r204 31 33 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.965 $Y=1.765
+ $X2=1.965 $Y2=2.4
r205 28 82 19.4347 $w=1.5e-07 $l=2.72e-07 $layer=POLY_cond $X=1.63 $Y=1.22
+ $X2=1.63 $Y2=1.492
r206 28 30 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.63 $Y=1.22
+ $X2=1.63 $Y2=0.74
r207 25 81 19.4347 $w=1.5e-07 $l=2.73e-07 $layer=POLY_cond $X=1.515 $Y=1.765
+ $X2=1.515 $Y2=1.492
r208 25 27 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.515 $Y=1.765
+ $X2=1.515 $Y2=2.4
r209 21 81 49.6176 $w=3.06e-07 $l=3.15e-07 $layer=POLY_cond $X=1.2 $Y=1.492
+ $X2=1.515 $Y2=1.492
r210 21 79 21.2647 $w=3.06e-07 $l=1.35e-07 $layer=POLY_cond $X=1.2 $Y=1.492
+ $X2=1.065 $Y2=1.492
r211 21 23 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.2 $Y=1.4 $X2=1.2
+ $Y2=0.74
r212 18 79 19.4347 $w=1.5e-07 $l=2.73e-07 $layer=POLY_cond $X=1.065 $Y=1.765
+ $X2=1.065 $Y2=1.492
r213 18 20 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.065 $Y=1.765
+ $X2=1.065 $Y2=2.4
r214 17 40 7.1379 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=0.705 $Y=1.475
+ $X2=0.615 $Y2=1.475
r215 16 79 26.7213 $w=3.06e-07 $l=9.81326e-08 $layer=POLY_cond $X=0.975 $Y=1.475
+ $X2=1.065 $Y2=1.492
r216 16 17 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=0.975 $Y=1.475
+ $X2=0.705 $Y2=1.475
r217 13 40 114.876 $w=1.8e-07 $l=2.9e-07 $layer=POLY_cond $X=0.615 $Y=1.765
+ $X2=0.615 $Y2=1.475
r218 13 15 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.615 $Y=1.765
+ $X2=0.615 $Y2=2.4
r219 4 53 600 $w=1.7e-07 $l=2.48948e-07 $layer=licon1_PDIFF $count=1 $X=3.51
+ $Y=1.96 $X2=3.66 $Y2=2.145
r220 3 75 182 $w=1.7e-07 $l=5.55608e-07 $layer=licon1_NDIFF $count=1 $X=5.75
+ $Y=0.615 $X2=5.89 $Y2=1.105
r221 2 69 182 $w=1.7e-07 $l=4.29651e-07 $layer=licon1_NDIFF $count=1 $X=3.975
+ $Y=0.54 $X2=4.14 $Y2=0.895
r222 1 65 182 $w=1.7e-07 $l=5.60647e-07 $layer=licon1_NDIFF $count=1 $X=3.055
+ $Y=0.47 $X2=3.195 $Y2=0.965
r223 1 57 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=3.055
+ $Y=0.47 $X2=3.195 $Y2=0.615
.ends

.subckt PM_SKY130_FD_SC_HS__A211O_4%B1 1 3 6 8 10 13 15 18 23 24
c96 18 0 1.35305e-19 $X=2.94 $Y=1.635
c97 13 0 7.83994e-20 $X=4.375 $Y=0.935
c98 8 0 6.11229e-20 $X=4.36 $Y=1.885
r99 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.35
+ $Y=1.635 $X2=4.35 $Y2=1.635
r100 24 34 6.74519 $w=4.16e-07 $l=2.995e-07 $layer=LI1_cond $X=4.08 $Y=2.035
+ $X2=4.24 $Y2=1.805
r101 23 34 4.10577 $w=4.16e-07 $l=1.4e-07 $layer=LI1_cond $X=4.24 $Y=1.665
+ $X2=4.24 $Y2=1.805
r102 23 30 0.879808 $w=4.16e-07 $l=3e-08 $layer=LI1_cond $X=4.24 $Y=1.665
+ $X2=4.24 $Y2=1.635
r103 18 21 6.12235 $w=3.18e-07 $l=1.7e-07 $layer=LI1_cond $X=2.945 $Y=1.635
+ $X2=2.945 $Y2=1.805
r104 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.94
+ $Y=1.635 $X2=2.94 $Y2=1.635
r105 16 21 4.44149 $w=1.7e-07 $l=1.6e-07 $layer=LI1_cond $X=3.105 $Y=1.805
+ $X2=2.945 $Y2=1.805
r106 15 34 6.01746 $w=1.7e-07 $l=2.75e-07 $layer=LI1_cond $X=3.965 $Y=1.805
+ $X2=4.24 $Y2=1.805
r107 15 16 56.107 $w=1.68e-07 $l=8.6e-07 $layer=LI1_cond $X=3.965 $Y=1.805
+ $X2=3.105 $Y2=1.805
r108 11 29 38.5562 $w=2.99e-07 $l=1.77059e-07 $layer=POLY_cond $X=4.375 $Y=1.47
+ $X2=4.35 $Y2=1.635
r109 11 13 274.33 $w=1.5e-07 $l=5.35e-07 $layer=POLY_cond $X=4.375 $Y=1.47
+ $X2=4.375 $Y2=0.935
r110 8 29 52.2586 $w=2.99e-07 $l=2.54951e-07 $layer=POLY_cond $X=4.36 $Y=1.885
+ $X2=4.35 $Y2=1.635
r111 8 10 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=4.36 $Y=1.885
+ $X2=4.36 $Y2=2.46
r112 4 19 38.5562 $w=2.99e-07 $l=1.83916e-07 $layer=POLY_cond $X=2.98 $Y=1.47
+ $X2=2.94 $Y2=1.635
r113 4 6 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=2.98 $Y=1.47 $X2=2.98
+ $Y2=0.79
r114 1 19 52.2586 $w=2.99e-07 $l=2.52488e-07 $layer=POLY_cond $X=2.935 $Y=1.885
+ $X2=2.94 $Y2=1.635
r115 1 3 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=2.935 $Y=1.885
+ $X2=2.935 $Y2=2.46
.ends

.subckt PM_SKY130_FD_SC_HS__A211O_4%C1 3 6 7 9 11 12 14 15 17 18 27
c63 18 0 5.16691e-20 $X=3.6 $Y=1.295
c64 15 0 1.3059e-19 $X=3.9 $Y=1.29
c65 7 0 7.25396e-20 $X=3.435 $Y=1.885
c66 3 0 1.44395e-19 $X=3.41 $Y=0.79
r67 26 27 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=3.885 $Y=1.455
+ $X2=3.9 $Y2=1.455
r68 24 26 47.2125 $w=3.3e-07 $l=2.7e-07 $layer=POLY_cond $X=3.615 $Y=1.455
+ $X2=3.885 $Y2=1.455
r69 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.615
+ $Y=1.455 $X2=3.615 $Y2=1.455
r70 22 24 31.475 $w=3.3e-07 $l=1.8e-07 $layer=POLY_cond $X=3.435 $Y=1.455
+ $X2=3.615 $Y2=1.455
r71 20 22 4.37153 $w=3.3e-07 $l=2.5e-08 $layer=POLY_cond $X=3.41 $Y=1.455
+ $X2=3.435 $Y2=1.455
r72 18 25 5.5876 $w=3.28e-07 $l=1.6e-07 $layer=LI1_cond $X=3.615 $Y=1.295
+ $X2=3.615 $Y2=1.455
r73 15 27 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.9 $Y=1.29 $X2=3.9
+ $Y2=1.455
r74 15 17 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=3.9 $Y=1.29 $X2=3.9
+ $Y2=0.86
r75 12 14 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=3.885 $Y=1.885
+ $X2=3.885 $Y2=2.46
r76 11 12 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=3.885 $Y=1.795
+ $X2=3.885 $Y2=1.885
r77 10 26 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=3.885 $Y=1.62
+ $X2=3.885 $Y2=1.455
r78 10 11 68.0242 $w=1.8e-07 $l=1.75e-07 $layer=POLY_cond $X=3.885 $Y=1.62
+ $X2=3.885 $Y2=1.795
r79 7 9 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=3.435 $Y=1.885
+ $X2=3.435 $Y2=2.46
r80 6 7 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=3.435 $Y=1.795 $X2=3.435
+ $Y2=1.885
r81 5 22 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=3.435 $Y=1.62
+ $X2=3.435 $Y2=1.455
r82 5 6 68.0242 $w=1.8e-07 $l=1.75e-07 $layer=POLY_cond $X=3.435 $Y=1.62
+ $X2=3.435 $Y2=1.795
r83 1 20 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.41 $Y=1.29
+ $X2=3.41 $Y2=1.455
r84 1 3 256.383 $w=1.5e-07 $l=5e-07 $layer=POLY_cond $X=3.41 $Y=1.29 $X2=3.41
+ $Y2=0.79
.ends

.subckt PM_SKY130_FD_SC_HS__A211O_4%A1 1 3 6 8 10 13 15 16 17 26
c52 17 0 8.78532e-20 $X=6 $Y=1.665
c53 13 0 1.54739e-19 $X=6.105 $Y=0.935
c54 8 0 2.23913e-19 $X=6.07 $Y=1.885
c55 6 0 1.25287e-19 $X=5.675 $Y=0.935
c56 1 0 1.60917e-19 $X=5.62 $Y=1.885
r57 26 27 4.34794 $w=3.88e-07 $l=3.5e-08 $layer=POLY_cond $X=6.07 $Y=1.667
+ $X2=6.105 $Y2=1.667
r58 24 26 46.5851 $w=3.88e-07 $l=3.75e-07 $layer=POLY_cond $X=5.695 $Y=1.667
+ $X2=6.07 $Y2=1.667
r59 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.695
+ $Y=1.615 $X2=5.695 $Y2=1.615
r60 22 24 2.48454 $w=3.88e-07 $l=2e-08 $layer=POLY_cond $X=5.675 $Y=1.667
+ $X2=5.695 $Y2=1.667
r61 21 22 6.83247 $w=3.88e-07 $l=5.5e-08 $layer=POLY_cond $X=5.62 $Y=1.667
+ $X2=5.675 $Y2=1.667
r62 17 25 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=6 $Y=1.615
+ $X2=5.695 $Y2=1.615
r63 16 25 6.11144 $w=3.28e-07 $l=1.75e-07 $layer=LI1_cond $X=5.52 $Y=1.615
+ $X2=5.695 $Y2=1.615
r64 15 16 16.7628 $w=3.28e-07 $l=4.8e-07 $layer=LI1_cond $X=5.04 $Y=1.615
+ $X2=5.52 $Y2=1.615
r65 11 27 25.1189 $w=1.5e-07 $l=2.17e-07 $layer=POLY_cond $X=6.105 $Y=1.45
+ $X2=6.105 $Y2=1.667
r66 11 13 264.074 $w=1.5e-07 $l=5.15e-07 $layer=POLY_cond $X=6.105 $Y=1.45
+ $X2=6.105 $Y2=0.935
r67 8 26 25.1189 $w=1.5e-07 $l=2.18e-07 $layer=POLY_cond $X=6.07 $Y=1.885
+ $X2=6.07 $Y2=1.667
r68 8 10 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=6.07 $Y=1.885
+ $X2=6.07 $Y2=2.46
r69 4 22 25.1189 $w=1.5e-07 $l=2.17e-07 $layer=POLY_cond $X=5.675 $Y=1.45
+ $X2=5.675 $Y2=1.667
r70 4 6 264.074 $w=1.5e-07 $l=5.15e-07 $layer=POLY_cond $X=5.675 $Y=1.45
+ $X2=5.675 $Y2=0.935
r71 1 21 25.1189 $w=1.5e-07 $l=2.18e-07 $layer=POLY_cond $X=5.62 $Y=1.885
+ $X2=5.62 $Y2=1.667
r72 1 3 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=5.62 $Y=1.885
+ $X2=5.62 $Y2=2.46
.ends

.subckt PM_SKY130_FD_SC_HS__A211O_4%A2 2 3 5 6 7 11 12 14 15 16 18 22 24 26
c67 24 0 1.25287e-19 $X=5.04 $Y=0.555
c68 22 0 3.8172e-19 $X=6.535 $Y=0.935
r69 29 31 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.155 $Y=0.34
+ $X2=5.155 $Y2=0.505
r70 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.155
+ $Y=0.34 $X2=5.155 $Y2=0.34
r71 26 29 24.4806 $w=3.3e-07 $l=1.4e-07 $layer=POLY_cond $X=5.155 $Y=0.2
+ $X2=5.155 $Y2=0.34
r72 24 30 8.27445 $w=3.17e-07 $l=2.15e-07 $layer=LI1_cond $X=5.122 $Y=0.555
+ $X2=5.122 $Y2=0.34
r73 22 23 230.745 $w=1.5e-07 $l=4.5e-07 $layer=POLY_cond $X=6.535 $Y=0.935
+ $X2=6.535 $Y2=1.385
r74 19 22 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=6.535 $Y=0.275
+ $X2=6.535 $Y2=0.935
r75 16 18 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=6.52 $Y=1.885
+ $X2=6.52 $Y2=2.46
r76 15 16 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=6.52 $Y=1.795 $X2=6.52
+ $Y2=1.885
r77 14 23 37.1337 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=6.52 $Y=1.475 $X2=6.52
+ $Y2=1.385
r78 14 15 124.387 $w=1.8e-07 $l=3.2e-07 $layer=POLY_cond $X=6.52 $Y=1.475
+ $X2=6.52 $Y2=1.795
r79 13 26 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.32 $Y=0.2
+ $X2=5.155 $Y2=0.2
r80 12 19 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=6.46 $Y=0.2
+ $X2=6.535 $Y2=0.275
r81 12 13 584.553 $w=1.5e-07 $l=1.14e-06 $layer=POLY_cond $X=6.46 $Y=0.2
+ $X2=5.32 $Y2=0.2
r82 11 31 220.489 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=5.245 $Y=0.935
+ $X2=5.245 $Y2=0.505
r83 9 11 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=5.245 $Y=1.33
+ $X2=5.245 $Y2=0.935
r84 6 9 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.17 $Y=1.405
+ $X2=5.245 $Y2=1.33
r85 6 7 135.883 $w=1.5e-07 $l=2.65e-07 $layer=POLY_cond $X=5.17 $Y=1.405
+ $X2=4.905 $Y2=1.405
r86 3 5 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=4.815 $Y=1.885
+ $X2=4.815 $Y2=2.46
r87 2 3 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=4.815 $Y=1.795 $X2=4.815
+ $Y2=1.885
r88 1 7 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=4.815 $Y=1.48
+ $X2=4.905 $Y2=1.405
r89 1 2 122.444 $w=1.8e-07 $l=3.15e-07 $layer=POLY_cond $X=4.815 $Y=1.48
+ $X2=4.815 $Y2=1.795
.ends

.subckt PM_SKY130_FD_SC_HS__A211O_4%VPWR 1 2 3 4 5 16 18 22 26 28 32 38 42 45 46
+ 47 49 62 63 69 72 75
r93 75 76 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r94 72 73 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r95 70 73 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.16 $Y2=3.33
r96 69 70 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r97 67 70 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=1.2 $Y2=3.33
r98 66 67 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r99 62 63 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r100 60 63 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6 $Y=3.33 $X2=6.96
+ $Y2=3.33
r101 60 76 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6 $Y=3.33 $X2=5.04
+ $Y2=3.33
r102 59 60 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r103 57 75 13.399 $w=1.7e-07 $l=3.38e-07 $layer=LI1_cond $X=5.555 $Y=3.33
+ $X2=5.217 $Y2=3.33
r104 57 59 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=5.555 $Y=3.33
+ $X2=6 $Y2=3.33
r105 56 76 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=5.04 $Y2=3.33
r106 55 56 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r107 53 73 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=2.16 $Y2=3.33
r108 52 55 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=2.64 $Y=3.33
+ $X2=4.56 $Y2=3.33
r109 52 53 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r110 50 72 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.275 $Y=3.33
+ $X2=2.19 $Y2=3.33
r111 50 52 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=2.275 $Y=3.33
+ $X2=2.64 $Y2=3.33
r112 49 75 13.399 $w=1.7e-07 $l=3.37e-07 $layer=LI1_cond $X=4.88 $Y=3.33
+ $X2=5.217 $Y2=3.33
r113 49 55 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=4.88 $Y=3.33
+ $X2=4.56 $Y2=3.33
r114 47 56 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.56 $Y2=3.33
r115 47 53 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=2.64 $Y2=3.33
r116 45 59 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=6.13 $Y=3.33 $X2=6
+ $Y2=3.33
r117 45 46 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.13 $Y=3.33
+ $X2=6.295 $Y2=3.33
r118 44 62 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=6.46 $Y=3.33 $X2=6.96
+ $Y2=3.33
r119 44 46 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.46 $Y=3.33
+ $X2=6.295 $Y2=3.33
r120 40 46 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.295 $Y=3.245
+ $X2=6.295 $Y2=3.33
r121 40 42 30.3826 $w=3.28e-07 $l=8.7e-07 $layer=LI1_cond $X=6.295 $Y=3.245
+ $X2=6.295 $Y2=2.375
r122 36 75 2.78459 $w=6.75e-07 $l=8.5e-08 $layer=LI1_cond $X=5.217 $Y=3.245
+ $X2=5.217 $Y2=3.33
r123 36 38 13.467 $w=6.73e-07 $l=7.6e-07 $layer=LI1_cond $X=5.217 $Y=3.245
+ $X2=5.217 $Y2=2.485
r124 32 35 54.1497 $w=1.68e-07 $l=8.3e-07 $layer=LI1_cond $X=2.19 $Y=1.985
+ $X2=2.19 $Y2=2.815
r125 30 72 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.19 $Y=3.245
+ $X2=2.19 $Y2=3.33
r126 30 35 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=2.19 $Y=3.245
+ $X2=2.19 $Y2=2.815
r127 29 69 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.375 $Y=3.33
+ $X2=1.25 $Y2=3.33
r128 28 72 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.105 $Y=3.33
+ $X2=2.19 $Y2=3.33
r129 28 29 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=2.105 $Y=3.33
+ $X2=1.375 $Y2=3.33
r130 24 69 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.25 $Y=3.245
+ $X2=1.25 $Y2=3.33
r131 24 26 47.0197 $w=2.48e-07 $l=1.02e-06 $layer=LI1_cond $X=1.25 $Y=3.245
+ $X2=1.25 $Y2=2.225
r132 23 66 3.89925 $w=1.7e-07 $l=2.38e-07 $layer=LI1_cond $X=0.475 $Y=3.33
+ $X2=0.237 $Y2=3.33
r133 22 69 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.125 $Y=3.33
+ $X2=1.25 $Y2=3.33
r134 22 23 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=1.125 $Y=3.33
+ $X2=0.475 $Y2=3.33
r135 18 21 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=0.35 $Y=1.985
+ $X2=0.35 $Y2=2.815
r136 16 66 3.24391 $w=2.5e-07 $l=1.49579e-07 $layer=LI1_cond $X=0.35 $Y=3.245
+ $X2=0.237 $Y2=3.33
r137 16 21 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=0.35 $Y=3.245
+ $X2=0.35 $Y2=2.815
r138 5 42 300 $w=1.7e-07 $l=4.84226e-07 $layer=licon1_PDIFF $count=2 $X=6.145
+ $Y=1.96 $X2=6.295 $Y2=2.375
r139 4 38 150 $w=1.7e-07 $l=7.3357e-07 $layer=licon1_PDIFF $count=4 $X=4.89
+ $Y=1.96 $X2=5.39 $Y2=2.485
r140 3 35 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=2.04
+ $Y=1.84 $X2=2.19 $Y2=2.815
r141 3 32 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=2.04
+ $Y=1.84 $X2=2.19 $Y2=1.985
r142 2 26 300 $w=1.7e-07 $l=4.53845e-07 $layer=licon1_PDIFF $count=2 $X=1.14
+ $Y=1.84 $X2=1.29 $Y2=2.225
r143 1 21 400 $w=1.7e-07 $l=1.03562e-06 $layer=licon1_PDIFF $count=1 $X=0.265
+ $Y=1.84 $X2=0.39 $Y2=2.815
r144 1 18 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.265
+ $Y=1.84 $X2=0.39 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HS__A211O_4%X 1 2 3 4 14 17 21 22 23 27 31 35 37 39 43
+ 44 50 52
r71 49 52 0.128611 $w=4.63e-07 $l=5e-09 $layer=LI1_cond $X=1.562 $Y=0.96
+ $X2=1.562 $Y2=0.965
r72 44 50 2.39545 $w=4.65e-07 $l=8.5e-08 $layer=LI1_cond $X=1.562 $Y=1.325
+ $X2=1.562 $Y2=1.24
r73 44 50 0.385832 $w=4.63e-07 $l=1.5e-08 $layer=LI1_cond $X=1.562 $Y=1.225
+ $X2=1.562 $Y2=1.24
r74 43 49 2.99104 $w=3.17e-07 $l=8.5e-08 $layer=LI1_cond $X=1.562 $Y=0.875
+ $X2=1.562 $Y2=0.96
r75 43 44 6.17331 $w=4.63e-07 $l=2.4e-07 $layer=LI1_cond $X=1.562 $Y=0.985
+ $X2=1.562 $Y2=1.225
r76 43 52 0.514442 $w=4.63e-07 $l=2e-08 $layer=LI1_cond $X=1.562 $Y=0.985
+ $X2=1.562 $Y2=0.965
r77 39 41 7.58852 $w=1.88e-07 $l=1.3e-07 $layer=LI1_cond $X=2.275 $Y=0.745
+ $X2=2.275 $Y2=0.875
r78 36 43 3.66292 $w=1.7e-07 $l=2.33e-07 $layer=LI1_cond $X=1.795 $Y=0.875
+ $X2=1.562 $Y2=0.875
r79 35 41 1.386 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=2.18 $Y=0.875 $X2=2.275
+ $Y2=0.875
r80 35 36 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=2.18 $Y=0.875
+ $X2=1.795 $Y2=0.875
r81 31 33 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=1.74 $Y=1.985
+ $X2=1.74 $Y2=2.815
r82 29 31 3.31764 $w=3.28e-07 $l=9.5e-08 $layer=LI1_cond $X=1.74 $Y=1.89
+ $X2=1.74 $Y2=1.985
r83 25 43 2.99104 $w=3.17e-07 $l=1.84673e-07 $layer=LI1_cond $X=1.415 $Y=0.79
+ $X2=1.562 $Y2=0.875
r84 25 27 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=1.415 $Y=0.79
+ $X2=1.415 $Y2=0.515
r85 24 37 2.76166 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.925 $Y=1.805
+ $X2=0.8 $Y2=1.805
r86 23 29 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.575 $Y=1.805
+ $X2=1.74 $Y2=1.89
r87 23 24 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=1.575 $Y=1.805
+ $X2=0.925 $Y2=1.805
r88 21 44 6.53816 $w=1.7e-07 $l=2.32e-07 $layer=LI1_cond $X=1.33 $Y=1.325
+ $X2=1.562 $Y2=1.325
r89 21 22 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=1.33 $Y=1.325
+ $X2=0.925 $Y2=1.325
r90 17 19 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=0.8 $Y=1.985 $X2=0.8
+ $Y2=2.815
r91 15 37 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.8 $Y=1.89 $X2=0.8
+ $Y2=1.805
r92 15 17 4.37928 $w=2.48e-07 $l=9.5e-08 $layer=LI1_cond $X=0.8 $Y=1.89 $X2=0.8
+ $Y2=1.985
r93 14 37 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.8 $Y=1.72 $X2=0.8
+ $Y2=1.805
r94 13 22 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.8 $Y=1.41
+ $X2=0.925 $Y2=1.325
r95 13 14 14.2903 $w=2.48e-07 $l=3.1e-07 $layer=LI1_cond $X=0.8 $Y=1.41 $X2=0.8
+ $Y2=1.72
r96 4 33 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=1.59
+ $Y=1.84 $X2=1.74 $Y2=2.815
r97 4 31 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=1.59
+ $Y=1.84 $X2=1.74 $Y2=1.985
r98 3 19 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=0.69
+ $Y=1.84 $X2=0.84 $Y2=2.815
r99 3 17 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=0.69
+ $Y=1.84 $X2=0.84 $Y2=1.985
r100 2 39 182 $w=1.7e-07 $l=4.3946e-07 $layer=licon1_NDIFF $count=1 $X=2.135
+ $Y=0.37 $X2=2.275 $Y2=0.745
r101 1 52 182 $w=1.7e-07 $l=6.61306e-07 $layer=licon1_NDIFF $count=1 $X=1.275
+ $Y=0.37 $X2=1.415 $Y2=0.965
r102 1 27 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=1.275
+ $Y=0.37 $X2=1.415 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__A211O_4%A_517_392# 1 2 3 4 13 15 16 19 21 25 27 29
+ 31 33 41 42
c71 42 0 2.37887e-20 $X=5.82 $Y=2.035
c72 29 0 4.75553e-20 $X=6.77 $Y=2.12
c73 27 0 6.73012e-21 $X=6.58 $Y=2.035
c74 25 0 3.06756e-19 $X=5.845 $Y=2.465
r75 46 47 3.8299 $w=2.78e-07 $l=8.5e-08 $layer=LI1_cond $X=5.82 $Y=2.145
+ $X2=5.82 $Y2=2.23
r76 45 46 1.23476 $w=2.78e-07 $l=3e-08 $layer=LI1_cond $X=5.82 $Y=2.115 $X2=5.82
+ $Y2=2.145
r77 42 45 3.29269 $w=2.78e-07 $l=8e-08 $layer=LI1_cond $X=5.82 $Y=2.035 $X2=5.82
+ $Y2=2.115
r78 33 36 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=2.71 $Y=2.485 $X2=2.71
+ $Y2=2.565
r79 29 49 2.96985 $w=2.8e-07 $l=1.01735e-07 $layer=LI1_cond $X=6.77 $Y=2.12
+ $X2=6.745 $Y2=2.03
r80 29 31 28.6053 $w=2.78e-07 $l=6.95e-07 $layer=LI1_cond $X=6.77 $Y=2.12
+ $X2=6.77 $Y2=2.815
r81 28 42 3.65648 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=5.96 $Y=2.035
+ $X2=5.82 $Y2=2.035
r82 27 49 4.39021 $w=1.7e-07 $l=1.67481e-07 $layer=LI1_cond $X=6.58 $Y=2.035
+ $X2=6.745 $Y2=2.03
r83 27 28 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=6.58 $Y=2.035
+ $X2=5.96 $Y2=2.035
r84 25 47 11.5244 $w=2.33e-07 $l=2.35e-07 $layer=LI1_cond $X=5.842 $Y=2.465
+ $X2=5.842 $Y2=2.23
r85 22 39 4.68908 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=4.71 $Y=2.145
+ $X2=4.565 $Y2=2.145
r86 21 46 3.65648 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=5.68 $Y=2.145
+ $X2=5.82 $Y2=2.145
r87 21 22 63.2834 $w=1.68e-07 $l=9.7e-07 $layer=LI1_cond $X=5.68 $Y=2.145
+ $X2=4.71 $Y2=2.145
r88 17 41 3.70735 $w=2.5e-07 $l=1.03078e-07 $layer=LI1_cond $X=4.605 $Y=2.57
+ $X2=4.565 $Y2=2.485
r89 17 19 13.4675 $w=2.08e-07 $l=2.55e-07 $layer=LI1_cond $X=4.605 $Y=2.57
+ $X2=4.605 $Y2=2.825
r90 16 41 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.565 $Y=2.4
+ $X2=4.565 $Y2=2.485
r91 15 39 2.74877 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=4.565 $Y=2.23
+ $X2=4.565 $Y2=2.145
r92 15 16 6.7557 $w=2.88e-07 $l=1.7e-07 $layer=LI1_cond $X=4.565 $Y=2.23
+ $X2=4.565 $Y2=2.4
r93 14 33 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.875 $Y=2.485
+ $X2=2.71 $Y2=2.485
r94 13 41 2.76166 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=4.42 $Y=2.485
+ $X2=4.565 $Y2=2.485
r95 13 14 100.797 $w=1.68e-07 $l=1.545e-06 $layer=LI1_cond $X=4.42 $Y=2.485
+ $X2=2.875 $Y2=2.485
r96 4 49 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=6.595
+ $Y=1.96 $X2=6.745 $Y2=2.105
r97 4 31 400 $w=1.7e-07 $l=9.26971e-07 $layer=licon1_PDIFF $count=1 $X=6.595
+ $Y=1.96 $X2=6.745 $Y2=2.815
r98 3 45 600 $w=1.7e-07 $l=2.17428e-07 $layer=licon1_PDIFF $count=1 $X=5.695
+ $Y=1.96 $X2=5.845 $Y2=2.115
r99 3 25 300 $w=1.7e-07 $l=5.7513e-07 $layer=licon1_PDIFF $count=2 $X=5.695
+ $Y=1.96 $X2=5.845 $Y2=2.465
r100 2 41 600 $w=1.7e-07 $l=5.95294e-07 $layer=licon1_PDIFF $count=1 $X=4.435
+ $Y=1.96 $X2=4.585 $Y2=2.485
r101 2 39 600 $w=1.7e-07 $l=2.48948e-07 $layer=licon1_PDIFF $count=1 $X=4.435
+ $Y=1.96 $X2=4.585 $Y2=2.145
r102 2 19 600 $w=1.7e-07 $l=9.37003e-07 $layer=licon1_PDIFF $count=1 $X=4.435
+ $Y=1.96 $X2=4.585 $Y2=2.825
r103 1 36 600 $w=1.7e-07 $l=6.64568e-07 $layer=licon1_PDIFF $count=1 $X=2.585
+ $Y=1.96 $X2=2.71 $Y2=2.565
.ends

.subckt PM_SKY130_FD_SC_HS__A211O_4%A_602_392# 1 2 11
r14 8 11 41.9489 $w=2.48e-07 $l=9.1e-07 $layer=LI1_cond $X=3.21 $Y=2.865
+ $X2=4.12 $Y2=2.865
r15 2 11 600 $w=1.7e-07 $l=9.41608e-07 $layer=licon1_PDIFF $count=1 $X=3.96
+ $Y=1.96 $X2=4.12 $Y2=2.825
r16 1 8 600 $w=1.7e-07 $l=9.59805e-07 $layer=licon1_PDIFF $count=1 $X=3.01
+ $Y=1.96 $X2=3.21 $Y2=2.825
.ends

.subckt PM_SKY130_FD_SC_HS__A211O_4%VGND 1 2 3 4 5 6 21 23 27 31 37 41 45 47 48
+ 49 50 51 52 58 63 68 82 84 87 90 93
r101 93 94 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r102 87 88 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r103 84 85 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r104 81 82 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=0 $X2=6.96
+ $Y2=0
r105 79 82 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=0 $X2=6.96
+ $Y2=0
r106 78 79 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.48 $Y=0 $X2=6.48
+ $Y2=0
r107 76 79 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=5.04 $Y=0
+ $X2=6.48 $Y2=0
r108 76 94 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=4.56
+ $Y2=0
r109 75 78 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=5.04 $Y=0 $X2=6.48
+ $Y2=0
r110 75 76 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r111 73 93 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.755 $Y=0 $X2=4.59
+ $Y2=0
r112 73 75 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=4.755 $Y=0
+ $X2=5.04 $Y2=0
r113 72 94 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=4.56
+ $Y2=0
r114 71 72 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r115 69 90 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.79 $Y=0 $X2=3.625
+ $Y2=0
r116 69 71 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=3.79 $Y=0 $X2=4.08
+ $Y2=0
r117 68 93 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.425 $Y=0 $X2=4.59
+ $Y2=0
r118 68 71 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=4.425 $Y=0 $X2=4.08
+ $Y2=0
r119 67 88 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=2.64
+ $Y2=0
r120 66 67 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r121 64 87 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.87 $Y=0 $X2=2.705
+ $Y2=0
r122 64 66 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=2.87 $Y=0 $X2=3.12
+ $Y2=0
r123 63 90 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.46 $Y=0 $X2=3.625
+ $Y2=0
r124 63 66 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=3.46 $Y=0 $X2=3.12
+ $Y2=0
r125 62 88 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r126 62 85 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.68
+ $Y2=0
r127 61 62 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r128 59 84 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.01 $Y=0 $X2=1.845
+ $Y2=0
r129 59 61 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=2.01 $Y=0 $X2=2.16
+ $Y2=0
r130 58 87 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.54 $Y=0 $X2=2.705
+ $Y2=0
r131 58 61 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=2.54 $Y=0 $X2=2.16
+ $Y2=0
r132 56 85 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r133 55 56 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r134 52 72 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.08
+ $Y2=0
r135 52 67 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=3.12
+ $Y2=0
r136 52 90 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r137 50 78 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=6.585 $Y=0
+ $X2=6.48 $Y2=0
r138 50 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.585 $Y=0 $X2=6.75
+ $Y2=0
r139 49 81 3.22941 $w=1.7e-07 $l=4.5e-08 $layer=LI1_cond $X=6.915 $Y=0 $X2=6.96
+ $Y2=0
r140 49 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.915 $Y=0 $X2=6.75
+ $Y2=0
r141 47 55 6.52406 $w=1.68e-07 $l=1e-07 $layer=LI1_cond $X=0.82 $Y=0 $X2=0.72
+ $Y2=0
r142 47 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.82 $Y=0 $X2=0.985
+ $Y2=0
r143 43 51 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.75 $Y=0.085
+ $X2=6.75 $Y2=0
r144 43 45 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=6.75 $Y=0.085
+ $X2=6.75 $Y2=0.76
r145 39 93 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.59 $Y=0.085
+ $X2=4.59 $Y2=0
r146 39 41 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=4.59 $Y=0.085
+ $X2=4.59 $Y2=0.765
r147 35 90 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.625 $Y=0.085
+ $X2=3.625 $Y2=0
r148 35 37 18.5089 $w=3.28e-07 $l=5.3e-07 $layer=LI1_cond $X=3.625 $Y=0.085
+ $X2=3.625 $Y2=0.615
r149 31 33 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=2.705 $Y=0.515
+ $X2=2.705 $Y2=0.855
r150 29 87 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.705 $Y=0.085
+ $X2=2.705 $Y2=0
r151 29 31 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=2.705 $Y=0.085
+ $X2=2.705 $Y2=0.515
r152 25 84 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.845 $Y=0.085
+ $X2=1.845 $Y2=0
r153 25 27 15.3659 $w=3.28e-07 $l=4.4e-07 $layer=LI1_cond $X=1.845 $Y=0.085
+ $X2=1.845 $Y2=0.525
r154 24 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.15 $Y=0 $X2=0.985
+ $Y2=0
r155 23 84 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.68 $Y=0 $X2=1.845
+ $Y2=0
r156 23 24 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=1.68 $Y=0 $X2=1.15
+ $Y2=0
r157 19 48 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.985 $Y=0.085
+ $X2=0.985 $Y2=0
r158 19 21 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=0.985 $Y=0.085
+ $X2=0.985 $Y2=0.515
r159 6 45 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=6.61
+ $Y=0.615 $X2=6.75 $Y2=0.76
r160 5 41 182 $w=1.7e-07 $l=2.08567e-07 $layer=licon1_NDIFF $count=1 $X=4.45
+ $Y=0.615 $X2=4.59 $Y2=0.765
r161 4 37 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=3.485
+ $Y=0.47 $X2=3.625 $Y2=0.615
r162 3 33 182 $w=1.7e-07 $l=5.50568e-07 $layer=licon1_NDIFF $count=1 $X=2.565
+ $Y=0.37 $X2=2.705 $Y2=0.855
r163 3 31 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=2.565
+ $Y=0.37 $X2=2.705 $Y2=0.515
r164 2 27 182 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_NDIFF $count=1 $X=1.705
+ $Y=0.37 $X2=1.845 $Y2=0.525
r165 1 21 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.86
+ $Y=0.37 $X2=0.985 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__A211O_4%A_1064_123# 1 2 7 11 13
c23 13 0 2.7959e-19 $X=6.32 $Y=1.11
c24 11 0 1.39955e-19 $X=6.32 $Y=0.845
r25 11 16 3.40825 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.32 $Y=0.845
+ $X2=6.32 $Y2=0.72
r26 11 13 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=6.32 $Y=0.845
+ $X2=6.32 $Y2=1.11
r27 7 16 3.40825 $w=1.7e-07 $l=1.03078e-07 $layer=LI1_cond $X=6.235 $Y=0.76
+ $X2=6.32 $Y2=0.72
r28 7 9 50.5615 $w=1.68e-07 $l=7.75e-07 $layer=LI1_cond $X=6.235 $Y=0.76
+ $X2=5.46 $Y2=0.76
r29 2 16 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=6.18
+ $Y=0.615 $X2=6.32 $Y2=0.76
r30 2 13 182 $w=1.7e-07 $l=5.60647e-07 $layer=licon1_NDIFF $count=1 $X=6.18
+ $Y=0.615 $X2=6.32 $Y2=1.11
r31 1 9 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=5.32
+ $Y=0.615 $X2=5.46 $Y2=0.76
.ends

