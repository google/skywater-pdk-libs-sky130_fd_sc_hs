* File: sky130_fd_sc_hs__nand2b_4.pex.spice
* Created: Thu Aug 27 20:50:47 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HS__NAND2B_4%A_N 3 5 7 8 10 12 13 14 15 16 19 22
c53 8 0 7.22234e-20 $X=1.53 $Y=1.65
r54 24 25 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=0.27
+ $Y=1.465 $X2=0.27 $Y2=1.465
r55 21 22 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=0.95
+ $Y=1.465 $X2=0.95 $Y2=1.465
r56 19 21 47.1095 $w=4.25e-07 $l=3.6e-07 $layer=POLY_cond $X=0.59 $Y=1.512
+ $X2=0.95 $Y2=1.512
r57 16 22 5.73121 $w=4.78e-07 $l=2.3e-07 $layer=LI1_cond $X=0.72 $Y=1.54
+ $X2=0.95 $Y2=1.54
r58 16 25 11.2132 $w=4.78e-07 $l=4.5e-07 $layer=LI1_cond $X=0.72 $Y=1.54
+ $X2=0.27 $Y2=1.54
r59 15 25 0.747549 $w=4.78e-07 $l=3e-08 $layer=LI1_cond $X=0.24 $Y=1.54 $X2=0.27
+ $Y2=1.54
r60 13 21 17.0118 $w=4.25e-07 $l=1.3e-07 $layer=POLY_cond $X=1.08 $Y=1.512
+ $X2=0.95 $Y2=1.512
r61 13 14 11.5413 $w=2.87e-07 $l=9.94987e-08 $layer=POLY_cond $X=1.08 $Y=1.512
+ $X2=1.17 $Y2=1.532
r62 10 12 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=1.62 $Y=1.765
+ $X2=1.62 $Y2=2.26
r63 9 14 11.5413 $w=2.87e-07 $l=1.56665e-07 $layer=POLY_cond $X=1.26 $Y=1.65
+ $X2=1.17 $Y2=1.532
r64 8 10 26.9307 $w=1.5e-07 $l=1.53542e-07 $layer=POLY_cond $X=1.53 $Y=1.65
+ $X2=1.62 $Y2=1.765
r65 8 9 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=1.53 $Y=1.65 $X2=1.26
+ $Y2=1.65
r66 5 14 14.8601 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=1.17 $Y=1.765
+ $X2=1.17 $Y2=1.532
r67 5 7 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=1.17 $Y=1.765 $X2=1.17
+ $Y2=2.26
r68 1 19 9.81448 $w=4.25e-07 $l=7.5e-08 $layer=POLY_cond $X=0.515 $Y=1.512
+ $X2=0.59 $Y2=1.512
r69 1 24 32.0606 $w=4.25e-07 $l=2.45e-07 $layer=POLY_cond $X=0.515 $Y=1.512
+ $X2=0.27 $Y2=1.512
r70 1 3 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=0.515 $Y=1.3 $X2=0.515
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HS__NAND2B_4%A_31_74# 1 2 7 9 10 11 12 14 15 17 18 20 21
+ 23 24 26 29 31 32 35 38 46 49 50 56
r117 56 57 1.50312 $w=4.81e-07 $l=1.5e-08 $layer=POLY_cond $X=2.985 $Y=1.475
+ $X2=3 $Y2=1.475
r118 47 56 7.51559 $w=4.81e-07 $l=7.5e-08 $layer=POLY_cond $X=2.91 $Y=1.475
+ $X2=2.985 $Y2=1.475
r119 47 54 47.5988 $w=4.81e-07 $l=4.75e-07 $layer=POLY_cond $X=2.91 $Y=1.475
+ $X2=2.435 $Y2=1.475
r120 46 47 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=2.91
+ $Y=1.515 $X2=2.91 $Y2=1.515
r121 44 54 20.5426 $w=4.81e-07 $l=2.05e-07 $layer=POLY_cond $X=2.23 $Y=1.475
+ $X2=2.435 $Y2=1.475
r122 44 52 7.51559 $w=4.81e-07 $l=7.5e-08 $layer=POLY_cond $X=2.23 $Y=1.475
+ $X2=2.155 $Y2=1.475
r123 43 46 31.3464 $w=2.48e-07 $l=6.8e-07 $layer=LI1_cond $X=2.23 $Y=1.555
+ $X2=2.91 $Y2=1.555
r124 43 44 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=2.23
+ $Y=1.515 $X2=2.23 $Y2=1.515
r125 41 50 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.455 $Y=1.555
+ $X2=1.37 $Y2=1.555
r126 41 43 35.7257 $w=2.48e-07 $l=7.75e-07 $layer=LI1_cond $X=1.455 $Y=1.555
+ $X2=2.23 $Y2=1.555
r127 39 50 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.37 $Y=1.68
+ $X2=1.37 $Y2=1.555
r128 39 49 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=1.37 $Y=1.68
+ $X2=1.37 $Y2=1.95
r129 38 50 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.37 $Y=1.43
+ $X2=1.37 $Y2=1.555
r130 37 38 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=1.37 $Y=1.13 $X2=1.37
+ $Y2=1.43
r131 35 49 7.36219 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=1.395 $Y=2.115
+ $X2=1.395 $Y2=1.95
r132 31 37 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.285 $Y=1.045
+ $X2=1.37 $Y2=1.13
r133 31 32 58.7166 $w=1.68e-07 $l=9e-07 $layer=LI1_cond $X=1.285 $Y=1.045
+ $X2=0.385 $Y2=1.045
r134 27 32 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.26 $Y=0.96
+ $X2=0.385 $Y2=1.045
r135 27 29 20.5135 $w=2.48e-07 $l=4.45e-07 $layer=LI1_cond $X=0.26 $Y=0.96
+ $X2=0.26 $Y2=0.515
r136 24 57 30.4321 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=3 $Y=1.185 $X2=3
+ $Y2=1.475
r137 24 26 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=3 $Y=1.185 $X2=3
+ $Y2=0.74
r138 21 56 30.4321 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=2.985 $Y=1.765
+ $X2=2.985 $Y2=1.475
r139 21 23 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.985 $Y=1.765
+ $X2=2.985 $Y2=2.4
r140 18 54 30.4321 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=2.435 $Y=1.185
+ $X2=2.435 $Y2=1.475
r141 18 20 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=2.435 $Y=1.185
+ $X2=2.435 $Y2=0.74
r142 15 52 30.4321 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=2.155 $Y=1.765
+ $X2=2.155 $Y2=1.475
r143 15 17 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.155 $Y=1.765
+ $X2=2.155 $Y2=2.4
r144 12 52 15.0312 $w=4.81e-07 $l=3.57211e-07 $layer=POLY_cond $X=2.005 $Y=1.185
+ $X2=2.155 $Y2=1.475
r145 12 14 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=2.005 $Y=1.185
+ $X2=2.005 $Y2=0.74
r146 10 12 32.422 $w=4.81e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.93 $Y=1.26
+ $X2=2.005 $Y2=1.185
r147 10 11 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=1.93 $Y=1.26
+ $X2=1.65 $Y2=1.26
r148 7 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.575 $Y=1.185
+ $X2=1.65 $Y2=1.26
r149 7 9 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=1.575 $Y=1.185
+ $X2=1.575 $Y2=0.74
r150 2 35 300 $w=1.7e-07 $l=3.4187e-07 $layer=licon1_PDIFF $count=2 $X=1.245
+ $Y=1.84 $X2=1.395 $Y2=2.115
r151 1 29 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.155
+ $Y=0.37 $X2=0.3 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__NAND2B_4%B 3 5 6 9 13 15 17 18 20 23 30 31 32 44 48
+ 56
c80 15 0 1.73061e-19 $X=4.735 $Y=1.765
c81 9 0 1.04617e-19 $X=3.93 $Y=0.74
r82 46 47 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.37
+ $Y=1.465 $X2=5.37 $Y2=1.465
r83 44 46 14.1369 $w=3.58e-07 $l=1.05e-07 $layer=POLY_cond $X=5.265 $Y=1.532
+ $X2=5.37 $Y2=1.532
r84 43 44 8.07821 $w=3.58e-07 $l=6e-08 $layer=POLY_cond $X=5.205 $Y=1.532
+ $X2=5.265 $Y2=1.532
r85 42 43 63.2793 $w=3.58e-07 $l=4.7e-07 $layer=POLY_cond $X=4.735 $Y=1.532
+ $X2=5.205 $Y2=1.532
r86 41 48 5.8558 $w=4.78e-07 $l=2.35e-07 $layer=LI1_cond $X=4.69 $Y=1.54
+ $X2=4.925 $Y2=1.54
r87 40 42 6.05866 $w=3.58e-07 $l=4.5e-08 $layer=POLY_cond $X=4.69 $Y=1.532
+ $X2=4.735 $Y2=1.532
r88 40 41 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=4.69
+ $Y=1.465 $X2=4.69 $Y2=1.465
r89 38 40 44.4302 $w=3.58e-07 $l=3.3e-07 $layer=POLY_cond $X=4.36 $Y=1.532
+ $X2=4.69 $Y2=1.532
r90 32 47 3.73775 $w=4.78e-07 $l=1.5e-07 $layer=LI1_cond $X=5.52 $Y=1.54
+ $X2=5.37 $Y2=1.54
r91 31 47 8.22304 $w=4.78e-07 $l=3.3e-07 $layer=LI1_cond $X=5.04 $Y=1.54
+ $X2=5.37 $Y2=1.54
r92 31 48 2.8656 $w=4.78e-07 $l=1.15e-07 $layer=LI1_cond $X=5.04 $Y=1.54
+ $X2=4.925 $Y2=1.54
r93 30 41 3.23938 $w=4.78e-07 $l=1.3e-07 $layer=LI1_cond $X=4.56 $Y=1.54
+ $X2=4.69 $Y2=1.54
r94 30 56 4.04332 $w=4.78e-07 $l=1.15e-07 $layer=LI1_cond $X=4.56 $Y=1.54
+ $X2=4.445 $Y2=1.54
r95 28 38 47.1229 $w=3.58e-07 $l=3.5e-07 $layer=POLY_cond $X=4.01 $Y=1.532
+ $X2=4.36 $Y2=1.532
r96 28 36 10.7709 $w=3.58e-07 $l=8e-08 $layer=POLY_cond $X=4.01 $Y=1.532
+ $X2=3.93 $Y2=1.532
r97 27 56 15.1913 $w=3.28e-07 $l=4.35e-07 $layer=LI1_cond $X=4.01 $Y=1.465
+ $X2=4.445 $Y2=1.465
r98 27 28 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=4.01
+ $Y=1.465 $X2=4.01 $Y2=1.465
r99 21 44 23.1716 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=5.265 $Y=1.3
+ $X2=5.265 $Y2=1.532
r100 21 23 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=5.265 $Y=1.3
+ $X2=5.265 $Y2=0.74
r101 18 43 23.1716 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=5.205 $Y=1.765
+ $X2=5.205 $Y2=1.532
r102 18 20 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=5.205 $Y=1.765
+ $X2=5.205 $Y2=2.4
r103 15 42 23.1716 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=4.735 $Y=1.765
+ $X2=4.735 $Y2=1.532
r104 15 17 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=4.735 $Y=1.765
+ $X2=4.735 $Y2=2.4
r105 11 38 23.1716 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=4.36 $Y=1.3
+ $X2=4.36 $Y2=1.532
r106 11 13 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=4.36 $Y=1.3
+ $X2=4.36 $Y2=0.74
r107 7 36 23.1716 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=3.93 $Y=1.3
+ $X2=3.93 $Y2=1.532
r108 7 9 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=3.93 $Y=1.3 $X2=3.93
+ $Y2=0.74
r109 5 36 10.4746 $w=3.58e-07 $l=1.03199e-07 $layer=POLY_cond $X=3.855 $Y=1.465
+ $X2=3.93 $Y2=1.532
r110 5 6 61.2015 $w=3.3e-07 $l=3.5e-07 $layer=POLY_cond $X=3.855 $Y=1.465
+ $X2=3.505 $Y2=1.465
r111 1 6 32.1775 $w=3.3e-07 $l=1.98997e-07 $layer=POLY_cond $X=3.43 $Y=1.3
+ $X2=3.505 $Y2=1.465
r112 1 3 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=3.43 $Y=1.3 $X2=3.43
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HS__NAND2B_4%VPWR 1 2 3 4 15 19 23 25 30 31 32 34 47 53
+ 58 69 72
r60 71 72 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r61 67 69 12.4766 $w=1.093e-06 $l=8.5e-08 $layer=LI1_cond $X=4.56 $Y=2.867
+ $X2=4.645 $Y2=2.867
r62 67 68 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r63 65 67 0.891324 $w=1.093e-06 $l=8e-08 $layer=LI1_cond $X=4.48 $Y=2.867
+ $X2=4.56 $Y2=2.867
r64 63 68 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.56 $Y2=3.33
r65 62 65 9.80457 $w=1.093e-06 $l=8.8e-07 $layer=LI1_cond $X=3.6 $Y=2.867
+ $X2=4.48 $Y2=2.867
r66 62 63 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r67 60 62 4.34521 $w=1.093e-06 $l=3.9e-07 $layer=LI1_cond $X=3.21 $Y=2.867
+ $X2=3.6 $Y2=2.867
r68 57 63 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=3.6 $Y2=3.33
r69 56 60 1.00274 $w=1.093e-06 $l=9e-08 $layer=LI1_cond $X=3.12 $Y=2.867
+ $X2=3.21 $Y2=2.867
r70 56 58 12.3651 $w=1.093e-06 $l=7.5e-08 $layer=LI1_cond $X=3.12 $Y=2.867
+ $X2=3.045 $Y2=2.867
r71 56 57 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r72 53 54 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r73 51 72 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=5.52 $Y2=3.33
r74 51 68 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=4.56 $Y2=3.33
r75 50 69 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=5.04 $Y=3.33
+ $X2=4.645 $Y2=3.33
r76 50 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r77 47 71 4.2442 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=5.315 $Y=3.33
+ $X2=5.537 $Y2=3.33
r78 47 50 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=5.315 $Y=3.33
+ $X2=5.04 $Y2=3.33
r79 45 58 57.738 $w=1.68e-07 $l=8.85e-07 $layer=LI1_cond $X=2.16 $Y=3.33
+ $X2=3.045 $Y2=3.33
r80 45 46 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r81 42 46 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r82 42 54 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=0.72 $Y2=3.33
r83 41 42 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r84 39 53 12.8484 $w=1.7e-07 $l=3.13e-07 $layer=LI1_cond $X=1.06 $Y=3.33
+ $X2=0.747 $Y2=3.33
r85 39 41 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=1.06 $Y=3.33
+ $X2=1.68 $Y2=3.33
r86 37 54 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r87 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r88 34 53 12.8484 $w=1.7e-07 $l=3.12e-07 $layer=LI1_cond $X=0.435 $Y=3.33
+ $X2=0.747 $Y2=3.33
r89 34 36 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=0.435 $Y=3.33
+ $X2=0.24 $Y2=3.33
r90 32 57 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.88 $Y=3.33
+ $X2=3.12 $Y2=3.33
r91 32 46 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=2.88 $Y=3.33
+ $X2=2.16 $Y2=3.33
r92 30 41 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=1.765 $Y=3.33
+ $X2=1.68 $Y2=3.33
r93 30 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.765 $Y=3.33
+ $X2=1.93 $Y2=3.33
r94 29 45 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=2.095 $Y=3.33
+ $X2=2.16 $Y2=3.33
r95 29 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.095 $Y=3.33
+ $X2=1.93 $Y2=3.33
r96 25 28 28.3056 $w=2.83e-07 $l=7e-07 $layer=LI1_cond $X=5.457 $Y=2.115
+ $X2=5.457 $Y2=2.815
r97 23 71 3.15447 $w=2.85e-07 $l=1.18427e-07 $layer=LI1_cond $X=5.457 $Y=3.245
+ $X2=5.537 $Y2=3.33
r98 23 28 17.3877 $w=2.83e-07 $l=4.3e-07 $layer=LI1_cond $X=5.457 $Y=3.245
+ $X2=5.457 $Y2=2.815
r99 19 22 27.938 $w=3.28e-07 $l=8e-07 $layer=LI1_cond $X=1.93 $Y=2.015 $X2=1.93
+ $Y2=2.815
r100 17 31 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.93 $Y=3.245
+ $X2=1.93 $Y2=3.33
r101 17 22 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=1.93 $Y=3.245
+ $X2=1.93 $Y2=2.815
r102 13 53 2.61429 $w=6.25e-07 $l=8.5e-08 $layer=LI1_cond $X=0.747 $Y=3.245
+ $X2=0.747 $Y2=3.33
r103 13 15 21.6251 $w=6.23e-07 $l=1.13e-06 $layer=LI1_cond $X=0.747 $Y=3.245
+ $X2=0.747 $Y2=2.115
r104 4 28 400 $w=1.7e-07 $l=1.04964e-06 $layer=licon1_PDIFF $count=1 $X=5.28
+ $Y=1.84 $X2=5.435 $Y2=2.815
r105 4 25 400 $w=1.7e-07 $l=3.43875e-07 $layer=licon1_PDIFF $count=1 $X=5.28
+ $Y=1.84 $X2=5.435 $Y2=2.115
r106 3 65 150 $w=1.7e-07 $l=1.6789e-06 $layer=licon1_PDIFF $count=4 $X=3.06
+ $Y=1.84 $X2=4.48 $Y2=2.405
r107 3 60 150 $w=1.7e-07 $l=6.3559e-07 $layer=licon1_PDIFF $count=4 $X=3.06
+ $Y=1.84 $X2=3.21 $Y2=2.405
r108 2 22 600 $w=1.7e-07 $l=1.08616e-06 $layer=licon1_PDIFF $count=1 $X=1.695
+ $Y=1.84 $X2=1.93 $Y2=2.815
r109 2 19 300 $w=1.7e-07 $l=3.10403e-07 $layer=licon1_PDIFF $count=2 $X=1.695
+ $Y=1.84 $X2=1.93 $Y2=2.015
r110 1 15 150 $w=1.7e-07 $l=6.07124e-07 $layer=licon1_PDIFF $count=4 $X=0.455
+ $Y=1.84 $X2=0.94 $Y2=2.115
.ends

.subckt PM_SKY130_FD_SC_HS__NAND2B_4%Y 1 2 3 4 15 17 18 19 21 25 27 29 32 33 35
+ 37 41 44 45 50 57 59
c81 37 0 1.73061e-19 $X=4.98 $Y=2.815
c82 18 0 7.22234e-20 $X=1.885 $Y=1.175
r83 50 57 1.34452 $w=2.98e-07 $l=3.5e-08 $layer=LI1_cond $X=4.045 $Y=2 $X2=4.08
+ $Y2=2
r84 45 59 4.74082 $w=2.98e-07 $l=9e-08 $layer=LI1_cond $X=4.105 $Y=2 $X2=4.195
+ $Y2=2
r85 45 57 0.960369 $w=2.98e-07 $l=2.5e-08 $layer=LI1_cond $X=4.105 $Y=2 $X2=4.08
+ $Y2=2
r86 45 50 0.960369 $w=2.98e-07 $l=2.5e-08 $layer=LI1_cond $X=4.02 $Y=2 $X2=4.045
+ $Y2=2
r87 44 51 6.12828 $w=3e-07 $l=1.85e-07 $layer=LI1_cond $X=3.47 $Y=2 $X2=3.655
+ $Y2=2
r88 44 45 13.4452 $w=2.98e-07 $l=3.5e-07 $layer=LI1_cond $X=3.67 $Y=2 $X2=4.02
+ $Y2=2
r89 44 51 0.576222 $w=2.98e-07 $l=1.5e-08 $layer=LI1_cond $X=3.67 $Y=2 $X2=3.655
+ $Y2=2
r90 35 43 2.77883 $w=3.3e-07 $l=1e-07 $layer=LI1_cond $X=4.98 $Y=2.15 $X2=4.98
+ $Y2=2.05
r91 35 37 23.2235 $w=3.28e-07 $l=6.65e-07 $layer=LI1_cond $X=4.98 $Y=2.15
+ $X2=4.98 $Y2=2.815
r92 33 43 4.58506 $w=2e-07 $l=1.65e-07 $layer=LI1_cond $X=4.815 $Y=2.05 $X2=4.98
+ $Y2=2.05
r93 33 59 34.3818 $w=1.98e-07 $l=6.2e-07 $layer=LI1_cond $X=4.815 $Y=2.05
+ $X2=4.195 $Y2=2.05
r94 32 44 0.599429 $w=3.7e-07 $l=1.5e-07 $layer=LI1_cond $X=3.47 $Y=1.85
+ $X2=3.47 $Y2=2
r95 31 32 18.3768 $w=3.68e-07 $l=5.9e-07 $layer=LI1_cond $X=3.47 $Y=1.26
+ $X2=3.47 $Y2=1.85
r96 30 41 8.5188 $w=1.7e-07 $l=1.63e-07 $layer=LI1_cond $X=2.88 $Y=1.175
+ $X2=2.717 $Y2=1.175
r97 29 31 8.10976 $w=1.7e-07 $l=2.23495e-07 $layer=LI1_cond $X=3.285 $Y=1.175
+ $X2=3.47 $Y2=1.26
r98 29 30 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=3.285 $Y=1.175
+ $X2=2.88 $Y2=1.175
r99 28 40 5.29536 $w=3e-07 $l=3.05e-07 $layer=LI1_cond $X=2.875 $Y=2 $X2=2.57
+ $Y2=2
r100 27 44 6.12828 $w=3e-07 $l=1.85e-07 $layer=LI1_cond $X=3.285 $Y=2 $X2=3.47
+ $Y2=2
r101 27 28 15.7501 $w=2.98e-07 $l=4.1e-07 $layer=LI1_cond $X=3.285 $Y=2
+ $X2=2.875 $Y2=2
r102 23 41 0.848899 $w=3.25e-07 $l=8.5e-08 $layer=LI1_cond $X=2.717 $Y=1.09
+ $X2=2.717 $Y2=1.175
r103 23 25 9.57414 $w=3.23e-07 $l=2.7e-07 $layer=LI1_cond $X=2.717 $Y=1.09
+ $X2=2.717 $Y2=0.82
r104 19 40 2.60428 $w=6.1e-07 $l=1.5e-07 $layer=LI1_cond $X=2.57 $Y=2.15
+ $X2=2.57 $Y2=2
r105 19 21 5.19608 $w=6.08e-07 $l=2.65e-07 $layer=LI1_cond $X=2.57 $Y=2.15
+ $X2=2.57 $Y2=2.415
r106 17 41 8.5188 $w=1.7e-07 $l=1.62e-07 $layer=LI1_cond $X=2.555 $Y=1.175
+ $X2=2.717 $Y2=1.175
r107 17 18 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.555 $Y=1.175
+ $X2=1.885 $Y2=1.175
r108 13 18 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=1.755 $Y=1.09
+ $X2=1.885 $Y2=1.175
r109 13 15 11.9677 $w=2.58e-07 $l=2.7e-07 $layer=LI1_cond $X=1.755 $Y=1.09
+ $X2=1.755 $Y2=0.82
r110 4 43 400 $w=1.7e-07 $l=3.49821e-07 $layer=licon1_PDIFF $count=1 $X=4.81
+ $Y=1.84 $X2=4.98 $Y2=2.115
r111 4 37 400 $w=1.7e-07 $l=1.05659e-06 $layer=licon1_PDIFF $count=1 $X=4.81
+ $Y=1.84 $X2=4.98 $Y2=2.815
r112 3 40 300 $w=1.7e-07 $l=6.11269e-07 $layer=licon1_PDIFF $count=2 $X=2.23
+ $Y=1.84 $X2=2.76 $Y2=2.015
r113 3 21 150 $w=1.7e-07 $l=7.97104e-07 $layer=licon1_PDIFF $count=4 $X=2.23
+ $Y=1.84 $X2=2.76 $Y2=2.415
r114 2 25 182 $w=1.7e-07 $l=5.47037e-07 $layer=licon1_NDIFF $count=1 $X=2.51
+ $Y=0.37 $X2=2.725 $Y2=0.82
r115 1 15 182 $w=1.7e-07 $l=5.15267e-07 $layer=licon1_NDIFF $count=1 $X=1.65
+ $Y=0.37 $X2=1.79 $Y2=0.82
.ends

.subckt PM_SKY130_FD_SC_HS__NAND2B_4%VGND 1 2 3 12 16 18 22 24 26 31 38 39 42 45
+ 48
r69 49 51 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=4.56
+ $Y2=0
r70 48 51 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r71 48 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r72 46 51 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.56
+ $Y2=0
r73 45 46 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r74 42 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r75 39 49 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=5.04
+ $Y2=0
r76 38 39 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r77 36 48 13.2917 $w=1.7e-07 $l=3.33e-07 $layer=LI1_cond $X=5.145 $Y=0 $X2=4.812
+ $Y2=0
r78 36 38 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=5.145 $Y=0 $X2=5.52
+ $Y2=0
r79 35 43 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r80 34 35 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r81 32 42 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.895 $Y=0 $X2=0.73
+ $Y2=0
r82 32 34 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.895 $Y=0 $X2=1.2
+ $Y2=0
r83 31 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.55 $Y=0 $X2=3.715
+ $Y2=0
r84 31 34 153.316 $w=1.68e-07 $l=2.35e-06 $layer=LI1_cond $X=3.55 $Y=0 $X2=1.2
+ $Y2=0
r85 29 43 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r86 28 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r87 26 42 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.565 $Y=0 $X2=0.73
+ $Y2=0
r88 26 28 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.565 $Y=0 $X2=0.24
+ $Y2=0
r89 24 46 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=2.88 $Y=0 $X2=3.6
+ $Y2=0
r90 24 35 0.468274 $w=4.9e-07 $l=1.68e-06 $layer=MET1_cond $X=2.88 $Y=0 $X2=1.2
+ $Y2=0
r91 20 48 2.7522 $w=6.65e-07 $l=8.5e-08 $layer=LI1_cond $X=4.812 $Y=0.085
+ $X2=4.812 $Y2=0
r92 20 22 9.71252 $w=6.63e-07 $l=5.4e-07 $layer=LI1_cond $X=4.812 $Y=0.085
+ $X2=4.812 $Y2=0.625
r93 19 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.88 $Y=0 $X2=3.715
+ $Y2=0
r94 18 48 13.2917 $w=1.7e-07 $l=3.32e-07 $layer=LI1_cond $X=4.48 $Y=0 $X2=4.812
+ $Y2=0
r95 18 19 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=4.48 $Y=0 $X2=3.88
+ $Y2=0
r96 14 45 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.715 $Y=0.085
+ $X2=3.715 $Y2=0
r97 14 16 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=3.715 $Y=0.085
+ $X2=3.715 $Y2=0.495
r98 10 42 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.73 $Y=0.085
+ $X2=0.73 $Y2=0
r99 10 12 16.9374 $w=3.28e-07 $l=4.85e-07 $layer=LI1_cond $X=0.73 $Y=0.085
+ $X2=0.73 $Y2=0.57
r100 3 22 91 $w=1.7e-07 $l=7.31471e-07 $layer=licon1_NDIFF $count=2 $X=4.435
+ $Y=0.37 $X2=5.05 $Y2=0.625
r101 2 16 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=3.505
+ $Y=0.37 $X2=3.715 $Y2=0.495
r102 1 12 182 $w=1.7e-07 $l=2.60768e-07 $layer=licon1_NDIFF $count=1 $X=0.59
+ $Y=0.37 $X2=0.73 $Y2=0.57
.ends

.subckt PM_SKY130_FD_SC_HS__NAND2B_4%A_243_74# 1 2 3 4 5 18 20 21 24 26 31 32 33
+ 36 38 42 44 45
c88 38 0 1.19111e-20 $X=5.315 $Y=1.045
c89 26 0 9.27061e-20 $X=3.05 $Y=0.34
r90 48 49 3.66686 $w=3.28e-07 $l=1.05e-07 $layer=LI1_cond $X=4.145 $Y=0.94
+ $X2=4.145 $Y2=1.045
r91 45 48 3.66686 $w=3.28e-07 $l=1.05e-07 $layer=LI1_cond $X=4.145 $Y=0.835
+ $X2=4.145 $Y2=0.94
r92 45 46 3.51899 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=4.145 $Y=0.835
+ $X2=4.145 $Y2=0.75
r93 40 42 15.5405 $w=3.28e-07 $l=4.45e-07 $layer=LI1_cond $X=5.48 $Y=0.96
+ $X2=5.48 $Y2=0.515
r94 39 49 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.31 $Y=1.045
+ $X2=4.145 $Y2=1.045
r95 38 40 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=5.315 $Y=1.045
+ $X2=5.48 $Y2=0.96
r96 38 39 65.5668 $w=1.68e-07 $l=1.005e-06 $layer=LI1_cond $X=5.315 $Y=1.045
+ $X2=4.31 $Y2=1.045
r97 36 46 11.3028 $w=2.58e-07 $l=2.55e-07 $layer=LI1_cond $X=4.18 $Y=0.495
+ $X2=4.18 $Y2=0.75
r98 32 45 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.98 $Y=0.835
+ $X2=4.145 $Y2=0.835
r99 32 33 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=3.98 $Y=0.835 $X2=3.38
+ $Y2=0.835
r100 29 33 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.215 $Y=0.75
+ $X2=3.38 $Y2=0.835
r101 29 31 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=3.215 $Y=0.75
+ $X2=3.215 $Y2=0.495
r102 28 31 2.44458 $w=3.28e-07 $l=7e-08 $layer=LI1_cond $X=3.215 $Y=0.425
+ $X2=3.215 $Y2=0.495
r103 27 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.385 $Y=0.34
+ $X2=2.22 $Y2=0.34
r104 26 28 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.05 $Y=0.34
+ $X2=3.215 $Y2=0.425
r105 26 27 43.385 $w=1.68e-07 $l=6.65e-07 $layer=LI1_cond $X=3.05 $Y=0.34
+ $X2=2.385 $Y2=0.34
r106 22 44 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.22 $Y=0.425
+ $X2=2.22 $Y2=0.34
r107 22 24 2.44458 $w=3.28e-07 $l=7e-08 $layer=LI1_cond $X=2.22 $Y=0.425
+ $X2=2.22 $Y2=0.495
r108 20 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.055 $Y=0.34
+ $X2=2.22 $Y2=0.34
r109 20 21 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=2.055 $Y=0.34
+ $X2=1.455 $Y2=0.34
r110 16 21 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=1.325 $Y=0.425
+ $X2=1.455 $Y2=0.34
r111 16 18 6.42709 $w=2.58e-07 $l=1.45e-07 $layer=LI1_cond $X=1.325 $Y=0.425
+ $X2=1.325 $Y2=0.57
r112 5 42 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=5.34
+ $Y=0.37 $X2=5.48 $Y2=0.515
r113 4 48 182 $w=1.7e-07 $l=6.3616e-07 $layer=licon1_NDIFF $count=1 $X=4.005
+ $Y=0.37 $X2=4.145 $Y2=0.94
r114 4 36 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=4.005
+ $Y=0.37 $X2=4.145 $Y2=0.495
r115 3 31 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=3.075
+ $Y=0.37 $X2=3.215 $Y2=0.495
r116 2 24 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=2.08
+ $Y=0.37 $X2=2.22 $Y2=0.495
r117 1 18 182 $w=1.7e-07 $l=2.62678e-07 $layer=licon1_NDIFF $count=1 $X=1.215
+ $Y=0.37 $X2=1.36 $Y2=0.57
.ends

