* File: sky130_fd_sc_hs__xnor2_2.spice
* Created: Tue Sep  1 20:25:16 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hs__xnor2_2.pex.spice"
.subckt sky130_fd_sc_hs__xnor2_2  VNB VPB A B VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* B	B
* A	A
* VPB	VPB
* VNB	VNB
MM1011 A_151_74# N_A_M1011_g N_VGND_M1011_s VNB NLOWVT L=0.15 W=0.74 AD=0.0888
+ AS=0.25 PD=0.98 PS=2.44 NRD=10.536 NRS=21.888 M=1 R=4.93333 SA=75000.3
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1010 N_A_133_368#_M1010_d N_B_M1010_g A_151_74# VNB NLOWVT L=0.15 W=0.74
+ AD=0.206875 AS=0.0888 PD=2.05 PS=0.98 NRD=0 NRS=10.536 M=1 R=4.93333
+ SA=75000.6 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1001 N_Y_M1001_d N_A_133_368#_M1001_g N_A_340_107#_M1001_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.2004 AS=0.197775 PD=1.335 PS=2.05 NRD=17.832 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75002.9 A=0.111 P=1.78 MULT=1
MM1014 N_Y_M1001_d N_A_133_368#_M1014_g N_A_340_107#_M1014_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.2004 AS=0.1036 PD=1.335 PS=1.02 NRD=18.648 NRS=0 M=1 R=4.93333
+ SA=75000.8 SB=75002.3 A=0.111 P=1.78 MULT=1
MM1004 N_VGND_M1004_d N_A_M1004_g N_A_340_107#_M1014_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1912 AS=0.1036 PD=1.365 PS=1.02 NRD=32.976 NRS=0 M=1 R=4.93333 SA=75001.3
+ SB=75001.9 A=0.111 P=1.78 MULT=1
MM1000 N_A_340_107#_M1000_d N_B_M1000_g N_VGND_M1004_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.111 AS=0.1912 PD=1.04 PS=1.365 NRD=0 NRS=32.976 M=1 R=4.93333 SA=75001.9
+ SB=75001.3 A=0.111 P=1.78 MULT=1
MM1002 N_A_340_107#_M1000_d N_B_M1002_g N_VGND_M1002_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.111 AS=0.1958 PD=1.04 PS=1.375 NRD=0 NRS=33.984 M=1 R=4.93333 SA=75002.3
+ SB=75000.8 A=0.111 P=1.78 MULT=1
MM1005 N_VGND_M1002_s N_A_M1005_g N_A_340_107#_M1005_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1958 AS=0.20355 PD=1.375 PS=2.05 NRD=33.984 NRS=0 M=1 R=4.93333
+ SA=75002.9 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1015 N_A_133_368#_M1015_d N_A_M1015_g N_VPWR_M1015_s VPB PSHORT L=0.15 W=1
+ AD=0.1725 AS=0.4177 PD=1.345 PS=3.02 NRD=5.8903 NRS=19.6803 M=1 R=6.66667
+ SA=75000.3 SB=75004.4 A=0.15 P=2.3 MULT=1
MM1003 N_VPWR_M1003_d N_B_M1003_g N_A_133_368#_M1015_d VPB PSHORT L=0.15 W=1
+ AD=0.425684 AS=0.1725 PD=1.83019 PS=1.345 NRD=15.7403 NRS=6.8753 M=1 R=6.66667
+ SA=75000.8 SB=75003.9 A=0.15 P=2.3 MULT=1
MM1012 N_Y_M1012_d N_A_133_368#_M1012_g N_VPWR_M1003_d VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.476766 PD=1.42 PS=2.04981 NRD=1.7533 NRS=7.0329 M=1 R=7.46667
+ SA=75001.6 SB=75002.9 A=0.168 P=2.54 MULT=1
MM1013 N_Y_M1012_d N_A_133_368#_M1013_g N_VPWR_M1013_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.27625 PD=1.42 PS=1.68 NRD=1.7533 NRS=17.5724 M=1 R=7.46667
+ SA=75002.1 SB=75002.5 A=0.168 P=2.54 MULT=1
MM1008 N_VPWR_M1013_s N_A_M1008_g N_A_638_368#_M1008_s VPB PSHORT L=0.15 W=1.12
+ AD=0.27625 AS=0.2823 PD=1.68 PS=1.69 NRD=17.5724 NRS=18.4589 M=1 R=7.46667
+ SA=75002.7 SB=75001.8 A=0.168 P=2.54 MULT=1
MM1006 N_Y_M1006_d N_B_M1006_g N_A_638_368#_M1008_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.2823 PD=1.42 PS=1.69 NRD=1.7533 NRS=18.4589 M=1 R=7.46667
+ SA=75003.3 SB=75001.2 A=0.168 P=2.54 MULT=1
MM1007 N_Y_M1006_d N_B_M1007_g N_A_638_368#_M1007_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.196 PD=1.42 PS=1.47 NRD=1.7533 NRS=10.5395 M=1 R=7.46667
+ SA=75003.8 SB=75000.8 A=0.168 P=2.54 MULT=1
MM1009 N_VPWR_M1009_d N_A_M1009_g N_A_638_368#_M1007_s VPB PSHORT L=0.15 W=1.12
+ AD=0.3864 AS=0.196 PD=2.93 PS=1.47 NRD=10.5395 NRS=1.7533 M=1 R=7.46667
+ SA=75004.3 SB=75000.3 A=0.168 P=2.54 MULT=1
DX16_noxref VNB VPB NWDIODE A=10.5276 P=15.04
*
.include "sky130_fd_sc_hs__xnor2_2.pxi.spice"
*
.ends
*
*
