* File: sky130_fd_sc_hs__o221ai_2.pxi.spice
* Created: Thu Aug 27 20:59:44 2020
* 
x_PM_SKY130_FD_SC_HS__O221AI_2%C1 N_C1_M1015_g N_C1_c_96_n N_C1_M1018_g
+ N_C1_M1016_g N_C1_c_97_n N_C1_M1019_g C1 N_C1_c_94_n N_C1_c_95_n
+ PM_SKY130_FD_SC_HS__O221AI_2%C1
x_PM_SKY130_FD_SC_HS__O221AI_2%B1 N_B1_c_135_n N_B1_M1012_g N_B1_c_136_n
+ N_B1_M1007_g N_B1_c_137_n N_B1_M1013_g N_B1_M1011_g N_B1_c_151_p N_B1_c_139_n
+ B1 B1 B1 N_B1_c_140_n PM_SKY130_FD_SC_HS__O221AI_2%B1
x_PM_SKY130_FD_SC_HS__O221AI_2%B2 N_B2_c_222_n N_B2_M1005_g N_B2_M1001_g
+ N_B2_c_223_n N_B2_M1014_g N_B2_M1004_g B2 N_B2_c_220_n N_B2_c_221_n
+ PM_SKY130_FD_SC_HS__O221AI_2%B2
x_PM_SKY130_FD_SC_HS__O221AI_2%A1 N_A1_M1003_g N_A1_c_270_n N_A1_M1000_g
+ N_A1_c_271_n N_A1_M1009_g N_A1_M1017_g N_A1_c_273_n N_A1_c_290_p N_A1_c_285_n
+ A1 N_A1_c_274_n PM_SKY130_FD_SC_HS__O221AI_2%A1
x_PM_SKY130_FD_SC_HS__O221AI_2%A2 N_A2_M1002_g N_A2_c_353_n N_A2_M1008_g
+ N_A2_c_354_n N_A2_M1010_g N_A2_M1006_g A2 N_A2_c_351_n N_A2_c_352_n
+ PM_SKY130_FD_SC_HS__O221AI_2%A2
x_PM_SKY130_FD_SC_HS__O221AI_2%VPWR N_VPWR_M1018_s N_VPWR_M1019_s N_VPWR_M1013_s
+ N_VPWR_M1009_d N_VPWR_c_404_n N_VPWR_c_405_n N_VPWR_c_406_n N_VPWR_c_407_n
+ N_VPWR_c_408_n VPWR N_VPWR_c_409_n N_VPWR_c_410_n N_VPWR_c_411_n
+ N_VPWR_c_412_n N_VPWR_c_413_n N_VPWR_c_403_n PM_SKY130_FD_SC_HS__O221AI_2%VPWR
x_PM_SKY130_FD_SC_HS__O221AI_2%Y N_Y_M1015_d N_Y_M1018_d N_Y_M1005_d N_Y_M1008_d
+ N_Y_c_487_n N_Y_c_502_n N_Y_c_477_n N_Y_c_491_n Y Y Y Y Y Y
+ PM_SKY130_FD_SC_HS__O221AI_2%Y
x_PM_SKY130_FD_SC_HS__O221AI_2%A_376_368# N_A_376_368#_M1012_d
+ N_A_376_368#_M1014_s N_A_376_368#_c_535_n N_A_376_368#_c_536_n
+ N_A_376_368#_c_537_n PM_SKY130_FD_SC_HS__O221AI_2%A_376_368#
x_PM_SKY130_FD_SC_HS__O221AI_2%A_776_368# N_A_776_368#_M1000_s
+ N_A_776_368#_M1010_s N_A_776_368#_c_563_n N_A_776_368#_c_571_n
+ N_A_776_368#_c_564_n PM_SKY130_FD_SC_HS__O221AI_2%A_776_368#
x_PM_SKY130_FD_SC_HS__O221AI_2%A_27_74# N_A_27_74#_M1015_s N_A_27_74#_M1016_s
+ N_A_27_74#_M1007_d N_A_27_74#_M1004_s N_A_27_74#_c_593_n N_A_27_74#_c_594_n
+ N_A_27_74#_c_595_n N_A_27_74#_c_596_n N_A_27_74#_c_597_n N_A_27_74#_c_598_n
+ N_A_27_74#_c_633_p N_A_27_74#_c_599_n N_A_27_74#_c_618_n N_A_27_74#_c_600_n
+ PM_SKY130_FD_SC_HS__O221AI_2%A_27_74#
x_PM_SKY130_FD_SC_HS__O221AI_2%A_311_85# N_A_311_85#_M1007_s N_A_311_85#_M1001_d
+ N_A_311_85#_M1011_s N_A_311_85#_M1002_d N_A_311_85#_M1017_s
+ N_A_311_85#_c_644_n N_A_311_85#_c_645_n N_A_311_85#_c_646_n
+ N_A_311_85#_c_659_n N_A_311_85#_c_647_n N_A_311_85#_c_670_n
+ N_A_311_85#_c_648_n N_A_311_85#_c_649_n N_A_311_85#_c_650_n
+ N_A_311_85#_c_651_n N_A_311_85#_c_652_n N_A_311_85#_c_653_n
+ N_A_311_85#_c_654_n PM_SKY130_FD_SC_HS__O221AI_2%A_311_85#
x_PM_SKY130_FD_SC_HS__O221AI_2%VGND N_VGND_M1003_d N_VGND_M1006_s N_VGND_c_723_n
+ N_VGND_c_724_n VGND N_VGND_c_725_n N_VGND_c_726_n N_VGND_c_727_n
+ N_VGND_c_728_n N_VGND_c_729_n N_VGND_c_730_n PM_SKY130_FD_SC_HS__O221AI_2%VGND
cc_1 VNB N_C1_M1015_g 0.0274728f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_2 VNB N_C1_M1016_g 0.025282f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=0.74
cc_3 VNB N_C1_c_94_n 0.00617983f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.465
cc_4 VNB N_C1_c_95_n 0.0979341f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=1.532
cc_5 VNB N_B1_c_135_n 0.0331326f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.3
cc_6 VNB N_B1_c_136_n 0.0215291f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_7 VNB N_B1_c_137_n 0.0268444f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=2.4
cc_8 VNB N_B1_M1011_g 0.021044f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=1.765
cc_9 VNB N_B1_c_139_n 0.00167757f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.465
cc_10 VNB N_B1_c_140_n 0.0119268f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_B2_M1001_g 0.0192446f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=2.4
cc_12 VNB N_B2_M1004_g 0.0206166f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=2.4
cc_13 VNB N_B2_c_220_n 8.29228e-19 $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=1.532
cc_14 VNB N_B2_c_221_n 0.0331819f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=1.532
cc_15 VNB N_A1_M1003_g 0.0211602f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_16 VNB N_A1_c_270_n 0.0270041f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=1.765
cc_17 VNB N_A1_c_271_n 0.0288661f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=1.3
cc_18 VNB N_A1_M1017_g 0.0288546f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=2.4
cc_19 VNB N_A1_c_273_n 0.00167078f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.532
cc_20 VNB N_A1_c_274_n 0.0202222f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A2_M1002_g 0.0219922f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_22 VNB N_A2_M1006_g 0.0214811f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=2.4
cc_23 VNB N_A2_c_351_n 0.00139482f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=1.532
cc_24 VNB N_A2_c_352_n 0.036617f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=1.532
cc_25 VNB N_VPWR_c_403_n 0.243291f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB Y 0.00220761f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.465
cc_27 VNB N_A_27_74#_c_593_n 0.0275751f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_28 VNB N_A_27_74#_c_594_n 0.00664238f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.532
cc_29 VNB N_A_27_74#_c_595_n 0.00931596f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.465
cc_30 VNB N_A_27_74#_c_596_n 0.0062256f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=1.532
cc_31 VNB N_A_27_74#_c_597_n 0.0143267f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=1.532
cc_32 VNB N_A_27_74#_c_598_n 0.00353358f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.465
cc_33 VNB N_A_27_74#_c_599_n 0.0147249f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_27_74#_c_600_n 0.00157355f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_311_85#_c_644_n 0.00367062f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.465
cc_36 VNB N_A_311_85#_c_645_n 0.00702435f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.532
cc_37 VNB N_A_311_85#_c_646_n 0.00454744f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=1.532
cc_38 VNB N_A_311_85#_c_647_n 0.0135463f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.665
cc_39 VNB N_A_311_85#_c_648_n 0.00924121f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_311_85#_c_649_n 0.00789247f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_311_85#_c_650_n 0.00316307f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_311_85#_c_651_n 0.0148853f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_311_85#_c_652_n 0.0249008f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_311_85#_c_653_n 0.00238018f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_A_311_85#_c_654_n 0.00312418f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_VGND_c_723_n 0.0108406f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=0.74
cc_47 VNB N_VGND_c_724_n 0.00891632f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=2.4
cc_48 VNB N_VGND_c_725_n 0.0937136f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.532
cc_49 VNB N_VGND_c_726_n 0.0189057f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_VGND_c_727_n 0.0178712f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_VGND_c_728_n 0.34449f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_VGND_c_729_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_VGND_c_730_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VPB N_C1_c_96_n 0.0175845f $X=-0.19 $Y=1.66 $X2=0.545 $Y2=1.765
cc_55 VPB N_C1_c_97_n 0.0170243f $X=-0.19 $Y=1.66 $X2=0.995 $Y2=1.765
cc_56 VPB N_C1_c_94_n 0.0106053f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.465
cc_57 VPB N_C1_c_95_n 0.0139891f $X=-0.19 $Y=1.66 $X2=0.925 $Y2=1.532
cc_58 VPB N_B1_c_135_n 0.0282484f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.3
cc_59 VPB N_B1_c_137_n 0.026612f $X=-0.19 $Y=1.66 $X2=0.545 $Y2=2.4
cc_60 VPB N_B1_c_139_n 0.00252244f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.465
cc_61 VPB N_B1_c_140_n 0.00289424f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_62 VPB N_B2_c_222_n 0.014851f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.3
cc_63 VPB N_B2_c_223_n 0.0152444f $X=-0.19 $Y=1.66 $X2=0.925 $Y2=1.3
cc_64 VPB N_B2_c_220_n 0.00305195f $X=-0.19 $Y=1.66 $X2=0.545 $Y2=1.532
cc_65 VPB N_B2_c_221_n 0.0199107f $X=-0.19 $Y=1.66 $X2=0.925 $Y2=1.532
cc_66 VPB N_A1_c_270_n 0.0266274f $X=-0.19 $Y=1.66 $X2=0.545 $Y2=1.765
cc_67 VPB N_A1_c_271_n 0.0279928f $X=-0.19 $Y=1.66 $X2=0.925 $Y2=1.3
cc_68 VPB N_A1_c_273_n 0.00266333f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.532
cc_69 VPB N_A1_c_274_n 0.020571f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_70 VPB N_A2_c_353_n 0.0152057f $X=-0.19 $Y=1.66 $X2=0.545 $Y2=1.765
cc_71 VPB N_A2_c_354_n 0.0148813f $X=-0.19 $Y=1.66 $X2=0.925 $Y2=1.3
cc_72 VPB N_A2_c_351_n 0.00283822f $X=-0.19 $Y=1.66 $X2=0.545 $Y2=1.532
cc_73 VPB N_A2_c_352_n 0.0201893f $X=-0.19 $Y=1.66 $X2=0.925 $Y2=1.532
cc_74 VPB N_VPWR_c_404_n 0.011928f $X=-0.19 $Y=1.66 $X2=0.995 $Y2=2.4
cc_75 VPB N_VPWR_c_405_n 0.0488362f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_76 VPB N_VPWR_c_406_n 0.00888536f $X=-0.19 $Y=1.66 $X2=0.545 $Y2=1.532
cc_77 VPB N_VPWR_c_407_n 0.0121872f $X=-0.19 $Y=1.66 $X2=0.995 $Y2=1.532
cc_78 VPB N_VPWR_c_408_n 0.0387973f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_79 VPB N_VPWR_c_409_n 0.0185562f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_80 VPB N_VPWR_c_410_n 0.0401022f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_81 VPB N_VPWR_c_411_n 0.0389463f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_82 VPB N_VPWR_c_412_n 0.02096f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_83 VPB N_VPWR_c_413_n 0.00631492f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_84 VPB N_VPWR_c_403_n 0.0735095f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_85 VPB Y 0.00126282f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.465
cc_86 VPB Y 0.00216998f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_87 VPB N_A_376_368#_c_535_n 0.00310533f $X=-0.19 $Y=1.66 $X2=0.545 $Y2=2.4
cc_88 VPB N_A_376_368#_c_536_n 0.00247979f $X=-0.19 $Y=1.66 $X2=0.925 $Y2=0.74
cc_89 VPB N_A_376_368#_c_537_n 0.00248006f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_90 VPB N_A_776_368#_c_563_n 0.00480458f $X=-0.19 $Y=1.66 $X2=0.545 $Y2=2.4
cc_91 VPB N_A_776_368#_c_564_n 0.00248006f $X=-0.19 $Y=1.66 $X2=0.995 $Y2=2.4
cc_92 N_C1_M1016_g N_B1_c_135_n 2.45528e-19 $X=0.925 $Y=0.74 $X2=-0.19
+ $Y2=-0.245
cc_93 N_C1_c_97_n N_B1_c_135_n 0.0138862f $X=0.995 $Y=1.765 $X2=-0.19 $Y2=-0.245
cc_94 N_C1_c_95_n N_B1_c_135_n 0.00819054f $X=0.925 $Y=1.532 $X2=-0.19
+ $Y2=-0.245
cc_95 N_C1_c_97_n N_B1_c_140_n 0.00361726f $X=0.995 $Y=1.765 $X2=0 $Y2=0
cc_96 N_C1_c_95_n N_B1_c_140_n 0.00668078f $X=0.925 $Y=1.532 $X2=0 $Y2=0
cc_97 N_C1_c_96_n N_VPWR_c_405_n 0.00700598f $X=0.545 $Y=1.765 $X2=0 $Y2=0
cc_98 N_C1_c_94_n N_VPWR_c_405_n 0.0222392f $X=0.27 $Y=1.465 $X2=0 $Y2=0
cc_99 N_C1_c_95_n N_VPWR_c_405_n 0.0013689f $X=0.925 $Y=1.532 $X2=0 $Y2=0
cc_100 N_C1_c_96_n N_VPWR_c_409_n 0.00445602f $X=0.545 $Y=1.765 $X2=0 $Y2=0
cc_101 N_C1_c_97_n N_VPWR_c_409_n 0.00415318f $X=0.995 $Y=1.765 $X2=0 $Y2=0
cc_102 N_C1_c_96_n N_VPWR_c_412_n 4.49144e-19 $X=0.545 $Y=1.765 $X2=0 $Y2=0
cc_103 N_C1_c_97_n N_VPWR_c_412_n 0.00863491f $X=0.995 $Y=1.765 $X2=0 $Y2=0
cc_104 N_C1_c_96_n N_VPWR_c_403_n 0.00861209f $X=0.545 $Y=1.765 $X2=0 $Y2=0
cc_105 N_C1_c_97_n N_VPWR_c_403_n 0.00817726f $X=0.995 $Y=1.765 $X2=0 $Y2=0
cc_106 N_C1_c_97_n N_Y_c_477_n 0.0182839f $X=0.995 $Y=1.765 $X2=0 $Y2=0
cc_107 N_C1_M1015_g Y 0.00526147f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_108 N_C1_c_96_n Y 0.0118459f $X=0.545 $Y=1.765 $X2=0 $Y2=0
cc_109 N_C1_M1016_g Y 0.0147581f $X=0.925 $Y=0.74 $X2=0 $Y2=0
cc_110 N_C1_c_97_n Y 7.33691e-19 $X=0.995 $Y=1.765 $X2=0 $Y2=0
cc_111 N_C1_c_94_n Y 0.0360521f $X=0.27 $Y=1.465 $X2=0 $Y2=0
cc_112 N_C1_c_95_n Y 0.031229f $X=0.925 $Y=1.532 $X2=0 $Y2=0
cc_113 N_C1_c_96_n Y 0.00797844f $X=0.545 $Y=1.765 $X2=0 $Y2=0
cc_114 N_C1_c_97_n Y 0.00499464f $X=0.995 $Y=1.765 $X2=0 $Y2=0
cc_115 N_C1_M1015_g N_A_27_74#_c_593_n 0.00161118f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_116 N_C1_c_94_n N_A_27_74#_c_593_n 0.0215684f $X=0.27 $Y=1.465 $X2=0 $Y2=0
cc_117 N_C1_c_95_n N_A_27_74#_c_593_n 0.00196285f $X=0.925 $Y=1.532 $X2=0 $Y2=0
cc_118 N_C1_M1015_g N_A_27_74#_c_594_n 0.0139957f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_119 N_C1_M1016_g N_A_27_74#_c_594_n 0.0132617f $X=0.925 $Y=0.74 $X2=0 $Y2=0
cc_120 N_C1_M1016_g N_A_27_74#_c_598_n 0.00162302f $X=0.925 $Y=0.74 $X2=0 $Y2=0
cc_121 N_C1_c_95_n N_A_27_74#_c_598_n 0.00149613f $X=0.925 $Y=1.532 $X2=0 $Y2=0
cc_122 N_C1_M1016_g N_A_311_85#_c_646_n 5.96586e-19 $X=0.925 $Y=0.74 $X2=0 $Y2=0
cc_123 N_C1_M1015_g N_VGND_c_725_n 0.00278271f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_124 N_C1_M1016_g N_VGND_c_725_n 0.00278271f $X=0.925 $Y=0.74 $X2=0 $Y2=0
cc_125 N_C1_M1015_g N_VGND_c_728_n 0.00357086f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_126 N_C1_M1016_g N_VGND_c_728_n 0.00358427f $X=0.925 $Y=0.74 $X2=0 $Y2=0
cc_127 N_B1_c_135_n N_B2_c_222_n 0.0364391f $X=1.805 $Y=1.765 $X2=-0.19
+ $Y2=-0.245
cc_128 N_B1_c_151_p N_B2_c_222_n 0.00877506f $X=3.075 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_129 N_B1_c_140_n N_B2_c_222_n 0.0106898f $X=2.275 $Y=1.735 $X2=-0.19
+ $Y2=-0.245
cc_130 N_B1_c_136_n N_B2_M1001_g 0.0167366f $X=1.915 $Y=1.29 $X2=0 $Y2=0
cc_131 N_B1_c_137_n N_B2_c_223_n 0.0387809f $X=3.255 $Y=1.765 $X2=0 $Y2=0
cc_132 N_B1_c_151_p N_B2_c_223_n 0.0110248f $X=3.075 $Y=2.035 $X2=0 $Y2=0
cc_133 N_B1_c_139_n N_B2_c_223_n 0.00380443f $X=3.24 $Y=1.515 $X2=0 $Y2=0
cc_134 N_B1_c_140_n N_B2_c_223_n 8.75562e-19 $X=2.275 $Y=1.735 $X2=0 $Y2=0
cc_135 N_B1_M1011_g N_B2_M1004_g 0.0194733f $X=3.33 $Y=0.795 $X2=0 $Y2=0
cc_136 N_B1_c_137_n N_B2_c_220_n 0.00149884f $X=3.255 $Y=1.765 $X2=0 $Y2=0
cc_137 N_B1_c_151_p N_B2_c_220_n 0.0224724f $X=3.075 $Y=2.035 $X2=0 $Y2=0
cc_138 N_B1_c_139_n N_B2_c_220_n 0.0266359f $X=3.24 $Y=1.515 $X2=0 $Y2=0
cc_139 N_B1_c_140_n N_B2_c_220_n 0.0259253f $X=2.275 $Y=1.735 $X2=0 $Y2=0
cc_140 N_B1_c_135_n N_B2_c_221_n 0.0307043f $X=1.805 $Y=1.765 $X2=0 $Y2=0
cc_141 N_B1_c_137_n N_B2_c_221_n 0.0225823f $X=3.255 $Y=1.765 $X2=0 $Y2=0
cc_142 N_B1_c_151_p N_B2_c_221_n 0.00526911f $X=3.075 $Y=2.035 $X2=0 $Y2=0
cc_143 N_B1_c_139_n N_B2_c_221_n 0.0016488f $X=3.24 $Y=1.515 $X2=0 $Y2=0
cc_144 N_B1_c_140_n N_B2_c_221_n 0.0140197f $X=2.275 $Y=1.735 $X2=0 $Y2=0
cc_145 N_B1_M1011_g N_A1_M1003_g 0.0172352f $X=3.33 $Y=0.795 $X2=0 $Y2=0
cc_146 N_B1_c_137_n N_A1_c_270_n 0.0562037f $X=3.255 $Y=1.765 $X2=0 $Y2=0
cc_147 N_B1_c_151_p N_A1_c_270_n 6.60789e-19 $X=3.075 $Y=2.035 $X2=0 $Y2=0
cc_148 N_B1_c_139_n N_A1_c_270_n 0.00213389f $X=3.24 $Y=1.515 $X2=0 $Y2=0
cc_149 N_B1_c_137_n N_A1_c_273_n 0.00215343f $X=3.255 $Y=1.765 $X2=0 $Y2=0
cc_150 N_B1_c_139_n N_A1_c_273_n 0.0360504f $X=3.24 $Y=1.515 $X2=0 $Y2=0
cc_151 N_B1_c_137_n N_A1_c_285_n 6.74604e-19 $X=3.255 $Y=1.765 $X2=0 $Y2=0
cc_152 N_B1_c_151_p N_A1_c_285_n 0.0118527f $X=3.075 $Y=2.035 $X2=0 $Y2=0
cc_153 N_B1_c_140_n N_VPWR_M1019_s 0.0123684f $X=2.275 $Y=1.735 $X2=0 $Y2=0
cc_154 N_B1_c_151_p N_VPWR_M1013_s 0.0019941f $X=3.075 $Y=2.035 $X2=0 $Y2=0
cc_155 N_B1_c_139_n N_VPWR_M1013_s 0.00113608f $X=3.24 $Y=1.515 $X2=0 $Y2=0
cc_156 N_B1_c_137_n N_VPWR_c_406_n 0.00344761f $X=3.255 $Y=1.765 $X2=0 $Y2=0
cc_157 N_B1_c_135_n N_VPWR_c_410_n 0.00444353f $X=1.805 $Y=1.765 $X2=0 $Y2=0
cc_158 N_B1_c_137_n N_VPWR_c_410_n 0.00444353f $X=3.255 $Y=1.765 $X2=0 $Y2=0
cc_159 N_B1_c_135_n N_VPWR_c_412_n 0.00196266f $X=1.805 $Y=1.765 $X2=0 $Y2=0
cc_160 N_B1_c_135_n N_VPWR_c_403_n 0.00859247f $X=1.805 $Y=1.765 $X2=0 $Y2=0
cc_161 N_B1_c_137_n N_VPWR_c_403_n 0.00857817f $X=3.255 $Y=1.765 $X2=0 $Y2=0
cc_162 N_B1_c_151_p N_Y_M1005_d 0.00426668f $X=3.075 $Y=2.035 $X2=0 $Y2=0
cc_163 N_B1_c_137_n N_Y_c_487_n 0.0156632f $X=3.255 $Y=1.765 $X2=0 $Y2=0
cc_164 N_B1_c_151_p N_Y_c_487_n 0.0167062f $X=3.075 $Y=2.035 $X2=0 $Y2=0
cc_165 N_B1_c_135_n N_Y_c_477_n 0.016416f $X=1.805 $Y=1.765 $X2=0 $Y2=0
cc_166 N_B1_c_140_n N_Y_c_477_n 0.0618215f $X=2.275 $Y=1.735 $X2=0 $Y2=0
cc_167 N_B1_c_137_n N_Y_c_491_n 7.44665e-19 $X=3.255 $Y=1.765 $X2=0 $Y2=0
cc_168 N_B1_c_151_p N_Y_c_491_n 0.0618215f $X=3.075 $Y=2.035 $X2=0 $Y2=0
cc_169 N_B1_c_140_n Y 0.0337483f $X=2.275 $Y=1.735 $X2=0 $Y2=0
cc_170 N_B1_c_140_n N_A_376_368#_M1012_d 0.00245767f $X=2.275 $Y=1.735 $X2=-0.19
+ $Y2=-0.245
cc_171 N_B1_c_151_p N_A_376_368#_M1014_s 0.00964917f $X=3.075 $Y=2.035 $X2=0
+ $Y2=0
cc_172 N_B1_c_139_n N_A_376_368#_M1014_s 0.00144886f $X=3.24 $Y=1.515 $X2=0
+ $Y2=0
cc_173 N_B1_c_135_n N_A_376_368#_c_536_n 0.00603755f $X=1.805 $Y=1.765 $X2=0
+ $Y2=0
cc_174 N_B1_c_137_n N_A_376_368#_c_537_n 0.00591159f $X=3.255 $Y=1.765 $X2=0
+ $Y2=0
cc_175 N_B1_c_136_n N_A_27_74#_c_594_n 5.53247e-19 $X=1.915 $Y=1.29 $X2=0 $Y2=0
cc_176 N_B1_c_136_n N_A_27_74#_c_596_n 0.00501983f $X=1.915 $Y=1.29 $X2=0 $Y2=0
cc_177 N_B1_c_135_n N_A_27_74#_c_597_n 0.00561567f $X=1.805 $Y=1.765 $X2=0 $Y2=0
cc_178 N_B1_c_136_n N_A_27_74#_c_597_n 0.0133087f $X=1.915 $Y=1.29 $X2=0 $Y2=0
cc_179 N_B1_c_140_n N_A_27_74#_c_597_n 0.0599647f $X=2.275 $Y=1.735 $X2=0 $Y2=0
cc_180 N_B1_c_140_n N_A_27_74#_c_598_n 0.0205272f $X=2.275 $Y=1.735 $X2=0 $Y2=0
cc_181 N_B1_c_137_n N_A_27_74#_c_599_n 0.00138414f $X=3.255 $Y=1.765 $X2=0 $Y2=0
cc_182 N_B1_M1011_g N_A_27_74#_c_599_n 0.00232271f $X=3.33 $Y=0.795 $X2=0 $Y2=0
cc_183 N_B1_c_139_n N_A_27_74#_c_599_n 0.0178644f $X=3.24 $Y=1.515 $X2=0 $Y2=0
cc_184 N_B1_c_140_n N_A_27_74#_c_599_n 0.00496728f $X=2.275 $Y=1.735 $X2=0 $Y2=0
cc_185 N_B1_M1011_g N_A_27_74#_c_618_n 0.0046047f $X=3.33 $Y=0.795 $X2=0 $Y2=0
cc_186 N_B1_c_140_n N_A_27_74#_c_600_n 0.0156866f $X=2.275 $Y=1.735 $X2=0 $Y2=0
cc_187 N_B1_c_136_n N_A_311_85#_c_644_n 0.00631411f $X=1.915 $Y=1.29 $X2=0 $Y2=0
cc_188 N_B1_c_136_n N_A_311_85#_c_645_n 0.00817976f $X=1.915 $Y=1.29 $X2=0 $Y2=0
cc_189 N_B1_c_136_n N_A_311_85#_c_646_n 0.0032816f $X=1.915 $Y=1.29 $X2=0 $Y2=0
cc_190 N_B1_c_136_n N_A_311_85#_c_659_n 5.66812e-19 $X=1.915 $Y=1.29 $X2=0 $Y2=0
cc_191 N_B1_M1011_g N_A_311_85#_c_659_n 5.11849e-19 $X=3.33 $Y=0.795 $X2=0 $Y2=0
cc_192 N_B1_M1011_g N_A_311_85#_c_647_n 0.01343f $X=3.33 $Y=0.795 $X2=0 $Y2=0
cc_193 N_B1_c_136_n N_VGND_c_725_n 8.82278e-19 $X=1.915 $Y=1.29 $X2=0 $Y2=0
cc_194 N_B1_M1011_g N_VGND_c_725_n 8.63546e-19 $X=3.33 $Y=0.795 $X2=0 $Y2=0
cc_195 N_B2_c_222_n N_VPWR_c_410_n 0.00278271f $X=2.29 $Y=1.765 $X2=0 $Y2=0
cc_196 N_B2_c_223_n N_VPWR_c_410_n 0.00278271f $X=2.755 $Y=1.765 $X2=0 $Y2=0
cc_197 N_B2_c_222_n N_VPWR_c_403_n 0.00354355f $X=2.29 $Y=1.765 $X2=0 $Y2=0
cc_198 N_B2_c_223_n N_VPWR_c_403_n 0.0035448f $X=2.755 $Y=1.765 $X2=0 $Y2=0
cc_199 N_B2_c_223_n N_Y_c_487_n 0.0094057f $X=2.755 $Y=1.765 $X2=0 $Y2=0
cc_200 N_B2_c_222_n N_Y_c_477_n 0.0101212f $X=2.29 $Y=1.765 $X2=0 $Y2=0
cc_201 N_B2_c_222_n N_Y_c_491_n 9.47616e-19 $X=2.29 $Y=1.765 $X2=0 $Y2=0
cc_202 N_B2_c_223_n N_Y_c_491_n 0.00550771f $X=2.755 $Y=1.765 $X2=0 $Y2=0
cc_203 N_B2_c_222_n N_A_376_368#_c_535_n 0.00927258f $X=2.29 $Y=1.765 $X2=0
+ $Y2=0
cc_204 N_B2_c_223_n N_A_376_368#_c_535_n 0.00955976f $X=2.755 $Y=1.765 $X2=0
+ $Y2=0
cc_205 N_B2_c_222_n N_A_376_368#_c_536_n 4.3059e-19 $X=2.29 $Y=1.765 $X2=0 $Y2=0
cc_206 N_B2_c_223_n N_A_376_368#_c_537_n 5.05939e-19 $X=2.755 $Y=1.765 $X2=0
+ $Y2=0
cc_207 N_B2_M1001_g N_A_27_74#_c_599_n 0.0155704f $X=2.345 $Y=0.795 $X2=0 $Y2=0
cc_208 N_B2_M1004_g N_A_27_74#_c_599_n 0.0127188f $X=2.775 $Y=0.795 $X2=0 $Y2=0
cc_209 N_B2_c_220_n N_A_27_74#_c_599_n 0.0247257f $X=2.685 $Y=1.515 $X2=0 $Y2=0
cc_210 N_B2_c_221_n N_A_27_74#_c_599_n 0.00127221f $X=2.755 $Y=1.557 $X2=0 $Y2=0
cc_211 N_B2_M1001_g N_A_311_85#_c_644_n 5.66812e-19 $X=2.345 $Y=0.795 $X2=0
+ $Y2=0
cc_212 N_B2_M1001_g N_A_311_85#_c_645_n 0.00817976f $X=2.345 $Y=0.795 $X2=0
+ $Y2=0
cc_213 N_B2_M1001_g N_A_311_85#_c_659_n 0.00603381f $X=2.345 $Y=0.795 $X2=0
+ $Y2=0
cc_214 N_B2_M1004_g N_A_311_85#_c_659_n 0.00647806f $X=2.775 $Y=0.795 $X2=0
+ $Y2=0
cc_215 N_B2_M1004_g N_A_311_85#_c_647_n 0.00866507f $X=2.775 $Y=0.795 $X2=0
+ $Y2=0
cc_216 N_B2_M1001_g N_A_311_85#_c_653_n 0.00221614f $X=2.345 $Y=0.795 $X2=0
+ $Y2=0
cc_217 N_B2_M1004_g N_A_311_85#_c_653_n 0.00221614f $X=2.775 $Y=0.795 $X2=0
+ $Y2=0
cc_218 N_B2_M1001_g N_VGND_c_725_n 8.82278e-19 $X=2.345 $Y=0.795 $X2=0 $Y2=0
cc_219 N_B2_M1004_g N_VGND_c_725_n 8.82278e-19 $X=2.775 $Y=0.795 $X2=0 $Y2=0
cc_220 N_A1_M1003_g N_A2_M1002_g 0.0242339f $X=3.76 $Y=0.795 $X2=0 $Y2=0
cc_221 N_A1_c_270_n N_A2_c_353_n 0.038752f $X=3.805 $Y=1.765 $X2=0 $Y2=0
cc_222 N_A1_c_273_n N_A2_c_353_n 0.00381853f $X=3.81 $Y=1.515 $X2=0 $Y2=0
cc_223 N_A1_c_290_p N_A2_c_353_n 0.0144349f $X=4.925 $Y=2.035 $X2=0 $Y2=0
cc_224 N_A1_c_271_n N_A2_c_354_n 0.025819f $X=5.205 $Y=1.765 $X2=0 $Y2=0
cc_225 N_A1_c_290_p N_A2_c_354_n 0.0184179f $X=4.925 $Y=2.035 $X2=0 $Y2=0
cc_226 N_A1_c_274_n N_A2_c_354_n 0.00556549f $X=5.28 $Y=1.515 $X2=0 $Y2=0
cc_227 N_A1_M1017_g N_A2_M1006_g 0.0286785f $X=5.26 $Y=0.795 $X2=0 $Y2=0
cc_228 N_A1_c_270_n N_A2_c_351_n 0.00109273f $X=3.805 $Y=1.765 $X2=0 $Y2=0
cc_229 N_A1_c_271_n N_A2_c_351_n 3.16521e-19 $X=5.205 $Y=1.765 $X2=0 $Y2=0
cc_230 N_A1_c_273_n N_A2_c_351_n 0.0176718f $X=3.81 $Y=1.515 $X2=0 $Y2=0
cc_231 N_A1_c_290_p N_A2_c_351_n 0.0220806f $X=4.925 $Y=2.035 $X2=0 $Y2=0
cc_232 N_A1_c_274_n N_A2_c_351_n 0.0272575f $X=5.28 $Y=1.515 $X2=0 $Y2=0
cc_233 N_A1_c_270_n N_A2_c_352_n 0.021408f $X=3.805 $Y=1.765 $X2=0 $Y2=0
cc_234 N_A1_c_271_n N_A2_c_352_n 0.0190431f $X=5.205 $Y=1.765 $X2=0 $Y2=0
cc_235 N_A1_c_273_n N_A2_c_352_n 0.00214653f $X=3.81 $Y=1.515 $X2=0 $Y2=0
cc_236 N_A1_c_290_p N_A2_c_352_n 0.00131029f $X=4.925 $Y=2.035 $X2=0 $Y2=0
cc_237 N_A1_c_274_n N_A2_c_352_n 0.00426734f $X=5.28 $Y=1.515 $X2=0 $Y2=0
cc_238 N_A1_c_273_n N_VPWR_M1013_s 0.00113133f $X=3.81 $Y=1.515 $X2=0 $Y2=0
cc_239 N_A1_c_285_n N_VPWR_M1013_s 0.00209749f $X=3.975 $Y=2.035 $X2=0 $Y2=0
cc_240 N_A1_c_274_n N_VPWR_M1009_d 0.00549103f $X=5.28 $Y=1.515 $X2=0 $Y2=0
cc_241 N_A1_c_270_n N_VPWR_c_406_n 0.00344761f $X=3.805 $Y=1.765 $X2=0 $Y2=0
cc_242 N_A1_c_271_n N_VPWR_c_408_n 0.0167564f $X=5.205 $Y=1.765 $X2=0 $Y2=0
cc_243 N_A1_c_274_n N_VPWR_c_408_n 0.0268099f $X=5.28 $Y=1.515 $X2=0 $Y2=0
cc_244 N_A1_c_270_n N_VPWR_c_411_n 0.00444353f $X=3.805 $Y=1.765 $X2=0 $Y2=0
cc_245 N_A1_c_271_n N_VPWR_c_411_n 0.0044313f $X=5.205 $Y=1.765 $X2=0 $Y2=0
cc_246 N_A1_c_270_n N_VPWR_c_403_n 0.00857817f $X=3.805 $Y=1.765 $X2=0 $Y2=0
cc_247 N_A1_c_271_n N_VPWR_c_403_n 0.00856421f $X=5.205 $Y=1.765 $X2=0 $Y2=0
cc_248 N_A1_c_290_p N_Y_M1008_d 0.00381027f $X=4.925 $Y=2.035 $X2=0 $Y2=0
cc_249 N_A1_c_270_n N_Y_c_487_n 0.0156643f $X=3.805 $Y=1.765 $X2=0 $Y2=0
cc_250 N_A1_c_290_p N_Y_c_487_n 0.0385649f $X=4.925 $Y=2.035 $X2=0 $Y2=0
cc_251 N_A1_c_285_n N_Y_c_487_n 0.0167062f $X=3.975 $Y=2.035 $X2=0 $Y2=0
cc_252 N_A1_c_270_n N_Y_c_502_n 7.43872e-19 $X=3.805 $Y=1.765 $X2=0 $Y2=0
cc_253 N_A1_c_273_n N_A_776_368#_M1000_s 0.00146091f $X=3.81 $Y=1.515 $X2=-0.19
+ $Y2=-0.245
cc_254 N_A1_c_290_p N_A_776_368#_M1000_s 0.0096159f $X=4.925 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_255 N_A1_c_285_n N_A_776_368#_M1000_s 4.10458e-19 $X=3.975 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_256 N_A1_c_290_p N_A_776_368#_M1010_s 0.00226438f $X=4.925 $Y=2.035 $X2=0
+ $Y2=0
cc_257 N_A1_c_274_n N_A_776_368#_M1010_s 0.00349324f $X=5.28 $Y=1.515 $X2=0
+ $Y2=0
cc_258 N_A1_c_271_n N_A_776_368#_c_563_n 0.00319436f $X=5.205 $Y=1.765 $X2=0
+ $Y2=0
cc_259 N_A1_c_271_n N_A_776_368#_c_571_n 0.00630539f $X=5.205 $Y=1.765 $X2=0
+ $Y2=0
cc_260 N_A1_c_290_p N_A_776_368#_c_571_n 0.00411595f $X=4.925 $Y=2.035 $X2=0
+ $Y2=0
cc_261 N_A1_c_274_n N_A_776_368#_c_571_n 0.0143966f $X=5.28 $Y=1.515 $X2=0 $Y2=0
cc_262 N_A1_c_270_n N_A_776_368#_c_564_n 0.00591159f $X=3.805 $Y=1.765 $X2=0
+ $Y2=0
cc_263 N_A1_M1003_g N_A_311_85#_c_647_n 0.00322639f $X=3.76 $Y=0.795 $X2=0 $Y2=0
cc_264 N_A1_M1003_g N_A_311_85#_c_670_n 0.0083539f $X=3.76 $Y=0.795 $X2=0 $Y2=0
cc_265 N_A1_M1003_g N_A_311_85#_c_648_n 0.0116199f $X=3.76 $Y=0.795 $X2=0 $Y2=0
cc_266 N_A1_c_270_n N_A_311_85#_c_648_n 9.75223e-19 $X=3.805 $Y=1.765 $X2=0
+ $Y2=0
cc_267 N_A1_c_273_n N_A_311_85#_c_648_n 0.0205962f $X=3.81 $Y=1.515 $X2=0 $Y2=0
cc_268 N_A1_M1003_g N_A_311_85#_c_649_n 8.73939e-19 $X=3.76 $Y=0.795 $X2=0 $Y2=0
cc_269 N_A1_c_270_n N_A_311_85#_c_649_n 3.08675e-19 $X=3.805 $Y=1.765 $X2=0
+ $Y2=0
cc_270 N_A1_c_273_n N_A_311_85#_c_649_n 0.0055933f $X=3.81 $Y=1.515 $X2=0 $Y2=0
cc_271 N_A1_M1017_g N_A_311_85#_c_650_n 9.38284e-19 $X=5.26 $Y=0.795 $X2=0 $Y2=0
cc_272 N_A1_c_271_n N_A_311_85#_c_651_n 0.00130872f $X=5.205 $Y=1.765 $X2=0
+ $Y2=0
cc_273 N_A1_M1017_g N_A_311_85#_c_651_n 0.012834f $X=5.26 $Y=0.795 $X2=0 $Y2=0
cc_274 N_A1_c_274_n N_A_311_85#_c_651_n 0.0599533f $X=5.28 $Y=1.515 $X2=0 $Y2=0
cc_275 N_A1_M1017_g N_A_311_85#_c_652_n 0.0014977f $X=5.26 $Y=0.795 $X2=0 $Y2=0
cc_276 N_A1_M1003_g N_VGND_c_723_n 0.00335812f $X=3.76 $Y=0.795 $X2=0 $Y2=0
cc_277 N_A1_M1017_g N_VGND_c_724_n 0.0121211f $X=5.26 $Y=0.795 $X2=0 $Y2=0
cc_278 N_A1_M1003_g N_VGND_c_725_n 0.00462669f $X=3.76 $Y=0.795 $X2=0 $Y2=0
cc_279 N_A1_M1017_g N_VGND_c_727_n 0.00447026f $X=5.26 $Y=0.795 $X2=0 $Y2=0
cc_280 N_A1_M1003_g N_VGND_c_728_n 0.00440294f $X=3.76 $Y=0.795 $X2=0 $Y2=0
cc_281 N_A1_M1017_g N_VGND_c_728_n 0.00443817f $X=5.26 $Y=0.795 $X2=0 $Y2=0
cc_282 N_A2_c_353_n N_VPWR_c_411_n 0.00278271f $X=4.305 $Y=1.765 $X2=0 $Y2=0
cc_283 N_A2_c_354_n N_VPWR_c_411_n 0.00278257f $X=4.755 $Y=1.765 $X2=0 $Y2=0
cc_284 N_A2_c_353_n N_VPWR_c_403_n 0.00354337f $X=4.305 $Y=1.765 $X2=0 $Y2=0
cc_285 N_A2_c_354_n N_VPWR_c_403_n 0.00353905f $X=4.755 $Y=1.765 $X2=0 $Y2=0
cc_286 N_A2_c_353_n N_Y_c_487_n 0.0100747f $X=4.305 $Y=1.765 $X2=0 $Y2=0
cc_287 N_A2_c_354_n N_Y_c_487_n 8.55285e-19 $X=4.755 $Y=1.765 $X2=0 $Y2=0
cc_288 N_A2_c_353_n N_Y_c_502_n 0.00453488f $X=4.305 $Y=1.765 $X2=0 $Y2=0
cc_289 N_A2_c_354_n N_Y_c_502_n 0.00107601f $X=4.755 $Y=1.765 $X2=0 $Y2=0
cc_290 N_A2_c_353_n N_A_776_368#_c_563_n 0.00951383f $X=4.305 $Y=1.765 $X2=0
+ $Y2=0
cc_291 N_A2_c_354_n N_A_776_368#_c_563_n 0.0125077f $X=4.755 $Y=1.765 $X2=0
+ $Y2=0
cc_292 N_A2_c_353_n N_A_776_368#_c_571_n 6.70277e-19 $X=4.305 $Y=1.765 $X2=0
+ $Y2=0
cc_293 N_A2_c_354_n N_A_776_368#_c_571_n 0.00778115f $X=4.755 $Y=1.765 $X2=0
+ $Y2=0
cc_294 N_A2_c_353_n N_A_776_368#_c_564_n 5.05939e-19 $X=4.305 $Y=1.765 $X2=0
+ $Y2=0
cc_295 N_A2_M1002_g N_A_311_85#_c_670_n 6.11774e-19 $X=4.29 $Y=0.795 $X2=0 $Y2=0
cc_296 N_A2_M1002_g N_A_311_85#_c_648_n 0.0176332f $X=4.29 $Y=0.795 $X2=0 $Y2=0
cc_297 N_A2_c_351_n N_A_311_85#_c_648_n 0.00251202f $X=4.51 $Y=1.515 $X2=0 $Y2=0
cc_298 N_A2_M1002_g N_A_311_85#_c_650_n 4.62671e-19 $X=4.29 $Y=0.795 $X2=0 $Y2=0
cc_299 N_A2_M1006_g N_A_311_85#_c_650_n 0.00846178f $X=4.77 $Y=0.795 $X2=0 $Y2=0
cc_300 N_A2_M1006_g N_A_311_85#_c_651_n 0.0162346f $X=4.77 $Y=0.795 $X2=0 $Y2=0
cc_301 N_A2_M1006_g N_A_311_85#_c_654_n 0.0011955f $X=4.77 $Y=0.795 $X2=0 $Y2=0
cc_302 N_A2_c_351_n N_A_311_85#_c_654_n 0.025376f $X=4.51 $Y=1.515 $X2=0 $Y2=0
cc_303 N_A2_c_352_n N_A_311_85#_c_654_n 0.00118721f $X=4.755 $Y=1.557 $X2=0
+ $Y2=0
cc_304 N_A2_M1002_g N_VGND_c_723_n 0.00231397f $X=4.29 $Y=0.795 $X2=0 $Y2=0
cc_305 N_A2_M1006_g N_VGND_c_724_n 0.0039639f $X=4.77 $Y=0.795 $X2=0 $Y2=0
cc_306 N_A2_M1002_g N_VGND_c_726_n 0.00537957f $X=4.29 $Y=0.795 $X2=0 $Y2=0
cc_307 N_A2_M1006_g N_VGND_c_726_n 0.00523995f $X=4.77 $Y=0.795 $X2=0 $Y2=0
cc_308 N_A2_M1002_g N_VGND_c_728_n 0.00528353f $X=4.29 $Y=0.795 $X2=0 $Y2=0
cc_309 N_A2_M1006_g N_VGND_c_728_n 0.00528353f $X=4.77 $Y=0.795 $X2=0 $Y2=0
cc_310 N_VPWR_M1013_s N_Y_c_487_n 0.0129983f $X=3.33 $Y=1.84 $X2=0 $Y2=0
cc_311 N_VPWR_c_406_n N_Y_c_487_n 0.0232685f $X=3.53 $Y=2.805 $X2=0 $Y2=0
cc_312 N_VPWR_M1019_s N_Y_c_477_n 0.0143738f $X=1.07 $Y=1.84 $X2=0 $Y2=0
cc_313 N_VPWR_c_412_n N_Y_c_477_n 0.0454461f $X=1.58 $Y=2.795 $X2=0 $Y2=0
cc_314 N_VPWR_c_405_n Y 0.0224263f $X=0.32 $Y=2.115 $X2=0 $Y2=0
cc_315 N_VPWR_c_405_n Y 0.0462534f $X=0.32 $Y=2.115 $X2=0 $Y2=0
cc_316 N_VPWR_c_409_n Y 0.0110241f $X=1.055 $Y=3.33 $X2=0 $Y2=0
cc_317 N_VPWR_c_412_n Y 0.024726f $X=1.58 $Y=2.795 $X2=0 $Y2=0
cc_318 N_VPWR_c_403_n Y 0.00909194f $X=5.52 $Y=3.33 $X2=0 $Y2=0
cc_319 N_VPWR_c_410_n N_A_376_368#_c_535_n 0.042287f $X=3.365 $Y=3.33 $X2=0
+ $Y2=0
cc_320 N_VPWR_c_403_n N_A_376_368#_c_535_n 0.0238254f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_321 N_VPWR_c_410_n N_A_376_368#_c_536_n 0.0227333f $X=3.365 $Y=3.33 $X2=0
+ $Y2=0
cc_322 N_VPWR_c_412_n N_A_376_368#_c_536_n 0.0219394f $X=1.58 $Y=2.795 $X2=0
+ $Y2=0
cc_323 N_VPWR_c_403_n N_A_376_368#_c_536_n 0.0125508f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_324 N_VPWR_c_406_n N_A_376_368#_c_537_n 0.0214404f $X=3.53 $Y=2.805 $X2=0
+ $Y2=0
cc_325 N_VPWR_c_410_n N_A_376_368#_c_537_n 0.0227333f $X=3.365 $Y=3.33 $X2=0
+ $Y2=0
cc_326 N_VPWR_c_403_n N_A_376_368#_c_537_n 0.0125508f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_327 N_VPWR_c_408_n N_A_776_368#_c_563_n 0.0119239f $X=5.48 $Y=2.455 $X2=0
+ $Y2=0
cc_328 N_VPWR_c_411_n N_A_776_368#_c_563_n 0.0626347f $X=5.315 $Y=3.33 $X2=0
+ $Y2=0
cc_329 N_VPWR_c_403_n N_A_776_368#_c_563_n 0.0347026f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_330 N_VPWR_c_406_n N_A_776_368#_c_564_n 0.0214404f $X=3.53 $Y=2.805 $X2=0
+ $Y2=0
cc_331 N_VPWR_c_411_n N_A_776_368#_c_564_n 0.0227333f $X=5.315 $Y=3.33 $X2=0
+ $Y2=0
cc_332 N_VPWR_c_403_n N_A_776_368#_c_564_n 0.0125508f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_333 N_Y_c_477_n N_A_376_368#_M1012_d 0.00468385f $X=2.365 $Y=2.512 $X2=-0.19
+ $Y2=-0.245
cc_334 N_Y_c_487_n N_A_376_368#_M1014_s 0.00497012f $X=4.365 $Y=2.375 $X2=0
+ $Y2=0
cc_335 N_Y_M1005_d N_A_376_368#_c_535_n 0.00214188f $X=2.365 $Y=1.84 $X2=0 $Y2=0
cc_336 N_Y_c_487_n N_A_376_368#_c_535_n 0.0041825f $X=4.365 $Y=2.375 $X2=0 $Y2=0
cc_337 N_Y_c_477_n N_A_376_368#_c_535_n 0.0046334f $X=2.365 $Y=2.512 $X2=0 $Y2=0
cc_338 N_Y_c_491_n N_A_376_368#_c_535_n 0.015762f $X=2.695 $Y=2.512 $X2=0 $Y2=0
cc_339 N_Y_c_477_n N_A_376_368#_c_536_n 0.0183658f $X=2.365 $Y=2.512 $X2=0 $Y2=0
cc_340 N_Y_c_487_n N_A_376_368#_c_537_n 0.0195451f $X=4.365 $Y=2.375 $X2=0 $Y2=0
cc_341 N_Y_c_487_n N_A_776_368#_M1000_s 0.00497922f $X=4.365 $Y=2.375 $X2=-0.19
+ $Y2=-0.245
cc_342 N_Y_M1008_d N_A_776_368#_c_563_n 0.00222494f $X=4.38 $Y=1.84 $X2=0 $Y2=0
cc_343 N_Y_c_487_n N_A_776_368#_c_563_n 0.0041825f $X=4.365 $Y=2.375 $X2=0 $Y2=0
cc_344 N_Y_c_502_n N_A_776_368#_c_563_n 0.0140094f $X=4.49 $Y=2.46 $X2=0 $Y2=0
cc_345 N_Y_c_487_n N_A_776_368#_c_571_n 0.0123817f $X=4.365 $Y=2.375 $X2=0 $Y2=0
cc_346 N_Y_c_502_n N_A_776_368#_c_571_n 0.0184049f $X=4.49 $Y=2.46 $X2=0 $Y2=0
cc_347 N_Y_c_487_n N_A_776_368#_c_564_n 0.0195451f $X=4.365 $Y=2.375 $X2=0 $Y2=0
cc_348 Y N_A_27_74#_c_593_n 0.00119776f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_349 N_Y_M1015_d N_A_27_74#_c_594_n 0.00176461f $X=0.57 $Y=0.37 $X2=0 $Y2=0
cc_350 Y N_A_27_74#_c_594_n 0.0143448f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_351 Y N_A_27_74#_c_598_n 0.00902371f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_352 N_A_27_74#_c_597_n N_A_311_85#_M1007_s 0.00343588f $X=2.045 $Y=1.095
+ $X2=-0.19 $Y2=-0.245
cc_353 N_A_27_74#_c_599_n N_A_311_85#_M1001_d 0.00184993f $X=2.895 $Y=1.095
+ $X2=0 $Y2=0
cc_354 N_A_27_74#_c_596_n N_A_311_85#_c_644_n 0.0260161f $X=1.14 $Y=0.515 $X2=0
+ $Y2=0
cc_355 N_A_27_74#_c_597_n N_A_311_85#_c_644_n 0.0198855f $X=2.045 $Y=1.095 $X2=0
+ $Y2=0
cc_356 N_A_27_74#_c_597_n N_A_311_85#_c_645_n 0.00390898f $X=2.045 $Y=1.095
+ $X2=0 $Y2=0
cc_357 N_A_27_74#_c_633_p N_A_311_85#_c_645_n 0.0127861f $X=2.13 $Y=0.885 $X2=0
+ $Y2=0
cc_358 N_A_27_74#_c_599_n N_A_311_85#_c_645_n 0.00390898f $X=2.895 $Y=1.095
+ $X2=0 $Y2=0
cc_359 N_A_27_74#_c_594_n N_A_311_85#_c_646_n 0.0128665f $X=1.055 $Y=0.34 $X2=0
+ $Y2=0
cc_360 N_A_27_74#_c_599_n N_A_311_85#_c_659_n 0.0154602f $X=2.895 $Y=1.095 $X2=0
+ $Y2=0
cc_361 N_A_27_74#_c_599_n N_A_311_85#_c_647_n 0.00376163f $X=2.895 $Y=1.095
+ $X2=0 $Y2=0
cc_362 N_A_27_74#_c_618_n N_A_311_85#_c_647_n 0.0265061f $X=3.085 $Y=0.68 $X2=0
+ $Y2=0
cc_363 N_A_27_74#_c_599_n N_A_311_85#_c_649_n 0.00749835f $X=2.895 $Y=1.095
+ $X2=0 $Y2=0
cc_364 N_A_27_74#_c_594_n N_VGND_c_725_n 0.0614387f $X=1.055 $Y=0.34 $X2=0 $Y2=0
cc_365 N_A_27_74#_c_595_n N_VGND_c_725_n 0.0179217f $X=0.365 $Y=0.34 $X2=0 $Y2=0
cc_366 N_A_27_74#_c_594_n N_VGND_c_728_n 0.0342887f $X=1.055 $Y=0.34 $X2=0 $Y2=0
cc_367 N_A_27_74#_c_595_n N_VGND_c_728_n 0.00971942f $X=0.365 $Y=0.34 $X2=0
+ $Y2=0
cc_368 N_A_311_85#_c_648_n N_VGND_M1003_d 0.00313482f $X=4.38 $Y=1.095 $X2=-0.19
+ $Y2=-0.245
cc_369 N_A_311_85#_c_651_n N_VGND_M1006_s 0.00251857f $X=5.39 $Y=1.095 $X2=0
+ $Y2=0
cc_370 N_A_311_85#_c_647_n N_VGND_c_723_n 0.0144041f $X=3.46 $Y=0.34 $X2=0 $Y2=0
cc_371 N_A_311_85#_c_648_n N_VGND_c_723_n 0.0199169f $X=4.38 $Y=1.095 $X2=0
+ $Y2=0
cc_372 N_A_311_85#_c_650_n N_VGND_c_723_n 0.00158095f $X=4.545 $Y=0.57 $X2=0
+ $Y2=0
cc_373 N_A_311_85#_c_650_n N_VGND_c_724_n 0.0163623f $X=4.545 $Y=0.57 $X2=0
+ $Y2=0
cc_374 N_A_311_85#_c_651_n N_VGND_c_724_n 0.0185548f $X=5.39 $Y=1.095 $X2=0
+ $Y2=0
cc_375 N_A_311_85#_c_652_n N_VGND_c_724_n 0.0156043f $X=5.475 $Y=0.57 $X2=0
+ $Y2=0
cc_376 N_A_311_85#_c_645_n N_VGND_c_725_n 0.0340834f $X=2.395 $Y=0.34 $X2=0
+ $Y2=0
cc_377 N_A_311_85#_c_646_n N_VGND_c_725_n 0.0233304f $X=1.865 $Y=0.34 $X2=0
+ $Y2=0
cc_378 N_A_311_85#_c_647_n N_VGND_c_725_n 0.0652108f $X=3.46 $Y=0.34 $X2=0 $Y2=0
cc_379 N_A_311_85#_c_653_n N_VGND_c_725_n 0.0233304f $X=2.56 $Y=0.34 $X2=0 $Y2=0
cc_380 N_A_311_85#_c_650_n N_VGND_c_726_n 0.0119397f $X=4.545 $Y=0.57 $X2=0
+ $Y2=0
cc_381 N_A_311_85#_c_652_n N_VGND_c_727_n 0.0092394f $X=5.475 $Y=0.57 $X2=0
+ $Y2=0
cc_382 N_A_311_85#_c_645_n N_VGND_c_728_n 0.0199188f $X=2.395 $Y=0.34 $X2=0
+ $Y2=0
cc_383 N_A_311_85#_c_646_n N_VGND_c_728_n 0.0127683f $X=1.865 $Y=0.34 $X2=0
+ $Y2=0
cc_384 N_A_311_85#_c_647_n N_VGND_c_728_n 0.0373458f $X=3.46 $Y=0.34 $X2=0 $Y2=0
cc_385 N_A_311_85#_c_650_n N_VGND_c_728_n 0.0116912f $X=4.545 $Y=0.57 $X2=0
+ $Y2=0
cc_386 N_A_311_85#_c_652_n N_VGND_c_728_n 0.0090278f $X=5.475 $Y=0.57 $X2=0
+ $Y2=0
cc_387 N_A_311_85#_c_653_n N_VGND_c_728_n 0.0127683f $X=2.56 $Y=0.34 $X2=0 $Y2=0
