* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hs__a41o_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
M1000 VPWR a_113_98# X VPB pshort w=1.12e+06u l=150000u
+  ad=2.6382e+12p pd=1.979e+07u as=6.72e+11p ps=5.68e+06u
M1001 X a_113_98# VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1002 VGND a_113_98# X VNB nlowvt w=740000u l=150000u
+  ad=1.5409e+12p pd=1.26e+07u as=4.144e+11p ps=4.08e+06u
M1003 VPWR a_113_98# X VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_1205_74# A4 VGND VNB nlowvt w=740000u l=150000u
+  ad=6.216e+11p pd=6.12e+06u as=0p ps=0u
M1005 VPWR A1 a_27_392# VPB pshort w=1e+06u l=150000u
+  ad=0p pd=0u as=2.035e+12p ps=1.607e+07u
M1006 a_27_392# B1 a_113_98# VPB pshort w=1e+06u l=150000u
+  ad=0p pd=0u as=3.5e+11p ps=2.7e+06u
M1007 a_1205_74# A3 a_1010_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=4.144e+11p ps=4.08e+06u
M1008 a_27_392# A1 VPWR VPB pshort w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 X a_113_98# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_113_98# B1 a_27_392# VPB pshort w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_751_74# A2 a_1010_74# VNB nlowvt w=740000u l=150000u
+  ad=6.216e+11p pd=6.12e+06u as=0p ps=0u
M1012 a_113_98# B1 VGND VNB nlowvt w=740000u l=150000u
+  ad=4.144e+11p pd=4.08e+06u as=0p ps=0u
M1013 a_113_98# A1 a_751_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_751_74# A1 a_113_98# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VGND A4 a_1205_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VGND a_113_98# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 VGND B1 a_113_98# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_1010_74# A3 a_1205_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VPWR A3 a_27_392# VPB pshort w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_27_392# A4 VPWR VPB pshort w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_27_392# A3 VPWR VPB pshort w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 VPWR A4 a_27_392# VPB pshort w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 X a_113_98# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 a_27_392# A2 VPWR VPB pshort w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 VPWR A2 a_27_392# VPB pshort w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 a_1010_74# A2 a_751_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 X a_113_98# VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
