* File: sky130_fd_sc_hs__nor4bb_1.pxi.spice
* Created: Thu Aug 27 20:55:29 2020
* 
x_PM_SKY130_FD_SC_HS__NOR4BB_1%C_N N_C_N_c_75_n N_C_N_M1009_g N_C_N_c_72_n
+ N_C_N_M1001_g C_N N_C_N_c_74_n PM_SKY130_FD_SC_HS__NOR4BB_1%C_N
x_PM_SKY130_FD_SC_HS__NOR4BB_1%A N_A_M1011_g N_A_c_98_n N_A_M1000_g A A
+ N_A_c_99_n PM_SKY130_FD_SC_HS__NOR4BB_1%A
x_PM_SKY130_FD_SC_HS__NOR4BB_1%B N_B_M1010_g N_B_c_132_n N_B_M1004_g B
+ N_B_c_133_n PM_SKY130_FD_SC_HS__NOR4BB_1%B
x_PM_SKY130_FD_SC_HS__NOR4BB_1%A_27_112# N_A_27_112#_M1001_s N_A_27_112#_M1009_s
+ N_A_27_112#_c_162_n N_A_27_112#_M1007_g N_A_27_112#_M1008_g
+ N_A_27_112#_c_164_n N_A_27_112#_c_168_n N_A_27_112#_c_165_n
+ N_A_27_112#_c_170_n N_A_27_112#_c_171_n N_A_27_112#_c_172_n
+ N_A_27_112#_c_173_n N_A_27_112#_c_166_n PM_SKY130_FD_SC_HS__NOR4BB_1%A_27_112#
x_PM_SKY130_FD_SC_HS__NOR4BB_1%A_611_244# N_A_611_244#_M1002_d
+ N_A_611_244#_M1003_d N_A_611_244#_M1006_g N_A_611_244#_c_259_n
+ N_A_611_244#_M1005_g N_A_611_244#_c_268_n N_A_611_244#_c_269_n
+ N_A_611_244#_c_260_n N_A_611_244#_c_261_n N_A_611_244#_c_262_n
+ N_A_611_244#_c_271_n N_A_611_244#_c_285_n N_A_611_244#_c_263_n
+ N_A_611_244#_c_264_n N_A_611_244#_c_265_n N_A_611_244#_c_266_n
+ PM_SKY130_FD_SC_HS__NOR4BB_1%A_611_244#
x_PM_SKY130_FD_SC_HS__NOR4BB_1%D_N N_D_N_c_333_n N_D_N_M1003_g N_D_N_M1002_g D_N
+ N_D_N_c_335_n PM_SKY130_FD_SC_HS__NOR4BB_1%D_N
x_PM_SKY130_FD_SC_HS__NOR4BB_1%VPWR N_VPWR_M1009_d N_VPWR_M1003_s N_VPWR_c_364_n
+ VPWR N_VPWR_c_365_n N_VPWR_c_366_n N_VPWR_c_363_n N_VPWR_c_368_n
+ N_VPWR_c_369_n N_VPWR_c_370_n PM_SKY130_FD_SC_HS__NOR4BB_1%VPWR
x_PM_SKY130_FD_SC_HS__NOR4BB_1%Y N_Y_M1011_d N_Y_M1008_d N_Y_M1006_d N_Y_c_412_n
+ N_Y_c_413_n N_Y_c_435_n N_Y_c_427_n N_Y_c_429_n N_Y_c_414_n Y N_Y_c_415_n
+ PM_SKY130_FD_SC_HS__NOR4BB_1%Y
x_PM_SKY130_FD_SC_HS__NOR4BB_1%VGND N_VGND_M1001_d N_VGND_M1010_d N_VGND_M1005_d
+ N_VGND_c_469_n N_VGND_c_470_n N_VGND_c_471_n N_VGND_c_472_n VGND
+ N_VGND_c_473_n N_VGND_c_474_n N_VGND_c_475_n N_VGND_c_476_n N_VGND_c_477_n
+ N_VGND_c_478_n PM_SKY130_FD_SC_HS__NOR4BB_1%VGND
cc_1 VNB N_C_N_c_72_n 0.0235244f $X=-0.19 $Y=-0.245 $X2=0.76 $Y2=1.22
cc_2 VNB C_N 0.00873016f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_3 VNB N_C_N_c_74_n 0.0958354f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.492
cc_4 VNB N_A_M1011_g 0.0275783f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.26
cc_5 VNB N_A_c_98_n 0.0360234f $X=-0.19 $Y=-0.245 $X2=0.76 $Y2=0.835
cc_6 VNB N_A_c_99_n 0.00391014f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.295
cc_7 VNB N_B_M1010_g 0.0292581f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.26
cc_8 VNB N_B_c_132_n 0.030975f $X=-0.19 $Y=-0.245 $X2=0.76 $Y2=0.835
cc_9 VNB N_B_c_133_n 0.00558343f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.492
cc_10 VNB N_A_27_112#_c_162_n 0.0270436f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_11 VNB N_A_27_112#_M1008_g 0.0288172f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.492
cc_12 VNB N_A_27_112#_c_164_n 0.013952f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.295
cc_13 VNB N_A_27_112#_c_165_n 0.00208657f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_27_112#_c_166_n 0.00361275f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_611_244#_c_259_n 0.0193467f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.385
cc_16 VNB N_A_611_244#_c_260_n 0.0042639f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.385
cc_17 VNB N_A_611_244#_c_261_n 0.00913271f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_611_244#_c_262_n 0.0244614f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_611_244#_c_263_n 0.0657569f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_611_244#_c_264_n 0.00488535f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_611_244#_c_265_n 0.0130414f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_611_244#_c_266_n 0.0186936f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_D_N_c_333_n 0.0212115f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.765
cc_24 VNB N_D_N_M1002_g 0.0388469f $X=-0.19 $Y=-0.245 $X2=0.76 $Y2=0.835
cc_25 VNB N_D_N_c_335_n 0.00237576f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.492
cc_26 VNB N_VPWR_c_363_n 0.203486f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_Y_c_412_n 0.00280366f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.492
cc_28 VNB N_Y_c_413_n 0.00582747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_Y_c_414_n 0.00264733f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_Y_c_415_n 0.00280529f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_469_n 0.0233407f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.492
cc_32 VNB N_VGND_c_470_n 0.0223553f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_471_n 0.0295327f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_472_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_473_n 0.0196163f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_474_n 0.0202692f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_475_n 0.284156f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_476_n 0.0185359f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_477_n 0.0209009f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_478_n 0.0148108f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VPB N_C_N_c_75_n 0.0230455f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.765
cc_42 VPB N_C_N_c_74_n 0.0101023f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.492
cc_43 VPB N_A_c_98_n 0.0338497f $X=-0.19 $Y=1.66 $X2=0.76 $Y2=0.835
cc_44 VPB N_A_c_99_n 0.0018347f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.295
cc_45 VPB N_B_c_132_n 0.0316325f $X=-0.19 $Y=1.66 $X2=0.76 $Y2=0.835
cc_46 VPB N_B_c_133_n 0.0040518f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.492
cc_47 VPB N_A_27_112#_c_162_n 0.0292215f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.21
cc_48 VPB N_A_27_112#_c_168_n 0.00395509f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_49 VPB N_A_27_112#_c_165_n 4.28226e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_50 VPB N_A_27_112#_c_170_n 0.010553f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_51 VPB N_A_27_112#_c_171_n 0.00136445f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_52 VPB N_A_27_112#_c_172_n 0.0056417f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_53 VPB N_A_27_112#_c_173_n 0.0457101f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_54 VPB N_A_27_112#_c_166_n 0.00289395f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_55 VPB N_A_611_244#_M1006_g 0.0101464f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.385
cc_56 VPB N_A_611_244#_c_268_n 0.0351197f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.295
cc_57 VPB N_A_611_244#_c_269_n 0.0131585f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_58 VPB N_A_611_244#_c_260_n 0.0754522f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.385
cc_59 VPB N_A_611_244#_c_271_n 0.0416965f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_60 VPB N_A_611_244#_c_263_n 0.006841f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_61 VPB N_A_611_244#_c_266_n 0.0210419f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_62 VPB N_D_N_c_333_n 0.0556681f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.765
cc_63 VPB N_D_N_c_335_n 0.00161194f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.492
cc_64 VPB N_VPWR_c_364_n 0.0110696f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.385
cc_65 VPB N_VPWR_c_365_n 0.0716443f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_66 VPB N_VPWR_c_366_n 0.0191515f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_67 VPB N_VPWR_c_363_n 0.0754283f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_68 VPB N_VPWR_c_368_n 0.020284f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_69 VPB N_VPWR_c_369_n 0.0297663f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_70 VPB N_VPWR_c_370_n 0.00420575f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_71 VPB N_Y_c_413_n 0.00167527f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_72 N_C_N_c_72_n N_A_M1011_g 0.0167728f $X=0.76 $Y=1.22 $X2=0 $Y2=0
cc_73 N_C_N_c_74_n N_A_c_98_n 0.0160801f $X=0.505 $Y=1.492 $X2=0 $Y2=0
cc_74 N_C_N_c_75_n N_A_c_99_n 0.00155563f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_75 N_C_N_c_74_n N_A_c_99_n 0.00112291f $X=0.505 $Y=1.492 $X2=0 $Y2=0
cc_76 N_C_N_c_72_n N_A_27_112#_c_164_n 0.00666781f $X=0.76 $Y=1.22 $X2=0 $Y2=0
cc_77 C_N N_A_27_112#_c_164_n 0.0264607f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_78 N_C_N_c_74_n N_A_27_112#_c_164_n 0.00931158f $X=0.505 $Y=1.492 $X2=0 $Y2=0
cc_79 N_C_N_c_75_n N_A_27_112#_c_168_n 7.7421e-19 $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_80 N_C_N_c_75_n N_A_27_112#_c_173_n 0.0435186f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_81 C_N N_A_27_112#_c_173_n 0.0191865f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_82 N_C_N_c_74_n N_A_27_112#_c_173_n 0.00394142f $X=0.505 $Y=1.492 $X2=0 $Y2=0
cc_83 N_C_N_c_75_n N_A_27_112#_c_166_n 0.00216635f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_84 N_C_N_c_72_n N_A_27_112#_c_166_n 0.00678818f $X=0.76 $Y=1.22 $X2=0 $Y2=0
cc_85 C_N N_A_27_112#_c_166_n 0.0267372f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_86 N_C_N_c_74_n N_A_27_112#_c_166_n 0.0290046f $X=0.505 $Y=1.492 $X2=0 $Y2=0
cc_87 N_C_N_c_75_n N_VPWR_c_363_n 0.00462577f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_88 N_C_N_c_75_n N_VPWR_c_368_n 0.00309432f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_89 N_C_N_c_72_n N_VGND_c_469_n 0.0108888f $X=0.76 $Y=1.22 $X2=0 $Y2=0
cc_90 N_C_N_c_72_n N_VGND_c_471_n 0.00390814f $X=0.76 $Y=1.22 $X2=0 $Y2=0
cc_91 N_C_N_c_72_n N_VGND_c_475_n 0.00487769f $X=0.76 $Y=1.22 $X2=0 $Y2=0
cc_92 N_A_M1011_g N_B_M1010_g 0.0212654f $X=1.395 $Y=0.74 $X2=0 $Y2=0
cc_93 N_A_c_98_n N_B_c_132_n 0.0814761f $X=1.49 $Y=1.765 $X2=0 $Y2=0
cc_94 N_A_c_98_n N_B_c_133_n 3.37032e-19 $X=1.49 $Y=1.765 $X2=0 $Y2=0
cc_95 N_A_c_98_n N_A_27_112#_c_168_n 0.0179061f $X=1.49 $Y=1.765 $X2=0 $Y2=0
cc_96 N_A_c_99_n N_A_27_112#_c_168_n 0.0119677f $X=1.24 $Y=1.515 $X2=0 $Y2=0
cc_97 N_A_c_98_n N_A_27_112#_c_173_n 3.11412e-19 $X=1.49 $Y=1.765 $X2=0 $Y2=0
cc_98 N_A_M1011_g N_A_27_112#_c_166_n 0.00110337f $X=1.395 $Y=0.74 $X2=0 $Y2=0
cc_99 N_A_c_98_n N_A_27_112#_c_166_n 0.0129014f $X=1.49 $Y=1.765 $X2=0 $Y2=0
cc_100 N_A_c_99_n N_A_27_112#_c_166_n 0.0411462f $X=1.24 $Y=1.515 $X2=0 $Y2=0
cc_101 N_A_c_99_n N_VPWR_M1009_d 0.0124807f $X=1.24 $Y=1.515 $X2=-0.19
+ $Y2=-0.245
cc_102 N_A_c_98_n N_VPWR_c_365_n 0.00322368f $X=1.49 $Y=1.765 $X2=0 $Y2=0
cc_103 N_A_c_98_n N_VPWR_c_363_n 0.00409691f $X=1.49 $Y=1.765 $X2=0 $Y2=0
cc_104 N_A_c_98_n N_VPWR_c_369_n 0.00857215f $X=1.49 $Y=1.765 $X2=0 $Y2=0
cc_105 N_A_M1011_g N_Y_c_412_n 0.00670807f $X=1.395 $Y=0.74 $X2=0 $Y2=0
cc_106 N_A_M1011_g N_Y_c_413_n 0.00508657f $X=1.395 $Y=0.74 $X2=0 $Y2=0
cc_107 N_A_c_98_n N_Y_c_413_n 0.0101944f $X=1.49 $Y=1.765 $X2=0 $Y2=0
cc_108 N_A_c_99_n N_Y_c_413_n 0.035499f $X=1.24 $Y=1.515 $X2=0 $Y2=0
cc_109 N_A_M1011_g N_Y_c_414_n 0.0041358f $X=1.395 $Y=0.74 $X2=0 $Y2=0
cc_110 N_A_c_98_n N_Y_c_414_n 0.00478726f $X=1.49 $Y=1.765 $X2=0 $Y2=0
cc_111 N_A_M1011_g N_VGND_c_469_n 0.00970997f $X=1.395 $Y=0.74 $X2=0 $Y2=0
cc_112 N_A_c_98_n N_VGND_c_469_n 0.00151797f $X=1.49 $Y=1.765 $X2=0 $Y2=0
cc_113 N_A_c_99_n N_VGND_c_469_n 0.0145292f $X=1.24 $Y=1.515 $X2=0 $Y2=0
cc_114 N_A_M1011_g N_VGND_c_475_n 0.00825771f $X=1.395 $Y=0.74 $X2=0 $Y2=0
cc_115 N_A_M1011_g N_VGND_c_476_n 0.00434272f $X=1.395 $Y=0.74 $X2=0 $Y2=0
cc_116 N_A_M1011_g N_VGND_c_477_n 4.31196e-19 $X=1.395 $Y=0.74 $X2=0 $Y2=0
cc_117 N_B_c_132_n N_A_27_112#_c_162_n 0.0509632f $X=1.91 $Y=1.765 $X2=0 $Y2=0
cc_118 N_B_c_133_n N_A_27_112#_c_162_n 0.00260445f $X=2.08 $Y=1.515 $X2=0 $Y2=0
cc_119 N_B_M1010_g N_A_27_112#_M1008_g 0.0132106f $X=1.895 $Y=0.74 $X2=0 $Y2=0
cc_120 N_B_c_132_n N_A_27_112#_c_168_n 0.0123771f $X=1.91 $Y=1.765 $X2=0 $Y2=0
cc_121 N_B_c_132_n N_A_27_112#_c_165_n 4.32175e-19 $X=1.91 $Y=1.765 $X2=0 $Y2=0
cc_122 N_B_c_133_n N_A_27_112#_c_165_n 0.0251458f $X=2.08 $Y=1.515 $X2=0 $Y2=0
cc_123 N_B_c_132_n N_A_27_112#_c_171_n 0.00143563f $X=1.91 $Y=1.765 $X2=0 $Y2=0
cc_124 N_B_c_133_n N_A_27_112#_c_171_n 0.00439118f $X=2.08 $Y=1.515 $X2=0 $Y2=0
cc_125 N_B_c_132_n N_VPWR_c_365_n 0.00322368f $X=1.91 $Y=1.765 $X2=0 $Y2=0
cc_126 N_B_c_132_n N_VPWR_c_363_n 0.00407249f $X=1.91 $Y=1.765 $X2=0 $Y2=0
cc_127 N_B_M1010_g N_Y_c_412_n 0.00282538f $X=1.895 $Y=0.74 $X2=0 $Y2=0
cc_128 N_B_M1010_g N_Y_c_413_n 0.00817586f $X=1.895 $Y=0.74 $X2=0 $Y2=0
cc_129 N_B_c_132_n N_Y_c_413_n 0.0064313f $X=1.91 $Y=1.765 $X2=0 $Y2=0
cc_130 N_B_c_133_n N_Y_c_413_n 0.0324919f $X=2.08 $Y=1.515 $X2=0 $Y2=0
cc_131 N_B_c_132_n N_Y_c_427_n 0.0221043f $X=1.91 $Y=1.765 $X2=0 $Y2=0
cc_132 N_B_c_133_n N_Y_c_427_n 0.0189046f $X=2.08 $Y=1.515 $X2=0 $Y2=0
cc_133 N_B_M1010_g N_Y_c_429_n 0.019134f $X=1.895 $Y=0.74 $X2=0 $Y2=0
cc_134 N_B_c_132_n N_Y_c_429_n 0.00155505f $X=1.91 $Y=1.765 $X2=0 $Y2=0
cc_135 N_B_c_133_n N_Y_c_429_n 0.0161271f $X=2.08 $Y=1.515 $X2=0 $Y2=0
cc_136 N_B_M1010_g N_Y_c_414_n 8.5887e-19 $X=1.895 $Y=0.74 $X2=0 $Y2=0
cc_137 N_B_M1010_g N_VGND_c_475_n 0.00753637f $X=1.895 $Y=0.74 $X2=0 $Y2=0
cc_138 N_B_M1010_g N_VGND_c_476_n 0.00383152f $X=1.895 $Y=0.74 $X2=0 $Y2=0
cc_139 N_B_M1010_g N_VGND_c_477_n 0.00911669f $X=1.895 $Y=0.74 $X2=0 $Y2=0
cc_140 N_A_27_112#_c_162_n N_A_611_244#_M1006_g 0.0387322f $X=2.575 $Y=1.765
+ $X2=0 $Y2=0
cc_141 N_A_27_112#_c_168_n N_A_611_244#_M1006_g 0.0127304f $X=3.625 $Y=2.645
+ $X2=0 $Y2=0
cc_142 N_A_27_112#_c_170_n N_A_611_244#_M1006_g 0.00751738f $X=3.625 $Y=1.805
+ $X2=0 $Y2=0
cc_143 N_A_27_112#_c_172_n N_A_611_244#_M1006_g 0.00171644f $X=3.71 $Y=2.56
+ $X2=0 $Y2=0
cc_144 N_A_27_112#_M1008_g N_A_611_244#_c_259_n 0.0198165f $X=2.74 $Y=0.74 $X2=0
+ $Y2=0
cc_145 N_A_27_112#_c_168_n N_A_611_244#_c_268_n 0.00364013f $X=3.625 $Y=2.645
+ $X2=0 $Y2=0
cc_146 N_A_27_112#_c_162_n N_A_611_244#_c_269_n 0.00222188f $X=2.575 $Y=1.765
+ $X2=0 $Y2=0
cc_147 N_A_27_112#_c_168_n N_A_611_244#_c_260_n 0.010494f $X=3.625 $Y=2.645
+ $X2=0 $Y2=0
cc_148 N_A_27_112#_c_170_n N_A_611_244#_c_260_n 0.00914877f $X=3.625 $Y=1.805
+ $X2=0 $Y2=0
cc_149 N_A_27_112#_c_172_n N_A_611_244#_c_260_n 0.0195706f $X=3.71 $Y=2.56 $X2=0
+ $Y2=0
cc_150 N_A_27_112#_c_170_n N_A_611_244#_c_261_n 0.00230969f $X=3.625 $Y=1.805
+ $X2=0 $Y2=0
cc_151 N_A_27_112#_M1008_g N_A_611_244#_c_285_n 0.00151227f $X=2.74 $Y=0.74
+ $X2=0 $Y2=0
cc_152 N_A_27_112#_c_165_n N_A_611_244#_c_285_n 0.0114575f $X=2.65 $Y=1.515
+ $X2=0 $Y2=0
cc_153 N_A_27_112#_c_170_n N_A_611_244#_c_285_n 0.0410022f $X=3.625 $Y=1.805
+ $X2=0 $Y2=0
cc_154 N_A_27_112#_c_162_n N_A_611_244#_c_263_n 0.00235515f $X=2.575 $Y=1.765
+ $X2=0 $Y2=0
cc_155 N_A_27_112#_M1008_g N_A_611_244#_c_263_n 0.0261067f $X=2.74 $Y=0.74 $X2=0
+ $Y2=0
cc_156 N_A_27_112#_c_165_n N_A_611_244#_c_263_n 0.00260664f $X=2.65 $Y=1.515
+ $X2=0 $Y2=0
cc_157 N_A_27_112#_c_170_n N_A_611_244#_c_263_n 0.0091046f $X=3.625 $Y=1.805
+ $X2=0 $Y2=0
cc_158 N_A_27_112#_c_170_n N_A_611_244#_c_264_n 0.0094058f $X=3.625 $Y=1.805
+ $X2=0 $Y2=0
cc_159 N_A_27_112#_c_170_n N_D_N_c_333_n 0.00265843f $X=3.625 $Y=1.805 $X2=-0.19
+ $Y2=-0.245
cc_160 N_A_27_112#_c_172_n N_D_N_c_333_n 0.004149f $X=3.71 $Y=2.56 $X2=-0.19
+ $Y2=-0.245
cc_161 N_A_27_112#_c_170_n N_D_N_c_335_n 0.00529505f $X=3.625 $Y=1.805 $X2=0
+ $Y2=0
cc_162 N_A_27_112#_c_168_n N_VPWR_M1009_d 0.0267619f $X=3.625 $Y=2.645 $X2=-0.19
+ $Y2=-0.245
cc_163 N_A_27_112#_c_173_n N_VPWR_M1009_d 0.0147071f $X=0.28 $Y=1.985 $X2=-0.19
+ $Y2=-0.245
cc_164 N_A_27_112#_c_168_n N_VPWR_c_364_n 0.0143758f $X=3.625 $Y=2.645 $X2=0
+ $Y2=0
cc_165 N_A_27_112#_c_172_n N_VPWR_c_364_n 0.0346722f $X=3.71 $Y=2.56 $X2=0 $Y2=0
cc_166 N_A_27_112#_c_162_n N_VPWR_c_365_n 0.00322368f $X=2.575 $Y=1.765 $X2=0
+ $Y2=0
cc_167 N_A_27_112#_c_168_n N_VPWR_c_365_n 0.0421091f $X=3.625 $Y=2.645 $X2=0
+ $Y2=0
cc_168 N_A_27_112#_c_162_n N_VPWR_c_363_n 0.00408387f $X=2.575 $Y=1.765 $X2=0
+ $Y2=0
cc_169 N_A_27_112#_c_168_n N_VPWR_c_363_n 0.069632f $X=3.625 $Y=2.645 $X2=0
+ $Y2=0
cc_170 N_A_27_112#_c_173_n N_VPWR_c_363_n 0.0171245f $X=0.28 $Y=1.985 $X2=0
+ $Y2=0
cc_171 N_A_27_112#_c_173_n N_VPWR_c_368_n 0.0112837f $X=0.28 $Y=1.985 $X2=0
+ $Y2=0
cc_172 N_A_27_112#_c_168_n N_VPWR_c_369_n 0.0427245f $X=3.625 $Y=2.645 $X2=0
+ $Y2=0
cc_173 N_A_27_112#_c_173_n N_VPWR_c_369_n 0.0103275f $X=0.28 $Y=1.985 $X2=0
+ $Y2=0
cc_174 N_A_27_112#_c_168_n A_313_368# 0.00425335f $X=3.625 $Y=2.645 $X2=-0.19
+ $Y2=-0.245
cc_175 N_A_27_112#_c_168_n A_397_368# 0.0124101f $X=3.625 $Y=2.645 $X2=-0.19
+ $Y2=-0.245
cc_176 N_A_27_112#_c_168_n A_530_368# 0.00892815f $X=3.625 $Y=2.645 $X2=-0.19
+ $Y2=-0.245
cc_177 N_A_27_112#_c_170_n A_530_368# 0.00214741f $X=3.625 $Y=1.805 $X2=-0.19
+ $Y2=-0.245
cc_178 N_A_27_112#_c_171_n A_530_368# 0.00117868f $X=2.815 $Y=1.805 $X2=-0.19
+ $Y2=-0.245
cc_179 N_A_27_112#_c_168_n N_Y_M1006_d 0.00643825f $X=3.625 $Y=2.645 $X2=0 $Y2=0
cc_180 N_A_27_112#_c_170_n N_Y_M1006_d 0.00309907f $X=3.625 $Y=1.805 $X2=0 $Y2=0
cc_181 N_A_27_112#_c_168_n N_Y_c_435_n 0.00996222f $X=3.625 $Y=2.645 $X2=0 $Y2=0
cc_182 N_A_27_112#_c_162_n N_Y_c_427_n 0.0204949f $X=2.575 $Y=1.765 $X2=0 $Y2=0
cc_183 N_A_27_112#_c_168_n N_Y_c_427_n 0.102213f $X=3.625 $Y=2.645 $X2=0 $Y2=0
cc_184 N_A_27_112#_c_170_n N_Y_c_427_n 0.0393727f $X=3.625 $Y=1.805 $X2=0 $Y2=0
cc_185 N_A_27_112#_c_171_n N_Y_c_427_n 0.0207922f $X=2.815 $Y=1.805 $X2=0 $Y2=0
cc_186 N_A_27_112#_c_172_n N_Y_c_427_n 0.0258892f $X=3.71 $Y=2.56 $X2=0 $Y2=0
cc_187 N_A_27_112#_c_162_n N_Y_c_429_n 9.45731e-19 $X=2.575 $Y=1.765 $X2=0 $Y2=0
cc_188 N_A_27_112#_M1008_g N_Y_c_429_n 0.0166532f $X=2.74 $Y=0.74 $X2=0 $Y2=0
cc_189 N_A_27_112#_c_165_n N_Y_c_429_n 0.0145929f $X=2.65 $Y=1.515 $X2=0 $Y2=0
cc_190 N_A_27_112#_c_170_n N_Y_c_429_n 0.00614593f $X=3.625 $Y=1.805 $X2=0 $Y2=0
cc_191 N_A_27_112#_M1008_g N_Y_c_415_n 0.00282724f $X=2.74 $Y=0.74 $X2=0 $Y2=0
cc_192 N_A_27_112#_c_164_n N_VGND_c_469_n 0.0271305f $X=0.605 $Y=0.845 $X2=0
+ $Y2=0
cc_193 N_A_27_112#_c_166_n N_VGND_c_469_n 0.00887541f $X=0.445 $Y=1.82 $X2=0
+ $Y2=0
cc_194 N_A_27_112#_c_164_n N_VGND_c_471_n 0.0104931f $X=0.605 $Y=0.845 $X2=0
+ $Y2=0
cc_195 N_A_27_112#_M1008_g N_VGND_c_473_n 0.00383152f $X=2.74 $Y=0.74 $X2=0
+ $Y2=0
cc_196 N_A_27_112#_M1008_g N_VGND_c_475_n 0.00753637f $X=2.74 $Y=0.74 $X2=0
+ $Y2=0
cc_197 N_A_27_112#_c_164_n N_VGND_c_475_n 0.0187574f $X=0.605 $Y=0.845 $X2=0
+ $Y2=0
cc_198 N_A_27_112#_M1008_g N_VGND_c_477_n 0.00923995f $X=2.74 $Y=0.74 $X2=0
+ $Y2=0
cc_199 N_A_611_244#_c_260_n N_D_N_c_333_n 0.0188632f $X=3.665 $Y=3.035 $X2=-0.19
+ $Y2=-0.245
cc_200 N_A_611_244#_c_261_n N_D_N_c_333_n 0.00483947f $X=4.355 $Y=1.175
+ $X2=-0.19 $Y2=-0.245
cc_201 N_A_611_244#_c_271_n N_D_N_c_333_n 0.0142271f $X=4.52 $Y=2.265 $X2=-0.19
+ $Y2=-0.245
cc_202 N_A_611_244#_c_263_n N_D_N_c_333_n 0.0150445f $X=3.575 $Y=1.385 $X2=-0.19
+ $Y2=-0.245
cc_203 N_A_611_244#_c_266_n N_D_N_c_333_n 0.00983191f $X=4.52 $Y=2.1 $X2=-0.19
+ $Y2=-0.245
cc_204 N_A_611_244#_c_261_n N_D_N_M1002_g 0.0130612f $X=4.355 $Y=1.175 $X2=0
+ $Y2=0
cc_205 N_A_611_244#_c_262_n N_D_N_M1002_g 0.0150412f $X=4.52 $Y=0.835 $X2=0
+ $Y2=0
cc_206 N_A_611_244#_c_263_n N_D_N_M1002_g 0.00455351f $X=3.575 $Y=1.385 $X2=0
+ $Y2=0
cc_207 N_A_611_244#_c_264_n N_D_N_M1002_g 0.00101533f $X=3.74 $Y=1.32 $X2=0
+ $Y2=0
cc_208 N_A_611_244#_c_265_n N_D_N_M1002_g 0.00508894f $X=4.52 $Y=1.175 $X2=0
+ $Y2=0
cc_209 N_A_611_244#_c_266_n N_D_N_M1002_g 0.0128589f $X=4.52 $Y=2.1 $X2=0 $Y2=0
cc_210 N_A_611_244#_c_261_n N_D_N_c_335_n 0.0260399f $X=4.355 $Y=1.175 $X2=0
+ $Y2=0
cc_211 N_A_611_244#_c_263_n N_D_N_c_335_n 0.00435647f $X=3.575 $Y=1.385 $X2=0
+ $Y2=0
cc_212 N_A_611_244#_c_264_n N_D_N_c_335_n 0.00674841f $X=3.74 $Y=1.32 $X2=0
+ $Y2=0
cc_213 N_A_611_244#_c_266_n N_D_N_c_335_n 0.0250404f $X=4.52 $Y=2.1 $X2=0 $Y2=0
cc_214 N_A_611_244#_c_260_n N_VPWR_c_364_n 0.0129397f $X=3.665 $Y=3.035 $X2=0
+ $Y2=0
cc_215 N_A_611_244#_c_271_n N_VPWR_c_364_n 0.034469f $X=4.52 $Y=2.265 $X2=0
+ $Y2=0
cc_216 N_A_611_244#_c_269_n N_VPWR_c_365_n 0.0169667f $X=3.22 $Y=3.11 $X2=0
+ $Y2=0
cc_217 N_A_611_244#_c_271_n N_VPWR_c_366_n 0.0145938f $X=4.52 $Y=2.265 $X2=0
+ $Y2=0
cc_218 N_A_611_244#_c_268_n N_VPWR_c_363_n 0.0160334f $X=3.59 $Y=3.11 $X2=0
+ $Y2=0
cc_219 N_A_611_244#_c_269_n N_VPWR_c_363_n 0.0063013f $X=3.22 $Y=3.11 $X2=0
+ $Y2=0
cc_220 N_A_611_244#_c_271_n N_VPWR_c_363_n 0.0120466f $X=4.52 $Y=2.265 $X2=0
+ $Y2=0
cc_221 N_A_611_244#_M1006_g N_Y_c_427_n 0.0139841f $X=3.145 $Y=2.4 $X2=0 $Y2=0
cc_222 N_A_611_244#_c_260_n N_Y_c_427_n 0.00257284f $X=3.665 $Y=3.035 $X2=0
+ $Y2=0
cc_223 N_A_611_244#_c_259_n N_Y_c_429_n 0.00812308f $X=3.24 $Y=1.22 $X2=0 $Y2=0
cc_224 N_A_611_244#_c_285_n N_Y_c_429_n 0.0108526f $X=3.575 $Y=1.385 $X2=0 $Y2=0
cc_225 N_A_611_244#_c_263_n N_Y_c_429_n 0.00290188f $X=3.575 $Y=1.385 $X2=0
+ $Y2=0
cc_226 N_A_611_244#_c_259_n N_Y_c_415_n 0.00814444f $X=3.24 $Y=1.22 $X2=0 $Y2=0
cc_227 N_A_611_244#_c_261_n N_VGND_M1005_d 0.00472896f $X=4.355 $Y=1.175 $X2=0
+ $Y2=0
cc_228 N_A_611_244#_c_264_n N_VGND_M1005_d 0.00214094f $X=3.74 $Y=1.32 $X2=0
+ $Y2=0
cc_229 N_A_611_244#_c_259_n N_VGND_c_470_n 0.0174322f $X=3.24 $Y=1.22 $X2=0
+ $Y2=0
cc_230 N_A_611_244#_c_262_n N_VGND_c_470_n 0.0144669f $X=4.52 $Y=0.835 $X2=0
+ $Y2=0
cc_231 N_A_611_244#_c_285_n N_VGND_c_470_n 0.00873167f $X=3.575 $Y=1.385 $X2=0
+ $Y2=0
cc_232 N_A_611_244#_c_263_n N_VGND_c_470_n 0.00475493f $X=3.575 $Y=1.385 $X2=0
+ $Y2=0
cc_233 N_A_611_244#_c_264_n N_VGND_c_470_n 0.0500172f $X=3.74 $Y=1.32 $X2=0
+ $Y2=0
cc_234 N_A_611_244#_c_259_n N_VGND_c_473_n 0.00383287f $X=3.24 $Y=1.22 $X2=0
+ $Y2=0
cc_235 N_A_611_244#_c_262_n N_VGND_c_474_n 0.00816527f $X=4.52 $Y=0.835 $X2=0
+ $Y2=0
cc_236 N_A_611_244#_c_259_n N_VGND_c_475_n 0.00661688f $X=3.24 $Y=1.22 $X2=0
+ $Y2=0
cc_237 N_A_611_244#_c_262_n N_VGND_c_475_n 0.0106525f $X=4.52 $Y=0.835 $X2=0
+ $Y2=0
cc_238 N_A_611_244#_c_259_n N_VGND_c_477_n 6.14575e-19 $X=3.24 $Y=1.22 $X2=0
+ $Y2=0
cc_239 N_D_N_c_333_n N_VPWR_c_364_n 0.0081869f $X=4.295 $Y=2.045 $X2=0 $Y2=0
cc_240 N_D_N_c_335_n N_VPWR_c_364_n 0.0116968f $X=4.18 $Y=1.615 $X2=0 $Y2=0
cc_241 N_D_N_c_333_n N_VPWR_c_366_n 0.00445602f $X=4.295 $Y=2.045 $X2=0 $Y2=0
cc_242 N_D_N_c_333_n N_VPWR_c_363_n 0.00861878f $X=4.295 $Y=2.045 $X2=0 $Y2=0
cc_243 N_D_N_M1002_g N_VGND_c_470_n 0.0124771f $X=4.305 $Y=0.835 $X2=0 $Y2=0
cc_244 N_D_N_M1002_g N_VGND_c_474_n 0.0043356f $X=4.305 $Y=0.835 $X2=0 $Y2=0
cc_245 N_D_N_M1002_g N_VGND_c_475_n 0.00487769f $X=4.305 $Y=0.835 $X2=0 $Y2=0
cc_246 A_313_368# N_Y_c_413_n 0.00264145f $X=1.565 $Y=1.84 $X2=0.545 $Y2=0.845
cc_247 A_313_368# N_Y_c_435_n 0.00193973f $X=1.565 $Y=1.84 $X2=0.545 $Y2=0.845
cc_248 A_313_368# N_Y_c_427_n 0.00167087f $X=1.565 $Y=1.84 $X2=0.69 $Y2=1.82
cc_249 A_397_368# N_Y_c_427_n 0.0168674f $X=1.985 $Y=1.84 $X2=0.69 $Y2=1.82
cc_250 A_530_368# N_Y_c_427_n 0.00756005f $X=2.65 $Y=1.84 $X2=0.69 $Y2=1.82
cc_251 N_Y_c_429_n N_VGND_M1010_d 0.0220163f $X=2.86 $Y=0.965 $X2=0 $Y2=0
cc_252 N_Y_c_412_n N_VGND_c_469_n 0.0206398f $X=1.61 $Y=0.515 $X2=0 $Y2=0
cc_253 N_Y_c_414_n N_VGND_c_469_n 0.0109738f $X=1.61 $Y=0.965 $X2=0 $Y2=0
cc_254 N_Y_c_429_n N_VGND_c_470_n 0.00348012f $X=2.86 $Y=0.965 $X2=0 $Y2=0
cc_255 N_Y_c_415_n N_VGND_c_470_n 0.0439579f $X=3.025 $Y=0.515 $X2=0 $Y2=0
cc_256 N_Y_c_415_n N_VGND_c_473_n 0.0164719f $X=3.025 $Y=0.515 $X2=0 $Y2=0
cc_257 N_Y_c_412_n N_VGND_c_475_n 0.0119984f $X=1.61 $Y=0.515 $X2=0 $Y2=0
cc_258 N_Y_c_415_n N_VGND_c_475_n 0.013457f $X=3.025 $Y=0.515 $X2=0 $Y2=0
cc_259 N_Y_c_412_n N_VGND_c_476_n 0.0145639f $X=1.61 $Y=0.515 $X2=0 $Y2=0
cc_260 N_Y_c_412_n N_VGND_c_477_n 0.0146527f $X=1.61 $Y=0.515 $X2=0 $Y2=0
cc_261 N_Y_c_429_n N_VGND_c_477_n 0.0449771f $X=2.86 $Y=0.965 $X2=0 $Y2=0
cc_262 N_Y_c_415_n N_VGND_c_477_n 0.0146682f $X=3.025 $Y=0.515 $X2=0 $Y2=0
