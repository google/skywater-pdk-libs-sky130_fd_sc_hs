* File: sky130_fd_sc_hs__nand4b_2.pex.spice
* Created: Tue Sep  1 20:10:13 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HS__NAND4B_2%A_N 3 6 7 9 10 11 18 19
c33 18 0 1.48501e-19 $X=0.82 $Y=1.345
r34 17 19 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=0.82 $Y=1.345
+ $X2=0.895 $Y2=1.345
r35 17 18 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.82
+ $Y=1.345 $X2=0.82 $Y2=1.345
r36 14 17 56.8299 $w=3.3e-07 $l=3.25e-07 $layer=POLY_cond $X=0.495 $Y=1.345
+ $X2=0.82 $Y2=1.345
r37 11 18 3.49225 $w=3.28e-07 $l=1e-07 $layer=LI1_cond $X=0.72 $Y=1.345 $X2=0.82
+ $Y2=1.345
r38 10 11 16.7628 $w=3.28e-07 $l=4.8e-07 $layer=LI1_cond $X=0.24 $Y=1.345
+ $X2=0.72 $Y2=1.345
r39 7 9 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=0.895 $Y=1.765
+ $X2=0.895 $Y2=2.34
r40 6 7 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=0.895 $Y=1.675 $X2=0.895
+ $Y2=1.765
r41 5 19 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=0.895 $Y=1.51
+ $X2=0.895 $Y2=1.345
r42 5 6 64.1371 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=0.895 $Y=1.51
+ $X2=0.895 $Y2=1.675
r43 1 14 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.495 $Y=1.18
+ $X2=0.495 $Y2=1.345
r44 1 3 251.255 $w=1.5e-07 $l=4.9e-07 $layer=POLY_cond $X=0.495 $Y=1.18
+ $X2=0.495 $Y2=0.69
.ends

.subckt PM_SKY130_FD_SC_HS__NAND4B_2%A_27_74# 1 2 7 9 12 14 16 19 23 25 26 29 33
+ 34 36 38 44
c86 44 0 1.48501e-19 $X=1.885 $Y=1.557
c87 19 0 9.65687e-20 $X=1.945 $Y=0.74
c88 12 0 4.22696e-20 $X=1.485 $Y=0.74
r89 44 45 7.712 $w=3.75e-07 $l=6e-08 $layer=POLY_cond $X=1.885 $Y=1.557
+ $X2=1.945 $Y2=1.557
r90 41 42 6.42667 $w=3.75e-07 $l=5e-08 $layer=POLY_cond $X=1.435 $Y=1.557
+ $X2=1.485 $Y2=1.557
r91 39 44 42.416 $w=3.75e-07 $l=3.3e-07 $layer=POLY_cond $X=1.555 $Y=1.557
+ $X2=1.885 $Y2=1.557
r92 39 42 8.99733 $w=3.75e-07 $l=7e-08 $layer=POLY_cond $X=1.555 $Y=1.557
+ $X2=1.485 $Y2=1.557
r93 38 39 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.555
+ $Y=1.515 $X2=1.555 $Y2=1.515
r94 36 38 9.29987 $w=4.3e-07 $l=2.67047e-07 $layer=LI1_cond $X=1.24 $Y=1.35
+ $X2=1.437 $Y2=1.515
r95 35 36 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=1.24 $Y=1.01
+ $X2=1.24 $Y2=1.35
r96 33 38 7.09302 $w=4.3e-07 $l=3.87329e-07 $layer=LI1_cond $X=1.155 $Y=1.765
+ $X2=1.437 $Y2=1.515
r97 33 34 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=1.155 $Y=1.765
+ $X2=0.835 $Y2=1.765
r98 29 31 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=0.67 $Y=1.985
+ $X2=0.67 $Y2=2.695
r99 27 34 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.67 $Y=1.85
+ $X2=0.835 $Y2=1.765
r100 27 29 4.71454 $w=3.28e-07 $l=1.35e-07 $layer=LI1_cond $X=0.67 $Y=1.85
+ $X2=0.67 $Y2=1.985
r101 25 35 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.155 $Y=0.925
+ $X2=1.24 $Y2=1.01
r102 25 26 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=1.155 $Y=0.925
+ $X2=0.365 $Y2=0.925
r103 21 26 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.24 $Y=0.84
+ $X2=0.365 $Y2=0.925
r104 21 23 7.37564 $w=2.48e-07 $l=1.6e-07 $layer=LI1_cond $X=0.24 $Y=0.84
+ $X2=0.24 $Y2=0.68
r105 17 45 24.2915 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.945 $Y=1.35
+ $X2=1.945 $Y2=1.557
r106 17 19 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.945 $Y=1.35
+ $X2=1.945 $Y2=0.74
r107 14 44 24.2915 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=1.885 $Y=1.765
+ $X2=1.885 $Y2=1.557
r108 14 16 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.885 $Y=1.765
+ $X2=1.885 $Y2=2.4
r109 10 42 24.2915 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.485 $Y=1.35
+ $X2=1.485 $Y2=1.557
r110 10 12 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.485 $Y=1.35
+ $X2=1.485 $Y2=0.74
r111 7 41 24.2915 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=1.435 $Y=1.765
+ $X2=1.435 $Y2=1.557
r112 7 9 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.435 $Y=1.765
+ $X2=1.435 $Y2=2.4
r113 2 31 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=0.525
+ $Y=1.84 $X2=0.67 $Y2=2.695
r114 2 29 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.525
+ $Y=1.84 $X2=0.67 $Y2=1.985
r115 1 23 182 $w=1.7e-07 $l=3.75566e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.68
.ends

.subckt PM_SKY130_FD_SC_HS__NAND4B_2%B 3 5 7 10 12 14 15 20 22
c59 12 0 6.34043e-20 $X=3.15 $Y=1.765
c60 3 0 3.91537e-20 $X=2.375 $Y=0.74
r61 22 23 24.7008 $w=3.61e-07 $l=1.85e-07 $layer=POLY_cond $X=2.965 $Y=1.557
+ $X2=3.15 $Y2=1.557
r62 21 22 35.3823 $w=3.61e-07 $l=2.65e-07 $layer=POLY_cond $X=2.7 $Y=1.557
+ $X2=2.965 $Y2=1.557
r63 19 21 36.7175 $w=3.61e-07 $l=2.75e-07 $layer=POLY_cond $X=2.425 $Y=1.557
+ $X2=2.7 $Y2=1.557
r64 19 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.425
+ $Y=1.515 $X2=2.425 $Y2=1.515
r65 17 19 6.6759 $w=3.61e-07 $l=5e-08 $layer=POLY_cond $X=2.375 $Y=1.557
+ $X2=2.425 $Y2=1.557
r66 15 20 7.10226 $w=4.28e-07 $l=2.65e-07 $layer=LI1_cond $X=2.16 $Y=1.565
+ $X2=2.425 $Y2=1.565
r67 12 23 23.3725 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=3.15 $Y=1.765
+ $X2=3.15 $Y2=1.557
r68 12 14 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.15 $Y=1.765
+ $X2=3.15 $Y2=2.4
r69 8 22 23.3725 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.965 $Y=1.35
+ $X2=2.965 $Y2=1.557
r70 8 10 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.965 $Y=1.35
+ $X2=2.965 $Y2=0.74
r71 5 21 23.3725 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=2.7 $Y=1.765 $X2=2.7
+ $Y2=1.557
r72 5 7 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.7 $Y=1.765 $X2=2.7
+ $Y2=2.4
r73 1 17 23.3725 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.375 $Y=1.35
+ $X2=2.375 $Y2=1.557
r74 1 3 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.375 $Y=1.35
+ $X2=2.375 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HS__NAND4B_2%C 1 3 6 8 10 13 15 16 24
c57 16 0 6.34043e-20 $X=4.08 $Y=1.665
c58 8 0 1.20111e-19 $X=4.15 $Y=1.765
r59 22 24 18.075 $w=3.2e-07 $l=1.2e-07 $layer=POLY_cond $X=4.03 $Y=1.557
+ $X2=4.15 $Y2=1.557
r60 22 23 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.03
+ $Y=1.515 $X2=4.03 $Y2=1.515
r61 20 22 11.2969 $w=3.2e-07 $l=7.5e-08 $layer=POLY_cond $X=3.955 $Y=1.557
+ $X2=4.03 $Y2=1.557
r62 19 20 38.4094 $w=3.2e-07 $l=2.55e-07 $layer=POLY_cond $X=3.7 $Y=1.557
+ $X2=3.955 $Y2=1.557
r63 16 23 1.34005 $w=4.28e-07 $l=5e-08 $layer=LI1_cond $X=4.08 $Y=1.565 $X2=4.03
+ $Y2=1.565
r64 15 23 11.5244 $w=4.28e-07 $l=4.3e-07 $layer=LI1_cond $X=3.6 $Y=1.565
+ $X2=4.03 $Y2=1.565
r65 11 24 35.3969 $w=3.2e-07 $l=3.22289e-07 $layer=POLY_cond $X=4.385 $Y=1.35
+ $X2=4.15 $Y2=1.557
r66 11 13 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=4.385 $Y=1.35
+ $X2=4.385 $Y2=0.79
r67 8 24 20.4921 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=4.15 $Y=1.765
+ $X2=4.15 $Y2=1.557
r68 8 10 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=4.15 $Y=1.765
+ $X2=4.15 $Y2=2.4
r69 4 20 20.4921 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.955 $Y=1.35
+ $X2=3.955 $Y2=1.557
r70 4 6 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=3.955 $Y=1.35
+ $X2=3.955 $Y2=0.79
r71 1 19 20.4921 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=3.7 $Y=1.765 $X2=3.7
+ $Y2=1.557
r72 1 3 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.7 $Y=1.765 $X2=3.7
+ $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_HS__NAND4B_2%D 1 3 6 8 10 13 15 16 17 26
c46 17 0 1.20111e-19 $X=5.52 $Y=1.665
r47 26 27 1.95935 $w=3.69e-07 $l=1.5e-08 $layer=POLY_cond $X=5.25 $Y=1.557
+ $X2=5.265 $Y2=1.557
r48 24 26 45.065 $w=3.69e-07 $l=3.45e-07 $layer=POLY_cond $X=4.905 $Y=1.557
+ $X2=5.25 $Y2=1.557
r49 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.905
+ $Y=1.515 $X2=4.905 $Y2=1.515
r50 22 24 11.7561 $w=3.69e-07 $l=9e-08 $layer=POLY_cond $X=4.815 $Y=1.557
+ $X2=4.905 $Y2=1.557
r51 21 22 1.95935 $w=3.69e-07 $l=1.5e-08 $layer=POLY_cond $X=4.8 $Y=1.557
+ $X2=4.815 $Y2=1.557
r52 16 17 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=5.04 $Y=1.565
+ $X2=5.52 $Y2=1.565
r53 16 25 3.61813 $w=4.28e-07 $l=1.35e-07 $layer=LI1_cond $X=5.04 $Y=1.565
+ $X2=4.905 $Y2=1.565
r54 15 25 9.24634 $w=4.28e-07 $l=3.45e-07 $layer=LI1_cond $X=4.56 $Y=1.565
+ $X2=4.905 $Y2=1.565
r55 11 27 23.9013 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=5.265 $Y=1.35
+ $X2=5.265 $Y2=1.557
r56 11 13 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=5.265 $Y=1.35
+ $X2=5.265 $Y2=0.79
r57 8 26 23.9013 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=5.25 $Y=1.765
+ $X2=5.25 $Y2=1.557
r58 8 10 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=5.25 $Y=1.765
+ $X2=5.25 $Y2=2.4
r59 4 22 23.9013 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.815 $Y=1.35
+ $X2=4.815 $Y2=1.557
r60 4 6 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=4.815 $Y=1.35
+ $X2=4.815 $Y2=0.79
r61 1 21 23.9013 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=4.8 $Y=1.765 $X2=4.8
+ $Y2=1.557
r62 1 3 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=4.8 $Y=1.765 $X2=4.8
+ $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_HS__NAND4B_2%VPWR 1 2 3 4 5 18 24 28 32 34 36 41 42 43
+ 45 50 59 63 69 72 75 79
r75 78 79 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r76 75 76 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r77 72 73 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r78 69 70 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r79 67 79 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=5.52 $Y2=3.33
r80 67 76 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=4.56 $Y2=3.33
r81 66 67 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r82 64 75 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.65 $Y=3.33
+ $X2=4.485 $Y2=3.33
r83 64 66 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=4.65 $Y=3.33
+ $X2=5.04 $Y2=3.33
r84 63 78 4.31409 $w=1.7e-07 $l=2e-07 $layer=LI1_cond $X=5.36 $Y=3.33 $X2=5.56
+ $Y2=3.33
r85 63 66 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=5.36 $Y=3.33 $X2=5.04
+ $Y2=3.33
r86 62 76 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=4.56 $Y2=3.33
r87 61 62 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r88 59 75 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.32 $Y=3.33
+ $X2=4.485 $Y2=3.33
r89 59 61 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=4.32 $Y=3.33
+ $X2=4.08 $Y2=3.33
r90 58 62 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=4.08 $Y2=3.33
r91 57 58 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r92 55 72 12.4999 $w=1.7e-07 $l=2.98e-07 $layer=LI1_cond $X=2.59 $Y=3.33
+ $X2=2.292 $Y2=3.33
r93 55 57 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=2.59 $Y=3.33
+ $X2=3.12 $Y2=3.33
r94 54 73 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r95 54 70 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r96 53 54 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r97 51 69 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.37 $Y=3.33
+ $X2=1.205 $Y2=3.33
r98 51 53 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=1.37 $Y=3.33
+ $X2=1.68 $Y2=3.33
r99 50 72 12.4999 $w=1.7e-07 $l=2.97e-07 $layer=LI1_cond $X=1.995 $Y=3.33
+ $X2=2.292 $Y2=3.33
r100 50 53 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=1.995 $Y=3.33
+ $X2=1.68 $Y2=3.33
r101 48 70 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r102 47 48 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r103 45 69 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.04 $Y=3.33
+ $X2=1.205 $Y2=3.33
r104 45 47 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=1.04 $Y=3.33
+ $X2=0.72 $Y2=3.33
r105 43 58 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.88 $Y=3.33
+ $X2=3.12 $Y2=3.33
r106 43 73 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=2.88 $Y=3.33
+ $X2=2.16 $Y2=3.33
r107 41 57 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=3.26 $Y=3.33
+ $X2=3.12 $Y2=3.33
r108 41 42 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.26 $Y=3.33
+ $X2=3.425 $Y2=3.33
r109 40 61 31.9679 $w=1.68e-07 $l=4.9e-07 $layer=LI1_cond $X=3.59 $Y=3.33
+ $X2=4.08 $Y2=3.33
r110 40 42 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.59 $Y=3.33
+ $X2=3.425 $Y2=3.33
r111 36 39 28.3056 $w=2.83e-07 $l=7e-07 $layer=LI1_cond $X=5.502 $Y=2.115
+ $X2=5.502 $Y2=2.815
r112 34 78 3.08458 $w=2.85e-07 $l=1.1025e-07 $layer=LI1_cond $X=5.502 $Y=3.245
+ $X2=5.56 $Y2=3.33
r113 34 39 17.3877 $w=2.83e-07 $l=4.3e-07 $layer=LI1_cond $X=5.502 $Y=3.245
+ $X2=5.502 $Y2=2.815
r114 30 75 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.485 $Y=3.245
+ $X2=4.485 $Y2=3.33
r115 30 32 29.1603 $w=3.28e-07 $l=8.35e-07 $layer=LI1_cond $X=4.485 $Y=3.245
+ $X2=4.485 $Y2=2.41
r116 26 42 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.425 $Y=3.245
+ $X2=3.425 $Y2=3.33
r117 26 28 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=3.425 $Y=3.245
+ $X2=3.425 $Y2=2.415
r118 22 72 2.50116 $w=5.95e-07 $l=8.5e-08 $layer=LI1_cond $X=2.292 $Y=3.245
+ $X2=2.292 $Y2=3.33
r119 22 24 15.8807 $w=5.93e-07 $l=7.9e-07 $layer=LI1_cond $X=2.292 $Y=3.245
+ $X2=2.292 $Y2=2.455
r120 18 21 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=1.205 $Y=2.105
+ $X2=1.205 $Y2=2.785
r121 16 69 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.205 $Y=3.245
+ $X2=1.205 $Y2=3.33
r122 16 21 16.0644 $w=3.28e-07 $l=4.6e-07 $layer=LI1_cond $X=1.205 $Y=3.245
+ $X2=1.205 $Y2=2.785
r123 5 39 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=5.325
+ $Y=1.84 $X2=5.475 $Y2=2.815
r124 5 36 400 $w=1.7e-07 $l=3.4187e-07 $layer=licon1_PDIFF $count=1 $X=5.325
+ $Y=1.84 $X2=5.475 $Y2=2.115
r125 4 32 300 $w=1.7e-07 $l=6.87823e-07 $layer=licon1_PDIFF $count=2 $X=4.225
+ $Y=1.84 $X2=4.485 $Y2=2.41
r126 3 28 300 $w=1.7e-07 $l=6.67552e-07 $layer=licon1_PDIFF $count=2 $X=3.225
+ $Y=1.84 $X2=3.425 $Y2=2.415
r127 2 24 150 $w=1.7e-07 $l=8.33637e-07 $layer=licon1_PDIFF $count=4 $X=1.96
+ $Y=1.84 $X2=2.475 $Y2=2.455
r128 1 21 600 $w=1.7e-07 $l=1.05598e-06 $layer=licon1_PDIFF $count=1 $X=0.97
+ $Y=1.84 $X2=1.205 $Y2=2.785
r129 1 18 300 $w=1.7e-07 $l=3.64005e-07 $layer=licon1_PDIFF $count=2 $X=0.97
+ $Y=1.84 $X2=1.205 $Y2=2.105
.ends

.subckt PM_SKY130_FD_SC_HS__NAND4B_2%Y 1 2 3 4 5 16 18 20 22 26 28 32 34 36 38
+ 41 49 55 58 59
c102 22 0 4.22696e-20 $X=3.005 $Y=1.095
r103 58 59 18.5393 $w=2.28e-07 $l=3.7e-07 $layer=LI1_cond $X=3.12 $Y=1.295
+ $X2=3.12 $Y2=1.665
r104 53 58 5.76222 $w=2.28e-07 $l=1.15e-07 $layer=LI1_cond $X=3.12 $Y=1.18
+ $X2=3.12 $Y2=1.295
r105 50 59 7.76646 $w=2.28e-07 $l=1.55e-07 $layer=LI1_cond $X=3.12 $Y=1.82
+ $X2=3.12 $Y2=1.665
r106 49 50 7.34574 $w=4.73e-07 $l=1.65e-07 $layer=LI1_cond $X=2.997 $Y=1.985
+ $X2=2.997 $Y2=1.82
r107 41 43 4.1616 $w=3.58e-07 $l=1.3e-07 $layer=LI1_cond $X=1.715 $Y=0.965
+ $X2=1.715 $Y2=1.095
r108 36 57 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.025 $Y=2.12
+ $X2=5.025 $Y2=2.035
r109 36 38 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=5.025 $Y=2.12
+ $X2=5.025 $Y2=2.815
r110 35 55 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.09 $Y=2.035
+ $X2=3.925 $Y2=2.035
r111 34 57 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.86 $Y=2.035
+ $X2=5.025 $Y2=2.035
r112 34 35 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=4.86 $Y=2.035
+ $X2=4.09 $Y2=2.035
r113 30 55 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.925 $Y=2.12
+ $X2=3.925 $Y2=2.035
r114 30 32 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=3.925 $Y=2.12
+ $X2=3.925 $Y2=2.815
r115 28 55 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.76 $Y=2.035
+ $X2=3.925 $Y2=2.035
r116 28 29 34.2513 $w=1.68e-07 $l=5.25e-07 $layer=LI1_cond $X=3.76 $Y=2.035
+ $X2=3.235 $Y2=2.035
r117 26 52 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=2.925 $Y=2.815
+ $X2=2.925 $Y2=2.12
r118 23 43 5.14255 $w=1.7e-07 $l=1.8e-07 $layer=LI1_cond $X=1.895 $Y=1.095
+ $X2=1.715 $Y2=1.095
r119 22 53 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=3.005 $Y=1.095
+ $X2=3.12 $Y2=1.18
r120 22 23 72.4171 $w=1.68e-07 $l=1.11e-06 $layer=LI1_cond $X=3.005 $Y=1.095
+ $X2=1.895 $Y2=1.095
r121 21 46 4.26175 $w=1.7e-07 $l=1.61071e-07 $layer=LI1_cond $X=1.825 $Y=2.035
+ $X2=1.687 $Y2=1.985
r122 20 52 3.26684 $w=4.73e-07 $l=8.5e-08 $layer=LI1_cond $X=2.997 $Y=2.035
+ $X2=2.997 $Y2=2.12
r123 20 29 6.83586 $w=1.7e-07 $l=2.38e-07 $layer=LI1_cond $X=2.997 $Y=2.035
+ $X2=3.235 $Y2=2.035
r124 20 49 1.25903 $w=4.73e-07 $l=5e-08 $layer=LI1_cond $X=2.997 $Y=2.035
+ $X2=2.997 $Y2=1.985
r125 20 21 61 $w=1.68e-07 $l=9.35e-07 $layer=LI1_cond $X=2.76 $Y=2.035 $X2=1.825
+ $Y2=2.035
r126 16 46 3.0603 $w=2.75e-07 $l=1.35e-07 $layer=LI1_cond $X=1.687 $Y=2.12
+ $X2=1.687 $Y2=1.985
r127 16 18 29.1254 $w=2.73e-07 $l=6.95e-07 $layer=LI1_cond $X=1.687 $Y=2.12
+ $X2=1.687 $Y2=2.815
r128 5 57 400 $w=1.7e-07 $l=2.59374e-07 $layer=licon1_PDIFF $count=1 $X=4.875
+ $Y=1.84 $X2=5.025 $Y2=2.035
r129 5 38 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=4.875
+ $Y=1.84 $X2=5.025 $Y2=2.815
r130 4 55 400 $w=1.7e-07 $l=2.59374e-07 $layer=licon1_PDIFF $count=1 $X=3.775
+ $Y=1.84 $X2=3.925 $Y2=2.035
r131 4 32 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=3.775
+ $Y=1.84 $X2=3.925 $Y2=2.815
r132 3 49 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=2.775
+ $Y=1.84 $X2=2.925 $Y2=1.985
r133 3 26 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=2.775
+ $Y=1.84 $X2=2.925 $Y2=2.815
r134 2 46 400 $w=1.7e-07 $l=2.38485e-07 $layer=licon1_PDIFF $count=1 $X=1.51
+ $Y=1.84 $X2=1.66 $Y2=2.015
r135 2 18 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=1.51
+ $Y=1.84 $X2=1.66 $Y2=2.815
r136 1 41 182 $w=1.7e-07 $l=6.68019e-07 $layer=licon1_NDIFF $count=1 $X=1.56
+ $Y=0.37 $X2=1.715 $Y2=0.965
.ends

.subckt PM_SKY130_FD_SC_HS__NAND4B_2%VGND 1 2 9 13 15 17 22 32 33 36 39
r56 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r57 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r58 33 40 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=5.04
+ $Y2=0
r59 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r60 30 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.195 $Y=0 $X2=5.03
+ $Y2=0
r61 30 32 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=5.195 $Y=0 $X2=5.52
+ $Y2=0
r62 29 40 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=5.04
+ $Y2=0
r63 28 29 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r64 26 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r65 25 28 219.209 $w=1.68e-07 $l=3.36e-06 $layer=LI1_cond $X=1.2 $Y=0 $X2=4.56
+ $Y2=0
r66 25 26 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r67 23 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.875 $Y=0 $X2=0.71
+ $Y2=0
r68 23 25 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.875 $Y=0 $X2=1.2
+ $Y2=0
r69 22 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.865 $Y=0 $X2=5.03
+ $Y2=0
r70 22 28 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=4.865 $Y=0 $X2=4.56
+ $Y2=0
r71 20 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r72 19 20 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r73 17 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.545 $Y=0 $X2=0.71
+ $Y2=0
r74 17 19 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.545 $Y=0 $X2=0.24
+ $Y2=0
r75 15 29 0.468274 $w=4.9e-07 $l=1.68e-06 $layer=MET1_cond $X=2.88 $Y=0 $X2=4.56
+ $Y2=0
r76 15 26 0.468274 $w=4.9e-07 $l=1.68e-06 $layer=MET1_cond $X=2.88 $Y=0 $X2=1.2
+ $Y2=0
r77 11 39 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.03 $Y=0.085
+ $X2=5.03 $Y2=0
r78 11 13 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=5.03 $Y=0.085
+ $X2=5.03 $Y2=0.58
r79 7 36 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.71 $Y=0.085 $X2=0.71
+ $Y2=0
r80 7 9 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=0.71 $Y=0.085 $X2=0.71
+ $Y2=0.55
r81 2 13 182 $w=1.7e-07 $l=2.19089e-07 $layer=licon1_NDIFF $count=1 $X=4.89
+ $Y=0.42 $X2=5.03 $Y2=0.58
r82 1 9 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=0.57 $Y=0.37
+ $X2=0.71 $Y2=0.55
.ends

.subckt PM_SKY130_FD_SC_HS__NAND4B_2%A_225_74# 1 2 3 10 16 23 24
c37 16 0 9.65687e-20 $X=2.2 $Y=0.49
c38 10 0 3.91537e-20 $X=2.075 $Y=0.49
r39 23 24 8.85254 $w=2.43e-07 $l=1.65e-07 $layer=LI1_cond $X=3.18 $Y=0.717
+ $X2=3.015 $Y2=0.717
r40 19 20 7.37564 $w=2.48e-07 $l=1.6e-07 $layer=LI1_cond $X=2.2 $Y=0.595 $X2=2.2
+ $Y2=0.755
r41 16 19 4.84026 $w=2.48e-07 $l=1.05e-07 $layer=LI1_cond $X=2.2 $Y=0.49 $X2=2.2
+ $Y2=0.595
r42 15 20 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.325 $Y=0.755
+ $X2=2.2 $Y2=0.755
r43 15 24 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=2.325 $Y=0.755
+ $X2=3.015 $Y2=0.755
r44 10 16 0.0129374 $w=2.8e-07 $l=1.25e-07 $layer=LI1_cond $X=2.075 $Y=0.49
+ $X2=2.2 $Y2=0.49
r45 10 12 33.1327 $w=2.78e-07 $l=8.05e-07 $layer=LI1_cond $X=2.075 $Y=0.49
+ $X2=1.27 $Y2=0.49
r46 3 23 182 $w=1.7e-07 $l=4.09054e-07 $layer=licon1_NDIFF $count=1 $X=3.04
+ $Y=0.37 $X2=3.18 $Y2=0.715
r47 2 19 182 $w=1.7e-07 $l=2.86575e-07 $layer=licon1_NDIFF $count=1 $X=2.02
+ $Y=0.37 $X2=2.16 $Y2=0.595
r48 1 12 182 $w=1.7e-07 $l=2.20907e-07 $layer=licon1_NDIFF $count=1 $X=1.125
+ $Y=0.37 $X2=1.27 $Y2=0.53
.ends

.subckt PM_SKY130_FD_SC_HS__NAND4B_2%A_490_74# 1 2 7 11 16
r27 14 16 8.85254 $w=2.43e-07 $l=1.65e-07 $layer=LI1_cond $X=2.67 $Y=0.377
+ $X2=2.835 $Y2=0.377
r28 9 11 5.41299 $w=3.28e-07 $l=1.55e-07 $layer=LI1_cond $X=4.17 $Y=0.425
+ $X2=4.17 $Y2=0.58
r29 7 9 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.005 $Y=0.34
+ $X2=4.17 $Y2=0.425
r30 7 16 76.3316 $w=1.68e-07 $l=1.17e-06 $layer=LI1_cond $X=4.005 $Y=0.34
+ $X2=2.835 $Y2=0.34
r31 2 11 182 $w=1.7e-07 $l=2.19089e-07 $layer=licon1_NDIFF $count=1 $X=4.03
+ $Y=0.42 $X2=4.17 $Y2=0.58
r32 1 14 182 $w=1.7e-07 $l=2.41454e-07 $layer=licon1_NDIFF $count=1 $X=2.45
+ $Y=0.37 $X2=2.67 $Y2=0.415
.ends

.subckt PM_SKY130_FD_SC_HS__NAND4B_2%A_719_123# 1 2 3 10 13 14 17 19 21 23 26
r42 21 28 3.40825 $w=2.5e-07 $l=1.25e-07 $layer=LI1_cond $X=5.52 $Y=0.93
+ $X2=5.52 $Y2=1.055
r43 21 23 16.8257 $w=2.48e-07 $l=3.65e-07 $layer=LI1_cond $X=5.52 $Y=0.93
+ $X2=5.52 $Y2=0.565
r44 20 26 4.08801 $w=2.5e-07 $l=9.5e-08 $layer=LI1_cond $X=4.695 $Y=1.055
+ $X2=4.6 $Y2=1.055
r45 19 28 3.40825 $w=2.5e-07 $l=1.25e-07 $layer=LI1_cond $X=5.395 $Y=1.055
+ $X2=5.52 $Y2=1.055
r46 19 20 32.2684 $w=2.48e-07 $l=7e-07 $layer=LI1_cond $X=5.395 $Y=1.055
+ $X2=4.695 $Y2=1.055
r47 15 26 2.34704 $w=1.9e-07 $l=1.25e-07 $layer=LI1_cond $X=4.6 $Y=0.93 $X2=4.6
+ $Y2=1.055
r48 15 17 21.3062 $w=1.88e-07 $l=3.65e-07 $layer=LI1_cond $X=4.6 $Y=0.93 $X2=4.6
+ $Y2=0.565
r49 13 26 4.08801 $w=2.5e-07 $l=9.5e-08 $layer=LI1_cond $X=4.505 $Y=1.055
+ $X2=4.6 $Y2=1.055
r50 13 14 31.3464 $w=2.48e-07 $l=6.8e-07 $layer=LI1_cond $X=4.505 $Y=1.055
+ $X2=3.825 $Y2=1.055
r51 10 14 6.81649 $w=2.5e-07 $l=1.76777e-07 $layer=LI1_cond $X=3.7 $Y=0.93
+ $X2=3.825 $Y2=1.055
r52 10 12 2.196 $w=2.5e-07 $l=4.5e-08 $layer=LI1_cond $X=3.7 $Y=0.93 $X2=3.7
+ $Y2=0.885
r53 3 28 182 $w=1.7e-07 $l=6.61306e-07 $layer=licon1_NDIFF $count=1 $X=5.34
+ $Y=0.42 $X2=5.48 $Y2=1.015
r54 3 23 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=5.34
+ $Y=0.42 $X2=5.48 $Y2=0.565
r55 2 26 182 $w=1.7e-07 $l=6.61306e-07 $layer=licon1_NDIFF $count=1 $X=4.46
+ $Y=0.42 $X2=4.6 $Y2=1.015
r56 2 17 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=4.46
+ $Y=0.42 $X2=4.6 $Y2=0.565
r57 1 12 182 $w=1.7e-07 $l=3.34739e-07 $layer=licon1_NDIFF $count=1 $X=3.595
+ $Y=0.615 $X2=3.74 $Y2=0.885
.ends

