* NGSPICE file created from sky130_fd_sc_hs__dlrbn_1.ext - technology: sky130A

.subckt sky130_fd_sc_hs__dlrbn_1 D GATE_N RESET_B VGND VNB VPB VPWR Q Q_N
M1000 VPWR a_889_92# a_1437_112# VPB pshort w=840000u l=150000u
+  ad=2.32665e+12p pd=1.625e+07u as=2.31e+11p ps=2.23e+06u
M1001 a_608_74# a_27_424# VGND VNB nlowvt w=640000u l=150000u
+  ad=1.536e+11p pd=1.76e+06u as=1.4043e+12p ps=1.104e+07u
M1002 a_686_74# a_231_74# a_608_74# VNB nlowvt w=640000u l=150000u
+  ad=3.835e+11p pd=2.53e+06u as=0p ps=0u
M1003 a_231_74# GATE_N VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1004 Q a_889_92# VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=3.248e+11p pd=2.82e+06u as=0p ps=0u
M1005 VPWR a_231_74# a_373_74# VPB pshort w=840000u l=150000u
+  ad=0p pd=0u as=3.83e+11p ps=2.88e+06u
M1006 VGND RESET_B a_1133_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=1.776e+11p ps=1.96e+06u
M1007 VPWR RESET_B a_889_92# VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=3.472e+11p ps=2.86e+06u
M1008 a_611_392# a_27_424# VPWR VPB pshort w=1e+06u l=150000u
+  ad=2.7e+11p pd=2.54e+06u as=0p ps=0u
M1009 VGND D a_27_424# VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=1.5675e+11p ps=1.67e+06u
M1010 VGND a_889_92# a_1437_112# VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=1.925e+11p ps=1.8e+06u
M1011 a_841_118# a_373_74# a_686_74# VNB nlowvt w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=0p ps=0u
M1012 a_686_74# a_373_74# a_611_392# VPB pshort w=1e+06u l=150000u
+  ad=3.328e+11p pd=2.77e+06u as=0p ps=0u
M1013 VGND a_231_74# a_373_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1014 a_1133_74# a_686_74# a_889_92# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1015 a_231_74# GATE_N VPWR VPB pshort w=840000u l=150000u
+  ad=2.478e+11p pd=2.27e+06u as=0p ps=0u
M1016 VPWR a_889_92# a_802_508# VPB pshort w=420000u l=150000u
+  ad=0p pd=0u as=2.247e+11p ps=1.91e+06u
M1017 a_889_92# a_686_74# VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 Q a_889_92# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1019 VPWR D a_27_424# VPB pshort w=840000u l=150000u
+  ad=0p pd=0u as=2.478e+11p ps=2.27e+06u
M1020 Q_N a_1437_112# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1021 a_802_508# a_231_74# a_686_74# VPB pshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 VGND a_889_92# a_841_118# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 Q_N a_1437_112# VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=3.304e+11p pd=2.83e+06u as=0p ps=0u
.ends

