* File: sky130_fd_sc_hs__mux4_1.pex.spice
* Created: Thu Aug 27 20:49:32 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HS__MUX4_1%A0 1 3 6 8 12
c29 12 0 4.25082e-20 $X=1.155 $Y=1.38
r30 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.155
+ $Y=1.38 $X2=1.155 $Y2=1.38
r31 8 12 9.95292 $w=3.28e-07 $l=2.85e-07 $layer=LI1_cond $X=1.155 $Y=1.665
+ $X2=1.155 $Y2=1.38
r32 4 11 38.5562 $w=2.99e-07 $l=2.05122e-07 $layer=POLY_cond $X=1.245 $Y=1.215
+ $X2=1.155 $Y2=1.38
r33 4 6 269.202 $w=1.5e-07 $l=5.25e-07 $layer=POLY_cond $X=1.245 $Y=1.215
+ $X2=1.245 $Y2=0.69
r34 1 11 52.2586 $w=2.99e-07 $l=2.7157e-07 $layer=POLY_cond $X=1.2 $Y=1.63
+ $X2=1.155 $Y2=1.38
r35 1 3 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=1.2 $Y=1.63 $X2=1.2
+ $Y2=2.205
.ends

.subckt PM_SKY130_FD_SC_HS__MUX4_1%A_27_74# 1 2 9 11 13 16 17 19 22 28 30 33 36
+ 37 39 42 45 49 50 53 54 56 59 61 62 63 65 66 67 69 71 78
c180 67 0 1.99713e-19 $X=1.695 $Y=1.2
c181 63 0 6.3344e-20 $X=1.615 $Y=0.945
c182 53 0 1.11609e-19 $X=4.665 $Y=1.445
c183 50 0 1.18946e-20 $X=4.245 $Y=1.285
c184 49 0 1.11257e-19 $X=4.245 $Y=1.285
c185 17 0 1.88063e-19 $X=5.25 $Y=1.86
r186 66 74 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.695 $Y=1.365
+ $X2=1.695 $Y2=1.2
r187 65 67 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=1.695 $Y=1.365
+ $X2=1.695 $Y2=1.2
r188 65 66 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.695
+ $Y=1.365 $X2=1.695 $Y2=1.365
r189 61 62 6.78944 $w=4.43e-07 $l=8.5e-08 $layer=LI1_cond $X=0.332 $Y=2.035
+ $X2=0.332 $Y2=1.95
r190 56 57 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.175
+ $Y=1.61 $X2=5.175 $Y2=1.61
r191 54 56 14.8421 $w=3.28e-07 $l=4.25e-07 $layer=LI1_cond $X=4.75 $Y=1.61
+ $X2=5.175 $Y2=1.61
r192 53 54 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.665 $Y=1.445
+ $X2=4.75 $Y2=1.61
r193 52 71 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.665 $Y=1.045
+ $X2=4.665 $Y2=0.96
r194 52 53 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=4.665 $Y=1.045
+ $X2=4.665 $Y2=1.445
r195 50 78 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.245 $Y=1.285
+ $X2=4.245 $Y2=1.12
r196 49 50 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.245
+ $Y=1.285 $X2=4.245 $Y2=1.285
r197 47 71 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=4.245 $Y=0.96
+ $X2=4.665 $Y2=0.96
r198 47 49 8.3814 $w=3.28e-07 $l=2.4e-07 $layer=LI1_cond $X=4.245 $Y=1.045
+ $X2=4.245 $Y2=1.285
r199 46 69 2.76166 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.79 $Y=0.96
+ $X2=2.625 $Y2=0.96
r200 45 47 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=4.08 $Y=0.96
+ $X2=4.245 $Y2=0.96
r201 45 46 84.1604 $w=1.68e-07 $l=1.29e-06 $layer=LI1_cond $X=4.08 $Y=0.96
+ $X2=2.79 $Y2=0.96
r202 42 43 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.625
+ $Y=1.285 $X2=2.625 $Y2=1.285
r203 40 69 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.625 $Y=1.045
+ $X2=2.625 $Y2=0.96
r204 40 42 8.3814 $w=3.28e-07 $l=2.4e-07 $layer=LI1_cond $X=2.625 $Y=1.045
+ $X2=2.625 $Y2=1.285
r205 39 69 3.70735 $w=2.5e-07 $l=1.18427e-07 $layer=LI1_cond $X=2.545 $Y=0.875
+ $X2=2.625 $Y2=0.96
r206 38 39 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=2.545 $Y=0.425
+ $X2=2.545 $Y2=0.875
r207 36 38 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.46 $Y=0.34
+ $X2=2.545 $Y2=0.425
r208 36 37 49.5829 $w=1.68e-07 $l=7.6e-07 $layer=LI1_cond $X=2.46 $Y=0.34
+ $X2=1.7 $Y2=0.34
r209 34 63 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.615 $Y=1.03
+ $X2=1.615 $Y2=0.945
r210 34 67 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=1.615 $Y=1.03
+ $X2=1.615 $Y2=1.2
r211 33 63 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.615 $Y=0.86
+ $X2=1.615 $Y2=0.945
r212 32 37 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.615 $Y=0.425
+ $X2=1.7 $Y2=0.34
r213 32 33 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=1.615 $Y=0.425
+ $X2=1.615 $Y2=0.86
r214 31 59 2.79892 $w=1.7e-07 $l=1.68e-07 $layer=LI1_cond $X=0.445 $Y=0.945
+ $X2=0.277 $Y2=0.945
r215 30 63 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.53 $Y=0.945
+ $X2=1.615 $Y2=0.945
r216 30 31 70.7861 $w=1.68e-07 $l=1.085e-06 $layer=LI1_cond $X=1.53 $Y=0.945
+ $X2=0.445 $Y2=0.945
r217 26 61 3.54797 $w=4.43e-07 $l=1.37e-07 $layer=LI1_cond $X=0.332 $Y=2.172
+ $X2=0.332 $Y2=2.035
r218 26 28 14.0624 $w=4.43e-07 $l=5.43e-07 $layer=LI1_cond $X=0.332 $Y=2.172
+ $X2=0.332 $Y2=2.715
r219 24 59 3.67481 $w=2.52e-07 $l=1.19143e-07 $layer=LI1_cond $X=0.195 $Y=1.03
+ $X2=0.277 $Y2=0.945
r220 24 62 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=0.195 $Y=1.03
+ $X2=0.195 $Y2=1.95
r221 20 59 3.67481 $w=2.52e-07 $l=8.5e-08 $layer=LI1_cond $X=0.277 $Y=0.86
+ $X2=0.277 $Y2=0.945
r222 20 22 11.8684 $w=3.33e-07 $l=3.45e-07 $layer=LI1_cond $X=0.277 $Y=0.86
+ $X2=0.277 $Y2=0.515
r223 17 57 52.2586 $w=2.99e-07 $l=2.85044e-07 $layer=POLY_cond $X=5.25 $Y=1.86
+ $X2=5.175 $Y2=1.61
r224 17 19 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=5.25 $Y=1.86
+ $X2=5.25 $Y2=2.435
r225 16 78 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=4.155 $Y=0.69
+ $X2=4.155 $Y2=1.12
r226 11 43 70.0964 $w=2.77e-07 $l=3.5242e-07 $layer=POLY_cond $X=2.61 $Y=1.63
+ $X2=2.625 $Y2=1.285
r227 11 13 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=2.61 $Y=1.63
+ $X2=2.61 $Y2=2.205
r228 9 74 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=1.635 $Y=0.69
+ $X2=1.635 $Y2=1.2
r229 2 61 400 $w=1.7e-07 $l=2.57488e-07 $layer=licon1_PDIFF $count=1 $X=0.245
+ $Y=1.84 $X2=0.39 $Y2=2.035
r230 2 28 400 $w=1.7e-07 $l=9.44722e-07 $layer=licon1_PDIFF $count=1 $X=0.245
+ $Y=1.84 $X2=0.39 $Y2=2.715
r231 1 22 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__MUX4_1%A1 3 5 7 8 9 14
r34 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.165
+ $Y=1.38 $X2=3.165 $Y2=1.38
r35 8 9 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=3.165 $Y=1.665
+ $X2=3.165 $Y2=2.035
r36 8 14 9.95292 $w=3.28e-07 $l=2.85e-07 $layer=LI1_cond $X=3.165 $Y=1.665
+ $X2=3.165 $Y2=1.38
r37 5 13 52.2586 $w=2.99e-07 $l=2.7157e-07 $layer=POLY_cond $X=3.12 $Y=1.63
+ $X2=3.165 $Y2=1.38
r38 5 7 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=3.12 $Y=1.63 $X2=3.12
+ $Y2=2.205
r39 1 13 38.5562 $w=2.99e-07 $l=2.05122e-07 $layer=POLY_cond $X=3.075 $Y=1.215
+ $X2=3.165 $Y2=1.38
r40 1 3 269.202 $w=1.5e-07 $l=5.25e-07 $layer=POLY_cond $X=3.075 $Y=1.215
+ $X2=3.075 $Y2=0.69
.ends

.subckt PM_SKY130_FD_SC_HS__MUX4_1%A2 1 3 6 8 9 14
r34 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.705
+ $Y=1.38 $X2=3.705 $Y2=1.38
r35 8 9 11.5244 $w=3.68e-07 $l=3.7e-07 $layer=LI1_cond $X=3.685 $Y=1.665
+ $X2=3.685 $Y2=2.035
r36 8 14 8.87693 $w=3.68e-07 $l=2.85e-07 $layer=LI1_cond $X=3.685 $Y=1.665
+ $X2=3.685 $Y2=1.38
r37 4 13 38.5562 $w=2.99e-07 $l=1.92678e-07 $layer=POLY_cond $X=3.765 $Y=1.215
+ $X2=3.705 $Y2=1.38
r38 4 6 269.202 $w=1.5e-07 $l=5.25e-07 $layer=POLY_cond $X=3.765 $Y=1.215
+ $X2=3.765 $Y2=0.69
r39 1 13 52.2586 $w=2.99e-07 $l=2.66927e-07 $layer=POLY_cond $X=3.74 $Y=1.63
+ $X2=3.705 $Y2=1.38
r40 1 3 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=3.74 $Y=1.63 $X2=3.74
+ $Y2=2.205
.ends

.subckt PM_SKY130_FD_SC_HS__MUX4_1%S0 3 5 8 9 11 12 13 14 15 18 21 22 27 28 29
+ 31 32 34 35 37 38 41 43 47
c135 37 0 1.25715e-19 $X=2.16 $Y=1.085
c136 32 0 1.11257e-19 $X=4.82 $Y=1.085
c137 11 0 1.37343e-19 $X=2.16 $Y=1.175
c138 8 0 4.25082e-20 $X=0.615 $Y=2.34
r139 46 47 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.615
+ $Y=1.38 $X2=0.615 $Y2=1.38
r140 43 47 8.87693 $w=3.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.635 $Y=1.665
+ $X2=0.635 $Y2=1.38
r141 39 41 48.7128 $w=1.5e-07 $l=9.5e-08 $layer=POLY_cond $X=4.725 $Y=1.16
+ $X2=4.82 $Y2=1.16
r142 32 41 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.82 $Y=1.085
+ $X2=4.82 $Y2=1.16
r143 32 34 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=4.82 $Y=1.085
+ $X2=4.82 $Y2=0.69
r144 30 39 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.725 $Y=1.235
+ $X2=4.725 $Y2=1.16
r145 30 31 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=4.725 $Y=1.235
+ $X2=4.725 $Y2=1.69
r146 28 31 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.65 $Y=1.765
+ $X2=4.725 $Y2=1.69
r147 28 29 161.521 $w=1.5e-07 $l=3.15e-07 $layer=POLY_cond $X=4.65 $Y=1.765
+ $X2=4.335 $Y2=1.765
r148 25 27 294.84 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=4.245 $Y=3.01
+ $X2=4.245 $Y2=2.435
r149 24 29 26.9307 $w=1.5e-07 $l=1.32571e-07 $layer=POLY_cond $X=4.245 $Y=1.86
+ $X2=4.335 $Y2=1.765
r150 24 27 294.84 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=4.245 $Y=1.86
+ $X2=4.245 $Y2=2.435
r151 23 38 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=2.25 $Y=3.15 $X2=2.16
+ $Y2=3.15
r152 22 25 26.9307 $w=1.5e-07 $l=1.79444e-07 $layer=POLY_cond $X=4.155 $Y=3.15
+ $X2=4.245 $Y2=3.01
r153 22 23 976.819 $w=1.5e-07 $l=1.905e-06 $layer=POLY_cond $X=4.155 $Y=3.15
+ $X2=2.25 $Y2=3.15
r154 21 37 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=2.175 $Y=0.69
+ $X2=2.175 $Y2=1.085
r155 16 18 294.84 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=2.16 $Y=2.78
+ $X2=2.16 $Y2=2.205
r156 15 18 294.84 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=2.16 $Y=1.63
+ $X2=2.16 $Y2=2.205
r157 14 38 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=2.16 $Y=3.075
+ $X2=2.16 $Y2=3.15
r158 13 16 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=2.16 $Y=2.87 $X2=2.16
+ $Y2=2.78
r159 13 14 79.6855 $w=1.8e-07 $l=2.05e-07 $layer=POLY_cond $X=2.16 $Y=2.87
+ $X2=2.16 $Y2=3.075
r160 12 15 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=2.16 $Y=1.54 $X2=2.16
+ $Y2=1.63
r161 11 37 37.1337 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=2.16 $Y=1.175
+ $X2=2.16 $Y2=1.085
r162 11 12 141.879 $w=1.8e-07 $l=3.65e-07 $layer=POLY_cond $X=2.16 $Y=1.175
+ $X2=2.16 $Y2=1.54
r163 10 35 7.1379 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=0.705 $Y=3.15
+ $X2=0.615 $Y2=3.15
r164 9 38 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=2.07 $Y=3.15 $X2=2.16
+ $Y2=3.15
r165 9 10 699.926 $w=1.5e-07 $l=1.365e-06 $layer=POLY_cond $X=2.07 $Y=3.15
+ $X2=0.705 $Y2=3.15
r166 6 35 93.4966 $w=1.8e-07 $l=2.35e-07 $layer=POLY_cond $X=0.615 $Y=2.915
+ $X2=0.615 $Y2=3.15
r167 6 8 294.84 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=0.615 $Y=2.915
+ $X2=0.615 $Y2=2.34
r168 5 46 75.4537 $w=2.88e-07 $l=3.92428e-07 $layer=POLY_cond $X=0.615 $Y=1.765
+ $X2=0.6 $Y2=1.38
r169 5 8 294.84 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=0.615 $Y=1.765
+ $X2=0.615 $Y2=2.34
r170 1 46 38.6342 $w=2.88e-07 $l=2.11069e-07 $layer=POLY_cond $X=0.495 $Y=1.215
+ $X2=0.6 $Y2=1.38
r171 1 3 269.202 $w=1.5e-07 $l=5.25e-07 $layer=POLY_cond $X=0.495 $Y=1.215
+ $X2=0.495 $Y2=0.69
.ends

.subckt PM_SKY130_FD_SC_HS__MUX4_1%A3 1 3 4 5 6 8 9
c40 9 0 4.73862e-20 $X=6 $Y=1.665
c41 5 0 1.11609e-19 $X=5.285 $Y=1.16
r42 11 13 41.3143 $w=5.25e-07 $l=4.5e-07 $layer=POLY_cond $X=5.887 $Y=1.16
+ $X2=5.887 $Y2=1.61
r43 9 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.015
+ $Y=1.61 $X2=6.015 $Y2=1.61
r44 6 13 50.382 $w=5.25e-07 $l=3.41687e-07 $layer=POLY_cond $X=5.67 $Y=1.86
+ $X2=5.887 $Y2=1.61
r45 6 8 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=5.67 $Y=1.86 $X2=5.67
+ $Y2=2.435
r46 4 11 32.6451 $w=1.5e-07 $l=2.77e-07 $layer=POLY_cond $X=5.61 $Y=1.16
+ $X2=5.887 $Y2=1.16
r47 4 5 166.649 $w=1.5e-07 $l=3.25e-07 $layer=POLY_cond $X=5.61 $Y=1.16
+ $X2=5.285 $Y2=1.16
r48 1 5 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.21 $Y=1.085
+ $X2=5.285 $Y2=1.16
r49 1 3 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=5.21 $Y=1.085
+ $X2=5.21 $Y2=0.69
.ends

.subckt PM_SKY130_FD_SC_HS__MUX4_1%A_1396_99# 1 2 9 12 13 15 16 18 23 28 30 32
+ 34 37
c67 13 0 2.10579e-19 $X=7.18 $Y=1.885
r68 34 36 17.4812 $w=5.43e-07 $l=5.15e-07 $layer=LI1_cond $X=8.137 $Y=0.665
+ $X2=8.137 $Y2=1.18
r69 31 32 10.4914 $w=1.83e-07 $l=1.75e-07 $layer=LI1_cond $X=7.942 $Y=1.775
+ $X2=7.942 $Y2=1.95
r70 30 36 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=7.95 $Y=1.445
+ $X2=7.95 $Y2=1.18
r71 29 37 16.6118 $w=3.3e-07 $l=9.5e-08 $layer=POLY_cond $X=7.795 $Y=1.61
+ $X2=7.795 $Y2=1.515
r72 28 31 8.13117 $w=4.03e-07 $l=1.65e-07 $layer=LI1_cond $X=7.832 $Y=1.61
+ $X2=7.832 $Y2=1.775
r73 28 30 8.6688 $w=4.03e-07 $l=1.65e-07 $layer=LI1_cond $X=7.832 $Y=1.61
+ $X2=7.832 $Y2=1.445
r74 28 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.795
+ $Y=1.61 $X2=7.795 $Y2=1.61
r75 23 32 7.96936 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=8.015 $Y=2.115
+ $X2=8.015 $Y2=1.95
r76 17 18 6.66866 $w=1.5e-07 $l=1.45e-07 $layer=POLY_cond $X=7.27 $Y=1.515
+ $X2=7.125 $Y2=1.515
r77 16 37 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.63 $Y=1.515
+ $X2=7.795 $Y2=1.515
r78 16 17 184.596 $w=1.5e-07 $l=3.6e-07 $layer=POLY_cond $X=7.63 $Y=1.515
+ $X2=7.27 $Y2=1.515
r79 13 15 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=7.18 $Y=1.885
+ $X2=7.18 $Y2=2.46
r80 12 13 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=7.18 $Y=1.795 $X2=7.18
+ $Y2=1.885
r81 11 18 18.8402 $w=1.65e-07 $l=9.87421e-08 $layer=POLY_cond $X=7.18 $Y=1.59
+ $X2=7.125 $Y2=1.515
r82 11 12 79.6855 $w=1.8e-07 $l=2.05e-07 $layer=POLY_cond $X=7.18 $Y=1.59
+ $X2=7.18 $Y2=1.795
r83 7 18 18.8402 $w=1.65e-07 $l=1.04283e-07 $layer=POLY_cond $X=7.055 $Y=1.44
+ $X2=7.125 $Y2=1.515
r84 7 9 253.819 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=7.055 $Y=1.44
+ $X2=7.055 $Y2=0.945
r85 2 23 300 $w=1.7e-07 $l=2.41868e-07 $layer=licon1_PDIFF $count=2 $X=7.87
+ $Y=1.935 $X2=8.015 $Y2=2.115
r86 1 34 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=8.1
+ $Y=0.52 $X2=8.245 $Y2=0.665
.ends

.subckt PM_SKY130_FD_SC_HS__MUX4_1%S1 4 6 7 9 10 11 12 14 18 20 21 25
c78 20 0 4.73862e-20 $X=6.655 $Y=1.49
c79 12 0 7.34196e-20 $X=8.29 $Y=1.86
c80 4 0 1.50188e-19 $X=6.615 $Y=0.945
r81 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.37
+ $Y=1.515 $X2=8.37 $Y2=1.515
r82 21 25 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=8.37 $Y=1.665
+ $X2=8.37 $Y2=1.515
r83 19 20 60.4563 $w=1.8e-07 $l=1.5e-07 $layer=POLY_cond $X=6.655 $Y=1.34
+ $X2=6.655 $Y2=1.49
r84 16 24 38.7751 $w=2.77e-07 $l=2.06325e-07 $layer=POLY_cond $X=8.46 $Y=1.35
+ $X2=8.367 $Y2=1.515
r85 16 18 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=8.46 $Y=1.35
+ $X2=8.46 $Y2=0.84
r86 15 18 299.968 $w=1.5e-07 $l=5.85e-07 $layer=POLY_cond $X=8.46 $Y=0.255
+ $X2=8.46 $Y2=0.84
r87 12 24 70.0964 $w=2.77e-07 $l=3.81563e-07 $layer=POLY_cond $X=8.29 $Y=1.86
+ $X2=8.367 $Y2=1.515
r88 12 14 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=8.29 $Y=1.86
+ $X2=8.29 $Y2=2.435
r89 10 15 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=8.385 $Y=0.18
+ $X2=8.46 $Y2=0.255
r90 10 11 869.138 $w=1.5e-07 $l=1.695e-06 $layer=POLY_cond $X=8.385 $Y=0.18
+ $X2=6.69 $Y2=0.18
r91 7 9 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=6.68 $Y=1.885
+ $X2=6.68 $Y2=2.46
r92 6 7 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=6.68 $Y=1.795 $X2=6.68
+ $Y2=1.885
r93 6 20 118.556 $w=1.8e-07 $l=3.05e-07 $layer=POLY_cond $X=6.68 $Y=1.795
+ $X2=6.68 $Y2=1.49
r94 4 19 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=6.615 $Y=0.945
+ $X2=6.615 $Y2=1.34
r95 1 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=6.615 $Y=0.255
+ $X2=6.69 $Y2=0.18
r96 1 4 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=6.615 $Y=0.255
+ $X2=6.615 $Y2=0.945
.ends

.subckt PM_SKY130_FD_SC_HS__MUX4_1%A_1338_125# 1 2 9 11 13 14 17 20 21 23 24 25
+ 27 31
c77 24 0 7.34196e-20 $X=8.745 $Y=2.035
c78 14 0 1.50188e-19 $X=6.955 $Y=1.285
r79 31 34 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=8.91 $Y=1.515
+ $X2=8.91 $Y2=1.68
r80 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.91
+ $Y=1.515 $X2=8.91 $Y2=1.515
r81 27 34 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=8.83 $Y=1.95 $X2=8.83
+ $Y2=1.68
r82 24 27 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.745 $Y=2.035
+ $X2=8.83 $Y2=1.95
r83 24 25 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=8.745 $Y=2.035
+ $X2=8.52 $Y2=2.035
r84 22 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.435 $Y=2.12
+ $X2=8.52 $Y2=2.035
r85 22 23 51.2139 $w=1.68e-07 $l=7.85e-07 $layer=LI1_cond $X=8.435 $Y=2.12
+ $X2=8.435 $Y2=2.905
r86 20 23 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.35 $Y=2.99
+ $X2=8.435 $Y2=2.905
r87 20 21 80.246 $w=1.68e-07 $l=1.23e-06 $layer=LI1_cond $X=8.35 $Y=2.99
+ $X2=7.12 $Y2=2.99
r88 17 19 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=6.955 $Y=2.105
+ $X2=6.955 $Y2=2.815
r89 15 21 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=6.955 $Y=2.905
+ $X2=7.12 $Y2=2.99
r90 15 19 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=6.955 $Y=2.905
+ $X2=6.955 $Y2=2.815
r91 14 29 6.41518 $w=3.3e-07 $l=1.76125e-07 $layer=LI1_cond $X=6.955 $Y=1.285
+ $X2=6.932 $Y2=1.12
r92 14 17 28.6365 $w=3.28e-07 $l=8.2e-07 $layer=LI1_cond $X=6.955 $Y=1.285
+ $X2=6.955 $Y2=2.105
r93 11 32 50.0734 $w=3.74e-07 $l=3.05369e-07 $layer=POLY_cond $X=9.08 $Y=1.765
+ $X2=8.957 $Y2=1.515
r94 11 13 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=9.08 $Y=1.765
+ $X2=9.08 $Y2=2.4
r95 7 32 39.1188 $w=3.74e-07 $l=1.98167e-07 $layer=POLY_cond $X=9.03 $Y=1.35
+ $X2=8.957 $Y2=1.515
r96 7 9 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=9.03 $Y=1.35 $X2=9.03
+ $Y2=0.79
r97 2 19 400 $w=1.7e-07 $l=9.4975e-07 $layer=licon1_PDIFF $count=1 $X=6.755
+ $Y=1.96 $X2=6.955 $Y2=2.815
r98 2 17 400 $w=1.7e-07 $l=2.62678e-07 $layer=licon1_PDIFF $count=1 $X=6.755
+ $Y=1.96 $X2=6.955 $Y2=2.105
r99 1 29 182 $w=1.7e-07 $l=5.6285e-07 $layer=licon1_NDIFF $count=1 $X=6.69
+ $Y=0.625 $X2=6.835 $Y2=1.12
.ends

.subckt PM_SKY130_FD_SC_HS__MUX4_1%VPWR 1 2 3 4 15 21 25 29 32 33 35 36 37 49 56
+ 63 64 67 70
c92 25 0 1.88063e-19 $X=5.895 $Y=2.775
r93 70 71 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r94 67 68 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r95 64 71 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.36 $Y=3.33
+ $X2=8.88 $Y2=3.33
r96 63 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.36 $Y=3.33
+ $X2=9.36 $Y2=3.33
r97 61 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.02 $Y=3.33
+ $X2=8.855 $Y2=3.33
r98 61 63 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=9.02 $Y=3.33
+ $X2=9.36 $Y2=3.33
r99 60 71 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=3.33
+ $X2=8.88 $Y2=3.33
r100 60 68 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=8.4 $Y=3.33 $X2=6
+ $Y2=3.33
r101 59 60 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=8.4 $Y=3.33 $X2=8.4
+ $Y2=3.33
r102 57 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.06 $Y=3.33
+ $X2=5.895 $Y2=3.33
r103 57 59 152.663 $w=1.68e-07 $l=2.34e-06 $layer=LI1_cond $X=6.06 $Y=3.33
+ $X2=8.4 $Y2=3.33
r104 56 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.69 $Y=3.33
+ $X2=8.855 $Y2=3.33
r105 56 59 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=8.69 $Y=3.33
+ $X2=8.4 $Y2=3.33
r106 55 68 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=3.33 $X2=6
+ $Y2=3.33
r107 54 55 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r108 51 54 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=3.6 $Y=3.33
+ $X2=5.52 $Y2=3.33
r109 51 52 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r110 49 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.73 $Y=3.33
+ $X2=5.895 $Y2=3.33
r111 49 54 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=5.73 $Y=3.33
+ $X2=5.52 $Y2=3.33
r112 48 52 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=3.6 $Y2=3.33
r113 47 48 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r114 45 48 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=3.12 $Y2=3.33
r115 44 47 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=1.2 $Y=3.33
+ $X2=3.12 $Y2=3.33
r116 44 45 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r117 41 45 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r118 40 41 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r119 37 55 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=4.8 $Y=3.33
+ $X2=5.52 $Y2=3.33
r120 37 52 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=4.8 $Y=3.33
+ $X2=3.6 $Y2=3.33
r121 35 47 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=3.265 $Y=3.33
+ $X2=3.12 $Y2=3.33
r122 35 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.265 $Y=3.33
+ $X2=3.43 $Y2=3.33
r123 34 51 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=3.595 $Y=3.33
+ $X2=3.6 $Y2=3.33
r124 34 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.595 $Y=3.33
+ $X2=3.43 $Y2=3.33
r125 32 40 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=0.725 $Y=3.33
+ $X2=0.72 $Y2=3.33
r126 32 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.725 $Y=3.33
+ $X2=0.89 $Y2=3.33
r127 31 44 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=1.055 $Y=3.33
+ $X2=1.2 $Y2=3.33
r128 31 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.055 $Y=3.33
+ $X2=0.89 $Y2=3.33
r129 27 70 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.855 $Y=3.245
+ $X2=8.855 $Y2=3.33
r130 27 29 27.5888 $w=3.28e-07 $l=7.9e-07 $layer=LI1_cond $X=8.855 $Y=3.245
+ $X2=8.855 $Y2=2.455
r131 23 67 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.895 $Y=3.245
+ $X2=5.895 $Y2=3.33
r132 23 25 16.4136 $w=3.28e-07 $l=4.7e-07 $layer=LI1_cond $X=5.895 $Y=3.245
+ $X2=5.895 $Y2=2.775
r133 19 36 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.43 $Y=3.245
+ $X2=3.43 $Y2=3.33
r134 19 21 14.1436 $w=3.28e-07 $l=4.05e-07 $layer=LI1_cond $X=3.43 $Y=3.245
+ $X2=3.43 $Y2=2.84
r135 15 18 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=0.89 $Y=2.035
+ $X2=0.89 $Y2=2.715
r136 13 33 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.89 $Y=3.245
+ $X2=0.89 $Y2=3.33
r137 13 18 18.5089 $w=3.28e-07 $l=5.3e-07 $layer=LI1_cond $X=0.89 $Y=3.245
+ $X2=0.89 $Y2=2.715
r138 4 29 300 $w=1.7e-07 $l=7.24707e-07 $layer=licon1_PDIFF $count=2 $X=8.365
+ $Y=1.935 $X2=8.855 $Y2=2.455
r139 3 25 600 $w=1.7e-07 $l=9.11921e-07 $layer=licon1_PDIFF $count=1 $X=5.745
+ $Y=1.935 $X2=5.895 $Y2=2.775
r140 2 21 600 $w=1.7e-07 $l=1.24698e-06 $layer=licon1_PDIFF $count=1 $X=3.195
+ $Y=1.705 $X2=3.43 $Y2=2.84
r141 1 18 600 $w=1.7e-07 $l=9.69858e-07 $layer=licon1_PDIFF $count=1 $X=0.69
+ $Y=1.84 $X2=0.89 $Y2=2.715
r142 1 15 300 $w=1.7e-07 $l=2.81069e-07 $layer=licon1_PDIFF $count=2 $X=0.69
+ $Y=1.84 $X2=0.89 $Y2=2.035
.ends

.subckt PM_SKY130_FD_SC_HS__MUX4_1%A_342_74# 1 2 3 4 16 17 20 21 22 24 25 26 28
+ 30 33 38 42 45 46 47 51 52 54 55
c142 52 0 1.25754e-19 $X=6.455 $Y=2.42
c143 33 0 1.17971e-19 $X=6.455 $Y=2.815
c144 30 0 9.26086e-20 $X=6.455 $Y=2.115
c145 21 0 5.47968e-20 $X=5.35 $Y=2.99
r146 54 55 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=7.27 $Y=0.77
+ $X2=7.105 $Y2=0.77
r147 47 49 3.22021 $w=5.18e-07 $l=1.4e-07 $layer=LI1_cond $X=2.29 $Y=2.42
+ $X2=2.29 $Y2=2.56
r148 45 46 9.6413 $w=5.18e-07 $l=1.65e-07 $layer=LI1_cond $X=2.29 $Y=1.85
+ $X2=2.29 $Y2=1.685
r149 40 42 4.10641 $w=4.33e-07 $l=1.55e-07 $layer=LI1_cond $X=1.96 $Y=0.812
+ $X2=2.115 $Y2=0.812
r150 38 55 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=6.575 $Y=0.7
+ $X2=7.105 $Y2=0.7
r151 35 38 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.49 $Y=0.785
+ $X2=6.575 $Y2=0.7
r152 35 51 76.0053 $w=1.68e-07 $l=1.165e-06 $layer=LI1_cond $X=6.49 $Y=0.785
+ $X2=6.49 $Y2=1.95
r153 31 52 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.455 $Y=2.505
+ $X2=6.455 $Y2=2.42
r154 31 33 10.826 $w=3.28e-07 $l=3.1e-07 $layer=LI1_cond $X=6.455 $Y=2.505
+ $X2=6.455 $Y2=2.815
r155 30 51 7.49019 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=6.455 $Y=2.115
+ $X2=6.455 $Y2=1.95
r156 28 52 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.455 $Y=2.335
+ $X2=6.455 $Y2=2.42
r157 28 30 7.68295 $w=3.28e-07 $l=2.2e-07 $layer=LI1_cond $X=6.455 $Y=2.335
+ $X2=6.455 $Y2=2.115
r158 25 52 3.80956 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.29 $Y=2.42
+ $X2=6.455 $Y2=2.42
r159 25 26 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=6.29 $Y=2.42
+ $X2=5.55 $Y2=2.42
r160 23 26 6.87494 $w=1.7e-07 $l=1.36015e-07 $layer=LI1_cond $X=5.45 $Y=2.505
+ $X2=5.55 $Y2=2.42
r161 23 24 22.1818 $w=1.98e-07 $l=4e-07 $layer=LI1_cond $X=5.45 $Y=2.505
+ $X2=5.45 $Y2=2.905
r162 21 24 6.87494 $w=1.7e-07 $l=1.36015e-07 $layer=LI1_cond $X=5.35 $Y=2.99
+ $X2=5.45 $Y2=2.905
r163 21 22 86.7701 $w=1.68e-07 $l=1.33e-06 $layer=LI1_cond $X=5.35 $Y=2.99
+ $X2=4.02 $Y2=2.99
r164 20 22 6.9898 $w=1.7e-07 $l=1.49579e-07 $layer=LI1_cond $X=3.907 $Y=2.905
+ $X2=4.02 $Y2=2.99
r165 19 20 20.4879 $w=2.23e-07 $l=4e-07 $layer=LI1_cond $X=3.907 $Y=2.505
+ $X2=3.907 $Y2=2.905
r166 18 47 7.40362 $w=1.7e-07 $l=2.6e-07 $layer=LI1_cond $X=2.55 $Y=2.42
+ $X2=2.29 $Y2=2.42
r167 17 19 6.9898 $w=1.7e-07 $l=1.4854e-07 $layer=LI1_cond $X=3.795 $Y=2.42
+ $X2=3.907 $Y2=2.505
r168 17 18 81.2246 $w=1.68e-07 $l=1.245e-06 $layer=LI1_cond $X=3.795 $Y=2.42
+ $X2=2.55 $Y2=2.42
r169 16 47 1.95513 $w=5.18e-07 $l=8.5e-08 $layer=LI1_cond $X=2.29 $Y=2.335
+ $X2=2.29 $Y2=2.42
r170 15 45 2.18514 $w=5.18e-07 $l=9.5e-08 $layer=LI1_cond $X=2.29 $Y=1.945
+ $X2=2.29 $Y2=1.85
r171 15 16 8.97059 $w=5.18e-07 $l=3.9e-07 $layer=LI1_cond $X=2.29 $Y=1.945
+ $X2=2.29 $Y2=2.335
r172 13 42 6.29128 $w=1.7e-07 $l=2.18e-07 $layer=LI1_cond $X=2.115 $Y=1.03
+ $X2=2.115 $Y2=0.812
r173 13 46 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=2.115 $Y=1.03
+ $X2=2.115 $Y2=1.685
r174 4 33 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=6.31
+ $Y=1.96 $X2=6.455 $Y2=2.815
r175 4 30 400 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_PDIFF $count=1 $X=6.31
+ $Y=1.96 $X2=6.455 $Y2=2.115
r176 3 49 400 $w=1.7e-07 $l=9.26971e-07 $layer=licon1_PDIFF $count=1 $X=2.235
+ $Y=1.705 $X2=2.385 $Y2=2.56
r177 3 45 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=2.235
+ $Y=1.705 $X2=2.385 $Y2=1.85
r178 2 54 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=7.13
+ $Y=0.625 $X2=7.27 $Y2=0.77
r179 1 40 182 $w=1.7e-07 $l=5.50999e-07 $layer=licon1_NDIFF $count=1 $X=1.71
+ $Y=0.37 $X2=1.96 $Y2=0.81
.ends

.subckt PM_SKY130_FD_SC_HS__MUX4_1%A_846_74# 1 2 3 4 13 18 19 20 21 24 25 27 30
+ 31 33 39 42 46 47 50 53 55
c122 46 0 1.18946e-20 $X=5.165 $Y=2.365
r123 51 53 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=7.375 $Y=1.19
+ $X2=7.61 $Y2=1.19
r124 44 46 10.6559 $w=7.38e-07 $l=1.4e-07 $layer=LI1_cond $X=5.025 $Y=2.365
+ $X2=5.165 $Y2=2.365
r125 42 53 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.61 $Y=1.105
+ $X2=7.61 $Y2=1.19
r126 41 42 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=7.61 $Y=0.435
+ $X2=7.61 $Y2=1.105
r127 39 55 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=7.455 $Y=2.11
+ $X2=7.455 $Y2=1.945
r128 35 51 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.375 $Y=1.275
+ $X2=7.375 $Y2=1.19
r129 35 55 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=7.375 $Y=1.275
+ $X2=7.375 $Y2=1.945
r130 33 41 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.525 $Y=0.35
+ $X2=7.61 $Y2=0.435
r131 33 50 67.8503 $w=1.68e-07 $l=1.04e-06 $layer=LI1_cond $X=7.525 $Y=0.35
+ $X2=6.485 $Y2=0.35
r132 32 49 4.10122 $w=1.8e-07 $l=1.25e-07 $layer=LI1_cond $X=6.235 $Y=0.355
+ $X2=6.11 $Y2=0.355
r133 31 50 5.59224 $w=1.78e-07 $l=9e-08 $layer=LI1_cond $X=6.395 $Y=0.355
+ $X2=6.485 $Y2=0.355
r134 31 32 9.85859 $w=1.78e-07 $l=1.6e-07 $layer=LI1_cond $X=6.395 $Y=0.355
+ $X2=6.235 $Y2=0.355
r135 28 30 13.1378 $w=2.48e-07 $l=2.85e-07 $layer=LI1_cond $X=6.11 $Y=1.105
+ $X2=6.11 $Y2=0.82
r136 27 49 2.95288 $w=2.5e-07 $l=9e-08 $layer=LI1_cond $X=6.11 $Y=0.445 $X2=6.11
+ $Y2=0.355
r137 27 30 17.2866 $w=2.48e-07 $l=3.75e-07 $layer=LI1_cond $X=6.11 $Y=0.445
+ $X2=6.11 $Y2=0.82
r138 26 47 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.68 $Y=1.19
+ $X2=5.595 $Y2=1.19
r139 25 28 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=5.985 $Y=1.19
+ $X2=6.11 $Y2=1.105
r140 25 26 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=5.985 $Y=1.19
+ $X2=5.68 $Y2=1.19
r141 23 47 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.595 $Y=1.275
+ $X2=5.595 $Y2=1.19
r142 23 24 46.9733 $w=1.68e-07 $l=7.2e-07 $layer=LI1_cond $X=5.595 $Y=1.275
+ $X2=5.595 $Y2=1.995
r143 21 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.51 $Y=2.08
+ $X2=5.595 $Y2=1.995
r144 21 46 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=5.51 $Y=2.08
+ $X2=5.165 $Y2=2.08
r145 19 47 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.51 $Y=1.19
+ $X2=5.595 $Y2=1.19
r146 19 20 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=5.51 $Y=1.19
+ $X2=5.09 $Y2=1.19
r147 18 20 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.005 $Y=1.105
+ $X2=5.09 $Y2=1.19
r148 17 18 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=5.005 $Y=0.705
+ $X2=5.005 $Y2=1.105
r149 13 17 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.92 $Y=0.54
+ $X2=5.005 $Y2=0.705
r150 13 15 15.1913 $w=3.28e-07 $l=4.35e-07 $layer=LI1_cond $X=4.92 $Y=0.54
+ $X2=4.485 $Y2=0.54
r151 4 39 300 $w=1.7e-07 $l=2.64575e-07 $layer=licon1_PDIFF $count=2 $X=7.255
+ $Y=1.96 $X2=7.455 $Y2=2.11
r152 3 44 150 $w=1.7e-07 $l=7.74112e-07 $layer=licon1_PDIFF $count=4 $X=4.32
+ $Y=1.935 $X2=5.025 $Y2=2.08
r153 2 49 182 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_NDIFF $count=1 $X=5.995
+ $Y=0.215 $X2=6.15 $Y2=0.36
r154 2 30 182 $w=1.7e-07 $l=6.78086e-07 $layer=licon1_NDIFF $count=1 $X=5.995
+ $Y=0.215 $X2=6.15 $Y2=0.82
r155 1 15 182 $w=1.7e-07 $l=3.29204e-07 $layer=licon1_NDIFF $count=1 $X=4.23
+ $Y=0.37 $X2=4.485 $Y2=0.54
.ends

.subckt PM_SKY130_FD_SC_HS__MUX4_1%X 1 2 7 8 9 10 11 12 13 30
r20 22 30 1.50814 $w=4.03e-07 $l=5.3e-08 $layer=LI1_cond $X=9.282 $Y=0.978
+ $X2=9.282 $Y2=0.925
r21 13 45 7.30194 $w=2.63e-07 $l=1.65e-07 $layer=LI1_cond $X=9.352 $Y=2.725
+ $X2=9.352 $Y2=2.56
r22 12 45 7.44286 $w=2.38e-07 $l=1.55e-07 $layer=LI1_cond $X=9.365 $Y=2.405
+ $X2=9.365 $Y2=2.56
r23 11 12 17.7668 $w=2.38e-07 $l=3.7e-07 $layer=LI1_cond $X=9.365 $Y=2.035
+ $X2=9.365 $Y2=2.405
r24 10 11 17.7668 $w=2.38e-07 $l=3.7e-07 $layer=LI1_cond $X=9.365 $Y=1.665
+ $X2=9.365 $Y2=2.035
r25 9 10 17.7668 $w=2.38e-07 $l=3.7e-07 $layer=LI1_cond $X=9.365 $Y=1.295
+ $X2=9.365 $Y2=1.665
r26 9 42 5.52212 $w=2.38e-07 $l=1.15e-07 $layer=LI1_cond $X=9.365 $Y=1.295
+ $X2=9.365 $Y2=1.18
r27 8 42 7.19001 $w=4.03e-07 $l=1.86e-07 $layer=LI1_cond $X=9.282 $Y=0.994
+ $X2=9.282 $Y2=1.18
r28 8 22 0.455286 $w=4.03e-07 $l=1.6e-08 $layer=LI1_cond $X=9.282 $Y=0.994
+ $X2=9.282 $Y2=0.978
r29 8 30 0.455286 $w=4.03e-07 $l=1.6e-08 $layer=LI1_cond $X=9.282 $Y=0.909
+ $X2=9.282 $Y2=0.925
r30 8 27 9.78865 $w=4.03e-07 $l=3.44e-07 $layer=LI1_cond $X=9.282 $Y=0.909
+ $X2=9.282 $Y2=0.565
r31 7 27 0.284554 $w=4.03e-07 $l=1e-08 $layer=LI1_cond $X=9.282 $Y=0.555
+ $X2=9.282 $Y2=0.565
r32 2 13 600 $w=1.7e-07 $l=9.59375e-07 $layer=licon1_PDIFF $count=1 $X=9.155
+ $Y=1.84 $X2=9.31 $Y2=2.725
r33 1 27 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=9.105
+ $Y=0.42 $X2=9.245 $Y2=0.565
.ends

.subckt PM_SKY130_FD_SC_HS__MUX4_1%VGND 1 2 3 4 17 21 25 29 32 33 34 36 44 57 58
+ 61 64 67
r83 67 68 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=5.52 $Y=0
+ $X2=5.52 $Y2=0
r84 64 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r85 61 62 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r86 57 58 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.36 $Y=0 $X2=9.36
+ $Y2=0
r87 55 58 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=8.4 $Y=0 $X2=9.36
+ $Y2=0
r88 55 68 0.802756 $w=4.9e-07 $l=2.88e-06 $layer=MET1_cond $X=8.4 $Y=0 $X2=5.52
+ $Y2=0
r89 54 55 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=8.4 $Y=0
+ $X2=8.4 $Y2=0
r90 52 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.59 $Y=0 $X2=5.425
+ $Y2=0
r91 52 54 183.326 $w=1.68e-07 $l=2.81e-06 $layer=LI1_cond $X=5.59 $Y=0 $X2=8.4
+ $Y2=0
r92 51 68 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=5.52
+ $Y2=0
r93 50 51 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r94 48 65 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=3.6
+ $Y2=0
r95 47 50 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=4.08 $Y=0 $X2=5.04
+ $Y2=0
r96 47 48 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r97 45 64 12.4404 $w=1.7e-07 $l=2.95e-07 $layer=LI1_cond $X=3.715 $Y=0 $X2=3.42
+ $Y2=0
r98 45 47 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=3.715 $Y=0 $X2=4.08
+ $Y2=0
r99 44 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.26 $Y=0 $X2=5.425
+ $Y2=0
r100 44 50 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=5.26 $Y=0 $X2=5.04
+ $Y2=0
r101 43 65 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=3.6
+ $Y2=0
r102 42 43 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.12 $Y=0
+ $X2=3.12 $Y2=0
r103 40 43 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=1.2 $Y=0 $X2=3.12
+ $Y2=0
r104 40 62 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r105 39 42 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=1.2 $Y=0 $X2=3.12
+ $Y2=0
r106 39 40 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r107 37 61 9.6488 $w=1.7e-07 $l=1.95e-07 $layer=LI1_cond $X=1.09 $Y=0 $X2=0.895
+ $Y2=0
r108 37 39 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=1.09 $Y=0 $X2=1.2
+ $Y2=0
r109 36 64 12.4404 $w=1.7e-07 $l=2.95e-07 $layer=LI1_cond $X=3.125 $Y=0 $X2=3.42
+ $Y2=0
r110 36 42 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=3.125 $Y=0 $X2=3.12
+ $Y2=0
r111 34 51 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=4.8 $Y=0 $X2=5.04
+ $Y2=0
r112 34 48 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=4.8 $Y=0 $X2=4.08
+ $Y2=0
r113 32 54 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=8.58 $Y=0 $X2=8.4
+ $Y2=0
r114 32 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.58 $Y=0 $X2=8.745
+ $Y2=0
r115 31 57 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=8.91 $Y=0 $X2=9.36
+ $Y2=0
r116 31 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.91 $Y=0 $X2=8.745
+ $Y2=0
r117 27 33 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.745 $Y=0.085
+ $X2=8.745 $Y2=0
r118 27 29 20.2551 $w=3.28e-07 $l=5.8e-07 $layer=LI1_cond $X=8.745 $Y=0.085
+ $X2=8.745 $Y2=0.665
r119 23 67 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.425 $Y=0.085
+ $X2=5.425 $Y2=0
r120 23 25 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=5.425 $Y=0.085
+ $X2=5.425 $Y2=0.495
r121 19 64 2.48142 $w=5.9e-07 $l=8.5e-08 $layer=LI1_cond $X=3.42 $Y=0.085
+ $X2=3.42 $Y2=0
r122 19 21 8.71718 $w=5.88e-07 $l=4.3e-07 $layer=LI1_cond $X=3.42 $Y=0.085
+ $X2=3.42 $Y2=0.515
r123 15 61 1.39532 $w=3.9e-07 $l=8.5e-08 $layer=LI1_cond $X=0.895 $Y=0.085
+ $X2=0.895 $Y2=0
r124 15 17 13.7407 $w=3.88e-07 $l=4.65e-07 $layer=LI1_cond $X=0.895 $Y=0.085
+ $X2=0.895 $Y2=0.55
r125 4 29 91 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=2 $X=8.535
+ $Y=0.52 $X2=8.745 $Y2=0.665
r126 3 25 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=5.285
+ $Y=0.37 $X2=5.425 $Y2=0.495
r127 2 21 182 $w=1.7e-07 $l=3.34739e-07 $layer=licon1_NDIFF $count=1 $X=3.15
+ $Y=0.37 $X2=3.42 $Y2=0.515
r128 1 17 182 $w=1.7e-07 $l=4.05123e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.37 $X2=0.895 $Y2=0.55
.ends

