* File: sky130_fd_sc_hs__a222oi_2.pex.spice
* Created: Tue Sep  1 19:51:00 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HS__A222OI_2%C2 2 3 5 8 10 12 15 17 18 20 21 22 25 26 28
+ 32
c93 25 0 1.11993e-19 $X=1.96 $Y=1.295
r94 33 40 6.84127 $w=4.08e-07 $l=1.65e-07 $layer=LI1_cond $X=0.63 $Y=1.33
+ $X2=0.63 $Y2=1.495
r95 32 35 40.7132 $w=3.4e-07 $l=1.65e-07 $layer=POLY_cond $X=0.585 $Y=1.33
+ $X2=0.585 $Y2=1.495
r96 32 34 46.3065 $w=3.4e-07 $l=1.65e-07 $layer=POLY_cond $X=0.585 $Y=1.33
+ $X2=0.585 $Y2=1.165
r97 32 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.59
+ $Y=1.33 $X2=0.59 $Y2=1.33
r98 28 33 0.983793 $w=4.08e-07 $l=3.5e-08 $layer=LI1_cond $X=0.63 $Y=1.295
+ $X2=0.63 $Y2=1.33
r99 25 26 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.96
+ $Y=1.295 $X2=1.96 $Y2=1.295
r100 23 25 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.96 $Y=1.665
+ $X2=1.96 $Y2=1.295
r101 21 23 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.795 $Y=1.75
+ $X2=1.96 $Y2=1.665
r102 21 22 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.795 $Y=1.75
+ $X2=0.835 $Y2=1.75
r103 20 22 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=0.72 $Y=1.665
+ $X2=0.835 $Y2=1.75
r104 20 40 8.51806 $w=2.28e-07 $l=1.7e-07 $layer=LI1_cond $X=0.72 $Y=1.665
+ $X2=0.72 $Y2=1.495
r105 18 26 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.96 $Y=1.635
+ $X2=1.96 $Y2=1.295
r106 17 26 41.8716 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.96 $Y=1.13
+ $X2=1.96 $Y2=1.295
r107 15 17 141.387 $w=1.5e-07 $l=4.4e-07 $layer=POLY_cond $X=1.9 $Y=0.69 $X2=1.9
+ $Y2=1.13
r108 10 18 43.19 $w=2.79e-07 $l=2.85044e-07 $layer=POLY_cond $X=1.885 $Y=1.885
+ $X2=1.96 $Y2=1.635
r109 10 12 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=1.885 $Y=1.885
+ $X2=1.885 $Y2=2.46
r110 8 34 243.564 $w=1.5e-07 $l=4.75e-07 $layer=POLY_cond $X=0.61 $Y=0.69
+ $X2=0.61 $Y2=1.165
r111 3 5 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=0.505 $Y=1.885
+ $X2=0.505 $Y2=2.46
r112 2 3 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=0.505 $Y=1.795
+ $X2=0.505 $Y2=1.885
r113 2 35 116.613 $w=1.8e-07 $l=3e-07 $layer=POLY_cond $X=0.505 $Y=1.795
+ $X2=0.505 $Y2=1.495
.ends

.subckt PM_SKY130_FD_SC_HS__A222OI_2%C1 1 3 6 9 11 12 14 17 21 23 31
r62 30 31 6.12014 $w=3.3e-07 $l=3.5e-08 $layer=POLY_cond $X=1.435 $Y=1.33
+ $X2=1.47 $Y2=1.33
r63 28 30 46.3382 $w=3.3e-07 $l=2.65e-07 $layer=POLY_cond $X=1.17 $Y=1.33
+ $X2=1.435 $Y2=1.33
r64 25 28 22.732 $w=3.3e-07 $l=1.3e-07 $layer=POLY_cond $X=1.04 $Y=1.33 $X2=1.17
+ $Y2=1.33
r65 23 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.17
+ $Y=1.33 $X2=1.17 $Y2=1.33
r66 19 21 43.5851 $w=1.5e-07 $l=8.5e-08 $layer=POLY_cond $X=0.955 $Y=1.81
+ $X2=1.04 $Y2=1.81
r67 15 31 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.47 $Y=1.165
+ $X2=1.47 $Y2=1.33
r68 15 17 243.564 $w=1.5e-07 $l=4.75e-07 $layer=POLY_cond $X=1.47 $Y=1.165
+ $X2=1.47 $Y2=0.69
r69 12 14 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=1.435 $Y=1.885
+ $X2=1.435 $Y2=2.46
r70 11 12 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=1.435 $Y=1.795
+ $X2=1.435 $Y2=1.885
r71 10 30 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.435 $Y=1.495
+ $X2=1.435 $Y2=1.33
r72 10 11 116.613 $w=1.8e-07 $l=3e-07 $layer=POLY_cond $X=1.435 $Y=1.495
+ $X2=1.435 $Y2=1.795
r73 9 21 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.04 $Y=1.735
+ $X2=1.04 $Y2=1.81
r74 8 25 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.04 $Y=1.495
+ $X2=1.04 $Y2=1.33
r75 8 9 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=1.04 $Y=1.495 $X2=1.04
+ $Y2=1.735
r76 4 25 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.04 $Y=1.165
+ $X2=1.04 $Y2=1.33
r77 4 6 243.564 $w=1.5e-07 $l=4.75e-07 $layer=POLY_cond $X=1.04 $Y=1.165
+ $X2=1.04 $Y2=0.69
r78 1 19 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.955 $Y=1.885
+ $X2=0.955 $Y2=1.81
r79 1 3 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=0.955 $Y=1.885
+ $X2=0.955 $Y2=2.46
.ends

.subckt PM_SKY130_FD_SC_HS__A222OI_2%B1 3 5 7 8 10 13 15 16 17 18 20 24 27 34
c94 18 0 8.44867e-20 $X=3.235 $Y=2.035
c95 13 0 4.20912e-19 $X=4.4 $Y=0.69
c96 8 0 2.94511e-19 $X=4.385 $Y=1.885
c97 3 0 2.78e-19 $X=2.89 $Y=0.69
r98 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.84
+ $Y=1.635 $X2=2.84 $Y2=1.635
r99 27 34 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.15 $Y=1.635
+ $X2=3.065 $Y2=1.635
r100 27 34 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=3.05 $Y=1.635
+ $X2=3.065 $Y2=1.635
r101 27 32 7.33373 $w=3.28e-07 $l=2.1e-07 $layer=LI1_cond $X=3.05 $Y=1.635
+ $X2=2.84 $Y2=1.635
r102 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.31
+ $Y=1.615 $X2=4.31 $Y2=1.615
r103 21 24 4.1907 $w=3.28e-07 $l=1.2e-07 $layer=LI1_cond $X=4.19 $Y=1.615
+ $X2=4.31 $Y2=1.615
r104 19 21 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.19 $Y=1.78
+ $X2=4.19 $Y2=1.615
r105 19 20 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=4.19 $Y=1.78
+ $X2=4.19 $Y2=1.95
r106 17 20 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.105 $Y=2.035
+ $X2=4.19 $Y2=1.95
r107 17 18 56.7594 $w=1.68e-07 $l=8.7e-07 $layer=LI1_cond $X=4.105 $Y=2.035
+ $X2=3.235 $Y2=2.035
r108 16 18 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.15 $Y=1.95
+ $X2=3.235 $Y2=2.035
r109 15 27 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.15 $Y=1.8
+ $X2=3.15 $Y2=1.635
r110 15 16 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=3.15 $Y=1.8 $X2=3.15
+ $Y2=1.95
r111 11 25 38.5916 $w=2.93e-07 $l=2.05122e-07 $layer=POLY_cond $X=4.4 $Y=1.45
+ $X2=4.31 $Y2=1.615
r112 11 13 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=4.4 $Y=1.45 $X2=4.4
+ $Y2=0.69
r113 8 25 55.8646 $w=2.93e-07 $l=3.05205e-07 $layer=POLY_cond $X=4.385 $Y=1.885
+ $X2=4.31 $Y2=1.615
r114 8 10 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=4.385 $Y=1.885
+ $X2=4.385 $Y2=2.46
r115 5 31 51.2457 $w=3.23e-07 $l=2.91548e-07 $layer=POLY_cond $X=2.945 $Y=1.885
+ $X2=2.855 $Y2=1.635
r116 5 7 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=2.945 $Y=1.885
+ $X2=2.945 $Y2=2.46
r117 1 31 38.5615 $w=3.23e-07 $l=1.81659e-07 $layer=POLY_cond $X=2.89 $Y=1.47
+ $X2=2.855 $Y2=1.635
r118 1 3 399.957 $w=1.5e-07 $l=7.8e-07 $layer=POLY_cond $X=2.89 $Y=1.47 $X2=2.89
+ $Y2=0.69
.ends

.subckt PM_SKY130_FD_SC_HS__A222OI_2%B2 3 6 7 9 11 12 14 15 17 18 24 25
c66 24 0 1.25492e-19 $X=3.57 $Y=1.425
c67 15 0 7.65804e-20 $X=3.97 $Y=1.09
r68 23 25 39.3323 $w=3.37e-07 $l=2.75e-07 $layer=POLY_cond $X=3.57 $Y=1.34
+ $X2=3.845 $Y2=1.34
r69 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.57
+ $Y=1.425 $X2=3.57 $Y2=1.425
r70 21 23 25.0297 $w=3.37e-07 $l=1.75e-07 $layer=POLY_cond $X=3.395 $Y=1.34
+ $X2=3.57 $Y2=1.34
r71 18 24 8.3814 $w=3.28e-07 $l=2.4e-07 $layer=LI1_cond $X=3.57 $Y=1.665
+ $X2=3.57 $Y2=1.425
r72 15 25 17.8783 $w=3.37e-07 $l=3.06186e-07 $layer=POLY_cond $X=3.97 $Y=1.09
+ $X2=3.845 $Y2=1.34
r73 15 17 128.533 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=3.97 $Y=1.09 $X2=3.97
+ $Y2=0.69
r74 12 14 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=3.845 $Y=1.885
+ $X2=3.845 $Y2=2.46
r75 11 12 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=3.845 $Y=1.795
+ $X2=3.845 $Y2=1.885
r76 10 25 17.4215 $w=1.8e-07 $l=2.5e-07 $layer=POLY_cond $X=3.845 $Y=1.59
+ $X2=3.845 $Y2=1.34
r77 10 11 79.6855 $w=1.8e-07 $l=2.05e-07 $layer=POLY_cond $X=3.845 $Y=1.59
+ $X2=3.845 $Y2=1.795
r78 7 9 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=3.395 $Y=1.885
+ $X2=3.395 $Y2=2.46
r79 6 7 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=3.395 $Y=1.795 $X2=3.395
+ $Y2=1.885
r80 5 21 17.4215 $w=1.8e-07 $l=2.5e-07 $layer=POLY_cond $X=3.395 $Y=1.59
+ $X2=3.395 $Y2=1.34
r81 5 6 79.6855 $w=1.8e-07 $l=2.05e-07 $layer=POLY_cond $X=3.395 $Y=1.59
+ $X2=3.395 $Y2=1.795
r82 1 21 10.727 $w=3.37e-07 $l=7.5e-08 $layer=POLY_cond $X=3.32 $Y=1.34
+ $X2=3.395 $Y2=1.34
r83 1 3 292.277 $w=1.5e-07 $l=5.7e-07 $layer=POLY_cond $X=3.32 $Y=1.26 $X2=3.32
+ $Y2=0.69
.ends

.subckt PM_SKY130_FD_SC_HS__A222OI_2%A1 3 5 7 10 12 14 16 17 18 20 25 27 32
c87 18 0 5.31033e-20 $X=5.115 $Y=2.035
c88 5 0 1.51266e-19 $X=4.835 $Y=1.885
r89 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.29
+ $Y=1.615 $X2=6.29 $Y2=1.615
r90 27 32 10.1275 $w=3.28e-07 $l=2.9e-07 $layer=LI1_cond $X=6 $Y=1.615 $X2=6.29
+ $Y2=1.615
r91 27 33 1.04768 $w=3.28e-07 $l=3e-08 $layer=LI1_cond $X=6 $Y=1.615 $X2=5.97
+ $Y2=1.615
r92 22 25 6.28605 $w=3.28e-07 $l=1.8e-07 $layer=LI1_cond $X=4.85 $Y=1.615
+ $X2=5.03 $Y2=1.615
r93 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.85
+ $Y=1.615 $X2=4.85 $Y2=1.615
r94 19 33 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.97 $Y=1.78
+ $X2=5.97 $Y2=1.615
r95 19 20 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=5.97 $Y=1.78
+ $X2=5.97 $Y2=1.95
r96 17 20 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.885 $Y=2.035
+ $X2=5.97 $Y2=1.95
r97 17 18 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=5.885 $Y=2.035
+ $X2=5.115 $Y2=2.035
r98 16 18 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.03 $Y=1.95
+ $X2=5.115 $Y2=2.035
r99 15 25 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.03 $Y=1.78
+ $X2=5.03 $Y2=1.615
r100 15 16 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=5.03 $Y=1.78
+ $X2=5.03 $Y2=1.95
r101 12 31 55.8646 $w=2.93e-07 $l=3.05205e-07 $layer=POLY_cond $X=6.215 $Y=1.885
+ $X2=6.29 $Y2=1.615
r102 12 14 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=6.215 $Y=1.885
+ $X2=6.215 $Y2=2.46
r103 8 31 38.5916 $w=2.93e-07 $l=2.05122e-07 $layer=POLY_cond $X=6.2 $Y=1.45
+ $X2=6.29 $Y2=1.615
r104 8 10 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=6.2 $Y=1.45 $X2=6.2
+ $Y2=0.69
r105 5 23 55.8646 $w=2.93e-07 $l=2.77399e-07 $layer=POLY_cond $X=4.835 $Y=1.885
+ $X2=4.85 $Y2=1.615
r106 5 7 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=4.835 $Y=1.885
+ $X2=4.835 $Y2=2.46
r107 1 23 38.5916 $w=2.93e-07 $l=1.74714e-07 $layer=POLY_cond $X=4.83 $Y=1.45
+ $X2=4.85 $Y2=1.615
r108 1 3 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=4.83 $Y=1.45 $X2=4.83
+ $Y2=0.69
.ends

.subckt PM_SKY130_FD_SC_HS__A222OI_2%A2 1 3 6 8 10 13 15 22
r56 22 23 0.617949 $w=3.9e-07 $l=5e-09 $layer=POLY_cond $X=5.765 $Y=1.667
+ $X2=5.77 $Y2=1.667
r57 20 22 36.459 $w=3.9e-07 $l=2.95e-07 $layer=POLY_cond $X=5.47 $Y=1.667
+ $X2=5.765 $Y2=1.667
r58 18 20 17.3026 $w=3.9e-07 $l=1.4e-07 $layer=POLY_cond $X=5.33 $Y=1.667
+ $X2=5.47 $Y2=1.667
r59 17 18 1.85385 $w=3.9e-07 $l=1.5e-08 $layer=POLY_cond $X=5.315 $Y=1.667
+ $X2=5.33 $Y2=1.667
r60 15 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.47
+ $Y=1.615 $X2=5.47 $Y2=1.615
r61 11 23 25.2441 $w=1.5e-07 $l=2.17e-07 $layer=POLY_cond $X=5.77 $Y=1.45
+ $X2=5.77 $Y2=1.667
r62 11 13 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=5.77 $Y=1.45
+ $X2=5.77 $Y2=0.69
r63 8 22 25.2441 $w=1.5e-07 $l=2.18e-07 $layer=POLY_cond $X=5.765 $Y=1.885
+ $X2=5.765 $Y2=1.667
r64 8 10 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=5.765 $Y=1.885
+ $X2=5.765 $Y2=2.46
r65 4 18 25.2441 $w=1.5e-07 $l=2.17e-07 $layer=POLY_cond $X=5.33 $Y=1.45
+ $X2=5.33 $Y2=1.667
r66 4 6 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=5.33 $Y=1.45 $X2=5.33
+ $Y2=0.69
r67 1 17 25.2441 $w=1.5e-07 $l=2.18e-07 $layer=POLY_cond $X=5.315 $Y=1.885
+ $X2=5.315 $Y2=1.667
r68 1 3 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=5.315 $Y=1.885
+ $X2=5.315 $Y2=2.46
.ends

.subckt PM_SKY130_FD_SC_HS__A222OI_2%Y 1 2 3 4 5 6 7 23 25 26 30 32 37 40 42 43
+ 46 48 52 55 57 58 61 67 68 69
c148 48 0 1.28994e-19 $X=6.32 $Y=1.195
c149 42 0 7.65804e-20 $X=4.45 $Y=1.005
r150 68 69 15.2287 $w=2.78e-07 $l=3.7e-07 $layer=LI1_cond $X=0.225 $Y=2.405
+ $X2=0.225 $Y2=2.775
r151 68 73 9.4665 $w=2.78e-07 $l=2.3e-07 $layer=LI1_cond $X=0.225 $Y=2.405
+ $X2=0.225 $Y2=2.175
r152 67 73 4.06715 $w=2.25e-07 $l=1.28e-07 $layer=LI1_cond $X=0.225 $Y=2.047
+ $X2=0.225 $Y2=2.175
r153 57 58 9.38152 $w=2.13e-07 $l=1.65e-07 $layer=LI1_cond $X=1.255 $Y=0.887
+ $X2=1.09 $Y2=0.887
r154 50 52 26.3732 $w=2.58e-07 $l=5.95e-07 $layer=LI1_cond $X=6.45 $Y=1.11
+ $X2=6.45 $Y2=0.515
r155 49 65 3.33486 $w=1.7e-07 $l=1.33e-07 $layer=LI1_cond $X=4.715 $Y=1.195
+ $X2=4.582 $Y2=1.195
r156 48 50 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=6.32 $Y=1.195
+ $X2=6.45 $Y2=1.11
r157 48 49 104.711 $w=1.68e-07 $l=1.605e-06 $layer=LI1_cond $X=6.32 $Y=1.195
+ $X2=4.715 $Y2=1.195
r158 44 46 17.6128 $w=2.63e-07 $l=4.05e-07 $layer=LI1_cond $X=4.582 $Y=0.92
+ $X2=4.582 $Y2=0.515
r159 43 63 8.98989 $w=2.97e-07 $l=2.11069e-07 $layer=LI1_cond $X=2.84 $Y=1.005
+ $X2=2.675 $Y2=1.11
r160 42 65 8.2628 $w=2.63e-07 $l=1.9e-07 $layer=LI1_cond $X=4.582 $Y=1.005
+ $X2=4.582 $Y2=1.195
r161 42 44 3.69652 $w=2.63e-07 $l=8.5e-08 $layer=LI1_cond $X=4.582 $Y=1.005
+ $X2=4.582 $Y2=0.92
r162 42 43 105.037 $w=1.68e-07 $l=1.61e-06 $layer=LI1_cond $X=4.45 $Y=1.005
+ $X2=2.84 $Y2=1.005
r163 38 63 0.0633028 $w=3.3e-07 $l=1.9e-07 $layer=LI1_cond $X=2.675 $Y=0.92
+ $X2=2.675 $Y2=1.11
r164 38 40 14.1436 $w=3.28e-07 $l=4.05e-07 $layer=LI1_cond $X=2.675 $Y=0.92
+ $X2=2.675 $Y2=0.515
r165 37 61 2.96976 $w=3.2e-07 $l=1.8775e-07 $layer=LI1_cond $X=2.38 $Y=2.005
+ $X2=2.23 $Y2=2.09
r166 36 63 12.1178 $w=2.97e-07 $l=3.78253e-07 $layer=LI1_cond $X=2.38 $Y=1.3
+ $X2=2.675 $Y2=1.11
r167 36 37 45.9947 $w=1.68e-07 $l=7.05e-07 $layer=LI1_cond $X=2.38 $Y=1.3
+ $X2=2.38 $Y2=2.005
r168 33 55 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.325 $Y=2.09
+ $X2=1.195 $Y2=2.09
r169 32 61 3.69268 $w=1.7e-07 $l=2.35e-07 $layer=LI1_cond $X=1.995 $Y=2.09
+ $X2=2.23 $Y2=2.09
r170 32 33 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.995 $Y=2.09
+ $X2=1.325 $Y2=2.09
r171 28 55 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=1.195 $Y=2.175
+ $X2=1.195 $Y2=2.09
r172 28 30 17.5083 $w=2.58e-07 $l=3.95e-07 $layer=LI1_cond $X=1.195 $Y=2.175
+ $X2=1.195 $Y2=2.57
r173 27 67 2.36881 $w=1.7e-07 $l=1.60062e-07 $layer=LI1_cond $X=0.365 $Y=2.09
+ $X2=0.225 $Y2=2.047
r174 26 55 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.065 $Y=2.09
+ $X2=1.195 $Y2=2.09
r175 26 27 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=1.065 $Y=2.09
+ $X2=0.365 $Y2=2.09
r176 25 58 54.4759 $w=1.68e-07 $l=8.35e-07 $layer=LI1_cond $X=0.255 $Y=0.91
+ $X2=1.09 $Y2=0.91
r177 23 67 4.06715 $w=2.25e-07 $l=1.52033e-07 $layer=LI1_cond $X=0.17 $Y=1.92
+ $X2=0.225 $Y2=2.047
r178 22 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.17 $Y=0.995
+ $X2=0.255 $Y2=0.91
r179 22 23 60.3476 $w=1.68e-07 $l=9.25e-07 $layer=LI1_cond $X=0.17 $Y=0.995
+ $X2=0.17 $Y2=1.92
r180 7 61 300 $w=1.7e-07 $l=2.93428e-07 $layer=licon1_PDIFF $count=2 $X=1.96
+ $Y=1.96 $X2=2.16 $Y2=2.17
r181 6 55 600 $w=1.7e-07 $l=2.20624e-07 $layer=licon1_PDIFF $count=1 $X=1.03
+ $Y=1.96 $X2=1.195 $Y2=2.09
r182 6 30 600 $w=1.7e-07 $l=6.87568e-07 $layer=licon1_PDIFF $count=1 $X=1.03
+ $Y=1.96 $X2=1.195 $Y2=2.57
r183 5 67 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.96 $X2=0.28 $Y2=2.105
r184 5 69 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.96 $X2=0.28 $Y2=2.815
r185 4 52 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=6.275
+ $Y=0.37 $X2=6.415 $Y2=0.515
r186 3 46 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=4.475
+ $Y=0.37 $X2=4.615 $Y2=0.515
r187 2 40 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=2.53
+ $Y=0.37 $X2=2.675 $Y2=0.515
r188 1 57 182 $w=1.7e-07 $l=5.60647e-07 $layer=licon1_NDIFF $count=1 $X=1.115
+ $Y=0.37 $X2=1.255 $Y2=0.865
.ends

.subckt PM_SKY130_FD_SC_HS__A222OI_2%A_116_392# 1 2 3 4 15 17 18 21 27 29 32 33
r59 31 33 5.06676 $w=4.43e-07 $l=1.65e-07 $layer=LI1_cond $X=3.17 $Y=2.852
+ $X2=3.335 $Y2=2.852
r60 31 32 8.86124 $w=4.43e-07 $l=1.65e-07 $layer=LI1_cond $X=3.17 $Y=2.852
+ $X2=3.005 $Y2=2.852
r61 27 33 27.2396 $w=3.28e-07 $l=7.8e-07 $layer=LI1_cond $X=4.115 $Y=2.815
+ $X2=3.335 $Y2=2.815
r62 24 29 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.825 $Y=2.99
+ $X2=1.66 $Y2=2.99
r63 24 32 76.984 $w=1.68e-07 $l=1.18e-06 $layer=LI1_cond $X=1.825 $Y=2.99
+ $X2=3.005 $Y2=2.99
r64 19 29 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.66 $Y=2.905
+ $X2=1.66 $Y2=2.99
r65 19 21 16.5882 $w=3.28e-07 $l=4.75e-07 $layer=LI1_cond $X=1.66 $Y=2.905
+ $X2=1.66 $Y2=2.43
r66 17 29 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.495 $Y=2.99
+ $X2=1.66 $Y2=2.99
r67 17 18 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=1.495 $Y=2.99
+ $X2=0.895 $Y2=2.99
r68 13 18 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.73 $Y=2.905
+ $X2=0.895 $Y2=2.99
r69 13 15 16.5882 $w=3.28e-07 $l=4.75e-07 $layer=LI1_cond $X=0.73 $Y=2.905
+ $X2=0.73 $Y2=2.43
r70 4 27 600 $w=1.7e-07 $l=9.47497e-07 $layer=licon1_PDIFF $count=1 $X=3.92
+ $Y=1.96 $X2=4.115 $Y2=2.815
r71 3 31 600 $w=1.7e-07 $l=9.16938e-07 $layer=licon1_PDIFF $count=1 $X=3.02
+ $Y=1.96 $X2=3.17 $Y2=2.805
r72 2 21 300 $w=1.7e-07 $l=5.39815e-07 $layer=licon1_PDIFF $count=2 $X=1.51
+ $Y=1.96 $X2=1.66 $Y2=2.43
r73 1 15 300 $w=1.7e-07 $l=5.39815e-07 $layer=licon1_PDIFF $count=2 $X=0.58
+ $Y=1.96 $X2=0.73 $Y2=2.43
.ends

.subckt PM_SKY130_FD_SC_HS__A222OI_2%A_515_392# 1 2 3 4 5 18 22 24 30 34 38 40
+ 44 48 50 52 54
c78 50 0 3.20286e-19 $X=4.61 $Y=2.465
r79 42 54 3.48018 $w=3e-07 $l=9.5e-08 $layer=LI1_cond $X=6.44 $Y=2.29 $X2=6.44
+ $Y2=2.385
r80 42 44 7.15912 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=6.44 $Y=2.29
+ $X2=6.44 $Y2=2.085
r81 41 52 6.03773 $w=1.9e-07 $l=1.15e-07 $layer=LI1_cond $X=5.655 $Y=2.385
+ $X2=5.54 $Y2=2.385
r82 40 54 3.02843 $w=1.9e-07 $l=1.65e-07 $layer=LI1_cond $X=6.275 $Y=2.385
+ $X2=6.44 $Y2=2.385
r83 40 41 36.1914 $w=1.88e-07 $l=6.2e-07 $layer=LI1_cond $X=6.275 $Y=2.385
+ $X2=5.655 $Y2=2.385
r84 36 52 0.664496 $w=2.3e-07 $l=9.5e-08 $layer=LI1_cond $X=5.54 $Y=2.48
+ $X2=5.54 $Y2=2.385
r85 36 38 16.7856 $w=2.28e-07 $l=3.35e-07 $layer=LI1_cond $X=5.54 $Y=2.48
+ $X2=5.54 $Y2=2.815
r86 35 50 4.39947 $w=1.9e-07 $l=3.745e-07 $layer=LI1_cond $X=4.775 $Y=2.385
+ $X2=4.445 $Y2=2.29
r87 34 52 6.03773 $w=1.9e-07 $l=1.15e-07 $layer=LI1_cond $X=5.425 $Y=2.385
+ $X2=5.54 $Y2=2.385
r88 34 35 37.9426 $w=1.88e-07 $l=6.5e-07 $layer=LI1_cond $X=5.425 $Y=2.385
+ $X2=4.775 $Y2=2.385
r89 28 50 1.88912 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=4.61 $Y=2.29
+ $X2=4.445 $Y2=2.29
r90 28 30 6.11144 $w=3.28e-07 $l=1.75e-07 $layer=LI1_cond $X=4.61 $Y=2.29
+ $X2=4.61 $Y2=2.115
r91 25 48 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.805 $Y=2.375
+ $X2=2.72 $Y2=2.375
r92 25 27 53.1711 $w=1.68e-07 $l=8.15e-07 $layer=LI1_cond $X=2.805 $Y=2.375
+ $X2=3.62 $Y2=2.375
r93 24 50 4.39947 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.445 $Y=2.375
+ $X2=4.445 $Y2=2.29
r94 24 27 53.8235 $w=1.68e-07 $l=8.25e-07 $layer=LI1_cond $X=4.445 $Y=2.375
+ $X2=3.62 $Y2=2.375
r95 20 48 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.72 $Y=2.46 $X2=2.72
+ $Y2=2.375
r96 20 22 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=2.72 $Y=2.46
+ $X2=2.72 $Y2=2.57
r97 16 48 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.72 $Y=2.29 $X2=2.72
+ $Y2=2.375
r98 16 18 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=2.72 $Y=2.29
+ $X2=2.72 $Y2=2.135
r99 5 54 300 $w=1.7e-07 $l=5.65044e-07 $layer=licon1_PDIFF $count=2 $X=6.29
+ $Y=1.96 $X2=6.44 $Y2=2.455
r100 5 44 600 $w=1.7e-07 $l=2.03101e-07 $layer=licon1_PDIFF $count=1 $X=6.29
+ $Y=1.96 $X2=6.44 $Y2=2.085
r101 4 52 600 $w=1.7e-07 $l=4.94343e-07 $layer=licon1_PDIFF $count=1 $X=5.39
+ $Y=1.96 $X2=5.54 $Y2=2.385
r102 4 38 600 $w=1.7e-07 $l=9.26971e-07 $layer=licon1_PDIFF $count=1 $X=5.39
+ $Y=1.96 $X2=5.54 $Y2=2.815
r103 3 50 300 $w=1.7e-07 $l=5.7513e-07 $layer=licon1_PDIFF $count=2 $X=4.46
+ $Y=1.96 $X2=4.61 $Y2=2.465
r104 3 30 600 $w=1.7e-07 $l=2.17428e-07 $layer=licon1_PDIFF $count=1 $X=4.46
+ $Y=1.96 $X2=4.61 $Y2=2.115
r105 2 27 600 $w=1.7e-07 $l=4.84226e-07 $layer=licon1_PDIFF $count=1 $X=3.47
+ $Y=1.96 $X2=3.62 $Y2=2.375
r106 1 22 600 $w=1.7e-07 $l=6.78638e-07 $layer=licon1_PDIFF $count=1 $X=2.575
+ $Y=1.96 $X2=2.72 $Y2=2.57
r107 1 18 600 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=2.575
+ $Y=1.96 $X2=2.72 $Y2=2.135
.ends

.subckt PM_SKY130_FD_SC_HS__A222OI_2%VPWR 1 2 9 13 15 17 25 32 33 36 39
r71 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r72 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r73 33 40 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=3.33 $X2=6
+ $Y2=3.33
r74 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r75 30 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.155 $Y=3.33
+ $X2=5.99 $Y2=3.33
r76 30 32 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=6.155 $Y=3.33
+ $X2=6.48 $Y2=3.33
r77 29 40 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=3.33 $X2=6
+ $Y2=3.33
r78 29 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=5.04 $Y2=3.33
r79 28 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r80 26 36 9.14399 $w=1.7e-07 $l=1.8e-07 $layer=LI1_cond $X=5.255 $Y=3.33
+ $X2=5.075 $Y2=3.33
r81 26 28 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=5.255 $Y=3.33
+ $X2=5.52 $Y2=3.33
r82 25 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.825 $Y=3.33
+ $X2=5.99 $Y2=3.33
r83 25 28 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=5.825 $Y=3.33
+ $X2=5.52 $Y2=3.33
r84 24 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=5.04 $Y2=3.33
r85 23 24 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r86 19 23 281.84 $w=1.68e-07 $l=4.32e-06 $layer=LI1_cond $X=0.24 $Y=3.33
+ $X2=4.56 $Y2=3.33
r87 19 20 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r88 17 36 9.14399 $w=1.7e-07 $l=1.8e-07 $layer=LI1_cond $X=4.895 $Y=3.33
+ $X2=5.075 $Y2=3.33
r89 17 23 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=4.895 $Y=3.33
+ $X2=4.56 $Y2=3.33
r90 15 24 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=3.36 $Y=3.33
+ $X2=4.56 $Y2=3.33
r91 15 20 0.869652 $w=4.9e-07 $l=3.12e-06 $layer=MET1_cond $X=3.36 $Y=3.33
+ $X2=0.24 $Y2=3.33
r92 11 39 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.99 $Y=3.245
+ $X2=5.99 $Y2=3.33
r93 11 13 16.7628 $w=3.28e-07 $l=4.8e-07 $layer=LI1_cond $X=5.99 $Y=3.245
+ $X2=5.99 $Y2=2.765
r94 7 36 1.16013 $w=3.6e-07 $l=8.5e-08 $layer=LI1_cond $X=5.075 $Y=3.245
+ $X2=5.075 $Y2=3.33
r95 7 9 15.3659 $w=3.58e-07 $l=4.8e-07 $layer=LI1_cond $X=5.075 $Y=3.245
+ $X2=5.075 $Y2=2.765
r96 2 13 600 $w=1.7e-07 $l=8.76798e-07 $layer=licon1_PDIFF $count=1 $X=5.84
+ $Y=1.96 $X2=5.99 $Y2=2.765
r97 1 9 600 $w=1.7e-07 $l=8.83657e-07 $layer=licon1_PDIFF $count=1 $X=4.91
+ $Y=1.96 $X2=5.075 $Y2=2.765
.ends

.subckt PM_SKY130_FD_SC_HS__A222OI_2%VGND 1 2 3 4 13 15 19 23 25 27 35 40 50 51
+ 57 61 67
r89 67 68 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r90 61 64 9.60369 $w=3.88e-07 $l=3.25e-07 $layer=LI1_cond $X=3.645 $Y=0
+ $X2=3.645 $Y2=0.325
r91 61 62 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r92 57 58 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r93 54 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r94 51 68 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.48 $Y=0 $X2=5.52
+ $Y2=0
r95 50 51 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.48 $Y=0 $X2=6.48
+ $Y2=0
r96 48 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.715 $Y=0 $X2=5.55
+ $Y2=0
r97 48 50 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=5.715 $Y=0 $X2=6.48
+ $Y2=0
r98 47 68 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=5.52
+ $Y2=0
r99 46 47 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r100 44 47 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=5.04
+ $Y2=0
r101 44 62 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=3.6
+ $Y2=0
r102 43 46 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=4.08 $Y=0 $X2=5.04
+ $Y2=0
r103 43 44 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r104 41 61 5.6248 $w=1.7e-07 $l=1.95e-07 $layer=LI1_cond $X=3.84 $Y=0 $X2=3.645
+ $Y2=0
r105 41 43 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=3.84 $Y=0 $X2=4.08
+ $Y2=0
r106 40 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.385 $Y=0 $X2=5.55
+ $Y2=0
r107 40 46 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=5.385 $Y=0 $X2=5.04
+ $Y2=0
r108 39 58 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=2.16
+ $Y2=0
r109 38 39 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r110 36 57 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.28 $Y=0 $X2=2.115
+ $Y2=0
r111 36 38 54.8021 $w=1.68e-07 $l=8.4e-07 $layer=LI1_cond $X=2.28 $Y=0 $X2=3.12
+ $Y2=0
r112 35 61 5.6248 $w=1.7e-07 $l=1.95e-07 $layer=LI1_cond $X=3.45 $Y=0 $X2=3.645
+ $Y2=0
r113 35 38 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=3.45 $Y=0 $X2=3.12
+ $Y2=0
r114 34 58 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r115 33 34 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r116 31 34 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r117 31 55 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r118 30 33 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r119 30 31 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r120 28 54 5.06789 $w=1.7e-07 $l=2.4e-07 $layer=LI1_cond $X=0.48 $Y=0 $X2=0.24
+ $Y2=0
r121 28 30 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=0.48 $Y=0 $X2=0.72
+ $Y2=0
r122 27 57 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.95 $Y=0 $X2=2.115
+ $Y2=0
r123 27 33 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=1.95 $Y=0 $X2=1.68
+ $Y2=0
r124 25 62 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=3.36 $Y=0 $X2=3.6
+ $Y2=0
r125 25 39 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=3.36 $Y=0
+ $X2=3.12 $Y2=0
r126 21 67 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.55 $Y=0.085
+ $X2=5.55 $Y2=0
r127 21 23 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=5.55 $Y=0.085
+ $X2=5.55 $Y2=0.515
r128 17 57 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.115 $Y=0.085
+ $X2=2.115 $Y2=0
r129 17 19 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=2.115 $Y=0.085
+ $X2=2.115 $Y2=0.515
r130 13 54 2.9985 $w=3.65e-07 $l=1.09864e-07 $layer=LI1_cond $X=0.297 $Y=0.085
+ $X2=0.24 $Y2=0
r131 13 15 12.7874 $w=3.63e-07 $l=4.05e-07 $layer=LI1_cond $X=0.297 $Y=0.085
+ $X2=0.297 $Y2=0.49
r132 4 23 182 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=1 $X=5.405
+ $Y=0.37 $X2=5.55 $Y2=0.515
r133 3 64 182 $w=1.7e-07 $l=2.7157e-07 $layer=licon1_NDIFF $count=1 $X=3.395
+ $Y=0.37 $X2=3.645 $Y2=0.325
r134 2 19 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.975
+ $Y=0.37 $X2=2.115 $Y2=0.515
r135 1 15 182 $w=1.7e-07 $l=2.20907e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.345 $X2=0.295 $Y2=0.49
.ends

.subckt PM_SKY130_FD_SC_HS__A222OI_2%A_137_74# 1 2 7
r13 11 13 4.96172 $w=1.88e-07 $l=8.5e-08 $layer=LI1_cond $X=1.685 $Y=0.61
+ $X2=1.685 $Y2=0.695
r14 7 11 7.03324 $w=2.6e-07 $l=1.71026e-07 $layer=LI1_cond $X=1.59 $Y=0.48
+ $X2=1.685 $Y2=0.61
r15 7 9 33.9084 $w=2.58e-07 $l=7.65e-07 $layer=LI1_cond $X=1.59 $Y=0.48
+ $X2=0.825 $Y2=0.48
r16 2 13 182 $w=1.7e-07 $l=3.88748e-07 $layer=licon1_NDIFF $count=1 $X=1.545
+ $Y=0.37 $X2=1.685 $Y2=0.695
r17 1 9 182 $w=1.7e-07 $l=2.08567e-07 $layer=licon1_NDIFF $count=1 $X=0.685
+ $Y=0.37 $X2=0.825 $Y2=0.52
.ends

.subckt PM_SKY130_FD_SC_HS__A222OI_2%A_593_74# 1 2 7 10 15
c26 15 0 1.66006e-19 $X=4.185 $Y=0.55
c27 10 0 1.66006e-19 $X=3.105 $Y=0.55
r28 15 17 5.30124 $w=2.48e-07 $l=1.15e-07 $layer=LI1_cond $X=4.145 $Y=0.55
+ $X2=4.145 $Y2=0.665
r29 10 12 5.30124 $w=2.48e-07 $l=1.15e-07 $layer=LI1_cond $X=3.145 $Y=0.55
+ $X2=3.145 $Y2=0.665
r30 8 12 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.27 $Y=0.665
+ $X2=3.145 $Y2=0.665
r31 7 17 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.02 $Y=0.665
+ $X2=4.145 $Y2=0.665
r32 7 8 48.9305 $w=1.68e-07 $l=7.5e-07 $layer=LI1_cond $X=4.02 $Y=0.665 $X2=3.27
+ $Y2=0.665
r33 2 15 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=4.045 $Y=0.37
+ $X2=4.185 $Y2=0.55
r34 1 10 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=2.965 $Y=0.37
+ $X2=3.105 $Y2=0.55
.ends

.subckt PM_SKY130_FD_SC_HS__A222OI_2%A_981_74# 1 2 9 11 12 13 15
c24 9 0 1.25912e-19 $X=5.05 $Y=0.495
r25 13 18 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.025 $Y=0.77
+ $X2=6.025 $Y2=0.855
r26 13 15 12.6769 $w=2.48e-07 $l=2.75e-07 $layer=LI1_cond $X=6.025 $Y=0.77
+ $X2=6.025 $Y2=0.495
r27 11 18 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.9 $Y=0.855
+ $X2=6.025 $Y2=0.855
r28 11 12 44.6898 $w=1.68e-07 $l=6.85e-07 $layer=LI1_cond $X=5.9 $Y=0.855
+ $X2=5.215 $Y2=0.855
r29 7 12 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=5.05 $Y=0.77
+ $X2=5.215 $Y2=0.855
r30 7 9 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=5.05 $Y=0.77 $X2=5.05
+ $Y2=0.495
r31 2 18 182 $w=1.7e-07 $l=5.50568e-07 $layer=licon1_NDIFF $count=1 $X=5.845
+ $Y=0.37 $X2=5.985 $Y2=0.855
r32 2 15 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=5.845
+ $Y=0.37 $X2=5.985 $Y2=0.495
r33 1 9 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=4.905
+ $Y=0.37 $X2=5.05 $Y2=0.495
.ends

