* File: sky130_fd_sc_hs__o31a_1.pxi.spice
* Created: Thu Aug 27 21:02:28 2020
* 
x_PM_SKY130_FD_SC_HS__O31A_1%A_84_48# N_A_84_48#_M1004_d N_A_84_48#_M1001_d
+ N_A_84_48#_M1009_g N_A_84_48#_c_61_n N_A_84_48#_M1002_g N_A_84_48#_c_62_n
+ N_A_84_48#_c_77_p N_A_84_48#_c_111_p N_A_84_48#_c_69_n N_A_84_48#_c_70_n
+ N_A_84_48#_c_63_n N_A_84_48#_c_64_n N_A_84_48#_c_65_n N_A_84_48#_c_88_p
+ N_A_84_48#_c_66_n PM_SKY130_FD_SC_HS__O31A_1%A_84_48#
x_PM_SKY130_FD_SC_HS__O31A_1%A1 N_A1_M1008_g N_A1_c_135_n N_A1_M1000_g A1
+ N_A1_c_136_n PM_SKY130_FD_SC_HS__O31A_1%A1
x_PM_SKY130_FD_SC_HS__O31A_1%A2 N_A2_M1006_g N_A2_c_168_n N_A2_M1007_g A2
+ N_A2_c_169_n PM_SKY130_FD_SC_HS__O31A_1%A2
x_PM_SKY130_FD_SC_HS__O31A_1%A3 N_A3_c_197_n N_A3_M1001_g N_A3_M1003_g A3
+ N_A3_c_199_n PM_SKY130_FD_SC_HS__O31A_1%A3
x_PM_SKY130_FD_SC_HS__O31A_1%B1 N_B1_c_229_n N_B1_M1005_g N_B1_M1004_g B1
+ N_B1_c_231_n PM_SKY130_FD_SC_HS__O31A_1%B1
x_PM_SKY130_FD_SC_HS__O31A_1%X N_X_M1009_s N_X_M1002_s N_X_c_255_n N_X_c_256_n X
+ X X X N_X_c_257_n PM_SKY130_FD_SC_HS__O31A_1%X
x_PM_SKY130_FD_SC_HS__O31A_1%VPWR N_VPWR_M1002_d N_VPWR_M1005_d N_VPWR_c_280_n
+ N_VPWR_c_281_n N_VPWR_c_282_n N_VPWR_c_283_n VPWR N_VPWR_c_284_n
+ N_VPWR_c_285_n N_VPWR_c_279_n N_VPWR_c_287_n PM_SKY130_FD_SC_HS__O31A_1%VPWR
x_PM_SKY130_FD_SC_HS__O31A_1%VGND N_VGND_M1009_d N_VGND_M1006_d N_VGND_c_318_n
+ N_VGND_c_319_n N_VGND_c_320_n N_VGND_c_321_n VGND N_VGND_c_322_n
+ N_VGND_c_323_n N_VGND_c_324_n N_VGND_c_325_n PM_SKY130_FD_SC_HS__O31A_1%VGND
x_PM_SKY130_FD_SC_HS__O31A_1%A_230_94# N_A_230_94#_M1008_d N_A_230_94#_M1003_d
+ N_A_230_94#_c_357_n N_A_230_94#_c_358_n N_A_230_94#_c_359_n
+ N_A_230_94#_c_360_n PM_SKY130_FD_SC_HS__O31A_1%A_230_94#
cc_1 VNB N_A_84_48#_M1009_g 0.030112f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_2 VNB N_A_84_48#_c_61_n 0.0344604f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=1.765
cc_3 VNB N_A_84_48#_c_62_n 2.46719e-19 $X=-0.19 $Y=-0.245 $X2=0.71 $Y2=1.95
cc_4 VNB N_A_84_48#_c_63_n 0.0233423f $X=-0.19 $Y=-0.245 $X2=3.08 $Y2=0.615
cc_5 VNB N_A_84_48#_c_64_n 0.0253498f $X=-0.19 $Y=-0.245 $X2=3.17 $Y2=1.95
cc_6 VNB N_A_84_48#_c_65_n 0.0026276f $X=-0.19 $Y=-0.245 $X2=0.71 $Y2=1.485
cc_7 VNB N_A_84_48#_c_66_n 0.0137511f $X=-0.19 $Y=-0.245 $X2=3.085 $Y2=1.13
cc_8 VNB N_A1_M1008_g 0.026484f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A1_c_135_n 0.0243423f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A1_c_136_n 0.00495499f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=2.4
cc_11 VNB N_A2_M1006_g 0.0247917f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A2_c_168_n 0.0338774f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A2_c_169_n 0.00206174f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=2.4
cc_14 VNB N_A3_c_197_n 0.0263889f $X=-0.19 $Y=-0.245 $X2=2.87 $Y2=0.47
cc_15 VNB N_A3_M1003_g 0.0277067f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A3_c_199_n 0.00182951f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=2.4
cc_17 VNB N_B1_c_229_n 0.0266141f $X=-0.19 $Y=-0.245 $X2=2.87 $Y2=0.47
cc_18 VNB N_B1_M1004_g 0.0287531f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_B1_c_231_n 0.00535768f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=2.4
cc_20 VNB N_X_c_255_n 0.0265914f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_21 VNB N_X_c_256_n 0.0139041f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=2.4
cc_22 VNB N_X_c_257_n 0.0249534f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.485
cc_23 VNB N_VPWR_c_279_n 0.143779f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.485
cc_24 VNB N_VGND_c_318_n 0.0212254f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_25 VNB N_VGND_c_319_n 0.0189386f $X=-0.19 $Y=-0.245 $X2=0.71 $Y2=1.95
cc_26 VNB N_VGND_c_320_n 0.023893f $X=-0.19 $Y=-0.245 $X2=2.36 $Y2=2.12
cc_27 VNB N_VGND_c_321_n 0.00702069f $X=-0.19 $Y=-0.245 $X2=2.36 $Y2=2.375
cc_28 VNB N_VGND_c_322_n 0.0189171f $X=-0.19 $Y=-0.245 $X2=2.36 $Y2=2.715
cc_29 VNB N_VGND_c_323_n 0.0370094f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_324_n 0.227175f $X=-0.19 $Y=-0.245 $X2=0.71 $Y2=1.485
cc_31 VNB N_VGND_c_325_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=2.36 $Y2=2.035
cc_32 VNB N_A_230_94#_c_357_n 0.00335993f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_33 VNB N_A_230_94#_c_358_n 0.0191055f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=1.765
cc_34 VNB N_A_230_94#_c_359_n 0.0070898f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=2.4
cc_35 VNB N_A_230_94#_c_360_n 0.00330195f $X=-0.19 $Y=-0.245 $X2=0.71 $Y2=1.95
cc_36 VPB N_A_84_48#_c_61_n 0.0298916f $X=-0.19 $Y=1.66 $X2=0.515 $Y2=1.765
cc_37 VPB N_A_84_48#_c_62_n 0.00288338f $X=-0.19 $Y=1.66 $X2=0.71 $Y2=1.95
cc_38 VPB N_A_84_48#_c_69_n 0.00500809f $X=-0.19 $Y=1.66 $X2=2.36 $Y2=2.375
cc_39 VPB N_A_84_48#_c_70_n 0.0082934f $X=-0.19 $Y=1.66 $X2=3.085 $Y2=2.035
cc_40 VPB N_A_84_48#_c_64_n 0.0125422f $X=-0.19 $Y=1.66 $X2=3.17 $Y2=1.95
cc_41 VPB N_A1_c_135_n 0.0273748f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_42 VPB N_A1_c_136_n 0.00329379f $X=-0.19 $Y=1.66 $X2=0.515 $Y2=2.4
cc_43 VPB N_A2_c_168_n 0.0213052f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_44 VPB N_A2_c_169_n 0.0032264f $X=-0.19 $Y=1.66 $X2=0.515 $Y2=2.4
cc_45 VPB N_A3_c_197_n 0.0285229f $X=-0.19 $Y=1.66 $X2=2.87 $Y2=0.47
cc_46 VPB N_A3_c_199_n 0.00238263f $X=-0.19 $Y=1.66 $X2=0.515 $Y2=2.4
cc_47 VPB N_B1_c_229_n 0.0299966f $X=-0.19 $Y=1.66 $X2=2.87 $Y2=0.47
cc_48 VPB N_B1_c_231_n 0.00374395f $X=-0.19 $Y=1.66 $X2=0.515 $Y2=2.4
cc_49 VPB X 0.0143414f $X=-0.19 $Y=1.66 $X2=0.71 $Y2=1.65
cc_50 VPB X 0.0420589f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_51 VPB N_X_c_257_n 0.00757469f $X=-0.19 $Y=1.66 $X2=0.59 $Y2=1.485
cc_52 VPB N_VPWR_c_280_n 0.0165678f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.74
cc_53 VPB N_VPWR_c_281_n 0.0294894f $X=-0.19 $Y=1.66 $X2=0.515 $Y2=2.4
cc_54 VPB N_VPWR_c_282_n 0.0501782f $X=-0.19 $Y=1.66 $X2=2.195 $Y2=2.035
cc_55 VPB N_VPWR_c_283_n 0.00603306f $X=-0.19 $Y=1.66 $X2=0.795 $Y2=2.035
cc_56 VPB N_VPWR_c_284_n 0.0191572f $X=-0.19 $Y=1.66 $X2=2.36 $Y2=2.375
cc_57 VPB N_VPWR_c_285_n 0.0120081f $X=-0.19 $Y=1.66 $X2=0.59 $Y2=1.485
cc_58 VPB N_VPWR_c_279_n 0.100285f $X=-0.19 $Y=1.66 $X2=0.59 $Y2=1.485
cc_59 VPB N_VPWR_c_287_n 0.00891827f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_60 N_A_84_48#_M1009_g N_A1_M1008_g 0.0209698f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_61 N_A_84_48#_c_61_n N_A1_M1008_g 0.00145529f $X=0.515 $Y=1.765 $X2=0 $Y2=0
cc_62 N_A_84_48#_c_65_n N_A1_M1008_g 6.58026e-19 $X=0.71 $Y=1.485 $X2=0 $Y2=0
cc_63 N_A_84_48#_c_61_n N_A1_c_135_n 0.0385042f $X=0.515 $Y=1.765 $X2=0 $Y2=0
cc_64 N_A_84_48#_c_62_n N_A1_c_135_n 0.0036717f $X=0.71 $Y=1.95 $X2=0 $Y2=0
cc_65 N_A_84_48#_c_77_p N_A1_c_135_n 0.0166347f $X=2.195 $Y=2.035 $X2=0 $Y2=0
cc_66 N_A_84_48#_c_65_n N_A1_c_135_n 0.00170526f $X=0.71 $Y=1.485 $X2=0 $Y2=0
cc_67 N_A_84_48#_c_61_n N_A1_c_136_n 3.43766e-19 $X=0.515 $Y=1.765 $X2=0 $Y2=0
cc_68 N_A_84_48#_c_62_n N_A1_c_136_n 0.0102298f $X=0.71 $Y=1.95 $X2=0 $Y2=0
cc_69 N_A_84_48#_c_77_p N_A1_c_136_n 0.0235257f $X=2.195 $Y=2.035 $X2=0 $Y2=0
cc_70 N_A_84_48#_c_65_n N_A1_c_136_n 0.0240984f $X=0.71 $Y=1.485 $X2=0 $Y2=0
cc_71 N_A_84_48#_c_77_p N_A2_c_168_n 0.015854f $X=2.195 $Y=2.035 $X2=0 $Y2=0
cc_72 N_A_84_48#_c_69_n N_A2_c_168_n 0.00351095f $X=2.36 $Y=2.375 $X2=0 $Y2=0
cc_73 N_A_84_48#_c_77_p N_A2_c_169_n 0.0217893f $X=2.195 $Y=2.035 $X2=0 $Y2=0
cc_74 N_A_84_48#_c_77_p N_A3_c_197_n 0.0122632f $X=2.195 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_75 N_A_84_48#_c_69_n N_A3_c_197_n 0.0151658f $X=2.36 $Y=2.375 $X2=-0.19
+ $Y2=-0.245
cc_76 N_A_84_48#_c_88_p N_A3_c_197_n 0.00122754f $X=2.36 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_77 N_A_84_48#_c_77_p N_A3_c_199_n 0.0104762f $X=2.195 $Y=2.035 $X2=0 $Y2=0
cc_78 N_A_84_48#_c_88_p N_A3_c_199_n 0.0131798f $X=2.36 $Y=2.035 $X2=0 $Y2=0
cc_79 N_A_84_48#_c_69_n N_B1_c_229_n 0.00945062f $X=2.36 $Y=2.375 $X2=-0.19
+ $Y2=-0.245
cc_80 N_A_84_48#_c_70_n N_B1_c_229_n 0.017672f $X=3.085 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_81 N_A_84_48#_c_64_n N_B1_c_229_n 0.0127548f $X=3.17 $Y=1.95 $X2=-0.19
+ $Y2=-0.245
cc_82 N_A_84_48#_c_63_n N_B1_M1004_g 0.0132958f $X=3.08 $Y=0.615 $X2=0 $Y2=0
cc_83 N_A_84_48#_c_64_n N_B1_M1004_g 0.00714331f $X=3.17 $Y=1.95 $X2=0 $Y2=0
cc_84 N_A_84_48#_c_70_n N_B1_c_231_n 0.0243966f $X=3.085 $Y=2.035 $X2=0 $Y2=0
cc_85 N_A_84_48#_c_64_n N_B1_c_231_n 0.0330212f $X=3.17 $Y=1.95 $X2=0 $Y2=0
cc_86 N_A_84_48#_M1009_g N_X_c_255_n 0.00805909f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_87 N_A_84_48#_M1009_g N_X_c_256_n 0.00272781f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_88 N_A_84_48#_c_65_n N_X_c_256_n 0.00138666f $X=0.71 $Y=1.485 $X2=0 $Y2=0
cc_89 N_A_84_48#_c_61_n X 0.0031072f $X=0.515 $Y=1.765 $X2=0 $Y2=0
cc_90 N_A_84_48#_c_62_n X 0.00567892f $X=0.71 $Y=1.95 $X2=0 $Y2=0
cc_91 N_A_84_48#_c_65_n X 0.00238236f $X=0.71 $Y=1.485 $X2=0 $Y2=0
cc_92 N_A_84_48#_c_61_n X 0.0131077f $X=0.515 $Y=1.765 $X2=0 $Y2=0
cc_93 N_A_84_48#_M1009_g N_X_c_257_n 0.0122939f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_94 N_A_84_48#_c_61_n N_X_c_257_n 0.00261936f $X=0.515 $Y=1.765 $X2=0 $Y2=0
cc_95 N_A_84_48#_c_62_n N_X_c_257_n 0.00525753f $X=0.71 $Y=1.95 $X2=0 $Y2=0
cc_96 N_A_84_48#_c_65_n N_X_c_257_n 0.0249901f $X=0.71 $Y=1.485 $X2=0 $Y2=0
cc_97 N_A_84_48#_c_62_n N_VPWR_M1002_d 0.00232437f $X=0.71 $Y=1.95 $X2=-0.19
+ $Y2=-0.245
cc_98 N_A_84_48#_c_77_p N_VPWR_M1002_d 0.0117909f $X=2.195 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_99 N_A_84_48#_c_111_p N_VPWR_M1002_d 0.00300113f $X=0.795 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_100 N_A_84_48#_c_70_n N_VPWR_M1005_d 0.0203419f $X=3.085 $Y=2.035 $X2=0 $Y2=0
cc_101 N_A_84_48#_c_64_n N_VPWR_M1005_d 0.0022761f $X=3.17 $Y=1.95 $X2=0 $Y2=0
cc_102 N_A_84_48#_c_61_n N_VPWR_c_280_n 0.0106903f $X=0.515 $Y=1.765 $X2=0 $Y2=0
cc_103 N_A_84_48#_c_77_p N_VPWR_c_280_n 0.0225812f $X=2.195 $Y=2.035 $X2=0 $Y2=0
cc_104 N_A_84_48#_c_111_p N_VPWR_c_280_n 0.0129456f $X=0.795 $Y=2.035 $X2=0
+ $Y2=0
cc_105 N_A_84_48#_c_69_n N_VPWR_c_281_n 0.0394066f $X=2.36 $Y=2.375 $X2=0 $Y2=0
cc_106 N_A_84_48#_c_70_n N_VPWR_c_281_n 0.0207131f $X=3.085 $Y=2.035 $X2=0 $Y2=0
cc_107 N_A_84_48#_c_69_n N_VPWR_c_282_n 0.0103753f $X=2.36 $Y=2.375 $X2=0 $Y2=0
cc_108 N_A_84_48#_c_61_n N_VPWR_c_284_n 0.00445602f $X=0.515 $Y=1.765 $X2=0
+ $Y2=0
cc_109 N_A_84_48#_c_61_n N_VPWR_c_279_n 0.00865246f $X=0.515 $Y=1.765 $X2=0
+ $Y2=0
cc_110 N_A_84_48#_c_69_n N_VPWR_c_279_n 0.0113454f $X=2.36 $Y=2.375 $X2=0 $Y2=0
cc_111 N_A_84_48#_c_77_p A_256_368# 0.0119045f $X=2.195 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_112 N_A_84_48#_c_77_p A_340_368# 0.0165158f $X=2.195 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_113 N_A_84_48#_M1009_g N_VGND_c_318_n 0.00946427f $X=0.495 $Y=0.74 $X2=0
+ $Y2=0
cc_114 N_A_84_48#_c_61_n N_VGND_c_318_n 0.00320573f $X=0.515 $Y=1.765 $X2=0
+ $Y2=0
cc_115 N_A_84_48#_c_65_n N_VGND_c_318_n 0.0140528f $X=0.71 $Y=1.485 $X2=0 $Y2=0
cc_116 N_A_84_48#_M1009_g N_VGND_c_322_n 0.00434272f $X=0.495 $Y=0.74 $X2=0
+ $Y2=0
cc_117 N_A_84_48#_c_63_n N_VGND_c_323_n 0.0107295f $X=3.08 $Y=0.615 $X2=0 $Y2=0
cc_118 N_A_84_48#_M1009_g N_VGND_c_324_n 0.00828717f $X=0.495 $Y=0.74 $X2=0
+ $Y2=0
cc_119 N_A_84_48#_c_63_n N_VGND_c_324_n 0.0117056f $X=3.08 $Y=0.615 $X2=0 $Y2=0
cc_120 N_A_84_48#_c_66_n N_A_230_94#_c_358_n 0.00795851f $X=3.085 $Y=1.13 $X2=0
+ $Y2=0
cc_121 N_A_84_48#_c_63_n N_A_230_94#_c_360_n 0.019893f $X=3.08 $Y=0.615 $X2=0
+ $Y2=0
cc_122 N_A1_M1008_g N_A2_M1006_g 0.022073f $X=1.075 $Y=0.79 $X2=0 $Y2=0
cc_123 N_A1_c_135_n N_A2_c_168_n 0.0840966f $X=1.205 $Y=1.765 $X2=0 $Y2=0
cc_124 N_A1_c_136_n N_A2_c_168_n 0.00209467f $X=1.13 $Y=1.515 $X2=0 $Y2=0
cc_125 N_A1_M1008_g N_A2_c_169_n 2.93475e-19 $X=1.075 $Y=0.79 $X2=0 $Y2=0
cc_126 N_A1_c_135_n N_A2_c_169_n 8.38018e-19 $X=1.205 $Y=1.765 $X2=0 $Y2=0
cc_127 N_A1_c_136_n N_A2_c_169_n 0.0320796f $X=1.13 $Y=1.515 $X2=0 $Y2=0
cc_128 N_A1_c_135_n X 8.16665e-19 $X=1.205 $Y=1.765 $X2=0 $Y2=0
cc_129 N_A1_c_135_n N_VPWR_c_280_n 0.00835009f $X=1.205 $Y=1.765 $X2=0 $Y2=0
cc_130 N_A1_c_135_n N_VPWR_c_282_n 0.0049405f $X=1.205 $Y=1.765 $X2=0 $Y2=0
cc_131 N_A1_c_135_n N_VPWR_c_279_n 0.00508379f $X=1.205 $Y=1.765 $X2=0 $Y2=0
cc_132 N_A1_M1008_g N_VGND_c_318_n 0.00744236f $X=1.075 $Y=0.79 $X2=0 $Y2=0
cc_133 N_A1_M1008_g N_VGND_c_320_n 0.00485498f $X=1.075 $Y=0.79 $X2=0 $Y2=0
cc_134 N_A1_M1008_g N_VGND_c_324_n 0.00514438f $X=1.075 $Y=0.79 $X2=0 $Y2=0
cc_135 N_A1_M1008_g N_A_230_94#_c_357_n 0.00590569f $X=1.075 $Y=0.79 $X2=0 $Y2=0
cc_136 N_A1_M1008_g N_A_230_94#_c_359_n 0.00247091f $X=1.075 $Y=0.79 $X2=0 $Y2=0
cc_137 N_A1_c_135_n N_A_230_94#_c_359_n 0.00109423f $X=1.205 $Y=1.765 $X2=0
+ $Y2=0
cc_138 N_A1_c_136_n N_A_230_94#_c_359_n 0.0133988f $X=1.13 $Y=1.515 $X2=0 $Y2=0
cc_139 N_A2_c_168_n N_A3_c_197_n 0.0649444f $X=1.625 $Y=1.765 $X2=-0.19
+ $Y2=-0.245
cc_140 N_A2_c_169_n N_A3_c_197_n 0.00194911f $X=1.67 $Y=1.465 $X2=-0.19
+ $Y2=-0.245
cc_141 N_A2_M1006_g N_A3_M1003_g 0.0169838f $X=1.58 $Y=0.79 $X2=0 $Y2=0
cc_142 N_A2_c_168_n N_A3_M1003_g 0.00168165f $X=1.625 $Y=1.765 $X2=0 $Y2=0
cc_143 N_A2_c_169_n N_A3_M1003_g 2.86174e-19 $X=1.67 $Y=1.465 $X2=0 $Y2=0
cc_144 N_A2_c_168_n N_A3_c_199_n 0.00116285f $X=1.625 $Y=1.765 $X2=0 $Y2=0
cc_145 N_A2_c_169_n N_A3_c_199_n 0.0279436f $X=1.67 $Y=1.465 $X2=0 $Y2=0
cc_146 N_A2_c_168_n N_VPWR_c_282_n 0.0049405f $X=1.625 $Y=1.765 $X2=0 $Y2=0
cc_147 N_A2_c_168_n N_VPWR_c_279_n 0.00508379f $X=1.625 $Y=1.765 $X2=0 $Y2=0
cc_148 N_A2_M1006_g N_VGND_c_319_n 0.0070805f $X=1.58 $Y=0.79 $X2=0 $Y2=0
cc_149 N_A2_M1006_g N_VGND_c_320_n 0.00507111f $X=1.58 $Y=0.79 $X2=0 $Y2=0
cc_150 N_A2_M1006_g N_VGND_c_324_n 0.00514438f $X=1.58 $Y=0.79 $X2=0 $Y2=0
cc_151 N_A2_M1006_g N_A_230_94#_c_357_n 0.00279704f $X=1.58 $Y=0.79 $X2=0 $Y2=0
cc_152 N_A2_M1006_g N_A_230_94#_c_358_n 0.0163236f $X=1.58 $Y=0.79 $X2=0 $Y2=0
cc_153 N_A2_c_168_n N_A_230_94#_c_358_n 0.001257f $X=1.625 $Y=1.765 $X2=0 $Y2=0
cc_154 N_A2_c_169_n N_A_230_94#_c_358_n 0.0249418f $X=1.67 $Y=1.465 $X2=0 $Y2=0
cc_155 N_A3_c_197_n N_B1_c_229_n 0.0379472f $X=2.135 $Y=1.765 $X2=-0.19
+ $Y2=-0.245
cc_156 N_A3_c_199_n N_B1_c_229_n 7.18891e-19 $X=2.21 $Y=1.515 $X2=-0.19
+ $Y2=-0.245
cc_157 N_A3_M1003_g N_B1_M1004_g 0.023509f $X=2.3 $Y=0.79 $X2=0 $Y2=0
cc_158 N_A3_c_197_n N_B1_c_231_n 0.00214941f $X=2.135 $Y=1.765 $X2=0 $Y2=0
cc_159 N_A3_c_199_n N_B1_c_231_n 0.0347535f $X=2.21 $Y=1.515 $X2=0 $Y2=0
cc_160 N_A3_c_197_n N_VPWR_c_281_n 0.00249115f $X=2.135 $Y=1.765 $X2=0 $Y2=0
cc_161 N_A3_c_197_n N_VPWR_c_282_n 0.00481822f $X=2.135 $Y=1.765 $X2=0 $Y2=0
cc_162 N_A3_c_197_n N_VPWR_c_279_n 0.00508379f $X=2.135 $Y=1.765 $X2=0 $Y2=0
cc_163 N_A3_M1003_g N_VGND_c_319_n 0.00716063f $X=2.3 $Y=0.79 $X2=0 $Y2=0
cc_164 N_A3_M1003_g N_VGND_c_323_n 0.00507111f $X=2.3 $Y=0.79 $X2=0 $Y2=0
cc_165 N_A3_M1003_g N_VGND_c_324_n 0.00514438f $X=2.3 $Y=0.79 $X2=0 $Y2=0
cc_166 N_A3_c_197_n N_A_230_94#_c_358_n 0.00118195f $X=2.135 $Y=1.765 $X2=0
+ $Y2=0
cc_167 N_A3_M1003_g N_A_230_94#_c_358_n 0.0165716f $X=2.3 $Y=0.79 $X2=0 $Y2=0
cc_168 N_A3_c_199_n N_A_230_94#_c_358_n 0.0202397f $X=2.21 $Y=1.515 $X2=0 $Y2=0
cc_169 N_A3_M1003_g N_A_230_94#_c_360_n 0.00275413f $X=2.3 $Y=0.79 $X2=0 $Y2=0
cc_170 N_B1_c_229_n N_VPWR_c_281_n 0.00922946f $X=2.675 $Y=1.765 $X2=0 $Y2=0
cc_171 N_B1_c_229_n N_VPWR_c_282_n 0.00361294f $X=2.675 $Y=1.765 $X2=0 $Y2=0
cc_172 N_B1_c_229_n N_VPWR_c_279_n 0.00419404f $X=2.675 $Y=1.765 $X2=0 $Y2=0
cc_173 N_B1_M1004_g N_VGND_c_323_n 0.00485498f $X=2.795 $Y=0.79 $X2=0 $Y2=0
cc_174 N_B1_M1004_g N_VGND_c_324_n 0.00514438f $X=2.795 $Y=0.79 $X2=0 $Y2=0
cc_175 N_B1_c_229_n N_A_230_94#_c_358_n 0.00101882f $X=2.675 $Y=1.765 $X2=0
+ $Y2=0
cc_176 N_B1_M1004_g N_A_230_94#_c_358_n 0.00247983f $X=2.795 $Y=0.79 $X2=0 $Y2=0
cc_177 N_B1_c_231_n N_A_230_94#_c_358_n 0.0141977f $X=2.75 $Y=1.515 $X2=0 $Y2=0
cc_178 N_B1_M1004_g N_A_230_94#_c_360_n 0.00594451f $X=2.795 $Y=0.79 $X2=0 $Y2=0
cc_179 X N_VPWR_c_280_n 0.0271803f $X=0.24 $Y=2.035 $X2=0 $Y2=0
cc_180 X N_VPWR_c_284_n 0.0163786f $X=0.24 $Y=2.035 $X2=0 $Y2=0
cc_181 X N_VPWR_c_279_n 0.0135239f $X=0.24 $Y=2.035 $X2=0 $Y2=0
cc_182 N_X_c_255_n N_VGND_c_318_n 0.0312028f $X=0.28 $Y=0.515 $X2=0 $Y2=0
cc_183 N_X_c_255_n N_VGND_c_322_n 0.0159025f $X=0.28 $Y=0.515 $X2=0 $Y2=0
cc_184 N_X_c_255_n N_VGND_c_324_n 0.0131064f $X=0.28 $Y=0.515 $X2=0 $Y2=0
cc_185 N_VGND_c_318_n N_A_230_94#_c_357_n 0.0190445f $X=0.78 $Y=0.515 $X2=0
+ $Y2=0
cc_186 N_VGND_c_319_n N_A_230_94#_c_357_n 0.00929705f $X=1.945 $Y=0.615 $X2=0
+ $Y2=0
cc_187 N_VGND_c_320_n N_A_230_94#_c_357_n 0.0105078f $X=1.765 $Y=0 $X2=0 $Y2=0
cc_188 N_VGND_c_324_n N_A_230_94#_c_357_n 0.0115086f $X=3.12 $Y=0 $X2=0 $Y2=0
cc_189 N_VGND_M1006_d N_A_230_94#_c_358_n 0.00923283f $X=1.655 $Y=0.47 $X2=0
+ $Y2=0
cc_190 N_VGND_c_319_n N_A_230_94#_c_358_n 0.0282971f $X=1.945 $Y=0.615 $X2=0
+ $Y2=0
cc_191 N_VGND_c_318_n N_A_230_94#_c_359_n 0.00760062f $X=0.78 $Y=0.515 $X2=0
+ $Y2=0
cc_192 N_VGND_c_319_n N_A_230_94#_c_360_n 0.00976671f $X=1.945 $Y=0.615 $X2=0
+ $Y2=0
cc_193 N_VGND_c_323_n N_A_230_94#_c_360_n 0.0103491f $X=3.12 $Y=0 $X2=0 $Y2=0
cc_194 N_VGND_c_324_n N_A_230_94#_c_360_n 0.0113354f $X=3.12 $Y=0 $X2=0 $Y2=0
