* File: sky130_fd_sc_hs__a221oi_2.pex.spice
* Created: Tue Sep  1 19:50:31 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HS__A221OI_2%C1 1 3 6 8 10 13 15 21 22
r46 22 23 1.9127 $w=3.78e-07 $l=1.5e-08 $layer=POLY_cond $X=0.945 $Y=1.557
+ $X2=0.96 $Y2=1.557
r47 20 22 24.8651 $w=3.78e-07 $l=1.95e-07 $layer=POLY_cond $X=0.75 $Y=1.557
+ $X2=0.945 $Y2=1.557
r48 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.75
+ $Y=1.515 $X2=0.75 $Y2=1.515
r49 18 20 30.6032 $w=3.78e-07 $l=2.4e-07 $layer=POLY_cond $X=0.51 $Y=1.557
+ $X2=0.75 $Y2=1.557
r50 17 18 1.9127 $w=3.78e-07 $l=1.5e-08 $layer=POLY_cond $X=0.495 $Y=1.557
+ $X2=0.51 $Y2=1.557
r51 15 21 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=0.75 $Y=1.665
+ $X2=0.75 $Y2=1.515
r52 11 23 24.4846 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.96 $Y=1.35
+ $X2=0.96 $Y2=1.557
r53 11 13 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=0.96 $Y=1.35
+ $X2=0.96 $Y2=0.74
r54 8 22 24.4846 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=0.945 $Y=1.765
+ $X2=0.945 $Y2=1.557
r55 8 10 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.945 $Y=1.765
+ $X2=0.945 $Y2=2.4
r56 4 18 24.4846 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.51 $Y=1.35
+ $X2=0.51 $Y2=1.557
r57 4 6 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=0.51 $Y=1.35 $X2=0.51
+ $Y2=0.74
r58 1 17 24.4846 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=0.495 $Y=1.765
+ $X2=0.495 $Y2=1.557
r59 1 3 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.495 $Y=1.765
+ $X2=0.495 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_HS__A221OI_2%B1 3 5 7 8 10 13 16 17 18 23 25
c95 13 0 1.99054e-19 $X=2.83 $Y=0.74
c96 5 0 1.53182e-20 $X=1.395 $Y=1.765
r97 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.85
+ $Y=1.515 $X2=2.85 $Y2=1.515
r98 25 37 7.02022 $w=6.43e-07 $l=3.7e-07 $layer=LI1_cond $X=2.88 $Y=1.665
+ $X2=2.88 $Y2=2.035
r99 25 32 2.84603 $w=6.43e-07 $l=1.5e-07 $layer=LI1_cond $X=2.88 $Y=1.665
+ $X2=2.88 $Y2=1.515
r100 20 23 4.60977 $w=2.48e-07 $l=1e-07 $layer=LI1_cond $X=1.41 $Y=1.555
+ $X2=1.51 $Y2=1.555
r101 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.41
+ $Y=1.515 $X2=1.41 $Y2=1.515
r102 17 37 8.76525 $w=1.7e-07 $l=3.55e-07 $layer=LI1_cond $X=2.525 $Y=2.035
+ $X2=2.88 $Y2=2.035
r103 17 18 60.6738 $w=1.68e-07 $l=9.3e-07 $layer=LI1_cond $X=2.525 $Y=2.035
+ $X2=1.595 $Y2=2.035
r104 16 18 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.51 $Y=1.95
+ $X2=1.595 $Y2=2.035
r105 15 23 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.51 $Y=1.68
+ $X2=1.51 $Y2=1.555
r106 15 16 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=1.51 $Y=1.68
+ $X2=1.51 $Y2=1.95
r107 11 31 38.5562 $w=2.99e-07 $l=1.74714e-07 $layer=POLY_cond $X=2.83 $Y=1.35
+ $X2=2.85 $Y2=1.515
r108 11 13 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.83 $Y=1.35
+ $X2=2.83 $Y2=0.74
r109 8 31 52.2586 $w=2.99e-07 $l=2.85044e-07 $layer=POLY_cond $X=2.775 $Y=1.765
+ $X2=2.85 $Y2=1.515
r110 8 10 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.775 $Y=1.765
+ $X2=2.775 $Y2=2.4
r111 5 21 52.2586 $w=2.99e-07 $l=2.57391e-07 $layer=POLY_cond $X=1.395 $Y=1.765
+ $X2=1.41 $Y2=1.515
r112 5 7 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.395 $Y=1.765
+ $X2=1.395 $Y2=2.4
r113 1 21 38.5562 $w=2.99e-07 $l=1.74714e-07 $layer=POLY_cond $X=1.39 $Y=1.35
+ $X2=1.41 $Y2=1.515
r114 1 3 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.39 $Y=1.35 $X2=1.39
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HS__A221OI_2%B2 3 5 7 8 10 13 15 21 22
c52 3 0 1.69771e-19 $X=1.86 $Y=0.74
r53 22 23 10.0978 $w=3.58e-07 $l=7.5e-08 $layer=POLY_cond $X=2.325 $Y=1.557
+ $X2=2.4 $Y2=1.557
r54 20 22 28.9469 $w=3.58e-07 $l=2.15e-07 $layer=POLY_cond $X=2.11 $Y=1.557
+ $X2=2.325 $Y2=1.557
r55 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.11
+ $Y=1.515 $X2=2.11 $Y2=1.515
r56 18 20 31.6397 $w=3.58e-07 $l=2.35e-07 $layer=POLY_cond $X=1.875 $Y=1.557
+ $X2=2.11 $Y2=1.557
r57 17 18 2.01955 $w=3.58e-07 $l=1.5e-08 $layer=POLY_cond $X=1.86 $Y=1.557
+ $X2=1.875 $Y2=1.557
r58 15 21 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=2.11 $Y=1.665
+ $X2=2.11 $Y2=1.515
r59 11 23 23.1716 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.4 $Y=1.35 $X2=2.4
+ $Y2=1.557
r60 11 13 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.4 $Y=1.35 $X2=2.4
+ $Y2=0.74
r61 8 22 23.1716 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=2.325 $Y=1.765
+ $X2=2.325 $Y2=1.557
r62 8 10 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.325 $Y=1.765
+ $X2=2.325 $Y2=2.4
r63 5 18 23.1716 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=1.875 $Y=1.765
+ $X2=1.875 $Y2=1.557
r64 5 7 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.875 $Y=1.765
+ $X2=1.875 $Y2=2.4
r65 1 17 23.1716 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.86 $Y=1.35
+ $X2=1.86 $Y2=1.557
r66 1 3 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.86 $Y=1.35 $X2=1.86
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HS__A221OI_2%A1 3 5 7 10 12 14 17 18 20 21 22 23 24 25
c78 22 0 1.26728e-19 $X=4.98 $Y=1.78
c79 5 0 1.07574e-19 $X=3.745 $Y=1.765
c80 3 0 1.63824e-19 $X=3.3 $Y=0.74
r81 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.14
+ $Y=1.515 $X2=5.14 $Y2=1.515
r82 25 34 12.5122 $w=3.48e-07 $l=3.8e-07 $layer=LI1_cond $X=5.52 $Y=1.605
+ $X2=5.14 $Y2=1.605
r83 24 35 2.59474 $w=3.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.98 $Y=1.605
+ $X2=5.065 $Y2=1.605
r84 24 34 1.48171 $w=3.48e-07 $l=4.5e-08 $layer=LI1_cond $X=5.095 $Y=1.605
+ $X2=5.14 $Y2=1.605
r85 24 35 0.987808 $w=3.48e-07 $l=3e-08 $layer=LI1_cond $X=5.095 $Y=1.605
+ $X2=5.065 $Y2=1.605
r86 22 24 5.34211 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=4.98 $Y=1.78
+ $X2=4.98 $Y2=1.605
r87 22 23 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=4.98 $Y=1.78
+ $X2=4.98 $Y2=1.95
r88 20 23 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.895 $Y=2.035
+ $X2=4.98 $Y2=1.95
r89 20 21 75.6791 $w=1.68e-07 $l=1.16e-06 $layer=LI1_cond $X=4.895 $Y=2.035
+ $X2=3.735 $Y2=2.035
r90 18 31 23.7606 $w=3.55e-07 $l=1.75e-07 $layer=POLY_cond $X=3.57 $Y=1.557
+ $X2=3.745 $Y2=1.557
r91 18 29 36.6592 $w=3.55e-07 $l=2.7e-07 $layer=POLY_cond $X=3.57 $Y=1.557
+ $X2=3.3 $Y2=1.557
r92 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.57
+ $Y=1.515 $X2=3.57 $Y2=1.515
r93 15 21 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.57 $Y=1.95
+ $X2=3.735 $Y2=2.035
r94 15 17 15.1913 $w=3.28e-07 $l=4.35e-07 $layer=LI1_cond $X=3.57 $Y=1.95
+ $X2=3.57 $Y2=1.515
r95 12 33 52.2586 $w=2.99e-07 $l=2.7157e-07 $layer=POLY_cond $X=5.095 $Y=1.765
+ $X2=5.14 $Y2=1.515
r96 12 14 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=5.095 $Y=1.765
+ $X2=5.095 $Y2=2.4
r97 8 33 38.5562 $w=2.99e-07 $l=2.05122e-07 $layer=POLY_cond $X=5.05 $Y=1.35
+ $X2=5.14 $Y2=1.515
r98 8 10 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=5.05 $Y=1.35 $X2=5.05
+ $Y2=0.74
r99 5 31 22.9692 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=3.745 $Y=1.765
+ $X2=3.745 $Y2=1.557
r100 5 7 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.745 $Y=1.765
+ $X2=3.745 $Y2=2.4
r101 1 29 22.9692 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.3 $Y=1.35 $X2=3.3
+ $Y2=1.557
r102 1 3 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=3.3 $Y=1.35 $X2=3.3
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HS__A221OI_2%A2 3 5 7 10 12 14 15 16 24
c52 16 0 1.07574e-19 $X=4.56 $Y=1.665
c53 12 0 1.26728e-19 $X=4.645 $Y=1.765
r54 24 25 3.22193 $w=3.74e-07 $l=2.5e-08 $layer=POLY_cond $X=4.62 $Y=1.557
+ $X2=4.645 $Y2=1.557
r55 22 24 52.8396 $w=3.74e-07 $l=4.1e-07 $layer=POLY_cond $X=4.21 $Y=1.557
+ $X2=4.62 $Y2=1.557
r56 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.21
+ $Y=1.515 $X2=4.21 $Y2=1.515
r57 20 22 1.93316 $w=3.74e-07 $l=1.5e-08 $layer=POLY_cond $X=4.195 $Y=1.557
+ $X2=4.21 $Y2=1.557
r58 19 20 9.66578 $w=3.74e-07 $l=7.5e-08 $layer=POLY_cond $X=4.12 $Y=1.557
+ $X2=4.195 $Y2=1.557
r59 16 23 11.5244 $w=3.48e-07 $l=3.5e-07 $layer=LI1_cond $X=4.56 $Y=1.605
+ $X2=4.21 $Y2=1.605
r60 15 23 4.2805 $w=3.48e-07 $l=1.3e-07 $layer=LI1_cond $X=4.08 $Y=1.605
+ $X2=4.21 $Y2=1.605
r61 12 25 24.2268 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=4.645 $Y=1.765
+ $X2=4.645 $Y2=1.557
r62 12 14 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=4.645 $Y=1.765
+ $X2=4.645 $Y2=2.4
r63 8 24 24.2268 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.62 $Y=1.35
+ $X2=4.62 $Y2=1.557
r64 8 10 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=4.62 $Y=1.35 $X2=4.62
+ $Y2=0.74
r65 5 20 24.2268 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=4.195 $Y=1.765
+ $X2=4.195 $Y2=1.557
r66 5 7 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=4.195 $Y=1.765
+ $X2=4.195 $Y2=2.4
r67 1 19 24.2268 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.12 $Y=1.35
+ $X2=4.12 $Y2=1.557
r68 1 3 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=4.12 $Y=1.35 $X2=4.12
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HS__A221OI_2%A_29_368# 1 2 3 4 15 17 18 21 29 31 34 35
r50 33 35 4.83021 $w=4.43e-07 $l=1.65e-07 $layer=LI1_cond $X=2.1 $Y=2.852
+ $X2=2.265 $Y2=2.852
r51 33 34 6.78944 $w=4.43e-07 $l=8.5e-08 $layer=LI1_cond $X=2.1 $Y=2.852
+ $X2=2.015 $Y2=2.852
r52 29 35 24.2013 $w=3.48e-07 $l=7.35e-07 $layer=LI1_cond $X=3 $Y=2.805
+ $X2=2.265 $Y2=2.805
r53 26 31 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.255 $Y=2.99
+ $X2=1.17 $Y2=2.99
r54 26 34 49.5829 $w=1.68e-07 $l=7.6e-07 $layer=LI1_cond $X=1.255 $Y=2.99
+ $X2=2.015 $Y2=2.99
r55 21 24 52.1925 $w=1.68e-07 $l=8e-07 $layer=LI1_cond $X=1.17 $Y=2.015 $X2=1.17
+ $Y2=2.815
r56 19 31 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.17 $Y=2.905
+ $X2=1.17 $Y2=2.99
r57 19 24 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=1.17 $Y=2.905 $X2=1.17
+ $Y2=2.815
r58 17 31 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.085 $Y=2.99
+ $X2=1.17 $Y2=2.99
r59 17 18 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=1.085 $Y=2.99
+ $X2=0.355 $Y2=2.99
r60 13 18 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.23 $Y=2.905
+ $X2=0.355 $Y2=2.99
r61 13 15 20.744 $w=2.48e-07 $l=4.5e-07 $layer=LI1_cond $X=0.23 $Y=2.905
+ $X2=0.23 $Y2=2.455
r62 4 29 600 $w=1.7e-07 $l=1.03729e-06 $layer=licon1_PDIFF $count=1 $X=2.85
+ $Y=1.84 $X2=3 $Y2=2.805
r63 3 33 600 $w=1.7e-07 $l=1.03729e-06 $layer=licon1_PDIFF $count=1 $X=1.95
+ $Y=1.84 $X2=2.1 $Y2=2.805
r64 2 24 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=1.02
+ $Y=1.84 $X2=1.17 $Y2=2.815
r65 2 21 400 $w=1.7e-07 $l=2.38485e-07 $layer=licon1_PDIFF $count=1 $X=1.02
+ $Y=1.84 $X2=1.17 $Y2=2.015
r66 1 15 300 $w=1.7e-07 $l=6.74611e-07 $layer=licon1_PDIFF $count=2 $X=0.145
+ $Y=1.84 $X2=0.27 $Y2=2.455
.ends

.subckt PM_SKY130_FD_SC_HS__A221OI_2%Y 1 2 3 4 5 18 20 22 23 28 30 34 36 40 43
+ 46 47 48 49 50
r93 49 50 16.7217 $w=2.53e-07 $l=3.7e-07 $layer=LI1_cond $X=0.252 $Y=1.295
+ $X2=0.252 $Y2=1.665
r94 44 50 12.8802 $w=2.53e-07 $l=2.85e-07 $layer=LI1_cond $X=0.252 $Y=1.95
+ $X2=0.252 $Y2=1.665
r95 42 49 5.19729 $w=2.53e-07 $l=1.15e-07 $layer=LI1_cond $X=0.252 $Y=1.18
+ $X2=0.252 $Y2=1.295
r96 42 43 3.64284 $w=2.55e-07 $l=8.5e-08 $layer=LI1_cond $X=0.252 $Y=1.18
+ $X2=0.252 $Y2=1.095
r97 38 40 26.5062 $w=2.48e-07 $l=5.75e-07 $layer=LI1_cond $X=5.305 $Y=1.09
+ $X2=5.305 $Y2=0.515
r98 37 48 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=3.18 $Y=1.175
+ $X2=3.065 $Y2=1.175
r99 36 38 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=5.18 $Y=1.175
+ $X2=5.305 $Y2=1.09
r100 36 37 130.481 $w=1.68e-07 $l=2e-06 $layer=LI1_cond $X=5.18 $Y=1.175
+ $X2=3.18 $Y2=1.175
r101 32 48 0.280307 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.065 $Y=1.09
+ $X2=3.065 $Y2=1.175
r102 32 34 28.8111 $w=2.28e-07 $l=5.75e-07 $layer=LI1_cond $X=3.065 $Y=1.09
+ $X2=3.065 $Y2=0.515
r103 31 47 5.16603 $w=1.7e-07 $l=1.03078e-07 $layer=LI1_cond $X=1.26 $Y=1.175
+ $X2=1.175 $Y2=1.135
r104 30 48 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=2.95 $Y=1.175
+ $X2=3.065 $Y2=1.175
r105 30 31 110.257 $w=1.68e-07 $l=1.69e-06 $layer=LI1_cond $X=2.95 $Y=1.175
+ $X2=1.26 $Y2=1.175
r106 26 47 1.34256 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.175 $Y=1.01
+ $X2=1.175 $Y2=1.135
r107 26 28 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=1.175 $Y=1.01
+ $X2=1.175 $Y2=0.515
r108 23 44 7.17723 $w=1.7e-07 $l=1.65118e-07 $layer=LI1_cond $X=0.38 $Y=2.035
+ $X2=0.252 $Y2=1.95
r109 22 46 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.555 $Y=2.035
+ $X2=0.72 $Y2=2.035
r110 22 23 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=0.555 $Y=2.035
+ $X2=0.38 $Y2=2.035
r111 21 43 2.83584 $w=1.7e-07 $l=1.28e-07 $layer=LI1_cond $X=0.38 $Y=1.095
+ $X2=0.252 $Y2=1.095
r112 20 47 5.16603 $w=1.7e-07 $l=1.03078e-07 $layer=LI1_cond $X=1.09 $Y=1.095
+ $X2=1.175 $Y2=1.135
r113 20 21 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=1.09 $Y=1.095
+ $X2=0.38 $Y2=1.095
r114 16 43 3.64284 $w=2.55e-07 $l=8.5e-08 $layer=LI1_cond $X=0.252 $Y=1.01
+ $X2=0.252 $Y2=1.095
r115 16 18 22.371 $w=2.53e-07 $l=4.95e-07 $layer=LI1_cond $X=0.252 $Y=1.01
+ $X2=0.252 $Y2=0.515
r116 5 46 300 $w=1.7e-07 $l=2.85307e-07 $layer=licon1_PDIFF $count=2 $X=0.57
+ $Y=1.84 $X2=0.72 $Y2=2.06
r117 4 40 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=5.125
+ $Y=0.37 $X2=5.265 $Y2=0.515
r118 3 34 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.905
+ $Y=0.37 $X2=3.045 $Y2=0.515
r119 2 28 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.035
+ $Y=0.37 $X2=1.175 $Y2=0.515
r120 1 18 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.17
+ $Y=0.37 $X2=0.295 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__A221OI_2%A_294_368# 1 2 3 4 13 19 23 29 31
c57 13 0 1.53182e-20 $X=3.805 $Y=2.375
r58 23 26 4.32166 $w=3.58e-07 $l=1.35e-07 $layer=LI1_cond $X=1.635 $Y=2.375
+ $X2=1.635 $Y2=2.51
r59 20 29 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.135 $Y=2.375
+ $X2=3.97 $Y2=2.375
r60 19 31 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.705 $Y=2.375
+ $X2=4.87 $Y2=2.375
r61 19 20 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=4.705 $Y=2.375
+ $X2=4.135 $Y2=2.375
r62 14 23 5.14255 $w=1.7e-07 $l=1.8e-07 $layer=LI1_cond $X=1.815 $Y=2.375
+ $X2=1.635 $Y2=2.375
r63 14 16 47.9519 $w=1.68e-07 $l=7.35e-07 $layer=LI1_cond $X=1.815 $Y=2.375
+ $X2=2.55 $Y2=2.375
r64 13 29 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.805 $Y=2.375
+ $X2=3.97 $Y2=2.375
r65 13 16 81.877 $w=1.68e-07 $l=1.255e-06 $layer=LI1_cond $X=3.805 $Y=2.375
+ $X2=2.55 $Y2=2.375
r66 4 31 300 $w=1.7e-07 $l=6.20484e-07 $layer=licon1_PDIFF $count=2 $X=4.72
+ $Y=1.84 $X2=4.87 $Y2=2.39
r67 3 29 300 $w=1.7e-07 $l=6.20484e-07 $layer=licon1_PDIFF $count=2 $X=3.82
+ $Y=1.84 $X2=3.97 $Y2=2.39
r68 2 16 600 $w=1.7e-07 $l=6.05372e-07 $layer=licon1_PDIFF $count=1 $X=2.4
+ $Y=1.84 $X2=2.55 $Y2=2.375
r69 1 26 600 $w=1.7e-07 $l=7.47964e-07 $layer=licon1_PDIFF $count=1 $X=1.47
+ $Y=1.84 $X2=1.635 $Y2=2.51
.ends

.subckt PM_SKY130_FD_SC_HS__A221OI_2%VPWR 1 2 3 12 16 20 25 26 28 29 30 31 32 33
+ 50
r65 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r66 47 50 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=5.52 $Y2=3.33
r67 46 47 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r68 44 47 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=5.04 $Y2=3.33
r69 43 44 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r70 41 44 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=4.08 $Y2=3.33
r71 40 41 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r72 36 40 187.893 $w=1.68e-07 $l=2.88e-06 $layer=LI1_cond $X=0.24 $Y=3.33
+ $X2=3.12 $Y2=3.33
r73 36 37 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r74 33 41 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.88 $Y=3.33
+ $X2=3.12 $Y2=3.33
r75 33 37 0.73586 $w=4.9e-07 $l=2.64e-06 $layer=MET1_cond $X=2.88 $Y=3.33
+ $X2=0.24 $Y2=3.33
r76 31 46 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=5.235 $Y=3.33
+ $X2=5.04 $Y2=3.33
r77 31 32 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.235 $Y=3.33
+ $X2=5.36 $Y2=3.33
r78 30 49 2.51176 $w=1.7e-07 $l=3.5e-08 $layer=LI1_cond $X=5.485 $Y=3.33
+ $X2=5.52 $Y2=3.33
r79 30 32 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.485 $Y=3.33
+ $X2=5.36 $Y2=3.33
r80 28 43 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=4.335 $Y=3.33
+ $X2=4.08 $Y2=3.33
r81 28 29 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.335 $Y=3.33
+ $X2=4.42 $Y2=3.33
r82 27 46 34.9037 $w=1.68e-07 $l=5.35e-07 $layer=LI1_cond $X=4.505 $Y=3.33
+ $X2=5.04 $Y2=3.33
r83 27 29 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.505 $Y=3.33
+ $X2=4.42 $Y2=3.33
r84 25 40 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=3.355 $Y=3.33
+ $X2=3.12 $Y2=3.33
r85 25 26 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.355 $Y=3.33
+ $X2=3.48 $Y2=3.33
r86 24 43 30.9893 $w=1.68e-07 $l=4.75e-07 $layer=LI1_cond $X=3.605 $Y=3.33
+ $X2=4.08 $Y2=3.33
r87 24 26 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.605 $Y=3.33
+ $X2=3.48 $Y2=3.33
r88 20 23 32.2684 $w=2.48e-07 $l=7e-07 $layer=LI1_cond $X=5.36 $Y=2.115 $X2=5.36
+ $Y2=2.815
r89 18 32 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.36 $Y=3.245
+ $X2=5.36 $Y2=3.33
r90 18 23 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=5.36 $Y=3.245
+ $X2=5.36 $Y2=2.815
r91 14 29 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.42 $Y=3.245
+ $X2=4.42 $Y2=3.33
r92 14 16 28.7059 $w=1.68e-07 $l=4.4e-07 $layer=LI1_cond $X=4.42 $Y=3.245
+ $X2=4.42 $Y2=2.805
r93 10 26 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.48 $Y=3.245
+ $X2=3.48 $Y2=3.33
r94 10 12 20.283 $w=2.48e-07 $l=4.4e-07 $layer=LI1_cond $X=3.48 $Y=3.245
+ $X2=3.48 $Y2=2.805
r95 3 23 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=5.17
+ $Y=1.84 $X2=5.32 $Y2=2.815
r96 3 20 400 $w=1.7e-07 $l=3.4187e-07 $layer=licon1_PDIFF $count=1 $X=5.17
+ $Y=1.84 $X2=5.32 $Y2=2.115
r97 2 16 600 $w=1.7e-07 $l=1.03729e-06 $layer=licon1_PDIFF $count=1 $X=4.27
+ $Y=1.84 $X2=4.42 $Y2=2.805
r98 1 12 600 $w=1.7e-07 $l=1.0256e-06 $layer=licon1_PDIFF $count=1 $X=3.395
+ $Y=1.84 $X2=3.52 $Y2=2.805
.ends

.subckt PM_SKY130_FD_SC_HS__A221OI_2%VGND 1 2 3 12 16 20 23 24 25 27 32 48 49 52
+ 55
r74 55 56 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r75 52 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r76 48 49 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r77 46 49 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=5.52
+ $Y2=0
r78 45 48 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=4.56 $Y=0 $X2=5.52
+ $Y2=0
r79 45 46 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r80 43 46 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=4.56
+ $Y2=0
r81 42 43 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r82 40 56 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=2.16
+ $Y2=0
r83 39 42 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=2.64 $Y=0 $X2=4.08
+ $Y2=0
r84 39 40 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r85 37 55 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=2.28 $Y=0 $X2=2.11
+ $Y2=0
r86 37 39 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=2.28 $Y=0 $X2=2.64
+ $Y2=0
r87 36 56 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r88 36 53 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=0.72
+ $Y2=0
r89 35 36 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r90 33 52 8.9695 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=0.91 $Y=0 $X2=0.735
+ $Y2=0
r91 33 35 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=0.91 $Y=0 $X2=1.68
+ $Y2=0
r92 32 55 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=1.94 $Y=0 $X2=2.11
+ $Y2=0
r93 32 35 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=1.94 $Y=0 $X2=1.68
+ $Y2=0
r94 30 53 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r95 29 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r96 27 52 8.9695 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=0.56 $Y=0 $X2=0.735
+ $Y2=0
r97 27 29 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=0.56 $Y=0 $X2=0.24
+ $Y2=0
r98 25 43 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=2.88 $Y=0 $X2=4.08
+ $Y2=0
r99 25 40 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.88 $Y=0 $X2=2.64
+ $Y2=0
r100 23 42 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=4.2 $Y=0 $X2=4.08
+ $Y2=0
r101 23 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.2 $Y=0 $X2=4.365
+ $Y2=0
r102 22 45 1.95722 $w=1.68e-07 $l=3e-08 $layer=LI1_cond $X=4.53 $Y=0 $X2=4.56
+ $Y2=0
r103 22 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.53 $Y=0 $X2=4.365
+ $Y2=0
r104 18 24 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.365 $Y=0.085
+ $X2=4.365 $Y2=0
r105 18 20 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=4.365 $Y=0.085
+ $X2=4.365 $Y2=0.495
r106 14 55 0.987631 $w=3.4e-07 $l=8.5e-08 $layer=LI1_cond $X=2.11 $Y=0.085
+ $X2=2.11 $Y2=0
r107 14 16 13.8971 $w=3.38e-07 $l=4.1e-07 $layer=LI1_cond $X=2.11 $Y=0.085
+ $X2=2.11 $Y2=0.495
r108 10 52 1.07557 $w=3.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.735 $Y=0.085
+ $X2=0.735 $Y2=0
r109 10 12 19.4269 $w=3.48e-07 $l=5.9e-07 $layer=LI1_cond $X=0.735 $Y=0.085
+ $X2=0.735 $Y2=0.675
r110 3 20 182 $w=1.7e-07 $l=2.23942e-07 $layer=licon1_NDIFF $count=1 $X=4.195
+ $Y=0.37 $X2=4.365 $Y2=0.495
r111 2 16 182 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_NDIFF $count=1 $X=1.935
+ $Y=0.37 $X2=2.11 $Y2=0.495
r112 1 12 182 $w=1.7e-07 $l=3.72525e-07 $layer=licon1_NDIFF $count=1 $X=0.585
+ $Y=0.37 $X2=0.735 $Y2=0.675
.ends

.subckt PM_SKY130_FD_SC_HS__A221OI_2%A_293_74# 1 2 7 9 11 15
c28 15 0 1.63824e-19 $X=2.615 $Y=0.495
c29 9 0 1.69771e-19 $X=1.605 $Y=0.495
r30 13 15 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=2.615 $Y=0.75
+ $X2=2.615 $Y2=0.495
r31 12 18 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.77 $Y=0.835
+ $X2=1.605 $Y2=0.835
r32 11 13 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.45 $Y=0.835
+ $X2=2.615 $Y2=0.75
r33 11 12 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=2.45 $Y=0.835
+ $X2=1.77 $Y2=0.835
r34 7 18 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.605 $Y=0.75 $X2=1.605
+ $Y2=0.835
r35 7 9 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=1.605 $Y=0.75
+ $X2=1.605 $Y2=0.495
r36 2 15 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=2.475
+ $Y=0.37 $X2=2.615 $Y2=0.495
r37 1 18 182 $w=1.7e-07 $l=5.30401e-07 $layer=licon1_NDIFF $count=1 $X=1.465
+ $Y=0.37 $X2=1.605 $Y2=0.835
r38 1 9 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=1.465
+ $Y=0.37 $X2=1.605 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_HS__A221OI_2%A_675_74# 1 2 7 9 11 16
c27 16 0 1.99054e-19 $X=4.03 $Y=0.625
r28 14 16 9.28002 $w=5.88e-07 $l=1.25e-07 $layer=LI1_cond $X=3.905 $Y=0.625
+ $X2=4.03 $Y2=0.625
r29 9 18 2.71916 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.85 $Y=0.75 $X2=4.85
+ $Y2=0.835
r30 9 11 9.79577 $w=2.98e-07 $l=2.55e-07 $layer=LI1_cond $X=4.85 $Y=0.75
+ $X2=4.85 $Y2=0.495
r31 7 18 4.79851 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=4.7 $Y=0.835 $X2=4.85
+ $Y2=0.835
r32 7 16 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.7 $Y=0.835 $X2=4.03
+ $Y2=0.835
r33 2 18 182 $w=1.7e-07 $l=5.30401e-07 $layer=licon1_NDIFF $count=1 $X=4.695
+ $Y=0.37 $X2=4.835 $Y2=0.835
r34 2 11 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=4.695
+ $Y=0.37 $X2=4.835 $Y2=0.495
r35 1 14 45.5 $w=1.7e-07 $l=5.89194e-07 $layer=licon1_NDIFF $count=4 $X=3.375
+ $Y=0.37 $X2=3.905 $Y2=0.495
.ends

