* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hs__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
X0 a_1468_493# a_1518_203# VPWR VPB sky130_fd_pr__pfet_01v8 w=420000u l=150000u
X1 VGND a_1266_74# a_1864_409# VNB sky130_fd_pr__nfet_01v8_lvt w=550000u l=150000u
X2 VGND a_306_74# a_490_366# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X3 a_30_78# a_306_74# a_695_457# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X4 a_830_359# a_490_366# a_1266_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X5 VGND a_695_457# a_830_359# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X6 VPWR a_1266_74# a_1864_409# VPB sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X7 a_306_74# CLK VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X8 a_695_457# a_306_74# a_785_457# VPB sky130_fd_pr__pfet_01v8 w=420000u l=150000u
X9 VPWR RESET_B a_695_457# VPB sky130_fd_pr__pfet_01v8 w=420000u l=150000u
X10 Q a_1864_409# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X11 VPWR D a_30_78# VPB sky130_fd_pr__pfet_01v8 w=420000u l=150000u
X12 a_306_74# CLK VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X13 a_1266_74# a_490_366# a_1468_493# VPB sky130_fd_pr__pfet_01v8 w=420000u l=150000u
X14 a_695_457# a_490_366# a_816_138# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X15 Q a_1864_409# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X16 VGND RESET_B a_1656_81# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X17 a_785_457# a_830_359# VPWR VPB sky130_fd_pr__pfet_01v8 w=420000u l=150000u
X18 a_1518_203# a_1266_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=420000u l=150000u
X19 a_1656_81# a_1266_74# a_1518_203# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X20 a_894_138# RESET_B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X21 VPWR a_695_457# a_830_359# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=150000u
X22 a_30_78# a_490_366# a_695_457# VPB sky130_fd_pr__pfet_01v8 w=420000u l=150000u
X23 VPWR a_306_74# a_490_366# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X24 a_117_78# RESET_B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X25 a_30_78# D a_117_78# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X26 a_830_359# a_306_74# a_1266_74# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=150000u
X27 a_1476_81# a_1518_203# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X28 a_816_138# a_830_359# a_894_138# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X29 a_30_78# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8 w=420000u l=150000u
X30 VPWR RESET_B a_1518_203# VPB sky130_fd_pr__pfet_01v8 w=420000u l=150000u
X31 a_1266_74# a_306_74# a_1476_81# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
.ends
