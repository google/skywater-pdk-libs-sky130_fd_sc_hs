* NGSPICE file created from sky130_fd_sc_hs__dlxtn_2.ext - technology: sky130A

.subckt sky130_fd_sc_hs__dlxtn_2 D GATE_N VGND VNB VPB VPWR Q
M1000 Q a_842_405# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.516e+11p pd=2.16e+06u as=1.54015e+12p ps=1.207e+07u
M1001 a_669_392# a_232_82# a_658_79# VNB nlowvt w=640000u l=150000u
+  ad=2.803e+11p pd=2.53e+06u as=1.536e+11p ps=1.76e+06u
M1002 a_658_79# a_27_120# VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1003 a_232_82# GATE_N VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1004 a_232_82# GATE_N VPWR VPB pshort w=840000u l=150000u
+  ad=2.478e+11p pd=2.27e+06u as=2.00335e+12p ps=1.509e+07u
M1005 VGND a_842_405# a_875_139# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1006 VPWR a_232_82# a_369_392# VPB pshort w=840000u l=150000u
+  ad=0p pd=0u as=2.478e+11p ps=2.27e+06u
M1007 Q a_842_405# VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=3.864e+11p pd=2.93e+06u as=0p ps=0u
M1008 VPWR D a_27_120# VPB pshort w=840000u l=150000u
+  ad=0p pd=0u as=2.478e+11p ps=2.27e+06u
M1009 VGND a_232_82# a_369_392# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1010 a_791_503# a_232_82# a_669_392# VPB pshort w=420000u l=150000u
+  ad=1.134e+11p pd=1.38e+06u as=4.05175e+11p ps=2.92e+06u
M1011 VPWR a_842_405# Q VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VGND a_842_405# Q VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VPWR a_842_405# a_791_503# VPB pshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_842_405# a_669_392# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1015 a_875_139# a_369_392# a_669_392# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_585_392# a_27_120# VPWR VPB pshort w=1e+06u l=150000u
+  ad=2.7e+11p pd=2.54e+06u as=0p ps=0u
M1017 VGND D a_27_120# VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=1.5675e+11p ps=1.67e+06u
M1018 a_669_392# a_369_392# a_585_392# VPB pshort w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_842_405# a_669_392# VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=3.304e+11p pd=2.83e+06u as=0p ps=0u
.ends

