* File: sky130_fd_sc_hs__dfrtn_1.pxi.spice
* Created: Thu Aug 27 20:38:30 2020
* 
x_PM_SKY130_FD_SC_HS__DFRTN_1%D N_D_c_240_n N_D_c_247_n N_D_c_248_n N_D_c_249_n
+ N_D_M1008_g N_D_M1029_g N_D_c_242_n N_D_c_243_n D D D N_D_c_244_n N_D_c_245_n
+ PM_SKY130_FD_SC_HS__DFRTN_1%D
x_PM_SKY130_FD_SC_HS__DFRTN_1%RESET_B N_RESET_B_M1024_g N_RESET_B_c_291_n
+ N_RESET_B_c_292_n N_RESET_B_M1007_g N_RESET_B_M1015_g N_RESET_B_c_293_n
+ N_RESET_B_c_294_n N_RESET_B_M1022_g N_RESET_B_M1012_g N_RESET_B_c_295_n
+ N_RESET_B_c_296_n N_RESET_B_M1025_g N_RESET_B_c_280_n N_RESET_B_c_281_n
+ N_RESET_B_c_282_n N_RESET_B_c_283_n N_RESET_B_c_284_n N_RESET_B_c_285_n
+ RESET_B N_RESET_B_c_286_n N_RESET_B_c_287_n N_RESET_B_c_288_n
+ N_RESET_B_c_289_n N_RESET_B_c_290_n PM_SKY130_FD_SC_HS__DFRTN_1%RESET_B
x_PM_SKY130_FD_SC_HS__DFRTN_1%CLK_N N_CLK_N_c_478_n N_CLK_N_M1027_g
+ N_CLK_N_c_479_n N_CLK_N_M1017_g CLK_N PM_SKY130_FD_SC_HS__DFRTN_1%CLK_N
x_PM_SKY130_FD_SC_HS__DFRTN_1%A_507_368# N_A_507_368#_M1010_d
+ N_A_507_368#_M1009_d N_A_507_368#_c_514_n N_A_507_368#_M1013_g
+ N_A_507_368#_c_535_n N_A_507_368#_c_536_n N_A_507_368#_c_537_n
+ N_A_507_368#_M1016_g N_A_507_368#_c_515_n N_A_507_368#_c_539_n
+ N_A_507_368#_M1011_g N_A_507_368#_c_516_n N_A_507_368#_c_517_n
+ N_A_507_368#_c_518_n N_A_507_368#_M1021_g N_A_507_368#_c_519_n
+ N_A_507_368#_c_520_n N_A_507_368#_c_541_n N_A_507_368#_c_542_n
+ N_A_507_368#_c_521_n N_A_507_368#_c_522_n N_A_507_368#_c_523_n
+ N_A_507_368#_c_551_n N_A_507_368#_c_563_p N_A_507_368#_c_524_n
+ N_A_507_368#_c_525_n N_A_507_368#_c_526_n N_A_507_368#_c_527_n
+ N_A_507_368#_c_553_n N_A_507_368#_c_554_n N_A_507_368#_c_528_n
+ N_A_507_368#_c_529_n N_A_507_368#_c_530_n N_A_507_368#_c_531_n
+ N_A_507_368#_c_532_n N_A_507_368#_c_533_n N_A_507_368#_c_534_n
+ PM_SKY130_FD_SC_HS__DFRTN_1%A_507_368#
x_PM_SKY130_FD_SC_HS__DFRTN_1%A_856_304# N_A_856_304#_M1019_d
+ N_A_856_304#_M1018_d N_A_856_304#_c_721_n N_A_856_304#_c_722_n
+ N_A_856_304#_M1004_g N_A_856_304#_M1026_g N_A_856_304#_c_714_n
+ N_A_856_304#_c_715_n N_A_856_304#_c_716_n N_A_856_304#_c_723_n
+ N_A_856_304#_c_717_n N_A_856_304#_c_718_n N_A_856_304#_c_719_n
+ N_A_856_304#_c_745_n N_A_856_304#_c_746_n N_A_856_304#_c_720_n
+ PM_SKY130_FD_SC_HS__DFRTN_1%A_856_304#
x_PM_SKY130_FD_SC_HS__DFRTN_1%A_714_127# N_A_714_127#_M1013_d
+ N_A_714_127#_M1014_d N_A_714_127#_M1022_d N_A_714_127#_M1019_g
+ N_A_714_127#_c_813_n N_A_714_127#_M1018_g N_A_714_127#_c_814_n
+ N_A_714_127#_c_815_n N_A_714_127#_c_816_n N_A_714_127#_c_822_n
+ N_A_714_127#_c_823_n N_A_714_127#_c_824_n N_A_714_127#_c_825_n
+ N_A_714_127#_c_817_n N_A_714_127#_c_827_n N_A_714_127#_c_818_n
+ N_A_714_127#_c_828_n PM_SKY130_FD_SC_HS__DFRTN_1%A_714_127#
x_PM_SKY130_FD_SC_HS__DFRTN_1%A_300_74# N_A_300_74#_M1027_d N_A_300_74#_M1017_d
+ N_A_300_74#_c_947_n N_A_300_74#_M1009_g N_A_300_74#_c_931_n
+ N_A_300_74#_M1010_g N_A_300_74#_c_932_n N_A_300_74#_c_933_n
+ N_A_300_74#_c_934_n N_A_300_74#_c_949_n N_A_300_74#_c_950_n
+ N_A_300_74#_c_951_n N_A_300_74#_M1014_g N_A_300_74#_M1030_g
+ N_A_300_74#_c_936_n N_A_300_74#_c_937_n N_A_300_74#_M1005_g
+ N_A_300_74#_c_952_n N_A_300_74#_M1006_g N_A_300_74#_c_939_n
+ N_A_300_74#_c_940_n N_A_300_74#_c_941_n N_A_300_74#_c_955_n
+ N_A_300_74#_c_956_n N_A_300_74#_c_942_n N_A_300_74#_c_943_n
+ N_A_300_74#_c_959_n N_A_300_74#_c_960_n N_A_300_74#_c_944_n
+ N_A_300_74#_c_945_n N_A_300_74#_c_946_n PM_SKY130_FD_SC_HS__DFRTN_1%A_300_74#
x_PM_SKY130_FD_SC_HS__DFRTN_1%A_1598_93# N_A_1598_93#_M1002_d
+ N_A_1598_93#_M1025_d N_A_1598_93#_M1000_g N_A_1598_93#_c_1141_n
+ N_A_1598_93#_M1023_g N_A_1598_93#_c_1142_n N_A_1598_93#_c_1143_n
+ N_A_1598_93#_c_1144_n N_A_1598_93#_c_1138_n N_A_1598_93#_c_1146_n
+ N_A_1598_93#_c_1139_n PM_SKY130_FD_SC_HS__DFRTN_1%A_1598_93#
x_PM_SKY130_FD_SC_HS__DFRTN_1%A_1266_119# N_A_1266_119#_M1005_d
+ N_A_1266_119#_M1011_d N_A_1266_119#_c_1226_n N_A_1266_119#_M1002_g
+ N_A_1266_119#_c_1227_n N_A_1266_119#_c_1237_n N_A_1266_119#_c_1238_n
+ N_A_1266_119#_M1031_g N_A_1266_119#_c_1228_n N_A_1266_119#_c_1239_n
+ N_A_1266_119#_c_1229_n N_A_1266_119#_M1020_g N_A_1266_119#_c_1240_n
+ N_A_1266_119#_M1003_g N_A_1266_119#_c_1230_n N_A_1266_119#_c_1266_n
+ N_A_1266_119#_c_1241_n N_A_1266_119#_c_1231_n N_A_1266_119#_c_1232_n
+ N_A_1266_119#_c_1233_n N_A_1266_119#_c_1243_n N_A_1266_119#_c_1274_n
+ N_A_1266_119#_c_1234_n N_A_1266_119#_c_1235_n
+ PM_SKY130_FD_SC_HS__DFRTN_1%A_1266_119#
x_PM_SKY130_FD_SC_HS__DFRTN_1%A_1934_94# N_A_1934_94#_M1020_s
+ N_A_1934_94#_M1003_s N_A_1934_94#_c_1364_n N_A_1934_94#_M1028_g
+ N_A_1934_94#_c_1365_n N_A_1934_94#_M1001_g N_A_1934_94#_c_1371_n
+ N_A_1934_94#_c_1372_n N_A_1934_94#_c_1366_n N_A_1934_94#_c_1367_n
+ N_A_1934_94#_c_1368_n N_A_1934_94#_c_1369_n
+ PM_SKY130_FD_SC_HS__DFRTN_1%A_1934_94#
x_PM_SKY130_FD_SC_HS__DFRTN_1%VPWR N_VPWR_M1008_s N_VPWR_M1007_d N_VPWR_M1009_s
+ N_VPWR_M1004_d N_VPWR_M1018_s N_VPWR_M1023_d N_VPWR_M1031_d N_VPWR_M1003_d
+ N_VPWR_c_1425_n N_VPWR_c_1426_n N_VPWR_c_1427_n N_VPWR_c_1428_n
+ N_VPWR_c_1429_n N_VPWR_c_1430_n N_VPWR_c_1431_n N_VPWR_c_1432_n
+ N_VPWR_c_1433_n N_VPWR_c_1434_n N_VPWR_c_1435_n N_VPWR_c_1436_n
+ N_VPWR_c_1437_n N_VPWR_c_1438_n VPWR N_VPWR_c_1439_n N_VPWR_c_1440_n
+ N_VPWR_c_1441_n N_VPWR_c_1442_n N_VPWR_c_1443_n N_VPWR_c_1424_n
+ N_VPWR_c_1445_n N_VPWR_c_1446_n N_VPWR_c_1447_n N_VPWR_c_1448_n
+ N_VPWR_c_1449_n PM_SKY130_FD_SC_HS__DFRTN_1%VPWR
x_PM_SKY130_FD_SC_HS__DFRTN_1%A_33_74# N_A_33_74#_M1029_s N_A_33_74#_M1013_s
+ N_A_33_74#_M1008_d N_A_33_74#_M1014_s N_A_33_74#_c_1558_n N_A_33_74#_c_1564_n
+ N_A_33_74#_c_1565_n N_A_33_74#_c_1566_n N_A_33_74#_c_1559_n
+ N_A_33_74#_c_1560_n N_A_33_74#_c_1634_n N_A_33_74#_c_1568_n
+ N_A_33_74#_c_1569_n N_A_33_74#_c_1561_n N_A_33_74#_c_1642_n
+ N_A_33_74#_c_1562_n PM_SKY130_FD_SC_HS__DFRTN_1%A_33_74#
x_PM_SKY130_FD_SC_HS__DFRTN_1%Q N_Q_M1028_d N_Q_M1001_d N_Q_c_1675_n
+ N_Q_c_1676_n Q Q Q Q N_Q_c_1677_n PM_SKY130_FD_SC_HS__DFRTN_1%Q
x_PM_SKY130_FD_SC_HS__DFRTN_1%VGND N_VGND_M1024_d N_VGND_M1010_s N_VGND_M1015_d
+ N_VGND_M1000_d N_VGND_M1020_d N_VGND_c_1703_n N_VGND_c_1704_n N_VGND_c_1705_n
+ N_VGND_c_1706_n N_VGND_c_1707_n VGND N_VGND_c_1708_n N_VGND_c_1709_n
+ N_VGND_c_1710_n N_VGND_c_1711_n N_VGND_c_1712_n N_VGND_c_1713_n
+ N_VGND_c_1714_n N_VGND_c_1715_n N_VGND_c_1716_n N_VGND_c_1717_n
+ N_VGND_c_1718_n N_VGND_c_1719_n PM_SKY130_FD_SC_HS__DFRTN_1%VGND
cc_1 VNB N_D_c_240_n 0.00193067f $X=-0.19 $Y=-0.245 $X2=0.36 $Y2=1.92
cc_2 VNB N_D_M1029_g 0.027501f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=0.58
cc_3 VNB N_D_c_242_n 0.0345854f $X=-0.19 $Y=-0.245 $X2=0.352 $Y2=1.11
cc_4 VNB N_D_c_243_n 0.0230272f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.63
cc_5 VNB N_D_c_244_n 0.0385312f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.125
cc_6 VNB N_D_c_245_n 0.00478024f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.125
cc_7 VNB N_RESET_B_M1024_g 0.044437f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=2.07
cc_8 VNB N_RESET_B_M1015_g 0.0385765f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.11
cc_9 VNB N_RESET_B_M1012_g 0.034399f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_10 VNB N_RESET_B_c_280_n 0.0201687f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.125
cc_11 VNB N_RESET_B_c_281_n 0.00278029f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.125
cc_12 VNB N_RESET_B_c_282_n 0.013881f $X=-0.19 $Y=-0.245 $X2=0.237 $Y2=1.125
cc_13 VNB N_RESET_B_c_283_n 5.71827e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_RESET_B_c_284_n 6.54175e-19 $X=-0.19 $Y=-0.245 $X2=0.237 $Y2=2.035
cc_15 VNB N_RESET_B_c_285_n 0.00357755f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_RESET_B_c_286_n 0.0286105f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_RESET_B_c_287_n 0.0157912f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_RESET_B_c_288_n 0.00223158f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_RESET_B_c_289_n 0.0154637f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_RESET_B_c_290_n 0.00440073f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_CLK_N_c_478_n 0.0208002f $X=-0.19 $Y=-0.245 $X2=0.36 $Y2=1.63
cc_22 VNB N_CLK_N_c_479_n 0.0400688f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=2.375
cc_23 VNB CLK_N 0.00545876f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=2.75
cc_24 VNB N_A_507_368#_c_514_n 0.0488801f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=0.58
cc_25 VNB N_A_507_368#_c_515_n 0.0165317f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_507_368#_c_516_n 0.0171653f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_507_368#_c_517_n 0.0191633f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_507_368#_c_518_n 0.0231425f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.125
cc_29 VNB N_A_507_368#_c_519_n 0.0018344f $X=-0.19 $Y=-0.245 $X2=0.237 $Y2=1.295
cc_30 VNB N_A_507_368#_c_520_n 0.00885409f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_507_368#_c_521_n 0.00308204f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_507_368#_c_522_n 0.0147543f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_507_368#_c_523_n 0.00195044f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_507_368#_c_524_n 0.0039155f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_507_368#_c_525_n 0.0193653f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_507_368#_c_526_n 0.00260538f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_507_368#_c_527_n 0.00739636f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_507_368#_c_528_n 0.00166696f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_507_368#_c_529_n 0.0294493f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_507_368#_c_530_n 0.00474842f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_507_368#_c_531_n 0.00605204f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_507_368#_c_532_n 0.0458542f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_507_368#_c_533_n 0.00628108f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_507_368#_c_534_n 0.0169284f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_A_856_304#_M1026_g 0.0297395f $X=-0.19 $Y=-0.245 $X2=0.352 $Y2=1.11
cc_46 VNB N_A_856_304#_c_714_n 0.0155687f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_856_304#_c_715_n 0.00162463f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=1.995
cc_48 VNB N_A_856_304#_c_716_n 0.00112198f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_49 VNB N_A_856_304#_c_717_n 0.00277557f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_A_856_304#_c_718_n 0.0171047f $X=-0.19 $Y=-0.245 $X2=0.237 $Y2=1.295
cc_51 VNB N_A_856_304#_c_719_n 0.00207547f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_A_856_304#_c_720_n 0.0021497f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_A_714_127#_M1019_g 0.0201455f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.11
cc_54 VNB N_A_714_127#_c_813_n 0.0093697f $X=-0.19 $Y=-0.245 $X2=0.352 $Y2=1.11
cc_55 VNB N_A_714_127#_c_814_n 0.0216047f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_A_714_127#_c_815_n 0.0014057f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_57 VNB N_A_714_127#_c_816_n 0.00663354f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_A_714_127#_c_817_n 0.00306892f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_A_714_127#_c_818_n 3.87698e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_A_300_74#_c_931_n 0.019408f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=0.58
cc_61 VNB N_A_300_74#_c_932_n 0.024949f $X=-0.19 $Y=-0.245 $X2=0.352 $Y2=0.96
cc_62 VNB N_A_300_74#_c_933_n 0.00502702f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.63
cc_63 VNB N_A_300_74#_c_934_n 0.0835617f $X=-0.19 $Y=-0.245 $X2=0.36 $Y2=1.995
cc_64 VNB N_A_300_74#_M1030_g 0.0270717f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.125
cc_65 VNB N_A_300_74#_c_936_n 0.150233f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.125
cc_66 VNB N_A_300_74#_c_937_n 0.0116916f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.125
cc_67 VNB N_A_300_74#_M1005_g 0.030044f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_A_300_74#_c_939_n 0.0371644f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_A_300_74#_c_940_n 0.0103095f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_A_300_74#_c_941_n 0.0066402f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_A_300_74#_c_942_n 0.00453807f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_A_300_74#_c_943_n 0.00454971f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_A_300_74#_c_944_n 0.0161152f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_A_300_74#_c_945_n 0.00265148f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_A_300_74#_c_946_n 0.018162f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_A_1598_93#_M1000_g 0.0473326f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=0.58
cc_77 VNB N_A_1598_93#_c_1138_n 0.0107986f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_A_1598_93#_c_1139_n 0.0121095f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VNB N_A_1266_119#_c_1226_n 0.0202606f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=2.75
cc_80 VNB N_A_1266_119#_c_1227_n 0.00226217f $X=-0.19 $Y=-0.245 $X2=0.525
+ $Y2=0.58
cc_81 VNB N_A_1266_119#_c_1228_n 0.0586053f $X=-0.19 $Y=-0.245 $X2=0.27
+ $Y2=1.465
cc_82 VNB N_A_1266_119#_c_1229_n 0.0219742f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=1.995
cc_83 VNB N_A_1266_119#_c_1230_n 0.00948676f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_84 VNB N_A_1266_119#_c_1231_n 0.00100139f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_85 VNB N_A_1266_119#_c_1232_n 0.0107396f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_86 VNB N_A_1266_119#_c_1233_n 0.0235899f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_87 VNB N_A_1266_119#_c_1234_n 5.53899e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_88 VNB N_A_1266_119#_c_1235_n 0.024655f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_89 VNB N_A_1934_94#_c_1364_n 0.0213736f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=2.75
cc_90 VNB N_A_1934_94#_c_1365_n 0.0409762f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=0.58
cc_91 VNB N_A_1934_94#_c_1366_n 0.00180273f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=1.995
cc_92 VNB N_A_1934_94#_c_1367_n 2.65185e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_93 VNB N_A_1934_94#_c_1368_n 0.0106069f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.125
cc_94 VNB N_A_1934_94#_c_1369_n 0.00429191f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_95 VNB N_VPWR_c_1424_n 0.462217f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_96 VNB N_A_33_74#_c_1558_n 0.0122231f $X=-0.19 $Y=-0.245 $X2=0.352 $Y2=1.11
cc_97 VNB N_A_33_74#_c_1559_n 8.35165e-19 $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_98 VNB N_A_33_74#_c_1560_n 0.00632162f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.95
cc_99 VNB N_A_33_74#_c_1561_n 0.0216357f $X=-0.19 $Y=-0.245 $X2=0.237 $Y2=1.665
cc_100 VNB N_A_33_74#_c_1562_n 0.00670563f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_101 VNB N_Q_c_1675_n 0.0243417f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=0.58
cc_102 VNB N_Q_c_1676_n 0.00719696f $X=-0.19 $Y=-0.245 $X2=0.352 $Y2=0.96
cc_103 VNB N_Q_c_1677_n 0.0236409f $X=-0.19 $Y=-0.245 $X2=0.237 $Y2=1.295
cc_104 VNB N_VGND_c_1703_n 0.0093175f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_105 VNB N_VGND_c_1704_n 0.0115761f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_106 VNB N_VGND_c_1705_n 0.00866422f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_107 VNB N_VGND_c_1706_n 0.0246564f $X=-0.19 $Y=-0.245 $X2=0.237 $Y2=1.125
cc_108 VNB N_VGND_c_1707_n 0.017712f $X=-0.19 $Y=-0.245 $X2=0.237 $Y2=1.665
cc_109 VNB N_VGND_c_1708_n 0.0309922f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_110 VNB N_VGND_c_1709_n 0.0194767f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_111 VNB N_VGND_c_1710_n 0.067058f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_112 VNB N_VGND_c_1711_n 0.0716605f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_113 VNB N_VGND_c_1712_n 0.0470737f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_114 VNB N_VGND_c_1713_n 0.0198148f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_115 VNB N_VGND_c_1714_n 0.606817f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_116 VNB N_VGND_c_1715_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_117 VNB N_VGND_c_1716_n 0.00631443f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_118 VNB N_VGND_c_1717_n 0.0043699f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_119 VNB N_VGND_c_1718_n 0.00846329f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_120 VNB N_VGND_c_1719_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_121 VPB N_D_c_240_n 0.0175703f $X=-0.19 $Y=1.66 $X2=0.36 $Y2=1.92
cc_122 VPB N_D_c_247_n 0.0220469f $X=-0.19 $Y=1.66 $X2=0.5 $Y2=2.07
cc_123 VPB N_D_c_248_n 0.0222831f $X=-0.19 $Y=1.66 $X2=0.5 $Y2=2.375
cc_124 VPB N_D_c_249_n 0.0276024f $X=-0.19 $Y=1.66 $X2=0.5 $Y2=2.465
cc_125 VPB N_D_c_245_n 0.0217648f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.125
cc_126 VPB N_RESET_B_c_291_n 0.0394534f $X=-0.19 $Y=1.66 $X2=0.5 $Y2=2.75
cc_127 VPB N_RESET_B_c_292_n 0.0220066f $X=-0.19 $Y=1.66 $X2=0.5 $Y2=2.75
cc_128 VPB N_RESET_B_c_293_n 0.0376165f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.465
cc_129 VPB N_RESET_B_c_294_n 0.0257859f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.63
cc_130 VPB N_RESET_B_c_295_n 0.0283395f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_131 VPB N_RESET_B_c_296_n 0.0223436f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_132 VPB N_RESET_B_c_280_n 0.0167338f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.125
cc_133 VPB N_RESET_B_c_281_n 0.00350731f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.125
cc_134 VPB N_RESET_B_c_282_n 0.00673887f $X=-0.19 $Y=1.66 $X2=0.237 $Y2=1.125
cc_135 VPB N_RESET_B_c_283_n 5.68911e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_136 VPB N_RESET_B_c_284_n 6.35107e-19 $X=-0.19 $Y=1.66 $X2=0.237 $Y2=2.035
cc_137 VPB N_RESET_B_c_285_n 0.00257552f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_138 VPB N_RESET_B_c_286_n 0.00580778f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_139 VPB N_RESET_B_c_287_n 0.0106707f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_140 VPB N_RESET_B_c_288_n 0.00127854f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_141 VPB N_RESET_B_c_289_n 0.0112707f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_142 VPB N_RESET_B_c_290_n 0.00294651f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_143 VPB N_CLK_N_c_479_n 0.0252199f $X=-0.19 $Y=1.66 $X2=0.5 $Y2=2.375
cc_144 VPB N_A_507_368#_c_535_n 0.0236638f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.11
cc_145 VPB N_A_507_368#_c_536_n 0.0157267f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.465
cc_146 VPB N_A_507_368#_c_537_n 0.0207289f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.63
cc_147 VPB N_A_507_368#_c_515_n 0.00582876f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_148 VPB N_A_507_368#_c_539_n 0.0310581f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.21
cc_149 VPB N_A_507_368#_c_519_n 0.00333529f $X=-0.19 $Y=1.66 $X2=0.237 $Y2=1.295
cc_150 VPB N_A_507_368#_c_541_n 0.00484614f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_151 VPB N_A_507_368#_c_542_n 0.0306901f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_152 VPB N_A_856_304#_c_721_n 0.0285873f $X=-0.19 $Y=1.66 $X2=0.525 $Y2=0.96
cc_153 VPB N_A_856_304#_c_722_n 0.0214741f $X=-0.19 $Y=1.66 $X2=0.525 $Y2=0.58
cc_154 VPB N_A_856_304#_c_723_n 0.00690074f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.125
cc_155 VPB N_A_856_304#_c_717_n 0.00138754f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_156 VPB N_A_856_304#_c_718_n 0.0180227f $X=-0.19 $Y=1.66 $X2=0.237 $Y2=1.295
cc_157 VPB N_A_856_304#_c_720_n 0.00306186f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_158 VPB N_A_714_127#_c_813_n 0.0340256f $X=-0.19 $Y=1.66 $X2=0.352 $Y2=1.11
cc_159 VPB N_A_714_127#_c_814_n 0.017529f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_160 VPB N_A_714_127#_c_816_n 0.00499466f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_161 VPB N_A_714_127#_c_822_n 0.00622025f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_162 VPB N_A_714_127#_c_823_n 0.017859f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.125
cc_163 VPB N_A_714_127#_c_824_n 0.0126793f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_164 VPB N_A_714_127#_c_825_n 0.0137564f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_165 VPB N_A_714_127#_c_817_n 0.00436057f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_166 VPB N_A_714_127#_c_827_n 0.00568939f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_167 VPB N_A_714_127#_c_828_n 0.00346183f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_168 VPB N_A_300_74#_c_947_n 0.0214657f $X=-0.19 $Y=1.66 $X2=0.5 $Y2=2.75
cc_169 VPB N_A_300_74#_c_933_n 0.037939f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.63
cc_170 VPB N_A_300_74#_c_949_n 0.0322163f $X=-0.19 $Y=1.66 $X2=0.5 $Y2=1.995
cc_171 VPB N_A_300_74#_c_950_n 0.00953795f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_172 VPB N_A_300_74#_c_951_n 0.0192231f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.21
cc_173 VPB N_A_300_74#_c_952_n 0.0178649f $X=-0.19 $Y=1.66 $X2=0.237 $Y2=1.665
cc_174 VPB N_A_300_74#_c_939_n 0.0152429f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_175 VPB N_A_300_74#_c_940_n 0.00751241f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_176 VPB N_A_300_74#_c_955_n 0.0322371f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_177 VPB N_A_300_74#_c_956_n 0.0087286f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_178 VPB N_A_300_74#_c_942_n 0.0021356f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_179 VPB N_A_300_74#_c_943_n 0.0168815f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_180 VPB N_A_300_74#_c_959_n 0.00232654f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_181 VPB N_A_300_74#_c_960_n 0.0463369f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_182 VPB N_A_300_74#_c_945_n 0.00280482f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_183 VPB N_A_300_74#_c_946_n 0.0167017f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_184 VPB N_A_1598_93#_M1000_g 0.01871f $X=-0.19 $Y=1.66 $X2=0.525 $Y2=0.58
cc_185 VPB N_A_1598_93#_c_1141_n 0.0544767f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_186 VPB N_A_1598_93#_c_1142_n 0.00706063f $X=-0.19 $Y=1.66 $X2=0.352 $Y2=1.11
cc_187 VPB N_A_1598_93#_c_1143_n 0.00257348f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.21
cc_188 VPB N_A_1598_93#_c_1144_n 0.00961486f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.95
cc_189 VPB N_A_1598_93#_c_1138_n 0.00471733f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_190 VPB N_A_1598_93#_c_1146_n 0.00400474f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.125
cc_191 VPB N_A_1266_119#_c_1227_n 0.023609f $X=-0.19 $Y=1.66 $X2=0.525 $Y2=0.58
cc_192 VPB N_A_1266_119#_c_1237_n 0.0201446f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_193 VPB N_A_1266_119#_c_1238_n 0.0231244f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.11
cc_194 VPB N_A_1266_119#_c_1239_n 0.059564f $X=-0.19 $Y=1.66 $X2=0.36 $Y2=1.995
cc_195 VPB N_A_1266_119#_c_1240_n 0.0184812f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_196 VPB N_A_1266_119#_c_1241_n 0.00674641f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_197 VPB N_A_1266_119#_c_1232_n 0.0132664f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_198 VPB N_A_1266_119#_c_1243_n 0.00103675f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_199 VPB N_A_1266_119#_c_1234_n 5.52803e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_200 VPB N_A_1934_94#_c_1365_n 0.0302218f $X=-0.19 $Y=1.66 $X2=0.525 $Y2=0.58
cc_201 VPB N_A_1934_94#_c_1371_n 0.00268013f $X=-0.19 $Y=1.66 $X2=0.352 $Y2=0.96
cc_202 VPB N_A_1934_94#_c_1372_n 0.00754272f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.465
cc_203 VPB N_A_1934_94#_c_1367_n 0.0059282f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_204 VPB N_VPWR_c_1425_n 0.0117486f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_205 VPB N_VPWR_c_1426_n 0.0301445f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.125
cc_206 VPB N_VPWR_c_1427_n 0.00577735f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_207 VPB N_VPWR_c_1428_n 0.0120309f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_208 VPB N_VPWR_c_1429_n 0.0102968f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_209 VPB N_VPWR_c_1430_n 0.0196495f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_210 VPB N_VPWR_c_1431_n 0.0127233f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_211 VPB N_VPWR_c_1432_n 0.00931072f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_212 VPB N_VPWR_c_1433_n 0.0161288f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_213 VPB N_VPWR_c_1434_n 0.00977211f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_214 VPB N_VPWR_c_1435_n 0.0619705f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_215 VPB N_VPWR_c_1436_n 0.00614127f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_216 VPB N_VPWR_c_1437_n 0.0193312f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_217 VPB N_VPWR_c_1438_n 0.0047828f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_218 VPB N_VPWR_c_1439_n 0.0175706f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_219 VPB N_VPWR_c_1440_n 0.0214173f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_220 VPB N_VPWR_c_1441_n 0.0598398f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_221 VPB N_VPWR_c_1442_n 0.0209223f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_222 VPB N_VPWR_c_1443_n 0.0197908f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_223 VPB N_VPWR_c_1424_n 0.137623f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_224 VPB N_VPWR_c_1445_n 0.00614589f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_225 VPB N_VPWR_c_1446_n 0.00614127f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_226 VPB N_VPWR_c_1447_n 0.00614127f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_227 VPB N_VPWR_c_1448_n 0.00614127f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_228 VPB N_VPWR_c_1449_n 0.0047828f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_229 VPB N_A_33_74#_c_1558_n 0.00638159f $X=-0.19 $Y=1.66 $X2=0.352 $Y2=1.11
cc_230 VPB N_A_33_74#_c_1564_n 0.00391661f $X=-0.19 $Y=1.66 $X2=0.36 $Y2=1.995
cc_231 VPB N_A_33_74#_c_1565_n 0.00826827f $X=-0.19 $Y=1.66 $X2=0.5 $Y2=1.995
cc_232 VPB N_A_33_74#_c_1566_n 0.00856541f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_233 VPB N_A_33_74#_c_1559_n 0.00114288f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_234 VPB N_A_33_74#_c_1568_n 0.0074189f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_235 VPB N_A_33_74#_c_1569_n 0.0105105f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.125
cc_236 VPB Q 0.00930674f $X=-0.19 $Y=1.66 $X2=0.352 $Y2=1.11
cc_237 VPB Q 0.0416636f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.95
cc_238 VPB N_Q_c_1677_n 0.00772285f $X=-0.19 $Y=1.66 $X2=0.237 $Y2=1.295
cc_239 N_D_M1029_g N_RESET_B_M1024_g 0.0435282f $X=0.525 $Y=0.58 $X2=0 $Y2=0
cc_240 N_D_c_244_n N_RESET_B_M1024_g 0.00520474f $X=0.27 $Y=1.125 $X2=0 $Y2=0
cc_241 N_D_c_240_n N_RESET_B_c_291_n 0.00462577f $X=0.36 $Y=1.92 $X2=0 $Y2=0
cc_242 N_D_c_247_n N_RESET_B_c_291_n 0.0120295f $X=0.5 $Y=2.07 $X2=0 $Y2=0
cc_243 N_D_c_248_n N_RESET_B_c_292_n 0.0120295f $X=0.5 $Y=2.375 $X2=0 $Y2=0
cc_244 N_D_c_249_n N_RESET_B_c_292_n 0.00873326f $X=0.5 $Y=2.465 $X2=0 $Y2=0
cc_245 N_D_c_244_n N_RESET_B_c_286_n 0.00843167f $X=0.27 $Y=1.125 $X2=0 $Y2=0
cc_246 N_D_c_247_n N_VPWR_c_1426_n 0.00199186f $X=0.5 $Y=2.07 $X2=0 $Y2=0
cc_247 N_D_c_249_n N_VPWR_c_1426_n 0.0120884f $X=0.5 $Y=2.465 $X2=0 $Y2=0
cc_248 N_D_c_245_n N_VPWR_c_1426_n 0.0140568f $X=0.27 $Y=1.125 $X2=0 $Y2=0
cc_249 N_D_c_249_n N_VPWR_c_1439_n 0.00413917f $X=0.5 $Y=2.465 $X2=0 $Y2=0
cc_250 N_D_c_249_n N_VPWR_c_1424_n 0.00853987f $X=0.5 $Y=2.465 $X2=0 $Y2=0
cc_251 N_D_c_247_n N_A_33_74#_c_1558_n 0.00493271f $X=0.5 $Y=2.07 $X2=0 $Y2=0
cc_252 N_D_c_248_n N_A_33_74#_c_1558_n 0.00297569f $X=0.5 $Y=2.375 $X2=0 $Y2=0
cc_253 N_D_M1029_g N_A_33_74#_c_1558_n 0.00857134f $X=0.525 $Y=0.58 $X2=0 $Y2=0
cc_254 N_D_c_242_n N_A_33_74#_c_1558_n 0.00517676f $X=0.352 $Y=1.11 $X2=0 $Y2=0
cc_255 N_D_c_244_n N_A_33_74#_c_1558_n 0.00670016f $X=0.27 $Y=1.125 $X2=0 $Y2=0
cc_256 N_D_c_245_n N_A_33_74#_c_1558_n 0.0866708f $X=0.27 $Y=1.125 $X2=0 $Y2=0
cc_257 N_D_c_248_n N_A_33_74#_c_1564_n 0.00295199f $X=0.5 $Y=2.375 $X2=0 $Y2=0
cc_258 N_D_c_249_n N_A_33_74#_c_1564_n 0.00329762f $X=0.5 $Y=2.465 $X2=0 $Y2=0
cc_259 N_D_c_248_n N_A_33_74#_c_1566_n 0.0128044f $X=0.5 $Y=2.375 $X2=0 $Y2=0
cc_260 N_D_M1029_g N_A_33_74#_c_1561_n 0.0152419f $X=0.525 $Y=0.58 $X2=0 $Y2=0
cc_261 N_D_c_242_n N_A_33_74#_c_1561_n 0.0040449f $X=0.352 $Y=1.11 $X2=0 $Y2=0
cc_262 N_D_c_245_n N_A_33_74#_c_1561_n 0.0188861f $X=0.27 $Y=1.125 $X2=0 $Y2=0
cc_263 N_D_M1029_g N_VGND_c_1708_n 0.00291649f $X=0.525 $Y=0.58 $X2=0 $Y2=0
cc_264 N_D_M1029_g N_VGND_c_1714_n 0.00362587f $X=0.525 $Y=0.58 $X2=0 $Y2=0
cc_265 N_RESET_B_M1024_g N_CLK_N_c_478_n 0.0270985f $X=0.915 $Y=0.58 $X2=-0.19
+ $Y2=-0.245
cc_266 N_RESET_B_c_291_n N_CLK_N_c_479_n 0.0266963f $X=0.95 $Y=2.375 $X2=0 $Y2=0
cc_267 N_RESET_B_c_292_n N_CLK_N_c_479_n 0.0130184f $X=0.95 $Y=2.465 $X2=0 $Y2=0
cc_268 N_RESET_B_c_280_n N_CLK_N_c_479_n 0.0146119f $X=4.895 $Y=1.665 $X2=0
+ $Y2=0
cc_269 N_RESET_B_c_281_n N_CLK_N_c_479_n 0.00153261f $X=1.345 $Y=1.665 $X2=0
+ $Y2=0
cc_270 N_RESET_B_c_286_n N_CLK_N_c_479_n 0.0201394f $X=0.975 $Y=1.515 $X2=0
+ $Y2=0
cc_271 N_RESET_B_c_290_n N_CLK_N_c_479_n 0.00400589f $X=1.2 $Y=1.665 $X2=0 $Y2=0
cc_272 N_RESET_B_M1024_g CLK_N 8.20196e-19 $X=0.915 $Y=0.58 $X2=0 $Y2=0
cc_273 N_RESET_B_c_280_n CLK_N 0.0106116f $X=4.895 $Y=1.665 $X2=0 $Y2=0
cc_274 N_RESET_B_c_290_n CLK_N 0.0160113f $X=1.2 $Y=1.665 $X2=0 $Y2=0
cc_275 N_RESET_B_c_280_n N_A_507_368#_c_535_n 0.0025283f $X=4.895 $Y=1.665 $X2=0
+ $Y2=0
cc_276 N_RESET_B_c_282_n N_A_507_368#_c_515_n 0.00221676f $X=8.255 $Y=1.665
+ $X2=0 $Y2=0
cc_277 N_RESET_B_c_282_n N_A_507_368#_c_517_n 0.00405791f $X=8.255 $Y=1.665
+ $X2=0 $Y2=0
cc_278 N_RESET_B_c_280_n N_A_507_368#_c_519_n 0.0231711f $X=4.895 $Y=1.665 $X2=0
+ $Y2=0
cc_279 N_RESET_B_c_280_n N_A_507_368#_c_520_n 0.0202117f $X=4.895 $Y=1.665 $X2=0
+ $Y2=0
cc_280 N_RESET_B_c_280_n N_A_507_368#_c_541_n 0.0253267f $X=4.895 $Y=1.665 $X2=0
+ $Y2=0
cc_281 N_RESET_B_c_280_n N_A_507_368#_c_542_n 0.00464699f $X=4.895 $Y=1.665
+ $X2=0 $Y2=0
cc_282 N_RESET_B_M1015_g N_A_507_368#_c_523_n 0.00114254f $X=4.895 $Y=0.845
+ $X2=0 $Y2=0
cc_283 N_RESET_B_M1015_g N_A_507_368#_c_551_n 0.0113412f $X=4.895 $Y=0.845 $X2=0
+ $Y2=0
cc_284 N_RESET_B_M1015_g N_A_507_368#_c_524_n 0.00400898f $X=4.895 $Y=0.845
+ $X2=0 $Y2=0
cc_285 N_RESET_B_c_282_n N_A_507_368#_c_553_n 0.00155657f $X=8.255 $Y=1.665
+ $X2=0 $Y2=0
cc_286 N_RESET_B_c_282_n N_A_507_368#_c_554_n 0.0169144f $X=8.255 $Y=1.665 $X2=0
+ $Y2=0
cc_287 N_RESET_B_c_282_n N_A_507_368#_c_529_n 0.011489f $X=8.255 $Y=1.665 $X2=0
+ $Y2=0
cc_288 N_RESET_B_c_282_n N_A_507_368#_c_533_n 0.00501712f $X=8.255 $Y=1.665
+ $X2=0 $Y2=0
cc_289 N_RESET_B_c_293_n N_A_856_304#_c_721_n 0.0123779f $X=4.91 $Y=2.375 $X2=0
+ $Y2=0
cc_290 N_RESET_B_c_294_n N_A_856_304#_c_722_n 0.0240847f $X=4.91 $Y=2.465 $X2=0
+ $Y2=0
cc_291 N_RESET_B_M1015_g N_A_856_304#_M1026_g 0.0423195f $X=4.895 $Y=0.845 $X2=0
+ $Y2=0
cc_292 N_RESET_B_c_288_n N_A_856_304#_M1026_g 0.00110316f $X=4.985 $Y=1.635
+ $X2=0 $Y2=0
cc_293 N_RESET_B_M1015_g N_A_856_304#_c_714_n 0.0119822f $X=4.895 $Y=0.845 $X2=0
+ $Y2=0
cc_294 N_RESET_B_c_280_n N_A_856_304#_c_714_n 0.00880086f $X=4.895 $Y=1.665
+ $X2=0 $Y2=0
cc_295 N_RESET_B_c_282_n N_A_856_304#_c_714_n 0.014851f $X=8.255 $Y=1.665 $X2=0
+ $Y2=0
cc_296 N_RESET_B_c_283_n N_A_856_304#_c_714_n 0.00289579f $X=5.185 $Y=1.665
+ $X2=0 $Y2=0
cc_297 N_RESET_B_c_287_n N_A_856_304#_c_714_n 0.0041539f $X=4.985 $Y=1.635 $X2=0
+ $Y2=0
cc_298 N_RESET_B_c_288_n N_A_856_304#_c_714_n 0.0227858f $X=4.985 $Y=1.635 $X2=0
+ $Y2=0
cc_299 N_RESET_B_c_280_n N_A_856_304#_c_717_n 0.0276574f $X=4.895 $Y=1.665 $X2=0
+ $Y2=0
cc_300 N_RESET_B_c_283_n N_A_856_304#_c_717_n 5.41012e-19 $X=5.185 $Y=1.665
+ $X2=0 $Y2=0
cc_301 N_RESET_B_c_287_n N_A_856_304#_c_717_n 3.43048e-19 $X=4.985 $Y=1.635
+ $X2=0 $Y2=0
cc_302 N_RESET_B_c_280_n N_A_856_304#_c_718_n 0.00299097f $X=4.895 $Y=1.665
+ $X2=0 $Y2=0
cc_303 N_RESET_B_c_287_n N_A_856_304#_c_718_n 0.0423195f $X=4.985 $Y=1.635 $X2=0
+ $Y2=0
cc_304 N_RESET_B_M1015_g N_A_856_304#_c_719_n 0.00114614f $X=4.895 $Y=0.845
+ $X2=0 $Y2=0
cc_305 N_RESET_B_c_287_n N_A_856_304#_c_719_n 5.12513e-19 $X=4.985 $Y=1.635
+ $X2=0 $Y2=0
cc_306 N_RESET_B_c_288_n N_A_856_304#_c_719_n 0.0184766f $X=4.985 $Y=1.635 $X2=0
+ $Y2=0
cc_307 N_RESET_B_c_282_n N_A_856_304#_c_745_n 0.00468242f $X=8.255 $Y=1.665
+ $X2=0 $Y2=0
cc_308 N_RESET_B_c_282_n N_A_856_304#_c_746_n 0.00919057f $X=8.255 $Y=1.665
+ $X2=0 $Y2=0
cc_309 N_RESET_B_c_282_n N_A_856_304#_c_720_n 0.0226321f $X=8.255 $Y=1.665 $X2=0
+ $Y2=0
cc_310 N_RESET_B_c_282_n N_A_714_127#_c_813_n 0.00611789f $X=8.255 $Y=1.665
+ $X2=0 $Y2=0
cc_311 N_RESET_B_c_282_n N_A_714_127#_c_814_n 0.00272004f $X=8.255 $Y=1.665
+ $X2=0 $Y2=0
cc_312 N_RESET_B_c_283_n N_A_714_127#_c_814_n 0.00140145f $X=5.185 $Y=1.665
+ $X2=0 $Y2=0
cc_313 N_RESET_B_c_287_n N_A_714_127#_c_814_n 0.0214999f $X=4.985 $Y=1.635 $X2=0
+ $Y2=0
cc_314 N_RESET_B_c_288_n N_A_714_127#_c_814_n 0.00169603f $X=4.985 $Y=1.635
+ $X2=0 $Y2=0
cc_315 N_RESET_B_c_280_n N_A_714_127#_c_816_n 0.0180232f $X=4.895 $Y=1.665 $X2=0
+ $Y2=0
cc_316 N_RESET_B_c_293_n N_A_714_127#_c_823_n 0.0133901f $X=4.91 $Y=2.375 $X2=0
+ $Y2=0
cc_317 N_RESET_B_c_280_n N_A_714_127#_c_823_n 0.0198714f $X=4.895 $Y=1.665 $X2=0
+ $Y2=0
cc_318 N_RESET_B_c_283_n N_A_714_127#_c_823_n 0.00176425f $X=5.185 $Y=1.665
+ $X2=0 $Y2=0
cc_319 N_RESET_B_c_288_n N_A_714_127#_c_823_n 0.017712f $X=4.985 $Y=1.635 $X2=0
+ $Y2=0
cc_320 N_RESET_B_c_293_n N_A_714_127#_c_824_n 0.00748522f $X=4.91 $Y=2.375 $X2=0
+ $Y2=0
cc_321 N_RESET_B_c_294_n N_A_714_127#_c_824_n 0.0121385f $X=4.91 $Y=2.465 $X2=0
+ $Y2=0
cc_322 N_RESET_B_c_293_n N_A_714_127#_c_825_n 0.00501433f $X=4.91 $Y=2.375 $X2=0
+ $Y2=0
cc_323 N_RESET_B_c_282_n N_A_714_127#_c_825_n 0.0084368f $X=8.255 $Y=1.665 $X2=0
+ $Y2=0
cc_324 N_RESET_B_c_283_n N_A_714_127#_c_825_n 0.00133381f $X=5.185 $Y=1.665
+ $X2=0 $Y2=0
cc_325 N_RESET_B_c_287_n N_A_714_127#_c_825_n 0.00325305f $X=4.985 $Y=1.635
+ $X2=0 $Y2=0
cc_326 N_RESET_B_c_293_n N_A_714_127#_c_817_n 0.00674835f $X=4.91 $Y=2.375 $X2=0
+ $Y2=0
cc_327 N_RESET_B_c_282_n N_A_714_127#_c_817_n 0.0166072f $X=8.255 $Y=1.665 $X2=0
+ $Y2=0
cc_328 N_RESET_B_c_283_n N_A_714_127#_c_817_n 0.00259167f $X=5.185 $Y=1.665
+ $X2=0 $Y2=0
cc_329 N_RESET_B_c_287_n N_A_714_127#_c_817_n 5.08278e-19 $X=4.985 $Y=1.635
+ $X2=0 $Y2=0
cc_330 N_RESET_B_c_288_n N_A_714_127#_c_817_n 0.0191898f $X=4.985 $Y=1.635 $X2=0
+ $Y2=0
cc_331 N_RESET_B_c_280_n N_A_714_127#_c_818_n 0.00271395f $X=4.895 $Y=1.665
+ $X2=0 $Y2=0
cc_332 N_RESET_B_c_280_n N_A_300_74#_c_932_n 8.18829e-19 $X=4.895 $Y=1.665 $X2=0
+ $Y2=0
cc_333 N_RESET_B_c_280_n N_A_300_74#_c_933_n 0.00594403f $X=4.895 $Y=1.665 $X2=0
+ $Y2=0
cc_334 N_RESET_B_c_280_n N_A_300_74#_c_934_n 0.0172561f $X=4.895 $Y=1.665 $X2=0
+ $Y2=0
cc_335 N_RESET_B_M1015_g N_A_300_74#_c_936_n 0.00816399f $X=4.895 $Y=0.845 $X2=0
+ $Y2=0
cc_336 N_RESET_B_c_280_n N_A_300_74#_c_939_n 0.00887879f $X=4.895 $Y=1.665 $X2=0
+ $Y2=0
cc_337 N_RESET_B_c_280_n N_A_300_74#_c_940_n 0.00376569f $X=4.895 $Y=1.665 $X2=0
+ $Y2=0
cc_338 N_RESET_B_c_282_n N_A_300_74#_c_955_n 2.3419e-19 $X=8.255 $Y=1.665 $X2=0
+ $Y2=0
cc_339 N_RESET_B_c_291_n N_A_300_74#_c_956_n 0.00152784f $X=0.95 $Y=2.375 $X2=0
+ $Y2=0
cc_340 N_RESET_B_c_280_n N_A_300_74#_c_956_n 0.0164168f $X=4.895 $Y=1.665 $X2=0
+ $Y2=0
cc_341 N_RESET_B_c_280_n N_A_300_74#_c_942_n 0.0248558f $X=4.895 $Y=1.665 $X2=0
+ $Y2=0
cc_342 N_RESET_B_c_281_n N_A_300_74#_c_942_n 0.00197244f $X=1.345 $Y=1.665 $X2=0
+ $Y2=0
cc_343 N_RESET_B_c_290_n N_A_300_74#_c_942_n 0.00326944f $X=1.2 $Y=1.665 $X2=0
+ $Y2=0
cc_344 N_RESET_B_c_282_n N_A_300_74#_c_943_n 0.0603286f $X=8.255 $Y=1.665 $X2=0
+ $Y2=0
cc_345 N_RESET_B_c_282_n N_A_300_74#_c_960_n 0.00727375f $X=8.255 $Y=1.665 $X2=0
+ $Y2=0
cc_346 N_RESET_B_M1024_g N_A_300_74#_c_944_n 0.00104412f $X=0.915 $Y=0.58 $X2=0
+ $Y2=0
cc_347 N_RESET_B_c_280_n N_A_300_74#_c_944_n 0.0062195f $X=4.895 $Y=1.665 $X2=0
+ $Y2=0
cc_348 N_RESET_B_c_282_n N_A_300_74#_c_945_n 0.0194318f $X=8.255 $Y=1.665 $X2=0
+ $Y2=0
cc_349 N_RESET_B_c_282_n N_A_300_74#_c_946_n 0.00169661f $X=8.255 $Y=1.665 $X2=0
+ $Y2=0
cc_350 N_RESET_B_M1012_g N_A_1598_93#_M1000_g 0.0206165f $X=8.605 $Y=0.805 $X2=0
+ $Y2=0
cc_351 N_RESET_B_c_295_n N_A_1598_93#_M1000_g 0.0068596f $X=8.62 $Y=2.375 $X2=0
+ $Y2=0
cc_352 N_RESET_B_c_282_n N_A_1598_93#_M1000_g 0.00903792f $X=8.255 $Y=1.665
+ $X2=0 $Y2=0
cc_353 N_RESET_B_c_284_n N_A_1598_93#_M1000_g 0.00140024f $X=8.4 $Y=1.665 $X2=0
+ $Y2=0
cc_354 N_RESET_B_c_285_n N_A_1598_93#_M1000_g 0.00248623f $X=8.4 $Y=1.665 $X2=0
+ $Y2=0
cc_355 N_RESET_B_c_289_n N_A_1598_93#_M1000_g 0.0174849f $X=8.545 $Y=1.63 $X2=0
+ $Y2=0
cc_356 N_RESET_B_c_295_n N_A_1598_93#_c_1141_n 0.0255241f $X=8.62 $Y=2.375 $X2=0
+ $Y2=0
cc_357 N_RESET_B_c_296_n N_A_1598_93#_c_1141_n 0.0102544f $X=8.62 $Y=2.465 $X2=0
+ $Y2=0
cc_358 N_RESET_B_c_285_n N_A_1598_93#_c_1141_n 2.32727e-19 $X=8.4 $Y=1.665 $X2=0
+ $Y2=0
cc_359 N_RESET_B_c_295_n N_A_1598_93#_c_1142_n 0.0179198f $X=8.62 $Y=2.375 $X2=0
+ $Y2=0
cc_360 N_RESET_B_c_282_n N_A_1598_93#_c_1142_n 0.00534563f $X=8.255 $Y=1.665
+ $X2=0 $Y2=0
cc_361 N_RESET_B_c_284_n N_A_1598_93#_c_1142_n 0.00307024f $X=8.4 $Y=1.665 $X2=0
+ $Y2=0
cc_362 N_RESET_B_c_285_n N_A_1598_93#_c_1142_n 0.0292669f $X=8.4 $Y=1.665 $X2=0
+ $Y2=0
cc_363 N_RESET_B_c_289_n N_A_1598_93#_c_1142_n 0.00342754f $X=8.545 $Y=1.63
+ $X2=0 $Y2=0
cc_364 N_RESET_B_c_295_n N_A_1598_93#_c_1143_n 0.00121111f $X=8.62 $Y=2.375
+ $X2=0 $Y2=0
cc_365 N_RESET_B_c_296_n N_A_1598_93#_c_1143_n 0.0107743f $X=8.62 $Y=2.465 $X2=0
+ $Y2=0
cc_366 N_RESET_B_c_295_n N_A_1598_93#_c_1138_n 2.15799e-19 $X=8.62 $Y=2.375
+ $X2=0 $Y2=0
cc_367 N_RESET_B_c_289_n N_A_1598_93#_c_1138_n 0.00106075f $X=8.545 $Y=1.63
+ $X2=0 $Y2=0
cc_368 N_RESET_B_c_295_n N_A_1598_93#_c_1146_n 0.00567658f $X=8.62 $Y=2.375
+ $X2=0 $Y2=0
cc_369 N_RESET_B_c_285_n N_A_1598_93#_c_1146_n 0.00239474f $X=8.4 $Y=1.665 $X2=0
+ $Y2=0
cc_370 N_RESET_B_M1012_g N_A_1598_93#_c_1139_n 0.00117144f $X=8.605 $Y=0.805
+ $X2=0 $Y2=0
cc_371 N_RESET_B_M1012_g N_A_1266_119#_c_1226_n 0.0535388f $X=8.605 $Y=0.805
+ $X2=0 $Y2=0
cc_372 N_RESET_B_c_295_n N_A_1266_119#_c_1227_n 0.0166298f $X=8.62 $Y=2.375
+ $X2=0 $Y2=0
cc_373 N_RESET_B_c_296_n N_A_1266_119#_c_1237_n 0.0166298f $X=8.62 $Y=2.465
+ $X2=0 $Y2=0
cc_374 N_RESET_B_c_296_n N_A_1266_119#_c_1238_n 0.00943438f $X=8.62 $Y=2.465
+ $X2=0 $Y2=0
cc_375 N_RESET_B_c_282_n N_A_1266_119#_c_1232_n 0.0247374f $X=8.255 $Y=1.665
+ $X2=0 $Y2=0
cc_376 N_RESET_B_c_284_n N_A_1266_119#_c_1232_n 0.00232289f $X=8.4 $Y=1.665
+ $X2=0 $Y2=0
cc_377 N_RESET_B_c_285_n N_A_1266_119#_c_1232_n 0.0115131f $X=8.4 $Y=1.665 $X2=0
+ $Y2=0
cc_378 N_RESET_B_M1012_g N_A_1266_119#_c_1233_n 0.0144298f $X=8.605 $Y=0.805
+ $X2=0 $Y2=0
cc_379 N_RESET_B_c_282_n N_A_1266_119#_c_1233_n 0.0108617f $X=8.255 $Y=1.665
+ $X2=0 $Y2=0
cc_380 N_RESET_B_c_284_n N_A_1266_119#_c_1233_n 0.0025054f $X=8.4 $Y=1.665 $X2=0
+ $Y2=0
cc_381 N_RESET_B_c_285_n N_A_1266_119#_c_1233_n 0.0302597f $X=8.4 $Y=1.665 $X2=0
+ $Y2=0
cc_382 N_RESET_B_c_289_n N_A_1266_119#_c_1233_n 0.0041539f $X=8.545 $Y=1.63
+ $X2=0 $Y2=0
cc_383 N_RESET_B_M1012_g N_A_1266_119#_c_1234_n 0.00109666f $X=8.605 $Y=0.805
+ $X2=0 $Y2=0
cc_384 N_RESET_B_c_284_n N_A_1266_119#_c_1234_n 0.00111187f $X=8.4 $Y=1.665
+ $X2=0 $Y2=0
cc_385 N_RESET_B_c_285_n N_A_1266_119#_c_1234_n 0.0199249f $X=8.4 $Y=1.665 $X2=0
+ $Y2=0
cc_386 N_RESET_B_c_289_n N_A_1266_119#_c_1234_n 4.14158e-19 $X=8.545 $Y=1.63
+ $X2=0 $Y2=0
cc_387 N_RESET_B_c_285_n N_A_1266_119#_c_1235_n 0.0011399f $X=8.4 $Y=1.665 $X2=0
+ $Y2=0
cc_388 N_RESET_B_c_289_n N_A_1266_119#_c_1235_n 0.0207482f $X=8.545 $Y=1.63
+ $X2=0 $Y2=0
cc_389 N_RESET_B_c_292_n N_VPWR_c_1426_n 5.0378e-19 $X=0.95 $Y=2.465 $X2=0 $Y2=0
cc_390 N_RESET_B_c_292_n N_VPWR_c_1427_n 0.00350285f $X=0.95 $Y=2.465 $X2=0
+ $Y2=0
cc_391 N_RESET_B_c_294_n N_VPWR_c_1429_n 0.00569538f $X=4.91 $Y=2.465 $X2=0
+ $Y2=0
cc_392 N_RESET_B_c_294_n N_VPWR_c_1430_n 0.00445602f $X=4.91 $Y=2.465 $X2=0
+ $Y2=0
cc_393 N_RESET_B_c_293_n N_VPWR_c_1431_n 4.0961e-19 $X=4.91 $Y=2.375 $X2=0 $Y2=0
cc_394 N_RESET_B_c_294_n N_VPWR_c_1431_n 0.00389322f $X=4.91 $Y=2.465 $X2=0
+ $Y2=0
cc_395 N_RESET_B_c_296_n N_VPWR_c_1432_n 0.00722976f $X=8.62 $Y=2.465 $X2=0
+ $Y2=0
cc_396 N_RESET_B_c_292_n N_VPWR_c_1439_n 0.00445602f $X=0.95 $Y=2.465 $X2=0
+ $Y2=0
cc_397 N_RESET_B_c_296_n N_VPWR_c_1442_n 0.00445602f $X=8.62 $Y=2.465 $X2=0
+ $Y2=0
cc_398 N_RESET_B_c_292_n N_VPWR_c_1424_n 0.00895384f $X=0.95 $Y=2.465 $X2=0
+ $Y2=0
cc_399 N_RESET_B_c_294_n N_VPWR_c_1424_n 0.00900367f $X=4.91 $Y=2.465 $X2=0
+ $Y2=0
cc_400 N_RESET_B_c_296_n N_VPWR_c_1424_n 0.00896557f $X=8.62 $Y=2.465 $X2=0
+ $Y2=0
cc_401 N_RESET_B_M1024_g N_A_33_74#_c_1558_n 0.0120626f $X=0.915 $Y=0.58 $X2=0
+ $Y2=0
cc_402 N_RESET_B_c_291_n N_A_33_74#_c_1558_n 0.00946659f $X=0.95 $Y=2.375 $X2=0
+ $Y2=0
cc_403 N_RESET_B_c_281_n N_A_33_74#_c_1558_n 0.00111707f $X=1.345 $Y=1.665 $X2=0
+ $Y2=0
cc_404 N_RESET_B_c_286_n N_A_33_74#_c_1558_n 0.00280068f $X=0.975 $Y=1.515 $X2=0
+ $Y2=0
cc_405 N_RESET_B_c_290_n N_A_33_74#_c_1558_n 0.0317714f $X=1.2 $Y=1.665 $X2=0
+ $Y2=0
cc_406 N_RESET_B_c_291_n N_A_33_74#_c_1564_n 4.6202e-19 $X=0.95 $Y=2.375 $X2=0
+ $Y2=0
cc_407 N_RESET_B_c_292_n N_A_33_74#_c_1564_n 0.0098481f $X=0.95 $Y=2.465 $X2=0
+ $Y2=0
cc_408 N_RESET_B_c_280_n N_A_33_74#_c_1565_n 0.0109181f $X=4.895 $Y=1.665 $X2=0
+ $Y2=0
cc_409 N_RESET_B_c_281_n N_A_33_74#_c_1565_n 0.00321192f $X=1.345 $Y=1.665 $X2=0
+ $Y2=0
cc_410 N_RESET_B_c_290_n N_A_33_74#_c_1565_n 0.00106938f $X=1.2 $Y=1.665 $X2=0
+ $Y2=0
cc_411 N_RESET_B_c_291_n N_A_33_74#_c_1566_n 0.0155155f $X=0.95 $Y=2.375 $X2=0
+ $Y2=0
cc_412 N_RESET_B_c_281_n N_A_33_74#_c_1566_n 0.00427024f $X=1.345 $Y=1.665 $X2=0
+ $Y2=0
cc_413 N_RESET_B_c_286_n N_A_33_74#_c_1566_n 0.00216774f $X=0.975 $Y=1.515 $X2=0
+ $Y2=0
cc_414 N_RESET_B_c_290_n N_A_33_74#_c_1566_n 0.0120416f $X=1.2 $Y=1.665 $X2=0
+ $Y2=0
cc_415 N_RESET_B_c_280_n N_A_33_74#_c_1559_n 0.0232185f $X=4.895 $Y=1.665 $X2=0
+ $Y2=0
cc_416 N_RESET_B_c_280_n N_A_33_74#_c_1568_n 0.00625408f $X=4.895 $Y=1.665 $X2=0
+ $Y2=0
cc_417 N_RESET_B_M1024_g N_A_33_74#_c_1561_n 0.00390091f $X=0.915 $Y=0.58 $X2=0
+ $Y2=0
cc_418 N_RESET_B_M1024_g N_VGND_c_1703_n 0.00554804f $X=0.915 $Y=0.58 $X2=0
+ $Y2=0
cc_419 N_RESET_B_c_286_n N_VGND_c_1703_n 0.00170814f $X=0.975 $Y=1.515 $X2=0
+ $Y2=0
cc_420 N_RESET_B_c_290_n N_VGND_c_1703_n 0.00881738f $X=1.2 $Y=1.665 $X2=0 $Y2=0
cc_421 N_RESET_B_M1015_g N_VGND_c_1705_n 0.00323567f $X=4.895 $Y=0.845 $X2=0
+ $Y2=0
cc_422 N_RESET_B_M1012_g N_VGND_c_1706_n 0.0103576f $X=8.605 $Y=0.805 $X2=0
+ $Y2=0
cc_423 N_RESET_B_M1024_g N_VGND_c_1708_n 0.00461464f $X=0.915 $Y=0.58 $X2=0
+ $Y2=0
cc_424 N_RESET_B_M1012_g N_VGND_c_1712_n 0.0035863f $X=8.605 $Y=0.805 $X2=0
+ $Y2=0
cc_425 N_RESET_B_M1024_g N_VGND_c_1714_n 0.00908835f $X=0.915 $Y=0.58 $X2=0
+ $Y2=0
cc_426 N_RESET_B_M1015_g N_VGND_c_1714_n 9.53055e-19 $X=4.895 $Y=0.845 $X2=0
+ $Y2=0
cc_427 N_RESET_B_M1012_g N_VGND_c_1714_n 0.00401353f $X=8.605 $Y=0.805 $X2=0
+ $Y2=0
cc_428 N_CLK_N_c_479_n N_A_300_74#_c_931_n 0.00127467f $X=1.455 $Y=1.765 $X2=0
+ $Y2=0
cc_429 N_CLK_N_c_479_n N_A_300_74#_c_939_n 0.0179035f $X=1.455 $Y=1.765 $X2=0
+ $Y2=0
cc_430 CLK_N N_A_300_74#_c_939_n 0.00127888f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_431 N_CLK_N_c_479_n N_A_300_74#_c_956_n 0.0111842f $X=1.455 $Y=1.765 $X2=0
+ $Y2=0
cc_432 CLK_N N_A_300_74#_c_956_n 0.00883408f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_433 N_CLK_N_c_478_n N_A_300_74#_c_942_n 0.00345144f $X=1.425 $Y=1.22 $X2=0
+ $Y2=0
cc_434 N_CLK_N_c_479_n N_A_300_74#_c_942_n 0.00385024f $X=1.455 $Y=1.765 $X2=0
+ $Y2=0
cc_435 CLK_N N_A_300_74#_c_942_n 0.0290384f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_436 N_CLK_N_c_478_n N_A_300_74#_c_944_n 0.010507f $X=1.425 $Y=1.22 $X2=0
+ $Y2=0
cc_437 N_CLK_N_c_479_n N_A_300_74#_c_944_n 0.00128681f $X=1.455 $Y=1.765 $X2=0
+ $Y2=0
cc_438 CLK_N N_A_300_74#_c_944_n 0.0220074f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_439 N_CLK_N_c_479_n N_VPWR_c_1427_n 0.0201177f $X=1.455 $Y=1.765 $X2=0 $Y2=0
cc_440 N_CLK_N_c_479_n N_VPWR_c_1428_n 0.0109122f $X=1.455 $Y=1.765 $X2=0 $Y2=0
cc_441 N_CLK_N_c_479_n N_VPWR_c_1440_n 0.00429299f $X=1.455 $Y=1.765 $X2=0 $Y2=0
cc_442 N_CLK_N_c_479_n N_VPWR_c_1424_n 0.00435647f $X=1.455 $Y=1.765 $X2=0 $Y2=0
cc_443 N_CLK_N_c_479_n N_A_33_74#_c_1564_n 7.91415e-19 $X=1.455 $Y=1.765 $X2=0
+ $Y2=0
cc_444 N_CLK_N_c_479_n N_A_33_74#_c_1565_n 0.0153107f $X=1.455 $Y=1.765 $X2=0
+ $Y2=0
cc_445 N_CLK_N_c_479_n N_A_33_74#_c_1566_n 0.00386276f $X=1.455 $Y=1.765 $X2=0
+ $Y2=0
cc_446 N_CLK_N_c_478_n N_VGND_c_1703_n 0.00334184f $X=1.425 $Y=1.22 $X2=0 $Y2=0
cc_447 N_CLK_N_c_478_n N_VGND_c_1704_n 0.00301319f $X=1.425 $Y=1.22 $X2=0 $Y2=0
cc_448 N_CLK_N_c_478_n N_VGND_c_1709_n 0.00433139f $X=1.425 $Y=1.22 $X2=0 $Y2=0
cc_449 N_CLK_N_c_478_n N_VGND_c_1714_n 0.00822407f $X=1.425 $Y=1.22 $X2=0 $Y2=0
cc_450 N_A_507_368#_c_535_n N_A_856_304#_c_721_n 0.021338f $X=3.92 $Y=2.015
+ $X2=0 $Y2=0
cc_451 N_A_507_368#_c_542_n N_A_856_304#_c_721_n 9.74447e-19 $X=3.55 $Y=1.94
+ $X2=0 $Y2=0
cc_452 N_A_507_368#_c_536_n N_A_856_304#_c_722_n 0.011728f $X=4.01 $Y=2.375
+ $X2=0 $Y2=0
cc_453 N_A_507_368#_c_537_n N_A_856_304#_c_722_n 0.0306548f $X=4.01 $Y=2.465
+ $X2=0 $Y2=0
cc_454 N_A_507_368#_c_523_n N_A_856_304#_M1026_g 0.00605388f $X=4.38 $Y=0.79
+ $X2=0 $Y2=0
cc_455 N_A_507_368#_c_551_n N_A_856_304#_M1026_g 0.00705941f $X=5.525 $Y=0.875
+ $X2=0 $Y2=0
cc_456 N_A_507_368#_c_563_p N_A_856_304#_M1026_g 0.00110234f $X=4.465 $Y=0.875
+ $X2=0 $Y2=0
cc_457 N_A_507_368#_c_551_n N_A_856_304#_c_714_n 0.072849f $X=5.525 $Y=0.875
+ $X2=0 $Y2=0
cc_458 N_A_507_368#_c_551_n N_A_856_304#_c_715_n 0.0110644f $X=5.525 $Y=0.875
+ $X2=0 $Y2=0
cc_459 N_A_507_368#_c_563_p N_A_856_304#_c_715_n 0.00128608f $X=4.465 $Y=0.875
+ $X2=0 $Y2=0
cc_460 N_A_507_368#_c_525_n N_A_856_304#_c_716_n 0.0206843f $X=6.365 $Y=0.34
+ $X2=0 $Y2=0
cc_461 N_A_507_368#_c_539_n N_A_856_304#_c_723_n 9.21729e-19 $X=6.81 $Y=1.885
+ $X2=0 $Y2=0
cc_462 N_A_507_368#_c_563_p N_A_856_304#_c_717_n 0.00382995f $X=4.465 $Y=0.875
+ $X2=0 $Y2=0
cc_463 N_A_507_368#_c_542_n N_A_856_304#_c_718_n 0.00112285f $X=3.55 $Y=1.94
+ $X2=0 $Y2=0
cc_464 N_A_507_368#_c_563_p N_A_856_304#_c_718_n 7.16239e-19 $X=4.465 $Y=0.875
+ $X2=0 $Y2=0
cc_465 N_A_507_368#_c_539_n N_A_856_304#_c_720_n 0.00175018f $X=6.81 $Y=1.885
+ $X2=0 $Y2=0
cc_466 N_A_507_368#_c_521_n N_A_714_127#_M1013_d 0.00383506f $X=3.62 $Y=1.245
+ $X2=-0.19 $Y2=-0.245
cc_467 N_A_507_368#_c_524_n N_A_714_127#_M1019_g 0.00745398f $X=5.61 $Y=0.79
+ $X2=0 $Y2=0
cc_468 N_A_507_368#_c_525_n N_A_714_127#_M1019_g 0.00330666f $X=6.365 $Y=0.34
+ $X2=0 $Y2=0
cc_469 N_A_507_368#_c_514_n N_A_714_127#_c_815_n 0.00127496f $X=3.495 $Y=0.525
+ $X2=0 $Y2=0
cc_470 N_A_507_368#_c_521_n N_A_714_127#_c_815_n 0.0329256f $X=3.62 $Y=1.245
+ $X2=0 $Y2=0
cc_471 N_A_507_368#_c_522_n N_A_714_127#_c_815_n 0.0171416f $X=4.295 $Y=0.36
+ $X2=0 $Y2=0
cc_472 N_A_507_368#_c_514_n N_A_714_127#_c_816_n 2.00396e-19 $X=3.495 $Y=0.525
+ $X2=0 $Y2=0
cc_473 N_A_507_368#_c_535_n N_A_714_127#_c_816_n 0.00696166f $X=3.92 $Y=2.015
+ $X2=0 $Y2=0
cc_474 N_A_507_368#_c_520_n N_A_714_127#_c_816_n 0.0130477f $X=3.535 $Y=1.33
+ $X2=0 $Y2=0
cc_475 N_A_507_368#_c_541_n N_A_714_127#_c_816_n 0.0191101f $X=3.55 $Y=1.94
+ $X2=0 $Y2=0
cc_476 N_A_507_368#_c_542_n N_A_714_127#_c_816_n 5.90768e-19 $X=3.55 $Y=1.94
+ $X2=0 $Y2=0
cc_477 N_A_507_368#_c_521_n N_A_714_127#_c_816_n 0.0117841f $X=3.62 $Y=1.245
+ $X2=0 $Y2=0
cc_478 N_A_507_368#_c_536_n N_A_714_127#_c_822_n 0.00667108f $X=4.01 $Y=2.375
+ $X2=0 $Y2=0
cc_479 N_A_507_368#_c_537_n N_A_714_127#_c_822_n 0.00514831f $X=4.01 $Y=2.465
+ $X2=0 $Y2=0
cc_480 N_A_507_368#_c_535_n N_A_714_127#_c_823_n 0.00168553f $X=3.92 $Y=2.015
+ $X2=0 $Y2=0
cc_481 N_A_507_368#_c_536_n N_A_714_127#_c_823_n 0.00296904f $X=4.01 $Y=2.375
+ $X2=0 $Y2=0
cc_482 N_A_507_368#_c_537_n N_A_714_127#_c_827_n 0.0123127f $X=4.01 $Y=2.465
+ $X2=0 $Y2=0
cc_483 N_A_507_368#_c_541_n N_A_714_127#_c_827_n 0.00390957f $X=3.55 $Y=1.94
+ $X2=0 $Y2=0
cc_484 N_A_507_368#_c_542_n N_A_714_127#_c_827_n 0.00649417f $X=3.55 $Y=1.94
+ $X2=0 $Y2=0
cc_485 N_A_507_368#_c_535_n N_A_714_127#_c_828_n 0.00328163f $X=3.92 $Y=2.015
+ $X2=0 $Y2=0
cc_486 N_A_507_368#_c_536_n N_A_714_127#_c_828_n 0.00229797f $X=4.01 $Y=2.375
+ $X2=0 $Y2=0
cc_487 N_A_507_368#_c_541_n N_A_714_127#_c_828_n 0.00711067f $X=3.55 $Y=1.94
+ $X2=0 $Y2=0
cc_488 N_A_507_368#_c_519_n N_A_300_74#_c_947_n 0.00325649f $X=2.807 $Y=1.775
+ $X2=0 $Y2=0
cc_489 N_A_507_368#_c_530_n N_A_300_74#_c_931_n 0.00886276f $X=2.76 $Y=1.14
+ $X2=0 $Y2=0
cc_490 N_A_507_368#_c_531_n N_A_300_74#_c_931_n 5.05212e-19 $X=3.54 $Y=0.36
+ $X2=0 $Y2=0
cc_491 N_A_507_368#_c_532_n N_A_300_74#_c_931_n 0.0040039f $X=3.54 $Y=0.36 $X2=0
+ $Y2=0
cc_492 N_A_507_368#_c_519_n N_A_300_74#_c_932_n 0.0163301f $X=2.807 $Y=1.775
+ $X2=0 $Y2=0
cc_493 N_A_507_368#_c_520_n N_A_300_74#_c_932_n 0.00207366f $X=3.535 $Y=1.33
+ $X2=0 $Y2=0
cc_494 N_A_507_368#_c_530_n N_A_300_74#_c_932_n 0.00654739f $X=2.76 $Y=1.14
+ $X2=0 $Y2=0
cc_495 N_A_507_368#_c_519_n N_A_300_74#_c_933_n 0.00702611f $X=2.807 $Y=1.775
+ $X2=0 $Y2=0
cc_496 N_A_507_368#_c_541_n N_A_300_74#_c_933_n 0.017658f $X=3.55 $Y=1.94 $X2=0
+ $Y2=0
cc_497 N_A_507_368#_c_542_n N_A_300_74#_c_933_n 0.018134f $X=3.55 $Y=1.94 $X2=0
+ $Y2=0
cc_498 N_A_507_368#_c_514_n N_A_300_74#_c_934_n 0.0126901f $X=3.495 $Y=0.525
+ $X2=0 $Y2=0
cc_499 N_A_507_368#_c_535_n N_A_300_74#_c_934_n 0.00965271f $X=3.92 $Y=2.015
+ $X2=0 $Y2=0
cc_500 N_A_507_368#_c_520_n N_A_300_74#_c_934_n 0.0203333f $X=3.535 $Y=1.33
+ $X2=0 $Y2=0
cc_501 N_A_507_368#_c_541_n N_A_300_74#_c_934_n 0.00602473f $X=3.55 $Y=1.94
+ $X2=0 $Y2=0
cc_502 N_A_507_368#_c_542_n N_A_300_74#_c_934_n 0.0175066f $X=3.55 $Y=1.94 $X2=0
+ $Y2=0
cc_503 N_A_507_368#_c_521_n N_A_300_74#_c_934_n 0.00192412f $X=3.62 $Y=1.245
+ $X2=0 $Y2=0
cc_504 N_A_507_368#_c_522_n N_A_300_74#_c_934_n 0.00209574f $X=4.295 $Y=0.36
+ $X2=0 $Y2=0
cc_505 N_A_507_368#_c_536_n N_A_300_74#_c_949_n 0.00718348f $X=4.01 $Y=2.375
+ $X2=0 $Y2=0
cc_506 N_A_507_368#_c_541_n N_A_300_74#_c_949_n 0.00364965f $X=3.55 $Y=1.94
+ $X2=0 $Y2=0
cc_507 N_A_507_368#_c_542_n N_A_300_74#_c_949_n 0.0178863f $X=3.55 $Y=1.94 $X2=0
+ $Y2=0
cc_508 N_A_507_368#_c_537_n N_A_300_74#_c_951_n 0.0101748f $X=4.01 $Y=2.465
+ $X2=0 $Y2=0
cc_509 N_A_507_368#_c_514_n N_A_300_74#_M1030_g 0.0068834f $X=3.495 $Y=0.525
+ $X2=0 $Y2=0
cc_510 N_A_507_368#_c_521_n N_A_300_74#_M1030_g 0.00180495f $X=3.62 $Y=1.245
+ $X2=0 $Y2=0
cc_511 N_A_507_368#_c_522_n N_A_300_74#_M1030_g 0.0173102f $X=4.295 $Y=0.36
+ $X2=0 $Y2=0
cc_512 N_A_507_368#_c_523_n N_A_300_74#_M1030_g 0.00309568f $X=4.38 $Y=0.79
+ $X2=0 $Y2=0
cc_513 N_A_507_368#_c_522_n N_A_300_74#_c_936_n 0.004367f $X=4.295 $Y=0.36 $X2=0
+ $Y2=0
cc_514 N_A_507_368#_c_551_n N_A_300_74#_c_936_n 0.00973035f $X=5.525 $Y=0.875
+ $X2=0 $Y2=0
cc_515 N_A_507_368#_c_525_n N_A_300_74#_c_936_n 0.00676815f $X=6.365 $Y=0.34
+ $X2=0 $Y2=0
cc_516 N_A_507_368#_c_526_n N_A_300_74#_c_936_n 0.0041995f $X=5.695 $Y=0.34
+ $X2=0 $Y2=0
cc_517 N_A_507_368#_c_514_n N_A_300_74#_c_937_n 0.0100071f $X=3.495 $Y=0.525
+ $X2=0 $Y2=0
cc_518 N_A_507_368#_c_516_n N_A_300_74#_M1005_g 0.00954257f $X=6.9 $Y=1.29 $X2=0
+ $Y2=0
cc_519 N_A_507_368#_c_524_n N_A_300_74#_M1005_g 8.97611e-19 $X=5.61 $Y=0.79
+ $X2=0 $Y2=0
cc_520 N_A_507_368#_c_525_n N_A_300_74#_M1005_g 0.0169375f $X=6.365 $Y=0.34
+ $X2=0 $Y2=0
cc_521 N_A_507_368#_c_527_n N_A_300_74#_M1005_g 0.0152469f $X=6.45 $Y=1.125
+ $X2=0 $Y2=0
cc_522 N_A_507_368#_c_554_n N_A_300_74#_M1005_g 8.5704e-19 $X=7.08 $Y=1.29 $X2=0
+ $Y2=0
cc_523 N_A_507_368#_c_539_n N_A_300_74#_c_952_n 0.00540267f $X=6.81 $Y=1.885
+ $X2=0 $Y2=0
cc_524 N_A_507_368#_c_519_n N_A_300_74#_c_940_n 0.00175358f $X=2.807 $Y=1.775
+ $X2=0 $Y2=0
cc_525 N_A_507_368#_c_520_n N_A_300_74#_c_941_n 0.00557643f $X=3.535 $Y=1.33
+ $X2=0 $Y2=0
cc_526 N_A_507_368#_c_539_n N_A_300_74#_c_955_n 0.00223241f $X=6.81 $Y=1.885
+ $X2=0 $Y2=0
cc_527 N_A_507_368#_c_515_n N_A_300_74#_c_943_n 0.00883406f $X=6.81 $Y=1.795
+ $X2=0 $Y2=0
cc_528 N_A_507_368#_c_539_n N_A_300_74#_c_943_n 0.00783008f $X=6.81 $Y=1.885
+ $X2=0 $Y2=0
cc_529 N_A_507_368#_c_517_n N_A_300_74#_c_943_n 0.00107089f $X=7.6 $Y=1.2 $X2=0
+ $Y2=0
cc_530 N_A_507_368#_c_553_n N_A_300_74#_c_943_n 8.672e-19 $X=6.535 $Y=1.21 $X2=0
+ $Y2=0
cc_531 N_A_507_368#_c_554_n N_A_300_74#_c_943_n 0.0348735f $X=7.08 $Y=1.29 $X2=0
+ $Y2=0
cc_532 N_A_507_368#_c_528_n N_A_300_74#_c_943_n 0.00717074f $X=7.255 $Y=1.29
+ $X2=0 $Y2=0
cc_533 N_A_507_368#_c_529_n N_A_300_74#_c_943_n 0.00892364f $X=7.255 $Y=1.29
+ $X2=0 $Y2=0
cc_534 N_A_507_368#_c_533_n N_A_300_74#_c_943_n 0.00691585f $X=6.75 $Y=1.29
+ $X2=0 $Y2=0
cc_535 N_A_507_368#_c_534_n N_A_300_74#_c_943_n 6.09268e-19 $X=7.42 $Y=1.29
+ $X2=0 $Y2=0
cc_536 N_A_507_368#_c_539_n N_A_300_74#_c_959_n 0.00250118f $X=6.81 $Y=1.885
+ $X2=0 $Y2=0
cc_537 N_A_507_368#_c_515_n N_A_300_74#_c_960_n 0.00562911f $X=6.81 $Y=1.795
+ $X2=0 $Y2=0
cc_538 N_A_507_368#_c_539_n N_A_300_74#_c_960_n 0.0130552f $X=6.81 $Y=1.885
+ $X2=0 $Y2=0
cc_539 N_A_507_368#_c_517_n N_A_300_74#_c_960_n 0.00873909f $X=7.6 $Y=1.2 $X2=0
+ $Y2=0
cc_540 N_A_507_368#_c_534_n N_A_300_74#_c_960_n 0.00582183f $X=7.42 $Y=1.29
+ $X2=0 $Y2=0
cc_541 N_A_507_368#_c_515_n N_A_300_74#_c_945_n 0.00134609f $X=6.81 $Y=1.795
+ $X2=0 $Y2=0
cc_542 N_A_507_368#_c_553_n N_A_300_74#_c_945_n 0.00994746f $X=6.535 $Y=1.21
+ $X2=0 $Y2=0
cc_543 N_A_507_368#_c_515_n N_A_300_74#_c_946_n 0.0215527f $X=6.81 $Y=1.795
+ $X2=0 $Y2=0
cc_544 N_A_507_368#_c_553_n N_A_300_74#_c_946_n 0.00106755f $X=6.535 $Y=1.21
+ $X2=0 $Y2=0
cc_545 N_A_507_368#_c_518_n N_A_1598_93#_M1000_g 0.0413341f $X=7.675 $Y=1.125
+ $X2=0 $Y2=0
cc_546 N_A_507_368#_c_534_n N_A_1598_93#_M1000_g 0.00246675f $X=7.42 $Y=1.29
+ $X2=0 $Y2=0
cc_547 N_A_507_368#_c_527_n N_A_1266_119#_M1005_d 0.0153989f $X=6.45 $Y=1.125
+ $X2=-0.19 $Y2=-0.245
cc_548 N_A_507_368#_c_553_n N_A_1266_119#_M1005_d 0.00269935f $X=6.535 $Y=1.21
+ $X2=-0.19 $Y2=-0.245
cc_549 N_A_507_368#_c_533_n N_A_1266_119#_M1005_d 0.0025788f $X=6.75 $Y=1.29
+ $X2=-0.19 $Y2=-0.245
cc_550 N_A_507_368#_c_516_n N_A_1266_119#_c_1266_n 0.0198469f $X=6.9 $Y=1.29
+ $X2=0 $Y2=0
cc_551 N_A_507_368#_c_518_n N_A_1266_119#_c_1266_n 0.0148493f $X=7.675 $Y=1.125
+ $X2=0 $Y2=0
cc_552 N_A_507_368#_c_527_n N_A_1266_119#_c_1266_n 0.0266855f $X=6.45 $Y=1.125
+ $X2=0 $Y2=0
cc_553 N_A_507_368#_c_533_n N_A_1266_119#_c_1266_n 0.0553581f $X=6.75 $Y=1.29
+ $X2=0 $Y2=0
cc_554 N_A_507_368#_c_539_n N_A_1266_119#_c_1241_n 0.00416251f $X=6.81 $Y=1.885
+ $X2=0 $Y2=0
cc_555 N_A_507_368#_c_518_n N_A_1266_119#_c_1231_n 0.00779099f $X=7.675 $Y=1.125
+ $X2=0 $Y2=0
cc_556 N_A_507_368#_c_528_n N_A_1266_119#_c_1232_n 0.0080525f $X=7.255 $Y=1.29
+ $X2=0 $Y2=0
cc_557 N_A_507_368#_c_534_n N_A_1266_119#_c_1232_n 6.25344e-19 $X=7.42 $Y=1.29
+ $X2=0 $Y2=0
cc_558 N_A_507_368#_c_517_n N_A_1266_119#_c_1274_n 0.00534427f $X=7.6 $Y=1.2
+ $X2=0 $Y2=0
cc_559 N_A_507_368#_c_528_n N_A_1266_119#_c_1274_n 0.00890259f $X=7.255 $Y=1.29
+ $X2=0 $Y2=0
cc_560 N_A_507_368#_c_537_n N_VPWR_c_1429_n 0.00177436f $X=4.01 $Y=2.465 $X2=0
+ $Y2=0
cc_561 N_A_507_368#_c_539_n N_VPWR_c_1435_n 0.00445972f $X=6.81 $Y=1.885 $X2=0
+ $Y2=0
cc_562 N_A_507_368#_c_537_n N_VPWR_c_1441_n 0.00325612f $X=4.01 $Y=2.465 $X2=0
+ $Y2=0
cc_563 N_A_507_368#_c_537_n N_VPWR_c_1424_n 0.00502377f $X=4.01 $Y=2.465 $X2=0
+ $Y2=0
cc_564 N_A_507_368#_c_539_n N_VPWR_c_1424_n 0.00863862f $X=6.81 $Y=1.885 $X2=0
+ $Y2=0
cc_565 N_A_507_368#_c_519_n N_A_33_74#_c_1559_n 0.0290839f $X=2.807 $Y=1.775
+ $X2=0 $Y2=0
cc_566 N_A_507_368#_c_530_n N_A_33_74#_c_1559_n 0.0572975f $X=2.76 $Y=1.14 $X2=0
+ $Y2=0
cc_567 N_A_507_368#_M1010_d N_A_33_74#_c_1560_n 0.010153f $X=2.55 $Y=0.5 $X2=0
+ $Y2=0
cc_568 N_A_507_368#_c_520_n N_A_33_74#_c_1560_n 0.00683052f $X=3.535 $Y=1.33
+ $X2=0 $Y2=0
cc_569 N_A_507_368#_c_530_n N_A_33_74#_c_1560_n 0.0215648f $X=2.76 $Y=1.14 $X2=0
+ $Y2=0
cc_570 N_A_507_368#_c_531_n N_A_33_74#_c_1560_n 0.00549888f $X=3.54 $Y=0.36
+ $X2=0 $Y2=0
cc_571 N_A_507_368#_c_532_n N_A_33_74#_c_1560_n 0.00192524f $X=3.54 $Y=0.36
+ $X2=0 $Y2=0
cc_572 N_A_507_368#_M1009_d N_A_33_74#_c_1568_n 0.0117553f $X=2.535 $Y=1.84
+ $X2=0 $Y2=0
cc_573 N_A_507_368#_c_519_n N_A_33_74#_c_1568_n 0.0210739f $X=2.807 $Y=1.775
+ $X2=0 $Y2=0
cc_574 N_A_507_368#_c_541_n N_A_33_74#_c_1568_n 0.0306116f $X=3.55 $Y=1.94 $X2=0
+ $Y2=0
cc_575 N_A_507_368#_c_514_n N_A_33_74#_c_1562_n 0.00101545f $X=3.495 $Y=0.525
+ $X2=0 $Y2=0
cc_576 N_A_507_368#_c_520_n N_A_33_74#_c_1562_n 0.0195074f $X=3.535 $Y=1.33
+ $X2=0 $Y2=0
cc_577 N_A_507_368#_c_521_n N_A_33_74#_c_1562_n 0.0156696f $X=3.62 $Y=1.245
+ $X2=0 $Y2=0
cc_578 N_A_507_368#_c_530_n N_A_33_74#_c_1562_n 0.00785713f $X=2.76 $Y=1.14
+ $X2=0 $Y2=0
cc_579 N_A_507_368#_c_531_n N_A_33_74#_c_1562_n 0.0181046f $X=3.54 $Y=0.36 $X2=0
+ $Y2=0
cc_580 N_A_507_368#_c_532_n N_A_33_74#_c_1562_n 0.00611936f $X=3.54 $Y=0.36
+ $X2=0 $Y2=0
cc_581 N_A_507_368#_c_551_n N_VGND_M1015_d 0.0158358f $X=5.525 $Y=0.875 $X2=0
+ $Y2=0
cc_582 N_A_507_368#_c_524_n N_VGND_M1015_d 0.00465623f $X=5.61 $Y=0.79 $X2=0
+ $Y2=0
cc_583 N_A_507_368#_c_532_n N_VGND_c_1704_n 0.0024897f $X=3.54 $Y=0.36 $X2=0
+ $Y2=0
cc_584 N_A_507_368#_c_522_n N_VGND_c_1705_n 0.00810195f $X=4.295 $Y=0.36 $X2=0
+ $Y2=0
cc_585 N_A_507_368#_c_523_n N_VGND_c_1705_n 0.00489725f $X=4.38 $Y=0.79 $X2=0
+ $Y2=0
cc_586 N_A_507_368#_c_551_n N_VGND_c_1705_n 0.0260579f $X=5.525 $Y=0.875 $X2=0
+ $Y2=0
cc_587 N_A_507_368#_c_524_n N_VGND_c_1705_n 0.0153511f $X=5.61 $Y=0.79 $X2=0
+ $Y2=0
cc_588 N_A_507_368#_c_526_n N_VGND_c_1705_n 0.0150385f $X=5.695 $Y=0.34 $X2=0
+ $Y2=0
cc_589 N_A_507_368#_c_518_n N_VGND_c_1706_n 0.00102171f $X=7.675 $Y=1.125 $X2=0
+ $Y2=0
cc_590 N_A_507_368#_c_522_n N_VGND_c_1710_n 0.0496784f $X=4.295 $Y=0.36 $X2=0
+ $Y2=0
cc_591 N_A_507_368#_c_531_n N_VGND_c_1710_n 0.0427221f $X=3.54 $Y=0.36 $X2=0
+ $Y2=0
cc_592 N_A_507_368#_c_532_n N_VGND_c_1710_n 0.012631f $X=3.54 $Y=0.36 $X2=0
+ $Y2=0
cc_593 N_A_507_368#_c_518_n N_VGND_c_1711_n 0.00332223f $X=7.675 $Y=1.125 $X2=0
+ $Y2=0
cc_594 N_A_507_368#_c_525_n N_VGND_c_1711_n 0.0548435f $X=6.365 $Y=0.34 $X2=0
+ $Y2=0
cc_595 N_A_507_368#_c_526_n N_VGND_c_1711_n 0.0116199f $X=5.695 $Y=0.34 $X2=0
+ $Y2=0
cc_596 N_A_507_368#_c_514_n N_VGND_c_1714_n 0.00735925f $X=3.495 $Y=0.525 $X2=0
+ $Y2=0
cc_597 N_A_507_368#_c_518_n N_VGND_c_1714_n 0.00477801f $X=7.675 $Y=1.125 $X2=0
+ $Y2=0
cc_598 N_A_507_368#_c_522_n N_VGND_c_1714_n 0.0272206f $X=4.295 $Y=0.36 $X2=0
+ $Y2=0
cc_599 N_A_507_368#_c_551_n N_VGND_c_1714_n 0.0237285f $X=5.525 $Y=0.875 $X2=0
+ $Y2=0
cc_600 N_A_507_368#_c_525_n N_VGND_c_1714_n 0.0291469f $X=6.365 $Y=0.34 $X2=0
+ $Y2=0
cc_601 N_A_507_368#_c_526_n N_VGND_c_1714_n 0.00583764f $X=5.695 $Y=0.34 $X2=0
+ $Y2=0
cc_602 N_A_507_368#_c_531_n N_VGND_c_1714_n 0.0224006f $X=3.54 $Y=0.36 $X2=0
+ $Y2=0
cc_603 N_A_507_368#_c_532_n N_VGND_c_1714_n 0.00994116f $X=3.54 $Y=0.36 $X2=0
+ $Y2=0
cc_604 N_A_507_368#_c_563_p A_850_127# 0.00165194f $X=4.465 $Y=0.875 $X2=-0.19
+ $Y2=-0.245
cc_605 N_A_507_368#_c_551_n A_922_127# 0.00179164f $X=5.525 $Y=0.875 $X2=-0.19
+ $Y2=-0.245
cc_606 N_A_856_304#_c_714_n N_A_714_127#_M1019_g 0.013473f $X=5.865 $Y=1.215
+ $X2=0 $Y2=0
cc_607 N_A_856_304#_c_716_n N_A_714_127#_M1019_g 0.011387f $X=6.03 $Y=0.76 $X2=0
+ $Y2=0
cc_608 N_A_856_304#_c_745_n N_A_714_127#_M1019_g 3.84191e-19 $X=6.03 $Y=1.215
+ $X2=0 $Y2=0
cc_609 N_A_856_304#_c_720_n N_A_714_127#_M1019_g 0.00824116f $X=6.282 $Y=1.97
+ $X2=0 $Y2=0
cc_610 N_A_856_304#_c_723_n N_A_714_127#_c_813_n 4.6813e-19 $X=6.11 $Y=2.815
+ $X2=0 $Y2=0
cc_611 N_A_856_304#_c_746_n N_A_714_127#_c_813_n 0.00710477f $X=6.11 $Y=2.135
+ $X2=0 $Y2=0
cc_612 N_A_856_304#_c_720_n N_A_714_127#_c_813_n 0.0157335f $X=6.282 $Y=1.97
+ $X2=0 $Y2=0
cc_613 N_A_856_304#_c_714_n N_A_714_127#_c_814_n 0.00228823f $X=5.865 $Y=1.215
+ $X2=0 $Y2=0
cc_614 N_A_856_304#_M1026_g N_A_714_127#_c_815_n 2.5148e-19 $X=4.535 $Y=0.845
+ $X2=0 $Y2=0
cc_615 N_A_856_304#_c_721_n N_A_714_127#_c_816_n 0.00221106f $X=4.4 $Y=2.375
+ $X2=0 $Y2=0
cc_616 N_A_856_304#_M1026_g N_A_714_127#_c_816_n 0.00103829f $X=4.535 $Y=0.845
+ $X2=0 $Y2=0
cc_617 N_A_856_304#_c_715_n N_A_714_127#_c_816_n 0.00755217f $X=4.61 $Y=1.215
+ $X2=0 $Y2=0
cc_618 N_A_856_304#_c_717_n N_A_714_127#_c_816_n 0.0186696f $X=4.445 $Y=1.685
+ $X2=0 $Y2=0
cc_619 N_A_856_304#_c_718_n N_A_714_127#_c_816_n 0.00494708f $X=4.445 $Y=1.685
+ $X2=0 $Y2=0
cc_620 N_A_856_304#_c_719_n N_A_714_127#_c_816_n 0.00936947f $X=4.445 $Y=1.52
+ $X2=0 $Y2=0
cc_621 N_A_856_304#_c_721_n N_A_714_127#_c_822_n 0.00167493f $X=4.4 $Y=2.375
+ $X2=0 $Y2=0
cc_622 N_A_856_304#_c_722_n N_A_714_127#_c_822_n 3.29789e-19 $X=4.4 $Y=2.465
+ $X2=0 $Y2=0
cc_623 N_A_856_304#_c_721_n N_A_714_127#_c_823_n 0.0162018f $X=4.4 $Y=2.375
+ $X2=0 $Y2=0
cc_624 N_A_856_304#_c_717_n N_A_714_127#_c_823_n 0.0232433f $X=4.445 $Y=1.685
+ $X2=0 $Y2=0
cc_625 N_A_856_304#_c_718_n N_A_714_127#_c_823_n 0.00103212f $X=4.445 $Y=1.685
+ $X2=0 $Y2=0
cc_626 N_A_856_304#_c_721_n N_A_714_127#_c_824_n 0.00127637f $X=4.4 $Y=2.375
+ $X2=0 $Y2=0
cc_627 N_A_856_304#_c_722_n N_A_714_127#_c_824_n 3.90246e-19 $X=4.4 $Y=2.465
+ $X2=0 $Y2=0
cc_628 N_A_856_304#_c_746_n N_A_714_127#_c_825_n 0.0103534f $X=6.11 $Y=2.135
+ $X2=0 $Y2=0
cc_629 N_A_856_304#_c_714_n N_A_714_127#_c_817_n 0.0234898f $X=5.865 $Y=1.215
+ $X2=0 $Y2=0
cc_630 N_A_856_304#_c_720_n N_A_714_127#_c_817_n 0.0399258f $X=6.282 $Y=1.97
+ $X2=0 $Y2=0
cc_631 N_A_856_304#_c_722_n N_A_714_127#_c_827_n 0.00152047f $X=4.4 $Y=2.465
+ $X2=0 $Y2=0
cc_632 N_A_856_304#_M1026_g N_A_714_127#_c_818_n 5.79331e-19 $X=4.535 $Y=0.845
+ $X2=0 $Y2=0
cc_633 N_A_856_304#_M1026_g N_A_300_74#_c_934_n 0.00462129f $X=4.535 $Y=0.845
+ $X2=0 $Y2=0
cc_634 N_A_856_304#_c_715_n N_A_300_74#_c_934_n 0.00147567f $X=4.61 $Y=1.215
+ $X2=0 $Y2=0
cc_635 N_A_856_304#_c_718_n N_A_300_74#_c_934_n 9.12797e-19 $X=4.445 $Y=1.685
+ $X2=0 $Y2=0
cc_636 N_A_856_304#_c_719_n N_A_300_74#_c_934_n 7.03563e-19 $X=4.445 $Y=1.52
+ $X2=0 $Y2=0
cc_637 N_A_856_304#_M1026_g N_A_300_74#_M1030_g 0.0464456f $X=4.535 $Y=0.845
+ $X2=0 $Y2=0
cc_638 N_A_856_304#_M1026_g N_A_300_74#_c_936_n 0.00815681f $X=4.535 $Y=0.845
+ $X2=0 $Y2=0
cc_639 N_A_856_304#_c_716_n N_A_300_74#_M1005_g 0.00547135f $X=6.03 $Y=0.76
+ $X2=0 $Y2=0
cc_640 N_A_856_304#_c_745_n N_A_300_74#_M1005_g 0.00198105f $X=6.03 $Y=1.215
+ $X2=0 $Y2=0
cc_641 N_A_856_304#_c_720_n N_A_300_74#_M1005_g 0.00421803f $X=6.282 $Y=1.97
+ $X2=0 $Y2=0
cc_642 N_A_856_304#_c_746_n N_A_300_74#_c_943_n 0.013462f $X=6.11 $Y=2.135 $X2=0
+ $Y2=0
cc_643 N_A_856_304#_c_746_n N_A_300_74#_c_945_n 0.0229541f $X=6.11 $Y=2.135
+ $X2=0 $Y2=0
cc_644 N_A_856_304#_c_720_n N_A_300_74#_c_945_n 0.0236964f $X=6.282 $Y=1.97
+ $X2=0 $Y2=0
cc_645 N_A_856_304#_c_746_n N_A_300_74#_c_946_n 0.00343033f $X=6.11 $Y=2.135
+ $X2=0 $Y2=0
cc_646 N_A_856_304#_c_722_n N_VPWR_c_1429_n 0.011809f $X=4.4 $Y=2.465 $X2=0
+ $Y2=0
cc_647 N_A_856_304#_c_723_n N_VPWR_c_1431_n 0.0241513f $X=6.11 $Y=2.815 $X2=0
+ $Y2=0
cc_648 N_A_856_304#_c_723_n N_VPWR_c_1435_n 0.0315916f $X=6.11 $Y=2.815 $X2=0
+ $Y2=0
cc_649 N_A_856_304#_c_722_n N_VPWR_c_1441_n 0.00413917f $X=4.4 $Y=2.465 $X2=0
+ $Y2=0
cc_650 N_A_856_304#_c_722_n N_VPWR_c_1424_n 0.00855067f $X=4.4 $Y=2.465 $X2=0
+ $Y2=0
cc_651 N_A_856_304#_c_723_n N_VPWR_c_1424_n 0.0261488f $X=6.11 $Y=2.815 $X2=0
+ $Y2=0
cc_652 N_A_856_304#_c_714_n N_VGND_M1015_d 0.00417413f $X=5.865 $Y=1.215 $X2=0
+ $Y2=0
cc_653 N_A_856_304#_M1026_g N_VGND_c_1714_n 9.24014e-19 $X=4.535 $Y=0.845 $X2=0
+ $Y2=0
cc_654 N_A_714_127#_c_816_n N_A_300_74#_c_934_n 0.023636f $X=3.97 $Y=2.02 $X2=0
+ $Y2=0
cc_655 N_A_714_127#_c_818_n N_A_300_74#_c_934_n 0.00240424f $X=4 $Y=1.075 $X2=0
+ $Y2=0
cc_656 N_A_714_127#_c_822_n N_A_300_74#_c_949_n 0.00130581f $X=3.97 $Y=2.52
+ $X2=0 $Y2=0
cc_657 N_A_714_127#_c_827_n N_A_300_74#_c_949_n 4.01822e-19 $X=3.97 $Y=2.75
+ $X2=0 $Y2=0
cc_658 N_A_714_127#_c_822_n N_A_300_74#_c_951_n 4.17088e-19 $X=3.97 $Y=2.52
+ $X2=0 $Y2=0
cc_659 N_A_714_127#_c_827_n N_A_300_74#_c_951_n 0.00615847f $X=3.97 $Y=2.75
+ $X2=0 $Y2=0
cc_660 N_A_714_127#_c_815_n N_A_300_74#_M1030_g 0.00380092f $X=3.96 $Y=0.855
+ $X2=0 $Y2=0
cc_661 N_A_714_127#_c_816_n N_A_300_74#_M1030_g 0.00146855f $X=3.97 $Y=2.02
+ $X2=0 $Y2=0
cc_662 N_A_714_127#_c_818_n N_A_300_74#_M1030_g 0.00289954f $X=4 $Y=1.075 $X2=0
+ $Y2=0
cc_663 N_A_714_127#_M1019_g N_A_300_74#_c_936_n 0.00882199f $X=5.815 $Y=0.965
+ $X2=0 $Y2=0
cc_664 N_A_714_127#_M1019_g N_A_300_74#_M1005_g 0.0106687f $X=5.815 $Y=0.965
+ $X2=0 $Y2=0
cc_665 N_A_714_127#_c_813_n N_A_300_74#_c_945_n 4.20447e-19 $X=5.88 $Y=1.885
+ $X2=0 $Y2=0
cc_666 N_A_714_127#_c_813_n N_A_300_74#_c_946_n 0.0214083f $X=5.88 $Y=1.885
+ $X2=0 $Y2=0
cc_667 N_A_714_127#_c_825_n N_VPWR_M1018_s 0.00509503f $X=5.53 $Y=2.02 $X2=0
+ $Y2=0
cc_668 N_A_714_127#_c_817_n N_VPWR_M1018_s 0.00133386f $X=5.53 $Y=1.635 $X2=0
+ $Y2=0
cc_669 N_A_714_127#_c_823_n N_VPWR_c_1429_n 0.0172889f $X=4.97 $Y=2.105 $X2=0
+ $Y2=0
cc_670 N_A_714_127#_c_824_n N_VPWR_c_1429_n 0.0180054f $X=5.135 $Y=2.75 $X2=0
+ $Y2=0
cc_671 N_A_714_127#_c_827_n N_VPWR_c_1429_n 0.017479f $X=3.97 $Y=2.75 $X2=0
+ $Y2=0
cc_672 N_A_714_127#_c_824_n N_VPWR_c_1430_n 0.0145938f $X=5.135 $Y=2.75 $X2=0
+ $Y2=0
cc_673 N_A_714_127#_c_813_n N_VPWR_c_1431_n 0.0143441f $X=5.88 $Y=1.885 $X2=0
+ $Y2=0
cc_674 N_A_714_127#_c_814_n N_VPWR_c_1431_n 0.00226768f $X=5.74 $Y=1.635 $X2=0
+ $Y2=0
cc_675 N_A_714_127#_c_824_n N_VPWR_c_1431_n 0.0477416f $X=5.135 $Y=2.75 $X2=0
+ $Y2=0
cc_676 N_A_714_127#_c_825_n N_VPWR_c_1431_n 0.0166816f $X=5.53 $Y=2.02 $X2=0
+ $Y2=0
cc_677 N_A_714_127#_c_813_n N_VPWR_c_1435_n 0.00413917f $X=5.88 $Y=1.885 $X2=0
+ $Y2=0
cc_678 N_A_714_127#_c_827_n N_VPWR_c_1441_n 0.0183913f $X=3.97 $Y=2.75 $X2=0
+ $Y2=0
cc_679 N_A_714_127#_c_813_n N_VPWR_c_1424_n 0.00822528f $X=5.88 $Y=1.885 $X2=0
+ $Y2=0
cc_680 N_A_714_127#_c_824_n N_VPWR_c_1424_n 0.0120466f $X=5.135 $Y=2.75 $X2=0
+ $Y2=0
cc_681 N_A_714_127#_c_827_n N_VPWR_c_1424_n 0.0151919f $X=3.97 $Y=2.75 $X2=0
+ $Y2=0
cc_682 N_A_714_127#_c_822_n N_A_33_74#_c_1568_n 0.00642724f $X=3.97 $Y=2.52
+ $X2=0 $Y2=0
cc_683 N_A_714_127#_c_822_n N_A_33_74#_c_1569_n 0.00132593f $X=3.97 $Y=2.52
+ $X2=0 $Y2=0
cc_684 N_A_714_127#_c_827_n N_A_33_74#_c_1569_n 0.0315489f $X=3.97 $Y=2.75 $X2=0
+ $Y2=0
cc_685 N_A_300_74#_c_960_n N_A_1598_93#_M1000_g 0.0139991f $X=7.475 $Y=1.86
+ $X2=0 $Y2=0
cc_686 N_A_300_74#_c_952_n N_A_1598_93#_c_1141_n 0.0275569f $X=7.66 $Y=2.465
+ $X2=0 $Y2=0
cc_687 N_A_300_74#_c_955_n N_A_1598_93#_c_1141_n 0.0185966f $X=7.515 $Y=2.16
+ $X2=0 $Y2=0
cc_688 N_A_300_74#_c_943_n N_A_1266_119#_c_1266_n 0.00277079f $X=7.31 $Y=1.715
+ $X2=0 $Y2=0
cc_689 N_A_300_74#_c_955_n N_A_1266_119#_c_1241_n 9.05598e-19 $X=7.515 $Y=2.16
+ $X2=0 $Y2=0
cc_690 N_A_300_74#_c_959_n N_A_1266_119#_c_1241_n 0.0103637f $X=7.475 $Y=1.86
+ $X2=0 $Y2=0
cc_691 N_A_300_74#_c_952_n N_A_1266_119#_c_1232_n 0.00314472f $X=7.66 $Y=2.465
+ $X2=0 $Y2=0
cc_692 N_A_300_74#_c_955_n N_A_1266_119#_c_1232_n 0.0046061f $X=7.515 $Y=2.16
+ $X2=0 $Y2=0
cc_693 N_A_300_74#_c_943_n N_A_1266_119#_c_1232_n 0.01265f $X=7.31 $Y=1.715
+ $X2=0 $Y2=0
cc_694 N_A_300_74#_c_959_n N_A_1266_119#_c_1232_n 0.0415019f $X=7.475 $Y=1.86
+ $X2=0 $Y2=0
cc_695 N_A_300_74#_c_960_n N_A_1266_119#_c_1232_n 0.0057575f $X=7.475 $Y=1.86
+ $X2=0 $Y2=0
cc_696 N_A_300_74#_c_952_n N_A_1266_119#_c_1243_n 0.0157277f $X=7.66 $Y=2.465
+ $X2=0 $Y2=0
cc_697 N_A_300_74#_c_955_n N_A_1266_119#_c_1243_n 0.00213739f $X=7.515 $Y=2.16
+ $X2=0 $Y2=0
cc_698 N_A_300_74#_c_959_n N_A_1266_119#_c_1243_n 0.010457f $X=7.475 $Y=1.86
+ $X2=0 $Y2=0
cc_699 N_A_300_74#_c_956_n N_VPWR_M1009_s 0.00470783f $X=1.935 $Y=1.982 $X2=0
+ $Y2=0
cc_700 N_A_300_74#_c_947_n N_VPWR_c_1428_n 0.0215013f $X=2.46 $Y=1.765 $X2=0
+ $Y2=0
cc_701 N_A_300_74#_c_952_n N_VPWR_c_1432_n 0.00171173f $X=7.66 $Y=2.465 $X2=0
+ $Y2=0
cc_702 N_A_300_74#_c_952_n N_VPWR_c_1435_n 0.00323148f $X=7.66 $Y=2.465 $X2=0
+ $Y2=0
cc_703 N_A_300_74#_c_947_n N_VPWR_c_1441_n 0.00413917f $X=2.46 $Y=1.765 $X2=0
+ $Y2=0
cc_704 N_A_300_74#_c_951_n N_VPWR_c_1441_n 0.00444483f $X=3.56 $Y=2.465 $X2=0
+ $Y2=0
cc_705 N_A_300_74#_c_947_n N_VPWR_c_1424_n 0.00420259f $X=2.46 $Y=1.765 $X2=0
+ $Y2=0
cc_706 N_A_300_74#_c_949_n N_VPWR_c_1424_n 0.00132957f $X=3.485 $Y=2.39 $X2=0
+ $Y2=0
cc_707 N_A_300_74#_c_951_n N_VPWR_c_1424_n 0.00859578f $X=3.56 $Y=2.465 $X2=0
+ $Y2=0
cc_708 N_A_300_74#_c_952_n N_VPWR_c_1424_n 0.00410412f $X=7.66 $Y=2.465 $X2=0
+ $Y2=0
cc_709 N_A_300_74#_M1017_d N_A_33_74#_c_1565_n 0.00817345f $X=1.53 $Y=1.84 $X2=0
+ $Y2=0
cc_710 N_A_300_74#_c_939_n N_A_33_74#_c_1565_n 0.00352376f $X=2.37 $Y=1.515
+ $X2=0 $Y2=0
cc_711 N_A_300_74#_c_956_n N_A_33_74#_c_1565_n 0.0459311f $X=1.935 $Y=1.982
+ $X2=0 $Y2=0
cc_712 N_A_300_74#_c_947_n N_A_33_74#_c_1559_n 0.0190515f $X=2.46 $Y=1.765 $X2=0
+ $Y2=0
cc_713 N_A_300_74#_c_931_n N_A_33_74#_c_1559_n 0.018377f $X=2.475 $Y=1.35 $X2=0
+ $Y2=0
cc_714 N_A_300_74#_c_933_n N_A_33_74#_c_1559_n 0.00136931f $X=3.07 $Y=2.315
+ $X2=0 $Y2=0
cc_715 N_A_300_74#_c_939_n N_A_33_74#_c_1559_n 0.00654167f $X=2.37 $Y=1.515
+ $X2=0 $Y2=0
cc_716 N_A_300_74#_c_940_n N_A_33_74#_c_1559_n 0.0106567f $X=2.46 $Y=1.557 $X2=0
+ $Y2=0
cc_717 N_A_300_74#_c_956_n N_A_33_74#_c_1559_n 0.0152428f $X=1.935 $Y=1.982
+ $X2=0 $Y2=0
cc_718 N_A_300_74#_c_942_n N_A_33_74#_c_1559_n 0.058464f $X=2.08 $Y=1.515 $X2=0
+ $Y2=0
cc_719 N_A_300_74#_c_944_n N_A_33_74#_c_1559_n 0.0166618f $X=1.64 $Y=0.515 $X2=0
+ $Y2=0
cc_720 N_A_300_74#_c_931_n N_A_33_74#_c_1560_n 0.00737917f $X=2.475 $Y=1.35
+ $X2=0 $Y2=0
cc_721 N_A_300_74#_c_932_n N_A_33_74#_c_1560_n 0.00235036f $X=2.995 $Y=1.47
+ $X2=0 $Y2=0
cc_722 N_A_300_74#_c_931_n N_A_33_74#_c_1634_n 0.006364f $X=2.475 $Y=1.35 $X2=0
+ $Y2=0
cc_723 N_A_300_74#_c_944_n N_A_33_74#_c_1634_n 0.0153439f $X=1.64 $Y=0.515 $X2=0
+ $Y2=0
cc_724 N_A_300_74#_c_947_n N_A_33_74#_c_1568_n 0.0048384f $X=2.46 $Y=1.765 $X2=0
+ $Y2=0
cc_725 N_A_300_74#_c_949_n N_A_33_74#_c_1568_n 0.0126174f $X=3.485 $Y=2.39 $X2=0
+ $Y2=0
cc_726 N_A_300_74#_c_950_n N_A_33_74#_c_1568_n 0.00908322f $X=3.145 $Y=2.39
+ $X2=0 $Y2=0
cc_727 N_A_300_74#_c_951_n N_A_33_74#_c_1568_n 5.42424e-19 $X=3.56 $Y=2.465
+ $X2=0 $Y2=0
cc_728 N_A_300_74#_c_947_n N_A_33_74#_c_1569_n 0.0109581f $X=2.46 $Y=1.765 $X2=0
+ $Y2=0
cc_729 N_A_300_74#_c_951_n N_A_33_74#_c_1569_n 0.00384622f $X=3.56 $Y=2.465
+ $X2=0 $Y2=0
cc_730 N_A_300_74#_c_947_n N_A_33_74#_c_1642_n 0.00905898f $X=2.46 $Y=1.765
+ $X2=0 $Y2=0
cc_731 N_A_300_74#_c_931_n N_A_33_74#_c_1562_n 0.00302447f $X=2.475 $Y=1.35
+ $X2=0 $Y2=0
cc_732 N_A_300_74#_c_941_n N_A_33_74#_c_1562_n 0.00132089f $X=3.07 $Y=1.47 $X2=0
+ $Y2=0
cc_733 N_A_300_74#_c_942_n N_VGND_M1010_s 0.00302838f $X=2.08 $Y=1.515 $X2=0
+ $Y2=0
cc_734 N_A_300_74#_c_944_n N_VGND_M1010_s 0.00711052f $X=1.64 $Y=0.515 $X2=0
+ $Y2=0
cc_735 N_A_300_74#_c_944_n N_VGND_c_1703_n 0.018056f $X=1.64 $Y=0.515 $X2=0
+ $Y2=0
cc_736 N_A_300_74#_c_931_n N_VGND_c_1704_n 0.00401707f $X=2.475 $Y=1.35 $X2=0
+ $Y2=0
cc_737 N_A_300_74#_c_944_n N_VGND_c_1704_n 0.0203575f $X=1.64 $Y=0.515 $X2=0
+ $Y2=0
cc_738 N_A_300_74#_c_936_n N_VGND_c_1705_n 0.0251635f $X=6.18 $Y=0.18 $X2=0
+ $Y2=0
cc_739 N_A_300_74#_c_944_n N_VGND_c_1709_n 0.0188466f $X=1.64 $Y=0.515 $X2=0
+ $Y2=0
cc_740 N_A_300_74#_c_931_n N_VGND_c_1710_n 0.00374483f $X=2.475 $Y=1.35 $X2=0
+ $Y2=0
cc_741 N_A_300_74#_c_937_n N_VGND_c_1710_n 0.0279684f $X=4.25 $Y=0.18 $X2=0
+ $Y2=0
cc_742 N_A_300_74#_c_936_n N_VGND_c_1711_n 0.0230598f $X=6.18 $Y=0.18 $X2=0
+ $Y2=0
cc_743 N_A_300_74#_c_931_n N_VGND_c_1714_n 0.00505379f $X=2.475 $Y=1.35 $X2=0
+ $Y2=0
cc_744 N_A_300_74#_c_936_n N_VGND_c_1714_n 0.0470713f $X=6.18 $Y=0.18 $X2=0
+ $Y2=0
cc_745 N_A_300_74#_c_937_n N_VGND_c_1714_n 0.00563078f $X=4.25 $Y=0.18 $X2=0
+ $Y2=0
cc_746 N_A_300_74#_c_944_n N_VGND_c_1714_n 0.0192545f $X=1.64 $Y=0.515 $X2=0
+ $Y2=0
cc_747 N_A_1598_93#_c_1138_n N_A_1266_119#_c_1226_n 0.0048734f $X=9.475 $Y=1.965
+ $X2=0 $Y2=0
cc_748 N_A_1598_93#_c_1139_n N_A_1266_119#_c_1226_n 0.00750942f $X=9.475
+ $Y=0.765 $X2=0 $Y2=0
cc_749 N_A_1598_93#_c_1144_n N_A_1266_119#_c_1227_n 0.00514416f $X=9.39 $Y=2.05
+ $X2=0 $Y2=0
cc_750 N_A_1598_93#_c_1146_n N_A_1266_119#_c_1227_n 0.00291268f $X=8.865 $Y=2.15
+ $X2=0 $Y2=0
cc_751 N_A_1598_93#_c_1143_n N_A_1266_119#_c_1237_n 0.00130111f $X=8.845 $Y=2.75
+ $X2=0 $Y2=0
cc_752 N_A_1598_93#_c_1144_n N_A_1266_119#_c_1237_n 0.00755711f $X=9.39 $Y=2.05
+ $X2=0 $Y2=0
cc_753 N_A_1598_93#_c_1146_n N_A_1266_119#_c_1237_n 0.015254f $X=8.865 $Y=2.15
+ $X2=0 $Y2=0
cc_754 N_A_1598_93#_c_1143_n N_A_1266_119#_c_1238_n 0.0111813f $X=8.845 $Y=2.75
+ $X2=0 $Y2=0
cc_755 N_A_1598_93#_c_1144_n N_A_1266_119#_c_1228_n 6.15368e-19 $X=9.39 $Y=2.05
+ $X2=0 $Y2=0
cc_756 N_A_1598_93#_c_1138_n N_A_1266_119#_c_1228_n 0.0128412f $X=9.475 $Y=1.965
+ $X2=0 $Y2=0
cc_757 N_A_1598_93#_c_1139_n N_A_1266_119#_c_1228_n 8.36802e-19 $X=9.475
+ $Y=0.765 $X2=0 $Y2=0
cc_758 N_A_1598_93#_c_1144_n N_A_1266_119#_c_1239_n 0.0109475f $X=9.39 $Y=2.05
+ $X2=0 $Y2=0
cc_759 N_A_1598_93#_c_1138_n N_A_1266_119#_c_1239_n 0.00680794f $X=9.475
+ $Y=1.965 $X2=0 $Y2=0
cc_760 N_A_1598_93#_c_1138_n N_A_1266_119#_c_1229_n 7.21124e-19 $X=9.475
+ $Y=1.965 $X2=0 $Y2=0
cc_761 N_A_1598_93#_c_1139_n N_A_1266_119#_c_1229_n 7.36949e-19 $X=9.475
+ $Y=0.765 $X2=0 $Y2=0
cc_762 N_A_1598_93#_c_1144_n N_A_1266_119#_c_1240_n 3.81375e-19 $X=9.39 $Y=2.05
+ $X2=0 $Y2=0
cc_763 N_A_1598_93#_c_1139_n N_A_1266_119#_c_1230_n 0.0071021f $X=9.475 $Y=0.765
+ $X2=0 $Y2=0
cc_764 N_A_1598_93#_M1000_g N_A_1266_119#_c_1266_n 0.00369318f $X=8.065 $Y=0.805
+ $X2=0 $Y2=0
cc_765 N_A_1598_93#_M1000_g N_A_1266_119#_c_1231_n 0.00375809f $X=8.065 $Y=0.805
+ $X2=0 $Y2=0
cc_766 N_A_1598_93#_M1000_g N_A_1266_119#_c_1232_n 0.0199131f $X=8.065 $Y=0.805
+ $X2=0 $Y2=0
cc_767 N_A_1598_93#_c_1141_n N_A_1266_119#_c_1232_n 0.00132521f $X=8.08 $Y=2.465
+ $X2=0 $Y2=0
cc_768 N_A_1598_93#_c_1142_n N_A_1266_119#_c_1232_n 0.0293641f $X=8.68 $Y=2.15
+ $X2=0 $Y2=0
cc_769 N_A_1598_93#_M1000_g N_A_1266_119#_c_1233_n 0.0157592f $X=8.065 $Y=0.805
+ $X2=0 $Y2=0
cc_770 N_A_1598_93#_c_1142_n N_A_1266_119#_c_1233_n 0.0023008f $X=8.68 $Y=2.15
+ $X2=0 $Y2=0
cc_771 N_A_1598_93#_c_1146_n N_A_1266_119#_c_1233_n 0.00676946f $X=8.865 $Y=2.15
+ $X2=0 $Y2=0
cc_772 N_A_1598_93#_c_1141_n N_A_1266_119#_c_1243_n 0.00189609f $X=8.08 $Y=2.465
+ $X2=0 $Y2=0
cc_773 N_A_1598_93#_c_1144_n N_A_1266_119#_c_1234_n 0.0128235f $X=9.39 $Y=2.05
+ $X2=0 $Y2=0
cc_774 N_A_1598_93#_c_1138_n N_A_1266_119#_c_1234_n 0.0502151f $X=9.475 $Y=1.965
+ $X2=0 $Y2=0
cc_775 N_A_1598_93#_c_1146_n N_A_1266_119#_c_1234_n 0.0110236f $X=8.865 $Y=2.15
+ $X2=0 $Y2=0
cc_776 N_A_1598_93#_c_1139_n N_A_1266_119#_c_1234_n 0.0121056f $X=9.475 $Y=0.765
+ $X2=0 $Y2=0
cc_777 N_A_1598_93#_c_1138_n N_A_1266_119#_c_1235_n 0.0103445f $X=9.475 $Y=1.965
+ $X2=0 $Y2=0
cc_778 N_A_1598_93#_c_1143_n N_A_1934_94#_c_1371_n 0.00529924f $X=8.845 $Y=2.75
+ $X2=0 $Y2=0
cc_779 N_A_1598_93#_c_1146_n N_A_1934_94#_c_1371_n 9.63229e-19 $X=8.865 $Y=2.15
+ $X2=0 $Y2=0
cc_780 N_A_1598_93#_c_1138_n N_A_1934_94#_c_1366_n 0.0270211f $X=9.475 $Y=1.965
+ $X2=0 $Y2=0
cc_781 N_A_1598_93#_c_1139_n N_A_1934_94#_c_1366_n 0.0315201f $X=9.475 $Y=0.765
+ $X2=0 $Y2=0
cc_782 N_A_1598_93#_c_1144_n N_A_1934_94#_c_1367_n 0.0140451f $X=9.39 $Y=2.05
+ $X2=0 $Y2=0
cc_783 N_A_1598_93#_c_1138_n N_A_1934_94#_c_1367_n 0.0238206f $X=9.475 $Y=1.965
+ $X2=0 $Y2=0
cc_784 N_A_1598_93#_c_1138_n N_A_1934_94#_c_1369_n 0.0278717f $X=9.475 $Y=1.965
+ $X2=0 $Y2=0
cc_785 N_A_1598_93#_c_1141_n N_VPWR_c_1432_n 0.0154036f $X=8.08 $Y=2.465 $X2=0
+ $Y2=0
cc_786 N_A_1598_93#_c_1142_n N_VPWR_c_1432_n 0.0267292f $X=8.68 $Y=2.15 $X2=0
+ $Y2=0
cc_787 N_A_1598_93#_c_1143_n N_VPWR_c_1432_n 0.0304142f $X=8.845 $Y=2.75 $X2=0
+ $Y2=0
cc_788 N_A_1598_93#_c_1143_n N_VPWR_c_1433_n 0.0309026f $X=8.845 $Y=2.75 $X2=0
+ $Y2=0
cc_789 N_A_1598_93#_c_1144_n N_VPWR_c_1433_n 0.0121819f $X=9.39 $Y=2.05 $X2=0
+ $Y2=0
cc_790 N_A_1598_93#_c_1141_n N_VPWR_c_1435_n 0.00413917f $X=8.08 $Y=2.465 $X2=0
+ $Y2=0
cc_791 N_A_1598_93#_c_1143_n N_VPWR_c_1442_n 0.014552f $X=8.845 $Y=2.75 $X2=0
+ $Y2=0
cc_792 N_A_1598_93#_c_1141_n N_VPWR_c_1424_n 0.0085536f $X=8.08 $Y=2.465 $X2=0
+ $Y2=0
cc_793 N_A_1598_93#_c_1143_n N_VPWR_c_1424_n 0.0119791f $X=8.845 $Y=2.75 $X2=0
+ $Y2=0
cc_794 N_A_1598_93#_M1000_g N_VGND_c_1706_n 0.00889071f $X=8.065 $Y=0.805 $X2=0
+ $Y2=0
cc_795 N_A_1598_93#_c_1139_n N_VGND_c_1706_n 0.0110474f $X=9.475 $Y=0.765 $X2=0
+ $Y2=0
cc_796 N_A_1598_93#_M1000_g N_VGND_c_1711_n 0.0035863f $X=8.065 $Y=0.805 $X2=0
+ $Y2=0
cc_797 N_A_1598_93#_c_1139_n N_VGND_c_1712_n 0.0112924f $X=9.475 $Y=0.765 $X2=0
+ $Y2=0
cc_798 N_A_1598_93#_M1000_g N_VGND_c_1714_n 0.00401353f $X=8.065 $Y=0.805 $X2=0
+ $Y2=0
cc_799 N_A_1598_93#_c_1139_n N_VGND_c_1714_n 0.0158807f $X=9.475 $Y=0.765 $X2=0
+ $Y2=0
cc_800 N_A_1266_119#_c_1229_n N_A_1934_94#_c_1364_n 0.0160558f $X=10.03 $Y=1.125
+ $X2=0 $Y2=0
cc_801 N_A_1266_119#_c_1239_n N_A_1934_94#_c_1365_n 0.00551483f $X=9.965 $Y=1.97
+ $X2=0 $Y2=0
cc_802 N_A_1266_119#_c_1240_n N_A_1934_94#_c_1365_n 0.0170234f $X=10.04 $Y=2.045
+ $X2=0 $Y2=0
cc_803 N_A_1266_119#_c_1237_n N_A_1934_94#_c_1371_n 0.00273194f $X=9.07 $Y=2.375
+ $X2=0 $Y2=0
cc_804 N_A_1266_119#_c_1238_n N_A_1934_94#_c_1371_n 0.0015885f $X=9.07 $Y=2.465
+ $X2=0 $Y2=0
cc_805 N_A_1266_119#_c_1239_n N_A_1934_94#_c_1371_n 0.00292339f $X=9.965 $Y=1.97
+ $X2=0 $Y2=0
cc_806 N_A_1266_119#_c_1240_n N_A_1934_94#_c_1371_n 0.00167606f $X=10.04
+ $Y=2.045 $X2=0 $Y2=0
cc_807 N_A_1266_119#_c_1240_n N_A_1934_94#_c_1372_n 0.00842612f $X=10.04
+ $Y=2.045 $X2=0 $Y2=0
cc_808 N_A_1266_119#_c_1226_n N_A_1934_94#_c_1366_n 0.00140435f $X=8.995
+ $Y=1.125 $X2=0 $Y2=0
cc_809 N_A_1266_119#_c_1228_n N_A_1934_94#_c_1366_n 0.0161335f $X=9.955 $Y=1.2
+ $X2=0 $Y2=0
cc_810 N_A_1266_119#_c_1229_n N_A_1934_94#_c_1366_n 0.010444f $X=10.03 $Y=1.125
+ $X2=0 $Y2=0
cc_811 N_A_1266_119#_c_1237_n N_A_1934_94#_c_1367_n 0.00438224f $X=9.07 $Y=2.375
+ $X2=0 $Y2=0
cc_812 N_A_1266_119#_c_1239_n N_A_1934_94#_c_1367_n 0.0166743f $X=9.965 $Y=1.97
+ $X2=0 $Y2=0
cc_813 N_A_1266_119#_c_1240_n N_A_1934_94#_c_1367_n 0.00434926f $X=10.04
+ $Y=2.045 $X2=0 $Y2=0
cc_814 N_A_1266_119#_c_1228_n N_A_1934_94#_c_1368_n 0.00434645f $X=9.955 $Y=1.2
+ $X2=0 $Y2=0
cc_815 N_A_1266_119#_c_1239_n N_A_1934_94#_c_1368_n 0.00425121f $X=9.965 $Y=1.97
+ $X2=0 $Y2=0
cc_816 N_A_1266_119#_c_1232_n N_VPWR_c_1432_n 8.41136e-19 $X=7.815 $Y=2.535
+ $X2=0 $Y2=0
cc_817 N_A_1266_119#_c_1243_n N_VPWR_c_1432_n 0.0157089f $X=7.435 $Y=2.7 $X2=0
+ $Y2=0
cc_818 N_A_1266_119#_c_1238_n N_VPWR_c_1433_n 0.00729942f $X=9.07 $Y=2.465 $X2=0
+ $Y2=0
cc_819 N_A_1266_119#_c_1239_n N_VPWR_c_1433_n 0.00128121f $X=9.965 $Y=1.97 $X2=0
+ $Y2=0
cc_820 N_A_1266_119#_c_1240_n N_VPWR_c_1433_n 0.00366284f $X=10.04 $Y=2.045
+ $X2=0 $Y2=0
cc_821 N_A_1266_119#_c_1240_n N_VPWR_c_1434_n 0.00784561f $X=10.04 $Y=2.045
+ $X2=0 $Y2=0
cc_822 N_A_1266_119#_c_1241_n N_VPWR_c_1435_n 0.0150066f $X=7.435 $Y=2.7 $X2=0
+ $Y2=0
cc_823 N_A_1266_119#_c_1243_n N_VPWR_c_1435_n 0.00884848f $X=7.435 $Y=2.7 $X2=0
+ $Y2=0
cc_824 N_A_1266_119#_c_1240_n N_VPWR_c_1437_n 0.00445602f $X=10.04 $Y=2.045
+ $X2=0 $Y2=0
cc_825 N_A_1266_119#_c_1238_n N_VPWR_c_1442_n 0.00445602f $X=9.07 $Y=2.465 $X2=0
+ $Y2=0
cc_826 N_A_1266_119#_c_1238_n N_VPWR_c_1424_n 0.00900303f $X=9.07 $Y=2.465 $X2=0
+ $Y2=0
cc_827 N_A_1266_119#_c_1240_n N_VPWR_c_1424_n 0.00862274f $X=10.04 $Y=2.045
+ $X2=0 $Y2=0
cc_828 N_A_1266_119#_c_1241_n N_VPWR_c_1424_n 0.0187253f $X=7.435 $Y=2.7 $X2=0
+ $Y2=0
cc_829 N_A_1266_119#_c_1243_n N_VPWR_c_1424_n 0.013677f $X=7.435 $Y=2.7 $X2=0
+ $Y2=0
cc_830 N_A_1266_119#_c_1243_n A_1547_508# 0.00356592f $X=7.435 $Y=2.7 $X2=-0.19
+ $Y2=-0.245
cc_831 N_A_1266_119#_c_1228_n N_Q_c_1675_n 2.48707e-19 $X=9.955 $Y=1.2 $X2=0
+ $Y2=0
cc_832 N_A_1266_119#_c_1239_n Q 6.01794e-19 $X=9.965 $Y=1.97 $X2=0 $Y2=0
cc_833 N_A_1266_119#_c_1240_n Q 4.02579e-19 $X=10.04 $Y=2.045 $X2=0 $Y2=0
cc_834 N_A_1266_119#_c_1226_n N_VGND_c_1706_n 0.00147671f $X=8.995 $Y=1.125
+ $X2=0 $Y2=0
cc_835 N_A_1266_119#_c_1266_n N_VGND_c_1706_n 0.0196844f $X=7.73 $Y=0.79 $X2=0
+ $Y2=0
cc_836 N_A_1266_119#_c_1233_n N_VGND_c_1706_n 0.0254301f $X=8.92 $Y=1.21 $X2=0
+ $Y2=0
cc_837 N_A_1266_119#_c_1229_n N_VGND_c_1707_n 0.0072589f $X=10.03 $Y=1.125 $X2=0
+ $Y2=0
cc_838 N_A_1266_119#_c_1266_n N_VGND_c_1711_n 0.0212446f $X=7.73 $Y=0.79 $X2=0
+ $Y2=0
cc_839 N_A_1266_119#_c_1226_n N_VGND_c_1712_n 0.00414396f $X=8.995 $Y=1.125
+ $X2=0 $Y2=0
cc_840 N_A_1266_119#_c_1229_n N_VGND_c_1712_n 0.00486718f $X=10.03 $Y=1.125
+ $X2=0 $Y2=0
cc_841 N_A_1266_119#_c_1226_n N_VGND_c_1714_n 0.00477801f $X=8.995 $Y=1.125
+ $X2=0 $Y2=0
cc_842 N_A_1266_119#_c_1229_n N_VGND_c_1714_n 0.00514438f $X=10.03 $Y=1.125
+ $X2=0 $Y2=0
cc_843 N_A_1266_119#_c_1266_n N_VGND_c_1714_n 0.0353228f $X=7.73 $Y=0.79 $X2=0
+ $Y2=0
cc_844 N_A_1266_119#_c_1266_n A_1550_119# 0.00494929f $X=7.73 $Y=0.79 $X2=-0.19
+ $Y2=-0.245
cc_845 N_A_1266_119#_c_1231_n A_1550_119# 6.55526e-19 $X=7.815 $Y=1.125
+ $X2=-0.19 $Y2=-0.245
cc_846 N_A_1934_94#_c_1372_n N_VPWR_c_1433_n 0.0346921f $X=9.815 $Y=2.815 $X2=0
+ $Y2=0
cc_847 N_A_1934_94#_c_1365_n N_VPWR_c_1434_n 0.00845898f $X=10.545 $Y=1.765
+ $X2=0 $Y2=0
cc_848 N_A_1934_94#_c_1367_n N_VPWR_c_1434_n 0.0341417f $X=9.815 $Y=2.27 $X2=0
+ $Y2=0
cc_849 N_A_1934_94#_c_1368_n N_VPWR_c_1434_n 0.0104409f $X=10.48 $Y=1.485 $X2=0
+ $Y2=0
cc_850 N_A_1934_94#_c_1372_n N_VPWR_c_1437_n 0.0145919f $X=9.815 $Y=2.815 $X2=0
+ $Y2=0
cc_851 N_A_1934_94#_c_1365_n N_VPWR_c_1443_n 0.00445602f $X=10.545 $Y=1.765
+ $X2=0 $Y2=0
cc_852 N_A_1934_94#_c_1365_n N_VPWR_c_1424_n 0.00861717f $X=10.545 $Y=1.765
+ $X2=0 $Y2=0
cc_853 N_A_1934_94#_c_1372_n N_VPWR_c_1424_n 0.0120459f $X=9.815 $Y=2.815 $X2=0
+ $Y2=0
cc_854 N_A_1934_94#_c_1364_n N_Q_c_1675_n 0.00640271f $X=10.54 $Y=1.32 $X2=0
+ $Y2=0
cc_855 N_A_1934_94#_c_1364_n N_Q_c_1676_n 0.00241276f $X=10.54 $Y=1.32 $X2=0
+ $Y2=0
cc_856 N_A_1934_94#_c_1366_n N_Q_c_1676_n 5.13862e-19 $X=9.815 $Y=0.745 $X2=0
+ $Y2=0
cc_857 N_A_1934_94#_c_1368_n N_Q_c_1676_n 0.00188005f $X=10.48 $Y=1.485 $X2=0
+ $Y2=0
cc_858 N_A_1934_94#_c_1365_n Q 0.0049232f $X=10.545 $Y=1.765 $X2=0 $Y2=0
cc_859 N_A_1934_94#_c_1367_n Q 0.0072771f $X=9.815 $Y=2.27 $X2=0 $Y2=0
cc_860 N_A_1934_94#_c_1368_n Q 7.18422e-19 $X=10.48 $Y=1.485 $X2=0 $Y2=0
cc_861 N_A_1934_94#_c_1365_n Q 0.0126267f $X=10.545 $Y=1.765 $X2=0 $Y2=0
cc_862 N_A_1934_94#_c_1364_n N_Q_c_1677_n 0.0040915f $X=10.54 $Y=1.32 $X2=0
+ $Y2=0
cc_863 N_A_1934_94#_c_1365_n N_Q_c_1677_n 0.0119541f $X=10.545 $Y=1.765 $X2=0
+ $Y2=0
cc_864 N_A_1934_94#_c_1368_n N_Q_c_1677_n 0.0262114f $X=10.48 $Y=1.485 $X2=0
+ $Y2=0
cc_865 N_A_1934_94#_c_1364_n N_VGND_c_1707_n 0.00292117f $X=10.54 $Y=1.32 $X2=0
+ $Y2=0
cc_866 N_A_1934_94#_c_1365_n N_VGND_c_1707_n 0.00216466f $X=10.545 $Y=1.765
+ $X2=0 $Y2=0
cc_867 N_A_1934_94#_c_1366_n N_VGND_c_1707_n 0.024751f $X=9.815 $Y=0.745 $X2=0
+ $Y2=0
cc_868 N_A_1934_94#_c_1368_n N_VGND_c_1707_n 0.0194281f $X=10.48 $Y=1.485 $X2=0
+ $Y2=0
cc_869 N_A_1934_94#_c_1366_n N_VGND_c_1712_n 0.00541117f $X=9.815 $Y=0.745 $X2=0
+ $Y2=0
cc_870 N_A_1934_94#_c_1364_n N_VGND_c_1713_n 0.00485341f $X=10.54 $Y=1.32 $X2=0
+ $Y2=0
cc_871 N_A_1934_94#_c_1364_n N_VGND_c_1714_n 0.00514438f $X=10.54 $Y=1.32 $X2=0
+ $Y2=0
cc_872 N_A_1934_94#_c_1366_n N_VGND_c_1714_n 0.00809617f $X=9.815 $Y=0.745 $X2=0
+ $Y2=0
cc_873 N_VPWR_c_1426_n N_A_33_74#_c_1564_n 0.0309025f $X=0.275 $Y=2.75 $X2=0
+ $Y2=0
cc_874 N_VPWR_c_1427_n N_A_33_74#_c_1564_n 0.0124773f $X=1.225 $Y=2.775 $X2=0
+ $Y2=0
cc_875 N_VPWR_c_1439_n N_A_33_74#_c_1564_n 0.0110241f $X=1.06 $Y=3.33 $X2=0
+ $Y2=0
cc_876 N_VPWR_c_1424_n N_A_33_74#_c_1564_n 0.00909194f $X=10.8 $Y=3.33 $X2=0
+ $Y2=0
cc_877 N_VPWR_M1007_d N_A_33_74#_c_1565_n 0.00265359f $X=1.025 $Y=2.54 $X2=0
+ $Y2=0
cc_878 N_VPWR_M1009_s N_A_33_74#_c_1565_n 0.0057427f $X=2.09 $Y=1.84 $X2=0 $Y2=0
cc_879 N_VPWR_c_1427_n N_A_33_74#_c_1565_n 0.00799774f $X=1.225 $Y=2.775 $X2=0
+ $Y2=0
cc_880 N_VPWR_c_1428_n N_A_33_74#_c_1565_n 0.0205174f $X=2.235 $Y=2.82 $X2=0
+ $Y2=0
cc_881 N_VPWR_c_1424_n N_A_33_74#_c_1565_n 0.0237962f $X=10.8 $Y=3.33 $X2=0
+ $Y2=0
cc_882 N_VPWR_M1007_d N_A_33_74#_c_1566_n 0.0047622f $X=1.025 $Y=2.54 $X2=0
+ $Y2=0
cc_883 N_VPWR_c_1427_n N_A_33_74#_c_1566_n 0.0131939f $X=1.225 $Y=2.775 $X2=0
+ $Y2=0
cc_884 N_VPWR_c_1424_n N_A_33_74#_c_1566_n 5.66126e-19 $X=10.8 $Y=3.33 $X2=0
+ $Y2=0
cc_885 N_VPWR_c_1424_n N_A_33_74#_c_1568_n 0.0226376f $X=10.8 $Y=3.33 $X2=0
+ $Y2=0
cc_886 N_VPWR_c_1441_n N_A_33_74#_c_1569_n 0.011048f $X=4.46 $Y=3.33 $X2=0 $Y2=0
cc_887 N_VPWR_c_1424_n N_A_33_74#_c_1569_n 0.00915249f $X=10.8 $Y=3.33 $X2=0
+ $Y2=0
cc_888 N_VPWR_c_1428_n N_A_33_74#_c_1642_n 0.00111477f $X=2.235 $Y=2.82 $X2=0
+ $Y2=0
cc_889 N_VPWR_c_1424_n N_A_33_74#_c_1642_n 0.00355367f $X=10.8 $Y=3.33 $X2=0
+ $Y2=0
cc_890 N_VPWR_c_1434_n Q 0.0581843f $X=10.315 $Y=2.265 $X2=0 $Y2=0
cc_891 N_VPWR_c_1443_n Q 0.0154862f $X=10.8 $Y=3.33 $X2=0 $Y2=0
cc_892 N_VPWR_c_1424_n Q 0.0127853f $X=10.8 $Y=3.33 $X2=0 $Y2=0
cc_893 N_A_33_74#_c_1561_n A_120_74# 0.00489958f $X=0.625 $Y=0.57 $X2=-0.19
+ $Y2=-0.245
cc_894 N_A_33_74#_c_1559_n N_VGND_M1010_s 0.00460265f $X=2.42 $Y=2.315 $X2=0
+ $Y2=0
cc_895 N_A_33_74#_c_1634_n N_VGND_M1010_s 0.00196634f $X=2.505 $Y=0.72 $X2=0
+ $Y2=0
cc_896 N_A_33_74#_c_1558_n N_VGND_c_1703_n 9.42187e-19 $X=0.625 $Y=2.18 $X2=0
+ $Y2=0
cc_897 N_A_33_74#_c_1561_n N_VGND_c_1703_n 0.0120647f $X=0.625 $Y=0.57 $X2=0
+ $Y2=0
cc_898 N_A_33_74#_c_1634_n N_VGND_c_1704_n 9.594e-19 $X=2.505 $Y=0.72 $X2=0
+ $Y2=0
cc_899 N_A_33_74#_c_1561_n N_VGND_c_1708_n 0.0239076f $X=0.625 $Y=0.57 $X2=0
+ $Y2=0
cc_900 N_A_33_74#_c_1560_n N_VGND_c_1710_n 0.00887637f $X=3.115 $Y=0.72 $X2=0
+ $Y2=0
cc_901 N_A_33_74#_c_1634_n N_VGND_c_1710_n 0.0023627f $X=2.505 $Y=0.72 $X2=0
+ $Y2=0
cc_902 N_A_33_74#_c_1560_n N_VGND_c_1714_n 0.0152481f $X=3.115 $Y=0.72 $X2=0
+ $Y2=0
cc_903 N_A_33_74#_c_1634_n N_VGND_c_1714_n 0.00469507f $X=2.505 $Y=0.72 $X2=0
+ $Y2=0
cc_904 N_A_33_74#_c_1561_n N_VGND_c_1714_n 0.0198316f $X=0.625 $Y=0.57 $X2=0
+ $Y2=0
cc_905 N_Q_c_1675_n N_VGND_c_1707_n 0.0261897f $X=10.755 $Y=0.605 $X2=0 $Y2=0
cc_906 N_Q_c_1675_n N_VGND_c_1713_n 0.0118258f $X=10.755 $Y=0.605 $X2=0 $Y2=0
cc_907 N_Q_c_1675_n N_VGND_c_1714_n 0.0126447f $X=10.755 $Y=0.605 $X2=0 $Y2=0
