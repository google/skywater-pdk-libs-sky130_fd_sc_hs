* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hs__einvn_2 A TE_B VGND VNB VPB VPWR Z
M1000 VGND a_115_464# a_231_74# VNB nlowvt w=740000u l=150000u
+  ad=3.269e+11p pd=3.45e+06u as=6.176e+11p ps=6.17e+06u
M1001 a_231_74# A Z VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1002 VPWR TE_B a_227_368# VPB pshort w=1.12e+06u l=150000u
+  ad=5.216e+11p pd=4.7e+06u as=9.968e+11p ps=8.5e+06u
M1003 a_231_74# a_115_464# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_227_368# TE_B VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 Z A a_227_368# VPB pshort w=1.12e+06u l=150000u
+  ad=3.36e+11p pd=2.84e+06u as=0p ps=0u
M1006 a_227_368# A Z VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_115_464# TE_B VPWR VPB pshort w=640000u l=150000u
+  ad=1.856e+11p pd=1.86e+06u as=0p ps=0u
M1008 Z A a_231_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_115_464# TE_B VGND VNB nlowvt w=420000u l=150000u
+  ad=1.197e+11p pd=1.41e+06u as=0p ps=0u
.ends
