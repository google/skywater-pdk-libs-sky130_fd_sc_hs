# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_hs__a32o_4
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_hs__a32o_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  8.160000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.635000 1.450000 6.115000 1.780000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.440000 1.470000 5.350000 1.790000 ;
        RECT 5.180000 1.790000 5.350000 1.950000 ;
        RECT 5.180000 1.950000 6.595000 2.120000 ;
        RECT 6.425000 1.440000 6.825000 1.770000 ;
        RECT 6.425000 1.770000 6.595000 1.950000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.065000 1.450000 8.035000 1.780000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.005000 1.450000 3.715000 1.780000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.505000 1.450000 2.835000 1.780000 ;
        RECT 2.570000 0.255000 4.415000 0.425000 ;
        RECT 2.570000 0.425000 2.740000 1.450000 ;
        RECT 4.085000 0.425000 4.415000 0.585000 ;
    END
  END B2
  PIN X
    ANTENNADIFFAREA  1.097500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 0.930000 1.900000 1.180000 ;
        RECT 0.125000 1.180000 0.355000 1.480000 ;
        RECT 0.125000 1.480000 0.815000 1.650000 ;
        RECT 0.565000 1.650000 0.815000 1.850000 ;
        RECT 0.565000 1.850000 1.795000 2.020000 ;
        RECT 0.565000 2.020000 0.815000 2.980000 ;
        RECT 0.615000 0.410000 0.820000 0.930000 ;
        RECT 1.515000 2.020000 1.795000 3.000000 ;
        RECT 1.570000 0.430000 1.900000 0.930000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 8.160000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 8.160000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 8.160000 0.085000 ;
      RECT 0.000000  3.245000 8.160000 3.415000 ;
      RECT 0.115000  0.085000 0.445000 0.760000 ;
      RECT 0.115000  1.820000 0.365000 3.245000 ;
      RECT 0.985000  1.350000 2.185000 1.680000 ;
      RECT 0.990000  0.085000 1.400000 0.760000 ;
      RECT 1.015000  2.190000 1.345000 3.245000 ;
      RECT 1.965000  2.290000 2.295000 3.245000 ;
      RECT 2.015000  1.680000 2.185000 1.950000 ;
      RECT 2.015000  1.950000 4.355000 2.120000 ;
      RECT 2.070000  0.085000 2.400000 1.180000 ;
      RECT 2.525000  2.290000 2.855000 2.905000 ;
      RECT 2.525000  2.905000 4.925000 3.075000 ;
      RECT 2.910000  0.595000 3.240000 0.755000 ;
      RECT 2.910000  0.755000 4.180000 0.925000 ;
      RECT 2.910000  0.925000 3.240000 1.210000 ;
      RECT 3.025000  2.120000 3.355000 2.735000 ;
      RECT 3.420000  1.095000 3.750000 1.110000 ;
      RECT 3.420000  1.110000 6.130000 1.280000 ;
      RECT 3.525000  2.290000 3.855000 2.905000 ;
      RECT 3.885000  1.280000 4.055000 1.950000 ;
      RECT 4.025000  2.120000 4.355000 2.735000 ;
      RECT 4.350000  0.755000 4.755000 0.940000 ;
      RECT 4.585000  0.085000 4.755000 0.755000 ;
      RECT 4.595000  1.960000 4.925000 2.290000 ;
      RECT 4.595000  2.290000 7.095000 2.460000 ;
      RECT 4.595000  2.460000 4.925000 2.905000 ;
      RECT 4.940000  0.255000 6.990000 0.425000 ;
      RECT 4.940000  0.425000 5.190000 0.940000 ;
      RECT 5.210000  2.630000 5.615000 3.245000 ;
      RECT 5.370000  0.595000 6.560000 0.765000 ;
      RECT 5.370000  0.765000 5.620000 0.940000 ;
      RECT 5.785000  2.460000 6.115000 2.900000 ;
      RECT 5.800000  0.935000 6.130000 1.110000 ;
      RECT 6.285000  2.630000 6.645000 3.245000 ;
      RECT 6.310000  0.765000 6.560000 1.270000 ;
      RECT 6.740000  0.425000 6.990000 1.100000 ;
      RECT 6.740000  1.100000 8.045000 1.270000 ;
      RECT 6.765000  1.950000 8.045000 2.120000 ;
      RECT 6.765000  2.120000 7.095000 2.290000 ;
      RECT 6.815000  2.460000 7.095000 3.000000 ;
      RECT 7.190000  0.085000 7.545000 0.920000 ;
      RECT 7.265000  2.290000 7.545000 3.245000 ;
      RECT 7.715000  0.590000 8.045000 1.100000 ;
      RECT 7.715000  2.120000 8.045000 2.980000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
      RECT 7.835000 -0.085000 8.005000 0.085000 ;
      RECT 7.835000  3.245000 8.005000 3.415000 ;
  END
END sky130_fd_sc_hs__a32o_4
