* File: sky130_fd_sc_hs__a21boi_2.pxi.spice
* Created: Tue Sep  1 19:49:22 2020
* 
x_PM_SKY130_FD_SC_HS__A21BOI_2%B1_N N_B1_N_c_80_n N_B1_N_M1012_g N_B1_N_M1002_g
+ N_B1_N_c_82_n B1_N PM_SKY130_FD_SC_HS__A21BOI_2%B1_N
x_PM_SKY130_FD_SC_HS__A21BOI_2%A_62_94# N_A_62_94#_M1002_s N_A_62_94#_M1012_d
+ N_A_62_94#_M1003_g N_A_62_94#_c_118_n N_A_62_94#_M1005_g N_A_62_94#_M1009_g
+ N_A_62_94#_c_112_n N_A_62_94#_c_113_n N_A_62_94#_c_121_n N_A_62_94#_M1006_g
+ N_A_62_94#_c_114_n N_A_62_94#_c_115_n N_A_62_94#_c_116_n N_A_62_94#_c_122_n
+ N_A_62_94#_c_123_n N_A_62_94#_c_117_n N_A_62_94#_c_124_n
+ PM_SKY130_FD_SC_HS__A21BOI_2%A_62_94#
x_PM_SKY130_FD_SC_HS__A21BOI_2%A1 N_A1_c_192_n N_A1_M1007_g N_A1_M1000_g
+ N_A1_c_193_n N_A1_M1008_g N_A1_M1011_g A1 N_A1_c_190_n N_A1_c_191_n
+ PM_SKY130_FD_SC_HS__A21BOI_2%A1
x_PM_SKY130_FD_SC_HS__A21BOI_2%A2 N_A2_c_250_n N_A2_M1001_g N_A2_c_246_n
+ N_A2_M1004_g N_A2_c_247_n N_A2_M1013_g N_A2_c_251_n N_A2_M1010_g A2
+ N_A2_c_249_n PM_SKY130_FD_SC_HS__A21BOI_2%A2
x_PM_SKY130_FD_SC_HS__A21BOI_2%VPWR N_VPWR_M1012_s N_VPWR_M1007_d N_VPWR_M1001_s
+ N_VPWR_c_288_n N_VPWR_c_289_n N_VPWR_c_290_n N_VPWR_c_291_n VPWR
+ N_VPWR_c_292_n N_VPWR_c_293_n N_VPWR_c_294_n N_VPWR_c_287_n N_VPWR_c_296_n
+ N_VPWR_c_297_n PM_SKY130_FD_SC_HS__A21BOI_2%VPWR
x_PM_SKY130_FD_SC_HS__A21BOI_2%A_241_368# N_A_241_368#_M1005_s
+ N_A_241_368#_M1006_s N_A_241_368#_M1008_s N_A_241_368#_M1010_d
+ N_A_241_368#_c_341_n N_A_241_368#_c_342_n N_A_241_368#_c_343_n
+ N_A_241_368#_c_344_n N_A_241_368#_c_360_n N_A_241_368#_c_361_n
+ N_A_241_368#_c_345_n N_A_241_368#_c_346_n N_A_241_368#_c_347_n
+ N_A_241_368#_c_348_n PM_SKY130_FD_SC_HS__A21BOI_2%A_241_368#
x_PM_SKY130_FD_SC_HS__A21BOI_2%Y N_Y_M1003_d N_Y_M1000_s N_Y_M1005_d N_Y_c_401_n
+ N_Y_c_402_n N_Y_c_403_n N_Y_c_404_n N_Y_c_405_n Y N_Y_c_406_n N_Y_c_407_n
+ PM_SKY130_FD_SC_HS__A21BOI_2%Y
x_PM_SKY130_FD_SC_HS__A21BOI_2%VGND N_VGND_M1002_d N_VGND_M1009_s N_VGND_M1004_d
+ N_VGND_c_458_n N_VGND_c_459_n N_VGND_c_460_n N_VGND_c_461_n N_VGND_c_462_n
+ N_VGND_c_463_n VGND N_VGND_c_464_n N_VGND_c_465_n N_VGND_c_466_n
+ N_VGND_c_467_n N_VGND_c_468_n PM_SKY130_FD_SC_HS__A21BOI_2%VGND
x_PM_SKY130_FD_SC_HS__A21BOI_2%A_436_74# N_A_436_74#_M1000_d N_A_436_74#_M1011_d
+ N_A_436_74#_M1013_s N_A_436_74#_c_517_n N_A_436_74#_c_518_n
+ N_A_436_74#_c_530_n N_A_436_74#_c_524_n N_A_436_74#_c_519_n
+ N_A_436_74#_c_520_n PM_SKY130_FD_SC_HS__A21BOI_2%A_436_74#
cc_1 VNB N_B1_N_c_80_n 0.0117911f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.885
cc_2 VNB N_B1_N_M1002_g 0.0389049f $X=-0.19 $Y=-0.245 $X2=0.65 $Y2=0.79
cc_3 VNB N_B1_N_c_82_n 0.0255356f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.615
cc_4 VNB B1_N 0.0085963f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_5 VNB N_A_62_94#_M1003_g 0.0238777f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.615
cc_6 VNB N_A_62_94#_M1009_g 0.0256721f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_7 VNB N_A_62_94#_c_112_n 0.0154846f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_A_62_94#_c_113_n 0.0485631f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A_62_94#_c_114_n 0.0274788f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_62_94#_c_115_n 0.00519287f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_62_94#_c_116_n 0.00946887f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_62_94#_c_117_n 0.0170134f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A1_M1000_g 0.0246159f $X=-0.19 $Y=-0.245 $X2=0.65 $Y2=0.79
cc_14 VNB N_A1_M1011_g 0.0222596f $X=-0.19 $Y=-0.245 $X2=0.31 $Y2=1.615
cc_15 VNB N_A1_c_190_n 0.00102877f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A1_c_191_n 0.0535786f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A2_c_246_n 0.0168884f $X=-0.19 $Y=-0.245 $X2=0.65 $Y2=1.45
cc_18 VNB N_A2_c_247_n 0.0224993f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB A2 0.00752679f $X=-0.19 $Y=-0.245 $X2=0.31 $Y2=1.615
cc_20 VNB N_A2_c_249_n 0.0681622f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_VPWR_c_287_n 0.183584f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_Y_c_401_n 0.00178908f $X=-0.19 $Y=-0.245 $X2=0.31 $Y2=1.615
cc_23 VNB N_Y_c_402_n 0.00252401f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_Y_c_403_n 0.00316101f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_Y_c_404_n 0.00314005f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_Y_c_405_n 0.00402553f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_Y_c_406_n 0.00185509f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_Y_c_407_n 0.0220781f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_458_n 0.00948899f $X=-0.19 $Y=-0.245 $X2=0.31 $Y2=1.615
cc_30 VNB N_VGND_c_459_n 0.0151736f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_460_n 0.0117687f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_461_n 0.00396467f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_462_n 0.0247362f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_463_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_464_n 0.0382181f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_465_n 0.0178682f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_466_n 0.267893f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_467_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_468_n 0.00604233f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_436_74#_c_517_n 0.00820512f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_41 VNB N_A_436_74#_c_518_n 0.00160668f $X=-0.19 $Y=-0.245 $X2=0.31 $Y2=1.615
cc_42 VNB N_A_436_74#_c_519_n 0.0159805f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_436_74#_c_520_n 0.0207145f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VPB N_B1_N_c_80_n 0.0377352f $X=-0.19 $Y=1.66 $X2=0.585 $Y2=1.885
cc_45 VPB N_B1_N_c_82_n 0.0189871f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.615
cc_46 VPB B1_N 0.00521552f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_47 VPB N_A_62_94#_c_118_n 0.017108f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_48 VPB N_A_62_94#_c_112_n 0.0111815f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_49 VPB N_A_62_94#_c_113_n 0.00624366f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_50 VPB N_A_62_94#_c_121_n 0.0145849f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_51 VPB N_A_62_94#_c_122_n 0.00332341f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_52 VPB N_A_62_94#_c_123_n 0.0105928f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_53 VPB N_A_62_94#_c_124_n 0.00608507f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_54 VPB N_A1_c_192_n 0.0153302f $X=-0.19 $Y=1.66 $X2=0.585 $Y2=1.885
cc_55 VPB N_A1_c_193_n 0.0153972f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=1.615
cc_56 VPB N_A1_c_190_n 0.00361438f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_57 VPB N_A1_c_191_n 0.01263f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_58 VPB N_A2_c_250_n 0.0148084f $X=-0.19 $Y=1.66 $X2=0.585 $Y2=1.885
cc_59 VPB N_A2_c_251_n 0.0188573f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_60 VPB N_A2_c_249_n 0.0150151f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_61 VPB N_VPWR_c_288_n 0.013204f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_62 VPB N_VPWR_c_289_n 0.0517348f $X=-0.19 $Y=1.66 $X2=0.31 $Y2=1.615
cc_63 VPB N_VPWR_c_290_n 0.00329129f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_64 VPB N_VPWR_c_291_n 0.00329222f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_65 VPB N_VPWR_c_292_n 0.0519976f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_66 VPB N_VPWR_c_293_n 0.0164465f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_67 VPB N_VPWR_c_294_n 0.0177091f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_68 VPB N_VPWR_c_287_n 0.0813562f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_69 VPB N_VPWR_c_296_n 0.00601644f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_70 VPB N_VPWR_c_297_n 0.00638264f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_71 VPB N_A_241_368#_c_341_n 0.0114607f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_72 VPB N_A_241_368#_c_342_n 0.00524063f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_73 VPB N_A_241_368#_c_343_n 0.00449591f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_74 VPB N_A_241_368#_c_344_n 0.00321012f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_75 VPB N_A_241_368#_c_345_n 0.00180921f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_76 VPB N_A_241_368#_c_346_n 0.0175888f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_77 VPB N_A_241_368#_c_347_n 0.043203f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_78 VPB N_A_241_368#_c_348_n 0.0049323f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_79 N_B1_N_M1002_g N_A_62_94#_M1003_g 0.0146457f $X=0.65 $Y=0.79 $X2=0 $Y2=0
cc_80 N_B1_N_c_80_n N_A_62_94#_c_113_n 0.0146457f $X=0.585 $Y=1.885 $X2=0 $Y2=0
cc_81 N_B1_N_M1002_g N_A_62_94#_c_114_n 4.61877e-19 $X=0.65 $Y=0.79 $X2=0 $Y2=0
cc_82 N_B1_N_c_80_n N_A_62_94#_c_115_n 0.0022655f $X=0.585 $Y=1.885 $X2=0 $Y2=0
cc_83 N_B1_N_M1002_g N_A_62_94#_c_115_n 0.019447f $X=0.65 $Y=0.79 $X2=0 $Y2=0
cc_84 N_B1_N_c_82_n N_A_62_94#_c_116_n 0.00681442f $X=0.495 $Y=1.615 $X2=0 $Y2=0
cc_85 B1_N N_A_62_94#_c_116_n 0.0172883f $X=0.155 $Y=1.58 $X2=0 $Y2=0
cc_86 N_B1_N_c_80_n N_A_62_94#_c_122_n 0.00518959f $X=0.585 $Y=1.885 $X2=0 $Y2=0
cc_87 N_B1_N_c_80_n N_A_62_94#_c_123_n 0.00991534f $X=0.585 $Y=1.885 $X2=0 $Y2=0
cc_88 N_B1_N_M1002_g N_A_62_94#_c_117_n 0.00745999f $X=0.65 $Y=0.79 $X2=0 $Y2=0
cc_89 B1_N N_A_62_94#_c_117_n 0.0101785f $X=0.155 $Y=1.58 $X2=0 $Y2=0
cc_90 N_B1_N_c_80_n N_A_62_94#_c_124_n 0.00965756f $X=0.585 $Y=1.885 $X2=0 $Y2=0
cc_91 B1_N N_A_62_94#_c_124_n 0.00592225f $X=0.155 $Y=1.58 $X2=0 $Y2=0
cc_92 N_B1_N_c_80_n N_VPWR_c_289_n 0.00850665f $X=0.585 $Y=1.885 $X2=0 $Y2=0
cc_93 N_B1_N_c_82_n N_VPWR_c_289_n 0.00577732f $X=0.495 $Y=1.615 $X2=0 $Y2=0
cc_94 B1_N N_VPWR_c_289_n 0.0209147f $X=0.155 $Y=1.58 $X2=0 $Y2=0
cc_95 N_B1_N_c_80_n N_VPWR_c_292_n 0.00445602f $X=0.585 $Y=1.885 $X2=0 $Y2=0
cc_96 N_B1_N_c_80_n N_VPWR_c_287_n 0.00866122f $X=0.585 $Y=1.885 $X2=0 $Y2=0
cc_97 N_B1_N_c_80_n N_A_241_368#_c_341_n 0.00142885f $X=0.585 $Y=1.885 $X2=0
+ $Y2=0
cc_98 N_B1_N_c_80_n N_A_241_368#_c_343_n 0.00293173f $X=0.585 $Y=1.885 $X2=0
+ $Y2=0
cc_99 N_B1_N_M1002_g N_VGND_c_458_n 0.00577735f $X=0.65 $Y=0.79 $X2=0 $Y2=0
cc_100 N_B1_N_M1002_g N_VGND_c_462_n 0.00507111f $X=0.65 $Y=0.79 $X2=0 $Y2=0
cc_101 N_B1_N_M1002_g N_VGND_c_466_n 0.00514438f $X=0.65 $Y=0.79 $X2=0 $Y2=0
cc_102 N_A_62_94#_c_121_n N_A1_c_192_n 0.00928675f $X=2.005 $Y=1.765 $X2=-0.19
+ $Y2=-0.245
cc_103 N_A_62_94#_c_112_n N_A1_c_190_n 5.73974e-19 $X=1.93 $Y=1.69 $X2=0 $Y2=0
cc_104 N_A_62_94#_c_112_n N_A1_c_191_n 0.00739224f $X=1.93 $Y=1.69 $X2=0 $Y2=0
cc_105 N_A_62_94#_c_113_n N_A1_c_191_n 0.00305683f $X=1.645 $Y=1.69 $X2=0 $Y2=0
cc_106 N_A_62_94#_c_122_n N_VPWR_c_289_n 0.069074f $X=0.81 $Y=2.105 $X2=0 $Y2=0
cc_107 N_A_62_94#_c_118_n N_VPWR_c_292_n 0.00278271f $X=1.555 $Y=1.765 $X2=0
+ $Y2=0
cc_108 N_A_62_94#_c_121_n N_VPWR_c_292_n 0.00278271f $X=2.005 $Y=1.765 $X2=0
+ $Y2=0
cc_109 N_A_62_94#_c_123_n N_VPWR_c_292_n 0.0145938f $X=0.81 $Y=2.815 $X2=0 $Y2=0
cc_110 N_A_62_94#_c_118_n N_VPWR_c_287_n 0.00358624f $X=1.555 $Y=1.765 $X2=0
+ $Y2=0
cc_111 N_A_62_94#_c_121_n N_VPWR_c_287_n 0.00353907f $X=2.005 $Y=1.765 $X2=0
+ $Y2=0
cc_112 N_A_62_94#_c_123_n N_VPWR_c_287_n 0.0120466f $X=0.81 $Y=2.815 $X2=0 $Y2=0
cc_113 N_A_62_94#_c_118_n N_A_241_368#_c_341_n 0.00807154f $X=1.555 $Y=1.765
+ $X2=0 $Y2=0
cc_114 N_A_62_94#_c_113_n N_A_241_368#_c_341_n 0.00240798f $X=1.645 $Y=1.69
+ $X2=0 $Y2=0
cc_115 N_A_62_94#_c_117_n N_A_241_368#_c_341_n 0.0194066f $X=0.89 $Y=1.65 $X2=0
+ $Y2=0
cc_116 N_A_62_94#_c_124_n N_A_241_368#_c_341_n 0.0812758f $X=0.81 $Y=1.94 $X2=0
+ $Y2=0
cc_117 N_A_62_94#_c_118_n N_A_241_368#_c_342_n 0.0136535f $X=1.555 $Y=1.765
+ $X2=0 $Y2=0
cc_118 N_A_62_94#_c_121_n N_A_241_368#_c_342_n 0.012504f $X=2.005 $Y=1.765 $X2=0
+ $Y2=0
cc_119 N_A_62_94#_c_123_n N_A_241_368#_c_343_n 0.00613236f $X=0.81 $Y=2.815
+ $X2=0 $Y2=0
cc_120 N_A_62_94#_M1003_g N_Y_c_401_n 3.92313e-19 $X=1.14 $Y=0.74 $X2=0 $Y2=0
cc_121 N_A_62_94#_M1009_g N_Y_c_401_n 3.92313e-19 $X=1.57 $Y=0.74 $X2=0 $Y2=0
cc_122 N_A_62_94#_M1003_g N_Y_c_402_n 4.14962e-19 $X=1.14 $Y=0.74 $X2=0 $Y2=0
cc_123 N_A_62_94#_c_113_n N_Y_c_402_n 0.00101398f $X=1.645 $Y=1.69 $X2=0 $Y2=0
cc_124 N_A_62_94#_c_117_n N_Y_c_402_n 0.0131103f $X=0.89 $Y=1.65 $X2=0 $Y2=0
cc_125 N_A_62_94#_c_118_n N_Y_c_403_n 0.0120829f $X=1.555 $Y=1.765 $X2=0 $Y2=0
cc_126 N_A_62_94#_c_112_n N_Y_c_403_n 0.0149807f $X=1.93 $Y=1.69 $X2=0 $Y2=0
cc_127 N_A_62_94#_c_113_n N_Y_c_403_n 0.0107456f $X=1.645 $Y=1.69 $X2=0 $Y2=0
cc_128 N_A_62_94#_c_121_n N_Y_c_403_n 0.0107007f $X=2.005 $Y=1.765 $X2=0 $Y2=0
cc_129 N_A_62_94#_c_117_n N_Y_c_403_n 0.0153964f $X=0.89 $Y=1.65 $X2=0 $Y2=0
cc_130 N_A_62_94#_c_124_n N_Y_c_403_n 0.00462354f $X=0.81 $Y=1.94 $X2=0 $Y2=0
cc_131 N_A_62_94#_M1009_g N_Y_c_406_n 0.0126976f $X=1.57 $Y=0.74 $X2=0 $Y2=0
cc_132 N_A_62_94#_M1003_g N_Y_c_407_n 5.22898e-19 $X=1.14 $Y=0.74 $X2=0 $Y2=0
cc_133 N_A_62_94#_M1009_g N_Y_c_407_n 0.0124603f $X=1.57 $Y=0.74 $X2=0 $Y2=0
cc_134 N_A_62_94#_c_112_n N_Y_c_407_n 0.00782278f $X=1.93 $Y=1.69 $X2=0 $Y2=0
cc_135 N_A_62_94#_c_113_n N_Y_c_407_n 0.00363407f $X=1.645 $Y=1.69 $X2=0 $Y2=0
cc_136 N_A_62_94#_c_117_n N_Y_c_407_n 0.0113438f $X=0.89 $Y=1.65 $X2=0 $Y2=0
cc_137 N_A_62_94#_c_117_n N_VGND_M1002_d 0.00188126f $X=0.89 $Y=1.65 $X2=-0.19
+ $Y2=-0.245
cc_138 N_A_62_94#_M1003_g N_VGND_c_458_n 0.0113786f $X=1.14 $Y=0.74 $X2=0 $Y2=0
cc_139 N_A_62_94#_M1009_g N_VGND_c_458_n 5.01478e-19 $X=1.57 $Y=0.74 $X2=0 $Y2=0
cc_140 N_A_62_94#_c_114_n N_VGND_c_458_n 0.00121634f $X=0.435 $Y=0.615 $X2=0
+ $Y2=0
cc_141 N_A_62_94#_c_115_n N_VGND_c_458_n 0.00265802f $X=0.805 $Y=1.195 $X2=0
+ $Y2=0
cc_142 N_A_62_94#_c_117_n N_VGND_c_458_n 0.0192874f $X=0.89 $Y=1.65 $X2=0 $Y2=0
cc_143 N_A_62_94#_M1003_g N_VGND_c_459_n 0.00383152f $X=1.14 $Y=0.74 $X2=0 $Y2=0
cc_144 N_A_62_94#_M1009_g N_VGND_c_459_n 0.00383152f $X=1.57 $Y=0.74 $X2=0 $Y2=0
cc_145 N_A_62_94#_M1003_g N_VGND_c_460_n 4.62684e-19 $X=1.14 $Y=0.74 $X2=0 $Y2=0
cc_146 N_A_62_94#_M1009_g N_VGND_c_460_n 0.0117356f $X=1.57 $Y=0.74 $X2=0 $Y2=0
cc_147 N_A_62_94#_c_114_n N_VGND_c_462_n 0.00787252f $X=0.435 $Y=0.615 $X2=0
+ $Y2=0
cc_148 N_A_62_94#_M1003_g N_VGND_c_466_n 0.0075754f $X=1.14 $Y=0.74 $X2=0 $Y2=0
cc_149 N_A_62_94#_M1009_g N_VGND_c_466_n 0.0075754f $X=1.57 $Y=0.74 $X2=0 $Y2=0
cc_150 N_A_62_94#_c_114_n N_VGND_c_466_n 0.0085887f $X=0.435 $Y=0.615 $X2=0
+ $Y2=0
cc_151 N_A_62_94#_M1009_g N_A_436_74#_c_517_n 6.92543e-19 $X=1.57 $Y=0.74 $X2=0
+ $Y2=0
cc_152 N_A1_c_193_n N_A2_c_250_n 0.00908185f $X=2.905 $Y=1.765 $X2=-0.19
+ $Y2=-0.245
cc_153 N_A1_M1011_g N_A2_c_246_n 0.0123753f $X=2.95 $Y=0.74 $X2=0 $Y2=0
cc_154 N_A1_M1011_g A2 0.00134497f $X=2.95 $Y=0.74 $X2=0 $Y2=0
cc_155 N_A1_c_190_n A2 0.00804954f $X=2.65 $Y=1.485 $X2=0 $Y2=0
cc_156 N_A1_c_191_n A2 3.7708e-19 $X=2.905 $Y=1.542 $X2=0 $Y2=0
cc_157 N_A1_M1011_g N_A2_c_249_n 0.0135068f $X=2.95 $Y=0.74 $X2=0 $Y2=0
cc_158 N_A1_c_190_n N_A2_c_249_n 6.70895e-19 $X=2.65 $Y=1.485 $X2=0 $Y2=0
cc_159 N_A1_c_191_n N_A2_c_249_n 0.0147294f $X=2.905 $Y=1.542 $X2=0 $Y2=0
cc_160 N_A1_c_192_n N_VPWR_c_290_n 0.0109842f $X=2.455 $Y=1.765 $X2=0 $Y2=0
cc_161 N_A1_c_193_n N_VPWR_c_290_n 0.0116643f $X=2.905 $Y=1.765 $X2=0 $Y2=0
cc_162 N_A1_c_193_n N_VPWR_c_291_n 5.87505e-19 $X=2.905 $Y=1.765 $X2=0 $Y2=0
cc_163 N_A1_c_192_n N_VPWR_c_292_n 0.00413917f $X=2.455 $Y=1.765 $X2=0 $Y2=0
cc_164 N_A1_c_193_n N_VPWR_c_293_n 0.00413917f $X=2.905 $Y=1.765 $X2=0 $Y2=0
cc_165 N_A1_c_192_n N_VPWR_c_287_n 0.0081781f $X=2.455 $Y=1.765 $X2=0 $Y2=0
cc_166 N_A1_c_193_n N_VPWR_c_287_n 0.0081781f $X=2.905 $Y=1.765 $X2=0 $Y2=0
cc_167 N_A1_c_192_n N_A_241_368#_c_342_n 0.00125031f $X=2.455 $Y=1.765 $X2=0
+ $Y2=0
cc_168 N_A1_c_192_n N_A_241_368#_c_344_n 0.00272065f $X=2.455 $Y=1.765 $X2=0
+ $Y2=0
cc_169 N_A1_c_192_n N_A_241_368#_c_360_n 0.00564091f $X=2.455 $Y=1.765 $X2=0
+ $Y2=0
cc_170 N_A1_c_192_n N_A_241_368#_c_361_n 0.0157383f $X=2.455 $Y=1.765 $X2=0
+ $Y2=0
cc_171 N_A1_c_193_n N_A_241_368#_c_361_n 0.0171849f $X=2.905 $Y=1.765 $X2=0
+ $Y2=0
cc_172 N_A1_c_190_n N_A_241_368#_c_361_n 0.0225224f $X=2.65 $Y=1.485 $X2=0 $Y2=0
cc_173 N_A1_c_191_n N_A_241_368#_c_361_n 0.00121734f $X=2.905 $Y=1.542 $X2=0
+ $Y2=0
cc_174 N_A1_c_193_n N_A_241_368#_c_348_n 0.00949056f $X=2.905 $Y=1.765 $X2=0
+ $Y2=0
cc_175 N_A1_c_190_n N_A_241_368#_c_348_n 0.00384606f $X=2.65 $Y=1.485 $X2=0
+ $Y2=0
cc_176 N_A1_c_191_n N_A_241_368#_c_348_n 3.5928e-19 $X=2.905 $Y=1.542 $X2=0
+ $Y2=0
cc_177 N_A1_c_192_n N_Y_c_403_n 2.64799e-19 $X=2.455 $Y=1.765 $X2=0 $Y2=0
cc_178 N_A1_c_190_n N_Y_c_403_n 0.011574f $X=2.65 $Y=1.485 $X2=0 $Y2=0
cc_179 N_A1_c_191_n N_Y_c_403_n 0.00273312f $X=2.905 $Y=1.542 $X2=0 $Y2=0
cc_180 N_A1_M1000_g N_Y_c_404_n 0.0126181f $X=2.52 $Y=0.74 $X2=0 $Y2=0
cc_181 N_A1_c_190_n N_Y_c_404_n 0.00619439f $X=2.65 $Y=1.485 $X2=0 $Y2=0
cc_182 N_A1_c_191_n N_Y_c_404_n 0.00328281f $X=2.905 $Y=1.542 $X2=0 $Y2=0
cc_183 N_A1_M1000_g N_Y_c_405_n 0.0103649f $X=2.52 $Y=0.74 $X2=0 $Y2=0
cc_184 N_A1_M1011_g N_Y_c_405_n 0.00672659f $X=2.95 $Y=0.74 $X2=0 $Y2=0
cc_185 N_A1_c_190_n N_Y_c_405_n 0.0200194f $X=2.65 $Y=1.485 $X2=0 $Y2=0
cc_186 N_A1_c_191_n N_Y_c_405_n 7.50363e-19 $X=2.905 $Y=1.542 $X2=0 $Y2=0
cc_187 N_A1_M1000_g N_Y_c_407_n 0.00689063f $X=2.52 $Y=0.74 $X2=0 $Y2=0
cc_188 N_A1_c_190_n N_Y_c_407_n 0.00638885f $X=2.65 $Y=1.485 $X2=0 $Y2=0
cc_189 N_A1_c_191_n N_Y_c_407_n 0.00143746f $X=2.905 $Y=1.542 $X2=0 $Y2=0
cc_190 N_A1_M1000_g N_VGND_c_460_n 0.00714008f $X=2.52 $Y=0.74 $X2=0 $Y2=0
cc_191 N_A1_M1011_g N_VGND_c_461_n 6.35276e-19 $X=2.95 $Y=0.74 $X2=0 $Y2=0
cc_192 N_A1_M1000_g N_VGND_c_464_n 0.00291649f $X=2.52 $Y=0.74 $X2=0 $Y2=0
cc_193 N_A1_M1011_g N_VGND_c_464_n 0.00291649f $X=2.95 $Y=0.74 $X2=0 $Y2=0
cc_194 N_A1_M1000_g N_VGND_c_466_n 0.0036412f $X=2.52 $Y=0.74 $X2=0 $Y2=0
cc_195 N_A1_M1011_g N_VGND_c_466_n 0.00359219f $X=2.95 $Y=0.74 $X2=0 $Y2=0
cc_196 N_A1_M1000_g N_A_436_74#_c_517_n 0.01124f $X=2.52 $Y=0.74 $X2=0 $Y2=0
cc_197 N_A1_M1011_g N_A_436_74#_c_517_n 0.0142063f $X=2.95 $Y=0.74 $X2=0 $Y2=0
cc_198 N_A2_c_250_n N_VPWR_c_290_n 5.35985e-19 $X=3.355 $Y=1.765 $X2=0 $Y2=0
cc_199 N_A2_c_250_n N_VPWR_c_291_n 0.013448f $X=3.355 $Y=1.765 $X2=0 $Y2=0
cc_200 N_A2_c_251_n N_VPWR_c_291_n 0.0166899f $X=3.825 $Y=1.765 $X2=0 $Y2=0
cc_201 N_A2_c_250_n N_VPWR_c_293_n 0.00413917f $X=3.355 $Y=1.765 $X2=0 $Y2=0
cc_202 N_A2_c_251_n N_VPWR_c_294_n 0.00413917f $X=3.825 $Y=1.765 $X2=0 $Y2=0
cc_203 N_A2_c_250_n N_VPWR_c_287_n 0.0081781f $X=3.355 $Y=1.765 $X2=0 $Y2=0
cc_204 N_A2_c_251_n N_VPWR_c_287_n 0.00821187f $X=3.825 $Y=1.765 $X2=0 $Y2=0
cc_205 N_A2_c_250_n N_A_241_368#_c_346_n 0.00993732f $X=3.355 $Y=1.765 $X2=0
+ $Y2=0
cc_206 N_A2_c_251_n N_A_241_368#_c_346_n 0.0109805f $X=3.825 $Y=1.765 $X2=0
+ $Y2=0
cc_207 A2 N_A_241_368#_c_346_n 0.0334689f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_208 N_A2_c_249_n N_A_241_368#_c_346_n 0.0157657f $X=3.81 $Y=1.492 $X2=0 $Y2=0
cc_209 N_A2_c_251_n N_A_241_368#_c_347_n 0.00808878f $X=3.825 $Y=1.765 $X2=0
+ $Y2=0
cc_210 N_A2_c_250_n N_A_241_368#_c_348_n 0.00667324f $X=3.355 $Y=1.765 $X2=0
+ $Y2=0
cc_211 N_A2_c_246_n N_Y_c_405_n 4.34981e-19 $X=3.38 $Y=1.22 $X2=0 $Y2=0
cc_212 N_A2_c_246_n N_VGND_c_461_n 0.00768902f $X=3.38 $Y=1.22 $X2=0 $Y2=0
cc_213 N_A2_c_247_n N_VGND_c_461_n 0.010528f $X=3.81 $Y=1.22 $X2=0 $Y2=0
cc_214 N_A2_c_246_n N_VGND_c_464_n 0.00383152f $X=3.38 $Y=1.22 $X2=0 $Y2=0
cc_215 N_A2_c_247_n N_VGND_c_465_n 0.00383152f $X=3.81 $Y=1.22 $X2=0 $Y2=0
cc_216 N_A2_c_246_n N_VGND_c_466_n 0.00384065f $X=3.38 $Y=1.22 $X2=0 $Y2=0
cc_217 N_A2_c_247_n N_VGND_c_466_n 0.00387675f $X=3.81 $Y=1.22 $X2=0 $Y2=0
cc_218 N_A2_c_246_n N_A_436_74#_c_524_n 0.00985057f $X=3.38 $Y=1.22 $X2=0 $Y2=0
cc_219 N_A2_c_247_n N_A_436_74#_c_524_n 0.0141214f $X=3.81 $Y=1.22 $X2=0 $Y2=0
cc_220 A2 N_A_436_74#_c_524_n 0.0271317f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_221 N_A2_c_249_n N_A_436_74#_c_524_n 6.30401e-19 $X=3.81 $Y=1.492 $X2=0 $Y2=0
cc_222 N_A2_c_247_n N_A_436_74#_c_519_n 7.92899e-19 $X=3.81 $Y=1.22 $X2=0 $Y2=0
cc_223 N_A2_c_247_n N_A_436_74#_c_520_n 0.00159319f $X=3.81 $Y=1.22 $X2=0 $Y2=0
cc_224 N_VPWR_c_290_n N_A_241_368#_c_342_n 0.0125885f $X=2.68 $Y=2.375 $X2=0
+ $Y2=0
cc_225 N_VPWR_c_292_n N_A_241_368#_c_342_n 0.0584986f $X=2.515 $Y=3.33 $X2=0
+ $Y2=0
cc_226 N_VPWR_c_287_n N_A_241_368#_c_342_n 0.0327208f $X=4.08 $Y=3.33 $X2=0
+ $Y2=0
cc_227 N_VPWR_c_292_n N_A_241_368#_c_343_n 0.0179217f $X=2.515 $Y=3.33 $X2=0
+ $Y2=0
cc_228 N_VPWR_c_287_n N_A_241_368#_c_343_n 0.00971942f $X=4.08 $Y=3.33 $X2=0
+ $Y2=0
cc_229 N_VPWR_c_290_n N_A_241_368#_c_360_n 0.0405146f $X=2.68 $Y=2.375 $X2=0
+ $Y2=0
cc_230 N_VPWR_M1007_d N_A_241_368#_c_361_n 0.00360966f $X=2.53 $Y=1.84 $X2=0
+ $Y2=0
cc_231 N_VPWR_c_290_n N_A_241_368#_c_361_n 0.0171813f $X=2.68 $Y=2.375 $X2=0
+ $Y2=0
cc_232 N_VPWR_c_290_n N_A_241_368#_c_345_n 0.0449718f $X=2.68 $Y=2.375 $X2=0
+ $Y2=0
cc_233 N_VPWR_c_293_n N_A_241_368#_c_345_n 0.00749631f $X=3.415 $Y=3.33 $X2=0
+ $Y2=0
cc_234 N_VPWR_c_287_n N_A_241_368#_c_345_n 0.0062048f $X=4.08 $Y=3.33 $X2=0
+ $Y2=0
cc_235 N_VPWR_M1001_s N_A_241_368#_c_346_n 0.00218982f $X=3.43 $Y=1.84 $X2=0
+ $Y2=0
cc_236 N_VPWR_c_291_n N_A_241_368#_c_346_n 0.0188085f $X=3.59 $Y=2.145 $X2=0
+ $Y2=0
cc_237 N_VPWR_c_291_n N_A_241_368#_c_347_n 0.0619908f $X=3.59 $Y=2.145 $X2=0
+ $Y2=0
cc_238 N_VPWR_c_294_n N_A_241_368#_c_347_n 0.011066f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_239 N_VPWR_c_287_n N_A_241_368#_c_347_n 0.00915947f $X=4.08 $Y=3.33 $X2=0
+ $Y2=0
cc_240 N_VPWR_c_291_n N_A_241_368#_c_348_n 0.0601953f $X=3.59 $Y=2.145 $X2=0
+ $Y2=0
cc_241 N_A_241_368#_c_342_n N_Y_M1005_d 0.00197722f $X=2.115 $Y=2.99 $X2=0 $Y2=0
cc_242 N_A_241_368#_c_341_n N_Y_c_402_n 6.70242e-19 $X=1.33 $Y=1.985 $X2=0 $Y2=0
cc_243 N_A_241_368#_c_341_n N_Y_c_403_n 0.0613813f $X=1.33 $Y=1.985 $X2=0 $Y2=0
cc_244 N_A_241_368#_c_342_n N_Y_c_403_n 0.0160777f $X=2.115 $Y=2.99 $X2=0 $Y2=0
cc_245 N_A_241_368#_c_344_n N_Y_c_403_n 0.0120471f $X=2.215 $Y=2.12 $X2=0 $Y2=0
cc_246 N_A_241_368#_c_344_n N_Y_c_404_n 0.00127772f $X=2.215 $Y=2.12 $X2=0 $Y2=0
cc_247 N_A_241_368#_c_344_n N_Y_c_407_n 0.00783425f $X=2.215 $Y=2.12 $X2=0 $Y2=0
cc_248 N_A_241_368#_c_346_n N_A_436_74#_c_530_n 0.00103389f $X=3.965 $Y=1.805
+ $X2=0 $Y2=0
cc_249 N_A_241_368#_c_348_n N_A_436_74#_c_530_n 0.00450741f $X=3.13 $Y=1.805
+ $X2=0 $Y2=0
cc_250 N_A_241_368#_c_346_n N_A_436_74#_c_519_n 0.00969915f $X=3.965 $Y=1.805
+ $X2=0 $Y2=0
cc_251 N_Y_c_407_n N_VGND_M1009_s 0.00288199f $X=2.275 $Y=1.195 $X2=0 $Y2=0
cc_252 N_Y_c_401_n N_VGND_c_458_n 0.0218329f $X=1.355 $Y=0.515 $X2=0 $Y2=0
cc_253 N_Y_c_401_n N_VGND_c_459_n 0.00749631f $X=1.355 $Y=0.515 $X2=0 $Y2=0
cc_254 N_Y_c_401_n N_VGND_c_460_n 0.0171736f $X=1.355 $Y=0.515 $X2=0 $Y2=0
cc_255 N_Y_c_405_n N_VGND_c_460_n 0.0011882f $X=2.735 $Y=0.91 $X2=0 $Y2=0
cc_256 N_Y_c_407_n N_VGND_c_460_n 0.023479f $X=2.275 $Y=1.195 $X2=0 $Y2=0
cc_257 N_Y_c_401_n N_VGND_c_466_n 0.0062048f $X=1.355 $Y=0.515 $X2=0 $Y2=0
cc_258 N_Y_c_404_n N_A_436_74#_M1000_d 0.00174919f $X=2.57 $Y=1.065 $X2=-0.19
+ $Y2=-0.245
cc_259 N_Y_c_407_n N_A_436_74#_M1000_d 0.00213669f $X=2.275 $Y=1.195 $X2=-0.19
+ $Y2=-0.245
cc_260 N_Y_M1000_s N_A_436_74#_c_517_n 0.00178571f $X=2.595 $Y=0.37 $X2=0 $Y2=0
cc_261 N_Y_c_405_n N_A_436_74#_c_517_n 0.0162079f $X=2.735 $Y=0.91 $X2=0 $Y2=0
cc_262 N_Y_c_407_n N_A_436_74#_c_517_n 0.0153378f $X=2.275 $Y=1.195 $X2=0 $Y2=0
cc_263 N_VGND_c_460_n N_A_436_74#_c_517_n 0.0202776f $X=1.785 $Y=0.645 $X2=0
+ $Y2=0
cc_264 N_VGND_c_464_n N_A_436_74#_c_517_n 0.038121f $X=3.43 $Y=0 $X2=0 $Y2=0
cc_265 N_VGND_c_466_n N_A_436_74#_c_517_n 0.0321651f $X=4.08 $Y=0 $X2=0 $Y2=0
cc_266 N_VGND_c_461_n N_A_436_74#_c_518_n 0.00985092f $X=3.595 $Y=0.55 $X2=0
+ $Y2=0
cc_267 N_VGND_c_464_n N_A_436_74#_c_518_n 0.00760167f $X=3.43 $Y=0 $X2=0 $Y2=0
cc_268 N_VGND_c_466_n N_A_436_74#_c_518_n 0.00628491f $X=4.08 $Y=0 $X2=0 $Y2=0
cc_269 N_VGND_M1004_d N_A_436_74#_c_524_n 0.00328934f $X=3.455 $Y=0.37 $X2=0
+ $Y2=0
cc_270 N_VGND_c_461_n N_A_436_74#_c_524_n 0.0167019f $X=3.595 $Y=0.55 $X2=0
+ $Y2=0
cc_271 N_VGND_c_466_n N_A_436_74#_c_524_n 0.0116543f $X=4.08 $Y=0 $X2=0 $Y2=0
cc_272 N_VGND_c_461_n N_A_436_74#_c_520_n 0.0121972f $X=3.595 $Y=0.55 $X2=0
+ $Y2=0
cc_273 N_VGND_c_465_n N_A_436_74#_c_520_n 0.011066f $X=4.08 $Y=0 $X2=0 $Y2=0
cc_274 N_VGND_c_466_n N_A_436_74#_c_520_n 0.00915947f $X=4.08 $Y=0 $X2=0 $Y2=0
