* File: sky130_fd_sc_hs__a21oi_1.pxi.spice
* Created: Thu Aug 27 20:25:09 2020
* 
x_PM_SKY130_FD_SC_HS__A21OI_1%A2 N_A2_c_36_n N_A2_M1001_g N_A2_c_37_n
+ N_A2_M1005_g A2 PM_SKY130_FD_SC_HS__A21OI_1%A2
x_PM_SKY130_FD_SC_HS__A21OI_1%A1 N_A1_M1002_g N_A1_c_59_n N_A1_M1004_g A1
+ N_A1_c_60_n PM_SKY130_FD_SC_HS__A21OI_1%A1
x_PM_SKY130_FD_SC_HS__A21OI_1%B1 N_B1_c_91_n N_B1_M1003_g N_B1_c_92_n
+ N_B1_M1000_g B1 PM_SKY130_FD_SC_HS__A21OI_1%B1
x_PM_SKY130_FD_SC_HS__A21OI_1%A_29_368# N_A_29_368#_M1001_s N_A_29_368#_M1004_d
+ N_A_29_368#_c_115_n N_A_29_368#_c_116_n N_A_29_368#_c_121_n
+ N_A_29_368#_c_117_n PM_SKY130_FD_SC_HS__A21OI_1%A_29_368#
x_PM_SKY130_FD_SC_HS__A21OI_1%VPWR N_VPWR_M1001_d N_VPWR_c_141_n VPWR
+ N_VPWR_c_142_n N_VPWR_c_143_n N_VPWR_c_140_n N_VPWR_c_145_n
+ PM_SKY130_FD_SC_HS__A21OI_1%VPWR
x_PM_SKY130_FD_SC_HS__A21OI_1%Y N_Y_M1002_d N_Y_M1000_d N_Y_c_165_n N_Y_c_166_n
+ N_Y_c_169_n N_Y_c_170_n N_Y_c_167_n Y Y Y PM_SKY130_FD_SC_HS__A21OI_1%Y
x_PM_SKY130_FD_SC_HS__A21OI_1%VGND N_VGND_M1005_s N_VGND_M1003_d N_VGND_c_201_n
+ N_VGND_c_202_n N_VGND_c_203_n N_VGND_c_204_n VGND N_VGND_c_205_n
+ N_VGND_c_206_n PM_SKY130_FD_SC_HS__A21OI_1%VGND
cc_1 VNB N_A2_c_36_n 0.0669347f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.765
cc_2 VNB N_A2_c_37_n 0.0204319f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=1.22
cc_3 VNB A2 0.00894107f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_4 VNB N_A1_M1002_g 0.0248365f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.4
cc_5 VNB N_A1_c_59_n 0.0236943f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=0.74
cc_6 VNB N_A1_c_60_n 0.00959608f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.295
cc_7 VNB N_B1_c_91_n 0.0209416f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.765
cc_8 VNB N_B1_c_92_n 0.0665189f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=1.22
cc_9 VNB B1 0.00662327f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_10 VNB N_VPWR_c_140_n 0.0840719f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_Y_c_165_n 0.00320135f $X=-0.19 $Y=-0.245 $X2=0.345 $Y2=1.385
cc_12 VNB N_Y_c_166_n 0.0035645f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.295
cc_13 VNB N_Y_c_167_n 0.00543429f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_VGND_c_201_n 0.0125057f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_15 VNB N_VGND_c_202_n 0.0350088f $X=-0.19 $Y=-0.245 $X2=0.345 $Y2=1.385
cc_16 VNB N_VGND_c_203_n 0.0107718f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.385
cc_17 VNB N_VGND_c_204_n 0.0358154f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_VGND_c_205_n 0.0319078f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_VGND_c_206_n 0.146074f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VPB N_A2_c_36_n 0.0309207f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.765
cc_21 VPB N_A1_c_59_n 0.0270859f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=0.74
cc_22 VPB N_A1_c_60_n 0.00422406f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.295
cc_23 VPB N_B1_c_92_n 0.027762f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=1.22
cc_24 VPB N_A_29_368#_c_115_n 0.0191639f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.21
cc_25 VPB N_A_29_368#_c_116_n 0.0314243f $X=-0.19 $Y=1.66 $X2=0.345 $Y2=1.385
cc_26 VPB N_A_29_368#_c_117_n 0.0025758f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_27 VPB N_VPWR_c_141_n 0.00981021f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=0.74
cc_28 VPB N_VPWR_c_142_n 0.0179929f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.385
cc_29 VPB N_VPWR_c_143_n 0.0303755f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_30 VPB N_VPWR_c_140_n 0.0551234f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_31 VPB N_VPWR_c_145_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_32 VPB N_Y_c_166_n 3.49014e-19 $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.295
cc_33 VPB N_Y_c_169_n 0.00934184f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_34 VPB N_Y_c_170_n 0.00104144f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_35 VPB Y 0.043203f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_36 N_A2_c_37_n N_A1_M1002_g 0.0428684f $X=0.51 $Y=1.22 $X2=0 $Y2=0
cc_37 A2 N_A1_M1002_g 6.23327e-19 $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_38 N_A2_c_36_n N_A1_c_59_n 0.0687299f $X=0.495 $Y=1.765 $X2=0 $Y2=0
cc_39 N_A2_c_36_n N_A1_c_60_n 0.00846493f $X=0.495 $Y=1.765 $X2=0 $Y2=0
cc_40 A2 N_A1_c_60_n 0.0162065f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_41 N_A2_c_36_n N_A_29_368#_c_115_n 0.00788863f $X=0.495 $Y=1.765 $X2=0 $Y2=0
cc_42 A2 N_A_29_368#_c_115_n 0.0196638f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_43 N_A2_c_36_n N_A_29_368#_c_116_n 9.60518e-19 $X=0.495 $Y=1.765 $X2=0 $Y2=0
cc_44 N_A2_c_36_n N_A_29_368#_c_121_n 0.0186687f $X=0.495 $Y=1.765 $X2=0 $Y2=0
cc_45 N_A2_c_36_n N_VPWR_c_141_n 0.00342349f $X=0.495 $Y=1.765 $X2=0 $Y2=0
cc_46 N_A2_c_36_n N_VPWR_c_142_n 0.00460063f $X=0.495 $Y=1.765 $X2=0 $Y2=0
cc_47 N_A2_c_36_n N_VPWR_c_140_n 0.00911302f $X=0.495 $Y=1.765 $X2=0 $Y2=0
cc_48 N_A2_c_37_n N_Y_c_165_n 0.0026419f $X=0.51 $Y=1.22 $X2=0 $Y2=0
cc_49 N_A2_c_36_n N_VGND_c_202_n 0.00199271f $X=0.495 $Y=1.765 $X2=0 $Y2=0
cc_50 N_A2_c_37_n N_VGND_c_202_n 0.0167319f $X=0.51 $Y=1.22 $X2=0 $Y2=0
cc_51 A2 N_VGND_c_202_n 0.024157f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_52 N_A2_c_37_n N_VGND_c_205_n 0.00383152f $X=0.51 $Y=1.22 $X2=0 $Y2=0
cc_53 N_A2_c_37_n N_VGND_c_206_n 0.0075694f $X=0.51 $Y=1.22 $X2=0 $Y2=0
cc_54 N_A1_M1002_g N_B1_c_91_n 0.0197297f $X=0.87 $Y=0.74 $X2=-0.19 $Y2=-0.245
cc_55 N_A1_c_59_n N_B1_c_92_n 0.0472655f $X=0.975 $Y=1.765 $X2=0 $Y2=0
cc_56 N_A1_c_60_n N_B1_c_92_n 3.93518e-19 $X=0.96 $Y=1.515 $X2=0 $Y2=0
cc_57 N_A1_c_59_n N_A_29_368#_c_115_n 7.74545e-19 $X=0.975 $Y=1.765 $X2=0 $Y2=0
cc_58 N_A1_c_59_n N_A_29_368#_c_121_n 2.05924e-19 $X=0.975 $Y=1.765 $X2=0 $Y2=0
cc_59 N_A1_c_60_n N_A_29_368#_c_121_n 0.0155105f $X=0.96 $Y=1.515 $X2=0 $Y2=0
cc_60 N_A1_c_59_n N_A_29_368#_c_117_n 0.0190842f $X=0.975 $Y=1.765 $X2=0 $Y2=0
cc_61 N_A1_c_60_n N_A_29_368#_c_117_n 0.0111003f $X=0.96 $Y=1.515 $X2=0 $Y2=0
cc_62 N_A1_c_59_n N_VPWR_c_141_n 0.00342349f $X=0.975 $Y=1.765 $X2=0 $Y2=0
cc_63 N_A1_c_59_n N_VPWR_c_143_n 0.00460063f $X=0.975 $Y=1.765 $X2=0 $Y2=0
cc_64 N_A1_c_59_n N_VPWR_c_140_n 0.00907925f $X=0.975 $Y=1.765 $X2=0 $Y2=0
cc_65 N_A1_M1002_g N_Y_c_165_n 0.0117918f $X=0.87 $Y=0.74 $X2=0 $Y2=0
cc_66 N_A1_M1002_g N_Y_c_166_n 0.00323848f $X=0.87 $Y=0.74 $X2=0 $Y2=0
cc_67 N_A1_c_59_n N_Y_c_166_n 0.00226362f $X=0.975 $Y=1.765 $X2=0 $Y2=0
cc_68 N_A1_c_60_n N_Y_c_166_n 0.0284774f $X=0.96 $Y=1.515 $X2=0 $Y2=0
cc_69 N_A1_c_59_n N_Y_c_170_n 0.00331133f $X=0.975 $Y=1.765 $X2=0 $Y2=0
cc_70 N_A1_c_60_n N_Y_c_170_n 0.00500939f $X=0.96 $Y=1.515 $X2=0 $Y2=0
cc_71 N_A1_M1002_g N_Y_c_167_n 0.00444011f $X=0.87 $Y=0.74 $X2=0 $Y2=0
cc_72 N_A1_c_59_n N_Y_c_167_n 0.00620958f $X=0.975 $Y=1.765 $X2=0 $Y2=0
cc_73 N_A1_c_60_n N_Y_c_167_n 0.0109718f $X=0.96 $Y=1.515 $X2=0 $Y2=0
cc_74 N_A1_M1002_g N_VGND_c_202_n 0.00236525f $X=0.87 $Y=0.74 $X2=0 $Y2=0
cc_75 N_A1_M1002_g N_VGND_c_205_n 0.00434272f $X=0.87 $Y=0.74 $X2=0 $Y2=0
cc_76 N_A1_M1002_g N_VGND_c_206_n 0.00821699f $X=0.87 $Y=0.74 $X2=0 $Y2=0
cc_77 N_B1_c_92_n N_A_29_368#_c_117_n 0.012717f $X=1.425 $Y=1.765 $X2=0 $Y2=0
cc_78 N_B1_c_92_n N_VPWR_c_143_n 0.00445602f $X=1.425 $Y=1.765 $X2=0 $Y2=0
cc_79 N_B1_c_92_n N_VPWR_c_140_n 0.00861895f $X=1.425 $Y=1.765 $X2=0 $Y2=0
cc_80 N_B1_c_91_n N_Y_c_165_n 0.0038671f $X=1.41 $Y=1.22 $X2=0 $Y2=0
cc_81 N_B1_c_91_n N_Y_c_166_n 0.00108982f $X=1.41 $Y=1.22 $X2=0 $Y2=0
cc_82 N_B1_c_92_n N_Y_c_166_n 0.0164374f $X=1.425 $Y=1.765 $X2=0 $Y2=0
cc_83 B1 N_Y_c_166_n 0.0252697f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_84 N_B1_c_92_n N_Y_c_169_n 0.0182813f $X=1.425 $Y=1.765 $X2=0 $Y2=0
cc_85 B1 N_Y_c_169_n 0.0212273f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_86 N_B1_c_92_n N_Y_c_170_n 0.00366405f $X=1.425 $Y=1.765 $X2=0 $Y2=0
cc_87 N_B1_c_91_n N_Y_c_167_n 0.0131024f $X=1.41 $Y=1.22 $X2=0 $Y2=0
cc_88 N_B1_c_92_n Y 0.00715325f $X=1.425 $Y=1.765 $X2=0 $Y2=0
cc_89 N_B1_c_91_n N_VGND_c_204_n 0.0075574f $X=1.41 $Y=1.22 $X2=0 $Y2=0
cc_90 N_B1_c_92_n N_VGND_c_204_n 0.00166151f $X=1.425 $Y=1.765 $X2=0 $Y2=0
cc_91 B1 N_VGND_c_204_n 0.0200189f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_92 N_B1_c_91_n N_VGND_c_205_n 0.00461464f $X=1.41 $Y=1.22 $X2=0 $Y2=0
cc_93 N_B1_c_91_n N_VGND_c_206_n 0.00913518f $X=1.41 $Y=1.22 $X2=0 $Y2=0
cc_94 N_A_29_368#_c_121_n N_VPWR_M1001_d 0.00452124f $X=0.833 $Y=2.107 $X2=-0.19
+ $Y2=1.66
cc_95 N_A_29_368#_c_117_n N_VPWR_M1001_d 2.02994e-19 $X=1.2 $Y=2.225 $X2=-0.19
+ $Y2=1.66
cc_96 N_A_29_368#_c_116_n N_VPWR_c_141_n 0.0248659f $X=0.27 $Y=2.4 $X2=0 $Y2=0
cc_97 N_A_29_368#_c_121_n N_VPWR_c_141_n 0.0171441f $X=0.833 $Y=2.107 $X2=0
+ $Y2=0
cc_98 N_A_29_368#_c_117_n N_VPWR_c_141_n 0.0257042f $X=1.2 $Y=2.225 $X2=0 $Y2=0
cc_99 N_A_29_368#_c_116_n N_VPWR_c_142_n 0.0130739f $X=0.27 $Y=2.4 $X2=0 $Y2=0
cc_100 N_A_29_368#_c_117_n N_VPWR_c_143_n 0.0130321f $X=1.2 $Y=2.225 $X2=0 $Y2=0
cc_101 N_A_29_368#_c_116_n N_VPWR_c_140_n 0.0108215f $X=0.27 $Y=2.4 $X2=0 $Y2=0
cc_102 N_A_29_368#_c_117_n N_VPWR_c_140_n 0.0107539f $X=1.2 $Y=2.225 $X2=0 $Y2=0
cc_103 N_A_29_368#_M1004_d N_Y_c_170_n 0.00148214f $X=1.05 $Y=1.84 $X2=0 $Y2=0
cc_104 N_A_29_368#_c_117_n N_Y_c_170_n 0.00780925f $X=1.2 $Y=2.225 $X2=0 $Y2=0
cc_105 N_A_29_368#_c_117_n Y 0.0641597f $X=1.2 $Y=2.225 $X2=0 $Y2=0
cc_106 N_VPWR_c_143_n Y 0.011066f $X=1.68 $Y=3.33 $X2=0 $Y2=0
cc_107 N_VPWR_c_140_n Y 0.00915947f $X=1.68 $Y=3.33 $X2=0 $Y2=0
cc_108 N_Y_c_165_n N_VGND_c_202_n 0.0222599f $X=1.105 $Y=0.515 $X2=0 $Y2=0
cc_109 N_Y_c_165_n N_VGND_c_204_n 0.0184459f $X=1.105 $Y=0.515 $X2=0 $Y2=0
cc_110 N_Y_c_167_n N_VGND_c_204_n 7.76044e-19 $X=1.155 $Y=1.18 $X2=0 $Y2=0
cc_111 N_Y_c_165_n N_VGND_c_205_n 0.0163488f $X=1.105 $Y=0.515 $X2=0 $Y2=0
cc_112 N_Y_c_165_n N_VGND_c_206_n 0.0134757f $X=1.105 $Y=0.515 $X2=0 $Y2=0
