* NGSPICE file created from sky130_fd_sc_hs__nand4bb_4.ext - technology: sky130A

.subckt sky130_fd_sc_hs__nand4bb_4 A_N B_N C D VGND VNB VPB VPWR Y
M1000 a_374_74# a_27_114# Y VNB nlowvt w=740000u l=150000u
+  ad=1.0508e+12p pd=1.024e+07u as=4.921e+11p ps=4.29e+06u
M1001 Y a_232_114# VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=2.744e+12p pd=2.282e+07u as=3.9592e+12p ps=3.104e+07u
M1002 a_828_74# a_232_114# a_374_74# VNB nlowvt w=740000u l=150000u
+  ad=9.53e+11p pd=8.52e+06u as=0p ps=0u
M1003 a_1229_74# D VGND VNB nlowvt w=740000u l=150000u
+  ad=1.0434e+12p pd=1.022e+07u as=9.049e+11p ps=7.36e+06u
M1004 VPWR a_232_114# Y VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_374_74# a_27_114# Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 Y C VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_374_74# a_232_114# a_828_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VGND D a_1229_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 Y C VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 Y D VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 Y a_27_114# a_374_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VPWR C Y VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VGND D a_1229_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 VPWR C Y VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VPWR D Y VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 Y D VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_828_74# a_232_114# a_374_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 VPWR D Y VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VGND A_N a_27_114# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1020 Y a_27_114# VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 VPWR a_27_114# Y VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_232_114# B_N VGND VNB nlowvt w=740000u l=150000u
+  ad=2.368e+11p pd=2.12e+06u as=0p ps=0u
M1023 a_828_74# C a_1229_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 a_828_74# C a_1229_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 a_27_114# A_N VPWR VPB pshort w=840000u l=150000u
+  ad=2.52e+11p pd=2.28e+06u as=0p ps=0u
M1026 VPWR A_N a_27_114# VPB pshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 Y a_27_114# VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1028 a_374_74# a_232_114# a_828_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1029 a_232_114# B_N VPWR VPB pshort w=840000u l=150000u
+  ad=2.52e+11p pd=2.28e+06u as=0p ps=0u
M1030 VPWR a_27_114# Y VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1031 Y a_27_114# a_374_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1032 VPWR B_N a_232_114# VPB pshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1033 Y a_232_114# VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1034 a_1229_74# D VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1035 VPWR a_232_114# Y VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1036 a_1229_74# C a_828_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1037 a_1229_74# C a_828_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

