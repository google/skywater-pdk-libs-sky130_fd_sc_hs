* File: sky130_fd_sc_hs__a2111oi_2.pex.spice
* Created: Thu Aug 27 20:23:00 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HS__A2111OI_2%D1 1 3 6 8 10 11 12 18
c39 18 0 5.54777e-20 $X=1.13 $Y=1.515
c40 12 0 5.55949e-20 $X=1.2 $Y=1.665
c41 8 0 4.66136e-20 $X=1.145 $Y=1.765
r42 18 20 1.93316 $w=3.74e-07 $l=1.5e-08 $layer=POLY_cond $X=1.13 $Y=1.557
+ $X2=1.145 $Y2=1.557
r43 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.13
+ $Y=1.515 $X2=1.13 $Y2=1.515
r44 16 18 11.5989 $w=3.74e-07 $l=9e-08 $layer=POLY_cond $X=1.04 $Y=1.557
+ $X2=1.13 $Y2=1.557
r45 15 16 44.4626 $w=3.74e-07 $l=3.45e-07 $layer=POLY_cond $X=0.695 $Y=1.557
+ $X2=1.04 $Y2=1.557
r46 12 19 1.87607 $w=4.28e-07 $l=7e-08 $layer=LI1_cond $X=1.2 $Y=1.565 $X2=1.13
+ $Y2=1.565
r47 11 19 10.9884 $w=4.28e-07 $l=4.1e-07 $layer=LI1_cond $X=0.72 $Y=1.565
+ $X2=1.13 $Y2=1.565
r48 8 20 24.2268 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=1.145 $Y=1.765
+ $X2=1.145 $Y2=1.557
r49 8 10 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.145 $Y=1.765
+ $X2=1.145 $Y2=2.4
r50 4 16 24.2268 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.04 $Y=1.35
+ $X2=1.04 $Y2=1.557
r51 4 6 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.04 $Y=1.35 $X2=1.04
+ $Y2=0.74
r52 1 15 24.2268 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=0.695 $Y=1.765
+ $X2=0.695 $Y2=1.557
r53 1 3 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.695 $Y=1.765
+ $X2=0.695 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_HS__A2111OI_2%C1 3 5 7 8 10 11 12 13 20
c43 13 0 4.66136e-20 $X=2.64 $Y=1.665
c44 5 0 5.55949e-20 $X=1.595 $Y=1.765
c45 3 0 7.82037e-20 $X=1.58 $Y=0.74
r46 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.67
+ $Y=1.515 $X2=1.67 $Y2=1.515
r47 18 20 12.4655 $w=2.9e-07 $l=7.5e-08 $layer=POLY_cond $X=1.595 $Y=1.557
+ $X2=1.67 $Y2=1.557
r48 17 18 2.4931 $w=2.9e-07 $l=1.5e-08 $layer=POLY_cond $X=1.58 $Y=1.557
+ $X2=1.595 $Y2=1.557
r49 12 13 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=2.16 $Y=1.565
+ $X2=2.64 $Y2=1.565
r50 11 12 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=1.68 $Y=1.565
+ $X2=2.16 $Y2=1.565
r51 11 21 0.26801 $w=4.28e-07 $l=1e-08 $layer=LI1_cond $X=1.68 $Y=1.565 $X2=1.67
+ $Y2=1.565
r52 8 20 62.3276 $w=2.9e-07 $l=4.67574e-07 $layer=POLY_cond $X=2.045 $Y=1.765
+ $X2=1.67 $Y2=1.557
r53 8 10 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.045 $Y=1.765
+ $X2=2.045 $Y2=2.4
r54 5 18 18.1727 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=1.595 $Y=1.765
+ $X2=1.595 $Y2=1.557
r55 5 7 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.595 $Y=1.765
+ $X2=1.595 $Y2=2.4
r56 1 17 18.1727 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.58 $Y=1.35
+ $X2=1.58 $Y2=1.557
r57 1 3 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.58 $Y=1.35 $X2=1.58
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HS__A2111OI_2%B1 1 3 4 5 6 8 9 11 12 13 18
c49 9 0 6.23122e-20 $X=3.465 $Y=1.765
r50 18 20 7.423 $w=4.87e-07 $l=7.5e-08 $layer=POLY_cond $X=3.39 $Y=1.475
+ $X2=3.465 $Y2=1.475
r51 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.39
+ $Y=1.385 $X2=3.39 $Y2=1.385
r52 16 18 37.115 $w=4.87e-07 $l=3.75e-07 $layer=POLY_cond $X=3.015 $Y=1.475
+ $X2=3.39 $Y2=1.475
r53 13 19 6.54089 $w=3.68e-07 $l=2.1e-07 $layer=LI1_cond $X=3.6 $Y=1.365
+ $X2=3.39 $Y2=1.365
r54 12 19 8.40972 $w=3.68e-07 $l=2.7e-07 $layer=LI1_cond $X=3.12 $Y=1.365
+ $X2=3.39 $Y2=1.365
r55 9 20 30.7438 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=3.465 $Y=1.765
+ $X2=3.465 $Y2=1.475
r56 9 11 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.465 $Y=1.765
+ $X2=3.465 $Y2=2.4
r57 6 16 30.7438 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=3.015 $Y=1.765
+ $X2=3.015 $Y2=1.475
r58 6 8 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.015 $Y=1.765
+ $X2=3.015 $Y2=2.4
r59 4 16 34.1696 $w=4.87e-07 $l=2.56076e-07 $layer=POLY_cond $X=2.925 $Y=1.26
+ $X2=3.015 $Y2=1.475
r60 4 5 374.319 $w=1.5e-07 $l=7.3e-07 $layer=POLY_cond $X=2.925 $Y=1.26
+ $X2=2.195 $Y2=1.26
r61 1 5 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.12 $Y=1.185
+ $X2=2.195 $Y2=1.26
r62 1 3 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=2.12 $Y=1.185
+ $X2=2.12 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HS__A2111OI_2%A1 1 3 6 8 10 13 15 16 24
c55 16 0 1.73537e-19 $X=4.56 $Y=1.665
c56 8 0 9.91077e-21 $X=4.365 $Y=1.765
r57 24 25 1.9127 $w=3.78e-07 $l=1.5e-08 $layer=POLY_cond $X=4.365 $Y=1.557
+ $X2=4.38 $Y2=1.557
r58 22 24 29.9656 $w=3.78e-07 $l=2.35e-07 $layer=POLY_cond $X=4.13 $Y=1.557
+ $X2=4.365 $Y2=1.557
r59 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.13
+ $Y=1.515 $X2=4.13 $Y2=1.515
r60 20 22 22.9524 $w=3.78e-07 $l=1.8e-07 $layer=POLY_cond $X=3.95 $Y=1.557
+ $X2=4.13 $Y2=1.557
r61 19 20 4.46296 $w=3.78e-07 $l=3.5e-08 $layer=POLY_cond $X=3.915 $Y=1.557
+ $X2=3.95 $Y2=1.557
r62 16 23 11.5244 $w=4.28e-07 $l=4.3e-07 $layer=LI1_cond $X=4.56 $Y=1.565
+ $X2=4.13 $Y2=1.565
r63 15 23 1.34005 $w=4.28e-07 $l=5e-08 $layer=LI1_cond $X=4.08 $Y=1.565 $X2=4.13
+ $Y2=1.565
r64 11 25 24.4846 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.38 $Y=1.35
+ $X2=4.38 $Y2=1.557
r65 11 13 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=4.38 $Y=1.35
+ $X2=4.38 $Y2=0.74
r66 8 24 24.4846 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=4.365 $Y=1.765
+ $X2=4.365 $Y2=1.557
r67 8 10 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=4.365 $Y=1.765
+ $X2=4.365 $Y2=2.4
r68 4 20 24.4846 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.95 $Y=1.35
+ $X2=3.95 $Y2=1.557
r69 4 6 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=3.95 $Y=1.35 $X2=3.95
+ $Y2=0.74
r70 1 19 24.4846 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=3.915 $Y=1.765
+ $X2=3.915 $Y2=1.557
r71 1 3 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.915 $Y=1.765
+ $X2=3.915 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_HS__A2111OI_2%A2 3 5 7 10 12 14 15 21 22
c38 21 0 9.91077e-21 $X=5.015 $Y=1.515
c39 5 0 1.11225e-19 $X=4.815 $Y=1.765
c40 3 0 2.06049e-19 $X=4.81 $Y=0.74
r41 22 23 1.94879 $w=3.71e-07 $l=1.5e-08 $layer=POLY_cond $X=5.25 $Y=1.557
+ $X2=5.265 $Y2=1.557
r42 20 22 30.531 $w=3.71e-07 $l=2.35e-07 $layer=POLY_cond $X=5.015 $Y=1.557
+ $X2=5.25 $Y2=1.557
r43 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.015
+ $Y=1.515 $X2=5.015 $Y2=1.515
r44 18 20 25.9838 $w=3.71e-07 $l=2e-07 $layer=POLY_cond $X=4.815 $Y=1.557
+ $X2=5.015 $Y2=1.557
r45 17 18 0.649596 $w=3.71e-07 $l=5e-09 $layer=POLY_cond $X=4.81 $Y=1.557
+ $X2=4.815 $Y2=1.557
r46 15 21 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=5.015 $Y=1.665
+ $X2=5.015 $Y2=1.515
r47 12 23 24.032 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=5.265 $Y=1.765
+ $X2=5.265 $Y2=1.557
r48 12 14 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=5.265 $Y=1.765
+ $X2=5.265 $Y2=2.4
r49 8 22 24.032 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=5.25 $Y=1.35 $X2=5.25
+ $Y2=1.557
r50 8 10 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=5.25 $Y=1.35 $X2=5.25
+ $Y2=0.74
r51 5 18 24.032 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=4.815 $Y=1.765
+ $X2=4.815 $Y2=1.557
r52 5 7 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=4.815 $Y=1.765
+ $X2=4.815 $Y2=2.4
r53 1 17 24.032 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.81 $Y=1.35 $X2=4.81
+ $Y2=1.557
r54 1 3 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=4.81 $Y=1.35 $X2=4.81
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HS__A2111OI_2%A_69_368# 1 2 3 12 14 15 18 22 26 28
c36 18 0 5.54777e-20 $X=1.37 $Y=2.115
c37 1 0 1.93692e-19 $X=0.345 $Y=1.84
r38 24 26 20.744 $w=2.48e-07 $l=4.5e-07 $layer=LI1_cond $X=2.31 $Y=2.905
+ $X2=2.31 $Y2=2.455
r39 23 28 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.455 $Y=2.99
+ $X2=1.37 $Y2=2.99
r40 22 24 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=2.185 $Y=2.99
+ $X2=2.31 $Y2=2.905
r41 22 23 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=2.185 $Y=2.99
+ $X2=1.455 $Y2=2.99
r42 18 21 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=1.37 $Y=2.115 $X2=1.37
+ $Y2=2.815
r43 16 28 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.37 $Y=2.905
+ $X2=1.37 $Y2=2.99
r44 16 21 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=1.37 $Y=2.905 $X2=1.37
+ $Y2=2.815
r45 14 28 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.285 $Y=2.99
+ $X2=1.37 $Y2=2.99
r46 14 15 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=1.285 $Y=2.99
+ $X2=0.555 $Y2=2.99
r47 10 15 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.43 $Y=2.905
+ $X2=0.555 $Y2=2.99
r48 10 12 20.744 $w=2.48e-07 $l=4.5e-07 $layer=LI1_cond $X=0.43 $Y=2.905
+ $X2=0.43 $Y2=2.455
r49 3 26 300 $w=1.7e-07 $l=6.85912e-07 $layer=licon1_PDIFF $count=2 $X=2.12
+ $Y=1.84 $X2=2.27 $Y2=2.455
r50 2 21 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=1.22
+ $Y=1.84 $X2=1.37 $Y2=2.815
r51 2 18 400 $w=1.7e-07 $l=3.4187e-07 $layer=licon1_PDIFF $count=1 $X=1.22
+ $Y=1.84 $X2=1.37 $Y2=2.115
r52 1 12 300 $w=1.7e-07 $l=6.74611e-07 $layer=licon1_PDIFF $count=2 $X=0.345
+ $Y=1.84 $X2=0.47 $Y2=2.455
.ends

.subckt PM_SKY130_FD_SC_HS__A2111OI_2%Y 1 2 3 4 13 14 15 16 21 23 27 29 34 35 36
+ 39 44 45
c73 39 0 4.44094e-20 $X=4.165 $Y=0.872
c74 36 0 7.82037e-20 $X=2.335 $Y=0.872
c75 16 0 1.93692e-19 $X=0.355 $Y=2.035
r76 44 45 18.5393 $w=2.28e-07 $l=3.7e-07 $layer=LI1_cond $X=0.24 $Y=1.295
+ $X2=0.24 $Y2=1.665
r77 39 42 2.72396 $w=3.28e-07 $l=7.8e-08 $layer=LI1_cond $X=4.165 $Y=0.872
+ $X2=4.165 $Y2=0.95
r78 36 37 7.78772 $w=3.28e-07 $l=2.23e-07 $layer=LI1_cond $X=2.335 $Y=0.872
+ $X2=2.335 $Y2=1.095
r79 32 45 14.2803 $w=2.28e-07 $l=2.85e-07 $layer=LI1_cond $X=0.24 $Y=1.95
+ $X2=0.24 $Y2=1.665
r80 31 44 5.76222 $w=2.28e-07 $l=1.15e-07 $layer=LI1_cond $X=0.24 $Y=1.18
+ $X2=0.24 $Y2=1.295
r81 30 36 3.54104 $w=2.05e-07 $l=1.65e-07 $layer=LI1_cond $X=2.5 $Y=0.872
+ $X2=2.335 $Y2=0.872
r82 29 39 3.54104 $w=2.05e-07 $l=1.65e-07 $layer=LI1_cond $X=4 $Y=0.872
+ $X2=4.165 $Y2=0.872
r83 29 30 81.153 $w=2.03e-07 $l=1.5e-06 $layer=LI1_cond $X=4 $Y=0.872 $X2=2.5
+ $Y2=0.872
r84 25 36 3.5621 $w=3.28e-07 $l=1.02e-07 $layer=LI1_cond $X=2.335 $Y=0.77
+ $X2=2.335 $Y2=0.872
r85 25 27 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=2.335 $Y=0.77
+ $X2=2.335 $Y2=0.515
r86 24 35 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.49 $Y=1.095
+ $X2=1.325 $Y2=1.095
r87 23 37 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.17 $Y=1.095
+ $X2=2.335 $Y2=1.095
r88 23 24 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=2.17 $Y=1.095
+ $X2=1.49 $Y2=1.095
r89 19 35 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.325 $Y=1.01
+ $X2=1.325 $Y2=1.095
r90 19 21 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=1.325 $Y=1.01
+ $X2=1.325 $Y2=0.515
r91 16 32 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=0.355 $Y=2.035
+ $X2=0.24 $Y2=1.95
r92 15 34 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.755 $Y=2.035
+ $X2=0.92 $Y2=2.035
r93 15 16 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=0.755 $Y=2.035
+ $X2=0.355 $Y2=2.035
r94 14 31 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=0.355 $Y=1.095
+ $X2=0.24 $Y2=1.18
r95 13 35 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.16 $Y=1.095
+ $X2=1.325 $Y2=1.095
r96 13 14 52.5187 $w=1.68e-07 $l=8.05e-07 $layer=LI1_cond $X=1.16 $Y=1.095
+ $X2=0.355 $Y2=1.095
r97 4 34 300 $w=1.7e-07 $l=3.4187e-07 $layer=licon1_PDIFF $count=2 $X=0.77
+ $Y=1.84 $X2=0.92 $Y2=2.115
r98 3 42 182 $w=1.7e-07 $l=6.4622e-07 $layer=licon1_NDIFF $count=1 $X=4.025
+ $Y=0.37 $X2=4.165 $Y2=0.95
r99 2 27 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.195
+ $Y=0.37 $X2=2.335 $Y2=0.515
r100 1 21 91 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=2 $X=1.115
+ $Y=0.37 $X2=1.325 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__A2111OI_2%A_334_368# 1 2 9 14 16
r27 10 14 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.985 $Y=2.035
+ $X2=1.82 $Y2=2.035
r28 9 16 3.99177 $w=1.7e-07 $l=1.5411e-07 $layer=LI1_cond $X=3.075 $Y=2.035
+ $X2=3.2 $Y2=1.97
r29 9 10 71.1123 $w=1.68e-07 $l=1.09e-06 $layer=LI1_cond $X=3.075 $Y=2.035
+ $X2=1.985 $Y2=2.035
r30 2 16 300 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=2 $X=3.09
+ $Y=1.84 $X2=3.24 $Y2=1.985
r31 1 14 300 $w=1.7e-07 $l=3.4187e-07 $layer=licon1_PDIFF $count=2 $X=1.67
+ $Y=1.84 $X2=1.82 $Y2=2.115
.ends

.subckt PM_SKY130_FD_SC_HS__A2111OI_2%A_533_368# 1 2 3 4 15 17 18 19 22 23 27 29
+ 31 33 38
r58 31 40 3.1514 $w=2.5e-07 $l=1.5e-07 $layer=LI1_cond $X=5.53 $Y=2.12 $X2=5.53
+ $Y2=1.97
r59 31 33 12.9074 $w=2.48e-07 $l=2.8e-07 $layer=LI1_cond $X=5.53 $Y=2.12
+ $X2=5.53 $Y2=2.4
r60 30 38 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.675 $Y=2.035
+ $X2=4.55 $Y2=2.035
r61 29 40 3.99177 $w=1.7e-07 $l=1.5411e-07 $layer=LI1_cond $X=5.405 $Y=2.035
+ $X2=5.53 $Y2=1.97
r62 29 30 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=5.405 $Y=2.035
+ $X2=4.675 $Y2=2.035
r63 25 38 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.55 $Y=2.12
+ $X2=4.55 $Y2=2.035
r64 25 27 14.9818 $w=2.48e-07 $l=3.25e-07 $layer=LI1_cond $X=4.55 $Y=2.12
+ $X2=4.55 $Y2=2.445
r65 24 36 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.855 $Y=2.035
+ $X2=3.69 $Y2=2.035
r66 23 38 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.425 $Y=2.035
+ $X2=4.55 $Y2=2.035
r67 23 24 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=4.425 $Y=2.035
+ $X2=3.855 $Y2=2.035
r68 20 22 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=3.69 $Y=2.905 $X2=3.69
+ $Y2=2.815
r69 19 36 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.69 $Y=2.12 $X2=3.69
+ $Y2=2.035
r70 19 22 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=3.69 $Y=2.12
+ $X2=3.69 $Y2=2.815
r71 17 20 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.525 $Y=2.99
+ $X2=3.69 $Y2=2.905
r72 17 18 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=3.525 $Y=2.99
+ $X2=2.905 $Y2=2.99
r73 13 18 7.36005 $w=1.7e-07 $l=1.77482e-07 $layer=LI1_cond $X=2.765 $Y=2.905
+ $X2=2.905 $Y2=2.99
r74 13 15 18.5214 $w=2.78e-07 $l=4.5e-07 $layer=LI1_cond $X=2.765 $Y=2.905
+ $X2=2.765 $Y2=2.455
r75 4 40 600 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=5.34
+ $Y=1.84 $X2=5.49 $Y2=1.985
r76 4 33 300 $w=1.7e-07 $l=6.30555e-07 $layer=licon1_PDIFF $count=2 $X=5.34
+ $Y=1.84 $X2=5.49 $Y2=2.4
r77 3 38 600 $w=1.7e-07 $l=2.59374e-07 $layer=licon1_PDIFF $count=1 $X=4.44
+ $Y=1.84 $X2=4.59 $Y2=2.035
r78 3 27 300 $w=1.7e-07 $l=6.75851e-07 $layer=licon1_PDIFF $count=2 $X=4.44
+ $Y=1.84 $X2=4.59 $Y2=2.445
r79 2 36 400 $w=1.7e-07 $l=2.59374e-07 $layer=licon1_PDIFF $count=1 $X=3.54
+ $Y=1.84 $X2=3.69 $Y2=2.035
r80 2 22 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=3.54
+ $Y=1.84 $X2=3.69 $Y2=2.815
r81 1 15 300 $w=1.7e-07 $l=6.74611e-07 $layer=licon1_PDIFF $count=2 $X=2.665
+ $Y=1.84 $X2=2.79 $Y2=2.455
.ends

.subckt PM_SKY130_FD_SC_HS__A2111OI_2%VPWR 1 2 9 13 15 17 22 29 30 33 36
r59 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r60 33 34 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r61 30 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=5.04 $Y2=3.33
r62 29 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r63 27 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.205 $Y=3.33
+ $X2=5.04 $Y2=3.33
r64 27 29 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=5.205 $Y=3.33
+ $X2=5.52 $Y2=3.33
r65 26 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=5.04 $Y2=3.33
r66 26 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=4.08 $Y2=3.33
r67 25 26 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r68 23 33 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.225 $Y=3.33
+ $X2=4.14 $Y2=3.33
r69 23 25 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=4.225 $Y=3.33
+ $X2=4.56 $Y2=3.33
r70 22 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.875 $Y=3.33
+ $X2=5.04 $Y2=3.33
r71 22 25 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=4.875 $Y=3.33
+ $X2=4.56 $Y2=3.33
r72 19 20 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r73 17 33 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.055 $Y=3.33
+ $X2=4.14 $Y2=3.33
r74 17 19 248.893 $w=1.68e-07 $l=3.815e-06 $layer=LI1_cond $X=4.055 $Y=3.33
+ $X2=0.24 $Y2=3.33
r75 15 34 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=2.88 $Y=3.33
+ $X2=4.08 $Y2=3.33
r76 15 20 0.73586 $w=4.9e-07 $l=2.64e-06 $layer=MET1_cond $X=2.88 $Y=3.33
+ $X2=0.24 $Y2=3.33
r77 11 36 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.04 $Y=3.245
+ $X2=5.04 $Y2=3.33
r78 11 13 29.3349 $w=3.28e-07 $l=8.4e-07 $layer=LI1_cond $X=5.04 $Y=3.245
+ $X2=5.04 $Y2=2.405
r79 7 33 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.14 $Y=3.245 $X2=4.14
+ $Y2=3.33
r80 7 9 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=4.14 $Y=3.245 $X2=4.14
+ $Y2=2.455
r81 2 13 300 $w=1.7e-07 $l=6.3559e-07 $layer=licon1_PDIFF $count=2 $X=4.89
+ $Y=1.84 $X2=5.04 $Y2=2.405
r82 1 9 300 $w=1.7e-07 $l=6.85912e-07 $layer=licon1_PDIFF $count=2 $X=3.99
+ $Y=1.84 $X2=4.14 $Y2=2.455
.ends

.subckt PM_SKY130_FD_SC_HS__A2111OI_2%VGND 1 2 3 14 16 20 24 26 28 38 39 42 45
+ 48
r53 48 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r54 45 46 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r55 43 46 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r56 42 43 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r57 39 49 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=5.04
+ $Y2=0
r58 38 39 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r59 36 48 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=5.2 $Y=0 $X2=5.03
+ $Y2=0
r60 36 38 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=5.2 $Y=0 $X2=5.52
+ $Y2=0
r61 35 49 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=5.04
+ $Y2=0
r62 34 35 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r63 32 46 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.68
+ $Y2=0
r64 31 34 156.578 $w=1.68e-07 $l=2.4e-06 $layer=LI1_cond $X=2.16 $Y=0 $X2=4.56
+ $Y2=0
r65 31 32 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r66 29 45 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=2 $Y=0 $X2=1.83 $Y2=0
r67 29 31 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=2 $Y=0 $X2=2.16
+ $Y2=0
r68 28 48 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=4.86 $Y=0 $X2=5.03
+ $Y2=0
r69 28 34 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=4.86 $Y=0 $X2=4.56
+ $Y2=0
r70 26 35 0.468274 $w=4.9e-07 $l=1.68e-06 $layer=MET1_cond $X=2.88 $Y=0 $X2=4.56
+ $Y2=0
r71 26 32 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=2.88 $Y=0 $X2=2.16
+ $Y2=0
r72 22 48 0.987631 $w=3.4e-07 $l=8.5e-08 $layer=LI1_cond $X=5.03 $Y=0.085
+ $X2=5.03 $Y2=0
r73 22 24 19.9983 $w=3.38e-07 $l=5.9e-07 $layer=LI1_cond $X=5.03 $Y=0.085
+ $X2=5.03 $Y2=0.675
r74 18 45 0.987631 $w=3.4e-07 $l=8.5e-08 $layer=LI1_cond $X=1.83 $Y=0.085
+ $X2=1.83 $Y2=0
r75 18 20 19.9983 $w=3.38e-07 $l=5.9e-07 $layer=LI1_cond $X=1.83 $Y=0.085
+ $X2=1.83 $Y2=0.675
r76 17 42 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.99 $Y=0 $X2=0.825
+ $Y2=0
r77 16 45 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=1.66 $Y=0 $X2=1.83
+ $Y2=0
r78 16 17 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.66 $Y=0 $X2=0.99
+ $Y2=0
r79 12 42 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.825 $Y=0.085
+ $X2=0.825 $Y2=0
r80 12 14 20.6043 $w=3.28e-07 $l=5.9e-07 $layer=LI1_cond $X=0.825 $Y=0.085
+ $X2=0.825 $Y2=0.675
r81 3 24 182 $w=1.7e-07 $l=3.70473e-07 $layer=licon1_NDIFF $count=1 $X=4.885
+ $Y=0.37 $X2=5.03 $Y2=0.675
r82 2 20 182 $w=1.7e-07 $l=3.82623e-07 $layer=licon1_NDIFF $count=1 $X=1.655
+ $Y=0.37 $X2=1.83 $Y2=0.675
r83 1 14 182 $w=1.7e-07 $l=3.70473e-07 $layer=licon1_NDIFF $count=1 $X=0.68
+ $Y=0.37 $X2=0.825 $Y2=0.675
.ends

.subckt PM_SKY130_FD_SC_HS__A2111OI_2%A_722_74# 1 2 3 10 14 18 19 22
c30 14 0 1.6164e-19 $X=4.595 $Y=0.6
r31 20 22 22.8184 $w=2.48e-07 $l=4.95e-07 $layer=LI1_cond $X=5.505 $Y=1.01
+ $X2=5.505 $Y2=0.515
r32 18 20 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=5.38 $Y=1.095
+ $X2=5.505 $Y2=1.01
r33 18 19 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=5.38 $Y=1.095 $X2=4.68
+ $Y2=1.095
r34 15 19 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.595 $Y=1.01
+ $X2=4.68 $Y2=1.095
r35 15 17 2.93583 $w=1.68e-07 $l=4.5e-08 $layer=LI1_cond $X=4.595 $Y=1.01
+ $X2=4.595 $Y2=0.965
r36 14 25 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.595 $Y=0.6
+ $X2=4.595 $Y2=0.475
r37 14 17 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=4.595 $Y=0.6
+ $X2=4.595 $Y2=0.965
r38 10 25 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.51 $Y=0.475
+ $X2=4.595 $Y2=0.475
r39 10 12 35.7257 $w=2.48e-07 $l=7.75e-07 $layer=LI1_cond $X=4.51 $Y=0.475
+ $X2=3.735 $Y2=0.475
r40 3 22 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=5.325
+ $Y=0.37 $X2=5.465 $Y2=0.515
r41 2 25 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=4.455
+ $Y=0.37 $X2=4.595 $Y2=0.515
r42 2 17 182 $w=1.7e-07 $l=6.61306e-07 $layer=licon1_NDIFF $count=1 $X=4.455
+ $Y=0.37 $X2=4.595 $Y2=0.965
r43 1 12 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=3.61
+ $Y=0.37 $X2=3.735 $Y2=0.515
.ends

