* File: sky130_fd_sc_hs__a2bb2o_2.pxi.spice
* Created: Tue Sep  1 19:51:46 2020
* 
x_PM_SKY130_FD_SC_HS__A2BB2O_2%B1 N_B1_c_89_n N_B1_c_95_n N_B1_M1011_g
+ N_B1_c_90_n N_B1_M1008_g N_B1_c_91_n N_B1_c_92_n B1
+ PM_SKY130_FD_SC_HS__A2BB2O_2%B1
x_PM_SKY130_FD_SC_HS__A2BB2O_2%B2 N_B2_M1001_g N_B2_c_118_n N_B2_c_123_n
+ N_B2_M1012_g B2 B2 N_B2_c_120_n N_B2_c_121_n PM_SKY130_FD_SC_HS__A2BB2O_2%B2
x_PM_SKY130_FD_SC_HS__A2BB2O_2%A_293_333# N_A_293_333#_M1006_d
+ N_A_293_333#_M1003_s N_A_293_333#_c_160_n N_A_293_333#_M1002_g
+ N_A_293_333#_c_161_n N_A_293_333#_M1007_g N_A_293_333#_c_162_n
+ N_A_293_333#_c_163_n N_A_293_333#_c_164_n N_A_293_333#_c_165_n
+ N_A_293_333#_c_169_n N_A_293_333#_c_170_n N_A_293_333#_c_166_n
+ PM_SKY130_FD_SC_HS__A2BB2O_2%A_293_333#
x_PM_SKY130_FD_SC_HS__A2BB2O_2%A2_N N_A2_N_M1006_g N_A2_N_c_239_n N_A2_N_M1003_g
+ N_A2_N_c_240_n A2_N N_A2_N_c_242_n PM_SKY130_FD_SC_HS__A2BB2O_2%A2_N
x_PM_SKY130_FD_SC_HS__A2BB2O_2%A1_N N_A1_N_M1010_g N_A1_N_c_280_n N_A1_N_c_284_n
+ N_A1_N_M1013_g A1_N A1_N A1_N N_A1_N_c_282_n PM_SKY130_FD_SC_HS__A2BB2O_2%A1_N
x_PM_SKY130_FD_SC_HS__A2BB2O_2%A_221_74# N_A_221_74#_M1001_d N_A_221_74#_M1002_d
+ N_A_221_74#_M1000_g N_A_221_74#_c_336_n N_A_221_74#_M1004_g
+ N_A_221_74#_c_327_n N_A_221_74#_M1009_g N_A_221_74#_c_338_n
+ N_A_221_74#_M1005_g N_A_221_74#_c_329_n N_A_221_74#_c_330_n
+ N_A_221_74#_c_331_n N_A_221_74#_c_340_n N_A_221_74#_c_341_n
+ N_A_221_74#_c_342_n N_A_221_74#_c_414_p N_A_221_74#_c_332_n
+ N_A_221_74#_c_352_n N_A_221_74#_c_333_n N_A_221_74#_c_344_n
+ N_A_221_74#_c_334_n N_A_221_74#_c_335_n PM_SKY130_FD_SC_HS__A2BB2O_2%A_221_74#
x_PM_SKY130_FD_SC_HS__A2BB2O_2%A_61_392# N_A_61_392#_M1011_s N_A_61_392#_M1012_d
+ N_A_61_392#_c_438_n N_A_61_392#_c_439_n N_A_61_392#_c_440_n
+ N_A_61_392#_c_441_n PM_SKY130_FD_SC_HS__A2BB2O_2%A_61_392#
x_PM_SKY130_FD_SC_HS__A2BB2O_2%VPWR N_VPWR_M1011_d N_VPWR_M1013_d N_VPWR_M1005_s
+ N_VPWR_c_466_n N_VPWR_c_467_n N_VPWR_c_468_n N_VPWR_c_469_n VPWR
+ N_VPWR_c_470_n N_VPWR_c_471_n N_VPWR_c_465_n N_VPWR_c_473_n N_VPWR_c_474_n
+ N_VPWR_c_475_n PM_SKY130_FD_SC_HS__A2BB2O_2%VPWR
x_PM_SKY130_FD_SC_HS__A2BB2O_2%X N_X_M1000_d N_X_M1004_d X X X X X N_X_c_520_n
+ PM_SKY130_FD_SC_HS__A2BB2O_2%X
x_PM_SKY130_FD_SC_HS__A2BB2O_2%VGND N_VGND_M1008_s N_VGND_M1007_d N_VGND_M1010_d
+ N_VGND_M1009_s N_VGND_c_542_n N_VGND_c_543_n N_VGND_c_544_n N_VGND_c_545_n
+ N_VGND_c_546_n N_VGND_c_547_n N_VGND_c_548_n N_VGND_c_549_n VGND
+ N_VGND_c_550_n N_VGND_c_551_n N_VGND_c_552_n N_VGND_c_553_n N_VGND_c_554_n
+ PM_SKY130_FD_SC_HS__A2BB2O_2%VGND
cc_1 VNB N_B1_c_89_n 0.00936933f $X=-0.19 $Y=-0.245 $X2=0.655 $Y2=1.795
cc_2 VNB N_B1_c_90_n 0.0202425f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=1.22
cc_3 VNB N_B1_c_91_n 0.059209f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=1.385
cc_4 VNB N_B1_c_92_n 0.0104458f $X=-0.19 $Y=-0.245 $X2=0.655 $Y2=1.385
cc_5 VNB B1 0.0176299f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_6 VNB N_B2_c_118_n 0.00631214f $X=-0.19 $Y=-0.245 $X2=0.655 $Y2=2.46
cc_7 VNB B2 0.0143856f $X=-0.19 $Y=-0.245 $X2=0.655 $Y2=1.385
cc_8 VNB N_B2_c_120_n 0.0271287f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.385
cc_9 VNB N_B2_c_121_n 0.0176606f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_293_333#_c_160_n 0.0156766f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=0.74
cc_11 VNB N_A_293_333#_c_161_n 0.019625f $X=-0.19 $Y=-0.245 $X2=0.655 $Y2=1.385
cc_12 VNB N_A_293_333#_c_162_n 0.00604743f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_293_333#_c_163_n 0.0556188f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_293_333#_c_164_n 0.0105416f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.385
cc_15 VNB N_A_293_333#_c_165_n 0.00151515f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_293_333#_c_166_n 0.00187269f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A2_N_M1006_g 0.0284145f $X=-0.19 $Y=-0.245 $X2=0.655 $Y2=1.885
cc_18 VNB N_A2_N_c_239_n 7.20236e-19 $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=0.74
cc_19 VNB N_A2_N_c_240_n 0.00862154f $X=-0.19 $Y=-0.245 $X2=0.655 $Y2=1.385
cc_20 VNB A2_N 0.00534845f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_21 VNB N_A2_N_c_242_n 0.0279307f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.385
cc_22 VNB N_A1_N_M1010_g 0.0285108f $X=-0.19 $Y=-0.245 $X2=0.655 $Y2=1.885
cc_23 VNB N_A1_N_c_280_n 0.00501416f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=1.22
cc_24 VNB A1_N 0.00410784f $X=-0.19 $Y=-0.245 $X2=0.655 $Y2=1.385
cc_25 VNB N_A1_N_c_282_n 0.0318604f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.295
cc_26 VNB N_A_221_74#_M1000_g 0.0319619f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=1.385
cc_27 VNB N_A_221_74#_c_327_n 0.00628553f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.385
cc_28 VNB N_A_221_74#_M1009_g 0.0298511f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_221_74#_c_329_n 0.0052061f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_221_74#_c_330_n 0.00345942f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_221_74#_c_331_n 0.0032478f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_221_74#_c_332_n 0.0196001f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_221_74#_c_333_n 0.00114654f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_221_74#_c_334_n 0.00101052f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_221_74#_c_335_n 0.0403155f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_VPWR_c_465_n 0.203486f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_X_c_520_n 0.00240191f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_542_n 0.0344105f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.385
cc_39 VNB N_VGND_c_543_n 0.0150946f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.295
cc_40 VNB N_VGND_c_544_n 0.00604242f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_545_n 0.0427357f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_546_n 0.0113717f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_547_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_548_n 0.0215341f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_VGND_c_549_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_VGND_c_550_n 0.0164632f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_VGND_c_551_n 0.29594f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_VGND_c_552_n 0.0293947f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_VGND_c_553_n 0.0280857f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_VGND_c_554_n 0.00490766f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VPB N_B1_c_89_n 0.00967211f $X=-0.19 $Y=1.66 $X2=0.655 $Y2=1.795
cc_52 VPB N_B1_c_95_n 0.0248047f $X=-0.19 $Y=1.66 $X2=0.655 $Y2=1.885
cc_53 VPB N_B2_c_118_n 0.00675285f $X=-0.19 $Y=1.66 $X2=0.655 $Y2=2.46
cc_54 VPB N_B2_c_123_n 0.0202834f $X=-0.19 $Y=1.66 $X2=0.67 $Y2=1.22
cc_55 VPB N_A_293_333#_c_160_n 0.0369306f $X=-0.19 $Y=1.66 $X2=0.67 $Y2=0.74
cc_56 VPB N_A_293_333#_c_162_n 0.00107914f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_57 VPB N_A_293_333#_c_169_n 0.0200304f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_58 VPB N_A_293_333#_c_170_n 0.0105912f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_59 VPB N_A2_N_c_239_n 0.0282291f $X=-0.19 $Y=1.66 $X2=0.67 $Y2=0.74
cc_60 VPB N_A1_N_c_280_n 0.00285283f $X=-0.19 $Y=1.66 $X2=0.67 $Y2=1.22
cc_61 VPB N_A1_N_c_284_n 0.0185799f $X=-0.19 $Y=1.66 $X2=0.67 $Y2=0.74
cc_62 VPB A1_N 0.00306792f $X=-0.19 $Y=1.66 $X2=0.655 $Y2=1.385
cc_63 VPB N_A_221_74#_c_336_n 0.0161503f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.21
cc_64 VPB N_A_221_74#_c_327_n 0.00761409f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.385
cc_65 VPB N_A_221_74#_c_338_n 0.0171705f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.385
cc_66 VPB N_A_221_74#_c_329_n 0.00624556f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_67 VPB N_A_221_74#_c_340_n 0.0108125f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_68 VPB N_A_221_74#_c_341_n 0.0213935f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_69 VPB N_A_221_74#_c_342_n 0.00952536f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_70 VPB N_A_221_74#_c_332_n 0.0273555f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_71 VPB N_A_221_74#_c_344_n 0.00242448f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_72 VPB N_A_221_74#_c_334_n 0.00333408f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_73 VPB N_A_221_74#_c_335_n 0.0174015f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_74 VPB N_A_61_392#_c_438_n 0.0440661f $X=-0.19 $Y=1.66 $X2=0.565 $Y2=1.385
cc_75 VPB N_A_61_392#_c_439_n 0.015992f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.385
cc_76 VPB N_A_61_392#_c_440_n 0.00959065f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.385
cc_77 VPB N_A_61_392#_c_441_n 0.00290407f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.295
cc_78 VPB N_VPWR_c_466_n 0.00396467f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.385
cc_79 VPB N_VPWR_c_467_n 0.00614661f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_80 VPB N_VPWR_c_468_n 0.0177589f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.385
cc_81 VPB N_VPWR_c_469_n 0.0214006f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_82 VPB N_VPWR_c_470_n 0.0535977f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_83 VPB N_VPWR_c_471_n 0.0150312f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_84 VPB N_VPWR_c_465_n 0.0904416f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_85 VPB N_VPWR_c_473_n 0.0288171f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_86 VPB N_VPWR_c_474_n 0.00729535f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_87 VPB N_VPWR_c_475_n 0.00614127f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_88 VPB N_X_c_520_n 4.33269e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_89 N_B1_c_89_n N_B2_c_118_n 0.0084355f $X=0.655 $Y=1.795 $X2=0 $Y2=0
cc_90 N_B1_c_95_n N_B2_c_123_n 0.0276501f $X=0.655 $Y=1.885 $X2=0 $Y2=0
cc_91 N_B1_c_90_n B2 0.00732765f $X=0.67 $Y=1.22 $X2=0 $Y2=0
cc_92 N_B1_c_92_n B2 0.0141119f $X=0.655 $Y=1.385 $X2=0 $Y2=0
cc_93 B1 B2 0.0295948f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_94 N_B1_c_92_n N_B2_c_120_n 0.0396846f $X=0.655 $Y=1.385 $X2=0 $Y2=0
cc_95 N_B1_c_90_n N_B2_c_121_n 0.0396846f $X=0.67 $Y=1.22 $X2=0 $Y2=0
cc_96 N_B1_c_90_n N_A_221_74#_c_330_n 0.00179159f $X=0.67 $Y=1.22 $X2=0 $Y2=0
cc_97 N_B1_c_95_n N_A_61_392#_c_438_n 0.00846769f $X=0.655 $Y=1.885 $X2=0 $Y2=0
cc_98 N_B1_c_89_n N_A_61_392#_c_439_n 0.0071463f $X=0.655 $Y=1.795 $X2=0 $Y2=0
cc_99 N_B1_c_95_n N_A_61_392#_c_439_n 0.0110211f $X=0.655 $Y=1.885 $X2=0 $Y2=0
cc_100 N_B1_c_91_n N_A_61_392#_c_439_n 0.00184075f $X=0.565 $Y=1.385 $X2=0 $Y2=0
cc_101 N_B1_c_91_n N_A_61_392#_c_440_n 0.00493733f $X=0.565 $Y=1.385 $X2=0 $Y2=0
cc_102 B1 N_A_61_392#_c_440_n 0.0144344f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_103 N_B1_c_95_n N_VPWR_c_466_n 0.0190232f $X=0.655 $Y=1.885 $X2=0 $Y2=0
cc_104 N_B1_c_95_n N_VPWR_c_465_n 0.00821622f $X=0.655 $Y=1.885 $X2=0 $Y2=0
cc_105 N_B1_c_95_n N_VPWR_c_473_n 0.00413917f $X=0.655 $Y=1.885 $X2=0 $Y2=0
cc_106 N_B1_c_90_n N_VGND_c_542_n 0.0162081f $X=0.67 $Y=1.22 $X2=0 $Y2=0
cc_107 N_B1_c_91_n N_VGND_c_542_n 0.00663559f $X=0.565 $Y=1.385 $X2=0 $Y2=0
cc_108 B1 N_VGND_c_542_n 0.0125933f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_109 N_B1_c_90_n N_VGND_c_551_n 0.0075694f $X=0.67 $Y=1.22 $X2=0 $Y2=0
cc_110 N_B1_c_90_n N_VGND_c_552_n 0.00383152f $X=0.67 $Y=1.22 $X2=0 $Y2=0
cc_111 N_B2_c_118_n N_A_293_333#_c_160_n 0.0145534f $X=1.105 $Y=1.795 $X2=0
+ $Y2=0
cc_112 N_B2_c_123_n N_A_293_333#_c_160_n 0.00770144f $X=1.105 $Y=1.885 $X2=0
+ $Y2=0
cc_113 B2 N_A_293_333#_c_160_n 6.15159e-19 $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_114 N_B2_c_120_n N_A_293_333#_c_160_n 0.0215146f $X=1.12 $Y=1.385 $X2=0 $Y2=0
cc_115 B2 N_A_293_333#_c_161_n 7.52582e-19 $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_116 N_B2_c_121_n N_A_293_333#_c_161_n 0.0078714f $X=1.12 $Y=1.22 $X2=0 $Y2=0
cc_117 N_B2_c_121_n N_A_221_74#_c_330_n 0.00863182f $X=1.12 $Y=1.22 $X2=0 $Y2=0
cc_118 B2 N_A_221_74#_c_331_n 0.0168621f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_119 N_B2_c_120_n N_A_221_74#_c_331_n 4.33788e-19 $X=1.12 $Y=1.385 $X2=0 $Y2=0
cc_120 N_B2_c_121_n N_A_221_74#_c_331_n 0.00128434f $X=1.12 $Y=1.22 $X2=0 $Y2=0
cc_121 B2 N_A_221_74#_c_352_n 0.0176548f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_122 N_B2_c_120_n N_A_221_74#_c_352_n 0.00110623f $X=1.12 $Y=1.385 $X2=0 $Y2=0
cc_123 N_B2_c_121_n N_A_221_74#_c_352_n 0.00303924f $X=1.12 $Y=1.22 $X2=0 $Y2=0
cc_124 B2 N_A_221_74#_c_333_n 0.0147664f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_125 N_B2_c_120_n N_A_221_74#_c_333_n 4.94042e-19 $X=1.12 $Y=1.385 $X2=0 $Y2=0
cc_126 N_B2_c_118_n N_A_221_74#_c_334_n 0.00101298f $X=1.105 $Y=1.795 $X2=0
+ $Y2=0
cc_127 N_B2_c_123_n N_A_221_74#_c_334_n 2.62141e-19 $X=1.105 $Y=1.885 $X2=0
+ $Y2=0
cc_128 N_B2_c_118_n N_A_61_392#_c_439_n 0.00516691f $X=1.105 $Y=1.795 $X2=0
+ $Y2=0
cc_129 N_B2_c_123_n N_A_61_392#_c_439_n 0.00999603f $X=1.105 $Y=1.885 $X2=0
+ $Y2=0
cc_130 B2 N_A_61_392#_c_439_n 0.0542449f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_131 N_B2_c_120_n N_A_61_392#_c_439_n 0.00363229f $X=1.12 $Y=1.385 $X2=0 $Y2=0
cc_132 N_B2_c_123_n N_A_61_392#_c_441_n 0.00658191f $X=1.105 $Y=1.885 $X2=0
+ $Y2=0
cc_133 N_B2_c_123_n N_VPWR_c_466_n 0.0158814f $X=1.105 $Y=1.885 $X2=0 $Y2=0
cc_134 N_B2_c_123_n N_VPWR_c_470_n 0.00413917f $X=1.105 $Y=1.885 $X2=0 $Y2=0
cc_135 N_B2_c_123_n N_VPWR_c_465_n 0.0081781f $X=1.105 $Y=1.885 $X2=0 $Y2=0
cc_136 B2 N_VGND_c_542_n 0.00112687f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_137 N_B2_c_121_n N_VGND_c_542_n 0.00236525f $X=1.12 $Y=1.22 $X2=0 $Y2=0
cc_138 N_B2_c_121_n N_VGND_c_551_n 0.00821699f $X=1.12 $Y=1.22 $X2=0 $Y2=0
cc_139 N_B2_c_121_n N_VGND_c_552_n 0.00434272f $X=1.12 $Y=1.22 $X2=0 $Y2=0
cc_140 N_A_293_333#_c_162_n N_A2_N_M1006_g 0.00516264f $X=2.01 $Y=1.385 $X2=0
+ $Y2=0
cc_141 N_A_293_333#_c_164_n N_A2_N_M1006_g 0.0130552f $X=2.69 $Y=0.925 $X2=0
+ $Y2=0
cc_142 N_A_293_333#_c_166_n N_A2_N_M1006_g 4.84042e-19 $X=2.785 $Y=0.645 $X2=0
+ $Y2=0
cc_143 N_A_293_333#_c_169_n N_A2_N_c_239_n 0.00636618f $X=2.422 $Y=1.85 $X2=0
+ $Y2=0
cc_144 N_A_293_333#_c_170_n N_A2_N_c_239_n 0.00191916f $X=2.43 $Y=2.05 $X2=0
+ $Y2=0
cc_145 N_A_293_333#_c_162_n N_A2_N_c_240_n 0.00391824f $X=2.01 $Y=1.385 $X2=0
+ $Y2=0
cc_146 N_A_293_333#_c_163_n N_A2_N_c_240_n 0.00144075f $X=2.01 $Y=1.385 $X2=0
+ $Y2=0
cc_147 N_A_293_333#_c_162_n A2_N 0.0207819f $X=2.01 $Y=1.385 $X2=0 $Y2=0
cc_148 N_A_293_333#_c_163_n A2_N 0.00115534f $X=2.01 $Y=1.385 $X2=0 $Y2=0
cc_149 N_A_293_333#_c_164_n A2_N 0.027957f $X=2.69 $Y=0.925 $X2=0 $Y2=0
cc_150 N_A_293_333#_c_169_n A2_N 0.0145994f $X=2.422 $Y=1.85 $X2=0 $Y2=0
cc_151 N_A_293_333#_c_162_n N_A2_N_c_242_n 6.38029e-19 $X=2.01 $Y=1.385 $X2=0
+ $Y2=0
cc_152 N_A_293_333#_c_163_n N_A2_N_c_242_n 0.0192745f $X=2.01 $Y=1.385 $X2=0
+ $Y2=0
cc_153 N_A_293_333#_c_164_n N_A2_N_c_242_n 0.00432985f $X=2.69 $Y=0.925 $X2=0
+ $Y2=0
cc_154 N_A_293_333#_c_169_n N_A2_N_c_242_n 0.00431149f $X=2.422 $Y=1.85 $X2=0
+ $Y2=0
cc_155 N_A_293_333#_c_164_n N_A1_N_M1010_g 0.00160245f $X=2.69 $Y=0.925 $X2=0
+ $Y2=0
cc_156 N_A_293_333#_c_166_n N_A1_N_M1010_g 4.77224e-19 $X=2.785 $Y=0.645 $X2=0
+ $Y2=0
cc_157 N_A_293_333#_c_169_n A1_N 0.00824122f $X=2.422 $Y=1.85 $X2=0 $Y2=0
cc_158 N_A_293_333#_c_170_n A1_N 0.0085385f $X=2.43 $Y=2.05 $X2=0 $Y2=0
cc_159 N_A_293_333#_c_161_n N_A_221_74#_c_330_n 3.42943e-19 $X=1.57 $Y=1.22
+ $X2=0 $Y2=0
cc_160 N_A_293_333#_c_160_n N_A_221_74#_c_331_n 0.00295591f $X=1.555 $Y=1.885
+ $X2=0 $Y2=0
cc_161 N_A_293_333#_c_161_n N_A_221_74#_c_331_n 0.00645454f $X=1.57 $Y=1.22
+ $X2=0 $Y2=0
cc_162 N_A_293_333#_c_162_n N_A_221_74#_c_331_n 0.0167429f $X=2.01 $Y=1.385
+ $X2=0 $Y2=0
cc_163 N_A_293_333#_c_163_n N_A_221_74#_c_331_n 0.00314762f $X=2.01 $Y=1.385
+ $X2=0 $Y2=0
cc_164 N_A_293_333#_c_160_n N_A_221_74#_c_340_n 0.00984649f $X=1.555 $Y=1.885
+ $X2=0 $Y2=0
cc_165 N_A_293_333#_M1003_s N_A_221_74#_c_341_n 0.00273279f $X=2.305 $Y=1.89
+ $X2=0 $Y2=0
cc_166 N_A_293_333#_c_170_n N_A_221_74#_c_341_n 0.0200424f $X=2.43 $Y=2.05 $X2=0
+ $Y2=0
cc_167 N_A_293_333#_c_161_n N_A_221_74#_c_352_n 0.00866889f $X=1.57 $Y=1.22
+ $X2=0 $Y2=0
cc_168 N_A_293_333#_c_160_n N_A_221_74#_c_333_n 0.00773775f $X=1.555 $Y=1.885
+ $X2=0 $Y2=0
cc_169 N_A_293_333#_c_162_n N_A_221_74#_c_333_n 0.0122188f $X=2.01 $Y=1.385
+ $X2=0 $Y2=0
cc_170 N_A_293_333#_c_163_n N_A_221_74#_c_333_n 0.00855797f $X=2.01 $Y=1.385
+ $X2=0 $Y2=0
cc_171 N_A_293_333#_c_160_n N_A_221_74#_c_344_n 0.00206972f $X=1.555 $Y=1.885
+ $X2=0 $Y2=0
cc_172 N_A_293_333#_c_163_n N_A_221_74#_c_344_n 0.00552706f $X=2.01 $Y=1.385
+ $X2=0 $Y2=0
cc_173 N_A_293_333#_c_169_n N_A_221_74#_c_344_n 0.00156692f $X=2.422 $Y=1.85
+ $X2=0 $Y2=0
cc_174 N_A_293_333#_c_170_n N_A_221_74#_c_344_n 0.0333926f $X=2.43 $Y=2.05 $X2=0
+ $Y2=0
cc_175 N_A_293_333#_c_160_n N_A_221_74#_c_334_n 0.0143878f $X=1.555 $Y=1.885
+ $X2=0 $Y2=0
cc_176 N_A_293_333#_c_162_n N_A_221_74#_c_334_n 0.0100833f $X=2.01 $Y=1.385
+ $X2=0 $Y2=0
cc_177 N_A_293_333#_c_163_n N_A_221_74#_c_334_n 0.00263747f $X=2.01 $Y=1.385
+ $X2=0 $Y2=0
cc_178 N_A_293_333#_c_169_n N_A_221_74#_c_334_n 0.0141439f $X=2.422 $Y=1.85
+ $X2=0 $Y2=0
cc_179 N_A_293_333#_c_170_n N_A_221_74#_c_334_n 0.00616994f $X=2.43 $Y=2.05
+ $X2=0 $Y2=0
cc_180 N_A_293_333#_c_160_n N_A_61_392#_c_439_n 0.00138997f $X=1.555 $Y=1.885
+ $X2=0 $Y2=0
cc_181 N_A_293_333#_c_160_n N_A_61_392#_c_441_n 0.00335433f $X=1.555 $Y=1.885
+ $X2=0 $Y2=0
cc_182 N_A_293_333#_c_160_n N_VPWR_c_466_n 8.1496e-19 $X=1.555 $Y=1.885 $X2=0
+ $Y2=0
cc_183 N_A_293_333#_c_160_n N_VPWR_c_470_n 0.00410479f $X=1.555 $Y=1.885 $X2=0
+ $Y2=0
cc_184 N_A_293_333#_c_160_n N_VPWR_c_465_n 0.00749507f $X=1.555 $Y=1.885 $X2=0
+ $Y2=0
cc_185 N_A_293_333#_c_164_n N_X_c_520_n 0.0022519f $X=2.69 $Y=0.925 $X2=0 $Y2=0
cc_186 N_A_293_333#_c_164_n N_VGND_M1007_d 0.00336173f $X=2.69 $Y=0.925 $X2=0
+ $Y2=0
cc_187 N_A_293_333#_c_165_n N_VGND_M1007_d 0.00472124f $X=2.175 $Y=0.925 $X2=0
+ $Y2=0
cc_188 N_A_293_333#_c_166_n N_VGND_c_543_n 0.00792522f $X=2.785 $Y=0.645 $X2=0
+ $Y2=0
cc_189 N_A_293_333#_c_164_n N_VGND_c_544_n 0.00433169f $X=2.69 $Y=0.925 $X2=0
+ $Y2=0
cc_190 N_A_293_333#_c_166_n N_VGND_c_544_n 0.0176744f $X=2.785 $Y=0.645 $X2=0
+ $Y2=0
cc_191 N_A_293_333#_c_161_n N_VGND_c_551_n 0.00468239f $X=1.57 $Y=1.22 $X2=0
+ $Y2=0
cc_192 N_A_293_333#_c_164_n N_VGND_c_551_n 0.00606296f $X=2.69 $Y=0.925 $X2=0
+ $Y2=0
cc_193 N_A_293_333#_c_165_n N_VGND_c_551_n 9.1246e-19 $X=2.175 $Y=0.925 $X2=0
+ $Y2=0
cc_194 N_A_293_333#_c_166_n N_VGND_c_551_n 0.00656744f $X=2.785 $Y=0.645 $X2=0
+ $Y2=0
cc_195 N_A_293_333#_c_161_n N_VGND_c_552_n 0.00461464f $X=1.57 $Y=1.22 $X2=0
+ $Y2=0
cc_196 N_A_293_333#_c_161_n N_VGND_c_553_n 0.00585758f $X=1.57 $Y=1.22 $X2=0
+ $Y2=0
cc_197 N_A_293_333#_c_163_n N_VGND_c_553_n 0.00822318f $X=2.01 $Y=1.385 $X2=0
+ $Y2=0
cc_198 N_A_293_333#_c_164_n N_VGND_c_553_n 0.0226052f $X=2.69 $Y=0.925 $X2=0
+ $Y2=0
cc_199 N_A_293_333#_c_165_n N_VGND_c_553_n 0.0218905f $X=2.175 $Y=0.925 $X2=0
+ $Y2=0
cc_200 N_A_293_333#_c_166_n N_VGND_c_553_n 0.0141617f $X=2.785 $Y=0.645 $X2=0
+ $Y2=0
cc_201 N_A2_N_M1006_g N_A1_N_M1010_g 0.023397f $X=2.57 $Y=0.645 $X2=0 $Y2=0
cc_202 A2_N N_A1_N_M1010_g 0.00184827f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_203 N_A2_N_c_242_n N_A1_N_M1010_g 0.0115108f $X=2.55 $Y=1.345 $X2=0 $Y2=0
cc_204 N_A2_N_c_239_n N_A1_N_c_280_n 0.0092314f $X=2.655 $Y=1.815 $X2=0 $Y2=0
cc_205 N_A2_N_c_240_n N_A1_N_c_280_n 0.0054529f $X=2.655 $Y=1.66 $X2=0 $Y2=0
cc_206 N_A2_N_c_239_n N_A1_N_c_284_n 0.0584024f $X=2.655 $Y=1.815 $X2=0 $Y2=0
cc_207 N_A2_N_c_239_n A1_N 0.00273903f $X=2.655 $Y=1.815 $X2=0 $Y2=0
cc_208 N_A2_N_c_240_n A1_N 0.00242122f $X=2.655 $Y=1.66 $X2=0 $Y2=0
cc_209 A2_N A1_N 0.0262861f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_210 N_A2_N_c_242_n A1_N 6.48348e-19 $X=2.55 $Y=1.345 $X2=0 $Y2=0
cc_211 N_A2_N_c_240_n N_A1_N_c_282_n 0.0115108f $X=2.655 $Y=1.66 $X2=0 $Y2=0
cc_212 N_A2_N_c_239_n N_A_221_74#_c_341_n 0.0154956f $X=2.655 $Y=1.815 $X2=0
+ $Y2=0
cc_213 N_A2_N_c_239_n N_A_221_74#_c_344_n 0.00487538f $X=2.655 $Y=1.815 $X2=0
+ $Y2=0
cc_214 N_A2_N_c_239_n N_VPWR_c_467_n 3.7546e-19 $X=2.655 $Y=1.815 $X2=0 $Y2=0
cc_215 N_A2_N_c_239_n N_VPWR_c_470_n 0.00375243f $X=2.655 $Y=1.815 $X2=0 $Y2=0
cc_216 N_A2_N_c_239_n N_VPWR_c_465_n 0.00523671f $X=2.655 $Y=1.815 $X2=0 $Y2=0
cc_217 N_A2_N_M1006_g N_VGND_c_543_n 0.00383152f $X=2.57 $Y=0.645 $X2=0 $Y2=0
cc_218 N_A2_N_M1006_g N_VGND_c_544_n 5.49548e-19 $X=2.57 $Y=0.645 $X2=0 $Y2=0
cc_219 N_A2_N_M1006_g N_VGND_c_551_n 0.00382415f $X=2.57 $Y=0.645 $X2=0 $Y2=0
cc_220 N_A2_N_M1006_g N_VGND_c_553_n 0.00912161f $X=2.57 $Y=0.645 $X2=0 $Y2=0
cc_221 N_A1_N_M1010_g N_A_221_74#_M1000_g 0.0204801f $X=3 $Y=0.645 $X2=0 $Y2=0
cc_222 A1_N N_A_221_74#_M1000_g 0.001321f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_223 N_A1_N_c_282_n N_A_221_74#_M1000_g 0.0191691f $X=3.09 $Y=1.385 $X2=0
+ $Y2=0
cc_224 N_A1_N_c_284_n N_A_221_74#_c_336_n 0.0291524f $X=3.045 $Y=1.815 $X2=0
+ $Y2=0
cc_225 A1_N N_A_221_74#_c_336_n 0.00259969f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_226 N_A1_N_c_280_n N_A_221_74#_c_329_n 0.00754656f $X=3.045 $Y=1.725 $X2=0
+ $Y2=0
cc_227 A1_N N_A_221_74#_c_329_n 0.00165197f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_228 N_A1_N_c_284_n N_A_221_74#_c_341_n 0.00100688f $X=3.045 $Y=1.815 $X2=0
+ $Y2=0
cc_229 N_A1_N_c_284_n N_A_221_74#_c_342_n 0.0114471f $X=3.045 $Y=1.815 $X2=0
+ $Y2=0
cc_230 A1_N N_A_221_74#_c_342_n 0.0176909f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_231 A1_N N_VPWR_M1013_d 0.00389938f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_232 N_A1_N_c_284_n N_VPWR_c_467_n 0.00610303f $X=3.045 $Y=1.815 $X2=0 $Y2=0
cc_233 N_A1_N_c_284_n N_VPWR_c_470_n 0.00473462f $X=3.045 $Y=1.815 $X2=0 $Y2=0
cc_234 N_A1_N_c_284_n N_VPWR_c_465_n 0.00474795f $X=3.045 $Y=1.815 $X2=0 $Y2=0
cc_235 N_A1_N_M1010_g N_X_c_520_n 0.00152927f $X=3 $Y=0.645 $X2=0 $Y2=0
cc_236 N_A1_N_c_280_n N_X_c_520_n 2.76261e-19 $X=3.045 $Y=1.725 $X2=0 $Y2=0
cc_237 N_A1_N_c_284_n N_X_c_520_n 3.51282e-19 $X=3.045 $Y=1.815 $X2=0 $Y2=0
cc_238 A1_N N_X_c_520_n 0.0605438f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_239 N_A1_N_c_282_n N_X_c_520_n 0.00111347f $X=3.09 $Y=1.385 $X2=0 $Y2=0
cc_240 N_A1_N_M1010_g N_VGND_c_543_n 0.00383152f $X=3 $Y=0.645 $X2=0 $Y2=0
cc_241 N_A1_N_M1010_g N_VGND_c_544_n 0.0125324f $X=3 $Y=0.645 $X2=0 $Y2=0
cc_242 A1_N N_VGND_c_544_n 0.0146144f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_243 N_A1_N_c_282_n N_VGND_c_544_n 0.00123829f $X=3.09 $Y=1.385 $X2=0 $Y2=0
cc_244 N_A1_N_M1010_g N_VGND_c_551_n 0.00757637f $X=3 $Y=0.645 $X2=0 $Y2=0
cc_245 N_A1_N_M1010_g N_VGND_c_553_n 4.13238e-19 $X=3 $Y=0.645 $X2=0 $Y2=0
cc_246 N_A_221_74#_c_334_n N_A_61_392#_c_439_n 0.01368f $X=1.765 $Y=2.02 $X2=0
+ $Y2=0
cc_247 N_A_221_74#_c_340_n N_A_61_392#_c_441_n 0.0133878f $X=1.765 $Y=2.81 $X2=0
+ $Y2=0
cc_248 N_A_221_74#_c_334_n N_A_61_392#_c_441_n 0.0677988f $X=1.765 $Y=2.02 $X2=0
+ $Y2=0
cc_249 N_A_221_74#_c_342_n N_VPWR_M1013_d 0.0098464f $X=4.09 $Y=2.405 $X2=0
+ $Y2=0
cc_250 N_A_221_74#_c_342_n N_VPWR_M1005_s 0.00327359f $X=4.09 $Y=2.405 $X2=0
+ $Y2=0
cc_251 N_A_221_74#_c_332_n N_VPWR_M1005_s 0.00367736f $X=4.255 $Y=1.515 $X2=0
+ $Y2=0
cc_252 N_A_221_74#_c_336_n N_VPWR_c_467_n 0.0106187f $X=3.555 $Y=1.765 $X2=0
+ $Y2=0
cc_253 N_A_221_74#_c_338_n N_VPWR_c_467_n 0.00127018f $X=4.005 $Y=1.765 $X2=0
+ $Y2=0
cc_254 N_A_221_74#_c_341_n N_VPWR_c_467_n 0.0100491f $X=2.75 $Y=2.895 $X2=0
+ $Y2=0
cc_255 N_A_221_74#_c_342_n N_VPWR_c_467_n 0.0215778f $X=4.09 $Y=2.405 $X2=0
+ $Y2=0
cc_256 N_A_221_74#_c_336_n N_VPWR_c_468_n 0.00413917f $X=3.555 $Y=1.765 $X2=0
+ $Y2=0
cc_257 N_A_221_74#_c_338_n N_VPWR_c_468_n 0.00413917f $X=4.005 $Y=1.765 $X2=0
+ $Y2=0
cc_258 N_A_221_74#_c_336_n N_VPWR_c_469_n 0.00127141f $X=3.555 $Y=1.765 $X2=0
+ $Y2=0
cc_259 N_A_221_74#_c_338_n N_VPWR_c_469_n 0.0106215f $X=4.005 $Y=1.765 $X2=0
+ $Y2=0
cc_260 N_A_221_74#_c_342_n N_VPWR_c_469_n 0.0237488f $X=4.09 $Y=2.405 $X2=0
+ $Y2=0
cc_261 N_A_221_74#_c_340_n N_VPWR_c_470_n 0.0159103f $X=1.765 $Y=2.81 $X2=0
+ $Y2=0
cc_262 N_A_221_74#_c_341_n N_VPWR_c_470_n 0.0396437f $X=2.75 $Y=2.895 $X2=0
+ $Y2=0
cc_263 N_A_221_74#_c_336_n N_VPWR_c_465_n 0.00414505f $X=3.555 $Y=1.765 $X2=0
+ $Y2=0
cc_264 N_A_221_74#_c_338_n N_VPWR_c_465_n 0.00414505f $X=4.005 $Y=1.765 $X2=0
+ $Y2=0
cc_265 N_A_221_74#_c_340_n N_VPWR_c_465_n 0.0130733f $X=1.765 $Y=2.81 $X2=0
+ $Y2=0
cc_266 N_A_221_74#_c_341_n N_VPWR_c_465_n 0.0346145f $X=2.75 $Y=2.895 $X2=0
+ $Y2=0
cc_267 N_A_221_74#_c_342_n N_VPWR_c_465_n 0.0291572f $X=4.09 $Y=2.405 $X2=0
+ $Y2=0
cc_268 N_A_221_74#_c_414_p A_546_378# 0.00569187f $X=2.92 $Y=2.405 $X2=-0.19
+ $Y2=-0.245
cc_269 N_A_221_74#_c_342_n N_X_M1004_d 0.00556519f $X=4.09 $Y=2.405 $X2=0 $Y2=0
cc_270 N_A_221_74#_M1000_g N_X_c_520_n 0.030377f $X=3.54 $Y=0.74 $X2=0 $Y2=0
cc_271 N_A_221_74#_c_336_n N_X_c_520_n 0.0103241f $X=3.555 $Y=1.765 $X2=0 $Y2=0
cc_272 N_A_221_74#_c_327_n N_X_c_520_n 0.0114285f $X=3.895 $Y=1.605 $X2=0 $Y2=0
cc_273 N_A_221_74#_M1009_g N_X_c_520_n 0.0223512f $X=3.97 $Y=0.74 $X2=0 $Y2=0
cc_274 N_A_221_74#_c_338_n N_X_c_520_n 6.44513e-19 $X=4.005 $Y=1.765 $X2=0 $Y2=0
cc_275 N_A_221_74#_c_329_n N_X_c_520_n 0.00632342f $X=3.555 $Y=1.605 $X2=0 $Y2=0
cc_276 N_A_221_74#_c_342_n N_X_c_520_n 0.0260598f $X=4.09 $Y=2.405 $X2=0 $Y2=0
cc_277 N_A_221_74#_c_332_n N_X_c_520_n 0.0385107f $X=4.255 $Y=1.515 $X2=0 $Y2=0
cc_278 N_A_221_74#_c_335_n N_X_c_520_n 0.0102738f $X=4.005 $Y=1.557 $X2=0 $Y2=0
cc_279 N_A_221_74#_c_330_n N_VGND_c_542_n 0.0225615f $X=1.3 $Y=0.495 $X2=0 $Y2=0
cc_280 N_A_221_74#_M1000_g N_VGND_c_544_n 0.00687023f $X=3.54 $Y=0.74 $X2=0
+ $Y2=0
cc_281 N_A_221_74#_M1009_g N_VGND_c_545_n 0.00647412f $X=3.97 $Y=0.74 $X2=0
+ $Y2=0
cc_282 N_A_221_74#_c_332_n N_VGND_c_545_n 0.0181982f $X=4.255 $Y=1.515 $X2=0
+ $Y2=0
cc_283 N_A_221_74#_c_335_n N_VGND_c_545_n 0.00190129f $X=4.005 $Y=1.557 $X2=0
+ $Y2=0
cc_284 N_A_221_74#_M1000_g N_VGND_c_548_n 0.00315306f $X=3.54 $Y=0.74 $X2=0
+ $Y2=0
cc_285 N_A_221_74#_M1009_g N_VGND_c_548_n 0.00434272f $X=3.97 $Y=0.74 $X2=0
+ $Y2=0
cc_286 N_A_221_74#_M1000_g N_VGND_c_551_n 0.00437087f $X=3.54 $Y=0.74 $X2=0
+ $Y2=0
cc_287 N_A_221_74#_M1009_g N_VGND_c_551_n 0.00825283f $X=3.97 $Y=0.74 $X2=0
+ $Y2=0
cc_288 N_A_221_74#_c_330_n N_VGND_c_551_n 0.0145687f $X=1.3 $Y=0.495 $X2=0 $Y2=0
cc_289 N_A_221_74#_c_352_n N_VGND_c_551_n 0.00533986f $X=1.367 $Y=1.01 $X2=0
+ $Y2=0
cc_290 N_A_221_74#_c_330_n N_VGND_c_552_n 0.017649f $X=1.3 $Y=0.495 $X2=0 $Y2=0
cc_291 N_A_221_74#_c_330_n N_VGND_c_553_n 0.00170296f $X=1.3 $Y=0.495 $X2=0
+ $Y2=0
cc_292 N_A_61_392#_c_438_n N_VPWR_c_466_n 0.0617165f $X=0.43 $Y=2.105 $X2=0
+ $Y2=0
cc_293 N_A_61_392#_c_439_n N_VPWR_c_466_n 0.021739f $X=1.245 $Y=1.805 $X2=0
+ $Y2=0
cc_294 N_A_61_392#_c_441_n N_VPWR_c_466_n 0.0599532f $X=1.33 $Y=2.105 $X2=0
+ $Y2=0
cc_295 N_A_61_392#_c_441_n N_VPWR_c_470_n 0.00749631f $X=1.33 $Y=2.105 $X2=0
+ $Y2=0
cc_296 N_A_61_392#_c_438_n N_VPWR_c_465_n 0.00915947f $X=0.43 $Y=2.105 $X2=0
+ $Y2=0
cc_297 N_A_61_392#_c_441_n N_VPWR_c_465_n 0.0062048f $X=1.33 $Y=2.105 $X2=0
+ $Y2=0
cc_298 N_A_61_392#_c_438_n N_VPWR_c_473_n 0.011066f $X=0.43 $Y=2.105 $X2=0 $Y2=0
cc_299 N_X_c_520_n N_VGND_c_544_n 0.0460212f $X=3.755 $Y=0.515 $X2=0 $Y2=0
cc_300 N_X_c_520_n N_VGND_c_545_n 0.030619f $X=3.755 $Y=0.515 $X2=0 $Y2=0
cc_301 N_X_c_520_n N_VGND_c_548_n 0.0188635f $X=3.755 $Y=0.515 $X2=0 $Y2=0
cc_302 N_X_c_520_n N_VGND_c_551_n 0.0152542f $X=3.755 $Y=0.515 $X2=0 $Y2=0
