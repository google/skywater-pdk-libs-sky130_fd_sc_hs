# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_hs__a211o_1
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_hs__a211o_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.840000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.045000 1.450000 2.755000 1.780000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.585000 1.450000 1.835000 1.780000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.045000 0.255000 2.875000 0.570000 ;
        RECT 2.045000 0.570000 2.275000 0.670000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.385000 0.255000 3.715000 0.670000 ;
    END
  END C1
  PIN X
    ANTENNADIFFAREA  0.504100 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.435000 1.075000 1.130000 ;
        RECT 0.085000 1.130000 0.255000 1.820000 ;
        RECT 0.085000 1.820000 0.435000 2.980000 ;
        RECT 0.825000 0.345000 1.075000 0.435000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 3.840000 0.085000 ;
        RECT 1.255000  0.085000 1.705000 0.940000 ;
        RECT 2.780000  0.740000 3.215000 0.910000 ;
        RECT 3.045000  0.085000 3.215000 0.740000 ;
      LAYER mcon ;
        RECT 0.155000 -0.085000 0.325000 0.085000 ;
        RECT 0.635000 -0.085000 0.805000 0.085000 ;
        RECT 1.115000 -0.085000 1.285000 0.085000 ;
        RECT 1.595000 -0.085000 1.765000 0.085000 ;
        RECT 2.075000 -0.085000 2.245000 0.085000 ;
        RECT 2.555000 -0.085000 2.725000 0.085000 ;
        RECT 3.035000 -0.085000 3.205000 0.085000 ;
        RECT 3.515000 -0.085000 3.685000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.245000 3.840000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 3.245000 3.840000 3.415000 ;
        RECT 0.635000 1.820000 0.885000 3.245000 ;
        RECT 1.885000 2.290000 2.085000 3.245000 ;
      LAYER mcon ;
        RECT 0.155000 3.245000 0.325000 3.415000 ;
        RECT 0.635000 3.245000 0.805000 3.415000 ;
        RECT 1.115000 3.245000 1.285000 3.415000 ;
        RECT 1.595000 3.245000 1.765000 3.415000 ;
        RECT 2.075000 3.245000 2.245000 3.415000 ;
        RECT 2.555000 3.245000 2.725000 3.415000 ;
        RECT 3.035000 3.245000 3.205000 3.415000 ;
        RECT 3.515000 3.245000 3.685000 3.415000 ;
      LAYER met1 ;
        RECT 0.000000 3.085000 3.840000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.425000 1.400000 1.415000 1.650000 ;
      RECT 1.245000 1.110000 3.540000 1.280000 ;
      RECT 1.245000 1.280000 1.415000 1.400000 ;
      RECT 1.355000 1.950000 2.615000 2.120000 ;
      RECT 1.355000 2.120000 1.685000 2.980000 ;
      RECT 2.280000 0.840000 2.610000 1.080000 ;
      RECT 2.280000 1.080000 3.540000 1.110000 ;
      RECT 2.285000 2.120000 2.615000 2.980000 ;
      RECT 3.125000 1.280000 3.540000 2.980000 ;
  END
END sky130_fd_sc_hs__a211o_1
