* File: sky130_fd_sc_hs__o31a_1.spice
* Created: Thu Aug 27 21:02:28 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hs__o31a_1.pex.spice"
.subckt sky130_fd_sc_hs__o31a_1  VNB VPB A1 A2 A3 B1 X VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* X	X
* B1	B1
* A3	A3
* A2	A2
* A1	A1
* VPB	VPB
* VNB	VNB
MM1009 N_VGND_M1009_d N_A_84_48#_M1009_g N_X_M1009_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.166607 AS=0.2109 PD=1.25478 PS=2.05 NRD=11.34 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75002.3 A=0.111 P=1.78 MULT=1
MM1008 N_A_230_94#_M1008_d N_A1_M1008_g N_VGND_M1009_d VNB NLOWVT L=0.15 W=0.64
+ AD=0.1136 AS=0.144093 PD=0.995 PS=1.08522 NRD=0 NRS=15.468 M=1 R=4.26667
+ SA=75000.8 SB=75002 A=0.096 P=1.58 MULT=1
MM1006 N_VGND_M1006_d N_A2_M1006_g N_A_230_94#_M1008_d VNB NLOWVT L=0.15 W=0.64
+ AD=0.1824 AS=0.1136 PD=1.21 PS=0.995 NRD=28.116 NRS=14.052 M=1 R=4.26667
+ SA=75001.3 SB=75001.5 A=0.096 P=1.58 MULT=1
MM1003 N_A_230_94#_M1003_d N_A3_M1003_g N_VGND_M1006_d VNB NLOWVT L=0.15 W=0.64
+ AD=0.1104 AS=0.1824 PD=0.985 PS=1.21 NRD=12.18 NRS=26.244 M=1 R=4.26667
+ SA=75002 SB=75000.8 A=0.096 P=1.58 MULT=1
MM1004 N_A_84_48#_M1004_d N_B1_M1004_g N_A_230_94#_M1003_d VNB NLOWVT L=0.15
+ W=0.64 AD=0.2272 AS=0.1104 PD=1.99 PS=0.985 NRD=13.116 NRS=0 M=1 R=4.26667
+ SA=75002.5 SB=75000.3 A=0.096 P=1.58 MULT=1
MM1002 N_VPWR_M1002_d N_A_84_48#_M1002_g N_X_M1002_s VPB PSHORT L=0.15 W=1.12
+ AD=0.307155 AS=0.3304 PD=1.75396 PS=2.83 NRD=22.4186 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75002.2 A=0.168 P=2.54 MULT=1
MM1000 A_256_368# N_A1_M1000_g N_VPWR_M1002_d VPB PSHORT L=0.15 W=1 AD=0.135
+ AS=0.274245 PD=1.27 PS=1.56604 NRD=15.7403 NRS=26.595 M=1 R=6.66667 SA=75000.9
+ SB=75001.8 A=0.15 P=2.3 MULT=1
MM1007 A_340_368# N_A2_M1007_g A_256_368# VPB PSHORT L=0.15 W=1 AD=0.18 AS=0.135
+ PD=1.36 PS=1.27 NRD=24.6053 NRS=15.7403 M=1 R=6.66667 SA=75001.3 SB=75001.3
+ A=0.15 P=2.3 MULT=1
MM1001 N_A_84_48#_M1001_d N_A3_M1001_g A_340_368# VPB PSHORT L=0.15 W=1
+ AD=0.203696 AS=0.18 PD=1.51087 PS=1.36 NRD=1.9503 NRS=24.6053 M=1 R=6.66667
+ SA=75001.8 SB=75000.8 A=0.15 P=2.3 MULT=1
MM1005 N_VPWR_M1005_d N_B1_M1005_g N_A_84_48#_M1001_d VPB PSHORT L=0.15 W=0.84
+ AD=0.399 AS=0.171104 PD=2.63 PS=1.26913 NRD=2.3443 NRS=23.837 M=1 R=5.6
+ SA=75002.4 SB=75000.4 A=0.126 P=1.98 MULT=1
DX10_noxref VNB VPB NWDIODE A=6.9564 P=11.2
*
.include "sky130_fd_sc_hs__o31a_1.pxi.spice"
*
.ends
*
*
