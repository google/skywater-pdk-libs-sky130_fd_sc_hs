* File: sky130_fd_sc_hs__a211oi_2.pxi.spice
* Created: Tue Sep  1 19:48:47 2020
* 
x_PM_SKY130_FD_SC_HS__A211OI_2%A1 N_A1_c_79_n N_A1_M1000_g N_A1_c_75_n
+ N_A1_M1008_g N_A1_c_80_n N_A1_M1001_g N_A1_c_76_n N_A1_M1011_g A1 N_A1_c_78_n
+ PM_SKY130_FD_SC_HS__A211OI_2%A1
x_PM_SKY130_FD_SC_HS__A211OI_2%A2 N_A2_M1002_g N_A2_c_126_n N_A2_M1004_g
+ N_A2_c_127_n N_A2_M1006_g N_A2_M1005_g A2 A2 A2 N_A2_c_125_n
+ PM_SKY130_FD_SC_HS__A211OI_2%A2
x_PM_SKY130_FD_SC_HS__A211OI_2%B1 N_B1_c_178_n N_B1_M1003_g N_B1_c_181_n
+ N_B1_M1009_g N_B1_c_182_n N_B1_M1010_g B1 B1 N_B1_c_180_n
+ PM_SKY130_FD_SC_HS__A211OI_2%B1
x_PM_SKY130_FD_SC_HS__A211OI_2%C1 N_C1_c_224_n N_C1_M1007_g N_C1_c_227_n
+ N_C1_M1012_g N_C1_c_228_n N_C1_M1013_g C1 C1 N_C1_c_226_n
+ PM_SKY130_FD_SC_HS__A211OI_2%C1
x_PM_SKY130_FD_SC_HS__A211OI_2%VPWR N_VPWR_M1000_s N_VPWR_M1001_s N_VPWR_M1006_s
+ N_VPWR_c_258_n N_VPWR_c_259_n N_VPWR_c_260_n N_VPWR_c_261_n VPWR
+ N_VPWR_c_262_n N_VPWR_c_263_n N_VPWR_c_264_n N_VPWR_c_257_n N_VPWR_c_266_n
+ N_VPWR_c_267_n PM_SKY130_FD_SC_HS__A211OI_2%VPWR
x_PM_SKY130_FD_SC_HS__A211OI_2%A_114_368# N_A_114_368#_M1000_d
+ N_A_114_368#_M1004_d N_A_114_368#_M1009_d N_A_114_368#_c_317_n
+ N_A_114_368#_c_318_n N_A_114_368#_c_327_n N_A_114_368#_c_319_n
+ N_A_114_368#_c_333_n N_A_114_368#_c_320_n N_A_114_368#_c_338_n
+ N_A_114_368#_c_339_n N_A_114_368#_c_335_n N_A_114_368#_c_321_n
+ PM_SKY130_FD_SC_HS__A211OI_2%A_114_368#
x_PM_SKY130_FD_SC_HS__A211OI_2%A_497_368# N_A_497_368#_M1009_s
+ N_A_497_368#_M1010_s N_A_497_368#_M1013_s N_A_497_368#_c_366_n
+ N_A_497_368#_c_367_n N_A_497_368#_c_368_n N_A_497_368#_c_378_n
+ N_A_497_368#_c_369_n N_A_497_368#_c_370_n N_A_497_368#_c_371_n
+ PM_SKY130_FD_SC_HS__A211OI_2%A_497_368#
x_PM_SKY130_FD_SC_HS__A211OI_2%Y N_Y_M1008_d N_Y_M1003_d N_Y_M1012_d N_Y_c_468_p
+ N_Y_c_409_n N_Y_c_410_n N_Y_c_432_n N_Y_c_414_n N_Y_c_437_n N_Y_c_411_n Y Y
+ N_Y_c_412_n N_Y_c_415_n Y Y PM_SKY130_FD_SC_HS__A211OI_2%Y
x_PM_SKY130_FD_SC_HS__A211OI_2%A_38_74# N_A_38_74#_M1008_s N_A_38_74#_M1011_s
+ N_A_38_74#_M1005_d N_A_38_74#_c_486_n N_A_38_74#_c_487_n N_A_38_74#_c_488_n
+ N_A_38_74#_c_498_n N_A_38_74#_c_499_n N_A_38_74#_c_502_n N_A_38_74#_c_489_n
+ N_A_38_74#_c_490_n PM_SKY130_FD_SC_HS__A211OI_2%A_38_74#
x_PM_SKY130_FD_SC_HS__A211OI_2%VGND N_VGND_M1002_s N_VGND_M1003_s N_VGND_M1007_d
+ N_VGND_c_531_n N_VGND_c_532_n N_VGND_c_533_n N_VGND_c_534_n N_VGND_c_535_n
+ N_VGND_c_536_n N_VGND_c_537_n N_VGND_c_538_n VGND N_VGND_c_539_n
+ N_VGND_c_540_n N_VGND_c_541_n N_VGND_c_542_n PM_SKY130_FD_SC_HS__A211OI_2%VGND
cc_1 VNB N_A1_c_75_n 0.0208392f $X=-0.19 $Y=-0.245 $X2=0.53 $Y2=1.22
cc_2 VNB N_A1_c_76_n 0.0152841f $X=-0.19 $Y=-0.245 $X2=0.96 $Y2=1.22
cc_3 VNB A1 0.0221259f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_4 VNB N_A1_c_78_n 0.0814724f $X=-0.19 $Y=-0.245 $X2=0.945 $Y2=1.492
cc_5 VNB N_A2_M1002_g 0.0227439f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.4
cc_6 VNB N_A2_M1005_g 0.0274828f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_7 VNB A2 0.0102109f $X=-0.19 $Y=-0.245 $X2=0.325 $Y2=1.385
cc_8 VNB N_A2_c_125_n 0.0406811f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_B1_c_178_n 0.02217f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.765
cc_10 VNB B1 0.00938409f $X=-0.19 $Y=-0.245 $X2=0.96 $Y2=0.74
cc_11 VNB N_B1_c_180_n 0.0642394f $X=-0.19 $Y=-0.245 $X2=0.325 $Y2=1.385
cc_12 VNB N_C1_c_224_n 0.0238441f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.765
cc_13 VNB C1 0.049094f $X=-0.19 $Y=-0.245 $X2=0.96 $Y2=0.74
cc_14 VNB N_C1_c_226_n 0.0682866f $X=-0.19 $Y=-0.245 $X2=0.325 $Y2=1.385
cc_15 VNB N_VPWR_c_257_n 0.203486f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_Y_c_409_n 0.0283899f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_Y_c_410_n 9.77343e-19 $X=-0.19 $Y=-0.245 $X2=0.325 $Y2=1.492
cc_18 VNB N_Y_c_411_n 0.00657274f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_Y_c_412_n 0.00205455f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB Y 0.00994006f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_38_74#_c_486_n 0.022879f $X=-0.19 $Y=-0.245 $X2=0.96 $Y2=0.74
cc_22 VNB N_A_38_74#_c_487_n 0.00450214f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_38_74#_c_488_n 0.00975702f $X=-0.19 $Y=-0.245 $X2=0.325 $Y2=1.492
cc_24 VNB N_A_38_74#_c_489_n 0.00230074f $X=-0.19 $Y=-0.245 $X2=0.302 $Y2=1.295
cc_25 VNB N_A_38_74#_c_490_n 0.00655536f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_VGND_c_531_n 0.00523743f $X=-0.19 $Y=-0.245 $X2=0.96 $Y2=0.74
cc_27 VNB N_VGND_c_532_n 0.0102131f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_533_n 0.0344107f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.492
cc_29 VNB N_VGND_c_534_n 0.0364374f $X=-0.19 $Y=-0.245 $X2=0.96 $Y2=1.492
cc_30 VNB N_VGND_c_535_n 0.00307831f $X=-0.19 $Y=-0.245 $X2=0.302 $Y2=1.295
cc_31 VNB N_VGND_c_536_n 0.00142485f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_537_n 0.0253857f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_538_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_539_n 0.022637f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_540_n 0.0247369f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_541_n 0.302138f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_542_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VPB N_A1_c_79_n 0.0176569f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.765
cc_39 VPB N_A1_c_80_n 0.0152251f $X=-0.19 $Y=1.66 $X2=0.945 $Y2=1.765
cc_40 VPB N_A1_c_78_n 0.0165004f $X=-0.19 $Y=1.66 $X2=0.945 $Y2=1.492
cc_41 VPB N_A2_c_126_n 0.015104f $X=-0.19 $Y=1.66 $X2=0.53 $Y2=0.74
cc_42 VPB N_A2_c_127_n 0.0177914f $X=-0.19 $Y=1.66 $X2=0.945 $Y2=2.4
cc_43 VPB A2 0.0112392f $X=-0.19 $Y=1.66 $X2=0.325 $Y2=1.385
cc_44 VPB N_A2_c_125_n 0.0223461f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_45 VPB N_B1_c_181_n 0.0170299f $X=-0.19 $Y=1.66 $X2=0.53 $Y2=1.22
cc_46 VPB N_B1_c_182_n 0.0141404f $X=-0.19 $Y=1.66 $X2=0.945 $Y2=1.765
cc_47 VPB N_B1_c_180_n 0.0131907f $X=-0.19 $Y=1.66 $X2=0.325 $Y2=1.385
cc_48 VPB N_C1_c_227_n 0.0141404f $X=-0.19 $Y=1.66 $X2=0.53 $Y2=1.22
cc_49 VPB N_C1_c_228_n 0.0181207f $X=-0.19 $Y=1.66 $X2=0.945 $Y2=1.765
cc_50 VPB N_C1_c_226_n 0.0160642f $X=-0.19 $Y=1.66 $X2=0.325 $Y2=1.385
cc_51 VPB N_VPWR_c_258_n 0.0103331f $X=-0.19 $Y=1.66 $X2=0.96 $Y2=1.22
cc_52 VPB N_VPWR_c_259_n 0.0572609f $X=-0.19 $Y=1.66 $X2=0.96 $Y2=0.74
cc_53 VPB N_VPWR_c_260_n 0.00271781f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.492
cc_54 VPB N_VPWR_c_261_n 0.0110015f $X=-0.19 $Y=1.66 $X2=0.302 $Y2=1.295
cc_55 VPB N_VPWR_c_262_n 0.0185253f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_56 VPB N_VPWR_c_263_n 0.0164465f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_57 VPB N_VPWR_c_264_n 0.0631895f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_58 VPB N_VPWR_c_257_n 0.0828734f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_59 VPB N_VPWR_c_266_n 0.00601644f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_60 VPB N_VPWR_c_267_n 0.00614127f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_61 VPB N_A_114_368#_c_317_n 0.00493179f $X=-0.19 $Y=1.66 $X2=0.96 $Y2=1.22
cc_62 VPB N_A_114_368#_c_318_n 0.00216998f $X=-0.19 $Y=1.66 $X2=0.96 $Y2=0.74
cc_63 VPB N_A_114_368#_c_319_n 0.00180921f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.492
cc_64 VPB N_A_114_368#_c_320_n 0.00918628f $X=-0.19 $Y=1.66 $X2=0.302 $Y2=1.295
cc_65 VPB N_A_114_368#_c_321_n 0.0110589f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_66 VPB N_A_497_368#_c_366_n 0.00465684f $X=-0.19 $Y=1.66 $X2=0.96 $Y2=0.74
cc_67 VPB N_A_497_368#_c_367_n 0.00259172f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_68 VPB N_A_497_368#_c_368_n 0.00430699f $X=-0.19 $Y=1.66 $X2=0.325 $Y2=1.492
cc_69 VPB N_A_497_368#_c_369_n 0.0124466f $X=-0.19 $Y=1.66 $X2=0.945 $Y2=1.492
cc_70 VPB N_A_497_368#_c_370_n 0.0436631f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_71 VPB N_A_497_368#_c_371_n 0.00123754f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_72 VPB N_Y_c_414_n 0.0115233f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.492
cc_73 VPB N_Y_c_415_n 0.00179554f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_74 VPB Y 0.00118476f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_75 N_A1_c_76_n N_A2_M1002_g 0.0209092f $X=0.96 $Y=1.22 $X2=0 $Y2=0
cc_76 N_A1_c_80_n N_A2_c_126_n 0.0248293f $X=0.945 $Y=1.765 $X2=0 $Y2=0
cc_77 N_A1_c_80_n A2 4.36825e-19 $X=0.945 $Y=1.765 $X2=0 $Y2=0
cc_78 A1 A2 0.00383248f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_79 N_A1_c_78_n A2 0.00867206f $X=0.945 $Y=1.492 $X2=0 $Y2=0
cc_80 N_A1_c_78_n N_A2_c_125_n 0.0258954f $X=0.945 $Y=1.492 $X2=0 $Y2=0
cc_81 N_A1_c_79_n N_VPWR_c_259_n 0.00877831f $X=0.495 $Y=1.765 $X2=0 $Y2=0
cc_82 A1 N_VPWR_c_259_n 0.0139183f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_83 N_A1_c_78_n N_VPWR_c_259_n 0.00145147f $X=0.945 $Y=1.492 $X2=0 $Y2=0
cc_84 N_A1_c_79_n N_VPWR_c_260_n 5.66285e-19 $X=0.495 $Y=1.765 $X2=0 $Y2=0
cc_85 N_A1_c_80_n N_VPWR_c_260_n 0.011741f $X=0.945 $Y=1.765 $X2=0 $Y2=0
cc_86 N_A1_c_79_n N_VPWR_c_262_n 0.00445602f $X=0.495 $Y=1.765 $X2=0 $Y2=0
cc_87 N_A1_c_80_n N_VPWR_c_262_n 0.00413917f $X=0.945 $Y=1.765 $X2=0 $Y2=0
cc_88 N_A1_c_79_n N_VPWR_c_257_n 0.0086105f $X=0.495 $Y=1.765 $X2=0 $Y2=0
cc_89 N_A1_c_80_n N_VPWR_c_257_n 0.00817726f $X=0.945 $Y=1.765 $X2=0 $Y2=0
cc_90 N_A1_c_79_n N_A_114_368#_c_317_n 0.00420119f $X=0.495 $Y=1.765 $X2=0 $Y2=0
cc_91 N_A1_c_80_n N_A_114_368#_c_317_n 0.00285814f $X=0.945 $Y=1.765 $X2=0 $Y2=0
cc_92 N_A1_c_78_n N_A_114_368#_c_317_n 0.00317782f $X=0.945 $Y=1.492 $X2=0 $Y2=0
cc_93 N_A1_c_79_n N_A_114_368#_c_318_n 0.0100425f $X=0.495 $Y=1.765 $X2=0 $Y2=0
cc_94 N_A1_c_80_n N_A_114_368#_c_318_n 0.00627629f $X=0.945 $Y=1.765 $X2=0 $Y2=0
cc_95 N_A1_c_80_n N_A_114_368#_c_327_n 0.0171849f $X=0.945 $Y=1.765 $X2=0 $Y2=0
cc_96 N_A1_c_76_n N_Y_c_409_n 0.00842504f $X=0.96 $Y=1.22 $X2=0 $Y2=0
cc_97 N_A1_c_78_n N_Y_c_409_n 0.0101657f $X=0.945 $Y=1.492 $X2=0 $Y2=0
cc_98 N_A1_c_75_n N_Y_c_410_n 0.00262654f $X=0.53 $Y=1.22 $X2=0 $Y2=0
cc_99 A1 N_Y_c_410_n 0.00656158f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_100 N_A1_c_78_n N_Y_c_410_n 0.00850071f $X=0.945 $Y=1.492 $X2=0 $Y2=0
cc_101 N_A1_c_75_n N_A_38_74#_c_486_n 0.00776833f $X=0.53 $Y=1.22 $X2=0 $Y2=0
cc_102 N_A1_c_76_n N_A_38_74#_c_486_n 6.58694e-19 $X=0.96 $Y=1.22 $X2=0 $Y2=0
cc_103 A1 N_A_38_74#_c_486_n 0.0260993f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_104 N_A1_c_78_n N_A_38_74#_c_486_n 0.00193135f $X=0.945 $Y=1.492 $X2=0 $Y2=0
cc_105 N_A1_c_75_n N_A_38_74#_c_487_n 0.0100245f $X=0.53 $Y=1.22 $X2=0 $Y2=0
cc_106 N_A1_c_76_n N_A_38_74#_c_487_n 0.00969779f $X=0.96 $Y=1.22 $X2=0 $Y2=0
cc_107 N_A1_c_75_n N_A_38_74#_c_488_n 0.00282152f $X=0.53 $Y=1.22 $X2=0 $Y2=0
cc_108 N_A1_c_76_n N_A_38_74#_c_498_n 0.00211217f $X=0.96 $Y=1.22 $X2=0 $Y2=0
cc_109 N_A1_c_75_n N_A_38_74#_c_499_n 5.88012e-19 $X=0.53 $Y=1.22 $X2=0 $Y2=0
cc_110 N_A1_c_76_n N_A_38_74#_c_499_n 0.00482477f $X=0.96 $Y=1.22 $X2=0 $Y2=0
cc_111 N_A1_c_75_n N_VGND_c_534_n 0.00278247f $X=0.53 $Y=1.22 $X2=0 $Y2=0
cc_112 N_A1_c_76_n N_VGND_c_534_n 0.00278247f $X=0.96 $Y=1.22 $X2=0 $Y2=0
cc_113 N_A1_c_75_n N_VGND_c_541_n 0.00357198f $X=0.53 $Y=1.22 $X2=0 $Y2=0
cc_114 N_A1_c_76_n N_VGND_c_541_n 0.00353524f $X=0.96 $Y=1.22 $X2=0 $Y2=0
cc_115 A2 N_B1_c_180_n 9.22828e-19 $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_116 N_A2_c_126_n N_VPWR_c_260_n 0.0116098f $X=1.395 $Y=1.765 $X2=0 $Y2=0
cc_117 N_A2_c_127_n N_VPWR_c_260_n 5.35985e-19 $X=1.845 $Y=1.765 $X2=0 $Y2=0
cc_118 N_A2_c_126_n N_VPWR_c_261_n 5.02548e-19 $X=1.395 $Y=1.765 $X2=0 $Y2=0
cc_119 N_A2_c_127_n N_VPWR_c_261_n 0.0109013f $X=1.845 $Y=1.765 $X2=0 $Y2=0
cc_120 N_A2_c_126_n N_VPWR_c_263_n 0.00413917f $X=1.395 $Y=1.765 $X2=0 $Y2=0
cc_121 N_A2_c_127_n N_VPWR_c_263_n 0.00413917f $X=1.845 $Y=1.765 $X2=0 $Y2=0
cc_122 N_A2_c_126_n N_VPWR_c_257_n 0.00817726f $X=1.395 $Y=1.765 $X2=0 $Y2=0
cc_123 N_A2_c_127_n N_VPWR_c_257_n 0.00817726f $X=1.845 $Y=1.765 $X2=0 $Y2=0
cc_124 N_A2_c_126_n N_A_114_368#_c_327_n 0.0126342f $X=1.395 $Y=1.765 $X2=0
+ $Y2=0
cc_125 A2 N_A_114_368#_c_327_n 0.0300496f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_126 N_A2_c_125_n N_A_114_368#_c_327_n 4.42778e-19 $X=1.845 $Y=1.557 $X2=0
+ $Y2=0
cc_127 N_A2_c_126_n N_A_114_368#_c_319_n 0.0034769f $X=1.395 $Y=1.765 $X2=0
+ $Y2=0
cc_128 N_A2_c_127_n N_A_114_368#_c_319_n 0.00526412f $X=1.845 $Y=1.765 $X2=0
+ $Y2=0
cc_129 N_A2_c_127_n N_A_114_368#_c_333_n 0.0189628f $X=1.845 $Y=1.765 $X2=0
+ $Y2=0
cc_130 A2 N_A_114_368#_c_333_n 0.0407594f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_131 A2 N_A_114_368#_c_335_n 0.0148009f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_132 N_A2_c_125_n N_A_114_368#_c_335_n 0.00104579f $X=1.845 $Y=1.557 $X2=0
+ $Y2=0
cc_133 N_A2_c_127_n N_A_497_368#_c_368_n 5.94256e-19 $X=1.845 $Y=1.765 $X2=0
+ $Y2=0
cc_134 N_A2_M1002_g N_Y_c_409_n 0.010666f $X=1.39 $Y=0.74 $X2=0 $Y2=0
cc_135 N_A2_M1005_g N_Y_c_409_n 0.0127668f $X=1.86 $Y=0.74 $X2=0 $Y2=0
cc_136 A2 N_Y_c_409_n 0.0907992f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_137 N_A2_c_125_n N_Y_c_409_n 0.00518776f $X=1.845 $Y=1.557 $X2=0 $Y2=0
cc_138 N_A2_M1005_g N_Y_c_412_n 0.00261336f $X=1.86 $Y=0.74 $X2=0 $Y2=0
cc_139 N_A2_c_127_n N_Y_c_415_n 0.00295863f $X=1.845 $Y=1.765 $X2=0 $Y2=0
cc_140 A2 N_Y_c_415_n 0.00421358f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_141 N_A2_M1005_g Y 0.0042677f $X=1.86 $Y=0.74 $X2=0 $Y2=0
cc_142 A2 Y 0.0189927f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_143 N_A2_c_125_n Y 0.00101046f $X=1.845 $Y=1.557 $X2=0 $Y2=0
cc_144 N_A2_M1002_g N_A_38_74#_c_487_n 9.71323e-19 $X=1.39 $Y=0.74 $X2=0 $Y2=0
cc_145 N_A2_M1002_g N_A_38_74#_c_502_n 0.0100656f $X=1.39 $Y=0.74 $X2=0 $Y2=0
cc_146 N_A2_M1005_g N_A_38_74#_c_502_n 0.0100792f $X=1.86 $Y=0.74 $X2=0 $Y2=0
cc_147 N_A2_M1005_g N_A_38_74#_c_490_n 9.08649e-19 $X=1.86 $Y=0.74 $X2=0 $Y2=0
cc_148 N_A2_M1002_g N_VGND_c_531_n 0.00236272f $X=1.39 $Y=0.74 $X2=0 $Y2=0
cc_149 N_A2_M1005_g N_VGND_c_531_n 0.00186481f $X=1.86 $Y=0.74 $X2=0 $Y2=0
cc_150 N_A2_M1005_g N_VGND_c_532_n 0.00282671f $X=1.86 $Y=0.74 $X2=0 $Y2=0
cc_151 N_A2_M1002_g N_VGND_c_534_n 0.00281141f $X=1.39 $Y=0.74 $X2=0 $Y2=0
cc_152 N_A2_M1002_g N_VGND_c_536_n 0.00347646f $X=1.39 $Y=0.74 $X2=0 $Y2=0
cc_153 N_A2_M1005_g N_VGND_c_536_n 0.00378394f $X=1.86 $Y=0.74 $X2=0 $Y2=0
cc_154 N_A2_M1005_g N_VGND_c_539_n 0.00329872f $X=1.86 $Y=0.74 $X2=0 $Y2=0
cc_155 N_A2_M1002_g N_VGND_c_541_n 0.00365164f $X=1.39 $Y=0.74 $X2=0 $Y2=0
cc_156 N_A2_M1005_g N_VGND_c_541_n 0.00433324f $X=1.86 $Y=0.74 $X2=0 $Y2=0
cc_157 N_B1_c_178_n N_C1_c_224_n 0.00764828f $X=2.84 $Y=1.22 $X2=-0.19
+ $Y2=-0.245
cc_158 B1 N_C1_c_224_n 0.00527496f $X=3.515 $Y=1.21 $X2=-0.19 $Y2=-0.245
cc_159 N_B1_c_182_n N_C1_c_227_n 0.0228756f $X=3.305 $Y=1.765 $X2=0 $Y2=0
cc_160 B1 C1 0.0231228f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_161 B1 N_C1_c_226_n 0.0122116f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_162 N_B1_c_180_n N_C1_c_226_n 0.032889f $X=3.26 $Y=1.385 $X2=0 $Y2=0
cc_163 N_B1_c_181_n N_VPWR_c_261_n 0.0017223f $X=2.855 $Y=1.765 $X2=0 $Y2=0
cc_164 N_B1_c_181_n N_VPWR_c_264_n 0.00278257f $X=2.855 $Y=1.765 $X2=0 $Y2=0
cc_165 N_B1_c_182_n N_VPWR_c_264_n 0.00278271f $X=3.305 $Y=1.765 $X2=0 $Y2=0
cc_166 N_B1_c_181_n N_VPWR_c_257_n 0.00358623f $X=2.855 $Y=1.765 $X2=0 $Y2=0
cc_167 N_B1_c_182_n N_VPWR_c_257_n 0.00353907f $X=3.305 $Y=1.765 $X2=0 $Y2=0
cc_168 N_B1_c_181_n N_A_114_368#_c_320_n 0.012519f $X=2.855 $Y=1.765 $X2=0 $Y2=0
cc_169 N_B1_c_182_n N_A_114_368#_c_338_n 0.00192129f $X=3.305 $Y=1.765 $X2=0
+ $Y2=0
cc_170 N_B1_c_182_n N_A_114_368#_c_339_n 0.00566256f $X=3.305 $Y=1.765 $X2=0
+ $Y2=0
cc_171 N_B1_c_181_n N_A_114_368#_c_321_n 0.00342267f $X=2.855 $Y=1.765 $X2=0
+ $Y2=0
cc_172 N_B1_c_181_n N_A_497_368#_c_366_n 0.00651743f $X=2.855 $Y=1.765 $X2=0
+ $Y2=0
cc_173 N_B1_c_182_n N_A_497_368#_c_366_n 4.50629e-19 $X=3.305 $Y=1.765 $X2=0
+ $Y2=0
cc_174 N_B1_c_181_n N_A_497_368#_c_367_n 0.00879888f $X=2.855 $Y=1.765 $X2=0
+ $Y2=0
cc_175 N_B1_c_182_n N_A_497_368#_c_367_n 0.0128006f $X=3.305 $Y=1.765 $X2=0
+ $Y2=0
cc_176 N_B1_c_181_n N_A_497_368#_c_368_n 0.00262441f $X=2.855 $Y=1.765 $X2=0
+ $Y2=0
cc_177 N_B1_c_182_n N_A_497_368#_c_378_n 0.00443298f $X=3.305 $Y=1.765 $X2=0
+ $Y2=0
cc_178 N_B1_c_178_n N_Y_c_432_n 0.0151832f $X=2.84 $Y=1.22 $X2=0 $Y2=0
cc_179 N_B1_c_181_n N_Y_c_414_n 0.00773257f $X=2.855 $Y=1.765 $X2=0 $Y2=0
cc_180 N_B1_c_182_n N_Y_c_414_n 0.0109522f $X=3.305 $Y=1.765 $X2=0 $Y2=0
cc_181 B1 N_Y_c_414_n 0.0538531f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_182 N_B1_c_180_n N_Y_c_414_n 0.0178899f $X=3.26 $Y=1.385 $X2=0 $Y2=0
cc_183 N_B1_c_182_n N_Y_c_437_n 9.44162e-19 $X=3.305 $Y=1.765 $X2=0 $Y2=0
cc_184 N_B1_c_178_n N_Y_c_411_n 8.86064e-19 $X=2.84 $Y=1.22 $X2=0 $Y2=0
cc_185 B1 N_Y_c_411_n 0.0505593f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_186 N_B1_c_180_n N_Y_c_411_n 0.00472374f $X=3.26 $Y=1.385 $X2=0 $Y2=0
cc_187 N_B1_c_178_n N_Y_c_412_n 0.00783386f $X=2.84 $Y=1.22 $X2=0 $Y2=0
cc_188 B1 N_Y_c_412_n 0.005464f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_189 B1 Y 0.0176772f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_190 N_B1_c_180_n Y 0.0168492f $X=3.26 $Y=1.385 $X2=0 $Y2=0
cc_191 N_B1_c_178_n N_A_38_74#_c_489_n 0.00298356f $X=2.84 $Y=1.22 $X2=0 $Y2=0
cc_192 N_B1_c_178_n N_A_38_74#_c_490_n 0.00172044f $X=2.84 $Y=1.22 $X2=0 $Y2=0
cc_193 N_B1_c_178_n N_VGND_c_532_n 0.010855f $X=2.84 $Y=1.22 $X2=0 $Y2=0
cc_194 N_B1_c_178_n N_VGND_c_537_n 0.00383152f $X=2.84 $Y=1.22 $X2=0 $Y2=0
cc_195 N_B1_c_178_n N_VGND_c_541_n 0.00386893f $X=2.84 $Y=1.22 $X2=0 $Y2=0
cc_196 N_C1_c_227_n N_VPWR_c_264_n 0.00278271f $X=3.755 $Y=1.765 $X2=0 $Y2=0
cc_197 N_C1_c_228_n N_VPWR_c_264_n 0.00278271f $X=4.205 $Y=1.765 $X2=0 $Y2=0
cc_198 N_C1_c_227_n N_VPWR_c_257_n 0.00353907f $X=3.755 $Y=1.765 $X2=0 $Y2=0
cc_199 N_C1_c_228_n N_VPWR_c_257_n 0.00357579f $X=4.205 $Y=1.765 $X2=0 $Y2=0
cc_200 N_C1_c_227_n N_A_497_368#_c_378_n 0.0062909f $X=3.755 $Y=1.765 $X2=0
+ $Y2=0
cc_201 N_C1_c_227_n N_A_497_368#_c_369_n 0.0128006f $X=3.755 $Y=1.765 $X2=0
+ $Y2=0
cc_202 N_C1_c_228_n N_A_497_368#_c_369_n 0.0136604f $X=4.205 $Y=1.765 $X2=0
+ $Y2=0
cc_203 N_C1_c_228_n N_A_497_368#_c_370_n 0.00807045f $X=4.205 $Y=1.765 $X2=0
+ $Y2=0
cc_204 C1 N_A_497_368#_c_370_n 0.0160108f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_205 N_C1_c_227_n N_Y_c_414_n 0.0100928f $X=3.755 $Y=1.765 $X2=0 $Y2=0
cc_206 N_C1_c_228_n N_Y_c_414_n 0.00418463f $X=4.205 $Y=1.765 $X2=0 $Y2=0
cc_207 C1 N_Y_c_414_n 0.0151664f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_208 N_C1_c_226_n N_Y_c_414_n 0.0158572f $X=4.13 $Y=1.385 $X2=0 $Y2=0
cc_209 N_C1_c_227_n N_Y_c_437_n 0.0100465f $X=3.755 $Y=1.765 $X2=0 $Y2=0
cc_210 N_C1_c_228_n N_Y_c_437_n 0.00925235f $X=4.205 $Y=1.765 $X2=0 $Y2=0
cc_211 N_C1_c_224_n N_Y_c_411_n 0.00641f $X=3.71 $Y=1.22 $X2=0 $Y2=0
cc_212 N_C1_c_224_n N_VGND_c_533_n 0.0153376f $X=3.71 $Y=1.22 $X2=0 $Y2=0
cc_213 C1 N_VGND_c_533_n 0.0108734f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_214 N_C1_c_226_n N_VGND_c_533_n 0.00776363f $X=4.13 $Y=1.385 $X2=0 $Y2=0
cc_215 N_C1_c_224_n N_VGND_c_537_n 0.00383152f $X=3.71 $Y=1.22 $X2=0 $Y2=0
cc_216 N_C1_c_224_n N_VGND_c_541_n 0.00760466f $X=3.71 $Y=1.22 $X2=0 $Y2=0
cc_217 N_VPWR_c_259_n N_A_114_368#_c_317_n 0.0207081f $X=0.27 $Y=1.985 $X2=0
+ $Y2=0
cc_218 N_VPWR_c_259_n N_A_114_368#_c_318_n 0.0564818f $X=0.27 $Y=1.985 $X2=0
+ $Y2=0
cc_219 N_VPWR_c_260_n N_A_114_368#_c_318_n 0.0462948f $X=1.17 $Y=2.375 $X2=0
+ $Y2=0
cc_220 N_VPWR_c_262_n N_A_114_368#_c_318_n 0.0110241f $X=1.005 $Y=3.33 $X2=0
+ $Y2=0
cc_221 N_VPWR_c_257_n N_A_114_368#_c_318_n 0.00909194f $X=4.56 $Y=3.33 $X2=0
+ $Y2=0
cc_222 N_VPWR_M1001_s N_A_114_368#_c_327_n 0.00414387f $X=1.02 $Y=1.84 $X2=0
+ $Y2=0
cc_223 N_VPWR_c_260_n N_A_114_368#_c_327_n 0.0171814f $X=1.17 $Y=2.375 $X2=0
+ $Y2=0
cc_224 N_VPWR_c_260_n N_A_114_368#_c_319_n 0.0449718f $X=1.17 $Y=2.375 $X2=0
+ $Y2=0
cc_225 N_VPWR_c_261_n N_A_114_368#_c_319_n 0.0378067f $X=2.07 $Y=2.485 $X2=0
+ $Y2=0
cc_226 N_VPWR_c_263_n N_A_114_368#_c_319_n 0.00749631f $X=1.905 $Y=3.33 $X2=0
+ $Y2=0
cc_227 N_VPWR_c_257_n N_A_114_368#_c_319_n 0.0062048f $X=4.56 $Y=3.33 $X2=0
+ $Y2=0
cc_228 N_VPWR_M1006_s N_A_114_368#_c_333_n 0.00687715f $X=1.92 $Y=1.84 $X2=0
+ $Y2=0
cc_229 N_VPWR_c_261_n N_A_114_368#_c_333_n 0.0227209f $X=2.07 $Y=2.485 $X2=0
+ $Y2=0
cc_230 N_VPWR_c_261_n N_A_497_368#_c_366_n 0.0340127f $X=2.07 $Y=2.485 $X2=0
+ $Y2=0
cc_231 N_VPWR_c_264_n N_A_497_368#_c_367_n 0.0409869f $X=4.56 $Y=3.33 $X2=0
+ $Y2=0
cc_232 N_VPWR_c_257_n N_A_497_368#_c_367_n 0.0231342f $X=4.56 $Y=3.33 $X2=0
+ $Y2=0
cc_233 N_VPWR_c_261_n N_A_497_368#_c_368_n 0.0121617f $X=2.07 $Y=2.485 $X2=0
+ $Y2=0
cc_234 N_VPWR_c_264_n N_A_497_368#_c_368_n 0.0235908f $X=4.56 $Y=3.33 $X2=0
+ $Y2=0
cc_235 N_VPWR_c_257_n N_A_497_368#_c_368_n 0.0127585f $X=4.56 $Y=3.33 $X2=0
+ $Y2=0
cc_236 N_VPWR_c_264_n N_A_497_368#_c_369_n 0.0640155f $X=4.56 $Y=3.33 $X2=0
+ $Y2=0
cc_237 N_VPWR_c_257_n N_A_497_368#_c_369_n 0.0357926f $X=4.56 $Y=3.33 $X2=0
+ $Y2=0
cc_238 N_VPWR_c_264_n N_A_497_368#_c_371_n 0.0121867f $X=4.56 $Y=3.33 $X2=0
+ $Y2=0
cc_239 N_VPWR_c_257_n N_A_497_368#_c_371_n 0.00660921f $X=4.56 $Y=3.33 $X2=0
+ $Y2=0
cc_240 N_A_114_368#_c_320_n N_A_497_368#_M1009_s 0.00723035f $X=2.965 $Y=2.145
+ $X2=-0.19 $Y2=1.66
cc_241 N_A_114_368#_c_320_n N_A_497_368#_c_366_n 0.0219791f $X=2.965 $Y=2.145
+ $X2=0 $Y2=0
cc_242 N_A_114_368#_M1009_d N_A_497_368#_c_367_n 0.00197722f $X=2.93 $Y=1.84
+ $X2=0 $Y2=0
cc_243 N_A_114_368#_c_320_n N_A_497_368#_c_367_n 0.00286566f $X=2.965 $Y=2.145
+ $X2=0 $Y2=0
cc_244 N_A_114_368#_c_339_n N_A_497_368#_c_367_n 0.0151087f $X=3.08 $Y=2.57
+ $X2=0 $Y2=0
cc_245 N_A_114_368#_c_338_n N_A_497_368#_c_378_n 0.0117758f $X=3.105 $Y=2.23
+ $X2=0 $Y2=0
cc_246 N_A_114_368#_c_339_n N_A_497_368#_c_378_n 0.0324485f $X=3.08 $Y=2.57
+ $X2=0 $Y2=0
cc_247 N_A_114_368#_c_317_n N_Y_c_410_n 0.00556109f $X=0.68 $Y=2.12 $X2=0 $Y2=0
cc_248 N_A_114_368#_M1009_d N_Y_c_414_n 0.00197722f $X=2.93 $Y=1.84 $X2=0 $Y2=0
cc_249 N_A_114_368#_c_320_n N_Y_c_414_n 0.0101332f $X=2.965 $Y=2.145 $X2=0 $Y2=0
cc_250 N_A_114_368#_c_338_n N_Y_c_414_n 0.0162234f $X=3.105 $Y=2.23 $X2=0 $Y2=0
cc_251 N_A_114_368#_c_320_n N_Y_c_415_n 0.016109f $X=2.965 $Y=2.145 $X2=0 $Y2=0
cc_252 N_A_497_368#_c_369_n N_Y_M1012_d 0.00197722f $X=4.345 $Y=2.99 $X2=0 $Y2=0
cc_253 N_A_497_368#_M1010_s N_Y_c_414_n 0.00247267f $X=3.38 $Y=1.84 $X2=0 $Y2=0
cc_254 N_A_497_368#_c_378_n N_Y_c_414_n 0.0136682f $X=3.53 $Y=2.225 $X2=0 $Y2=0
cc_255 N_A_497_368#_c_370_n N_Y_c_414_n 0.00501285f $X=4.43 $Y=1.985 $X2=0 $Y2=0
cc_256 N_A_497_368#_c_378_n N_Y_c_437_n 0.0439674f $X=3.53 $Y=2.225 $X2=0 $Y2=0
cc_257 N_A_497_368#_c_369_n N_Y_c_437_n 0.0160777f $X=4.345 $Y=2.99 $X2=0 $Y2=0
cc_258 N_A_497_368#_c_370_n N_Y_c_437_n 0.0566253f $X=4.43 $Y=1.985 $X2=0 $Y2=0
cc_259 N_A_497_368#_M1009_s N_Y_c_415_n 0.00335686f $X=2.485 $Y=1.84 $X2=0 $Y2=0
cc_260 N_Y_c_409_n N_A_38_74#_M1011_s 0.00176461f $X=2.525 $Y=1.175 $X2=0 $Y2=0
cc_261 N_Y_c_409_n N_A_38_74#_M1005_d 0.00265093f $X=2.525 $Y=1.175 $X2=0 $Y2=0
cc_262 N_Y_M1008_d N_A_38_74#_c_487_n 0.00193374f $X=0.605 $Y=0.37 $X2=0 $Y2=0
cc_263 N_Y_c_468_p N_A_38_74#_c_487_n 0.0104673f $X=0.745 $Y=0.8 $X2=0 $Y2=0
cc_264 N_Y_c_409_n N_A_38_74#_c_487_n 0.00270072f $X=2.525 $Y=1.175 $X2=0 $Y2=0
cc_265 N_Y_c_409_n N_A_38_74#_c_498_n 0.0153397f $X=2.525 $Y=1.175 $X2=0 $Y2=0
cc_266 N_Y_c_409_n N_A_38_74#_c_502_n 0.0352288f $X=2.525 $Y=1.175 $X2=0 $Y2=0
cc_267 N_Y_c_409_n N_A_38_74#_c_489_n 0.0199765f $X=2.525 $Y=1.175 $X2=0 $Y2=0
cc_268 N_Y_c_412_n N_A_38_74#_c_489_n 0.00424281f $X=2.64 $Y=1.26 $X2=0 $Y2=0
cc_269 N_Y_c_409_n N_VGND_M1002_s 0.00219516f $X=2.525 $Y=1.175 $X2=-0.19
+ $Y2=-0.245
cc_270 N_Y_c_409_n N_VGND_M1003_s 4.19828e-19 $X=2.525 $Y=1.175 $X2=0 $Y2=0
cc_271 N_Y_c_412_n N_VGND_M1003_s 0.00661954f $X=2.64 $Y=1.26 $X2=0 $Y2=0
cc_272 N_Y_c_409_n N_VGND_c_532_n 0.00278236f $X=2.525 $Y=1.175 $X2=0 $Y2=0
cc_273 N_Y_c_432_n N_VGND_c_532_n 0.00174615f $X=2.96 $Y=0.925 $X2=0 $Y2=0
cc_274 N_Y_c_411_n N_VGND_c_532_n 0.0145467f $X=3.425 $Y=0.495 $X2=0 $Y2=0
cc_275 N_Y_c_412_n N_VGND_c_532_n 0.0135866f $X=2.64 $Y=1.26 $X2=0 $Y2=0
cc_276 N_Y_c_411_n N_VGND_c_533_n 0.0273043f $X=3.425 $Y=0.495 $X2=0 $Y2=0
cc_277 N_Y_c_411_n N_VGND_c_537_n 0.0304615f $X=3.425 $Y=0.495 $X2=0 $Y2=0
cc_278 N_Y_c_432_n N_VGND_c_541_n 0.0050789f $X=2.96 $Y=0.925 $X2=0 $Y2=0
cc_279 N_Y_c_411_n N_VGND_c_541_n 0.0234693f $X=3.425 $Y=0.495 $X2=0 $Y2=0
cc_280 N_Y_c_412_n N_VGND_c_541_n 6.18724e-19 $X=2.64 $Y=1.26 $X2=0 $Y2=0
cc_281 N_A_38_74#_c_502_n N_VGND_M1002_s 0.00413472f $X=1.99 $Y=0.835 $X2=-0.19
+ $Y2=-0.245
cc_282 N_A_38_74#_c_487_n N_VGND_c_531_n 0.00579606f $X=1.01 $Y=0.34 $X2=0 $Y2=0
cc_283 N_A_38_74#_c_490_n N_VGND_c_532_n 0.0231522f $X=2.075 $Y=0.495 $X2=0
+ $Y2=0
cc_284 N_A_38_74#_c_487_n N_VGND_c_534_n 0.0511653f $X=1.01 $Y=0.34 $X2=0 $Y2=0
cc_285 N_A_38_74#_c_488_n N_VGND_c_534_n 0.0235688f $X=0.48 $Y=0.34 $X2=0 $Y2=0
cc_286 N_A_38_74#_c_502_n N_VGND_c_534_n 0.00197156f $X=1.99 $Y=0.835 $X2=0
+ $Y2=0
cc_287 N_A_38_74#_c_487_n N_VGND_c_536_n 0.00517005f $X=1.01 $Y=0.34 $X2=0 $Y2=0
cc_288 N_A_38_74#_c_502_n N_VGND_c_536_n 0.0181541f $X=1.99 $Y=0.835 $X2=0 $Y2=0
cc_289 N_A_38_74#_c_490_n N_VGND_c_536_n 0.0105553f $X=2.075 $Y=0.495 $X2=0
+ $Y2=0
cc_290 N_A_38_74#_c_502_n N_VGND_c_539_n 0.00197884f $X=1.99 $Y=0.835 $X2=0
+ $Y2=0
cc_291 N_A_38_74#_c_490_n N_VGND_c_539_n 0.011905f $X=2.075 $Y=0.495 $X2=0 $Y2=0
cc_292 N_A_38_74#_c_487_n N_VGND_c_541_n 0.0283816f $X=1.01 $Y=0.34 $X2=0 $Y2=0
cc_293 N_A_38_74#_c_488_n N_VGND_c_541_n 0.0127152f $X=0.48 $Y=0.34 $X2=0 $Y2=0
cc_294 N_A_38_74#_c_502_n N_VGND_c_541_n 0.00846746f $X=1.99 $Y=0.835 $X2=0
+ $Y2=0
cc_295 N_A_38_74#_c_490_n N_VGND_c_541_n 0.00922555f $X=2.075 $Y=0.495 $X2=0
+ $Y2=0
