* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hs__a2111oi_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
X0 Y D1 a_29_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X1 Y B1 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X2 a_853_368# B1 a_474_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X3 VPWR A2 a_853_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X4 VGND A2 a_1228_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X5 Y D1 a_29_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X6 a_474_368# B1 a_853_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X7 a_474_368# C1 a_29_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X8 a_853_368# B1 a_474_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X9 a_474_368# C1 a_29_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X10 a_853_368# A1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X11 a_1228_74# A2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X12 VGND D1 Y VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X13 a_853_368# A1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X14 a_29_368# D1 Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X15 a_853_368# A2 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X16 a_853_368# A2 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X17 VGND C1 Y VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X18 a_1228_74# A1 Y VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X19 a_29_368# D1 Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X20 Y D1 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X21 a_29_368# C1 a_474_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X22 a_1228_74# A1 Y VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X23 a_29_368# C1 a_474_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X24 Y C1 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X25 a_474_368# B1 a_853_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X26 VGND B1 Y VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X27 Y A1 a_1228_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X28 VPWR A1 a_853_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X29 a_1228_74# A2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X30 VPWR A1 a_853_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X31 VGND A2 a_1228_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X32 Y A1 a_1228_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X33 VPWR A2 a_853_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
.ends
