/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */

`ifndef SKY130_FD_SC_HS__A2BB2O_TB_V
`define SKY130_FD_SC_HS__A2BB2O_TB_V

/**
 * a2bb2o: 2-input AND, both inputs inverted, into first input, and
 *         2-input AND into 2nd input of 2-input OR.
 *
 *         X = ((!A1 & !A2) | (B1 & B2))
 *
 * Autogenerated test bench.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none

`include "sky130_fd_sc_hs__a2bb2o.v"

module top();

    // Inputs are registered
    reg A1_N;
    reg A2_N;
    reg B1;
    reg B2;
    reg VPWR;
    reg VGND;

    // Outputs are wires
    wire X;

    initial
    begin
        // Initial state is x for all inputs.
        A1_N = 1'bX;
        A2_N = 1'bX;
        B1   = 1'bX;
        B2   = 1'bX;
        VGND = 1'bX;
        VPWR = 1'bX;

        #20   A1_N = 1'b0;
        #40   A2_N = 1'b0;
        #60   B1   = 1'b0;
        #80   B2   = 1'b0;
        #100  VGND = 1'b0;
        #120  VPWR = 1'b0;
        #140  A1_N = 1'b1;
        #160  A2_N = 1'b1;
        #180  B1   = 1'b1;
        #200  B2   = 1'b1;
        #220  VGND = 1'b1;
        #240  VPWR = 1'b1;
        #260  A1_N = 1'b0;
        #280  A2_N = 1'b0;
        #300  B1   = 1'b0;
        #320  B2   = 1'b0;
        #340  VGND = 1'b0;
        #360  VPWR = 1'b0;
        #380  VPWR = 1'b1;
        #400  VGND = 1'b1;
        #420  B2   = 1'b1;
        #440  B1   = 1'b1;
        #460  A2_N = 1'b1;
        #480  A1_N = 1'b1;
        #500  VPWR = 1'bx;
        #520  VGND = 1'bx;
        #540  B2   = 1'bx;
        #560  B1   = 1'bx;
        #580  A2_N = 1'bx;
        #600  A1_N = 1'bx;
    end

    sky130_fd_sc_hs__a2bb2o dut (.A1_N(A1_N), .A2_N(A2_N), .B1(B1), .B2(B2), .VPWR(VPWR), .VGND(VGND), .X(X));

endmodule

`default_nettype wire
`endif  // SKY130_FD_SC_HS__A2BB2O_TB_V
