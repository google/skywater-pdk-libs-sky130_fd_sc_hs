/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */

`ifndef SKY130_FD_SC_HS__SDFXBP_TB_V
`define SKY130_FD_SC_HS__SDFXBP_TB_V

/**
 * sdfxbp: Scan delay flop, non-inverted clock, complementary outputs.
 *
 * Autogenerated test bench.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none

`include "sky130_fd_sc_hs__sdfxbp.v"

module top();

    // Inputs are registered
    reg D;
    reg SCD;
    reg SCE;
    reg VPWR;
    reg VGND;

    // Outputs are wires
    wire Q;
    wire Q_N;

    initial
    begin
        // Initial state is x for all inputs.
        D    = 1'bX;
        SCD  = 1'bX;
        SCE  = 1'bX;
        VGND = 1'bX;
        VPWR = 1'bX;

        #20   D    = 1'b0;
        #40   SCD  = 1'b0;
        #60   SCE  = 1'b0;
        #80   VGND = 1'b0;
        #100  VPWR = 1'b0;
        #120  D    = 1'b1;
        #140  SCD  = 1'b1;
        #160  SCE  = 1'b1;
        #180  VGND = 1'b1;
        #200  VPWR = 1'b1;
        #220  D    = 1'b0;
        #240  SCD  = 1'b0;
        #260  SCE  = 1'b0;
        #280  VGND = 1'b0;
        #300  VPWR = 1'b0;
        #320  VPWR = 1'b1;
        #340  VGND = 1'b1;
        #360  SCE  = 1'b1;
        #380  SCD  = 1'b1;
        #400  D    = 1'b1;
        #420  VPWR = 1'bx;
        #440  VGND = 1'bx;
        #460  SCE  = 1'bx;
        #480  SCD  = 1'bx;
        #500  D    = 1'bx;
    end

    // Create a clock
    reg CLK;
    initial
    begin
        CLK = 1'b0;
    end

    always
    begin
        #5 CLK = ~CLK;
    end

    sky130_fd_sc_hs__sdfxbp dut (.D(D), .SCD(SCD), .SCE(SCE), .VPWR(VPWR), .VGND(VGND), .Q(Q), .Q_N(Q_N), .CLK(CLK));

endmodule

`default_nettype wire
`endif  // SKY130_FD_SC_HS__SDFXBP_TB_V
