# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_hs__clkbuf_8
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__clkbuf_8 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.280000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.462000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.350000 1.095000 1.780000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  1.841700 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.615000 0.350000 1.945000 0.850000 ;
        RECT 1.615000 0.850000 4.880000 1.020000 ;
        RECT 1.615000 1.690000 5.155000 1.860000 ;
        RECT 1.615000 1.860000 1.880000 2.980000 ;
        RECT 2.585000 1.860000 2.845000 2.980000 ;
        RECT 2.615000 0.350000 2.865000 0.850000 ;
        RECT 3.415000 1.860000 3.680000 2.980000 ;
        RECT 3.555000 0.350000 3.725000 0.850000 ;
        RECT 4.385000 1.860000 4.645000 2.980000 ;
        RECT 4.485000 0.350000 4.655000 0.850000 ;
        RECT 4.710000 1.020000 4.880000 1.180000 ;
        RECT 4.710000 1.180000 5.155000 1.690000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 5.280000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 5.280000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.280000 0.085000 ;
      RECT 0.000000  3.245000 5.280000 3.415000 ;
      RECT 0.115000  0.085000 0.445000 0.810000 ;
      RECT 0.115000  1.950000 0.445000 3.245000 ;
      RECT 0.615000  0.350000 0.945000 0.980000 ;
      RECT 0.615000  0.980000 1.445000 1.150000 ;
      RECT 0.615000  1.950000 1.445000 2.120000 ;
      RECT 0.615000  2.120000 0.945000 2.980000 ;
      RECT 1.115000  0.085000 1.445000 0.810000 ;
      RECT 1.115000  2.290000 1.445000 3.245000 ;
      RECT 1.275000  1.150000 1.445000 1.190000 ;
      RECT 1.275000  1.190000 4.515000 1.520000 ;
      RECT 1.275000  1.520000 1.445000 1.950000 ;
      RECT 2.065000  2.030000 2.395000 3.245000 ;
      RECT 2.115000  0.085000 2.445000 0.680000 ;
      RECT 3.045000  0.085000 3.375000 0.680000 ;
      RECT 3.045000  2.030000 3.215000 3.245000 ;
      RECT 3.865000  2.030000 4.195000 3.245000 ;
      RECT 3.905000  0.085000 4.305000 0.680000 ;
      RECT 4.830000  2.030000 5.160000 3.245000 ;
      RECT 4.835000  0.085000 5.165000 0.680000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
  END
END sky130_fd_sc_hs__clkbuf_8
END LIBRARY
