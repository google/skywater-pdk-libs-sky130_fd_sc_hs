* File: sky130_fd_sc_hs__dfrtp_2.spice
* Created: Tue Sep  1 20:00:03 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hs__dfrtp_2.pex.spice"
.subckt sky130_fd_sc_hs__dfrtp_2  VNB VPB D RESET_B CLK VPWR Q VGND
* 
* VGND	VGND
* Q	Q
* VPWR	VPWR
* CLK	CLK
* RESET_B	RESET_B
* D	D
* VPB	VPB
* VNB	VNB
MM1030 A_117_78# N_D_M1030_g N_A_30_78#_M1030_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.0504 AS=0.1197 PD=0.66 PS=1.41 NRD=18.564 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1018 N_VGND_M1018_d N_RESET_B_M1018_g A_117_78# VNB NLOWVT L=0.15 W=0.42
+ AD=0.1197 AS=0.0504 PD=1.41 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75000.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1000 N_VGND_M1000_d N_CLK_M1000_g N_A_306_74#_M1000_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1554 AS=0.2109 PD=1.16 PS=2.05 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75000.8 A=0.111 P=1.78 MULT=1
MM1019 N_A_490_362#_M1019_d N_A_306_74#_M1019_g N_VGND_M1000_d VNB NLOWVT L=0.15
+ W=0.74 AD=0.2109 AS=0.1554 PD=2.05 PS=1.16 NRD=0 NRS=11.34 M=1 R=4.93333
+ SA=75000.8 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1029 N_A_696_457#_M1029_d N_A_306_74#_M1029_g N_A_30_78#_M1029_s VNB NLOWVT
+ L=0.15 W=0.42 AD=0.0735 AS=0.1197 PD=0.77 PS=1.41 NRD=19.992 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75003.7 A=0.063 P=1.14 MULT=1
MM1028 A_817_138# N_A_490_362#_M1028_g N_A_696_457#_M1029_d VNB NLOWVT L=0.15
+ W=0.42 AD=0.0504 AS=0.0735 PD=0.66 PS=0.77 NRD=18.564 NRS=0 M=1 R=2.8
+ SA=75000.7 SB=75003.2 A=0.063 P=1.14 MULT=1
MM1015 A_895_138# N_A_837_359#_M1015_g A_817_138# VNB NLOWVT L=0.15 W=0.42
+ AD=0.0504 AS=0.0504 PD=0.66 PS=0.66 NRD=18.564 NRS=18.564 M=1 R=2.8 SA=75001.1
+ SB=75002.8 A=0.063 P=1.14 MULT=1
MM1001 N_VGND_M1001_d N_RESET_B_M1001_g A_895_138# VNB NLOWVT L=0.15 W=0.42
+ AD=0.255829 AS=0.0504 PD=1.33241 PS=0.66 NRD=158.316 NRS=18.564 M=1 R=2.8
+ SA=75001.5 SB=75002.4 A=0.063 P=1.14 MULT=1
MM1025 N_A_837_359#_M1025_d N_A_696_457#_M1025_g N_VGND_M1001_d VNB NLOWVT
+ L=0.15 W=0.74 AD=0.12025 AS=0.450746 PD=1.065 PS=2.34759 NRD=0 NRS=89.856 M=1
+ R=4.93333 SA=75001.7 SB=75002 A=0.111 P=1.78 MULT=1
MM1003 N_A_1271_74#_M1003_d N_A_490_362#_M1003_g N_A_837_359#_M1025_d VNB NLOWVT
+ L=0.15 W=0.74 AD=0.292172 AS=0.12025 PD=2.09241 PS=1.065 NRD=4.044 NRS=7.296
+ M=1 R=4.93333 SA=75002.2 SB=75001.5 A=0.111 P=1.78 MULT=1
MM1032 A_1481_81# N_A_306_74#_M1032_g N_A_1271_74#_M1003_d VNB NLOWVT L=0.15
+ W=0.42 AD=0.0504 AS=0.165828 PD=0.66 PS=1.18759 NRD=18.564 NRS=47.136 M=1
+ R=2.8 SA=75002.8 SB=75001.5 A=0.063 P=1.14 MULT=1
MM1010 N_VGND_M1010_d N_A_1525_212#_M1010_g A_1481_81# VNB NLOWVT L=0.15 W=0.42
+ AD=0.0777 AS=0.0504 PD=0.79 PS=0.66 NRD=12.852 NRS=18.564 M=1 R=2.8 SA=75003.2
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1023 A_1663_81# N_RESET_B_M1023_g N_VGND_M1010_d VNB NLOWVT L=0.15 W=0.42
+ AD=0.0504 AS=0.0777 PD=0.66 PS=0.79 NRD=18.564 NRS=12.852 M=1 R=2.8 SA=75003.7
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1024 N_A_1525_212#_M1024_d N_A_1271_74#_M1024_g A_1663_81# VNB NLOWVT L=0.15
+ W=0.42 AD=0.1176 AS=0.0504 PD=1.4 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8
+ SA=75004.1 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1022 N_A_1921_409#_M1022_d N_A_1271_74#_M1022_g N_VGND_M1022_s VNB NLOWVT
+ L=0.15 W=0.74 AD=0.2109 AS=0.2072 PD=2.05 PS=2.04 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1031 N_Q_M1031_d N_A_1921_409#_M1031_g N_VGND_M1031_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.2109 PD=1.02 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1033 N_Q_M1031_d N_A_1921_409#_M1033_g N_VGND_M1033_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.2072 PD=1.02 PS=2.04 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.6
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1016 N_A_30_78#_M1016_d N_D_M1016_g N_VPWR_M1016_s VPB PSHORT L=0.15 W=0.42
+ AD=0.063 AS=0.1197 PD=0.72 PS=1.41 NRD=4.6886 NRS=4.6886 M=1 R=2.8 SA=75000.2
+ SB=75000.7 A=0.063 P=1.14 MULT=1
MM1017 N_VPWR_M1017_d N_RESET_B_M1017_g N_A_30_78#_M1016_d VPB PSHORT L=0.15
+ W=0.42 AD=0.1176 AS=0.063 PD=1.4 PS=0.72 NRD=4.6886 NRS=4.6886 M=1 R=2.8
+ SA=75000.7 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1007 N_VPWR_M1007_d N_CLK_M1007_g N_A_306_74#_M1007_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.3136 PD=1.42 PS=2.8 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1012 N_A_490_362#_M1012_d N_A_306_74#_M1012_g N_VPWR_M1007_d VPB PSHORT L=0.15
+ W=1.12 AD=0.3136 AS=0.168 PD=2.8 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.7 SB=75000.2 A=0.168 P=2.54 MULT=1
MM1005 N_A_696_457#_M1005_d N_A_490_362#_M1005_g N_A_30_78#_M1005_s VPB PSHORT
+ L=0.15 W=0.42 AD=0.063 AS=0.1218 PD=0.72 PS=1.42 NRD=4.6886 NRS=4.6886 M=1
+ R=2.8 SA=75000.2 SB=75001.7 A=0.063 P=1.14 MULT=1
MM1008 A_786_457# N_A_306_74#_M1008_g N_A_696_457#_M1005_d VPB PSHORT L=0.15
+ W=0.42 AD=0.0567 AS=0.063 PD=0.69 PS=0.72 NRD=37.5088 NRS=4.6886 M=1 R=2.8
+ SA=75000.7 SB=75001.3 A=0.063 P=1.14 MULT=1
MM1027 N_VPWR_M1027_d N_A_837_359#_M1027_g A_786_457# VPB PSHORT L=0.15 W=0.42
+ AD=0.1393 AS=0.0567 PD=1.17 PS=0.69 NRD=129.764 NRS=37.5088 M=1 R=2.8
+ SA=75001.1 SB=75000.8 A=0.063 P=1.14 MULT=1
MM1020 N_A_696_457#_M1020_d N_RESET_B_M1020_g N_VPWR_M1027_d VPB PSHORT L=0.15
+ W=0.42 AD=0.1239 AS=0.1393 PD=1.43 PS=1.17 NRD=4.6886 NRS=129.764 M=1 R=2.8
+ SA=75001.7 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1013 N_A_837_359#_M1013_d N_A_696_457#_M1013_g N_VPWR_M1013_s VPB PSHORT
+ L=0.15 W=1 AD=0.184062 AS=0.295 PD=1.43 PS=2.59 NRD=11.8003 NRS=1.9503 M=1
+ R=6.66667 SA=75000.2 SB=75001.5 A=0.15 P=2.3 MULT=1
MM1021 N_A_1271_74#_M1021_d N_A_306_74#_M1021_g N_A_837_359#_M1013_d VPB PSHORT
+ L=0.15 W=1 AD=0.319665 AS=0.184062 PD=2.57746 PS=1.43 NRD=10.8153 NRS=2.9353
+ M=1 R=6.66667 SA=75000.7 SB=75001.3 A=0.15 P=2.3 MULT=1
MM1026 A_1478_493# N_A_490_362#_M1026_g N_A_1271_74#_M1021_d VPB PSHORT L=0.15
+ W=0.42 AD=0.0567 AS=0.13426 PD=0.69 PS=1.08254 NRD=37.5088 NRS=4.6886 M=1
+ R=2.8 SA=75001.3 SB=75002.4 A=0.063 P=1.14 MULT=1
MM1011 N_VPWR_M1011_d N_A_1525_212#_M1011_g A_1478_493# VPB PSHORT L=0.15 W=0.42
+ AD=0.0735 AS=0.0567 PD=0.77 PS=0.69 NRD=4.6886 NRS=37.5088 M=1 R=2.8
+ SA=75001.7 SB=75002 A=0.063 P=1.14 MULT=1
MM1009 N_A_1525_212#_M1009_d N_RESET_B_M1009_g N_VPWR_M1011_d VPB PSHORT L=0.15
+ W=0.42 AD=0.1176 AS=0.0735 PD=0.98 PS=0.77 NRD=65.6601 NRS=28.1316 M=1 R=2.8
+ SA=75002.2 SB=75001.5 A=0.063 P=1.14 MULT=1
MM1014 N_VPWR_M1014_d N_A_1271_74#_M1014_g N_A_1525_212#_M1009_d VPB PSHORT
+ L=0.15 W=0.42 AD=0.1092 AS=0.1176 PD=0.85 PS=0.98 NRD=44.5417 NRS=65.6601 M=1
+ R=2.8 SA=75002.9 SB=75000.8 A=0.063 P=1.14 MULT=1
MM1002 N_A_1921_409#_M1002_d N_A_1271_74#_M1002_g N_VPWR_M1014_d VPB PSHORT
+ L=0.15 W=0.84 AD=0.2478 AS=0.2184 PD=2.27 PS=1.7 NRD=2.3443 NRS=14.0658 M=1
+ R=5.6 SA=75001.9 SB=75000.2 A=0.126 P=1.98 MULT=1
MM1004 N_Q_M1004_d N_A_1921_409#_M1004_g N_VPWR_M1004_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.3584 PD=1.42 PS=2.88 NRD=1.7533 NRS=6.1464 M=1 R=7.46667
+ SA=75000.2 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1006 N_Q_M1004_d N_A_1921_409#_M1006_g N_VPWR_M1006_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.3304 PD=1.42 PS=2.83 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.7 SB=75000.2 A=0.168 P=2.54 MULT=1
DX34_noxref VNB VPB NWDIODE A=22.7157 P=27.73
c_115 VNB 0 8.65509e-20 $X=0 $Y=0
c_242 VPB 0 1.21261e-19 $X=0 $Y=3.085
c_1690 A_1478_493# 0 1.15577e-19 $X=7.39 $Y=2.465
*
.include "sky130_fd_sc_hs__dfrtp_2.pxi.spice"
*
.ends
*
*
