* File: sky130_fd_sc_hs__nand2b_2.pex.spice
* Created: Thu Aug 27 20:50:36 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HS__NAND2B_2%A_N 3 5 7 8 12
c28 12 0 1.50161e-19 $X=0.405 $Y=1.515
c29 5 0 1.52201e-19 $X=0.505 $Y=1.765
r30 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.405
+ $Y=1.515 $X2=0.405 $Y2=1.515
r31 8 12 4.42216 $w=4.28e-07 $l=1.65e-07 $layer=LI1_cond $X=0.24 $Y=1.565
+ $X2=0.405 $Y2=1.565
r32 5 11 52.4661 $w=2.95e-07 $l=2.93684e-07 $layer=POLY_cond $X=0.505 $Y=1.765
+ $X2=0.41 $Y2=1.515
r33 5 7 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=0.505 $Y=1.765
+ $X2=0.505 $Y2=2.34
r34 1 11 38.578 $w=2.95e-07 $l=2.03101e-07 $layer=POLY_cond $X=0.495 $Y=1.35
+ $X2=0.41 $Y2=1.515
r35 1 3 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.495 $Y=1.35
+ $X2=0.495 $Y2=0.69
.ends

.subckt PM_SKY130_FD_SC_HS__NAND2B_2%A_27_74# 1 2 7 10 11 13 16 18 21 22 24 27
+ 29 30 33 37 38 39 41 42 44 48
c99 48 0 1.50161e-19 $X=0.97 $Y=1.305
c100 41 0 3.18194e-19 $X=0.89 $Y=1.47
c101 30 0 2.21113e-19 $X=1.97 $Y=1.395
r102 48 51 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=0.97 $Y=1.305
+ $X2=0.97 $Y2=1.395
r103 47 48 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.97
+ $Y=1.305 $X2=0.97 $Y2=1.305
r104 45 47 9.02113 $w=2.84e-07 $l=2.1e-07 $layer=LI1_cond $X=0.97 $Y=1.095
+ $X2=0.97 $Y2=1.305
r105 41 47 9.03839 $w=2.84e-07 $l=2.0106e-07 $layer=LI1_cond $X=0.89 $Y=1.47
+ $X2=0.97 $Y2=1.305
r106 41 42 31.3155 $w=1.68e-07 $l=4.8e-07 $layer=LI1_cond $X=0.89 $Y=1.47
+ $X2=0.89 $Y2=1.95
r107 40 44 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.445 $Y=2.035
+ $X2=0.28 $Y2=2.035
r108 39 42 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.805 $Y=2.035
+ $X2=0.89 $Y2=1.95
r109 39 40 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=0.805 $Y=2.035
+ $X2=0.445 $Y2=2.035
r110 37 45 3.73949 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.805 $Y=1.095
+ $X2=0.97 $Y2=1.095
r111 37 38 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=0.805 $Y=1.095
+ $X2=0.445 $Y2=1.095
r112 31 38 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.28 $Y=1.01
+ $X2=0.445 $Y2=1.095
r113 31 33 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=0.28 $Y=1.01
+ $X2=0.28 $Y2=0.515
r114 25 30 18.8402 $w=1.65e-07 $l=8.87412e-08 $layer=POLY_cond $X=2 $Y=1.32
+ $X2=1.97 $Y2=1.395
r115 25 27 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=2 $Y=1.32 $X2=2
+ $Y2=0.74
r116 22 24 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.955 $Y=1.765
+ $X2=1.955 $Y2=2.4
r117 21 22 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=1.955 $Y=1.675
+ $X2=1.955 $Y2=1.765
r118 20 30 18.8402 $w=1.65e-07 $l=8.21584e-08 $layer=POLY_cond $X=1.955 $Y=1.47
+ $X2=1.97 $Y2=1.395
r119 20 21 79.6855 $w=1.8e-07 $l=2.05e-07 $layer=POLY_cond $X=1.955 $Y=1.47
+ $X2=1.955 $Y2=1.675
r120 19 29 13.2179 $w=1.5e-07 $l=1.15e-07 $layer=POLY_cond $X=1.645 $Y=1.395
+ $X2=1.53 $Y2=1.395
r121 18 30 6.66866 $w=1.5e-07 $l=1.05e-07 $layer=POLY_cond $X=1.865 $Y=1.395
+ $X2=1.97 $Y2=1.395
r122 18 19 112.809 $w=1.5e-07 $l=2.2e-07 $layer=POLY_cond $X=1.865 $Y=1.395
+ $X2=1.645 $Y2=1.395
r123 14 29 10.9219 $w=1.5e-07 $l=9.28709e-08 $layer=POLY_cond $X=1.57 $Y=1.32
+ $X2=1.53 $Y2=1.395
r124 14 16 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=1.57 $Y=1.32
+ $X2=1.57 $Y2=0.74
r125 11 13 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.505 $Y=1.765
+ $X2=1.505 $Y2=2.4
r126 10 11 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=1.505 $Y=1.675
+ $X2=1.505 $Y2=1.765
r127 9 29 10.9219 $w=1.8e-07 $l=8.66025e-08 $layer=POLY_cond $X=1.505 $Y=1.47
+ $X2=1.53 $Y2=1.395
r128 9 10 79.6855 $w=1.8e-07 $l=2.05e-07 $layer=POLY_cond $X=1.505 $Y=1.47
+ $X2=1.505 $Y2=1.675
r129 8 51 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.135 $Y=1.395
+ $X2=0.97 $Y2=1.395
r130 7 29 13.2179 $w=1.5e-07 $l=1.15e-07 $layer=POLY_cond $X=1.415 $Y=1.395
+ $X2=1.53 $Y2=1.395
r131 7 8 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=1.415 $Y=1.395
+ $X2=1.135 $Y2=1.395
r132 2 44 300 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.115
r133 1 33 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__NAND2B_2%B 1 3 6 8 10 13 15 21 22
c50 21 0 8.98252e-20 $X=2.61 $Y=1.515
r51 22 23 1.27513 $w=3.78e-07 $l=1e-08 $layer=POLY_cond $X=2.855 $Y=1.557
+ $X2=2.865 $Y2=1.557
r52 20 22 31.2407 $w=3.78e-07 $l=2.45e-07 $layer=POLY_cond $X=2.61 $Y=1.557
+ $X2=2.855 $Y2=1.557
r53 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.61
+ $Y=1.515 $X2=2.61 $Y2=1.515
r54 18 20 22.9524 $w=3.78e-07 $l=1.8e-07 $layer=POLY_cond $X=2.43 $Y=1.557
+ $X2=2.61 $Y2=1.557
r55 17 18 3.18783 $w=3.78e-07 $l=2.5e-08 $layer=POLY_cond $X=2.405 $Y=1.557
+ $X2=2.43 $Y2=1.557
r56 15 21 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=2.61 $Y=1.665
+ $X2=2.61 $Y2=1.515
r57 11 23 24.4846 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.865 $Y=1.35
+ $X2=2.865 $Y2=1.557
r58 11 13 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.865 $Y=1.35
+ $X2=2.865 $Y2=0.74
r59 8 22 24.4846 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=2.855 $Y=1.765
+ $X2=2.855 $Y2=1.557
r60 8 10 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.855 $Y=1.765
+ $X2=2.855 $Y2=2.4
r61 4 18 24.4846 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.43 $Y=1.35
+ $X2=2.43 $Y2=1.557
r62 4 6 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.43 $Y=1.35 $X2=2.43
+ $Y2=0.74
r63 1 17 24.4846 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=2.405 $Y=1.765
+ $X2=2.405 $Y2=1.557
r64 1 3 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.405 $Y=1.765
+ $X2=2.405 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_HS__NAND2B_2%VPWR 1 2 3 12 16 18 20 23 24 25 31 35 41 45
r47 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r48 41 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r49 39 45 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r50 39 42 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=2.16 $Y2=3.33
r51 38 39 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r52 36 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.345 $Y=3.33
+ $X2=2.18 $Y2=3.33
r53 36 38 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=2.345 $Y=3.33
+ $X2=2.64 $Y2=3.33
r54 35 44 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=2.915 $Y=3.33
+ $X2=3.137 $Y2=3.33
r55 35 38 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=2.915 $Y=3.33
+ $X2=2.64 $Y2=3.33
r56 31 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.015 $Y=3.33
+ $X2=2.18 $Y2=3.33
r57 31 33 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=2.015 $Y=3.33
+ $X2=1.68 $Y2=3.33
r58 28 29 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r59 25 42 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r60 25 29 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=0.72 $Y2=3.33
r61 25 33 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r62 23 28 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=0.725 $Y=3.33
+ $X2=0.72 $Y2=3.33
r63 23 24 9.31531 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=0.725 $Y=3.33
+ $X2=0.91 $Y2=3.33
r64 22 33 38.1658 $w=1.68e-07 $l=5.85e-07 $layer=LI1_cond $X=1.095 $Y=3.33
+ $X2=1.68 $Y2=3.33
r65 22 24 9.31531 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=1.095 $Y=3.33
+ $X2=0.91 $Y2=3.33
r66 18 44 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=3.08 $Y=3.245
+ $X2=3.137 $Y2=3.33
r67 18 20 15.3659 $w=3.28e-07 $l=4.4e-07 $layer=LI1_cond $X=3.08 $Y=3.245
+ $X2=3.08 $Y2=2.805
r68 14 41 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.18 $Y=3.245
+ $X2=2.18 $Y2=3.33
r69 14 16 15.3659 $w=3.28e-07 $l=4.4e-07 $layer=LI1_cond $X=2.18 $Y=3.245
+ $X2=2.18 $Y2=2.805
r70 10 24 1.24149 $w=3.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.91 $Y=3.245
+ $X2=0.91 $Y2=3.33
r71 10 12 26.1636 $w=3.68e-07 $l=8.4e-07 $layer=LI1_cond $X=0.91 $Y=3.245
+ $X2=0.91 $Y2=2.405
r72 3 20 600 $w=1.7e-07 $l=1.03729e-06 $layer=licon1_PDIFF $count=1 $X=2.93
+ $Y=1.84 $X2=3.08 $Y2=2.805
r73 2 16 600 $w=1.7e-07 $l=1.03729e-06 $layer=licon1_PDIFF $count=1 $X=2.03
+ $Y=1.84 $X2=2.18 $Y2=2.805
r74 1 12 300 $w=1.7e-07 $l=7.13092e-07 $layer=licon1_PDIFF $count=2 $X=0.58
+ $Y=1.84 $X2=0.915 $Y2=2.405
.ends

.subckt PM_SKY130_FD_SC_HS__NAND2B_2%Y 1 2 3 10 16 18 19 22 25 26
c43 26 0 1.91961e-19 $X=2.16 $Y=2.035
c44 19 0 1.31288e-19 $X=1.87 $Y=1.305
r45 26 29 2.49594 $w=2.3e-07 $l=1.9e-07 $layer=LI1_cond $X=2.16 $Y=2.01 $X2=2.16
+ $Y2=1.82
r46 25 29 7.76646 $w=2.28e-07 $l=1.55e-07 $layer=LI1_cond $X=2.16 $Y=1.665
+ $X2=2.16 $Y2=1.82
r47 24 25 13.7792 $w=2.28e-07 $l=2.75e-07 $layer=LI1_cond $X=2.16 $Y=1.39
+ $X2=2.16 $Y2=1.665
r48 20 26 3.9473 $w=3.15e-07 $l=1.43875e-07 $layer=LI1_cond $X=2.275 $Y=2.075
+ $X2=2.16 $Y2=2.01
r49 20 22 16.3647 $w=2.48e-07 $l=3.55e-07 $layer=LI1_cond $X=2.275 $Y=2.075
+ $X2=2.63 $Y2=2.075
r50 18 24 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=2.045 $Y=1.305
+ $X2=2.16 $Y2=1.39
r51 18 19 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=2.045 $Y=1.305
+ $X2=1.87 $Y2=1.305
r52 14 19 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.785 $Y=1.22
+ $X2=1.87 $Y2=1.305
r53 14 16 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=1.785 $Y=1.22
+ $X2=1.785 $Y2=0.825
r54 10 26 3.9473 $w=3.15e-07 $l=1.15e-07 $layer=LI1_cond $X=2.045 $Y=2.01
+ $X2=2.16 $Y2=2.01
r55 10 12 9.55315 $w=3.78e-07 $l=3.15e-07 $layer=LI1_cond $X=2.045 $Y=2.01
+ $X2=1.73 $Y2=2.01
r56 3 22 600 $w=1.7e-07 $l=3.4187e-07 $layer=licon1_PDIFF $count=1 $X=2.48
+ $Y=1.84 $X2=2.63 $Y2=2.115
r57 2 12 600 $w=1.7e-07 $l=2.33238e-07 $layer=licon1_PDIFF $count=1 $X=1.58
+ $Y=1.84 $X2=1.73 $Y2=2.01
r58 1 16 182 $w=1.7e-07 $l=5.20312e-07 $layer=licon1_NDIFF $count=1 $X=1.645
+ $Y=0.37 $X2=1.785 $Y2=0.825
.ends

.subckt PM_SKY130_FD_SC_HS__NAND2B_2%VGND 1 2 9 13 15 17 22 29 30 33 36
c40 1 0 1.65994e-19 $X=0.57 $Y=0.37
r41 36 37 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r42 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r43 30 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=2.64
+ $Y2=0
r44 29 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r45 27 36 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.73 $Y=0 $X2=2.645
+ $Y2=0
r46 27 29 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=2.73 $Y=0 $X2=3.12
+ $Y2=0
r47 26 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r48 25 26 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r49 23 33 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=0.875 $Y=0 $X2=0.745
+ $Y2=0
r50 23 25 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.875 $Y=0 $X2=1.2
+ $Y2=0
r51 22 36 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.56 $Y=0 $X2=2.645
+ $Y2=0
r52 22 25 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=2.56 $Y=0 $X2=1.2
+ $Y2=0
r53 20 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r54 19 20 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r55 17 33 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=0.615 $Y=0 $X2=0.745
+ $Y2=0
r56 17 19 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=0.615 $Y=0 $X2=0.24
+ $Y2=0
r57 15 37 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.64
+ $Y2=0
r58 15 26 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r59 11 36 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.645 $Y=0.085
+ $X2=2.645 $Y2=0
r60 11 13 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=2.645 $Y=0.085
+ $X2=2.645 $Y2=0.515
r61 7 33 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=0.745 $Y=0.085
+ $X2=0.745 $Y2=0
r62 7 9 26.1516 $w=2.58e-07 $l=5.9e-07 $layer=LI1_cond $X=0.745 $Y=0.085
+ $X2=0.745 $Y2=0.675
r63 2 13 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.505
+ $Y=0.37 $X2=2.645 $Y2=0.515
r64 1 9 182 $w=1.7e-07 $l=3.68409e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.37 $X2=0.71 $Y2=0.675
.ends

.subckt PM_SKY130_FD_SC_HS__NAND2B_2%A_242_74# 1 2 3 13 15 16 17 18 19 22 26 29
+ 30 31
r80 29 31 80.8984 $w=1.68e-07 $l=1.24e-06 $layer=LI1_cond $X=3.16 $Y=2.37
+ $X2=3.16 $Y2=1.13
r81 24 31 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=3.08 $Y=0.965
+ $X2=3.08 $Y2=1.13
r82 24 26 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=3.08 $Y=0.965
+ $X2=3.08 $Y2=0.515
r83 20 22 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=2.215 $Y=0.425
+ $X2=2.215 $Y2=0.515
r84 18 20 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.05 $Y=0.34
+ $X2=2.215 $Y2=0.425
r85 18 19 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=2.05 $Y=0.34
+ $X2=1.52 $Y2=0.34
r86 16 29 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.075 $Y=2.455
+ $X2=3.16 $Y2=2.37
r87 16 17 104.385 $w=1.68e-07 $l=1.6e-06 $layer=LI1_cond $X=3.075 $Y=2.455
+ $X2=1.475 $Y2=2.455
r88 15 17 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.39 $Y=2.37
+ $X2=1.475 $Y2=2.455
r89 15 30 91.3369 $w=1.68e-07 $l=1.4e-06 $layer=LI1_cond $X=1.39 $Y=2.37
+ $X2=1.39 $Y2=0.97
r90 11 30 7.49019 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=1.355 $Y=0.805
+ $X2=1.355 $Y2=0.97
r91 11 13 10.1275 $w=3.28e-07 $l=2.9e-07 $layer=LI1_cond $X=1.355 $Y=0.805
+ $X2=1.355 $Y2=0.515
r92 10 19 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.355 $Y=0.425
+ $X2=1.52 $Y2=0.34
r93 10 13 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=1.355 $Y=0.425
+ $X2=1.355 $Y2=0.515
r94 3 26 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.94
+ $Y=0.37 $X2=3.08 $Y2=0.515
r95 2 22 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.075
+ $Y=0.37 $X2=2.215 $Y2=0.515
r96 1 13 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=1.21
+ $Y=0.37 $X2=1.355 $Y2=0.515
.ends

