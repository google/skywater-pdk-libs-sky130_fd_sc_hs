* File: sky130_fd_sc_hs__ebufn_8.spice
* Created: Tue Sep  1 20:04:15 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hs__ebufn_8.pex.spice"
.subckt sky130_fd_sc_hs__ebufn_8  VNB VPB TE_B A Z VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* Z	Z
* A	A
* TE_B	TE_B
* VPB	VPB
* VNB	VNB
MM1005 N_A_27_74#_M1005_d N_A_84_48#_M1005_g N_Z_M1005_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.2109 AS=0.1036 PD=2.05 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75007 A=0.111 P=1.78 MULT=1
MM1009 N_A_27_74#_M1009_d N_A_84_48#_M1009_g N_Z_M1005_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.11285 AS=0.1036 PD=1.045 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.6 SB=75006.5 A=0.111 P=1.78 MULT=1
MM1011 N_A_27_74#_M1009_d N_A_84_48#_M1011_g N_Z_M1011_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.11285 AS=0.1036 PD=1.045 PS=1.02 NRD=4.044 NRS=0 M=1 R=4.93333
+ SA=75001.1 SB=75006.1 A=0.111 P=1.78 MULT=1
MM1029 N_A_27_74#_M1029_d N_A_84_48#_M1029_g N_Z_M1011_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1295 AS=0.1036 PD=1.09 PS=1.02 NRD=11.34 NRS=0 M=1 R=4.93333
+ SA=75001.5 SB=75005.6 A=0.111 P=1.78 MULT=1
MM1032 N_A_27_74#_M1029_d N_A_84_48#_M1032_g N_Z_M1032_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1295 AS=0.1295 PD=1.09 PS=1.09 NRD=0 NRS=11.34 M=1 R=4.93333
+ SA=75002 SB=75005.1 A=0.111 P=1.78 MULT=1
MM1033 N_A_27_74#_M1033_d N_A_84_48#_M1033_g N_Z_M1032_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.13505 AS=0.1295 PD=1.105 PS=1.09 NRD=11.34 NRS=0 M=1 R=4.93333
+ SA=75002.5 SB=75004.6 A=0.111 P=1.78 MULT=1
MM1034 N_A_27_74#_M1033_d N_A_84_48#_M1034_g N_Z_M1034_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.13505 AS=0.12395 PD=1.105 PS=1.075 NRD=2.424 NRS=8.916 M=1
+ R=4.93333 SA=75003 SB=75004.1 A=0.111 P=1.78 MULT=1
MM1036 N_A_27_74#_M1036_d N_A_84_48#_M1036_g N_Z_M1034_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.12395 PD=1.02 PS=1.075 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75003.5 SB=75003.6 A=0.111 P=1.78 MULT=1
MM1001 N_A_27_74#_M1036_d N_A_833_48#_M1001_g N_VGND_M1001_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75004
+ SB=75003.2 A=0.111 P=1.78 MULT=1
MM1003 N_A_27_74#_M1003_d N_A_833_48#_M1003_g N_VGND_M1001_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75004.4 SB=75002.8 A=0.111 P=1.78 MULT=1
MM1004 N_A_27_74#_M1003_d N_A_833_48#_M1004_g N_VGND_M1004_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75004.8 SB=75002.4 A=0.111 P=1.78 MULT=1
MM1012 N_A_27_74#_M1012_d N_A_833_48#_M1012_g N_VGND_M1004_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75005.2 SB=75001.9 A=0.111 P=1.78 MULT=1
MM1025 N_A_27_74#_M1012_d N_A_833_48#_M1025_g N_VGND_M1025_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75005.7 SB=75001.5 A=0.111 P=1.78 MULT=1
MM1027 N_A_27_74#_M1027_d N_A_833_48#_M1027_g N_VGND_M1025_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75006.1 SB=75001.1 A=0.111 P=1.78 MULT=1
MM1035 N_A_27_74#_M1027_d N_A_833_48#_M1035_g N_VGND_M1035_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75006.5 SB=75000.6 A=0.111 P=1.78 MULT=1
MM1037 N_A_27_74#_M1037_d N_A_833_48#_M1037_g N_VGND_M1035_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.2109 AS=0.1036 PD=2.05 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75007
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1031 N_VGND_M1031_d N_TE_B_M1031_g N_A_833_48#_M1031_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.2109 PD=1.02 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75001.1 A=0.111 P=1.78 MULT=1
MM1008 N_A_84_48#_M1008_d N_A_M1008_g N_VGND_M1031_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.6
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1018 N_A_84_48#_M1008_d N_A_M1018_g N_VGND_M1018_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.2146 PD=1.02 PS=2.06 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.1
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1006 N_A_28_368#_M1006_d N_A_84_48#_M1006_g N_Z_M1006_s VPB PSHORT L=0.15
+ W=1.12 AD=0.3304 AS=0.168 PD=2.83 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75007.6 A=0.168 P=2.54 MULT=1
MM1010 N_A_28_368#_M1010_d N_A_84_48#_M1010_g N_Z_M1006_s VPB PSHORT L=0.15
+ W=1.12 AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.7 SB=75007.1 A=0.168 P=2.54 MULT=1
MM1013 N_A_28_368#_M1010_d N_A_84_48#_M1013_g N_Z_M1013_s VPB PSHORT L=0.15
+ W=1.12 AD=0.168 AS=0.196 PD=1.42 PS=1.47 NRD=1.7533 NRS=10.5395 M=1 R=7.46667
+ SA=75001.1 SB=75006.7 A=0.168 P=2.54 MULT=1
MM1014 N_A_28_368#_M1014_d N_A_84_48#_M1014_g N_Z_M1013_s VPB PSHORT L=0.15
+ W=1.12 AD=0.168 AS=0.196 PD=1.42 PS=1.47 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.6 SB=75006.2 A=0.168 P=2.54 MULT=1
MM1015 N_A_28_368#_M1014_d N_A_84_48#_M1015_g N_Z_M1015_s VPB PSHORT L=0.15
+ W=1.12 AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75002.1 SB=75005.7 A=0.168 P=2.54 MULT=1
MM1017 N_A_28_368#_M1017_d N_A_84_48#_M1017_g N_Z_M1015_s VPB PSHORT L=0.15
+ W=1.12 AD=0.196 AS=0.168 PD=1.47 PS=1.42 NRD=10.5395 NRS=1.7533 M=1 R=7.46667
+ SA=75002.5 SB=75005.3 A=0.168 P=2.54 MULT=1
MM1019 N_A_28_368#_M1017_d N_A_84_48#_M1019_g N_Z_M1019_s VPB PSHORT L=0.15
+ W=1.12 AD=0.196 AS=0.1876 PD=1.47 PS=1.455 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75003 SB=75004.8 A=0.168 P=2.54 MULT=1
MM1020 N_A_28_368#_M1020_d N_A_84_48#_M1020_g N_Z_M1019_s VPB PSHORT L=0.15
+ W=1.12 AD=0.1764 AS=0.1876 PD=1.435 PS=1.455 NRD=4.3931 NRS=7.8997 M=1
+ R=7.46667 SA=75003.5 SB=75004.3 A=0.168 P=2.54 MULT=1
MM1016 N_A_28_368#_M1020_d N_TE_B_M1016_g N_VPWR_M1016_s VPB PSHORT L=0.15
+ W=1.12 AD=0.1764 AS=0.224 PD=1.435 PS=1.52 NRD=1.7533 NRS=10.5395 M=1
+ R=7.46667 SA=75004 SB=75003.8 A=0.168 P=2.54 MULT=1
MM1021 N_A_28_368#_M1021_d N_TE_B_M1021_g N_VPWR_M1016_s VPB PSHORT L=0.15
+ W=1.12 AD=0.168 AS=0.224 PD=1.42 PS=1.52 NRD=1.7533 NRS=10.5395 M=1 R=7.46667
+ SA=75004.5 SB=75003.3 A=0.168 P=2.54 MULT=1
MM1022 N_A_28_368#_M1021_d N_TE_B_M1022_g N_VPWR_M1022_s VPB PSHORT L=0.15
+ W=1.12 AD=0.168 AS=0.224 PD=1.42 PS=1.52 NRD=1.7533 NRS=10.5395 M=1 R=7.46667
+ SA=75005 SB=75002.8 A=0.168 P=2.54 MULT=1
MM1023 N_A_28_368#_M1023_d N_TE_B_M1023_g N_VPWR_M1022_s VPB PSHORT L=0.15
+ W=1.12 AD=0.168 AS=0.224 PD=1.42 PS=1.52 NRD=1.7533 NRS=10.5395 M=1 R=7.46667
+ SA=75005.5 SB=75002.3 A=0.168 P=2.54 MULT=1
MM1024 N_A_28_368#_M1023_d N_TE_B_M1024_g N_VPWR_M1024_s VPB PSHORT L=0.15
+ W=1.12 AD=0.168 AS=0.224 PD=1.42 PS=1.52 NRD=1.7533 NRS=10.5395 M=1 R=7.46667
+ SA=75006 SB=75001.8 A=0.168 P=2.54 MULT=1
MM1026 N_A_28_368#_M1026_d N_TE_B_M1026_g N_VPWR_M1024_s VPB PSHORT L=0.15
+ W=1.12 AD=0.168 AS=0.224 PD=1.42 PS=1.52 NRD=1.7533 NRS=10.5395 M=1 R=7.46667
+ SA=75006.5 SB=75001.3 A=0.168 P=2.54 MULT=1
MM1028 N_A_28_368#_M1026_d N_TE_B_M1028_g N_VPWR_M1028_s VPB PSHORT L=0.15
+ W=1.12 AD=0.168 AS=0.28785 PD=1.42 PS=1.76 NRD=0 NRS=35.5191 M=1 R=7.46667
+ SA=75007 SB=75000.8 A=0.168 P=2.54 MULT=1
MM1030 N_A_28_368#_M1030_d N_TE_B_M1030_g N_VPWR_M1028_s VPB PSHORT L=0.15
+ W=1.12 AD=0.3304 AS=0.28785 PD=2.83 PS=1.76 NRD=0 NRS=35.5191 M=1 R=7.46667
+ SA=75007.6 SB=75000.2 A=0.168 P=2.54 MULT=1
MM1002 N_VPWR_M1002_d N_TE_B_M1002_g N_A_833_48#_M1002_s VPB PSHORT L=0.15
+ W=1.12 AD=0.196 AS=0.5712 PD=1.47 PS=3.26 NRD=1.7533 NRS=21.0987 M=1 R=7.46667
+ SA=75000.4 SB=75001.2 A=0.168 P=2.54 MULT=1
MM1000 N_A_84_48#_M1000_d N_A_M1000_g N_VPWR_M1002_d VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.196 PD=1.42 PS=1.47 NRD=1.7533 NRS=10.5395 M=1 R=7.46667
+ SA=75000.9 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1007 N_A_84_48#_M1000_d N_A_M1007_g N_VPWR_M1007_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.3304 PD=1.42 PS=2.83 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.4 SB=75000.2 A=0.168 P=2.54 MULT=1
DX38_noxref VNB VPB NWDIODE A=20.3484 P=25.6
c_117 VNB 0 8.42804e-20 $X=0 $Y=0
*
.include "sky130_fd_sc_hs__ebufn_8.pxi.spice"
*
.ends
*
*
