* File: sky130_fd_sc_hs__nor4bb_4.pxi.spice
* Created: Tue Sep  1 20:12:52 2020
* 
x_PM_SKY130_FD_SC_HS__NOR4BB_4%B N_B_c_185_n N_B_M1010_g N_B_M1001_g N_B_M1020_g
+ N_B_c_195_n N_B_M1012_g N_B_c_196_n N_B_M1015_g N_B_M1028_g N_B_c_197_n
+ N_B_M1027_g N_B_M1034_g N_B_c_190_n N_B_c_199_n N_B_c_191_n N_B_c_192_n B
+ N_B_c_193_n PM_SKY130_FD_SC_HS__NOR4BB_4%B
x_PM_SKY130_FD_SC_HS__NOR4BB_4%A N_A_c_305_n N_A_M1011_g N_A_c_313_n N_A_M1021_g
+ N_A_c_314_n N_A_M1022_g N_A_c_306_n N_A_M1017_g N_A_c_315_n N_A_M1024_g
+ N_A_c_307_n N_A_M1023_g N_A_c_308_n N_A_M1033_g N_A_c_309_n N_A_M1031_g
+ N_A_c_310_n A A N_A_c_311_n N_A_c_312_n PM_SKY130_FD_SC_HS__NOR4BB_4%A
x_PM_SKY130_FD_SC_HS__NOR4BB_4%A_864_48# N_A_864_48#_M1025_d N_A_864_48#_M1000_d
+ N_A_864_48#_M1009_g N_A_864_48#_c_414_n N_A_864_48#_M1007_g
+ N_A_864_48#_c_415_n N_A_864_48#_M1013_g N_A_864_48#_M1014_g
+ N_A_864_48#_M1035_g N_A_864_48#_c_402_n N_A_864_48#_M1032_g
+ N_A_864_48#_c_417_n N_A_864_48#_M1037_g N_A_864_48#_c_403_n
+ N_A_864_48#_M1036_g N_A_864_48#_c_404_n N_A_864_48#_c_405_n
+ N_A_864_48#_c_430_n N_A_864_48#_c_406_n N_A_864_48#_c_420_n
+ N_A_864_48#_c_438_p N_A_864_48#_c_489_p N_A_864_48#_c_516_p
+ N_A_864_48#_c_421_n N_A_864_48#_c_422_n N_A_864_48#_c_407_n
+ N_A_864_48#_c_408_n N_A_864_48#_c_409_n N_A_864_48#_c_410_n
+ N_A_864_48#_c_424_n N_A_864_48#_c_411_n N_A_864_48#_c_425_n
+ N_A_864_48#_c_426_n N_A_864_48#_c_412_n N_A_864_48#_c_413_n
+ PM_SKY130_FD_SC_HS__NOR4BB_4%A_864_48#
x_PM_SKY130_FD_SC_HS__NOR4BB_4%A_1162_48# N_A_1162_48#_M1008_d
+ N_A_1162_48#_M1026_d N_A_1162_48#_M1004_g N_A_1162_48#_c_581_n
+ N_A_1162_48#_c_602_n N_A_1162_48#_M1002_g N_A_1162_48#_c_582_n
+ N_A_1162_48#_c_583_n N_A_1162_48#_c_604_n N_A_1162_48#_M1006_g
+ N_A_1162_48#_M1005_g N_A_1162_48#_c_585_n N_A_1162_48#_c_586_n
+ N_A_1162_48#_M1018_g N_A_1162_48#_c_605_n N_A_1162_48#_M1016_g
+ N_A_1162_48#_c_606_n N_A_1162_48#_M1019_g N_A_1162_48#_c_587_n
+ N_A_1162_48#_M1030_g N_A_1162_48#_c_588_n N_A_1162_48#_c_589_n
+ N_A_1162_48#_c_590_n N_A_1162_48#_c_591_n N_A_1162_48#_c_592_n
+ N_A_1162_48#_c_638_n N_A_1162_48#_c_739_p N_A_1162_48#_c_740_p
+ N_A_1162_48#_c_593_n N_A_1162_48#_c_594_n N_A_1162_48#_c_595_n
+ N_A_1162_48#_c_596_n N_A_1162_48#_c_597_n N_A_1162_48#_c_608_n
+ N_A_1162_48#_c_609_n N_A_1162_48#_c_610_n N_A_1162_48#_c_598_n
+ N_A_1162_48#_c_599_n N_A_1162_48#_c_600_n
+ PM_SKY130_FD_SC_HS__NOR4BB_4%A_1162_48#
x_PM_SKY130_FD_SC_HS__NOR4BB_4%C_N N_C_N_c_775_n N_C_N_M1000_g N_C_N_M1025_g
+ N_C_N_c_776_n N_C_N_M1003_g C_N C_N N_C_N_c_774_n
+ PM_SKY130_FD_SC_HS__NOR4BB_4%C_N
x_PM_SKY130_FD_SC_HS__NOR4BB_4%D_N N_D_N_c_823_n N_D_N_c_824_n N_D_N_M1026_g
+ N_D_N_c_825_n N_D_N_c_826_n N_D_N_M1029_g N_D_N_M1008_g D_N N_D_N_c_822_n
+ PM_SKY130_FD_SC_HS__NOR4BB_4%D_N
x_PM_SKY130_FD_SC_HS__NOR4BB_4%A_27_368# N_A_27_368#_M1010_d N_A_27_368#_M1012_d
+ N_A_27_368#_M1027_d N_A_27_368#_M1013_d N_A_27_368#_M1037_d
+ N_A_27_368#_c_863_n N_A_27_368#_c_870_n N_A_27_368#_c_876_n
+ N_A_27_368#_c_878_n N_A_27_368#_c_942_p N_A_27_368#_c_864_n
+ N_A_27_368#_c_865_n N_A_27_368#_c_866_n N_A_27_368#_c_867_n
+ N_A_27_368#_c_868_n N_A_27_368#_c_886_n PM_SKY130_FD_SC_HS__NOR4BB_4%A_27_368#
x_PM_SKY130_FD_SC_HS__NOR4BB_4%A_116_368# N_A_116_368#_M1010_s
+ N_A_116_368#_M1022_s N_A_116_368#_M1033_s N_A_116_368#_M1015_s
+ N_A_116_368#_c_965_n N_A_116_368#_c_949_n N_A_116_368#_c_970_n
+ N_A_116_368#_c_983_n N_A_116_368#_c_950_n N_A_116_368#_c_951_n
+ N_A_116_368#_c_952_n N_A_116_368#_c_953_n N_A_116_368#_c_954_n
+ N_A_116_368#_c_976_n PM_SKY130_FD_SC_HS__NOR4BB_4%A_116_368#
x_PM_SKY130_FD_SC_HS__NOR4BB_4%VPWR N_VPWR_M1021_d N_VPWR_M1024_d N_VPWR_M1000_s
+ N_VPWR_M1003_s N_VPWR_M1029_s N_VPWR_c_1011_n N_VPWR_c_1012_n N_VPWR_c_1013_n
+ N_VPWR_c_1014_n N_VPWR_c_1015_n N_VPWR_c_1016_n N_VPWR_c_1017_n VPWR
+ N_VPWR_c_1018_n N_VPWR_c_1019_n N_VPWR_c_1020_n N_VPWR_c_1021_n
+ N_VPWR_c_1022_n N_VPWR_c_1023_n N_VPWR_c_1024_n N_VPWR_c_1025_n
+ N_VPWR_c_1010_n PM_SKY130_FD_SC_HS__NOR4BB_4%VPWR
x_PM_SKY130_FD_SC_HS__NOR4BB_4%A_897_349# N_A_897_349#_M1007_s
+ N_A_897_349#_M1032_s N_A_897_349#_M1006_s N_A_897_349#_M1019_s
+ N_A_897_349#_c_1125_n N_A_897_349#_c_1127_n N_A_897_349#_c_1134_n
+ N_A_897_349#_c_1139_n N_A_897_349#_c_1140_n
+ PM_SKY130_FD_SC_HS__NOR4BB_4%A_897_349#
x_PM_SKY130_FD_SC_HS__NOR4BB_4%Y N_Y_M1001_d N_Y_M1017_s N_Y_M1031_s N_Y_M1028_d
+ N_Y_M1009_s N_Y_M1035_s N_Y_M1005_s N_Y_M1030_s N_Y_M1002_d N_Y_M1016_d
+ N_Y_c_1159_n N_Y_c_1176_n N_Y_c_1160_n N_Y_c_1161_n N_Y_c_1207_n N_Y_c_1162_n
+ N_Y_c_1181_n N_Y_c_1163_n N_Y_c_1187_n N_Y_c_1164_n N_Y_c_1222_n N_Y_c_1165_n
+ N_Y_c_1166_n N_Y_c_1167_n N_Y_c_1168_n N_Y_c_1169_n N_Y_c_1174_n N_Y_c_1170_n
+ N_Y_c_1171_n N_Y_c_1268_n N_Y_c_1212_n N_Y_c_1189_n N_Y_c_1194_n N_Y_c_1239_n
+ N_Y_c_1172_n N_Y_c_1280_n Y Y N_Y_c_1284_n PM_SKY130_FD_SC_HS__NOR4BB_4%Y
x_PM_SKY130_FD_SC_HS__NOR4BB_4%VGND N_VGND_M1001_s N_VGND_M1011_d N_VGND_M1023_d
+ N_VGND_M1020_s N_VGND_M1034_s N_VGND_M1014_d N_VGND_M1004_d N_VGND_M1018_d
+ N_VGND_M1036_d N_VGND_M1008_s N_VGND_c_1342_n N_VGND_c_1343_n N_VGND_c_1344_n
+ N_VGND_c_1345_n N_VGND_c_1346_n N_VGND_c_1347_n N_VGND_c_1348_n
+ N_VGND_c_1349_n N_VGND_c_1350_n N_VGND_c_1351_n N_VGND_c_1352_n
+ N_VGND_c_1353_n N_VGND_c_1354_n N_VGND_c_1355_n N_VGND_c_1356_n
+ N_VGND_c_1357_n N_VGND_c_1358_n VGND N_VGND_c_1359_n N_VGND_c_1360_n
+ N_VGND_c_1361_n N_VGND_c_1362_n N_VGND_c_1363_n N_VGND_c_1364_n
+ N_VGND_c_1365_n N_VGND_c_1366_n N_VGND_c_1367_n N_VGND_c_1368_n
+ N_VGND_c_1369_n N_VGND_c_1370_n N_VGND_c_1371_n N_VGND_c_1372_n
+ PM_SKY130_FD_SC_HS__NOR4BB_4%VGND
cc_1 VNB N_B_c_185_n 0.039028f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.765
cc_2 VNB N_B_M1001_g 0.028848f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=0.74
cc_3 VNB N_B_M1020_g 0.0200116f $X=-0.19 $Y=-0.245 $X2=2.985 $Y2=0.74
cc_4 VNB N_B_M1028_g 0.0195717f $X=-0.19 $Y=-0.245 $X2=3.465 $Y2=0.74
cc_5 VNB N_B_M1034_g 0.0192847f $X=-0.19 $Y=-0.245 $X2=3.965 $Y2=0.74
cc_6 VNB N_B_c_190_n 0.0213295f $X=-0.19 $Y=-0.245 $X2=1.085 $Y2=1.485
cc_7 VNB N_B_c_191_n 0.00430013f $X=-0.19 $Y=-0.245 $X2=2.89 $Y2=1.42
cc_8 VNB N_B_c_192_n 8.17781e-19 $X=-0.19 $Y=-0.245 $X2=3.755 $Y2=1.42
cc_9 VNB N_B_c_193_n 0.0554281f $X=-0.19 $Y=-0.245 $X2=3.95 $Y2=1.462
cc_10 VNB N_A_c_305_n 0.0181504f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.765
cc_11 VNB N_A_c_306_n 0.0182597f $X=-0.19 $Y=-0.245 $X2=2.985 $Y2=0.74
cc_12 VNB N_A_c_307_n 0.0181432f $X=-0.19 $Y=-0.245 $X2=3.45 $Y2=2.305
cc_13 VNB N_A_c_308_n 0.018196f $X=-0.19 $Y=-0.245 $X2=3.465 $Y2=0.74
cc_14 VNB N_A_c_309_n 0.0185456f $X=-0.19 $Y=-0.245 $X2=3.95 $Y2=1.67
cc_15 VNB N_A_c_310_n 0.0220391f $X=-0.19 $Y=-0.245 $X2=3.965 $Y2=0.74
cc_16 VNB N_A_c_311_n 0.0785707f $X=-0.19 $Y=-0.245 $X2=0.43 $Y2=1.485
cc_17 VNB N_A_c_312_n 0.00664843f $X=-0.19 $Y=-0.245 $X2=2.72 $Y2=1.795
cc_18 VNB N_A_864_48#_M1009_g 0.019288f $X=-0.19 $Y=-0.245 $X2=2.985 $Y2=0.74
cc_19 VNB N_A_864_48#_M1014_g 0.0203284f $X=-0.19 $Y=-0.245 $X2=3.465 $Y2=0.74
cc_20 VNB N_A_864_48#_M1035_g 0.0200078f $X=-0.19 $Y=-0.245 $X2=3.95 $Y2=2.305
cc_21 VNB N_A_864_48#_c_402_n 0.0153424f $X=-0.19 $Y=-0.245 $X2=3.965 $Y2=1.255
cc_22 VNB N_A_864_48#_c_403_n 0.0187743f $X=-0.19 $Y=-0.245 $X2=0.43 $Y2=1.485
cc_23 VNB N_A_864_48#_c_404_n 0.0157565f $X=-0.19 $Y=-0.245 $X2=3.075 $Y2=1.42
cc_24 VNB N_A_864_48#_c_405_n 0.0116141f $X=-0.19 $Y=-0.245 $X2=3.075 $Y2=1.42
cc_25 VNB N_A_864_48#_c_406_n 4.22572e-19 $X=-0.19 $Y=-0.245 $X2=2.805 $Y2=1.42
cc_26 VNB N_A_864_48#_c_407_n 8.64312e-19 $X=-0.19 $Y=-0.245 $X2=3.465 $Y2=1.462
cc_27 VNB N_A_864_48#_c_408_n 0.0358637f $X=-0.19 $Y=-0.245 $X2=3.755 $Y2=1.462
cc_28 VNB N_A_864_48#_c_409_n 0.0136884f $X=-0.19 $Y=-0.245 $X2=3.95 $Y2=1.462
cc_29 VNB N_A_864_48#_c_410_n 0.0033037f $X=-0.19 $Y=-0.245 $X2=3.965 $Y2=1.462
cc_30 VNB N_A_864_48#_c_411_n 0.00567519f $X=-0.19 $Y=-0.245 $X2=1.2 $Y2=1.795
cc_31 VNB N_A_864_48#_c_412_n 0.03166f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_864_48#_c_413_n 0.0313862f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_1162_48#_M1004_g 0.0200448f $X=-0.19 $Y=-0.245 $X2=2.985 $Y2=0.74
cc_34 VNB N_A_1162_48#_c_581_n 0.00769317f $X=-0.19 $Y=-0.245 $X2=3 $Y2=1.67
cc_35 VNB N_A_1162_48#_c_582_n 0.0111044f $X=-0.19 $Y=-0.245 $X2=3.45 $Y2=2.305
cc_36 VNB N_A_1162_48#_c_583_n 0.00757305f $X=-0.19 $Y=-0.245 $X2=3.465 $Y2=0.74
cc_37 VNB N_A_1162_48#_M1005_g 0.0190494f $X=-0.19 $Y=-0.245 $X2=3.965 $Y2=1.255
cc_38 VNB N_A_1162_48#_c_585_n 0.00968014f $X=-0.19 $Y=-0.245 $X2=3.965 $Y2=0.74
cc_39 VNB N_A_1162_48#_c_586_n 0.0202067f $X=-0.19 $Y=-0.245 $X2=1.085 $Y2=1.485
cc_40 VNB N_A_1162_48#_c_587_n 0.0207538f $X=-0.19 $Y=-0.245 $X2=3.075 $Y2=1.42
cc_41 VNB N_A_1162_48#_c_588_n 0.00621828f $X=-0.19 $Y=-0.245 $X2=3.755 $Y2=1.42
cc_42 VNB N_A_1162_48#_c_589_n 0.00286548f $X=-0.19 $Y=-0.245 $X2=3.755 $Y2=1.42
cc_43 VNB N_A_1162_48#_c_590_n 0.00580254f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_1162_48#_c_591_n 0.0755506f $X=-0.19 $Y=-0.245 $X2=0.452 $Y2=1.485
cc_45 VNB N_A_1162_48#_c_592_n 0.00400717f $X=-0.19 $Y=-0.245 $X2=3 $Y2=1.462
cc_46 VNB N_A_1162_48#_c_593_n 0.0148872f $X=-0.19 $Y=-0.245 $X2=3.95 $Y2=1.462
cc_47 VNB N_A_1162_48#_c_594_n 0.00244505f $X=-0.19 $Y=-0.245 $X2=3.965
+ $Y2=1.462
cc_48 VNB N_A_1162_48#_c_595_n 0.0159898f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A_1162_48#_c_596_n 0.0186198f $X=-0.19 $Y=-0.245 $X2=1.2 $Y2=1.665
cc_50 VNB N_A_1162_48#_c_597_n 0.00413971f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_A_1162_48#_c_598_n 0.0305002f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_A_1162_48#_c_599_n 0.0181746f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_A_1162_48#_c_600_n 0.00907668f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_C_N_M1025_g 0.0446979f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=0.74
cc_55 VNB C_N 0.0121798f $X=-0.19 $Y=-0.245 $X2=3 $Y2=1.67
cc_56 VNB N_C_N_c_774_n 0.0152698f $X=-0.19 $Y=-0.245 $X2=3.465 $Y2=1.255
cc_57 VNB N_D_N_M1008_g 0.0429595f $X=-0.19 $Y=-0.245 $X2=3 $Y2=2.305
cc_58 VNB D_N 0.00304223f $X=-0.19 $Y=-0.245 $X2=3.45 $Y2=1.67
cc_59 VNB N_D_N_c_822_n 0.0389064f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_VPWR_c_1010_n 0.462217f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_Y_c_1159_n 0.00240191f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_Y_c_1160_n 0.00271729f $X=-0.19 $Y=-0.245 $X2=2.89 $Y2=1.42
cc_63 VNB N_Y_c_1161_n 0.00280753f $X=-0.19 $Y=-0.245 $X2=3.075 $Y2=1.42
cc_64 VNB N_Y_c_1162_n 0.00226043f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_Y_c_1163_n 0.00252795f $X=-0.19 $Y=-0.245 $X2=2.985 $Y2=1.462
cc_66 VNB N_Y_c_1164_n 0.00280455f $X=-0.19 $Y=-0.245 $X2=3.95 $Y2=1.462
cc_67 VNB N_Y_c_1165_n 0.00252744f $X=-0.19 $Y=-0.245 $X2=1.2 $Y2=1.795
cc_68 VNB N_Y_c_1166_n 0.00293083f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_Y_c_1167_n 0.00336665f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_Y_c_1168_n 0.00834913f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_Y_c_1169_n 6.82525e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_Y_c_1170_n 0.00240268f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_Y_c_1171_n 0.00126073f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_Y_c_1172_n 0.00235498f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB Y 0.00280987f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_VGND_c_1342_n 0.0122168f $X=-0.19 $Y=-0.245 $X2=0.43 $Y2=1.485
cc_77 VNB N_VGND_c_1343_n 0.0489892f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_VGND_c_1344_n 0.00836159f $X=-0.19 $Y=-0.245 $X2=3.075 $Y2=1.42
cc_79 VNB N_VGND_c_1345_n 0.0186948f $X=-0.19 $Y=-0.245 $X2=3.075 $Y2=1.42
cc_80 VNB N_VGND_c_1346_n 0.00831619f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_81 VNB N_VGND_c_1347_n 0.0183451f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_82 VNB N_VGND_c_1348_n 0.00502317f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_83 VNB N_VGND_c_1349_n 0.0167762f $X=-0.19 $Y=-0.245 $X2=2.985 $Y2=1.462
cc_84 VNB N_VGND_c_1350_n 0.00277973f $X=-0.19 $Y=-0.245 $X2=3.465 $Y2=1.462
cc_85 VNB N_VGND_c_1351_n 0.0185368f $X=-0.19 $Y=-0.245 $X2=3.95 $Y2=1.462
cc_86 VNB N_VGND_c_1352_n 0.00508214f $X=-0.19 $Y=-0.245 $X2=1.2 $Y2=1.665
cc_87 VNB N_VGND_c_1353_n 0.0167762f $X=-0.19 $Y=-0.245 $X2=1.2 $Y2=1.795
cc_88 VNB N_VGND_c_1354_n 0.0076926f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_89 VNB N_VGND_c_1355_n 0.0186948f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_90 VNB N_VGND_c_1356_n 0.0110414f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_91 VNB N_VGND_c_1357_n 0.0111595f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_92 VNB N_VGND_c_1358_n 0.0133782f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_93 VNB N_VGND_c_1359_n 0.0186948f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_94 VNB N_VGND_c_1360_n 0.018682f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_95 VNB N_VGND_c_1361_n 0.0331435f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_96 VNB N_VGND_c_1362_n 0.0173128f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_97 VNB N_VGND_c_1363_n 0.56772f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_98 VNB N_VGND_c_1364_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_99 VNB N_VGND_c_1365_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_100 VNB N_VGND_c_1366_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_101 VNB N_VGND_c_1367_n 0.00604233f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_102 VNB N_VGND_c_1368_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_103 VNB N_VGND_c_1369_n 0.00616716f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_104 VNB N_VGND_c_1370_n 0.0113485f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_105 VNB N_VGND_c_1371_n 0.0104829f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_106 VNB N_VGND_c_1372_n 0.00750435f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_107 VPB N_B_c_185_n 0.0314713f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.765
cc_108 VPB N_B_c_195_n 0.0147015f $X=-0.19 $Y=1.66 $X2=3 $Y2=1.67
cc_109 VPB N_B_c_196_n 0.0145691f $X=-0.19 $Y=1.66 $X2=3.45 $Y2=1.67
cc_110 VPB N_B_c_197_n 0.0150201f $X=-0.19 $Y=1.66 $X2=3.95 $Y2=1.67
cc_111 VPB N_B_c_190_n 0.00142531f $X=-0.19 $Y=1.66 $X2=1.085 $Y2=1.485
cc_112 VPB N_B_c_199_n 0.0114519f $X=-0.19 $Y=1.66 $X2=2.72 $Y2=1.795
cc_113 VPB N_B_c_191_n 0.00290786f $X=-0.19 $Y=1.66 $X2=2.89 $Y2=1.42
cc_114 VPB N_B_c_192_n 3.23044e-19 $X=-0.19 $Y=1.66 $X2=3.755 $Y2=1.42
cc_115 VPB N_B_c_193_n 0.0345899f $X=-0.19 $Y=1.66 $X2=3.95 $Y2=1.462
cc_116 VPB N_A_c_313_n 0.0166277f $X=-0.19 $Y=1.66 $X2=0.565 $Y2=1.32
cc_117 VPB N_A_c_314_n 0.0148198f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_118 VPB N_A_c_315_n 0.0155955f $X=-0.19 $Y=1.66 $X2=3 $Y2=2.305
cc_119 VPB N_A_c_308_n 0.0257012f $X=-0.19 $Y=1.66 $X2=3.465 $Y2=0.74
cc_120 VPB N_A_c_311_n 0.0191276f $X=-0.19 $Y=1.66 $X2=0.43 $Y2=1.485
cc_121 VPB N_A_864_48#_c_414_n 0.0144781f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_122 VPB N_A_864_48#_c_415_n 0.0153682f $X=-0.19 $Y=1.66 $X2=3 $Y2=2.305
cc_123 VPB N_A_864_48#_c_402_n 0.02489f $X=-0.19 $Y=1.66 $X2=3.965 $Y2=1.255
cc_124 VPB N_A_864_48#_c_417_n 0.018222f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_125 VPB N_A_864_48#_c_404_n 0.0158639f $X=-0.19 $Y=1.66 $X2=3.075 $Y2=1.42
cc_126 VPB N_A_864_48#_c_405_n 0.00860839f $X=-0.19 $Y=1.66 $X2=3.075 $Y2=1.42
cc_127 VPB N_A_864_48#_c_420_n 0.00308062f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_128 VPB N_A_864_48#_c_421_n 0.00841225f $X=-0.19 $Y=1.66 $X2=0.452 $Y2=1.485
cc_129 VPB N_A_864_48#_c_422_n 0.00121417f $X=-0.19 $Y=1.66 $X2=2.985 $Y2=1.462
cc_130 VPB N_A_864_48#_c_407_n 0.0023849f $X=-0.19 $Y=1.66 $X2=3.465 $Y2=1.462
cc_131 VPB N_A_864_48#_c_424_n 0.00568661f $X=-0.19 $Y=1.66 $X2=1.2 $Y2=1.485
cc_132 VPB N_A_864_48#_c_425_n 0.00239217f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_133 VPB N_A_864_48#_c_426_n 0.0186483f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_134 VPB N_A_864_48#_c_412_n 0.0217304f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_135 VPB N_A_1162_48#_c_581_n 7.11257e-19 $X=-0.19 $Y=1.66 $X2=3 $Y2=1.67
cc_136 VPB N_A_1162_48#_c_602_n 0.0196116f $X=-0.19 $Y=1.66 $X2=3 $Y2=2.305
cc_137 VPB N_A_1162_48#_c_583_n 6.92077e-19 $X=-0.19 $Y=1.66 $X2=3.465 $Y2=0.74
cc_138 VPB N_A_1162_48#_c_604_n 0.0191294f $X=-0.19 $Y=1.66 $X2=3.465 $Y2=0.74
cc_139 VPB N_A_1162_48#_c_605_n 0.0140991f $X=-0.19 $Y=1.66 $X2=0.43 $Y2=1.485
cc_140 VPB N_A_1162_48#_c_606_n 0.0163215f $X=-0.19 $Y=1.66 $X2=1.315 $Y2=1.795
cc_141 VPB N_A_1162_48#_c_591_n 0.0141641f $X=-0.19 $Y=1.66 $X2=0.452 $Y2=1.485
cc_142 VPB N_A_1162_48#_c_608_n 0.00216998f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_143 VPB N_A_1162_48#_c_609_n 0.0137844f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_144 VPB N_A_1162_48#_c_610_n 0.00176996f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_145 VPB N_A_1162_48#_c_599_n 0.013841f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_146 VPB N_C_N_c_775_n 0.0174096f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.765
cc_147 VPB N_C_N_c_776_n 0.0156052f $X=-0.19 $Y=1.66 $X2=2.985 $Y2=1.255
cc_148 VPB C_N 0.00798441f $X=-0.19 $Y=1.66 $X2=3 $Y2=1.67
cc_149 VPB N_C_N_c_774_n 0.0543254f $X=-0.19 $Y=1.66 $X2=3.465 $Y2=1.255
cc_150 VPB N_D_N_c_823_n 0.00940528f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.4
cc_151 VPB N_D_N_c_824_n 0.0214216f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.4
cc_152 VPB N_D_N_c_825_n 0.00996055f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_153 VPB N_D_N_c_826_n 0.0237077f $X=-0.19 $Y=1.66 $X2=2.985 $Y2=1.255
cc_154 VPB D_N 8.33115e-19 $X=-0.19 $Y=1.66 $X2=3.45 $Y2=1.67
cc_155 VPB N_D_N_c_822_n 0.0163849f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_156 VPB N_A_27_368#_c_863_n 0.0315989f $X=-0.19 $Y=1.66 $X2=3.465 $Y2=1.255
cc_157 VPB N_A_27_368#_c_864_n 6.86314e-19 $X=-0.19 $Y=1.66 $X2=0.43 $Y2=1.485
cc_158 VPB N_A_27_368#_c_865_n 0.057648f $X=-0.19 $Y=1.66 $X2=0.43 $Y2=1.485
cc_159 VPB N_A_27_368#_c_866_n 0.00299413f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_160 VPB N_A_27_368#_c_867_n 9.30091e-19 $X=-0.19 $Y=1.66 $X2=3.075 $Y2=1.42
cc_161 VPB N_A_27_368#_c_868_n 0.0223071f $X=-0.19 $Y=1.66 $X2=3.755 $Y2=1.42
cc_162 VPB N_A_116_368#_c_949_n 0.00216476f $X=-0.19 $Y=1.66 $X2=3.465 $Y2=0.74
cc_163 VPB N_A_116_368#_c_950_n 3.2727e-19 $X=-0.19 $Y=1.66 $X2=3.95 $Y2=2.305
cc_164 VPB N_A_116_368#_c_951_n 0.0130805f $X=-0.19 $Y=1.66 $X2=3.965 $Y2=1.255
cc_165 VPB N_A_116_368#_c_952_n 0.00300498f $X=-0.19 $Y=1.66 $X2=3.965 $Y2=0.74
cc_166 VPB N_A_116_368#_c_953_n 3.27053e-19 $X=-0.19 $Y=1.66 $X2=1.085 $Y2=1.485
cc_167 VPB N_A_116_368#_c_954_n 0.00289021f $X=-0.19 $Y=1.66 $X2=0.43 $Y2=1.485
cc_168 VPB N_VPWR_c_1011_n 0.00590893f $X=-0.19 $Y=1.66 $X2=3.465 $Y2=1.255
cc_169 VPB N_VPWR_c_1012_n 0.00614703f $X=-0.19 $Y=1.66 $X2=3.95 $Y2=1.67
cc_170 VPB N_VPWR_c_1013_n 0.0065445f $X=-0.19 $Y=1.66 $X2=3.965 $Y2=0.74
cc_171 VPB N_VPWR_c_1014_n 0.0184891f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_172 VPB N_VPWR_c_1015_n 0.00886271f $X=-0.19 $Y=1.66 $X2=0.43 $Y2=1.485
cc_173 VPB N_VPWR_c_1016_n 0.0120106f $X=-0.19 $Y=1.66 $X2=2.72 $Y2=1.795
cc_174 VPB N_VPWR_c_1017_n 0.0351405f $X=-0.19 $Y=1.66 $X2=2.89 $Y2=1.42
cc_175 VPB N_VPWR_c_1018_n 0.0325002f $X=-0.19 $Y=1.66 $X2=3.755 $Y2=1.42
cc_176 VPB N_VPWR_c_1019_n 0.0175706f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_177 VPB N_VPWR_c_1020_n 0.148862f $X=-0.19 $Y=1.66 $X2=0.452 $Y2=1.485
cc_178 VPB N_VPWR_c_1021_n 0.0185253f $X=-0.19 $Y=1.66 $X2=3.965 $Y2=1.462
cc_179 VPB N_VPWR_c_1022_n 0.00614151f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_180 VPB N_VPWR_c_1023_n 0.00691093f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_181 VPB N_VPWR_c_1024_n 0.00614589f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_182 VPB N_VPWR_c_1025_n 0.00324402f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_183 VPB N_VPWR_c_1010_n 0.133222f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_184 VPB N_Y_c_1174_n 0.00488297f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_185 N_B_M1001_g N_A_c_305_n 0.0115403f $X=0.565 $Y=0.74 $X2=-0.19 $Y2=-0.245
cc_186 N_B_c_185_n N_A_c_313_n 0.0320099f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_187 N_B_c_190_n N_A_c_313_n 0.00206195f $X=1.085 $Y=1.485 $X2=0 $Y2=0
cc_188 N_B_c_199_n N_A_c_314_n 0.00598814f $X=2.72 $Y=1.795 $X2=0 $Y2=0
cc_189 N_B_c_199_n N_A_c_315_n 0.00674481f $X=2.72 $Y=1.795 $X2=0 $Y2=0
cc_190 N_B_c_195_n N_A_c_308_n 0.0341835f $X=3 $Y=1.67 $X2=0 $Y2=0
cc_191 N_B_c_199_n N_A_c_308_n 0.0153288f $X=2.72 $Y=1.795 $X2=0 $Y2=0
cc_192 N_B_c_191_n N_A_c_308_n 0.00661169f $X=2.89 $Y=1.42 $X2=0 $Y2=0
cc_193 N_B_c_193_n N_A_c_308_n 0.015851f $X=3.95 $Y=1.462 $X2=0 $Y2=0
cc_194 N_B_M1020_g N_A_c_309_n 0.0121945f $X=2.985 $Y=0.74 $X2=0 $Y2=0
cc_195 N_B_c_199_n N_A_c_310_n 0.00418282f $X=2.72 $Y=1.795 $X2=0 $Y2=0
cc_196 N_B_c_185_n N_A_c_311_n 0.0264328f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_197 N_B_c_190_n N_A_c_311_n 0.0412963f $X=1.085 $Y=1.485 $X2=0 $Y2=0
cc_198 N_B_c_199_n N_A_c_311_n 0.0147463f $X=2.72 $Y=1.795 $X2=0 $Y2=0
cc_199 N_B_M1020_g N_A_c_312_n 3.59919e-19 $X=2.985 $Y=0.74 $X2=0 $Y2=0
cc_200 N_B_c_190_n N_A_c_312_n 0.0170371f $X=1.085 $Y=1.485 $X2=0 $Y2=0
cc_201 N_B_c_199_n N_A_c_312_n 0.0749231f $X=2.72 $Y=1.795 $X2=0 $Y2=0
cc_202 N_B_c_191_n N_A_c_312_n 0.0183579f $X=2.89 $Y=1.42 $X2=0 $Y2=0
cc_203 N_B_M1034_g N_A_864_48#_M1009_g 0.0247844f $X=3.965 $Y=0.74 $X2=0 $Y2=0
cc_204 N_B_c_197_n N_A_864_48#_c_414_n 0.00838353f $X=3.95 $Y=1.67 $X2=0 $Y2=0
cc_205 N_B_c_192_n N_A_864_48#_c_430_n 0.0131687f $X=3.755 $Y=1.42 $X2=0 $Y2=0
cc_206 N_B_c_193_n N_A_864_48#_c_430_n 0.00149213f $X=3.95 $Y=1.462 $X2=0 $Y2=0
cc_207 N_B_c_192_n N_A_864_48#_c_412_n 0.00123555f $X=3.755 $Y=1.42 $X2=0 $Y2=0
cc_208 N_B_c_193_n N_A_864_48#_c_412_n 0.0247844f $X=3.95 $Y=1.462 $X2=0 $Y2=0
cc_209 N_B_c_185_n N_A_27_368#_c_863_n 0.00979381f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_210 N_B_c_185_n N_A_27_368#_c_870_n 0.014025f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_211 N_B_c_195_n N_A_27_368#_c_870_n 0.0146606f $X=3 $Y=1.67 $X2=0 $Y2=0
cc_212 N_B_c_190_n N_A_27_368#_c_870_n 0.0369916f $X=1.085 $Y=1.485 $X2=0 $Y2=0
cc_213 N_B_c_199_n N_A_27_368#_c_870_n 0.0750254f $X=2.72 $Y=1.795 $X2=0 $Y2=0
cc_214 N_B_c_191_n N_A_27_368#_c_870_n 0.0118777f $X=2.89 $Y=1.42 $X2=0 $Y2=0
cc_215 N_B_c_192_n N_A_27_368#_c_870_n 0.00492396f $X=3.755 $Y=1.42 $X2=0 $Y2=0
cc_216 N_B_c_195_n N_A_27_368#_c_876_n 0.00664619f $X=3 $Y=1.67 $X2=0 $Y2=0
cc_217 N_B_c_196_n N_A_27_368#_c_876_n 0.00508464f $X=3.45 $Y=1.67 $X2=0 $Y2=0
cc_218 N_B_c_196_n N_A_27_368#_c_878_n 0.0133259f $X=3.45 $Y=1.67 $X2=0 $Y2=0
cc_219 N_B_c_197_n N_A_27_368#_c_878_n 0.0145383f $X=3.95 $Y=1.67 $X2=0 $Y2=0
cc_220 N_B_c_192_n N_A_27_368#_c_878_n 0.0345575f $X=3.755 $Y=1.42 $X2=0 $Y2=0
cc_221 N_B_c_193_n N_A_27_368#_c_878_n 0.00758128f $X=3.95 $Y=1.462 $X2=0 $Y2=0
cc_222 N_B_c_197_n N_A_27_368#_c_864_n 0.00610799f $X=3.95 $Y=1.67 $X2=0 $Y2=0
cc_223 N_B_c_197_n N_A_27_368#_c_866_n 7.99395e-19 $X=3.95 $Y=1.67 $X2=0 $Y2=0
cc_224 N_B_c_185_n N_A_27_368#_c_868_n 0.010049f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_225 N_B_c_190_n N_A_27_368#_c_868_n 0.0160704f $X=1.085 $Y=1.485 $X2=0 $Y2=0
cc_226 N_B_c_195_n N_A_27_368#_c_886_n 0.00527979f $X=3 $Y=1.67 $X2=0 $Y2=0
cc_227 N_B_c_196_n N_A_27_368#_c_886_n 0.00527418f $X=3.45 $Y=1.67 $X2=0 $Y2=0
cc_228 N_B_c_197_n N_A_27_368#_c_886_n 9.80037e-19 $X=3.95 $Y=1.67 $X2=0 $Y2=0
cc_229 N_B_c_192_n N_A_27_368#_c_886_n 0.0218087f $X=3.755 $Y=1.42 $X2=0 $Y2=0
cc_230 N_B_c_193_n N_A_27_368#_c_886_n 0.00650717f $X=3.95 $Y=1.462 $X2=0 $Y2=0
cc_231 N_B_c_199_n N_A_116_368#_M1022_s 0.00198204f $X=2.72 $Y=1.795 $X2=0 $Y2=0
cc_232 N_B_c_199_n N_A_116_368#_M1033_s 0.00131601f $X=2.72 $Y=1.795 $X2=0 $Y2=0
cc_233 N_B_c_191_n N_A_116_368#_M1033_s 0.00255839f $X=2.89 $Y=1.42 $X2=0 $Y2=0
cc_234 N_B_c_195_n N_A_116_368#_c_950_n 0.00221804f $X=3 $Y=1.67 $X2=0 $Y2=0
cc_235 N_B_c_195_n N_A_116_368#_c_951_n 0.0119646f $X=3 $Y=1.67 $X2=0 $Y2=0
cc_236 N_B_c_196_n N_A_116_368#_c_951_n 0.0122229f $X=3.45 $Y=1.67 $X2=0 $Y2=0
cc_237 N_B_c_197_n N_A_116_368#_c_951_n 0.00243878f $X=3.95 $Y=1.67 $X2=0 $Y2=0
cc_238 N_B_c_196_n N_A_116_368#_c_953_n 0.00471804f $X=3.45 $Y=1.67 $X2=0 $Y2=0
cc_239 N_B_c_197_n N_A_116_368#_c_953_n 0.00973697f $X=3.95 $Y=1.67 $X2=0 $Y2=0
cc_240 N_B_c_185_n N_A_116_368#_c_954_n 0.00229911f $X=0.505 $Y=1.765 $X2=0
+ $Y2=0
cc_241 N_B_c_190_n N_VPWR_M1021_d 0.00204483f $X=1.085 $Y=1.485 $X2=-0.19
+ $Y2=-0.245
cc_242 N_B_c_199_n N_VPWR_M1021_d 7.14335e-19 $X=2.72 $Y=1.795 $X2=-0.19
+ $Y2=-0.245
cc_243 N_B_c_199_n N_VPWR_M1024_d 0.00294109f $X=2.72 $Y=1.795 $X2=0 $Y2=0
cc_244 N_B_c_185_n N_VPWR_c_1018_n 0.00445602f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_245 N_B_c_195_n N_VPWR_c_1020_n 7.74126e-19 $X=3 $Y=1.67 $X2=0 $Y2=0
cc_246 N_B_c_196_n N_VPWR_c_1020_n 7.74126e-19 $X=3.45 $Y=1.67 $X2=0 $Y2=0
cc_247 N_B_c_197_n N_VPWR_c_1020_n 0.00467123f $X=3.95 $Y=1.67 $X2=0 $Y2=0
cc_248 N_B_c_185_n N_VPWR_c_1010_n 0.0086236f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_249 N_B_c_197_n N_VPWR_c_1010_n 0.00464368f $X=3.95 $Y=1.67 $X2=0 $Y2=0
cc_250 N_B_M1001_g N_Y_c_1159_n 0.00637485f $X=0.565 $Y=0.74 $X2=0 $Y2=0
cc_251 N_B_c_190_n N_Y_c_1176_n 0.0159768f $X=1.085 $Y=1.485 $X2=0 $Y2=0
cc_252 N_B_M1001_g N_Y_c_1160_n 0.00370932f $X=0.565 $Y=0.74 $X2=0 $Y2=0
cc_253 N_B_c_190_n N_Y_c_1160_n 0.0265437f $X=1.085 $Y=1.485 $X2=0 $Y2=0
cc_254 N_B_M1020_g N_Y_c_1162_n 0.00541476f $X=2.985 $Y=0.74 $X2=0 $Y2=0
cc_255 N_B_M1028_g N_Y_c_1162_n 4.79174e-19 $X=3.465 $Y=0.74 $X2=0 $Y2=0
cc_256 N_B_M1020_g N_Y_c_1181_n 0.0127242f $X=2.985 $Y=0.74 $X2=0 $Y2=0
cc_257 N_B_M1028_g N_Y_c_1181_n 0.0123838f $X=3.465 $Y=0.74 $X2=0 $Y2=0
cc_258 N_B_c_192_n N_Y_c_1181_n 0.0432892f $X=3.755 $Y=1.42 $X2=0 $Y2=0
cc_259 N_B_c_193_n N_Y_c_1181_n 0.00336308f $X=3.95 $Y=1.462 $X2=0 $Y2=0
cc_260 N_B_M1028_g N_Y_c_1163_n 2.39553e-19 $X=3.465 $Y=0.74 $X2=0 $Y2=0
cc_261 N_B_M1034_g N_Y_c_1163_n 0.00300429f $X=3.965 $Y=0.74 $X2=0 $Y2=0
cc_262 N_B_M1034_g N_Y_c_1187_n 0.0163097f $X=3.965 $Y=0.74 $X2=0 $Y2=0
cc_263 N_B_c_192_n N_Y_c_1187_n 0.00383088f $X=3.755 $Y=1.42 $X2=0 $Y2=0
cc_264 N_B_M1020_g N_Y_c_1189_n 0.00149831f $X=2.985 $Y=0.74 $X2=0 $Y2=0
cc_265 N_B_M1028_g N_Y_c_1189_n 3.42471e-19 $X=3.465 $Y=0.74 $X2=0 $Y2=0
cc_266 N_B_c_199_n N_Y_c_1189_n 0.00173114f $X=2.72 $Y=1.795 $X2=0 $Y2=0
cc_267 N_B_c_191_n N_Y_c_1189_n 0.0137221f $X=2.89 $Y=1.42 $X2=0 $Y2=0
cc_268 N_B_c_192_n N_Y_c_1189_n 0.00119318f $X=3.755 $Y=1.42 $X2=0 $Y2=0
cc_269 N_B_c_192_n N_Y_c_1194_n 0.020017f $X=3.755 $Y=1.42 $X2=0 $Y2=0
cc_270 N_B_c_193_n N_Y_c_1194_n 0.00396026f $X=3.95 $Y=1.462 $X2=0 $Y2=0
cc_271 N_B_c_185_n N_VGND_c_1343_n 0.00420326f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_272 N_B_M1001_g N_VGND_c_1343_n 0.0184904f $X=0.565 $Y=0.74 $X2=0 $Y2=0
cc_273 N_B_c_190_n N_VGND_c_1343_n 0.0138849f $X=1.085 $Y=1.485 $X2=0 $Y2=0
cc_274 N_B_M1020_g N_VGND_c_1347_n 0.00456932f $X=2.985 $Y=0.74 $X2=0 $Y2=0
cc_275 N_B_M1020_g N_VGND_c_1348_n 0.00195929f $X=2.985 $Y=0.74 $X2=0 $Y2=0
cc_276 N_B_M1028_g N_VGND_c_1348_n 0.00870655f $X=3.465 $Y=0.74 $X2=0 $Y2=0
cc_277 N_B_M1034_g N_VGND_c_1348_n 4.36693e-19 $X=3.965 $Y=0.74 $X2=0 $Y2=0
cc_278 N_B_M1028_g N_VGND_c_1349_n 0.00383152f $X=3.465 $Y=0.74 $X2=0 $Y2=0
cc_279 N_B_M1034_g N_VGND_c_1349_n 0.00383152f $X=3.965 $Y=0.74 $X2=0 $Y2=0
cc_280 N_B_M1028_g N_VGND_c_1350_n 4.31571e-19 $X=3.465 $Y=0.74 $X2=0 $Y2=0
cc_281 N_B_M1034_g N_VGND_c_1350_n 0.00862521f $X=3.965 $Y=0.74 $X2=0 $Y2=0
cc_282 N_B_M1001_g N_VGND_c_1359_n 0.00434272f $X=0.565 $Y=0.74 $X2=0 $Y2=0
cc_283 N_B_M1001_g N_VGND_c_1363_n 0.00824032f $X=0.565 $Y=0.74 $X2=0 $Y2=0
cc_284 N_B_M1020_g N_VGND_c_1363_n 0.00889961f $X=2.985 $Y=0.74 $X2=0 $Y2=0
cc_285 N_B_M1028_g N_VGND_c_1363_n 0.00758198f $X=3.465 $Y=0.74 $X2=0 $Y2=0
cc_286 N_B_M1034_g N_VGND_c_1363_n 0.00758198f $X=3.965 $Y=0.74 $X2=0 $Y2=0
cc_287 N_A_c_313_n N_A_27_368#_c_870_n 0.0124477f $X=1.005 $Y=1.765 $X2=0 $Y2=0
cc_288 N_A_c_314_n N_A_27_368#_c_870_n 0.0110058f $X=1.505 $Y=1.765 $X2=0 $Y2=0
cc_289 N_A_c_315_n N_A_27_368#_c_870_n 0.0111989f $X=1.955 $Y=1.765 $X2=0 $Y2=0
cc_290 N_A_c_308_n N_A_27_368#_c_870_n 0.0114366f $X=2.495 $Y=1.765 $X2=0 $Y2=0
cc_291 N_A_c_311_n N_A_27_368#_c_870_n 4.73237e-19 $X=2.07 $Y=1.385 $X2=0 $Y2=0
cc_292 N_A_c_313_n N_A_27_368#_c_868_n 0.00159209f $X=1.005 $Y=1.765 $X2=0 $Y2=0
cc_293 N_A_c_308_n N_A_27_368#_c_886_n 0.00159206f $X=2.495 $Y=1.765 $X2=0 $Y2=0
cc_294 N_A_c_313_n N_A_116_368#_c_965_n 0.00923282f $X=1.005 $Y=1.765 $X2=0
+ $Y2=0
cc_295 N_A_c_314_n N_A_116_368#_c_965_n 0.00988709f $X=1.505 $Y=1.765 $X2=0
+ $Y2=0
cc_296 N_A_c_314_n N_A_116_368#_c_949_n 0.00454039f $X=1.505 $Y=1.765 $X2=0
+ $Y2=0
cc_297 N_A_c_315_n N_A_116_368#_c_949_n 0.00586411f $X=1.955 $Y=1.765 $X2=0
+ $Y2=0
cc_298 N_A_c_308_n N_A_116_368#_c_949_n 5.75503e-19 $X=2.495 $Y=1.765 $X2=0
+ $Y2=0
cc_299 N_A_c_315_n N_A_116_368#_c_970_n 0.00942648f $X=1.955 $Y=1.765 $X2=0
+ $Y2=0
cc_300 N_A_c_308_n N_A_116_368#_c_970_n 0.0100808f $X=2.495 $Y=1.765 $X2=0 $Y2=0
cc_301 N_A_c_308_n N_A_116_368#_c_950_n 0.00497595f $X=2.495 $Y=1.765 $X2=0
+ $Y2=0
cc_302 N_A_c_308_n N_A_116_368#_c_952_n 0.0027197f $X=2.495 $Y=1.765 $X2=0 $Y2=0
cc_303 N_A_c_313_n N_A_116_368#_c_954_n 0.00630231f $X=1.005 $Y=1.765 $X2=0
+ $Y2=0
cc_304 N_A_c_314_n N_A_116_368#_c_954_n 6.00298e-19 $X=1.505 $Y=1.765 $X2=0
+ $Y2=0
cc_305 N_A_c_315_n N_A_116_368#_c_976_n 4.11408e-19 $X=1.955 $Y=1.765 $X2=0
+ $Y2=0
cc_306 N_A_c_313_n N_VPWR_c_1011_n 0.00452824f $X=1.005 $Y=1.765 $X2=0 $Y2=0
cc_307 N_A_c_314_n N_VPWR_c_1011_n 0.00658099f $X=1.505 $Y=1.765 $X2=0 $Y2=0
cc_308 N_A_c_315_n N_VPWR_c_1011_n 4.17603e-19 $X=1.955 $Y=1.765 $X2=0 $Y2=0
cc_309 N_A_c_315_n N_VPWR_c_1012_n 0.0032886f $X=1.955 $Y=1.765 $X2=0 $Y2=0
cc_310 N_A_c_308_n N_VPWR_c_1012_n 0.00632774f $X=2.495 $Y=1.765 $X2=0 $Y2=0
cc_311 N_A_c_313_n N_VPWR_c_1018_n 0.00445602f $X=1.005 $Y=1.765 $X2=0 $Y2=0
cc_312 N_A_c_314_n N_VPWR_c_1019_n 0.00413917f $X=1.505 $Y=1.765 $X2=0 $Y2=0
cc_313 N_A_c_315_n N_VPWR_c_1019_n 0.00445602f $X=1.955 $Y=1.765 $X2=0 $Y2=0
cc_314 N_A_c_308_n N_VPWR_c_1020_n 0.00413917f $X=2.495 $Y=1.765 $X2=0 $Y2=0
cc_315 N_A_c_313_n N_VPWR_c_1010_n 0.00437274f $X=1.005 $Y=1.765 $X2=0 $Y2=0
cc_316 N_A_c_314_n N_VPWR_c_1010_n 0.00398641f $X=1.505 $Y=1.765 $X2=0 $Y2=0
cc_317 N_A_c_315_n N_VPWR_c_1010_n 0.00437098f $X=1.955 $Y=1.765 $X2=0 $Y2=0
cc_318 N_A_c_308_n N_VPWR_c_1010_n 0.00403443f $X=2.495 $Y=1.765 $X2=0 $Y2=0
cc_319 N_A_c_305_n N_Y_c_1159_n 0.00784719f $X=0.995 $Y=1.22 $X2=0 $Y2=0
cc_320 N_A_c_306_n N_Y_c_1159_n 4.2483e-19 $X=1.52 $Y=1.22 $X2=0 $Y2=0
cc_321 N_A_c_305_n N_Y_c_1176_n 0.0097007f $X=0.995 $Y=1.22 $X2=0 $Y2=0
cc_322 N_A_c_306_n N_Y_c_1176_n 0.0115834f $X=1.52 $Y=1.22 $X2=0 $Y2=0
cc_323 N_A_c_311_n N_Y_c_1176_n 0.00520288f $X=2.07 $Y=1.385 $X2=0 $Y2=0
cc_324 N_A_c_312_n N_Y_c_1176_n 0.00872056f $X=2.33 $Y=1.385 $X2=0 $Y2=0
cc_325 N_A_c_305_n N_Y_c_1160_n 0.00336331f $X=0.995 $Y=1.22 $X2=0 $Y2=0
cc_326 N_A_c_306_n N_Y_c_1160_n 5.61187e-19 $X=1.52 $Y=1.22 $X2=0 $Y2=0
cc_327 N_A_c_306_n N_Y_c_1161_n 2.72399e-19 $X=1.52 $Y=1.22 $X2=0 $Y2=0
cc_328 N_A_c_307_n N_Y_c_1161_n 0.00733959f $X=1.995 $Y=1.22 $X2=0 $Y2=0
cc_329 N_A_c_309_n N_Y_c_1161_n 6.72946e-19 $X=2.535 $Y=1.22 $X2=0 $Y2=0
cc_330 N_A_c_307_n N_Y_c_1207_n 0.0091168f $X=1.995 $Y=1.22 $X2=0 $Y2=0
cc_331 N_A_c_309_n N_Y_c_1207_n 0.0138617f $X=2.535 $Y=1.22 $X2=0 $Y2=0
cc_332 N_A_c_310_n N_Y_c_1207_n 0.0013216f $X=2.405 $Y=1.385 $X2=0 $Y2=0
cc_333 N_A_c_312_n N_Y_c_1207_n 0.0379485f $X=2.33 $Y=1.385 $X2=0 $Y2=0
cc_334 N_A_c_309_n N_Y_c_1162_n 2.29378e-19 $X=2.535 $Y=1.22 $X2=0 $Y2=0
cc_335 N_A_c_307_n N_Y_c_1212_n 7.17169e-19 $X=1.995 $Y=1.22 $X2=0 $Y2=0
cc_336 N_A_c_311_n N_Y_c_1212_n 0.00101923f $X=2.07 $Y=1.385 $X2=0 $Y2=0
cc_337 N_A_c_312_n N_Y_c_1212_n 0.0243104f $X=2.33 $Y=1.385 $X2=0 $Y2=0
cc_338 N_A_c_305_n N_VGND_c_1344_n 0.00357681f $X=0.995 $Y=1.22 $X2=0 $Y2=0
cc_339 N_A_c_306_n N_VGND_c_1344_n 0.00209449f $X=1.52 $Y=1.22 $X2=0 $Y2=0
cc_340 N_A_c_306_n N_VGND_c_1345_n 0.00460063f $X=1.52 $Y=1.22 $X2=0 $Y2=0
cc_341 N_A_c_307_n N_VGND_c_1345_n 0.00434272f $X=1.995 $Y=1.22 $X2=0 $Y2=0
cc_342 N_A_c_307_n N_VGND_c_1346_n 0.00365613f $X=1.995 $Y=1.22 $X2=0 $Y2=0
cc_343 N_A_c_309_n N_VGND_c_1346_n 0.00204108f $X=2.535 $Y=1.22 $X2=0 $Y2=0
cc_344 N_A_c_309_n N_VGND_c_1347_n 0.00461464f $X=2.535 $Y=1.22 $X2=0 $Y2=0
cc_345 N_A_c_305_n N_VGND_c_1359_n 0.00434272f $X=0.995 $Y=1.22 $X2=0 $Y2=0
cc_346 N_A_c_305_n N_VGND_c_1363_n 0.00445807f $X=0.995 $Y=1.22 $X2=0 $Y2=0
cc_347 N_A_c_306_n N_VGND_c_1363_n 0.00463677f $X=1.52 $Y=1.22 $X2=0 $Y2=0
cc_348 N_A_c_307_n N_VGND_c_1363_n 0.00446267f $X=1.995 $Y=1.22 $X2=0 $Y2=0
cc_349 N_A_c_309_n N_VGND_c_1363_n 0.00463984f $X=2.535 $Y=1.22 $X2=0 $Y2=0
cc_350 N_A_864_48#_M1035_g N_A_1162_48#_M1004_g 0.0183805f $X=5.395 $Y=0.74
+ $X2=0 $Y2=0
cc_351 N_A_864_48#_c_402_n N_A_1162_48#_c_581_n 0.0125304f $X=5.48 $Y=1.67 $X2=0
+ $Y2=0
cc_352 N_A_864_48#_c_406_n N_A_1162_48#_c_581_n 3.39552e-19 $X=5.27 $Y=1.585
+ $X2=0 $Y2=0
cc_353 N_A_864_48#_c_402_n N_A_1162_48#_c_602_n 0.0384046f $X=5.48 $Y=1.67 $X2=0
+ $Y2=0
cc_354 N_A_864_48#_c_438_p N_A_1162_48#_c_602_n 0.0147903f $X=7.4 $Y=2.31 $X2=0
+ $Y2=0
cc_355 N_A_864_48#_c_438_p N_A_1162_48#_c_604_n 0.0107759f $X=7.4 $Y=2.31 $X2=0
+ $Y2=0
cc_356 N_A_864_48#_c_438_p N_A_1162_48#_c_605_n 0.0107391f $X=7.4 $Y=2.31 $X2=0
+ $Y2=0
cc_357 N_A_864_48#_c_417_n N_A_1162_48#_c_606_n 0.00918158f $X=8.095 $Y=1.67
+ $X2=0 $Y2=0
cc_358 N_A_864_48#_c_438_p N_A_1162_48#_c_606_n 0.0131369f $X=7.4 $Y=2.31 $X2=0
+ $Y2=0
cc_359 N_A_864_48#_c_422_n N_A_1162_48#_c_606_n 0.00159297f $X=7.57 $Y=1.81
+ $X2=0 $Y2=0
cc_360 N_A_864_48#_c_403_n N_A_1162_48#_c_587_n 0.0105422f $X=8.11 $Y=1.22 $X2=0
+ $Y2=0
cc_361 N_A_864_48#_c_405_n N_A_1162_48#_c_587_n 2.49057e-19 $X=8.095 $Y=1.445
+ $X2=0 $Y2=0
cc_362 N_A_864_48#_c_402_n N_A_1162_48#_c_588_n 0.00831798f $X=5.48 $Y=1.67
+ $X2=0 $Y2=0
cc_363 N_A_864_48#_c_405_n N_A_1162_48#_c_590_n 0.0183882f $X=8.095 $Y=1.445
+ $X2=0 $Y2=0
cc_364 N_A_864_48#_c_438_p N_A_1162_48#_c_590_n 0.00348077f $X=7.4 $Y=2.31 $X2=0
+ $Y2=0
cc_365 N_A_864_48#_c_421_n N_A_1162_48#_c_590_n 0.0624317f $X=8.545 $Y=1.81
+ $X2=0 $Y2=0
cc_366 N_A_864_48#_c_422_n N_A_1162_48#_c_590_n 0.014319f $X=7.57 $Y=1.81 $X2=0
+ $Y2=0
cc_367 N_A_864_48#_c_407_n N_A_1162_48#_c_590_n 0.0156389f $X=8.71 $Y=1.385
+ $X2=0 $Y2=0
cc_368 N_A_864_48#_c_410_n N_A_1162_48#_c_590_n 0.0114279f $X=8.875 $Y=1.275
+ $X2=0 $Y2=0
cc_369 N_A_864_48#_c_413_n N_A_1162_48#_c_590_n 0.0133498f $X=8.545 $Y=1.385
+ $X2=0 $Y2=0
cc_370 N_A_864_48#_c_405_n N_A_1162_48#_c_591_n 0.0244702f $X=8.095 $Y=1.445
+ $X2=0 $Y2=0
cc_371 N_A_864_48#_c_421_n N_A_1162_48#_c_591_n 0.00567282f $X=8.545 $Y=1.81
+ $X2=0 $Y2=0
cc_372 N_A_864_48#_c_422_n N_A_1162_48#_c_591_n 0.00426736f $X=7.57 $Y=1.81
+ $X2=0 $Y2=0
cc_373 N_A_864_48#_c_403_n N_A_1162_48#_c_592_n 0.0061889f $X=8.11 $Y=1.22 $X2=0
+ $Y2=0
cc_374 N_A_864_48#_c_410_n N_A_1162_48#_c_592_n 0.00288052f $X=8.875 $Y=1.275
+ $X2=0 $Y2=0
cc_375 N_A_864_48#_c_413_n N_A_1162_48#_c_592_n 0.00361137f $X=8.545 $Y=1.385
+ $X2=0 $Y2=0
cc_376 N_A_864_48#_c_408_n N_A_1162_48#_c_638_n 0.00213653f $X=8.71 $Y=1.385
+ $X2=0 $Y2=0
cc_377 N_A_864_48#_c_409_n N_A_1162_48#_c_638_n 0.0165488f $X=9.26 $Y=1.275
+ $X2=0 $Y2=0
cc_378 N_A_864_48#_c_410_n N_A_1162_48#_c_638_n 0.0274729f $X=8.875 $Y=1.275
+ $X2=0 $Y2=0
cc_379 N_A_864_48#_c_413_n N_A_1162_48#_c_638_n 0.00611177f $X=8.545 $Y=1.385
+ $X2=0 $Y2=0
cc_380 N_A_864_48#_M1025_d N_A_1162_48#_c_593_n 0.0031664f $X=9.28 $Y=0.37 $X2=0
+ $Y2=0
cc_381 N_A_864_48#_c_411_n N_A_1162_48#_c_593_n 0.0147399f $X=9.42 $Y=0.835
+ $X2=0 $Y2=0
cc_382 N_A_864_48#_c_411_n N_A_1162_48#_c_595_n 0.0348053f $X=9.42 $Y=0.835
+ $X2=0 $Y2=0
cc_383 N_A_864_48#_c_409_n N_A_1162_48#_c_597_n 0.0084327f $X=9.26 $Y=1.275
+ $X2=0 $Y2=0
cc_384 N_A_864_48#_c_411_n N_A_1162_48#_c_597_n 0.00702742f $X=9.42 $Y=0.835
+ $X2=0 $Y2=0
cc_385 N_A_864_48#_c_424_n N_A_1162_48#_c_610_n 0.00214236f $X=9.3 $Y=2.115
+ $X2=0 $Y2=0
cc_386 N_A_864_48#_c_424_n N_C_N_c_775_n 0.0126899f $X=9.3 $Y=2.115 $X2=-0.19
+ $Y2=-0.245
cc_387 N_A_864_48#_c_425_n N_C_N_c_775_n 8.94338e-19 $X=9.41 $Y=2.265 $X2=-0.19
+ $Y2=-0.245
cc_388 N_A_864_48#_c_407_n N_C_N_M1025_g 0.00108093f $X=8.71 $Y=1.385 $X2=0
+ $Y2=0
cc_389 N_A_864_48#_c_408_n N_C_N_M1025_g 0.0167074f $X=8.71 $Y=1.385 $X2=0 $Y2=0
cc_390 N_A_864_48#_c_409_n N_C_N_M1025_g 0.0157095f $X=9.26 $Y=1.275 $X2=0 $Y2=0
cc_391 N_A_864_48#_c_411_n N_C_N_M1025_g 0.0143653f $X=9.42 $Y=0.835 $X2=0 $Y2=0
cc_392 N_A_864_48#_c_424_n N_C_N_c_776_n 0.00289837f $X=9.3 $Y=2.115 $X2=0 $Y2=0
cc_393 N_A_864_48#_c_425_n N_C_N_c_776_n 0.00988129f $X=9.41 $Y=2.265 $X2=0
+ $Y2=0
cc_394 N_A_864_48#_c_407_n C_N 0.0132892f $X=8.71 $Y=1.385 $X2=0 $Y2=0
cc_395 N_A_864_48#_c_409_n C_N 0.0398912f $X=9.26 $Y=1.275 $X2=0 $Y2=0
cc_396 N_A_864_48#_c_424_n C_N 0.0377554f $X=9.3 $Y=2.115 $X2=0 $Y2=0
cc_397 N_A_864_48#_c_426_n C_N 0.00983292f $X=8.71 $Y=1.81 $X2=0 $Y2=0
cc_398 N_A_864_48#_c_407_n N_C_N_c_774_n 0.00126063f $X=8.71 $Y=1.385 $X2=0
+ $Y2=0
cc_399 N_A_864_48#_c_408_n N_C_N_c_774_n 0.00121877f $X=8.71 $Y=1.385 $X2=0
+ $Y2=0
cc_400 N_A_864_48#_c_409_n N_C_N_c_774_n 0.00542909f $X=9.26 $Y=1.275 $X2=0
+ $Y2=0
cc_401 N_A_864_48#_c_424_n N_C_N_c_774_n 0.0069495f $X=9.3 $Y=2.115 $X2=0 $Y2=0
cc_402 N_A_864_48#_c_426_n N_C_N_c_774_n 0.0069332f $X=8.71 $Y=1.81 $X2=0 $Y2=0
cc_403 N_A_864_48#_c_424_n N_D_N_c_824_n 2.32272e-19 $X=9.3 $Y=2.115 $X2=0 $Y2=0
cc_404 N_A_864_48#_c_420_n N_A_27_368#_M1013_d 0.00872108f $X=5.27 $Y=2.225
+ $X2=0 $Y2=0
cc_405 N_A_864_48#_c_489_p N_A_27_368#_M1013_d 0.00433073f $X=5.355 $Y=2.31
+ $X2=0 $Y2=0
cc_406 N_A_864_48#_c_421_n N_A_27_368#_M1037_d 0.00420989f $X=8.545 $Y=1.81
+ $X2=0 $Y2=0
cc_407 N_A_864_48#_c_414_n N_A_27_368#_c_864_n 0.00612425f $X=4.41 $Y=1.67 $X2=0
+ $Y2=0
cc_408 N_A_864_48#_c_414_n N_A_27_368#_c_865_n 0.0118236f $X=4.41 $Y=1.67 $X2=0
+ $Y2=0
cc_409 N_A_864_48#_c_415_n N_A_27_368#_c_865_n 0.00831966f $X=4.86 $Y=1.67 $X2=0
+ $Y2=0
cc_410 N_A_864_48#_c_402_n N_A_27_368#_c_865_n 0.00832028f $X=5.48 $Y=1.67 $X2=0
+ $Y2=0
cc_411 N_A_864_48#_c_417_n N_A_27_368#_c_865_n 0.0134012f $X=8.095 $Y=1.67 $X2=0
+ $Y2=0
cc_412 N_A_864_48#_c_417_n N_A_27_368#_c_867_n 0.00360154f $X=8.095 $Y=1.67
+ $X2=0 $Y2=0
cc_413 N_A_864_48#_c_421_n N_A_27_368#_c_867_n 0.0213159f $X=8.545 $Y=1.81 $X2=0
+ $Y2=0
cc_414 N_A_864_48#_c_426_n N_A_27_368#_c_867_n 0.00980595f $X=8.71 $Y=1.81 $X2=0
+ $Y2=0
cc_415 N_A_864_48#_c_424_n N_VPWR_M1000_s 0.00205208f $X=9.3 $Y=2.115 $X2=0
+ $Y2=0
cc_416 N_A_864_48#_c_426_n N_VPWR_M1000_s 0.00258952f $X=8.71 $Y=1.81 $X2=0
+ $Y2=0
cc_417 N_A_864_48#_c_417_n N_VPWR_c_1013_n 0.00138416f $X=8.095 $Y=1.67 $X2=0
+ $Y2=0
cc_418 N_A_864_48#_c_424_n N_VPWR_c_1013_n 0.0150888f $X=9.3 $Y=2.115 $X2=0
+ $Y2=0
cc_419 N_A_864_48#_c_425_n N_VPWR_c_1013_n 0.0226017f $X=9.41 $Y=2.265 $X2=0
+ $Y2=0
cc_420 N_A_864_48#_c_426_n N_VPWR_c_1013_n 0.00757359f $X=8.71 $Y=1.81 $X2=0
+ $Y2=0
cc_421 N_A_864_48#_c_425_n N_VPWR_c_1014_n 0.0121397f $X=9.41 $Y=2.265 $X2=0
+ $Y2=0
cc_422 N_A_864_48#_c_424_n N_VPWR_c_1015_n 0.00695425f $X=9.3 $Y=2.115 $X2=0
+ $Y2=0
cc_423 N_A_864_48#_c_425_n N_VPWR_c_1015_n 0.0500942f $X=9.41 $Y=2.265 $X2=0
+ $Y2=0
cc_424 N_A_864_48#_c_414_n N_VPWR_c_1020_n 7.74126e-19 $X=4.41 $Y=1.67 $X2=0
+ $Y2=0
cc_425 N_A_864_48#_c_415_n N_VPWR_c_1020_n 7.74126e-19 $X=4.86 $Y=1.67 $X2=0
+ $Y2=0
cc_426 N_A_864_48#_c_402_n N_VPWR_c_1020_n 7.74126e-19 $X=5.48 $Y=1.67 $X2=0
+ $Y2=0
cc_427 N_A_864_48#_c_417_n N_VPWR_c_1020_n 7.74126e-19 $X=8.095 $Y=1.67 $X2=0
+ $Y2=0
cc_428 N_A_864_48#_c_425_n N_VPWR_c_1010_n 0.0100153f $X=9.41 $Y=2.265 $X2=0
+ $Y2=0
cc_429 N_A_864_48#_c_438_p N_A_897_349#_M1032_s 0.00907897f $X=7.4 $Y=2.31 $X2=0
+ $Y2=0
cc_430 N_A_864_48#_c_438_p N_A_897_349#_M1006_s 0.00417719f $X=7.4 $Y=2.31 $X2=0
+ $Y2=0
cc_431 N_A_864_48#_c_438_p N_A_897_349#_M1019_s 0.00359897f $X=7.4 $Y=2.31 $X2=0
+ $Y2=0
cc_432 N_A_864_48#_c_516_p N_A_897_349#_M1019_s 0.00549419f $X=7.485 $Y=2.225
+ $X2=0 $Y2=0
cc_433 N_A_864_48#_c_421_n N_A_897_349#_M1019_s 0.00835454f $X=8.545 $Y=1.81
+ $X2=0 $Y2=0
cc_434 N_A_864_48#_c_422_n N_A_897_349#_M1019_s 0.00122878f $X=7.57 $Y=1.81
+ $X2=0 $Y2=0
cc_435 N_A_864_48#_c_414_n N_A_897_349#_c_1125_n 0.00197554f $X=4.41 $Y=1.67
+ $X2=0 $Y2=0
cc_436 N_A_864_48#_c_415_n N_A_897_349#_c_1125_n 4.23958e-19 $X=4.86 $Y=1.67
+ $X2=0 $Y2=0
cc_437 N_A_864_48#_c_414_n N_A_897_349#_c_1127_n 0.00857957f $X=4.41 $Y=1.67
+ $X2=0 $Y2=0
cc_438 N_A_864_48#_c_415_n N_A_897_349#_c_1127_n 0.0130166f $X=4.86 $Y=1.67
+ $X2=0 $Y2=0
cc_439 N_A_864_48#_c_402_n N_A_897_349#_c_1127_n 0.00105625f $X=5.48 $Y=1.67
+ $X2=0 $Y2=0
cc_440 N_A_864_48#_c_430_n N_A_897_349#_c_1127_n 0.0218087f $X=5.185 $Y=1.42
+ $X2=0 $Y2=0
cc_441 N_A_864_48#_c_420_n N_A_897_349#_c_1127_n 0.018465f $X=5.27 $Y=2.225
+ $X2=0 $Y2=0
cc_442 N_A_864_48#_c_489_p N_A_897_349#_c_1127_n 0.00748036f $X=5.355 $Y=2.31
+ $X2=0 $Y2=0
cc_443 N_A_864_48#_c_412_n N_A_897_349#_c_1127_n 0.00642829f $X=4.97 $Y=1.42
+ $X2=0 $Y2=0
cc_444 N_A_864_48#_c_415_n N_A_897_349#_c_1134_n 0.0127765f $X=4.86 $Y=1.67
+ $X2=0 $Y2=0
cc_445 N_A_864_48#_c_402_n N_A_897_349#_c_1134_n 0.00932878f $X=5.48 $Y=1.67
+ $X2=0 $Y2=0
cc_446 N_A_864_48#_c_438_p N_A_897_349#_c_1134_n 0.117458f $X=7.4 $Y=2.31 $X2=0
+ $Y2=0
cc_447 N_A_864_48#_c_489_p N_A_897_349#_c_1134_n 0.0132166f $X=5.355 $Y=2.31
+ $X2=0 $Y2=0
cc_448 N_A_864_48#_c_421_n N_A_897_349#_c_1134_n 0.004886f $X=8.545 $Y=1.81
+ $X2=0 $Y2=0
cc_449 N_A_864_48#_c_417_n N_A_897_349#_c_1139_n 0.00188661f $X=8.095 $Y=1.67
+ $X2=0 $Y2=0
cc_450 N_A_864_48#_c_417_n N_A_897_349#_c_1140_n 0.00563621f $X=8.095 $Y=1.67
+ $X2=0 $Y2=0
cc_451 N_A_864_48#_c_438_p N_A_897_349#_c_1140_n 0.0131549f $X=7.4 $Y=2.31 $X2=0
+ $Y2=0
cc_452 N_A_864_48#_c_516_p N_A_897_349#_c_1140_n 0.0110665f $X=7.485 $Y=2.225
+ $X2=0 $Y2=0
cc_453 N_A_864_48#_c_421_n N_A_897_349#_c_1140_n 0.0174376f $X=8.545 $Y=1.81
+ $X2=0 $Y2=0
cc_454 N_A_864_48#_c_438_p N_Y_M1002_d 0.00395925f $X=7.4 $Y=2.31 $X2=0 $Y2=0
cc_455 N_A_864_48#_c_438_p N_Y_M1016_d 0.00382413f $X=7.4 $Y=2.31 $X2=0 $Y2=0
cc_456 N_A_864_48#_M1009_g N_Y_c_1187_n 0.0152126f $X=4.395 $Y=0.74 $X2=0 $Y2=0
cc_457 N_A_864_48#_c_430_n N_Y_c_1187_n 0.0106151f $X=5.185 $Y=1.42 $X2=0 $Y2=0
cc_458 N_A_864_48#_M1009_g N_Y_c_1164_n 0.00300817f $X=4.395 $Y=0.74 $X2=0 $Y2=0
cc_459 N_A_864_48#_M1014_g N_Y_c_1164_n 0.00794599f $X=4.895 $Y=0.74 $X2=0 $Y2=0
cc_460 N_A_864_48#_M1035_g N_Y_c_1164_n 8.40071e-19 $X=5.395 $Y=0.74 $X2=0 $Y2=0
cc_461 N_A_864_48#_M1014_g N_Y_c_1222_n 0.0113806f $X=4.895 $Y=0.74 $X2=0 $Y2=0
cc_462 N_A_864_48#_M1035_g N_Y_c_1222_n 0.0158551f $X=5.395 $Y=0.74 $X2=0 $Y2=0
cc_463 N_A_864_48#_c_404_n N_Y_c_1222_n 0.0031198f $X=5.32 $Y=1.42 $X2=0 $Y2=0
cc_464 N_A_864_48#_c_430_n N_Y_c_1222_n 0.0226228f $X=5.185 $Y=1.42 $X2=0 $Y2=0
cc_465 N_A_864_48#_c_406_n N_Y_c_1222_n 0.0111559f $X=5.27 $Y=1.585 $X2=0 $Y2=0
cc_466 N_A_864_48#_M1035_g N_Y_c_1165_n 4.59389e-19 $X=5.395 $Y=0.74 $X2=0 $Y2=0
cc_467 N_A_864_48#_M1035_g N_Y_c_1166_n 0.00381103f $X=5.395 $Y=0.74 $X2=0 $Y2=0
cc_468 N_A_864_48#_c_402_n N_Y_c_1166_n 0.00223065f $X=5.48 $Y=1.67 $X2=0 $Y2=0
cc_469 N_A_864_48#_c_406_n N_Y_c_1166_n 0.00348532f $X=5.27 $Y=1.585 $X2=0 $Y2=0
cc_470 N_A_864_48#_c_402_n N_Y_c_1168_n 0.00721851f $X=5.48 $Y=1.67 $X2=0 $Y2=0
cc_471 N_A_864_48#_c_406_n N_Y_c_1168_n 0.0143906f $X=5.27 $Y=1.585 $X2=0 $Y2=0
cc_472 N_A_864_48#_c_402_n N_Y_c_1169_n 0.00184597f $X=5.48 $Y=1.67 $X2=0 $Y2=0
cc_473 N_A_864_48#_c_406_n N_Y_c_1169_n 0.00304405f $X=5.27 $Y=1.585 $X2=0 $Y2=0
cc_474 N_A_864_48#_c_420_n N_Y_c_1169_n 0.00868733f $X=5.27 $Y=2.225 $X2=0 $Y2=0
cc_475 N_A_864_48#_c_438_p N_Y_c_1169_n 0.0170404f $X=7.4 $Y=2.31 $X2=0 $Y2=0
cc_476 N_A_864_48#_c_438_p N_Y_c_1174_n 0.0505044f $X=7.4 $Y=2.31 $X2=0 $Y2=0
cc_477 N_A_864_48#_c_422_n N_Y_c_1174_n 0.00799568f $X=7.57 $Y=1.81 $X2=0 $Y2=0
cc_478 N_A_864_48#_M1014_g N_Y_c_1239_n 7.32094e-19 $X=4.895 $Y=0.74 $X2=0 $Y2=0
cc_479 N_A_864_48#_c_430_n N_Y_c_1239_n 0.024044f $X=5.185 $Y=1.42 $X2=0 $Y2=0
cc_480 N_A_864_48#_c_412_n N_Y_c_1239_n 0.00396026f $X=4.97 $Y=1.42 $X2=0 $Y2=0
cc_481 N_A_864_48#_M1009_g N_VGND_c_1350_n 0.00873943f $X=4.395 $Y=0.74 $X2=0
+ $Y2=0
cc_482 N_A_864_48#_M1014_g N_VGND_c_1350_n 4.55829e-19 $X=4.895 $Y=0.74 $X2=0
+ $Y2=0
cc_483 N_A_864_48#_M1009_g N_VGND_c_1351_n 0.00383152f $X=4.395 $Y=0.74 $X2=0
+ $Y2=0
cc_484 N_A_864_48#_M1014_g N_VGND_c_1351_n 0.00434272f $X=4.895 $Y=0.74 $X2=0
+ $Y2=0
cc_485 N_A_864_48#_M1014_g N_VGND_c_1352_n 0.00383319f $X=4.895 $Y=0.74 $X2=0
+ $Y2=0
cc_486 N_A_864_48#_M1035_g N_VGND_c_1352_n 0.00875509f $X=5.395 $Y=0.74 $X2=0
+ $Y2=0
cc_487 N_A_864_48#_M1035_g N_VGND_c_1353_n 0.00383152f $X=5.395 $Y=0.74 $X2=0
+ $Y2=0
cc_488 N_A_864_48#_M1035_g N_VGND_c_1354_n 4.65366e-19 $X=5.395 $Y=0.74 $X2=0
+ $Y2=0
cc_489 N_A_864_48#_c_403_n N_VGND_c_1357_n 0.00399234f $X=8.11 $Y=1.22 $X2=0
+ $Y2=0
cc_490 N_A_864_48#_c_413_n N_VGND_c_1357_n 8.39687e-19 $X=8.545 $Y=1.385 $X2=0
+ $Y2=0
cc_491 N_A_864_48#_c_403_n N_VGND_c_1360_n 0.00461464f $X=8.11 $Y=1.22 $X2=0
+ $Y2=0
cc_492 N_A_864_48#_M1009_g N_VGND_c_1363_n 0.00758198f $X=4.395 $Y=0.74 $X2=0
+ $Y2=0
cc_493 N_A_864_48#_M1014_g N_VGND_c_1363_n 0.00821377f $X=4.895 $Y=0.74 $X2=0
+ $Y2=0
cc_494 N_A_864_48#_M1035_g N_VGND_c_1363_n 0.00758168f $X=5.395 $Y=0.74 $X2=0
+ $Y2=0
cc_495 N_A_864_48#_c_403_n N_VGND_c_1363_n 0.00912873f $X=8.11 $Y=1.22 $X2=0
+ $Y2=0
cc_496 N_A_1162_48#_c_593_n N_C_N_M1025_g 0.0163041f $X=9.755 $Y=0.34 $X2=0
+ $Y2=0
cc_497 N_A_1162_48#_c_595_n N_C_N_M1025_g 0.00439827f $X=9.84 $Y=1.11 $X2=0
+ $Y2=0
cc_498 N_A_1162_48#_c_597_n N_C_N_M1025_g 7.16704e-19 $X=9.925 $Y=1.195 $X2=0
+ $Y2=0
cc_499 N_A_1162_48#_c_596_n C_N 0.00178939f $X=10.665 $Y=1.195 $X2=0 $Y2=0
cc_500 N_A_1162_48#_c_597_n C_N 0.0114792f $X=9.925 $Y=1.195 $X2=0 $Y2=0
cc_501 N_A_1162_48#_c_610_n N_C_N_c_774_n 4.18443e-19 $X=10.395 $Y=2.035 $X2=0
+ $Y2=0
cc_502 N_A_1162_48#_c_610_n N_D_N_c_823_n 4.33562e-19 $X=10.395 $Y=2.035 $X2=0
+ $Y2=0
cc_503 N_A_1162_48#_c_608_n N_D_N_c_824_n 0.0106101f $X=10.31 $Y=2.265 $X2=0
+ $Y2=0
cc_504 N_A_1162_48#_c_610_n N_D_N_c_824_n 0.00534188f $X=10.395 $Y=2.035 $X2=0
+ $Y2=0
cc_505 N_A_1162_48#_c_609_n N_D_N_c_825_n 0.00497176f $X=10.755 $Y=2.035 $X2=0
+ $Y2=0
cc_506 N_A_1162_48#_c_608_n N_D_N_c_826_n 0.0067581f $X=10.31 $Y=2.265 $X2=0
+ $Y2=0
cc_507 N_A_1162_48#_c_609_n N_D_N_c_826_n 0.0144943f $X=10.755 $Y=2.035 $X2=0
+ $Y2=0
cc_508 N_A_1162_48#_c_593_n N_D_N_M1008_g 5.08672e-19 $X=9.755 $Y=0.34 $X2=0
+ $Y2=0
cc_509 N_A_1162_48#_c_595_n N_D_N_M1008_g 0.00266659f $X=9.84 $Y=1.11 $X2=0
+ $Y2=0
cc_510 N_A_1162_48#_c_596_n N_D_N_M1008_g 0.0199401f $X=10.665 $Y=1.195 $X2=0
+ $Y2=0
cc_511 N_A_1162_48#_c_598_n N_D_N_M1008_g 0.00160885f $X=10.76 $Y=0.515 $X2=0
+ $Y2=0
cc_512 N_A_1162_48#_c_599_n N_D_N_M1008_g 0.0110911f $X=10.84 $Y=1.95 $X2=0
+ $Y2=0
cc_513 N_A_1162_48#_c_596_n D_N 0.0247729f $X=10.665 $Y=1.195 $X2=0 $Y2=0
cc_514 N_A_1162_48#_c_609_n D_N 0.00438543f $X=10.755 $Y=2.035 $X2=0 $Y2=0
cc_515 N_A_1162_48#_c_610_n D_N 0.0210537f $X=10.395 $Y=2.035 $X2=0 $Y2=0
cc_516 N_A_1162_48#_c_599_n D_N 0.0162242f $X=10.84 $Y=1.95 $X2=0 $Y2=0
cc_517 N_A_1162_48#_c_596_n N_D_N_c_822_n 0.00832055f $X=10.665 $Y=1.195 $X2=0
+ $Y2=0
cc_518 N_A_1162_48#_c_610_n N_D_N_c_822_n 7.12326e-19 $X=10.395 $Y=2.035 $X2=0
+ $Y2=0
cc_519 N_A_1162_48#_c_599_n N_D_N_c_822_n 0.010436f $X=10.84 $Y=1.95 $X2=0 $Y2=0
cc_520 N_A_1162_48#_c_602_n N_A_27_368#_c_865_n 0.00789801f $X=5.93 $Y=1.67
+ $X2=0 $Y2=0
cc_521 N_A_1162_48#_c_604_n N_A_27_368#_c_865_n 0.0079556f $X=6.38 $Y=1.67 $X2=0
+ $Y2=0
cc_522 N_A_1162_48#_c_605_n N_A_27_368#_c_865_n 0.0079556f $X=6.84 $Y=1.67 $X2=0
+ $Y2=0
cc_523 N_A_1162_48#_c_606_n N_A_27_368#_c_865_n 0.00858719f $X=7.29 $Y=1.67
+ $X2=0 $Y2=0
cc_524 N_A_1162_48#_c_609_n N_VPWR_M1029_s 0.00165994f $X=10.755 $Y=2.035 $X2=0
+ $Y2=0
cc_525 N_A_1162_48#_c_608_n N_VPWR_c_1015_n 0.0548333f $X=10.31 $Y=2.265 $X2=0
+ $Y2=0
cc_526 N_A_1162_48#_c_610_n N_VPWR_c_1015_n 0.00141269f $X=10.395 $Y=2.035 $X2=0
+ $Y2=0
cc_527 N_A_1162_48#_c_608_n N_VPWR_c_1017_n 0.0462948f $X=10.31 $Y=2.265 $X2=0
+ $Y2=0
cc_528 N_A_1162_48#_c_609_n N_VPWR_c_1017_n 0.0257228f $X=10.755 $Y=2.035 $X2=0
+ $Y2=0
cc_529 N_A_1162_48#_c_602_n N_VPWR_c_1020_n 7.74126e-19 $X=5.93 $Y=1.67 $X2=0
+ $Y2=0
cc_530 N_A_1162_48#_c_604_n N_VPWR_c_1020_n 7.74126e-19 $X=6.38 $Y=1.67 $X2=0
+ $Y2=0
cc_531 N_A_1162_48#_c_605_n N_VPWR_c_1020_n 7.74126e-19 $X=6.84 $Y=1.67 $X2=0
+ $Y2=0
cc_532 N_A_1162_48#_c_606_n N_VPWR_c_1020_n 7.74126e-19 $X=7.29 $Y=1.67 $X2=0
+ $Y2=0
cc_533 N_A_1162_48#_c_608_n N_VPWR_c_1021_n 0.0110241f $X=10.31 $Y=2.265 $X2=0
+ $Y2=0
cc_534 N_A_1162_48#_c_608_n N_VPWR_c_1010_n 0.00909194f $X=10.31 $Y=2.265 $X2=0
+ $Y2=0
cc_535 N_A_1162_48#_c_602_n N_A_897_349#_c_1134_n 0.008518f $X=5.93 $Y=1.67
+ $X2=0 $Y2=0
cc_536 N_A_1162_48#_c_604_n N_A_897_349#_c_1134_n 0.008518f $X=6.38 $Y=1.67
+ $X2=0 $Y2=0
cc_537 N_A_1162_48#_c_605_n N_A_897_349#_c_1134_n 0.00853169f $X=6.84 $Y=1.67
+ $X2=0 $Y2=0
cc_538 N_A_1162_48#_c_606_n N_A_897_349#_c_1134_n 0.00853169f $X=7.29 $Y=1.67
+ $X2=0 $Y2=0
cc_539 N_A_1162_48#_c_606_n N_A_897_349#_c_1140_n 0.0036122f $X=7.29 $Y=1.67
+ $X2=0 $Y2=0
cc_540 N_A_1162_48#_M1004_g N_Y_c_1165_n 0.0029934f $X=5.885 $Y=0.74 $X2=0 $Y2=0
cc_541 N_A_1162_48#_M1004_g N_Y_c_1166_n 0.00287639f $X=5.885 $Y=0.74 $X2=0
+ $Y2=0
cc_542 N_A_1162_48#_c_581_n N_Y_c_1167_n 0.00811005f $X=5.93 $Y=1.58 $X2=0 $Y2=0
cc_543 N_A_1162_48#_c_588_n N_Y_c_1167_n 0.00990124f $X=5.915 $Y=1.33 $X2=0
+ $Y2=0
cc_544 N_A_1162_48#_c_581_n N_Y_c_1169_n 0.00355452f $X=5.93 $Y=1.58 $X2=0 $Y2=0
cc_545 N_A_1162_48#_c_602_n N_Y_c_1169_n 0.0113893f $X=5.93 $Y=1.67 $X2=0 $Y2=0
cc_546 N_A_1162_48#_c_582_n N_Y_c_1169_n 7.49892e-19 $X=6.29 $Y=1.33 $X2=0 $Y2=0
cc_547 N_A_1162_48#_c_583_n N_Y_c_1169_n 0.00329097f $X=6.38 $Y=1.58 $X2=0 $Y2=0
cc_548 N_A_1162_48#_c_604_n N_Y_c_1169_n 0.00559319f $X=6.38 $Y=1.67 $X2=0 $Y2=0
cc_549 N_A_1162_48#_c_605_n N_Y_c_1169_n 2.52756e-19 $X=6.84 $Y=1.67 $X2=0 $Y2=0
cc_550 N_A_1162_48#_c_590_n N_Y_c_1169_n 0.00295342f $X=8.205 $Y=1.39 $X2=0
+ $Y2=0
cc_551 N_A_1162_48#_c_591_n N_Y_c_1169_n 8.52083e-19 $X=7.63 $Y=1.39 $X2=0 $Y2=0
cc_552 N_A_1162_48#_c_604_n N_Y_c_1174_n 0.0128445f $X=6.38 $Y=1.67 $X2=0 $Y2=0
cc_553 N_A_1162_48#_c_585_n N_Y_c_1174_n 0.00126853f $X=6.75 $Y=1.33 $X2=0 $Y2=0
cc_554 N_A_1162_48#_c_605_n N_Y_c_1174_n 0.0135953f $X=6.84 $Y=1.67 $X2=0 $Y2=0
cc_555 N_A_1162_48#_c_606_n N_Y_c_1174_n 0.00391611f $X=7.29 $Y=1.67 $X2=0 $Y2=0
cc_556 N_A_1162_48#_c_590_n N_Y_c_1174_n 0.034623f $X=8.205 $Y=1.39 $X2=0 $Y2=0
cc_557 N_A_1162_48#_c_591_n N_Y_c_1174_n 0.00782875f $X=7.63 $Y=1.39 $X2=0 $Y2=0
cc_558 N_A_1162_48#_M1005_g N_Y_c_1170_n 0.00592975f $X=6.395 $Y=0.74 $X2=0
+ $Y2=0
cc_559 N_A_1162_48#_c_586_n N_Y_c_1170_n 0.0128221f $X=6.825 $Y=1.225 $X2=0
+ $Y2=0
cc_560 N_A_1162_48#_M1004_g N_Y_c_1171_n 4.17689e-19 $X=5.885 $Y=0.74 $X2=0
+ $Y2=0
cc_561 N_A_1162_48#_M1005_g N_Y_c_1171_n 0.00448642f $X=6.395 $Y=0.74 $X2=0
+ $Y2=0
cc_562 N_A_1162_48#_c_585_n N_Y_c_1171_n 0.00297174f $X=6.75 $Y=1.33 $X2=0 $Y2=0
cc_563 N_A_1162_48#_c_586_n N_Y_c_1171_n 0.00378048f $X=6.825 $Y=1.225 $X2=0
+ $Y2=0
cc_564 N_A_1162_48#_c_589_n N_Y_c_1171_n 0.00143354f $X=6.38 $Y=1.33 $X2=0 $Y2=0
cc_565 N_A_1162_48#_c_590_n N_Y_c_1171_n 0.00574535f $X=8.205 $Y=1.39 $X2=0
+ $Y2=0
cc_566 N_A_1162_48#_c_586_n N_Y_c_1268_n 0.0126093f $X=6.825 $Y=1.225 $X2=0
+ $Y2=0
cc_567 N_A_1162_48#_c_587_n N_Y_c_1268_n 0.0124766f $X=7.655 $Y=1.225 $X2=0
+ $Y2=0
cc_568 N_A_1162_48#_c_590_n N_Y_c_1268_n 0.0631748f $X=8.205 $Y=1.39 $X2=0 $Y2=0
cc_569 N_A_1162_48#_c_591_n N_Y_c_1268_n 0.0118441f $X=7.63 $Y=1.39 $X2=0 $Y2=0
cc_570 N_A_1162_48#_c_581_n N_Y_c_1172_n 9.83931e-19 $X=5.93 $Y=1.58 $X2=0 $Y2=0
cc_571 N_A_1162_48#_c_582_n N_Y_c_1172_n 0.00678571f $X=6.29 $Y=1.33 $X2=0 $Y2=0
cc_572 N_A_1162_48#_c_583_n N_Y_c_1172_n 0.00462284f $X=6.38 $Y=1.58 $X2=0 $Y2=0
cc_573 N_A_1162_48#_c_585_n N_Y_c_1172_n 0.00420978f $X=6.75 $Y=1.33 $X2=0 $Y2=0
cc_574 N_A_1162_48#_c_588_n N_Y_c_1172_n 7.03201e-19 $X=5.915 $Y=1.33 $X2=0
+ $Y2=0
cc_575 N_A_1162_48#_c_589_n N_Y_c_1172_n 0.00873822f $X=6.38 $Y=1.33 $X2=0 $Y2=0
cc_576 N_A_1162_48#_c_590_n N_Y_c_1172_n 0.0145093f $X=8.205 $Y=1.39 $X2=0 $Y2=0
cc_577 N_A_1162_48#_c_591_n N_Y_c_1172_n 5.3629e-19 $X=7.63 $Y=1.39 $X2=0 $Y2=0
cc_578 N_A_1162_48#_M1005_g N_Y_c_1280_n 0.00174725f $X=6.395 $Y=0.74 $X2=0
+ $Y2=0
cc_579 N_A_1162_48#_c_585_n N_Y_c_1280_n 0.00115804f $X=6.75 $Y=1.33 $X2=0 $Y2=0
cc_580 N_A_1162_48#_c_586_n N_Y_c_1280_n 0.00101451f $X=6.825 $Y=1.225 $X2=0
+ $Y2=0
cc_581 N_A_1162_48#_c_587_n Y 0.0128049f $X=7.655 $Y=1.225 $X2=0 $Y2=0
cc_582 N_A_1162_48#_c_587_n N_Y_c_1284_n 7.18118e-19 $X=7.655 $Y=1.225 $X2=0
+ $Y2=0
cc_583 N_A_1162_48#_c_590_n N_Y_c_1284_n 0.0229387f $X=8.205 $Y=1.39 $X2=0 $Y2=0
cc_584 N_A_1162_48#_c_591_n N_Y_c_1284_n 0.00134042f $X=7.63 $Y=1.39 $X2=0 $Y2=0
cc_585 N_A_1162_48#_c_592_n N_VGND_M1036_d 0.00353466f $X=8.29 $Y=1.225 $X2=0
+ $Y2=0
cc_586 N_A_1162_48#_c_638_n N_VGND_M1036_d 0.0207416f $X=8.92 $Y=0.935 $X2=0
+ $Y2=0
cc_587 N_A_1162_48#_c_739_p N_VGND_M1036_d 0.00270595f $X=8.375 $Y=0.935 $X2=0
+ $Y2=0
cc_588 N_A_1162_48#_c_740_p N_VGND_M1036_d 0.0115019f $X=9.005 $Y=0.85 $X2=0
+ $Y2=0
cc_589 N_A_1162_48#_c_594_n N_VGND_M1036_d 7.01469e-19 $X=9.09 $Y=0.34 $X2=0
+ $Y2=0
cc_590 N_A_1162_48#_M1004_g N_VGND_c_1352_n 4.39057e-19 $X=5.885 $Y=0.74 $X2=0
+ $Y2=0
cc_591 N_A_1162_48#_M1004_g N_VGND_c_1353_n 0.00413917f $X=5.885 $Y=0.74 $X2=0
+ $Y2=0
cc_592 N_A_1162_48#_M1004_g N_VGND_c_1354_n 0.0124606f $X=5.885 $Y=0.74 $X2=0
+ $Y2=0
cc_593 N_A_1162_48#_c_582_n N_VGND_c_1354_n 0.00448541f $X=6.29 $Y=1.33 $X2=0
+ $Y2=0
cc_594 N_A_1162_48#_M1005_g N_VGND_c_1354_n 0.00601529f $X=6.395 $Y=0.74 $X2=0
+ $Y2=0
cc_595 N_A_1162_48#_M1005_g N_VGND_c_1355_n 0.00434272f $X=6.395 $Y=0.74 $X2=0
+ $Y2=0
cc_596 N_A_1162_48#_c_586_n N_VGND_c_1355_n 0.00434272f $X=6.825 $Y=1.225 $X2=0
+ $Y2=0
cc_597 N_A_1162_48#_c_586_n N_VGND_c_1356_n 0.00251551f $X=6.825 $Y=1.225 $X2=0
+ $Y2=0
cc_598 N_A_1162_48#_c_587_n N_VGND_c_1356_n 0.00251551f $X=7.655 $Y=1.225 $X2=0
+ $Y2=0
cc_599 N_A_1162_48#_c_638_n N_VGND_c_1357_n 0.0297517f $X=8.92 $Y=0.935 $X2=0
+ $Y2=0
cc_600 N_A_1162_48#_c_739_p N_VGND_c_1357_n 0.0117442f $X=8.375 $Y=0.935 $X2=0
+ $Y2=0
cc_601 N_A_1162_48#_c_740_p N_VGND_c_1357_n 0.0202451f $X=9.005 $Y=0.85 $X2=0
+ $Y2=0
cc_602 N_A_1162_48#_c_594_n N_VGND_c_1357_n 0.0154073f $X=9.09 $Y=0.34 $X2=0
+ $Y2=0
cc_603 N_A_1162_48#_c_593_n N_VGND_c_1358_n 0.0152482f $X=9.755 $Y=0.34 $X2=0
+ $Y2=0
cc_604 N_A_1162_48#_c_595_n N_VGND_c_1358_n 0.041427f $X=9.84 $Y=1.11 $X2=0
+ $Y2=0
cc_605 N_A_1162_48#_c_596_n N_VGND_c_1358_n 0.0301874f $X=10.665 $Y=1.195 $X2=0
+ $Y2=0
cc_606 N_A_1162_48#_c_598_n N_VGND_c_1358_n 0.023562f $X=10.76 $Y=0.515 $X2=0
+ $Y2=0
cc_607 N_A_1162_48#_c_587_n N_VGND_c_1360_n 0.00434272f $X=7.655 $Y=1.225 $X2=0
+ $Y2=0
cc_608 N_A_1162_48#_c_593_n N_VGND_c_1361_n 0.05453f $X=9.755 $Y=0.34 $X2=0
+ $Y2=0
cc_609 N_A_1162_48#_c_594_n N_VGND_c_1361_n 0.0121867f $X=9.09 $Y=0.34 $X2=0
+ $Y2=0
cc_610 N_A_1162_48#_c_598_n N_VGND_c_1362_n 0.0115122f $X=10.76 $Y=0.515 $X2=0
+ $Y2=0
cc_611 N_A_1162_48#_M1004_g N_VGND_c_1363_n 0.00818158f $X=5.885 $Y=0.74 $X2=0
+ $Y2=0
cc_612 N_A_1162_48#_M1005_g N_VGND_c_1363_n 0.00820805f $X=6.395 $Y=0.74 $X2=0
+ $Y2=0
cc_613 N_A_1162_48#_c_586_n N_VGND_c_1363_n 0.00822865f $X=6.825 $Y=1.225 $X2=0
+ $Y2=0
cc_614 N_A_1162_48#_c_587_n N_VGND_c_1363_n 0.00823191f $X=7.655 $Y=1.225 $X2=0
+ $Y2=0
cc_615 N_A_1162_48#_c_638_n N_VGND_c_1363_n 0.00702258f $X=8.92 $Y=0.935 $X2=0
+ $Y2=0
cc_616 N_A_1162_48#_c_739_p N_VGND_c_1363_n 6.0824e-19 $X=8.375 $Y=0.935 $X2=0
+ $Y2=0
cc_617 N_A_1162_48#_c_593_n N_VGND_c_1363_n 0.0309211f $X=9.755 $Y=0.34 $X2=0
+ $Y2=0
cc_618 N_A_1162_48#_c_594_n N_VGND_c_1363_n 0.00660921f $X=9.09 $Y=0.34 $X2=0
+ $Y2=0
cc_619 N_A_1162_48#_c_598_n N_VGND_c_1363_n 0.0095288f $X=10.76 $Y=0.515 $X2=0
+ $Y2=0
cc_620 N_C_N_c_776_n N_D_N_c_824_n 0.0119213f $X=9.635 $Y=2.045 $X2=0 $Y2=0
cc_621 C_N D_N 0.0209957f $X=9.755 $Y=1.58 $X2=0 $Y2=0
cc_622 N_C_N_M1025_g N_D_N_c_822_n 0.00189327f $X=9.205 $Y=0.74 $X2=0 $Y2=0
cc_623 C_N N_D_N_c_822_n 0.00589106f $X=9.755 $Y=1.58 $X2=0 $Y2=0
cc_624 N_C_N_c_774_n N_D_N_c_822_n 0.0187596f $X=9.26 $Y=1.695 $X2=0 $Y2=0
cc_625 N_C_N_c_775_n N_A_27_368#_c_865_n 6.10827e-19 $X=9.185 $Y=2.045 $X2=0
+ $Y2=0
cc_626 N_C_N_c_775_n N_A_27_368#_c_867_n 0.0031691f $X=9.185 $Y=2.045 $X2=0
+ $Y2=0
cc_627 N_C_N_c_775_n N_VPWR_c_1013_n 0.0106474f $X=9.185 $Y=2.045 $X2=0 $Y2=0
cc_628 N_C_N_c_776_n N_VPWR_c_1013_n 5.79063e-19 $X=9.635 $Y=2.045 $X2=0 $Y2=0
cc_629 N_C_N_c_775_n N_VPWR_c_1014_n 0.00429299f $X=9.185 $Y=2.045 $X2=0 $Y2=0
cc_630 N_C_N_c_776_n N_VPWR_c_1014_n 0.00445602f $X=9.635 $Y=2.045 $X2=0 $Y2=0
cc_631 N_C_N_c_776_n N_VPWR_c_1015_n 0.00505864f $X=9.635 $Y=2.045 $X2=0 $Y2=0
cc_632 C_N N_VPWR_c_1015_n 0.0116692f $X=9.755 $Y=1.58 $X2=0 $Y2=0
cc_633 N_C_N_c_775_n N_VPWR_c_1010_n 0.00847721f $X=9.185 $Y=2.045 $X2=0 $Y2=0
cc_634 N_C_N_c_776_n N_VPWR_c_1010_n 0.00857673f $X=9.635 $Y=2.045 $X2=0 $Y2=0
cc_635 N_C_N_M1025_g N_VGND_c_1357_n 0.00175002f $X=9.205 $Y=0.74 $X2=0 $Y2=0
cc_636 N_C_N_M1025_g N_VGND_c_1361_n 0.00278271f $X=9.205 $Y=0.74 $X2=0 $Y2=0
cc_637 N_C_N_M1025_g N_VGND_c_1363_n 0.00363426f $X=9.205 $Y=0.74 $X2=0 $Y2=0
cc_638 N_D_N_c_824_n N_VPWR_c_1015_n 0.00505454f $X=10.085 $Y=2.045 $X2=0 $Y2=0
cc_639 N_D_N_c_824_n N_VPWR_c_1017_n 6.2661e-19 $X=10.085 $Y=2.045 $X2=0 $Y2=0
cc_640 N_D_N_c_826_n N_VPWR_c_1017_n 0.0127617f $X=10.535 $Y=2.045 $X2=0 $Y2=0
cc_641 N_D_N_c_824_n N_VPWR_c_1021_n 0.00445602f $X=10.085 $Y=2.045 $X2=0 $Y2=0
cc_642 N_D_N_c_826_n N_VPWR_c_1021_n 0.00413917f $X=10.535 $Y=2.045 $X2=0 $Y2=0
cc_643 N_D_N_c_824_n N_VPWR_c_1010_n 0.00857673f $X=10.085 $Y=2.045 $X2=0 $Y2=0
cc_644 N_D_N_c_826_n N_VPWR_c_1010_n 0.00817726f $X=10.535 $Y=2.045 $X2=0 $Y2=0
cc_645 N_D_N_M1008_g N_VGND_c_1358_n 0.0146102f $X=10.545 $Y=0.74 $X2=0 $Y2=0
cc_646 N_D_N_M1008_g N_VGND_c_1362_n 0.00383152f $X=10.545 $Y=0.74 $X2=0 $Y2=0
cc_647 N_D_N_M1008_g N_VGND_c_1363_n 0.00761198f $X=10.545 $Y=0.74 $X2=0 $Y2=0
cc_648 N_A_27_368#_c_870_n N_A_116_368#_M1010_s 0.00624689f $X=3.06 $Y=2.135
+ $X2=-0.19 $Y2=1.66
cc_649 N_A_27_368#_c_870_n N_A_116_368#_M1022_s 0.00385275f $X=3.06 $Y=2.135
+ $X2=0 $Y2=0
cc_650 N_A_27_368#_c_870_n N_A_116_368#_M1033_s 0.00510511f $X=3.06 $Y=2.135
+ $X2=0 $Y2=0
cc_651 N_A_27_368#_c_878_n N_A_116_368#_M1015_s 0.00448384f $X=4.09 $Y=1.84
+ $X2=0 $Y2=0
cc_652 N_A_27_368#_c_870_n N_A_116_368#_c_965_n 0.0368632f $X=3.06 $Y=2.135
+ $X2=0 $Y2=0
cc_653 N_A_27_368#_c_870_n N_A_116_368#_c_970_n 0.0398412f $X=3.06 $Y=2.135
+ $X2=0 $Y2=0
cc_654 N_A_27_368#_c_870_n N_A_116_368#_c_983_n 0.0188865f $X=3.06 $Y=2.135
+ $X2=0 $Y2=0
cc_655 N_A_27_368#_c_876_n N_A_116_368#_c_951_n 0.0206353f $X=3.225 $Y=2.57
+ $X2=0 $Y2=0
cc_656 N_A_27_368#_c_866_n N_A_116_368#_c_951_n 0.0137714f $X=4.26 $Y=2.99 $X2=0
+ $Y2=0
cc_657 N_A_27_368#_c_878_n N_A_116_368#_c_953_n 0.0202249f $X=4.09 $Y=1.84 $X2=0
+ $Y2=0
cc_658 N_A_27_368#_c_864_n N_A_116_368#_c_953_n 0.052749f $X=4.175 $Y=2.72 $X2=0
+ $Y2=0
cc_659 N_A_27_368#_c_863_n N_A_116_368#_c_954_n 0.0165499f $X=0.28 $Y=2.815
+ $X2=0 $Y2=0
cc_660 N_A_27_368#_c_870_n N_A_116_368#_c_954_n 0.0200687f $X=3.06 $Y=2.135
+ $X2=0 $Y2=0
cc_661 N_A_27_368#_c_870_n N_A_116_368#_c_976_n 0.0154051f $X=3.06 $Y=2.135
+ $X2=0 $Y2=0
cc_662 N_A_27_368#_c_870_n N_VPWR_M1021_d 0.00483954f $X=3.06 $Y=2.135 $X2=-0.19
+ $Y2=1.66
cc_663 N_A_27_368#_c_870_n N_VPWR_M1024_d 0.00594772f $X=3.06 $Y=2.135 $X2=0
+ $Y2=0
cc_664 N_A_27_368#_c_865_n N_VPWR_c_1013_n 0.0100323f $X=8.205 $Y=2.99 $X2=0
+ $Y2=0
cc_665 N_A_27_368#_c_867_n N_VPWR_c_1013_n 0.027995f $X=8.325 $Y=2.23 $X2=0
+ $Y2=0
cc_666 N_A_27_368#_c_863_n N_VPWR_c_1018_n 0.0145938f $X=0.28 $Y=2.815 $X2=0
+ $Y2=0
cc_667 N_A_27_368#_c_865_n N_VPWR_c_1020_n 0.274203f $X=8.205 $Y=2.99 $X2=0
+ $Y2=0
cc_668 N_A_27_368#_c_866_n N_VPWR_c_1020_n 0.0121867f $X=4.26 $Y=2.99 $X2=0
+ $Y2=0
cc_669 N_A_27_368#_M1013_d N_VPWR_c_1010_n 0.00281977f $X=4.935 $Y=1.745 $X2=0
+ $Y2=0
cc_670 N_A_27_368#_c_863_n N_VPWR_c_1010_n 0.0120466f $X=0.28 $Y=2.815 $X2=0
+ $Y2=0
cc_671 N_A_27_368#_c_865_n N_VPWR_c_1010_n 0.159396f $X=8.205 $Y=2.99 $X2=0
+ $Y2=0
cc_672 N_A_27_368#_c_866_n N_VPWR_c_1010_n 0.00660921f $X=4.26 $Y=2.99 $X2=0
+ $Y2=0
cc_673 N_A_27_368#_c_864_n N_A_897_349#_c_1125_n 0.0113397f $X=4.175 $Y=2.72
+ $X2=0 $Y2=0
cc_674 N_A_27_368#_c_865_n N_A_897_349#_c_1125_n 0.0207779f $X=8.205 $Y=2.99
+ $X2=0 $Y2=0
cc_675 N_A_27_368#_c_942_p N_A_897_349#_c_1127_n 0.011926f $X=4.175 $Y=1.925
+ $X2=0 $Y2=0
cc_676 N_A_27_368#_c_864_n N_A_897_349#_c_1127_n 0.0400918f $X=4.175 $Y=2.72
+ $X2=0 $Y2=0
cc_677 N_A_27_368#_M1013_d N_A_897_349#_c_1134_n 0.0137248f $X=4.935 $Y=1.745
+ $X2=0 $Y2=0
cc_678 N_A_27_368#_c_865_n N_A_897_349#_c_1134_n 0.180357f $X=8.205 $Y=2.99
+ $X2=0 $Y2=0
cc_679 N_A_27_368#_c_865_n N_A_897_349#_c_1139_n 0.0188891f $X=8.205 $Y=2.99
+ $X2=0 $Y2=0
cc_680 N_A_27_368#_c_878_n N_Y_c_1187_n 0.00250275f $X=4.09 $Y=1.84 $X2=0 $Y2=0
cc_681 N_A_27_368#_c_942_p N_Y_c_1187_n 0.00481666f $X=4.175 $Y=1.925 $X2=0
+ $Y2=0
cc_682 N_A_116_368#_c_965_n N_VPWR_M1021_d 0.00495301f $X=1.645 $Y=2.475
+ $X2=-0.19 $Y2=1.66
cc_683 N_A_116_368#_c_970_n N_VPWR_M1024_d 0.00609612f $X=2.635 $Y=2.475 $X2=0
+ $Y2=0
cc_684 N_A_116_368#_c_965_n N_VPWR_c_1011_n 0.0195803f $X=1.645 $Y=2.475 $X2=0
+ $Y2=0
cc_685 N_A_116_368#_c_949_n N_VPWR_c_1011_n 0.0167923f $X=1.73 $Y=2.815 $X2=0
+ $Y2=0
cc_686 N_A_116_368#_c_954_n N_VPWR_c_1011_n 0.0101711f $X=0.78 $Y=2.475 $X2=0
+ $Y2=0
cc_687 N_A_116_368#_c_949_n N_VPWR_c_1012_n 0.00979415f $X=1.73 $Y=2.815 $X2=0
+ $Y2=0
cc_688 N_A_116_368#_c_970_n N_VPWR_c_1012_n 0.0228229f $X=2.635 $Y=2.475 $X2=0
+ $Y2=0
cc_689 N_A_116_368#_c_950_n N_VPWR_c_1012_n 0.0118017f $X=2.76 $Y=2.905 $X2=0
+ $Y2=0
cc_690 N_A_116_368#_c_952_n N_VPWR_c_1012_n 0.0126878f $X=2.885 $Y=2.99 $X2=0
+ $Y2=0
cc_691 N_A_116_368#_c_954_n N_VPWR_c_1018_n 0.0144443f $X=0.78 $Y=2.475 $X2=0
+ $Y2=0
cc_692 N_A_116_368#_c_949_n N_VPWR_c_1019_n 0.0109113f $X=1.73 $Y=2.815 $X2=0
+ $Y2=0
cc_693 N_A_116_368#_c_951_n N_VPWR_c_1020_n 0.0670515f $X=3.56 $Y=2.99 $X2=0
+ $Y2=0
cc_694 N_A_116_368#_c_952_n N_VPWR_c_1020_n 0.0179317f $X=2.885 $Y=2.99 $X2=0
+ $Y2=0
cc_695 N_A_116_368#_c_965_n N_VPWR_c_1010_n 0.0128064f $X=1.645 $Y=2.475 $X2=0
+ $Y2=0
cc_696 N_A_116_368#_c_949_n N_VPWR_c_1010_n 0.0090481f $X=1.73 $Y=2.815 $X2=0
+ $Y2=0
cc_697 N_A_116_368#_c_970_n N_VPWR_c_1010_n 0.0129506f $X=2.635 $Y=2.475 $X2=0
+ $Y2=0
cc_698 N_A_116_368#_c_951_n N_VPWR_c_1010_n 0.0381961f $X=3.56 $Y=2.99 $X2=0
+ $Y2=0
cc_699 N_A_116_368#_c_952_n N_VPWR_c_1010_n 0.0097213f $X=2.885 $Y=2.99 $X2=0
+ $Y2=0
cc_700 N_A_116_368#_c_954_n N_VPWR_c_1010_n 0.0119886f $X=0.78 $Y=2.475 $X2=0
+ $Y2=0
cc_701 N_A_897_349#_c_1134_n N_Y_M1002_d 0.0038712f $X=7.76 $Y=2.65 $X2=4.395
+ $Y2=0.74
cc_702 N_A_897_349#_c_1134_n N_Y_M1016_d 0.0038712f $X=7.76 $Y=2.65 $X2=0 $Y2=0
cc_703 N_A_897_349#_M1006_s N_Y_c_1174_n 0.00213169f $X=6.455 $Y=1.745 $X2=8.71
+ $Y2=2.115
cc_704 N_Y_c_1176_n N_VGND_M1011_d 0.00675773f $X=1.615 $Y=0.925 $X2=0 $Y2=0
cc_705 N_Y_c_1207_n N_VGND_M1023_d 0.00565919f $X=2.665 $Y=0.925 $X2=0 $Y2=0
cc_706 N_Y_c_1181_n N_VGND_M1020_s 0.00425479f $X=3.595 $Y=1 $X2=0 $Y2=0
cc_707 N_Y_c_1187_n N_VGND_M1034_s 0.00520194f $X=4.515 $Y=1 $X2=0 $Y2=0
cc_708 N_Y_c_1222_n N_VGND_M1014_d 0.0046331f $X=5.525 $Y=1 $X2=0 $Y2=0
cc_709 N_Y_c_1268_n N_VGND_M1018_d 0.0142442f $X=7.705 $Y=0.97 $X2=0 $Y2=0
cc_710 N_Y_c_1159_n N_VGND_c_1343_n 0.0191389f $X=0.78 $Y=0.515 $X2=0 $Y2=0
cc_711 N_Y_c_1160_n N_VGND_c_1343_n 0.0124832f $X=0.945 $Y=0.925 $X2=0 $Y2=0
cc_712 N_Y_c_1159_n N_VGND_c_1344_n 0.0127977f $X=0.78 $Y=0.515 $X2=0 $Y2=0
cc_713 N_Y_c_1176_n N_VGND_c_1344_n 0.0207693f $X=1.615 $Y=0.925 $X2=0 $Y2=0
cc_714 N_Y_c_1161_n N_VGND_c_1344_n 0.0140622f $X=1.78 $Y=0.515 $X2=0 $Y2=0
cc_715 N_Y_c_1161_n N_VGND_c_1345_n 0.0145323f $X=1.78 $Y=0.515 $X2=0 $Y2=0
cc_716 N_Y_c_1161_n N_VGND_c_1346_n 0.0127977f $X=1.78 $Y=0.515 $X2=0 $Y2=0
cc_717 N_Y_c_1207_n N_VGND_c_1346_n 0.021963f $X=2.665 $Y=0.925 $X2=0 $Y2=0
cc_718 N_Y_c_1162_n N_VGND_c_1346_n 0.00129215f $X=2.75 $Y=0.515 $X2=0 $Y2=0
cc_719 N_Y_c_1162_n N_VGND_c_1347_n 0.011054f $X=2.75 $Y=0.515 $X2=0 $Y2=0
cc_720 N_Y_c_1162_n N_VGND_c_1348_n 0.0149945f $X=2.75 $Y=0.515 $X2=0 $Y2=0
cc_721 N_Y_c_1181_n N_VGND_c_1348_n 0.0193595f $X=3.595 $Y=1 $X2=0 $Y2=0
cc_722 N_Y_c_1163_n N_VGND_c_1348_n 0.0148853f $X=3.68 $Y=0.515 $X2=0 $Y2=0
cc_723 N_Y_c_1163_n N_VGND_c_1349_n 0.011066f $X=3.68 $Y=0.515 $X2=0 $Y2=0
cc_724 N_Y_c_1163_n N_VGND_c_1350_n 0.0155793f $X=3.68 $Y=0.515 $X2=0 $Y2=0
cc_725 N_Y_c_1187_n N_VGND_c_1350_n 0.0170777f $X=4.515 $Y=1 $X2=0 $Y2=0
cc_726 N_Y_c_1164_n N_VGND_c_1350_n 0.0156118f $X=4.68 $Y=0.515 $X2=0 $Y2=0
cc_727 N_Y_c_1164_n N_VGND_c_1351_n 0.0145639f $X=4.68 $Y=0.515 $X2=0 $Y2=0
cc_728 N_Y_c_1164_n N_VGND_c_1352_n 0.0156118f $X=4.68 $Y=0.515 $X2=0 $Y2=0
cc_729 N_Y_c_1222_n N_VGND_c_1352_n 0.0209867f $X=5.525 $Y=1 $X2=0 $Y2=0
cc_730 N_Y_c_1165_n N_VGND_c_1352_n 0.0148853f $X=5.61 $Y=0.515 $X2=0 $Y2=0
cc_731 N_Y_c_1165_n N_VGND_c_1353_n 0.011066f $X=5.61 $Y=0.515 $X2=0 $Y2=0
cc_732 N_Y_c_1165_n N_VGND_c_1354_n 0.0219581f $X=5.61 $Y=0.515 $X2=0 $Y2=0
cc_733 N_Y_c_1166_n N_VGND_c_1354_n 0.00244646f $X=5.65 $Y=1.3 $X2=0 $Y2=0
cc_734 N_Y_c_1167_n N_VGND_c_1354_n 0.0263348f $X=5.99 $Y=1.385 $X2=0 $Y2=0
cc_735 N_Y_c_1170_n N_VGND_c_1354_n 0.0208274f $X=6.61 $Y=0.515 $X2=0 $Y2=0
cc_736 N_Y_c_1171_n N_VGND_c_1354_n 0.00329837f $X=6.53 $Y=1.3 $X2=0 $Y2=0
cc_737 N_Y_c_1170_n N_VGND_c_1355_n 0.0145106f $X=6.61 $Y=0.515 $X2=0 $Y2=0
cc_738 N_Y_c_1170_n N_VGND_c_1356_n 0.0132454f $X=6.61 $Y=0.515 $X2=0 $Y2=0
cc_739 N_Y_c_1268_n N_VGND_c_1356_n 0.0400561f $X=7.705 $Y=0.97 $X2=0 $Y2=0
cc_740 Y N_VGND_c_1356_n 0.0132454f $X=7.835 $Y=0.47 $X2=0 $Y2=0
cc_741 Y N_VGND_c_1357_n 0.0145404f $X=7.835 $Y=0.47 $X2=0 $Y2=0
cc_742 N_Y_c_1159_n N_VGND_c_1359_n 0.0144922f $X=0.78 $Y=0.515 $X2=0 $Y2=0
cc_743 Y N_VGND_c_1360_n 0.0146023f $X=7.835 $Y=0.47 $X2=0 $Y2=0
cc_744 N_Y_c_1159_n N_VGND_c_1363_n 0.0118826f $X=0.78 $Y=0.515 $X2=0 $Y2=0
cc_745 N_Y_c_1176_n N_VGND_c_1363_n 0.0108249f $X=1.615 $Y=0.925 $X2=0 $Y2=0
cc_746 N_Y_c_1161_n N_VGND_c_1363_n 0.0119861f $X=1.78 $Y=0.515 $X2=0 $Y2=0
cc_747 N_Y_c_1207_n N_VGND_c_1363_n 0.0125718f $X=2.665 $Y=0.925 $X2=0 $Y2=0
cc_748 N_Y_c_1162_n N_VGND_c_1363_n 0.00914017f $X=2.75 $Y=0.515 $X2=0 $Y2=0
cc_749 N_Y_c_1163_n N_VGND_c_1363_n 0.00915947f $X=3.68 $Y=0.515 $X2=0 $Y2=0
cc_750 N_Y_c_1164_n N_VGND_c_1363_n 0.0119984f $X=4.68 $Y=0.515 $X2=0 $Y2=0
cc_751 N_Y_c_1165_n N_VGND_c_1363_n 0.00915947f $X=5.61 $Y=0.515 $X2=0 $Y2=0
cc_752 N_Y_c_1170_n N_VGND_c_1363_n 0.0118899f $X=6.61 $Y=0.515 $X2=0 $Y2=0
cc_753 Y N_VGND_c_1363_n 0.0120134f $X=7.835 $Y=0.47 $X2=0 $Y2=0
