* NGSPICE file created from sky130_fd_sc_hs__or3_2.ext - technology: sky130A

.subckt sky130_fd_sc_hs__or3_2 A B C VGND VNB VPB VPWR X
M1000 VGND a_27_74# X VNB nlowvt w=740000u l=150000u
+  ad=9.725e+11p pd=7.09e+06u as=2.072e+11p ps=2.04e+06u
M1001 a_150_392# C a_27_74# VPB pshort w=1e+06u l=150000u
+  ad=2.7e+11p pd=2.54e+06u as=2.95e+11p ps=2.59e+06u
M1002 X a_27_74# VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=3.36e+11p pd=2.84e+06u as=8.782e+11p ps=6.09e+06u
M1003 VPWR a_27_74# X VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 VPWR A a_234_392# VPB pshort w=1e+06u l=150000u
+  ad=0p pd=0u as=4.2e+11p ps=2.84e+06u
M1005 a_234_392# B a_150_392# VPB pshort w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VGND A a_27_74# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=4.064e+11p ps=3.83e+06u
M1007 X a_27_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_27_74# B VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VGND C a_27_74# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

