* NGSPICE file created from sky130_fd_sc_hs__or2_1.ext - technology: sky130A

.subckt sky130_fd_sc_hs__or2_1 A B VGND VNB VPB VPWR X
M1000 a_152_368# B a_63_368# VPB pshort w=840000u l=150000u
+  ad=2.268e+11p pd=2.22e+06u as=2.478e+11p ps=2.27e+06u
M1001 X a_63_368# VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=3.304e+11p pd=2.83e+06u as=6.692e+11p ps=3.52e+06u
M1002 X a_63_368# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=5.7345e+11p ps=4.42e+06u
M1003 VPWR A a_152_368# VPB pshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 VGND A a_63_368# VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=2.6125e+11p ps=2.05e+06u
M1005 a_63_368# B VGND VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

