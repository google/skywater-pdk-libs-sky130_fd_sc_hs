* File: sky130_fd_sc_hs__a22oi_4.pex.spice
* Created: Thu Aug 27 20:27:28 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HS__A22OI_4%B2 1 3 6 10 12 14 17 19 21 24 26 28 29 30 31
+ 46 47
c83 47 0 1.91457e-19 $X=1.87 $Y=1.557
c84 46 0 1.48228e-20 $X=1.79 $Y=1.515
c85 26 0 9.9816e-20 $X=1.925 $Y=1.765
c86 24 0 8.01953e-20 $X=1.87 $Y=0.74
r87 47 48 7.2038 $w=3.68e-07 $l=5.5e-08 $layer=POLY_cond $X=1.87 $Y=1.557
+ $X2=1.925 $Y2=1.557
r88 45 47 10.4783 $w=3.68e-07 $l=8e-08 $layer=POLY_cond $X=1.79 $Y=1.557
+ $X2=1.87 $Y2=1.557
r89 45 46 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.79
+ $Y=1.515 $X2=1.79 $Y2=1.515
r90 43 45 41.2582 $w=3.68e-07 $l=3.15e-07 $layer=POLY_cond $X=1.475 $Y=1.557
+ $X2=1.79 $Y2=1.557
r91 42 43 4.58424 $w=3.68e-07 $l=3.5e-08 $layer=POLY_cond $X=1.44 $Y=1.557
+ $X2=1.475 $Y2=1.557
r92 41 42 54.356 $w=3.68e-07 $l=4.15e-07 $layer=POLY_cond $X=1.025 $Y=1.557
+ $X2=1.44 $Y2=1.557
r93 40 41 1.96467 $w=3.68e-07 $l=1.5e-08 $layer=POLY_cond $X=1.01 $Y=1.557
+ $X2=1.025 $Y2=1.557
r94 38 40 31.4348 $w=3.68e-07 $l=2.4e-07 $layer=POLY_cond $X=0.77 $Y=1.557
+ $X2=1.01 $Y2=1.557
r95 38 39 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.77
+ $Y=1.515 $X2=0.77 $Y2=1.515
r96 36 38 24.8859 $w=3.68e-07 $l=1.9e-07 $layer=POLY_cond $X=0.58 $Y=1.557
+ $X2=0.77 $Y2=1.557
r97 35 36 0.654891 $w=3.68e-07 $l=5e-09 $layer=POLY_cond $X=0.575 $Y=1.557
+ $X2=0.58 $Y2=1.557
r98 31 46 2.94811 $w=4.28e-07 $l=1.1e-07 $layer=LI1_cond $X=1.68 $Y=1.565
+ $X2=1.79 $Y2=1.565
r99 30 31 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=1.2 $Y=1.565
+ $X2=1.68 $Y2=1.565
r100 30 39 11.5244 $w=4.28e-07 $l=4.3e-07 $layer=LI1_cond $X=1.2 $Y=1.565
+ $X2=0.77 $Y2=1.565
r101 29 39 1.34005 $w=4.28e-07 $l=5e-08 $layer=LI1_cond $X=0.72 $Y=1.565
+ $X2=0.77 $Y2=1.565
r102 26 48 23.8357 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=1.925 $Y=1.765
+ $X2=1.925 $Y2=1.557
r103 26 28 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.925 $Y=1.765
+ $X2=1.925 $Y2=2.4
r104 22 47 23.8357 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.87 $Y=1.35
+ $X2=1.87 $Y2=1.557
r105 22 24 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.87 $Y=1.35
+ $X2=1.87 $Y2=0.74
r106 19 43 23.8357 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=1.475 $Y=1.765
+ $X2=1.475 $Y2=1.557
r107 19 21 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.475 $Y=1.765
+ $X2=1.475 $Y2=2.4
r108 15 42 23.8357 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.44 $Y=1.35
+ $X2=1.44 $Y2=1.557
r109 15 17 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.44 $Y=1.35
+ $X2=1.44 $Y2=0.74
r110 12 41 23.8357 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=1.025 $Y=1.765
+ $X2=1.025 $Y2=1.557
r111 12 14 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.025 $Y=1.765
+ $X2=1.025 $Y2=2.4
r112 8 40 23.8357 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.01 $Y=1.35
+ $X2=1.01 $Y2=1.557
r113 8 10 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.01 $Y=1.35
+ $X2=1.01 $Y2=0.74
r114 4 36 23.8357 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.58 $Y=1.35
+ $X2=0.58 $Y2=1.557
r115 4 6 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=0.58 $Y=1.35 $X2=0.58
+ $Y2=0.74
r116 1 35 23.8357 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=0.575 $Y=1.765
+ $X2=0.575 $Y2=1.557
r117 1 3 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.575 $Y=1.765
+ $X2=0.575 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_HS__A22OI_4%B1 3 5 7 10 12 14 17 19 21 24 26 28 29 30 45
c97 30 0 9.9816e-20 $X=3.12 $Y=1.665
c98 5 0 1.48228e-20 $X=2.375 $Y=1.765
c99 3 0 1.9142e-19 $X=2.3 $Y=0.74
r100 45 46 16.5573 $w=3.93e-07 $l=1.35e-07 $layer=POLY_cond $X=3.59 $Y=1.542
+ $X2=3.725 $Y2=1.542
r101 44 45 38.6336 $w=3.93e-07 $l=3.15e-07 $layer=POLY_cond $X=3.275 $Y=1.542
+ $X2=3.59 $Y2=1.542
r102 43 44 14.1043 $w=3.93e-07 $l=1.15e-07 $layer=POLY_cond $X=3.16 $Y=1.542
+ $X2=3.275 $Y2=1.542
r103 41 43 6.13232 $w=3.93e-07 $l=5e-08 $layer=POLY_cond $X=3.11 $Y=1.542
+ $X2=3.16 $Y2=1.542
r104 41 42 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=3.11
+ $Y=1.515 $X2=3.11 $Y2=1.515
r105 39 41 34.9542 $w=3.93e-07 $l=2.85e-07 $layer=POLY_cond $X=2.825 $Y=1.542
+ $X2=3.11 $Y2=1.542
r106 38 39 11.6514 $w=3.93e-07 $l=9.5e-08 $layer=POLY_cond $X=2.73 $Y=1.542
+ $X2=2.825 $Y2=1.542
r107 36 38 36.7939 $w=3.93e-07 $l=3e-07 $layer=POLY_cond $X=2.43 $Y=1.542
+ $X2=2.73 $Y2=1.542
r108 36 37 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=2.43
+ $Y=1.515 $X2=2.43 $Y2=1.515
r109 34 36 6.74555 $w=3.93e-07 $l=5.5e-08 $layer=POLY_cond $X=2.375 $Y=1.542
+ $X2=2.43 $Y2=1.542
r110 33 34 9.19847 $w=3.93e-07 $l=7.5e-08 $layer=POLY_cond $X=2.3 $Y=1.542
+ $X2=2.375 $Y2=1.542
r111 30 42 0.26801 $w=4.28e-07 $l=1e-08 $layer=LI1_cond $X=3.12 $Y=1.565
+ $X2=3.11 $Y2=1.565
r112 29 42 12.5965 $w=4.28e-07 $l=4.7e-07 $layer=LI1_cond $X=2.64 $Y=1.565
+ $X2=3.11 $Y2=1.565
r113 29 37 5.62821 $w=4.28e-07 $l=2.1e-07 $layer=LI1_cond $X=2.64 $Y=1.565
+ $X2=2.43 $Y2=1.565
r114 26 46 25.4309 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=3.725 $Y=1.765
+ $X2=3.725 $Y2=1.542
r115 26 28 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.725 $Y=1.765
+ $X2=3.725 $Y2=2.4
r116 22 45 25.4309 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=3.59 $Y=1.32
+ $X2=3.59 $Y2=1.542
r117 22 24 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=3.59 $Y=1.32
+ $X2=3.59 $Y2=0.74
r118 19 44 25.4309 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=3.275 $Y=1.765
+ $X2=3.275 $Y2=1.542
r119 19 21 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.275 $Y=1.765
+ $X2=3.275 $Y2=2.4
r120 15 43 25.4309 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=3.16 $Y=1.32
+ $X2=3.16 $Y2=1.542
r121 15 17 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=3.16 $Y=1.32
+ $X2=3.16 $Y2=0.74
r122 12 39 25.4309 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=2.825 $Y=1.765
+ $X2=2.825 $Y2=1.542
r123 12 14 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.825 $Y=1.765
+ $X2=2.825 $Y2=2.4
r124 8 38 25.4309 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=2.73 $Y=1.32
+ $X2=2.73 $Y2=1.542
r125 8 10 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=2.73 $Y=1.32
+ $X2=2.73 $Y2=0.74
r126 5 34 25.4309 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=2.375 $Y=1.765
+ $X2=2.375 $Y2=1.542
r127 5 7 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.375 $Y=1.765
+ $X2=2.375 $Y2=2.4
r128 1 33 25.4309 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=2.3 $Y=1.32 $X2=2.3
+ $Y2=1.542
r129 1 3 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=2.3 $Y=1.32 $X2=2.3
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HS__A22OI_4%A1 1 3 4 8 10 12 15 17 19 22 24 26 29 31 33
+ 34 35 50
c90 50 0 3.11837e-19 $X=5.755 $Y=1.557
c91 35 0 1.97869e-19 $X=5.52 $Y=1.665
c92 24 0 1.34612e-19 $X=5.755 $Y=1.765
c93 4 0 9.91884e-20 $X=4.465 $Y=1.575
r94 50 51 10.0417 $w=3.6e-07 $l=7.5e-08 $layer=POLY_cond $X=5.755 $Y=1.557
+ $X2=5.83 $Y2=1.557
r95 48 50 46.1917 $w=3.6e-07 $l=3.45e-07 $layer=POLY_cond $X=5.41 $Y=1.557
+ $X2=5.755 $Y2=1.557
r96 48 49 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.41
+ $Y=1.515 $X2=5.41 $Y2=1.515
r97 46 48 1.33889 $w=3.6e-07 $l=1e-08 $layer=POLY_cond $X=5.4 $Y=1.557 $X2=5.41
+ $Y2=1.557
r98 45 46 43.5139 $w=3.6e-07 $l=3.25e-07 $layer=POLY_cond $X=5.075 $Y=1.557
+ $X2=5.4 $Y2=1.557
r99 44 49 9.11234 $w=4.28e-07 $l=3.4e-07 $layer=LI1_cond $X=5.07 $Y=1.565
+ $X2=5.41 $Y2=1.565
r100 43 45 0.669444 $w=3.6e-07 $l=5e-09 $layer=POLY_cond $X=5.07 $Y=1.557
+ $X2=5.075 $Y2=1.557
r101 43 44 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.07
+ $Y=1.515 $X2=5.07 $Y2=1.515
r102 41 43 13.3889 $w=3.6e-07 $l=1e-07 $layer=POLY_cond $X=4.97 $Y=1.557
+ $X2=5.07 $Y2=1.557
r103 40 41 46.1917 $w=3.6e-07 $l=3.45e-07 $layer=POLY_cond $X=4.625 $Y=1.557
+ $X2=4.97 $Y2=1.557
r104 39 40 11.3806 $w=3.6e-07 $l=8.5e-08 $layer=POLY_cond $X=4.54 $Y=1.557
+ $X2=4.625 $Y2=1.557
r105 35 49 2.94811 $w=4.28e-07 $l=1.1e-07 $layer=LI1_cond $X=5.52 $Y=1.565
+ $X2=5.41 $Y2=1.565
r106 34 44 0.80403 $w=4.28e-07 $l=3e-08 $layer=LI1_cond $X=5.04 $Y=1.565
+ $X2=5.07 $Y2=1.565
r107 33 34 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=4.56 $Y=1.565
+ $X2=5.04 $Y2=1.565
r108 27 51 23.3057 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=5.83 $Y=1.35
+ $X2=5.83 $Y2=1.557
r109 27 29 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=5.83 $Y=1.35
+ $X2=5.83 $Y2=0.74
r110 24 50 23.3057 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=5.755 $Y=1.765
+ $X2=5.755 $Y2=1.557
r111 24 26 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=5.755 $Y=1.765
+ $X2=5.755 $Y2=2.4
r112 20 46 23.3057 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=5.4 $Y=1.35
+ $X2=5.4 $Y2=1.557
r113 20 22 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=5.4 $Y=1.35 $X2=5.4
+ $Y2=0.74
r114 17 45 23.3057 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=5.075 $Y=1.765
+ $X2=5.075 $Y2=1.557
r115 17 19 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=5.075 $Y=1.765
+ $X2=5.075 $Y2=2.4
r116 13 41 23.3057 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.97 $Y=1.35
+ $X2=4.97 $Y2=1.557
r117 13 15 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=4.97 $Y=1.35
+ $X2=4.97 $Y2=0.74
r118 10 40 23.3057 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=4.625 $Y=1.765
+ $X2=4.625 $Y2=1.557
r119 10 12 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=4.625 $Y=1.765
+ $X2=4.625 $Y2=2.4
r120 6 39 23.3057 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.54 $Y=1.35
+ $X2=4.54 $Y2=1.557
r121 6 8 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=4.54 $Y=1.35 $X2=4.54
+ $Y2=0.74
r122 5 31 7.1379 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=4.265 $Y=1.575
+ $X2=4.175 $Y2=1.575
r123 4 39 26.8603 $w=3.6e-07 $l=8.35165e-08 $layer=POLY_cond $X=4.465 $Y=1.575
+ $X2=4.54 $Y2=1.557
r124 4 5 102.553 $w=1.5e-07 $l=2e-07 $layer=POLY_cond $X=4.465 $Y=1.575
+ $X2=4.265 $Y2=1.575
r125 1 31 76.0046 $w=1.8e-07 $l=1.9e-07 $layer=POLY_cond $X=4.175 $Y=1.765
+ $X2=4.175 $Y2=1.575
r126 1 3 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=4.175 $Y=1.765
+ $X2=4.175 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_HS__A22OI_4%A2 1 3 6 8 10 13 15 17 20 24 26 28 29 30 31
+ 46 47
c78 47 0 1.97869e-19 $X=7.55 $Y=1.557
c79 46 0 1.34612e-19 $X=7.3 $Y=1.515
c80 6 0 2.04552e-19 $X=6.26 $Y=0.74
r81 47 48 0.651351 $w=3.7e-07 $l=5e-09 $layer=POLY_cond $X=7.55 $Y=1.557
+ $X2=7.555 $Y2=1.557
r82 45 47 32.5676 $w=3.7e-07 $l=2.5e-07 $layer=POLY_cond $X=7.3 $Y=1.557
+ $X2=7.55 $Y2=1.557
r83 45 46 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=7.3
+ $Y=1.515 $X2=7.3 $Y2=1.515
r84 43 45 23.4486 $w=3.7e-07 $l=1.8e-07 $layer=POLY_cond $X=7.12 $Y=1.557
+ $X2=7.3 $Y2=1.557
r85 42 43 1.95405 $w=3.7e-07 $l=1.5e-08 $layer=POLY_cond $X=7.105 $Y=1.557
+ $X2=7.12 $Y2=1.557
r86 41 42 54.0622 $w=3.7e-07 $l=4.15e-07 $layer=POLY_cond $X=6.69 $Y=1.557
+ $X2=7.105 $Y2=1.557
r87 40 41 4.55946 $w=3.7e-07 $l=3.5e-08 $layer=POLY_cond $X=6.655 $Y=1.557
+ $X2=6.69 $Y2=1.557
r88 38 40 48.8514 $w=3.7e-07 $l=3.75e-07 $layer=POLY_cond $X=6.28 $Y=1.557
+ $X2=6.655 $Y2=1.557
r89 38 39 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.28
+ $Y=1.515 $X2=6.28 $Y2=1.515
r90 36 38 2.60541 $w=3.7e-07 $l=2e-08 $layer=POLY_cond $X=6.26 $Y=1.557 $X2=6.28
+ $Y2=1.557
r91 35 36 7.16487 $w=3.7e-07 $l=5.5e-08 $layer=POLY_cond $X=6.205 $Y=1.557
+ $X2=6.26 $Y2=1.557
r92 31 46 9.11234 $w=4.28e-07 $l=3.4e-07 $layer=LI1_cond $X=6.96 $Y=1.565
+ $X2=7.3 $Y2=1.565
r93 30 31 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=6.48 $Y=1.565
+ $X2=6.96 $Y2=1.565
r94 30 39 5.3602 $w=4.28e-07 $l=2e-07 $layer=LI1_cond $X=6.48 $Y=1.565 $X2=6.28
+ $Y2=1.565
r95 29 39 7.50428 $w=4.28e-07 $l=2.8e-07 $layer=LI1_cond $X=6 $Y=1.565 $X2=6.28
+ $Y2=1.565
r96 26 48 23.9667 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=7.555 $Y=1.765
+ $X2=7.555 $Y2=1.557
r97 26 28 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=7.555 $Y=1.765
+ $X2=7.555 $Y2=2.4
r98 22 47 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=7.55 $Y=1.35
+ $X2=7.55 $Y2=1.557
r99 22 24 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=7.55 $Y=1.35
+ $X2=7.55 $Y2=0.74
r100 18 43 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=7.12 $Y=1.35
+ $X2=7.12 $Y2=1.557
r101 18 20 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=7.12 $Y=1.35
+ $X2=7.12 $Y2=0.74
r102 15 42 23.9667 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=7.105 $Y=1.765
+ $X2=7.105 $Y2=1.557
r103 15 17 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=7.105 $Y=1.765
+ $X2=7.105 $Y2=2.4
r104 11 41 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=6.69 $Y=1.35
+ $X2=6.69 $Y2=1.557
r105 11 13 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=6.69 $Y=1.35
+ $X2=6.69 $Y2=0.74
r106 8 40 23.9667 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=6.655 $Y=1.765
+ $X2=6.655 $Y2=1.557
r107 8 10 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=6.655 $Y=1.765
+ $X2=6.655 $Y2=2.4
r108 4 36 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=6.26 $Y=1.35
+ $X2=6.26 $Y2=1.557
r109 4 6 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=6.26 $Y=1.35 $X2=6.26
+ $Y2=0.74
r110 1 35 23.9667 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=6.205 $Y=1.765
+ $X2=6.205 $Y2=1.557
r111 1 3 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=6.205 $Y=1.765
+ $X2=6.205 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_HS__A22OI_4%A_45_368# 1 2 3 4 5 6 7 8 9 30 34 35 38 40
+ 44 46 50 52 54 57 58 62 64 68 70 74 76 78 80 82 83 84 88 90 92
c150 90 0 1.16853e-19 $X=5.98 $Y=2.035
c151 58 0 1.94984e-19 $X=4.765 $Y=2.035
r152 78 94 3.1514 $w=2.5e-07 $l=1.5e-07 $layer=LI1_cond $X=7.82 $Y=2.12 $X2=7.82
+ $Y2=1.97
r153 78 80 12.9074 $w=2.48e-07 $l=2.8e-07 $layer=LI1_cond $X=7.82 $Y=2.12
+ $X2=7.82 $Y2=2.4
r154 77 92 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.965 $Y=2.035
+ $X2=6.88 $Y2=2.035
r155 76 94 3.99177 $w=1.7e-07 $l=1.5411e-07 $layer=LI1_cond $X=7.695 $Y=2.035
+ $X2=7.82 $Y2=1.97
r156 76 77 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=7.695 $Y=2.035
+ $X2=6.965 $Y2=2.035
r157 72 92 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.88 $Y=2.12
+ $X2=6.88 $Y2=2.035
r158 72 74 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=6.88 $Y=2.12
+ $X2=6.88 $Y2=2.465
r159 71 90 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.065 $Y=2.035
+ $X2=5.94 $Y2=2.035
r160 70 92 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.795 $Y=2.035
+ $X2=6.88 $Y2=2.035
r161 70 71 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=6.795 $Y=2.035
+ $X2=6.065 $Y2=2.035
r162 66 90 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.94 $Y=2.12
+ $X2=5.94 $Y2=2.035
r163 66 68 15.9037 $w=2.48e-07 $l=3.45e-07 $layer=LI1_cond $X=5.94 $Y=2.12
+ $X2=5.94 $Y2=2.465
r164 65 88 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.015 $Y=2.035
+ $X2=4.89 $Y2=2.035
r165 64 90 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.815 $Y=2.035
+ $X2=5.94 $Y2=2.035
r166 64 65 52.1925 $w=1.68e-07 $l=8e-07 $layer=LI1_cond $X=5.815 $Y=2.035
+ $X2=5.015 $Y2=2.035
r167 60 88 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.89 $Y=2.12
+ $X2=4.89 $Y2=2.035
r168 60 62 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=4.89 $Y=2.12
+ $X2=4.89 $Y2=2.415
r169 59 86 3.99177 $w=1.7e-07 $l=1.5411e-07 $layer=LI1_cond $X=4.035 $Y=2.035
+ $X2=3.91 $Y2=1.97
r170 58 88 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.765 $Y=2.035
+ $X2=4.89 $Y2=2.035
r171 58 59 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=4.765 $Y=2.035
+ $X2=4.035 $Y2=2.035
r172 55 57 23.2793 $w=2.48e-07 $l=5.05e-07 $layer=LI1_cond $X=3.91 $Y=2.905
+ $X2=3.91 $Y2=2.4
r173 54 86 3.1514 $w=2.5e-07 $l=1.5e-07 $layer=LI1_cond $X=3.91 $Y=2.12 $X2=3.91
+ $Y2=1.97
r174 54 57 12.9074 $w=2.48e-07 $l=2.8e-07 $layer=LI1_cond $X=3.91 $Y=2.12
+ $X2=3.91 $Y2=2.4
r175 53 84 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.215 $Y=2.99
+ $X2=3.05 $Y2=2.99
r176 52 55 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=3.785 $Y=2.99
+ $X2=3.91 $Y2=2.905
r177 52 53 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=3.785 $Y=2.99
+ $X2=3.215 $Y2=2.99
r178 48 84 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.05 $Y=2.905
+ $X2=3.05 $Y2=2.99
r179 48 50 18.5089 $w=3.28e-07 $l=5.3e-07 $layer=LI1_cond $X=3.05 $Y=2.905
+ $X2=3.05 $Y2=2.375
r180 47 83 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.315 $Y=2.99
+ $X2=2.15 $Y2=2.99
r181 46 84 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.885 $Y=2.99
+ $X2=3.05 $Y2=2.99
r182 46 47 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=2.885 $Y=2.99
+ $X2=2.315 $Y2=2.99
r183 42 83 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.15 $Y=2.905
+ $X2=2.15 $Y2=2.99
r184 42 44 18.5089 $w=3.28e-07 $l=5.3e-07 $layer=LI1_cond $X=2.15 $Y=2.905
+ $X2=2.15 $Y2=2.375
r185 41 82 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.415 $Y=2.99
+ $X2=1.25 $Y2=2.99
r186 40 83 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.985 $Y=2.99
+ $X2=2.15 $Y2=2.99
r187 40 41 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=1.985 $Y=2.99
+ $X2=1.415 $Y2=2.99
r188 36 82 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.25 $Y=2.905
+ $X2=1.25 $Y2=2.99
r189 36 38 18.5089 $w=3.28e-07 $l=5.3e-07 $layer=LI1_cond $X=1.25 $Y=2.905
+ $X2=1.25 $Y2=2.375
r190 34 82 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.085 $Y=2.99
+ $X2=1.25 $Y2=2.99
r191 34 35 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=1.085 $Y=2.99
+ $X2=0.435 $Y2=2.99
r192 30 33 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=0.31 $Y=1.985
+ $X2=0.31 $Y2=2.815
r193 28 35 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.31 $Y=2.905
+ $X2=0.435 $Y2=2.99
r194 28 33 4.14879 $w=2.48e-07 $l=9e-08 $layer=LI1_cond $X=0.31 $Y=2.905
+ $X2=0.31 $Y2=2.815
r195 9 94 600 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=7.63
+ $Y=1.84 $X2=7.78 $Y2=1.985
r196 9 80 300 $w=1.7e-07 $l=6.30555e-07 $layer=licon1_PDIFF $count=2 $X=7.63
+ $Y=1.84 $X2=7.78 $Y2=2.4
r197 8 92 600 $w=1.7e-07 $l=2.59374e-07 $layer=licon1_PDIFF $count=1 $X=6.73
+ $Y=1.84 $X2=6.88 $Y2=2.035
r198 8 74 300 $w=1.7e-07 $l=6.95971e-07 $layer=licon1_PDIFF $count=2 $X=6.73
+ $Y=1.84 $X2=6.88 $Y2=2.465
r199 7 90 600 $w=1.7e-07 $l=2.59374e-07 $layer=licon1_PDIFF $count=1 $X=5.83
+ $Y=1.84 $X2=5.98 $Y2=2.035
r200 7 68 300 $w=1.7e-07 $l=6.95971e-07 $layer=licon1_PDIFF $count=2 $X=5.83
+ $Y=1.84 $X2=5.98 $Y2=2.465
r201 6 88 600 $w=1.7e-07 $l=2.59374e-07 $layer=licon1_PDIFF $count=1 $X=4.7
+ $Y=1.84 $X2=4.85 $Y2=2.035
r202 6 62 300 $w=1.7e-07 $l=6.45659e-07 $layer=licon1_PDIFF $count=2 $X=4.7
+ $Y=1.84 $X2=4.85 $Y2=2.415
r203 5 86 600 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=3.8
+ $Y=1.84 $X2=3.95 $Y2=1.985
r204 5 57 300 $w=1.7e-07 $l=6.30555e-07 $layer=licon1_PDIFF $count=2 $X=3.8
+ $Y=1.84 $X2=3.95 $Y2=2.4
r205 4 50 300 $w=1.7e-07 $l=6.05372e-07 $layer=licon1_PDIFF $count=2 $X=2.9
+ $Y=1.84 $X2=3.05 $Y2=2.375
r206 3 44 300 $w=1.7e-07 $l=6.05372e-07 $layer=licon1_PDIFF $count=2 $X=2
+ $Y=1.84 $X2=2.15 $Y2=2.375
r207 2 38 300 $w=1.7e-07 $l=6.05372e-07 $layer=licon1_PDIFF $count=2 $X=1.1
+ $Y=1.84 $X2=1.25 $Y2=2.375
r208 1 33 400 $w=1.7e-07 $l=1.03562e-06 $layer=licon1_PDIFF $count=1 $X=0.225
+ $Y=1.84 $X2=0.35 $Y2=2.815
r209 1 30 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.225
+ $Y=1.84 $X2=0.35 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HS__A22OI_4%Y 1 2 3 4 5 6 7 8 25 27 29 33 35 39 43 45 46
+ 47 52 54 60 62 64 66 67 69 70
c114 67 0 9.91884e-20 $X=5.45 $Y=0.95
c115 66 0 4.29123e-20 $X=5.615 $Y=0.95
c116 46 0 8.01953e-20 $X=2.68 $Y=1.095
c117 35 0 1.91457e-19 $X=2.515 $Y=2.035
r118 74 75 2.90031 $w=6.52e-07 $l=1.55e-07 $layer=LI1_cond $X=3.375 $Y=1.145
+ $X2=3.53 $Y2=1.145
r119 69 70 8.9816 $w=6.52e-07 $l=4.8e-07 $layer=LI1_cond $X=3.6 $Y=1.145
+ $X2=4.08 $Y2=1.145
r120 69 75 1.30982 $w=6.52e-07 $l=7e-08 $layer=LI1_cond $X=3.6 $Y=1.145 $X2=3.53
+ $Y2=1.145
r121 66 67 5.88189 $w=3.58e-07 $l=1.65e-07 $layer=LI1_cond $X=5.615 $Y=0.95
+ $X2=5.45 $Y2=0.95
r122 56 67 28.6053 $w=2.78e-07 $l=6.95e-07 $layer=LI1_cond $X=4.755 $Y=0.99
+ $X2=5.45 $Y2=0.99
r123 54 70 6.20325 $w=6.52e-07 $l=2.04573e-07 $layer=LI1_cond $X=4.195 $Y=0.99
+ $X2=4.08 $Y2=1.145
r124 54 56 23.0489 $w=2.78e-07 $l=5.6e-07 $layer=LI1_cond $X=4.195 $Y=0.99
+ $X2=4.755 $Y2=0.99
r125 52 64 4.81226 $w=1.85e-07 $l=9.21954e-08 $layer=LI1_cond $X=3.53 $Y=1.95
+ $X2=3.515 $Y2=2.035
r126 51 75 8.85584 $w=1.7e-07 $l=3.75e-07 $layer=LI1_cond $X=3.53 $Y=1.52
+ $X2=3.53 $Y2=1.145
r127 51 52 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=3.53 $Y=1.52
+ $X2=3.53 $Y2=1.95
r128 48 62 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.685 $Y=2.035
+ $X2=2.6 $Y2=2.035
r129 47 64 1.64875 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=3.415 $Y=2.035
+ $X2=3.515 $Y2=2.035
r130 47 48 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=3.415 $Y=2.035
+ $X2=2.685 $Y2=2.035
r131 45 74 10.7048 $w=6.52e-07 $l=1.88348e-07 $layer=LI1_cond $X=3.21 $Y=1.095
+ $X2=3.375 $Y2=1.145
r132 45 46 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=3.21 $Y=1.095
+ $X2=2.68 $Y2=1.095
r133 41 62 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.6 $Y=2.12 $X2=2.6
+ $Y2=2.035
r134 41 43 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=2.6 $Y=2.12 $X2=2.6
+ $Y2=2.57
r135 37 46 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.515 $Y=1.01
+ $X2=2.68 $Y2=1.095
r136 37 39 8.73063 $w=3.28e-07 $l=2.5e-07 $layer=LI1_cond $X=2.515 $Y=1.01
+ $X2=2.515 $Y2=0.76
r137 36 60 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.785 $Y=2.035
+ $X2=1.7 $Y2=2.035
r138 35 62 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.515 $Y=2.035
+ $X2=2.6 $Y2=2.035
r139 35 36 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=2.515 $Y=2.035
+ $X2=1.785 $Y2=2.035
r140 31 60 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.7 $Y=2.12 $X2=1.7
+ $Y2=2.035
r141 31 33 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=1.7 $Y=2.12 $X2=1.7
+ $Y2=2.57
r142 30 58 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.885 $Y=2.035
+ $X2=0.76 $Y2=2.035
r143 29 60 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.615 $Y=2.035
+ $X2=1.7 $Y2=2.035
r144 29 30 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=1.615 $Y=2.035
+ $X2=0.885 $Y2=2.035
r145 25 58 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.76 $Y=2.12
+ $X2=0.76 $Y2=2.035
r146 25 27 20.744 $w=2.48e-07 $l=4.5e-07 $layer=LI1_cond $X=0.76 $Y=2.12
+ $X2=0.76 $Y2=2.57
r147 8 64 300 $w=1.7e-07 $l=3.4187e-07 $layer=licon1_PDIFF $count=2 $X=3.35
+ $Y=1.84 $X2=3.5 $Y2=2.115
r148 7 62 600 $w=1.7e-07 $l=2.59374e-07 $layer=licon1_PDIFF $count=1 $X=2.45
+ $Y=1.84 $X2=2.6 $Y2=2.035
r149 7 43 600 $w=1.7e-07 $l=8.01499e-07 $layer=licon1_PDIFF $count=1 $X=2.45
+ $Y=1.84 $X2=2.6 $Y2=2.57
r150 6 60 600 $w=1.7e-07 $l=2.59374e-07 $layer=licon1_PDIFF $count=1 $X=1.55
+ $Y=1.84 $X2=1.7 $Y2=2.035
r151 6 33 600 $w=1.7e-07 $l=8.01499e-07 $layer=licon1_PDIFF $count=1 $X=1.55
+ $Y=1.84 $X2=1.7 $Y2=2.57
r152 5 58 600 $w=1.7e-07 $l=2.59374e-07 $layer=licon1_PDIFF $count=1 $X=0.65
+ $Y=1.84 $X2=0.8 $Y2=2.035
r153 5 27 600 $w=1.7e-07 $l=8.01499e-07 $layer=licon1_PDIFF $count=1 $X=0.65
+ $Y=1.84 $X2=0.8 $Y2=2.57
r154 4 66 182 $w=1.7e-07 $l=6.4622e-07 $layer=licon1_NDIFF $count=1 $X=5.475
+ $Y=0.37 $X2=5.615 $Y2=0.95
r155 3 56 182 $w=1.7e-07 $l=6.4622e-07 $layer=licon1_NDIFF $count=1 $X=4.615
+ $Y=0.37 $X2=4.755 $Y2=0.95
r156 2 74 182 $w=1.7e-07 $l=6.0597e-07 $layer=licon1_NDIFF $count=1 $X=3.235
+ $Y=0.37 $X2=3.375 $Y2=0.91
r157 1 39 182 $w=1.7e-07 $l=4.54643e-07 $layer=licon1_NDIFF $count=1 $X=2.375
+ $Y=0.37 $X2=2.515 $Y2=0.76
.ends

.subckt PM_SKY130_FD_SC_HS__A22OI_4%VPWR 1 2 3 4 15 19 23 27 30 31 33 34 35 44
+ 48 58 59 62 65
r101 65 66 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r102 62 63 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r103 58 59 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r104 56 59 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=7.92 $Y2=3.33
r105 56 66 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=6.48 $Y2=3.33
r106 55 56 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r107 53 65 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.595 $Y=3.33
+ $X2=6.43 $Y2=3.33
r108 53 55 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=6.595 $Y=3.33
+ $X2=6.96 $Y2=3.33
r109 52 66 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=3.33 $X2=6.48
+ $Y2=3.33
r110 52 63 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=3.33 $X2=5.52
+ $Y2=3.33
r111 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r112 49 62 10.7288 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=5.645 $Y=3.33
+ $X2=5.415 $Y2=3.33
r113 49 51 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=5.645 $Y=3.33
+ $X2=6 $Y2=3.33
r114 48 65 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.265 $Y=3.33
+ $X2=6.43 $Y2=3.33
r115 48 51 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=6.265 $Y=3.33
+ $X2=6 $Y2=3.33
r116 47 63 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=5.52 $Y2=3.33
r117 46 47 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r118 44 62 10.7288 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=5.185 $Y=3.33
+ $X2=5.415 $Y2=3.33
r119 44 46 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=5.185 $Y=3.33
+ $X2=5.04 $Y2=3.33
r120 38 42 250.524 $w=1.68e-07 $l=3.84e-06 $layer=LI1_cond $X=0.24 $Y=3.33
+ $X2=4.08 $Y2=3.33
r121 38 39 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r122 35 47 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=5.04 $Y2=3.33
r123 35 39 1.07034 $w=4.9e-07 $l=3.84e-06 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=0.24 $Y2=3.33
r124 35 42 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r125 33 55 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=7.165 $Y=3.33
+ $X2=6.96 $Y2=3.33
r126 33 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.165 $Y=3.33
+ $X2=7.33 $Y2=3.33
r127 32 58 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=7.495 $Y=3.33
+ $X2=7.92 $Y2=3.33
r128 32 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.495 $Y=3.33
+ $X2=7.33 $Y2=3.33
r129 30 42 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=4.235 $Y=3.33
+ $X2=4.08 $Y2=3.33
r130 30 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.235 $Y=3.33
+ $X2=4.4 $Y2=3.33
r131 29 46 30.9893 $w=1.68e-07 $l=4.75e-07 $layer=LI1_cond $X=4.565 $Y=3.33
+ $X2=5.04 $Y2=3.33
r132 29 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.565 $Y=3.33
+ $X2=4.4 $Y2=3.33
r133 25 34 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.33 $Y=3.245
+ $X2=7.33 $Y2=3.33
r134 25 27 30.3826 $w=3.28e-07 $l=8.7e-07 $layer=LI1_cond $X=7.33 $Y=3.245
+ $X2=7.33 $Y2=2.375
r135 21 65 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.43 $Y=3.245
+ $X2=6.43 $Y2=3.33
r136 21 23 30.3826 $w=3.28e-07 $l=8.7e-07 $layer=LI1_cond $X=6.43 $Y=3.245
+ $X2=6.43 $Y2=2.375
r137 17 62 1.85547 $w=4.6e-07 $l=8.5e-08 $layer=LI1_cond $X=5.415 $Y=3.245
+ $X2=5.415 $Y2=3.33
r138 17 19 22.6215 $w=4.58e-07 $l=8.7e-07 $layer=LI1_cond $X=5.415 $Y=3.245
+ $X2=5.415 $Y2=2.375
r139 13 31 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.4 $Y=3.245 $X2=4.4
+ $Y2=3.33
r140 13 15 30.3826 $w=3.28e-07 $l=8.7e-07 $layer=LI1_cond $X=4.4 $Y=3.245
+ $X2=4.4 $Y2=2.375
r141 4 27 300 $w=1.7e-07 $l=6.05372e-07 $layer=licon1_PDIFF $count=2 $X=7.18
+ $Y=1.84 $X2=7.33 $Y2=2.375
r142 3 23 300 $w=1.7e-07 $l=6.05372e-07 $layer=licon1_PDIFF $count=2 $X=6.28
+ $Y=1.84 $X2=6.43 $Y2=2.375
r143 2 19 300 $w=1.7e-07 $l=6.54217e-07 $layer=licon1_PDIFF $count=2 $X=5.15
+ $Y=1.84 $X2=5.415 $Y2=2.375
r144 1 15 300 $w=1.7e-07 $l=6.05372e-07 $layer=licon1_PDIFF $count=2 $X=4.25
+ $Y=1.84 $X2=4.4 $Y2=2.375
.ends

.subckt PM_SKY130_FD_SC_HS__A22OI_4%A_48_74# 1 2 3 4 5 18 20 21 24 26 32 33 36
+ 38 39
r66 34 43 10.9604 $w=1.68e-07 $l=1.68e-07 $layer=LI1_cond $X=2.945 $Y=0.427
+ $X2=2.945 $Y2=0.595
r67 34 39 5.67594 $w=1.68e-07 $l=8.7e-08 $layer=LI1_cond $X=2.945 $Y=0.427
+ $X2=2.945 $Y2=0.34
r68 34 36 25.8882 $w=3.43e-07 $l=7.75e-07 $layer=LI1_cond $X=3.03 $Y=0.427
+ $X2=3.805 $Y2=0.427
r69 32 39 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.86 $Y=0.34
+ $X2=2.945 $Y2=0.34
r70 32 33 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=2.86 $Y=0.34 $X2=2.17
+ $Y2=0.34
r71 29 31 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=2.085 $Y=1.01
+ $X2=2.085 $Y2=0.515
r72 28 33 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.085 $Y=0.425
+ $X2=2.17 $Y2=0.34
r73 28 31 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=2.085 $Y=0.425
+ $X2=2.085 $Y2=0.515
r74 27 38 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.31 $Y=1.095
+ $X2=1.185 $Y2=1.095
r75 26 29 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2 $Y=1.095
+ $X2=2.085 $Y2=1.01
r76 26 27 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=2 $Y=1.095 $X2=1.31
+ $Y2=1.095
r77 22 38 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.185 $Y=1.01
+ $X2=1.185 $Y2=1.095
r78 22 24 22.8184 $w=2.48e-07 $l=4.95e-07 $layer=LI1_cond $X=1.185 $Y=1.01
+ $X2=1.185 $Y2=0.515
r79 20 38 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.06 $Y=1.095
+ $X2=1.185 $Y2=1.095
r80 20 21 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=1.06 $Y=1.095
+ $X2=0.45 $Y2=1.095
r81 16 21 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.325 $Y=1.01
+ $X2=0.45 $Y2=1.095
r82 16 18 22.8184 $w=2.48e-07 $l=4.95e-07 $layer=LI1_cond $X=0.325 $Y=1.01
+ $X2=0.325 $Y2=0.515
r83 5 36 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=3.665
+ $Y=0.37 $X2=3.805 $Y2=0.515
r84 4 43 182 $w=1.7e-07 $l=2.86575e-07 $layer=licon1_NDIFF $count=1 $X=2.805
+ $Y=0.37 $X2=2.945 $Y2=0.595
r85 3 31 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.945
+ $Y=0.37 $X2=2.085 $Y2=0.515
r86 2 24 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.085
+ $Y=0.37 $X2=1.225 $Y2=0.515
r87 1 18 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.24
+ $Y=0.37 $X2=0.365 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__A22OI_4%VGND 1 2 3 4 15 19 23 27 30 31 33 34 35 37
+ 42 58 59 62 65
c94 19 0 1.9142e-19 $X=1.655 $Y=0.675
r95 65 66 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r96 62 63 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r97 58 59 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.92 $Y=0 $X2=7.92
+ $Y2=0
r98 56 59 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.96 $Y=0 $X2=7.92
+ $Y2=0
r99 55 56 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.96 $Y=0 $X2=6.96
+ $Y2=0
r100 53 56 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6 $Y=0 $X2=6.96
+ $Y2=0
r101 52 53 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=6 $Y=0 $X2=6
+ $Y2=0
r102 50 66 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.68
+ $Y2=0
r103 49 52 250.524 $w=1.68e-07 $l=3.84e-06 $layer=LI1_cond $X=2.16 $Y=0 $X2=6
+ $Y2=0
r104 49 50 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=2.16 $Y=0
+ $X2=2.16 $Y2=0
r105 47 65 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.82 $Y=0 $X2=1.655
+ $Y2=0
r106 47 49 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=1.82 $Y=0 $X2=2.16
+ $Y2=0
r107 46 66 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=1.68
+ $Y2=0
r108 46 63 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r109 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r110 43 62 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.88 $Y=0 $X2=0.755
+ $Y2=0
r111 43 45 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=0.88 $Y=0 $X2=1.2
+ $Y2=0
r112 42 65 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.49 $Y=0 $X2=1.655
+ $Y2=0
r113 42 45 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=1.49 $Y=0 $X2=1.2
+ $Y2=0
r114 40 63 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r115 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r116 37 62 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.63 $Y=0 $X2=0.755
+ $Y2=0
r117 37 39 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=0.63 $Y=0 $X2=0.24
+ $Y2=0
r118 35 53 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=4.08 $Y=0 $X2=6
+ $Y2=0
r119 35 50 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=4.08 $Y=0
+ $X2=2.16 $Y2=0
r120 33 55 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=7.17 $Y=0 $X2=6.96
+ $Y2=0
r121 33 34 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.17 $Y=0 $X2=7.295
+ $Y2=0
r122 32 58 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=7.42 $Y=0 $X2=7.92
+ $Y2=0
r123 32 34 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.42 $Y=0 $X2=7.295
+ $Y2=0
r124 30 52 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=6.31 $Y=0 $X2=6
+ $Y2=0
r125 30 31 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.31 $Y=0 $X2=6.435
+ $Y2=0
r126 29 55 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=6.56 $Y=0 $X2=6.96
+ $Y2=0
r127 29 31 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.56 $Y=0 $X2=6.435
+ $Y2=0
r128 25 34 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=7.295 $Y=0.085
+ $X2=7.295 $Y2=0
r129 25 27 23.5098 $w=2.48e-07 $l=5.1e-07 $layer=LI1_cond $X=7.295 $Y=0.085
+ $X2=7.295 $Y2=0.595
r130 21 31 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.435 $Y=0.085
+ $X2=6.435 $Y2=0
r131 21 23 23.5098 $w=2.48e-07 $l=5.1e-07 $layer=LI1_cond $X=6.435 $Y=0.085
+ $X2=6.435 $Y2=0.595
r132 17 65 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.655 $Y=0.085
+ $X2=1.655 $Y2=0
r133 17 19 20.6043 $w=3.28e-07 $l=5.9e-07 $layer=LI1_cond $X=1.655 $Y=0.085
+ $X2=1.655 $Y2=0.675
r134 13 62 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.755 $Y=0.085
+ $X2=0.755 $Y2=0
r135 13 15 27.1977 $w=2.48e-07 $l=5.9e-07 $layer=LI1_cond $X=0.755 $Y=0.085
+ $X2=0.755 $Y2=0.675
r136 4 27 182 $w=1.7e-07 $l=2.86575e-07 $layer=licon1_NDIFF $count=1 $X=7.195
+ $Y=0.37 $X2=7.335 $Y2=0.595
r137 3 23 182 $w=1.7e-07 $l=2.86575e-07 $layer=licon1_NDIFF $count=1 $X=6.335
+ $Y=0.37 $X2=6.475 $Y2=0.595
r138 2 19 182 $w=1.7e-07 $l=3.68409e-07 $layer=licon1_NDIFF $count=1 $X=1.515
+ $Y=0.37 $X2=1.655 $Y2=0.675
r139 1 15 182 $w=1.7e-07 $l=3.68409e-07 $layer=licon1_NDIFF $count=1 $X=0.655
+ $Y=0.37 $X2=0.795 $Y2=0.675
.ends

.subckt PM_SKY130_FD_SC_HS__A22OI_4%A_840_74# 1 2 3 4 5 16 20 24 25 28 30 34 39
+ 42
c62 20 0 1.6164e-19 $X=6.045 $Y=0.6
r63 37 39 6.46688 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=4.325 $Y=0.515
+ $X2=4.49 $Y2=0.515
r64 32 34 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=7.765 $Y=1.01
+ $X2=7.765 $Y2=0.515
r65 31 42 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.99 $Y=1.095
+ $X2=6.865 $Y2=1.095
r66 30 32 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=7.6 $Y=1.095
+ $X2=7.765 $Y2=1.01
r67 30 31 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=7.6 $Y=1.095
+ $X2=6.99 $Y2=1.095
r68 26 42 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.865 $Y=1.01
+ $X2=6.865 $Y2=1.095
r69 26 28 22.8184 $w=2.48e-07 $l=4.95e-07 $layer=LI1_cond $X=6.865 $Y=1.01
+ $X2=6.865 $Y2=0.515
r70 24 42 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.74 $Y=1.095
+ $X2=6.865 $Y2=1.095
r71 24 25 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=6.74 $Y=1.095
+ $X2=6.13 $Y2=1.095
r72 21 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.045 $Y=1.01
+ $X2=6.13 $Y2=1.095
r73 21 23 2.93583 $w=1.68e-07 $l=4.5e-08 $layer=LI1_cond $X=6.045 $Y=1.01
+ $X2=6.045 $Y2=0.965
r74 20 41 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.045 $Y=0.6
+ $X2=6.045 $Y2=0.475
r75 20 23 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=6.045 $Y=0.6
+ $X2=6.045 $Y2=0.965
r76 19 39 32.0379 $w=2.48e-07 $l=6.95e-07 $layer=LI1_cond $X=5.185 $Y=0.475
+ $X2=4.49 $Y2=0.475
r77 16 41 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.96 $Y=0.475
+ $X2=6.045 $Y2=0.475
r78 16 19 35.7257 $w=2.48e-07 $l=7.75e-07 $layer=LI1_cond $X=5.96 $Y=0.475
+ $X2=5.185 $Y2=0.475
r79 5 34 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=7.625
+ $Y=0.37 $X2=7.765 $Y2=0.515
r80 4 28 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=6.765
+ $Y=0.37 $X2=6.905 $Y2=0.515
r81 3 41 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=5.905
+ $Y=0.37 $X2=6.045 $Y2=0.515
r82 3 23 182 $w=1.7e-07 $l=6.61306e-07 $layer=licon1_NDIFF $count=1 $X=5.905
+ $Y=0.37 $X2=6.045 $Y2=0.965
r83 2 19 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=5.045
+ $Y=0.37 $X2=5.185 $Y2=0.515
r84 1 37 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=4.2
+ $Y=0.37 $X2=4.325 $Y2=0.515
.ends

