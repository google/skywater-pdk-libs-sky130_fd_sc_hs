* NGSPICE file created from sky130_fd_sc_hs__or4_4.ext - technology: sky130A

.subckt sky130_fd_sc_hs__or4_4 A B C D VGND VNB VPB VPWR X
M1000 VPWR A a_588_392# VPB pshort w=1e+06u l=150000u
+  ad=1.2968e+12p pd=1.11e+07u as=6.2e+11p ps=5.24e+06u
M1001 a_588_392# A VPWR VPB pshort w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1002 VGND a_83_264# X VNB nlowvt w=740000u l=150000u
+  ad=2.2402e+12p pd=1.413e+07u as=6.549e+11p ps=4.73e+06u
M1003 a_83_264# B VGND VNB nlowvt w=740000u l=150000u
+  ad=4.662e+11p pd=4.22e+06u as=0p ps=0u
M1004 X a_83_264# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VGND D a_83_264# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VGND a_83_264# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 X a_83_264# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_962_392# C a_499_392# VPB pshort w=1e+06u l=150000u
+  ad=6.5e+11p pd=5.3e+06u as=9.9e+11p ps=7.98e+06u
M1009 a_499_392# B a_588_392# VPB pshort w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VPWR a_83_264# X VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=6.72e+11p ps=5.68e+06u
M1011 X a_83_264# VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 X a_83_264# VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VGND A a_83_264# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_83_264# D a_962_392# VPB pshort w=1e+06u l=150000u
+  ad=3e+11p pd=2.6e+06u as=0p ps=0u
M1015 a_83_264# C VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VPWR a_83_264# X VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_962_392# D a_83_264# VPB pshort w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_499_392# C a_962_392# VPB pshort w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_588_392# B a_499_392# VPB pshort w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

