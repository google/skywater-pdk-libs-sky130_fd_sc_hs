# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_hs__a21boi_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.320000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.558000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.485000 1.320000 2.815000 1.780000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.558000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.265000 1.220000 3.715000 1.550000 ;
        RECT 3.485000 1.180000 3.715000 1.220000 ;
    END
  END A2
  PIN B1_N
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.450000 0.475000 1.780000 ;
    END
  END B1_N
  PIN Y
    ANTENNADIFFAREA  0.750400 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.270000 0.350000 1.440000 0.980000 ;
        RECT 1.270000 0.980000 2.900000 1.150000 ;
        RECT 1.615000 1.150000 2.275000 1.410000 ;
        RECT 1.615000 1.410000 1.945000 2.735000 ;
        RECT 2.570000 0.770000 2.900000 0.980000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 4.320000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 4.320000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.320000 0.085000 ;
      RECT 0.000000  3.245000 4.320000 3.415000 ;
      RECT 0.195000  1.950000 0.445000 3.245000 ;
      RECT 0.270000  0.450000 0.520000 1.110000 ;
      RECT 0.270000  1.110000 0.975000 1.280000 ;
      RECT 0.645000  1.940000 0.975000 2.980000 ;
      RECT 0.760000  0.085000 1.090000 0.940000 ;
      RECT 0.805000  1.280000 0.975000 1.320000 ;
      RECT 0.805000  1.320000 1.395000 1.650000 ;
      RECT 0.805000  1.650000 0.975000 1.940000 ;
      RECT 1.165000  1.820000 1.415000 2.905000 ;
      RECT 1.165000  2.905000 2.315000 3.075000 ;
      RECT 1.620000  0.085000 1.950000 0.810000 ;
      RECT 2.115000  1.820000 2.315000 1.950000 ;
      RECT 2.115000  1.950000 3.215000 2.120000 ;
      RECT 2.115000  2.120000 2.315000 2.905000 ;
      RECT 2.140000  0.350000 3.250000 0.600000 ;
      RECT 2.515000  2.290000 2.845000 3.245000 ;
      RECT 3.045000  1.720000 4.215000 1.890000 ;
      RECT 3.045000  1.890000 3.215000 1.950000 ;
      RECT 3.045000  2.120000 3.215000 2.980000 ;
      RECT 3.080000  0.600000 3.250000 0.840000 ;
      RECT 3.080000  0.840000 4.190000 1.010000 ;
      RECT 3.080000  1.010000 3.250000 1.050000 ;
      RECT 3.415000  2.060000 3.765000 3.245000 ;
      RECT 3.430000  0.085000 3.760000 0.670000 ;
      RECT 3.940000  0.350000 4.190000 0.840000 ;
      RECT 3.940000  1.010000 4.190000 1.130000 ;
      RECT 3.965000  1.890000 4.215000 2.980000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
  END
END sky130_fd_sc_hs__a21boi_2
