* File: sky130_fd_sc_hs__nand2_4.pex.spice
* Created: Tue Sep  1 20:08:42 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HS__NAND2_4%B 3 5 7 10 14 16 18 21 28 29 30 42 44 52
c60 42 0 1.62664e-19 $X=1.77 $Y=1.557
r61 42 43 2.05983 $w=3.51e-07 $l=1.5e-08 $layer=POLY_cond $X=1.77 $Y=1.557
+ $X2=1.785 $Y2=1.557
r62 40 42 10.2991 $w=3.51e-07 $l=7.5e-08 $layer=POLY_cond $X=1.695 $Y=1.557
+ $X2=1.77 $Y2=1.557
r63 40 41 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.695
+ $Y=1.515 $X2=1.695 $Y2=1.515
r64 38 40 46.6895 $w=3.51e-07 $l=3.4e-07 $layer=POLY_cond $X=1.355 $Y=1.557
+ $X2=1.695 $Y2=1.557
r65 37 38 59.0484 $w=3.51e-07 $l=4.3e-07 $layer=POLY_cond $X=0.925 $Y=1.557
+ $X2=1.355 $Y2=1.557
r66 34 35 2.05983 $w=3.51e-07 $l=1.5e-08 $layer=POLY_cond $X=0.495 $Y=1.557
+ $X2=0.51 $Y2=1.557
r67 30 41 12.4625 $w=4.28e-07 $l=4.65e-07 $layer=LI1_cond $X=2.16 $Y=1.565
+ $X2=1.695 $Y2=1.565
r68 29 41 0.402015 $w=4.28e-07 $l=1.5e-08 $layer=LI1_cond $X=1.68 $Y=1.565
+ $X2=1.695 $Y2=1.565
r69 29 44 4.42216 $w=4.28e-07 $l=1.65e-07 $layer=LI1_cond $X=1.68 $Y=1.565
+ $X2=1.515 $Y2=1.565
r70 28 44 8.44232 $w=4.28e-07 $l=3.15e-07 $layer=LI1_cond $X=1.2 $Y=1.565
+ $X2=1.515 $Y2=1.565
r71 28 52 3.73456 $w=4.28e-07 $l=1.15e-07 $layer=LI1_cond $X=1.2 $Y=1.565
+ $X2=1.085 $Y2=1.565
r72 26 37 34.3305 $w=3.51e-07 $l=2.5e-07 $layer=POLY_cond $X=0.675 $Y=1.557
+ $X2=0.925 $Y2=1.557
r73 26 35 22.6581 $w=3.51e-07 $l=1.65e-07 $layer=POLY_cond $X=0.675 $Y=1.557
+ $X2=0.51 $Y2=1.557
r74 25 52 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=0.675 $Y=1.515
+ $X2=1.085 $Y2=1.515
r75 25 26 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.675
+ $Y=1.515 $X2=0.675 $Y2=1.515
r76 19 43 22.6971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.785 $Y=1.35
+ $X2=1.785 $Y2=1.557
r77 19 21 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.785 $Y=1.35
+ $X2=1.785 $Y2=0.74
r78 16 42 22.6971 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=1.77 $Y=1.765
+ $X2=1.77 $Y2=1.557
r79 16 18 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.77 $Y=1.765
+ $X2=1.77 $Y2=2.4
r80 12 38 22.6971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.355 $Y=1.35
+ $X2=1.355 $Y2=1.557
r81 12 14 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.355 $Y=1.35
+ $X2=1.355 $Y2=0.74
r82 8 37 22.6971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.925 $Y=1.35
+ $X2=0.925 $Y2=1.557
r83 8 10 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=0.925 $Y=1.35
+ $X2=0.925 $Y2=0.74
r84 5 35 22.6971 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=0.51 $Y=1.765
+ $X2=0.51 $Y2=1.557
r85 5 7 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.51 $Y=1.765
+ $X2=0.51 $Y2=2.4
r86 1 34 22.6971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.495 $Y=1.35
+ $X2=0.495 $Y2=1.557
r87 1 3 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=0.495 $Y=1.35
+ $X2=0.495 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HS__NAND2_4%A 3 5 7 10 12 13 16 18 20 23 26 27 28 29 30
+ 31 37
c69 37 0 1.62664e-19 $X=3.63 $Y=1.515
c70 3 0 1.84535e-19 $X=2.255 $Y=0.74
r71 41 43 14.2563 $w=3.55e-07 $l=1.05e-07 $layer=POLY_cond $X=2.61 $Y=1.557
+ $X2=2.715 $Y2=1.557
r72 41 42 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.61
+ $Y=1.515 $X2=2.61 $Y2=1.515
r73 39 41 46.1634 $w=3.55e-07 $l=3.4e-07 $layer=POLY_cond $X=2.27 $Y=1.557
+ $X2=2.61 $Y2=1.557
r74 38 39 2.03662 $w=3.55e-07 $l=1.5e-08 $layer=POLY_cond $X=2.255 $Y=1.557
+ $X2=2.27 $Y2=1.557
r75 36 37 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.63
+ $Y=1.515 $X2=3.63 $Y2=1.515
r76 31 37 0.80403 $w=4.28e-07 $l=3e-08 $layer=LI1_cond $X=3.6 $Y=1.565 $X2=3.63
+ $Y2=1.565
r77 30 31 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=3.12 $Y=1.565
+ $X2=3.6 $Y2=1.565
r78 29 30 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=2.64 $Y=1.565
+ $X2=3.12 $Y2=1.565
r79 29 42 0.80403 $w=4.28e-07 $l=3e-08 $layer=LI1_cond $X=2.64 $Y=1.565 $X2=2.61
+ $Y2=1.565
r80 27 36 7.86876 $w=3.3e-07 $l=4.5e-08 $layer=POLY_cond $X=3.675 $Y=1.515
+ $X2=3.63 $Y2=1.515
r81 27 28 5.03009 $w=3.3e-07 $l=1.08995e-07 $layer=POLY_cond $X=3.675 $Y=1.515
+ $X2=3.765 $Y2=1.557
r82 25 36 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=3.29 $Y=1.515
+ $X2=3.63 $Y2=1.515
r83 25 26 10.1687 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=3.29 $Y=1.515
+ $X2=3.215 $Y2=1.515
r84 21 28 37.0704 $w=1.5e-07 $l=2.14369e-07 $layer=POLY_cond $X=3.78 $Y=1.35
+ $X2=3.765 $Y2=1.557
r85 21 23 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=3.78 $Y=1.35
+ $X2=3.78 $Y2=0.74
r86 18 28 37.0704 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=3.765 $Y=1.765
+ $X2=3.765 $Y2=1.557
r87 18 20 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.765 $Y=1.765
+ $X2=3.765 $Y2=2.4
r88 14 26 16.9349 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.215 $Y=1.35
+ $X2=3.215 $Y2=1.515
r89 14 16 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=3.215 $Y=1.35
+ $X2=3.215 $Y2=0.74
r90 13 43 10.495 $w=3.55e-07 $l=9.3675e-08 $layer=POLY_cond $X=2.79 $Y=1.515
+ $X2=2.715 $Y2=1.557
r91 12 26 10.1687 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=3.14 $Y=1.515
+ $X2=3.215 $Y2=1.515
r92 12 13 61.2015 $w=3.3e-07 $l=3.5e-07 $layer=POLY_cond $X=3.14 $Y=1.515
+ $X2=2.79 $Y2=1.515
r93 8 43 22.9692 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.715 $Y=1.35
+ $X2=2.715 $Y2=1.557
r94 8 10 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.715 $Y=1.35
+ $X2=2.715 $Y2=0.74
r95 5 39 22.9692 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=2.27 $Y=1.765
+ $X2=2.27 $Y2=1.557
r96 5 7 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.27 $Y=1.765
+ $X2=2.27 $Y2=2.4
r97 1 38 22.9692 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.255 $Y=1.35
+ $X2=2.255 $Y2=1.557
r98 1 3 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.255 $Y=1.35
+ $X2=2.255 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HS__NAND2_4%VPWR 1 2 3 10 12 18 20 22 25 26 27 36 48
r37 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r38 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r39 42 48 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.08 $Y2=3.33
r40 41 42 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r41 38 41 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=2.16 $Y=3.33
+ $X2=3.6 $Y2=3.33
r42 36 47 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=3.875 $Y=3.33
+ $X2=4.097 $Y2=3.33
r43 36 41 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=3.875 $Y=3.33
+ $X2=3.6 $Y2=3.33
r44 34 35 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r45 32 35 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.68 $Y2=3.33
r46 32 45 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r47 31 34 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.72 $Y=3.33 $X2=1.68
+ $Y2=3.33
r48 31 32 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r49 29 44 4.73185 $w=1.7e-07 $l=2.23e-07 $layer=LI1_cond $X=0.445 $Y=3.33
+ $X2=0.222 $Y2=3.33
r50 29 31 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=0.445 $Y=3.33
+ $X2=0.72 $Y2=3.33
r51 27 42 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=3.6 $Y2=3.33
r52 27 35 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.68 $Y2=3.33
r53 27 38 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r54 26 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.995 $Y=3.33
+ $X2=2.16 $Y2=3.33
r55 25 34 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=1.83 $Y=3.33 $X2=1.68
+ $Y2=3.33
r56 25 26 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.83 $Y=3.33
+ $X2=1.995 $Y2=3.33
r57 20 47 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=4.04 $Y=3.245
+ $X2=4.097 $Y2=3.33
r58 20 22 28.8111 $w=3.28e-07 $l=8.25e-07 $layer=LI1_cond $X=4.04 $Y=3.245
+ $X2=4.04 $Y2=2.42
r59 16 26 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.995 $Y=3.245
+ $X2=1.995 $Y2=3.33
r60 16 18 28.8111 $w=3.28e-07 $l=8.25e-07 $layer=LI1_cond $X=1.995 $Y=3.245
+ $X2=1.995 $Y2=2.42
r61 12 15 27.938 $w=3.28e-07 $l=8e-07 $layer=LI1_cond $X=0.28 $Y=2.015 $X2=0.28
+ $Y2=2.815
r62 10 44 3.03433 $w=3.3e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.28 $Y=3.245
+ $X2=0.222 $Y2=3.33
r63 10 15 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=0.28 $Y=3.245
+ $X2=0.28 $Y2=2.815
r64 3 22 300 $w=1.7e-07 $l=6.72607e-07 $layer=licon1_PDIFF $count=2 $X=3.84
+ $Y=1.84 $X2=4.04 $Y2=2.42
r65 2 18 300 $w=1.7e-07 $l=6.50692e-07 $layer=licon1_PDIFF $count=2 $X=1.845
+ $Y=1.84 $X2=1.995 $Y2=2.42
r66 1 15 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.815
r67 1 12 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.015
.ends

.subckt PM_SKY130_FD_SC_HS__NAND2_4%Y 1 2 3 4 17 19 20 23 25 27 37 40 46 47 50
+ 51
r66 50 51 18.5393 $w=2.28e-07 $l=3.7e-07 $layer=LI1_cond $X=4.08 $Y=1.295
+ $X2=4.08 $Y2=1.665
r67 49 51 14.2803 $w=2.28e-07 $l=2.85e-07 $layer=LI1_cond $X=4.08 $Y=1.95
+ $X2=4.08 $Y2=1.665
r68 48 50 5.76222 $w=2.28e-07 $l=1.15e-07 $layer=LI1_cond $X=4.08 $Y=1.18
+ $X2=4.08 $Y2=1.295
r69 45 46 13.0168 $w=1.028e-06 $l=1.65e-07 $layer=LI1_cond $X=3.54 $Y=2.465
+ $X2=3.705 $Y2=2.465
r70 42 45 8.29126 $w=1.028e-06 $l=7e-07 $layer=LI1_cond $X=2.84 $Y=2.465
+ $X2=3.54 $Y2=2.465
r71 39 42 4.08641 $w=1.028e-06 $l=3.45e-07 $layer=LI1_cond $X=2.495 $Y=2.465
+ $X2=2.84 $Y2=2.465
r72 39 40 13.0168 $w=1.028e-06 $l=1.65e-07 $layer=LI1_cond $X=2.495 $Y=2.465
+ $X2=2.33 $Y2=2.465
r73 37 40 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.66 $Y=2.035
+ $X2=2.33 $Y2=2.035
r74 36 37 12.4245 $w=1.028e-06 $l=1.15e-07 $layer=LI1_cond $X=1.545 $Y=2.465
+ $X2=1.66 $Y2=2.465
r75 33 36 4.85631 $w=1.028e-06 $l=4.1e-07 $layer=LI1_cond $X=1.135 $Y=2.465
+ $X2=1.545 $Y2=2.465
r76 30 33 4.73786 $w=1.028e-06 $l=4e-07 $layer=LI1_cond $X=0.735 $Y=2.465
+ $X2=1.135 $Y2=2.465
r77 27 49 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=3.965 $Y=2.035
+ $X2=4.08 $Y2=1.95
r78 27 46 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=3.965 $Y=2.035
+ $X2=3.705 $Y2=2.035
r79 26 47 9.31531 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=3.705 $Y=1.095
+ $X2=3.52 $Y2=1.095
r80 25 48 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=3.965 $Y=1.095
+ $X2=4.08 $Y2=1.18
r81 25 26 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=3.965 $Y=1.095
+ $X2=3.705 $Y2=1.095
r82 21 47 1.24149 $w=3.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.52 $Y=1.01 $X2=3.52
+ $Y2=1.095
r83 21 23 7.0081 $w=3.68e-07 $l=2.25e-07 $layer=LI1_cond $X=3.52 $Y=1.01
+ $X2=3.52 $Y2=0.785
r84 19 47 9.31531 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=3.335 $Y=1.095
+ $X2=3.52 $Y2=1.095
r85 19 20 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.335 $Y=1.095
+ $X2=2.665 $Y2=1.095
r86 15 20 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.5 $Y=1.01
+ $X2=2.665 $Y2=1.095
r87 15 17 7.85757 $w=3.28e-07 $l=2.25e-07 $layer=LI1_cond $X=2.5 $Y=1.01 $X2=2.5
+ $Y2=0.785
r88 4 45 200 $w=1.7e-07 $l=1.47678e-06 $layer=licon1_PDIFF $count=3 $X=2.345
+ $Y=1.84 $X2=3.54 $Y2=2.47
r89 4 42 200 $w=1.7e-07 $l=1.19718e-06 $layer=licon1_PDIFF $count=3 $X=2.345
+ $Y=1.84 $X2=2.84 $Y2=2.815
r90 4 42 200 $w=1.7e-07 $l=6.17373e-07 $layer=licon1_PDIFF $count=3 $X=2.345
+ $Y=1.84 $X2=2.84 $Y2=2.115
r91 4 39 200 $w=1.7e-07 $l=7.00999e-07 $layer=licon1_PDIFF $count=3 $X=2.345
+ $Y=1.84 $X2=2.495 $Y2=2.47
r92 3 36 266.667 $w=1.7e-07 $l=1.23548e-06 $layer=licon1_PDIFF $count=2 $X=0.585
+ $Y=1.84 $X2=1.545 $Y2=2.47
r93 3 33 266.667 $w=1.7e-07 $l=1.21937e-06 $layer=licon1_PDIFF $count=2 $X=0.585
+ $Y=1.84 $X2=1.135 $Y2=2.815
r94 3 33 266.667 $w=1.7e-07 $l=6.7361e-07 $layer=licon1_PDIFF $count=2 $X=0.585
+ $Y=1.84 $X2=1.135 $Y2=2.115
r95 3 30 266.667 $w=1.7e-07 $l=7.00999e-07 $layer=licon1_PDIFF $count=2 $X=0.585
+ $Y=1.84 $X2=0.735 $Y2=2.47
r96 2 23 182 $w=1.7e-07 $l=5.17373e-07 $layer=licon1_NDIFF $count=1 $X=3.29
+ $Y=0.37 $X2=3.52 $Y2=0.785
r97 1 17 182 $w=1.7e-07 $l=4.92722e-07 $layer=licon1_NDIFF $count=1 $X=2.33
+ $Y=0.37 $X2=2.5 $Y2=0.785
.ends

.subckt PM_SKY130_FD_SC_HS__NAND2_4%A_27_74# 1 2 3 4 5 18 20 21 24 26 32 33 36
+ 38 42 44 45
r68 40 42 6.9845 $w=3.28e-07 $l=2e-07 $layer=LI1_cond $X=4.04 $Y=0.425 $X2=4.04
+ $Y2=0.625
r69 39 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.165 $Y=0.34 $X2=3
+ $Y2=0.34
r70 38 40 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.875 $Y=0.34
+ $X2=4.04 $Y2=0.425
r71 38 39 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=3.875 $Y=0.34
+ $X2=3.165 $Y2=0.34
r72 34 45 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3 $Y=0.425 $X2=3
+ $Y2=0.34
r73 34 36 6.9845 $w=3.28e-07 $l=2e-07 $layer=LI1_cond $X=3 $Y=0.425 $X2=3
+ $Y2=0.625
r74 32 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.835 $Y=0.34 $X2=3
+ $Y2=0.34
r75 32 33 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.835 $Y=0.34
+ $X2=2.165 $Y2=0.34
r76 29 31 22.8184 $w=2.48e-07 $l=4.95e-07 $layer=LI1_cond $X=2.04 $Y=1.01
+ $X2=2.04 $Y2=0.515
r77 28 33 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=2.04 $Y=0.425
+ $X2=2.165 $Y2=0.34
r78 28 31 4.14879 $w=2.48e-07 $l=9e-08 $layer=LI1_cond $X=2.04 $Y=0.425 $X2=2.04
+ $Y2=0.515
r79 27 44 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.225 $Y=1.095
+ $X2=1.14 $Y2=1.095
r80 26 29 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.915 $Y=1.095
+ $X2=2.04 $Y2=1.01
r81 26 27 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.915 $Y=1.095
+ $X2=1.225 $Y2=1.095
r82 22 44 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.14 $Y=1.01 $X2=1.14
+ $Y2=1.095
r83 22 24 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=1.14 $Y=1.01
+ $X2=1.14 $Y2=0.515
r84 20 44 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.055 $Y=1.095
+ $X2=1.14 $Y2=1.095
r85 20 21 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.055 $Y=1.095
+ $X2=0.365 $Y2=1.095
r86 16 21 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.24 $Y=1.01
+ $X2=0.365 $Y2=1.095
r87 16 18 22.8184 $w=2.48e-07 $l=4.95e-07 $layer=LI1_cond $X=0.24 $Y=1.01
+ $X2=0.24 $Y2=0.515
r88 5 42 182 $w=1.7e-07 $l=3.34963e-07 $layer=licon1_NDIFF $count=1 $X=3.855
+ $Y=0.37 $X2=4.04 $Y2=0.625
r89 4 36 182 $w=1.7e-07 $l=3.44347e-07 $layer=licon1_NDIFF $count=1 $X=2.79
+ $Y=0.37 $X2=3 $Y2=0.625
r90 3 31 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.86
+ $Y=0.37 $X2=2 $Y2=0.515
r91 2 24 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1 $Y=0.37
+ $X2=1.14 $Y2=0.515
r92 1 18 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__NAND2_4%VGND 1 2 9 13 15 17 22 29 30 33 36
c50 13 0 1.84535e-19 $X=1.57 $Y=0.625
r51 36 37 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r52 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r53 29 30 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r54 27 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.735 $Y=0 $X2=1.57
+ $Y2=0
r55 27 29 152.989 $w=1.68e-07 $l=2.345e-06 $layer=LI1_cond $X=1.735 $Y=0
+ $X2=4.08 $Y2=0
r56 26 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=1.68
+ $Y2=0
r57 26 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r58 25 26 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r59 23 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.875 $Y=0 $X2=0.71
+ $Y2=0
r60 23 25 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.875 $Y=0 $X2=1.2
+ $Y2=0
r61 22 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.405 $Y=0 $X2=1.57
+ $Y2=0
r62 22 25 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=1.405 $Y=0 $X2=1.2
+ $Y2=0
r63 20 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r64 19 20 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r65 17 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.545 $Y=0 $X2=0.71
+ $Y2=0
r66 17 19 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.545 $Y=0 $X2=0.24
+ $Y2=0
r67 15 30 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=2.16 $Y=0 $X2=4.08
+ $Y2=0
r68 15 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.68
+ $Y2=0
r69 11 36 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.57 $Y=0.085
+ $X2=1.57 $Y2=0
r70 11 13 18.8582 $w=3.28e-07 $l=5.4e-07 $layer=LI1_cond $X=1.57 $Y=0.085
+ $X2=1.57 $Y2=0.625
r71 7 33 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.71 $Y=0.085 $X2=0.71
+ $Y2=0
r72 7 9 18.8582 $w=3.28e-07 $l=5.4e-07 $layer=LI1_cond $X=0.71 $Y=0.085 $X2=0.71
+ $Y2=0.625
r73 2 13 182 $w=1.7e-07 $l=3.17372e-07 $layer=licon1_NDIFF $count=1 $X=1.43
+ $Y=0.37 $X2=1.57 $Y2=0.625
r74 1 9 182 $w=1.7e-07 $l=3.17372e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.37 $X2=0.71 $Y2=0.625
.ends

