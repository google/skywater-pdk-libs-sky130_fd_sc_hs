* File: sky130_fd_sc_hs__sdfsbp_1.pex.spice
* Created: Tue Sep  1 20:22:57 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HS__SDFSBP_1%A_27_74# 1 2 9 11 13 16 19 22 24 28 29 33
+ 36 37
c78 33 0 1.30292e-19 $X=1.96 $Y=1.995
c79 29 0 2.93935e-19 $X=0.975 $Y=1.115
c80 24 0 1.64248e-19 $X=1.795 $Y=2.375
c81 9 0 1.50564e-19 $X=1.065 $Y=0.58
r82 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.96
+ $Y=1.995 $X2=1.96 $Y2=1.995
r83 31 33 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=1.92 $Y=2.29
+ $X2=1.92 $Y2=1.995
r84 29 39 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.975 $Y=1.115
+ $X2=0.975 $Y2=0.95
r85 28 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.975
+ $Y=1.115 $X2=0.975 $Y2=1.115
r86 26 36 0.695019 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=0.445 $Y=1.115
+ $X2=0.28 $Y2=1.115
r87 26 28 18.5089 $w=3.28e-07 $l=5.3e-07 $layer=LI1_cond $X=0.445 $Y=1.115
+ $X2=0.975 $Y2=1.115
r88 25 37 2.53056 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.365 $Y=2.375
+ $X2=0.24 $Y2=2.375
r89 24 31 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.795 $Y=2.375
+ $X2=1.92 $Y2=2.29
r90 24 25 93.2941 $w=1.68e-07 $l=1.43e-06 $layer=LI1_cond $X=1.795 $Y=2.375
+ $X2=0.365 $Y2=2.375
r91 20 37 3.91525 $w=2.35e-07 $l=8.5e-08 $layer=LI1_cond $X=0.24 $Y=2.46
+ $X2=0.24 $Y2=2.375
r92 20 22 0.230489 $w=2.48e-07 $l=5e-09 $layer=LI1_cond $X=0.24 $Y=2.46 $X2=0.24
+ $Y2=2.465
r93 19 37 3.91525 $w=2.35e-07 $l=9.21954e-08 $layer=LI1_cond $X=0.225 $Y=2.29
+ $X2=0.24 $Y2=2.375
r94 18 36 5.99569 $w=2.75e-07 $l=1.90526e-07 $layer=LI1_cond $X=0.225 $Y=1.28
+ $X2=0.28 $Y2=1.115
r95 18 19 52.9076 $w=2.18e-07 $l=1.01e-06 $layer=LI1_cond $X=0.225 $Y=1.28
+ $X2=0.225 $Y2=2.29
r96 14 36 5.99569 $w=2.75e-07 $l=1.65e-07 $layer=LI1_cond $X=0.28 $Y=0.95
+ $X2=0.28 $Y2=1.115
r97 14 16 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=0.28 $Y=0.95
+ $X2=0.28 $Y2=0.58
r98 11 34 52.2586 $w=2.99e-07 $l=2.7157e-07 $layer=POLY_cond $X=2.005 $Y=2.245
+ $X2=1.96 $Y2=1.995
r99 11 13 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=2.005 $Y=2.245
+ $X2=2.005 $Y2=2.64
r100 9 39 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=1.065 $Y=0.58
+ $X2=1.065 $Y2=0.95
r101 2 22 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=2.32 $X2=0.28 $Y2=2.465
r102 1 16 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_HS__SDFSBP_1%SCE 2 5 7 9 10 12 17 19 20 23 24 28 33 39
c78 39 0 1.89796e-19 $X=0.67 $Y=1.535
c79 24 0 1.10806e-19 $X=1.96 $Y=1.425
c80 23 0 1.50331e-19 $X=1.96 $Y=1.425
r81 31 33 29.4556 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.505 $Y=1.685
+ $X2=0.67 $Y2=1.685
r82 30 31 1.78519 $w=2.7e-07 $l=1e-08 $layer=POLY_cond $X=0.495 $Y=1.685
+ $X2=0.505 $Y2=1.685
r83 28 39 4.53993 $w=3.28e-07 $l=1.3e-07 $layer=LI1_cond $X=0.67 $Y=1.665
+ $X2=0.67 $Y2=1.535
r84 28 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.67
+ $Y=1.685 $X2=0.67 $Y2=1.685
r85 24 37 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.96 $Y=1.425
+ $X2=1.96 $Y2=1.26
r86 23 26 5.07075 $w=2.48e-07 $l=1.1e-07 $layer=LI1_cond $X=1.92 $Y=1.425
+ $X2=1.92 $Y2=1.535
r87 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.96
+ $Y=1.425 $X2=1.96 $Y2=1.425
r88 21 39 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.835 $Y=1.535
+ $X2=0.67 $Y2=1.535
r89 20 26 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.795 $Y=1.535
+ $X2=1.92 $Y2=1.535
r90 20 21 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.795 $Y=1.535
+ $X2=0.835 $Y2=1.535
r91 17 37 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=1.885 $Y=0.58
+ $X2=1.885 $Y2=1.26
r92 13 33 53.5556 $w=2.7e-07 $l=3.73497e-07 $layer=POLY_cond $X=0.97 $Y=1.85
+ $X2=0.67 $Y2=1.685
r93 13 19 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=0.97 $Y=1.85
+ $X2=0.97 $Y2=2.09
r94 10 19 60.25 $w=1.8e-07 $l=1.55e-07 $layer=POLY_cond $X=0.955 $Y=2.245
+ $X2=0.955 $Y2=2.09
r95 10 12 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=0.955 $Y=2.245
+ $X2=0.955 $Y2=2.64
r96 7 9 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=0.505 $Y=2.245
+ $X2=0.505 $Y2=2.64
r97 3 30 16.5046 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.495 $Y=1.52
+ $X2=0.495 $Y2=1.685
r98 3 5 482 $w=1.5e-07 $l=9.4e-07 $layer=POLY_cond $X=0.495 $Y=1.52 $X2=0.495
+ $Y2=0.58
r99 2 7 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=0.505 $Y=2.155 $X2=0.505
+ $Y2=2.245
r100 1 31 12.2893 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=0.505 $Y=1.85
+ $X2=0.505 $Y2=1.685
r101 1 2 118.556 $w=1.8e-07 $l=3.05e-07 $layer=POLY_cond $X=0.505 $Y=1.85
+ $X2=0.505 $Y2=2.155
.ends

.subckt PM_SKY130_FD_SC_HS__SDFSBP_1%D 1 3 6 8 12
c34 1 0 2.35667e-19 $X=1.375 $Y=2.245
r35 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.42
+ $Y=1.955 $X2=1.42 $Y2=1.955
r36 8 12 7.68295 $w=3.28e-07 $l=2.2e-07 $layer=LI1_cond $X=1.2 $Y=1.955 $X2=1.42
+ $Y2=1.955
r37 4 11 38.6342 $w=2.88e-07 $l=1.81659e-07 $layer=POLY_cond $X=1.455 $Y=1.79
+ $X2=1.42 $Y2=1.955
r38 4 6 620.447 $w=1.5e-07 $l=1.21e-06 $layer=POLY_cond $X=1.455 $Y=1.79
+ $X2=1.455 $Y2=0.58
r39 1 11 59.5544 $w=2.88e-07 $l=3.11689e-07 $layer=POLY_cond $X=1.375 $Y=2.245
+ $X2=1.42 $Y2=1.955
r40 1 3 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=1.375 $Y=2.245
+ $X2=1.375 $Y2=2.64
.ends

.subckt PM_SKY130_FD_SC_HS__SDFSBP_1%SCD 1 3 4 6 7 8 9 10 11
c43 9 0 6.91441e-20 $X=2.64 $Y=1.295
c44 8 0 1.50331e-19 $X=2.597 $Y=1.918
c45 4 0 2.9454e-19 $X=2.425 $Y=2.245
r46 11 19 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=2.665
+ $Y=1.985 $X2=2.665 $Y2=1.985
r47 10 11 16.9004 $w=2.08e-07 $l=3.2e-07 $layer=LI1_cond $X=2.66 $Y=1.665
+ $X2=2.66 $Y2=1.985
r48 9 10 19.5411 $w=2.08e-07 $l=3.7e-07 $layer=LI1_cond $X=2.66 $Y=1.295
+ $X2=2.66 $Y2=1.665
r49 9 16 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=2.665
+ $Y=1.305 $X2=2.665 $Y2=1.305
r50 8 19 8.81262 $w=4.65e-07 $l=7.04131e-08 $layer=POLY_cond $X=2.597 $Y=1.918
+ $X2=2.59 $Y2=1.985
r51 7 16 10.4119 $w=4.65e-07 $l=1.10535e-07 $layer=POLY_cond $X=2.597 $Y=1.372
+ $X2=2.515 $Y2=1.305
r52 7 8 65.3032 $w=4.65e-07 $l=5.46e-07 $layer=POLY_cond $X=2.597 $Y=1.372
+ $X2=2.597 $Y2=1.918
r53 4 19 51.3137 $w=3.77e-07 $l=3.32415e-07 $layer=POLY_cond $X=2.425 $Y=2.245
+ $X2=2.59 $Y2=1.985
r54 4 6 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=2.425 $Y=2.245
+ $X2=2.425 $Y2=2.64
r55 1 16 77.4558 $w=3.42e-07 $l=5.46992e-07 $layer=POLY_cond $X=2.275 $Y=0.865
+ $X2=2.515 $Y2=1.305
r56 1 3 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=2.275 $Y=0.865
+ $X2=2.275 $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_HS__SDFSBP_1%CLK 1 3 4 6 7
c32 4 0 6.91441e-20 $X=3.515 $Y=1.765
c33 1 0 9.27061e-20 $X=3.33 $Y=1.22
r34 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.38
+ $Y=1.385 $X2=3.38 $Y2=1.385
r35 7 11 6.85236 $w=3.68e-07 $l=2.2e-07 $layer=LI1_cond $X=3.6 $Y=1.365 $X2=3.38
+ $Y2=1.365
r36 4 10 76.492 $w=2.75e-07 $l=4.29302e-07 $layer=POLY_cond $X=3.515 $Y=1.765
+ $X2=3.41 $Y2=1.385
r37 4 6 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.515 $Y=1.765
+ $X2=3.515 $Y2=2.4
r38 1 10 38.8084 $w=2.75e-07 $l=2.0106e-07 $layer=POLY_cond $X=3.33 $Y=1.22
+ $X2=3.41 $Y2=1.385
r39 1 3 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=3.33 $Y=1.22 $X2=3.33
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HS__SDFSBP_1%A_781_74# 1 2 7 9 14 18 22 25 29 31 32 33
+ 34 35 37 42 43 44 47 48 49 51 52 53 55 56 59 62 63 69 74
c210 74 0 1.55309e-19 $X=8.825 $Y=1.795
c211 55 0 3.2241e-19 $X=8.745 $Y=1.95
c212 51 0 1.38387e-19 $X=7.36 $Y=2.905
c213 32 0 9.27061e-20 $X=4.21 $Y=0.34
r214 68 69 30.474 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=5.5 $Y=1.855
+ $X2=5.425 $Y2=1.855
r215 63 74 66.3205 $w=3.3e-07 $l=2.8e-07 $layer=POLY_cond $X=8.825 $Y=1.515
+ $X2=8.825 $Y2=1.795
r216 63 73 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=8.825 $Y=1.515
+ $X2=8.825 $Y2=1.35
r217 62 65 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=8.825 $Y=1.515
+ $X2=8.825 $Y2=1.68
r218 62 63 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.825
+ $Y=1.515 $X2=8.825 $Y2=1.515
r219 59 68 25.3549 $w=3.3e-07 $l=1.45e-07 $layer=POLY_cond $X=5.645 $Y=1.855
+ $X2=5.5 $Y2=1.855
r220 58 60 16.8553 $w=2.28e-07 $l=3.15e-07 $layer=LI1_cond $X=5.675 $Y=1.855
+ $X2=5.675 $Y2=2.17
r221 58 59 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.645
+ $Y=1.855 $X2=5.645 $Y2=1.855
r222 55 65 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=8.745 $Y=1.95
+ $X2=8.745 $Y2=1.68
r223 52 55 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.66 $Y=2.035
+ $X2=8.745 $Y2=1.95
r224 52 53 79.2674 $w=1.68e-07 $l=1.215e-06 $layer=LI1_cond $X=8.66 $Y=2.035
+ $X2=7.445 $Y2=2.035
r225 50 53 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.36 $Y=2.12
+ $X2=7.445 $Y2=2.035
r226 50 51 51.2139 $w=1.68e-07 $l=7.85e-07 $layer=LI1_cond $X=7.36 $Y=2.12
+ $X2=7.36 $Y2=2.905
r227 48 51 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.275 $Y=2.99
+ $X2=7.36 $Y2=2.905
r228 48 49 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=7.275 $Y=2.99
+ $X2=6.765 $Y2=2.99
r229 47 49 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.68 $Y=2.905
+ $X2=6.765 $Y2=2.99
r230 46 47 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=6.68 $Y=2.255
+ $X2=6.68 $Y2=2.905
r231 45 60 2.45823 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=5.81 $Y=2.17
+ $X2=5.675 $Y2=2.17
r232 44 46 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.595 $Y=2.17
+ $X2=6.68 $Y2=2.255
r233 44 45 51.2139 $w=1.68e-07 $l=7.85e-07 $layer=LI1_cond $X=6.595 $Y=2.17
+ $X2=5.81 $Y2=2.17
r234 42 60 5.36411 $w=2.28e-07 $l=1.07121e-07 $layer=LI1_cond $X=5.725 $Y=2.255
+ $X2=5.675 $Y2=2.17
r235 42 43 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=5.725 $Y=2.255
+ $X2=5.725 $Y2=2.905
r236 40 56 61.6524 $w=1.68e-07 $l=9.45e-07 $layer=LI1_cond $X=4.945 $Y=0.425
+ $X2=4.945 $Y2=1.37
r237 38 67 37.5797 $w=2.95e-07 $l=2.3e-07 $layer=POLY_cond $X=4.925 $Y=1.535
+ $X2=4.925 $Y2=1.765
r238 37 38 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.925
+ $Y=1.535 $X2=4.925 $Y2=1.535
r239 35 56 7.33542 $w=2.68e-07 $l=1.35e-07 $layer=LI1_cond $X=4.895 $Y=1.505
+ $X2=4.895 $Y2=1.37
r240 35 37 1.28049 $w=2.68e-07 $l=3e-08 $layer=LI1_cond $X=4.895 $Y=1.505
+ $X2=4.895 $Y2=1.535
r241 33 43 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.64 $Y=2.99
+ $X2=5.725 $Y2=2.905
r242 33 34 83.8342 $w=1.68e-07 $l=1.285e-06 $layer=LI1_cond $X=5.64 $Y=2.99
+ $X2=4.355 $Y2=2.99
r243 31 40 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.86 $Y=0.34
+ $X2=4.945 $Y2=0.425
r244 31 32 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=4.86 $Y=0.34
+ $X2=4.21 $Y2=0.34
r245 27 34 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=4.23 $Y=2.905
+ $X2=4.355 $Y2=2.99
r246 27 29 6.45368 $w=2.48e-07 $l=1.4e-07 $layer=LI1_cond $X=4.23 $Y=2.905
+ $X2=4.23 $Y2=2.765
r247 23 32 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.045 $Y=0.425
+ $X2=4.21 $Y2=0.34
r248 23 25 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=4.045 $Y=0.425
+ $X2=4.045 $Y2=0.505
r249 22 74 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=8.9 $Y=2.08 $X2=8.9
+ $Y2=1.795
r250 18 73 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=8.735 $Y=0.69
+ $X2=8.735 $Y2=1.35
r251 12 68 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.5 $Y=1.69
+ $X2=5.5 $Y2=1.855
r252 12 14 569.17 $w=1.5e-07 $l=1.11e-06 $layer=POLY_cond $X=5.5 $Y=1.69 $X2=5.5
+ $Y2=0.58
r253 11 67 18.5736 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.09 $Y=1.765
+ $X2=4.925 $Y2=1.765
r254 11 69 171.777 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=5.09 $Y=1.765
+ $X2=5.425 $Y2=1.765
r255 7 67 89.2288 $w=2.95e-07 $l=5.04108e-07 $layer=POLY_cond $X=4.985 $Y=2.24
+ $X2=4.925 $Y2=1.765
r256 7 9 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=4.985 $Y=2.24
+ $X2=4.985 $Y2=2.525
r257 2 29 600 $w=1.7e-07 $l=9.97184e-07 $layer=licon1_PDIFF $count=1 $X=4.04
+ $Y=1.84 $X2=4.19 $Y2=2.765
r258 1 25 91 $w=1.7e-07 $l=1.96214e-07 $layer=licon1_NDIFF $count=2 $X=3.905
+ $Y=0.37 $X2=4.045 $Y2=0.505
.ends

.subckt PM_SKY130_FD_SC_HS__SDFSBP_1%A_1163_48# 1 2 7 9 10 11 12 14 16 17 19 26
+ 33
c75 12 0 6.11079e-20 $X=6.11 $Y=2.24
r76 35 37 41.0924 $w=3.3e-07 $l=2.35e-07 $layer=POLY_cond $X=5.89 $Y=1.065
+ $X2=6.125 $Y2=1.065
r77 33 37 34.0979 $w=3.3e-07 $l=1.95e-07 $layer=POLY_cond $X=6.32 $Y=1.065
+ $X2=6.125 $Y2=1.065
r78 32 33 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.32
+ $Y=1.065 $X2=6.32 $Y2=1.065
r79 24 26 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=7.02 $Y=1.915 $X2=7.02
+ $Y2=2.515
r80 21 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.215
+ $Y=1.8 $X2=6.215 $Y2=1.8
r81 19 24 6.9898 $w=2.25e-07 $l=1.49579e-07 $layer=LI1_cond $X=6.935 $Y=1.802
+ $X2=7.02 $Y2=1.915
r82 19 21 36.8782 $w=2.23e-07 $l=7.2e-07 $layer=LI1_cond $X=6.935 $Y=1.802
+ $X2=6.215 $Y2=1.802
r83 17 32 3.99273 $w=3.3e-07 $l=1.33492e-07 $layer=LI1_cond $X=6.263 $Y=0.957
+ $X2=6.32 $Y2=1.065
r84 17 29 15.4164 $w=3.3e-07 $l=6.79219e-07 $layer=LI1_cond $X=6.263 $Y=0.957
+ $X2=6.765 $Y2=0.54
r85 16 22 38.7084 $w=3.43e-07 $l=1.98997e-07 $layer=POLY_cond $X=6.125 $Y=1.635
+ $X2=6.2 $Y2=1.8
r86 15 37 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.125 $Y=1.23
+ $X2=6.125 $Y2=1.065
r87 15 16 207.67 $w=1.5e-07 $l=4.05e-07 $layer=POLY_cond $X=6.125 $Y=1.23
+ $X2=6.125 $Y2=1.635
r88 12 14 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=6.11 $Y=2.24 $X2=6.11
+ $Y2=2.525
r89 11 12 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=6.11 $Y=2.15 $X2=6.11
+ $Y2=2.24
r90 10 22 34.0194 $w=3.43e-07 $l=2.05122e-07 $layer=POLY_cond $X=6.11 $Y=1.965
+ $X2=6.2 $Y2=1.8
r91 10 11 71.9113 $w=1.8e-07 $l=1.85e-07 $layer=POLY_cond $X=6.11 $Y=1.965
+ $X2=6.11 $Y2=2.15
r92 7 35 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.89 $Y=0.9 $X2=5.89
+ $Y2=1.065
r93 7 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=5.89 $Y=0.9 $X2=5.89
+ $Y2=0.58
r94 2 26 600 $w=1.7e-07 $l=2.64575e-07 $layer=licon1_PDIFF $count=1 $X=6.87
+ $Y=2.315 $X2=7.02 $Y2=2.515
r95 1 29 182 $w=1.7e-07 $l=2.31409e-07 $layer=licon1_NDIFF $count=1 $X=6.62
+ $Y=0.37 $X2=6.765 $Y2=0.54
.ends

.subckt PM_SKY130_FD_SC_HS__SDFSBP_1%A_995_74# 1 2 7 8 9 11 14 16 18 19 21 24 27
+ 28 30 34 35 38 40 43
c137 27 0 6.11079e-20 $X=5.285 $Y=2.37
c138 8 0 1.19047e-19 $X=6.795 $Y=2.15
r139 43 45 3.42456 $w=2.85e-07 $l=8e-08 $layer=LI1_cond $X=6.917 $Y=1.355
+ $X2=6.917 $Y2=1.435
r140 43 44 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.89
+ $Y=1.355 $X2=6.89 $Y2=1.355
r141 35 49 42.2056 $w=3.94e-07 $l=3.45e-07 $layer=POLY_cond $X=8 $Y=1.39
+ $X2=8.345 $Y2=1.39
r142 35 47 9.17513 $w=3.94e-07 $l=7.5e-08 $layer=POLY_cond $X=8 $Y=1.39
+ $X2=7.925 $Y2=1.39
r143 34 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8
+ $Y=1.285 $X2=8 $Y2=1.285
r144 32 34 7.33373 $w=3.28e-07 $l=2.1e-07 $layer=LI1_cond $X=8 $Y=1.075 $X2=8
+ $Y2=1.285
r145 31 43 15.6246 $w=2.85e-07 $l=4.51298e-07 $layer=LI1_cond $X=7.11 $Y=0.99
+ $X2=6.917 $Y2=1.355
r146 30 32 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=7.835 $Y=0.99
+ $X2=8 $Y2=1.075
r147 30 31 47.2995 $w=1.68e-07 $l=7.25e-07 $layer=LI1_cond $X=7.835 $Y=0.99
+ $X2=7.11 $Y2=0.99
r148 29 40 2.11342 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.45 $Y=1.435
+ $X2=5.325 $Y2=1.435
r149 28 45 3.76007 $w=1.7e-07 $l=1.92e-07 $layer=LI1_cond $X=6.725 $Y=1.435
+ $X2=6.917 $Y2=1.435
r150 28 29 83.1818 $w=1.68e-07 $l=1.275e-06 $layer=LI1_cond $X=6.725 $Y=1.435
+ $X2=5.45 $Y2=1.435
r151 27 38 8.98601 $w=3.28e-07 $l=1.8e-07 $layer=LI1_cond $X=5.285 $Y=2.37
+ $X2=5.285 $Y2=2.55
r152 26 40 4.3182 $w=2.1e-07 $l=1.03078e-07 $layer=LI1_cond $X=5.285 $Y=1.52
+ $X2=5.325 $Y2=1.435
r153 26 27 55.4545 $w=1.68e-07 $l=8.5e-07 $layer=LI1_cond $X=5.285 $Y=1.52
+ $X2=5.285 $Y2=2.37
r154 22 40 4.3182 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=5.325 $Y=1.35
+ $X2=5.325 $Y2=1.435
r155 22 24 35.4952 $w=2.48e-07 $l=7.7e-07 $layer=LI1_cond $X=5.325 $Y=1.35
+ $X2=5.325 $Y2=0.58
r156 19 49 25.4929 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=8.345 $Y=1.12
+ $X2=8.345 $Y2=1.39
r157 19 21 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=8.345 $Y=1.12
+ $X2=8.345 $Y2=0.69
r158 16 47 25.4929 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=7.925 $Y=1.66
+ $X2=7.925 $Y2=1.39
r159 16 18 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=7.925 $Y=1.66
+ $X2=7.925 $Y2=2.235
r160 12 44 38.5662 $w=2.97e-07 $l=2.09105e-07 $layer=POLY_cond $X=6.98 $Y=1.19
+ $X2=6.88 $Y2=1.355
r161 12 14 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=6.98 $Y=1.19
+ $X2=6.98 $Y2=0.58
r162 9 11 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=6.795 $Y=2.24
+ $X2=6.795 $Y2=2.525
r163 8 9 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=6.795 $Y=2.15 $X2=6.795
+ $Y2=2.24
r164 7 44 48.8089 $w=2.97e-07 $l=2.94449e-07 $layer=POLY_cond $X=6.795 $Y=1.61
+ $X2=6.88 $Y2=1.355
r165 7 8 209.903 $w=1.8e-07 $l=5.4e-07 $layer=POLY_cond $X=6.795 $Y=1.61
+ $X2=6.795 $Y2=2.15
r166 2 38 600 $w=1.7e-07 $l=3.28786e-07 $layer=licon1_PDIFF $count=1 $X=5.06
+ $Y=2.315 $X2=5.285 $Y2=2.55
r167 1 24 182 $w=1.7e-07 $l=4.01497e-07 $layer=licon1_NDIFF $count=1 $X=4.975
+ $Y=0.37 $X2=5.285 $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_HS__SDFSBP_1%SET_B 3 6 7 9 10 12 13 14 20 21 23 24 25 27
+ 28 31 33 34 39 42 43 47
c156 43 0 1.19047e-19 $X=7.46 $Y=1.41
c157 28 0 1.8354e-19 $X=10.75 $Y=1.42
c158 14 0 7.13225e-20 $X=10.31 $Y=0.94
c159 13 0 1.94471e-19 $X=10.55 $Y=0.94
c160 7 0 2.22931e-19 $X=7.385 $Y=2.24
r161 42 45 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=7.46 $Y=1.41
+ $X2=7.46 $Y2=1.575
r162 42 44 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=7.46 $Y=1.41
+ $X2=7.46 $Y2=1.245
r163 42 43 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.46
+ $Y=1.41 $X2=7.46 $Y2=1.41
r164 39 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.84 $Y=1.665
+ $X2=9.84 $Y2=1.665
r165 37 43 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=7.46 $Y=1.665
+ $X2=7.46 $Y2=1.41
r166 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=1.665
+ $X2=7.44 $Y2=1.665
r167 34 36 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=7.585 $Y=1.665
+ $X2=7.44 $Y2=1.665
r168 33 39 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=9.695 $Y=1.665
+ $X2=9.84 $Y2=1.665
r169 33 34 2.61138 $w=1.4e-07 $l=2.11e-06 $layer=MET1_cond $X=9.695 $Y=1.665
+ $X2=7.585 $Y2=1.665
r170 31 53 37.3291 $w=2.28e-07 $l=7.45e-07 $layer=LI1_cond $X=10.585 $Y=1.665
+ $X2=9.84 $Y2=1.665
r171 30 31 2.85155 $w=2.3e-07 $l=1.65e-07 $layer=LI1_cond $X=10.75 $Y=1.665
+ $X2=10.585 $Y2=1.665
r172 28 47 45.6753 $w=4e-07 $l=1.65e-07 $layer=POLY_cond $X=10.75 $Y=1.42
+ $X2=10.75 $Y2=1.255
r173 27 30 8.55602 $w=3.28e-07 $l=2.45e-07 $layer=LI1_cond $X=10.75 $Y=1.42
+ $X2=10.75 $Y2=1.665
r174 27 28 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=10.75
+ $Y=1.42 $X2=10.75 $Y2=1.42
r175 24 25 37.8919 $w=4e-07 $l=1.5e-07 $layer=POLY_cond $X=10.765 $Y=1.775
+ $X2=10.765 $Y2=1.925
r176 21 23 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=10.89 $Y=2.465
+ $X2=10.89 $Y2=2.75
r177 20 21 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=10.89 $Y=2.375
+ $X2=10.89 $Y2=2.465
r178 20 25 174.919 $w=1.8e-07 $l=4.5e-07 $layer=POLY_cond $X=10.89 $Y=2.375
+ $X2=10.89 $Y2=1.925
r179 17 28 4.86635 $w=4e-07 $l=3.5e-08 $layer=POLY_cond $X=10.75 $Y=1.455
+ $X2=10.75 $Y2=1.42
r180 17 24 44.4923 $w=4e-07 $l=3.2e-07 $layer=POLY_cond $X=10.75 $Y=1.455
+ $X2=10.75 $Y2=1.775
r181 15 47 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=10.625 $Y=1.015
+ $X2=10.625 $Y2=1.255
r182 13 15 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=10.55 $Y=0.94
+ $X2=10.625 $Y2=1.015
r183 13 14 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=10.55 $Y=0.94
+ $X2=10.31 $Y2=0.94
r184 10 14 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=10.235 $Y=0.865
+ $X2=10.31 $Y2=0.94
r185 10 12 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=10.235 $Y=0.865
+ $X2=10.235 $Y2=0.58
r186 7 9 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=7.385 $Y=2.24
+ $X2=7.385 $Y2=2.525
r187 6 7 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=7.385 $Y=2.15 $X2=7.385
+ $Y2=2.24
r188 6 45 223.508 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=7.385 $Y=2.15
+ $X2=7.385 $Y2=1.575
r189 3 44 340.989 $w=1.5e-07 $l=6.65e-07 $layer=POLY_cond $X=7.37 $Y=0.58
+ $X2=7.37 $Y2=1.245
.ends

.subckt PM_SKY130_FD_SC_HS__SDFSBP_1%A_594_74# 1 2 7 9 10 12 13 16 17 19 20 23
+ 25 27 28 32 37 38 41 45 47 51 54 56 57 61 64 66 67
c180 57 0 2.88662e-20 $X=3.885 $Y=1.905
c181 45 0 1.51361e-19 $X=9.44 $Y=1.72
c182 37 0 1.7105e-19 $X=9.44 $Y=2.37
c183 16 0 1.84863e-19 $X=4.475 $Y=3.075
r184 66 67 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=3.29 $Y=1.985
+ $X2=3.455 $Y2=1.985
r185 61 62 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.05
+ $Y=1.385 $X2=4.05 $Y2=1.385
r186 59 61 15.1913 $w=3.28e-07 $l=4.35e-07 $layer=LI1_cond $X=4.05 $Y=1.82
+ $X2=4.05 $Y2=1.385
r187 57 59 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.885 $Y=1.905
+ $X2=4.05 $Y2=1.82
r188 57 67 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=3.885 $Y=1.905
+ $X2=3.455 $Y2=1.905
r189 56 66 6.46067 $w=3.28e-07 $l=1.85e-07 $layer=LI1_cond $X=3.105 $Y=1.985
+ $X2=3.29 $Y2=1.985
r190 54 56 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.02 $Y=1.82
+ $X2=3.105 $Y2=1.985
r191 54 64 52.8449 $w=1.68e-07 $l=8.1e-07 $layer=LI1_cond $X=3.02 $Y=1.82
+ $X2=3.02 $Y2=1.01
r192 49 64 7.21712 $w=2.63e-07 $l=1.32e-07 $layer=LI1_cond $X=3.067 $Y=0.878
+ $X2=3.067 $Y2=1.01
r193 49 51 16.2212 $w=2.63e-07 $l=3.73e-07 $layer=LI1_cond $X=3.067 $Y=0.878
+ $X2=3.067 $Y2=0.505
r194 43 45 69.2234 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=9.305 $Y=1.72
+ $X2=9.44 $Y2=1.72
r195 35 47 81.8353 $w=1.8e-07 $l=2.05e-07 $layer=POLY_cond $X=9.44 $Y=2.945
+ $X2=9.44 $Y2=3.15
r196 35 37 294.84 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=9.44 $Y=2.945
+ $X2=9.44 $Y2=2.37
r197 34 45 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=9.44 $Y=1.795
+ $X2=9.44 $Y2=1.72
r198 34 37 294.84 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=9.44 $Y=1.795
+ $X2=9.44 $Y2=2.37
r199 30 43 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=9.305 $Y=1.645
+ $X2=9.305 $Y2=1.72
r200 30 32 546.096 $w=1.5e-07 $l=1.065e-06 $layer=POLY_cond $X=9.305 $Y=1.645
+ $X2=9.305 $Y2=0.58
r201 29 41 7.1379 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=5.68 $Y=3.15 $X2=5.59
+ $Y2=3.15
r202 28 47 7.1379 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=9.35 $Y=3.15 $X2=9.44
+ $Y2=3.15
r203 28 29 1881.85 $w=1.5e-07 $l=3.67e-06 $layer=POLY_cond $X=9.35 $Y=3.15
+ $X2=5.68 $Y2=3.15
r204 25 41 105.158 $w=1.8e-07 $l=2.65e-07 $layer=POLY_cond $X=5.59 $Y=2.885
+ $X2=5.59 $Y2=3.15
r205 25 27 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=5.59 $Y=2.885
+ $X2=5.59 $Y2=2.6
r206 21 23 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=4.9 $Y=0.98 $X2=4.9
+ $Y2=0.58
r207 19 41 7.1379 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=5.5 $Y=3.15 $X2=5.59
+ $Y2=3.15
r208 19 20 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=5.5 $Y=3.15
+ $X2=4.55 $Y2=3.15
r209 18 38 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.55 $Y=1.055
+ $X2=4.475 $Y2=1.055
r210 17 21 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.825 $Y=1.055
+ $X2=4.9 $Y2=0.98
r211 17 18 141.011 $w=1.5e-07 $l=2.75e-07 $layer=POLY_cond $X=4.825 $Y=1.055
+ $X2=4.55 $Y2=1.055
r212 16 20 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.475 $Y=3.075
+ $X2=4.55 $Y2=3.15
r213 15 16 781.968 $w=1.5e-07 $l=1.525e-06 $layer=POLY_cond $X=4.475 $Y=1.55
+ $X2=4.475 $Y2=3.075
r214 13 15 84.6064 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.475 $Y=1.385
+ $X2=4.475 $Y2=1.55
r215 13 38 169.213 $w=1.5e-07 $l=3.3e-07 $layer=POLY_cond $X=4.475 $Y=1.385
+ $X2=4.475 $Y2=1.055
r216 13 62 60.3271 $w=3.3e-07 $l=3.45e-07 $layer=POLY_cond $X=4.4 $Y=1.385
+ $X2=4.055 $Y2=1.385
r217 10 62 90.2669 $w=2.13e-07 $l=4.08901e-07 $layer=POLY_cond $X=3.965 $Y=1.765
+ $X2=3.905 $Y2=1.385
r218 10 12 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.965 $Y=1.765
+ $X2=3.965 $Y2=2.4
r219 7 62 41.6143 $w=2.13e-07 $l=1.98997e-07 $layer=POLY_cond $X=3.83 $Y=1.22
+ $X2=3.905 $Y2=1.385
r220 7 9 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=3.83 $Y=1.22 $X2=3.83
+ $Y2=0.74
r221 2 66 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=3.15
+ $Y=1.84 $X2=3.29 $Y2=1.985
r222 1 51 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=2.97
+ $Y=0.37 $X2=3.115 $Y2=0.505
.ends

.subckt PM_SKY130_FD_SC_HS__SDFSBP_1%A_1924_48# 1 2 9 11 12 13 14 16 17 18 21 22
+ 24 28 31 32 33 36 38 39 41 42 46 48
c136 42 0 7.13225e-20 $X=9.785 $Y=0.985
c137 31 0 1.8354e-19 $X=11.31 $Y=1.3
c138 28 0 1.94471e-19 $X=11.23 $Y=0.58
r139 45 46 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.785
+ $Y=1.065 $X2=9.785 $Y2=1.065
r140 42 45 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=9.785 $Y=0.985
+ $X2=9.785 $Y2=1.065
r141 40 41 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=12.15 $Y=1.47
+ $X2=12.15 $Y2=2.18
r142 38 41 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=12.065 $Y=2.265
+ $X2=12.15 $Y2=2.18
r143 38 39 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=12.065 $Y=2.265
+ $X2=11.75 $Y2=2.265
r144 34 39 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=11.625 $Y=2.35
+ $X2=11.75 $Y2=2.265
r145 34 36 18.4391 $w=2.48e-07 $l=4e-07 $layer=LI1_cond $X=11.625 $Y=2.35
+ $X2=11.625 $Y2=2.75
r146 32 40 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=12.065 $Y=1.385
+ $X2=12.15 $Y2=1.47
r147 32 33 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=12.065 $Y=1.385
+ $X2=11.395 $Y2=1.385
r148 31 33 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=11.31 $Y=1.3
+ $X2=11.395 $Y2=1.385
r149 30 48 3.70735 $w=2.5e-07 $l=1.18427e-07 $layer=LI1_cond $X=11.31 $Y=1.07
+ $X2=11.23 $Y2=0.985
r150 30 31 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=11.31 $Y=1.07
+ $X2=11.31 $Y2=1.3
r151 26 48 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=11.23 $Y=0.9
+ $X2=11.23 $Y2=0.985
r152 26 28 11.1752 $w=3.28e-07 $l=3.2e-07 $layer=LI1_cond $X=11.23 $Y=0.9
+ $X2=11.23 $Y2=0.58
r153 25 42 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.95 $Y=0.985
+ $X2=9.785 $Y2=0.985
r154 24 48 2.76166 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.065 $Y=0.985
+ $X2=11.23 $Y2=0.985
r155 24 25 72.7433 $w=1.68e-07 $l=1.115e-06 $layer=LI1_cond $X=11.065 $Y=0.985
+ $X2=9.95 $Y2=0.985
r156 20 46 33.2236 $w=3.3e-07 $l=1.9e-07 $layer=POLY_cond $X=9.785 $Y=1.255
+ $X2=9.785 $Y2=1.065
r157 20 21 43.5886 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=9.825 $Y=1.255
+ $X2=9.825 $Y2=1.405
r158 17 46 6.12014 $w=3.3e-07 $l=3.5e-08 $layer=POLY_cond $X=9.785 $Y=1.03
+ $X2=9.785 $Y2=1.065
r159 17 18 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=9.785 $Y=1.03
+ $X2=9.785 $Y2=0.865
r160 14 22 89.6095 $w=1.8e-07 $l=2.25e-07 $layer=POLY_cond $X=10.44 $Y=2.465
+ $X2=10.44 $Y2=2.24
r161 14 16 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=10.44 $Y=2.465
+ $X2=10.44 $Y2=2.75
r162 12 22 7.1379 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=10.35 $Y=2.24
+ $X2=10.44 $Y2=2.24
r163 12 13 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=10.35 $Y=2.24
+ $X2=10.03 $Y2=2.24
r164 11 13 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=9.955 $Y=2.165
+ $X2=10.03 $Y2=2.24
r165 11 21 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=9.955 $Y=2.165
+ $X2=9.955 $Y2=1.405
r166 9 18 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=9.695 $Y=0.58
+ $X2=9.695 $Y2=0.865
r167 2 36 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=11.525
+ $Y=2.54 $X2=11.665 $Y2=2.75
r168 1 28 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=11.09
+ $Y=0.37 $X2=11.23 $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_HS__SDFSBP_1%A_1762_74# 1 2 3 10 12 14 16 17 19 22 24 25
+ 26 28 29 33 35 37 40 42 43 46 47 51 53 57 59 63 67 68 71 76 77
c194 68 0 3.56881e-20 $X=9.212 $Y=1.85
c195 47 0 1.92388e-19 $X=13.14 $Y=1.79
r196 76 77 10.7321 $w=3.28e-07 $l=2.3e-07 $layer=LI1_cond $X=11.115 $Y=2.75
+ $X2=11.115 $Y2=2.52
r197 71 73 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=10.085 $Y=2.035
+ $X2=10.085 $Y2=2.18
r198 67 69 0.688026 $w=3.33e-07 $l=2e-08 $layer=LI1_cond $X=9.212 $Y=2.015
+ $X2=9.212 $Y2=2.035
r199 67 68 8.46614 $w=3.33e-07 $l=1.65e-07 $layer=LI1_cond $X=9.212 $Y=2.015
+ $X2=9.212 $Y2=1.85
r200 65 68 52.1925 $w=1.68e-07 $l=8e-07 $layer=LI1_cond $X=9.295 $Y=1.05
+ $X2=9.295 $Y2=1.85
r201 63 65 17.5613 $w=5.93e-07 $l=5.35e-07 $layer=LI1_cond $X=9.082 $Y=0.515
+ $X2=9.082 $Y2=1.05
r202 59 60 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=11.73
+ $Y=1.805 $X2=11.73 $Y2=1.805
r203 57 81 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=11.195 $Y=1.805
+ $X2=11.195 $Y2=2.18
r204 57 59 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=11.28 $Y=1.805
+ $X2=11.73 $Y2=1.805
r205 55 81 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=11.195 $Y=2.265
+ $X2=11.195 $Y2=2.18
r206 55 77 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=11.195 $Y=2.265
+ $X2=11.195 $Y2=2.52
r207 54 73 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.17 $Y=2.18
+ $X2=10.085 $Y2=2.18
r208 53 81 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=11.11 $Y=2.18
+ $X2=11.195 $Y2=2.18
r209 53 54 61.3262 $w=1.68e-07 $l=9.4e-07 $layer=LI1_cond $X=11.11 $Y=2.18
+ $X2=10.17 $Y2=2.18
r210 52 69 4.71304 $w=1.7e-07 $l=1.68e-07 $layer=LI1_cond $X=9.38 $Y=2.035
+ $X2=9.212 $Y2=2.035
r211 51 71 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10 $Y=2.035
+ $X2=10.085 $Y2=2.035
r212 51 52 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=10 $Y=2.035
+ $X2=9.38 $Y2=2.035
r213 47 48 57.9764 $w=2.12e-07 $l=2.55e-07 $layer=POLY_cond $X=13.14 $Y=1.79
+ $X2=13.395 $Y2=1.79
r214 43 60 11.3783 $w=3.55e-07 $l=7e-08 $layer=POLY_cond $X=11.8 $Y=1.792
+ $X2=11.73 $Y2=1.792
r215 43 44 13.5596 $w=3.55e-07 $l=1.30457e-07 $layer=POLY_cond $X=11.8 $Y=1.792
+ $X2=11.89 $Y2=1.885
r216 42 60 57.7042 $w=3.55e-07 $l=3.55e-07 $layer=POLY_cond $X=11.375 $Y=1.792
+ $X2=11.73 $Y2=1.792
r217 38 40 146.138 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=11.015 $Y=0.94
+ $X2=11.3 $Y2=0.94
r218 35 48 10.9192 $w=1.5e-07 $l=1.5e-07 $layer=POLY_cond $X=13.395 $Y=1.94
+ $X2=13.395 $Y2=1.79
r219 35 37 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=13.395 $Y=1.94
+ $X2=13.395 $Y2=2.435
r220 31 47 10.9192 $w=1.5e-07 $l=1.75e-07 $layer=POLY_cond $X=13.14 $Y=1.615
+ $X2=13.14 $Y2=1.79
r221 31 33 423.032 $w=1.5e-07 $l=8.25e-07 $layer=POLY_cond $X=13.14 $Y=1.615
+ $X2=13.14 $Y2=0.79
r222 30 46 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=12.47 $Y=1.69
+ $X2=12.395 $Y2=1.69
r223 29 47 21.2379 $w=2.12e-07 $l=1.32288e-07 $layer=POLY_cond $X=13.065 $Y=1.69
+ $X2=13.14 $Y2=1.79
r224 29 30 305.096 $w=1.5e-07 $l=5.95e-07 $layer=POLY_cond $X=13.065 $Y=1.69
+ $X2=12.47 $Y2=1.69
r225 26 46 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=12.395 $Y=1.765
+ $X2=12.395 $Y2=1.69
r226 26 28 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=12.395 $Y=1.765
+ $X2=12.395 $Y2=2.4
r227 24 46 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=12.32 $Y=1.69
+ $X2=12.395 $Y2=1.69
r228 24 25 87.1702 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=12.32 $Y=1.69
+ $X2=12.15 $Y2=1.69
r229 20 25 24.0479 $w=2.99e-07 $l=1.06066e-07 $layer=POLY_cond $X=12.075
+ $Y=1.615 $X2=12.15 $Y2=1.69
r230 20 44 29.8227 $w=2.99e-07 $l=3.505e-07 $layer=POLY_cond $X=12.075 $Y=1.615
+ $X2=11.89 $Y2=1.885
r231 20 22 448.67 $w=1.5e-07 $l=8.75e-07 $layer=POLY_cond $X=12.075 $Y=1.615
+ $X2=12.075 $Y2=0.74
r232 17 19 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=11.89 $Y=2.465
+ $X2=11.89 $Y2=2.75
r233 16 17 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=11.89 $Y=2.375
+ $X2=11.89 $Y2=2.465
r234 15 44 14.6425 $w=1.8e-07 $l=2.1e-07 $layer=POLY_cond $X=11.89 $Y=2.095
+ $X2=11.89 $Y2=1.885
r235 15 16 108.839 $w=1.8e-07 $l=2.8e-07 $layer=POLY_cond $X=11.89 $Y=2.095
+ $X2=11.89 $Y2=2.375
r236 14 42 33.1523 $w=3.55e-07 $l=2.11197e-07 $layer=POLY_cond $X=11.3 $Y=1.615
+ $X2=11.375 $Y2=1.792
r237 13 40 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=11.3 $Y=1.015
+ $X2=11.3 $Y2=0.94
r238 13 14 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=11.3 $Y=1.015 $X2=11.3
+ $Y2=1.615
r239 10 38 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=11.015 $Y=0.865
+ $X2=11.015 $Y2=0.94
r240 10 12 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=11.015 $Y=0.865
+ $X2=11.015 $Y2=0.58
r241 3 76 600 $w=1.7e-07 $l=2.74955e-07 $layer=licon1_PDIFF $count=1 $X=10.965
+ $Y=2.54 $X2=11.115 $Y2=2.75
r242 2 67 600 $w=1.7e-07 $l=2.98831e-07 $layer=licon1_PDIFF $count=1 $X=8.975
+ $Y=1.87 $X2=9.21 $Y2=2.015
r243 1 63 91 $w=1.7e-07 $l=3.44964e-07 $layer=licon1_NDIFF $count=2 $X=8.81
+ $Y=0.37 $X2=9.09 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__SDFSBP_1%A_2556_94# 1 2 7 9 12 14 15 16 18 22
r45 26 27 19.3931 $w=3.46e-07 $l=5.5e-07 $layer=LI1_cond $X=13.047 $Y=0.835
+ $X2=13.047 $Y2=1.385
r46 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=13.62
+ $Y=1.385 $X2=13.62 $Y2=1.385
r47 20 27 1.00354 $w=3.3e-07 $l=2.08e-07 $layer=LI1_cond $X=13.255 $Y=1.385
+ $X2=13.047 $Y2=1.385
r48 20 22 12.7467 $w=3.28e-07 $l=3.65e-07 $layer=LI1_cond $X=13.255 $Y=1.385
+ $X2=13.62 $Y2=1.385
r49 16 27 6.77755 $w=3.46e-07 $l=2.02287e-07 $layer=LI1_cond $X=13.13 $Y=1.55
+ $X2=13.047 $Y2=1.385
r50 16 18 28.1196 $w=2.48e-07 $l=6.1e-07 $layer=LI1_cond $X=13.13 $Y=1.55
+ $X2=13.13 $Y2=2.16
r51 14 23 33.2236 $w=3.3e-07 $l=1.9e-07 $layer=POLY_cond $X=13.81 $Y=1.385
+ $X2=13.62 $Y2=1.385
r52 14 15 66.2869 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=13.9 $Y=1.385
+ $X2=13.9 $Y2=1.22
r53 12 15 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=13.905 $Y=0.74
+ $X2=13.905 $Y2=1.22
r54 7 14 149.859 $w=1.8e-07 $l=3.8e-07 $layer=POLY_cond $X=13.9 $Y=1.765
+ $X2=13.9 $Y2=1.385
r55 7 9 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=13.9 $Y=1.765
+ $X2=13.9 $Y2=2.4
r56 2 18 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=13.03
+ $Y=2.015 $X2=13.17 $Y2=2.16
r57 1 26 182 $w=1.7e-07 $l=4.31451e-07 $layer=licon1_NDIFF $count=1 $X=12.78
+ $Y=0.47 $X2=12.925 $Y2=0.835
.ends

.subckt PM_SKY130_FD_SC_HS__SDFSBP_1%VPWR 1 2 3 4 5 6 7 8 27 31 33 37 41 45 49
+ 53 57 60 61 63 64 66 67 68 70 75 102 109 116 117 120 123 126 129 132
c160 117 0 9.63842e-20 $X=14.16 $Y=3.33
c161 37 0 2.13729e-19 $X=3.74 $Y=2.78
r162 132 133 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.68 $Y=3.33
+ $X2=13.68 $Y2=3.33
r163 129 130 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=12.24 $Y=3.33
+ $X2=12.24 $Y2=3.33
r164 126 127 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r165 124 127 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.6 $Y2=3.33
r166 123 124 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r167 120 121 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r168 117 133 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=14.16 $Y=3.33
+ $X2=13.68 $Y2=3.33
r169 116 117 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=14.16 $Y=3.33
+ $X2=14.16 $Y2=3.33
r170 114 132 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=13.785 $Y=3.33
+ $X2=13.62 $Y2=3.33
r171 114 116 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=13.785 $Y=3.33
+ $X2=14.16 $Y2=3.33
r172 113 133 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=13.2 $Y=3.33
+ $X2=13.68 $Y2=3.33
r173 113 130 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=13.2 $Y=3.33
+ $X2=12.24 $Y2=3.33
r174 112 113 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=13.2 $Y=3.33
+ $X2=13.2 $Y2=3.33
r175 110 129 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12.28 $Y=3.33
+ $X2=12.115 $Y2=3.33
r176 110 112 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=12.28 $Y=3.33
+ $X2=13.2 $Y2=3.33
r177 109 132 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=13.455 $Y=3.33
+ $X2=13.62 $Y2=3.33
r178 109 112 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=13.455 $Y=3.33
+ $X2=13.2 $Y2=3.33
r179 108 130 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.76 $Y=3.33
+ $X2=12.24 $Y2=3.33
r180 107 108 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=11.76 $Y=3.33
+ $X2=11.76 $Y2=3.33
r181 105 108 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=10.8 $Y=3.33
+ $X2=11.76 $Y2=3.33
r182 104 107 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=10.8 $Y=3.33
+ $X2=11.76 $Y2=3.33
r183 104 105 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=10.8 $Y=3.33
+ $X2=10.8 $Y2=3.33
r184 102 129 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.95 $Y=3.33
+ $X2=12.115 $Y2=3.33
r185 102 107 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=11.95 $Y=3.33
+ $X2=11.76 $Y2=3.33
r186 101 105 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.32 $Y=3.33
+ $X2=10.8 $Y2=3.33
r187 100 101 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=10.32 $Y=3.33
+ $X2=10.32 $Y2=3.33
r188 98 101 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=7.92 $Y=3.33
+ $X2=10.32 $Y2=3.33
r189 97 100 156.578 $w=1.68e-07 $l=2.4e-06 $layer=LI1_cond $X=7.92 $Y=3.33
+ $X2=10.32 $Y2=3.33
r190 97 98 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r191 95 98 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=7.92 $Y2=3.33
r192 94 95 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r193 91 94 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=6.48 $Y=3.33
+ $X2=7.44 $Y2=3.33
r194 91 92 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r195 89 92 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=3.33 $X2=6.48
+ $Y2=3.33
r196 88 89 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r197 86 89 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=6 $Y2=3.33
r198 86 127 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=3.6 $Y2=3.33
r199 85 88 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=4.08 $Y=3.33 $X2=6
+ $Y2=3.33
r200 85 86 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r201 83 126 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.905 $Y=3.33
+ $X2=3.74 $Y2=3.33
r202 83 85 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=3.905 $Y=3.33
+ $X2=4.08 $Y2=3.33
r203 82 124 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r204 81 82 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r205 79 82 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.16 $Y2=3.33
r206 79 121 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r207 78 81 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.2 $Y=3.33 $X2=2.16
+ $Y2=3.33
r208 78 79 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r209 76 120 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.895 $Y=3.33
+ $X2=0.73 $Y2=3.33
r210 76 78 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.895 $Y=3.33
+ $X2=1.2 $Y2=3.33
r211 75 123 7.34436 $w=1.7e-07 $l=1.32e-07 $layer=LI1_cond $X=2.555 $Y=3.33
+ $X2=2.687 $Y2=3.33
r212 75 81 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=2.555 $Y=3.33
+ $X2=2.16 $Y2=3.33
r213 73 121 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r214 72 73 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r215 70 120 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.565 $Y=3.33
+ $X2=0.73 $Y2=3.33
r216 70 72 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.565 $Y=3.33
+ $X2=0.24 $Y2=3.33
r217 68 95 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=7.2 $Y=3.33
+ $X2=7.44 $Y2=3.33
r218 68 92 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=7.2 $Y=3.33
+ $X2=6.48 $Y2=3.33
r219 66 100 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=10.58 $Y=3.33
+ $X2=10.32 $Y2=3.33
r220 66 67 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.58 $Y=3.33
+ $X2=10.665 $Y2=3.33
r221 65 104 3.26203 $w=1.68e-07 $l=5e-08 $layer=LI1_cond $X=10.75 $Y=3.33
+ $X2=10.8 $Y2=3.33
r222 65 67 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.75 $Y=3.33
+ $X2=10.665 $Y2=3.33
r223 63 94 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=7.615 $Y=3.33
+ $X2=7.44 $Y2=3.33
r224 63 64 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.615 $Y=3.33
+ $X2=7.7 $Y2=3.33
r225 62 97 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=7.785 $Y=3.33
+ $X2=7.92 $Y2=3.33
r226 62 64 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.785 $Y=3.33
+ $X2=7.7 $Y2=3.33
r227 60 88 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=6.175 $Y=3.33
+ $X2=6 $Y2=3.33
r228 60 61 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.175 $Y=3.33
+ $X2=6.3 $Y2=3.33
r229 59 91 3.58824 $w=1.68e-07 $l=5.5e-08 $layer=LI1_cond $X=6.425 $Y=3.33
+ $X2=6.48 $Y2=3.33
r230 59 61 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.425 $Y=3.33
+ $X2=6.3 $Y2=3.33
r231 55 132 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=13.62 $Y=3.245
+ $X2=13.62 $Y2=3.33
r232 55 57 37.8909 $w=3.28e-07 $l=1.085e-06 $layer=LI1_cond $X=13.62 $Y=3.245
+ $X2=13.62 $Y2=2.16
r233 51 129 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=12.115 $Y=3.245
+ $X2=12.115 $Y2=3.33
r234 51 53 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=12.115 $Y=3.245
+ $X2=12.115 $Y2=2.75
r235 47 67 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.665 $Y=3.245
+ $X2=10.665 $Y2=3.33
r236 47 49 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=10.665 $Y=3.245
+ $X2=10.665 $Y2=2.75
r237 43 64 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.7 $Y=3.245 $X2=7.7
+ $Y2=3.33
r238 43 45 46.9733 $w=1.68e-07 $l=7.2e-07 $layer=LI1_cond $X=7.7 $Y=3.245
+ $X2=7.7 $Y2=2.525
r239 39 61 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.3 $Y=3.245
+ $X2=6.3 $Y2=3.33
r240 39 41 30.194 $w=2.48e-07 $l=6.55e-07 $layer=LI1_cond $X=6.3 $Y=3.245
+ $X2=6.3 $Y2=2.59
r241 35 126 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.74 $Y=3.245
+ $X2=3.74 $Y2=3.33
r242 35 37 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=3.74 $Y=3.245
+ $X2=3.74 $Y2=2.78
r243 34 123 7.34436 $w=1.7e-07 $l=1.33e-07 $layer=LI1_cond $X=2.82 $Y=3.33
+ $X2=2.687 $Y2=3.33
r244 33 126 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.575 $Y=3.33
+ $X2=3.74 $Y2=3.33
r245 33 34 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=3.575 $Y=3.33
+ $X2=2.82 $Y2=3.33
r246 29 123 0.195364 $w=2.65e-07 $l=8.5e-08 $layer=LI1_cond $X=2.687 $Y=3.245
+ $X2=2.687 $Y2=3.33
r247 29 31 18.2651 $w=2.63e-07 $l=4.2e-07 $layer=LI1_cond $X=2.687 $Y=3.245
+ $X2=2.687 $Y2=2.825
r248 25 120 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.73 $Y=3.245
+ $X2=0.73 $Y2=3.33
r249 25 27 15.3659 $w=3.28e-07 $l=4.4e-07 $layer=LI1_cond $X=0.73 $Y=3.245
+ $X2=0.73 $Y2=2.805
r250 8 57 300 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=2 $X=13.47
+ $Y=2.015 $X2=13.62 $Y2=2.16
r251 7 53 600 $w=1.7e-07 $l=2.74955e-07 $layer=licon1_PDIFF $count=1 $X=11.965
+ $Y=2.54 $X2=12.115 $Y2=2.75
r252 6 49 600 $w=1.7e-07 $l=2.74955e-07 $layer=licon1_PDIFF $count=1 $X=10.515
+ $Y=2.54 $X2=10.665 $Y2=2.75
r253 5 45 600 $w=1.7e-07 $l=3.28634e-07 $layer=licon1_PDIFF $count=1 $X=7.46
+ $Y=2.315 $X2=7.7 $Y2=2.525
r254 4 41 600 $w=1.7e-07 $l=3.43875e-07 $layer=licon1_PDIFF $count=1 $X=6.185
+ $Y=2.315 $X2=6.34 $Y2=2.59
r255 3 37 600 $w=1.7e-07 $l=1.01223e-06 $layer=licon1_PDIFF $count=1 $X=3.59
+ $Y=1.84 $X2=3.74 $Y2=2.78
r256 2 31 600 $w=1.7e-07 $l=5.77321e-07 $layer=licon1_PDIFF $count=1 $X=2.5
+ $Y=2.32 $X2=2.655 $Y2=2.825
r257 1 27 600 $w=1.7e-07 $l=5.54955e-07 $layer=licon1_PDIFF $count=1 $X=0.58
+ $Y=2.32 $X2=0.73 $Y2=2.805
.ends

.subckt PM_SKY130_FD_SC_HS__SDFSBP_1%A_290_464# 1 2 3 4 13 19 21 22 23 26 28 29
+ 31 34 37 39 40 41 48 50
c122 26 0 1.9349e-19 $X=2.3 $Y=2.32
c123 22 0 4.07687e-19 $X=1.835 $Y=1.005
r124 45 48 3.49225 $w=3.28e-07 $l=1e-07 $layer=LI1_cond $X=4.505 $Y=0.76
+ $X2=4.605 $Y2=0.76
r125 41 43 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=3.71 $Y=2.295
+ $X2=3.71 $Y2=2.405
r126 35 50 3.67481 $w=2.52e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.757 $Y=2.38
+ $X2=4.672 $Y2=2.295
r127 35 37 4.64417 $w=3.33e-07 $l=1.35e-07 $layer=LI1_cond $X=4.757 $Y=2.38
+ $X2=4.757 $Y2=2.515
r128 34 50 3.67481 $w=2.52e-07 $l=2.05144e-07 $layer=LI1_cond $X=4.505 $Y=2.21
+ $X2=4.672 $Y2=2.295
r129 33 45 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.505 $Y=0.925
+ $X2=4.505 $Y2=0.76
r130 33 34 83.8342 $w=1.68e-07 $l=1.285e-06 $layer=LI1_cond $X=4.505 $Y=0.925
+ $X2=4.505 $Y2=2.21
r131 32 41 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.795 $Y=2.295
+ $X2=3.71 $Y2=2.295
r132 31 50 2.79892 $w=1.7e-07 $l=2.52e-07 $layer=LI1_cond $X=4.42 $Y=2.295
+ $X2=4.672 $Y2=2.295
r133 31 32 40.7754 $w=1.68e-07 $l=6.25e-07 $layer=LI1_cond $X=4.42 $Y=2.295
+ $X2=3.795 $Y2=2.295
r134 30 40 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.385 $Y=2.405
+ $X2=2.3 $Y2=2.405
r135 29 43 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.625 $Y=2.405
+ $X2=3.71 $Y2=2.405
r136 29 30 80.8984 $w=1.68e-07 $l=1.24e-06 $layer=LI1_cond $X=3.625 $Y=2.405
+ $X2=2.385 $Y2=2.405
r137 27 40 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.3 $Y=2.49 $X2=2.3
+ $Y2=2.405
r138 27 28 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=2.3 $Y=2.49 $X2=2.3
+ $Y2=2.63
r139 26 40 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.3 $Y=2.32 $X2=2.3
+ $Y2=2.405
r140 25 26 80.246 $w=1.68e-07 $l=1.23e-06 $layer=LI1_cond $X=2.3 $Y=1.09 $X2=2.3
+ $Y2=2.32
r141 23 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.215 $Y=2.715
+ $X2=2.3 $Y2=2.63
r142 23 39 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=2.215 $Y=2.715
+ $X2=1.945 $Y2=2.715
r143 21 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.215 $Y=1.005
+ $X2=2.3 $Y2=1.09
r144 21 22 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=2.215 $Y=1.005
+ $X2=1.835 $Y2=1.005
r145 17 22 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.67 $Y=0.92
+ $X2=1.835 $Y2=1.005
r146 17 19 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=1.67 $Y=0.92
+ $X2=1.67 $Y2=0.58
r147 13 39 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=1.78 $Y=2.795
+ $X2=1.945 $Y2=2.795
r148 13 15 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=1.78 $Y=2.795
+ $X2=1.69 $Y2=2.795
r149 4 37 600 $w=1.7e-07 $l=2.58844e-07 $layer=licon1_PDIFF $count=1 $X=4.625
+ $Y=2.315 $X2=4.76 $Y2=2.515
r150 3 15 600 $w=1.7e-07 $l=5.82774e-07 $layer=licon1_PDIFF $count=1 $X=1.45
+ $Y=2.32 $X2=1.69 $Y2=2.795
r151 2 48 182 $w=1.7e-07 $l=4.56782e-07 $layer=licon1_NDIFF $count=1 $X=4.46
+ $Y=0.37 $X2=4.605 $Y2=0.76
r152 1 19 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.53
+ $Y=0.37 $X2=1.67 $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_HS__SDFSBP_1%A_1600_347# 1 2 7 9 16
c36 9 0 2.64934e-19 $X=8.15 $Y=2.435
r37 9 12 2.96841 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=8.15 $Y=2.435
+ $X2=8.15 $Y2=2.52
r38 8 9 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.315 $Y=2.435
+ $X2=8.15 $Y2=2.435
r39 7 16 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=9.58 $Y=2.435
+ $X2=9.705 $Y2=2.435
r40 7 8 82.5294 $w=1.68e-07 $l=1.265e-06 $layer=LI1_cond $X=9.58 $Y=2.435
+ $X2=8.315 $Y2=2.435
r41 2 16 600 $w=1.7e-07 $l=7.11056e-07 $layer=licon1_PDIFF $count=1 $X=9.515
+ $Y=1.87 $X2=9.665 $Y2=2.51
r42 1 12 600 $w=1.7e-07 $l=8.56723e-07 $layer=licon1_PDIFF $count=1 $X=8
+ $Y=1.735 $X2=8.15 $Y2=2.52
.ends

.subckt PM_SKY130_FD_SC_HS__SDFSBP_1%A_1712_374# 1 2 7 11 14
c34 14 0 1.1962e-19 $X=8.695 $Y=2.855
r35 14 16 4.71454 $w=3.28e-07 $l=1.35e-07 $layer=LI1_cond $X=8.695 $Y=2.855
+ $X2=8.695 $Y2=2.99
r36 9 11 5.41299 $w=3.28e-07 $l=1.55e-07 $layer=LI1_cond $X=10.215 $Y=2.905
+ $X2=10.215 $Y2=2.75
r37 8 16 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.86 $Y=2.99
+ $X2=8.695 $Y2=2.99
r38 7 9 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=10.05 $Y=2.99
+ $X2=10.215 $Y2=2.905
r39 7 8 77.6364 $w=1.68e-07 $l=1.19e-06 $layer=LI1_cond $X=10.05 $Y=2.99
+ $X2=8.86 $Y2=2.99
r40 2 11 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=10.075
+ $Y=2.54 $X2=10.215 $Y2=2.75
r41 1 14 600 $w=1.7e-07 $l=1.05033e-06 $layer=licon1_PDIFF $count=1 $X=8.56
+ $Y=1.87 $X2=8.695 $Y2=2.855
.ends

.subckt PM_SKY130_FD_SC_HS__SDFSBP_1%Q_N 1 2 9 11 15 16 17 28
c35 15 0 1.92388e-19 $X=12.577 $Y=1.82
r36 21 28 1.01485 $w=4.93e-07 $l=4.2e-08 $layer=LI1_cond $X=12.372 $Y=0.883
+ $X2=12.372 $Y2=0.925
r37 17 30 9.94566 $w=4.93e-07 $l=1.84e-07 $layer=LI1_cond $X=12.372 $Y=0.946
+ $X2=12.372 $Y2=1.13
r38 17 28 0.507427 $w=4.93e-07 $l=2.1e-08 $layer=LI1_cond $X=12.372 $Y=0.946
+ $X2=12.372 $Y2=0.925
r39 17 21 0.53159 $w=4.93e-07 $l=2.2e-08 $layer=LI1_cond $X=12.372 $Y=0.861
+ $X2=12.372 $Y2=0.883
r40 16 17 8.36047 $w=4.93e-07 $l=3.46e-07 $layer=LI1_cond $X=12.372 $Y=0.515
+ $X2=12.372 $Y2=0.861
r41 15 30 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=12.535 $Y=1.82
+ $X2=12.535 $Y2=1.13
r42 11 13 37.5109 $w=2.53e-07 $l=8.3e-07 $layer=LI1_cond $X=12.577 $Y=1.985
+ $X2=12.577 $Y2=2.815
r43 9 15 7.02311 $w=2.53e-07 $l=1.27e-07 $layer=LI1_cond $X=12.577 $Y=1.947
+ $X2=12.577 $Y2=1.82
r44 9 11 1.71737 $w=2.53e-07 $l=3.8e-08 $layer=LI1_cond $X=12.577 $Y=1.947
+ $X2=12.577 $Y2=1.985
r45 2 13 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=12.47
+ $Y=1.84 $X2=12.62 $Y2=2.815
r46 2 11 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=12.47
+ $Y=1.84 $X2=12.62 $Y2=1.985
r47 1 16 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=12.15
+ $Y=0.37 $X2=12.29 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__SDFSBP_1%Q 1 2 7 8 9 10 11 12 13
r14 12 13 12.7285 $w=3.33e-07 $l=3.7e-07 $layer=LI1_cond $X=14.122 $Y=2.405
+ $X2=14.122 $Y2=2.775
r15 11 12 14.4485 $w=3.33e-07 $l=4.2e-07 $layer=LI1_cond $X=14.122 $Y=1.985
+ $X2=14.122 $Y2=2.405
r16 10 11 11.0084 $w=3.33e-07 $l=3.2e-07 $layer=LI1_cond $X=14.122 $Y=1.665
+ $X2=14.122 $Y2=1.985
r17 9 10 12.7285 $w=3.33e-07 $l=3.7e-07 $layer=LI1_cond $X=14.122 $Y=1.295
+ $X2=14.122 $Y2=1.665
r18 8 9 12.7285 $w=3.33e-07 $l=3.7e-07 $layer=LI1_cond $X=14.122 $Y=0.925
+ $X2=14.122 $Y2=1.295
r19 7 8 14.1045 $w=3.33e-07 $l=4.1e-07 $layer=LI1_cond $X=14.122 $Y=0.515
+ $X2=14.122 $Y2=0.925
r20 2 13 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=13.975
+ $Y=1.84 $X2=14.125 $Y2=2.815
r21 2 11 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=13.975
+ $Y=1.84 $X2=14.125 $Y2=1.985
r22 1 7 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=13.98
+ $Y=0.37 $X2=14.12 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__SDFSBP_1%VGND 1 2 3 4 5 6 7 8 27 31 35 39 43 47 52
+ 53 55 56 57 59 71 89 94 99 109 110 113 116 121 124 127 135 138
r145 138 139 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.68 $Y=0
+ $X2=13.68 $Y2=0
r146 135 136 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.76 $Y=0
+ $X2=11.76 $Y2=0
r147 128 130 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.32 $Y=0
+ $X2=10.8 $Y2=0
r148 127 132 10.098 $w=6.08e-07 $l=5.15e-07 $layer=LI1_cond $X=10.59 $Y=0
+ $X2=10.59 $Y2=0.515
r149 127 130 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.8 $Y=0
+ $X2=10.8 $Y2=0
r150 127 128 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=10.32 $Y=0
+ $X2=10.32 $Y2=0
r151 123 124 11.5563 $w=8.18e-07 $l=1.65e-07 $layer=LI1_cond $X=8.13 $Y=0.325
+ $X2=8.295 $Y2=0.325
r152 119 123 3.06313 $w=8.18e-07 $l=2.1e-07 $layer=LI1_cond $X=7.92 $Y=0.325
+ $X2=8.13 $Y2=0.325
r153 119 121 15.2758 $w=8.18e-07 $l=4.2e-07 $layer=LI1_cond $X=7.92 $Y=0.325
+ $X2=7.5 $Y2=0.325
r154 119 120 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=0
+ $X2=7.92 $Y2=0
r155 116 117 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r156 113 114 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0
+ $X2=0.72 $Y2=0
r157 110 139 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=14.16 $Y=0
+ $X2=13.68 $Y2=0
r158 109 110 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=14.16 $Y=0
+ $X2=14.16 $Y2=0
r159 107 138 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=13.785 $Y=0
+ $X2=13.62 $Y2=0
r160 107 109 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=13.785 $Y=0
+ $X2=14.16 $Y2=0
r161 106 139 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=13.2 $Y=0
+ $X2=13.68 $Y2=0
r162 105 106 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=13.2 $Y=0
+ $X2=13.2 $Y2=0
r163 103 106 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=12.24 $Y=0
+ $X2=13.2 $Y2=0
r164 103 136 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.24 $Y=0
+ $X2=11.76 $Y2=0
r165 102 105 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=12.24 $Y=0
+ $X2=13.2 $Y2=0
r166 102 103 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=12.24 $Y=0
+ $X2=12.24 $Y2=0
r167 100 135 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.955 $Y=0
+ $X2=11.79 $Y2=0
r168 100 102 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=11.955 $Y=0
+ $X2=12.24 $Y2=0
r169 99 138 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=13.455 $Y=0
+ $X2=13.62 $Y2=0
r170 99 105 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=13.455 $Y=0
+ $X2=13.2 $Y2=0
r171 98 136 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.28 $Y=0
+ $X2=11.76 $Y2=0
r172 98 130 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.28 $Y=0
+ $X2=10.8 $Y2=0
r173 97 98 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.28 $Y=0
+ $X2=11.28 $Y2=0
r174 95 127 8.42348 $w=1.7e-07 $l=3.05e-07 $layer=LI1_cond $X=10.895 $Y=0
+ $X2=10.59 $Y2=0
r175 95 97 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=10.895 $Y=0
+ $X2=11.28 $Y2=0
r176 94 135 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.625 $Y=0
+ $X2=11.79 $Y2=0
r177 94 97 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=11.625 $Y=0
+ $X2=11.28 $Y2=0
r178 93 128 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=8.4 $Y=0
+ $X2=10.32 $Y2=0
r179 93 120 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=0 $X2=7.92
+ $Y2=0
r180 92 124 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=8.4 $Y=0
+ $X2=8.295 $Y2=0
r181 92 93 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r182 89 127 8.42348 $w=1.7e-07 $l=3.05e-07 $layer=LI1_cond $X=10.285 $Y=0
+ $X2=10.59 $Y2=0
r183 89 92 122.979 $w=1.68e-07 $l=1.885e-06 $layer=LI1_cond $X=10.285 $Y=0
+ $X2=8.4 $Y2=0
r184 88 120 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=0
+ $X2=7.92 $Y2=0
r185 87 121 3.91444 $w=1.68e-07 $l=6e-08 $layer=LI1_cond $X=7.44 $Y=0 $X2=7.5
+ $Y2=0
r186 87 88 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=7.44 $Y=0 $X2=7.44
+ $Y2=0
r187 84 87 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=6.48 $Y=0 $X2=7.44
+ $Y2=0
r188 84 85 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6.48 $Y=0 $X2=6.48
+ $Y2=0
r189 81 85 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=0 $X2=6.48
+ $Y2=0
r190 80 81 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6 $Y=0 $X2=6
+ $Y2=0
r191 78 81 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=4.08 $Y=0 $X2=6
+ $Y2=0
r192 78 117 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=3.6
+ $Y2=0
r193 77 80 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=4.08 $Y=0 $X2=6
+ $Y2=0
r194 77 78 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.08 $Y=0
+ $X2=4.08 $Y2=0
r195 75 116 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.71 $Y=0
+ $X2=3.545 $Y2=0
r196 75 77 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=3.71 $Y=0 $X2=4.08
+ $Y2=0
r197 74 117 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=3.6
+ $Y2=0
r198 73 74 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r199 71 116 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.38 $Y=0
+ $X2=3.545 $Y2=0
r200 71 73 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=3.38 $Y=0 $X2=3.12
+ $Y2=0
r201 70 74 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=3.12
+ $Y2=0
r202 69 70 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r203 67 70 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r204 67 114 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r205 66 69 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r206 66 67 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r207 64 113 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.945 $Y=0
+ $X2=0.78 $Y2=0
r208 64 66 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.945 $Y=0 $X2=1.2
+ $Y2=0
r209 62 114 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0
+ $X2=0.72 $Y2=0
r210 61 62 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r211 59 113 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.615 $Y=0
+ $X2=0.78 $Y2=0
r212 59 61 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=0.615 $Y=0
+ $X2=0.24 $Y2=0
r213 57 88 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=7.2 $Y=0 $X2=7.44
+ $Y2=0
r214 57 85 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=7.2 $Y=0 $X2=6.48
+ $Y2=0
r215 55 80 1.30481 $w=1.68e-07 $l=2e-08 $layer=LI1_cond $X=6.02 $Y=0 $X2=6 $Y2=0
r216 55 56 8.9695 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=6.02 $Y=0 $X2=6.195
+ $Y2=0
r217 54 84 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=6.37 $Y=0 $X2=6.48
+ $Y2=0
r218 54 56 8.9695 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=6.37 $Y=0 $X2=6.195
+ $Y2=0
r219 52 69 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=2.325 $Y=0
+ $X2=2.16 $Y2=0
r220 52 53 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.325 $Y=0 $X2=2.49
+ $Y2=0
r221 51 73 30.3369 $w=1.68e-07 $l=4.65e-07 $layer=LI1_cond $X=2.655 $Y=0
+ $X2=3.12 $Y2=0
r222 51 53 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.655 $Y=0 $X2=2.49
+ $Y2=0
r223 47 49 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=13.62 $Y=0.515
+ $X2=13.62 $Y2=0.885
r224 45 138 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=13.62 $Y=0.085
+ $X2=13.62 $Y2=0
r225 45 47 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=13.62 $Y=0.085
+ $X2=13.62 $Y2=0.515
r226 41 135 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=11.79 $Y=0.085
+ $X2=11.79 $Y2=0
r227 41 43 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=11.79 $Y=0.085
+ $X2=11.79 $Y2=0.515
r228 37 56 1.07557 $w=3.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.195 $Y=0.085
+ $X2=6.195 $Y2=0
r229 37 39 13.0061 $w=3.48e-07 $l=3.95e-07 $layer=LI1_cond $X=6.195 $Y=0.085
+ $X2=6.195 $Y2=0.48
r230 33 116 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.545 $Y=0.085
+ $X2=3.545 $Y2=0
r231 33 35 14.6675 $w=3.28e-07 $l=4.2e-07 $layer=LI1_cond $X=3.545 $Y=0.085
+ $X2=3.545 $Y2=0.505
r232 29 53 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.49 $Y=0.085
+ $X2=2.49 $Y2=0
r233 29 31 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=2.49 $Y=0.085
+ $X2=2.49 $Y2=0.55
r234 25 113 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.78 $Y=0.085
+ $X2=0.78 $Y2=0
r235 25 27 16.7628 $w=3.28e-07 $l=4.8e-07 $layer=LI1_cond $X=0.78 $Y=0.085
+ $X2=0.78 $Y2=0.565
r236 8 49 182 $w=1.7e-07 $l=5.83352e-07 $layer=licon1_NDIFF $count=1 $X=13.215
+ $Y=0.47 $X2=13.62 $Y2=0.885
r237 8 47 182 $w=1.7e-07 $l=4.26907e-07 $layer=licon1_NDIFF $count=1 $X=13.215
+ $Y=0.47 $X2=13.62 $Y2=0.515
r238 7 43 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=11.645
+ $Y=0.37 $X2=11.79 $Y2=0.515
r239 6 132 91 $w=1.7e-07 $l=5.57808e-07 $layer=licon1_NDIFF $count=2 $X=10.31
+ $Y=0.37 $X2=10.8 $Y2=0.515
r240 5 123 91 $w=1.7e-07 $l=7.78604e-07 $layer=licon1_NDIFF $count=2 $X=7.445
+ $Y=0.37 $X2=8.13 $Y2=0.57
r241 4 39 182 $w=1.7e-07 $l=2.79643e-07 $layer=licon1_NDIFF $count=1 $X=5.965
+ $Y=0.37 $X2=6.195 $Y2=0.48
r242 3 35 91 $w=1.7e-07 $l=1.96214e-07 $layer=licon1_NDIFF $count=2 $X=3.405
+ $Y=0.37 $X2=3.545 $Y2=0.505
r243 2 31 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=2.35 $Y=0.37
+ $X2=2.49 $Y2=0.55
r244 1 27 182 $w=1.7e-07 $l=2.91633e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.37 $X2=0.78 $Y2=0.565
.ends

