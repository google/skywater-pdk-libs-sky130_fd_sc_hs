* File: sky130_fd_sc_hs__nor4b_4.pex.spice
* Created: Tue Sep  1 20:12:33 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HS__NOR4B_4%D_N 1 3 4 6 7 9 10 11 16 18
r37 18 19 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=0.385
+ $Y=1.765 $X2=0.385 $Y2=1.765
r38 15 18 49.3614 $w=6.64e-07 $l=7.995e-07 $layer=POLY_cond $X=0.385 $Y=1.085
+ $X2=0.645 $Y2=1.765
r39 15 16 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=0.385
+ $Y=1.085 $X2=0.385 $Y2=1.085
r40 11 19 2.71163 $w=4.23e-07 $l=1e-07 $layer=LI1_cond $X=0.337 $Y=1.665
+ $X2=0.337 $Y2=1.765
r41 10 11 10.033 $w=4.23e-07 $l=3.7e-07 $layer=LI1_cond $X=0.337 $Y=1.295
+ $X2=0.337 $Y2=1.665
r42 10 16 5.69442 $w=4.23e-07 $l=2.1e-07 $layer=LI1_cond $X=0.337 $Y=1.295
+ $X2=0.337 $Y2=1.085
r43 7 15 41.5788 $w=6.64e-07 $l=6.58103e-07 $layer=POLY_cond $X=0.995 $Y=1.185
+ $X2=0.385 $Y2=1.085
r44 7 9 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=0.995 $Y=1.185
+ $X2=0.995 $Y2=0.74
r45 4 18 44.0784 $w=3.32e-07 $l=4.27668e-07 $layer=POLY_cond $X=0.955 $Y=2.045
+ $X2=0.645 $Y2=1.765
r46 4 6 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=0.955 $Y=2.045
+ $X2=0.955 $Y2=2.54
r47 1 18 44.0784 $w=3.32e-07 $l=3.42929e-07 $layer=POLY_cond $X=0.505 $Y=2.045
+ $X2=0.645 $Y2=1.765
r48 1 3 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=0.505 $Y=2.045
+ $X2=0.505 $Y2=2.54
.ends

.subckt PM_SKY130_FD_SC_HS__NOR4B_4%A_47_88# 1 2 9 13 15 17 18 20 23 27 29 31 32
+ 33 34 36 37 43 45 46 54 57 60
c122 34 0 1.227e-20 $X=3.365 $Y=1.765
c123 27 0 3.90676e-20 $X=2.88 $Y=0.74
c124 23 0 1.09607e-20 $X=2.45 $Y=0.74
r125 68 69 4.11463 $w=4.1e-07 $l=3.5e-08 $layer=POLY_cond $X=2.88 $Y=1.542
+ $X2=2.915 $Y2=1.542
r126 67 68 50.5512 $w=4.1e-07 $l=4.3e-07 $layer=POLY_cond $X=2.45 $Y=1.542
+ $X2=2.88 $Y2=1.542
r127 66 67 4.11463 $w=4.1e-07 $l=3.5e-08 $layer=POLY_cond $X=2.415 $Y=1.542
+ $X2=2.45 $Y2=1.542
r128 63 64 1.76341 $w=4.1e-07 $l=1.5e-08 $layer=POLY_cond $X=1.95 $Y=1.542
+ $X2=1.965 $Y2=1.542
r129 55 66 29.3902 $w=4.1e-07 $l=2.5e-07 $layer=POLY_cond $X=2.165 $Y=1.542
+ $X2=2.415 $Y2=1.542
r130 55 64 23.5122 $w=4.1e-07 $l=2e-07 $layer=POLY_cond $X=2.165 $Y=1.542
+ $X2=1.965 $Y2=1.542
r131 54 55 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=2.165
+ $Y=1.485 $X2=2.165 $Y2=1.485
r132 52 63 54.6659 $w=4.1e-07 $l=4.65e-07 $layer=POLY_cond $X=1.485 $Y=1.542
+ $X2=1.95 $Y2=1.542
r133 52 61 5.29024 $w=4.1e-07 $l=4.5e-08 $layer=POLY_cond $X=1.485 $Y=1.542
+ $X2=1.44 $Y2=1.542
r134 51 54 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=1.485 $Y=1.485
+ $X2=2.165 $Y2=1.485
r135 51 52 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.485
+ $Y=1.485 $X2=1.485 $Y2=1.485
r136 49 60 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.89 $Y=1.485
+ $X2=0.805 $Y2=1.485
r137 49 51 20.7789 $w=3.28e-07 $l=5.95e-07 $layer=LI1_cond $X=0.89 $Y=1.485
+ $X2=1.485 $Y2=1.485
r138 47 60 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.805 $Y=1.65
+ $X2=0.805 $Y2=1.485
r139 47 57 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=0.805 $Y=1.65
+ $X2=0.805 $Y2=2.1
r140 46 60 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.805 $Y=1.32
+ $X2=0.805 $Y2=1.485
r141 45 59 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.805 $Y=0.75
+ $X2=0.805 $Y2=0.585
r142 45 46 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=0.805 $Y=0.75
+ $X2=0.805 $Y2=1.32
r143 43 57 8.30336 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=0.73 $Y=2.265
+ $X2=0.73 $Y2=2.1
r144 37 59 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.72 $Y=0.585
+ $X2=0.805 $Y2=0.585
r145 37 39 9.7783 $w=3.28e-07 $l=2.8e-07 $layer=LI1_cond $X=0.72 $Y=0.585
+ $X2=0.44 $Y2=0.585
r146 34 36 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.365 $Y=1.765
+ $X2=3.365 $Y2=2.4
r147 33 69 30.9697 $w=4.1e-07 $l=1.46233e-07 $layer=POLY_cond $X=3.005 $Y=1.65
+ $X2=2.915 $Y2=1.542
r148 32 34 26.9307 $w=1.5e-07 $l=1.53542e-07 $layer=POLY_cond $X=3.275 $Y=1.65
+ $X2=3.365 $Y2=1.765
r149 32 33 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=3.275 $Y=1.65
+ $X2=3.005 $Y2=1.65
r150 29 69 26.4667 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=2.915 $Y=1.765
+ $X2=2.915 $Y2=1.542
r151 29 31 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.915 $Y=1.765
+ $X2=2.915 $Y2=2.4
r152 25 68 26.4667 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=2.88 $Y=1.32
+ $X2=2.88 $Y2=1.542
r153 25 27 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=2.88 $Y=1.32
+ $X2=2.88 $Y2=0.74
r154 21 67 26.4667 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=2.45 $Y=1.32
+ $X2=2.45 $Y2=1.542
r155 21 23 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=2.45 $Y=1.32
+ $X2=2.45 $Y2=0.74
r156 18 66 26.4667 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=2.415 $Y=1.765
+ $X2=2.415 $Y2=1.542
r157 18 20 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.415 $Y=1.765
+ $X2=2.415 $Y2=2.4
r158 15 64 26.4667 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=1.965 $Y=1.765
+ $X2=1.965 $Y2=1.542
r159 15 17 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.965 $Y=1.765
+ $X2=1.965 $Y2=2.4
r160 11 63 26.4667 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=1.95 $Y=1.32
+ $X2=1.95 $Y2=1.542
r161 11 13 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=1.95 $Y=1.32
+ $X2=1.95 $Y2=0.74
r162 7 61 26.4667 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=1.44 $Y=1.32
+ $X2=1.44 $Y2=1.542
r163 7 9 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=1.44 $Y=1.32 $X2=1.44
+ $Y2=0.74
r164 2 43 300 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=2 $X=0.58
+ $Y=2.12 $X2=0.73 $Y2=2.265
r165 1 59 182 $w=1.7e-07 $l=6.13229e-07 $layer=licon1_NDIFF $count=1 $X=0.235
+ $Y=0.44 $X2=0.78 $Y2=0.585
r166 1 39 182 $w=1.7e-07 $l=2.67862e-07 $layer=licon1_NDIFF $count=1 $X=0.235
+ $Y=0.44 $X2=0.44 $Y2=0.585
.ends

.subckt PM_SKY130_FD_SC_HS__NOR4B_4%C 1 3 4 5 6 8 9 11 12 14 15 17 18 20 21 22
+ 23 25 27 28 30 31 32 33 34
c95 28 0 7.8278e-20 $X=5.315 $Y=1.765
c96 23 0 1.8401e-19 $X=5.285 $Y=1.185
c97 12 0 9.04372e-20 $X=4.315 $Y=1.765
c98 1 0 5.58611e-20 $X=3.45 $Y=1.185
r99 47 48 1.35647 $w=5.33e-07 $l=1.5e-08 $layer=POLY_cond $X=4.84 $Y=1.475
+ $X2=4.855 $Y2=1.475
r100 45 47 6.78236 $w=5.33e-07 $l=7.5e-08 $layer=POLY_cond $X=4.765 $Y=1.475
+ $X2=4.84 $Y2=1.475
r101 45 46 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.765
+ $Y=1.515 $X2=4.765 $Y2=1.515
r102 43 45 40.6942 $w=5.33e-07 $l=4.5e-07 $layer=POLY_cond $X=4.315 $Y=1.475
+ $X2=4.765 $Y2=1.475
r103 41 43 20.7992 $w=5.33e-07 $l=2.3e-07 $layer=POLY_cond $X=4.085 $Y=1.475
+ $X2=4.315 $Y2=1.475
r104 41 42 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.085
+ $Y=1.515 $X2=4.085 $Y2=1.515
r105 39 41 18.5385 $w=5.33e-07 $l=2.05e-07 $layer=POLY_cond $X=3.88 $Y=1.475
+ $X2=4.085 $Y2=1.475
r106 38 39 5.87805 $w=5.33e-07 $l=6.5e-08 $layer=POLY_cond $X=3.815 $Y=1.475
+ $X2=3.88 $Y2=1.475
r107 34 46 7.37028 $w=4.28e-07 $l=2.75e-07 $layer=LI1_cond $X=5.04 $Y=1.565
+ $X2=4.765 $Y2=1.565
r108 33 46 5.4942 $w=4.28e-07 $l=2.05e-07 $layer=LI1_cond $X=4.56 $Y=1.565
+ $X2=4.765 $Y2=1.565
r109 33 42 12.7305 $w=4.28e-07 $l=4.75e-07 $layer=LI1_cond $X=4.56 $Y=1.565
+ $X2=4.085 $Y2=1.565
r110 32 42 0.134005 $w=4.28e-07 $l=5e-09 $layer=LI1_cond $X=4.08 $Y=1.565
+ $X2=4.085 $Y2=1.565
r111 28 30 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=5.315 $Y=1.765
+ $X2=5.315 $Y2=2.4
r112 27 28 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=5.315 $Y=1.675
+ $X2=5.315 $Y2=1.765
r113 26 31 18.8402 $w=1.65e-07 $l=7.88987e-08 $layer=POLY_cond $X=5.315 $Y=1.335
+ $X2=5.307 $Y2=1.26
r114 26 27 132.161 $w=1.8e-07 $l=3.4e-07 $layer=POLY_cond $X=5.315 $Y=1.335
+ $X2=5.315 $Y2=1.675
r115 23 31 18.8402 $w=1.65e-07 $l=8.52936e-08 $layer=POLY_cond $X=5.285 $Y=1.185
+ $X2=5.307 $Y2=1.26
r116 23 25 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=5.285 $Y=1.185
+ $X2=5.285 $Y2=0.74
r117 22 48 34.6507 $w=5.33e-07 $l=2.497e-07 $layer=POLY_cond $X=4.93 $Y=1.26
+ $X2=4.855 $Y2=1.475
r118 21 31 6.66866 $w=1.5e-07 $l=9.7e-08 $layer=POLY_cond $X=5.21 $Y=1.26
+ $X2=5.307 $Y2=1.26
r119 21 22 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=5.21 $Y=1.26
+ $X2=4.93 $Y2=1.26
r120 18 48 33.0303 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=4.855 $Y=1.185
+ $X2=4.855 $Y2=1.475
r121 18 20 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=4.855 $Y=1.185
+ $X2=4.855 $Y2=0.74
r122 15 47 33.0303 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=4.84 $Y=1.765
+ $X2=4.84 $Y2=1.475
r123 15 17 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=4.84 $Y=1.765
+ $X2=4.84 $Y2=2.4
r124 12 43 33.0303 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=4.315 $Y=1.765
+ $X2=4.315 $Y2=1.475
r125 12 14 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=4.315 $Y=1.765
+ $X2=4.315 $Y2=2.4
r126 9 39 33.0303 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=3.88 $Y=1.185
+ $X2=3.88 $Y2=1.475
r127 9 11 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=3.88 $Y=1.185
+ $X2=3.88 $Y2=0.74
r128 6 38 33.0303 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=3.815 $Y=1.765
+ $X2=3.815 $Y2=1.475
r129 6 8 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.815 $Y=1.765
+ $X2=3.815 $Y2=2.4
r130 4 38 36.0072 $w=5.33e-07 $l=2.56076e-07 $layer=POLY_cond $X=3.725 $Y=1.26
+ $X2=3.815 $Y2=1.475
r131 4 5 102.553 $w=1.5e-07 $l=2e-07 $layer=POLY_cond $X=3.725 $Y=1.26 $X2=3.525
+ $Y2=1.26
r132 1 5 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.45 $Y=1.185
+ $X2=3.525 $Y2=1.26
r133 1 3 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=3.45 $Y=1.185
+ $X2=3.45 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HS__NOR4B_4%B 3 5 7 10 12 14 17 19 21 24 26 28 29 30 31
+ 32 49
c94 32 0 1.743e-19 $X=7.44 $Y=1.665
c95 19 0 1.14315e-20 $X=7.325 $Y=1.765
r96 49 50 19.1479 $w=3.65e-07 $l=1.45e-07 $layer=POLY_cond $X=7.63 $Y=1.557
+ $X2=7.775 $Y2=1.557
r97 48 49 40.2767 $w=3.65e-07 $l=3.05e-07 $layer=POLY_cond $X=7.325 $Y=1.557
+ $X2=7.63 $Y2=1.557
r98 46 48 1.98082 $w=3.65e-07 $l=1.5e-08 $layer=POLY_cond $X=7.31 $Y=1.557
+ $X2=7.325 $Y2=1.557
r99 46 47 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=7.31
+ $Y=1.515 $X2=7.31 $Y2=1.515
r100 44 46 14.526 $w=3.65e-07 $l=1.1e-07 $layer=POLY_cond $X=7.2 $Y=1.557
+ $X2=7.31 $Y2=1.557
r101 43 44 49.5205 $w=3.65e-07 $l=3.75e-07 $layer=POLY_cond $X=6.825 $Y=1.557
+ $X2=7.2 $Y2=1.557
r102 42 43 16.5068 $w=3.65e-07 $l=1.25e-07 $layer=POLY_cond $X=6.7 $Y=1.557
+ $X2=6.825 $Y2=1.557
r103 41 42 49.5205 $w=3.65e-07 $l=3.75e-07 $layer=POLY_cond $X=6.325 $Y=1.557
+ $X2=6.7 $Y2=1.557
r104 39 41 4.62192 $w=3.65e-07 $l=3.5e-08 $layer=POLY_cond $X=6.29 $Y=1.557
+ $X2=6.325 $Y2=1.557
r105 39 40 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.29
+ $Y=1.515 $X2=6.29 $Y2=1.515
r106 37 39 11.8849 $w=3.65e-07 $l=9e-08 $layer=POLY_cond $X=6.2 $Y=1.557
+ $X2=6.29 $Y2=1.557
r107 32 47 3.48413 $w=4.28e-07 $l=1.3e-07 $layer=LI1_cond $X=7.44 $Y=1.565
+ $X2=7.31 $Y2=1.565
r108 31 47 9.38035 $w=4.28e-07 $l=3.5e-07 $layer=LI1_cond $X=6.96 $Y=1.565
+ $X2=7.31 $Y2=1.565
r109 30 31 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=6.48 $Y=1.565
+ $X2=6.96 $Y2=1.565
r110 30 40 5.09219 $w=4.28e-07 $l=1.9e-07 $layer=LI1_cond $X=6.48 $Y=1.565
+ $X2=6.29 $Y2=1.565
r111 29 40 7.77229 $w=4.28e-07 $l=2.9e-07 $layer=LI1_cond $X=6 $Y=1.565 $X2=6.29
+ $Y2=1.565
r112 26 50 23.6381 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=7.775 $Y=1.765
+ $X2=7.775 $Y2=1.557
r113 26 28 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=7.775 $Y=1.765
+ $X2=7.775 $Y2=2.4
r114 22 49 23.6381 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=7.63 $Y=1.35
+ $X2=7.63 $Y2=1.557
r115 22 24 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=7.63 $Y=1.35
+ $X2=7.63 $Y2=0.74
r116 19 48 23.6381 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=7.325 $Y=1.765
+ $X2=7.325 $Y2=1.557
r117 19 21 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=7.325 $Y=1.765
+ $X2=7.325 $Y2=2.4
r118 15 44 23.6381 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=7.2 $Y=1.35
+ $X2=7.2 $Y2=1.557
r119 15 17 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=7.2 $Y=1.35 $X2=7.2
+ $Y2=0.74
r120 12 43 23.6381 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=6.825 $Y=1.765
+ $X2=6.825 $Y2=1.557
r121 12 14 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=6.825 $Y=1.765
+ $X2=6.825 $Y2=2.4
r122 8 42 23.6381 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=6.7 $Y=1.35 $X2=6.7
+ $Y2=1.557
r123 8 10 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=6.7 $Y=1.35 $X2=6.7
+ $Y2=0.74
r124 5 41 23.6381 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=6.325 $Y=1.765
+ $X2=6.325 $Y2=1.557
r125 5 7 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=6.325 $Y=1.765
+ $X2=6.325 $Y2=2.4
r126 1 37 23.6381 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=6.2 $Y=1.35 $X2=6.2
+ $Y2=1.557
r127 1 3 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=6.2 $Y=1.35 $X2=6.2
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HS__NOR4B_4%A 3 5 7 10 12 14 17 19 21 24 26 28 29 30 31
+ 32 48
c82 48 0 2.47857e-19 $X=9.515 $Y=1.557
c83 32 0 1.14315e-20 $X=9.36 $Y=1.665
r84 48 49 7.8587 $w=3.68e-07 $l=6e-08 $layer=POLY_cond $X=9.515 $Y=1.557
+ $X2=9.575 $Y2=1.557
r85 46 48 23.5761 $w=3.68e-07 $l=1.8e-07 $layer=POLY_cond $X=9.335 $Y=1.557
+ $X2=9.515 $Y2=1.557
r86 46 47 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=9.335
+ $Y=1.515 $X2=9.335 $Y2=1.515
r87 44 46 27.5054 $w=3.68e-07 $l=2.1e-07 $layer=POLY_cond $X=9.125 $Y=1.557
+ $X2=9.335 $Y2=1.557
r88 43 44 5.23913 $w=3.68e-07 $l=4e-08 $layer=POLY_cond $X=9.085 $Y=1.557
+ $X2=9.125 $Y2=1.557
r89 42 43 53.7011 $w=3.68e-07 $l=4.1e-07 $layer=POLY_cond $X=8.675 $Y=1.557
+ $X2=9.085 $Y2=1.557
r90 41 42 2.61957 $w=3.68e-07 $l=2e-08 $layer=POLY_cond $X=8.655 $Y=1.557
+ $X2=8.675 $Y2=1.557
r91 39 41 44.5326 $w=3.68e-07 $l=3.4e-07 $layer=POLY_cond $X=8.315 $Y=1.557
+ $X2=8.655 $Y2=1.557
r92 39 40 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=8.315
+ $Y=1.515 $X2=8.315 $Y2=1.515
r93 37 39 11.788 $w=3.68e-07 $l=9e-08 $layer=POLY_cond $X=8.225 $Y=1.557
+ $X2=8.315 $Y2=1.557
r94 32 47 0.670025 $w=4.28e-07 $l=2.5e-08 $layer=LI1_cond $X=9.36 $Y=1.565
+ $X2=9.335 $Y2=1.565
r95 31 47 12.1945 $w=4.28e-07 $l=4.55e-07 $layer=LI1_cond $X=8.88 $Y=1.565
+ $X2=9.335 $Y2=1.565
r96 30 31 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=8.4 $Y=1.565
+ $X2=8.88 $Y2=1.565
r97 30 40 2.27808 $w=4.28e-07 $l=8.5e-08 $layer=LI1_cond $X=8.4 $Y=1.565
+ $X2=8.315 $Y2=1.565
r98 29 40 10.5864 $w=4.28e-07 $l=3.95e-07 $layer=LI1_cond $X=7.92 $Y=1.565
+ $X2=8.315 $Y2=1.565
r99 26 49 23.8357 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=9.575 $Y=1.765
+ $X2=9.575 $Y2=1.557
r100 26 28 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=9.575 $Y=1.765
+ $X2=9.575 $Y2=2.4
r101 22 48 23.8357 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=9.515 $Y=1.35
+ $X2=9.515 $Y2=1.557
r102 22 24 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=9.515 $Y=1.35
+ $X2=9.515 $Y2=0.74
r103 19 44 23.8357 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=9.125 $Y=1.765
+ $X2=9.125 $Y2=1.557
r104 19 21 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=9.125 $Y=1.765
+ $X2=9.125 $Y2=2.4
r105 15 43 23.8357 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=9.085 $Y=1.35
+ $X2=9.085 $Y2=1.557
r106 15 17 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=9.085 $Y=1.35
+ $X2=9.085 $Y2=0.74
r107 12 42 23.8357 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=8.675 $Y=1.765
+ $X2=8.675 $Y2=1.557
r108 12 14 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=8.675 $Y=1.765
+ $X2=8.675 $Y2=2.4
r109 8 41 23.8357 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=8.655 $Y=1.35
+ $X2=8.655 $Y2=1.557
r110 8 10 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=8.655 $Y=1.35
+ $X2=8.655 $Y2=0.74
r111 5 37 23.8357 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=8.225 $Y=1.765
+ $X2=8.225 $Y2=1.557
r112 5 7 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=8.225 $Y=1.765
+ $X2=8.225 $Y2=2.4
r113 1 37 23.8357 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=8.225 $Y=1.35
+ $X2=8.225 $Y2=1.557
r114 1 3 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=8.225 $Y=1.35
+ $X2=8.225 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HS__NOR4B_4%VPWR 1 2 3 4 13 15 19 23 27 29 31 36 44 51
+ 52 58 61 64
r104 64 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.36 $Y=3.33
+ $X2=9.36 $Y2=3.33
r105 61 62 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=3.33 $X2=8.4
+ $Y2=3.33
r106 58 59 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r107 55 56 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r108 52 65 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.84 $Y=3.33
+ $X2=9.36 $Y2=3.33
r109 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.84 $Y=3.33
+ $X2=9.84 $Y2=3.33
r110 49 64 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=9.515 $Y=3.33
+ $X2=9.39 $Y2=3.33
r111 49 51 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=9.515 $Y=3.33
+ $X2=9.84 $Y2=3.33
r112 48 65 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=3.33
+ $X2=9.36 $Y2=3.33
r113 48 62 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=3.33
+ $X2=8.4 $Y2=3.33
r114 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r115 45 61 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.535 $Y=3.33
+ $X2=8.41 $Y2=3.33
r116 45 47 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=8.535 $Y=3.33
+ $X2=8.88 $Y2=3.33
r117 44 64 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=9.265 $Y=3.33
+ $X2=9.39 $Y2=3.33
r118 44 47 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=9.265 $Y=3.33
+ $X2=8.88 $Y2=3.33
r119 43 62 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=3.33
+ $X2=8.4 $Y2=3.33
r120 42 43 1.32857 $w=1.7e-07 $l=1.19e-06 $layer=mcon $count=7 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r121 40 59 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r122 39 42 407.102 $w=1.68e-07 $l=6.24e-06 $layer=LI1_cond $X=1.68 $Y=3.33
+ $X2=7.92 $Y2=3.33
r123 39 40 1.32857 $w=1.7e-07 $l=1.19e-06 $layer=mcon $count=7 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r124 37 58 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=1.345 $Y=3.33
+ $X2=1.21 $Y2=3.33
r125 37 39 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=1.345 $Y=3.33
+ $X2=1.68 $Y2=3.33
r126 36 61 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.285 $Y=3.33
+ $X2=8.41 $Y2=3.33
r127 36 42 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=8.285 $Y=3.33
+ $X2=7.92 $Y2=3.33
r128 35 59 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r129 35 56 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r130 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r131 32 55 4.00981 $w=1.7e-07 $l=1.83e-07 $layer=LI1_cond $X=0.365 $Y=3.33
+ $X2=0.182 $Y2=3.33
r132 32 34 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=0.365 $Y=3.33
+ $X2=0.72 $Y2=3.33
r133 31 58 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=1.075 $Y=3.33
+ $X2=1.21 $Y2=3.33
r134 31 34 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=1.075 $Y=3.33
+ $X2=0.72 $Y2=3.33
r135 29 43 0.802756 $w=4.9e-07 $l=2.88e-06 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=7.92 $Y2=3.33
r136 29 40 0.936549 $w=4.9e-07 $l=3.36e-06 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=1.68 $Y2=3.33
r137 25 64 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=9.39 $Y=3.245
+ $X2=9.39 $Y2=3.33
r138 25 27 36.4172 $w=2.48e-07 $l=7.9e-07 $layer=LI1_cond $X=9.39 $Y=3.245
+ $X2=9.39 $Y2=2.455
r139 21 61 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=8.41 $Y=3.245
+ $X2=8.41 $Y2=3.33
r140 21 23 36.4172 $w=2.48e-07 $l=7.9e-07 $layer=LI1_cond $X=8.41 $Y=3.245
+ $X2=8.41 $Y2=2.455
r141 17 58 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.21 $Y=3.245
+ $X2=1.21 $Y2=3.33
r142 17 19 41.8294 $w=2.68e-07 $l=9.8e-07 $layer=LI1_cond $X=1.21 $Y=3.245
+ $X2=1.21 $Y2=2.265
r143 13 55 3.13335 $w=2.5e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.24 $Y=3.245
+ $X2=0.182 $Y2=3.33
r144 13 15 45.1758 $w=2.48e-07 $l=9.8e-07 $layer=LI1_cond $X=0.24 $Y=3.245
+ $X2=0.24 $Y2=2.265
r145 4 27 300 $w=1.7e-07 $l=6.85912e-07 $layer=licon1_PDIFF $count=2 $X=9.2
+ $Y=1.84 $X2=9.35 $Y2=2.455
r146 3 23 300 $w=1.7e-07 $l=6.85912e-07 $layer=licon1_PDIFF $count=2 $X=8.3
+ $Y=1.84 $X2=8.45 $Y2=2.455
r147 2 19 300 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=2 $X=1.03
+ $Y=2.12 $X2=1.18 $Y2=2.265
r148 1 15 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=2.12 $X2=0.28 $Y2=2.265
.ends

.subckt PM_SKY130_FD_SC_HS__NOR4B_4%A_319_368# 1 2 3 4 5 18 22 23 26 28 30 31 36
+ 41 42 44 45
c64 28 0 9.04372e-20 $X=3.475 $Y=2.99
r65 44 45 5.79692 $w=2.48e-07 $l=1e-07 $layer=LI1_cond $X=5.54 $Y=2.415 $X2=5.44
+ $Y2=2.415
r66 42 45 44.6898 $w=1.68e-07 $l=6.85e-07 $layer=LI1_cond $X=4.755 $Y=2.375
+ $X2=5.44 $Y2=2.375
r67 40 42 8.78489 $w=4.28e-07 $l=1.65e-07 $layer=LI1_cond $X=4.59 $Y=2.505
+ $X2=4.755 $Y2=2.505
r68 40 41 8.78489 $w=4.28e-07 $l=1.65e-07 $layer=LI1_cond $X=4.59 $Y=2.505
+ $X2=4.425 $Y2=2.505
r69 33 38 4.57959 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=3.755 $Y=2.405
+ $X2=3.615 $Y2=2.405
r70 33 41 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.755 $Y=2.405
+ $X2=4.425 $Y2=2.405
r71 30 38 2.78046 $w=2.8e-07 $l=8.5e-08 $layer=LI1_cond $X=3.615 $Y=2.49
+ $X2=3.615 $Y2=2.405
r72 30 31 17.0809 $w=2.78e-07 $l=4.15e-07 $layer=LI1_cond $X=3.615 $Y=2.49
+ $X2=3.615 $Y2=2.905
r73 29 36 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=2.805 $Y=2.99
+ $X2=2.665 $Y2=2.99
r74 28 31 7.36005 $w=1.7e-07 $l=1.77482e-07 $layer=LI1_cond $X=3.475 $Y=2.99
+ $X2=3.615 $Y2=2.905
r75 28 29 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.475 $Y=2.99
+ $X2=2.805 $Y2=2.99
r76 24 36 0.375625 $w=2.8e-07 $l=8.5e-08 $layer=LI1_cond $X=2.665 $Y=2.905
+ $X2=2.665 $Y2=2.99
r77 24 26 23.872 $w=2.78e-07 $l=5.8e-07 $layer=LI1_cond $X=2.665 $Y=2.905
+ $X2=2.665 $Y2=2.325
r78 22 36 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=2.525 $Y=2.99
+ $X2=2.665 $Y2=2.99
r79 22 23 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=2.525 $Y=2.99
+ $X2=1.825 $Y2=2.99
r80 18 21 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=1.7 $Y=1.985 $X2=1.7
+ $Y2=2.815
r81 16 23 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.7 $Y=2.905
+ $X2=1.825 $Y2=2.99
r82 16 21 4.14879 $w=2.48e-07 $l=9e-08 $layer=LI1_cond $X=1.7 $Y=2.905 $X2=1.7
+ $Y2=2.815
r83 5 44 600 $w=1.7e-07 $l=6.05372e-07 $layer=licon1_PDIFF $count=1 $X=5.39
+ $Y=1.84 $X2=5.54 $Y2=2.375
r84 4 40 600 $w=1.7e-07 $l=7.63479e-07 $layer=licon1_PDIFF $count=1 $X=4.39
+ $Y=1.84 $X2=4.59 $Y2=2.51
r85 3 38 300 $w=1.7e-07 $l=7.16083e-07 $layer=licon1_PDIFF $count=2 $X=3.44
+ $Y=1.84 $X2=3.59 $Y2=2.485
r86 2 26 300 $w=1.7e-07 $l=5.63627e-07 $layer=licon1_PDIFF $count=2 $X=2.49
+ $Y=1.84 $X2=2.66 $Y2=2.325
r87 1 21 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=1.595
+ $Y=1.84 $X2=1.74 $Y2=2.815
r88 1 18 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=1.595
+ $Y=1.84 $X2=1.74 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HS__NOR4B_4%Y 1 2 3 4 5 6 7 8 9 10 33 35 36 37 39 41 45
+ 47 51 53 57 59 63 65 66 69 71 75 77 81 83 87 91 94 99 106 107 108 109 110
c204 109 0 1.8401e-19 $X=5.52 $Y=1.295
c205 99 0 1.50238e-20 $X=3.625 $Y=1.095
c206 77 0 7.35572e-20 $X=8.275 $Y=1.095
c207 59 0 5.58611e-20 $X=4.905 $Y=1.095
c208 47 0 1.09607e-20 $X=3.5 $Y=1.385
c209 41 0 1.227e-20 $X=2.975 $Y=1.905
c210 35 0 2.40437e-20 $X=2.5 $Y=1.065
r211 109 110 18.5393 $w=2.28e-07 $l=3.7e-07 $layer=LI1_cond $X=5.52 $Y=1.295
+ $X2=5.52 $Y2=1.665
r212 105 110 14.2803 $w=2.28e-07 $l=2.85e-07 $layer=LI1_cond $X=5.52 $Y=1.95
+ $X2=5.52 $Y2=1.665
r213 104 109 5.76222 $w=2.28e-07 $l=1.15e-07 $layer=LI1_cond $X=5.52 $Y=1.18
+ $X2=5.52 $Y2=1.295
r214 99 100 13.3683 $w=2.48e-07 $l=2.9e-07 $layer=LI1_cond $X=3.625 $Y=1.095
+ $X2=3.625 $Y2=1.385
r215 97 98 2.26996 $w=3.28e-07 $l=6.5e-08 $layer=LI1_cond $X=3.14 $Y=1.97
+ $X2=3.14 $Y2=2.035
r216 94 97 2.26996 $w=3.28e-07 $l=6.5e-08 $layer=LI1_cond $X=3.14 $Y=1.905
+ $X2=3.14 $Y2=1.97
r217 91 92 11.1752 $w=3.28e-07 $l=3.2e-07 $layer=LI1_cond $X=2.665 $Y=1.065
+ $X2=2.665 $Y2=1.385
r218 85 87 22.8184 $w=2.48e-07 $l=4.95e-07 $layer=LI1_cond $X=9.34 $Y=1.01
+ $X2=9.34 $Y2=0.515
r219 84 108 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.525 $Y=1.095
+ $X2=8.4 $Y2=1.095
r220 83 85 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=9.215 $Y=1.095
+ $X2=9.34 $Y2=1.01
r221 83 84 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=9.215 $Y=1.095
+ $X2=8.525 $Y2=1.095
r222 79 108 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=8.4 $Y=1.01
+ $X2=8.4 $Y2=1.095
r223 79 81 22.8184 $w=2.48e-07 $l=4.95e-07 $layer=LI1_cond $X=8.4 $Y=1.01
+ $X2=8.4 $Y2=0.515
r224 78 107 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.58 $Y=1.095
+ $X2=7.415 $Y2=1.095
r225 77 108 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.275 $Y=1.095
+ $X2=8.4 $Y2=1.095
r226 77 78 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=8.275 $Y=1.095
+ $X2=7.58 $Y2=1.095
r227 73 107 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.415 $Y=1.01
+ $X2=7.415 $Y2=1.095
r228 73 75 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=7.415 $Y=1.01
+ $X2=7.415 $Y2=0.515
r229 72 106 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.58 $Y=1.095
+ $X2=6.415 $Y2=1.095
r230 71 107 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.25 $Y=1.095
+ $X2=7.415 $Y2=1.095
r231 71 72 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=7.25 $Y=1.095
+ $X2=6.58 $Y2=1.095
r232 67 106 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.415 $Y=1.01
+ $X2=6.415 $Y2=1.095
r233 67 69 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=6.415 $Y=1.01
+ $X2=6.415 $Y2=0.515
r234 66 104 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=5.635 $Y=1.095
+ $X2=5.52 $Y2=1.095
r235 65 106 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.25 $Y=1.095
+ $X2=6.415 $Y2=1.095
r236 65 66 40.123 $w=1.68e-07 $l=6.15e-07 $layer=LI1_cond $X=6.25 $Y=1.095
+ $X2=5.635 $Y2=1.095
r237 61 104 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=5.07 $Y=1.095
+ $X2=5.52 $Y2=1.095
r238 61 63 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=5.07 $Y=1.01
+ $X2=5.07 $Y2=0.515
r239 60 99 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.75 $Y=1.095
+ $X2=3.625 $Y2=1.095
r240 59 61 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=4.905 $Y=1.095
+ $X2=5.07 $Y2=1.095
r241 59 60 75.3529 $w=1.68e-07 $l=1.155e-06 $layer=LI1_cond $X=4.905 $Y=1.095
+ $X2=3.75 $Y2=1.095
r242 55 99 3.91831 $w=2.48e-07 $l=8.5e-08 $layer=LI1_cond $X=3.625 $Y=1.01
+ $X2=3.625 $Y2=1.095
r243 55 57 22.8184 $w=2.48e-07 $l=4.95e-07 $layer=LI1_cond $X=3.625 $Y=1.01
+ $X2=3.625 $Y2=0.515
r244 54 98 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.305 $Y=2.035
+ $X2=3.14 $Y2=2.035
r245 53 105 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=5.405 $Y=2.035
+ $X2=5.52 $Y2=1.95
r246 53 54 137.005 $w=1.68e-07 $l=2.1e-06 $layer=LI1_cond $X=5.405 $Y=2.035
+ $X2=3.305 $Y2=2.035
r247 49 98 2.96841 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=3.14 $Y=2.12
+ $X2=3.14 $Y2=2.035
r248 49 51 18.5089 $w=3.28e-07 $l=5.3e-07 $layer=LI1_cond $X=3.14 $Y=2.12
+ $X2=3.14 $Y2=2.65
r249 48 92 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.83 $Y=1.385
+ $X2=2.665 $Y2=1.385
r250 47 100 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.5 $Y=1.385
+ $X2=3.625 $Y2=1.385
r251 47 48 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.5 $Y=1.385
+ $X2=2.83 $Y2=1.385
r252 43 91 2.96841 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=2.665 $Y=0.98
+ $X2=2.665 $Y2=1.065
r253 43 45 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=2.665 $Y=0.98
+ $X2=2.665 $Y2=0.515
r254 42 90 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.355 $Y=1.905
+ $X2=2.19 $Y2=1.905
r255 41 94 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.975 $Y=1.905
+ $X2=3.14 $Y2=1.905
r256 41 42 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=2.975 $Y=1.905
+ $X2=2.355 $Y2=1.905
r257 37 90 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.19 $Y=1.99 $X2=2.19
+ $Y2=1.905
r258 37 39 23.0489 $w=3.28e-07 $l=6.6e-07 $layer=LI1_cond $X=2.19 $Y=1.99
+ $X2=2.19 $Y2=2.65
r259 35 91 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.5 $Y=1.065
+ $X2=2.665 $Y2=1.065
r260 35 36 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=2.5 $Y=1.065
+ $X2=1.82 $Y2=1.065
r261 31 36 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.695 $Y=0.98
+ $X2=1.82 $Y2=1.065
r262 31 33 21.4354 $w=2.48e-07 $l=4.65e-07 $layer=LI1_cond $X=1.695 $Y=0.98
+ $X2=1.695 $Y2=0.515
r263 10 97 400 $w=1.7e-07 $l=2.04939e-07 $layer=licon1_PDIFF $count=1 $X=2.99
+ $Y=1.84 $X2=3.14 $Y2=1.97
r264 10 51 400 $w=1.7e-07 $l=8.81816e-07 $layer=licon1_PDIFF $count=1 $X=2.99
+ $Y=1.84 $X2=3.14 $Y2=2.65
r265 9 90 400 $w=1.7e-07 $l=2.04939e-07 $layer=licon1_PDIFF $count=1 $X=2.04
+ $Y=1.84 $X2=2.19 $Y2=1.97
r266 9 39 400 $w=1.7e-07 $l=8.81816e-07 $layer=licon1_PDIFF $count=1 $X=2.04
+ $Y=1.84 $X2=2.19 $Y2=2.65
r267 8 87 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=9.16
+ $Y=0.37 $X2=9.3 $Y2=0.515
r268 7 81 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=8.3
+ $Y=0.37 $X2=8.44 $Y2=0.515
r269 6 75 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=7.275
+ $Y=0.37 $X2=7.415 $Y2=0.515
r270 5 69 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=6.275
+ $Y=0.37 $X2=6.415 $Y2=0.515
r271 4 63 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=4.93
+ $Y=0.37 $X2=5.07 $Y2=0.515
r272 3 57 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.525
+ $Y=0.37 $X2=3.665 $Y2=0.515
r273 2 45 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.525
+ $Y=0.37 $X2=2.665 $Y2=0.515
r274 1 33 91 $w=1.7e-07 $l=2.83373e-07 $layer=licon1_NDIFF $count=2 $X=1.515
+ $Y=0.37 $X2=1.735 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__NOR4B_4%A_778_368# 1 2 3 4 13 15 19 21 25 28 33 37
c60 13 0 7.8278e-20 $X=4.925 $Y=2.99
r61 33 35 7.85757 $w=3.28e-07 $l=2.25e-07 $layer=LI1_cond $X=5.09 $Y=2.765
+ $X2=5.09 $Y2=2.99
r62 28 30 7.33373 $w=3.28e-07 $l=2.1e-07 $layer=LI1_cond $X=4.09 $Y=2.78
+ $X2=4.09 $Y2=2.99
r63 23 25 20.744 $w=2.48e-07 $l=4.5e-07 $layer=LI1_cond $X=7.59 $Y=2.905
+ $X2=7.59 $Y2=2.455
r64 22 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.765 $Y=2.99
+ $X2=6.6 $Y2=2.99
r65 21 23 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=7.465 $Y=2.99
+ $X2=7.59 $Y2=2.905
r66 21 22 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=7.465 $Y=2.99
+ $X2=6.765 $Y2=2.99
r67 17 37 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.6 $Y=2.905 $X2=6.6
+ $Y2=2.99
r68 17 19 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=6.6 $Y=2.905 $X2=6.6
+ $Y2=2.455
r69 16 35 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.255 $Y=2.99
+ $X2=5.09 $Y2=2.99
r70 15 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.435 $Y=2.99
+ $X2=6.6 $Y2=2.99
r71 15 16 76.984 $w=1.68e-07 $l=1.18e-06 $layer=LI1_cond $X=6.435 $Y=2.99
+ $X2=5.255 $Y2=2.99
r72 14 30 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.255 $Y=2.99
+ $X2=4.09 $Y2=2.99
r73 13 35 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.925 $Y=2.99
+ $X2=5.09 $Y2=2.99
r74 13 14 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.925 $Y=2.99
+ $X2=4.255 $Y2=2.99
r75 4 25 300 $w=1.7e-07 $l=6.85912e-07 $layer=licon1_PDIFF $count=2 $X=7.4
+ $Y=1.84 $X2=7.55 $Y2=2.455
r76 3 19 300 $w=1.7e-07 $l=7.07972e-07 $layer=licon1_PDIFF $count=2 $X=6.4
+ $Y=1.84 $X2=6.6 $Y2=2.455
r77 2 33 600 $w=1.7e-07 $l=1.00871e-06 $layer=licon1_PDIFF $count=1 $X=4.915
+ $Y=1.84 $X2=5.09 $Y2=2.765
r78 1 28 600 $w=1.7e-07 $l=1.03518e-06 $layer=licon1_PDIFF $count=1 $X=3.89
+ $Y=1.84 $X2=4.09 $Y2=2.78
.ends

.subckt PM_SKY130_FD_SC_HS__NOR4B_4%A_1191_368# 1 2 3 4 5 18 22 24 28 30 34 36
+ 38 40 43 45 47 49
r71 38 51 3.1514 $w=2.5e-07 $l=1.5e-07 $layer=LI1_cond $X=9.84 $Y=2.12 $X2=9.84
+ $Y2=1.97
r72 38 40 12.9074 $w=2.48e-07 $l=2.8e-07 $layer=LI1_cond $X=9.84 $Y=2.12
+ $X2=9.84 $Y2=2.4
r73 37 49 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.065 $Y=2.035
+ $X2=8.9 $Y2=2.035
r74 36 51 3.99177 $w=1.7e-07 $l=1.5411e-07 $layer=LI1_cond $X=9.715 $Y=2.035
+ $X2=9.84 $Y2=1.97
r75 36 37 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=9.715 $Y=2.035
+ $X2=9.065 $Y2=2.035
r76 32 49 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.9 $Y=2.12 $X2=8.9
+ $Y2=2.035
r77 32 34 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=8.9 $Y=2.12 $X2=8.9
+ $Y2=2.815
r78 31 47 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=8.115 $Y=2.035 $X2=8
+ $Y2=2.035
r79 30 49 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.735 $Y=2.035
+ $X2=8.9 $Y2=2.035
r80 30 31 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=8.735 $Y=2.035
+ $X2=8.115 $Y2=2.035
r81 26 47 0.280307 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8 $Y=2.12 $X2=8
+ $Y2=2.035
r82 26 28 16.034 $w=2.28e-07 $l=3.2e-07 $layer=LI1_cond $X=8 $Y=2.12 $X2=8
+ $Y2=2.44
r83 25 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.265 $Y=2.035
+ $X2=7.1 $Y2=2.035
r84 24 47 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=7.885 $Y=2.035 $X2=8
+ $Y2=2.035
r85 24 25 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=7.885 $Y=2.035
+ $X2=7.265 $Y2=2.035
r86 20 45 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.1 $Y=2.12 $X2=7.1
+ $Y2=2.035
r87 20 22 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=7.1 $Y=2.12 $X2=7.1
+ $Y2=2.57
r88 19 43 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.265 $Y=2.035
+ $X2=6.1 $Y2=2.035
r89 18 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.935 $Y=2.035
+ $X2=7.1 $Y2=2.035
r90 18 19 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=6.935 $Y=2.035
+ $X2=6.265 $Y2=2.035
r91 5 51 600 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=9.65
+ $Y=1.84 $X2=9.8 $Y2=1.985
r92 5 40 300 $w=1.7e-07 $l=6.30555e-07 $layer=licon1_PDIFF $count=2 $X=9.65
+ $Y=1.84 $X2=9.8 $Y2=2.4
r93 4 49 400 $w=1.7e-07 $l=2.59374e-07 $layer=licon1_PDIFF $count=1 $X=8.75
+ $Y=1.84 $X2=8.9 $Y2=2.035
r94 4 34 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=8.75
+ $Y=1.84 $X2=8.9 $Y2=2.815
r95 3 47 600 $w=1.7e-07 $l=2.59374e-07 $layer=licon1_PDIFF $count=1 $X=7.85
+ $Y=1.84 $X2=8 $Y2=2.035
r96 3 28 300 $w=1.7e-07 $l=6.7082e-07 $layer=licon1_PDIFF $count=2 $X=7.85
+ $Y=1.84 $X2=8 $Y2=2.44
r97 2 45 600 $w=1.7e-07 $l=2.81069e-07 $layer=licon1_PDIFF $count=1 $X=6.9
+ $Y=1.84 $X2=7.1 $Y2=2.035
r98 2 22 600 $w=1.7e-07 $l=8.23954e-07 $layer=licon1_PDIFF $count=1 $X=6.9
+ $Y=1.84 $X2=7.1 $Y2=2.57
r99 1 43 300 $w=1.7e-07 $l=2.57488e-07 $layer=licon1_PDIFF $count=2 $X=5.955
+ $Y=1.84 $X2=6.1 $Y2=2.035
.ends

.subckt PM_SKY130_FD_SC_HS__NOR4B_4%VGND 1 2 3 4 5 6 7 8 9 30 34 38 42 46 50 54
+ 56 58 60 62 67 72 77 82 87 92 97 102 108 111 114 126 129 132 135 139
r136 138 139 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.84 $Y=0
+ $X2=9.84 $Y2=0
r137 135 136 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=0
+ $X2=8.88 $Y2=0
r138 132 133 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=0
+ $X2=7.92 $Y2=0
r139 129 130 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=0
+ $X2=6.96 $Y2=0
r140 126 127 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=0
+ $X2=5.52 $Y2=0
r141 119 121 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0
+ $X2=4.56 $Y2=0
r142 114 115 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0
+ $X2=3.12 $Y2=0
r143 111 112 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0
+ $X2=2.16 $Y2=0
r144 108 109 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r145 106 139 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.36 $Y=0
+ $X2=9.84 $Y2=0
r146 106 136 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.36 $Y=0
+ $X2=8.88 $Y2=0
r147 105 106 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.36 $Y=0
+ $X2=9.36 $Y2=0
r148 103 135 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.035 $Y=0
+ $X2=8.87 $Y2=0
r149 103 105 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=9.035 $Y=0
+ $X2=9.36 $Y2=0
r150 102 138 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=9.635 $Y=0
+ $X2=9.857 $Y2=0
r151 102 105 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=9.635 $Y=0
+ $X2=9.36 $Y2=0
r152 101 136 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=0
+ $X2=8.88 $Y2=0
r153 101 133 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=0
+ $X2=7.92 $Y2=0
r154 100 101 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r155 98 132 9.05715 $w=1.7e-07 $l=1.78e-07 $layer=LI1_cond $X=8.105 $Y=0
+ $X2=7.927 $Y2=0
r156 98 100 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=8.105 $Y=0 $X2=8.4
+ $Y2=0
r157 97 135 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.705 $Y=0
+ $X2=8.87 $Y2=0
r158 97 100 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=8.705 $Y=0
+ $X2=8.4 $Y2=0
r159 96 133 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=0
+ $X2=7.92 $Y2=0
r160 96 130 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=0
+ $X2=6.96 $Y2=0
r161 95 96 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=0 $X2=7.44
+ $Y2=0
r162 93 129 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.08 $Y=0
+ $X2=6.915 $Y2=0
r163 93 95 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=7.08 $Y=0 $X2=7.44
+ $Y2=0
r164 92 132 9.05715 $w=1.7e-07 $l=1.77e-07 $layer=LI1_cond $X=7.75 $Y=0
+ $X2=7.927 $Y2=0
r165 92 95 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=7.75 $Y=0 $X2=7.44
+ $Y2=0
r166 91 130 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=0
+ $X2=6.96 $Y2=0
r167 91 127 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.48 $Y=0
+ $X2=5.52 $Y2=0
r168 90 91 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.48 $Y=0 $X2=6.48
+ $Y2=0
r169 88 126 13.399 $w=1.7e-07 $l=3.38e-07 $layer=LI1_cond $X=6.08 $Y=0 $X2=5.742
+ $Y2=0
r170 88 90 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=6.08 $Y=0 $X2=6.48
+ $Y2=0
r171 87 129 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.75 $Y=0
+ $X2=6.915 $Y2=0
r172 87 90 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=6.75 $Y=0 $X2=6.48
+ $Y2=0
r173 83 85 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=4.735 $Y=0
+ $X2=5.04 $Y2=0
r174 82 126 13.399 $w=1.7e-07 $l=3.37e-07 $layer=LI1_cond $X=5.405 $Y=0
+ $X2=5.742 $Y2=0
r175 82 85 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=5.405 $Y=0
+ $X2=5.04 $Y2=0
r176 81 119 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.08
+ $Y2=0
r177 81 115 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=3.12
+ $Y2=0
r178 80 81 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r179 78 114 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.33 $Y=0
+ $X2=3.165 $Y2=0
r180 78 80 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=3.33 $Y=0 $X2=3.6
+ $Y2=0
r181 77 123 10.0292 $w=8.03e-07 $l=6.75e-07 $layer=LI1_cond $X=4.332 $Y=0
+ $X2=4.332 $Y2=0.675
r182 77 83 10.2506 $w=1.7e-07 $l=4.03e-07 $layer=LI1_cond $X=4.332 $Y=0
+ $X2=4.735 $Y2=0
r183 77 121 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r184 77 119 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r185 77 80 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=3.93 $Y=0 $X2=3.6
+ $Y2=0
r186 76 115 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0
+ $X2=3.12 $Y2=0
r187 76 112 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0
+ $X2=2.16 $Y2=0
r188 75 76 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r189 73 111 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.33 $Y=0
+ $X2=2.165 $Y2=0
r190 73 75 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=2.33 $Y=0 $X2=2.64
+ $Y2=0
r191 72 114 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3 $Y=0 $X2=3.165
+ $Y2=0
r192 72 75 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=3 $Y=0 $X2=2.64
+ $Y2=0
r193 71 112 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0
+ $X2=2.16 $Y2=0
r194 71 109 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r195 70 71 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r196 68 108 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.39 $Y=0
+ $X2=1.225 $Y2=0
r197 68 70 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=1.39 $Y=0 $X2=1.68
+ $Y2=0
r198 67 111 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2 $Y=0 $X2=2.165
+ $Y2=0
r199 67 70 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=2 $Y=0 $X2=1.68
+ $Y2=0
r200 65 109 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r201 64 65 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r202 62 108 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.06 $Y=0
+ $X2=1.225 $Y2=0
r203 62 64 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=1.06 $Y=0 $X2=0.72
+ $Y2=0
r204 60 127 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=0
+ $X2=5.52 $Y2=0
r205 60 121 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=0
+ $X2=4.56 $Y2=0
r206 60 85 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r207 56 138 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=9.8 $Y=0.085
+ $X2=9.857 $Y2=0
r208 56 58 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=9.8 $Y=0.085
+ $X2=9.8 $Y2=0.515
r209 52 135 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.87 $Y=0.085
+ $X2=8.87 $Y2=0
r210 52 54 19.382 $w=3.28e-07 $l=5.55e-07 $layer=LI1_cond $X=8.87 $Y=0.085
+ $X2=8.87 $Y2=0.64
r211 48 132 1.11826 $w=3.55e-07 $l=8.5e-08 $layer=LI1_cond $X=7.927 $Y=0.085
+ $X2=7.927 $Y2=0
r212 48 50 18.0171 $w=3.53e-07 $l=5.55e-07 $layer=LI1_cond $X=7.927 $Y=0.085
+ $X2=7.927 $Y2=0.64
r213 44 129 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.915 $Y=0.085
+ $X2=6.915 $Y2=0
r214 44 46 19.382 $w=3.28e-07 $l=5.55e-07 $layer=LI1_cond $X=6.915 $Y=0.085
+ $X2=6.915 $Y2=0.64
r215 40 126 2.78459 $w=6.75e-07 $l=8.5e-08 $layer=LI1_cond $X=5.742 $Y=0.085
+ $X2=5.742 $Y2=0
r216 40 42 10.4546 $w=6.73e-07 $l=5.9e-07 $layer=LI1_cond $X=5.742 $Y=0.085
+ $X2=5.742 $Y2=0.675
r217 36 114 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.165 $Y=0.085
+ $X2=3.165 $Y2=0
r218 36 38 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=3.165 $Y=0.085
+ $X2=3.165 $Y2=0.515
r219 32 111 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.165 $Y=0.085
+ $X2=2.165 $Y2=0
r220 32 34 18.8582 $w=3.28e-07 $l=5.4e-07 $layer=LI1_cond $X=2.165 $Y=0.085
+ $X2=2.165 $Y2=0.625
r221 28 108 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.225 $Y=0.085
+ $X2=1.225 $Y2=0
r222 28 30 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=1.225 $Y=0.085
+ $X2=1.225 $Y2=0.515
r223 9 58 91 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=2 $X=9.59
+ $Y=0.37 $X2=9.8 $Y2=0.515
r224 8 54 182 $w=1.7e-07 $l=3.32716e-07 $layer=licon1_NDIFF $count=1 $X=8.73
+ $Y=0.37 $X2=8.87 $Y2=0.64
r225 7 50 182 $w=1.7e-07 $l=3.63731e-07 $layer=licon1_NDIFF $count=1 $X=7.705
+ $Y=0.37 $X2=7.925 $Y2=0.64
r226 6 46 182 $w=1.7e-07 $l=3.32716e-07 $layer=licon1_NDIFF $count=1 $X=6.775
+ $Y=0.37 $X2=6.915 $Y2=0.64
r227 5 42 91 $w=1.7e-07 $l=7.62398e-07 $layer=licon1_NDIFF $count=2 $X=5.36
+ $Y=0.37 $X2=5.985 $Y2=0.675
r228 4 123 91 $w=1.7e-07 $l=8.23499e-07 $layer=licon1_NDIFF $count=2 $X=3.955
+ $Y=0.37 $X2=4.64 $Y2=0.675
r229 3 38 91 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=2 $X=2.955
+ $Y=0.37 $X2=3.165 $Y2=0.515
r230 2 34 182 $w=1.7e-07 $l=3.17372e-07 $layer=licon1_NDIFF $count=1 $X=2.025
+ $Y=0.37 $X2=2.165 $Y2=0.625
r231 1 30 91 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_NDIFF $count=2 $X=1.07
+ $Y=0.37 $X2=1.225 $Y2=0.515
.ends

