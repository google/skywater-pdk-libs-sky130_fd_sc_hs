* File: sky130_fd_sc_hs__o2bb2a_4.spice
* Created: Thu Aug 27 21:01:06 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hs__o2bb2a_4.pex.spice"
.subckt sky130_fd_sc_hs__o2bb2a_4  VNB VPB B1 B2 A2_N A1_N VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A1_N	A1_N
* A2_N	A2_N
* B2	B2
* B1	B1
* VPB	VPB
* VNB	VNB
MM1022 N_VGND_M1022_d N_B1_M1022_g N_A_27_74#_M1022_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.1344 AS=0.1824 PD=1.06 PS=1.85 NRD=13.116 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75002.7 A=0.096 P=1.58 MULT=1
MM1023 N_VGND_M1022_d N_B1_M1023_g N_A_27_74#_M1023_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.1344 AS=0.0896 PD=1.06 PS=0.92 NRD=13.116 NRS=0 M=1 R=4.26667 SA=75000.8
+ SB=75002.1 A=0.096 P=1.58 MULT=1
MM1004 N_A_27_74#_M1023_s N_B2_M1004_g N_VGND_M1004_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.0896 AS=0.112 PD=0.92 PS=0.99 NRD=0 NRS=13.116 M=1 R=4.26667 SA=75001.2
+ SB=75001.7 A=0.096 P=1.58 MULT=1
MM1006 N_A_27_74#_M1006_d N_B2_M1006_g N_VGND_M1004_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.0992 AS=0.112 PD=0.95 PS=0.99 NRD=2.808 NRS=0 M=1 R=4.26667 SA=75001.7
+ SB=75001.2 A=0.096 P=1.58 MULT=1
MM1001 N_A_27_74#_M1006_d N_A_476_48#_M1001_g N_A_310_392#_M1001_s VNB NLOWVT
+ L=0.15 W=0.64 AD=0.0992 AS=0.1008 PD=0.95 PS=0.955 NRD=2.808 NRS=0 M=1
+ R=4.26667 SA=75002.2 SB=75000.7 A=0.096 P=1.58 MULT=1
MM1020 N_A_27_74#_M1020_d N_A_476_48#_M1020_g N_A_310_392#_M1001_s VNB NLOWVT
+ L=0.15 W=0.64 AD=0.2048 AS=0.1008 PD=1.92 PS=0.955 NRD=6.552 NRS=6.552 M=1
+ R=4.26667 SA=75002.6 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1021 A_835_94# N_A2_N_M1021_g N_A_476_48#_M1021_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.0768 AS=0.1952 PD=0.88 PS=1.89 NRD=12.18 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75002.8 A=0.096 P=1.58 MULT=1
MM1008 N_VGND_M1008_d N_A1_N_M1008_g A_835_94# VNB NLOWVT L=0.15 W=0.64
+ AD=0.157032 AS=0.0768 PD=1.14087 PS=0.88 NRD=19.68 NRS=12.18 M=1 R=4.26667
+ SA=75000.6 SB=75002.4 A=0.096 P=1.58 MULT=1
MM1000 N_X_M1000_d N_A_310_392#_M1000_g N_VGND_M1008_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.15725 AS=0.181568 PD=1.165 PS=1.31913 NRD=12.156 NRS=17.016 M=1 R=4.93333
+ SA=75001.1 SB=75001.8 A=0.111 P=1.78 MULT=1
MM1002 N_X_M1000_d N_A_310_392#_M1002_g N_VGND_M1002_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.15725 AS=0.1295 PD=1.165 PS=1.09 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75001.7
+ SB=75001.2 A=0.111 P=1.78 MULT=1
MM1003 N_X_M1003_d N_A_310_392#_M1003_g N_VGND_M1002_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1295 PD=1.02 PS=1.09 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75002.2
+ SB=75000.7 A=0.111 P=1.78 MULT=1
MM1009 N_X_M1003_d N_A_310_392#_M1009_g N_VGND_M1009_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.2627 PD=1.02 PS=2.19 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75002.6
+ SB=75000.3 A=0.111 P=1.78 MULT=1
MM1007 N_VPWR_M1007_d N_B1_M1007_g N_A_41_392#_M1007_s VPB PSHORT L=0.15 W=1
+ AD=0.15 AS=0.295 PD=1.3 PS=2.59 NRD=1.9503 NRS=1.9503 M=1 R=6.66667 SA=75000.2
+ SB=75001.6 A=0.15 P=2.3 MULT=1
MM1015 N_VPWR_M1007_d N_B1_M1015_g N_A_41_392#_M1015_s VPB PSHORT L=0.15 W=1
+ AD=0.15 AS=0.15 PD=1.3 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=6.66667 SA=75000.7
+ SB=75001.1 A=0.15 P=2.3 MULT=1
MM1017 N_A_310_392#_M1017_d N_B2_M1017_g N_A_41_392#_M1015_s VPB PSHORT L=0.15
+ W=1 AD=0.15 AS=0.15 PD=1.3 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=6.66667
+ SA=75001.1 SB=75000.7 A=0.15 P=2.3 MULT=1
MM1019 N_A_310_392#_M1017_d N_B2_M1019_g N_A_41_392#_M1019_s VPB PSHORT L=0.15
+ W=1 AD=0.15 AS=0.295 PD=1.3 PS=2.59 NRD=1.9503 NRS=1.9503 M=1 R=6.66667
+ SA=75001.6 SB=75000.2 A=0.15 P=2.3 MULT=1
MM1010 N_A_310_392#_M1010_d N_A_476_48#_M1010_g N_VPWR_M1010_s VPB PSHORT L=0.15
+ W=0.84 AD=0.1554 AS=0.2478 PD=1.21 PS=2.27 NRD=3.5066 NRS=2.3443 M=1 R=5.6
+ SA=75000.2 SB=75004 A=0.126 P=1.98 MULT=1
MM1011 N_A_310_392#_M1010_d N_A_476_48#_M1011_g N_VPWR_M1011_s VPB PSHORT L=0.15
+ W=0.84 AD=0.1554 AS=0.2583 PD=1.21 PS=1.73 NRD=17.5724 NRS=59.1985 M=1 R=5.6
+ SA=75000.7 SB=75003.5 A=0.126 P=1.98 MULT=1
MM1014 N_A_476_48#_M1014_d N_A2_N_M1014_g N_VPWR_M1011_s VPB PSHORT L=0.15
+ W=0.84 AD=0.126 AS=0.2583 PD=1.14 PS=1.73 NRD=2.3443 NRS=59.1985 M=1 R=5.6
+ SA=75001.4 SB=75002.8 A=0.126 P=1.98 MULT=1
MM1018 N_VPWR_M1018_d N_A1_N_M1018_g N_A_476_48#_M1014_d VPB PSHORT L=0.15
+ W=0.84 AD=0.2322 AS=0.126 PD=1.48286 PS=1.14 NRD=51.9292 NRS=2.3443 M=1 R=5.6
+ SA=75001.8 SB=75002.4 A=0.126 P=1.98 MULT=1
MM1005 N_VPWR_M1018_d N_A_310_392#_M1005_g N_X_M1005_s VPB PSHORT L=0.15 W=1.12
+ AD=0.3096 AS=0.224 PD=1.97714 PS=1.52 NRD=17.5724 NRS=10.5395 M=1 R=7.46667
+ SA=75001.9 SB=75001.8 A=0.168 P=2.54 MULT=1
MM1012 N_VPWR_M1012_d N_A_310_392#_M1012_g N_X_M1005_s VPB PSHORT L=0.15 W=1.12
+ AD=0.196 AS=0.224 PD=1.47 PS=1.52 NRD=1.7533 NRS=10.5395 M=1 R=7.46667
+ SA=75002.4 SB=75001.2 A=0.168 P=2.54 MULT=1
MM1013 N_VPWR_M1012_d N_A_310_392#_M1013_g N_X_M1013_s VPB PSHORT L=0.15 W=1.12
+ AD=0.196 AS=0.1708 PD=1.47 PS=1.425 NRD=10.5395 NRS=1.7533 M=1 R=7.46667
+ SA=75002.9 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1016 N_VPWR_M1016_d N_A_310_392#_M1016_g N_X_M1013_s VPB PSHORT L=0.15 W=1.12
+ AD=0.3808 AS=0.1708 PD=2.92 PS=1.425 NRD=9.6727 NRS=2.6201 M=1 R=7.46667
+ SA=75003.4 SB=75000.3 A=0.168 P=2.54 MULT=1
DX24_noxref VNB VPB NWDIODE A=14.0988 P=18.88
c_68 VNB 0 1.74227e-19 $X=0 $Y=0
c_934 A_835_94# 0 2.65681e-20 $X=4.175 $Y=0.47
*
.include "sky130_fd_sc_hs__o2bb2a_4.pxi.spice"
*
.ends
*
*
