* File: sky130_fd_sc_hs__ebufn_2.pxi.spice
* Created: Tue Sep  1 20:04:03 2020
* 
x_PM_SKY130_FD_SC_HS__EBUFN_2%A_84_48# N_A_84_48#_M1001_d N_A_84_48#_M1002_d
+ N_A_84_48#_M1009_g N_A_84_48#_c_86_n N_A_84_48#_M1004_g N_A_84_48#_M1010_g
+ N_A_84_48#_c_87_n N_A_84_48#_M1005_g N_A_84_48#_c_81_n N_A_84_48#_c_88_n
+ N_A_84_48#_c_89_n N_A_84_48#_c_108_p N_A_84_48#_c_82_n N_A_84_48#_c_90_n
+ N_A_84_48#_c_83_n N_A_84_48#_c_91_n N_A_84_48#_c_84_n N_A_84_48#_c_85_n
+ PM_SKY130_FD_SC_HS__EBUFN_2%A_84_48#
x_PM_SKY130_FD_SC_HS__EBUFN_2%A_283_48# N_A_283_48#_M1011_s N_A_283_48#_M1006_s
+ N_A_283_48#_c_191_n N_A_283_48#_M1007_g N_A_283_48#_c_192_n
+ N_A_283_48#_c_193_n N_A_283_48#_c_194_n N_A_283_48#_M1008_g
+ N_A_283_48#_c_195_n N_A_283_48#_c_196_n N_A_283_48#_c_197_n
+ N_A_283_48#_c_201_n N_A_283_48#_c_202_n N_A_283_48#_c_198_n
+ N_A_283_48#_c_199_n PM_SKY130_FD_SC_HS__EBUFN_2%A_283_48#
x_PM_SKY130_FD_SC_HS__EBUFN_2%TE_B N_TE_B_c_270_n N_TE_B_M1000_g N_TE_B_c_263_n
+ N_TE_B_c_264_n N_TE_B_c_273_n N_TE_B_M1003_g N_TE_B_c_265_n N_TE_B_c_266_n
+ N_TE_B_M1006_g N_TE_B_M1011_g N_TE_B_c_268_n TE_B
+ PM_SKY130_FD_SC_HS__EBUFN_2%TE_B
x_PM_SKY130_FD_SC_HS__EBUFN_2%A N_A_M1001_g N_A_c_349_n N_A_M1002_g A
+ N_A_c_350_n PM_SKY130_FD_SC_HS__EBUFN_2%A
x_PM_SKY130_FD_SC_HS__EBUFN_2%A_33_368# N_A_33_368#_M1004_d N_A_33_368#_M1005_d
+ N_A_33_368#_M1003_d N_A_33_368#_c_379_n N_A_33_368#_c_380_n
+ N_A_33_368#_c_381_n N_A_33_368#_c_390_n N_A_33_368#_c_382_n
+ N_A_33_368#_c_383_n PM_SKY130_FD_SC_HS__EBUFN_2%A_33_368#
x_PM_SKY130_FD_SC_HS__EBUFN_2%Z N_Z_M1009_d N_Z_M1004_s N_Z_c_428_n N_Z_c_423_n
+ N_Z_c_435_n N_Z_c_424_n N_Z_c_426_n Z Z PM_SKY130_FD_SC_HS__EBUFN_2%Z
x_PM_SKY130_FD_SC_HS__EBUFN_2%VPWR N_VPWR_M1000_s N_VPWR_M1006_d N_VPWR_c_464_n
+ VPWR N_VPWR_c_465_n N_VPWR_c_466_n N_VPWR_c_467_n N_VPWR_c_463_n
+ N_VPWR_c_469_n N_VPWR_c_470_n PM_SKY130_FD_SC_HS__EBUFN_2%VPWR
x_PM_SKY130_FD_SC_HS__EBUFN_2%A_27_74# N_A_27_74#_M1009_s N_A_27_74#_M1010_s
+ N_A_27_74#_M1008_s N_A_27_74#_c_510_n N_A_27_74#_c_511_n N_A_27_74#_c_512_n
+ N_A_27_74#_c_513_n N_A_27_74#_c_514_n N_A_27_74#_c_515_n
+ PM_SKY130_FD_SC_HS__EBUFN_2%A_27_74#
x_PM_SKY130_FD_SC_HS__EBUFN_2%VGND N_VGND_M1007_d N_VGND_M1011_d N_VGND_c_551_n
+ N_VGND_c_552_n N_VGND_c_553_n N_VGND_c_554_n VGND N_VGND_c_555_n
+ N_VGND_c_556_n N_VGND_c_557_n N_VGND_c_558_n PM_SKY130_FD_SC_HS__EBUFN_2%VGND
cc_1 VNB N_A_84_48#_M1009_g 0.0267131f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_2 VNB N_A_84_48#_M1010_g 0.0219916f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=0.74
cc_3 VNB N_A_84_48#_c_81_n 0.006822f $X=-0.19 $Y=-0.245 $X2=1.965 $Y2=1.465
cc_4 VNB N_A_84_48#_c_82_n 0.0227309f $X=-0.19 $Y=-0.245 $X2=4.005 $Y2=0.515
cc_5 VNB N_A_84_48#_c_83_n 0.0131174f $X=-0.19 $Y=-0.245 $X2=4.022 $Y2=1.03
cc_6 VNB N_A_84_48#_c_84_n 0.0300599f $X=-0.19 $Y=-0.245 $X2=4.04 $Y2=1.95
cc_7 VNB N_A_84_48#_c_85_n 0.077667f $X=-0.19 $Y=-0.245 $X2=1.035 $Y2=1.532
cc_8 VNB N_A_283_48#_c_191_n 0.0157819f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.3
cc_9 VNB N_A_283_48#_c_192_n 0.0100196f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_283_48#_c_193_n 0.00785843f $X=-0.19 $Y=-0.245 $X2=0.535 $Y2=1.765
cc_11 VNB N_A_283_48#_c_194_n 0.0180733f $X=-0.19 $Y=-0.245 $X2=0.535 $Y2=2.4
cc_12 VNB N_A_283_48#_c_195_n 0.0317356f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=0.74
cc_13 VNB N_A_283_48#_c_196_n 0.00411221f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_283_48#_c_197_n 0.00429685f $X=-0.19 $Y=-0.245 $X2=1.04 $Y2=1.465
cc_15 VNB N_A_283_48#_c_198_n 0.0713883f $X=-0.19 $Y=-0.245 $X2=4.022 $Y2=0.848
cc_16 VNB N_A_283_48#_c_199_n 0.0105673f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_TE_B_c_263_n 0.00903142f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_TE_B_c_264_n 0.00498176f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_TE_B_c_265_n 0.0199833f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_20 VNB N_TE_B_c_266_n 0.0296471f $X=-0.19 $Y=-0.245 $X2=0.535 $Y2=1.765
cc_21 VNB N_TE_B_M1011_g 0.0337994f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=0.74
cc_22 VNB N_TE_B_c_268_n 0.0044442f $X=-0.19 $Y=-0.245 $X2=1.035 $Y2=1.765
cc_23 VNB TE_B 0.00265516f $X=-0.19 $Y=-0.245 $X2=1.035 $Y2=2.4
cc_24 VNB N_A_M1001_g 0.0382437f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_c_349_n 0.0294725f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_c_350_n 0.00603075f $X=-0.19 $Y=-0.245 $X2=0.535 $Y2=2.4
cc_27 VNB N_Z_c_423_n 0.00143713f $X=-0.19 $Y=-0.245 $X2=0.535 $Y2=2.4
cc_28 VNB N_Z_c_424_n 0.00185767f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_VPWR_c_463_n 0.183584f $X=-0.19 $Y=-0.245 $X2=2.135 $Y2=2.325
cc_30 VNB N_A_27_74#_c_510_n 0.0362285f $X=-0.19 $Y=-0.245 $X2=0.535 $Y2=2.4
cc_31 VNB N_A_27_74#_c_511_n 0.00655758f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=1.3
cc_32 VNB N_A_27_74#_c_512_n 0.00931596f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=0.74
cc_33 VNB N_A_27_74#_c_513_n 0.00423028f $X=-0.19 $Y=-0.245 $X2=1.035 $Y2=2.4
cc_34 VNB N_A_27_74#_c_514_n 0.00276453f $X=-0.19 $Y=-0.245 $X2=1.965 $Y2=1.465
cc_35 VNB N_A_27_74#_c_515_n 0.00206817f $X=-0.19 $Y=-0.245 $X2=1.04 $Y2=1.465
cc_36 VNB N_VGND_c_551_n 0.00563933f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_37 VNB N_VGND_c_552_n 0.0167127f $X=-0.19 $Y=-0.245 $X2=0.535 $Y2=2.4
cc_38 VNB N_VGND_c_553_n 0.0408183f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=0.74
cc_39 VNB N_VGND_c_554_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_555_n 0.039031f $X=-0.19 $Y=-0.245 $X2=1.035 $Y2=2.4
cc_41 VNB N_VGND_c_556_n 0.0199919f $X=-0.19 $Y=-0.245 $X2=4.04 $Y2=2.715
cc_42 VNB N_VGND_c_557_n 0.261479f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_558_n 0.00462376f $X=-0.19 $Y=-0.245 $X2=4.022 $Y2=1.03
cc_44 VPB N_A_84_48#_c_86_n 0.0189714f $X=-0.19 $Y=1.66 $X2=0.535 $Y2=1.765
cc_45 VPB N_A_84_48#_c_87_n 0.0152312f $X=-0.19 $Y=1.66 $X2=1.035 $Y2=1.765
cc_46 VPB N_A_84_48#_c_88_n 0.0011045f $X=-0.19 $Y=1.66 $X2=2.05 $Y2=2.24
cc_47 VPB N_A_84_48#_c_89_n 0.0124138f $X=-0.19 $Y=1.66 $X2=3.875 $Y2=2.325
cc_48 VPB N_A_84_48#_c_90_n 0.0204176f $X=-0.19 $Y=1.66 $X2=4.04 $Y2=2.715
cc_49 VPB N_A_84_48#_c_91_n 0.0174668f $X=-0.19 $Y=1.66 $X2=4.04 $Y2=2.035
cc_50 VPB N_A_84_48#_c_84_n 0.012594f $X=-0.19 $Y=1.66 $X2=4.04 $Y2=1.95
cc_51 VPB N_A_84_48#_c_85_n 0.0163843f $X=-0.19 $Y=1.66 $X2=1.035 $Y2=1.532
cc_52 VPB N_A_283_48#_c_197_n 0.00180087f $X=-0.19 $Y=1.66 $X2=1.04 $Y2=1.465
cc_53 VPB N_A_283_48#_c_201_n 0.00323268f $X=-0.19 $Y=1.66 $X2=1.04 $Y2=1.465
cc_54 VPB N_A_283_48#_c_202_n 0.00410054f $X=-0.19 $Y=1.66 $X2=2.05 $Y2=1.63
cc_55 VPB N_TE_B_c_270_n 0.0164274f $X=-0.19 $Y=1.66 $X2=3.865 $Y2=0.37
cc_56 VPB N_TE_B_c_263_n 0.0174936f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_57 VPB N_TE_B_c_264_n 0.00581755f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_58 VPB N_TE_B_c_273_n 0.0201064f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_59 VPB N_TE_B_c_265_n 0.0237703f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.74
cc_60 VPB N_TE_B_c_266_n 0.0290366f $X=-0.19 $Y=1.66 $X2=0.535 $Y2=1.765
cc_61 VPB N_TE_B_c_268_n 0.00450932f $X=-0.19 $Y=1.66 $X2=1.035 $Y2=1.765
cc_62 VPB N_A_c_349_n 0.0328271f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_63 VPB N_A_c_350_n 0.00490976f $X=-0.19 $Y=1.66 $X2=0.535 $Y2=2.4
cc_64 VPB N_A_33_368#_c_379_n 0.0297839f $X=-0.19 $Y=1.66 $X2=0.535 $Y2=2.4
cc_65 VPB N_A_33_368#_c_380_n 0.00297668f $X=-0.19 $Y=1.66 $X2=0.925 $Y2=1.3
cc_66 VPB N_A_33_368#_c_381_n 0.00983167f $X=-0.19 $Y=1.66 $X2=0.925 $Y2=0.74
cc_67 VPB N_A_33_368#_c_382_n 0.00249658f $X=-0.19 $Y=1.66 $X2=1.035 $Y2=2.4
cc_68 VPB N_A_33_368#_c_383_n 0.0092325f $X=-0.19 $Y=1.66 $X2=1.04 $Y2=1.465
cc_69 VPB N_Z_c_423_n 9.10919e-19 $X=-0.19 $Y=1.66 $X2=0.535 $Y2=2.4
cc_70 VPB N_Z_c_426_n 0.00202983f $X=-0.19 $Y=1.66 $X2=1.035 $Y2=2.4
cc_71 VPB Z 0.00417138f $X=-0.19 $Y=1.66 $X2=1.04 $Y2=1.465
cc_72 VPB N_VPWR_c_464_n 0.0191795f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.74
cc_73 VPB N_VPWR_c_465_n 0.0416792f $X=-0.19 $Y=1.66 $X2=0.535 $Y2=2.4
cc_74 VPB N_VPWR_c_466_n 0.0350409f $X=-0.19 $Y=1.66 $X2=1.035 $Y2=1.765
cc_75 VPB N_VPWR_c_467_n 0.0196898f $X=-0.19 $Y=1.66 $X2=3.875 $Y2=2.325
cc_76 VPB N_VPWR_c_463_n 0.0897536f $X=-0.19 $Y=1.66 $X2=2.135 $Y2=2.325
cc_77 VPB N_VPWR_c_469_n 0.0138344f $X=-0.19 $Y=1.66 $X2=4.005 $Y2=0.515
cc_78 VPB N_VPWR_c_470_n 0.00920679f $X=-0.19 $Y=1.66 $X2=4.12 $Y2=1.95
cc_79 N_A_84_48#_c_89_n N_A_283_48#_M1006_s 0.0124149f $X=3.875 $Y=2.325 $X2=0
+ $Y2=0
cc_80 N_A_84_48#_M1010_g N_A_283_48#_c_191_n 0.025089f $X=0.925 $Y=0.74 $X2=0
+ $Y2=0
cc_81 N_A_84_48#_c_81_n N_A_283_48#_c_192_n 0.00720366f $X=1.965 $Y=1.465 $X2=0
+ $Y2=0
cc_82 N_A_84_48#_c_81_n N_A_283_48#_c_193_n 0.00475854f $X=1.965 $Y=1.465 $X2=0
+ $Y2=0
cc_83 N_A_84_48#_c_85_n N_A_283_48#_c_193_n 0.00230752f $X=1.035 $Y=1.532 $X2=0
+ $Y2=0
cc_84 N_A_84_48#_c_81_n N_A_283_48#_c_195_n 0.00411929f $X=1.965 $Y=1.465 $X2=0
+ $Y2=0
cc_85 N_A_84_48#_c_81_n N_A_283_48#_c_196_n 0.00414715f $X=1.965 $Y=1.465 $X2=0
+ $Y2=0
cc_86 N_A_84_48#_c_81_n N_A_283_48#_c_197_n 0.0208807f $X=1.965 $Y=1.465 $X2=0
+ $Y2=0
cc_87 N_A_84_48#_c_88_n N_A_283_48#_c_197_n 0.00998417f $X=2.05 $Y=2.24 $X2=0
+ $Y2=0
cc_88 N_A_84_48#_c_88_n N_A_283_48#_c_201_n 0.0143326f $X=2.05 $Y=2.24 $X2=0
+ $Y2=0
cc_89 N_A_84_48#_c_89_n N_A_283_48#_c_201_n 0.0274686f $X=3.875 $Y=2.325 $X2=0
+ $Y2=0
cc_90 N_A_84_48#_c_89_n N_A_283_48#_c_202_n 0.0242025f $X=3.875 $Y=2.325 $X2=0
+ $Y2=0
cc_91 N_A_84_48#_c_87_n N_TE_B_c_270_n 0.0309437f $X=1.035 $Y=1.765 $X2=-0.19
+ $Y2=-0.245
cc_92 N_A_84_48#_c_88_n N_TE_B_c_270_n 0.00308504f $X=2.05 $Y=2.24 $X2=-0.19
+ $Y2=-0.245
cc_93 N_A_84_48#_c_108_p N_TE_B_c_270_n 0.0027244f $X=2.135 $Y=2.325 $X2=-0.19
+ $Y2=-0.245
cc_94 N_A_84_48#_c_81_n N_TE_B_c_263_n 0.0148711f $X=1.965 $Y=1.465 $X2=0 $Y2=0
cc_95 N_A_84_48#_c_88_n N_TE_B_c_263_n 0.00713319f $X=2.05 $Y=2.24 $X2=0 $Y2=0
cc_96 N_A_84_48#_c_81_n N_TE_B_c_264_n 0.0057255f $X=1.965 $Y=1.465 $X2=0 $Y2=0
cc_97 N_A_84_48#_c_88_n N_TE_B_c_264_n 7.29731e-19 $X=2.05 $Y=2.24 $X2=0 $Y2=0
cc_98 N_A_84_48#_c_85_n N_TE_B_c_264_n 0.00982968f $X=1.035 $Y=1.532 $X2=0 $Y2=0
cc_99 N_A_84_48#_c_88_n N_TE_B_c_273_n 0.0166373f $X=2.05 $Y=2.24 $X2=0 $Y2=0
cc_100 N_A_84_48#_c_89_n N_TE_B_c_273_n 0.0108355f $X=3.875 $Y=2.325 $X2=0 $Y2=0
cc_101 N_A_84_48#_c_108_p N_TE_B_c_273_n 0.00339691f $X=2.135 $Y=2.325 $X2=0
+ $Y2=0
cc_102 N_A_84_48#_c_89_n N_TE_B_c_265_n 0.00456525f $X=3.875 $Y=2.325 $X2=0
+ $Y2=0
cc_103 N_A_84_48#_c_89_n N_TE_B_c_266_n 0.0191734f $X=3.875 $Y=2.325 $X2=0 $Y2=0
cc_104 N_A_84_48#_c_91_n N_TE_B_c_266_n 0.00218744f $X=4.04 $Y=2.035 $X2=0 $Y2=0
cc_105 N_A_84_48#_c_82_n N_TE_B_M1011_g 2.21897e-19 $X=4.005 $Y=0.515 $X2=0
+ $Y2=0
cc_106 N_A_84_48#_c_81_n N_TE_B_c_268_n 0.00209232f $X=1.965 $Y=1.465 $X2=0
+ $Y2=0
cc_107 N_A_84_48#_c_88_n N_TE_B_c_268_n 0.0036274f $X=2.05 $Y=2.24 $X2=0 $Y2=0
cc_108 N_A_84_48#_c_89_n TE_B 0.00432473f $X=3.875 $Y=2.325 $X2=0 $Y2=0
cc_109 N_A_84_48#_c_82_n N_A_M1001_g 0.00575762f $X=4.005 $Y=0.515 $X2=0 $Y2=0
cc_110 N_A_84_48#_c_83_n N_A_M1001_g 0.00293996f $X=4.022 $Y=1.03 $X2=0 $Y2=0
cc_111 N_A_84_48#_c_84_n N_A_M1001_g 0.009227f $X=4.04 $Y=1.95 $X2=0 $Y2=0
cc_112 N_A_84_48#_c_89_n N_A_c_349_n 0.0155156f $X=3.875 $Y=2.325 $X2=0 $Y2=0
cc_113 N_A_84_48#_c_90_n N_A_c_349_n 0.00714186f $X=4.04 $Y=2.715 $X2=0 $Y2=0
cc_114 N_A_84_48#_c_83_n N_A_c_349_n 0.00160204f $X=4.022 $Y=1.03 $X2=0 $Y2=0
cc_115 N_A_84_48#_c_91_n N_A_c_349_n 0.00743535f $X=4.04 $Y=2.035 $X2=0 $Y2=0
cc_116 N_A_84_48#_c_84_n N_A_c_349_n 0.0131625f $X=4.04 $Y=1.95 $X2=0 $Y2=0
cc_117 N_A_84_48#_c_89_n N_A_c_350_n 0.0130245f $X=3.875 $Y=2.325 $X2=0 $Y2=0
cc_118 N_A_84_48#_c_83_n N_A_c_350_n 0.00112892f $X=4.022 $Y=1.03 $X2=0 $Y2=0
cc_119 N_A_84_48#_c_84_n N_A_c_350_n 0.0326295f $X=4.04 $Y=1.95 $X2=0 $Y2=0
cc_120 N_A_84_48#_c_89_n N_A_33_368#_M1003_d 0.00650959f $X=3.875 $Y=2.325 $X2=0
+ $Y2=0
cc_121 N_A_84_48#_c_86_n N_A_33_368#_c_379_n 0.0130723f $X=0.535 $Y=1.765 $X2=0
+ $Y2=0
cc_122 N_A_84_48#_c_87_n N_A_33_368#_c_379_n 2.69714e-19 $X=1.035 $Y=1.765 $X2=0
+ $Y2=0
cc_123 N_A_84_48#_c_86_n N_A_33_368#_c_380_n 0.011054f $X=0.535 $Y=1.765 $X2=0
+ $Y2=0
cc_124 N_A_84_48#_c_87_n N_A_33_368#_c_380_n 0.0126666f $X=1.035 $Y=1.765 $X2=0
+ $Y2=0
cc_125 N_A_84_48#_c_86_n N_A_33_368#_c_381_n 0.00262934f $X=0.535 $Y=1.765 $X2=0
+ $Y2=0
cc_126 N_A_84_48#_c_89_n N_A_33_368#_c_390_n 0.00538854f $X=3.875 $Y=2.325 $X2=0
+ $Y2=0
cc_127 N_A_84_48#_c_108_p N_A_33_368#_c_390_n 0.00878738f $X=2.135 $Y=2.325
+ $X2=0 $Y2=0
cc_128 N_A_84_48#_c_87_n N_A_33_368#_c_382_n 5.05939e-19 $X=1.035 $Y=1.765 $X2=0
+ $Y2=0
cc_129 N_A_84_48#_c_108_p N_A_33_368#_c_382_n 0.00326713f $X=2.135 $Y=2.325
+ $X2=0 $Y2=0
cc_130 N_A_84_48#_c_89_n N_A_33_368#_c_383_n 0.0211124f $X=3.875 $Y=2.325 $X2=0
+ $Y2=0
cc_131 N_A_84_48#_M1009_g N_Z_c_428_n 0.00439897f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_132 N_A_84_48#_M1010_g N_Z_c_428_n 0.00388974f $X=0.925 $Y=0.74 $X2=0 $Y2=0
cc_133 N_A_84_48#_M1009_g N_Z_c_423_n 0.00866774f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_134 N_A_84_48#_c_86_n N_Z_c_423_n 0.0021572f $X=0.535 $Y=1.765 $X2=0 $Y2=0
cc_135 N_A_84_48#_M1010_g N_Z_c_423_n 0.0025553f $X=0.925 $Y=0.74 $X2=0 $Y2=0
cc_136 N_A_84_48#_c_81_n N_Z_c_423_n 0.0249855f $X=1.965 $Y=1.465 $X2=0 $Y2=0
cc_137 N_A_84_48#_c_85_n N_Z_c_423_n 0.0349907f $X=1.035 $Y=1.532 $X2=0 $Y2=0
cc_138 N_A_84_48#_c_87_n N_Z_c_435_n 0.00727827f $X=1.035 $Y=1.765 $X2=0 $Y2=0
cc_139 N_A_84_48#_M1009_g N_Z_c_424_n 0.00379299f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_140 N_A_84_48#_M1010_g N_Z_c_424_n 0.00421865f $X=0.925 $Y=0.74 $X2=0 $Y2=0
cc_141 N_A_84_48#_c_85_n N_Z_c_424_n 0.00161894f $X=1.035 $Y=1.532 $X2=0 $Y2=0
cc_142 N_A_84_48#_c_86_n N_Z_c_426_n 0.0149681f $X=0.535 $Y=1.765 $X2=0 $Y2=0
cc_143 N_A_84_48#_c_87_n N_Z_c_426_n 0.00123972f $X=1.035 $Y=1.765 $X2=0 $Y2=0
cc_144 N_A_84_48#_c_81_n N_Z_c_426_n 0.0083655f $X=1.965 $Y=1.465 $X2=0 $Y2=0
cc_145 N_A_84_48#_c_85_n N_Z_c_426_n 0.00798369f $X=1.035 $Y=1.532 $X2=0 $Y2=0
cc_146 N_A_84_48#_c_87_n Z 0.0175719f $X=1.035 $Y=1.765 $X2=0 $Y2=0
cc_147 N_A_84_48#_c_81_n Z 0.0649368f $X=1.965 $Y=1.465 $X2=0 $Y2=0
cc_148 N_A_84_48#_c_88_n Z 0.0284331f $X=2.05 $Y=2.24 $X2=0 $Y2=0
cc_149 N_A_84_48#_c_85_n Z 0.00225694f $X=1.035 $Y=1.532 $X2=0 $Y2=0
cc_150 N_A_84_48#_c_88_n N_VPWR_M1000_s 0.00398828f $X=2.05 $Y=2.24 $X2=-0.19
+ $Y2=-0.245
cc_151 N_A_84_48#_c_108_p N_VPWR_M1000_s 0.00324468f $X=2.135 $Y=2.325 $X2=-0.19
+ $Y2=-0.245
cc_152 N_A_84_48#_c_89_n N_VPWR_M1006_d 0.0159751f $X=3.875 $Y=2.325 $X2=0 $Y2=0
cc_153 N_A_84_48#_c_89_n N_VPWR_c_464_n 0.0287575f $X=3.875 $Y=2.325 $X2=0 $Y2=0
cc_154 N_A_84_48#_c_90_n N_VPWR_c_464_n 0.0102171f $X=4.04 $Y=2.715 $X2=0 $Y2=0
cc_155 N_A_84_48#_c_86_n N_VPWR_c_465_n 0.00278257f $X=0.535 $Y=1.765 $X2=0
+ $Y2=0
cc_156 N_A_84_48#_c_87_n N_VPWR_c_465_n 0.00278271f $X=1.035 $Y=1.765 $X2=0
+ $Y2=0
cc_157 N_A_84_48#_c_90_n N_VPWR_c_467_n 0.0097982f $X=4.04 $Y=2.715 $X2=0 $Y2=0
cc_158 N_A_84_48#_c_86_n N_VPWR_c_463_n 0.00357873f $X=0.535 $Y=1.765 $X2=0
+ $Y2=0
cc_159 N_A_84_48#_c_87_n N_VPWR_c_463_n 0.00354798f $X=1.035 $Y=1.765 $X2=0
+ $Y2=0
cc_160 N_A_84_48#_c_90_n N_VPWR_c_463_n 0.0111907f $X=4.04 $Y=2.715 $X2=0 $Y2=0
cc_161 N_A_84_48#_M1009_g N_A_27_74#_c_510_n 0.0015901f $X=0.495 $Y=0.74 $X2=0
+ $Y2=0
cc_162 N_A_84_48#_M1009_g N_A_27_74#_c_511_n 0.0129836f $X=0.495 $Y=0.74 $X2=0
+ $Y2=0
cc_163 N_A_84_48#_M1010_g N_A_27_74#_c_511_n 0.013442f $X=0.925 $Y=0.74 $X2=0
+ $Y2=0
cc_164 N_A_84_48#_c_81_n N_A_27_74#_c_513_n 0.0582054f $X=1.965 $Y=1.465 $X2=0
+ $Y2=0
cc_165 N_A_84_48#_M1010_g N_A_27_74#_c_514_n 0.00109932f $X=0.925 $Y=0.74 $X2=0
+ $Y2=0
cc_166 N_A_84_48#_c_81_n N_A_27_74#_c_514_n 0.0285318f $X=1.965 $Y=1.465 $X2=0
+ $Y2=0
cc_167 N_A_84_48#_c_85_n N_A_27_74#_c_514_n 0.00400839f $X=1.035 $Y=1.532 $X2=0
+ $Y2=0
cc_168 N_A_84_48#_M1010_g N_VGND_c_551_n 2.65335e-19 $X=0.925 $Y=0.74 $X2=0
+ $Y2=0
cc_169 N_A_84_48#_c_82_n N_VGND_c_552_n 0.0259022f $X=4.005 $Y=0.515 $X2=0 $Y2=0
cc_170 N_A_84_48#_M1009_g N_VGND_c_555_n 0.00278271f $X=0.495 $Y=0.74 $X2=0
+ $Y2=0
cc_171 N_A_84_48#_M1010_g N_VGND_c_555_n 0.00278271f $X=0.925 $Y=0.74 $X2=0
+ $Y2=0
cc_172 N_A_84_48#_c_82_n N_VGND_c_556_n 0.0161257f $X=4.005 $Y=0.515 $X2=0 $Y2=0
cc_173 N_A_84_48#_M1009_g N_VGND_c_557_n 0.00357086f $X=0.495 $Y=0.74 $X2=0
+ $Y2=0
cc_174 N_A_84_48#_M1010_g N_VGND_c_557_n 0.00354644f $X=0.925 $Y=0.74 $X2=0
+ $Y2=0
cc_175 N_A_84_48#_c_82_n N_VGND_c_557_n 0.013291f $X=4.005 $Y=0.515 $X2=0 $Y2=0
cc_176 N_A_283_48#_c_192_n N_TE_B_c_263_n 0.0180315f $X=1.85 $Y=1.26 $X2=0 $Y2=0
cc_177 N_A_283_48#_c_193_n N_TE_B_c_264_n 0.0180315f $X=1.565 $Y=1.26 $X2=0
+ $Y2=0
cc_178 N_A_283_48#_c_197_n N_TE_B_c_273_n 0.0011225f $X=2.56 $Y=1.17 $X2=0 $Y2=0
cc_179 N_A_283_48#_c_201_n N_TE_B_c_273_n 0.00538263f $X=2.725 $Y=1.945 $X2=0
+ $Y2=0
cc_180 N_A_283_48#_c_195_n N_TE_B_c_265_n 0.0180315f $X=2.395 $Y=1.26 $X2=0
+ $Y2=0
cc_181 N_A_283_48#_c_197_n N_TE_B_c_265_n 0.0221236f $X=2.56 $Y=1.17 $X2=0 $Y2=0
cc_182 N_A_283_48#_c_202_n N_TE_B_c_265_n 0.0121482f $X=2.94 $Y=1.985 $X2=0
+ $Y2=0
cc_183 N_A_283_48#_c_199_n N_TE_B_c_265_n 0.00656082f $X=3.005 $Y=0.515 $X2=0
+ $Y2=0
cc_184 N_A_283_48#_c_195_n N_TE_B_c_266_n 8.25111e-19 $X=2.395 $Y=1.26 $X2=0
+ $Y2=0
cc_185 N_A_283_48#_c_197_n N_TE_B_c_266_n 0.00816918f $X=2.56 $Y=1.17 $X2=0
+ $Y2=0
cc_186 N_A_283_48#_c_202_n N_TE_B_c_266_n 0.0068896f $X=2.94 $Y=1.985 $X2=0
+ $Y2=0
cc_187 N_A_283_48#_c_199_n N_TE_B_c_266_n 8.67655e-19 $X=3.005 $Y=0.515 $X2=0
+ $Y2=0
cc_188 N_A_283_48#_c_197_n N_TE_B_M1011_g 0.00109888f $X=2.56 $Y=1.17 $X2=0
+ $Y2=0
cc_189 N_A_283_48#_c_198_n N_TE_B_M1011_g 0.0183842f $X=2.56 $Y=0.49 $X2=0 $Y2=0
cc_190 N_A_283_48#_c_199_n N_TE_B_M1011_g 0.00832294f $X=3.005 $Y=0.515 $X2=0
+ $Y2=0
cc_191 N_A_283_48#_c_196_n N_TE_B_c_268_n 0.0180315f $X=1.925 $Y=1.26 $X2=0
+ $Y2=0
cc_192 N_A_283_48#_c_197_n N_TE_B_c_268_n 8.76501e-19 $X=2.56 $Y=1.17 $X2=0
+ $Y2=0
cc_193 N_A_283_48#_c_197_n TE_B 0.0283543f $X=2.56 $Y=1.17 $X2=0 $Y2=0
cc_194 N_A_283_48#_c_202_n TE_B 0.011045f $X=2.94 $Y=1.985 $X2=0 $Y2=0
cc_195 N_A_283_48#_c_198_n TE_B 0.00125277f $X=2.56 $Y=0.49 $X2=0 $Y2=0
cc_196 N_A_283_48#_c_199_n TE_B 0.015386f $X=3.005 $Y=0.515 $X2=0 $Y2=0
cc_197 N_A_283_48#_c_202_n N_A_c_349_n 0.00105912f $X=2.94 $Y=1.985 $X2=0 $Y2=0
cc_198 N_A_283_48#_c_201_n N_A_33_368#_M1003_d 0.00498962f $X=2.725 $Y=1.945
+ $X2=0 $Y2=0
cc_199 N_A_283_48#_c_193_n Z 2.05626e-19 $X=1.565 $Y=1.26 $X2=0 $Y2=0
cc_200 N_A_283_48#_c_191_n N_A_27_74#_c_511_n 0.00148915f $X=1.49 $Y=1.185 $X2=0
+ $Y2=0
cc_201 N_A_283_48#_c_191_n N_A_27_74#_c_513_n 0.0147594f $X=1.49 $Y=1.185 $X2=0
+ $Y2=0
cc_202 N_A_283_48#_c_192_n N_A_27_74#_c_513_n 0.00230303f $X=1.85 $Y=1.26 $X2=0
+ $Y2=0
cc_203 N_A_283_48#_c_194_n N_A_27_74#_c_513_n 0.012029f $X=1.925 $Y=1.185 $X2=0
+ $Y2=0
cc_204 N_A_283_48#_c_195_n N_A_27_74#_c_513_n 0.00522989f $X=2.395 $Y=1.26 $X2=0
+ $Y2=0
cc_205 N_A_283_48#_c_197_n N_A_27_74#_c_513_n 0.00994473f $X=2.56 $Y=1.17 $X2=0
+ $Y2=0
cc_206 N_A_283_48#_c_198_n N_A_27_74#_c_513_n 0.0012571f $X=2.56 $Y=0.49 $X2=0
+ $Y2=0
cc_207 N_A_283_48#_c_199_n N_A_27_74#_c_513_n 0.00428282f $X=3.005 $Y=0.515
+ $X2=0 $Y2=0
cc_208 N_A_283_48#_c_191_n N_A_27_74#_c_515_n 6.17395e-19 $X=1.49 $Y=1.185 $X2=0
+ $Y2=0
cc_209 N_A_283_48#_c_194_n N_A_27_74#_c_515_n 0.00883931f $X=1.925 $Y=1.185
+ $X2=0 $Y2=0
cc_210 N_A_283_48#_c_198_n N_A_27_74#_c_515_n 0.00224515f $X=2.56 $Y=0.49 $X2=0
+ $Y2=0
cc_211 N_A_283_48#_c_199_n N_A_27_74#_c_515_n 0.0492585f $X=3.005 $Y=0.515 $X2=0
+ $Y2=0
cc_212 N_A_283_48#_c_191_n N_VGND_c_551_n 0.00803879f $X=1.49 $Y=1.185 $X2=0
+ $Y2=0
cc_213 N_A_283_48#_c_194_n N_VGND_c_551_n 0.00291064f $X=1.925 $Y=1.185 $X2=0
+ $Y2=0
cc_214 N_A_283_48#_c_199_n N_VGND_c_551_n 7.47461e-19 $X=3.005 $Y=0.515 $X2=0
+ $Y2=0
cc_215 N_A_283_48#_c_199_n N_VGND_c_552_n 0.0305673f $X=3.005 $Y=0.515 $X2=0
+ $Y2=0
cc_216 N_A_283_48#_c_194_n N_VGND_c_553_n 0.00434272f $X=1.925 $Y=1.185 $X2=0
+ $Y2=0
cc_217 N_A_283_48#_c_198_n N_VGND_c_553_n 0.00804684f $X=2.56 $Y=0.49 $X2=0
+ $Y2=0
cc_218 N_A_283_48#_c_199_n N_VGND_c_553_n 0.0371632f $X=3.005 $Y=0.515 $X2=0
+ $Y2=0
cc_219 N_A_283_48#_c_191_n N_VGND_c_555_n 0.00398535f $X=1.49 $Y=1.185 $X2=0
+ $Y2=0
cc_220 N_A_283_48#_c_191_n N_VGND_c_557_n 0.0078875f $X=1.49 $Y=1.185 $X2=0
+ $Y2=0
cc_221 N_A_283_48#_c_194_n N_VGND_c_557_n 0.00825333f $X=1.925 $Y=1.185 $X2=0
+ $Y2=0
cc_222 N_A_283_48#_c_198_n N_VGND_c_557_n 0.0114187f $X=2.56 $Y=0.49 $X2=0 $Y2=0
cc_223 N_A_283_48#_c_199_n N_VGND_c_557_n 0.0286628f $X=3.005 $Y=0.515 $X2=0
+ $Y2=0
cc_224 N_TE_B_M1011_g N_A_M1001_g 0.0255424f $X=3.22 $Y=0.69 $X2=0 $Y2=0
cc_225 TE_B N_A_M1001_g 9.57049e-19 $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_226 N_TE_B_c_266_n N_A_c_349_n 0.0455244f $X=3.165 $Y=1.765 $X2=0 $Y2=0
cc_227 TE_B N_A_c_349_n 3.46758e-19 $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_228 N_TE_B_c_266_n N_A_c_350_n 0.00518024f $X=3.165 $Y=1.765 $X2=0 $Y2=0
cc_229 TE_B N_A_c_350_n 0.0220909f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_230 N_TE_B_c_270_n N_A_33_368#_c_390_n 0.0112887f $X=1.535 $Y=1.765 $X2=0
+ $Y2=0
cc_231 N_TE_B_c_273_n N_A_33_368#_c_390_n 0.0100505f $X=2.155 $Y=1.765 $X2=0
+ $Y2=0
cc_232 N_TE_B_c_270_n N_A_33_368#_c_382_n 0.0125471f $X=1.535 $Y=1.765 $X2=0
+ $Y2=0
cc_233 N_TE_B_c_273_n N_A_33_368#_c_382_n 0.00168296f $X=2.155 $Y=1.765 $X2=0
+ $Y2=0
cc_234 N_TE_B_c_270_n N_A_33_368#_c_383_n 8.34906e-19 $X=1.535 $Y=1.765 $X2=0
+ $Y2=0
cc_235 N_TE_B_c_273_n N_A_33_368#_c_383_n 0.00567103f $X=2.155 $Y=1.765 $X2=0
+ $Y2=0
cc_236 N_TE_B_c_266_n N_A_33_368#_c_383_n 0.00978103f $X=3.165 $Y=1.765 $X2=0
+ $Y2=0
cc_237 N_TE_B_c_270_n N_Z_c_435_n 7.12084e-19 $X=1.535 $Y=1.765 $X2=0 $Y2=0
cc_238 N_TE_B_c_270_n Z 0.0192873f $X=1.535 $Y=1.765 $X2=0 $Y2=0
cc_239 N_TE_B_c_263_n Z 0.00370154f $X=2.065 $Y=1.65 $X2=0 $Y2=0
cc_240 N_TE_B_c_264_n Z 7.22718e-19 $X=1.625 $Y=1.65 $X2=0 $Y2=0
cc_241 N_TE_B_c_273_n Z 0.00120233f $X=2.155 $Y=1.765 $X2=0 $Y2=0
cc_242 N_TE_B_c_266_n N_VPWR_c_464_n 0.0225268f $X=3.165 $Y=1.765 $X2=0 $Y2=0
cc_243 N_TE_B_c_270_n N_VPWR_c_465_n 0.00317151f $X=1.535 $Y=1.765 $X2=0 $Y2=0
cc_244 N_TE_B_c_273_n N_VPWR_c_466_n 0.00318401f $X=2.155 $Y=1.765 $X2=0 $Y2=0
cc_245 N_TE_B_c_266_n N_VPWR_c_466_n 0.00443511f $X=3.165 $Y=1.765 $X2=0 $Y2=0
cc_246 N_TE_B_c_270_n N_VPWR_c_463_n 0.00396728f $X=1.535 $Y=1.765 $X2=0 $Y2=0
cc_247 N_TE_B_c_273_n N_VPWR_c_463_n 0.00401538f $X=2.155 $Y=1.765 $X2=0 $Y2=0
cc_248 N_TE_B_c_266_n N_VPWR_c_463_n 0.00460931f $X=3.165 $Y=1.765 $X2=0 $Y2=0
cc_249 N_TE_B_c_270_n N_VPWR_c_469_n 0.00196192f $X=1.535 $Y=1.765 $X2=0 $Y2=0
cc_250 N_TE_B_c_273_n N_VPWR_c_469_n 0.00374838f $X=2.155 $Y=1.765 $X2=0 $Y2=0
cc_251 N_TE_B_c_263_n N_A_27_74#_c_513_n 3.02853e-19 $X=2.065 $Y=1.65 $X2=0
+ $Y2=0
cc_252 N_TE_B_c_264_n N_A_27_74#_c_513_n 4.08485e-19 $X=1.625 $Y=1.65 $X2=0
+ $Y2=0
cc_253 N_TE_B_M1011_g N_VGND_c_552_n 0.00678145f $X=3.22 $Y=0.69 $X2=0 $Y2=0
cc_254 N_TE_B_M1011_g N_VGND_c_553_n 0.00432591f $X=3.22 $Y=0.69 $X2=0 $Y2=0
cc_255 N_TE_B_M1011_g N_VGND_c_557_n 0.00822267f $X=3.22 $Y=0.69 $X2=0 $Y2=0
cc_256 N_A_c_349_n N_VPWR_c_464_n 0.00544384f $X=3.815 $Y=1.765 $X2=0 $Y2=0
cc_257 N_A_c_349_n N_VPWR_c_467_n 0.00481995f $X=3.815 $Y=1.765 $X2=0 $Y2=0
cc_258 N_A_c_349_n N_VPWR_c_463_n 0.00508379f $X=3.815 $Y=1.765 $X2=0 $Y2=0
cc_259 N_A_M1001_g N_VGND_c_552_n 0.0072585f $X=3.79 $Y=0.69 $X2=0 $Y2=0
cc_260 N_A_c_349_n N_VGND_c_552_n 9.25785e-19 $X=3.815 $Y=1.765 $X2=0 $Y2=0
cc_261 N_A_c_350_n N_VGND_c_552_n 0.00897894f $X=3.7 $Y=1.515 $X2=0 $Y2=0
cc_262 N_A_M1001_g N_VGND_c_556_n 0.00434272f $X=3.79 $Y=0.69 $X2=0 $Y2=0
cc_263 N_A_M1001_g N_VGND_c_557_n 0.00825084f $X=3.79 $Y=0.69 $X2=0 $Y2=0
cc_264 N_A_33_368#_c_380_n N_Z_M1004_s 0.00250873f $X=1.145 $Y=2.99 $X2=0 $Y2=0
cc_265 N_A_33_368#_c_380_n N_Z_c_435_n 0.018923f $X=1.145 $Y=2.99 $X2=0 $Y2=0
cc_266 N_A_33_368#_M1005_d Z 0.00256509f $X=1.11 $Y=1.84 $X2=0 $Y2=0
cc_267 N_A_33_368#_c_390_n Z 0.00953391f $X=2.215 $Y=2.665 $X2=0 $Y2=0
cc_268 N_A_33_368#_c_382_n Z 0.0212627f $X=1.31 $Y=2.44 $X2=0 $Y2=0
cc_269 N_A_33_368#_c_390_n N_VPWR_M1000_s 0.0139846f $X=2.215 $Y=2.665 $X2=-0.19
+ $Y2=1.66
cc_270 N_A_33_368#_c_380_n N_VPWR_c_465_n 0.0423044f $X=1.145 $Y=2.99 $X2=0
+ $Y2=0
cc_271 N_A_33_368#_c_381_n N_VPWR_c_465_n 0.0236039f $X=0.475 $Y=2.99 $X2=0
+ $Y2=0
cc_272 N_A_33_368#_c_390_n N_VPWR_c_465_n 0.00341854f $X=2.215 $Y=2.665 $X2=0
+ $Y2=0
cc_273 N_A_33_368#_c_382_n N_VPWR_c_465_n 0.0234641f $X=1.31 $Y=2.44 $X2=0 $Y2=0
cc_274 N_A_33_368#_c_390_n N_VPWR_c_466_n 0.00341123f $X=2.215 $Y=2.665 $X2=0
+ $Y2=0
cc_275 N_A_33_368#_c_383_n N_VPWR_c_466_n 0.0140509f $X=2.38 $Y=2.665 $X2=0
+ $Y2=0
cc_276 N_A_33_368#_c_380_n N_VPWR_c_463_n 0.0238902f $X=1.145 $Y=2.99 $X2=0
+ $Y2=0
cc_277 N_A_33_368#_c_381_n N_VPWR_c_463_n 0.012761f $X=0.475 $Y=2.99 $X2=0 $Y2=0
cc_278 N_A_33_368#_c_390_n N_VPWR_c_463_n 0.0125902f $X=2.215 $Y=2.665 $X2=0
+ $Y2=0
cc_279 N_A_33_368#_c_382_n N_VPWR_c_463_n 0.0126878f $X=1.31 $Y=2.44 $X2=0 $Y2=0
cc_280 N_A_33_368#_c_383_n N_VPWR_c_463_n 0.0118378f $X=2.38 $Y=2.665 $X2=0
+ $Y2=0
cc_281 N_A_33_368#_c_390_n N_VPWR_c_469_n 0.0245475f $X=2.215 $Y=2.665 $X2=0
+ $Y2=0
cc_282 N_A_33_368#_c_382_n N_VPWR_c_469_n 0.0105977f $X=1.31 $Y=2.44 $X2=0 $Y2=0
cc_283 N_A_33_368#_c_383_n N_VPWR_c_469_n 0.00406395f $X=2.38 $Y=2.665 $X2=0
+ $Y2=0
cc_284 Z N_VPWR_M1000_s 0.0050653f $X=1.595 $Y=1.95 $X2=-0.19 $Y2=-0.245
cc_285 N_Z_c_428_n N_A_27_74#_c_510_n 0.0201328f $X=0.71 $Y=0.78 $X2=0 $Y2=0
cc_286 N_Z_M1009_d N_A_27_74#_c_511_n 0.00184993f $X=0.57 $Y=0.37 $X2=0 $Y2=0
cc_287 N_Z_c_428_n N_A_27_74#_c_511_n 0.0149881f $X=0.71 $Y=0.78 $X2=0 $Y2=0
cc_288 N_Z_c_424_n N_A_27_74#_c_514_n 0.00732422f $X=0.705 $Y=1.13 $X2=0 $Y2=0
cc_289 N_A_27_74#_c_513_n N_VGND_M1007_d 0.00181776f $X=1.975 $Y=1.045 $X2=-0.19
+ $Y2=-0.245
cc_290 N_A_27_74#_c_511_n N_VGND_c_551_n 0.0114567f $X=1.045 $Y=0.34 $X2=0 $Y2=0
cc_291 N_A_27_74#_c_513_n N_VGND_c_551_n 0.0153175f $X=1.975 $Y=1.045 $X2=0
+ $Y2=0
cc_292 N_A_27_74#_c_515_n N_VGND_c_551_n 0.0158413f $X=2.14 $Y=0.515 $X2=0 $Y2=0
cc_293 N_A_27_74#_c_515_n N_VGND_c_553_n 0.0109942f $X=2.14 $Y=0.515 $X2=0 $Y2=0
cc_294 N_A_27_74#_c_511_n N_VGND_c_555_n 0.0665295f $X=1.045 $Y=0.34 $X2=0 $Y2=0
cc_295 N_A_27_74#_c_512_n N_VGND_c_555_n 0.0179217f $X=0.365 $Y=0.34 $X2=0 $Y2=0
cc_296 N_A_27_74#_c_511_n N_VGND_c_557_n 0.0370229f $X=1.045 $Y=0.34 $X2=0 $Y2=0
cc_297 N_A_27_74#_c_512_n N_VGND_c_557_n 0.00971942f $X=0.365 $Y=0.34 $X2=0
+ $Y2=0
cc_298 N_A_27_74#_c_515_n N_VGND_c_557_n 0.00904371f $X=2.14 $Y=0.515 $X2=0
+ $Y2=0
