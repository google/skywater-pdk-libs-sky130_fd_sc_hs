* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hs__ebufn_2 A TE_B VGND VNB VPB VPWR Z
M1000 a_33_368# TE_B VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=1.0528e+12p pd=8.6e+06u as=1.0815e+12p ps=6.56e+06u
M1001 a_84_48# A VGND VNB nlowvt w=640000u l=150000u
+  ad=1.824e+11p pd=1.85e+06u as=4.797e+11p ps=4.17e+06u
M1002 a_84_48# A VPWR VPB pshort w=1e+06u l=150000u
+  ad=2.95e+11p pd=2.59e+06u as=0p ps=0u
M1003 VPWR TE_B a_33_368# VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_33_368# a_84_48# Z VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=3.92e+11p ps=2.94e+06u
M1005 Z a_84_48# a_33_368# VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VPWR TE_B a_283_48# VPB pshort w=1e+06u l=150000u
+  ad=0p pd=0u as=2.95e+11p ps=2.59e+06u
M1007 VGND a_283_48# a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=7.289e+11p ps=6.41e+06u
M1008 a_27_74# a_283_48# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 Z a_84_48# a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=2.072e+11p pd=2.04e+06u as=0p ps=0u
M1010 a_27_74# a_84_48# Z VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VGND TE_B a_283_48# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=1.824e+11p ps=1.85e+06u
.ends
