* File: sky130_fd_sc_hs__o41a_2.pex.spice
* Created: Tue Sep  1 20:19:16 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HS__O41A_2%A1 3 5 7 8 12
r25 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.43
+ $Y=1.515 $X2=0.43 $Y2=1.515
r26 8 12 5.09219 $w=4.28e-07 $l=1.9e-07 $layer=LI1_cond $X=0.24 $Y=1.565
+ $X2=0.43 $Y2=1.565
r27 5 11 52.2586 $w=2.99e-07 $l=2.85044e-07 $layer=POLY_cond $X=0.505 $Y=1.765
+ $X2=0.43 $Y2=1.515
r28 5 7 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.505 $Y=1.765
+ $X2=0.505 $Y2=2.4
r29 1 11 38.5562 $w=2.99e-07 $l=1.94808e-07 $layer=POLY_cond $X=0.495 $Y=1.35
+ $X2=0.43 $Y2=1.515
r30 1 3 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=0.495 $Y=1.35
+ $X2=0.495 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HS__O41A_2%A2 1 3 6 10 13 14 15
c35 1 0 1.89954e-19 $X=0.925 $Y=1.765
r36 14 15 9.21977 $w=4.78e-07 $l=3.7e-07 $layer=LI1_cond $X=1.075 $Y=2.405
+ $X2=1.075 $Y2=2.775
r37 14 20 6.10498 $w=4.78e-07 $l=2.45e-07 $layer=LI1_cond $X=1.075 $Y=2.405
+ $X2=1.075 $Y2=2.16
r38 13 20 3.11479 $w=4.78e-07 $l=1.25e-07 $layer=LI1_cond $X=1.075 $Y=2.035
+ $X2=1.075 $Y2=2.16
r39 13 27 4.04332 $w=4.78e-07 $l=1.15e-07 $layer=LI1_cond $X=1.075 $Y=2.035
+ $X2=1.075 $Y2=1.92
r40 10 27 14.1436 $w=3.28e-07 $l=4.05e-07 $layer=LI1_cond $X=1 $Y=1.515 $X2=1
+ $Y2=1.92
r41 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1 $Y=1.515
+ $X2=1 $Y2=1.515
r42 4 11 38.5562 $w=2.99e-07 $l=1.94808e-07 $layer=POLY_cond $X=1.065 $Y=1.35
+ $X2=1 $Y2=1.515
r43 4 6 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.065 $Y=1.35
+ $X2=1.065 $Y2=0.74
r44 1 11 52.2586 $w=2.99e-07 $l=2.85044e-07 $layer=POLY_cond $X=0.925 $Y=1.765
+ $X2=1 $Y2=1.515
r45 1 3 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.925 $Y=1.765
+ $X2=0.925 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_HS__O41A_2%A3 3 5 7 8 9 10 11
c35 5 0 1.367e-19 $X=1.495 $Y=1.765
r36 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.57
+ $Y=1.515 $X2=1.57 $Y2=1.515
r37 10 11 18.5393 $w=2.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.68 $Y=2.405
+ $X2=1.68 $Y2=2.775
r38 9 10 18.5393 $w=2.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.68 $Y=2.035
+ $X2=1.68 $Y2=2.405
r39 8 20 2.85155 $w=2.3e-07 $l=1.65e-07 $layer=LI1_cond $X=1.68 $Y=1.515
+ $X2=1.68 $Y2=1.68
r40 8 19 3.84148 $w=3.28e-07 $l=1.1e-07 $layer=LI1_cond $X=1.68 $Y=1.515
+ $X2=1.57 $Y2=1.515
r41 8 9 16.034 $w=2.28e-07 $l=3.2e-07 $layer=LI1_cond $X=1.68 $Y=1.715 $X2=1.68
+ $Y2=2.035
r42 8 20 1.75372 $w=2.28e-07 $l=3.5e-08 $layer=LI1_cond $X=1.68 $Y=1.715
+ $X2=1.68 $Y2=1.68
r43 5 18 52.2586 $w=2.99e-07 $l=2.85044e-07 $layer=POLY_cond $X=1.495 $Y=1.765
+ $X2=1.57 $Y2=1.515
r44 5 7 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.495 $Y=1.765
+ $X2=1.495 $Y2=2.4
r45 1 18 38.5562 $w=2.99e-07 $l=1.98997e-07 $layer=POLY_cond $X=1.495 $Y=1.35
+ $X2=1.57 $Y2=1.515
r46 1 3 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.495 $Y=1.35
+ $X2=1.495 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HS__O41A_2%A4 1 3 6 8 12
r28 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.14
+ $Y=1.515 $X2=2.14 $Y2=1.515
r29 8 12 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=2.14 $Y=1.665
+ $X2=2.14 $Y2=1.515
r30 4 11 38.5562 $w=2.99e-07 $l=2.05122e-07 $layer=POLY_cond $X=2.23 $Y=1.35
+ $X2=2.14 $Y2=1.515
r31 4 6 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.23 $Y=1.35 $X2=2.23
+ $Y2=0.74
r32 1 11 52.2586 $w=2.99e-07 $l=2.85044e-07 $layer=POLY_cond $X=2.065 $Y=1.765
+ $X2=2.14 $Y2=1.515
r33 1 3 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.065 $Y=1.765
+ $X2=2.065 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_HS__O41A_2%B1 1 3 6 8 9
c35 1 0 8.8899e-20 $X=2.635 $Y=1.765
r36 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.71
+ $Y=1.515 $X2=2.71 $Y2=1.515
r37 9 14 10.9884 $w=4.28e-07 $l=4.1e-07 $layer=LI1_cond $X=3.12 $Y=1.565
+ $X2=2.71 $Y2=1.565
r38 8 14 1.87607 $w=4.28e-07 $l=7e-08 $layer=LI1_cond $X=2.64 $Y=1.565 $X2=2.71
+ $Y2=1.565
r39 4 13 38.5562 $w=2.99e-07 $l=1.81659e-07 $layer=POLY_cond $X=2.675 $Y=1.35
+ $X2=2.71 $Y2=1.515
r40 4 6 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.675 $Y=1.35
+ $X2=2.675 $Y2=0.74
r41 1 13 52.2586 $w=2.99e-07 $l=2.85044e-07 $layer=POLY_cond $X=2.635 $Y=1.765
+ $X2=2.71 $Y2=1.515
r42 1 3 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=2.635 $Y=1.765
+ $X2=2.635 $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_HS__O41A_2%A_428_368# 1 2 9 11 13 16 18 20 21 23 25 29
+ 31 32 34 36 44
c78 36 0 8.8899e-20 $X=3.57 $Y=1.465
c79 21 0 1.367e-19 $X=2.29 $Y=2.12
r80 44 45 7.92329 $w=3.65e-07 $l=6e-08 $layer=POLY_cond $X=4.235 $Y=1.532
+ $X2=4.295 $Y2=1.532
r81 43 44 51.5014 $w=3.65e-07 $l=3.9e-07 $layer=POLY_cond $X=3.845 $Y=1.532
+ $X2=4.235 $Y2=1.532
r82 42 43 5.28219 $w=3.65e-07 $l=4e-08 $layer=POLY_cond $X=3.805 $Y=1.532
+ $X2=3.845 $Y2=1.532
r83 37 42 31.0329 $w=3.65e-07 $l=2.35e-07 $layer=POLY_cond $X=3.57 $Y=1.532
+ $X2=3.805 $Y2=1.532
r84 36 40 14.8553 $w=3.3e-07 $l=3.7e-07 $layer=LI1_cond $X=3.57 $Y=1.465
+ $X2=3.57 $Y2=1.095
r85 36 37 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.57
+ $Y=1.465 $X2=3.57 $Y2=1.465
r86 34 36 16.9374 $w=3.28e-07 $l=4.85e-07 $layer=LI1_cond $X=3.57 $Y=1.95
+ $X2=3.57 $Y2=1.465
r87 31 40 2.45823 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.405 $Y=1.095
+ $X2=3.57 $Y2=1.095
r88 31 32 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=3.405 $Y=1.095
+ $X2=3.125 $Y2=1.095
r89 27 32 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.96 $Y=1.01
+ $X2=3.125 $Y2=1.095
r90 27 29 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=2.96 $Y=1.01
+ $X2=2.96 $Y2=0.515
r91 26 39 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.455 $Y=2.035
+ $X2=2.29 $Y2=2.035
r92 25 34 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.405 $Y=2.035
+ $X2=3.57 $Y2=1.95
r93 25 26 61.9786 $w=1.68e-07 $l=9.5e-07 $layer=LI1_cond $X=3.405 $Y=2.035
+ $X2=2.455 $Y2=2.035
r94 21 39 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.29 $Y=2.12 $X2=2.29
+ $Y2=2.035
r95 21 23 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=2.29 $Y=2.12
+ $X2=2.29 $Y2=2.815
r96 18 45 23.6381 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=4.295 $Y=1.765
+ $X2=4.295 $Y2=1.532
r97 18 20 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=4.295 $Y=1.765
+ $X2=4.295 $Y2=2.4
r98 14 44 23.6381 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=4.235 $Y=1.3
+ $X2=4.235 $Y2=1.532
r99 14 16 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=4.235 $Y=1.3
+ $X2=4.235 $Y2=0.74
r100 11 43 23.6381 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=3.845 $Y=1.765
+ $X2=3.845 $Y2=1.532
r101 11 13 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.845 $Y=1.765
+ $X2=3.845 $Y2=2.4
r102 7 42 23.6381 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=3.805 $Y=1.3
+ $X2=3.805 $Y2=1.532
r103 7 9 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=3.805 $Y=1.3
+ $X2=3.805 $Y2=0.74
r104 2 39 300 $w=1.7e-07 $l=3.4187e-07 $layer=licon1_PDIFF $count=2 $X=2.14
+ $Y=1.84 $X2=2.29 $Y2=2.115
r105 2 23 600 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=2.14
+ $Y=1.84 $X2=2.29 $Y2=2.815
r106 1 29 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.75
+ $Y=0.37 $X2=2.89 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__O41A_2%VPWR 1 2 3 10 12 16 18 22 24 32 41 50
r48 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r49 38 39 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r50 36 50 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=4.56 $Y2=3.33
r51 36 46 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=3.6 $Y2=3.33
r52 35 36 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r53 33 35 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=3.78 $Y=3.33 $X2=4.08
+ $Y2=3.33
r54 32 49 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=4.355 $Y=3.33
+ $X2=4.577 $Y2=3.33
r55 32 35 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=4.355 $Y=3.33
+ $X2=4.08 $Y2=3.33
r56 31 46 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.6 $Y2=3.33
r57 30 31 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r58 28 39 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r59 27 30 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=0.72 $Y=3.33
+ $X2=2.64 $Y2=3.33
r60 27 28 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r61 25 38 4.73185 $w=1.7e-07 $l=2.23e-07 $layer=LI1_cond $X=0.445 $Y=3.33
+ $X2=0.222 $Y2=3.33
r62 25 27 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=0.445 $Y=3.33
+ $X2=0.72 $Y2=3.33
r63 24 33 12.2881 $w=1.7e-07 $l=5.43e-07 $layer=LI1_cond $X=3.237 $Y=3.33
+ $X2=3.78 $Y2=3.33
r64 24 46 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r65 24 41 10.7382 $w=1.083e-06 $l=9.55e-07 $layer=LI1_cond $X=3.237 $Y=3.33
+ $X2=3.237 $Y2=2.375
r66 24 30 3.58824 $w=1.68e-07 $l=5.5e-08 $layer=LI1_cond $X=2.695 $Y=3.33
+ $X2=2.64 $Y2=3.33
r67 22 31 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.4 $Y=3.33
+ $X2=2.64 $Y2=3.33
r68 22 28 0.468274 $w=4.9e-07 $l=1.68e-06 $layer=MET1_cond $X=2.4 $Y=3.33
+ $X2=0.72 $Y2=3.33
r69 18 21 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=4.52 $Y=1.985
+ $X2=4.52 $Y2=2.815
r70 16 49 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=4.52 $Y=3.245
+ $X2=4.577 $Y2=3.33
r71 16 21 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=4.52 $Y=3.245
+ $X2=4.52 $Y2=2.815
r72 12 15 24.4458 $w=3.28e-07 $l=7e-07 $layer=LI1_cond $X=0.28 $Y=2.115 $X2=0.28
+ $Y2=2.815
r73 10 38 3.03433 $w=3.3e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.28 $Y=3.245
+ $X2=0.222 $Y2=3.33
r74 10 15 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=0.28 $Y=3.245
+ $X2=0.28 $Y2=2.815
r75 3 21 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=4.37
+ $Y=1.84 $X2=4.52 $Y2=2.815
r76 3 18 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=4.37
+ $Y=1.84 $X2=4.52 $Y2=1.985
r77 2 41 300 $w=1.7e-07 $l=1.14158e-06 $layer=licon1_PDIFF $count=2 $X=2.71
+ $Y=1.84 $X2=3.615 $Y2=2.375
r78 2 41 150 $w=1.7e-07 $l=7.45922e-07 $layer=licon1_PDIFF $count=4 $X=2.71
+ $Y=1.84 $X2=3.215 $Y2=2.375
r79 1 15 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.815
r80 1 12 400 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.115
.ends

.subckt PM_SKY130_FD_SC_HS__O41A_2%X 1 2 9 11 13 17
r23 13 15 44.9047 $w=2.03e-07 $l=8.3e-07 $layer=LI1_cond $X=4.052 $Y=1.985
+ $X2=4.052 $Y2=2.815
r24 11 17 5.91863 $w=2.75e-07 $l=1.27789e-07 $layer=LI1_cond $X=4.052 $Y=1.41
+ $X2=4.025 $Y2=1.295
r25 11 13 31.1086 $w=2.03e-07 $l=5.75e-07 $layer=LI1_cond $X=4.052 $Y=1.41
+ $X2=4.052 $Y2=1.985
r26 7 17 12.5749 $w=3.3e-07 $l=3.32491e-07 $layer=LI1_cond $X=4.02 $Y=0.965
+ $X2=4.025 $Y2=1.295
r27 7 9 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=4.02 $Y=0.965 $X2=4.02
+ $Y2=0.515
r28 2 15 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=3.92
+ $Y=1.84 $X2=4.07 $Y2=2.815
r29 2 13 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=3.92
+ $Y=1.84 $X2=4.07 $Y2=1.985
r30 1 9 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.88
+ $Y=0.37 $X2=4.02 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__O41A_2%A_27_74# 1 2 3 12 14 15 18 20 24 26
c53 26 0 1.89954e-19 $X=1.28 $Y=1.095
r54 22 24 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=2.46 $Y=1.01
+ $X2=2.46 $Y2=0.515
r55 21 26 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.445 $Y=1.095
+ $X2=1.28 $Y2=1.095
r56 20 22 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.295 $Y=1.095
+ $X2=2.46 $Y2=1.01
r57 20 21 55.4545 $w=1.68e-07 $l=8.5e-07 $layer=LI1_cond $X=2.295 $Y=1.095
+ $X2=1.445 $Y2=1.095
r58 16 26 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.28 $Y=1.01 $X2=1.28
+ $Y2=1.095
r59 16 18 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=1.28 $Y=1.01
+ $X2=1.28 $Y2=0.515
r60 14 26 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.115 $Y=1.095
+ $X2=1.28 $Y2=1.095
r61 14 15 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.115 $Y=1.095
+ $X2=0.445 $Y2=1.095
r62 10 15 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.28 $Y=1.01
+ $X2=0.445 $Y2=1.095
r63 10 12 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=0.28 $Y=1.01
+ $X2=0.28 $Y2=0.515
r64 3 24 91 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_NDIFF $count=2 $X=2.305
+ $Y=0.37 $X2=2.46 $Y2=0.515
r65 2 18 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.14
+ $Y=0.37 $X2=1.28 $Y2=0.515
r66 1 12 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__O41A_2%VGND 1 2 3 4 15 17 21 25 27 29 31 33 38 46 52
+ 55 58 62
r61 61 62 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r62 58 59 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r63 55 56 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r64 53 56 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r65 52 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r66 50 62 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=4.56
+ $Y2=0
r67 50 59 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=3.6
+ $Y2=0
r68 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r69 47 58 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.685 $Y=0 $X2=3.52
+ $Y2=0
r70 47 49 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=3.685 $Y=0 $X2=4.08
+ $Y2=0
r71 46 61 4.01281 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=4.355 $Y=0 $X2=4.577
+ $Y2=0
r72 46 49 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=4.355 $Y=0 $X2=4.08
+ $Y2=0
r73 45 59 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=3.6
+ $Y2=0
r74 44 45 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r75 42 56 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.68
+ $Y2=0
r76 41 44 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=2.16 $Y=0 $X2=3.12
+ $Y2=0
r77 41 42 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r78 39 55 11.4275 $w=1.7e-07 $l=2.55e-07 $layer=LI1_cond $X=2.125 $Y=0 $X2=1.87
+ $Y2=0
r79 39 41 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=2.125 $Y=0 $X2=2.16
+ $Y2=0
r80 38 58 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.355 $Y=0 $X2=3.52
+ $Y2=0
r81 38 44 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=3.355 $Y=0 $X2=3.12
+ $Y2=0
r82 36 53 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r83 35 36 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r84 33 52 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.615 $Y=0 $X2=0.78
+ $Y2=0
r85 33 35 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=0.615 $Y=0 $X2=0.24
+ $Y2=0
r86 31 45 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=2.4 $Y=0 $X2=3.12
+ $Y2=0
r87 31 42 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.4 $Y=0 $X2=2.16
+ $Y2=0
r88 27 61 3.19941 $w=2.6e-07 $l=1.27609e-07 $layer=LI1_cond $X=4.485 $Y=0.085
+ $X2=4.577 $Y2=0
r89 27 29 18.1731 $w=2.58e-07 $l=4.1e-07 $layer=LI1_cond $X=4.485 $Y=0.085
+ $X2=4.485 $Y2=0.495
r90 23 58 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.52 $Y=0.085
+ $X2=3.52 $Y2=0
r91 23 25 19.9058 $w=3.28e-07 $l=5.7e-07 $layer=LI1_cond $X=3.52 $Y=0.085
+ $X2=3.52 $Y2=0.655
r92 19 55 2.12513 $w=5.1e-07 $l=8.5e-08 $layer=LI1_cond $X=1.87 $Y=0.085
+ $X2=1.87 $Y2=0
r93 19 21 12.4298 $w=5.08e-07 $l=5.3e-07 $layer=LI1_cond $X=1.87 $Y=0.085
+ $X2=1.87 $Y2=0.615
r94 18 52 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.945 $Y=0 $X2=0.78
+ $Y2=0
r95 17 55 11.4275 $w=1.7e-07 $l=2.55e-07 $layer=LI1_cond $X=1.615 $Y=0 $X2=1.87
+ $Y2=0
r96 17 18 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.615 $Y=0 $X2=0.945
+ $Y2=0
r97 13 52 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.78 $Y=0.085
+ $X2=0.78 $Y2=0
r98 13 15 17.8105 $w=3.28e-07 $l=5.1e-07 $layer=LI1_cond $X=0.78 $Y=0.085
+ $X2=0.78 $Y2=0.595
r99 4 29 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=4.31
+ $Y=0.37 $X2=4.45 $Y2=0.495
r100 3 25 182 $w=1.7e-07 $l=3.77492e-07 $layer=licon1_NDIFF $count=1 $X=3.375
+ $Y=0.37 $X2=3.59 $Y2=0.655
r101 2 21 182 $w=1.7e-07 $l=4.04351e-07 $layer=licon1_NDIFF $count=1 $X=1.57
+ $Y=0.37 $X2=1.87 $Y2=0.615
r102 1 15 182 $w=1.7e-07 $l=3.1285e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.37 $X2=0.78 $Y2=0.595
.ends

