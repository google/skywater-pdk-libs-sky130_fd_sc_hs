* NGSPICE file created from sky130_fd_sc_hs__buf_2.ext - technology: sky130A

.subckt sky130_fd_sc_hs__buf_2 A VGND VNB VPB VPWR X
M1000 VGND a_21_260# X VNB nlowvt w=740000u l=150000u
+  ad=5.216e+11p pd=4.39e+06u as=2.072e+11p ps=2.04e+06u
M1001 a_21_260# A VGND VNB nlowvt w=640000u l=150000u
+  ad=1.824e+11p pd=1.85e+06u as=0p ps=0u
M1002 X a_21_260# VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=3.36e+11p pd=2.84e+06u as=1.1764e+12p ps=6.6e+06u
M1003 VPWR a_21_260# X VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 X a_21_260# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_21_260# A VPWR VPB pshort w=1e+06u l=150000u
+  ad=3.2e+11p pd=2.64e+06u as=0p ps=0u
.ends

