* File: sky130_fd_sc_hs__fahcin_1.pex.spice
* Created: Tue Sep  1 20:05:57 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HS__FAHCIN_1%A 3 5 7 8 12
r30 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.71
+ $Y=1.515 $X2=0.71 $Y2=1.515
r31 8 12 5.96091 $w=2.88e-07 $l=1.5e-07 $layer=LI1_cond $X=0.69 $Y=1.665
+ $X2=0.69 $Y2=1.515
r32 5 11 49.8683 $w=3.94e-07 $l=3.10242e-07 $layer=POLY_cond $X=0.515 $Y=1.765
+ $X2=0.65 $Y2=1.515
r33 5 7 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.515 $Y=1.765
+ $X2=0.515 $Y2=2.4
r34 1 11 39.4698 $w=3.94e-07 $l=2.2798e-07 $layer=POLY_cond $X=0.5 $Y=1.35
+ $X2=0.65 $Y2=1.515
r35 1 3 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=0.5 $Y=1.35 $X2=0.5
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HS__FAHCIN_1%A_28_74# 1 2 3 4 13 15 18 22 26 30 32 33 35
+ 36 37 38 39 42 46 48
c105 33 0 1.71384e-19 $X=1.09 $Y=2.905
r106 51 52 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.28
+ $Y=1.465 $X2=1.28 $Y2=1.465
r107 49 51 12.2997 $w=3.67e-07 $l=3.7e-07 $layer=LI1_cond $X=1.225 $Y=1.095
+ $X2=1.225 $Y2=1.465
r108 44 46 21.8964 $w=2.48e-07 $l=4.75e-07 $layer=LI1_cond $X=3.81 $Y=2.905
+ $X2=3.81 $Y2=2.43
r109 40 42 5.76222 $w=2.48e-07 $l=1.25e-07 $layer=LI1_cond $X=2.71 $Y=0.425
+ $X2=2.71 $Y2=0.55
r110 38 40 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=2.585 $Y=0.34
+ $X2=2.71 $Y2=0.425
r111 38 39 84.4866 $w=1.68e-07 $l=1.295e-06 $layer=LI1_cond $X=2.585 $Y=0.34
+ $X2=1.29 $Y2=0.34
r112 36 44 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=3.685 $Y=2.99
+ $X2=3.81 $Y2=2.905
r113 36 37 163.754 $w=1.68e-07 $l=2.51e-06 $layer=LI1_cond $X=3.685 $Y=2.99
+ $X2=1.175 $Y2=2.99
r114 35 49 6.3706 $w=3.67e-07 $l=9.44722e-08 $layer=LI1_cond $X=1.205 $Y=1.01
+ $X2=1.225 $Y2=1.095
r115 34 39 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.205 $Y=0.425
+ $X2=1.29 $Y2=0.34
r116 34 35 38.1658 $w=1.68e-07 $l=5.85e-07 $layer=LI1_cond $X=1.205 $Y=0.425
+ $X2=1.205 $Y2=1.01
r117 33 37 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.09 $Y=2.905
+ $X2=1.175 $Y2=2.99
r118 32 51 9.03 $w=3.67e-07 $l=2.22486e-07 $layer=LI1_cond $X=1.09 $Y=1.63
+ $X2=1.225 $Y2=1.465
r119 32 33 83.1818 $w=1.68e-07 $l=1.275e-06 $layer=LI1_cond $X=1.09 $Y=1.63
+ $X2=1.09 $Y2=2.905
r120 31 48 3.35233 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.45 $Y=1.095
+ $X2=0.285 $Y2=1.095
r121 30 49 5.25812 $w=1.7e-07 $l=2.2e-07 $layer=LI1_cond $X=1.005 $Y=1.095
+ $X2=1.225 $Y2=1.095
r122 30 31 36.2086 $w=1.68e-07 $l=5.55e-07 $layer=LI1_cond $X=1.005 $Y=1.095
+ $X2=0.45 $Y2=1.095
r123 26 28 37.5109 $w=2.53e-07 $l=8.3e-07 $layer=LI1_cond $X=0.247 $Y=1.985
+ $X2=0.247 $Y2=2.815
r124 24 48 3.22182 $w=2.92e-07 $l=1.0225e-07 $layer=LI1_cond $X=0.247 $Y=1.18
+ $X2=0.285 $Y2=1.095
r125 24 26 36.381 $w=2.53e-07 $l=8.05e-07 $layer=LI1_cond $X=0.247 $Y=1.18
+ $X2=0.247 $Y2=1.985
r126 20 48 3.22182 $w=2.92e-07 $l=8.5e-08 $layer=LI1_cond $X=0.285 $Y=1.01
+ $X2=0.285 $Y2=1.095
r127 20 22 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=0.285 $Y=1.01
+ $X2=0.285 $Y2=0.515
r128 16 52 38.5347 $w=3.14e-07 $l=2.13014e-07 $layer=POLY_cond $X=1.41 $Y=1.3
+ $X2=1.3 $Y2=1.465
r129 16 18 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=1.41 $Y=1.3
+ $X2=1.41 $Y2=0.79
r130 13 52 59.2576 $w=3.14e-07 $l=3.44238e-07 $layer=POLY_cond $X=1.205 $Y=1.765
+ $X2=1.3 $Y2=1.465
r131 13 15 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=1.205 $Y=1.765
+ $X2=1.205 $Y2=2.34
r132 4 46 600 $w=1.7e-07 $l=6.27077e-07 $layer=licon1_PDIFF $count=1 $X=3.65
+ $Y=1.895 $X2=3.85 $Y2=2.43
r133 3 28 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=0.145
+ $Y=1.84 $X2=0.29 $Y2=2.815
r134 3 26 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.145
+ $Y=1.84 $X2=0.29 $Y2=1.985
r135 2 42 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=2.61 $Y=0.37
+ $X2=2.75 $Y2=0.55
r136 1 22 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.14
+ $Y=0.37 $X2=0.285 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__FAHCIN_1%A_492_48# 1 2 9 12 13 15 16 18 20 23 25 27
+ 30 32 34 35 36 40 41 43 44 48 50 53 59 61
c171 30 0 1.21008e-19 $X=6.09 $Y=0.725
c172 13 0 1.89903e-19 $X=2.55 $Y=2.015
c173 9 0 1.01566e-19 $X=2.535 $Y=0.69
r174 59 62 8.47192 $w=3.38e-07 $l=1.65e-07 $layer=LI1_cond $X=5.8 $Y=1.42
+ $X2=5.8 $Y2=1.585
r175 59 61 8.47192 $w=3.38e-07 $l=1.65e-07 $layer=LI1_cond $X=5.8 $Y=1.42
+ $X2=5.8 $Y2=1.255
r176 59 60 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.84
+ $Y=1.42 $X2=5.84 $Y2=1.42
r177 53 56 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=5.12 $Y=1.905
+ $X2=5.12 $Y2=2.055
r178 51 63 2.6208 $w=4.23e-07 $l=2.3e-08 $layer=POLY_cond $X=3.737 $Y=1.545
+ $X2=3.737 $Y2=1.522
r179 50 52 18.2271 $w=2.51e-07 $l=3.75e-07 $layer=LI1_cond $X=3.825 $Y=1.545
+ $X2=4.2 $Y2=1.545
r180 50 51 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.825
+ $Y=1.545 $X2=3.825 $Y2=1.545
r181 48 62 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=5.715 $Y=1.82
+ $X2=5.715 $Y2=1.585
r182 45 61 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=5.715 $Y=1.01
+ $X2=5.715 $Y2=1.255
r183 43 45 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.63 $Y=0.925
+ $X2=5.715 $Y2=1.01
r184 43 44 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=5.63 $Y=0.925
+ $X2=5.295 $Y2=0.925
r185 42 53 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.285 $Y=1.905
+ $X2=5.12 $Y2=1.905
r186 41 48 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.63 $Y=1.905
+ $X2=5.715 $Y2=1.82
r187 41 42 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=5.63 $Y=1.905
+ $X2=5.285 $Y2=1.905
r188 38 44 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=5.13 $Y=0.84
+ $X2=5.295 $Y2=0.925
r189 38 40 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=5.13 $Y=0.84
+ $X2=5.13 $Y2=0.585
r190 37 40 5.5876 $w=3.28e-07 $l=1.6e-07 $layer=LI1_cond $X=5.13 $Y=0.425
+ $X2=5.13 $Y2=0.585
r191 35 37 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.965 $Y=0.34
+ $X2=5.13 $Y2=0.425
r192 35 36 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=4.965 $Y=0.34
+ $X2=4.285 $Y2=0.34
r193 34 52 3.01842 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.2 $Y=1.38 $X2=4.2
+ $Y2=1.545
r194 33 36 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.2 $Y=0.425
+ $X2=4.285 $Y2=0.34
r195 33 34 62.3048 $w=1.68e-07 $l=9.55e-07 $layer=LI1_cond $X=4.2 $Y=0.425
+ $X2=4.2 $Y2=1.38
r196 28 60 39.2181 $w=3.8e-07 $l=2.38642e-07 $layer=POLY_cond $X=6.09 $Y=1.255
+ $X2=5.92 $Y2=1.42
r197 28 30 271.766 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=6.09 $Y=1.255
+ $X2=6.09 $Y2=0.725
r198 25 60 62.0497 $w=3.8e-07 $l=3.49964e-07 $layer=POLY_cond $X=5.91 $Y=1.765
+ $X2=5.92 $Y2=1.42
r199 25 27 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=5.91 $Y=1.765
+ $X2=5.91 $Y2=2.34
r200 21 63 37.4425 $w=4.23e-07 $l=1.82285e-07 $layer=POLY_cond $X=3.645 $Y=1.38
+ $X2=3.737 $Y2=1.522
r201 21 23 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=3.645 $Y=1.38
+ $X2=3.645 $Y2=0.915
r202 18 51 52.5976 $w=4.23e-07 $l=3.46663e-07 $layer=POLY_cond $X=3.575 $Y=1.82
+ $X2=3.737 $Y2=1.545
r203 18 20 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=3.575 $Y=1.82
+ $X2=3.575 $Y2=2.315
r204 17 32 2.09011 $w=2.85e-07 $l=9e-08 $layer=POLY_cond $X=2.64 $Y=1.522
+ $X2=2.55 $Y2=1.522
r205 16 63 12.1026 $w=2.85e-07 $l=2.52e-07 $layer=POLY_cond $X=3.485 $Y=1.522
+ $X2=3.737 $Y2=1.522
r206 16 17 177.856 $w=2.85e-07 $l=8.45e-07 $layer=POLY_cond $X=3.485 $Y=1.522
+ $X2=2.64 $Y2=1.522
r207 13 15 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=2.55 $Y=2.015
+ $X2=2.55 $Y2=2.51
r208 12 13 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=2.55 $Y=1.925
+ $X2=2.55 $Y2=2.015
r209 11 32 31.2989 $w=1.65e-07 $l=1.43e-07 $layer=POLY_cond $X=2.55 $Y=1.665
+ $X2=2.55 $Y2=1.522
r210 11 12 101.065 $w=1.8e-07 $l=2.6e-07 $layer=POLY_cond $X=2.55 $Y=1.665
+ $X2=2.55 $Y2=1.925
r211 7 32 31.2989 $w=1.65e-07 $l=1.49312e-07 $layer=POLY_cond $X=2.535 $Y=1.38
+ $X2=2.55 $Y2=1.522
r212 7 9 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=2.535 $Y=1.38
+ $X2=2.535 $Y2=0.69
r213 2 56 600 $w=1.7e-07 $l=2.78209e-07 $layer=licon1_PDIFF $count=1 $X=4.975
+ $Y=1.84 $X2=5.12 $Y2=2.055
r214 1 40 91 $w=1.7e-07 $l=2.41868e-07 $layer=licon1_NDIFF $count=2 $X=4.985
+ $Y=0.405 $X2=5.13 $Y2=0.585
.ends

.subckt PM_SKY130_FD_SC_HS__FAHCIN_1%B 1 3 4 6 7 8 9 10 11 12 13 15 18 20 22 25
+ 27 28 30 33 34 35 37 39 40 41
c142 27 0 1.27399e-19 $X=4.835 $Y=1.255
c143 18 0 3.79173e-20 $X=4.305 $Y=0.915
c144 13 0 2.07266e-20 $X=4.29 $Y=2.81
c145 7 0 9.05624e-20 $X=4.23 $Y=0.18
c146 4 0 9.51233e-20 $X=3.04 $Y=3.005
r147 44 45 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.04
+ $Y=1.42 $X2=5.04 $Y2=1.42
r148 41 45 4.36531 $w=3.28e-07 $l=1.25e-07 $layer=LI1_cond $X=5.04 $Y=1.295
+ $X2=5.04 $Y2=1.42
r149 39 44 37.5952 $w=3.3e-07 $l=2.15e-07 $layer=POLY_cond $X=5.255 $Y=1.42
+ $X2=5.04 $Y2=1.42
r150 39 40 66.2869 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=5.345 $Y=1.42
+ $X2=5.345 $Y2=1.255
r151 36 44 22.732 $w=3.3e-07 $l=1.3e-07 $layer=POLY_cond $X=4.91 $Y=1.42
+ $X2=5.04 $Y2=1.42
r152 36 37 5.03009 $w=3.3e-07 $l=1.67332e-07 $layer=POLY_cond $X=4.91 $Y=1.42
+ $X2=4.75 $Y2=1.435
r153 33 40 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=5.36 $Y=0.775
+ $X2=5.36 $Y2=1.255
r154 28 39 136.255 $w=1.8e-07 $l=3.45e-07 $layer=POLY_cond $X=5.345 $Y=1.765
+ $X2=5.345 $Y2=1.42
r155 28 30 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=5.345 $Y=1.765
+ $X2=5.345 $Y2=2.4
r156 27 37 37.0704 $w=1.5e-07 $l=2.18403e-07 $layer=POLY_cond $X=4.835 $Y=1.255
+ $X2=4.75 $Y2=1.435
r157 26 27 512.766 $w=1.5e-07 $l=1e-06 $layer=POLY_cond $X=4.835 $Y=0.255
+ $X2=4.835 $Y2=1.255
r158 24 37 37.0704 $w=1.5e-07 $l=1.83712e-07 $layer=POLY_cond $X=4.825 $Y=1.585
+ $X2=4.75 $Y2=1.435
r159 24 25 764.021 $w=1.5e-07 $l=1.49e-06 $layer=POLY_cond $X=4.825 $Y=1.585
+ $X2=4.825 $Y2=3.075
r160 23 34 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=4.38 $Y=3.15 $X2=4.29
+ $Y2=3.15
r161 22 25 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.75 $Y=3.15
+ $X2=4.825 $Y2=3.075
r162 22 23 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=4.75 $Y=3.15
+ $X2=4.38 $Y2=3.15
r163 21 35 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.38 $Y=0.18
+ $X2=4.305 $Y2=0.18
r164 20 26 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.76 $Y=0.18
+ $X2=4.835 $Y2=0.255
r165 20 21 194.851 $w=1.5e-07 $l=3.8e-07 $layer=POLY_cond $X=4.76 $Y=0.18
+ $X2=4.38 $Y2=0.18
r166 16 35 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.305 $Y=0.255
+ $X2=4.305 $Y2=0.18
r167 16 18 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.305 $Y=0.255
+ $X2=4.305 $Y2=0.915
r168 13 15 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=4.29 $Y=2.81
+ $X2=4.29 $Y2=2.315
r169 12 34 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=4.29 $Y=3.075
+ $X2=4.29 $Y2=3.15
r170 11 13 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=4.29 $Y=2.9 $X2=4.29
+ $Y2=2.81
r171 11 12 68.0242 $w=1.8e-07 $l=1.75e-07 $layer=POLY_cond $X=4.29 $Y=2.9
+ $X2=4.29 $Y2=3.075
r172 9 34 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=4.2 $Y=3.15 $X2=4.29
+ $Y2=3.15
r173 9 10 548.66 $w=1.5e-07 $l=1.07e-06 $layer=POLY_cond $X=4.2 $Y=3.15 $X2=3.13
+ $Y2=3.15
r174 7 35 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.23 $Y=0.18
+ $X2=4.305 $Y2=0.18
r175 7 8 610.191 $w=1.5e-07 $l=1.19e-06 $layer=POLY_cond $X=4.23 $Y=0.18
+ $X2=3.04 $Y2=0.18
r176 4 10 26.9307 $w=1.5e-07 $l=1.84594e-07 $layer=POLY_cond $X=3.04 $Y=3.005
+ $X2=3.13 $Y2=3.15
r177 4 6 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=3.04 $Y=3.005
+ $X2=3.04 $Y2=2.51
r178 1 8 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.965 $Y=0.255
+ $X2=3.04 $Y2=0.18
r179 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.965 $Y=0.255
+ $X2=2.965 $Y2=0.69
.ends

.subckt PM_SKY130_FD_SC_HS__FAHCIN_1%A_608_74# 1 2 7 9 10 12 16 17 18 19 21 22
+ 29 33 35 38 39 40 42 43 44 46 48 49 50 52 53 56 57 58 60 61 63 64 67 68 70 75
+ 79 85
c265 85 0 4.231e-20 $X=8.085 $Y=1.32
c266 70 0 1.05034e-19 $X=6.605 $Y=1.675
c267 67 0 2.07266e-20 $X=3.35 $Y=2.04
c268 63 0 2.11268e-20 $X=10.41 $Y=0.405
c269 35 0 3.79173e-20 $X=4.105 $Y=1.965
r270 76 85 30.6007 $w=3.3e-07 $l=1.75e-07 $layer=POLY_cond $X=7.91 $Y=1.32
+ $X2=8.085 $Y2=1.32
r271 75 78 8.51388 $w=2.88e-07 $l=1.65e-07 $layer=LI1_cond $X=7.89 $Y=1.32
+ $X2=7.89 $Y2=1.485
r272 75 76 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.91
+ $Y=1.32 $X2=7.91 $Y2=1.32
r273 70 73 8.79328 $w=2.48e-07 $l=1.65e-07 $layer=LI1_cond $X=6.605 $Y=1.675
+ $X2=6.605 $Y2=1.84
r274 70 71 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.605
+ $Y=1.675 $X2=6.605 $Y2=1.675
r275 63 64 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=10.41
+ $Y=0.405 $X2=10.41 $Y2=0.405
r276 61 63 37.5001 $w=3.13e-07 $l=1.025e-06 $layer=LI1_cond $X=9.385 $Y=0.412
+ $X2=10.41 $Y2=0.412
r277 59 61 7.64049 $w=3.15e-07 $l=1.95944e-07 $layer=LI1_cond $X=9.3 $Y=0.57
+ $X2=9.385 $Y2=0.412
r278 59 60 70.7861 $w=1.68e-07 $l=1.085e-06 $layer=LI1_cond $X=9.3 $Y=0.57
+ $X2=9.3 $Y2=1.655
r279 57 60 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.215 $Y=1.74
+ $X2=9.3 $Y2=1.655
r280 57 58 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=9.215 $Y=1.74
+ $X2=8.715 $Y2=1.74
r281 55 58 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.63 $Y=1.825
+ $X2=8.715 $Y2=1.74
r282 55 56 70.4599 $w=1.68e-07 $l=1.08e-06 $layer=LI1_cond $X=8.63 $Y=1.825
+ $X2=8.63 $Y2=2.905
r283 54 79 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.955 $Y=2.99
+ $X2=7.87 $Y2=2.99
r284 53 56 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.545 $Y=2.99
+ $X2=8.63 $Y2=2.905
r285 53 54 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=8.545 $Y=2.99
+ $X2=7.955 $Y2=2.99
r286 52 79 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.87 $Y=2.905
+ $X2=7.87 $Y2=2.99
r287 52 78 92.6417 $w=1.68e-07 $l=1.42e-06 $layer=LI1_cond $X=7.87 $Y=2.905
+ $X2=7.87 $Y2=1.485
r288 49 79 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.785 $Y=2.99
+ $X2=7.87 $Y2=2.99
r289 49 50 74.0481 $w=1.68e-07 $l=1.135e-06 $layer=LI1_cond $X=7.785 $Y=2.99
+ $X2=6.65 $Y2=2.99
r290 48 68 2.84813 $w=3.35e-07 $l=2.03101e-07 $layer=LI1_cond $X=6.565 $Y=2.39
+ $X2=6.4 $Y2=2.475
r291 48 73 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=6.565 $Y=2.39
+ $X2=6.565 $Y2=1.84
r292 46 50 9.23067 $w=1.7e-07 $l=2.89396e-07 $layer=LI1_cond $X=6.4 $Y=2.905
+ $X2=6.65 $Y2=2.99
r293 45 68 2.84813 $w=3.35e-07 $l=8.5e-08 $layer=LI1_cond $X=6.4 $Y=2.56 $X2=6.4
+ $Y2=2.475
r294 45 46 8.25294 $w=4.98e-07 $l=3.45e-07 $layer=LI1_cond $X=6.4 $Y=2.56
+ $X2=6.4 $Y2=2.905
r295 43 68 3.86674 $w=1.7e-07 $l=2.5e-07 $layer=LI1_cond $X=6.15 $Y=2.475
+ $X2=6.4 $Y2=2.475
r296 43 44 72.0909 $w=1.68e-07 $l=1.105e-06 $layer=LI1_cond $X=6.15 $Y=2.475
+ $X2=5.045 $Y2=2.475
r297 41 44 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.96 $Y=2.56
+ $X2=5.045 $Y2=2.475
r298 41 42 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=4.96 $Y=2.56
+ $X2=4.96 $Y2=2.905
r299 39 42 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.875 $Y=2.99
+ $X2=4.96 $Y2=2.905
r300 39 40 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=4.875 $Y=2.99
+ $X2=4.275 $Y2=2.99
r301 38 40 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.19 $Y=2.905
+ $X2=4.275 $Y2=2.99
r302 37 38 55.7807 $w=1.68e-07 $l=8.55e-07 $layer=LI1_cond $X=4.19 $Y=2.05
+ $X2=4.19 $Y2=2.905
r303 36 67 2.76166 $w=1.7e-07 $l=1.66493e-07 $layer=LI1_cond $X=3.515 $Y=1.965
+ $X2=3.35 $Y2=1.962
r304 35 37 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.105 $Y=1.965
+ $X2=4.19 $Y2=2.05
r305 35 36 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=4.105 $Y=1.965
+ $X2=3.515 $Y2=1.965
r306 31 67 3.70735 $w=2.5e-07 $l=1.20536e-07 $layer=LI1_cond $X=3.43 $Y=1.875
+ $X2=3.35 $Y2=1.962
r307 31 33 72.7433 $w=1.68e-07 $l=1.115e-06 $layer=LI1_cond $X=3.43 $Y=1.875
+ $X2=3.43 $Y2=0.76
r308 27 67 3.70735 $w=2.5e-07 $l=8.8e-08 $layer=LI1_cond $X=3.35 $Y=2.05
+ $X2=3.35 $Y2=1.962
r309 27 29 18.1597 $w=3.28e-07 $l=5.2e-07 $layer=LI1_cond $X=3.35 $Y=2.05
+ $X2=3.35 $Y2=2.57
r310 22 64 68.1959 $w=3.3e-07 $l=3.9e-07 $layer=POLY_cond $X=10.02 $Y=0.405
+ $X2=10.41 $Y2=0.405
r311 19 21 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=10.205 $Y=1.845
+ $X2=10.205 $Y2=2.34
r312 18 19 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=10.205 $Y=1.755
+ $X2=10.205 $Y2=1.845
r313 17 23 133.319 $w=1.5e-07 $l=2.6e-07 $layer=POLY_cond $X=10.205 $Y=1.47
+ $X2=9.945 $Y2=1.47
r314 17 18 81.629 $w=1.8e-07 $l=2.1e-07 $layer=POLY_cond $X=10.205 $Y=1.545
+ $X2=10.205 $Y2=1.755
r315 14 23 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=9.945 $Y=1.395
+ $X2=9.945 $Y2=1.47
r316 14 16 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=9.945 $Y=1.395
+ $X2=9.945 $Y2=1
r317 13 22 32.1775 $w=3.3e-07 $l=1.98997e-07 $layer=POLY_cond $X=9.945 $Y=0.57
+ $X2=10.02 $Y2=0.405
r318 13 16 220.489 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=9.945 $Y=0.57
+ $X2=9.945 $Y2=1
r319 10 85 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.085 $Y=1.155
+ $X2=8.085 $Y2=1.32
r320 10 12 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=8.085 $Y=1.155
+ $X2=8.085 $Y2=0.725
r321 7 71 51.1109 $w=3.27e-07 $l=2.92404e-07 $layer=POLY_cond $X=6.495 $Y=1.925
+ $X2=6.587 $Y2=1.675
r322 7 9 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=6.495 $Y=1.925
+ $X2=6.495 $Y2=2.42
r323 2 67 600 $w=1.7e-07 $l=2.58795e-07 $layer=licon1_PDIFF $count=1 $X=3.115
+ $Y=2.09 $X2=3.35 $Y2=2.04
r324 2 29 600 $w=1.7e-07 $l=5.85833e-07 $layer=licon1_PDIFF $count=1 $X=3.115
+ $Y=2.09 $X2=3.35 $Y2=2.57
r325 1 33 91 $w=1.7e-07 $l=5.51543e-07 $layer=licon1_NDIFF $count=2 $X=3.04
+ $Y=0.37 $X2=3.43 $Y2=0.76
.ends

.subckt PM_SKY130_FD_SC_HS__FAHCIN_1%A_430_418# 1 2 3 4 13 15 16 17 18 19 20 22
+ 23 25 26 28 33 37 39 41 42 43 44 45 46 49 53 58 62 63 66
c213 49 0 9.51233e-20 $X=2.16 $Y=2.035
c214 26 0 2.11268e-20 $X=10.89 $Y=1.43
c215 16 0 1.05034e-19 $X=7.205 $Y=1.195
r216 65 66 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.85
+ $Y=1.595 $X2=10.85 $Y2=1.595
r217 62 63 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=7.37
+ $Y=1.335 $X2=7.37 $Y2=1.335
r218 59 66 15.3659 $w=3.28e-07 $l=4.4e-07 $layer=LI1_cond $X=10.85 $Y=2.035
+ $X2=10.85 $Y2=1.595
r219 58 59 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.8 $Y=2.035
+ $X2=10.8 $Y2=2.035
r220 56 63 25.6098 $w=3.13e-07 $l=7e-07 $layer=LI1_cond $X=7.397 $Y=2.035
+ $X2=7.397 $Y2=1.335
r221 55 56 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=2.035
+ $X2=7.44 $Y2=2.035
r222 52 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=2.035
+ $X2=4.56 $Y2=2.035
r223 49 80 7.20241 $w=4.15e-07 $l=2.45e-07 $layer=LI1_cond $X=2.265 $Y=2.035
+ $X2=2.265 $Y2=2.28
r224 48 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=2.035
+ $X2=2.16 $Y2=2.035
r225 46 55 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=7.585 $Y=2.035
+ $X2=7.44 $Y2=2.035
r226 45 58 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=10.655 $Y=2.035
+ $X2=10.8 $Y2=2.035
r227 45 46 3.7995 $w=1.4e-07 $l=3.07e-06 $layer=MET1_cond $X=10.655 $Y=2.035
+ $X2=7.585 $Y2=2.035
r228 44 52 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.705 $Y=2.035
+ $X2=4.56 $Y2=2.035
r229 43 55 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=7.295 $Y=2.035
+ $X2=7.44 $Y2=2.035
r230 43 44 3.20544 $w=1.4e-07 $l=2.59e-06 $layer=MET1_cond $X=7.295 $Y=2.035
+ $X2=4.705 $Y2=2.035
r231 42 48 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.305 $Y=2.035
+ $X2=2.16 $Y2=2.035
r232 41 52 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.415 $Y=2.035
+ $X2=4.56 $Y2=2.035
r233 41 42 2.61138 $w=1.4e-07 $l=2.11e-06 $layer=MET1_cond $X=4.415 $Y=2.035
+ $X2=2.305 $Y2=2.035
r234 39 53 1.32974 $w=2.58e-07 $l=3e-08 $layer=LI1_cond $X=4.575 $Y=2.005
+ $X2=4.575 $Y2=2.035
r235 39 40 5.76222 $w=2.58e-07 $l=1.3e-07 $layer=LI1_cond $X=4.575 $Y=2.005
+ $X2=4.575 $Y2=1.875
r236 37 40 44.0233 $w=2.48e-07 $l=9.55e-07 $layer=LI1_cond $X=4.58 $Y=0.92
+ $X2=4.58 $Y2=1.875
r237 31 49 6.17653 $w=4.15e-07 $l=1.57003e-07 $layer=LI1_cond $X=2.29 $Y=1.89
+ $X2=2.265 $Y2=2.035
r238 31 33 51.1685 $w=2.48e-07 $l=1.11e-06 $layer=LI1_cond $X=2.29 $Y=1.89
+ $X2=2.29 $Y2=0.78
r239 30 62 68.1959 $w=3.3e-07 $l=3.9e-07 $layer=POLY_cond $X=7.37 $Y=1.725
+ $X2=7.37 $Y2=1.335
r240 29 62 11.366 $w=3.3e-07 $l=6.5e-08 $layer=POLY_cond $X=7.37 $Y=1.27
+ $X2=7.37 $Y2=1.335
r241 26 65 39.4698 $w=3.94e-07 $l=2.09105e-07 $layer=POLY_cond $X=10.89 $Y=1.43
+ $X2=10.79 $Y2=1.595
r242 26 28 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=10.89 $Y=1.43
+ $X2=10.89 $Y2=1
r243 23 65 49.8683 $w=3.94e-07 $l=3.10242e-07 $layer=POLY_cond $X=10.655
+ $Y=1.845 $X2=10.79 $Y2=1.595
r244 23 25 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=10.655 $Y=1.845
+ $X2=10.655 $Y2=2.34
r245 20 22 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=7.9 $Y=1.925
+ $X2=7.9 $Y2=2.42
r246 19 30 32.1775 $w=1.5e-07 $l=1.98997e-07 $layer=POLY_cond $X=7.535 $Y=1.8
+ $X2=7.37 $Y2=1.725
r247 18 20 26.9307 $w=1.5e-07 $l=1.63936e-07 $layer=POLY_cond $X=7.81 $Y=1.8
+ $X2=7.9 $Y2=1.925
r248 18 19 141.011 $w=1.5e-07 $l=2.75e-07 $layer=POLY_cond $X=7.81 $Y=1.8
+ $X2=7.535 $Y2=1.8
r249 16 29 32.1775 $w=1.5e-07 $l=1.98997e-07 $layer=POLY_cond $X=7.205 $Y=1.195
+ $X2=7.37 $Y2=1.27
r250 16 17 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=7.205 $Y=1.195
+ $X2=6.595 $Y2=1.195
r251 13 17 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=6.52 $Y=1.12
+ $X2=6.595 $Y2=1.195
r252 13 15 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=6.52 $Y=1.12
+ $X2=6.52 $Y2=0.725
r253 4 53 300 $w=1.7e-07 $l=2.26164e-07 $layer=licon1_PDIFF $count=2 $X=4.365
+ $Y=1.895 $X2=4.53 $Y2=2.04
r254 3 80 600 $w=1.7e-07 $l=2.61534e-07 $layer=licon1_PDIFF $count=1 $X=2.15
+ $Y=2.09 $X2=2.32 $Y2=2.28
r255 2 37 182 $w=1.7e-07 $l=3.9702e-07 $layer=licon1_NDIFF $count=1 $X=4.38
+ $Y=0.595 $X2=4.54 $Y2=0.92
r256 1 33 182 $w=1.7e-07 $l=4.68348e-07 $layer=licon1_NDIFF $count=1 $X=2.195
+ $Y=0.37 $X2=2.32 $Y2=0.78
.ends

.subckt PM_SKY130_FD_SC_HS__FAHCIN_1%CIN 1 3 4 6 7 9 10 12 13 20
r59 18 20 44.5028 $w=3.52e-07 $l=3.25e-07 $layer=POLY_cond $X=8.87 $Y=1.46
+ $X2=9.195 $Y2=1.46
r60 16 18 39.0256 $w=3.52e-07 $l=2.85e-07 $layer=POLY_cond $X=8.585 $Y=1.46
+ $X2=8.87 $Y2=1.46
r61 15 16 13.0085 $w=3.52e-07 $l=9.5e-08 $layer=POLY_cond $X=8.49 $Y=1.46
+ $X2=8.585 $Y2=1.46
r62 13 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.87
+ $Y=1.32 $X2=8.87 $Y2=1.32
r63 10 20 37.6562 $w=3.52e-07 $l=2.75e-07 $layer=POLY_cond $X=9.47 $Y=1.46
+ $X2=9.195 $Y2=1.46
r64 10 12 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=9.47 $Y=1.395
+ $X2=9.47 $Y2=0.95
r65 7 20 22.7654 $w=1.5e-07 $l=3.05e-07 $layer=POLY_cond $X=9.195 $Y=1.765
+ $X2=9.195 $Y2=1.46
r66 7 9 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=9.195 $Y=1.765
+ $X2=9.195 $Y2=2.4
r67 4 16 22.7654 $w=1.5e-07 $l=3.05e-07 $layer=POLY_cond $X=8.585 $Y=1.155
+ $X2=8.585 $Y2=1.46
r68 4 6 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=8.585 $Y=1.155
+ $X2=8.585 $Y2=0.725
r69 1 15 22.7654 $w=1.5e-07 $l=3.05e-07 $layer=POLY_cond $X=8.49 $Y=1.765
+ $X2=8.49 $Y2=1.46
r70 1 3 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=8.49 $Y=1.765
+ $X2=8.49 $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_HS__FAHCIN_1%A_1854_368# 1 2 3 10 12 13 15 19 22 27 28
+ 31 33 34 35 38 39 42 44
r95 42 48 9.98619 $w=3.62e-07 $l=7.5e-08 $layer=POLY_cond $X=11.7 $Y=1.557
+ $X2=11.775 $Y2=1.557
r96 42 46 31.2901 $w=3.62e-07 $l=2.35e-07 $layer=POLY_cond $X=11.7 $Y=1.557
+ $X2=11.465 $Y2=1.557
r97 41 44 6.63528 $w=3.28e-07 $l=1.9e-07 $layer=LI1_cond $X=11.7 $Y=1.515
+ $X2=11.89 $Y2=1.515
r98 41 42 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=11.7
+ $Y=1.515 $X2=11.7 $Y2=1.515
r99 37 39 8.98215 $w=3.33e-07 $l=1.8e-07 $layer=LI1_cond $X=10.975 $Y=2.907
+ $X2=11.155 $Y2=2.907
r100 37 38 8.81015 $w=3.33e-07 $l=1.75e-07 $layer=LI1_cond $X=10.975 $Y=2.907
+ $X2=10.8 $Y2=2.907
r101 34 35 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=9.64 $Y=1.995
+ $X2=9.64 $Y2=1.34
r102 33 34 7.30169 $w=4.68e-07 $l=8.5e-08 $layer=LI1_cond $X=9.49 $Y=2.08
+ $X2=9.49 $Y2=1.995
r103 30 44 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.89 $Y=1.68
+ $X2=11.89 $Y2=1.515
r104 30 31 79.9198 $w=1.68e-07 $l=1.225e-06 $layer=LI1_cond $X=11.89 $Y=1.68
+ $X2=11.89 $Y2=2.905
r105 28 31 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=11.805 $Y=2.99
+ $X2=11.89 $Y2=2.905
r106 28 39 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=11.805 $Y=2.99
+ $X2=11.155 $Y2=2.99
r107 27 38 70.1337 $w=1.68e-07 $l=1.075e-06 $layer=LI1_cond $X=9.725 $Y=2.99
+ $X2=10.8 $Y2=2.99
r108 20 35 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=9.72 $Y=1.175
+ $X2=9.72 $Y2=1.34
r109 20 22 12.2229 $w=3.28e-07 $l=3.5e-07 $layer=LI1_cond $X=9.72 $Y=1.175
+ $X2=9.72 $Y2=0.825
r110 17 27 8.97637 $w=1.7e-07 $l=2.74226e-07 $layer=LI1_cond $X=9.49 $Y=2.905
+ $X2=9.725 $Y2=2.99
r111 17 19 2.29036 $w=4.68e-07 $l=9e-08 $layer=LI1_cond $X=9.49 $Y=2.905
+ $X2=9.49 $Y2=2.815
r112 16 33 3.81727 $w=4.68e-07 $l=1.5e-07 $layer=LI1_cond $X=9.49 $Y=2.23
+ $X2=9.49 $Y2=2.08
r113 16 19 14.8874 $w=4.68e-07 $l=5.85e-07 $layer=LI1_cond $X=9.49 $Y=2.23
+ $X2=9.49 $Y2=2.815
r114 13 48 23.4391 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=11.775 $Y=1.765
+ $X2=11.775 $Y2=1.557
r115 13 15 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=11.775 $Y=1.765
+ $X2=11.775 $Y2=2.34
r116 10 46 23.4391 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=11.465 $Y=1.35
+ $X2=11.465 $Y2=1.557
r117 10 12 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=11.465 $Y=1.35
+ $X2=11.465 $Y2=0.92
r118 3 37 600 $w=1.7e-07 $l=1.1007e-06 $layer=licon1_PDIFF $count=1 $X=10.73
+ $Y=1.92 $X2=10.975 $Y2=2.905
r119 2 33 400 $w=1.7e-07 $l=3.05941e-07 $layer=licon1_PDIFF $count=1 $X=9.27
+ $Y=1.84 $X2=9.42 $Y2=2.08
r120 2 19 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=9.27
+ $Y=1.84 $X2=9.42 $Y2=2.815
r121 1 22 91 $w=1.7e-07 $l=3.2078e-07 $layer=licon1_NDIFF $count=2 $X=9.545
+ $Y=0.58 $X2=9.72 $Y2=0.825
.ends

.subckt PM_SKY130_FD_SC_HS__FAHCIN_1%A_2004_136# 1 2 7 9 10 12 15 18 19 20 22 23
+ 24 27 34
r83 33 34 3.56523 $w=5.18e-07 $l=1.55e-07 $layer=LI1_cond $X=10.675 $Y=1
+ $X2=10.83 $Y2=1
r84 30 33 6.55543 $w=5.18e-07 $l=2.85e-07 $layer=LI1_cond $X=10.39 $Y=1
+ $X2=10.675 $Y2=1
r85 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=12.285
+ $Y=1.515 $X2=12.285 $Y2=1.515
r86 25 27 13.7882 $w=2.78e-07 $l=3.35e-07 $layer=LI1_cond $X=12.285 $Y=1.18
+ $X2=12.285 $Y2=1.515
r87 23 25 7.36005 $w=1.7e-07 $l=1.77482e-07 $layer=LI1_cond $X=12.145 $Y=1.095
+ $X2=12.285 $Y2=1.18
r88 23 24 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=12.145 $Y=1.095
+ $X2=11.755 $Y2=1.095
r89 22 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=11.67 $Y=1.01
+ $X2=11.755 $Y2=1.095
r90 21 22 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=11.67 $Y=0.49
+ $X2=11.67 $Y2=1.01
r91 19 21 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=11.585 $Y=0.405
+ $X2=11.67 $Y2=0.49
r92 19 20 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=11.585 $Y=0.405
+ $X2=10.915 $Y2=0.405
r93 18 34 7.40362 $w=1.7e-07 $l=2.6e-07 $layer=LI1_cond $X=10.83 $Y=0.74
+ $X2=10.83 $Y2=1
r94 17 20 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=10.83 $Y=0.49
+ $X2=10.915 $Y2=0.405
r95 17 18 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=10.83 $Y=0.49
+ $X2=10.83 $Y2=0.74
r96 13 30 5.03516 $w=2.5e-07 $l=2.6e-07 $layer=LI1_cond $X=10.39 $Y=1.26
+ $X2=10.39 $Y2=1
r97 13 15 37.1087 $w=2.48e-07 $l=8.05e-07 $layer=LI1_cond $X=10.39 $Y=1.26
+ $X2=10.39 $Y2=2.065
r98 10 28 39.1188 $w=3.74e-07 $l=2.21743e-07 $layer=POLY_cond $X=12.465 $Y=1.35
+ $X2=12.332 $Y2=1.515
r99 10 12 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=12.465 $Y=1.35
+ $X2=12.465 $Y2=0.87
r100 7 28 50.0734 $w=3.74e-07 $l=3.05369e-07 $layer=POLY_cond $X=12.455 $Y=1.765
+ $X2=12.332 $Y2=1.515
r101 7 9 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=12.455 $Y=1.765
+ $X2=12.455 $Y2=2.4
r102 2 15 600 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=10.28
+ $Y=1.92 $X2=10.43 $Y2=2.065
r103 1 33 45.5 $w=1.7e-07 $l=7.23878e-07 $layer=licon1_NDIFF $count=4 $X=10.02
+ $Y=0.68 $X2=10.675 $Y2=0.825
.ends

.subckt PM_SKY130_FD_SC_HS__FAHCIN_1%VPWR 1 2 3 4 15 21 25 29 34 35 36 38 43 58
+ 67 68 71 74 77
r99 77 78 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.24 $Y=3.33
+ $X2=12.24 $Y2=3.33
r100 74 75 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r101 71 72 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r102 68 78 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.72 $Y=3.33
+ $X2=12.24 $Y2=3.33
r103 67 68 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.72 $Y=3.33
+ $X2=12.72 $Y2=3.33
r104 65 77 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=12.395 $Y=3.33
+ $X2=12.27 $Y2=3.33
r105 65 67 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=12.395 $Y=3.33
+ $X2=12.72 $Y2=3.33
r106 64 78 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.76 $Y=3.33
+ $X2=12.24 $Y2=3.33
r107 63 64 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=11.76 $Y=3.33
+ $X2=11.76 $Y2=3.33
r108 61 64 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=9.36 $Y=3.33
+ $X2=11.76 $Y2=3.33
r109 60 63 156.578 $w=1.68e-07 $l=2.4e-06 $layer=LI1_cond $X=9.36 $Y=3.33
+ $X2=11.76 $Y2=3.33
r110 60 61 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=9.36 $Y=3.33
+ $X2=9.36 $Y2=3.33
r111 58 77 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=12.145 $Y=3.33
+ $X2=12.27 $Y2=3.33
r112 58 63 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=12.145 $Y=3.33
+ $X2=11.76 $Y2=3.33
r113 57 61 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=3.33
+ $X2=9.36 $Y2=3.33
r114 56 57 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r115 54 75 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=3.33 $X2=5.52
+ $Y2=3.33
r116 53 56 187.893 $w=1.68e-07 $l=2.88e-06 $layer=LI1_cond $X=6 $Y=3.33 $X2=8.88
+ $Y2=3.33
r117 53 54 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=6 $Y=3.33
+ $X2=6 $Y2=3.33
r118 51 74 9.14399 $w=1.7e-07 $l=1.8e-07 $layer=LI1_cond $X=5.765 $Y=3.33
+ $X2=5.585 $Y2=3.33
r119 51 53 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=5.765 $Y=3.33
+ $X2=6 $Y2=3.33
r120 50 75 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=5.52 $Y2=3.33
r121 49 50 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r122 47 50 1.07034 $w=4.9e-07 $l=3.84e-06 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=5.04 $Y2=3.33
r123 47 72 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r124 46 49 250.524 $w=1.68e-07 $l=3.84e-06 $layer=LI1_cond $X=1.2 $Y=3.33
+ $X2=5.04 $Y2=3.33
r125 46 47 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r126 44 71 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.825 $Y=3.33
+ $X2=0.7 $Y2=3.33
r127 44 46 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=0.825 $Y=3.33
+ $X2=1.2 $Y2=3.33
r128 43 74 9.14399 $w=1.7e-07 $l=1.8e-07 $layer=LI1_cond $X=5.405 $Y=3.33
+ $X2=5.585 $Y2=3.33
r129 43 49 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=5.405 $Y=3.33
+ $X2=5.04 $Y2=3.33
r130 41 72 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r131 40 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r132 38 71 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.575 $Y=3.33
+ $X2=0.7 $Y2=3.33
r133 38 40 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=0.575 $Y=3.33
+ $X2=0.24 $Y2=3.33
r134 36 57 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=8.88 $Y2=3.33
r135 36 54 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=3.33 $X2=6
+ $Y2=3.33
r136 34 56 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=8.885 $Y=3.33
+ $X2=8.88 $Y2=3.33
r137 34 35 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.885 $Y=3.33
+ $X2=8.97 $Y2=3.33
r138 33 60 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=9.055 $Y=3.33
+ $X2=9.36 $Y2=3.33
r139 33 35 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.055 $Y=3.33
+ $X2=8.97 $Y2=3.33
r140 29 32 36.8782 $w=2.48e-07 $l=8e-07 $layer=LI1_cond $X=12.27 $Y=2.015
+ $X2=12.27 $Y2=2.815
r141 27 77 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=12.27 $Y=3.245
+ $X2=12.27 $Y2=3.33
r142 27 32 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=12.27 $Y=3.245
+ $X2=12.27 $Y2=2.815
r143 23 35 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.97 $Y=3.245
+ $X2=8.97 $Y2=3.33
r144 23 25 70.7861 $w=1.68e-07 $l=1.085e-06 $layer=LI1_cond $X=8.97 $Y=3.245
+ $X2=8.97 $Y2=2.16
r145 19 74 1.16013 $w=3.6e-07 $l=8.5e-08 $layer=LI1_cond $X=5.585 $Y=3.245
+ $X2=5.585 $Y2=3.33
r146 19 21 13.7653 $w=3.58e-07 $l=4.3e-07 $layer=LI1_cond $X=5.585 $Y=3.245
+ $X2=5.585 $Y2=2.815
r147 15 18 32.2684 $w=2.48e-07 $l=7e-07 $layer=LI1_cond $X=0.7 $Y=2.115 $X2=0.7
+ $Y2=2.815
r148 13 71 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.7 $Y=3.245
+ $X2=0.7 $Y2=3.33
r149 13 18 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=0.7 $Y=3.245 $X2=0.7
+ $Y2=2.815
r150 4 32 400 $w=1.7e-07 $l=1.1494e-06 $layer=licon1_PDIFF $count=1 $X=11.85
+ $Y=1.84 $X2=12.23 $Y2=2.815
r151 4 29 400 $w=1.7e-07 $l=4.59238e-07 $layer=licon1_PDIFF $count=1 $X=11.85
+ $Y=1.84 $X2=12.23 $Y2=2.015
r152 3 25 300 $w=1.7e-07 $l=5.41872e-07 $layer=licon1_PDIFF $count=2 $X=8.565
+ $Y=1.84 $X2=8.97 $Y2=2.16
r153 2 21 600 $w=1.7e-07 $l=1.05428e-06 $layer=licon1_PDIFF $count=1 $X=5.42
+ $Y=1.84 $X2=5.585 $Y2=2.815
r154 1 18 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=0.59
+ $Y=1.84 $X2=0.74 $Y2=2.815
r155 1 15 400 $w=1.7e-07 $l=3.4187e-07 $layer=licon1_PDIFF $count=1 $X=0.59
+ $Y=1.84 $X2=0.74 $Y2=2.115
.ends

.subckt PM_SKY130_FD_SC_HS__FAHCIN_1%A_256_368# 1 2 3 4 14 17 18 19 20 22 26 27
+ 28 31 34 35 39 41 46
c94 46 0 9.05624e-20 $X=3.09 $Y=1.005
c95 41 0 1.89903e-19 $X=2.817 $Y=2.045
c96 28 0 1.01566e-19 $X=3.175 $Y=0.34
r97 44 46 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=2.895 $Y=1.005
+ $X2=3.09 $Y2=1.005
r98 37 39 2.84554 $w=4.03e-07 $l=1e-07 $layer=LI1_cond $X=1.625 $Y=0.817
+ $X2=1.725 $Y2=0.817
r99 34 35 7.7063 $w=4.88e-07 $l=1.65e-07 $layer=LI1_cond $X=1.59 $Y=1.985
+ $X2=1.59 $Y2=1.82
r100 29 31 21.8964 $w=2.48e-07 $l=4.75e-07 $layer=LI1_cond $X=3.82 $Y=0.425
+ $X2=3.82 $Y2=0.9
r101 27 29 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=3.695 $Y=0.34
+ $X2=3.82 $Y2=0.425
r102 27 28 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=3.695 $Y=0.34
+ $X2=3.175 $Y2=0.34
r103 26 46 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.09 $Y=0.92
+ $X2=3.09 $Y2=1.005
r104 25 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.09 $Y=0.425
+ $X2=3.175 $Y2=0.34
r105 25 26 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=3.09 $Y=0.425
+ $X2=3.09 $Y2=0.92
r106 23 44 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.895 $Y=1.09
+ $X2=2.895 $Y2=1.005
r107 23 41 62.3048 $w=1.68e-07 $l=9.55e-07 $layer=LI1_cond $X=2.895 $Y=1.09
+ $X2=2.895 $Y2=2.045
r108 20 43 2.65806 $w=3.25e-07 $l=8.5e-08 $layer=LI1_cond $X=2.817 $Y=2.565
+ $X2=2.817 $Y2=2.65
r109 20 22 12.0563 $w=3.23e-07 $l=3.4e-07 $layer=LI1_cond $X=2.817 $Y=2.565
+ $X2=2.817 $Y2=2.225
r110 19 41 8.35379 $w=3.23e-07 $l=1.62e-07 $layer=LI1_cond $X=2.817 $Y=2.207
+ $X2=2.817 $Y2=2.045
r111 19 22 0.638276 $w=3.23e-07 $l=1.8e-08 $layer=LI1_cond $X=2.817 $Y=2.207
+ $X2=2.817 $Y2=2.225
r112 17 43 5.06595 $w=1.7e-07 $l=1.62e-07 $layer=LI1_cond $X=2.655 $Y=2.65
+ $X2=2.817 $Y2=2.65
r113 17 18 53.4973 $w=1.68e-07 $l=8.2e-07 $layer=LI1_cond $X=2.655 $Y=2.65
+ $X2=1.835 $Y2=2.65
r114 15 39 4.30998 $w=2.2e-07 $l=2.03e-07 $layer=LI1_cond $X=1.725 $Y=1.02
+ $X2=1.725 $Y2=0.817
r115 15 35 41.907 $w=2.18e-07 $l=8e-07 $layer=LI1_cond $X=1.725 $Y=1.02
+ $X2=1.725 $Y2=1.82
r116 14 18 9.14635 $w=1.7e-07 $l=2.84341e-07 $layer=LI1_cond $X=1.59 $Y=2.565
+ $X2=1.835 $Y2=2.65
r117 13 34 1.95278 $w=4.88e-07 $l=8e-08 $layer=LI1_cond $X=1.59 $Y=2.065
+ $X2=1.59 $Y2=1.985
r118 13 14 12.2049 $w=4.88e-07 $l=5e-07 $layer=LI1_cond $X=1.59 $Y=2.065
+ $X2=1.59 $Y2=2.565
r119 4 43 600 $w=1.7e-07 $l=6.48074e-07 $layer=licon1_PDIFF $count=1 $X=2.625
+ $Y=2.09 $X2=2.815 $Y2=2.65
r120 4 22 600 $w=1.7e-07 $l=2.48495e-07 $layer=licon1_PDIFF $count=1 $X=2.625
+ $Y=2.09 $X2=2.815 $Y2=2.225
r121 3 34 300 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=2 $X=1.28
+ $Y=1.84 $X2=1.43 $Y2=1.985
r122 2 31 182 $w=1.7e-07 $l=3.68409e-07 $layer=licon1_NDIFF $count=1 $X=3.72
+ $Y=0.595 $X2=3.86 $Y2=0.9
r123 1 37 182 $w=1.7e-07 $l=4.09054e-07 $layer=licon1_NDIFF $count=1 $X=1.485
+ $Y=0.47 $X2=1.625 $Y2=0.815
.ends

.subckt PM_SKY130_FD_SC_HS__FAHCIN_1%A_1197_368# 1 2 9 14 15 17
r37 15 17 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=6.225 $Y=1.82
+ $X2=6.225 $Y2=1.065
r38 14 15 10.8446 $w=3.38e-07 $l=2.35e-07 $layer=LI1_cond $X=6.14 $Y=2.055
+ $X2=6.14 $Y2=1.82
r39 7 17 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=6.305 $Y=0.9
+ $X2=6.305 $Y2=1.065
r40 7 9 12.2229 $w=3.28e-07 $l=3.5e-07 $layer=LI1_cond $X=6.305 $Y=0.9 $X2=6.305
+ $Y2=0.55
r41 2 14 600 $w=1.7e-07 $l=2.80134e-07 $layer=licon1_PDIFF $count=1 $X=5.985
+ $Y=1.84 $X2=6.135 $Y2=2.055
r42 1 9 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=6.165
+ $Y=0.405 $X2=6.305 $Y2=0.55
.ends

.subckt PM_SKY130_FD_SC_HS__FAHCIN_1%COUT 1 2 8 11 14 21 22
c47 14 0 1.63318e-19 $X=6.805 $Y=0.56
r48 21 22 9.43695 $w=5.43e-07 $l=4.3e-07 $layer=LI1_cond $X=7.44 $Y=0.712
+ $X2=7.87 $Y2=0.712
r49 21 26 6.14499 $w=5.43e-07 $l=2.8e-07 $layer=LI1_cond $X=7.44 $Y=0.712
+ $X2=7.16 $Y2=0.712
r50 17 26 1.97518 $w=5.43e-07 $l=9e-08 $layer=LI1_cond $X=7.07 $Y=0.712 $X2=7.16
+ $Y2=0.712
r51 17 18 20.3897 $w=4.28e-07 $l=5.98e-07 $layer=LI1_cond $X=6.855 $Y=0.712
+ $X2=6.855 $Y2=1.31
r52 14 17 4.07375 $w=4.28e-07 $l=1.52e-07 $layer=LI1_cond $X=6.855 $Y=0.56
+ $X2=6.855 $Y2=0.712
r53 9 20 2.94173 $w=3.3e-07 $l=1.25e-07 $layer=LI1_cond $X=7.07 $Y=2.5 $X2=6.945
+ $Y2=2.5
r54 9 11 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=7.07 $Y=2.5 $X2=7.5
+ $Y2=2.5
r55 8 20 4.82444 $w=1.7e-07 $l=1.83916e-07 $layer=LI1_cond $X=6.985 $Y=2.335
+ $X2=6.945 $Y2=2.5
r56 8 18 66.8717 $w=1.68e-07 $l=1.025e-06 $layer=LI1_cond $X=6.985 $Y=2.335
+ $X2=6.985 $Y2=1.31
r57 2 20 600 $w=1.7e-07 $l=6.5192e-07 $layer=licon1_PDIFF $count=1 $X=6.57 $Y=2
+ $X2=6.92 $Y2=2.5
r58 2 11 600 $w=1.7e-07 $l=1.15321e-06 $layer=licon1_PDIFF $count=1 $X=6.57 $Y=2
+ $X2=7.5 $Y2=2.5
r59 1 22 60.6667 $w=1.7e-07 $l=1.35028e-06 $layer=licon1_NDIFF $count=3 $X=6.595
+ $Y=0.405 $X2=7.87 $Y2=0.56
r60 1 26 60.6667 $w=1.7e-07 $l=6.37809e-07 $layer=licon1_NDIFF $count=3 $X=6.595
+ $Y=0.405 $X2=7.16 $Y2=0.56
r61 1 14 91 $w=1.7e-07 $l=2.76857e-07 $layer=licon1_NDIFF $count=2 $X=6.595
+ $Y=0.405 $X2=6.805 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HS__FAHCIN_1%A_1595_400# 1 2 7 9 13 17 18
r29 17 18 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=8.29 $Y=1.82
+ $X2=8.29 $Y2=1.065
r30 11 18 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=8.37 $Y=0.9
+ $X2=8.37 $Y2=1.065
r31 11 13 12.2229 $w=3.28e-07 $l=3.5e-07 $layer=LI1_cond $X=8.37 $Y=0.9 $X2=8.37
+ $Y2=0.55
r32 7 17 6.94937 $w=2.48e-07 $l=1.25e-07 $layer=LI1_cond $X=8.25 $Y=1.945
+ $X2=8.25 $Y2=1.82
r33 7 9 1.84391 $w=2.48e-07 $l=4e-08 $layer=LI1_cond $X=8.25 $Y=1.945 $X2=8.25
+ $Y2=1.985
r34 2 9 300 $w=1.7e-07 $l=2.42384e-07 $layer=licon1_PDIFF $count=2 $X=7.975 $Y=2
+ $X2=8.21 $Y2=1.985
r35 1 13 91 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=2 $X=8.16
+ $Y=0.405 $X2=8.37 $Y2=0.55
.ends

.subckt PM_SKY130_FD_SC_HS__FAHCIN_1%A_1967_384# 1 2 3 10 12 14 18 20 23 29 30
c50 20 0 8.64817e-20 $X=11.28 $Y=1.25
r51 29 30 8.83531 $w=4.38e-07 $l=1.65e-07 $layer=LI1_cond $X=11.415 $Y=2.015
+ $X2=11.415 $Y2=1.85
r52 22 29 1.44055 $w=4.38e-07 $l=5.5e-08 $layer=LI1_cond $X=11.415 $Y=2.07
+ $X2=11.415 $Y2=2.015
r53 22 23 8.64332 $w=4.38e-07 $l=3.3e-07 $layer=LI1_cond $X=11.415 $Y=2.07
+ $X2=11.415 $Y2=2.4
r54 20 27 7.81924 $w=3.22e-07 $l=1.49248e-07 $layer=LI1_cond $X=11.28 $Y=1.25
+ $X2=11.25 $Y2=1.115
r55 20 30 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=11.28 $Y=1.25
+ $X2=11.28 $Y2=1.85
r56 16 27 2.21818 $w=3.3e-07 $l=6e-08 $layer=LI1_cond $X=11.25 $Y=1.055
+ $X2=11.25 $Y2=1.115
r57 16 18 10.826 $w=3.28e-07 $l=3.1e-07 $layer=LI1_cond $X=11.25 $Y=1.055
+ $X2=11.25 $Y2=0.745
r58 15 25 3.40825 $w=1.7e-07 $l=1.19143e-07 $layer=LI1_cond $X=10.065 $Y=2.485
+ $X2=9.98 $Y2=2.567
r59 14 23 14.5445 $w=1.82e-07 $l=2.59037e-07 $layer=LI1_cond $X=11.195 $Y=2.485
+ $X2=11.415 $Y2=2.4
r60 14 15 73.7219 $w=1.68e-07 $l=1.13e-06 $layer=LI1_cond $X=11.195 $Y=2.485
+ $X2=10.065 $Y2=2.485
r61 10 25 3.40825 $w=1.7e-07 $l=1.67e-07 $layer=LI1_cond $X=9.98 $Y=2.4 $X2=9.98
+ $Y2=2.567
r62 10 12 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=9.98 $Y=2.4
+ $X2=9.98 $Y2=2.065
r63 3 29 300 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=2 $X=11.405
+ $Y=1.84 $X2=11.55 $Y2=2.015
r64 2 25 600 $w=1.7e-07 $l=7.18853e-07 $layer=licon1_PDIFF $count=1 $X=9.835
+ $Y=1.92 $X2=9.98 $Y2=2.57
r65 2 12 600 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=9.835
+ $Y=1.92 $X2=9.98 $Y2=2.065
r66 1 27 182 $w=1.7e-07 $l=5.59643e-07 $layer=licon1_NDIFF $count=1 $X=10.965
+ $Y=0.68 $X2=11.25 $Y2=1.115
r67 1 18 182 $w=1.7e-07 $l=3.15832e-07 $layer=licon1_NDIFF $count=1 $X=10.965
+ $Y=0.68 $X2=11.25 $Y2=0.745
.ends

.subckt PM_SKY130_FD_SC_HS__FAHCIN_1%SUM 1 2 7 8 9 10 11 12 13
r14 12 13 17.0562 $w=2.48e-07 $l=3.7e-07 $layer=LI1_cond $X=12.72 $Y=2.405
+ $X2=12.72 $Y2=2.775
r15 11 12 19.361 $w=2.48e-07 $l=4.2e-07 $layer=LI1_cond $X=12.72 $Y=1.985
+ $X2=12.72 $Y2=2.405
r16 10 11 14.7513 $w=2.48e-07 $l=3.2e-07 $layer=LI1_cond $X=12.72 $Y=1.665
+ $X2=12.72 $Y2=1.985
r17 9 10 17.0562 $w=2.48e-07 $l=3.7e-07 $layer=LI1_cond $X=12.72 $Y=1.295
+ $X2=12.72 $Y2=1.665
r18 9 26 9.21954 $w=2.48e-07 $l=2e-07 $layer=LI1_cond $X=12.72 $Y=1.295
+ $X2=12.72 $Y2=1.095
r19 8 44 5.50001 $w=4.18e-07 $l=1.8e-07 $layer=LI1_cond $X=12.68 $Y=0.84
+ $X2=12.68 $Y2=0.66
r20 8 26 7.83661 $w=2.48e-07 $l=1.7e-07 $layer=LI1_cond $X=12.72 $Y=0.925
+ $X2=12.72 $Y2=1.095
r21 7 44 3.66686 $w=3.28e-07 $l=1.05e-07 $layer=LI1_cond $X=12.68 $Y=0.555
+ $X2=12.68 $Y2=0.66
r22 2 13 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=12.53
+ $Y=1.84 $X2=12.68 $Y2=2.815
r23 2 11 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=12.53
+ $Y=1.84 $X2=12.68 $Y2=1.985
r24 1 44 182 $w=1.7e-07 $l=2.19089e-07 $layer=licon1_NDIFF $count=1 $X=12.54
+ $Y=0.5 $X2=12.68 $Y2=0.66
r25 1 26 182 $w=1.7e-07 $l=6.61306e-07 $layer=licon1_NDIFF $count=1 $X=12.54
+ $Y=0.5 $X2=12.68 $Y2=1.095
.ends

.subckt PM_SKY130_FD_SC_HS__FAHCIN_1%VGND 1 2 3 4 15 19 23 27 29 31 36 41 49 59
+ 60 63 66 69 72
c116 19 0 1.27399e-19 $X=5.715 $Y=0.55
r117 72 73 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.24 $Y=0
+ $X2=12.24 $Y2=0
r118 69 70 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=0 $X2=8.88
+ $Y2=0
r119 66 67 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r120 63 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r121 60 73 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.72 $Y=0
+ $X2=12.24 $Y2=0
r122 59 60 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.72 $Y=0
+ $X2=12.72 $Y2=0
r123 57 72 10.1275 $w=1.7e-07 $l=2.1e-07 $layer=LI1_cond $X=12.345 $Y=0
+ $X2=12.135 $Y2=0
r124 57 59 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=12.345 $Y=0
+ $X2=12.72 $Y2=0
r125 56 73 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.76 $Y=0
+ $X2=12.24 $Y2=0
r126 55 56 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=11.76 $Y=0
+ $X2=11.76 $Y2=0
r127 53 56 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=9.36 $Y=0
+ $X2=11.76 $Y2=0
r128 53 70 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.36 $Y=0 $X2=8.88
+ $Y2=0
r129 52 55 156.578 $w=1.68e-07 $l=2.4e-06 $layer=LI1_cond $X=9.36 $Y=0 $X2=11.76
+ $Y2=0
r130 52 53 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=9.36 $Y=0 $X2=9.36
+ $Y2=0
r131 50 69 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=9.045 $Y=0 $X2=8.875
+ $Y2=0
r132 50 52 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=9.045 $Y=0
+ $X2=9.36 $Y2=0
r133 49 72 10.1275 $w=1.7e-07 $l=2.1e-07 $layer=LI1_cond $X=11.925 $Y=0
+ $X2=12.135 $Y2=0
r134 49 55 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=11.925 $Y=0
+ $X2=11.76 $Y2=0
r135 48 70 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=0 $X2=8.88
+ $Y2=0
r136 47 48 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r137 45 67 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=0 $X2=5.52
+ $Y2=0
r138 44 47 156.578 $w=1.68e-07 $l=2.4e-06 $layer=LI1_cond $X=6 $Y=0 $X2=8.4
+ $Y2=0
r139 44 45 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=6 $Y=0 $X2=6 $Y2=0
r140 42 66 11.3601 $w=1.7e-07 $l=2.53e-07 $layer=LI1_cond $X=5.97 $Y=0 $X2=5.717
+ $Y2=0
r141 42 44 1.95722 $w=1.68e-07 $l=3e-08 $layer=LI1_cond $X=5.97 $Y=0 $X2=6 $Y2=0
r142 41 69 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=8.705 $Y=0 $X2=8.875
+ $Y2=0
r143 41 47 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=8.705 $Y=0 $X2=8.4
+ $Y2=0
r144 40 67 1.20413 $w=4.9e-07 $l=4.32e-06 $layer=MET1_cond $X=1.2 $Y=0 $X2=5.52
+ $Y2=0
r145 40 64 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r146 39 40 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r147 37 63 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.95 $Y=0 $X2=0.785
+ $Y2=0
r148 37 39 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=0.95 $Y=0 $X2=1.2
+ $Y2=0
r149 36 66 11.3601 $w=1.7e-07 $l=2.52e-07 $layer=LI1_cond $X=5.465 $Y=0
+ $X2=5.717 $Y2=0
r150 36 39 278.251 $w=1.68e-07 $l=4.265e-06 $layer=LI1_cond $X=5.465 $Y=0
+ $X2=1.2 $Y2=0
r151 34 64 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r152 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r153 31 63 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.62 $Y=0 $X2=0.785
+ $Y2=0
r154 31 33 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=0.62 $Y=0 $X2=0.24
+ $Y2=0
r155 29 48 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=6.48 $Y=0 $X2=8.4
+ $Y2=0
r156 29 45 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=0 $X2=6
+ $Y2=0
r157 25 72 1.60615 $w=4.2e-07 $l=8.5e-08 $layer=LI1_cond $X=12.135 $Y=0.085
+ $X2=12.135 $Y2=0
r158 25 27 15.3659 $w=4.18e-07 $l=5.6e-07 $layer=LI1_cond $X=12.135 $Y=0.085
+ $X2=12.135 $Y2=0.645
r159 21 69 0.987631 $w=3.4e-07 $l=8.5e-08 $layer=LI1_cond $X=8.875 $Y=0.085
+ $X2=8.875 $Y2=0
r160 21 23 15.7614 $w=3.38e-07 $l=4.65e-07 $layer=LI1_cond $X=8.875 $Y=0.085
+ $X2=8.875 $Y2=0.55
r161 17 66 2.09999 $w=5.05e-07 $l=8.5e-08 $layer=LI1_cond $X=5.717 $Y=0.085
+ $X2=5.717 $Y2=0
r162 17 19 11.0134 $w=5.03e-07 $l=4.65e-07 $layer=LI1_cond $X=5.717 $Y=0.085
+ $X2=5.717 $Y2=0.55
r163 13 63 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.785 $Y=0.085
+ $X2=0.785 $Y2=0
r164 13 15 20.6043 $w=3.28e-07 $l=5.9e-07 $layer=LI1_cond $X=0.785 $Y=0.085
+ $X2=0.785 $Y2=0.675
r165 4 27 182 $w=1.7e-07 $l=5.77062e-07 $layer=licon1_NDIFF $count=1 $X=11.54
+ $Y=0.6 $X2=12.095 $Y2=0.645
r166 3 23 91 $w=1.7e-07 $l=2.78209e-07 $layer=licon1_NDIFF $count=2 $X=8.66
+ $Y=0.405 $X2=8.875 $Y2=0.55
r167 2 19 182 $w=1.7e-07 $l=3.44964e-07 $layer=licon1_NDIFF $count=1 $X=5.435
+ $Y=0.405 $X2=5.715 $Y2=0.55
r168 1 15 182 $w=1.7e-07 $l=3.96327e-07 $layer=licon1_NDIFF $count=1 $X=0.575
+ $Y=0.37 $X2=0.785 $Y2=0.675
.ends

