* File: sky130_fd_sc_hs__o2111ai_4.pxi.spice
* Created: Tue Sep  1 20:13:29 2020
* 
x_PM_SKY130_FD_SC_HS__O2111AI_4%D1 N_D1_c_140_n N_D1_M1011_g N_D1_c_141_n
+ N_D1_M1013_g N_D1_c_146_n N_D1_M1020_g N_D1_c_142_n N_D1_M1030_g N_D1_c_147_n
+ N_D1_M1024_g N_D1_c_143_n N_D1_M1033_g D1 D1 D1 N_D1_c_145_n
+ PM_SKY130_FD_SC_HS__O2111AI_4%D1
x_PM_SKY130_FD_SC_HS__O2111AI_4%C1 N_C1_c_208_n N_C1_M1003_g N_C1_c_200_n
+ N_C1_M1000_g N_C1_c_201_n N_C1_M1008_g N_C1_c_209_n N_C1_M1022_g N_C1_c_202_n
+ N_C1_M1026_g N_C1_c_203_n N_C1_c_204_n N_C1_c_205_n N_C1_M1028_g C1
+ N_C1_c_207_n PM_SKY130_FD_SC_HS__O2111AI_4%C1
x_PM_SKY130_FD_SC_HS__O2111AI_4%B1 N_B1_c_286_n N_B1_M1002_g N_B1_c_276_n
+ N_B1_c_277_n N_B1_c_289_n N_B1_M1005_g N_B1_M1009_g N_B1_M1014_g N_B1_M1027_g
+ N_B1_c_281_n N_B1_M1032_g N_B1_c_283_n B1 B1 B1 B1 N_B1_c_285_n
+ PM_SKY130_FD_SC_HS__O2111AI_4%B1
x_PM_SKY130_FD_SC_HS__O2111AI_4%A1 N_A1_c_369_n N_A1_M1007_g N_A1_M1004_g
+ N_A1_c_370_n N_A1_M1010_g N_A1_M1006_g N_A1_c_371_n N_A1_M1015_g N_A1_M1012_g
+ N_A1_c_372_n N_A1_M1025_g N_A1_M1023_g A1 A1 A1 N_A1_c_373_n N_A1_c_368_n
+ PM_SKY130_FD_SC_HS__O2111AI_4%A1
x_PM_SKY130_FD_SC_HS__O2111AI_4%A2 N_A2_c_457_n N_A2_M1016_g N_A2_c_451_n
+ N_A2_M1001_g N_A2_c_458_n N_A2_M1017_g N_A2_c_452_n N_A2_M1018_g N_A2_c_459_n
+ N_A2_M1019_g N_A2_c_453_n N_A2_M1021_g N_A2_c_460_n N_A2_M1029_g N_A2_c_454_n
+ N_A2_M1031_g A2 A2 A2 A2 N_A2_c_455_n N_A2_c_456_n
+ PM_SKY130_FD_SC_HS__O2111AI_4%A2
x_PM_SKY130_FD_SC_HS__O2111AI_4%Y N_Y_M1011_s N_Y_M1030_s N_Y_M1020_d
+ N_Y_M1024_d N_Y_M1022_d N_Y_M1005_d N_Y_M1016_d N_Y_M1019_d N_Y_c_534_n
+ N_Y_c_551_n N_Y_c_554_n N_Y_c_535_n N_Y_c_537_n N_Y_c_538_n N_Y_c_536_n
+ N_Y_c_540_n N_Y_c_581_n N_Y_c_541_n N_Y_c_542_n N_Y_c_610_n N_Y_c_543_n
+ N_Y_c_544_n N_Y_c_545_n N_Y_c_614_n N_Y_c_618_n Y
+ PM_SKY130_FD_SC_HS__O2111AI_4%Y
x_PM_SKY130_FD_SC_HS__O2111AI_4%VPWR N_VPWR_M1020_s N_VPWR_M1003_s
+ N_VPWR_M1002_s N_VPWR_M1007_s N_VPWR_M1015_s N_VPWR_c_669_n N_VPWR_c_670_n
+ N_VPWR_c_671_n N_VPWR_c_672_n N_VPWR_c_673_n N_VPWR_c_674_n N_VPWR_c_675_n
+ N_VPWR_c_676_n N_VPWR_c_677_n VPWR N_VPWR_c_678_n N_VPWR_c_679_n
+ N_VPWR_c_680_n N_VPWR_c_681_n N_VPWR_c_668_n N_VPWR_c_683_n N_VPWR_c_684_n
+ N_VPWR_c_685_n PM_SKY130_FD_SC_HS__O2111AI_4%VPWR
x_PM_SKY130_FD_SC_HS__O2111AI_4%A_954_368# N_A_954_368#_M1007_d
+ N_A_954_368#_M1010_d N_A_954_368#_M1025_d N_A_954_368#_M1017_s
+ N_A_954_368#_M1029_s N_A_954_368#_c_767_n N_A_954_368#_c_776_n
+ N_A_954_368#_c_778_n N_A_954_368#_c_780_n N_A_954_368#_c_781_n
+ N_A_954_368#_c_768_n N_A_954_368#_c_769_n N_A_954_368#_c_792_n
+ N_A_954_368#_c_770_n N_A_954_368#_c_771_n N_A_954_368#_c_772_n
+ N_A_954_368#_c_773_n N_A_954_368#_c_774_n
+ PM_SKY130_FD_SC_HS__O2111AI_4%A_954_368#
x_PM_SKY130_FD_SC_HS__O2111AI_4%A_27_74# N_A_27_74#_M1011_d N_A_27_74#_M1013_d
+ N_A_27_74#_M1033_d N_A_27_74#_M1008_d N_A_27_74#_M1028_d N_A_27_74#_c_835_n
+ N_A_27_74#_c_836_n N_A_27_74#_c_837_n N_A_27_74#_c_838_n N_A_27_74#_c_839_n
+ PM_SKY130_FD_SC_HS__O2111AI_4%A_27_74#
x_PM_SKY130_FD_SC_HS__O2111AI_4%A_472_74# N_A_472_74#_M1000_s
+ N_A_472_74#_M1026_s N_A_472_74#_M1009_d N_A_472_74#_M1027_d
+ N_A_472_74#_c_882_n N_A_472_74#_c_883_n
+ PM_SKY130_FD_SC_HS__O2111AI_4%A_472_74#
x_PM_SKY130_FD_SC_HS__O2111AI_4%A_841_74# N_A_841_74#_M1009_s
+ N_A_841_74#_M1014_s N_A_841_74#_M1032_s N_A_841_74#_M1006_d
+ N_A_841_74#_M1023_d N_A_841_74#_M1018_d N_A_841_74#_M1031_d
+ N_A_841_74#_c_910_n N_A_841_74#_c_911_n N_A_841_74#_c_912_n
+ N_A_841_74#_c_913_n N_A_841_74#_c_914_n N_A_841_74#_c_915_n
+ N_A_841_74#_c_916_n N_A_841_74#_c_917_n N_A_841_74#_c_918_n
+ N_A_841_74#_c_919_n N_A_841_74#_c_920_n N_A_841_74#_c_921_n
+ N_A_841_74#_c_922_n N_A_841_74#_c_923_n N_A_841_74#_c_924_n
+ N_A_841_74#_c_925_n N_A_841_74#_c_926_n
+ PM_SKY130_FD_SC_HS__O2111AI_4%A_841_74#
x_PM_SKY130_FD_SC_HS__O2111AI_4%VGND N_VGND_M1004_s N_VGND_M1012_s
+ N_VGND_M1001_s N_VGND_M1021_s N_VGND_c_1018_n N_VGND_c_1019_n N_VGND_c_1020_n
+ N_VGND_c_1021_n VGND N_VGND_c_1022_n N_VGND_c_1023_n N_VGND_c_1024_n
+ N_VGND_c_1025_n N_VGND_c_1026_n N_VGND_c_1027_n N_VGND_c_1028_n
+ N_VGND_c_1029_n N_VGND_c_1030_n N_VGND_c_1031_n
+ PM_SKY130_FD_SC_HS__O2111AI_4%VGND
cc_1 VNB N_D1_c_140_n 0.0210761f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.185
cc_2 VNB N_D1_c_141_n 0.0155697f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=1.185
cc_3 VNB N_D1_c_142_n 0.015f $X=-0.19 $Y=-0.245 $X2=1.425 $Y2=1.185
cc_4 VNB N_D1_c_143_n 0.0151994f $X=-0.19 $Y=-0.245 $X2=1.855 $Y2=1.185
cc_5 VNB D1 0.0152189f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.58
cc_6 VNB N_D1_c_145_n 0.128767f $X=-0.19 $Y=-0.245 $X2=1.81 $Y2=1.475
cc_7 VNB N_C1_c_200_n 0.0154191f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=1.185
cc_8 VNB N_C1_c_201_n 0.0150343f $X=-0.19 $Y=-0.245 $X2=1.26 $Y2=1.765
cc_9 VNB N_C1_c_202_n 0.0150343f $X=-0.19 $Y=-0.245 $X2=1.81 $Y2=1.765
cc_10 VNB N_C1_c_203_n 0.0258382f $X=-0.19 $Y=-0.245 $X2=1.855 $Y2=1.185
cc_11 VNB N_C1_c_204_n 0.0733837f $X=-0.19 $Y=-0.245 $X2=1.855 $Y2=0.74
cc_12 VNB N_C1_c_205_n 0.0204573f $X=-0.19 $Y=-0.245 $X2=1.855 $Y2=0.74
cc_13 VNB C1 0.00693045f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=1.475
cc_14 VNB N_C1_c_207_n 0.0083658f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_B1_c_276_n 0.0138303f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=1.185
cc_16 VNB N_B1_c_277_n 0.00535301f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=0.74
cc_17 VNB N_B1_M1009_g 0.0326175f $X=-0.19 $Y=-0.245 $X2=1.81 $Y2=1.765
cc_18 VNB N_B1_M1014_g 0.0232165f $X=-0.19 $Y=-0.245 $X2=1.855 $Y2=0.74
cc_19 VNB N_B1_M1027_g 0.0230075f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.58
cc_20 VNB N_B1_c_281_n 0.0647671f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_B1_M1032_g 0.0244321f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.475
cc_22 VNB N_B1_c_283_n 0.00678423f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.515
cc_23 VNB B1 0.00643414f $X=-0.19 $Y=-0.245 $X2=1.185 $Y2=1.515
cc_24 VNB N_B1_c_285_n 0.0097572f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.565
cc_25 VNB N_A1_M1004_g 0.0237205f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=0.74
cc_26 VNB N_A1_M1006_g 0.021878f $X=-0.19 $Y=-0.245 $X2=1.81 $Y2=1.765
cc_27 VNB N_A1_M1012_g 0.0209643f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_28 VNB N_A1_M1023_g 0.0211601f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.515
cc_29 VNB N_A1_c_368_n 0.083687f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A2_c_451_n 0.0176036f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=1.185
cc_31 VNB N_A2_c_452_n 0.0175325f $X=-0.19 $Y=-0.245 $X2=1.425 $Y2=1.185
cc_32 VNB N_A2_c_453_n 0.0168814f $X=-0.19 $Y=-0.245 $X2=1.855 $Y2=1.185
cc_33 VNB N_A2_c_454_n 0.0218115f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A2_c_455_n 0.0037039f $X=-0.19 $Y=-0.245 $X2=1.2 $Y2=1.565
cc_35 VNB N_A2_c_456_n 0.11937f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_Y_c_534_n 0.00752994f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.475
cc_37 VNB N_Y_c_535_n 5.13074e-19 $X=-0.19 $Y=-0.245 $X2=1.185 $Y2=1.515
cc_38 VNB N_Y_c_536_n 0.00418294f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_VPWR_c_668_n 0.422413f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_27_74#_c_835_n 0.00813147f $X=-0.19 $Y=-0.245 $X2=1.855 $Y2=0.74
cc_41 VNB N_A_27_74#_c_836_n 0.00159969f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_27_74#_c_837_n 0.00288661f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_27_74#_c_838_n 0.012662f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.515
cc_44 VNB N_A_27_74#_c_839_n 0.036321f $X=-0.19 $Y=-0.245 $X2=1.185 $Y2=1.515
cc_45 VNB N_A_472_74#_c_882_n 0.002374f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_A_472_74#_c_883_n 0.0262662f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_841_74#_c_910_n 0.00382328f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_841_74#_c_911_n 0.00114016f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.515
cc_49 VNB N_A_841_74#_c_912_n 0.00279782f $X=-0.19 $Y=-0.245 $X2=1.185 $Y2=1.475
cc_50 VNB N_A_841_74#_c_913_n 0.00315816f $X=-0.19 $Y=-0.245 $X2=1.185 $Y2=1.515
cc_51 VNB N_A_841_74#_c_914_n 0.00178908f $X=-0.19 $Y=-0.245 $X2=1.855 $Y2=1.475
cc_52 VNB N_A_841_74#_c_915_n 0.00374231f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_A_841_74#_c_916_n 0.00206666f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_A_841_74#_c_917_n 0.00313208f $X=-0.19 $Y=-0.245 $X2=1.2 $Y2=1.565
cc_55 VNB N_A_841_74#_c_918_n 0.00253603f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_A_841_74#_c_919_n 0.0164817f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_A_841_74#_c_920_n 0.0266107f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_A_841_74#_c_921_n 0.00675567f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_A_841_74#_c_922_n 0.00250234f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_A_841_74#_c_923_n 0.00478213f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_A_841_74#_c_924_n 0.00126364f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_A_841_74#_c_925_n 0.00186907f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_A_841_74#_c_926_n 0.00172073f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_VGND_c_1018_n 0.00567996f $X=-0.19 $Y=-0.245 $X2=1.81 $Y2=2.4
cc_65 VNB N_VGND_c_1019_n 0.002601f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_66 VNB N_VGND_c_1020_n 0.00495983f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_VGND_c_1021_n 0.00334323f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.515
cc_68 VNB N_VGND_c_1022_n 0.162661f $X=-0.19 $Y=-0.245 $X2=1.185 $Y2=1.515
cc_69 VNB N_VGND_c_1023_n 0.0151736f $X=-0.19 $Y=-0.245 $X2=1.855 $Y2=1.475
cc_70 VNB N_VGND_c_1024_n 0.0169342f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.565
cc_71 VNB N_VGND_c_1025_n 0.0170944f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_VGND_c_1026_n 0.0173909f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_VGND_c_1027_n 0.525959f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_VGND_c_1028_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_VGND_c_1029_n 0.00604233f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_VGND_c_1030_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_VGND_c_1031_n 0.00604233f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VPB N_D1_c_146_n 0.0216043f $X=-0.19 $Y=1.66 $X2=1.26 $Y2=1.765
cc_79 VPB N_D1_c_147_n 0.0161232f $X=-0.19 $Y=1.66 $X2=1.81 $Y2=1.765
cc_80 VPB D1 0.0159123f $X=-0.19 $Y=1.66 $X2=1.115 $Y2=1.58
cc_81 VPB N_D1_c_145_n 0.0390354f $X=-0.19 $Y=1.66 $X2=1.81 $Y2=1.475
cc_82 VPB N_C1_c_208_n 0.0177341f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.185
cc_83 VPB N_C1_c_209_n 0.0177454f $X=-0.19 $Y=1.66 $X2=1.425 $Y2=1.185
cc_84 VPB N_C1_c_204_n 0.0338685f $X=-0.19 $Y=1.66 $X2=1.855 $Y2=0.74
cc_85 VPB C1 0.00143888f $X=-0.19 $Y=1.66 $X2=0.995 $Y2=1.475
cc_86 VPB N_B1_c_286_n 0.0163813f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.185
cc_87 VPB N_B1_c_276_n 0.011442f $X=-0.19 $Y=1.66 $X2=0.995 $Y2=1.185
cc_88 VPB N_B1_c_277_n 0.00553782f $X=-0.19 $Y=1.66 $X2=0.995 $Y2=0.74
cc_89 VPB N_B1_c_289_n 0.0214852f $X=-0.19 $Y=1.66 $X2=0.995 $Y2=0.74
cc_90 VPB N_B1_c_281_n 0.0517945f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_91 VPB N_B1_c_283_n 0.00438579f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.515
cc_92 VPB B1 0.0166777f $X=-0.19 $Y=1.66 $X2=1.185 $Y2=1.515
cc_93 VPB N_B1_c_285_n 0.00827427f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=1.565
cc_94 VPB N_A1_c_369_n 0.0207692f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.185
cc_95 VPB N_A1_c_370_n 0.0156298f $X=-0.19 $Y=1.66 $X2=1.26 $Y2=2.4
cc_96 VPB N_A1_c_371_n 0.0155127f $X=-0.19 $Y=1.66 $X2=1.81 $Y2=2.4
cc_97 VPB N_A1_c_372_n 0.0154299f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_98 VPB N_A1_c_373_n 0.00854133f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_99 VPB N_A1_c_368_n 0.047378f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_100 VPB N_A2_c_457_n 0.0151582f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.185
cc_101 VPB N_A2_c_458_n 0.0153208f $X=-0.19 $Y=1.66 $X2=1.26 $Y2=1.765
cc_102 VPB N_A2_c_459_n 0.0154263f $X=-0.19 $Y=1.66 $X2=1.81 $Y2=1.765
cc_103 VPB N_A2_c_460_n 0.0188241f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_104 VPB N_A2_c_455_n 0.012396f $X=-0.19 $Y=1.66 $X2=1.2 $Y2=1.565
cc_105 VPB N_A2_c_456_n 0.0507282f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_106 VPB N_Y_c_537_n 0.00257348f $X=-0.19 $Y=1.66 $X2=1.81 $Y2=1.475
cc_107 VPB N_Y_c_538_n 0.00459604f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=1.565
cc_108 VPB N_Y_c_536_n 0.00581265f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_109 VPB N_Y_c_540_n 0.00257348f $X=-0.19 $Y=1.66 $X2=0.72 $Y2=1.565
cc_110 VPB N_Y_c_541_n 0.0168372f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_111 VPB N_Y_c_542_n 0.0111346f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_112 VPB N_Y_c_543_n 0.0529354f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_113 VPB N_Y_c_544_n 0.0021196f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_114 VPB N_Y_c_545_n 2.51882e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_115 VPB N_VPWR_c_669_n 0.00899981f $X=-0.19 $Y=1.66 $X2=1.855 $Y2=0.74
cc_116 VPB N_VPWR_c_670_n 0.0116684f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_117 VPB N_VPWR_c_671_n 0.00900305f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.475
cc_118 VPB N_VPWR_c_672_n 0.00891904f $X=-0.19 $Y=1.66 $X2=1.185 $Y2=1.475
cc_119 VPB N_VPWR_c_673_n 0.00769929f $X=-0.19 $Y=1.66 $X2=1.425 $Y2=1.475
cc_120 VPB N_VPWR_c_674_n 0.0372801f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=1.565
cc_121 VPB N_VPWR_c_675_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_122 VPB N_VPWR_c_676_n 0.0186948f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.565
cc_123 VPB N_VPWR_c_677_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0.72 $Y2=1.565
cc_124 VPB N_VPWR_c_678_n 0.0186948f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_125 VPB N_VPWR_c_679_n 0.0600098f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_126 VPB N_VPWR_c_680_n 0.0206041f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_127 VPB N_VPWR_c_681_n 0.0625814f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_128 VPB N_VPWR_c_668_n 0.115774f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_129 VPB N_VPWR_c_683_n 0.0124767f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_130 VPB N_VPWR_c_684_n 0.0047828f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_131 VPB N_VPWR_c_685_n 0.00324402f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_132 VPB N_A_954_368#_c_767_n 0.0162776f $X=-0.19 $Y=1.66 $X2=1.855 $Y2=1.185
cc_133 VPB N_A_954_368#_c_768_n 0.00262732f $X=-0.19 $Y=1.66 $X2=1.185 $Y2=1.475
cc_134 VPB N_A_954_368#_c_769_n 0.0022931f $X=-0.19 $Y=1.66 $X2=1.185 $Y2=1.515
cc_135 VPB N_A_954_368#_c_770_n 0.0123062f $X=-0.19 $Y=1.66 $X2=1.855 $Y2=1.475
cc_136 VPB N_A_954_368#_c_771_n 0.0443668f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.565
cc_137 VPB N_A_954_368#_c_772_n 0.00331232f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_138 VPB N_A_954_368#_c_773_n 0.00257417f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_139 VPB N_A_954_368#_c_774_n 0.0022931f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_140 N_D1_c_147_n N_C1_c_208_n 0.0100458f $X=1.81 $Y=1.765 $X2=-0.19
+ $Y2=-0.245
cc_141 N_D1_c_143_n N_C1_c_200_n 0.0100279f $X=1.855 $Y=1.185 $X2=0 $Y2=0
cc_142 N_D1_c_145_n N_C1_c_204_n 0.0287625f $X=1.81 $Y=1.475 $X2=0 $Y2=0
cc_143 N_D1_c_145_n N_C1_c_207_n 0.0012731f $X=1.81 $Y=1.475 $X2=0 $Y2=0
cc_144 N_D1_c_140_n N_Y_c_534_n 0.00194106f $X=0.495 $Y=1.185 $X2=0 $Y2=0
cc_145 N_D1_c_141_n N_Y_c_534_n 0.0140453f $X=0.995 $Y=1.185 $X2=0 $Y2=0
cc_146 N_D1_c_142_n N_Y_c_534_n 0.0185273f $X=1.425 $Y=1.185 $X2=0 $Y2=0
cc_147 D1 N_Y_c_534_n 0.0486045f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_148 N_D1_c_145_n N_Y_c_534_n 0.00809939f $X=1.81 $Y=1.475 $X2=0 $Y2=0
cc_149 N_D1_c_146_n N_Y_c_551_n 0.0125195f $X=1.26 $Y=1.765 $X2=0 $Y2=0
cc_150 N_D1_c_147_n N_Y_c_551_n 0.012264f $X=1.81 $Y=1.765 $X2=0 $Y2=0
cc_151 N_D1_c_145_n N_Y_c_551_n 0.00788958f $X=1.81 $Y=1.475 $X2=0 $Y2=0
cc_152 N_D1_c_143_n N_Y_c_554_n 0.00436059f $X=1.855 $Y=1.185 $X2=0 $Y2=0
cc_153 N_D1_c_142_n N_Y_c_535_n 0.00135929f $X=1.425 $Y=1.185 $X2=0 $Y2=0
cc_154 N_D1_c_143_n N_Y_c_535_n 0.00141132f $X=1.855 $Y=1.185 $X2=0 $Y2=0
cc_155 D1 N_Y_c_535_n 0.0128263f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_156 N_D1_c_145_n N_Y_c_535_n 0.0259502f $X=1.81 $Y=1.475 $X2=0 $Y2=0
cc_157 N_D1_c_146_n N_Y_c_537_n 6.63386e-19 $X=1.26 $Y=1.765 $X2=0 $Y2=0
cc_158 N_D1_c_147_n N_Y_c_537_n 0.0109196f $X=1.81 $Y=1.765 $X2=0 $Y2=0
cc_159 N_D1_c_146_n N_Y_c_536_n 3.76014e-19 $X=1.26 $Y=1.765 $X2=0 $Y2=0
cc_160 N_D1_c_147_n N_Y_c_536_n 0.00452802f $X=1.81 $Y=1.765 $X2=0 $Y2=0
cc_161 D1 N_Y_c_536_n 0.0162205f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_162 N_D1_c_145_n N_Y_c_536_n 0.019f $X=1.81 $Y=1.475 $X2=0 $Y2=0
cc_163 N_D1_c_146_n N_Y_c_543_n 0.0115985f $X=1.26 $Y=1.765 $X2=0 $Y2=0
cc_164 N_D1_c_147_n N_Y_c_543_n 6.59344e-19 $X=1.81 $Y=1.765 $X2=0 $Y2=0
cc_165 D1 N_Y_c_543_n 0.10241f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_166 N_D1_c_145_n N_Y_c_543_n 0.00496069f $X=1.81 $Y=1.475 $X2=0 $Y2=0
cc_167 N_D1_c_146_n N_VPWR_c_669_n 0.00739417f $X=1.26 $Y=1.765 $X2=0 $Y2=0
cc_168 N_D1_c_147_n N_VPWR_c_669_n 0.00598632f $X=1.81 $Y=1.765 $X2=0 $Y2=0
cc_169 N_D1_c_146_n N_VPWR_c_674_n 0.00444483f $X=1.26 $Y=1.765 $X2=0 $Y2=0
cc_170 N_D1_c_147_n N_VPWR_c_678_n 0.00445602f $X=1.81 $Y=1.765 $X2=0 $Y2=0
cc_171 N_D1_c_146_n N_VPWR_c_668_n 0.00858941f $X=1.26 $Y=1.765 $X2=0 $Y2=0
cc_172 N_D1_c_147_n N_VPWR_c_668_n 0.00857881f $X=1.81 $Y=1.765 $X2=0 $Y2=0
cc_173 N_D1_c_140_n N_A_27_74#_c_835_n 0.0134011f $X=0.495 $Y=1.185 $X2=0 $Y2=0
cc_174 N_D1_c_141_n N_A_27_74#_c_835_n 0.0107985f $X=0.995 $Y=1.185 $X2=0 $Y2=0
cc_175 N_D1_c_142_n N_A_27_74#_c_835_n 0.0101492f $X=1.425 $Y=1.185 $X2=0 $Y2=0
cc_176 N_D1_c_143_n N_A_27_74#_c_835_n 0.0141739f $X=1.855 $Y=1.185 $X2=0 $Y2=0
cc_177 N_D1_c_145_n N_A_27_74#_c_835_n 3.08096e-19 $X=1.81 $Y=1.475 $X2=0 $Y2=0
cc_178 N_D1_c_140_n N_A_27_74#_c_839_n 0.0101315f $X=0.495 $Y=1.185 $X2=0 $Y2=0
cc_179 N_D1_c_141_n N_A_27_74#_c_839_n 8.60984e-19 $X=0.995 $Y=1.185 $X2=0 $Y2=0
cc_180 D1 N_A_27_74#_c_839_n 0.0234201f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_181 N_D1_c_145_n N_A_27_74#_c_839_n 0.00240493f $X=1.81 $Y=1.475 $X2=0 $Y2=0
cc_182 N_D1_c_140_n N_VGND_c_1022_n 0.00291626f $X=0.495 $Y=1.185 $X2=0 $Y2=0
cc_183 N_D1_c_141_n N_VGND_c_1022_n 0.00291649f $X=0.995 $Y=1.185 $X2=0 $Y2=0
cc_184 N_D1_c_142_n N_VGND_c_1022_n 0.00291649f $X=1.425 $Y=1.185 $X2=0 $Y2=0
cc_185 N_D1_c_143_n N_VGND_c_1022_n 0.00291649f $X=1.855 $Y=1.185 $X2=0 $Y2=0
cc_186 N_D1_c_140_n N_VGND_c_1027_n 0.00363419f $X=0.495 $Y=1.185 $X2=0 $Y2=0
cc_187 N_D1_c_141_n N_VGND_c_1027_n 0.00359779f $X=0.995 $Y=1.185 $X2=0 $Y2=0
cc_188 N_D1_c_142_n N_VGND_c_1027_n 0.00359121f $X=1.425 $Y=1.185 $X2=0 $Y2=0
cc_189 N_D1_c_143_n N_VGND_c_1027_n 0.00359219f $X=1.855 $Y=1.185 $X2=0 $Y2=0
cc_190 N_C1_c_209_n N_B1_c_286_n 0.0104167f $X=3.13 $Y=1.765 $X2=-0.19
+ $Y2=-0.245
cc_191 C1 N_B1_c_286_n 2.70636e-19 $X=3.995 $Y=1.58 $X2=-0.19 $Y2=-0.245
cc_192 C1 N_B1_c_276_n 0.00771269f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_193 N_C1_c_207_n N_B1_c_276_n 0.0106597f $X=3.965 $Y=1.54 $X2=0 $Y2=0
cc_194 N_C1_c_203_n N_B1_c_277_n 0.00883813f $X=3.5 $Y=1.26 $X2=0 $Y2=0
cc_195 N_C1_c_204_n N_B1_c_277_n 0.0111343f $X=3.22 $Y=1.26 $X2=0 $Y2=0
cc_196 C1 N_B1_c_277_n 7.93677e-19 $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_197 N_C1_c_207_n N_B1_c_277_n 0.00680233f $X=3.965 $Y=1.54 $X2=0 $Y2=0
cc_198 C1 N_B1_c_289_n 0.00237643f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_199 C1 N_B1_M1009_g 0.00178986f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_200 C1 N_B1_c_281_n 0.00151851f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_201 C1 N_B1_c_283_n 0.0092271f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_202 C1 B1 0.0281684f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_203 N_C1_c_200_n N_Y_c_535_n 9.37775e-19 $X=2.285 $Y=1.185 $X2=0 $Y2=0
cc_204 N_C1_c_204_n N_Y_c_535_n 2.73078e-19 $X=3.22 $Y=1.26 $X2=0 $Y2=0
cc_205 N_C1_c_207_n N_Y_c_535_n 0.00960541f $X=3.965 $Y=1.54 $X2=0 $Y2=0
cc_206 N_C1_c_208_n N_Y_c_537_n 0.0101743f $X=2.26 $Y=1.765 $X2=0 $Y2=0
cc_207 N_C1_c_208_n N_Y_c_538_n 0.0135553f $X=2.26 $Y=1.765 $X2=0 $Y2=0
cc_208 N_C1_c_209_n N_Y_c_538_n 0.0140508f $X=3.13 $Y=1.765 $X2=0 $Y2=0
cc_209 N_C1_c_204_n N_Y_c_538_n 0.0209171f $X=3.22 $Y=1.26 $X2=0 $Y2=0
cc_210 N_C1_c_207_n N_Y_c_538_n 0.0726736f $X=3.965 $Y=1.54 $X2=0 $Y2=0
cc_211 N_C1_c_208_n N_Y_c_536_n 0.00894692f $X=2.26 $Y=1.765 $X2=0 $Y2=0
cc_212 N_C1_c_204_n N_Y_c_536_n 0.00478153f $X=3.22 $Y=1.26 $X2=0 $Y2=0
cc_213 N_C1_c_207_n N_Y_c_536_n 0.00684868f $X=3.965 $Y=1.54 $X2=0 $Y2=0
cc_214 N_C1_c_209_n N_Y_c_540_n 0.0101743f $X=3.13 $Y=1.765 $X2=0 $Y2=0
cc_215 C1 N_Y_c_581_n 0.0150694f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_216 N_C1_c_207_n N_Y_c_581_n 0.0185458f $X=3.965 $Y=1.54 $X2=0 $Y2=0
cc_217 N_C1_c_209_n N_Y_c_544_n 0.00784674f $X=3.13 $Y=1.765 $X2=0 $Y2=0
cc_218 N_C1_c_203_n N_Y_c_544_n 0.00113801f $X=3.5 $Y=1.26 $X2=0 $Y2=0
cc_219 N_C1_c_204_n N_Y_c_544_n 4.80986e-19 $X=3.22 $Y=1.26 $X2=0 $Y2=0
cc_220 N_C1_c_207_n N_Y_c_544_n 0.028649f $X=3.965 $Y=1.54 $X2=0 $Y2=0
cc_221 C1 N_Y_c_545_n 4.10242e-19 $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_222 N_C1_c_208_n N_VPWR_c_670_n 0.00377044f $X=2.26 $Y=1.765 $X2=0 $Y2=0
cc_223 N_C1_c_209_n N_VPWR_c_670_n 0.00377044f $X=3.13 $Y=1.765 $X2=0 $Y2=0
cc_224 N_C1_c_209_n N_VPWR_c_676_n 0.00445602f $X=3.13 $Y=1.765 $X2=0 $Y2=0
cc_225 N_C1_c_208_n N_VPWR_c_678_n 0.00445602f $X=2.26 $Y=1.765 $X2=0 $Y2=0
cc_226 N_C1_c_208_n N_VPWR_c_668_n 0.00859788f $X=2.26 $Y=1.765 $X2=0 $Y2=0
cc_227 N_C1_c_209_n N_VPWR_c_668_n 0.00859788f $X=3.13 $Y=1.765 $X2=0 $Y2=0
cc_228 N_C1_c_200_n N_A_27_74#_c_838_n 0.0137455f $X=2.285 $Y=1.185 $X2=0 $Y2=0
cc_229 N_C1_c_201_n N_A_27_74#_c_838_n 0.0124572f $X=2.715 $Y=1.185 $X2=0 $Y2=0
cc_230 N_C1_c_202_n N_A_27_74#_c_838_n 0.0125299f $X=3.145 $Y=1.185 $X2=0 $Y2=0
cc_231 N_C1_c_203_n N_A_27_74#_c_838_n 0.00223574f $X=3.5 $Y=1.26 $X2=0 $Y2=0
cc_232 N_C1_c_204_n N_A_27_74#_c_838_n 0.00662756f $X=3.22 $Y=1.26 $X2=0 $Y2=0
cc_233 N_C1_c_205_n N_A_27_74#_c_838_n 0.0125731f $X=3.575 $Y=1.185 $X2=0 $Y2=0
cc_234 N_C1_c_207_n N_A_27_74#_c_838_n 0.136338f $X=3.965 $Y=1.54 $X2=0 $Y2=0
cc_235 N_C1_c_200_n N_A_472_74#_c_883_n 0.00382836f $X=2.285 $Y=1.185 $X2=0
+ $Y2=0
cc_236 N_C1_c_201_n N_A_472_74#_c_883_n 0.0114018f $X=2.715 $Y=1.185 $X2=0 $Y2=0
cc_237 N_C1_c_202_n N_A_472_74#_c_883_n 0.0114018f $X=3.145 $Y=1.185 $X2=0 $Y2=0
cc_238 N_C1_c_205_n N_A_472_74#_c_883_n 0.0149606f $X=3.575 $Y=1.185 $X2=0 $Y2=0
cc_239 N_C1_c_207_n N_A_472_74#_c_883_n 0.00760162f $X=3.965 $Y=1.54 $X2=0 $Y2=0
cc_240 N_C1_c_205_n N_A_841_74#_c_921_n 6.761e-19 $X=3.575 $Y=1.185 $X2=0 $Y2=0
cc_241 C1 N_A_841_74#_c_921_n 8.54022e-19 $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_242 N_C1_c_200_n N_VGND_c_1022_n 0.00433162f $X=2.285 $Y=1.185 $X2=0 $Y2=0
cc_243 N_C1_c_201_n N_VGND_c_1022_n 0.00291649f $X=2.715 $Y=1.185 $X2=0 $Y2=0
cc_244 N_C1_c_202_n N_VGND_c_1022_n 0.00291649f $X=3.145 $Y=1.185 $X2=0 $Y2=0
cc_245 N_C1_c_205_n N_VGND_c_1022_n 0.00291649f $X=3.575 $Y=1.185 $X2=0 $Y2=0
cc_246 N_C1_c_200_n N_VGND_c_1027_n 0.0044191f $X=2.285 $Y=1.185 $X2=0 $Y2=0
cc_247 N_C1_c_201_n N_VGND_c_1027_n 0.00359121f $X=2.715 $Y=1.185 $X2=0 $Y2=0
cc_248 N_C1_c_202_n N_VGND_c_1027_n 0.00359121f $X=3.145 $Y=1.185 $X2=0 $Y2=0
cc_249 N_C1_c_205_n N_VGND_c_1027_n 0.0036412f $X=3.575 $Y=1.185 $X2=0 $Y2=0
cc_250 B1 N_A1_c_369_n 2.97282e-19 $X=5.915 $Y=1.58 $X2=-0.19 $Y2=-0.245
cc_251 N_B1_M1032_g N_A1_M1004_g 0.0241978f $X=5.855 $Y=0.74 $X2=0 $Y2=0
cc_252 N_B1_c_281_n N_A1_c_373_n 2.81585e-19 $X=5.855 $Y=1.35 $X2=0 $Y2=0
cc_253 B1 N_A1_c_373_n 0.0381105f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_254 N_B1_M1032_g N_A1_c_368_n 0.0224536f $X=5.855 $Y=0.74 $X2=0 $Y2=0
cc_255 B1 N_A1_c_368_n 0.00429169f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_256 N_B1_c_286_n N_Y_c_540_n 0.0109304f $X=3.58 $Y=1.765 $X2=0 $Y2=0
cc_257 N_B1_c_286_n N_Y_c_581_n 0.0137395f $X=3.58 $Y=1.765 $X2=0 $Y2=0
cc_258 N_B1_c_276_n N_Y_c_581_n 0.0059407f $X=4.04 $Y=1.65 $X2=0 $Y2=0
cc_259 N_B1_c_289_n N_Y_c_581_n 0.0125195f $X=4.13 $Y=1.765 $X2=0 $Y2=0
cc_260 N_B1_c_286_n N_Y_c_541_n 6.63528e-19 $X=3.58 $Y=1.765 $X2=0 $Y2=0
cc_261 N_B1_c_289_n N_Y_c_541_n 0.0104f $X=4.13 $Y=1.765 $X2=0 $Y2=0
cc_262 N_B1_c_281_n N_Y_c_542_n 0.00847263f $X=5.855 $Y=1.35 $X2=0 $Y2=0
cc_263 B1 N_Y_c_542_n 0.127336f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_264 N_B1_c_286_n N_Y_c_544_n 0.00430581f $X=3.58 $Y=1.765 $X2=0 $Y2=0
cc_265 N_B1_c_277_n N_Y_c_544_n 3.70769e-19 $X=3.67 $Y=1.65 $X2=0 $Y2=0
cc_266 N_B1_c_289_n N_Y_c_544_n 0.00142903f $X=4.13 $Y=1.765 $X2=0 $Y2=0
cc_267 N_B1_c_289_n N_Y_c_545_n 7.26045e-19 $X=4.13 $Y=1.765 $X2=0 $Y2=0
cc_268 B1 N_Y_c_545_n 0.0066649f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_269 N_B1_c_285_n N_Y_c_545_n 0.00825538f $X=4.49 $Y=1.537 $X2=0 $Y2=0
cc_270 N_B1_c_286_n N_VPWR_c_671_n 0.00598632f $X=3.58 $Y=1.765 $X2=0 $Y2=0
cc_271 N_B1_c_289_n N_VPWR_c_671_n 0.00737447f $X=4.13 $Y=1.765 $X2=0 $Y2=0
cc_272 N_B1_c_286_n N_VPWR_c_676_n 0.00445602f $X=3.58 $Y=1.765 $X2=0 $Y2=0
cc_273 N_B1_c_289_n N_VPWR_c_679_n 0.00445602f $X=4.13 $Y=1.765 $X2=0 $Y2=0
cc_274 N_B1_c_286_n N_VPWR_c_668_n 0.00857881f $X=3.58 $Y=1.765 $X2=0 $Y2=0
cc_275 N_B1_c_289_n N_VPWR_c_668_n 0.00862599f $X=4.13 $Y=1.765 $X2=0 $Y2=0
cc_276 N_B1_c_289_n N_A_954_368#_c_767_n 0.00144273f $X=4.13 $Y=1.765 $X2=0
+ $Y2=0
cc_277 N_B1_c_277_n N_A_27_74#_c_838_n 0.00134885f $X=3.67 $Y=1.65 $X2=0 $Y2=0
cc_278 N_B1_M1009_g N_A_27_74#_c_838_n 6.87538e-19 $X=4.565 $Y=0.74 $X2=0 $Y2=0
cc_279 N_B1_M1027_g N_A_472_74#_c_882_n 0.00209099f $X=5.425 $Y=0.74 $X2=0 $Y2=0
cc_280 N_B1_M1032_g N_A_472_74#_c_882_n 0.00416883f $X=5.855 $Y=0.74 $X2=0 $Y2=0
cc_281 N_B1_M1009_g N_A_472_74#_c_883_n 0.0151398f $X=4.565 $Y=0.74 $X2=0 $Y2=0
cc_282 N_B1_M1014_g N_A_472_74#_c_883_n 0.0116171f $X=4.995 $Y=0.74 $X2=0 $Y2=0
cc_283 N_B1_M1027_g N_A_472_74#_c_883_n 0.0100664f $X=5.425 $Y=0.74 $X2=0 $Y2=0
cc_284 N_B1_M1027_g N_A_841_74#_c_910_n 0.0137239f $X=5.425 $Y=0.74 $X2=0 $Y2=0
cc_285 N_B1_c_281_n N_A_841_74#_c_910_n 0.00233808f $X=5.855 $Y=1.35 $X2=0 $Y2=0
cc_286 N_B1_M1032_g N_A_841_74#_c_910_n 0.0187194f $X=5.855 $Y=0.74 $X2=0 $Y2=0
cc_287 N_B1_M1009_g N_A_841_74#_c_911_n 2.36785e-19 $X=4.565 $Y=0.74 $X2=0 $Y2=0
cc_288 N_B1_M1014_g N_A_841_74#_c_911_n 0.00314204f $X=4.995 $Y=0.74 $X2=0 $Y2=0
cc_289 N_B1_c_281_n N_A_841_74#_c_911_n 0.00233553f $X=5.855 $Y=1.35 $X2=0 $Y2=0
cc_290 B1 N_A_841_74#_c_911_n 0.0738268f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_291 N_B1_M1032_g N_A_841_74#_c_912_n 0.00268885f $X=5.855 $Y=0.74 $X2=0 $Y2=0
cc_292 N_B1_M1009_g N_A_841_74#_c_921_n 0.00235917f $X=4.565 $Y=0.74 $X2=0 $Y2=0
cc_293 N_B1_c_283_n N_A_841_74#_c_921_n 0.006992f $X=4.13 $Y=1.67 $X2=0 $Y2=0
cc_294 B1 N_A_841_74#_c_921_n 0.0384622f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_295 N_B1_M1009_g N_A_841_74#_c_922_n 0.0104612f $X=4.565 $Y=0.74 $X2=0 $Y2=0
cc_296 N_B1_M1014_g N_A_841_74#_c_922_n 0.0104612f $X=4.995 $Y=0.74 $X2=0 $Y2=0
cc_297 N_B1_c_281_n N_A_841_74#_c_922_n 0.0022561f $X=5.855 $Y=1.35 $X2=0 $Y2=0
cc_298 B1 N_A_841_74#_c_923_n 0.0126236f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_299 N_B1_M1009_g N_VGND_c_1022_n 0.00291649f $X=4.565 $Y=0.74 $X2=0 $Y2=0
cc_300 N_B1_M1014_g N_VGND_c_1022_n 0.00291649f $X=4.995 $Y=0.74 $X2=0 $Y2=0
cc_301 N_B1_M1027_g N_VGND_c_1022_n 0.00291649f $X=5.425 $Y=0.74 $X2=0 $Y2=0
cc_302 N_B1_M1032_g N_VGND_c_1022_n 0.00433162f $X=5.855 $Y=0.74 $X2=0 $Y2=0
cc_303 N_B1_M1009_g N_VGND_c_1027_n 0.0036412f $X=4.565 $Y=0.74 $X2=0 $Y2=0
cc_304 N_B1_M1014_g N_VGND_c_1027_n 0.00359121f $X=4.995 $Y=0.74 $X2=0 $Y2=0
cc_305 N_B1_M1027_g N_VGND_c_1027_n 0.00359121f $X=5.425 $Y=0.74 $X2=0 $Y2=0
cc_306 N_B1_M1032_g N_VGND_c_1027_n 0.00449797f $X=5.855 $Y=0.74 $X2=0 $Y2=0
cc_307 N_A1_c_372_n N_A2_c_457_n 0.0256388f $X=7.625 $Y=1.765 $X2=-0.19
+ $Y2=-0.245
cc_308 N_A1_M1023_g N_A2_c_451_n 0.0131789f $X=7.715 $Y=0.74 $X2=0 $Y2=0
cc_309 N_A1_c_373_n N_A2_c_455_n 0.0381113f $X=7.47 $Y=1.515 $X2=0 $Y2=0
cc_310 N_A1_c_368_n N_A2_c_455_n 0.00370469f $X=7.625 $Y=1.542 $X2=0 $Y2=0
cc_311 N_A1_M1023_g N_A2_c_456_n 0.0174644f $X=7.715 $Y=0.74 $X2=0 $Y2=0
cc_312 N_A1_c_373_n N_A2_c_456_n 3.19861e-19 $X=7.47 $Y=1.515 $X2=0 $Y2=0
cc_313 N_A1_c_368_n N_A2_c_456_n 0.0126377f $X=7.625 $Y=1.542 $X2=0 $Y2=0
cc_314 N_A1_c_369_n N_Y_c_542_n 0.0156433f $X=6.26 $Y=1.765 $X2=0 $Y2=0
cc_315 N_A1_c_370_n N_Y_c_542_n 0.0108178f $X=6.725 $Y=1.765 $X2=0 $Y2=0
cc_316 N_A1_c_371_n N_Y_c_542_n 0.0107319f $X=7.175 $Y=1.765 $X2=0 $Y2=0
cc_317 N_A1_c_372_n N_Y_c_542_n 0.0127488f $X=7.625 $Y=1.765 $X2=0 $Y2=0
cc_318 N_A1_c_373_n N_Y_c_542_n 0.0921993f $X=7.47 $Y=1.515 $X2=0 $Y2=0
cc_319 N_A1_c_368_n N_Y_c_542_n 0.00572378f $X=7.625 $Y=1.542 $X2=0 $Y2=0
cc_320 N_A1_c_369_n N_VPWR_c_672_n 0.00324976f $X=6.26 $Y=1.765 $X2=0 $Y2=0
cc_321 N_A1_c_370_n N_VPWR_c_672_n 0.0041146f $X=6.725 $Y=1.765 $X2=0 $Y2=0
cc_322 N_A1_c_371_n N_VPWR_c_673_n 0.00379374f $X=7.175 $Y=1.765 $X2=0 $Y2=0
cc_323 N_A1_c_372_n N_VPWR_c_673_n 0.00224402f $X=7.625 $Y=1.765 $X2=0 $Y2=0
cc_324 N_A1_c_369_n N_VPWR_c_679_n 0.00460063f $X=6.26 $Y=1.765 $X2=0 $Y2=0
cc_325 N_A1_c_370_n N_VPWR_c_680_n 0.00445602f $X=6.725 $Y=1.765 $X2=0 $Y2=0
cc_326 N_A1_c_371_n N_VPWR_c_680_n 0.00445602f $X=7.175 $Y=1.765 $X2=0 $Y2=0
cc_327 N_A1_c_372_n N_VPWR_c_681_n 0.0044313f $X=7.625 $Y=1.765 $X2=0 $Y2=0
cc_328 N_A1_c_369_n N_VPWR_c_668_n 0.00912439f $X=6.26 $Y=1.765 $X2=0 $Y2=0
cc_329 N_A1_c_370_n N_VPWR_c_668_n 0.00857732f $X=6.725 $Y=1.765 $X2=0 $Y2=0
cc_330 N_A1_c_371_n N_VPWR_c_668_n 0.00857589f $X=7.175 $Y=1.765 $X2=0 $Y2=0
cc_331 N_A1_c_372_n N_VPWR_c_668_n 0.00853578f $X=7.625 $Y=1.765 $X2=0 $Y2=0
cc_332 N_A1_c_369_n N_A_954_368#_c_776_n 0.0129643f $X=6.26 $Y=1.765 $X2=0 $Y2=0
cc_333 N_A1_c_370_n N_A_954_368#_c_776_n 0.0118819f $X=6.725 $Y=1.765 $X2=0
+ $Y2=0
cc_334 N_A1_c_371_n N_A_954_368#_c_778_n 0.011796f $X=7.175 $Y=1.765 $X2=0 $Y2=0
cc_335 N_A1_c_372_n N_A_954_368#_c_778_n 0.011796f $X=7.625 $Y=1.765 $X2=0 $Y2=0
cc_336 N_A1_c_372_n N_A_954_368#_c_780_n 4.27055e-19 $X=7.625 $Y=1.765 $X2=0
+ $Y2=0
cc_337 N_A1_c_371_n N_A_954_368#_c_781_n 5.40974e-19 $X=7.175 $Y=1.765 $X2=0
+ $Y2=0
cc_338 N_A1_c_372_n N_A_954_368#_c_781_n 0.00574124f $X=7.625 $Y=1.765 $X2=0
+ $Y2=0
cc_339 N_A1_c_372_n N_A_954_368#_c_769_n 0.00328225f $X=7.625 $Y=1.765 $X2=0
+ $Y2=0
cc_340 N_A1_c_369_n N_A_954_368#_c_772_n 0.00145015f $X=6.26 $Y=1.765 $X2=0
+ $Y2=0
cc_341 N_A1_c_369_n N_A_954_368#_c_773_n 5.70119e-19 $X=6.26 $Y=1.765 $X2=0
+ $Y2=0
cc_342 N_A1_c_370_n N_A_954_368#_c_773_n 0.00744752f $X=6.725 $Y=1.765 $X2=0
+ $Y2=0
cc_343 N_A1_c_371_n N_A_954_368#_c_773_n 0.00730551f $X=7.175 $Y=1.765 $X2=0
+ $Y2=0
cc_344 N_A1_c_372_n N_A_954_368#_c_773_n 5.64076e-19 $X=7.625 $Y=1.765 $X2=0
+ $Y2=0
cc_345 N_A1_M1004_g N_A_841_74#_c_912_n 0.00654264f $X=6.355 $Y=0.74 $X2=0 $Y2=0
cc_346 N_A1_M1004_g N_A_841_74#_c_913_n 0.0115433f $X=6.355 $Y=0.74 $X2=0 $Y2=0
cc_347 N_A1_M1006_g N_A_841_74#_c_913_n 0.0135046f $X=6.855 $Y=0.74 $X2=0 $Y2=0
cc_348 N_A1_c_373_n N_A_841_74#_c_913_n 0.0510631f $X=7.47 $Y=1.515 $X2=0 $Y2=0
cc_349 N_A1_c_368_n N_A_841_74#_c_913_n 0.00418133f $X=7.625 $Y=1.542 $X2=0
+ $Y2=0
cc_350 N_A1_M1006_g N_A_841_74#_c_914_n 3.92313e-19 $X=6.855 $Y=0.74 $X2=0 $Y2=0
cc_351 N_A1_M1012_g N_A_841_74#_c_914_n 3.92313e-19 $X=7.285 $Y=0.74 $X2=0 $Y2=0
cc_352 N_A1_M1012_g N_A_841_74#_c_915_n 0.0131114f $X=7.285 $Y=0.74 $X2=0 $Y2=0
cc_353 N_A1_M1023_g N_A_841_74#_c_915_n 0.0173246f $X=7.715 $Y=0.74 $X2=0 $Y2=0
cc_354 N_A1_c_373_n N_A_841_74#_c_915_n 0.0362237f $X=7.47 $Y=1.515 $X2=0 $Y2=0
cc_355 N_A1_c_368_n N_A_841_74#_c_915_n 0.00238022f $X=7.625 $Y=1.542 $X2=0
+ $Y2=0
cc_356 N_A1_M1023_g N_A_841_74#_c_916_n 3.97481e-19 $X=7.715 $Y=0.74 $X2=0 $Y2=0
cc_357 N_A1_M1004_g N_A_841_74#_c_923_n 0.00524405f $X=6.355 $Y=0.74 $X2=0 $Y2=0
cc_358 N_A1_M1006_g N_A_841_74#_c_923_n 7.49986e-19 $X=6.855 $Y=0.74 $X2=0 $Y2=0
cc_359 N_A1_c_373_n N_A_841_74#_c_923_n 0.00162765f $X=7.47 $Y=1.515 $X2=0 $Y2=0
cc_360 N_A1_c_368_n N_A_841_74#_c_923_n 0.00545926f $X=7.625 $Y=1.542 $X2=0
+ $Y2=0
cc_361 N_A1_c_373_n N_A_841_74#_c_924_n 0.0146025f $X=7.47 $Y=1.515 $X2=0 $Y2=0
cc_362 N_A1_c_368_n N_A_841_74#_c_924_n 0.00254629f $X=7.625 $Y=1.542 $X2=0
+ $Y2=0
cc_363 N_A1_M1004_g N_VGND_c_1018_n 0.00560609f $X=6.355 $Y=0.74 $X2=0 $Y2=0
cc_364 N_A1_M1006_g N_VGND_c_1018_n 0.0102612f $X=6.855 $Y=0.74 $X2=0 $Y2=0
cc_365 N_A1_M1012_g N_VGND_c_1018_n 4.65668e-19 $X=7.285 $Y=0.74 $X2=0 $Y2=0
cc_366 N_A1_M1006_g N_VGND_c_1019_n 4.65668e-19 $X=6.855 $Y=0.74 $X2=0 $Y2=0
cc_367 N_A1_M1012_g N_VGND_c_1019_n 0.010248f $X=7.285 $Y=0.74 $X2=0 $Y2=0
cc_368 N_A1_M1023_g N_VGND_c_1019_n 0.0103688f $X=7.715 $Y=0.74 $X2=0 $Y2=0
cc_369 N_A1_M1004_g N_VGND_c_1022_n 0.00434272f $X=6.355 $Y=0.74 $X2=0 $Y2=0
cc_370 N_A1_M1006_g N_VGND_c_1023_n 0.00383152f $X=6.855 $Y=0.74 $X2=0 $Y2=0
cc_371 N_A1_M1012_g N_VGND_c_1023_n 0.00383152f $X=7.285 $Y=0.74 $X2=0 $Y2=0
cc_372 N_A1_M1023_g N_VGND_c_1024_n 0.00383152f $X=7.715 $Y=0.74 $X2=0 $Y2=0
cc_373 N_A1_M1004_g N_VGND_c_1027_n 0.0082143f $X=6.355 $Y=0.74 $X2=0 $Y2=0
cc_374 N_A1_M1006_g N_VGND_c_1027_n 0.0075754f $X=6.855 $Y=0.74 $X2=0 $Y2=0
cc_375 N_A1_M1012_g N_VGND_c_1027_n 0.0075754f $X=7.285 $Y=0.74 $X2=0 $Y2=0
cc_376 N_A1_M1023_g N_VGND_c_1027_n 0.00757637f $X=7.715 $Y=0.74 $X2=0 $Y2=0
cc_377 N_A2_c_457_n N_Y_c_542_n 0.0131451f $X=8.09 $Y=1.765 $X2=0 $Y2=0
cc_378 N_A2_c_455_n N_Y_c_542_n 0.026434f $X=9.405 $Y=1.515 $X2=0 $Y2=0
cc_379 N_A2_c_458_n N_Y_c_610_n 0.0122806f $X=8.575 $Y=1.765 $X2=0 $Y2=0
cc_380 N_A2_c_459_n N_Y_c_610_n 0.0154321f $X=9.075 $Y=1.765 $X2=0 $Y2=0
cc_381 N_A2_c_455_n N_Y_c_610_n 0.046015f $X=9.405 $Y=1.515 $X2=0 $Y2=0
cc_382 N_A2_c_456_n N_Y_c_610_n 0.00157789f $X=9.575 $Y=1.495 $X2=0 $Y2=0
cc_383 N_A2_c_458_n N_Y_c_614_n 0.00889139f $X=8.575 $Y=1.765 $X2=0 $Y2=0
cc_384 N_A2_c_459_n N_Y_c_614_n 4.54023e-19 $X=9.075 $Y=1.765 $X2=0 $Y2=0
cc_385 N_A2_c_455_n N_Y_c_614_n 0.0248048f $X=9.405 $Y=1.515 $X2=0 $Y2=0
cc_386 N_A2_c_456_n N_Y_c_614_n 0.00163693f $X=9.575 $Y=1.495 $X2=0 $Y2=0
cc_387 N_A2_c_460_n N_Y_c_618_n 0.0101384f $X=9.575 $Y=1.765 $X2=0 $Y2=0
cc_388 N_A2_c_455_n N_Y_c_618_n 0.0238641f $X=9.405 $Y=1.515 $X2=0 $Y2=0
cc_389 N_A2_c_456_n N_Y_c_618_n 0.00128027f $X=9.575 $Y=1.495 $X2=0 $Y2=0
cc_390 N_A2_c_457_n N_VPWR_c_681_n 0.00278271f $X=8.09 $Y=1.765 $X2=0 $Y2=0
cc_391 N_A2_c_458_n N_VPWR_c_681_n 0.00278271f $X=8.575 $Y=1.765 $X2=0 $Y2=0
cc_392 N_A2_c_459_n N_VPWR_c_681_n 0.00278257f $X=9.075 $Y=1.765 $X2=0 $Y2=0
cc_393 N_A2_c_460_n N_VPWR_c_681_n 0.00278271f $X=9.575 $Y=1.765 $X2=0 $Y2=0
cc_394 N_A2_c_457_n N_VPWR_c_668_n 0.00354367f $X=8.09 $Y=1.765 $X2=0 $Y2=0
cc_395 N_A2_c_458_n N_VPWR_c_668_n 0.00354611f $X=8.575 $Y=1.765 $X2=0 $Y2=0
cc_396 N_A2_c_459_n N_VPWR_c_668_n 0.00354744f $X=9.075 $Y=1.765 $X2=0 $Y2=0
cc_397 N_A2_c_460_n N_VPWR_c_668_n 0.00357778f $X=9.575 $Y=1.765 $X2=0 $Y2=0
cc_398 N_A2_c_457_n N_A_954_368#_c_768_n 0.0120121f $X=8.09 $Y=1.765 $X2=0 $Y2=0
cc_399 N_A2_c_458_n N_A_954_368#_c_768_n 0.0140488f $X=8.575 $Y=1.765 $X2=0
+ $Y2=0
cc_400 N_A2_c_457_n N_A_954_368#_c_769_n 0.00145169f $X=8.09 $Y=1.765 $X2=0
+ $Y2=0
cc_401 N_A2_c_459_n N_A_954_368#_c_792_n 0.00756708f $X=9.075 $Y=1.765 $X2=0
+ $Y2=0
cc_402 N_A2_c_460_n N_A_954_368#_c_792_n 8.49836e-19 $X=9.575 $Y=1.765 $X2=0
+ $Y2=0
cc_403 N_A2_c_459_n N_A_954_368#_c_770_n 0.0111147f $X=9.075 $Y=1.765 $X2=0
+ $Y2=0
cc_404 N_A2_c_460_n N_A_954_368#_c_770_n 0.0139779f $X=9.575 $Y=1.765 $X2=0
+ $Y2=0
cc_405 N_A2_c_460_n N_A_954_368#_c_771_n 0.010383f $X=9.575 $Y=1.765 $X2=0 $Y2=0
cc_406 N_A2_c_459_n N_A_954_368#_c_774_n 0.00193739f $X=9.075 $Y=1.765 $X2=0
+ $Y2=0
cc_407 N_A2_c_455_n N_A_841_74#_c_915_n 0.00320175f $X=9.405 $Y=1.515 $X2=0
+ $Y2=0
cc_408 N_A2_c_451_n N_A_841_74#_c_916_n 0.00930634f $X=8.145 $Y=1.225 $X2=0
+ $Y2=0
cc_409 N_A2_c_452_n N_A_841_74#_c_916_n 9.9103e-19 $X=8.645 $Y=1.225 $X2=0 $Y2=0
cc_410 N_A2_c_451_n N_A_841_74#_c_917_n 0.0115433f $X=8.145 $Y=1.225 $X2=0 $Y2=0
cc_411 N_A2_c_452_n N_A_841_74#_c_917_n 0.0136842f $X=8.645 $Y=1.225 $X2=0 $Y2=0
cc_412 N_A2_c_455_n N_A_841_74#_c_917_n 0.0510618f $X=9.405 $Y=1.515 $X2=0 $Y2=0
cc_413 N_A2_c_456_n N_A_841_74#_c_917_n 0.00472334f $X=9.575 $Y=1.495 $X2=0
+ $Y2=0
cc_414 N_A2_c_452_n N_A_841_74#_c_918_n 4.79304e-19 $X=8.645 $Y=1.225 $X2=0
+ $Y2=0
cc_415 N_A2_c_453_n N_A_841_74#_c_918_n 0.00351353f $X=9.155 $Y=1.225 $X2=0
+ $Y2=0
cc_416 N_A2_c_453_n N_A_841_74#_c_919_n 0.014803f $X=9.155 $Y=1.225 $X2=0 $Y2=0
cc_417 N_A2_c_454_n N_A_841_74#_c_919_n 0.0182356f $X=9.585 $Y=1.225 $X2=0 $Y2=0
cc_418 N_A2_c_455_n N_A_841_74#_c_919_n 0.035072f $X=9.405 $Y=1.515 $X2=0 $Y2=0
cc_419 N_A2_c_456_n N_A_841_74#_c_919_n 0.00308208f $X=9.575 $Y=1.495 $X2=0
+ $Y2=0
cc_420 N_A2_c_454_n N_A_841_74#_c_920_n 0.00159319f $X=9.585 $Y=1.225 $X2=0
+ $Y2=0
cc_421 N_A2_c_451_n N_A_841_74#_c_925_n 0.00155819f $X=8.145 $Y=1.225 $X2=0
+ $Y2=0
cc_422 N_A2_c_455_n N_A_841_74#_c_925_n 0.0220221f $X=9.405 $Y=1.515 $X2=0 $Y2=0
cc_423 N_A2_c_456_n N_A_841_74#_c_925_n 0.00219068f $X=9.575 $Y=1.495 $X2=0
+ $Y2=0
cc_424 N_A2_c_455_n N_A_841_74#_c_926_n 0.0214719f $X=9.405 $Y=1.515 $X2=0 $Y2=0
cc_425 N_A2_c_456_n N_A_841_74#_c_926_n 0.00520994f $X=9.575 $Y=1.495 $X2=0
+ $Y2=0
cc_426 N_A2_c_451_n N_VGND_c_1019_n 5.11853e-19 $X=8.145 $Y=1.225 $X2=0 $Y2=0
cc_427 N_A2_c_451_n N_VGND_c_1020_n 0.00413472f $X=8.145 $Y=1.225 $X2=0 $Y2=0
cc_428 N_A2_c_452_n N_VGND_c_1020_n 0.0105079f $X=8.645 $Y=1.225 $X2=0 $Y2=0
cc_429 N_A2_c_453_n N_VGND_c_1020_n 4.53659e-19 $X=9.155 $Y=1.225 $X2=0 $Y2=0
cc_430 N_A2_c_452_n N_VGND_c_1021_n 4.53659e-19 $X=8.645 $Y=1.225 $X2=0 $Y2=0
cc_431 N_A2_c_453_n N_VGND_c_1021_n 0.0104948f $X=9.155 $Y=1.225 $X2=0 $Y2=0
cc_432 N_A2_c_454_n N_VGND_c_1021_n 0.01328f $X=9.585 $Y=1.225 $X2=0 $Y2=0
cc_433 N_A2_c_451_n N_VGND_c_1024_n 0.00434272f $X=8.145 $Y=1.225 $X2=0 $Y2=0
cc_434 N_A2_c_452_n N_VGND_c_1025_n 0.00383152f $X=8.645 $Y=1.225 $X2=0 $Y2=0
cc_435 N_A2_c_453_n N_VGND_c_1025_n 0.00383152f $X=9.155 $Y=1.225 $X2=0 $Y2=0
cc_436 N_A2_c_454_n N_VGND_c_1026_n 0.00383152f $X=9.585 $Y=1.225 $X2=0 $Y2=0
cc_437 N_A2_c_451_n N_VGND_c_1027_n 0.00820816f $X=8.145 $Y=1.225 $X2=0 $Y2=0
cc_438 N_A2_c_452_n N_VGND_c_1027_n 0.00758285f $X=8.645 $Y=1.225 $X2=0 $Y2=0
cc_439 N_A2_c_453_n N_VGND_c_1027_n 0.00758285f $X=9.155 $Y=1.225 $X2=0 $Y2=0
cc_440 N_A2_c_454_n N_VGND_c_1027_n 0.00761198f $X=9.585 $Y=1.225 $X2=0 $Y2=0
cc_441 N_Y_c_551_n N_VPWR_M1020_s 0.00640259f $X=1.87 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_442 N_Y_c_538_n N_VPWR_M1003_s 0.00901236f $X=3.19 $Y=1.885 $X2=0 $Y2=0
cc_443 N_Y_c_581_n N_VPWR_M1002_s 0.00649593f $X=4.19 $Y=2.035 $X2=0 $Y2=0
cc_444 N_Y_c_542_n N_VPWR_M1007_s 0.00388867f $X=8.185 $Y=2.035 $X2=0 $Y2=0
cc_445 N_Y_c_542_n N_VPWR_M1015_s 0.00359847f $X=8.185 $Y=2.035 $X2=0 $Y2=0
cc_446 N_Y_c_551_n N_VPWR_c_669_n 0.0232685f $X=1.87 $Y=2.035 $X2=0 $Y2=0
cc_447 N_Y_c_537_n N_VPWR_c_669_n 0.0266809f $X=2.035 $Y=2.815 $X2=0 $Y2=0
cc_448 N_Y_c_543_n N_VPWR_c_669_n 0.0297756f $X=1.2 $Y=2.465 $X2=0 $Y2=0
cc_449 N_Y_c_537_n N_VPWR_c_670_n 0.0323945f $X=2.035 $Y=2.815 $X2=0 $Y2=0
cc_450 N_Y_c_538_n N_VPWR_c_670_n 0.0493032f $X=3.19 $Y=1.885 $X2=0 $Y2=0
cc_451 N_Y_c_540_n N_VPWR_c_670_n 0.0323945f $X=3.355 $Y=2.815 $X2=0 $Y2=0
cc_452 N_Y_c_540_n N_VPWR_c_671_n 0.0266809f $X=3.355 $Y=2.815 $X2=0 $Y2=0
cc_453 N_Y_c_581_n N_VPWR_c_671_n 0.0232685f $X=4.19 $Y=2.035 $X2=0 $Y2=0
cc_454 N_Y_c_541_n N_VPWR_c_671_n 0.0266809f $X=4.355 $Y=2.815 $X2=0 $Y2=0
cc_455 N_Y_c_543_n N_VPWR_c_674_n 0.0481755f $X=1.2 $Y=2.465 $X2=0 $Y2=0
cc_456 N_Y_c_540_n N_VPWR_c_676_n 0.014552f $X=3.355 $Y=2.815 $X2=0 $Y2=0
cc_457 N_Y_c_537_n N_VPWR_c_678_n 0.014552f $X=2.035 $Y=2.815 $X2=0 $Y2=0
cc_458 N_Y_c_541_n N_VPWR_c_679_n 0.0145938f $X=4.355 $Y=2.815 $X2=0 $Y2=0
cc_459 N_Y_c_537_n N_VPWR_c_668_n 0.0119791f $X=2.035 $Y=2.815 $X2=0 $Y2=0
cc_460 N_Y_c_540_n N_VPWR_c_668_n 0.0119791f $X=3.355 $Y=2.815 $X2=0 $Y2=0
cc_461 N_Y_c_541_n N_VPWR_c_668_n 0.0120466f $X=4.355 $Y=2.815 $X2=0 $Y2=0
cc_462 N_Y_c_543_n N_VPWR_c_668_n 0.0399762f $X=1.2 $Y=2.465 $X2=0 $Y2=0
cc_463 N_Y_c_542_n N_A_954_368#_M1007_d 0.0383262f $X=8.185 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_464 N_Y_c_542_n N_A_954_368#_M1010_d 0.00359365f $X=8.185 $Y=2.035 $X2=0
+ $Y2=0
cc_465 N_Y_c_542_n N_A_954_368#_M1025_d 0.00483883f $X=8.185 $Y=2.035 $X2=0
+ $Y2=0
cc_466 N_Y_c_610_n N_A_954_368#_M1017_s 0.00455969f $X=9.185 $Y=2.035 $X2=0
+ $Y2=0
cc_467 N_Y_c_541_n N_A_954_368#_c_767_n 0.0492197f $X=4.355 $Y=2.815 $X2=0 $Y2=0
cc_468 N_Y_c_542_n N_A_954_368#_c_767_n 0.145594f $X=8.185 $Y=2.035 $X2=0 $Y2=0
cc_469 N_Y_c_542_n N_A_954_368#_c_778_n 0.0317427f $X=8.185 $Y=2.035 $X2=0 $Y2=0
cc_470 N_Y_c_542_n N_A_954_368#_c_780_n 0.0174536f $X=8.185 $Y=2.035 $X2=0 $Y2=0
cc_471 N_Y_M1016_d N_A_954_368#_c_768_n 0.00234927f $X=8.165 $Y=1.84 $X2=0 $Y2=0
cc_472 N_Y_c_614_n N_A_954_368#_c_768_n 0.0177813f $X=8.35 $Y=2.115 $X2=0 $Y2=0
cc_473 N_Y_c_610_n N_A_954_368#_c_792_n 0.0202249f $X=9.185 $Y=2.035 $X2=0 $Y2=0
cc_474 N_Y_M1019_d N_A_954_368#_c_770_n 0.00250873f $X=9.15 $Y=1.84 $X2=0 $Y2=0
cc_475 N_Y_c_618_n N_A_954_368#_c_770_n 0.018923f $X=9.35 $Y=2.115 $X2=0 $Y2=0
cc_476 N_Y_c_618_n N_A_954_368#_c_771_n 0.0533059f $X=9.35 $Y=2.115 $X2=0 $Y2=0
cc_477 N_Y_c_542_n N_A_954_368#_c_773_n 0.0173542f $X=8.185 $Y=2.035 $X2=0 $Y2=0
cc_478 N_Y_c_534_n N_A_27_74#_M1013_d 0.00177442f $X=1.565 $Y=0.95 $X2=0 $Y2=0
cc_479 N_Y_M1011_s N_A_27_74#_c_835_n 0.00238148f $X=0.57 $Y=0.37 $X2=0 $Y2=0
cc_480 N_Y_M1030_s N_A_27_74#_c_835_n 0.00169014f $X=1.5 $Y=0.37 $X2=0 $Y2=0
cc_481 N_Y_c_534_n N_A_27_74#_c_835_n 0.0526342f $X=1.565 $Y=0.95 $X2=0 $Y2=0
cc_482 N_Y_c_554_n N_A_27_74#_c_835_n 0.0145945f $X=1.685 $Y=1.13 $X2=0 $Y2=0
cc_483 N_Y_c_554_n N_A_27_74#_c_837_n 0.0135821f $X=1.685 $Y=1.13 $X2=0 $Y2=0
cc_484 N_Y_c_536_n N_A_27_74#_c_837_n 0.00685376f $X=2.2 $Y=1.885 $X2=0 $Y2=0
cc_485 N_Y_c_538_n N_A_27_74#_c_838_n 2.54876e-19 $X=3.19 $Y=1.885 $X2=0 $Y2=0
cc_486 N_Y_c_536_n N_A_27_74#_c_838_n 0.00142628f $X=2.2 $Y=1.885 $X2=0 $Y2=0
cc_487 N_Y_c_534_n N_A_27_74#_c_839_n 0.0143359f $X=1.565 $Y=0.95 $X2=0 $Y2=0
cc_488 N_VPWR_c_679_n N_A_954_368#_c_767_n 0.0629185f $X=6.335 $Y=3.33 $X2=0
+ $Y2=0
cc_489 N_VPWR_c_668_n N_A_954_368#_c_767_n 0.0522437f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_490 N_VPWR_M1007_s N_A_954_368#_c_776_n 0.00434779f $X=6.335 $Y=1.84 $X2=0
+ $Y2=0
cc_491 N_VPWR_c_672_n N_A_954_368#_c_776_n 0.0156208f $X=6.5 $Y=2.805 $X2=0
+ $Y2=0
cc_492 N_VPWR_M1015_s N_A_954_368#_c_778_n 0.00428955f $X=7.25 $Y=1.84 $X2=0
+ $Y2=0
cc_493 N_VPWR_c_673_n N_A_954_368#_c_778_n 0.0136682f $X=7.4 $Y=2.805 $X2=0
+ $Y2=0
cc_494 N_VPWR_c_673_n N_A_954_368#_c_781_n 0.0178797f $X=7.4 $Y=2.805 $X2=0
+ $Y2=0
cc_495 N_VPWR_c_681_n N_A_954_368#_c_768_n 0.0422316f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_496 N_VPWR_c_668_n N_A_954_368#_c_768_n 0.0238179f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_497 N_VPWR_c_673_n N_A_954_368#_c_769_n 0.0119328f $X=7.4 $Y=2.805 $X2=0
+ $Y2=0
cc_498 N_VPWR_c_681_n N_A_954_368#_c_769_n 0.0236039f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_499 N_VPWR_c_668_n N_A_954_368#_c_769_n 0.012761f $X=9.84 $Y=3.33 $X2=0 $Y2=0
cc_500 N_VPWR_c_681_n N_A_954_368#_c_770_n 0.0621295f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_501 N_VPWR_c_668_n N_A_954_368#_c_770_n 0.0347335f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_502 N_VPWR_c_672_n N_A_954_368#_c_772_n 0.0147794f $X=6.5 $Y=2.805 $X2=0
+ $Y2=0
cc_503 N_VPWR_c_672_n N_A_954_368#_c_773_n 0.0234974f $X=6.5 $Y=2.805 $X2=0
+ $Y2=0
cc_504 N_VPWR_c_673_n N_A_954_368#_c_773_n 0.0228252f $X=7.4 $Y=2.805 $X2=0
+ $Y2=0
cc_505 N_VPWR_c_680_n N_A_954_368#_c_773_n 0.0145674f $X=7.315 $Y=3.33 $X2=0
+ $Y2=0
cc_506 N_VPWR_c_668_n N_A_954_368#_c_773_n 0.0119851f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_507 N_VPWR_c_681_n N_A_954_368#_c_774_n 0.0236039f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_508 N_VPWR_c_668_n N_A_954_368#_c_774_n 0.012761f $X=9.84 $Y=3.33 $X2=0 $Y2=0
cc_509 N_A_954_368#_c_771_n N_A_841_74#_c_919_n 0.00916738f $X=9.8 $Y=1.985
+ $X2=0 $Y2=0
cc_510 N_A_27_74#_c_838_n N_A_472_74#_M1000_s 0.00177476f $X=3.79 $Y=0.95
+ $X2=-0.19 $Y2=-0.245
cc_511 N_A_27_74#_c_838_n N_A_472_74#_M1026_s 0.00177476f $X=3.79 $Y=0.95 $X2=0
+ $Y2=0
cc_512 N_A_27_74#_M1008_d N_A_472_74#_c_883_n 0.00169036f $X=2.79 $Y=0.37 $X2=0
+ $Y2=0
cc_513 N_A_27_74#_M1028_d N_A_472_74#_c_883_n 0.00406362f $X=3.65 $Y=0.37 $X2=0
+ $Y2=0
cc_514 N_A_27_74#_c_836_n N_A_472_74#_c_883_n 0.0108703f $X=2.07 $Y=0.6 $X2=0
+ $Y2=0
cc_515 N_A_27_74#_c_838_n N_A_472_74#_c_883_n 0.0915637f $X=3.79 $Y=0.95 $X2=0
+ $Y2=0
cc_516 N_A_27_74#_c_838_n N_A_841_74#_c_921_n 0.0235569f $X=3.79 $Y=0.95 $X2=0
+ $Y2=0
cc_517 N_A_27_74#_c_835_n N_VGND_c_1022_n 0.0622328f $X=1.985 $Y=0.475 $X2=0
+ $Y2=0
cc_518 N_A_27_74#_c_836_n N_VGND_c_1022_n 0.00758556f $X=2.07 $Y=0.6 $X2=0 $Y2=0
cc_519 N_A_27_74#_c_839_n N_VGND_c_1022_n 0.0146502f $X=0.28 $Y=0.515 $X2=0
+ $Y2=0
cc_520 N_A_27_74#_c_835_n N_VGND_c_1027_n 0.052295f $X=1.985 $Y=0.475 $X2=0
+ $Y2=0
cc_521 N_A_27_74#_c_836_n N_VGND_c_1027_n 0.00627867f $X=2.07 $Y=0.6 $X2=0 $Y2=0
cc_522 N_A_27_74#_c_838_n N_VGND_c_1027_n 0.00825751f $X=3.79 $Y=0.95 $X2=0
+ $Y2=0
cc_523 N_A_27_74#_c_839_n N_VGND_c_1027_n 0.0120674f $X=0.28 $Y=0.515 $X2=0
+ $Y2=0
cc_524 N_A_472_74#_c_883_n N_A_841_74#_M1009_s 0.00406362f $X=5.475 $Y=0.515
+ $X2=-0.19 $Y2=-0.245
cc_525 N_A_472_74#_c_883_n N_A_841_74#_M1014_s 0.00195031f $X=5.475 $Y=0.515
+ $X2=0 $Y2=0
cc_526 N_A_472_74#_M1027_d N_A_841_74#_c_910_n 0.00178215f $X=5.5 $Y=0.37 $X2=0
+ $Y2=0
cc_527 N_A_472_74#_c_882_n N_A_841_74#_c_910_n 0.0165836f $X=5.64 $Y=0.515 $X2=0
+ $Y2=0
cc_528 N_A_472_74#_c_882_n N_A_841_74#_c_912_n 0.0144195f $X=5.64 $Y=0.515 $X2=0
+ $Y2=0
cc_529 N_A_472_74#_c_883_n N_A_841_74#_c_921_n 0.0209443f $X=5.475 $Y=0.515
+ $X2=0 $Y2=0
cc_530 N_A_472_74#_M1009_d N_A_841_74#_c_922_n 0.00191886f $X=4.64 $Y=0.37 $X2=0
+ $Y2=0
cc_531 N_A_472_74#_c_883_n N_A_841_74#_c_922_n 0.0460916f $X=5.475 $Y=0.515
+ $X2=0 $Y2=0
cc_532 N_A_472_74#_c_883_n N_VGND_c_1022_n 0.142867f $X=5.475 $Y=0.515 $X2=0
+ $Y2=0
cc_533 N_A_472_74#_c_883_n N_VGND_c_1027_n 0.120151f $X=5.475 $Y=0.515 $X2=0
+ $Y2=0
cc_534 N_A_841_74#_c_913_n N_VGND_M1004_s 0.00263002f $X=6.985 $Y=1.095
+ $X2=-0.19 $Y2=-0.245
cc_535 N_A_841_74#_c_915_n N_VGND_M1012_s 0.00184993f $X=7.845 $Y=1.095 $X2=0
+ $Y2=0
cc_536 N_A_841_74#_c_917_n N_VGND_M1001_s 0.00263002f $X=8.775 $Y=1.095 $X2=0
+ $Y2=0
cc_537 N_A_841_74#_c_919_n N_VGND_M1021_s 0.00184993f $X=9.715 $Y=1.095 $X2=0
+ $Y2=0
cc_538 N_A_841_74#_c_912_n N_VGND_c_1018_n 0.018426f $X=6.14 $Y=0.515 $X2=0
+ $Y2=0
cc_539 N_A_841_74#_c_913_n N_VGND_c_1018_n 0.0193036f $X=6.985 $Y=1.095 $X2=0
+ $Y2=0
cc_540 N_A_841_74#_c_914_n N_VGND_c_1018_n 0.017532f $X=7.07 $Y=0.515 $X2=0
+ $Y2=0
cc_541 N_A_841_74#_c_914_n N_VGND_c_1019_n 0.017532f $X=7.07 $Y=0.515 $X2=0
+ $Y2=0
cc_542 N_A_841_74#_c_915_n N_VGND_c_1019_n 0.0156953f $X=7.845 $Y=1.095 $X2=0
+ $Y2=0
cc_543 N_A_841_74#_c_916_n N_VGND_c_1019_n 0.0175734f $X=7.93 $Y=0.515 $X2=0
+ $Y2=0
cc_544 N_A_841_74#_c_916_n N_VGND_c_1020_n 0.0176914f $X=7.93 $Y=0.515 $X2=0
+ $Y2=0
cc_545 N_A_841_74#_c_917_n N_VGND_c_1020_n 0.0193036f $X=8.775 $Y=1.095 $X2=0
+ $Y2=0
cc_546 N_A_841_74#_c_918_n N_VGND_c_1020_n 0.0175734f $X=8.86 $Y=0.515 $X2=0
+ $Y2=0
cc_547 N_A_841_74#_c_918_n N_VGND_c_1021_n 0.0175734f $X=8.86 $Y=0.515 $X2=0
+ $Y2=0
cc_548 N_A_841_74#_c_919_n N_VGND_c_1021_n 0.0156953f $X=9.715 $Y=1.095 $X2=0
+ $Y2=0
cc_549 N_A_841_74#_c_920_n N_VGND_c_1021_n 0.0175734f $X=9.8 $Y=0.515 $X2=0
+ $Y2=0
cc_550 N_A_841_74#_c_912_n N_VGND_c_1022_n 0.0145639f $X=6.14 $Y=0.515 $X2=0
+ $Y2=0
cc_551 N_A_841_74#_c_914_n N_VGND_c_1023_n 0.00749631f $X=7.07 $Y=0.515 $X2=0
+ $Y2=0
cc_552 N_A_841_74#_c_916_n N_VGND_c_1024_n 0.0109942f $X=7.93 $Y=0.515 $X2=0
+ $Y2=0
cc_553 N_A_841_74#_c_918_n N_VGND_c_1025_n 0.011066f $X=8.86 $Y=0.515 $X2=0
+ $Y2=0
cc_554 N_A_841_74#_c_920_n N_VGND_c_1026_n 0.011066f $X=9.8 $Y=0.515 $X2=0 $Y2=0
cc_555 N_A_841_74#_c_912_n N_VGND_c_1027_n 0.0119984f $X=6.14 $Y=0.515 $X2=0
+ $Y2=0
cc_556 N_A_841_74#_c_914_n N_VGND_c_1027_n 0.0062048f $X=7.07 $Y=0.515 $X2=0
+ $Y2=0
cc_557 N_A_841_74#_c_916_n N_VGND_c_1027_n 0.00904371f $X=7.93 $Y=0.515 $X2=0
+ $Y2=0
cc_558 N_A_841_74#_c_918_n N_VGND_c_1027_n 0.00915947f $X=8.86 $Y=0.515 $X2=0
+ $Y2=0
cc_559 N_A_841_74#_c_920_n N_VGND_c_1027_n 0.00915947f $X=9.8 $Y=0.515 $X2=0
+ $Y2=0
cc_560 N_A_841_74#_c_922_n N_VGND_c_1027_n 0.00736333f $X=5.045 $Y=1.015 $X2=0
+ $Y2=0
