* File: sky130_fd_sc_hs__nor3_2.pex.spice
* Created: Tue Sep  1 20:11:32 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HS__NOR3_2%C 1 3 4 6 7 9 10 15
c40 15 0 8.80415e-20 $X=0.81 $Y=1.385
c41 7 0 3.88207e-20 $X=1.005 $Y=1.765
r42 15 17 20.4326 $w=4.6e-07 $l=1.95e-07 $layer=POLY_cond $X=0.81 $Y=1.492
+ $X2=1.005 $Y2=1.492
r43 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.81
+ $Y=1.385 $X2=0.81 $Y2=1.385
r44 10 16 2.80324 $w=3.68e-07 $l=9e-08 $layer=LI1_cond $X=0.79 $Y=1.295 $X2=0.79
+ $Y2=1.385
r45 7 17 29.3143 $w=1.5e-07 $l=2.73e-07 $layer=POLY_cond $X=1.005 $Y=1.765
+ $X2=1.005 $Y2=1.492
r46 7 9 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.005 $Y=1.765
+ $X2=1.005 $Y2=2.4
r47 4 15 31.9587 $w=4.6e-07 $l=4.19869e-07 $layer=POLY_cond $X=0.505 $Y=1.765
+ $X2=0.81 $Y2=1.492
r48 4 6 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.505 $Y=1.765
+ $X2=0.505 $Y2=2.4
r49 1 4 1.04783 $w=4.6e-07 $l=5.49977e-07 $layer=POLY_cond $X=0.495 $Y=1.22
+ $X2=0.505 $Y2=1.765
r50 1 3 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=0.495 $Y=1.22 $X2=0.495
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HS__NOR3_2%B 1 3 4 6 7 9 10 13 18
c63 13 0 1.08023e-19 $X=1.47 $Y=1.385
c64 1 0 1.72885e-19 $X=1.455 $Y=1.765
r65 23 28 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=3.09 $Y=1.385 $X2=3.09
+ $Y2=1.465
r66 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.09
+ $Y=1.385 $X2=3.09 $Y2=1.385
r67 18 23 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=3.09 $Y=1.295 $X2=3.09
+ $Y2=1.385
r68 13 16 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=1.47 $Y=1.385 $X2=1.47
+ $Y2=1.465
r69 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.47
+ $Y=1.385 $X2=1.47 $Y2=1.385
r70 11 16 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.635 $Y=1.465
+ $X2=1.47 $Y2=1.465
r71 10 28 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.925 $Y=1.465
+ $X2=3.09 $Y2=1.465
r72 10 11 84.1604 $w=1.68e-07 $l=1.29e-06 $layer=LI1_cond $X=2.925 $Y=1.465
+ $X2=1.635 $Y2=1.465
r73 7 22 72.5138 $w=3.05e-07 $l=4.50888e-07 $layer=POLY_cond $X=2.855 $Y=1.765
+ $X2=3.01 $Y2=1.385
r74 7 9 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.855 $Y=1.765
+ $X2=2.855 $Y2=2.4
r75 4 14 38.9026 $w=2.7e-07 $l=1.92678e-07 $layer=POLY_cond $X=1.53 $Y=1.22
+ $X2=1.47 $Y2=1.385
r76 4 6 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.53 $Y=1.22 $X2=1.53
+ $Y2=0.74
r77 1 14 77.2841 $w=2.7e-07 $l=3.87427e-07 $layer=POLY_cond $X=1.455 $Y=1.765
+ $X2=1.47 $Y2=1.385
r78 1 3 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.455 $Y=1.765
+ $X2=1.455 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_HS__NOR3_2%A 2 3 5 6 8 9 12 13 15 17 18 20 23 24 27
c62 2 0 1.08023e-19 $X=1.935 $Y=1.675
r63 27 28 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.815
+ $Y=0.475 $X2=2.815 $Y2=0.475
r64 24 28 5.44483 $w=6.68e-07 $l=3.05e-07 $layer=LI1_cond $X=3.12 $Y=0.645
+ $X2=2.815 $Y2=0.645
r65 22 27 35.3689 $w=4.45e-07 $l=2.83e-07 $layer=POLY_cond $X=2.757 $Y=0.758
+ $X2=2.757 $Y2=0.475
r66 22 23 53.9265 $w=4.45e-07 $l=2.22e-07 $layer=POLY_cond $X=2.757 $Y=0.758
+ $X2=2.757 $Y2=0.98
r67 17 20 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.61 $Y=1.185
+ $X2=2.61 $Y2=1.26
r68 17 23 105.117 $w=1.5e-07 $l=2.05e-07 $layer=POLY_cond $X=2.61 $Y=1.185
+ $X2=2.61 $Y2=0.98
r69 13 15 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.405 $Y=1.765
+ $X2=2.405 $Y2=2.4
r70 12 13 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=2.405 $Y=1.675
+ $X2=2.405 $Y2=1.765
r71 11 20 105.117 $w=1.5e-07 $l=2.05e-07 $layer=POLY_cond $X=2.405 $Y=1.26
+ $X2=2.61 $Y2=1.26
r72 11 12 132.161 $w=1.8e-07 $l=3.4e-07 $layer=POLY_cond $X=2.405 $Y=1.335
+ $X2=2.405 $Y2=1.675
r73 10 18 6.66866 $w=1.5e-07 $l=1.3e-07 $layer=POLY_cond $X=2.105 $Y=1.26
+ $X2=1.975 $Y2=1.26
r74 9 11 46.1489 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=2.315 $Y=1.26 $X2=2.405
+ $Y2=1.26
r75 9 10 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=2.315 $Y=1.26
+ $X2=2.105 $Y2=1.26
r76 6 18 18.8402 $w=1.65e-07 $l=9.87421e-08 $layer=POLY_cond $X=2.03 $Y=1.185
+ $X2=1.975 $Y2=1.26
r77 6 8 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=2.03 $Y=1.185
+ $X2=2.03 $Y2=0.74
r78 3 5 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.935 $Y=1.765
+ $X2=1.935 $Y2=2.4
r79 2 3 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=1.935 $Y=1.675 $X2=1.935
+ $Y2=1.765
r80 1 18 18.8402 $w=1.65e-07 $l=9.28709e-08 $layer=POLY_cond $X=1.935 $Y=1.335
+ $X2=1.975 $Y2=1.26
r81 1 2 132.161 $w=1.8e-07 $l=3.4e-07 $layer=POLY_cond $X=1.935 $Y=1.335
+ $X2=1.935 $Y2=1.675
.ends

.subckt PM_SKY130_FD_SC_HS__NOR3_2%A_27_368# 1 2 3 12 16 17 21 24 25 28
c48 25 0 7.12326e-20 $X=1.315 $Y=1.805
c49 1 0 1.80713e-19 $X=0.135 $Y=1.84
r50 28 30 34.1617 $w=2.78e-07 $l=8.3e-07 $layer=LI1_cond $X=3.105 $Y=1.985
+ $X2=3.105 $Y2=2.815
r51 26 28 3.91007 $w=2.78e-07 $l=9.5e-08 $layer=LI1_cond $X=3.105 $Y=1.89
+ $X2=3.105 $Y2=1.985
r52 24 26 7.36005 $w=1.7e-07 $l=1.77482e-07 $layer=LI1_cond $X=2.965 $Y=1.805
+ $X2=3.105 $Y2=1.89
r53 24 25 107.647 $w=1.68e-07 $l=1.65e-06 $layer=LI1_cond $X=2.965 $Y=1.805
+ $X2=1.315 $Y2=1.805
r54 21 23 54.1497 $w=1.68e-07 $l=8.3e-07 $layer=LI1_cond $X=1.23 $Y=1.985
+ $X2=1.23 $Y2=2.815
r55 19 23 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=1.23 $Y=2.905 $X2=1.23
+ $Y2=2.815
r56 18 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.23 $Y=1.89
+ $X2=1.315 $Y2=1.805
r57 18 21 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=1.23 $Y=1.89
+ $X2=1.23 $Y2=1.985
r58 16 19 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.145 $Y=2.99
+ $X2=1.23 $Y2=2.905
r59 16 17 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=1.145 $Y=2.99
+ $X2=0.445 $Y2=2.99
r60 12 15 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=0.28 $Y=2.145
+ $X2=0.28 $Y2=2.825
r61 10 17 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.28 $Y=2.905
+ $X2=0.445 $Y2=2.99
r62 10 15 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=0.28 $Y=2.905 $X2=0.28
+ $Y2=2.825
r63 3 30 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=2.93
+ $Y=1.84 $X2=3.08 $Y2=2.815
r64 3 28 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=2.93
+ $Y=1.84 $X2=3.08 $Y2=1.985
r65 2 23 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=1.08
+ $Y=1.84 $X2=1.23 $Y2=2.815
r66 2 21 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=1.08
+ $Y=1.84 $X2=1.23 $Y2=1.985
r67 1 15 400 $w=1.7e-07 $l=1.05501e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.825
r68 1 12 400 $w=1.7e-07 $l=3.70473e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.145
.ends

.subckt PM_SKY130_FD_SC_HS__NOR3_2%Y 1 2 3 10 12 16 22 24 25 26 27 42 48
c45 25 0 8.80415e-20 $X=0.24 $Y=0.925
c46 10 0 2.82366e-19 $X=0.615 $Y=1.805
r47 42 48 2.64102 $w=2.38e-07 $l=5.5e-08 $layer=LI1_cond $X=0.235 $Y=1.72
+ $X2=0.235 $Y2=1.665
r48 27 42 2.93484 $w=2.4e-07 $l=8.5e-08 $layer=LI1_cond $X=0.235 $Y=1.805
+ $X2=0.235 $Y2=1.72
r49 27 48 0.720277 $w=2.38e-07 $l=1.5e-08 $layer=LI1_cond $X=0.235 $Y=1.65
+ $X2=0.235 $Y2=1.665
r50 26 27 17.0466 $w=2.38e-07 $l=3.55e-07 $layer=LI1_cond $X=0.235 $Y=1.295
+ $X2=0.235 $Y2=1.65
r51 25 26 9.97569 $w=4.08e-07 $l=2.85e-07 $layer=LI1_cond $X=0.235 $Y=1.01
+ $X2=0.235 $Y2=1.295
r52 24 25 9.1582 $w=4.98e-07 $l=3.25e-07 $layer=LI1_cond $X=0.28 $Y=0.515
+ $X2=0.28 $Y2=0.84
r53 20 22 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=1.815 $Y=0.84
+ $X2=1.815 $Y2=0.515
r54 16 18 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=0.78 $Y=1.97
+ $X2=0.78 $Y2=2.65
r55 14 16 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=0.78 $Y=1.89 $X2=0.78
+ $Y2=1.97
r56 13 25 3.25423 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.445 $Y=0.925
+ $X2=0.28 $Y2=0.925
r57 12 20 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.65 $Y=0.925
+ $X2=1.815 $Y2=0.84
r58 12 13 78.615 $w=1.68e-07 $l=1.205e-06 $layer=LI1_cond $X=1.65 $Y=0.925
+ $X2=0.445 $Y2=0.925
r59 11 27 4.1433 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=0.355 $Y=1.805
+ $X2=0.235 $Y2=1.805
r60 10 14 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.615 $Y=1.805
+ $X2=0.78 $Y2=1.89
r61 10 11 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=0.615 $Y=1.805
+ $X2=0.355 $Y2=1.805
r62 3 18 400 $w=1.7e-07 $l=9.04489e-07 $layer=licon1_PDIFF $count=1 $X=0.58
+ $Y=1.84 $X2=0.78 $Y2=2.65
r63 3 16 400 $w=1.7e-07 $l=2.56905e-07 $layer=licon1_PDIFF $count=1 $X=0.58
+ $Y=1.84 $X2=0.78 $Y2=1.97
r64 2 22 91 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=2 $X=1.605
+ $Y=0.37 $X2=1.815 $Y2=0.515
r65 1 24 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__NOR3_2%A_306_368# 1 2 7 9 11 13 15
c27 9 0 3.88207e-20 $X=1.68 $Y=2.485
r28 13 20 2.78046 $w=2.8e-07 $l=8.5e-08 $layer=LI1_cond $X=2.655 $Y=2.23
+ $X2=2.655 $Y2=2.145
r29 13 15 10.4955 $w=2.78e-07 $l=2.55e-07 $layer=LI1_cond $X=2.655 $Y=2.23
+ $X2=2.655 $Y2=2.485
r30 12 18 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.845 $Y=2.145
+ $X2=1.68 $Y2=2.145
r31 11 20 4.57959 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=2.515 $Y=2.145
+ $X2=2.655 $Y2=2.145
r32 11 12 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.515 $Y=2.145
+ $X2=1.845 $Y2=2.145
r33 7 18 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.68 $Y=2.23 $X2=1.68
+ $Y2=2.145
r34 7 9 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=1.68 $Y=2.23 $X2=1.68
+ $Y2=2.485
r35 2 20 600 $w=1.7e-07 $l=3.72525e-07 $layer=licon1_PDIFF $count=1 $X=2.48
+ $Y=1.84 $X2=2.63 $Y2=2.145
r36 2 15 300 $w=1.7e-07 $l=7.16083e-07 $layer=licon1_PDIFF $count=2 $X=2.48
+ $Y=1.84 $X2=2.63 $Y2=2.485
r37 1 18 600 $w=1.7e-07 $l=3.72525e-07 $layer=licon1_PDIFF $count=1 $X=1.53
+ $Y=1.84 $X2=1.68 $Y2=2.145
r38 1 9 300 $w=1.7e-07 $l=7.16083e-07 $layer=licon1_PDIFF $count=2 $X=1.53
+ $Y=1.84 $X2=1.68 $Y2=2.485
.ends

.subckt PM_SKY130_FD_SC_HS__NOR3_2%VPWR 1 6 8 10 20 21 24
r36 24 25 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r37 21 25 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=2.16 $Y2=3.33
r38 20 21 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r39 18 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.345 $Y=3.33
+ $X2=2.18 $Y2=3.33
r40 18 20 50.5615 $w=1.68e-07 $l=7.75e-07 $layer=LI1_cond $X=2.345 $Y=3.33
+ $X2=3.12 $Y2=3.33
r41 12 16 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=0.24 $Y=3.33
+ $X2=1.68 $Y2=3.33
r42 12 13 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r43 10 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.015 $Y=3.33
+ $X2=2.18 $Y2=3.33
r44 10 16 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=2.015 $Y=3.33
+ $X2=1.68 $Y2=3.33
r45 8 25 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r46 8 13 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=0.24 $Y2=3.33
r47 8 16 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r48 4 24 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.18 $Y=3.245 $X2=2.18
+ $Y2=3.33
r49 4 6 26.5411 $w=3.28e-07 $l=7.6e-07 $layer=LI1_cond $X=2.18 $Y=3.245 $X2=2.18
+ $Y2=2.485
r50 1 6 300 $w=1.7e-07 $l=7.25034e-07 $layer=licon1_PDIFF $count=2 $X=2.01
+ $Y=1.84 $X2=2.18 $Y2=2.485
.ends

.subckt PM_SKY130_FD_SC_HS__NOR3_2%VGND 1 2 7 11 13 22 23 28 34 36
r35 36 37 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r36 33 34 11.0283 $w=7.33e-07 $l=1.65e-07 $layer=LI1_cond $X=1.315 $Y=0.282
+ $X2=1.48 $Y2=0.282
r37 30 33 1.87142 $w=7.33e-07 $l=1.15e-07 $layer=LI1_cond $X=1.2 $Y=0.282
+ $X2=1.315 $Y2=0.282
r38 30 31 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r39 27 31 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r40 26 30 7.81112 $w=7.33e-07 $l=4.8e-07 $layer=LI1_cond $X=0.72 $Y=0.282
+ $X2=1.2 $Y2=0.282
r41 26 28 10.0519 $w=7.33e-07 $l=1.05e-07 $layer=LI1_cond $X=0.72 $Y=0.282
+ $X2=0.615 $Y2=0.282
r42 26 27 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r43 23 37 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=2.16
+ $Y2=0
r44 22 23 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r45 20 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.48 $Y=0 $X2=2.315
+ $Y2=0
r46 20 22 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=2.48 $Y=0 $X2=3.12
+ $Y2=0
r47 18 27 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r48 17 28 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=0.24 $Y=0 $X2=0.615
+ $Y2=0
r49 17 18 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r50 13 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r51 13 31 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r52 9 36 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.315 $Y=0.085
+ $X2=2.315 $Y2=0
r53 9 11 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=2.315 $Y=0.085
+ $X2=2.315 $Y2=0.515
r54 7 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.15 $Y=0 $X2=2.315
+ $Y2=0
r55 7 34 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.15 $Y=0 $X2=1.48
+ $Y2=0
r56 2 11 91 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=2 $X=2.105
+ $Y=0.37 $X2=2.315 $Y2=0.515
r57 1 33 91 $w=1.7e-07 $l=8.14279e-07 $layer=licon1_NDIFF $count=2 $X=0.57
+ $Y=0.37 $X2=1.315 $Y2=0.515
.ends

