* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hs__nand2_2 A B VGND VNB VPB VPWR Y
M1000 Y A a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=2.442e+11p pd=2.14e+06u as=6.438e+11p ps=6.18e+06u
M1001 VPWR B Y VPB pshort w=1.12e+06u l=150000u
+  ad=1.008e+12p pd=8.52e+06u as=6.72e+11p ps=5.68e+06u
M1002 a_27_74# A Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1003 Y B VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_27_74# B VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.442e+11p ps=2.14e+06u
M1005 VGND B a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 Y A VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VPWR A Y VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
