* NGSPICE file created from sky130_fd_sc_hs__a32oi_1.ext - technology: sky130A

.subckt sky130_fd_sc_hs__a32oi_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
M1000 Y B1 a_119_74# VNB nlowvt w=740000u l=150000u
+  ad=6.068e+11p pd=3.12e+06u as=1.776e+11p ps=1.96e+06u
M1001 VGND A3 a_469_74# VNB nlowvt w=740000u l=150000u
+  ad=4.403e+11p pd=4.15e+06u as=3.108e+11p ps=2.32e+06u
M1002 a_119_74# B2 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1003 a_27_368# B1 Y VPB pshort w=1.12e+06u l=150000u
+  ad=1.1816e+12p pd=8.83e+06u as=3.92e+11p ps=2.94e+06u
M1004 Y B2 a_27_368# VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_27_368# A2 VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=1.0472e+12p ps=6.35e+06u
M1006 a_391_74# A1 Y VNB nlowvt w=740000u l=150000u
+  ad=1.776e+11p pd=1.96e+06u as=0p ps=0u
M1007 VPWR A3 a_27_368# VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VPWR A1 a_27_368# VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_469_74# A2 a_391_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

