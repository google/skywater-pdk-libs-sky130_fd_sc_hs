* File: sky130_fd_sc_hs__fah_2.pxi.spice
* Created: Thu Aug 27 20:46:17 2020
* 
x_PM_SKY130_FD_SC_HS__FAH_2%A_81_260# N_A_81_260#_M1017_s N_A_81_260#_M1015_s
+ N_A_81_260#_c_258_n N_A_81_260#_M1002_g N_A_81_260#_M1034_g
+ N_A_81_260#_c_260_n N_A_81_260#_c_261_n N_A_81_260#_c_262_n
+ N_A_81_260#_c_263_n N_A_81_260#_c_264_n PM_SKY130_FD_SC_HS__FAH_2%A_81_260#
x_PM_SKY130_FD_SC_HS__FAH_2%A N_A_c_316_n N_A_c_322_n N_A_M1015_g N_A_c_317_n
+ N_A_M1017_g N_A_c_318_n N_A_c_324_n N_A_M1030_g N_A_c_319_n N_A_M1005_g A
+ N_A_c_325_n N_A_c_320_n PM_SKY130_FD_SC_HS__FAH_2%A
x_PM_SKY130_FD_SC_HS__FAH_2%B N_B_M1006_g N_B_c_382_n N_B_M1010_g N_B_M1007_g
+ N_B_c_398_n N_B_M1024_g N_B_c_399_n N_B_M1000_g N_B_c_383_n N_B_c_384_n
+ N_B_M1033_g N_B_c_419_p N_B_c_464_p N_B_c_422_p N_B_c_386_n N_B_c_387_n
+ N_B_c_442_p N_B_c_447_p N_B_c_388_n N_B_c_448_p N_B_c_389_n N_B_c_390_n
+ N_B_c_391_n N_B_c_392_n N_B_c_393_n N_B_c_532_p N_B_c_571_p N_B_c_394_n B B
+ N_B_c_396_n PM_SKY130_FD_SC_HS__FAH_2%B
x_PM_SKY130_FD_SC_HS__FAH_2%A_481_379# N_A_481_379#_M1033_d N_A_481_379#_M1000_d
+ N_A_481_379#_c_602_n N_A_481_379#_M1003_g N_A_481_379#_c_603_n
+ N_A_481_379#_c_604_n N_A_481_379#_c_591_n N_A_481_379#_c_592_n
+ N_A_481_379#_M1008_g N_A_481_379#_c_593_n N_A_481_379#_c_594_n
+ N_A_481_379#_c_595_n N_A_481_379#_c_607_n N_A_481_379#_M1016_g
+ N_A_481_379#_c_608_n N_A_481_379#_c_609_n N_A_481_379#_M1025_g
+ N_A_481_379#_c_596_n N_A_481_379#_c_597_n N_A_481_379#_c_610_n
+ N_A_481_379#_c_598_n N_A_481_379#_c_599_n N_A_481_379#_c_600_n
+ N_A_481_379#_c_666_n N_A_481_379#_c_601_n N_A_481_379#_c_613_n
+ PM_SKY130_FD_SC_HS__FAH_2%A_481_379#
x_PM_SKY130_FD_SC_HS__FAH_2%A_514_424# N_A_514_424#_M1006_d N_A_514_424#_M1003_d
+ N_A_514_424#_c_758_n N_A_514_424#_M1012_g N_A_514_424#_M1020_g
+ N_A_514_424#_c_760_n N_A_514_424#_M1031_g N_A_514_424#_M1027_g
+ N_A_514_424#_c_796_n N_A_514_424#_c_762_n N_A_514_424#_c_802_n
+ N_A_514_424#_c_846_p N_A_514_424#_c_775_n N_A_514_424#_c_776_n
+ N_A_514_424#_c_806_n N_A_514_424#_c_777_n N_A_514_424#_c_809_n
+ N_A_514_424#_c_778_n N_A_514_424#_c_779_n N_A_514_424#_c_763_n
+ N_A_514_424#_c_764_n N_A_514_424#_c_781_n N_A_514_424#_c_782_n
+ N_A_514_424#_c_863_p N_A_514_424#_c_864_p N_A_514_424#_c_765_n
+ N_A_514_424#_c_766_n N_A_514_424#_c_841_n N_A_514_424#_c_783_n
+ N_A_514_424#_c_767_n N_A_514_424#_c_921_p N_A_514_424#_c_785_n
+ N_A_514_424#_c_768_n N_A_514_424#_c_769_n N_A_514_424#_c_770_n
+ N_A_514_424#_c_771_n PM_SKY130_FD_SC_HS__FAH_2%A_514_424#
x_PM_SKY130_FD_SC_HS__FAH_2%A_849_424# N_A_849_424#_M1007_d N_A_849_424#_M1016_d
+ N_A_849_424#_c_1004_n N_A_849_424#_M1019_g N_A_849_424#_c_1026_n
+ N_A_849_424#_c_1027_n N_A_849_424#_c_1028_n N_A_849_424#_M1004_g
+ N_A_849_424#_c_1029_n N_A_849_424#_c_1005_n N_A_849_424#_c_1006_n
+ N_A_849_424#_c_1007_n N_A_849_424#_M1009_g N_A_849_424#_c_1009_n
+ N_A_849_424#_c_1010_n N_A_849_424#_c_1032_n N_A_849_424#_M1013_g
+ N_A_849_424#_c_1011_n N_A_849_424#_c_1034_n N_A_849_424#_c_1012_n
+ N_A_849_424#_c_1035_n N_A_849_424#_c_1013_n N_A_849_424#_c_1037_n
+ N_A_849_424#_c_1014_n N_A_849_424#_c_1015_n N_A_849_424#_c_1016_n
+ N_A_849_424#_c_1017_n N_A_849_424#_c_1018_n N_A_849_424#_c_1198_p
+ N_A_849_424#_c_1019_n N_A_849_424#_c_1020_n N_A_849_424#_c_1021_n
+ N_A_849_424#_c_1022_n N_A_849_424#_c_1023_n N_A_849_424#_c_1039_n
+ N_A_849_424#_c_1024_n N_A_849_424#_c_1025_n
+ PM_SKY130_FD_SC_HS__FAH_2%A_849_424#
x_PM_SKY130_FD_SC_HS__FAH_2%A_1689_424# N_A_1689_424#_M1020_d
+ N_A_1689_424#_M1021_d N_A_1689_424#_M1004_d N_A_1689_424#_M1001_d
+ N_A_1689_424#_M1011_g N_A_1689_424#_c_1214_n N_A_1689_424#_M1032_g
+ N_A_1689_424#_c_1234_n N_A_1689_424#_c_1215_n N_A_1689_424#_c_1216_n
+ N_A_1689_424#_c_1217_n N_A_1689_424#_c_1293_p N_A_1689_424#_c_1223_n
+ N_A_1689_424#_c_1218_n N_A_1689_424#_c_1242_n N_A_1689_424#_c_1219_n
+ N_A_1689_424#_c_1220_n PM_SKY130_FD_SC_HS__FAH_2%A_1689_424#
x_PM_SKY130_FD_SC_HS__FAH_2%CI N_CI_M1021_g N_CI_c_1329_n N_CI_c_1330_n
+ N_CI_M1001_g N_CI_c_1331_n N_CI_c_1332_n CI PM_SKY130_FD_SC_HS__FAH_2%CI
x_PM_SKY130_FD_SC_HS__FAH_2%A_1451_424# N_A_1451_424#_M1019_d
+ N_A_1451_424#_M1012_d N_A_1451_424#_c_1381_n N_A_1451_424#_M1023_g
+ N_A_1451_424#_c_1372_n N_A_1451_424#_M1014_g N_A_1451_424#_c_1373_n
+ N_A_1451_424#_M1035_g N_A_1451_424#_c_1382_n N_A_1451_424#_M1026_g
+ N_A_1451_424#_c_1374_n N_A_1451_424#_c_1375_n N_A_1451_424#_c_1376_n
+ N_A_1451_424#_c_1377_n N_A_1451_424#_c_1378_n N_A_1451_424#_c_1379_n
+ N_A_1451_424#_c_1442_n N_A_1451_424#_c_1380_n
+ PM_SKY130_FD_SC_HS__FAH_2%A_1451_424#
x_PM_SKY130_FD_SC_HS__FAH_2%A_1895_424# N_A_1895_424#_M1009_d
+ N_A_1895_424#_M1031_d N_A_1895_424#_c_1511_n N_A_1895_424#_M1018_g
+ N_A_1895_424#_M1022_g N_A_1895_424#_c_1512_n N_A_1895_424#_M1028_g
+ N_A_1895_424#_M1029_g N_A_1895_424#_c_1524_n N_A_1895_424#_c_1513_n
+ N_A_1895_424#_c_1537_n N_A_1895_424#_c_1514_n N_A_1895_424#_c_1506_n
+ N_A_1895_424#_c_1507_n N_A_1895_424#_c_1508_n N_A_1895_424#_c_1517_n
+ N_A_1895_424#_c_1518_n N_A_1895_424#_c_1509_n N_A_1895_424#_c_1510_n
+ PM_SKY130_FD_SC_HS__FAH_2%A_1895_424#
x_PM_SKY130_FD_SC_HS__FAH_2%VPWR N_VPWR_M1002_s N_VPWR_M1015_d N_VPWR_M1000_s
+ N_VPWR_M1032_d N_VPWR_M1023_s N_VPWR_M1026_s N_VPWR_M1028_d N_VPWR_c_1628_n
+ N_VPWR_c_1629_n N_VPWR_c_1630_n N_VPWR_c_1631_n N_VPWR_c_1632_n
+ N_VPWR_c_1633_n N_VPWR_c_1634_n N_VPWR_c_1635_n VPWR N_VPWR_c_1636_n
+ N_VPWR_c_1637_n N_VPWR_c_1638_n N_VPWR_c_1639_n N_VPWR_c_1640_n
+ N_VPWR_c_1641_n N_VPWR_c_1642_n N_VPWR_c_1643_n N_VPWR_c_1644_n
+ N_VPWR_c_1645_n N_VPWR_c_1646_n N_VPWR_c_1627_n PM_SKY130_FD_SC_HS__FAH_2%VPWR
x_PM_SKY130_FD_SC_HS__FAH_2%A_114_368# N_A_114_368#_M1034_d N_A_114_368#_M1008_d
+ N_A_114_368#_M1002_d N_A_114_368#_M1010_d N_A_114_368#_c_1757_n
+ N_A_114_368#_c_1766_n N_A_114_368#_c_1758_n N_A_114_368#_c_1798_n
+ N_A_114_368#_c_1759_n N_A_114_368#_c_1760_n N_A_114_368#_c_1768_n
+ N_A_114_368#_c_1761_n N_A_114_368#_c_1762_n N_A_114_368#_c_1763_n
+ N_A_114_368#_c_1764_n PM_SKY130_FD_SC_HS__FAH_2%A_114_368#
x_PM_SKY130_FD_SC_HS__FAH_2%A_413_392# N_A_413_392#_M1005_d N_A_413_392#_M1025_d
+ N_A_413_392#_M1030_d N_A_413_392#_M1024_d N_A_413_392#_c_1864_n
+ N_A_413_392#_c_1871_n N_A_413_392#_c_1858_n N_A_413_392#_c_1865_n
+ N_A_413_392#_c_1866_n N_A_413_392#_c_1859_n N_A_413_392#_c_1860_n
+ N_A_413_392#_c_1867_n N_A_413_392#_c_1861_n N_A_413_392#_c_1862_n
+ N_A_413_392#_c_1863_n PM_SKY130_FD_SC_HS__FAH_2%A_413_392#
x_PM_SKY130_FD_SC_HS__FAH_2%A_2052_424# N_A_2052_424#_M1027_d
+ N_A_2052_424#_M1013_d N_A_2052_424#_c_1949_n N_A_2052_424#_c_1951_n
+ N_A_2052_424#_c_1946_n N_A_2052_424#_c_1947_n
+ PM_SKY130_FD_SC_HS__FAH_2%A_2052_424#
x_PM_SKY130_FD_SC_HS__FAH_2%COUT N_COUT_M1014_d N_COUT_M1023_d N_COUT_c_1985_n
+ COUT COUT COUT PM_SKY130_FD_SC_HS__FAH_2%COUT
x_PM_SKY130_FD_SC_HS__FAH_2%SUM N_SUM_M1022_s N_SUM_M1018_s N_SUM_c_2007_n
+ N_SUM_c_2010_n N_SUM_c_2011_n N_SUM_c_2008_n SUM PM_SKY130_FD_SC_HS__FAH_2%SUM
x_PM_SKY130_FD_SC_HS__FAH_2%VGND N_VGND_M1034_s N_VGND_M1017_d N_VGND_M1033_s
+ N_VGND_M1011_d N_VGND_M1014_s N_VGND_M1035_s N_VGND_M1029_d N_VGND_c_2043_n
+ N_VGND_c_2044_n N_VGND_c_2045_n N_VGND_c_2046_n N_VGND_c_2047_n
+ N_VGND_c_2048_n N_VGND_c_2049_n N_VGND_c_2050_n N_VGND_c_2051_n
+ N_VGND_c_2052_n N_VGND_c_2053_n N_VGND_c_2054_n N_VGND_c_2055_n VGND
+ N_VGND_c_2056_n N_VGND_c_2057_n N_VGND_c_2058_n N_VGND_c_2059_n
+ N_VGND_c_2060_n N_VGND_c_2061_n N_VGND_c_2062_n N_VGND_c_2063_n
+ PM_SKY130_FD_SC_HS__FAH_2%VGND
cc_1 VNB N_A_81_260#_c_258_n 0.0257256f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.765
cc_2 VNB N_A_81_260#_M1034_g 0.0304613f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=0.74
cc_3 VNB N_A_81_260#_c_260_n 9.71834e-19 $X=-0.19 $Y=-0.245 $X2=1.255 $Y2=2.105
cc_4 VNB N_A_81_260#_c_261_n 0.00383363f $X=-0.19 $Y=-0.245 $X2=1.31 $Y2=1.3
cc_5 VNB N_A_81_260#_c_262_n 0.0551545f $X=-0.19 $Y=-0.245 $X2=0.985 $Y2=1.465
cc_6 VNB N_A_81_260#_c_263_n 0.00341862f $X=-0.19 $Y=-0.245 $X2=1.31 $Y2=1.465
cc_7 VNB N_A_81_260#_c_264_n 0.014731f $X=-0.19 $Y=-0.245 $X2=1.54 $Y2=0.675
cc_8 VNB N_A_c_316_n 0.00208222f $X=-0.19 $Y=-0.245 $X2=1.12 $Y2=1.96
cc_9 VNB N_A_c_317_n 0.0212268f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_c_318_n 0.00228474f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.3
cc_11 VNB N_A_c_319_n 0.0158174f $X=-0.19 $Y=-0.245 $X2=0.532 $Y2=1.465
cc_12 VNB N_A_c_320_n 0.0675748f $X=-0.19 $Y=-0.245 $X2=0.985 $Y2=1.465
cc_13 VNB N_B_M1006_g 0.0215123f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_B_c_382_n 0.00584614f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_B_c_383_n 0.0295739f $X=-0.19 $Y=-0.245 $X2=1.215 $Y2=2.105
cc_16 VNB N_B_c_384_n 0.113621f $X=-0.19 $Y=-0.245 $X2=1.255 $Y2=2.105
cc_17 VNB N_B_M1033_g 0.0210016f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_B_c_386_n 0.00258973f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_B_c_387_n 0.0344524f $X=-0.19 $Y=-0.245 $X2=1.465 $Y2=1.12
cc_20 VNB N_B_c_388_n 0.00496422f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_B_c_389_n 0.00171296f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_B_c_390_n 0.0242761f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_B_c_391_n 8.6513e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_B_c_392_n 6.14813e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_B_c_393_n 0.00448366f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_B_c_394_n 0.0103395f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB B 8.20392e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_B_c_396_n 0.022256f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_481_379#_c_591_n 0.0141765f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_481_379#_c_592_n 0.0203544f $X=-0.19 $Y=-0.245 $X2=0.532 $Y2=1.465
cc_31 VNB N_A_481_379#_c_593_n 0.0388121f $X=-0.19 $Y=-0.245 $X2=1.215 $Y2=2.105
cc_32 VNB N_A_481_379#_c_594_n 0.0257093f $X=-0.19 $Y=-0.245 $X2=1.255 $Y2=2.105
cc_33 VNB N_A_481_379#_c_595_n 0.0164677f $X=-0.19 $Y=-0.245 $X2=1.255 $Y2=2.815
cc_34 VNB N_A_481_379#_c_596_n 0.0176523f $X=-0.19 $Y=-0.245 $X2=1.465 $Y2=1.12
cc_35 VNB N_A_481_379#_c_597_n 0.0198122f $X=-0.19 $Y=-0.245 $X2=0.985 $Y2=1.465
cc_36 VNB N_A_481_379#_c_598_n 0.00367338f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_481_379#_c_599_n 0.00946755f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_481_379#_c_600_n 0.00202061f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_481_379#_c_601_n 0.0196462f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_514_424#_c_758_n 0.0131556f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.765
cc_41 VNB N_A_514_424#_M1020_g 0.0292724f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=0.74
cc_42 VNB N_A_514_424#_c_760_n 0.0060955f $X=-0.19 $Y=-0.245 $X2=0.532 $Y2=1.465
cc_43 VNB N_A_514_424#_M1027_g 0.0302152f $X=-0.19 $Y=-0.245 $X2=1.215 $Y2=2.815
cc_44 VNB N_A_514_424#_c_762_n 0.00595314f $X=-0.19 $Y=-0.245 $X2=0.985
+ $Y2=1.465
cc_45 VNB N_A_514_424#_c_763_n 0.00239721f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_A_514_424#_c_764_n 0.0340035f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_514_424#_c_765_n 0.00246662f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_514_424#_c_766_n 5.08129e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A_514_424#_c_767_n 0.00320499f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_A_514_424#_c_768_n 0.00208667f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_A_514_424#_c_769_n 0.00500752f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_A_514_424#_c_770_n 0.00211508f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_A_514_424#_c_771_n 0.0243623f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_A_849_424#_c_1004_n 0.065048f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.765
cc_55 VNB N_A_849_424#_c_1005_n 0.0147053f $X=-0.19 $Y=-0.245 $X2=1.255
+ $Y2=2.105
cc_56 VNB N_A_849_424#_c_1006_n 0.0189045f $X=-0.19 $Y=-0.245 $X2=1.215
+ $Y2=2.815
cc_57 VNB N_A_849_424#_c_1007_n 0.00847401f $X=-0.19 $Y=-0.245 $X2=1.255
+ $Y2=2.815
cc_58 VNB N_A_849_424#_M1009_g 0.0263607f $X=-0.19 $Y=-0.245 $X2=1.31 $Y2=1.3
cc_59 VNB N_A_849_424#_c_1009_n 0.0297475f $X=-0.19 $Y=-0.245 $X2=0.985
+ $Y2=1.465
cc_60 VNB N_A_849_424#_c_1010_n 0.0157829f $X=-0.19 $Y=-0.245 $X2=1.215
+ $Y2=1.465
cc_61 VNB N_A_849_424#_c_1011_n 0.0183592f $X=-0.19 $Y=-0.245 $X2=0.985
+ $Y2=1.465
cc_62 VNB N_A_849_424#_c_1012_n 0.00487969f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_A_849_424#_c_1013_n 0.00435657f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_A_849_424#_c_1014_n 0.00393961f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_A_849_424#_c_1015_n 0.00329413f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_A_849_424#_c_1016_n 0.00409229f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_A_849_424#_c_1017_n 0.00717338f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_A_849_424#_c_1018_n 0.00596127f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_A_849_424#_c_1019_n 0.0104708f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_A_849_424#_c_1020_n 0.00246632f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_A_849_424#_c_1021_n 0.00570775f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_A_849_424#_c_1022_n 0.00359524f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_A_849_424#_c_1023_n 0.00469939f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_A_849_424#_c_1024_n 0.00658776f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_A_849_424#_c_1025_n 0.001369f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_A_1689_424#_M1011_g 0.0362251f $X=-0.19 $Y=-0.245 $X2=0.66 $Y2=1.465
cc_77 VNB N_A_1689_424#_c_1214_n 0.0237505f $X=-0.19 $Y=-0.245 $X2=1.215
+ $Y2=2.105
cc_78 VNB N_A_1689_424#_c_1215_n 0.0168712f $X=-0.19 $Y=-0.245 $X2=1.215
+ $Y2=1.465
cc_79 VNB N_A_1689_424#_c_1216_n 0.00586035f $X=-0.19 $Y=-0.245 $X2=1.31
+ $Y2=1.465
cc_80 VNB N_A_1689_424#_c_1217_n 0.00867081f $X=-0.19 $Y=-0.245 $X2=0.985
+ $Y2=1.465
cc_81 VNB N_A_1689_424#_c_1218_n 0.00690842f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_82 VNB N_A_1689_424#_c_1219_n 0.00578144f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_83 VNB N_A_1689_424#_c_1220_n 0.0197558f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_84 VNB N_CI_c_1329_n 0.0127735f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_85 VNB N_CI_c_1330_n 0.0187948f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_86 VNB N_CI_c_1331_n 0.0178059f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.4
cc_87 VNB N_CI_c_1332_n 0.0134725f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.3
cc_88 VNB CI 0.00489304f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=0.74
cc_89 VNB N_A_1451_424#_c_1372_n 0.0176257f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.3
cc_90 VNB N_A_1451_424#_c_1373_n 0.0171438f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_91 VNB N_A_1451_424#_c_1374_n 0.0420428f $X=-0.19 $Y=-0.245 $X2=1.215
+ $Y2=2.815
cc_92 VNB N_A_1451_424#_c_1375_n 0.0474858f $X=-0.19 $Y=-0.245 $X2=1.31 $Y2=1.12
cc_93 VNB N_A_1451_424#_c_1376_n 0.00755117f $X=-0.19 $Y=-0.245 $X2=0.985
+ $Y2=1.465
cc_94 VNB N_A_1451_424#_c_1377_n 0.0118556f $X=-0.19 $Y=-0.245 $X2=0.985
+ $Y2=1.465
cc_95 VNB N_A_1451_424#_c_1378_n 0.0151776f $X=-0.19 $Y=-0.245 $X2=1.465
+ $Y2=0.675
cc_96 VNB N_A_1451_424#_c_1379_n 0.00523245f $X=-0.19 $Y=-0.245 $X2=1.54
+ $Y2=0.675
cc_97 VNB N_A_1451_424#_c_1380_n 0.0180007f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_98 VNB N_A_1895_424#_M1022_g 0.0223658f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=0.74
cc_99 VNB N_A_1895_424#_M1029_g 0.0239451f $X=-0.19 $Y=-0.245 $X2=1.215
+ $Y2=2.815
cc_100 VNB N_A_1895_424#_c_1506_n 3.59478e-19 $X=-0.19 $Y=-0.245 $X2=1.54
+ $Y2=0.675
cc_101 VNB N_A_1895_424#_c_1507_n 0.00338173f $X=-0.19 $Y=-0.245 $X2=1.465
+ $Y2=1.12
cc_102 VNB N_A_1895_424#_c_1508_n 0.00326134f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_103 VNB N_A_1895_424#_c_1509_n 0.00320706f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_104 VNB N_A_1895_424#_c_1510_n 0.0618652f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_105 VNB N_VPWR_c_1627_n 0.601534f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_106 VNB N_A_114_368#_c_1757_n 0.00741748f $X=-0.19 $Y=-0.245 $X2=0.532
+ $Y2=1.465
cc_107 VNB N_A_114_368#_c_1758_n 0.0138891f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_108 VNB N_A_114_368#_c_1759_n 0.00340344f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_109 VNB N_A_114_368#_c_1760_n 0.00232803f $X=-0.19 $Y=-0.245 $X2=1.215
+ $Y2=1.465
cc_110 VNB N_A_114_368#_c_1761_n 0.0321667f $X=-0.19 $Y=-0.245 $X2=1.465
+ $Y2=1.12
cc_111 VNB N_A_114_368#_c_1762_n 0.0150676f $X=-0.19 $Y=-0.245 $X2=0.985
+ $Y2=1.465
cc_112 VNB N_A_114_368#_c_1763_n 0.0040707f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_113 VNB N_A_114_368#_c_1764_n 0.0232151f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_114 VNB N_A_413_392#_c_1858_n 9.33229e-19 $X=-0.19 $Y=-0.245 $X2=1.31
+ $Y2=1.12
cc_115 VNB N_A_413_392#_c_1859_n 0.0539803f $X=-0.19 $Y=-0.245 $X2=0.985
+ $Y2=1.465
cc_116 VNB N_A_413_392#_c_1860_n 0.0031605f $X=-0.19 $Y=-0.245 $X2=0.985
+ $Y2=1.465
cc_117 VNB N_A_413_392#_c_1861_n 0.00312637f $X=-0.19 $Y=-0.245 $X2=1.465
+ $Y2=0.675
cc_118 VNB N_A_413_392#_c_1862_n 0.00202458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_119 VNB N_A_413_392#_c_1863_n 0.0156939f $X=-0.19 $Y=-0.245 $X2=1.465
+ $Y2=1.12
cc_120 VNB N_A_2052_424#_c_1946_n 0.00355309f $X=-0.19 $Y=-0.245 $X2=1.215
+ $Y2=1.63
cc_121 VNB N_A_2052_424#_c_1947_n 0.0065492f $X=-0.19 $Y=-0.245 $X2=1.215
+ $Y2=2.815
cc_122 VNB N_COUT_c_1985_n 0.00303633f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.4
cc_123 VNB N_SUM_c_2007_n 0.00222347f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.4
cc_124 VNB N_SUM_c_2008_n 2.20818e-19 $X=-0.19 $Y=-0.245 $X2=1.215 $Y2=2.815
cc_125 VNB SUM 0.0421128f $X=-0.19 $Y=-0.245 $X2=1.255 $Y2=2.815
cc_126 VNB N_VGND_c_2043_n 0.0144549f $X=-0.19 $Y=-0.245 $X2=1.31 $Y2=1.12
cc_127 VNB N_VGND_c_2044_n 0.0273179f $X=-0.19 $Y=-0.245 $X2=0.985 $Y2=1.465
cc_128 VNB N_VGND_c_2045_n 0.0136114f $X=-0.19 $Y=-0.245 $X2=1.215 $Y2=1.465
cc_129 VNB N_VGND_c_2046_n 0.0176636f $X=-0.19 $Y=-0.245 $X2=1.54 $Y2=0.675
cc_130 VNB N_VGND_c_2047_n 0.0064467f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_131 VNB N_VGND_c_2048_n 0.0123668f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_132 VNB N_VGND_c_2049_n 0.012847f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_133 VNB N_VGND_c_2050_n 0.012003f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_134 VNB N_VGND_c_2051_n 0.0197038f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_135 VNB N_VGND_c_2052_n 0.0376514f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_136 VNB N_VGND_c_2053_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_137 VNB N_VGND_c_2054_n 0.106621f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_138 VNB N_VGND_c_2055_n 0.00477918f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_139 VNB N_VGND_c_2056_n 0.0998192f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_140 VNB N_VGND_c_2057_n 0.0198633f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_141 VNB N_VGND_c_2058_n 0.0172524f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_142 VNB N_VGND_c_2059_n 0.0171166f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_143 VNB N_VGND_c_2060_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_144 VNB N_VGND_c_2061_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_145 VNB N_VGND_c_2062_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_146 VNB N_VGND_c_2063_n 0.797122f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_147 VPB N_A_81_260#_c_258_n 0.0298194f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.765
cc_148 VPB N_A_81_260#_c_260_n 0.0179389f $X=-0.19 $Y=1.66 $X2=1.255 $Y2=2.105
cc_149 VPB N_A_c_316_n 0.00756744f $X=-0.19 $Y=1.66 $X2=1.12 $Y2=1.96
cc_150 VPB N_A_c_322_n 0.0255202f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_151 VPB N_A_c_318_n 0.00771209f $X=-0.19 $Y=1.66 $X2=0.585 $Y2=1.3
cc_152 VPB N_A_c_324_n 0.0229293f $X=-0.19 $Y=1.66 $X2=0.585 $Y2=0.74
cc_153 VPB N_A_c_325_n 0.00400445f $X=-0.19 $Y=1.66 $X2=0.985 $Y2=1.465
cc_154 VPB N_B_c_382_n 0.0493245f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_155 VPB N_B_c_398_n 0.0215473f $X=-0.19 $Y=1.66 $X2=0.585 $Y2=0.74
cc_156 VPB N_B_c_399_n 0.0180968f $X=-0.19 $Y=1.66 $X2=0.532 $Y2=1.465
cc_157 VPB N_B_c_384_n 0.0564647f $X=-0.19 $Y=1.66 $X2=1.255 $Y2=2.105
cc_158 VPB N_B_c_390_n 0.00521694f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_159 VPB N_B_c_392_n 0.00155578f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_160 VPB B 0.0035102f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_161 VPB N_A_481_379#_c_602_n 0.0184369f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.765
cc_162 VPB N_A_481_379#_c_603_n 0.0405885f $X=-0.19 $Y=1.66 $X2=0.585 $Y2=1.3
cc_163 VPB N_A_481_379#_c_604_n 0.0125754f $X=-0.19 $Y=1.66 $X2=0.585 $Y2=0.74
cc_164 VPB N_A_481_379#_c_591_n 0.0123522f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_165 VPB N_A_481_379#_c_595_n 0.0104813f $X=-0.19 $Y=1.66 $X2=1.255 $Y2=2.815
cc_166 VPB N_A_481_379#_c_607_n 0.018531f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_167 VPB N_A_481_379#_c_608_n 0.0666828f $X=-0.19 $Y=1.66 $X2=0.985 $Y2=1.465
cc_168 VPB N_A_481_379#_c_609_n 0.0149522f $X=-0.19 $Y=1.66 $X2=0.985 $Y2=1.465
cc_169 VPB N_A_481_379#_c_610_n 0.00975145f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_170 VPB N_A_481_379#_c_598_n 9.85156e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_171 VPB N_A_481_379#_c_601_n 0.0133658f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_172 VPB N_A_481_379#_c_613_n 0.00258507f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_173 VPB N_A_514_424#_c_758_n 0.0572427f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.765
cc_174 VPB N_A_514_424#_c_760_n 0.0494484f $X=-0.19 $Y=1.66 $X2=0.532 $Y2=1.465
cc_175 VPB N_A_514_424#_c_762_n 0.00618152f $X=-0.19 $Y=1.66 $X2=0.985 $Y2=1.465
cc_176 VPB N_A_514_424#_c_775_n 0.0114774f $X=-0.19 $Y=1.66 $X2=1.465 $Y2=0.675
cc_177 VPB N_A_514_424#_c_776_n 0.0017718f $X=-0.19 $Y=1.66 $X2=1.54 $Y2=0.675
cc_178 VPB N_A_514_424#_c_777_n 0.00546222f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_179 VPB N_A_514_424#_c_778_n 0.00958146f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_180 VPB N_A_514_424#_c_779_n 9.46358e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_181 VPB N_A_514_424#_c_763_n 0.00409879f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_182 VPB N_A_514_424#_c_781_n 0.00828456f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_183 VPB N_A_514_424#_c_782_n 0.00107913f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_184 VPB N_A_514_424#_c_783_n 0.00489604f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_185 VPB N_A_514_424#_c_767_n 0.00443824f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_186 VPB N_A_514_424#_c_785_n 0.00230964f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_187 VPB N_A_514_424#_c_768_n 0.00445955f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_188 VPB N_A_514_424#_c_770_n 0.00148142f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_189 VPB N_A_514_424#_c_771_n 0.0114979f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_190 VPB N_A_849_424#_c_1026_n 0.014381f $X=-0.19 $Y=1.66 $X2=0.585 $Y2=1.3
cc_191 VPB N_A_849_424#_c_1027_n 0.0160174f $X=-0.19 $Y=1.66 $X2=0.585 $Y2=0.74
cc_192 VPB N_A_849_424#_c_1028_n 0.0198383f $X=-0.19 $Y=1.66 $X2=0.585 $Y2=0.74
cc_193 VPB N_A_849_424#_c_1029_n 0.0438325f $X=-0.19 $Y=1.66 $X2=0.66 $Y2=1.465
cc_194 VPB N_A_849_424#_c_1005_n 0.00814155f $X=-0.19 $Y=1.66 $X2=1.255
+ $Y2=2.105
cc_195 VPB N_A_849_424#_c_1010_n 0.0129659f $X=-0.19 $Y=1.66 $X2=1.215 $Y2=1.465
cc_196 VPB N_A_849_424#_c_1032_n 0.0198066f $X=-0.19 $Y=1.66 $X2=1.31 $Y2=1.465
cc_197 VPB N_A_849_424#_c_1011_n 0.00918238f $X=-0.19 $Y=1.66 $X2=0.985
+ $Y2=1.465
cc_198 VPB N_A_849_424#_c_1034_n 0.0182908f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_199 VPB N_A_849_424#_c_1035_n 0.0282406f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_200 VPB N_A_849_424#_c_1013_n 0.0062303f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_201 VPB N_A_849_424#_c_1037_n 0.00228158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_202 VPB N_A_849_424#_c_1022_n 0.00456093f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_203 VPB N_A_849_424#_c_1039_n 0.00480806f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_204 VPB N_A_1689_424#_c_1214_n 0.0473341f $X=-0.19 $Y=1.66 $X2=1.215
+ $Y2=2.105
cc_205 VPB N_A_1689_424#_c_1217_n 0.0024247f $X=-0.19 $Y=1.66 $X2=0.985
+ $Y2=1.465
cc_206 VPB N_A_1689_424#_c_1223_n 0.0143153f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_207 VPB N_A_1689_424#_c_1219_n 0.00380673f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_208 VPB N_CI_c_1330_n 0.0426462f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_209 VPB CI 0.00348372f $X=-0.19 $Y=1.66 $X2=0.585 $Y2=0.74
cc_210 VPB N_A_1451_424#_c_1381_n 0.018531f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.765
cc_211 VPB N_A_1451_424#_c_1382_n 0.0148926f $X=-0.19 $Y=1.66 $X2=1.215 $Y2=1.63
cc_212 VPB N_A_1451_424#_c_1375_n 0.0137346f $X=-0.19 $Y=1.66 $X2=1.31 $Y2=1.12
cc_213 VPB N_A_1451_424#_c_1377_n 0.00750439f $X=-0.19 $Y=1.66 $X2=0.985
+ $Y2=1.465
cc_214 VPB N_A_1895_424#_c_1511_n 0.0148511f $X=-0.19 $Y=1.66 $X2=0.495
+ $Y2=1.765
cc_215 VPB N_A_1895_424#_c_1512_n 0.0175006f $X=-0.19 $Y=1.66 $X2=0.532
+ $Y2=1.465
cc_216 VPB N_A_1895_424#_c_1513_n 0.00201069f $X=-0.19 $Y=1.66 $X2=0.985
+ $Y2=1.465
cc_217 VPB N_A_1895_424#_c_1514_n 0.0125217f $X=-0.19 $Y=1.66 $X2=1.31 $Y2=1.465
cc_218 VPB N_A_1895_424#_c_1506_n 0.00132124f $X=-0.19 $Y=1.66 $X2=1.54
+ $Y2=0.675
cc_219 VPB N_A_1895_424#_c_1508_n 0.00315987f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_220 VPB N_A_1895_424#_c_1517_n 0.00336963f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_221 VPB N_A_1895_424#_c_1518_n 0.00657878f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_222 VPB N_A_1895_424#_c_1510_n 0.0161272f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_223 VPB N_VPWR_c_1628_n 0.0104293f $X=-0.19 $Y=1.66 $X2=1.31 $Y2=1.12
cc_224 VPB N_VPWR_c_1629_n 0.043308f $X=-0.19 $Y=1.66 $X2=0.985 $Y2=1.465
cc_225 VPB N_VPWR_c_1630_n 0.00869569f $X=-0.19 $Y=1.66 $X2=1.215 $Y2=1.465
cc_226 VPB N_VPWR_c_1631_n 0.0102397f $X=-0.19 $Y=1.66 $X2=1.465 $Y2=1.12
cc_227 VPB N_VPWR_c_1632_n 0.0102199f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_228 VPB N_VPWR_c_1633_n 0.0027459f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_229 VPB N_VPWR_c_1634_n 0.0103331f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_230 VPB N_VPWR_c_1635_n 0.0576732f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_231 VPB N_VPWR_c_1636_n 0.0328287f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_232 VPB N_VPWR_c_1637_n 0.103306f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_233 VPB N_VPWR_c_1638_n 0.110411f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_234 VPB N_VPWR_c_1639_n 0.0207068f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_235 VPB N_VPWR_c_1640_n 0.0177589f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_236 VPB N_VPWR_c_1641_n 0.0188912f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_237 VPB N_VPWR_c_1642_n 0.00614127f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_238 VPB N_VPWR_c_1643_n 0.00614127f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_239 VPB N_VPWR_c_1644_n 0.0152669f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_240 VPB N_VPWR_c_1645_n 0.00614248f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_241 VPB N_VPWR_c_1646_n 0.00601765f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_242 VPB N_VPWR_c_1627_n 0.165827f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_243 VPB N_A_114_368#_c_1757_n 0.00860109f $X=-0.19 $Y=1.66 $X2=0.532
+ $Y2=1.465
cc_244 VPB N_A_114_368#_c_1766_n 0.0117795f $X=-0.19 $Y=1.66 $X2=1.215 $Y2=2.105
cc_245 VPB N_A_114_368#_c_1760_n 0.00350404f $X=-0.19 $Y=1.66 $X2=1.215
+ $Y2=1.465
cc_246 VPB N_A_114_368#_c_1768_n 0.00389125f $X=-0.19 $Y=1.66 $X2=1.54 $Y2=0.675
cc_247 VPB N_A_413_392#_c_1864_n 7.85085e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_248 VPB N_A_413_392#_c_1865_n 0.0304019f $X=-0.19 $Y=1.66 $X2=1.31 $Y2=1.3
cc_249 VPB N_A_413_392#_c_1866_n 0.00238428f $X=-0.19 $Y=1.66 $X2=0.985
+ $Y2=1.465
cc_250 VPB N_A_413_392#_c_1867_n 0.00512971f $X=-0.19 $Y=1.66 $X2=1.31 $Y2=1.465
cc_251 VPB N_A_413_392#_c_1861_n 0.00575237f $X=-0.19 $Y=1.66 $X2=1.465
+ $Y2=0.675
cc_252 VPB N_A_2052_424#_c_1946_n 0.00391383f $X=-0.19 $Y=1.66 $X2=1.215
+ $Y2=1.63
cc_253 VPB N_SUM_c_2010_n 0.00169264f $X=-0.19 $Y=1.66 $X2=0.585 $Y2=0.74
cc_254 VPB N_SUM_c_2011_n 0.00226359f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_255 VPB N_SUM_c_2008_n 0.00117332f $X=-0.19 $Y=1.66 $X2=1.215 $Y2=2.815
cc_256 N_A_81_260#_c_260_n N_A_c_316_n 0.00797678f $X=1.255 $Y=2.105 $X2=0 $Y2=0
cc_257 N_A_81_260#_c_263_n N_A_c_316_n 4.048e-19 $X=1.31 $Y=1.465 $X2=0 $Y2=0
cc_258 N_A_81_260#_c_260_n N_A_c_322_n 0.0067129f $X=1.255 $Y=2.105 $X2=0 $Y2=0
cc_259 N_A_81_260#_c_261_n N_A_c_317_n 0.00420059f $X=1.31 $Y=1.3 $X2=0 $Y2=0
cc_260 N_A_81_260#_c_264_n N_A_c_317_n 0.0119793f $X=1.54 $Y=0.675 $X2=0 $Y2=0
cc_261 N_A_81_260#_c_260_n N_A_c_325_n 0.0096504f $X=1.255 $Y=2.105 $X2=0 $Y2=0
cc_262 N_A_81_260#_c_261_n N_A_c_325_n 5.90453e-19 $X=1.31 $Y=1.3 $X2=0 $Y2=0
cc_263 N_A_81_260#_c_262_n N_A_c_325_n 2.342e-19 $X=0.985 $Y=1.465 $X2=0 $Y2=0
cc_264 N_A_81_260#_c_263_n N_A_c_325_n 0.0256562f $X=1.31 $Y=1.465 $X2=0 $Y2=0
cc_265 N_A_81_260#_c_264_n N_A_c_325_n 0.00905679f $X=1.54 $Y=0.675 $X2=0 $Y2=0
cc_266 N_A_81_260#_c_261_n N_A_c_320_n 2.44171e-19 $X=1.31 $Y=1.3 $X2=0 $Y2=0
cc_267 N_A_81_260#_c_262_n N_A_c_320_n 0.0182968f $X=0.985 $Y=1.465 $X2=0 $Y2=0
cc_268 N_A_81_260#_c_263_n N_A_c_320_n 0.00761182f $X=1.31 $Y=1.465 $X2=0 $Y2=0
cc_269 N_A_81_260#_c_264_n N_A_c_320_n 0.00931944f $X=1.54 $Y=0.675 $X2=0 $Y2=0
cc_270 N_A_81_260#_c_258_n N_VPWR_c_1629_n 0.0095133f $X=0.495 $Y=1.765 $X2=0
+ $Y2=0
cc_271 N_A_81_260#_c_260_n N_VPWR_c_1630_n 0.0691069f $X=1.255 $Y=2.105 $X2=0
+ $Y2=0
cc_272 N_A_81_260#_c_258_n N_VPWR_c_1636_n 0.00445602f $X=0.495 $Y=1.765 $X2=0
+ $Y2=0
cc_273 N_A_81_260#_c_260_n N_VPWR_c_1636_n 0.011066f $X=1.255 $Y=2.105 $X2=0
+ $Y2=0
cc_274 N_A_81_260#_c_258_n N_VPWR_c_1627_n 0.0086574f $X=0.495 $Y=1.765 $X2=0
+ $Y2=0
cc_275 N_A_81_260#_c_260_n N_VPWR_c_1627_n 0.00915947f $X=1.255 $Y=2.105 $X2=0
+ $Y2=0
cc_276 N_A_81_260#_c_258_n N_A_114_368#_c_1757_n 0.0193504f $X=0.495 $Y=1.765
+ $X2=0 $Y2=0
cc_277 N_A_81_260#_c_260_n N_A_114_368#_c_1757_n 0.00800222f $X=1.255 $Y=2.105
+ $X2=0 $Y2=0
cc_278 N_A_81_260#_c_263_n N_A_114_368#_c_1757_n 0.0124434f $X=1.31 $Y=1.465
+ $X2=0 $Y2=0
cc_279 N_A_81_260#_c_258_n N_A_114_368#_c_1766_n 0.0175207f $X=0.495 $Y=1.765
+ $X2=0 $Y2=0
cc_280 N_A_81_260#_c_260_n N_A_114_368#_c_1766_n 0.0708045f $X=1.255 $Y=2.105
+ $X2=0 $Y2=0
cc_281 N_A_81_260#_M1034_g N_A_114_368#_c_1758_n 0.00131834f $X=0.585 $Y=0.74
+ $X2=0 $Y2=0
cc_282 N_A_81_260#_c_264_n N_A_114_368#_c_1758_n 0.0284815f $X=1.54 $Y=0.675
+ $X2=0 $Y2=0
cc_283 N_A_81_260#_c_258_n N_A_114_368#_c_1768_n 0.0202169f $X=0.495 $Y=1.765
+ $X2=0 $Y2=0
cc_284 N_A_81_260#_c_260_n N_A_114_368#_c_1768_n 0.0125537f $X=1.255 $Y=2.105
+ $X2=0 $Y2=0
cc_285 N_A_81_260#_c_263_n N_A_114_368#_c_1768_n 0.00424948f $X=1.31 $Y=1.465
+ $X2=0 $Y2=0
cc_286 N_A_81_260#_M1034_g N_A_114_368#_c_1761_n 0.00127632f $X=0.585 $Y=0.74
+ $X2=0 $Y2=0
cc_287 N_A_81_260#_c_260_n N_A_114_368#_c_1761_n 9.11644e-19 $X=1.255 $Y=2.105
+ $X2=0 $Y2=0
cc_288 N_A_81_260#_c_261_n N_A_114_368#_c_1761_n 0.0144711f $X=1.31 $Y=1.3 $X2=0
+ $Y2=0
cc_289 N_A_81_260#_c_262_n N_A_114_368#_c_1761_n 0.00631734f $X=0.985 $Y=1.465
+ $X2=0 $Y2=0
cc_290 N_A_81_260#_c_263_n N_A_114_368#_c_1761_n 0.0267146f $X=1.31 $Y=1.465
+ $X2=0 $Y2=0
cc_291 N_A_81_260#_c_264_n N_A_114_368#_c_1761_n 0.01337f $X=1.54 $Y=0.675 $X2=0
+ $Y2=0
cc_292 N_A_81_260#_c_258_n N_A_114_368#_c_1764_n 0.0111396f $X=0.495 $Y=1.765
+ $X2=0 $Y2=0
cc_293 N_A_81_260#_M1034_g N_A_114_368#_c_1764_n 0.019709f $X=0.585 $Y=0.74
+ $X2=0 $Y2=0
cc_294 N_A_81_260#_c_261_n N_A_114_368#_c_1764_n 0.00396224f $X=1.31 $Y=1.3
+ $X2=0 $Y2=0
cc_295 N_A_81_260#_c_262_n N_A_114_368#_c_1764_n 0.00852204f $X=0.985 $Y=1.465
+ $X2=0 $Y2=0
cc_296 N_A_81_260#_c_263_n N_A_114_368#_c_1764_n 0.0227862f $X=1.31 $Y=1.465
+ $X2=0 $Y2=0
cc_297 N_A_81_260#_c_264_n N_A_114_368#_c_1764_n 0.011112f $X=1.54 $Y=0.675
+ $X2=0 $Y2=0
cc_298 N_A_81_260#_c_258_n N_VGND_c_2044_n 3.98722e-19 $X=0.495 $Y=1.765 $X2=0
+ $Y2=0
cc_299 N_A_81_260#_M1034_g N_VGND_c_2044_n 0.0148971f $X=0.585 $Y=0.74 $X2=0
+ $Y2=0
cc_300 N_A_81_260#_c_264_n N_VGND_c_2045_n 0.0130628f $X=1.54 $Y=0.675 $X2=0
+ $Y2=0
cc_301 N_A_81_260#_M1034_g N_VGND_c_2052_n 0.00383152f $X=0.585 $Y=0.74 $X2=0
+ $Y2=0
cc_302 N_A_81_260#_c_264_n N_VGND_c_2052_n 0.0129877f $X=1.54 $Y=0.675 $X2=0
+ $Y2=0
cc_303 N_A_81_260#_M1034_g N_VGND_c_2063_n 0.00762539f $X=0.585 $Y=0.74 $X2=0
+ $Y2=0
cc_304 N_A_81_260#_c_264_n N_VGND_c_2063_n 0.0158921f $X=1.54 $Y=0.675 $X2=0
+ $Y2=0
cc_305 N_A_c_319_n N_B_M1006_g 0.0139617f $X=2.255 $Y=1.29 $X2=0 $Y2=0
cc_306 N_A_c_320_n N_B_c_389_n 2.91015e-19 $X=2.255 $Y=1.455 $X2=0 $Y2=0
cc_307 N_A_c_318_n N_B_c_390_n 0.0011792f $X=1.99 $Y=1.795 $X2=0 $Y2=0
cc_308 N_A_c_320_n N_B_c_390_n 0.0166544f $X=2.255 $Y=1.455 $X2=0 $Y2=0
cc_309 N_A_c_319_n N_B_c_391_n 3.87987e-19 $X=2.255 $Y=1.29 $X2=0 $Y2=0
cc_310 N_A_c_324_n N_A_481_379#_c_602_n 0.0189451f $X=1.99 $Y=1.885 $X2=0 $Y2=0
cc_311 N_A_c_324_n N_A_481_379#_c_604_n 0.00463694f $X=1.99 $Y=1.885 $X2=0 $Y2=0
cc_312 N_A_c_322_n N_VPWR_c_1630_n 0.0186866f $X=1.48 $Y=1.885 $X2=0 $Y2=0
cc_313 N_A_c_324_n N_VPWR_c_1630_n 0.00716177f $X=1.99 $Y=1.885 $X2=0 $Y2=0
cc_314 N_A_c_325_n N_VPWR_c_1630_n 0.0269294f $X=1.915 $Y=1.455 $X2=0 $Y2=0
cc_315 N_A_c_320_n N_VPWR_c_1630_n 8.09174e-19 $X=2.255 $Y=1.455 $X2=0 $Y2=0
cc_316 N_A_c_322_n N_VPWR_c_1636_n 0.00413917f $X=1.48 $Y=1.885 $X2=0 $Y2=0
cc_317 N_A_c_324_n N_VPWR_c_1637_n 0.00449387f $X=1.99 $Y=1.885 $X2=0 $Y2=0
cc_318 N_A_c_322_n N_VPWR_c_1627_n 0.00822528f $X=1.48 $Y=1.885 $X2=0 $Y2=0
cc_319 N_A_c_324_n N_VPWR_c_1627_n 0.00872565f $X=1.99 $Y=1.885 $X2=0 $Y2=0
cc_320 N_A_c_317_n N_A_114_368#_c_1761_n 0.00687655f $X=1.825 $Y=1.29 $X2=0
+ $Y2=0
cc_321 N_A_c_319_n N_A_114_368#_c_1761_n 0.00187082f $X=2.255 $Y=1.29 $X2=0
+ $Y2=0
cc_322 N_A_c_325_n N_A_114_368#_c_1761_n 0.0243406f $X=1.915 $Y=1.455 $X2=0
+ $Y2=0
cc_323 N_A_c_320_n N_A_114_368#_c_1761_n 0.0167594f $X=2.255 $Y=1.455 $X2=0
+ $Y2=0
cc_324 N_A_c_324_n N_A_413_392#_c_1864_n 0.00246973f $X=1.99 $Y=1.885 $X2=0
+ $Y2=0
cc_325 N_A_c_320_n N_A_413_392#_c_1864_n 0.00431505f $X=2.255 $Y=1.455 $X2=0
+ $Y2=0
cc_326 N_A_c_324_n N_A_413_392#_c_1871_n 0.00900274f $X=1.99 $Y=1.885 $X2=0
+ $Y2=0
cc_327 N_A_c_317_n N_A_413_392#_c_1858_n 6.32307e-19 $X=1.825 $Y=1.29 $X2=0
+ $Y2=0
cc_328 N_A_c_319_n N_A_413_392#_c_1858_n 0.00836151f $X=2.255 $Y=1.29 $X2=0
+ $Y2=0
cc_329 N_A_c_324_n N_A_413_392#_c_1866_n 0.00309192f $X=1.99 $Y=1.885 $X2=0
+ $Y2=0
cc_330 N_A_c_319_n N_A_413_392#_c_1860_n 0.0010929f $X=2.255 $Y=1.29 $X2=0 $Y2=0
cc_331 N_A_c_318_n N_A_413_392#_c_1861_n 0.00628793f $X=1.99 $Y=1.795 $X2=0
+ $Y2=0
cc_332 N_A_c_324_n N_A_413_392#_c_1861_n 0.00207727f $X=1.99 $Y=1.885 $X2=0
+ $Y2=0
cc_333 N_A_c_319_n N_A_413_392#_c_1861_n 0.00322503f $X=2.255 $Y=1.29 $X2=0
+ $Y2=0
cc_334 N_A_c_325_n N_A_413_392#_c_1861_n 0.0360454f $X=1.915 $Y=1.455 $X2=0
+ $Y2=0
cc_335 N_A_c_320_n N_A_413_392#_c_1861_n 0.0115321f $X=2.255 $Y=1.455 $X2=0
+ $Y2=0
cc_336 N_A_c_317_n N_A_413_392#_c_1862_n 0.00155092f $X=1.825 $Y=1.29 $X2=0
+ $Y2=0
cc_337 N_A_c_319_n N_A_413_392#_c_1862_n 0.00864538f $X=2.255 $Y=1.29 $X2=0
+ $Y2=0
cc_338 N_A_c_317_n N_VGND_c_2045_n 0.0105093f $X=1.825 $Y=1.29 $X2=0 $Y2=0
cc_339 N_A_c_319_n N_VGND_c_2045_n 9.5937e-19 $X=2.255 $Y=1.29 $X2=0 $Y2=0
cc_340 N_A_c_325_n N_VGND_c_2045_n 0.0029985f $X=1.915 $Y=1.455 $X2=0 $Y2=0
cc_341 N_A_c_320_n N_VGND_c_2045_n 0.0020495f $X=2.255 $Y=1.455 $X2=0 $Y2=0
cc_342 N_A_c_317_n N_VGND_c_2052_n 0.00392356f $X=1.825 $Y=1.29 $X2=0 $Y2=0
cc_343 N_A_c_319_n N_VGND_c_2056_n 0.00404525f $X=2.255 $Y=1.29 $X2=0 $Y2=0
cc_344 N_A_c_317_n N_VGND_c_2063_n 0.00418286f $X=1.825 $Y=1.29 $X2=0 $Y2=0
cc_345 N_A_c_319_n N_VGND_c_2063_n 0.00414967f $X=2.255 $Y=1.29 $X2=0 $Y2=0
cc_346 B N_A_481_379#_c_602_n 0.00337663f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_347 N_B_c_382_n N_A_481_379#_c_603_n 0.00435974f $X=3.56 $Y=2.045 $X2=0 $Y2=0
cc_348 B N_A_481_379#_c_603_n 0.0151394f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_349 N_B_c_390_n N_A_481_379#_c_604_n 0.0215523f $X=2.705 $Y=1.52 $X2=0 $Y2=0
cc_350 B N_A_481_379#_c_604_n 0.00162584f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_351 N_B_c_382_n N_A_481_379#_c_591_n 0.0206595f $X=3.56 $Y=2.045 $X2=0 $Y2=0
cc_352 N_B_c_389_n N_A_481_379#_c_591_n 0.00143137f $X=2.705 $Y=1.52 $X2=0 $Y2=0
cc_353 N_B_c_392_n N_A_481_379#_c_591_n 4.15056e-19 $X=3.605 $Y=1.795 $X2=0
+ $Y2=0
cc_354 N_B_c_393_n N_A_481_379#_c_591_n 0.00146447f $X=3.605 $Y=1.63 $X2=0 $Y2=0
cc_355 N_B_M1006_g N_A_481_379#_c_592_n 0.0108575f $X=2.685 $Y=0.845 $X2=0 $Y2=0
cc_356 N_B_c_419_p N_A_481_379#_c_592_n 0.0146196f $X=3.565 $Y=0.68 $X2=0 $Y2=0
cc_357 N_B_c_391_n N_A_481_379#_c_592_n 0.00126497f $X=2.725 $Y=1.355 $X2=0
+ $Y2=0
cc_358 N_B_c_393_n N_A_481_379#_c_592_n 0.00946779f $X=3.605 $Y=1.63 $X2=0 $Y2=0
cc_359 N_B_c_422_p N_A_481_379#_c_593_n 0.00420841f $X=4.405 $Y=0.68 $X2=0 $Y2=0
cc_360 N_B_c_387_n N_A_481_379#_c_593_n 0.0197433f $X=4.505 $Y=1.44 $X2=0 $Y2=0
cc_361 N_B_c_392_n N_A_481_379#_c_593_n 2.20813e-19 $X=3.605 $Y=1.795 $X2=0
+ $Y2=0
cc_362 N_B_c_393_n N_A_481_379#_c_593_n 0.0116988f $X=3.605 $Y=1.63 $X2=0 $Y2=0
cc_363 N_B_c_396_n N_A_481_379#_c_593_n 0.00172145f $X=4.505 $Y=1.275 $X2=0
+ $Y2=0
cc_364 N_B_M1006_g N_A_481_379#_c_594_n 0.00437192f $X=2.685 $Y=0.845 $X2=0
+ $Y2=0
cc_365 N_B_c_382_n N_A_481_379#_c_594_n 0.0179165f $X=3.56 $Y=2.045 $X2=0 $Y2=0
cc_366 N_B_c_419_p N_A_481_379#_c_594_n 6.57854e-19 $X=3.565 $Y=0.68 $X2=0 $Y2=0
cc_367 N_B_c_390_n N_A_481_379#_c_594_n 0.02131f $X=2.705 $Y=1.52 $X2=0 $Y2=0
cc_368 N_B_c_391_n N_A_481_379#_c_594_n 0.00143137f $X=2.725 $Y=1.355 $X2=0
+ $Y2=0
cc_369 N_B_c_392_n N_A_481_379#_c_594_n 8.89205e-19 $X=3.605 $Y=1.795 $X2=0
+ $Y2=0
cc_370 N_B_c_382_n N_A_481_379#_c_595_n 0.020571f $X=3.56 $Y=2.045 $X2=0 $Y2=0
cc_371 N_B_c_386_n N_A_481_379#_c_595_n 5.45615e-19 $X=4.505 $Y=1.44 $X2=0 $Y2=0
cc_372 N_B_c_392_n N_A_481_379#_c_595_n 3.81338e-19 $X=3.605 $Y=1.795 $X2=0
+ $Y2=0
cc_373 N_B_c_393_n N_A_481_379#_c_595_n 0.00149745f $X=3.605 $Y=1.63 $X2=0 $Y2=0
cc_374 N_B_c_382_n N_A_481_379#_c_607_n 0.0260793f $X=3.56 $Y=2.045 $X2=0 $Y2=0
cc_375 N_B_c_386_n N_A_481_379#_c_608_n 7.01095e-19 $X=4.505 $Y=1.44 $X2=0 $Y2=0
cc_376 N_B_c_387_n N_A_481_379#_c_608_n 0.0178647f $X=4.505 $Y=1.44 $X2=0 $Y2=0
cc_377 N_B_c_382_n N_A_481_379#_c_609_n 0.00234057f $X=3.56 $Y=2.045 $X2=0 $Y2=0
cc_378 N_B_c_387_n N_A_481_379#_c_596_n 0.00924236f $X=4.505 $Y=1.44 $X2=0 $Y2=0
cc_379 N_B_c_442_p N_A_481_379#_c_596_n 0.0025088f $X=5.265 $Y=0.68 $X2=0 $Y2=0
cc_380 N_B_c_396_n N_A_481_379#_c_596_n 3.56848e-19 $X=4.505 $Y=1.275 $X2=0
+ $Y2=0
cc_381 N_B_c_384_n N_A_481_379#_c_597_n 0.015925f $X=6.745 $Y=1.315 $X2=0 $Y2=0
cc_382 N_B_c_386_n N_A_481_379#_c_597_n 0.00146916f $X=4.505 $Y=1.44 $X2=0 $Y2=0
cc_383 N_B_c_442_p N_A_481_379#_c_597_n 0.0117513f $X=5.265 $Y=0.68 $X2=0 $Y2=0
cc_384 N_B_c_447_p N_A_481_379#_c_597_n 0.00659127f $X=5.35 $Y=0.92 $X2=0 $Y2=0
cc_385 N_B_c_448_p N_A_481_379#_c_597_n 0.00723096f $X=5.435 $Y=1.005 $X2=0
+ $Y2=0
cc_386 N_B_c_394_n N_A_481_379#_c_597_n 6.1072e-19 $X=6.04 $Y=1.005 $X2=0 $Y2=0
cc_387 N_B_c_396_n N_A_481_379#_c_597_n 0.0104779f $X=4.505 $Y=1.275 $X2=0 $Y2=0
cc_388 N_B_c_399_n N_A_481_379#_c_610_n 0.00904828f $X=6.655 $Y=1.765 $X2=0
+ $Y2=0
cc_389 N_B_c_384_n N_A_481_379#_c_610_n 0.0435266f $X=6.745 $Y=1.315 $X2=0 $Y2=0
cc_390 N_B_c_383_n N_A_481_379#_c_598_n 0.00940821f $X=7.05 $Y=1.315 $X2=0 $Y2=0
cc_391 N_B_c_384_n N_A_481_379#_c_598_n 0.0210249f $X=6.745 $Y=1.315 $X2=0 $Y2=0
cc_392 N_B_c_383_n N_A_481_379#_c_599_n 0.0139892f $X=7.05 $Y=1.315 $X2=0 $Y2=0
cc_393 N_B_c_384_n N_A_481_379#_c_599_n 0.00254469f $X=6.745 $Y=1.315 $X2=0
+ $Y2=0
cc_394 N_B_M1033_g N_A_481_379#_c_599_n 0.00786938f $X=7.125 $Y=0.74 $X2=0 $Y2=0
cc_395 N_B_M1033_g N_A_481_379#_c_600_n 0.0106204f $X=7.125 $Y=0.74 $X2=0 $Y2=0
cc_396 N_B_c_384_n N_A_481_379#_c_666_n 0.00131418f $X=6.745 $Y=1.315 $X2=0
+ $Y2=0
cc_397 N_B_c_384_n N_A_481_379#_c_601_n 0.0247303f $X=6.745 $Y=1.315 $X2=0 $Y2=0
cc_398 N_B_c_399_n N_A_481_379#_c_613_n 0.00780793f $X=6.655 $Y=1.765 $X2=0
+ $Y2=0
cc_399 N_B_c_384_n N_A_481_379#_c_613_n 3.62163e-19 $X=6.745 $Y=1.315 $X2=0
+ $Y2=0
cc_400 N_B_c_419_p N_A_514_424#_M1006_d 0.0118424f $X=3.565 $Y=0.68 $X2=-0.19
+ $Y2=-0.245
cc_401 N_B_c_464_p N_A_514_424#_M1006_d 8.24664e-19 $X=2.895 $Y=0.68 $X2=-0.19
+ $Y2=-0.245
cc_402 N_B_c_391_n N_A_514_424#_M1006_d 0.00490871f $X=2.725 $Y=1.355 $X2=-0.19
+ $Y2=-0.245
cc_403 B N_A_514_424#_M1003_d 0.0037536f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_404 N_B_c_399_n N_A_514_424#_c_758_n 0.0350095f $X=6.655 $Y=1.765 $X2=0 $Y2=0
cc_405 N_B_c_383_n N_A_514_424#_c_758_n 0.00728162f $X=7.05 $Y=1.315 $X2=0 $Y2=0
cc_406 N_B_c_384_n N_A_514_424#_c_758_n 0.00437122f $X=6.745 $Y=1.315 $X2=0
+ $Y2=0
cc_407 B N_A_514_424#_c_796_n 0.0184267f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_408 N_B_c_382_n N_A_514_424#_c_762_n 0.0111992f $X=3.56 $Y=2.045 $X2=0 $Y2=0
cc_409 N_B_c_389_n N_A_514_424#_c_762_n 0.0465238f $X=2.705 $Y=1.52 $X2=0 $Y2=0
cc_410 N_B_c_390_n N_A_514_424#_c_762_n 9.0699e-19 $X=2.705 $Y=1.52 $X2=0 $Y2=0
cc_411 N_B_c_392_n N_A_514_424#_c_762_n 0.0215497f $X=3.605 $Y=1.795 $X2=0 $Y2=0
cc_412 N_B_c_393_n N_A_514_424#_c_762_n 0.0185316f $X=3.605 $Y=1.63 $X2=0 $Y2=0
cc_413 N_B_c_382_n N_A_514_424#_c_802_n 0.0151103f $X=3.56 $Y=2.045 $X2=0 $Y2=0
cc_414 N_B_c_392_n N_A_514_424#_c_802_n 0.0040144f $X=3.605 $Y=1.795 $X2=0 $Y2=0
cc_415 N_B_c_398_n N_A_514_424#_c_775_n 0.0152167f $X=5.665 $Y=2.045 $X2=0 $Y2=0
cc_416 N_B_c_384_n N_A_514_424#_c_775_n 0.00256011f $X=6.745 $Y=1.315 $X2=0
+ $Y2=0
cc_417 N_B_c_399_n N_A_514_424#_c_806_n 0.0167834f $X=6.655 $Y=1.765 $X2=0 $Y2=0
cc_418 N_B_c_384_n N_A_514_424#_c_806_n 4.29596e-19 $X=6.745 $Y=1.315 $X2=0
+ $Y2=0
cc_419 N_B_c_399_n N_A_514_424#_c_777_n 5.49231e-19 $X=6.655 $Y=1.765 $X2=0
+ $Y2=0
cc_420 N_B_c_399_n N_A_514_424#_c_809_n 0.00185586f $X=6.655 $Y=1.765 $X2=0
+ $Y2=0
cc_421 N_B_c_399_n N_A_514_424#_c_779_n 5.39168e-19 $X=6.655 $Y=1.765 $X2=0
+ $Y2=0
cc_422 N_B_M1006_g N_A_514_424#_c_766_n 0.00115407f $X=2.685 $Y=0.845 $X2=0
+ $Y2=0
cc_423 N_B_c_419_p N_A_514_424#_c_766_n 0.0204713f $X=3.565 $Y=0.68 $X2=0 $Y2=0
cc_424 N_B_c_391_n N_A_514_424#_c_766_n 0.0465238f $X=2.725 $Y=1.355 $X2=0 $Y2=0
cc_425 N_B_c_393_n N_A_514_424#_c_766_n 0.010084f $X=3.605 $Y=1.63 $X2=0 $Y2=0
cc_426 N_B_c_398_n N_A_514_424#_c_783_n 0.00270588f $X=5.665 $Y=2.045 $X2=0
+ $Y2=0
cc_427 N_B_c_399_n N_A_514_424#_c_783_n 0.00554556f $X=6.655 $Y=1.765 $X2=0
+ $Y2=0
cc_428 N_B_c_384_n N_A_514_424#_c_783_n 8.28086e-19 $X=6.745 $Y=1.315 $X2=0
+ $Y2=0
cc_429 N_B_c_386_n N_A_849_424#_M1007_d 0.00517147f $X=4.505 $Y=1.44 $X2=-0.19
+ $Y2=-0.245
cc_430 N_B_c_442_p N_A_849_424#_M1007_d 0.0180031f $X=5.265 $Y=0.68 $X2=-0.19
+ $Y2=-0.245
cc_431 N_B_c_383_n N_A_849_424#_c_1004_n 0.0129921f $X=7.05 $Y=1.315 $X2=0 $Y2=0
cc_432 N_B_M1033_g N_A_849_424#_c_1004_n 0.0105359f $X=7.125 $Y=0.74 $X2=0 $Y2=0
cc_433 N_B_c_398_n N_A_849_424#_c_1013_n 0.00112071f $X=5.665 $Y=2.045 $X2=0
+ $Y2=0
cc_434 N_B_c_384_n N_A_849_424#_c_1013_n 0.00127148f $X=6.745 $Y=1.315 $X2=0
+ $Y2=0
cc_435 N_B_c_398_n N_A_849_424#_c_1037_n 0.00101863f $X=5.665 $Y=2.045 $X2=0
+ $Y2=0
cc_436 N_B_c_442_p N_A_849_424#_c_1014_n 0.0041436f $X=5.265 $Y=0.68 $X2=0 $Y2=0
cc_437 N_B_c_388_n N_A_849_424#_c_1014_n 0.0073604f $X=5.875 $Y=1.005 $X2=0
+ $Y2=0
cc_438 N_B_c_448_p N_A_849_424#_c_1014_n 0.010622f $X=5.435 $Y=1.005 $X2=0 $Y2=0
cc_439 N_B_c_384_n N_A_849_424#_c_1015_n 0.0416061f $X=6.745 $Y=1.315 $X2=0
+ $Y2=0
cc_440 N_B_c_388_n N_A_849_424#_c_1015_n 0.00940058f $X=5.875 $Y=1.005 $X2=0
+ $Y2=0
cc_441 N_B_c_394_n N_A_849_424#_c_1015_n 0.0231396f $X=6.04 $Y=1.005 $X2=0 $Y2=0
cc_442 N_B_c_384_n N_A_849_424#_c_1016_n 0.0159838f $X=6.745 $Y=1.315 $X2=0
+ $Y2=0
cc_443 N_B_M1033_g N_A_849_424#_c_1016_n 0.00285863f $X=7.125 $Y=0.74 $X2=0
+ $Y2=0
cc_444 N_B_c_394_n N_A_849_424#_c_1016_n 0.0123632f $X=6.04 $Y=1.005 $X2=0 $Y2=0
cc_445 N_B_c_383_n N_A_849_424#_c_1017_n 8.77712e-19 $X=7.05 $Y=1.315 $X2=0
+ $Y2=0
cc_446 N_B_c_384_n N_A_849_424#_c_1017_n 0.00740778f $X=6.745 $Y=1.315 $X2=0
+ $Y2=0
cc_447 N_B_c_384_n N_A_849_424#_c_1018_n 0.00232042f $X=6.745 $Y=1.315 $X2=0
+ $Y2=0
cc_448 N_B_c_394_n N_A_849_424#_c_1018_n 0.00838009f $X=6.04 $Y=1.005 $X2=0
+ $Y2=0
cc_449 N_B_M1033_g N_A_849_424#_c_1019_n 0.0144968f $X=7.125 $Y=0.74 $X2=0 $Y2=0
cc_450 N_B_c_383_n N_A_849_424#_c_1021_n 2.96363e-19 $X=7.05 $Y=1.315 $X2=0
+ $Y2=0
cc_451 N_B_c_386_n N_A_849_424#_c_1023_n 0.0502964f $X=4.505 $Y=1.44 $X2=0 $Y2=0
cc_452 N_B_c_387_n N_A_849_424#_c_1023_n 0.00283504f $X=4.505 $Y=1.44 $X2=0
+ $Y2=0
cc_453 N_B_c_442_p N_A_849_424#_c_1023_n 0.0263573f $X=5.265 $Y=0.68 $X2=0 $Y2=0
cc_454 N_B_c_448_p N_A_849_424#_c_1023_n 0.0126662f $X=5.435 $Y=1.005 $X2=0
+ $Y2=0
cc_455 N_B_c_396_n N_A_849_424#_c_1023_n 0.00128049f $X=4.505 $Y=1.275 $X2=0
+ $Y2=0
cc_456 N_B_c_386_n N_A_849_424#_c_1039_n 0.00685751f $X=4.505 $Y=1.44 $X2=0
+ $Y2=0
cc_457 N_B_c_384_n N_A_849_424#_c_1024_n 0.00492316f $X=6.745 $Y=1.315 $X2=0
+ $Y2=0
cc_458 N_B_c_388_n N_A_849_424#_c_1024_n 0.0130487f $X=5.875 $Y=1.005 $X2=0
+ $Y2=0
cc_459 N_B_c_398_n N_VPWR_c_1631_n 0.00208106f $X=5.665 $Y=2.045 $X2=0 $Y2=0
cc_460 N_B_c_399_n N_VPWR_c_1631_n 0.0130843f $X=6.655 $Y=1.765 $X2=0 $Y2=0
cc_461 N_B_c_382_n N_VPWR_c_1637_n 0.00280451f $X=3.56 $Y=2.045 $X2=0 $Y2=0
cc_462 N_B_c_398_n N_VPWR_c_1637_n 0.00280437f $X=5.665 $Y=2.045 $X2=0 $Y2=0
cc_463 N_B_c_399_n N_VPWR_c_1638_n 0.00413917f $X=6.655 $Y=1.765 $X2=0 $Y2=0
cc_464 N_B_c_382_n N_VPWR_c_1627_n 0.00360251f $X=3.56 $Y=2.045 $X2=0 $Y2=0
cc_465 N_B_c_398_n N_VPWR_c_1627_n 0.00363715f $X=5.665 $Y=2.045 $X2=0 $Y2=0
cc_466 N_B_c_399_n N_VPWR_c_1627_n 0.00818442f $X=6.655 $Y=1.765 $X2=0 $Y2=0
cc_467 N_B_c_422_p N_A_114_368#_M1008_d 0.017361f $X=4.405 $Y=0.68 $X2=0 $Y2=0
cc_468 N_B_c_393_n N_A_114_368#_M1008_d 0.00652478f $X=3.605 $Y=1.63 $X2=0 $Y2=0
cc_469 N_B_c_532_p N_A_114_368#_M1008_d 0.00199981f $X=3.65 $Y=0.68 $X2=0 $Y2=0
cc_470 N_B_c_382_n N_A_114_368#_c_1798_n 0.0091966f $X=3.56 $Y=2.045 $X2=0 $Y2=0
cc_471 N_B_c_392_n N_A_114_368#_c_1798_n 0.00964483f $X=3.605 $Y=1.795 $X2=0
+ $Y2=0
cc_472 N_B_c_422_p N_A_114_368#_c_1759_n 0.0252577f $X=4.405 $Y=0.68 $X2=0 $Y2=0
cc_473 N_B_c_386_n N_A_114_368#_c_1759_n 0.034324f $X=4.505 $Y=1.44 $X2=0 $Y2=0
cc_474 N_B_c_387_n N_A_114_368#_c_1759_n 8.57673e-19 $X=4.505 $Y=1.44 $X2=0
+ $Y2=0
cc_475 N_B_c_393_n N_A_114_368#_c_1759_n 0.0312978f $X=3.605 $Y=1.63 $X2=0 $Y2=0
cc_476 N_B_c_396_n N_A_114_368#_c_1759_n 0.00638897f $X=4.505 $Y=1.275 $X2=0
+ $Y2=0
cc_477 N_B_c_382_n N_A_114_368#_c_1760_n 0.00494839f $X=3.56 $Y=2.045 $X2=0
+ $Y2=0
cc_478 N_B_c_386_n N_A_114_368#_c_1760_n 0.00855772f $X=4.505 $Y=1.44 $X2=0
+ $Y2=0
cc_479 N_B_c_387_n N_A_114_368#_c_1760_n 6.92371e-19 $X=4.505 $Y=1.44 $X2=0
+ $Y2=0
cc_480 N_B_c_392_n N_A_114_368#_c_1760_n 0.0248017f $X=3.605 $Y=1.795 $X2=0
+ $Y2=0
cc_481 N_B_c_393_n N_A_114_368#_c_1760_n 0.0144589f $X=3.605 $Y=1.63 $X2=0 $Y2=0
cc_482 N_B_M1006_g N_A_114_368#_c_1761_n 0.00559595f $X=2.685 $Y=0.845 $X2=0
+ $Y2=0
cc_483 N_B_c_419_p N_A_114_368#_c_1761_n 0.0118231f $X=3.565 $Y=0.68 $X2=0 $Y2=0
cc_484 N_B_c_422_p N_A_114_368#_c_1761_n 0.00587363f $X=4.405 $Y=0.68 $X2=0
+ $Y2=0
cc_485 N_B_c_389_n N_A_114_368#_c_1761_n 0.0129237f $X=2.705 $Y=1.52 $X2=0 $Y2=0
cc_486 N_B_c_390_n N_A_114_368#_c_1761_n 0.00102947f $X=2.705 $Y=1.52 $X2=0
+ $Y2=0
cc_487 N_B_c_391_n N_A_114_368#_c_1761_n 0.0148095f $X=2.725 $Y=1.355 $X2=0
+ $Y2=0
cc_488 N_B_c_392_n N_A_114_368#_c_1761_n 0.00580183f $X=3.605 $Y=1.795 $X2=0
+ $Y2=0
cc_489 N_B_c_393_n N_A_114_368#_c_1761_n 0.0198691f $X=3.605 $Y=1.63 $X2=0 $Y2=0
cc_490 N_B_c_422_p N_A_114_368#_c_1763_n 0.00127969f $X=4.405 $Y=0.68 $X2=0
+ $Y2=0
cc_491 N_B_c_386_n N_A_114_368#_c_1763_n 0.00155876f $X=4.505 $Y=1.44 $X2=0
+ $Y2=0
cc_492 N_B_c_393_n N_A_114_368#_c_1763_n 0.00232151f $X=3.605 $Y=1.63 $X2=0
+ $Y2=0
cc_493 N_B_c_442_p N_A_413_392#_M1025_d 0.00253226f $X=5.265 $Y=0.68 $X2=0 $Y2=0
cc_494 N_B_c_447_p N_A_413_392#_M1025_d 0.0058378f $X=5.35 $Y=0.92 $X2=0 $Y2=0
cc_495 N_B_c_388_n N_A_413_392#_M1025_d 0.00563474f $X=5.875 $Y=1.005 $X2=0
+ $Y2=0
cc_496 B N_A_413_392#_c_1864_n 0.0299068f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_497 N_B_M1006_g N_A_413_392#_c_1858_n 0.00267229f $X=2.685 $Y=0.845 $X2=0
+ $Y2=0
cc_498 N_B_c_382_n N_A_413_392#_c_1865_n 0.0121547f $X=3.56 $Y=2.045 $X2=0 $Y2=0
cc_499 N_B_c_398_n N_A_413_392#_c_1865_n 0.0144452f $X=5.665 $Y=2.045 $X2=0
+ $Y2=0
cc_500 N_B_c_399_n N_A_413_392#_c_1865_n 5.96651e-19 $X=6.655 $Y=1.765 $X2=0
+ $Y2=0
cc_501 N_B_M1006_g N_A_413_392#_c_1859_n 0.00944525f $X=2.685 $Y=0.845 $X2=0
+ $Y2=0
cc_502 N_B_c_419_p N_A_413_392#_c_1859_n 0.0425031f $X=3.565 $Y=0.68 $X2=0 $Y2=0
cc_503 N_B_c_464_p N_A_413_392#_c_1859_n 0.0106895f $X=2.895 $Y=0.68 $X2=0 $Y2=0
cc_504 N_B_c_422_p N_A_413_392#_c_1859_n 0.0445932f $X=4.405 $Y=0.68 $X2=0 $Y2=0
cc_505 N_B_c_442_p N_A_413_392#_c_1859_n 0.0545925f $X=5.265 $Y=0.68 $X2=0 $Y2=0
cc_506 N_B_c_388_n N_A_413_392#_c_1859_n 0.00583807f $X=5.875 $Y=1.005 $X2=0
+ $Y2=0
cc_507 N_B_c_532_p N_A_413_392#_c_1859_n 0.0126899f $X=3.65 $Y=0.68 $X2=0 $Y2=0
cc_508 N_B_c_571_p N_A_413_392#_c_1859_n 0.011743f $X=4.5 $Y=0.68 $X2=0 $Y2=0
cc_509 N_B_c_396_n N_A_413_392#_c_1859_n 0.00632285f $X=4.505 $Y=1.275 $X2=0
+ $Y2=0
cc_510 N_B_c_398_n N_A_413_392#_c_1867_n 0.0119789f $X=5.665 $Y=2.045 $X2=0
+ $Y2=0
cc_511 N_B_c_399_n N_A_413_392#_c_1867_n 0.00323287f $X=6.655 $Y=1.765 $X2=0
+ $Y2=0
cc_512 N_B_M1006_g N_A_413_392#_c_1861_n 9.23558e-19 $X=2.685 $Y=0.845 $X2=0
+ $Y2=0
cc_513 N_B_c_389_n N_A_413_392#_c_1861_n 0.0299068f $X=2.705 $Y=1.52 $X2=0 $Y2=0
cc_514 N_B_c_390_n N_A_413_392#_c_1861_n 0.00198451f $X=2.705 $Y=1.52 $X2=0
+ $Y2=0
cc_515 N_B_c_391_n N_A_413_392#_c_1861_n 0.00583011f $X=2.725 $Y=1.355 $X2=0
+ $Y2=0
cc_516 N_B_c_390_n N_A_413_392#_c_1862_n 5.46617e-19 $X=2.705 $Y=1.52 $X2=0
+ $Y2=0
cc_517 N_B_c_391_n N_A_413_392#_c_1862_n 0.0149941f $X=2.725 $Y=1.355 $X2=0
+ $Y2=0
cc_518 N_B_c_384_n N_A_413_392#_c_1863_n 4.39176e-19 $X=6.745 $Y=1.315 $X2=0
+ $Y2=0
cc_519 N_B_c_442_p N_A_413_392#_c_1863_n 0.0132003f $X=5.265 $Y=0.68 $X2=0 $Y2=0
cc_520 N_B_c_388_n N_A_413_392#_c_1863_n 0.0216761f $X=5.875 $Y=1.005 $X2=0
+ $Y2=0
cc_521 N_B_c_394_n N_A_413_392#_c_1863_n 0.00465239f $X=6.04 $Y=1.005 $X2=0
+ $Y2=0
cc_522 N_B_c_384_n N_VGND_c_2046_n 0.0015889f $X=6.745 $Y=1.315 $X2=0 $Y2=0
cc_523 N_B_M1033_g N_VGND_c_2046_n 0.00162438f $X=7.125 $Y=0.74 $X2=0 $Y2=0
cc_524 N_B_M1033_g N_VGND_c_2054_n 0.00278271f $X=7.125 $Y=0.74 $X2=0 $Y2=0
cc_525 N_B_M1006_g N_VGND_c_2056_n 6.67145e-19 $X=2.685 $Y=0.845 $X2=0 $Y2=0
cc_526 N_B_c_396_n N_VGND_c_2056_n 6.67145e-19 $X=4.505 $Y=1.275 $X2=0 $Y2=0
cc_527 N_B_M1033_g N_VGND_c_2063_n 0.00363426f $X=7.125 $Y=0.74 $X2=0 $Y2=0
cc_528 N_A_481_379#_c_598_n N_A_514_424#_c_758_n 0.00403196f $X=6.88 $Y=1.76
+ $X2=0 $Y2=0
cc_529 N_A_481_379#_c_599_n N_A_514_424#_c_758_n 0.00321482f $X=7.34 $Y=1.19
+ $X2=0 $Y2=0
cc_530 N_A_481_379#_c_613_n N_A_514_424#_c_758_n 2.08723e-19 $X=6.88 $Y=1.845
+ $X2=0 $Y2=0
cc_531 N_A_481_379#_c_602_n N_A_514_424#_c_796_n 0.00354381f $X=2.495 $Y=2.045
+ $X2=0 $Y2=0
cc_532 N_A_481_379#_c_603_n N_A_514_424#_c_796_n 0.00694294f $X=3.08 $Y=1.97
+ $X2=0 $Y2=0
cc_533 N_A_481_379#_c_602_n N_A_514_424#_c_762_n 0.00585267f $X=2.495 $Y=2.045
+ $X2=0 $Y2=0
cc_534 N_A_481_379#_c_603_n N_A_514_424#_c_762_n 0.008304f $X=3.08 $Y=1.97 $X2=0
+ $Y2=0
cc_535 N_A_481_379#_c_591_n N_A_514_424#_c_762_n 0.0141386f $X=3.155 $Y=1.895
+ $X2=0 $Y2=0
cc_536 N_A_481_379#_c_592_n N_A_514_424#_c_762_n 5.7123e-19 $X=3.445 $Y=1.24
+ $X2=0 $Y2=0
cc_537 N_A_481_379#_c_594_n N_A_514_424#_c_762_n 0.00802156f $X=3.52 $Y=1.315
+ $X2=0 $Y2=0
cc_538 N_A_481_379#_c_607_n N_A_514_424#_c_802_n 0.0174179f $X=4.17 $Y=2.045
+ $X2=0 $Y2=0
cc_539 N_A_481_379#_c_608_n N_A_514_424#_c_802_n 0.00470179f $X=5.035 $Y=1.92
+ $X2=0 $Y2=0
cc_540 N_A_481_379#_c_609_n N_A_514_424#_c_802_n 2.66147e-19 $X=4.26 $Y=1.92
+ $X2=0 $Y2=0
cc_541 N_A_481_379#_c_610_n N_A_514_424#_c_802_n 5.67708e-19 $X=6.715 $Y=1.845
+ $X2=0 $Y2=0
cc_542 N_A_481_379#_c_666_n N_A_514_424#_c_802_n 0.0039703f $X=5.2 $Y=1.765
+ $X2=0 $Y2=0
cc_543 N_A_481_379#_c_610_n N_A_514_424#_c_775_n 0.0491708f $X=6.715 $Y=1.845
+ $X2=0 $Y2=0
cc_544 N_A_481_379#_c_610_n N_A_514_424#_c_776_n 0.0142489f $X=6.715 $Y=1.845
+ $X2=0 $Y2=0
cc_545 N_A_481_379#_M1000_d N_A_514_424#_c_806_n 0.01283f $X=6.73 $Y=1.84 $X2=0
+ $Y2=0
cc_546 N_A_481_379#_c_610_n N_A_514_424#_c_806_n 0.0116364f $X=6.715 $Y=1.845
+ $X2=0 $Y2=0
cc_547 N_A_481_379#_c_613_n N_A_514_424#_c_806_n 0.022063f $X=6.88 $Y=1.845
+ $X2=0 $Y2=0
cc_548 N_A_481_379#_c_613_n N_A_514_424#_c_777_n 0.0170323f $X=6.88 $Y=1.845
+ $X2=0 $Y2=0
cc_549 N_A_481_379#_c_592_n N_A_514_424#_c_766_n 0.00360634f $X=3.445 $Y=1.24
+ $X2=0 $Y2=0
cc_550 N_A_481_379#_c_594_n N_A_514_424#_c_766_n 0.00543558f $X=3.52 $Y=1.315
+ $X2=0 $Y2=0
cc_551 N_A_481_379#_c_603_n N_A_514_424#_c_841_n 4.93996e-19 $X=3.08 $Y=1.97
+ $X2=0 $Y2=0
cc_552 N_A_481_379#_c_610_n N_A_514_424#_c_783_n 0.0130347f $X=6.715 $Y=1.845
+ $X2=0 $Y2=0
cc_553 N_A_481_379#_c_598_n N_A_514_424#_c_767_n 0.0170323f $X=6.88 $Y=1.76
+ $X2=0 $Y2=0
cc_554 N_A_481_379#_c_599_n N_A_514_424#_c_767_n 0.0158838f $X=7.34 $Y=1.19
+ $X2=0 $Y2=0
cc_555 N_A_481_379#_c_598_n N_A_849_424#_c_1004_n 0.00127243f $X=6.88 $Y=1.76
+ $X2=0 $Y2=0
cc_556 N_A_481_379#_c_599_n N_A_849_424#_c_1004_n 0.00113702f $X=7.34 $Y=1.19
+ $X2=0 $Y2=0
cc_557 N_A_481_379#_c_600_n N_A_849_424#_c_1004_n 0.00164728f $X=7.34 $Y=0.795
+ $X2=0 $Y2=0
cc_558 N_A_481_379#_c_595_n N_A_849_424#_c_1013_n 0.00326584f $X=4.055 $Y=1.845
+ $X2=0 $Y2=0
cc_559 N_A_481_379#_c_607_n N_A_849_424#_c_1013_n 8.40069e-19 $X=4.17 $Y=2.045
+ $X2=0 $Y2=0
cc_560 N_A_481_379#_c_608_n N_A_849_424#_c_1013_n 0.0166124f $X=5.035 $Y=1.92
+ $X2=0 $Y2=0
cc_561 N_A_481_379#_c_609_n N_A_849_424#_c_1013_n 8.16755e-19 $X=4.26 $Y=1.92
+ $X2=0 $Y2=0
cc_562 N_A_481_379#_c_666_n N_A_849_424#_c_1013_n 0.0240014f $X=5.2 $Y=1.765
+ $X2=0 $Y2=0
cc_563 N_A_481_379#_c_601_n N_A_849_424#_c_1013_n 0.00895272f $X=5.2 $Y=1.765
+ $X2=0 $Y2=0
cc_564 N_A_481_379#_c_608_n N_A_849_424#_c_1037_n 0.0089554f $X=5.035 $Y=1.92
+ $X2=0 $Y2=0
cc_565 N_A_481_379#_c_666_n N_A_849_424#_c_1037_n 0.00848015f $X=5.2 $Y=1.765
+ $X2=0 $Y2=0
cc_566 N_A_481_379#_c_596_n N_A_849_424#_c_1014_n 0.0106363f $X=5.2 $Y=1.42
+ $X2=0 $Y2=0
cc_567 N_A_481_379#_c_610_n N_A_849_424#_c_1014_n 0.00808891f $X=6.715 $Y=1.845
+ $X2=0 $Y2=0
cc_568 N_A_481_379#_c_666_n N_A_849_424#_c_1014_n 0.0185209f $X=5.2 $Y=1.765
+ $X2=0 $Y2=0
cc_569 N_A_481_379#_c_601_n N_A_849_424#_c_1014_n 0.00413681f $X=5.2 $Y=1.765
+ $X2=0 $Y2=0
cc_570 N_A_481_379#_c_610_n N_A_849_424#_c_1015_n 0.0455979f $X=6.715 $Y=1.845
+ $X2=0 $Y2=0
cc_571 N_A_481_379#_c_598_n N_A_849_424#_c_1015_n 0.0131711f $X=6.88 $Y=1.76
+ $X2=0 $Y2=0
cc_572 N_A_481_379#_c_599_n N_A_849_424#_c_1016_n 0.0128646f $X=7.34 $Y=1.19
+ $X2=0 $Y2=0
cc_573 N_A_481_379#_c_600_n N_A_849_424#_c_1016_n 0.00469766f $X=7.34 $Y=0.795
+ $X2=0 $Y2=0
cc_574 N_A_481_379#_c_599_n N_A_849_424#_c_1017_n 0.0224706f $X=7.34 $Y=1.19
+ $X2=0 $Y2=0
cc_575 N_A_481_379#_M1033_d N_A_849_424#_c_1019_n 0.00243149f $X=7.2 $Y=0.37
+ $X2=0 $Y2=0
cc_576 N_A_481_379#_c_600_n N_A_849_424#_c_1019_n 0.0148603f $X=7.34 $Y=0.795
+ $X2=0 $Y2=0
cc_577 N_A_481_379#_c_598_n N_A_849_424#_c_1021_n 0.00880904f $X=6.88 $Y=1.76
+ $X2=0 $Y2=0
cc_578 N_A_481_379#_c_596_n N_A_849_424#_c_1023_n 0.00482183f $X=5.2 $Y=1.42
+ $X2=0 $Y2=0
cc_579 N_A_481_379#_c_597_n N_A_849_424#_c_1023_n 0.00644187f $X=5.2 $Y=1.255
+ $X2=0 $Y2=0
cc_580 N_A_481_379#_c_601_n N_A_849_424#_c_1023_n 0.00173932f $X=5.2 $Y=1.765
+ $X2=0 $Y2=0
cc_581 N_A_481_379#_c_607_n N_A_849_424#_c_1039_n 0.0049342f $X=4.17 $Y=2.045
+ $X2=0 $Y2=0
cc_582 N_A_481_379#_c_608_n N_A_849_424#_c_1039_n 0.016117f $X=5.035 $Y=1.92
+ $X2=0 $Y2=0
cc_583 N_A_481_379#_c_596_n N_A_849_424#_c_1024_n 2.7088e-19 $X=5.2 $Y=1.42
+ $X2=0 $Y2=0
cc_584 N_A_481_379#_c_610_n N_A_849_424#_c_1024_n 0.0100923f $X=6.715 $Y=1.845
+ $X2=0 $Y2=0
cc_585 N_A_481_379#_c_601_n N_A_849_424#_c_1024_n 0.00126796f $X=5.2 $Y=1.765
+ $X2=0 $Y2=0
cc_586 N_A_481_379#_c_599_n N_A_849_424#_c_1025_n 0.0141654f $X=7.34 $Y=1.19
+ $X2=0 $Y2=0
cc_587 N_A_481_379#_c_600_n N_A_849_424#_c_1025_n 0.0119023f $X=7.34 $Y=0.795
+ $X2=0 $Y2=0
cc_588 N_A_481_379#_c_610_n N_VPWR_M1000_s 0.00285282f $X=6.715 $Y=1.845 $X2=0
+ $Y2=0
cc_589 N_A_481_379#_c_602_n N_VPWR_c_1637_n 0.00280451f $X=2.495 $Y=2.045 $X2=0
+ $Y2=0
cc_590 N_A_481_379#_c_607_n N_VPWR_c_1637_n 0.00280451f $X=4.17 $Y=2.045 $X2=0
+ $Y2=0
cc_591 N_A_481_379#_c_602_n N_VPWR_c_1627_n 0.00359472f $X=2.495 $Y=2.045 $X2=0
+ $Y2=0
cc_592 N_A_481_379#_c_607_n N_VPWR_c_1627_n 0.00360251f $X=4.17 $Y=2.045 $X2=0
+ $Y2=0
cc_593 N_A_481_379#_c_607_n N_A_114_368#_c_1798_n 0.00792562f $X=4.17 $Y=2.045
+ $X2=0 $Y2=0
cc_594 N_A_481_379#_c_593_n N_A_114_368#_c_1759_n 0.00999031f $X=3.98 $Y=1.315
+ $X2=0 $Y2=0
cc_595 N_A_481_379#_c_595_n N_A_114_368#_c_1759_n 0.00111199f $X=4.055 $Y=1.845
+ $X2=0 $Y2=0
cc_596 N_A_481_379#_c_609_n N_A_114_368#_c_1759_n 4.8939e-19 $X=4.26 $Y=1.92
+ $X2=0 $Y2=0
cc_597 N_A_481_379#_c_595_n N_A_114_368#_c_1760_n 0.0145744f $X=4.055 $Y=1.845
+ $X2=0 $Y2=0
cc_598 N_A_481_379#_c_607_n N_A_114_368#_c_1760_n 0.00235568f $X=4.17 $Y=2.045
+ $X2=0 $Y2=0
cc_599 N_A_481_379#_c_609_n N_A_114_368#_c_1760_n 0.0106814f $X=4.26 $Y=1.92
+ $X2=0 $Y2=0
cc_600 N_A_481_379#_c_603_n N_A_114_368#_c_1761_n 0.00295089f $X=3.08 $Y=1.97
+ $X2=0 $Y2=0
cc_601 N_A_481_379#_c_604_n N_A_114_368#_c_1761_n 0.00303128f $X=2.57 $Y=1.97
+ $X2=0 $Y2=0
cc_602 N_A_481_379#_c_592_n N_A_114_368#_c_1761_n 0.00221413f $X=3.445 $Y=1.24
+ $X2=0 $Y2=0
cc_603 N_A_481_379#_c_593_n N_A_114_368#_c_1761_n 0.00869602f $X=3.98 $Y=1.315
+ $X2=0 $Y2=0
cc_604 N_A_481_379#_c_594_n N_A_114_368#_c_1761_n 0.0102793f $X=3.52 $Y=1.315
+ $X2=0 $Y2=0
cc_605 N_A_481_379#_c_593_n N_A_114_368#_c_1763_n 2.92053e-19 $X=3.98 $Y=1.315
+ $X2=0 $Y2=0
cc_606 N_A_481_379#_c_595_n N_A_114_368#_c_1763_n 8.60471e-19 $X=4.055 $Y=1.845
+ $X2=0 $Y2=0
cc_607 N_A_481_379#_c_602_n N_A_413_392#_c_1864_n 0.0047955f $X=2.495 $Y=2.045
+ $X2=0 $Y2=0
cc_608 N_A_481_379#_c_602_n N_A_413_392#_c_1865_n 0.0158167f $X=2.495 $Y=2.045
+ $X2=0 $Y2=0
cc_609 N_A_481_379#_c_607_n N_A_413_392#_c_1865_n 0.012141f $X=4.17 $Y=2.045
+ $X2=0 $Y2=0
cc_610 N_A_481_379#_c_592_n N_A_413_392#_c_1859_n 0.00629471f $X=3.445 $Y=1.24
+ $X2=0 $Y2=0
cc_611 N_A_481_379#_c_597_n N_A_413_392#_c_1859_n 0.00617956f $X=5.2 $Y=1.255
+ $X2=0 $Y2=0
cc_612 N_A_481_379#_c_604_n N_A_413_392#_c_1861_n 0.00160997f $X=2.57 $Y=1.97
+ $X2=0 $Y2=0
cc_613 N_A_481_379#_c_597_n N_A_413_392#_c_1863_n 0.00696738f $X=5.2 $Y=1.255
+ $X2=0 $Y2=0
cc_614 N_A_481_379#_c_592_n N_VGND_c_2056_n 6.67145e-19 $X=3.445 $Y=1.24 $X2=0
+ $Y2=0
cc_615 N_A_481_379#_c_597_n N_VGND_c_2056_n 6.67145e-19 $X=5.2 $Y=1.255 $X2=0
+ $Y2=0
cc_616 N_A_514_424#_c_802_n N_A_849_424#_M1016_d 0.0351341f $X=5.385 $Y=2.635
+ $X2=0 $Y2=0
cc_617 N_A_514_424#_c_846_p N_A_849_424#_M1016_d 0.00951037f $X=5.47 $Y=2.55
+ $X2=0 $Y2=0
cc_618 N_A_514_424#_c_776_n N_A_849_424#_M1016_d 0.0018675f $X=5.555 $Y=2.185
+ $X2=0 $Y2=0
cc_619 N_A_514_424#_M1020_g N_A_849_424#_c_1004_n 0.00114732f $X=8.625 $Y=0.715
+ $X2=0 $Y2=0
cc_620 N_A_514_424#_c_764_n N_A_849_424#_c_1004_n 0.00825234f $X=8.575 $Y=1.39
+ $X2=0 $Y2=0
cc_621 N_A_514_424#_c_778_n N_A_849_424#_c_1028_n 0.0173779f $X=8.48 $Y=2.99
+ $X2=0 $Y2=0
cc_622 N_A_514_424#_c_763_n N_A_849_424#_c_1028_n 0.0170565f $X=8.575 $Y=1.39
+ $X2=0 $Y2=0
cc_623 N_A_514_424#_c_763_n N_A_849_424#_c_1029_n 0.0163487f $X=8.575 $Y=1.39
+ $X2=0 $Y2=0
cc_624 N_A_514_424#_c_768_n N_A_849_424#_c_1029_n 0.0032852f $X=9.475 $Y=1.795
+ $X2=0 $Y2=0
cc_625 N_A_514_424#_c_760_n N_A_849_424#_c_1005_n 0.0196021f $X=9.4 $Y=2.045
+ $X2=0 $Y2=0
cc_626 N_A_514_424#_c_763_n N_A_849_424#_c_1005_n 0.00155904f $X=8.575 $Y=1.39
+ $X2=0 $Y2=0
cc_627 N_A_514_424#_c_769_n N_A_849_424#_c_1005_n 0.0032852f $X=9.41 $Y=1.63
+ $X2=0 $Y2=0
cc_628 N_A_514_424#_c_760_n N_A_849_424#_c_1006_n 0.0183232f $X=9.4 $Y=2.045
+ $X2=0 $Y2=0
cc_629 N_A_514_424#_c_769_n N_A_849_424#_c_1006_n 0.00914562f $X=9.41 $Y=1.63
+ $X2=0 $Y2=0
cc_630 N_A_514_424#_c_763_n N_A_849_424#_c_1007_n 3.57214e-19 $X=8.575 $Y=1.39
+ $X2=0 $Y2=0
cc_631 N_A_514_424#_c_764_n N_A_849_424#_c_1007_n 0.0196409f $X=8.575 $Y=1.39
+ $X2=0 $Y2=0
cc_632 N_A_514_424#_M1020_g N_A_849_424#_M1009_g 0.00954663f $X=8.625 $Y=0.715
+ $X2=0 $Y2=0
cc_633 N_A_514_424#_M1027_g N_A_849_424#_M1009_g 0.0123738f $X=10.285 $Y=0.715
+ $X2=0 $Y2=0
cc_634 N_A_514_424#_c_863_p N_A_849_424#_M1009_g 0.00838117f $X=10.085 $Y=0.68
+ $X2=0 $Y2=0
cc_635 N_A_514_424#_c_864_p N_A_849_424#_M1009_g 0.00334854f $X=9.415 $Y=0.68
+ $X2=0 $Y2=0
cc_636 N_A_514_424#_c_765_n N_A_849_424#_M1009_g 0.00131475f $X=10.17 $Y=1.355
+ $X2=0 $Y2=0
cc_637 N_A_514_424#_c_769_n N_A_849_424#_M1009_g 0.0131456f $X=9.41 $Y=1.63
+ $X2=0 $Y2=0
cc_638 N_A_514_424#_M1027_g N_A_849_424#_c_1009_n 0.0135199f $X=10.285 $Y=0.715
+ $X2=0 $Y2=0
cc_639 N_A_514_424#_c_863_p N_A_849_424#_c_1009_n 0.0040736f $X=10.085 $Y=0.68
+ $X2=0 $Y2=0
cc_640 N_A_514_424#_c_765_n N_A_849_424#_c_1009_n 8.02492e-19 $X=10.17 $Y=1.355
+ $X2=0 $Y2=0
cc_641 N_A_514_424#_c_770_n N_A_849_424#_c_1009_n 0.0020763f $X=10.375 $Y=1.52
+ $X2=0 $Y2=0
cc_642 N_A_514_424#_c_760_n N_A_849_424#_c_1010_n 0.0203607f $X=9.4 $Y=2.045
+ $X2=0 $Y2=0
cc_643 N_A_514_424#_c_768_n N_A_849_424#_c_1010_n 3.04548e-19 $X=9.475 $Y=1.795
+ $X2=0 $Y2=0
cc_644 N_A_514_424#_c_769_n N_A_849_424#_c_1010_n 0.00121181f $X=9.41 $Y=1.63
+ $X2=0 $Y2=0
cc_645 N_A_514_424#_c_771_n N_A_849_424#_c_1010_n 0.0135199f $X=10.375 $Y=1.52
+ $X2=0 $Y2=0
cc_646 N_A_514_424#_c_760_n N_A_849_424#_c_1032_n 0.0118269f $X=9.4 $Y=2.045
+ $X2=0 $Y2=0
cc_647 N_A_514_424#_c_781_n N_A_849_424#_c_1032_n 0.00202457f $X=9.405 $Y=2.99
+ $X2=0 $Y2=0
cc_648 N_A_514_424#_c_758_n N_A_849_424#_c_1011_n 0.0200325f $X=7.18 $Y=2.045
+ $X2=0 $Y2=0
cc_649 N_A_514_424#_c_767_n N_A_849_424#_c_1011_n 3.61457e-19 $X=7.34 $Y=1.795
+ $X2=0 $Y2=0
cc_650 N_A_514_424#_c_763_n N_A_849_424#_c_1034_n 0.00240428f $X=8.575 $Y=1.39
+ $X2=0 $Y2=0
cc_651 N_A_514_424#_c_764_n N_A_849_424#_c_1034_n 0.0189549f $X=8.575 $Y=1.39
+ $X2=0 $Y2=0
cc_652 N_A_514_424#_c_768_n N_A_849_424#_c_1012_n 0.00114375f $X=9.475 $Y=1.795
+ $X2=0 $Y2=0
cc_653 N_A_514_424#_c_769_n N_A_849_424#_c_1012_n 0.00376165f $X=9.41 $Y=1.63
+ $X2=0 $Y2=0
cc_654 N_A_514_424#_c_760_n N_A_849_424#_c_1035_n 0.00275525f $X=9.4 $Y=2.045
+ $X2=0 $Y2=0
cc_655 N_A_514_424#_c_782_n N_A_849_424#_c_1035_n 2.19183e-19 $X=9.49 $Y=2.905
+ $X2=0 $Y2=0
cc_656 N_A_514_424#_c_770_n N_A_849_424#_c_1035_n 0.00562228f $X=10.375 $Y=1.52
+ $X2=0 $Y2=0
cc_657 N_A_514_424#_c_771_n N_A_849_424#_c_1035_n 0.00483728f $X=10.375 $Y=1.52
+ $X2=0 $Y2=0
cc_658 N_A_514_424#_c_802_n N_A_849_424#_c_1037_n 0.0185318f $X=5.385 $Y=2.635
+ $X2=0 $Y2=0
cc_659 N_A_514_424#_c_846_p N_A_849_424#_c_1037_n 0.00639084f $X=5.47 $Y=2.55
+ $X2=0 $Y2=0
cc_660 N_A_514_424#_c_776_n N_A_849_424#_c_1037_n 0.0153044f $X=5.555 $Y=2.185
+ $X2=0 $Y2=0
cc_661 N_A_514_424#_c_758_n N_A_849_424#_c_1022_n 0.00180662f $X=7.18 $Y=2.045
+ $X2=0 $Y2=0
cc_662 N_A_514_424#_c_767_n N_A_849_424#_c_1022_n 0.0244767f $X=7.34 $Y=1.795
+ $X2=0 $Y2=0
cc_663 N_A_514_424#_c_802_n N_A_849_424#_c_1039_n 0.042919f $X=5.385 $Y=2.635
+ $X2=0 $Y2=0
cc_664 N_A_514_424#_c_864_p N_A_1689_424#_M1020_d 0.00252339f $X=9.415 $Y=0.68
+ $X2=-0.19 $Y2=-0.245
cc_665 N_A_514_424#_c_769_n N_A_1689_424#_M1020_d 0.00190212f $X=9.41 $Y=1.63
+ $X2=-0.19 $Y2=-0.245
cc_666 N_A_514_424#_c_763_n N_A_1689_424#_M1004_d 0.0177243f $X=8.575 $Y=1.39
+ $X2=0 $Y2=0
cc_667 N_A_514_424#_c_781_n N_A_1689_424#_M1004_d 0.0124929f $X=9.405 $Y=2.99
+ $X2=0 $Y2=0
cc_668 N_A_514_424#_c_785_n N_A_1689_424#_M1004_d 3.34869e-19 $X=8.607 $Y=2.99
+ $X2=0 $Y2=0
cc_669 N_A_514_424#_M1027_g N_A_1689_424#_M1011_g 0.0220276f $X=10.285 $Y=0.715
+ $X2=0 $Y2=0
cc_670 N_A_514_424#_c_765_n N_A_1689_424#_M1011_g 3.49739e-19 $X=10.17 $Y=1.355
+ $X2=0 $Y2=0
cc_671 N_A_514_424#_c_770_n N_A_1689_424#_M1011_g 2.87872e-19 $X=10.375 $Y=1.52
+ $X2=0 $Y2=0
cc_672 N_A_514_424#_c_771_n N_A_1689_424#_M1011_g 0.0171809f $X=10.375 $Y=1.52
+ $X2=0 $Y2=0
cc_673 N_A_514_424#_M1020_g N_A_1689_424#_c_1234_n 0.00572966f $X=8.625 $Y=0.715
+ $X2=0 $Y2=0
cc_674 N_A_514_424#_c_864_p N_A_1689_424#_c_1234_n 0.0144778f $X=9.415 $Y=0.68
+ $X2=0 $Y2=0
cc_675 N_A_514_424#_c_769_n N_A_1689_424#_c_1234_n 0.0436224f $X=9.41 $Y=1.63
+ $X2=0 $Y2=0
cc_676 N_A_514_424#_M1027_g N_A_1689_424#_c_1215_n 0.0128606f $X=10.285 $Y=0.715
+ $X2=0 $Y2=0
cc_677 N_A_514_424#_c_863_p N_A_1689_424#_c_1215_n 0.047342f $X=10.085 $Y=0.68
+ $X2=0 $Y2=0
cc_678 N_A_514_424#_c_864_p N_A_1689_424#_c_1215_n 0.00806988f $X=9.415 $Y=0.68
+ $X2=0 $Y2=0
cc_679 N_A_514_424#_M1020_g N_A_1689_424#_c_1216_n 0.00490006f $X=8.625 $Y=0.715
+ $X2=0 $Y2=0
cc_680 N_A_514_424#_c_768_n N_A_1689_424#_c_1218_n 0.0436224f $X=9.475 $Y=1.795
+ $X2=0 $Y2=0
cc_681 N_A_514_424#_c_760_n N_A_1689_424#_c_1242_n 0.0129686f $X=9.4 $Y=2.045
+ $X2=0 $Y2=0
cc_682 N_A_514_424#_c_781_n N_A_1689_424#_c_1242_n 0.0248568f $X=9.405 $Y=2.99
+ $X2=0 $Y2=0
cc_683 N_A_514_424#_c_782_n N_A_1689_424#_c_1242_n 0.0447254f $X=9.49 $Y=2.905
+ $X2=0 $Y2=0
cc_684 N_A_514_424#_M1020_g N_A_1689_424#_c_1219_n 0.0021401f $X=8.625 $Y=0.715
+ $X2=0 $Y2=0
cc_685 N_A_514_424#_c_760_n N_A_1689_424#_c_1219_n 0.00370778f $X=9.4 $Y=2.045
+ $X2=0 $Y2=0
cc_686 N_A_514_424#_c_763_n N_A_1689_424#_c_1219_n 0.115338f $X=8.575 $Y=1.39
+ $X2=0 $Y2=0
cc_687 N_A_514_424#_c_764_n N_A_1689_424#_c_1219_n 0.00183199f $X=8.575 $Y=1.39
+ $X2=0 $Y2=0
cc_688 N_A_514_424#_c_782_n N_A_1689_424#_c_1219_n 0.0073481f $X=9.49 $Y=2.905
+ $X2=0 $Y2=0
cc_689 N_A_514_424#_c_777_n N_A_1451_424#_M1012_d 0.00156777f $X=7.3 $Y=2.24
+ $X2=0 $Y2=0
cc_690 N_A_514_424#_c_809_n N_A_1451_424#_M1012_d 0.00992f $X=7.3 $Y=2.905 $X2=0
+ $Y2=0
cc_691 N_A_514_424#_c_778_n N_A_1451_424#_M1012_d 0.0157589f $X=8.48 $Y=2.99
+ $X2=0 $Y2=0
cc_692 N_A_514_424#_c_921_p N_A_1451_424#_M1012_d 0.00188126f $X=7.3 $Y=2.325
+ $X2=0 $Y2=0
cc_693 N_A_514_424#_M1020_g N_A_1451_424#_c_1376_n 0.0132473f $X=8.625 $Y=0.715
+ $X2=0 $Y2=0
cc_694 N_A_514_424#_c_763_n N_A_1451_424#_c_1376_n 0.00492931f $X=8.575 $Y=1.39
+ $X2=0 $Y2=0
cc_695 N_A_514_424#_c_764_n N_A_1451_424#_c_1376_n 0.00300137f $X=8.575 $Y=1.39
+ $X2=0 $Y2=0
cc_696 N_A_514_424#_c_758_n N_A_1451_424#_c_1377_n 0.00378564f $X=7.18 $Y=2.045
+ $X2=0 $Y2=0
cc_697 N_A_514_424#_M1020_g N_A_1451_424#_c_1377_n 0.00283903f $X=8.625 $Y=0.715
+ $X2=0 $Y2=0
cc_698 N_A_514_424#_c_777_n N_A_1451_424#_c_1377_n 0.00883155f $X=7.3 $Y=2.24
+ $X2=0 $Y2=0
cc_699 N_A_514_424#_c_809_n N_A_1451_424#_c_1377_n 0.0263235f $X=7.3 $Y=2.905
+ $X2=0 $Y2=0
cc_700 N_A_514_424#_c_778_n N_A_1451_424#_c_1377_n 0.0522285f $X=8.48 $Y=2.99
+ $X2=0 $Y2=0
cc_701 N_A_514_424#_c_763_n N_A_1451_424#_c_1377_n 0.0666571f $X=8.575 $Y=1.39
+ $X2=0 $Y2=0
cc_702 N_A_514_424#_c_764_n N_A_1451_424#_c_1377_n 0.00285755f $X=8.575 $Y=1.39
+ $X2=0 $Y2=0
cc_703 N_A_514_424#_c_767_n N_A_1451_424#_c_1377_n 4.09734e-19 $X=7.34 $Y=1.795
+ $X2=0 $Y2=0
cc_704 N_A_514_424#_c_921_p N_A_1451_424#_c_1377_n 0.0153274f $X=7.3 $Y=2.325
+ $X2=0 $Y2=0
cc_705 N_A_514_424#_M1020_g N_A_1451_424#_c_1378_n 0.00897056f $X=8.625 $Y=0.715
+ $X2=0 $Y2=0
cc_706 N_A_514_424#_M1027_g N_A_1451_424#_c_1378_n 0.00246693f $X=10.285
+ $Y=0.715 $X2=0 $Y2=0
cc_707 N_A_514_424#_c_763_n N_A_1451_424#_c_1378_n 0.00769204f $X=8.575 $Y=1.39
+ $X2=0 $Y2=0
cc_708 N_A_514_424#_c_863_p N_A_1451_424#_c_1378_n 0.0249927f $X=10.085 $Y=0.68
+ $X2=0 $Y2=0
cc_709 N_A_514_424#_c_765_n N_A_1451_424#_c_1378_n 0.0116545f $X=10.17 $Y=1.355
+ $X2=0 $Y2=0
cc_710 N_A_514_424#_c_769_n N_A_1451_424#_c_1378_n 0.0136154f $X=9.41 $Y=1.63
+ $X2=0 $Y2=0
cc_711 N_A_514_424#_c_770_n N_A_1451_424#_c_1378_n 0.00635749f $X=10.375 $Y=1.52
+ $X2=0 $Y2=0
cc_712 N_A_514_424#_c_771_n N_A_1451_424#_c_1378_n 0.00140296f $X=10.375 $Y=1.52
+ $X2=0 $Y2=0
cc_713 N_A_514_424#_c_763_n N_A_1451_424#_c_1379_n 5.09649e-19 $X=8.575 $Y=1.39
+ $X2=0 $Y2=0
cc_714 N_A_514_424#_c_863_p N_A_1895_424#_M1009_d 0.0129049f $X=10.085 $Y=0.68
+ $X2=-0.19 $Y2=-0.245
cc_715 N_A_514_424#_c_765_n N_A_1895_424#_M1009_d 0.00322197f $X=10.17 $Y=1.355
+ $X2=-0.19 $Y2=-0.245
cc_716 N_A_514_424#_c_781_n N_A_1895_424#_M1031_d 5.4799e-19 $X=9.405 $Y=2.99
+ $X2=0 $Y2=0
cc_717 N_A_514_424#_c_782_n N_A_1895_424#_M1031_d 0.0075045f $X=9.49 $Y=2.905
+ $X2=0 $Y2=0
cc_718 N_A_514_424#_c_782_n N_A_1895_424#_c_1524_n 0.0483622f $X=9.49 $Y=2.905
+ $X2=0 $Y2=0
cc_719 N_A_514_424#_M1027_g N_A_1895_424#_c_1507_n 9.60195e-19 $X=10.285
+ $Y=0.715 $X2=0 $Y2=0
cc_720 N_A_514_424#_c_863_p N_A_1895_424#_c_1507_n 0.0209502f $X=10.085 $Y=0.68
+ $X2=0 $Y2=0
cc_721 N_A_514_424#_c_765_n N_A_1895_424#_c_1507_n 0.0314353f $X=10.17 $Y=1.355
+ $X2=0 $Y2=0
cc_722 N_A_514_424#_c_769_n N_A_1895_424#_c_1507_n 0.0156657f $X=9.41 $Y=1.63
+ $X2=0 $Y2=0
cc_723 N_A_514_424#_c_760_n N_A_1895_424#_c_1508_n 0.00543807f $X=9.4 $Y=2.045
+ $X2=0 $Y2=0
cc_724 N_A_514_424#_c_768_n N_A_1895_424#_c_1508_n 0.0483622f $X=9.475 $Y=1.795
+ $X2=0 $Y2=0
cc_725 N_A_514_424#_c_769_n N_A_1895_424#_c_1508_n 0.0197285f $X=9.41 $Y=1.63
+ $X2=0 $Y2=0
cc_726 N_A_514_424#_c_770_n N_A_1895_424#_c_1508_n 0.0251734f $X=10.375 $Y=1.52
+ $X2=0 $Y2=0
cc_727 N_A_514_424#_c_771_n N_A_1895_424#_c_1508_n 2.83052e-19 $X=10.375 $Y=1.52
+ $X2=0 $Y2=0
cc_728 N_A_514_424#_c_781_n N_A_1895_424#_c_1517_n 0.00645303f $X=9.405 $Y=2.99
+ $X2=0 $Y2=0
cc_729 N_A_514_424#_c_806_n N_VPWR_M1000_s 0.00349181f $X=7.215 $Y=2.325 $X2=0
+ $Y2=0
cc_730 N_A_514_424#_c_783_n N_VPWR_M1000_s 0.00572595f $X=6.31 $Y=2.185 $X2=0
+ $Y2=0
cc_731 N_A_514_424#_c_758_n N_VPWR_c_1631_n 0.00158305f $X=7.18 $Y=2.045 $X2=0
+ $Y2=0
cc_732 N_A_514_424#_c_806_n N_VPWR_c_1631_n 0.0114382f $X=7.215 $Y=2.325 $X2=0
+ $Y2=0
cc_733 N_A_514_424#_c_809_n N_VPWR_c_1631_n 0.0079191f $X=7.3 $Y=2.905 $X2=0
+ $Y2=0
cc_734 N_A_514_424#_c_779_n N_VPWR_c_1631_n 0.00462202f $X=7.385 $Y=2.99 $X2=0
+ $Y2=0
cc_735 N_A_514_424#_c_783_n N_VPWR_c_1631_n 0.0110011f $X=6.31 $Y=2.185 $X2=0
+ $Y2=0
cc_736 N_A_514_424#_c_758_n N_VPWR_c_1638_n 0.00412574f $X=7.18 $Y=2.045 $X2=0
+ $Y2=0
cc_737 N_A_514_424#_c_760_n N_VPWR_c_1638_n 0.00278203f $X=9.4 $Y=2.045 $X2=0
+ $Y2=0
cc_738 N_A_514_424#_c_778_n N_VPWR_c_1638_n 0.0700431f $X=8.48 $Y=2.99 $X2=0
+ $Y2=0
cc_739 N_A_514_424#_c_779_n N_VPWR_c_1638_n 0.0120135f $X=7.385 $Y=2.99 $X2=0
+ $Y2=0
cc_740 N_A_514_424#_c_781_n N_VPWR_c_1638_n 0.0547801f $X=9.405 $Y=2.99 $X2=0
+ $Y2=0
cc_741 N_A_514_424#_c_785_n N_VPWR_c_1638_n 0.0182077f $X=8.607 $Y=2.99 $X2=0
+ $Y2=0
cc_742 N_A_514_424#_c_758_n N_VPWR_c_1627_n 0.00766989f $X=7.18 $Y=2.045 $X2=0
+ $Y2=0
cc_743 N_A_514_424#_c_760_n N_VPWR_c_1627_n 0.00360963f $X=9.4 $Y=2.045 $X2=0
+ $Y2=0
cc_744 N_A_514_424#_c_778_n N_VPWR_c_1627_n 0.040479f $X=8.48 $Y=2.99 $X2=0
+ $Y2=0
cc_745 N_A_514_424#_c_779_n N_VPWR_c_1627_n 0.00642149f $X=7.385 $Y=2.99 $X2=0
+ $Y2=0
cc_746 N_A_514_424#_c_781_n N_VPWR_c_1627_n 0.0311032f $X=9.405 $Y=2.99 $X2=0
+ $Y2=0
cc_747 N_A_514_424#_c_785_n N_VPWR_c_1627_n 0.00990325f $X=8.607 $Y=2.99 $X2=0
+ $Y2=0
cc_748 N_A_514_424#_c_802_n N_A_114_368#_M1010_d 0.00799774f $X=5.385 $Y=2.635
+ $X2=0 $Y2=0
cc_749 N_A_514_424#_c_762_n N_A_114_368#_c_1798_n 0.010078f $X=3.15 $Y=2.39
+ $X2=0 $Y2=0
cc_750 N_A_514_424#_c_802_n N_A_114_368#_c_1798_n 0.0285867f $X=5.385 $Y=2.635
+ $X2=0 $Y2=0
cc_751 N_A_514_424#_c_762_n N_A_114_368#_c_1761_n 0.0176866f $X=3.15 $Y=2.39
+ $X2=0 $Y2=0
cc_752 N_A_514_424#_c_766_n N_A_114_368#_c_1761_n 0.00841417f $X=3.23 $Y=1.02
+ $X2=0 $Y2=0
cc_753 N_A_514_424#_c_775_n N_A_413_392#_M1024_d 0.00328964f $X=6.225 $Y=2.185
+ $X2=0 $Y2=0
cc_754 N_A_514_424#_M1003_d N_A_413_392#_c_1865_n 0.0106552f $X=2.57 $Y=2.12
+ $X2=0 $Y2=0
cc_755 N_A_514_424#_c_796_n N_A_413_392#_c_1865_n 0.175584f $X=3.065 $Y=2.555
+ $X2=0 $Y2=0
cc_756 N_A_514_424#_c_802_n N_A_413_392#_c_1865_n 0.0112207f $X=5.385 $Y=2.635
+ $X2=0 $Y2=0
cc_757 N_A_514_424#_c_775_n N_A_413_392#_c_1865_n 0.00311653f $X=6.225 $Y=2.185
+ $X2=0 $Y2=0
cc_758 N_A_514_424#_c_775_n N_A_413_392#_c_1867_n 0.0218579f $X=6.225 $Y=2.185
+ $X2=0 $Y2=0
cc_759 N_A_514_424#_c_770_n N_A_2052_424#_c_1949_n 0.00572806f $X=10.375 $Y=1.52
+ $X2=0 $Y2=0
cc_760 N_A_514_424#_c_771_n N_A_2052_424#_c_1949_n 0.00521158f $X=10.375 $Y=1.52
+ $X2=0 $Y2=0
cc_761 N_A_514_424#_M1027_g N_A_2052_424#_c_1951_n 0.00128506f $X=10.285
+ $Y=0.715 $X2=0 $Y2=0
cc_762 N_A_514_424#_c_863_p N_A_2052_424#_c_1951_n 0.0133617f $X=10.085 $Y=0.68
+ $X2=0 $Y2=0
cc_763 N_A_514_424#_c_765_n N_A_2052_424#_c_1951_n 0.0170539f $X=10.17 $Y=1.355
+ $X2=0 $Y2=0
cc_764 N_A_514_424#_M1027_g N_A_2052_424#_c_1946_n 0.00128429f $X=10.285
+ $Y=0.715 $X2=0 $Y2=0
cc_765 N_A_514_424#_c_765_n N_A_2052_424#_c_1946_n 0.00659864f $X=10.17 $Y=1.355
+ $X2=0 $Y2=0
cc_766 N_A_514_424#_c_770_n N_A_2052_424#_c_1946_n 0.0250644f $X=10.375 $Y=1.52
+ $X2=0 $Y2=0
cc_767 N_A_514_424#_c_771_n N_A_2052_424#_c_1946_n 0.00218336f $X=10.375 $Y=1.52
+ $X2=0 $Y2=0
cc_768 N_A_514_424#_M1027_g N_A_2052_424#_c_1947_n 0.00150913f $X=10.285
+ $Y=0.715 $X2=0 $Y2=0
cc_769 N_A_514_424#_c_765_n N_A_2052_424#_c_1947_n 0.0128814f $X=10.17 $Y=1.355
+ $X2=0 $Y2=0
cc_770 N_A_514_424#_c_770_n N_A_2052_424#_c_1947_n 0.00318906f $X=10.375 $Y=1.52
+ $X2=0 $Y2=0
cc_771 N_A_514_424#_c_771_n N_A_2052_424#_c_1947_n 0.00363856f $X=10.375 $Y=1.52
+ $X2=0 $Y2=0
cc_772 N_A_514_424#_M1020_g N_VGND_c_2054_n 0.0055442f $X=8.625 $Y=0.715 $X2=0
+ $Y2=0
cc_773 N_A_514_424#_M1027_g N_VGND_c_2054_n 9.44495e-19 $X=10.285 $Y=0.715 $X2=0
+ $Y2=0
cc_774 N_A_514_424#_M1020_g N_VGND_c_2063_n 0.00537853f $X=8.625 $Y=0.715 $X2=0
+ $Y2=0
cc_775 N_A_849_424#_c_1032_n N_A_1689_424#_c_1214_n 0.0225262f $X=10.185
+ $Y=2.045 $X2=0 $Y2=0
cc_776 N_A_849_424#_c_1035_n N_A_1689_424#_c_1214_n 0.00275774f $X=10.185
+ $Y=1.97 $X2=0 $Y2=0
cc_777 N_A_849_424#_M1009_g N_A_1689_424#_c_1234_n 0.00584701f $X=9.455 $Y=0.715
+ $X2=0 $Y2=0
cc_778 N_A_849_424#_M1009_g N_A_1689_424#_c_1215_n 0.0128029f $X=9.455 $Y=0.715
+ $X2=0 $Y2=0
cc_779 N_A_849_424#_c_1029_n N_A_1689_424#_c_1242_n 0.0011642f $X=8.95 $Y=1.87
+ $X2=0 $Y2=0
cc_780 N_A_849_424#_c_1029_n N_A_1689_424#_c_1219_n 0.00936187f $X=8.95 $Y=1.87
+ $X2=0 $Y2=0
cc_781 N_A_849_424#_c_1005_n N_A_1689_424#_c_1219_n 0.0108539f $X=9.025 $Y=1.795
+ $X2=0 $Y2=0
cc_782 N_A_849_424#_c_1007_n N_A_1689_424#_c_1219_n 0.00731363f $X=9.1 $Y=1.315
+ $X2=0 $Y2=0
cc_783 N_A_849_424#_c_1019_n N_A_1451_424#_M1019_d 3.31987e-19 $X=7.675 $Y=0.34
+ $X2=-0.19 $Y2=-0.245
cc_784 N_A_849_424#_c_1025_n N_A_1451_424#_M1019_d 0.00955805f $X=7.822 $Y=1.275
+ $X2=-0.19 $Y2=-0.245
cc_785 N_A_849_424#_c_1004_n N_A_1451_424#_c_1376_n 7.93787e-19 $X=7.6 $Y=1.11
+ $X2=0 $Y2=0
cc_786 N_A_849_424#_c_1019_n N_A_1451_424#_c_1376_n 0.00311987f $X=7.675 $Y=0.34
+ $X2=0 $Y2=0
cc_787 N_A_849_424#_c_1025_n N_A_1451_424#_c_1376_n 0.0365201f $X=7.822 $Y=1.275
+ $X2=0 $Y2=0
cc_788 N_A_849_424#_c_1004_n N_A_1451_424#_c_1377_n 0.00977968f $X=7.6 $Y=1.11
+ $X2=0 $Y2=0
cc_789 N_A_849_424#_c_1026_n N_A_1451_424#_c_1377_n 0.0104179f $X=8.28 $Y=1.87
+ $X2=0 $Y2=0
cc_790 N_A_849_424#_c_1027_n N_A_1451_424#_c_1377_n 0.00985463f $X=8.045 $Y=1.87
+ $X2=0 $Y2=0
cc_791 N_A_849_424#_c_1028_n N_A_1451_424#_c_1377_n 0.00841885f $X=8.37 $Y=2.045
+ $X2=0 $Y2=0
cc_792 N_A_849_424#_c_1034_n N_A_1451_424#_c_1377_n 0.00631569f $X=8.37 $Y=1.87
+ $X2=0 $Y2=0
cc_793 N_A_849_424#_c_1021_n N_A_1451_424#_c_1377_n 0.0492509f $X=7.822 $Y=1.422
+ $X2=0 $Y2=0
cc_794 N_A_849_424#_c_1022_n N_A_1451_424#_c_1377_n 0.0238237f $X=7.88 $Y=1.44
+ $X2=0 $Y2=0
cc_795 N_A_849_424#_c_1025_n N_A_1451_424#_c_1377_n 0.0113824f $X=7.822 $Y=1.275
+ $X2=0 $Y2=0
cc_796 N_A_849_424#_c_1007_n N_A_1451_424#_c_1378_n 0.00420718f $X=9.1 $Y=1.315
+ $X2=0 $Y2=0
cc_797 N_A_849_424#_M1009_g N_A_1451_424#_c_1378_n 0.00473019f $X=9.455 $Y=0.715
+ $X2=0 $Y2=0
cc_798 N_A_849_424#_c_1009_n N_A_1451_424#_c_1378_n 0.003407f $X=9.85 $Y=1.315
+ $X2=0 $Y2=0
cc_799 N_A_849_424#_c_1025_n N_A_1451_424#_c_1379_n 0.00128282f $X=7.822
+ $Y=1.275 $X2=0 $Y2=0
cc_800 N_A_849_424#_c_1032_n N_A_1895_424#_c_1513_n 0.00447051f $X=10.185
+ $Y=2.045 $X2=0 $Y2=0
cc_801 N_A_849_424#_c_1035_n N_A_1895_424#_c_1513_n 0.00811102f $X=10.185
+ $Y=1.97 $X2=0 $Y2=0
cc_802 N_A_849_424#_c_1032_n N_A_1895_424#_c_1537_n 0.0165956f $X=10.185
+ $Y=2.045 $X2=0 $Y2=0
cc_803 N_A_849_424#_M1009_g N_A_1895_424#_c_1507_n 0.00265376f $X=9.455 $Y=0.715
+ $X2=0 $Y2=0
cc_804 N_A_849_424#_c_1009_n N_A_1895_424#_c_1507_n 0.00647484f $X=9.85 $Y=1.315
+ $X2=0 $Y2=0
cc_805 N_A_849_424#_M1009_g N_A_1895_424#_c_1508_n 5.45878e-19 $X=9.455 $Y=0.715
+ $X2=0 $Y2=0
cc_806 N_A_849_424#_c_1009_n N_A_1895_424#_c_1508_n 0.010022f $X=9.85 $Y=1.315
+ $X2=0 $Y2=0
cc_807 N_A_849_424#_c_1010_n N_A_1895_424#_c_1508_n 0.01798f $X=9.925 $Y=1.895
+ $X2=0 $Y2=0
cc_808 N_A_849_424#_c_1032_n N_A_1895_424#_c_1508_n 0.00125413f $X=10.185
+ $Y=2.045 $X2=0 $Y2=0
cc_809 N_A_849_424#_c_1035_n N_A_1895_424#_c_1508_n 0.00956941f $X=10.185
+ $Y=1.97 $X2=0 $Y2=0
cc_810 N_A_849_424#_c_1032_n N_A_1895_424#_c_1517_n 0.0022523f $X=10.185
+ $Y=2.045 $X2=0 $Y2=0
cc_811 N_A_849_424#_c_1028_n N_VPWR_c_1638_n 0.00278271f $X=8.37 $Y=2.045 $X2=0
+ $Y2=0
cc_812 N_A_849_424#_c_1032_n N_VPWR_c_1638_n 0.00317855f $X=10.185 $Y=2.045
+ $X2=0 $Y2=0
cc_813 N_A_849_424#_c_1028_n N_VPWR_c_1627_n 0.00363426f $X=8.37 $Y=2.045 $X2=0
+ $Y2=0
cc_814 N_A_849_424#_c_1032_n N_VPWR_c_1627_n 0.00400689f $X=10.185 $Y=2.045
+ $X2=0 $Y2=0
cc_815 N_A_849_424#_c_1013_n N_A_114_368#_c_1760_n 0.0121213f $X=4.85 $Y=2.1
+ $X2=0 $Y2=0
cc_816 N_A_849_424#_c_1039_n N_A_114_368#_c_1760_n 0.00179258f $X=4.85 $Y=2.225
+ $X2=0 $Y2=0
cc_817 N_A_849_424#_M1016_d N_A_413_392#_c_1865_n 0.0168757f $X=4.245 $Y=2.12
+ $X2=0 $Y2=0
cc_818 N_A_849_424#_c_1009_n N_A_2052_424#_c_1946_n 0.00441523f $X=9.85 $Y=1.315
+ $X2=0 $Y2=0
cc_819 N_A_849_424#_c_1032_n N_A_2052_424#_c_1946_n 0.00122247f $X=10.185
+ $Y=2.045 $X2=0 $Y2=0
cc_820 N_A_849_424#_c_1035_n N_A_2052_424#_c_1946_n 0.00287402f $X=10.185
+ $Y=1.97 $X2=0 $Y2=0
cc_821 N_A_849_424#_c_1017_n N_VGND_M1033_s 0.0041955f $X=6.835 $Y=0.935 $X2=0
+ $Y2=0
cc_822 N_A_849_424#_c_1198_p N_VGND_M1033_s 0.011619f $X=6.92 $Y=0.85 $X2=0
+ $Y2=0
cc_823 N_A_849_424#_c_1020_n N_VGND_M1033_s 7.1669e-19 $X=7.005 $Y=0.34 $X2=0
+ $Y2=0
cc_824 N_A_849_424#_c_1015_n N_VGND_c_2046_n 0.00109758f $X=6.375 $Y=1.44 $X2=0
+ $Y2=0
cc_825 N_A_849_424#_c_1017_n N_VGND_c_2046_n 0.00980311f $X=6.835 $Y=0.935 $X2=0
+ $Y2=0
cc_826 N_A_849_424#_c_1018_n N_VGND_c_2046_n 0.0155508f $X=6.545 $Y=0.935 $X2=0
+ $Y2=0
cc_827 N_A_849_424#_c_1198_p N_VGND_c_2046_n 0.0194818f $X=6.92 $Y=0.85 $X2=0
+ $Y2=0
cc_828 N_A_849_424#_c_1020_n N_VGND_c_2046_n 0.0148568f $X=7.005 $Y=0.34 $X2=0
+ $Y2=0
cc_829 N_A_849_424#_c_1004_n N_VGND_c_2054_n 9.63786e-19 $X=7.6 $Y=1.11 $X2=0
+ $Y2=0
cc_830 N_A_849_424#_M1009_g N_VGND_c_2054_n 9.44495e-19 $X=9.455 $Y=0.715 $X2=0
+ $Y2=0
cc_831 N_A_849_424#_c_1019_n N_VGND_c_2054_n 0.0548521f $X=7.675 $Y=0.34 $X2=0
+ $Y2=0
cc_832 N_A_849_424#_c_1020_n N_VGND_c_2054_n 0.0121867f $X=7.005 $Y=0.34 $X2=0
+ $Y2=0
cc_833 N_A_849_424#_c_1017_n N_VGND_c_2063_n 0.00621699f $X=6.835 $Y=0.935 $X2=0
+ $Y2=0
cc_834 N_A_849_424#_c_1018_n N_VGND_c_2063_n 6.09234e-19 $X=6.545 $Y=0.935 $X2=0
+ $Y2=0
cc_835 N_A_849_424#_c_1019_n N_VGND_c_2063_n 0.0311091f $X=7.675 $Y=0.34 $X2=0
+ $Y2=0
cc_836 N_A_849_424#_c_1020_n N_VGND_c_2063_n 0.00660921f $X=7.005 $Y=0.34 $X2=0
+ $Y2=0
cc_837 N_A_1689_424#_M1011_g N_CI_c_1329_n 0.00294053f $X=10.855 $Y=0.715 $X2=0
+ $Y2=0
cc_838 N_A_1689_424#_c_1217_n N_CI_c_1329_n 0.00449467f $X=11.075 $Y=1.635 $X2=0
+ $Y2=0
cc_839 N_A_1689_424#_c_1214_n N_CI_c_1330_n 0.0480095f $X=10.87 $Y=1.885 $X2=0
+ $Y2=0
cc_840 N_A_1689_424#_c_1217_n N_CI_c_1330_n 0.00409505f $X=11.075 $Y=1.635 $X2=0
+ $Y2=0
cc_841 N_A_1689_424#_c_1223_n N_CI_c_1330_n 0.0175476f $X=11.765 $Y=2.115 $X2=0
+ $Y2=0
cc_842 N_A_1689_424#_c_1220_n N_CI_c_1330_n 0.00369759f $X=11.11 $Y=0.715 $X2=0
+ $Y2=0
cc_843 N_A_1689_424#_M1011_g N_CI_c_1331_n 0.0190679f $X=10.855 $Y=0.715 $X2=0
+ $Y2=0
cc_844 N_A_1689_424#_c_1217_n N_CI_c_1331_n 0.00502896f $X=11.075 $Y=1.635 $X2=0
+ $Y2=0
cc_845 N_A_1689_424#_c_1220_n N_CI_c_1331_n 0.0231962f $X=11.11 $Y=0.715 $X2=0
+ $Y2=0
cc_846 N_A_1689_424#_c_1223_n N_CI_c_1332_n 0.00101041f $X=11.765 $Y=2.115 $X2=0
+ $Y2=0
cc_847 N_A_1689_424#_c_1220_n N_CI_c_1332_n 0.00141778f $X=11.11 $Y=0.715 $X2=0
+ $Y2=0
cc_848 N_A_1689_424#_c_1214_n CI 0.00114593f $X=10.87 $Y=1.885 $X2=0 $Y2=0
cc_849 N_A_1689_424#_c_1217_n CI 0.0209883f $X=11.075 $Y=1.635 $X2=0 $Y2=0
cc_850 N_A_1689_424#_c_1223_n CI 0.0327065f $X=11.765 $Y=2.115 $X2=0 $Y2=0
cc_851 N_A_1689_424#_c_1220_n CI 0.0156641f $X=11.11 $Y=0.715 $X2=0 $Y2=0
cc_852 N_A_1689_424#_c_1223_n N_A_1451_424#_c_1381_n 0.00421136f $X=11.765
+ $Y=2.115 $X2=0 $Y2=0
cc_853 N_A_1689_424#_c_1220_n N_A_1451_424#_c_1372_n 0.00510143f $X=11.11
+ $Y=0.715 $X2=0 $Y2=0
cc_854 N_A_1689_424#_c_1234_n N_A_1451_424#_c_1376_n 0.0237271f $X=8.91 $Y=0.54
+ $X2=0 $Y2=0
cc_855 N_A_1689_424#_c_1216_n N_A_1451_424#_c_1376_n 0.00148f $X=9.075 $Y=0.34
+ $X2=0 $Y2=0
cc_856 N_A_1689_424#_c_1218_n N_A_1451_424#_c_1377_n 5.98371e-19 $X=8.91
+ $Y=1.055 $X2=0 $Y2=0
cc_857 N_A_1689_424#_c_1219_n N_A_1451_424#_c_1377_n 0.0052908f $X=9.07 $Y=2.13
+ $X2=0 $Y2=0
cc_858 N_A_1689_424#_M1020_d N_A_1451_424#_c_1378_n 0.00668865f $X=8.7 $Y=0.395
+ $X2=0 $Y2=0
cc_859 N_A_1689_424#_M1011_g N_A_1451_424#_c_1378_n 0.00953662f $X=10.855
+ $Y=0.715 $X2=0 $Y2=0
cc_860 N_A_1689_424#_c_1214_n N_A_1451_424#_c_1378_n 0.00108239f $X=10.87
+ $Y=1.885 $X2=0 $Y2=0
cc_861 N_A_1689_424#_c_1234_n N_A_1451_424#_c_1378_n 0.0194893f $X=8.91 $Y=0.54
+ $X2=0 $Y2=0
cc_862 N_A_1689_424#_c_1215_n N_A_1451_424#_c_1378_n 0.0185981f $X=10.765
+ $Y=0.34 $X2=0 $Y2=0
cc_863 N_A_1689_424#_c_1218_n N_A_1451_424#_c_1378_n 0.0185795f $X=8.91 $Y=1.055
+ $X2=0 $Y2=0
cc_864 N_A_1689_424#_c_1220_n N_A_1451_424#_c_1378_n 0.0854708f $X=11.11
+ $Y=0.715 $X2=0 $Y2=0
cc_865 N_A_1689_424#_c_1234_n N_A_1451_424#_c_1379_n 3.44953e-19 $X=8.91 $Y=0.54
+ $X2=0 $Y2=0
cc_866 N_A_1689_424#_c_1218_n N_A_1451_424#_c_1379_n 3.44953e-19 $X=8.91
+ $Y=1.055 $X2=0 $Y2=0
cc_867 N_A_1689_424#_c_1220_n N_A_1451_424#_c_1442_n 7.34805e-19 $X=11.11
+ $Y=0.715 $X2=0 $Y2=0
cc_868 N_A_1689_424#_c_1220_n N_A_1451_424#_c_1380_n 0.0148352f $X=11.11
+ $Y=0.715 $X2=0 $Y2=0
cc_869 N_A_1689_424#_c_1215_n N_A_1895_424#_M1009_d 0.00633935f $X=10.765
+ $Y=0.34 $X2=-0.19 $Y2=-0.245
cc_870 N_A_1689_424#_M1001_d N_A_1895_424#_c_1537_n 0.00459945f $X=11.615
+ $Y=1.96 $X2=0 $Y2=0
cc_871 N_A_1689_424#_c_1214_n N_A_1895_424#_c_1537_n 0.0174486f $X=10.87
+ $Y=1.885 $X2=0 $Y2=0
cc_872 N_A_1689_424#_c_1293_p N_A_1895_424#_c_1537_n 0.0102889f $X=11.24
+ $Y=2.075 $X2=0 $Y2=0
cc_873 N_A_1689_424#_c_1223_n N_A_1895_424#_c_1537_n 0.0170132f $X=11.765
+ $Y=2.115 $X2=0 $Y2=0
cc_874 N_A_1689_424#_M1001_d N_A_1895_424#_c_1518_n 0.00800216f $X=11.615
+ $Y=1.96 $X2=0 $Y2=0
cc_875 N_A_1689_424#_c_1223_n N_A_1895_424#_c_1518_n 0.0104278f $X=11.765
+ $Y=2.115 $X2=0 $Y2=0
cc_876 N_A_1689_424#_c_1293_p N_VPWR_M1032_d 0.00689106f $X=11.24 $Y=2.075 $X2=0
+ $Y2=0
cc_877 N_A_1689_424#_c_1223_n N_VPWR_M1032_d 0.00324721f $X=11.765 $Y=2.115
+ $X2=0 $Y2=0
cc_878 N_A_1689_424#_c_1214_n N_VPWR_c_1638_n 0.00317855f $X=10.87 $Y=1.885
+ $X2=0 $Y2=0
cc_879 N_A_1689_424#_c_1214_n N_VPWR_c_1644_n 0.00448815f $X=10.87 $Y=1.885
+ $X2=0 $Y2=0
cc_880 N_A_1689_424#_c_1214_n N_VPWR_c_1627_n 0.00399413f $X=10.87 $Y=1.885
+ $X2=0 $Y2=0
cc_881 N_A_1689_424#_c_1215_n N_A_2052_424#_M1027_d 0.00431152f $X=10.765
+ $Y=0.34 $X2=-0.19 $Y2=-0.245
cc_882 N_A_1689_424#_c_1214_n N_A_2052_424#_c_1949_n 0.0111473f $X=10.87
+ $Y=1.885 $X2=0 $Y2=0
cc_883 N_A_1689_424#_M1011_g N_A_2052_424#_c_1951_n 0.00212364f $X=10.855
+ $Y=0.715 $X2=0 $Y2=0
cc_884 N_A_1689_424#_c_1215_n N_A_2052_424#_c_1951_n 0.0117801f $X=10.765
+ $Y=0.34 $X2=0 $Y2=0
cc_885 N_A_1689_424#_c_1220_n N_A_2052_424#_c_1951_n 0.00371604f $X=11.11
+ $Y=0.715 $X2=0 $Y2=0
cc_886 N_A_1689_424#_M1011_g N_A_2052_424#_c_1946_n 0.00556552f $X=10.855
+ $Y=0.715 $X2=0 $Y2=0
cc_887 N_A_1689_424#_c_1214_n N_A_2052_424#_c_1946_n 0.0167111f $X=10.87
+ $Y=1.885 $X2=0 $Y2=0
cc_888 N_A_1689_424#_c_1217_n N_A_2052_424#_c_1946_n 0.055213f $X=11.075
+ $Y=1.635 $X2=0 $Y2=0
cc_889 N_A_1689_424#_c_1293_p N_A_2052_424#_c_1946_n 0.00651472f $X=11.24
+ $Y=2.075 $X2=0 $Y2=0
cc_890 N_A_1689_424#_M1011_g N_A_2052_424#_c_1947_n 0.00466666f $X=10.855
+ $Y=0.715 $X2=0 $Y2=0
cc_891 N_A_1689_424#_c_1215_n N_A_2052_424#_c_1947_n 0.00160061f $X=10.765
+ $Y=0.34 $X2=0 $Y2=0
cc_892 N_A_1689_424#_c_1217_n N_A_2052_424#_c_1947_n 0.0101416f $X=11.075
+ $Y=1.635 $X2=0 $Y2=0
cc_893 N_A_1689_424#_c_1220_n N_A_2052_424#_c_1947_n 0.00415638f $X=11.11
+ $Y=0.715 $X2=0 $Y2=0
cc_894 N_A_1689_424#_c_1223_n COUT 0.00752309f $X=11.765 $Y=2.115 $X2=0 $Y2=0
cc_895 N_A_1689_424#_c_1220_n N_VGND_M1011_d 0.00733558f $X=11.11 $Y=0.715 $X2=0
+ $Y2=0
cc_896 N_A_1689_424#_M1011_g N_VGND_c_2047_n 9.38288e-19 $X=10.855 $Y=0.715
+ $X2=0 $Y2=0
cc_897 N_A_1689_424#_c_1215_n N_VGND_c_2047_n 0.0130541f $X=10.765 $Y=0.34 $X2=0
+ $Y2=0
cc_898 N_A_1689_424#_c_1220_n N_VGND_c_2047_n 0.0248266f $X=11.11 $Y=0.715 $X2=0
+ $Y2=0
cc_899 N_A_1689_424#_c_1220_n N_VGND_c_2048_n 0.0191013f $X=11.11 $Y=0.715 $X2=0
+ $Y2=0
cc_900 N_A_1689_424#_M1011_g N_VGND_c_2054_n 9.43124e-19 $X=10.855 $Y=0.715
+ $X2=0 $Y2=0
cc_901 N_A_1689_424#_c_1215_n N_VGND_c_2054_n 0.120865f $X=10.765 $Y=0.34 $X2=0
+ $Y2=0
cc_902 N_A_1689_424#_c_1216_n N_VGND_c_2054_n 0.0236566f $X=9.075 $Y=0.34 $X2=0
+ $Y2=0
cc_903 N_A_1689_424#_c_1220_n N_VGND_c_2054_n 0.00210799f $X=11.11 $Y=0.715
+ $X2=0 $Y2=0
cc_904 N_A_1689_424#_c_1220_n N_VGND_c_2057_n 0.0149664f $X=11.11 $Y=0.715 $X2=0
+ $Y2=0
cc_905 N_A_1689_424#_c_1215_n N_VGND_c_2063_n 0.070117f $X=10.765 $Y=0.34 $X2=0
+ $Y2=0
cc_906 N_A_1689_424#_c_1216_n N_VGND_c_2063_n 0.0128296f $X=9.075 $Y=0.34 $X2=0
+ $Y2=0
cc_907 N_A_1689_424#_c_1220_n N_VGND_c_2063_n 0.0204199f $X=11.11 $Y=0.715 $X2=0
+ $Y2=0
cc_908 CI N_A_1451_424#_c_1381_n 2.41345e-19 $X=11.675 $Y=1.58 $X2=0 $Y2=0
cc_909 N_CI_c_1330_n N_A_1451_424#_c_1374_n 0.00411358f $X=11.54 $Y=1.885 $X2=0
+ $Y2=0
cc_910 N_CI_c_1332_n N_A_1451_424#_c_1374_n 0.00673467f $X=11.505 $Y=1.26 $X2=0
+ $Y2=0
cc_911 CI N_A_1451_424#_c_1374_n 7.73815e-19 $X=11.675 $Y=1.58 $X2=0 $Y2=0
cc_912 N_CI_c_1330_n N_A_1451_424#_c_1375_n 0.00260536f $X=11.54 $Y=1.885 $X2=0
+ $Y2=0
cc_913 CI N_A_1451_424#_c_1375_n 0.00384117f $X=11.675 $Y=1.58 $X2=0 $Y2=0
cc_914 CI N_A_1451_424#_c_1378_n 0.00291244f $X=11.675 $Y=1.58 $X2=0 $Y2=0
cc_915 N_CI_c_1331_n N_A_1451_424#_c_1380_n 0.00175175f $X=11.505 $Y=1.11 $X2=0
+ $Y2=0
cc_916 N_CI_c_1332_n N_A_1451_424#_c_1380_n 0.00425048f $X=11.505 $Y=1.26 $X2=0
+ $Y2=0
cc_917 CI N_A_1451_424#_c_1380_n 0.006855f $X=11.675 $Y=1.58 $X2=0 $Y2=0
cc_918 N_CI_c_1330_n N_A_1895_424#_c_1537_n 0.0145452f $X=11.54 $Y=1.885 $X2=0
+ $Y2=0
cc_919 N_CI_c_1330_n N_A_1895_424#_c_1518_n 0.00857739f $X=11.54 $Y=1.885 $X2=0
+ $Y2=0
cc_920 N_CI_c_1330_n N_VPWR_c_1632_n 0.00814935f $X=11.54 $Y=1.885 $X2=0 $Y2=0
cc_921 N_CI_c_1330_n N_VPWR_c_1639_n 0.00317855f $X=11.54 $Y=1.885 $X2=0 $Y2=0
cc_922 N_CI_c_1330_n N_VPWR_c_1644_n 0.00448815f $X=11.54 $Y=1.885 $X2=0 $Y2=0
cc_923 N_CI_c_1330_n N_VPWR_c_1627_n 0.00402409f $X=11.54 $Y=1.885 $X2=0 $Y2=0
cc_924 N_CI_c_1330_n N_A_2052_424#_c_1949_n 0.0010181f $X=11.54 $Y=1.885 $X2=0
+ $Y2=0
cc_925 N_CI_c_1331_n N_VGND_c_2047_n 0.00401623f $X=11.505 $Y=1.11 $X2=0 $Y2=0
cc_926 N_CI_c_1331_n N_VGND_c_2048_n 0.00332406f $X=11.505 $Y=1.11 $X2=0 $Y2=0
cc_927 N_CI_c_1331_n N_VGND_c_2057_n 0.00469528f $X=11.505 $Y=1.11 $X2=0 $Y2=0
cc_928 N_CI_c_1331_n N_VGND_c_2063_n 0.00537853f $X=11.505 $Y=1.11 $X2=0 $Y2=0
cc_929 N_A_1451_424#_c_1378_n N_A_1895_424#_M1009_d 0.00961849f $X=12.095
+ $Y=0.925 $X2=-0.19 $Y2=-0.245
cc_930 N_A_1451_424#_c_1382_n N_A_1895_424#_c_1511_n 0.0377617f $X=12.98
+ $Y=1.765 $X2=0 $Y2=0
cc_931 N_A_1451_424#_c_1373_n N_A_1895_424#_M1022_g 0.0177055f $X=12.965 $Y=1.22
+ $X2=0 $Y2=0
cc_932 N_A_1451_424#_c_1375_n N_A_1895_424#_M1022_g 0.00334468f $X=12.965
+ $Y=1.492 $X2=0 $Y2=0
cc_933 N_A_1451_424#_c_1381_n N_A_1895_424#_c_1514_n 0.0174893f $X=12.53
+ $Y=1.765 $X2=0 $Y2=0
cc_934 N_A_1451_424#_c_1382_n N_A_1895_424#_c_1514_n 0.0159569f $X=12.98
+ $Y=1.765 $X2=0 $Y2=0
cc_935 N_A_1451_424#_c_1382_n N_A_1895_424#_c_1506_n 0.00666426f $X=12.98
+ $Y=1.765 $X2=0 $Y2=0
cc_936 N_A_1451_424#_c_1375_n N_A_1895_424#_c_1506_n 9.83334e-19 $X=12.965
+ $Y=1.492 $X2=0 $Y2=0
cc_937 N_A_1451_424#_c_1378_n N_A_1895_424#_c_1507_n 0.012893f $X=12.095
+ $Y=0.925 $X2=0 $Y2=0
cc_938 N_A_1451_424#_c_1381_n N_A_1895_424#_c_1518_n 0.00339403f $X=12.53
+ $Y=1.765 $X2=0 $Y2=0
cc_939 N_A_1451_424#_c_1375_n N_A_1895_424#_c_1509_n 0.00285281f $X=12.965
+ $Y=1.492 $X2=0 $Y2=0
cc_940 N_A_1451_424#_c_1375_n N_A_1895_424#_c_1510_n 0.0272512f $X=12.965
+ $Y=1.492 $X2=0 $Y2=0
cc_941 N_A_1451_424#_c_1381_n N_VPWR_c_1632_n 0.00974588f $X=12.53 $Y=1.765
+ $X2=0 $Y2=0
cc_942 N_A_1451_424#_c_1382_n N_VPWR_c_1632_n 0.00112373f $X=12.98 $Y=1.765
+ $X2=0 $Y2=0
cc_943 N_A_1451_424#_c_1381_n N_VPWR_c_1633_n 0.00112373f $X=12.53 $Y=1.765
+ $X2=0 $Y2=0
cc_944 N_A_1451_424#_c_1382_n N_VPWR_c_1633_n 0.00871578f $X=12.98 $Y=1.765
+ $X2=0 $Y2=0
cc_945 N_A_1451_424#_c_1381_n N_VPWR_c_1640_n 0.00413917f $X=12.53 $Y=1.765
+ $X2=0 $Y2=0
cc_946 N_A_1451_424#_c_1382_n N_VPWR_c_1640_n 0.00413917f $X=12.98 $Y=1.765
+ $X2=0 $Y2=0
cc_947 N_A_1451_424#_c_1381_n N_VPWR_c_1627_n 0.00403181f $X=12.53 $Y=1.765
+ $X2=0 $Y2=0
cc_948 N_A_1451_424#_c_1382_n N_VPWR_c_1627_n 0.00403181f $X=12.98 $Y=1.765
+ $X2=0 $Y2=0
cc_949 N_A_1451_424#_c_1378_n N_A_2052_424#_M1027_d 0.00464304f $X=12.095
+ $Y=0.925 $X2=-0.19 $Y2=-0.245
cc_950 N_A_1451_424#_c_1378_n N_A_2052_424#_c_1951_n 0.0107774f $X=12.095
+ $Y=0.925 $X2=0 $Y2=0
cc_951 N_A_1451_424#_c_1378_n N_A_2052_424#_c_1947_n 0.0106051f $X=12.095
+ $Y=0.925 $X2=0 $Y2=0
cc_952 N_A_1451_424#_c_1372_n N_COUT_c_1985_n 0.0165465f $X=12.535 $Y=1.22 $X2=0
+ $Y2=0
cc_953 N_A_1451_424#_c_1373_n N_COUT_c_1985_n 0.00285048f $X=12.965 $Y=1.22
+ $X2=0 $Y2=0
cc_954 N_A_1451_424#_c_1375_n N_COUT_c_1985_n 0.0199596f $X=12.965 $Y=1.492
+ $X2=0 $Y2=0
cc_955 N_A_1451_424#_c_1442_n N_COUT_c_1985_n 0.00150776f $X=12.24 $Y=0.925
+ $X2=0 $Y2=0
cc_956 N_A_1451_424#_c_1380_n N_COUT_c_1985_n 0.0419855f $X=12.24 $Y=0.925 $X2=0
+ $Y2=0
cc_957 N_A_1451_424#_c_1381_n COUT 0.014527f $X=12.53 $Y=1.765 $X2=0 $Y2=0
cc_958 N_A_1451_424#_c_1382_n COUT 0.00660289f $X=12.98 $Y=1.765 $X2=0 $Y2=0
cc_959 N_A_1451_424#_c_1375_n COUT 0.024684f $X=12.965 $Y=1.492 $X2=0 $Y2=0
cc_960 N_A_1451_424#_c_1378_n N_VGND_M1011_d 0.00119691f $X=12.095 $Y=0.925
+ $X2=0 $Y2=0
cc_961 N_A_1451_424#_c_1442_n N_VGND_M1014_s 0.0023149f $X=12.24 $Y=0.925 $X2=0
+ $Y2=0
cc_962 N_A_1451_424#_c_1380_n N_VGND_M1014_s 0.00530594f $X=12.24 $Y=0.925 $X2=0
+ $Y2=0
cc_963 N_A_1451_424#_c_1378_n N_VGND_c_2047_n 0.00140037f $X=12.095 $Y=0.925
+ $X2=0 $Y2=0
cc_964 N_A_1451_424#_c_1372_n N_VGND_c_2048_n 0.00875775f $X=12.535 $Y=1.22
+ $X2=0 $Y2=0
cc_965 N_A_1451_424#_c_1374_n N_VGND_c_2048_n 0.00109031f $X=12.44 $Y=1.385
+ $X2=0 $Y2=0
cc_966 N_A_1451_424#_c_1378_n N_VGND_c_2048_n 5.68876e-19 $X=12.095 $Y=0.925
+ $X2=0 $Y2=0
cc_967 N_A_1451_424#_c_1442_n N_VGND_c_2048_n 0.0024859f $X=12.24 $Y=0.925 $X2=0
+ $Y2=0
cc_968 N_A_1451_424#_c_1380_n N_VGND_c_2048_n 0.0233714f $X=12.24 $Y=0.925 $X2=0
+ $Y2=0
cc_969 N_A_1451_424#_c_1372_n N_VGND_c_2049_n 6.14817e-19 $X=12.535 $Y=1.22
+ $X2=0 $Y2=0
cc_970 N_A_1451_424#_c_1373_n N_VGND_c_2049_n 0.0143497f $X=12.965 $Y=1.22 $X2=0
+ $Y2=0
cc_971 N_A_1451_424#_c_1375_n N_VGND_c_2049_n 0.00155918f $X=12.965 $Y=1.492
+ $X2=0 $Y2=0
cc_972 N_A_1451_424#_c_1376_n N_VGND_c_2054_n 0.0203841f $X=8.225 $Y=1.04 $X2=0
+ $Y2=0
cc_973 N_A_1451_424#_c_1372_n N_VGND_c_2058_n 0.00434272f $X=12.535 $Y=1.22
+ $X2=0 $Y2=0
cc_974 N_A_1451_424#_c_1373_n N_VGND_c_2058_n 0.00383152f $X=12.965 $Y=1.22
+ $X2=0 $Y2=0
cc_975 N_A_1451_424#_c_1372_n N_VGND_c_2063_n 0.00825283f $X=12.535 $Y=1.22
+ $X2=0 $Y2=0
cc_976 N_A_1451_424#_c_1373_n N_VGND_c_2063_n 0.0075754f $X=12.965 $Y=1.22 $X2=0
+ $Y2=0
cc_977 N_A_1451_424#_c_1376_n N_VGND_c_2063_n 0.019286f $X=8.225 $Y=1.04 $X2=0
+ $Y2=0
cc_978 N_A_1451_424#_c_1380_n N_VGND_c_2063_n 0.00110717f $X=12.24 $Y=0.925
+ $X2=0 $Y2=0
cc_979 N_A_1895_424#_c_1537_n N_VPWR_M1032_d 0.0122082f $X=11.8 $Y=2.685 $X2=0
+ $Y2=0
cc_980 N_A_1895_424#_c_1514_n N_VPWR_M1023_s 0.0108986f $X=13.23 $Y=2.455 $X2=0
+ $Y2=0
cc_981 N_A_1895_424#_c_1514_n N_VPWR_M1026_s 0.00641412f $X=13.23 $Y=2.455 $X2=0
+ $Y2=0
cc_982 N_A_1895_424#_c_1506_n N_VPWR_M1026_s 0.00582265f $X=13.315 $Y=2.37 $X2=0
+ $Y2=0
cc_983 N_A_1895_424#_c_1514_n N_VPWR_c_1632_n 0.02153f $X=13.23 $Y=2.455 $X2=0
+ $Y2=0
cc_984 N_A_1895_424#_c_1518_n N_VPWR_c_1632_n 0.00475706f $X=11.885 $Y=2.455
+ $X2=0 $Y2=0
cc_985 N_A_1895_424#_c_1511_n N_VPWR_c_1633_n 0.00690587f $X=13.43 $Y=1.765
+ $X2=0 $Y2=0
cc_986 N_A_1895_424#_c_1512_n N_VPWR_c_1633_n 4.28852e-19 $X=13.89 $Y=1.765
+ $X2=0 $Y2=0
cc_987 N_A_1895_424#_c_1514_n N_VPWR_c_1633_n 0.0173772f $X=13.23 $Y=2.455 $X2=0
+ $Y2=0
cc_988 N_A_1895_424#_c_1512_n N_VPWR_c_1635_n 0.00806255f $X=13.89 $Y=1.765
+ $X2=0 $Y2=0
cc_989 N_A_1895_424#_c_1537_n N_VPWR_c_1638_n 0.0173595f $X=11.8 $Y=2.685 $X2=0
+ $Y2=0
cc_990 N_A_1895_424#_c_1517_n N_VPWR_c_1638_n 0.0146357f $X=9.91 $Y=2.685 $X2=0
+ $Y2=0
cc_991 N_A_1895_424#_c_1537_n N_VPWR_c_1639_n 0.00723205f $X=11.8 $Y=2.685 $X2=0
+ $Y2=0
cc_992 N_A_1895_424#_c_1518_n N_VPWR_c_1639_n 0.00376635f $X=11.885 $Y=2.455
+ $X2=0 $Y2=0
cc_993 N_A_1895_424#_c_1511_n N_VPWR_c_1641_n 0.00413917f $X=13.43 $Y=1.765
+ $X2=0 $Y2=0
cc_994 N_A_1895_424#_c_1512_n N_VPWR_c_1641_n 0.00394617f $X=13.89 $Y=1.765
+ $X2=0 $Y2=0
cc_995 N_A_1895_424#_c_1537_n N_VPWR_c_1644_n 0.0280851f $X=11.8 $Y=2.685 $X2=0
+ $Y2=0
cc_996 N_A_1895_424#_c_1511_n N_VPWR_c_1627_n 0.00723278f $X=13.43 $Y=1.765
+ $X2=0 $Y2=0
cc_997 N_A_1895_424#_c_1512_n N_VPWR_c_1627_n 0.00696441f $X=13.89 $Y=1.765
+ $X2=0 $Y2=0
cc_998 N_A_1895_424#_c_1537_n N_VPWR_c_1627_n 0.0405218f $X=11.8 $Y=2.685 $X2=0
+ $Y2=0
cc_999 N_A_1895_424#_c_1514_n N_VPWR_c_1627_n 0.0281946f $X=13.23 $Y=2.455 $X2=0
+ $Y2=0
cc_1000 N_A_1895_424#_c_1517_n N_VPWR_c_1627_n 0.0121141f $X=9.91 $Y=2.685 $X2=0
+ $Y2=0
cc_1001 N_A_1895_424#_c_1518_n N_VPWR_c_1627_n 0.00526389f $X=11.885 $Y=2.455
+ $X2=0 $Y2=0
cc_1002 N_A_1895_424#_c_1537_n N_A_2052_424#_M1013_d 0.0127788f $X=11.8 $Y=2.685
+ $X2=0 $Y2=0
cc_1003 N_A_1895_424#_c_1537_n N_A_2052_424#_c_1949_n 0.0334905f $X=11.8
+ $Y=2.685 $X2=0 $Y2=0
cc_1004 N_A_1895_424#_c_1513_n N_A_2052_424#_c_1946_n 7.68717e-19 $X=9.91
+ $Y=2.265 $X2=0 $Y2=0
cc_1005 N_A_1895_424#_c_1514_n N_COUT_M1023_d 0.00555567f $X=13.23 $Y=2.455
+ $X2=0 $Y2=0
cc_1006 N_A_1895_424#_M1022_g N_COUT_c_1985_n 3.16505e-19 $X=13.465 $Y=0.74
+ $X2=0 $Y2=0
cc_1007 N_A_1895_424#_c_1509_n N_COUT_c_1985_n 0.0102461f $X=13.445 $Y=1.465
+ $X2=0 $Y2=0
cc_1008 N_A_1895_424#_c_1510_n N_COUT_c_1985_n 2.11853e-19 $X=13.89 $Y=1.532
+ $X2=0 $Y2=0
cc_1009 N_A_1895_424#_c_1511_n COUT 3.90923e-19 $X=13.43 $Y=1.765 $X2=0 $Y2=0
cc_1010 N_A_1895_424#_c_1514_n COUT 0.0175546f $X=13.23 $Y=2.455 $X2=0 $Y2=0
cc_1011 N_A_1895_424#_c_1506_n COUT 0.026816f $X=13.315 $Y=2.37 $X2=0 $Y2=0
cc_1012 N_A_1895_424#_c_1509_n COUT 0.00398792f $X=13.445 $Y=1.465 $X2=0 $Y2=0
cc_1013 N_A_1895_424#_M1022_g N_SUM_c_2007_n 0.00545316f $X=13.465 $Y=0.74 $X2=0
+ $Y2=0
cc_1014 N_A_1895_424#_M1029_g N_SUM_c_2007_n 3.54397e-19 $X=13.905 $Y=0.74 $X2=0
+ $Y2=0
cc_1015 N_A_1895_424#_c_1511_n N_SUM_c_2010_n 0.0073959f $X=13.43 $Y=1.765 $X2=0
+ $Y2=0
cc_1016 N_A_1895_424#_c_1512_n N_SUM_c_2010_n 0.00217259f $X=13.89 $Y=1.765
+ $X2=0 $Y2=0
cc_1017 N_A_1895_424#_c_1506_n N_SUM_c_2010_n 0.040394f $X=13.315 $Y=2.37 $X2=0
+ $Y2=0
cc_1018 N_A_1895_424#_c_1510_n N_SUM_c_2010_n 0.00605575f $X=13.89 $Y=1.532
+ $X2=0 $Y2=0
cc_1019 N_A_1895_424#_c_1512_n N_SUM_c_2011_n 0.0143931f $X=13.89 $Y=1.765 $X2=0
+ $Y2=0
cc_1020 N_A_1895_424#_c_1514_n N_SUM_c_2011_n 0.0139285f $X=13.23 $Y=2.455 $X2=0
+ $Y2=0
cc_1021 N_A_1895_424#_c_1511_n N_SUM_c_2008_n 3.75863e-19 $X=13.43 $Y=1.765
+ $X2=0 $Y2=0
cc_1022 N_A_1895_424#_c_1512_n N_SUM_c_2008_n 0.00266312f $X=13.89 $Y=1.765
+ $X2=0 $Y2=0
cc_1023 N_A_1895_424#_c_1506_n N_SUM_c_2008_n 0.00875049f $X=13.315 $Y=2.37
+ $X2=0 $Y2=0
cc_1024 N_A_1895_424#_c_1509_n N_SUM_c_2008_n 0.00881172f $X=13.445 $Y=1.465
+ $X2=0 $Y2=0
cc_1025 N_A_1895_424#_c_1510_n N_SUM_c_2008_n 0.0188037f $X=13.89 $Y=1.532 $X2=0
+ $Y2=0
cc_1026 N_A_1895_424#_M1022_g SUM 0.00866623f $X=13.465 $Y=0.74 $X2=0 $Y2=0
cc_1027 N_A_1895_424#_M1029_g SUM 0.0220314f $X=13.905 $Y=0.74 $X2=0 $Y2=0
cc_1028 N_A_1895_424#_c_1509_n SUM 0.0176448f $X=13.445 $Y=1.465 $X2=0 $Y2=0
cc_1029 N_A_1895_424#_c_1510_n SUM 0.0218479f $X=13.89 $Y=1.532 $X2=0 $Y2=0
cc_1030 N_A_1895_424#_M1022_g N_VGND_c_2049_n 0.00585869f $X=13.465 $Y=0.74
+ $X2=0 $Y2=0
cc_1031 N_A_1895_424#_c_1509_n N_VGND_c_2049_n 0.00982041f $X=13.445 $Y=1.465
+ $X2=0 $Y2=0
cc_1032 N_A_1895_424#_c_1510_n N_VGND_c_2049_n 0.00149751f $X=13.89 $Y=1.532
+ $X2=0 $Y2=0
cc_1033 N_A_1895_424#_M1022_g N_VGND_c_2051_n 4.35221e-19 $X=13.465 $Y=0.74
+ $X2=0 $Y2=0
cc_1034 N_A_1895_424#_M1029_g N_VGND_c_2051_n 0.00835923f $X=13.905 $Y=0.74
+ $X2=0 $Y2=0
cc_1035 N_A_1895_424#_M1022_g N_VGND_c_2059_n 0.0043438f $X=13.465 $Y=0.74 $X2=0
+ $Y2=0
cc_1036 N_A_1895_424#_M1029_g N_VGND_c_2059_n 0.00383152f $X=13.905 $Y=0.74
+ $X2=0 $Y2=0
cc_1037 N_A_1895_424#_M1022_g N_VGND_c_2063_n 0.00820957f $X=13.465 $Y=0.74
+ $X2=0 $Y2=0
cc_1038 N_A_1895_424#_M1029_g N_VGND_c_2063_n 0.00375467f $X=13.905 $Y=0.74
+ $X2=0 $Y2=0
cc_1039 N_VPWR_c_1629_n N_A_114_368#_c_1766_n 0.0561756f $X=0.27 $Y=2.325 $X2=0
+ $Y2=0
cc_1040 N_VPWR_c_1636_n N_A_114_368#_c_1766_n 0.0145938f $X=1.54 $Y=3.33 $X2=0
+ $Y2=0
cc_1041 N_VPWR_c_1627_n N_A_114_368#_c_1766_n 0.0120466f $X=14.16 $Y=3.33 $X2=0
+ $Y2=0
cc_1042 N_VPWR_M1002_s N_A_114_368#_c_1768_n 0.00680795f $X=0.135 $Y=1.84 $X2=0
+ $Y2=0
cc_1043 N_VPWR_c_1629_n N_A_114_368#_c_1768_n 0.00195261f $X=0.27 $Y=2.325 $X2=0
+ $Y2=0
cc_1044 N_VPWR_c_1630_n N_A_114_368#_c_1761_n 0.00189778f $X=1.705 $Y=2.115
+ $X2=0 $Y2=0
cc_1045 N_VPWR_c_1631_n N_A_413_392#_c_1865_n 0.0129575f $X=6.43 $Y=2.745 $X2=0
+ $Y2=0
cc_1046 N_VPWR_c_1637_n N_A_413_392#_c_1865_n 0.216431f $X=6.265 $Y=3.33 $X2=0
+ $Y2=0
cc_1047 N_VPWR_c_1627_n N_A_413_392#_c_1865_n 0.134389f $X=14.16 $Y=3.33 $X2=0
+ $Y2=0
cc_1048 N_VPWR_c_1630_n N_A_413_392#_c_1866_n 0.0105843f $X=1.705 $Y=2.115 $X2=0
+ $Y2=0
cc_1049 N_VPWR_c_1637_n N_A_413_392#_c_1866_n 0.0215391f $X=6.265 $Y=3.33 $X2=0
+ $Y2=0
cc_1050 N_VPWR_c_1627_n N_A_413_392#_c_1866_n 0.0126858f $X=14.16 $Y=3.33 $X2=0
+ $Y2=0
cc_1051 N_VPWR_c_1631_n N_A_413_392#_c_1867_n 0.0222247f $X=6.43 $Y=2.745 $X2=0
+ $Y2=0
cc_1052 N_VPWR_c_1630_n N_A_413_392#_c_1861_n 0.00162355f $X=1.705 $Y=2.115
+ $X2=0 $Y2=0
cc_1053 N_VPWR_c_1635_n N_SUM_c_2010_n 0.0876529f $X=14.13 $Y=1.985 $X2=0 $Y2=0
cc_1054 N_VPWR_c_1633_n N_SUM_c_2011_n 0.0184122f $X=13.205 $Y=2.805 $X2=0 $Y2=0
cc_1055 N_VPWR_c_1641_n N_SUM_c_2011_n 0.0133438f $X=14.045 $Y=3.33 $X2=0 $Y2=0
cc_1056 N_VPWR_c_1627_n N_SUM_c_2011_n 0.0109062f $X=14.16 $Y=3.33 $X2=0 $Y2=0
cc_1057 N_VPWR_c_1635_n SUM 0.013979f $X=14.13 $Y=1.985 $X2=0 $Y2=0
cc_1058 N_A_114_368#_M1010_d N_A_413_392#_c_1865_n 0.00405827f $X=3.635 $Y=2.12
+ $X2=0 $Y2=0
cc_1059 N_A_114_368#_c_1761_n N_A_413_392#_c_1861_n 0.024605f $X=3.935 $Y=1.295
+ $X2=0 $Y2=0
cc_1060 N_A_114_368#_c_1761_n N_A_413_392#_c_1862_n 0.0101757f $X=3.935 $Y=1.295
+ $X2=0 $Y2=0
cc_1061 N_A_114_368#_c_1758_n N_VGND_c_2044_n 0.017529f $X=0.8 $Y=0.515 $X2=0
+ $Y2=0
cc_1062 N_A_114_368#_c_1761_n N_VGND_c_2044_n 9.72863e-19 $X=3.935 $Y=1.295
+ $X2=0 $Y2=0
cc_1063 N_A_114_368#_c_1762_n N_VGND_c_2044_n 0.00174148f $X=0.385 $Y=1.295
+ $X2=0 $Y2=0
cc_1064 N_A_114_368#_c_1764_n N_VGND_c_2044_n 0.0121491f $X=0.492 $Y=1.215 $X2=0
+ $Y2=0
cc_1065 N_A_114_368#_c_1761_n N_VGND_c_2045_n 0.00737634f $X=3.935 $Y=1.295
+ $X2=0 $Y2=0
cc_1066 N_A_114_368#_c_1758_n N_VGND_c_2052_n 0.0115122f $X=0.8 $Y=0.515 $X2=0
+ $Y2=0
cc_1067 N_A_114_368#_c_1758_n N_VGND_c_2063_n 0.0095288f $X=0.8 $Y=0.515 $X2=0
+ $Y2=0
cc_1068 N_A_413_392#_c_1858_n N_VGND_c_2045_n 0.0181851f $X=2.47 $Y=0.67 $X2=0
+ $Y2=0
cc_1069 N_A_413_392#_c_1860_n N_VGND_c_2045_n 0.014022f $X=2.555 $Y=0.34 $X2=0
+ $Y2=0
cc_1070 N_A_413_392#_c_1863_n N_VGND_c_2046_n 0.0195964f $X=5.77 $Y=0.34 $X2=0
+ $Y2=0
cc_1071 N_A_413_392#_c_1859_n N_VGND_c_2056_n 0.196447f $X=5.605 $Y=0.34 $X2=0
+ $Y2=0
cc_1072 N_A_413_392#_c_1860_n N_VGND_c_2056_n 0.0179217f $X=2.555 $Y=0.34 $X2=0
+ $Y2=0
cc_1073 N_A_413_392#_c_1863_n N_VGND_c_2056_n 0.0229596f $X=5.77 $Y=0.34 $X2=0
+ $Y2=0
cc_1074 N_A_413_392#_c_1859_n N_VGND_c_2063_n 0.114669f $X=5.605 $Y=0.34 $X2=0
+ $Y2=0
cc_1075 N_A_413_392#_c_1860_n N_VGND_c_2063_n 0.00971942f $X=2.555 $Y=0.34 $X2=0
+ $Y2=0
cc_1076 N_A_413_392#_c_1863_n N_VGND_c_2063_n 0.0126481f $X=5.77 $Y=0.34 $X2=0
+ $Y2=0
cc_1077 N_COUT_c_1985_n N_VGND_c_2048_n 0.0107203f $X=12.75 $Y=0.515 $X2=0 $Y2=0
cc_1078 N_COUT_c_1985_n N_VGND_c_2049_n 0.0294122f $X=12.75 $Y=0.515 $X2=0 $Y2=0
cc_1079 N_COUT_c_1985_n N_VGND_c_2058_n 0.0109942f $X=12.75 $Y=0.515 $X2=0 $Y2=0
cc_1080 N_COUT_c_1985_n N_VGND_c_2063_n 0.00904371f $X=12.75 $Y=0.515 $X2=0
+ $Y2=0
cc_1081 SUM N_VGND_M1029_d 0.00428496f $X=14.075 $Y=0.84 $X2=0 $Y2=0
cc_1082 N_SUM_c_2007_n N_VGND_c_2049_n 0.016738f $X=13.685 $Y=0.52 $X2=0 $Y2=0
cc_1083 SUM N_VGND_c_2049_n 0.0146948f $X=14.075 $Y=0.84 $X2=0 $Y2=0
cc_1084 N_SUM_c_2007_n N_VGND_c_2051_n 0.0108837f $X=13.685 $Y=0.52 $X2=0 $Y2=0
cc_1085 SUM N_VGND_c_2051_n 0.0229706f $X=14.075 $Y=0.84 $X2=0 $Y2=0
cc_1086 N_SUM_c_2007_n N_VGND_c_2059_n 0.011652f $X=13.685 $Y=0.52 $X2=0 $Y2=0
cc_1087 N_SUM_c_2007_n N_VGND_c_2063_n 0.00975232f $X=13.685 $Y=0.52 $X2=0 $Y2=0
cc_1088 SUM N_VGND_c_2063_n 0.00720744f $X=14.075 $Y=0.84 $X2=0 $Y2=0
