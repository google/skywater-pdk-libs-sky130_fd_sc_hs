* File: sky130_fd_sc_hs__nor4b_1.spice
* Created: Tue Sep  1 20:12:21 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hs__nor4b_1.pex.spice"
.subckt sky130_fd_sc_hs__nor4b_1  VNB VPB D_N A B C VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* C	C
* B	B
* A	A
* D_N	D_N
* VPB	VPB
* VNB	VNB
MM1008 N_VGND_M1008_d N_D_N_M1008_g N_A_57_368#_M1008_s VNB NLOWVT L=0.15 W=0.55
+ AD=0.11874 AS=0.15675 PD=0.989147 PS=1.67 NRD=15.264 NRS=0 M=1 R=3.66667
+ SA=75000.2 SB=75002.3 A=0.0825 P=1.4 MULT=1
MM1009 N_Y_M1009_d N_A_M1009_g N_VGND_M1008_d VNB NLOWVT L=0.15 W=0.74 AD=0.1036
+ AS=0.15976 PD=1.02 PS=1.33085 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75000.6
+ SB=75001.7 A=0.111 P=1.78 MULT=1
MM1006 N_VGND_M1006_d N_B_M1006_g N_Y_M1009_d VNB NLOWVT L=0.15 W=0.74 AD=0.1591
+ AS=0.1036 PD=1.17 PS=1.02 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75001.1 SB=75001.3
+ A=0.111 P=1.78 MULT=1
MM1001 N_Y_M1001_d N_C_M1001_g N_VGND_M1006_d VNB NLOWVT L=0.15 W=0.74 AD=0.1036
+ AS=0.1591 PD=1.02 PS=1.17 NRD=0 NRS=12.972 M=1 R=4.93333 SA=75001.6 SB=75000.7
+ A=0.111 P=1.78 MULT=1
MM1005 N_VGND_M1005_d N_A_57_368#_M1005_g N_Y_M1001_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.2627 AS=0.1036 PD=2.19 PS=1.02 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75002.1
+ SB=75000.3 A=0.111 P=1.78 MULT=1
MM1002 N_VPWR_M1002_d N_D_N_M1002_g N_A_57_368#_M1002_s VPB PSHORT L=0.15 W=0.84
+ AD=0.1866 AS=0.2478 PD=1.32 PS=2.27 NRD=30.4759 NRS=2.3443 M=1 R=5.6
+ SA=75000.2 SB=75002.4 A=0.126 P=1.98 MULT=1
MM1004 A_260_368# N_A_M1004_g N_VPWR_M1002_d VPB PSHORT L=0.15 W=1.12 AD=0.1512
+ AS=0.2488 PD=1.39 PS=1.76 NRD=14.0658 NRS=1.7533 M=1 R=7.46667 SA=75000.6
+ SB=75001.8 A=0.168 P=2.54 MULT=1
MM1007 A_344_368# N_B_M1007_g A_260_368# VPB PSHORT L=0.15 W=1.12 AD=0.2016
+ AS=0.1512 PD=1.48 PS=1.39 NRD=21.9852 NRS=14.0658 M=1 R=7.46667 SA=75001.1
+ SB=75001.4 A=0.168 P=2.54 MULT=1
MM1000 A_446_368# N_C_M1000_g A_344_368# VPB PSHORT L=0.15 W=1.12 AD=0.2352
+ AS=0.2016 PD=1.54 PS=1.48 NRD=27.2451 NRS=21.9852 M=1 R=7.46667 SA=75001.6
+ SB=75000.9 A=0.168 P=2.54 MULT=1
MM1003 N_Y_M1003_d N_A_57_368#_M1003_g A_446_368# VPB PSHORT L=0.15 W=1.12
+ AD=0.4648 AS=0.2352 PD=3.07 PS=1.54 NRD=22.852 NRS=27.2451 M=1 R=7.46667
+ SA=75002.1 SB=75000.3 A=0.168 P=2.54 MULT=1
DX10_noxref VNB VPB NWDIODE A=6.9564 P=11.2
*
.include "sky130_fd_sc_hs__nor4b_1.pxi.spice"
*
.ends
*
*
