* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hs__dfrbp_1 CLK D RESET_B VGND VNB VPB VPWR Q Q_N
M1000 a_38_78# D VPWR VPB pshort w=420000u l=150000u
+  ad=2.499e+11p pd=2.87e+06u as=2.03935e+12p ps=1.81e+07u
M1001 VPWR RESET_B a_38_78# VPB pshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1002 VGND CLK a_319_360# VNB nlowvt w=740000u l=150000u
+  ad=1.39535e+12p pd=1.224e+07u as=2.109e+11p ps=2.05e+06u
M1003 a_1434_74# a_319_360# a_1224_74# VNB nlowvt w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=4.33e+11p ps=3.08e+06u
M1004 a_841_401# a_706_463# VGND VNB nlowvt w=640000u l=150000u
+  ad=3.222e+11p pd=2.44e+06u as=0p ps=0u
M1005 VPWR a_841_401# a_796_463# VPB pshort w=420000u l=150000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1006 a_910_118# a_841_401# a_832_118# VNB nlowvt w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=1.008e+11p ps=1.32e+06u
M1007 a_1224_74# a_498_360# a_841_401# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VPWR a_1224_74# a_2026_424# VPB pshort w=840000u l=150000u
+  ad=0p pd=0u as=2.478e+11p ps=2.27e+06u
M1009 Q a_2026_424# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1010 Q a_2026_424# VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=3.304e+11p pd=2.83e+06u as=0p ps=0u
M1011 a_125_78# D a_38_78# VNB nlowvt w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=2.394e+11p ps=2.82e+06u
M1012 VGND a_1224_74# a_2026_424# VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=1.5675e+11p ps=1.67e+06u
M1013 a_498_360# a_319_360# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1014 Q_N a_1224_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.627e+11p pd=2.19e+06u as=0p ps=0u
M1015 a_1465_471# a_498_360# a_1224_74# VPB pshort w=420000u l=150000u
+  ad=1.134e+11p pd=1.38e+06u as=3.877e+11p ps=3.2e+06u
M1016 a_1482_48# RESET_B VPWR VPB pshort w=420000u l=150000u
+  ad=1.26e+11p pd=1.44e+06u as=0p ps=0u
M1017 VPWR CLK a_319_360# VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=3.304e+11p ps=2.83e+06u
M1018 a_832_118# a_498_360# a_706_463# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.47e+11p ps=1.54e+06u
M1019 VPWR a_1224_74# a_1482_48# VPB pshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_706_463# a_319_360# a_38_78# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_706_463# a_498_360# a_38_78# VPB pshort w=420000u l=150000u
+  ad=2.436e+11p pd=2.84e+06u as=0p ps=0u
M1022 VGND RESET_B a_910_118# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_498_360# a_319_360# VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=3.304e+11p pd=2.83e+06u as=0p ps=0u
M1024 Q_N a_1224_74# VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=6.888e+11p pd=3.47e+06u as=0p ps=0u
M1025 a_796_463# a_319_360# a_706_463# VPB pshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 VPWR a_1482_48# a_1465_471# VPB pshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 a_706_463# RESET_B VPWR VPB pshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1028 a_841_401# a_706_463# VPWR VPB pshort w=1e+06u l=150000u
+  ad=3e+11p pd=2.6e+06u as=0p ps=0u
M1029 VGND a_1482_48# a_1434_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1030 a_1624_74# RESET_B VGND VNB nlowvt w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=0p ps=0u
M1031 a_1482_48# a_1224_74# a_1624_74# VNB nlowvt w=420000u l=150000u
+  ad=1.197e+11p pd=1.41e+06u as=0p ps=0u
M1032 a_1224_74# a_319_360# a_841_401# VPB pshort w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1033 VGND RESET_B a_125_78# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
