* File: sky130_fd_sc_hs__maj3_4.spice
* Created: Tue Sep  1 20:07:29 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hs__maj3_4.pex.spice"
.subckt sky130_fd_sc_hs__maj3_4  VNB VPB B A C VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* C	C
* A	A
* B	B
* VPB	VPB
* VNB	VNB
MM1015 N_VGND_M1015_d N_A_M1015_g N_A_114_125#_M1015_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.1824 AS=0.174875 PD=1.85 PS=1.315 NRD=0 NRS=40.92 M=1 R=4.26667
+ SA=75000.2 SB=75005.8 A=0.096 P=1.58 MULT=1
MM1017 N_A_114_125#_M1015_s N_B_M1017_g N_A_219_392#_M1017_s VNB NLOWVT L=0.15
+ W=0.64 AD=0.174875 AS=0.0896 PD=1.315 PS=0.92 NRD=40.92 NRS=0 M=1 R=4.26667
+ SA=75000.8 SB=75005.2 A=0.096 P=1.58 MULT=1
MM1025 N_A_114_125#_M1025_d N_B_M1025_g N_A_219_392#_M1017_s VNB NLOWVT L=0.15
+ W=0.64 AD=0.112 AS=0.0896 PD=0.99 PS=0.92 NRD=13.116 NRS=0 M=1 R=4.26667
+ SA=75001.2 SB=75004.8 A=0.096 P=1.58 MULT=1
MM1022 N_VGND_M1022_d N_A_M1022_g N_A_114_125#_M1025_d VNB NLOWVT L=0.15 W=0.64
+ AD=0.0896 AS=0.112 PD=0.92 PS=0.99 NRD=0 NRS=0 M=1 R=4.26667 SA=75001.7
+ SB=75004.3 A=0.096 P=1.58 MULT=1
MM1005 N_VGND_M1022_d N_C_M1005_g N_A_504_125#_M1005_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.0896 AS=0.1088 PD=0.92 PS=0.98 NRD=0 NRS=5.616 M=1 R=4.26667 SA=75002.2
+ SB=75003.8 A=0.096 P=1.58 MULT=1
MM1001 N_A_219_392#_M1001_d N_B_M1001_g N_A_504_125#_M1005_s VNB NLOWVT L=0.15
+ W=0.64 AD=0.0896 AS=0.1088 PD=0.92 PS=0.98 NRD=0 NRS=5.616 M=1 R=4.26667
+ SA=75002.6 SB=75003.3 A=0.096 P=1.58 MULT=1
MM1026 N_A_219_392#_M1001_d N_B_M1026_g N_A_504_125#_M1026_s VNB NLOWVT L=0.15
+ W=0.64 AD=0.0896 AS=0.162087 PD=0.92 PS=1.32 NRD=0 NRS=37.164 M=1 R=4.26667
+ SA=75003.1 SB=75002.9 A=0.096 P=1.58 MULT=1
MM1018 N_VGND_M1018_d N_C_M1018_g N_A_504_125#_M1026_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.112 AS=0.162087 PD=0.99 PS=1.32 NRD=0 NRS=14.988 M=1 R=4.26667 SA=75002.4
+ SB=75002.9 A=0.096 P=1.58 MULT=1
MM1004 N_A_906_78#_M1004_d N_A_M1004_g N_VGND_M1018_d VNB NLOWVT L=0.15 W=0.64
+ AD=0.133137 AS=0.112 PD=1.205 PS=0.99 NRD=0 NRS=13.116 M=1 R=4.26667
+ SA=75002.9 SB=75002.4 A=0.096 P=1.58 MULT=1
MM1003 N_A_219_392#_M1003_d N_C_M1003_g N_A_906_78#_M1004_d VNB NLOWVT L=0.15
+ W=0.64 AD=0.0896 AS=0.133137 PD=0.92 PS=1.205 NRD=0 NRS=28.692 M=1 R=4.26667
+ SA=75003.1 SB=75002.9 A=0.096 P=1.58 MULT=1
MM1007 N_A_219_392#_M1003_d N_C_M1007_g N_A_906_78#_M1007_s VNB NLOWVT L=0.15
+ W=0.64 AD=0.0896 AS=0.0896 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75003.5 SB=75002.5 A=0.096 P=1.58 MULT=1
MM1008 N_A_906_78#_M1007_s N_A_M1008_g N_VGND_M1008_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.0896 AS=0.12007 PD=0.92 PS=1.02029 NRD=0 NRS=15.468 M=1 R=4.26667
+ SA=75003.9 SB=75002 A=0.096 P=1.58 MULT=1
MM1002 N_X_M1002_d N_A_219_392#_M1002_g N_VGND_M1008_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1184 AS=0.13883 PD=1.06 PS=1.17971 NRD=6.48 NRS=0 M=1 R=4.93333
+ SA=75003.9 SB=75001.5 A=0.111 P=1.78 MULT=1
MM1021 N_X_M1002_d N_A_219_392#_M1021_g N_VGND_M1021_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1184 AS=0.1036 PD=1.06 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75004.3
+ SB=75001.1 A=0.111 P=1.78 MULT=1
MM1023 N_X_M1023_d N_A_219_392#_M1023_g N_VGND_M1021_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75004.8
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1027 N_X_M1023_d N_A_219_392#_M1027_g N_VGND_M1027_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1962 PD=1.02 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333 SA=75005.2
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1019 N_A_119_392#_M1019_d N_A_M1019_g N_VPWR_M1019_s VPB PSHORT L=0.15 W=1
+ AD=0.175 AS=0.295 PD=1.35 PS=2.59 NRD=1.9503 NRS=1.9503 M=1 R=6.66667
+ SA=75000.2 SB=75007.4 A=0.15 P=2.3 MULT=1
MM1011 N_A_219_392#_M1011_d N_B_M1011_g N_A_119_392#_M1019_d VPB PSHORT L=0.15
+ W=1 AD=0.15 AS=0.175 PD=1.3 PS=1.35 NRD=1.9503 NRS=11.8003 M=1 R=6.66667
+ SA=75000.7 SB=75006.9 A=0.15 P=2.3 MULT=1
MM1016 N_A_219_392#_M1011_d N_B_M1016_g N_A_119_392#_M1016_s VPB PSHORT L=0.15
+ W=1 AD=0.15 AS=0.15 PD=1.3 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=6.66667
+ SA=75001.2 SB=75006.4 A=0.15 P=2.3 MULT=1
MM1020 N_A_119_392#_M1016_s N_A_M1020_g N_VPWR_M1020_s VPB PSHORT L=0.15 W=1
+ AD=0.15 AS=0.18 PD=1.3 PS=1.36 NRD=1.9503 NRS=2.9353 M=1 R=6.66667 SA=75001.6
+ SB=75006 A=0.15 P=2.3 MULT=1
MM1009 N_A_501_392#_M1009_d N_C_M1009_g N_VPWR_M1020_s VPB PSHORT L=0.15 W=1
+ AD=0.15 AS=0.18 PD=1.3 PS=1.36 NRD=1.9503 NRS=12.7853 M=1 R=6.66667 SA=75002.1
+ SB=75005.4 A=0.15 P=2.3 MULT=1
MM1012 N_A_501_392#_M1009_d N_B_M1012_g N_A_219_392#_M1012_s VPB PSHORT L=0.15
+ W=1 AD=0.15 AS=0.175 PD=1.3 PS=1.35 NRD=1.9503 NRS=11.8003 M=1 R=6.66667
+ SA=75002.6 SB=75005 A=0.15 P=2.3 MULT=1
MM1014 N_A_501_392#_M1014_d N_B_M1014_g N_A_219_392#_M1012_s VPB PSHORT L=0.15
+ W=1 AD=0.175 AS=0.175 PD=1.35 PS=1.35 NRD=11.8003 NRS=1.9503 M=1 R=6.66667
+ SA=75003.1 SB=75004.5 A=0.15 P=2.3 MULT=1
MM1013 N_A_501_392#_M1014_d N_C_M1013_g N_VPWR_M1013_s VPB PSHORT L=0.15 W=1
+ AD=0.175 AS=0.21 PD=1.35 PS=1.42 NRD=1.9503 NRS=11.8003 M=1 R=6.66667
+ SA=75003.6 SB=75004 A=0.15 P=2.3 MULT=1
MM1006 N_A_905_392#_M1006_d N_A_M1006_g N_VPWR_M1013_s VPB PSHORT L=0.15 W=1
+ AD=0.15 AS=0.21 PD=1.3 PS=1.42 NRD=1.9503 NRS=15.7403 M=1 R=6.66667 SA=75004.1
+ SB=75003.4 A=0.15 P=2.3 MULT=1
MM1010 N_A_219_392#_M1010_d N_C_M1010_g N_A_905_392#_M1006_d VPB PSHORT L=0.15
+ W=1 AD=0.15 AS=0.15 PD=1.3 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=6.66667
+ SA=75004.6 SB=75003 A=0.15 P=2.3 MULT=1
MM1024 N_A_219_392#_M1010_d N_C_M1024_g N_A_905_392#_M1024_s VPB PSHORT L=0.15
+ W=1 AD=0.15 AS=0.15 PD=1.3 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=6.66667 SA=75005
+ SB=75002.5 A=0.15 P=2.3 MULT=1
MM1029 N_A_905_392#_M1024_s N_A_M1029_g N_VPWR_M1029_s VPB PSHORT L=0.15 W=1
+ AD=0.15 AS=0.182453 PD=1.3 PS=1.39151 NRD=1.9503 NRS=1.9503 M=1 R=6.66667
+ SA=75005.5 SB=75002.1 A=0.15 P=2.3 MULT=1
MM1000 N_VPWR_M1029_s N_A_219_392#_M1000_g N_X_M1000_s VPB PSHORT L=0.15 W=1.12
+ AD=0.204347 AS=0.168 PD=1.55849 PS=1.42 NRD=11.426 NRS=1.7533 M=1 R=7.46667
+ SA=75005.4 SB=75001.6 A=0.168 P=2.54 MULT=1
MM1028 N_VPWR_M1028_d N_A_219_392#_M1028_g N_X_M1000_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75005.8 SB=75001.1 A=0.168 P=2.54 MULT=1
MM1030 N_VPWR_M1028_d N_A_219_392#_M1030_g N_X_M1030_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75006.3 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1031 N_VPWR_M1031_d N_A_219_392#_M1031_g N_X_M1030_s VPB PSHORT L=0.15 W=1.12
+ AD=0.3304 AS=0.168 PD=2.83 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75006.7 SB=75000.2 A=0.168 P=2.54 MULT=1
DX32_noxref VNB VPB NWDIODE A=15.8844 P=20.8
*
.include "sky130_fd_sc_hs__maj3_4.pxi.spice"
*
.ends
*
*
