* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hs__dlrbn_2 D GATE_N RESET_B VGND VNB VPB VPWR Q Q_N
M1000 a_1446_368# a_838_48# VPWR VPB pshort w=1e+06u l=150000u
+  ad=2.95e+11p pd=2.59e+06u as=2.8377e+12p ps=2.106e+07u
M1001 a_1066_74# a_670_74# a_838_48# VNB nlowvt w=740000u l=150000u
+  ad=1.776e+11p pd=1.96e+06u as=2.109e+11p ps=2.05e+06u
M1002 VGND RESET_B a_1066_74# VNB nlowvt w=740000u l=150000u
+  ad=1.80345e+12p pd=1.499e+07u as=0p ps=0u
M1003 Q a_838_48# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.072e+11p pd=2.04e+06u as=0p ps=0u
M1004 a_592_74# a_27_112# VGND VNB nlowvt w=640000u l=150000u
+  ad=1.536e+11p pd=1.76e+06u as=0p ps=0u
M1005 a_670_74# a_230_74# a_592_74# VNB nlowvt w=640000u l=150000u
+  ad=2.44e+11p pd=2.18e+06u as=0p ps=0u
M1006 a_230_74# GATE_N VPWR VPB pshort w=840000u l=150000u
+  ad=2.478e+11p pd=2.27e+06u as=0p ps=0u
M1007 a_670_74# a_363_74# a_595_392# VPB pshort w=1e+06u l=150000u
+  ad=3.478e+11p pd=2.8e+06u as=2.4e+11p ps=2.48e+06u
M1008 Q a_838_48# VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=3.36e+11p pd=2.84e+06u as=0p ps=0u
M1009 VPWR RESET_B a_838_48# VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=3.472e+11p ps=2.86e+06u
M1010 VPWR a_838_48# Q VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VPWR a_838_48# a_783_508# VPB pshort w=420000u l=150000u
+  ad=0p pd=0u as=1.995e+11p ps=1.79e+06u
M1012 a_230_74# GATE_N VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1013 Q_N a_1446_368# VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=3.36e+11p pd=2.84e+06u as=0p ps=0u
M1014 a_595_392# a_27_112# VPWR VPB pshort w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VGND D a_27_112# VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=1.5675e+11p ps=1.67e+06u
M1016 VPWR a_1446_368# Q_N VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_790_74# a_363_74# a_670_74# VNB nlowvt w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=0p ps=0u
M1018 a_1446_368# a_838_48# VGND VNB nlowvt w=640000u l=150000u
+  ad=1.824e+11p pd=1.85e+06u as=0p ps=0u
M1019 a_838_48# a_670_74# VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 VGND a_838_48# Q VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 VGND a_1446_368# Q_N VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.368e+11p ps=2.12e+06u
M1022 VPWR D a_27_112# VPB pshort w=840000u l=150000u
+  ad=0p pd=0u as=2.478e+11p ps=2.27e+06u
M1023 VPWR a_230_74# a_363_74# VPB pshort w=840000u l=150000u
+  ad=0p pd=0u as=3.83e+11p ps=2.88e+06u
M1024 a_783_508# a_230_74# a_670_74# VPB pshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 VGND a_230_74# a_363_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1026 VGND a_838_48# a_790_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 Q_N a_1446_368# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
