* File: sky130_fd_sc_hs__and4b_2.pex.spice
* Created: Tue Sep  1 19:56:07 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HS__AND4B_2%A_N 3 5 7 8 12
c28 3 0 6.09845e-20 $X=0.495 $Y=0.835
r29 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.29
+ $Y=1.465 $X2=0.29 $Y2=1.465
r30 8 12 6.9845 $w=3.28e-07 $l=2e-07 $layer=LI1_cond $X=0.29 $Y=1.665 $X2=0.29
+ $Y2=1.465
r31 5 11 56.2063 $w=3.85e-07 $l=3.65377e-07 $layer=POLY_cond $X=0.505 $Y=1.765
+ $X2=0.36 $Y2=1.465
r32 5 7 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=0.505 $Y=1.765
+ $X2=0.505 $Y2=2.26
r33 1 11 39.305 $w=3.85e-07 $l=2.22486e-07 $layer=POLY_cond $X=0.495 $Y=1.3
+ $X2=0.36 $Y2=1.465
r34 1 3 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=0.495 $Y=1.3
+ $X2=0.495 $Y2=0.835
.ends

.subckt PM_SKY130_FD_SC_HS__AND4B_2%A_186_48# 1 2 3 12 14 16 19 21 23 27 28 29
+ 30 34 38 41 43 48
c105 29 0 1.93659e-19 $X=1.78 $Y=1.045
r106 47 48 8.15885 $w=3.84e-07 $l=6.5e-08 $layer=POLY_cond $X=1.435 $Y=1.532
+ $X2=1.5 $Y2=1.532
r107 46 47 48.3255 $w=3.84e-07 $l=3.85e-07 $layer=POLY_cond $X=1.05 $Y=1.532
+ $X2=1.435 $Y2=1.532
r108 45 46 5.64844 $w=3.84e-07 $l=4.5e-08 $layer=POLY_cond $X=1.005 $Y=1.532
+ $X2=1.05 $Y2=1.532
r109 42 48 7.53125 $w=3.84e-07 $l=6e-08 $layer=POLY_cond $X=1.56 $Y=1.532
+ $X2=1.5 $Y2=1.532
r110 41 44 8.58894 $w=3.83e-07 $l=1.65e-07 $layer=LI1_cond $X=1.587 $Y=1.465
+ $X2=1.587 $Y2=1.63
r111 41 43 8.58894 $w=3.83e-07 $l=1.65e-07 $layer=LI1_cond $X=1.587 $Y=1.465
+ $X2=1.587 $Y2=1.3
r112 41 42 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.56
+ $Y=1.465 $X2=1.56 $Y2=1.465
r113 36 38 15.5405 $w=3.28e-07 $l=4.45e-07 $layer=LI1_cond $X=3.905 $Y=0.96
+ $X2=3.905 $Y2=0.515
r114 32 34 50.938 $w=2.48e-07 $l=1.105e-06 $layer=LI1_cond $X=2.355 $Y=2.075
+ $X2=3.46 $Y2=2.075
r115 30 32 26.5062 $w=2.48e-07 $l=5.75e-07 $layer=LI1_cond $X=1.78 $Y=2.075
+ $X2=2.355 $Y2=2.075
r116 28 36 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.74 $Y=1.045
+ $X2=3.905 $Y2=0.96
r117 28 29 127.872 $w=1.68e-07 $l=1.96e-06 $layer=LI1_cond $X=3.74 $Y=1.045
+ $X2=1.78 $Y2=1.045
r118 27 30 7.14316 $w=2.5e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.695 $Y=1.95
+ $X2=1.78 $Y2=2.075
r119 27 44 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=1.695 $Y=1.95
+ $X2=1.695 $Y2=1.63
r120 24 29 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.695 $Y=1.13
+ $X2=1.78 $Y2=1.045
r121 24 43 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=1.695 $Y=1.13
+ $X2=1.695 $Y2=1.3
r122 21 48 24.8669 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=1.5 $Y=1.765
+ $X2=1.5 $Y2=1.532
r123 21 23 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.5 $Y=1.765
+ $X2=1.5 $Y2=2.4
r124 17 47 24.8669 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=1.435 $Y=1.3
+ $X2=1.435 $Y2=1.532
r125 17 19 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=1.435 $Y=1.3
+ $X2=1.435 $Y2=0.74
r126 14 46 24.8669 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=1.05 $Y=1.765
+ $X2=1.05 $Y2=1.532
r127 14 16 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.05 $Y=1.765
+ $X2=1.05 $Y2=2.4
r128 10 45 24.8669 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=1.005 $Y=1.3
+ $X2=1.005 $Y2=1.532
r129 10 12 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=1.005 $Y=1.3
+ $X2=1.005 $Y2=0.74
r130 3 34 600 $w=1.7e-07 $l=2.66786e-07 $layer=licon1_PDIFF $count=1 $X=3.29
+ $Y=1.84 $X2=3.46 $Y2=2.035
r131 2 32 600 $w=1.7e-07 $l=2.63106e-07 $layer=licon1_PDIFF $count=1 $X=2.195
+ $Y=1.84 $X2=2.355 $Y2=2.035
r132 1 38 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.765
+ $Y=0.37 $X2=3.905 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__AND4B_2%D 1 3 6 8 12
c31 1 0 1.77991e-19 $X=2.12 $Y=1.765
r32 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.13
+ $Y=1.515 $X2=2.13 $Y2=1.515
r33 8 12 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=2.13 $Y=1.665
+ $X2=2.13 $Y2=1.515
r34 4 11 38.5562 $w=2.99e-07 $l=2.05122e-07 $layer=POLY_cond $X=2.22 $Y=1.35
+ $X2=2.13 $Y2=1.515
r35 4 6 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.22 $Y=1.35 $X2=2.22
+ $Y2=0.74
r36 1 11 52.2586 $w=2.99e-07 $l=2.54951e-07 $layer=POLY_cond $X=2.12 $Y=1.765
+ $X2=2.13 $Y2=1.515
r37 1 3 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=2.12 $Y=1.765
+ $X2=2.12 $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_HS__AND4B_2%C 1 3 6 8 12
r27 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.67
+ $Y=1.515 $X2=2.67 $Y2=1.515
r28 8 12 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=2.67 $Y=1.665
+ $X2=2.67 $Y2=1.515
r29 4 11 38.5562 $w=2.99e-07 $l=1.92678e-07 $layer=POLY_cond $X=2.61 $Y=1.35
+ $X2=2.67 $Y2=1.515
r30 4 6 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.61 $Y=1.35 $X2=2.61
+ $Y2=0.74
r31 1 11 52.2586 $w=2.99e-07 $l=2.85044e-07 $layer=POLY_cond $X=2.595 $Y=1.765
+ $X2=2.67 $Y2=1.515
r32 1 3 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=2.595 $Y=1.765
+ $X2=2.595 $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_HS__AND4B_2%B 3 5 7 8 12
r28 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.24
+ $Y=1.515 $X2=3.24 $Y2=1.515
r29 8 12 4.32166 $w=3.98e-07 $l=1.5e-07 $layer=LI1_cond $X=3.205 $Y=1.665
+ $X2=3.205 $Y2=1.515
r30 5 11 52.2586 $w=2.99e-07 $l=2.62202e-07 $layer=POLY_cond $X=3.215 $Y=1.765
+ $X2=3.24 $Y2=1.515
r31 5 7 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=3.215 $Y=1.765
+ $X2=3.215 $Y2=2.34
r32 1 11 38.5562 $w=2.99e-07 $l=2.05122e-07 $layer=POLY_cond $X=3.15 $Y=1.35
+ $X2=3.24 $Y2=1.515
r33 1 3 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=3.15 $Y=1.35 $X2=3.15
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HS__AND4B_2%A_27_112# 1 2 9 11 13 16 18 19 21 22 25 27
+ 33
r83 30 33 4.1907 $w=3.28e-07 $l=1.2e-07 $layer=LI1_cond $X=3.78 $Y=1.515 $X2=3.9
+ $Y2=1.515
r84 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.78
+ $Y=1.515 $X2=3.78 $Y2=1.515
r85 27 28 6.8562 $w=6.05e-07 $l=3.4e-07 $layer=LI1_cond $X=0.455 $Y=2.115
+ $X2=0.455 $Y2=2.455
r86 24 33 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.9 $Y=1.68 $X2=3.9
+ $Y2=1.515
r87 24 25 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=3.9 $Y=1.68 $X2=3.9
+ $Y2=2.37
r88 23 28 8.37032 $w=1.7e-07 $l=3.4e-07 $layer=LI1_cond $X=0.795 $Y=2.455
+ $X2=0.455 $Y2=2.455
r89 22 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.815 $Y=2.455
+ $X2=3.9 $Y2=2.37
r90 22 23 197.027 $w=1.68e-07 $l=3.02e-06 $layer=LI1_cond $X=3.815 $Y=2.455
+ $X2=0.795 $Y2=2.455
r91 21 27 10.3924 $w=6.05e-07 $l=3.27261e-07 $layer=LI1_cond $X=0.71 $Y=1.95
+ $X2=0.455 $Y2=2.115
r92 20 21 53.4973 $w=1.68e-07 $l=8.2e-07 $layer=LI1_cond $X=0.71 $Y=1.13
+ $X2=0.71 $Y2=1.95
r93 18 20 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.625 $Y=1.045
+ $X2=0.71 $Y2=1.13
r94 18 19 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=0.625 $Y=1.045
+ $X2=0.445 $Y2=1.045
r95 14 19 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.28 $Y=0.96
+ $X2=0.445 $Y2=1.045
r96 14 16 4.36531 $w=3.28e-07 $l=1.25e-07 $layer=LI1_cond $X=0.28 $Y=0.96
+ $X2=0.28 $Y2=0.835
r97 11 31 52.2586 $w=2.99e-07 $l=2.85044e-07 $layer=POLY_cond $X=3.705 $Y=1.765
+ $X2=3.78 $Y2=1.515
r98 11 13 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=3.705 $Y=1.765
+ $X2=3.705 $Y2=2.34
r99 7 31 38.5562 $w=2.99e-07 $l=2.05122e-07 $layer=POLY_cond $X=3.69 $Y=1.35
+ $X2=3.78 $Y2=1.515
r100 7 9 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=3.69 $Y=1.35 $X2=3.69
+ $Y2=0.74
r101 2 27 300 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.115
r102 1 16 182 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.56 $X2=0.28 $Y2=0.835
.ends

.subckt PM_SKY130_FD_SC_HS__AND4B_2%VPWR 1 2 3 4 17 19 23 27 29 31 34 35 36 42
+ 47 50 54
r54 53 54 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r55 50 51 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r56 48 51 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.68 $Y2=3.33
r57 47 48 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r58 45 54 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.08 $Y2=3.33
r59 44 45 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r60 42 53 4.96106 $w=1.7e-07 $l=2.35e-07 $layer=LI1_cond $X=3.85 $Y=3.33
+ $X2=4.085 $Y2=3.33
r61 42 44 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=3.85 $Y=3.33 $X2=3.6
+ $Y2=3.33
r62 41 45 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.6 $Y2=3.33
r63 40 41 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r64 38 50 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.975 $Y=3.33
+ $X2=1.81 $Y2=3.33
r65 38 40 43.385 $w=1.68e-07 $l=6.65e-07 $layer=LI1_cond $X=1.975 $Y=3.33
+ $X2=2.64 $Y2=3.33
r66 36 41 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r67 36 51 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.68 $Y2=3.33
r68 34 40 6.52406 $w=1.68e-07 $l=1e-07 $layer=LI1_cond $X=2.74 $Y=3.33 $X2=2.64
+ $Y2=3.33
r69 34 35 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.74 $Y=3.33
+ $X2=2.905 $Y2=3.33
r70 33 44 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=3.07 $Y=3.33 $X2=3.6
+ $Y2=3.33
r71 33 35 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.07 $Y=3.33
+ $X2=2.905 $Y2=3.33
r72 29 53 3.01886 $w=3.55e-07 $l=1.1025e-07 $layer=LI1_cond $X=4.027 $Y=3.245
+ $X2=4.085 $Y2=3.33
r73 29 31 14.2838 $w=3.53e-07 $l=4.4e-07 $layer=LI1_cond $X=4.027 $Y=3.245
+ $X2=4.027 $Y2=2.805
r74 25 35 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.905 $Y=3.245
+ $X2=2.905 $Y2=3.33
r75 25 27 15.3659 $w=3.28e-07 $l=4.4e-07 $layer=LI1_cond $X=2.905 $Y=3.245
+ $X2=2.905 $Y2=2.805
r76 21 50 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.81 $Y=3.245
+ $X2=1.81 $Y2=3.33
r77 21 23 15.3659 $w=3.28e-07 $l=4.4e-07 $layer=LI1_cond $X=1.81 $Y=3.245
+ $X2=1.81 $Y2=2.805
r78 20 47 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.98 $Y=3.33
+ $X2=0.815 $Y2=3.33
r79 19 50 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.645 $Y=3.33
+ $X2=1.81 $Y2=3.33
r80 19 20 43.385 $w=1.68e-07 $l=6.65e-07 $layer=LI1_cond $X=1.645 $Y=3.33
+ $X2=0.98 $Y2=3.33
r81 15 47 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.815 $Y=3.245
+ $X2=0.815 $Y2=3.33
r82 15 17 15.3659 $w=3.28e-07 $l=4.4e-07 $layer=LI1_cond $X=0.815 $Y=3.245
+ $X2=0.815 $Y2=2.805
r83 4 31 600 $w=1.7e-07 $l=1.08058e-06 $layer=licon1_PDIFF $count=1 $X=3.78
+ $Y=1.84 $X2=4.025 $Y2=2.805
r84 3 27 600 $w=1.7e-07 $l=1.0761e-06 $layer=licon1_PDIFF $count=1 $X=2.67
+ $Y=1.84 $X2=2.905 $Y2=2.805
r85 2 23 600 $w=1.7e-07 $l=1.0761e-06 $layer=licon1_PDIFF $count=1 $X=1.575
+ $Y=1.84 $X2=1.81 $Y2=2.805
r86 1 17 600 $w=1.7e-07 $l=1.0761e-06 $layer=licon1_PDIFF $count=1 $X=0.58
+ $Y=1.84 $X2=0.815 $Y2=2.805
.ends

.subckt PM_SKY130_FD_SC_HS__AND4B_2%X 1 2 9 12 13 14
c37 14 0 1.77991e-19 $X=1.2 $Y=2.035
c38 13 0 6.09845e-20 $X=1.22 $Y=1.13
r39 14 16 1.81965 $w=3.78e-07 $l=6e-08 $layer=LI1_cond $X=1.2 $Y=2.01 $X2=1.14
+ $Y2=2.01
r40 12 16 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.14 $Y=1.82 $X2=1.14
+ $Y2=2.01
r41 12 13 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.14 $Y=1.82 $X2=1.14
+ $Y2=1.13
r42 7 13 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=1.22 $Y=0.965
+ $X2=1.22 $Y2=1.13
r43 7 9 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=1.22 $Y=0.965 $X2=1.22
+ $Y2=0.515
r44 2 14 600 $w=1.7e-07 $l=2.33238e-07 $layer=licon1_PDIFF $count=1 $X=1.125
+ $Y=1.84 $X2=1.275 $Y2=2.01
r45 1 9 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.08
+ $Y=0.37 $X2=1.22 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__AND4B_2%VGND 1 2 9 13 15 17 22 29 30 33 36
r44 36 39 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r45 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r46 29 30 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r47 27 36 12.6759 $w=1.7e-07 $l=3.05e-07 $layer=LI1_cond $X=2.165 $Y=0 $X2=1.86
+ $Y2=0
r48 27 29 124.936 $w=1.68e-07 $l=1.915e-06 $layer=LI1_cond $X=2.165 $Y=0
+ $X2=4.08 $Y2=0
r49 26 39 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=1.68
+ $Y2=0
r50 26 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r51 25 26 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r52 23 33 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.875 $Y=0 $X2=0.75
+ $Y2=0
r53 23 25 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.875 $Y=0 $X2=1.2
+ $Y2=0
r54 22 36 12.6759 $w=1.7e-07 $l=3.05e-07 $layer=LI1_cond $X=1.555 $Y=0 $X2=1.86
+ $Y2=0
r55 22 25 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=1.555 $Y=0 $X2=1.2
+ $Y2=0
r56 20 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r57 19 20 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r58 17 33 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.625 $Y=0 $X2=0.75
+ $Y2=0
r59 17 19 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=0.625 $Y=0 $X2=0.24
+ $Y2=0
r60 15 30 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=2.16 $Y=0 $X2=4.08
+ $Y2=0
r61 15 39 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.68
+ $Y2=0
r62 15 36 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r63 11 36 2.55884 $w=6.1e-07 $l=8.5e-08 $layer=LI1_cond $X=1.86 $Y=0.085
+ $X2=1.86 $Y2=0
r64 11 13 10.5882 $w=6.08e-07 $l=5.4e-07 $layer=LI1_cond $X=1.86 $Y=0.085
+ $X2=1.86 $Y2=0.625
r65 7 33 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.75 $Y=0.085
+ $X2=0.75 $Y2=0
r66 7 9 24.8928 $w=2.48e-07 $l=5.4e-07 $layer=LI1_cond $X=0.75 $Y=0.085 $X2=0.75
+ $Y2=0.625
r67 2 13 91 $w=1.7e-07 $l=6.09303e-07 $layer=licon1_NDIFF $count=2 $X=1.51
+ $Y=0.37 $X2=2.005 $Y2=0.625
r68 1 9 182 $w=1.7e-07 $l=2.504e-07 $layer=licon1_NDIFF $count=1 $X=0.57 $Y=0.56
+ $X2=0.79 $Y2=0.625
.ends

