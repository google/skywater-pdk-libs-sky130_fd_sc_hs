# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_hs__xnor3_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__xnor3_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  8.640000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.955000 1.375000 1.315000 1.780000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.693000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.735000 1.350000 4.405000 1.780000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.381000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.845000 1.350000 7.175000 1.780000 ;
    END
  END C
  PIN X
    ANTENNADIFFAREA  0.543200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.750000 1.840000 8.095000 2.980000 ;
        RECT 7.765000 0.440000 8.095000 1.170000 ;
        RECT 7.925000 1.170000 8.095000 1.840000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 8.640000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 8.640000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 8.640000 0.085000 ;
      RECT 0.000000  3.245000 8.640000 3.415000 ;
      RECT 0.085000  0.385000 0.405000 1.065000 ;
      RECT 0.085000  1.065000 0.325000 2.290000 ;
      RECT 0.085000  2.290000 0.445000 2.885000 ;
      RECT 0.495000  1.235000 0.745000 1.950000 ;
      RECT 0.495000  1.950000 1.375000 2.120000 ;
      RECT 0.575000  1.035000 1.345000 1.205000 ;
      RECT 0.575000  1.205000 0.745000 1.235000 ;
      RECT 0.585000  0.085000 0.915000 0.865000 ;
      RECT 0.645000  2.305000 0.925000 3.245000 ;
      RECT 1.095000  0.255000 3.530000 0.425000 ;
      RECT 1.095000  0.425000 1.345000 1.035000 ;
      RECT 1.095000  2.120000 1.375000 2.905000 ;
      RECT 1.095000  2.905000 3.675000 3.075000 ;
      RECT 1.545000  1.165000 2.385000 1.380000 ;
      RECT 1.545000  1.380000 1.715000 2.565000 ;
      RECT 1.545000  2.565000 2.605000 2.735000 ;
      RECT 1.625000  0.595000 2.725000 0.615000 ;
      RECT 1.625000  0.615000 5.160000 0.765000 ;
      RECT 1.625000  0.765000 1.955000 0.995000 ;
      RECT 1.885000  1.550000 2.755000 1.720000 ;
      RECT 1.885000  1.720000 2.105000 2.395000 ;
      RECT 2.135000  0.935000 2.385000 1.165000 ;
      RECT 2.275000  1.890000 2.605000 2.565000 ;
      RECT 2.555000  0.765000 5.160000 0.785000 ;
      RECT 2.555000  0.955000 2.985000 1.285000 ;
      RECT 2.555000  1.285000 2.755000 1.550000 ;
      RECT 2.835000  1.875000 3.145000 2.370000 ;
      RECT 2.835000  2.370000 4.755000 2.395000 ;
      RECT 2.835000  2.395000 6.320000 2.540000 ;
      RECT 2.835000  2.540000 3.065000 2.620000 ;
      RECT 3.155000  1.375000 3.565000 1.705000 ;
      RECT 3.200000  0.425000 3.530000 0.445000 ;
      RECT 3.345000  2.710000 3.675000 2.905000 ;
      RECT 3.395000  0.955000 4.090000 1.125000 ;
      RECT 3.395000  1.125000 3.565000 1.375000 ;
      RECT 3.395000  1.705000 3.565000 1.950000 ;
      RECT 3.395000  1.950000 4.255000 2.200000 ;
      RECT 4.270000  0.085000 4.600000 0.445000 ;
      RECT 4.455000  2.735000 4.785000 3.245000 ;
      RECT 4.585000  0.785000 5.160000 0.965000 ;
      RECT 4.585000  0.965000 4.755000 2.370000 ;
      RECT 4.585000  2.540000 6.320000 2.565000 ;
      RECT 4.830000  0.350000 5.160000 0.615000 ;
      RECT 4.925000  1.135000 6.160000 1.305000 ;
      RECT 4.925000  1.305000 5.155000 1.975000 ;
      RECT 4.925000  1.975000 5.335000 2.225000 ;
      RECT 5.325000  1.475000 6.675000 1.805000 ;
      RECT 5.330000  0.255000 6.500000 0.425000 ;
      RECT 5.330000  0.425000 5.660000 0.965000 ;
      RECT 5.535000  2.735000 5.865000 2.905000 ;
      RECT 5.535000  2.905000 7.210000 3.075000 ;
      RECT 5.830000  0.595000 6.160000 1.135000 ;
      RECT 6.070000  1.975000 6.320000 2.395000 ;
      RECT 6.070000  2.565000 6.320000 2.735000 ;
      RECT 6.330000  0.425000 6.500000 0.660000 ;
      RECT 6.330000  0.660000 7.060000 0.830000 ;
      RECT 6.390000  1.000000 6.720000 1.170000 ;
      RECT 6.390000  1.170000 6.675000 1.475000 ;
      RECT 6.505000  1.805000 6.675000 1.950000 ;
      RECT 6.505000  1.950000 6.870000 2.500000 ;
      RECT 6.890000  0.830000 7.060000 1.010000 ;
      RECT 6.890000  1.010000 7.580000 1.180000 ;
      RECT 6.900000  0.085000 7.585000 0.490000 ;
      RECT 7.040000  1.950000 7.580000 2.120000 ;
      RECT 7.040000  2.120000 7.210000 2.905000 ;
      RECT 7.230000  0.490000 7.585000 0.840000 ;
      RECT 7.380000  2.290000 7.550000 3.245000 ;
      RECT 7.410000  1.180000 7.580000 1.340000 ;
      RECT 7.410000  1.340000 7.755000 1.670000 ;
      RECT 7.410000  1.670000 7.580000 1.950000 ;
      RECT 8.275000  0.085000 8.525000 1.250000 ;
      RECT 8.280000  1.820000 8.530000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  1.210000 0.325000 1.380000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  1.210000 1.765000 1.380000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  1.210000 2.725000 1.380000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  1.210000 5.125000 1.380000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
      RECT 7.835000 -0.085000 8.005000 0.085000 ;
      RECT 7.835000  3.245000 8.005000 3.415000 ;
      RECT 8.315000 -0.085000 8.485000 0.085000 ;
      RECT 8.315000  3.245000 8.485000 3.415000 ;
    LAYER met1 ;
      RECT 0.095000 1.180000 0.385000 1.225000 ;
      RECT 0.095000 1.225000 1.825000 1.365000 ;
      RECT 0.095000 1.365000 0.385000 1.410000 ;
      RECT 1.535000 1.180000 1.825000 1.225000 ;
      RECT 1.535000 1.365000 1.825000 1.410000 ;
      RECT 2.495000 1.180000 2.785000 1.225000 ;
      RECT 2.495000 1.225000 5.185000 1.365000 ;
      RECT 2.495000 1.365000 2.785000 1.410000 ;
      RECT 4.895000 1.180000 5.185000 1.225000 ;
      RECT 4.895000 1.365000 5.185000 1.410000 ;
  END
END sky130_fd_sc_hs__xnor3_2
END LIBRARY
