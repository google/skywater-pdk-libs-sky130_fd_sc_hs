* File: sky130_fd_sc_hs__nor2_4.pex.spice
* Created: Thu Aug 27 20:53:12 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HS__NOR2_4%A 1 3 4 6 7 9 10 12 13 15 16 18 19 20 21 22
+ 37
c69 37 0 3.08465e-20 $X=1.81 $Y=1.492
c70 16 0 6.46447e-20 $X=1.855 $Y=1.765
r71 37 38 5.11557 $w=4.24e-07 $l=4.5e-08 $layer=POLY_cond $X=1.81 $Y=1.492
+ $X2=1.855 $Y2=1.492
r72 35 37 20.4623 $w=4.24e-07 $l=1.8e-07 $layer=POLY_cond $X=1.63 $Y=1.492
+ $X2=1.81 $Y2=1.492
r73 35 36 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.63
+ $Y=1.385 $X2=1.63 $Y2=1.385
r74 33 35 25.5778 $w=4.24e-07 $l=2.25e-07 $layer=POLY_cond $X=1.405 $Y=1.492
+ $X2=1.63 $Y2=1.492
r75 32 33 51.1557 $w=4.24e-07 $l=4.5e-07 $layer=POLY_cond $X=0.955 $Y=1.492
+ $X2=1.405 $Y2=1.492
r76 30 32 39.2193 $w=4.24e-07 $l=3.45e-07 $layer=POLY_cond $X=0.61 $Y=1.492
+ $X2=0.955 $Y2=1.492
r77 30 31 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.61
+ $Y=1.385 $X2=0.61 $Y2=1.385
r78 28 30 10.2311 $w=4.24e-07 $l=9e-08 $layer=POLY_cond $X=0.52 $Y=1.492
+ $X2=0.61 $Y2=1.492
r79 27 28 1.70519 $w=4.24e-07 $l=1.5e-08 $layer=POLY_cond $X=0.505 $Y=1.492
+ $X2=0.52 $Y2=1.492
r80 22 36 1.55736 $w=3.68e-07 $l=5e-08 $layer=LI1_cond $X=1.68 $Y=1.365 $X2=1.63
+ $Y2=1.365
r81 21 36 13.3933 $w=3.68e-07 $l=4.3e-07 $layer=LI1_cond $X=1.2 $Y=1.365
+ $X2=1.63 $Y2=1.365
r82 20 21 14.9506 $w=3.68e-07 $l=4.8e-07 $layer=LI1_cond $X=0.72 $Y=1.365
+ $X2=1.2 $Y2=1.365
r83 20 31 3.42618 $w=3.68e-07 $l=1.1e-07 $layer=LI1_cond $X=0.72 $Y=1.365
+ $X2=0.61 $Y2=1.365
r84 19 31 11.5244 $w=3.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.24 $Y=1.365
+ $X2=0.61 $Y2=1.365
r85 16 38 27.2926 $w=1.5e-07 $l=2.73e-07 $layer=POLY_cond $X=1.855 $Y=1.765
+ $X2=1.855 $Y2=1.492
r86 16 18 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.855 $Y=1.765
+ $X2=1.855 $Y2=2.4
r87 13 37 27.2926 $w=1.5e-07 $l=2.72e-07 $layer=POLY_cond $X=1.81 $Y=1.22
+ $X2=1.81 $Y2=1.492
r88 13 15 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.81 $Y=1.22 $X2=1.81
+ $Y2=0.74
r89 10 33 27.2926 $w=1.5e-07 $l=2.73e-07 $layer=POLY_cond $X=1.405 $Y=1.765
+ $X2=1.405 $Y2=1.492
r90 10 12 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.405 $Y=1.765
+ $X2=1.405 $Y2=2.4
r91 7 32 27.2926 $w=1.5e-07 $l=2.73e-07 $layer=POLY_cond $X=0.955 $Y=1.765
+ $X2=0.955 $Y2=1.492
r92 7 9 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.955 $Y=1.765
+ $X2=0.955 $Y2=2.4
r93 4 28 27.2926 $w=1.5e-07 $l=2.72e-07 $layer=POLY_cond $X=0.52 $Y=1.22
+ $X2=0.52 $Y2=1.492
r94 4 6 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=0.52 $Y=1.22 $X2=0.52
+ $Y2=0.74
r95 1 27 27.2926 $w=1.5e-07 $l=2.73e-07 $layer=POLY_cond $X=0.505 $Y=1.765
+ $X2=0.505 $Y2=1.492
r96 1 3 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.505 $Y=1.765
+ $X2=0.505 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_HS__NOR2_4%B 1 3 4 6 7 9 10 12 13 15 16 18 19 20 21 33
r62 35 36 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=4.01
+ $Y=1.385 $X2=4.01 $Y2=1.385
r63 33 35 30.125 $w=4.08e-07 $l=2.55e-07 $layer=POLY_cond $X=3.755 $Y=1.492
+ $X2=4.01 $Y2=1.492
r64 31 33 50.2083 $w=4.08e-07 $l=4.25e-07 $layer=POLY_cond $X=3.33 $Y=1.492
+ $X2=3.755 $Y2=1.492
r65 31 32 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=3.33
+ $Y=1.385 $X2=3.33 $Y2=1.385
r66 29 31 8.86029 $w=4.08e-07 $l=7.5e-08 $layer=POLY_cond $X=3.255 $Y=1.492
+ $X2=3.33 $Y2=1.492
r67 28 29 59.0686 $w=4.08e-07 $l=5e-07 $layer=POLY_cond $X=2.755 $Y=1.492
+ $X2=3.255 $Y2=1.492
r68 27 28 1.77206 $w=4.08e-07 $l=1.5e-08 $layer=POLY_cond $X=2.74 $Y=1.492
+ $X2=2.755 $Y2=1.492
r69 26 27 51.3897 $w=4.08e-07 $l=4.35e-07 $layer=POLY_cond $X=2.305 $Y=1.492
+ $X2=2.74 $Y2=1.492
r70 25 26 1.77206 $w=4.08e-07 $l=1.5e-08 $layer=POLY_cond $X=2.29 $Y=1.492
+ $X2=2.305 $Y2=1.492
r71 21 36 2.1803 $w=3.68e-07 $l=7e-08 $layer=LI1_cond $X=4.08 $Y=1.365 $X2=4.01
+ $Y2=1.365
r72 20 36 12.7703 $w=3.68e-07 $l=4.1e-07 $layer=LI1_cond $X=3.6 $Y=1.365
+ $X2=4.01 $Y2=1.365
r73 20 32 8.40972 $w=3.68e-07 $l=2.7e-07 $layer=LI1_cond $X=3.6 $Y=1.365
+ $X2=3.33 $Y2=1.365
r74 19 32 6.54089 $w=3.68e-07 $l=2.1e-07 $layer=LI1_cond $X=3.12 $Y=1.365
+ $X2=3.33 $Y2=1.365
r75 16 33 26.3468 $w=1.5e-07 $l=2.73e-07 $layer=POLY_cond $X=3.755 $Y=1.765
+ $X2=3.755 $Y2=1.492
r76 16 18 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.755 $Y=1.765
+ $X2=3.755 $Y2=2.4
r77 13 29 26.3468 $w=1.5e-07 $l=2.73e-07 $layer=POLY_cond $X=3.255 $Y=1.765
+ $X2=3.255 $Y2=1.492
r78 13 15 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.255 $Y=1.765
+ $X2=3.255 $Y2=2.4
r79 10 28 26.3468 $w=1.5e-07 $l=2.73e-07 $layer=POLY_cond $X=2.755 $Y=1.765
+ $X2=2.755 $Y2=1.492
r80 10 12 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.755 $Y=1.765
+ $X2=2.755 $Y2=2.4
r81 7 27 26.3468 $w=1.5e-07 $l=2.72e-07 $layer=POLY_cond $X=2.74 $Y=1.22
+ $X2=2.74 $Y2=1.492
r82 7 9 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=2.74 $Y=1.22 $X2=2.74
+ $Y2=0.74
r83 4 26 26.3468 $w=1.5e-07 $l=2.73e-07 $layer=POLY_cond $X=2.305 $Y=1.765
+ $X2=2.305 $Y2=1.492
r84 4 6 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.305 $Y=1.765
+ $X2=2.305 $Y2=2.4
r85 1 25 26.3468 $w=1.5e-07 $l=2.72e-07 $layer=POLY_cond $X=2.29 $Y=1.22
+ $X2=2.29 $Y2=1.492
r86 1 3 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=2.29 $Y=1.22 $X2=2.29
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HS__NOR2_4%A_27_368# 1 2 3 4 5 18 22 23 26 30 35 38 39
+ 42 46 50 54 55
r76 50 53 34.1617 $w=2.78e-07 $l=8.3e-07 $layer=LI1_cond $X=4.005 $Y=1.985
+ $X2=4.005 $Y2=2.815
r77 48 53 3.70428 $w=2.78e-07 $l=9e-08 $layer=LI1_cond $X=4.005 $Y=2.905
+ $X2=4.005 $Y2=2.815
r78 47 55 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.195 $Y=2.99
+ $X2=3.03 $Y2=2.99
r79 46 48 7.36005 $w=1.7e-07 $l=1.77482e-07 $layer=LI1_cond $X=3.865 $Y=2.99
+ $X2=4.005 $Y2=2.905
r80 46 47 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.865 $Y=2.99
+ $X2=3.195 $Y2=2.99
r81 42 45 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=3.03 $Y=2.145
+ $X2=3.03 $Y2=2.825
r82 40 55 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.03 $Y=2.905
+ $X2=3.03 $Y2=2.99
r83 40 45 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=3.03 $Y=2.905 $X2=3.03
+ $Y2=2.825
r84 38 55 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.865 $Y=2.99
+ $X2=3.03 $Y2=2.99
r85 38 39 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.865 $Y=2.99
+ $X2=2.195 $Y2=2.99
r86 35 37 34.1617 $w=2.78e-07 $l=8.3e-07 $layer=LI1_cond $X=2.055 $Y=1.985
+ $X2=2.055 $Y2=2.815
r87 33 39 7.36005 $w=1.7e-07 $l=1.77482e-07 $layer=LI1_cond $X=2.055 $Y=2.905
+ $X2=2.195 $Y2=2.99
r88 33 37 3.70428 $w=2.78e-07 $l=9e-08 $layer=LI1_cond $X=2.055 $Y=2.905
+ $X2=2.055 $Y2=2.815
r89 32 35 3.91007 $w=2.78e-07 $l=9.5e-08 $layer=LI1_cond $X=2.055 $Y=1.89
+ $X2=2.055 $Y2=1.985
r90 31 54 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.345 $Y=1.805
+ $X2=1.18 $Y2=1.805
r91 30 32 7.36005 $w=1.7e-07 $l=1.77482e-07 $layer=LI1_cond $X=1.915 $Y=1.805
+ $X2=2.055 $Y2=1.89
r92 30 31 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=1.915 $Y=1.805
+ $X2=1.345 $Y2=1.805
r93 26 28 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=1.18 $Y=1.985
+ $X2=1.18 $Y2=2.815
r94 24 54 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.18 $Y=1.89 $X2=1.18
+ $Y2=1.805
r95 24 26 3.31764 $w=3.28e-07 $l=9.5e-08 $layer=LI1_cond $X=1.18 $Y=1.89
+ $X2=1.18 $Y2=1.985
r96 22 54 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.015 $Y=1.805
+ $X2=1.18 $Y2=1.805
r97 22 23 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=1.015 $Y=1.805
+ $X2=0.445 $Y2=1.805
r98 18 20 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=0.28 $Y=1.985
+ $X2=0.28 $Y2=2.815
r99 16 23 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.28 $Y=1.89
+ $X2=0.445 $Y2=1.805
r100 16 18 3.31764 $w=3.28e-07 $l=9.5e-08 $layer=LI1_cond $X=0.28 $Y=1.89
+ $X2=0.28 $Y2=1.985
r101 5 53 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=3.83
+ $Y=1.84 $X2=3.98 $Y2=2.815
r102 5 50 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=3.83
+ $Y=1.84 $X2=3.98 $Y2=1.985
r103 4 45 400 $w=1.7e-07 $l=1.08038e-06 $layer=licon1_PDIFF $count=1 $X=2.83
+ $Y=1.84 $X2=3.03 $Y2=2.825
r104 4 42 400 $w=1.7e-07 $l=3.9246e-07 $layer=licon1_PDIFF $count=1 $X=2.83
+ $Y=1.84 $X2=3.03 $Y2=2.145
r105 3 37 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=1.93
+ $Y=1.84 $X2=2.08 $Y2=2.815
r106 3 35 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=1.93
+ $Y=1.84 $X2=2.08 $Y2=1.985
r107 2 28 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=1.03
+ $Y=1.84 $X2=1.18 $Y2=2.815
r108 2 26 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=1.03
+ $Y=1.84 $X2=1.18 $Y2=1.985
r109 1 20 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.815
r110 1 18 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HS__NOR2_4%VPWR 1 2 11 15 17 19 26 27 30 33
r49 33 34 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r50 30 31 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r51 26 27 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r52 24 33 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.715 $Y=3.33
+ $X2=1.63 $Y2=3.33
r53 24 26 154.294 $w=1.68e-07 $l=2.365e-06 $layer=LI1_cond $X=1.715 $Y=3.33
+ $X2=4.08 $Y2=3.33
r54 23 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=1.68 $Y2=3.33
r55 23 31 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r56 22 23 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r57 20 30 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.815 $Y=3.33
+ $X2=0.73 $Y2=3.33
r58 20 22 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=0.815 $Y=3.33
+ $X2=1.2 $Y2=3.33
r59 19 33 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.545 $Y=3.33
+ $X2=1.63 $Y2=3.33
r60 19 22 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.545 $Y=3.33
+ $X2=1.2 $Y2=3.33
r61 17 27 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=4.08 $Y2=3.33
r62 17 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.68 $Y2=3.33
r63 13 33 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.63 $Y=3.245
+ $X2=1.63 $Y2=3.33
r64 13 15 66.5455 $w=1.68e-07 $l=1.02e-06 $layer=LI1_cond $X=1.63 $Y=3.245
+ $X2=1.63 $Y2=2.225
r65 9 30 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.73 $Y=3.245 $X2=0.73
+ $Y2=3.33
r66 9 11 66.5455 $w=1.68e-07 $l=1.02e-06 $layer=LI1_cond $X=0.73 $Y=3.245
+ $X2=0.73 $Y2=2.225
r67 2 15 300 $w=1.7e-07 $l=4.53845e-07 $layer=licon1_PDIFF $count=2 $X=1.48
+ $Y=1.84 $X2=1.63 $Y2=2.225
r68 1 11 300 $w=1.7e-07 $l=4.53845e-07 $layer=licon1_PDIFF $count=2 $X=0.58
+ $Y=1.84 $X2=0.73 $Y2=2.225
.ends

.subckt PM_SKY130_FD_SC_HS__NOR2_4%Y 1 2 3 4 13 17 21 23 24 27 31 35 41 42 43
c57 42 0 9.54912e-20 $X=2.53 $Y=1.805
r58 43 45 12.7875 $w=3.53e-07 $l=3.7e-07 $layer=LI1_cond $X=2.557 $Y=1.295
+ $X2=2.557 $Y2=0.925
r59 40 41 9.36207 $w=6.68e-07 $l=9.5e-08 $layer=LI1_cond $X=1.595 $Y=0.675
+ $X2=1.69 $Y2=0.675
r60 35 37 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=3.53 $Y=1.97
+ $X2=3.53 $Y2=2.65
r61 33 35 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=3.53 $Y=1.89 $X2=3.53
+ $Y2=1.97
r62 32 42 3.80956 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.695 $Y=1.805
+ $X2=2.53 $Y2=1.805
r63 31 33 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.365 $Y=1.805
+ $X2=3.53 $Y2=1.89
r64 31 32 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.365 $Y=1.805
+ $X2=2.695 $Y2=1.805
r65 27 29 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=2.53 $Y=1.97
+ $X2=2.53 $Y2=2.65
r66 25 42 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.53 $Y=1.89 $X2=2.53
+ $Y2=1.805
r67 25 27 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=2.53 $Y=1.89 $X2=2.53
+ $Y2=1.97
r68 24 42 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.53 $Y=1.72 $X2=2.53
+ $Y2=1.805
r69 23 43 4.04312 $w=3.53e-07 $l=1.27789e-07 $layer=LI1_cond $X=2.53 $Y=1.41
+ $X2=2.557 $Y2=1.295
r70 23 24 10.826 $w=3.28e-07 $l=3.1e-07 $layer=LI1_cond $X=2.53 $Y=1.41 $X2=2.53
+ $Y2=1.72
r71 19 45 3.00629 $w=3.53e-07 $l=9.97246e-08 $layer=LI1_cond $X=2.525 $Y=0.84
+ $X2=2.557 $Y2=0.925
r72 19 21 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=2.525 $Y=0.84
+ $X2=2.525 $Y2=0.515
r73 17 45 5.025 $w=1.7e-07 $l=1.97e-07 $layer=LI1_cond $X=2.36 $Y=0.925
+ $X2=2.557 $Y2=0.925
r74 17 41 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.36 $Y=0.925
+ $X2=1.69 $Y2=0.925
r75 13 40 4.28446 $w=6.68e-07 $l=2.4e-07 $layer=LI1_cond $X=1.355 $Y=0.675
+ $X2=1.595 $Y2=0.675
r76 13 15 3.65964 $w=6.68e-07 $l=2.05e-07 $layer=LI1_cond $X=1.355 $Y=0.675
+ $X2=1.15 $Y2=0.675
r77 4 37 400 $w=1.7e-07 $l=9.04489e-07 $layer=licon1_PDIFF $count=1 $X=3.33
+ $Y=1.84 $X2=3.53 $Y2=2.65
r78 4 35 400 $w=1.7e-07 $l=2.56905e-07 $layer=licon1_PDIFF $count=1 $X=3.33
+ $Y=1.84 $X2=3.53 $Y2=1.97
r79 3 29 400 $w=1.7e-07 $l=8.81816e-07 $layer=licon1_PDIFF $count=1 $X=2.38
+ $Y=1.84 $X2=2.53 $Y2=2.65
r80 3 27 400 $w=1.7e-07 $l=2.04939e-07 $layer=licon1_PDIFF $count=1 $X=2.38
+ $Y=1.84 $X2=2.53 $Y2=1.97
r81 2 21 91 $w=1.7e-07 $l=2.20907e-07 $layer=licon1_NDIFF $count=2 $X=2.365
+ $Y=0.37 $X2=2.525 $Y2=0.515
r82 1 40 91 $w=1.7e-07 $l=1.06536e-06 $layer=licon1_NDIFF $count=2 $X=0.595
+ $Y=0.37 $X2=1.595 $Y2=0.505
r83 1 15 45.5 $w=1.7e-07 $l=6.1883e-07 $layer=licon1_NDIFF $count=4 $X=0.595
+ $Y=0.37 $X2=1.15 $Y2=0.505
.ends

.subckt PM_SKY130_FD_SC_HS__NOR2_4%VGND 1 2 3 10 12 16 19 20 21 30 43 46
r34 45 46 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r35 43 45 0.477495 $w=1.022e-06 $l=4e-08 $layer=LI1_cond $X=4.04 $Y=0.462
+ $X2=4.08 $Y2=0.462
r36 41 46 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=4.08
+ $Y2=0
r37 40 43 10.9824 $w=1.022e-06 $l=9.2e-07 $layer=LI1_cond $X=3.12 $Y=0.462
+ $X2=4.04 $Y2=0.462
r38 40 41 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r39 38 40 1.96967 $w=1.022e-06 $l=1.65e-07 $layer=LI1_cond $X=2.955 $Y=0.462
+ $X2=3.12 $Y2=0.462
r40 35 36 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r41 33 41 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r42 32 33 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r43 30 38 12.137 $w=1.022e-06 $l=5.07281e-07 $layer=LI1_cond $X=2.86 $Y=0
+ $X2=2.955 $Y2=0.462
r44 30 32 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=2.86 $Y=0 $X2=2.64
+ $Y2=0
r45 28 29 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r46 26 29 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r47 26 36 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r48 25 28 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r49 25 26 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r50 23 35 4.97422 $w=1.7e-07 $l=2.35e-07 $layer=LI1_cond $X=0.47 $Y=0 $X2=0.235
+ $Y2=0
r51 23 25 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=0.47 $Y=0 $X2=0.72
+ $Y2=0
r52 21 33 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r53 21 29 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.68
+ $Y2=0
r54 19 28 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=1.86 $Y=0 $X2=1.68
+ $Y2=0
r55 19 20 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.86 $Y=0 $X2=2.025
+ $Y2=0
r56 18 32 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=2.19 $Y=0 $X2=2.64
+ $Y2=0
r57 18 20 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.19 $Y=0 $X2=2.025
+ $Y2=0
r58 14 20 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.025 $Y=0.085
+ $X2=2.025 $Y2=0
r59 14 16 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=2.025 $Y=0.085
+ $X2=2.025 $Y2=0.55
r60 10 35 3.0057 $w=3.55e-07 $l=1.09864e-07 $layer=LI1_cond $X=0.292 $Y=0.085
+ $X2=0.235 $Y2=0
r61 10 12 13.9592 $w=3.53e-07 $l=4.3e-07 $layer=LI1_cond $X=0.292 $Y=0.085
+ $X2=0.292 $Y2=0.515
r62 3 43 60.6667 $w=1.7e-07 $l=1.29074e-06 $layer=licon1_NDIFF $count=3 $X=2.815
+ $Y=0.37 $X2=4.04 $Y2=0.505
r63 3 38 60.6667 $w=1.7e-07 $l=1.96214e-07 $layer=licon1_NDIFF $count=3 $X=2.815
+ $Y=0.37 $X2=2.955 $Y2=0.505
r64 2 16 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=1.885 $Y=0.37
+ $X2=2.025 $Y2=0.55
r65 1 12 91 $w=1.7e-07 $l=2.31409e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.37 $X2=0.305 $Y2=0.515
.ends

