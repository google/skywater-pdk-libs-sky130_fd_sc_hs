# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_hs__nand4bb_1
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_hs__nand4bb_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.320000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A_N
    ANTENNAGATEAREA  0.208500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 0.255000 0.480000 0.670000 ;
    END
  END A_N
  PIN B_N
    ANTENNAGATEAREA  0.208500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605000 1.470000 1.315000 1.800000 ;
    END
  END B_N
  PIN C
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.985000 0.810000 3.315000 1.550000 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.485000 1.350000 3.885000 1.780000 ;
    END
  END D
  PIN Y
    ANTENNADIFFAREA  1.248650 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.675000 2.310000 3.095000 2.480000 ;
        RECT 1.675000 2.480000 2.005000 2.980000 ;
        RECT 1.720000 0.350000 3.655000 0.620000 ;
        RECT 2.525000 1.820000 3.095000 1.950000 ;
        RECT 2.525000 1.950000 4.225000 2.120000 ;
        RECT 2.525000 2.120000 3.095000 2.310000 ;
        RECT 2.765000 2.480000 3.095000 2.980000 ;
        RECT 3.485000 0.620000 3.655000 1.010000 ;
        RECT 3.485000 1.010000 4.225000 1.180000 ;
        RECT 3.765000 2.120000 4.225000 2.980000 ;
        RECT 4.055000 1.180000 4.225000 1.950000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 4.320000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 4.320000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.320000 0.085000 ;
      RECT 0.000000  3.245000 4.320000 3.415000 ;
      RECT 0.115000  0.840000 0.470000 1.130000 ;
      RECT 0.115000  1.130000 2.015000 1.300000 ;
      RECT 0.115000  1.300000 0.285000 1.970000 ;
      RECT 0.115000  1.970000 0.445000 2.850000 ;
      RECT 0.615000  1.970000 0.945000 3.245000 ;
      RECT 0.650000  0.085000 0.980000 0.960000 ;
      RECT 1.115000  1.970000 2.355000 2.140000 ;
      RECT 1.115000  2.140000 1.445000 2.850000 ;
      RECT 1.150000  0.630000 1.490000 0.790000 ;
      RECT 1.150000  0.790000 2.355000 0.960000 ;
      RECT 1.685000  1.300000 2.015000 1.550000 ;
      RECT 2.175000  2.650000 2.595000 3.245000 ;
      RECT 2.185000  0.960000 2.355000 1.220000 ;
      RECT 2.185000  1.220000 2.745000 1.550000 ;
      RECT 2.185000  1.550000 2.355000 1.970000 ;
      RECT 3.265000  2.290000 3.595000 3.245000 ;
      RECT 3.825000  0.085000 4.155000 0.840000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
  END
END sky130_fd_sc_hs__nand4bb_1
END LIBRARY
