* File: sky130_fd_sc_hs__dfxtp_1.pex.spice
* Created: Thu Aug 27 20:39:57 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HS__DFXTP_1%CLK 3 5 7 8 12
c33 5 0 1.5421e-19 $X=0.505 $Y=1.765
r34 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.34
+ $Y=1.465 $X2=0.34 $Y2=1.465
r35 8 12 6.06549 $w=3.78e-07 $l=2e-07 $layer=LI1_cond $X=0.315 $Y=1.665
+ $X2=0.315 $Y2=1.465
r36 5 11 57.3754 $w=3.5e-07 $l=3.54965e-07 $layer=POLY_cond $X=0.505 $Y=1.765
+ $X2=0.385 $Y2=1.465
r37 5 7 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.505 $Y=1.765
+ $X2=0.505 $Y2=2.4
r38 1 11 38.7839 $w=3.5e-07 $l=2.13014e-07 $layer=POLY_cond $X=0.495 $Y=1.3
+ $X2=0.385 $Y2=1.465
r39 1 3 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=0.495 $Y=1.3 $X2=0.495
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HS__DFXTP_1%A_27_74# 1 2 7 9 10 12 15 18 19 21 22 24 25
+ 30 31 35 37 39 41 42 43 46 49 50 52 53 54 56 57 58 59 62 65 67 68 71 73 76 77
+ 82 84 85 86
c278 84 0 6.36416e-20 $X=5.73 $Y=0.345
c279 76 0 1.82292e-19 $X=0.905 $Y=1.045
c280 19 0 1.86961e-19 $X=3.265 $Y=2.44
r281 85 94 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.73 $Y=0.345
+ $X2=5.73 $Y2=0.51
r282 84 86 8.74048 $w=2.53e-07 $l=1.65e-07 $layer=LI1_cond $X=5.73 $Y=0.382
+ $X2=5.565 $Y2=0.382
r283 84 85 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.73
+ $Y=0.345 $X2=5.73 $Y2=0.345
r284 79 81 9.2801 $w=4.58e-07 $l=1.65e-07 $layer=LI1_cond $X=0.905 $Y=1.385
+ $X2=0.905 $Y2=1.55
r285 79 80 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.97
+ $Y=1.385 $X2=0.97 $Y2=1.385
r286 76 79 8.84058 $w=4.58e-07 $l=3.4e-07 $layer=LI1_cond $X=0.905 $Y=1.045
+ $X2=0.905 $Y2=1.385
r287 76 77 7.19996 $w=4.58e-07 $l=8.5e-08 $layer=LI1_cond $X=0.905 $Y=1.045
+ $X2=0.905 $Y2=0.96
r288 73 86 59.0428 $w=1.68e-07 $l=9.05e-07 $layer=LI1_cond $X=4.66 $Y=0.34
+ $X2=5.565 $Y2=0.34
r289 70 73 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.575 $Y=0.425
+ $X2=4.66 $Y2=0.34
r290 70 71 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=4.575 $Y=0.425
+ $X2=4.575 $Y2=0.69
r291 69 82 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.76 $Y=0.775
+ $X2=3.675 $Y2=0.775
r292 68 71 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.49 $Y=0.775
+ $X2=4.575 $Y2=0.69
r293 68 69 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=4.49 $Y=0.775
+ $X2=3.76 $Y2=0.775
r294 66 82 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.675 $Y=0.86
+ $X2=3.675 $Y2=0.775
r295 66 67 58.0642 $w=1.68e-07 $l=8.9e-07 $layer=LI1_cond $X=3.675 $Y=0.86
+ $X2=3.675 $Y2=1.75
r296 65 82 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.675 $Y=0.69
+ $X2=3.675 $Y2=0.775
r297 64 65 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=3.675 $Y=0.445
+ $X2=3.675 $Y2=0.69
r298 62 91 40.9837 $w=3.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.215 $Y=1.915
+ $X2=3.215 $Y2=2.08
r299 62 90 46.7569 $w=3.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.215 $Y=1.915
+ $X2=3.215 $Y2=1.75
r300 61 62 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.235
+ $Y=1.915 $X2=3.235 $Y2=1.915
r301 59 67 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.59 $Y=1.915
+ $X2=3.675 $Y2=1.75
r302 59 61 12.3975 $w=3.28e-07 $l=3.55e-07 $layer=LI1_cond $X=3.59 $Y=1.915
+ $X2=3.235 $Y2=1.915
r303 57 64 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.59 $Y=0.36
+ $X2=3.675 $Y2=0.445
r304 57 58 61 $w=1.68e-07 $l=9.35e-07 $layer=LI1_cond $X=3.59 $Y=0.36 $X2=2.655
+ $Y2=0.36
r305 55 58 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.57 $Y=0.445
+ $X2=2.655 $Y2=0.36
r306 55 56 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=2.57 $Y=0.445
+ $X2=2.57 $Y2=0.73
r307 53 56 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.485 $Y=0.815
+ $X2=2.57 $Y2=0.73
r308 53 54 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.485 $Y=0.815
+ $X2=1.815 $Y2=0.815
r309 52 54 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.73 $Y=0.73
+ $X2=1.815 $Y2=0.815
r310 51 52 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.73 $Y=0.425
+ $X2=1.73 $Y2=0.73
r311 49 51 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.645 $Y=0.34
+ $X2=1.73 $Y2=0.425
r312 49 50 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=1.645 $Y=0.34
+ $X2=1.135 $Y2=0.34
r313 47 50 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.05 $Y=0.425
+ $X2=1.135 $Y2=0.34
r314 47 77 34.9037 $w=1.68e-07 $l=5.35e-07 $layer=LI1_cond $X=1.05 $Y=0.425
+ $X2=1.05 $Y2=0.96
r315 46 81 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=0.76 $Y=1.95 $X2=0.76
+ $Y2=1.55
r316 44 75 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.445 $Y=2.035
+ $X2=0.28 $Y2=2.035
r317 43 46 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.675 $Y=2.035
+ $X2=0.76 $Y2=1.95
r318 43 44 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=0.675 $Y=2.035
+ $X2=0.445 $Y2=2.035
r319 41 76 6.6364 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=0.675 $Y=1.045
+ $X2=0.905 $Y2=1.045
r320 41 42 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=0.675 $Y=1.045
+ $X2=0.365 $Y2=1.045
r321 37 75 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.28 $Y=2.12 $X2=0.28
+ $Y2=2.035
r322 37 39 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=0.28 $Y=2.12
+ $X2=0.28 $Y2=2.815
r323 33 42 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.24 $Y=0.96
+ $X2=0.365 $Y2=1.045
r324 33 35 20.5135 $w=2.48e-07 $l=4.45e-07 $layer=LI1_cond $X=0.24 $Y=0.96
+ $X2=0.24 $Y2=0.515
r325 30 94 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=5.765 $Y=0.83
+ $X2=5.765 $Y2=0.51
r326 28 30 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=5.765 $Y=1.69
+ $X2=5.765 $Y2=0.83
r327 26 31 7.1379 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=5.07 $Y=1.765 $X2=4.98
+ $Y2=1.765
r328 25 28 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.69 $Y=1.765
+ $X2=5.765 $Y2=1.69
r329 25 26 317.915 $w=1.5e-07 $l=6.2e-07 $layer=POLY_cond $X=5.69 $Y=1.765
+ $X2=5.07 $Y2=1.765
r330 22 31 110.989 $w=1.8e-07 $l=2.8e-07 $layer=POLY_cond $X=4.98 $Y=2.045
+ $X2=4.98 $Y2=1.765
r331 22 24 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=4.98 $Y=2.045
+ $X2=4.98 $Y2=2.54
r332 19 21 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=3.265 $Y=2.44
+ $X2=3.265 $Y2=2.725
r333 18 19 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=3.265 $Y=2.35
+ $X2=3.265 $Y2=2.44
r334 18 91 104.952 $w=1.8e-07 $l=2.7e-07 $layer=POLY_cond $X=3.265 $Y=2.35
+ $X2=3.265 $Y2=2.08
r335 15 90 469.181 $w=1.5e-07 $l=9.15e-07 $layer=POLY_cond $X=3.105 $Y=0.835
+ $X2=3.105 $Y2=1.75
r336 10 80 38.539 $w=3.04e-07 $l=2.1609e-07 $layer=POLY_cond $X=1.115 $Y=1.22
+ $X2=0.997 $Y2=1.385
r337 10 12 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.115 $Y=1.22
+ $X2=1.115 $Y2=0.74
r338 7 80 72.6278 $w=3.04e-07 $l=4.0045e-07 $layer=POLY_cond $X=0.955 $Y=1.765
+ $X2=0.997 $Y2=1.385
r339 7 9 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.955 $Y=1.765
+ $X2=0.955 $Y2=2.4
r340 2 75 400 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.115
r341 2 39 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.815
r342 1 35 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__DFXTP_1%D 1 3 4 6 7 14 15 22
r47 22 23 1.12427 $w=3.78e-07 $l=1e-08 $layer=LI1_cond $X=2.06 $Y=2.035 $X2=2.06
+ $Y2=2.025
r48 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.135
+ $Y=1.29 $X2=2.135 $Y2=1.29
r49 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.035
+ $Y=2.19 $X2=2.035 $Y2=2.19
r50 7 12 3.57864 $w=3.78e-07 $l=1.18e-07 $layer=LI1_cond $X=2.06 $Y=2.072
+ $X2=2.06 $Y2=2.19
r51 7 22 1.12212 $w=3.78e-07 $l=3.7e-08 $layer=LI1_cond $X=2.06 $Y=2.072
+ $X2=2.06 $Y2=2.035
r52 7 23 1.56403 $w=2.78e-07 $l=3.8e-08 $layer=LI1_cond $X=2.11 $Y=1.987
+ $X2=2.11 $Y2=2.025
r53 7 15 28.6876 $w=2.78e-07 $l=6.97e-07 $layer=LI1_cond $X=2.11 $Y=1.987
+ $X2=2.11 $Y2=1.29
r54 4 14 57.9147 $w=2.58e-07 $l=3.83732e-07 $layer=POLY_cond $X=2.445 $Y=1.125
+ $X2=2.135 $Y2=1.29
r55 4 6 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.445 $Y=1.125
+ $X2=2.445 $Y2=0.805
r56 1 11 50.1894 $w=3.66e-07 $l=3.03315e-07 $layer=POLY_cond $X=2.195 $Y=2.44
+ $X2=2.077 $Y2=2.19
r57 1 3 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=2.195 $Y=2.44 $X2=2.195
+ $Y2=2.725
.ends

.subckt PM_SKY130_FD_SC_HS__DFXTP_1%A_206_368# 1 2 9 10 11 14 15 17 20 22 24 25
+ 27 29 32 36 38 40 43 44 45 46 50 54 55 61 62 64 68 72 76 77 82
c235 77 0 1.78324e-19 $X=5.315 $Y=1.315
c236 62 0 1.82292e-19 $X=1.595 $Y=1.515
c237 54 0 1.5421e-19 $X=1.18 $Y=1.985
c238 40 0 1.86961e-19 $X=4.78 $Y=2.71
c239 25 0 1.31987e-20 $X=5.515 $Y=2.465
c240 20 0 2.31753e-20 $X=3.58 $Y=0.715
r241 77 85 32.3493 $w=3.3e-07 $l=1.85e-07 $layer=POLY_cond $X=5.315 $Y=1.315
+ $X2=5.13 $Y2=1.315
r242 76 79 5.20458 $w=3.08e-07 $l=1.4e-07 $layer=LI1_cond $X=5.325 $Y=1.315
+ $X2=5.325 $Y2=1.455
r243 76 77 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.315
+ $Y=1.315 $X2=5.315 $Y2=1.315
r244 72 73 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=4.865 $Y=2.71
+ $X2=4.865 $Y2=2.99
r245 68 70 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=3.375 $Y=2.71
+ $X2=3.375 $Y2=2.88
r246 64 66 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=2.165 $Y=2.71
+ $X2=2.165 $Y2=2.88
r247 62 83 39.3438 $w=3.3e-07 $l=2.25e-07 $layer=POLY_cond $X=1.595 $Y=1.515
+ $X2=1.595 $Y2=1.74
r248 62 82 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.595 $Y=1.515
+ $X2=1.595 $Y2=1.35
r249 61 62 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.595
+ $Y=1.515 $X2=1.595 $Y2=1.515
r250 58 61 7.15912 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=1.39 $Y=1.515
+ $X2=1.595 $Y2=1.515
r251 54 55 9.2801 $w=4.58e-07 $l=1.65e-07 $layer=LI1_cond $X=1.245 $Y=1.985
+ $X2=1.245 $Y2=1.82
r252 50 51 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.675
+ $Y=2.215 $X2=5.675 $Y2=2.215
r253 48 50 24.0965 $w=3.28e-07 $l=6.9e-07 $layer=LI1_cond $X=5.675 $Y=2.905
+ $X2=5.675 $Y2=2.215
r254 47 73 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.95 $Y=2.99
+ $X2=4.865 $Y2=2.99
r255 46 48 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=5.51 $Y=2.99
+ $X2=5.675 $Y2=2.905
r256 46 47 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=5.51 $Y=2.99
+ $X2=4.95 $Y2=2.99
r257 44 79 4.25403 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=5.17 $Y=1.455
+ $X2=5.325 $Y2=1.455
r258 44 45 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=5.17 $Y=1.455
+ $X2=4.95 $Y2=1.455
r259 43 72 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=4.865 $Y=2.625
+ $X2=4.865 $Y2=2.71
r260 42 45 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.865 $Y=1.54
+ $X2=4.95 $Y2=1.455
r261 42 43 70.7861 $w=1.68e-07 $l=1.085e-06 $layer=LI1_cond $X=4.865 $Y=1.54
+ $X2=4.865 $Y2=2.625
r262 41 68 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.46 $Y=2.71
+ $X2=3.375 $Y2=2.71
r263 40 72 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.78 $Y=2.71
+ $X2=4.865 $Y2=2.71
r264 40 41 86.1176 $w=1.68e-07 $l=1.32e-06 $layer=LI1_cond $X=4.78 $Y=2.71
+ $X2=3.46 $Y2=2.71
r265 39 66 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.25 $Y=2.88
+ $X2=2.165 $Y2=2.88
r266 38 70 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.29 $Y=2.88
+ $X2=3.375 $Y2=2.88
r267 38 39 67.8503 $w=1.68e-07 $l=1.04e-06 $layer=LI1_cond $X=3.29 $Y=2.88
+ $X2=2.25 $Y2=2.88
r268 37 57 5.73712 $w=1.7e-07 $l=2.7214e-07 $layer=LI1_cond $X=1.475 $Y=2.71
+ $X2=1.245 $Y2=2.802
r269 36 64 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.08 $Y=2.71
+ $X2=2.165 $Y2=2.71
r270 36 37 39.4706 $w=1.68e-07 $l=6.05e-07 $layer=LI1_cond $X=2.08 $Y=2.71
+ $X2=1.475 $Y2=2.71
r271 34 58 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.39 $Y=1.68
+ $X2=1.39 $Y2=1.515
r272 34 55 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=1.39 $Y=1.68
+ $X2=1.39 $Y2=1.82
r273 30 58 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.39 $Y=1.35
+ $X2=1.39 $Y2=1.515
r274 30 32 31.9679 $w=1.68e-07 $l=4.9e-07 $layer=LI1_cond $X=1.39 $Y=1.35
+ $X2=1.39 $Y2=0.86
r275 29 57 3.15363 $w=4.6e-07 $l=1.77e-07 $layer=LI1_cond $X=1.245 $Y=2.625
+ $X2=1.245 $Y2=2.802
r276 28 54 1.69011 $w=4.58e-07 $l=6.5e-08 $layer=LI1_cond $X=1.245 $Y=2.05
+ $X2=1.245 $Y2=1.985
r277 28 29 14.951 $w=4.58e-07 $l=5.75e-07 $layer=LI1_cond $X=1.245 $Y=2.05
+ $X2=1.245 $Y2=2.625
r278 25 51 50.1894 $w=3.66e-07 $l=3.02903e-07 $layer=POLY_cond $X=5.515 $Y=2.465
+ $X2=5.632 $Y2=2.215
r279 25 27 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=5.515 $Y=2.465
+ $X2=5.515 $Y2=2.75
r280 22 85 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.13 $Y=1.15
+ $X2=5.13 $Y2=1.315
r281 22 24 123.713 $w=1.5e-07 $l=3.85e-07 $layer=POLY_cond $X=5.13 $Y=1.15
+ $X2=5.13 $Y2=0.765
r282 18 20 235.872 $w=1.5e-07 $l=4.6e-07 $layer=POLY_cond $X=3.58 $Y=0.255
+ $X2=3.58 $Y2=0.715
r283 15 17 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=2.73 $Y=2.24
+ $X2=2.73 $Y2=2.525
r284 14 15 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=2.73 $Y=2.15 $X2=2.73
+ $Y2=2.24
r285 13 14 130.218 $w=1.8e-07 $l=3.35e-07 $layer=POLY_cond $X=2.73 $Y=1.815
+ $X2=2.73 $Y2=2.15
r286 12 83 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.76 $Y=1.74
+ $X2=1.595 $Y2=1.74
r287 11 13 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=2.64 $Y=1.74
+ $X2=2.73 $Y2=1.815
r288 11 12 451.234 $w=1.5e-07 $l=8.8e-07 $layer=POLY_cond $X=2.64 $Y=1.74
+ $X2=1.76 $Y2=1.74
r289 9 18 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.505 $Y=0.18
+ $X2=3.58 $Y2=0.255
r290 9 10 894.777 $w=1.5e-07 $l=1.745e-06 $layer=POLY_cond $X=3.505 $Y=0.18
+ $X2=1.76 $Y2=0.18
r291 7 10 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.685 $Y=0.255
+ $X2=1.76 $Y2=0.18
r292 7 82 561.479 $w=1.5e-07 $l=1.095e-06 $layer=POLY_cond $X=1.685 $Y=0.255
+ $X2=1.685 $Y2=1.35
r293 2 57 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=1.03
+ $Y=1.84 $X2=1.18 $Y2=2.815
r294 2 54 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=1.03
+ $Y=1.84 $X2=1.18 $Y2=1.985
r295 1 32 182 $w=1.7e-07 $l=5.81464e-07 $layer=licon1_NDIFF $count=1 $X=1.19
+ $Y=0.37 $X2=1.39 $Y2=0.86
.ends

.subckt PM_SKY130_FD_SC_HS__DFXTP_1%A_713_458# 1 2 9 14 16 17 18 22 26 28 35 36
+ 38 40
c96 28 0 1.54375e-19 $X=4.095 $Y=1.115
r97 35 36 8.58424 $w=2.73e-07 $l=1.65e-07 $layer=LI1_cond $X=4.472 $Y=2.29
+ $X2=4.472 $Y2=2.125
r98 32 40 28.8456 $w=2.59e-07 $l=1.55e-07 $layer=POLY_cond $X=4.095 $Y=1.25
+ $X2=3.94 $Y2=1.25
r99 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.095
+ $Y=1.25 $X2=4.095 $Y2=1.25
r100 28 31 4.71454 $w=3.28e-07 $l=1.35e-07 $layer=LI1_cond $X=4.095 $Y=1.115
+ $X2=4.095 $Y2=1.25
r101 24 26 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=4.915 $Y=1.03
+ $X2=4.915 $Y2=0.825
r102 23 38 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.61 $Y=1.115
+ $X2=4.525 $Y2=1.115
r103 22 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.83 $Y=1.115
+ $X2=4.915 $Y2=1.03
r104 22 23 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=4.83 $Y=1.115
+ $X2=4.61 $Y2=1.115
r105 20 38 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.525 $Y=1.2
+ $X2=4.525 $Y2=1.115
r106 20 36 60.3476 $w=1.68e-07 $l=9.25e-07 $layer=LI1_cond $X=4.525 $Y=1.2
+ $X2=4.525 $Y2=2.125
r107 19 28 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.26 $Y=1.115
+ $X2=4.095 $Y2=1.115
r108 18 38 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.44 $Y=1.115
+ $X2=4.525 $Y2=1.115
r109 18 19 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=4.44 $Y=1.115
+ $X2=4.26 $Y2=1.115
r110 16 17 51.0119 $w=1.95e-07 $l=1.5e-07 $layer=POLY_cond $X=3.662 $Y=2.29
+ $X2=3.662 $Y2=2.44
r111 12 40 15.5386 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.94 $Y=1.085
+ $X2=3.94 $Y2=1.25
r112 12 14 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=3.94 $Y=1.085
+ $X2=3.94 $Y2=0.715
r113 10 40 47.4556 $w=2.59e-07 $l=3.27261e-07 $layer=POLY_cond $X=3.685 $Y=1.415
+ $X2=3.94 $Y2=1.25
r114 10 16 448.67 $w=1.5e-07 $l=8.75e-07 $layer=POLY_cond $X=3.685 $Y=1.415
+ $X2=3.685 $Y2=2.29
r115 9 17 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=3.655 $Y=2.725
+ $X2=3.655 $Y2=2.44
r116 2 35 600 $w=1.7e-07 $l=2.36854e-07 $layer=licon1_PDIFF $count=1 $X=4.35
+ $Y=2.12 $X2=4.51 $Y2=2.29
r117 1 26 182 $w=1.7e-07 $l=5.4909e-07 $layer=licon1_NDIFF $count=1 $X=4.695
+ $Y=0.375 $X2=4.915 $Y2=0.825
.ends

.subckt PM_SKY130_FD_SC_HS__DFXTP_1%A_561_463# 1 2 7 9 11 14 17 19 20 21 22 26
+ 29 34 36 41
c120 17 0 1.31199e-19 $X=4.597 $Y=1.45
r121 37 41 24.2734 $w=2.78e-07 $l=1.4e-07 $layer=POLY_cond $X=4.135 $Y=1.835
+ $X2=4.275 $Y2=1.835
r122 36 39 8.48463 $w=2.98e-07 $l=1.65e-07 $layer=LI1_cond $X=4.12 $Y=1.79
+ $X2=4.12 $Y2=1.955
r123 36 37 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.135
+ $Y=1.79 $X2=4.135 $Y2=1.79
r124 33 34 8.47192 $w=3.38e-07 $l=1.65e-07 $layer=LI1_cond $X=2.955 $Y=2.455
+ $X2=3.12 $Y2=2.455
r125 30 33 3.72849 $w=3.38e-07 $l=1.1e-07 $layer=LI1_cond $X=2.845 $Y=2.455
+ $X2=2.955 $Y2=2.455
r126 29 39 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=4.055 $Y=2.285
+ $X2=4.055 $Y2=1.955
r127 24 26 27.3977 $w=2.63e-07 $l=6.3e-07 $layer=LI1_cond $X=3.287 $Y=1.41
+ $X2=3.287 $Y2=0.78
r128 22 29 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.97 $Y=2.37
+ $X2=4.055 $Y2=2.285
r129 22 34 55.4545 $w=1.68e-07 $l=8.5e-07 $layer=LI1_cond $X=3.97 $Y=2.37
+ $X2=3.12 $Y2=2.37
r130 20 24 7.24806 $w=1.7e-07 $l=1.69245e-07 $layer=LI1_cond $X=3.155 $Y=1.495
+ $X2=3.287 $Y2=1.41
r131 20 21 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=3.155 $Y=1.495
+ $X2=2.93 $Y2=1.495
r132 19 30 4.80115 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=2.845 $Y=2.285
+ $X2=2.845 $Y2=2.455
r133 18 21 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.845 $Y=1.58
+ $X2=2.93 $Y2=1.495
r134 18 19 45.9947 $w=1.68e-07 $l=7.05e-07 $layer=LI1_cond $X=2.845 $Y=1.58
+ $X2=2.845 $Y2=2.285
r135 16 17 51.0119 $w=1.95e-07 $l=1.5e-07 $layer=POLY_cond $X=4.597 $Y=1.3
+ $X2=4.597 $Y2=1.45
r136 14 16 333.298 $w=1.5e-07 $l=6.5e-07 $layer=POLY_cond $X=4.62 $Y=0.65
+ $X2=4.62 $Y2=1.3
r137 11 41 52.0144 $w=2.78e-07 $l=3.91152e-07 $layer=POLY_cond $X=4.575 $Y=1.625
+ $X2=4.275 $Y2=1.835
r138 11 17 89.734 $w=1.5e-07 $l=1.75e-07 $layer=POLY_cond $X=4.575 $Y=1.625
+ $X2=4.575 $Y2=1.45
r139 7 41 17.1848 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=4.275 $Y=2.045
+ $X2=4.275 $Y2=1.835
r140 7 9 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=4.275 $Y=2.045
+ $X2=4.275 $Y2=2.54
r141 2 33 600 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=2.805
+ $Y=2.315 $X2=2.955 $Y2=2.46
r142 1 26 182 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_NDIFF $count=1 $X=3.18
+ $Y=0.625 $X2=3.325 $Y2=0.78
.ends

.subckt PM_SKY130_FD_SC_HS__DFXTP_1%A_1210_314# 1 2 7 9 12 14 16 19 23 26 30 34
+ 36 38 39 43 44 45 47 49
c116 44 0 3.28719e-19 $X=6.215 $Y=1.735
c117 14 0 1.70354e-19 $X=7.655 $Y=1.765
c118 12 0 6.36416e-20 $X=6.18 $Y=0.83
r119 47 50 8.3232 $w=3.58e-07 $l=2.6e-07 $layer=LI1_cond $X=7.555 $Y=1.515
+ $X2=7.555 $Y2=1.775
r120 47 49 8.51103 $w=3.58e-07 $l=1.65e-07 $layer=LI1_cond $X=7.555 $Y=1.515
+ $X2=7.555 $Y2=1.35
r121 47 48 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.62
+ $Y=1.515 $X2=7.62 $Y2=1.515
r122 43 44 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.215
+ $Y=1.735 $X2=6.215 $Y2=1.735
r123 40 49 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=7.46 $Y=1.02
+ $X2=7.46 $Y2=1.35
r124 38 40 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.375 $Y=0.935
+ $X2=7.46 $Y2=1.02
r125 38 39 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=7.375 $Y=0.935
+ $X2=7.04 $Y2=0.935
r126 37 45 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.01 $Y=1.775
+ $X2=6.885 $Y2=1.775
r127 36 50 5.14255 $w=1.7e-07 $l=1.8e-07 $layer=LI1_cond $X=7.375 $Y=1.775
+ $X2=7.555 $Y2=1.775
r128 36 37 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=7.375 $Y=1.775
+ $X2=7.01 $Y2=1.775
r129 32 39 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=6.915 $Y=0.85
+ $X2=7.04 $Y2=0.935
r130 32 34 9.45003 $w=2.48e-07 $l=2.05e-07 $layer=LI1_cond $X=6.915 $Y=0.85
+ $X2=6.915 $Y2=0.645
r131 28 45 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.885 $Y=1.86
+ $X2=6.885 $Y2=1.775
r132 28 30 5.76222 $w=2.48e-07 $l=1.25e-07 $layer=LI1_cond $X=6.885 $Y=1.86
+ $X2=6.885 $Y2=1.985
r133 27 43 4.72267 $w=1.7e-07 $l=1.92678e-07 $layer=LI1_cond $X=6.38 $Y=1.775
+ $X2=6.215 $Y2=1.715
r134 26 45 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.76 $Y=1.775
+ $X2=6.885 $Y2=1.775
r135 26 27 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=6.76 $Y=1.775
+ $X2=6.38 $Y2=1.775
r136 23 44 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=6.215 $Y=2.075
+ $X2=6.215 $Y2=1.735
r137 22 44 39.6269 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.215 $Y=1.57
+ $X2=6.215 $Y2=1.735
r138 17 48 38.5562 $w=2.99e-07 $l=1.86145e-07 $layer=POLY_cond $X=7.665 $Y=1.35
+ $X2=7.62 $Y2=1.515
r139 17 19 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=7.665 $Y=1.35
+ $X2=7.665 $Y2=0.74
r140 14 48 52.2586 $w=2.99e-07 $l=2.66927e-07 $layer=POLY_cond $X=7.655 $Y=1.765
+ $X2=7.62 $Y2=1.515
r141 14 16 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=7.655 $Y=1.765
+ $X2=7.655 $Y2=2.4
r142 12 22 379.447 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=6.18 $Y=0.83
+ $X2=6.18 $Y2=1.57
r143 7 23 77.358 $w=2.43e-07 $l=4.25852e-07 $layer=POLY_cond $X=6.14 $Y=2.465
+ $X2=6.215 $Y2=2.075
r144 7 9 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=6.14 $Y=2.465 $X2=6.14
+ $Y2=2.75
r145 2 30 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=6.78
+ $Y=1.84 $X2=6.925 $Y2=1.985
r146 1 34 182 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_NDIFF $count=1 $X=6.81
+ $Y=0.37 $X2=6.955 $Y2=0.645
.ends

.subckt PM_SKY130_FD_SC_HS__DFXTP_1%A_1011_424# 1 2 7 8 9 11 14 18 20 24 25 27
+ 29 32 34 36
c102 36 0 1.31987e-20 $X=6.875 $Y=1.355
c103 34 0 1.70354e-19 $X=7.04 $Y=1.355
c104 29 0 1.71535e-19 $X=5.735 $Y=1.71
c105 25 0 1.78324e-19 $X=5.29 $Y=1.795
c106 24 0 1.57185e-19 $X=5.65 $Y=1.795
c107 14 0 2.87771e-20 $X=7.17 $Y=0.69
r108 34 36 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=7.04 $Y=1.355
+ $X2=6.875 $Y2=1.355
r109 34 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.04
+ $Y=1.355 $X2=7.04 $Y2=1.355
r110 31 32 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.82 $Y=1.315
+ $X2=5.735 $Y2=1.315
r111 31 36 68.8289 $w=1.68e-07 $l=1.055e-06 $layer=LI1_cond $X=5.82 $Y=1.315
+ $X2=6.875 $Y2=1.315
r112 28 32 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.735 $Y=1.4
+ $X2=5.735 $Y2=1.315
r113 28 29 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=5.735 $Y=1.4
+ $X2=5.735 $Y2=1.71
r114 27 32 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.735 $Y=1.23
+ $X2=5.735 $Y2=1.315
r115 26 27 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=5.735 $Y=0.98
+ $X2=5.735 $Y2=1.23
r116 24 29 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.65 $Y=1.795
+ $X2=5.735 $Y2=1.71
r117 24 25 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=5.65 $Y=1.795
+ $X2=5.29 $Y2=1.795
r118 20 26 7.14316 $w=2.5e-07 $l=1.62019e-07 $layer=LI1_cond $X=5.65 $Y=0.855
+ $X2=5.735 $Y2=0.98
r119 20 22 9.45003 $w=2.48e-07 $l=2.05e-07 $layer=LI1_cond $X=5.65 $Y=0.855
+ $X2=5.445 $Y2=0.855
r120 16 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.205 $Y=1.88
+ $X2=5.29 $Y2=1.795
r121 16 18 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=5.205 $Y=1.88
+ $X2=5.205 $Y2=2.48
r122 12 35 39.0103 $w=3.67e-07 $l=2.13014e-07 $layer=POLY_cond $X=7.17 $Y=1.19
+ $X2=7.06 $Y2=1.355
r123 12 14 256.383 $w=1.5e-07 $l=5e-07 $layer=POLY_cond $X=7.17 $Y=1.19 $X2=7.17
+ $Y2=0.69
r124 9 11 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=7.15 $Y=1.765
+ $X2=7.15 $Y2=2.26
r125 8 9 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=7.15 $Y=1.675 $X2=7.15
+ $Y2=1.765
r126 7 35 34.2012 $w=3.67e-07 $l=2.05122e-07 $layer=POLY_cond $X=7.15 $Y=1.52
+ $X2=7.06 $Y2=1.355
r127 7 8 60.25 $w=1.8e-07 $l=1.55e-07 $layer=POLY_cond $X=7.15 $Y=1.52 $X2=7.15
+ $Y2=1.675
r128 2 18 600 $w=1.7e-07 $l=4.28486e-07 $layer=licon1_PDIFF $count=1 $X=5.055
+ $Y=2.12 $X2=5.205 $Y2=2.48
r129 1 22 182 $w=1.7e-07 $l=4.28515e-07 $layer=licon1_NDIFF $count=1 $X=5.205
+ $Y=0.49 $X2=5.445 $Y2=0.815
.ends

.subckt PM_SKY130_FD_SC_HS__DFXTP_1%VPWR 1 2 3 4 5 20 24 28 31 32 33 35 40 52 58
+ 59 62 65 72 79
r99 79 80 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r100 72 75 9.7783 $w=3.28e-07 $l=2.8e-07 $layer=LI1_cond $X=3.965 $Y=3.05
+ $X2=3.965 $Y2=3.33
r101 62 63 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r102 59 80 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=3.33
+ $X2=7.44 $Y2=3.33
r103 58 59 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r104 56 79 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.54 $Y=3.33
+ $X2=7.375 $Y2=3.33
r105 56 58 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=7.54 $Y=3.33
+ $X2=7.92 $Y2=3.33
r106 55 80 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=7.44 $Y2=3.33
r107 54 55 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r108 52 79 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.21 $Y=3.33
+ $X2=7.375 $Y2=3.33
r109 52 54 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=7.21 $Y=3.33
+ $X2=6.96 $Y2=3.33
r110 51 55 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6 $Y=3.33 $X2=6.96
+ $Y2=3.33
r111 50 51 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r112 48 75 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.13 $Y=3.33
+ $X2=3.965 $Y2=3.33
r113 48 50 122 $w=1.68e-07 $l=1.87e-06 $layer=LI1_cond $X=4.13 $Y=3.33 $X2=6
+ $Y2=3.33
r114 46 47 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r115 44 47 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=3.6 $Y2=3.33
r116 44 69 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.68 $Y2=3.33
r117 43 46 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=2.16 $Y=3.33
+ $X2=3.6 $Y2=3.33
r118 43 44 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r119 41 43 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=1.91 $Y=3.33
+ $X2=2.16 $Y2=3.33
r120 40 75 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.8 $Y=3.33
+ $X2=3.965 $Y2=3.33
r121 40 46 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=3.8 $Y=3.33 $X2=3.6
+ $Y2=3.33
r122 39 69 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=1.68 $Y2=3.33
r123 39 63 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r124 38 39 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r125 36 62 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.815 $Y=3.33
+ $X2=0.73 $Y2=3.33
r126 36 38 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=0.815 $Y=3.33
+ $X2=1.2 $Y2=3.33
r127 35 41 4.71304 $w=1.7e-07 $l=1.68e-07 $layer=LI1_cond $X=1.742 $Y=3.33
+ $X2=1.91 $Y2=3.33
r128 35 69 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r129 35 65 9.63236 $w=3.33e-07 $l=2.8e-07 $layer=LI1_cond $X=1.742 $Y=3.33
+ $X2=1.742 $Y2=3.05
r130 35 38 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=1.575 $Y=3.33
+ $X2=1.2 $Y2=3.33
r131 33 51 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=6 $Y2=3.33
r132 33 47 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=3.6 $Y2=3.33
r133 33 75 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r134 31 50 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=6.2 $Y=3.33 $X2=6
+ $Y2=3.33
r135 31 32 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.2 $Y=3.33
+ $X2=6.365 $Y2=3.33
r136 30 54 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=6.53 $Y=3.33
+ $X2=6.96 $Y2=3.33
r137 30 32 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.53 $Y=3.33
+ $X2=6.365 $Y2=3.33
r138 26 79 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.375 $Y=3.245
+ $X2=7.375 $Y2=3.33
r139 26 28 38.764 $w=3.28e-07 $l=1.11e-06 $layer=LI1_cond $X=7.375 $Y=3.245
+ $X2=7.375 $Y2=2.135
r140 22 32 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.365 $Y=3.245
+ $X2=6.365 $Y2=3.33
r141 22 24 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=6.365 $Y=3.245
+ $X2=6.365 $Y2=2.75
r142 18 62 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.73 $Y=3.245
+ $X2=0.73 $Y2=3.33
r143 18 20 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=0.73 $Y=3.245
+ $X2=0.73 $Y2=2.455
r144 5 28 300 $w=1.7e-07 $l=3.62319e-07 $layer=licon1_PDIFF $count=2 $X=7.225
+ $Y=1.84 $X2=7.375 $Y2=2.135
r145 4 24 600 $w=1.7e-07 $l=2.74955e-07 $layer=licon1_PDIFF $count=1 $X=6.215
+ $Y=2.54 $X2=6.365 $Y2=2.75
r146 3 72 600 $w=1.7e-07 $l=6.41833e-07 $layer=licon1_PDIFF $count=1 $X=3.73
+ $Y=2.515 $X2=3.965 $Y2=3.05
r147 2 65 600 $w=1.7e-07 $l=6.03158e-07 $layer=licon1_PDIFF $count=1 $X=1.595
+ $Y=2.515 $X2=1.74 $Y2=3.05
r148 1 20 300 $w=1.7e-07 $l=6.85912e-07 $layer=licon1_PDIFF $count=2 $X=0.58
+ $Y=1.84 $X2=0.73 $Y2=2.455
.ends

.subckt PM_SKY130_FD_SC_HS__DFXTP_1%A_454_503# 1 2 9 11 13
r31 11 13 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=2.59 $Y=1.155
+ $X2=2.775 $Y2=1.155
r32 7 11 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.505 $Y=1.24
+ $X2=2.59 $Y2=1.155
r33 7 9 79.5936 $w=1.68e-07 $l=1.22e-06 $layer=LI1_cond $X=2.505 $Y=1.24
+ $X2=2.505 $Y2=2.46
r34 2 9 600 $w=1.7e-07 $l=2.61056e-07 $layer=licon1_PDIFF $count=1 $X=2.27
+ $Y=2.515 $X2=2.505 $Y2=2.46
r35 1 13 182 $w=1.7e-07 $l=6.75574e-07 $layer=licon1_NDIFF $count=1 $X=2.52
+ $Y=0.595 $X2=2.775 $Y2=1.155
.ends

.subckt PM_SKY130_FD_SC_HS__DFXTP_1%Q 1 2 9 14 15 16 17 28
c26 17 0 2.87771e-20 $X=7.835 $Y=0.84
r27 21 28 0.800308 $w=3.58e-07 $l=2.5e-08 $layer=LI1_cond $X=7.895 $Y=0.95
+ $X2=7.895 $Y2=0.925
r28 17 30 8.03084 $w=3.58e-07 $l=1.5e-07 $layer=LI1_cond $X=7.895 $Y=0.98
+ $X2=7.895 $Y2=1.13
r29 17 21 0.960369 $w=3.58e-07 $l=3e-08 $layer=LI1_cond $X=7.895 $Y=0.98
+ $X2=7.895 $Y2=0.95
r30 17 28 0.960369 $w=3.58e-07 $l=3e-08 $layer=LI1_cond $X=7.895 $Y=0.895
+ $X2=7.895 $Y2=0.925
r31 16 17 12.1647 $w=3.58e-07 $l=3.8e-07 $layer=LI1_cond $X=7.895 $Y=0.515
+ $X2=7.895 $Y2=0.895
r32 15 30 58.7166 $w=1.68e-07 $l=9e-07 $layer=LI1_cond $X=7.99 $Y=2.03 $X2=7.99
+ $Y2=1.13
r33 14 15 6.59029 $w=3.58e-07 $l=1.05e-07 $layer=LI1_cond $X=7.895 $Y=2.135
+ $X2=7.895 $Y2=2.03
r34 7 14 2.40092 $w=3.58e-07 $l=7.5e-08 $layer=LI1_cond $X=7.895 $Y=2.21
+ $X2=7.895 $Y2=2.135
r35 7 9 19.3674 $w=3.58e-07 $l=6.05e-07 $layer=LI1_cond $X=7.895 $Y=2.21
+ $X2=7.895 $Y2=2.815
r36 2 14 400 $w=1.7e-07 $l=3.62319e-07 $layer=licon1_PDIFF $count=1 $X=7.73
+ $Y=1.84 $X2=7.88 $Y2=2.135
r37 2 9 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=7.73
+ $Y=1.84 $X2=7.88 $Y2=2.815
r38 1 16 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=7.74
+ $Y=0.37 $X2=7.88 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__DFXTP_1%VGND 1 2 3 4 5 18 22 26 30 34 37 38 39 41 46
+ 51 63 69 70 73 76 79 82
r111 82 83 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=0 $X2=7.44
+ $Y2=0
r112 76 77 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r113 73 74 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r114 70 83 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=0 $X2=7.44
+ $Y2=0
r115 69 70 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=0 $X2=7.92
+ $Y2=0
r116 67 82 8.33247 $w=1.7e-07 $l=1.58e-07 $layer=LI1_cond $X=7.535 $Y=0
+ $X2=7.377 $Y2=0
r117 67 69 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=7.535 $Y=0
+ $X2=7.92 $Y2=0
r118 66 83 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=0 $X2=7.44
+ $Y2=0
r119 65 66 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.96 $Y=0 $X2=6.96
+ $Y2=0
r120 63 82 8.33247 $w=1.7e-07 $l=1.57e-07 $layer=LI1_cond $X=7.22 $Y=0 $X2=7.377
+ $Y2=0
r121 63 65 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=7.22 $Y=0 $X2=6.96
+ $Y2=0
r122 62 66 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6 $Y=0 $X2=6.96
+ $Y2=0
r123 61 62 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6 $Y=0 $X2=6 $Y2=0
r124 59 62 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=4.56 $Y=0 $X2=6
+ $Y2=0
r125 58 61 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=4.56 $Y=0 $X2=6
+ $Y2=0
r126 58 59 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r127 56 79 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.32 $Y=0 $X2=4.195
+ $Y2=0
r128 56 58 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=4.32 $Y=0 $X2=4.56
+ $Y2=0
r129 55 77 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=2.16
+ $Y2=0
r130 54 55 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r131 52 76 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.315 $Y=0 $X2=2.15
+ $Y2=0
r132 52 54 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=2.315 $Y=0
+ $X2=2.64 $Y2=0
r133 51 79 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.07 $Y=0 $X2=4.195
+ $Y2=0
r134 51 54 93.2941 $w=1.68e-07 $l=1.43e-06 $layer=LI1_cond $X=4.07 $Y=0 $X2=2.64
+ $Y2=0
r135 50 77 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r136 50 74 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=0.72
+ $Y2=0
r137 49 50 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r138 47 73 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.795 $Y=0 $X2=0.67
+ $Y2=0
r139 47 49 57.738 $w=1.68e-07 $l=8.85e-07 $layer=LI1_cond $X=0.795 $Y=0 $X2=1.68
+ $Y2=0
r140 46 76 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.985 $Y=0 $X2=2.15
+ $Y2=0
r141 46 49 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.985 $Y=0
+ $X2=1.68 $Y2=0
r142 44 74 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r143 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r144 41 73 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.545 $Y=0 $X2=0.67
+ $Y2=0
r145 41 43 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.545 $Y=0
+ $X2=0.24 $Y2=0
r146 39 59 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=4.56
+ $Y2=0
r147 39 55 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=4.08 $Y=0
+ $X2=2.64 $Y2=0
r148 39 79 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r149 37 61 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=6.23 $Y=0 $X2=6
+ $Y2=0
r150 37 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.23 $Y=0 $X2=6.395
+ $Y2=0
r151 36 65 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=6.56 $Y=0 $X2=6.96
+ $Y2=0
r152 36 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.56 $Y=0 $X2=6.395
+ $Y2=0
r153 32 82 0.751525 $w=3.15e-07 $l=8.5e-08 $layer=LI1_cond $X=7.377 $Y=0.085
+ $X2=7.377 $Y2=0
r154 32 34 15.7318 $w=3.13e-07 $l=4.3e-07 $layer=LI1_cond $X=7.377 $Y=0.085
+ $X2=7.377 $Y2=0.515
r155 28 38 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.395 $Y=0.085
+ $X2=6.395 $Y2=0
r156 28 30 26.0173 $w=3.28e-07 $l=7.45e-07 $layer=LI1_cond $X=6.395 $Y=0.085
+ $X2=6.395 $Y2=0.83
r157 24 79 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.195 $Y=0.085
+ $X2=4.195 $Y2=0
r158 24 26 12.4464 $w=2.48e-07 $l=2.7e-07 $layer=LI1_cond $X=4.195 $Y=0.085
+ $X2=4.195 $Y2=0.355
r159 20 76 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.15 $Y=0.085
+ $X2=2.15 $Y2=0
r160 20 22 13.6198 $w=3.28e-07 $l=3.9e-07 $layer=LI1_cond $X=2.15 $Y=0.085
+ $X2=2.15 $Y2=0.475
r161 16 73 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.67 $Y=0.085
+ $X2=0.67 $Y2=0
r162 16 18 22.3574 $w=2.48e-07 $l=4.85e-07 $layer=LI1_cond $X=0.67 $Y=0.085
+ $X2=0.67 $Y2=0.57
r163 5 34 182 $w=1.7e-07 $l=2.31409e-07 $layer=licon1_NDIFF $count=1 $X=7.245
+ $Y=0.37 $X2=7.415 $Y2=0.515
r164 4 30 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=6.255
+ $Y=0.62 $X2=6.395 $Y2=0.83
r165 3 26 182 $w=1.7e-07 $l=2.85307e-07 $layer=licon1_NDIFF $count=1 $X=4.015
+ $Y=0.505 $X2=4.235 $Y2=0.355
r166 2 22 182 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=1 $X=2.005
+ $Y=0.33 $X2=2.15 $Y2=0.475
r167 1 18 182 $w=1.7e-07 $l=2.60768e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.37 $X2=0.71 $Y2=0.57
.ends

