* File: sky130_fd_sc_hs__a21boi_4.pex.spice
* Created: Tue Sep  1 19:49:28 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HS__A21BOI_4%A1 1 3 6 8 10 13 15 17 20 22 24 27 29 30 31
+ 32 52
c81 32 0 3.82477e-20 $X=1.68 $Y=1.665
c82 22 0 3.82477e-20 $X=1.855 $Y=1.765
c83 20 0 9.07735e-20 $X=1.43 $Y=0.74
c84 6 0 1.44963e-19 $X=0.57 $Y=0.74
r85 52 53 0.651351 $w=3.7e-07 $l=5e-09 $layer=POLY_cond $X=1.855 $Y=1.557
+ $X2=1.86 $Y2=1.557
r86 50 52 33.2189 $w=3.7e-07 $l=2.55e-07 $layer=POLY_cond $X=1.6 $Y=1.557
+ $X2=1.855 $Y2=1.557
r87 50 51 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.6
+ $Y=1.515 $X2=1.6 $Y2=1.515
r88 48 50 22.1459 $w=3.7e-07 $l=1.7e-07 $layer=POLY_cond $X=1.43 $Y=1.557
+ $X2=1.6 $Y2=1.557
r89 47 48 3.25676 $w=3.7e-07 $l=2.5e-08 $layer=POLY_cond $X=1.405 $Y=1.557
+ $X2=1.43 $Y2=1.557
r90 46 51 11.1952 $w=3.48e-07 $l=3.4e-07 $layer=LI1_cond $X=1.26 $Y=1.605
+ $X2=1.6 $Y2=1.605
r91 45 47 18.8892 $w=3.7e-07 $l=1.45e-07 $layer=POLY_cond $X=1.26 $Y=1.557
+ $X2=1.405 $Y2=1.557
r92 45 46 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.26
+ $Y=1.515 $X2=1.26 $Y2=1.515
r93 43 45 33.8703 $w=3.7e-07 $l=2.6e-07 $layer=POLY_cond $X=1 $Y=1.557 $X2=1.26
+ $Y2=1.557
r94 42 43 5.86216 $w=3.7e-07 $l=4.5e-08 $layer=POLY_cond $X=0.955 $Y=1.557 $X2=1
+ $Y2=1.557
r95 40 42 4.55946 $w=3.7e-07 $l=3.5e-08 $layer=POLY_cond $X=0.92 $Y=1.557
+ $X2=0.955 $Y2=1.557
r96 40 41 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.92
+ $Y=1.515 $X2=0.92 $Y2=1.515
r97 38 40 45.5946 $w=3.7e-07 $l=3.5e-07 $layer=POLY_cond $X=0.57 $Y=1.557
+ $X2=0.92 $Y2=1.557
r98 37 38 8.46757 $w=3.7e-07 $l=6.5e-08 $layer=POLY_cond $X=0.505 $Y=1.557
+ $X2=0.57 $Y2=1.557
r99 32 51 2.63416 $w=3.48e-07 $l=8e-08 $layer=LI1_cond $X=1.68 $Y=1.605 $X2=1.6
+ $Y2=1.605
r100 31 46 1.97562 $w=3.48e-07 $l=6e-08 $layer=LI1_cond $X=1.2 $Y=1.605 $X2=1.26
+ $Y2=1.605
r101 31 41 9.21954 $w=3.48e-07 $l=2.8e-07 $layer=LI1_cond $X=1.2 $Y=1.605
+ $X2=0.92 $Y2=1.605
r102 30 41 6.58539 $w=3.48e-07 $l=2e-07 $layer=LI1_cond $X=0.72 $Y=1.605
+ $X2=0.92 $Y2=1.605
r103 29 30 15.8049 $w=3.48e-07 $l=4.8e-07 $layer=LI1_cond $X=0.24 $Y=1.605
+ $X2=0.72 $Y2=1.605
r104 25 53 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.86 $Y=1.35
+ $X2=1.86 $Y2=1.557
r105 25 27 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.86 $Y=1.35
+ $X2=1.86 $Y2=0.74
r106 22 52 23.9667 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=1.855 $Y=1.765
+ $X2=1.855 $Y2=1.557
r107 22 24 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.855 $Y=1.765
+ $X2=1.855 $Y2=2.4
r108 18 48 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.43 $Y=1.35
+ $X2=1.43 $Y2=1.557
r109 18 20 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.43 $Y=1.35
+ $X2=1.43 $Y2=0.74
r110 15 47 23.9667 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=1.405 $Y=1.765
+ $X2=1.405 $Y2=1.557
r111 15 17 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.405 $Y=1.765
+ $X2=1.405 $Y2=2.4
r112 11 43 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1 $Y=1.35 $X2=1
+ $Y2=1.557
r113 11 13 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1 $Y=1.35 $X2=1
+ $Y2=0.74
r114 8 42 23.9667 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=0.955 $Y=1.765
+ $X2=0.955 $Y2=1.557
r115 8 10 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.955 $Y=1.765
+ $X2=0.955 $Y2=2.4
r116 4 38 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.57 $Y=1.35
+ $X2=0.57 $Y2=1.557
r117 4 6 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=0.57 $Y=1.35 $X2=0.57
+ $Y2=0.74
r118 1 37 23.9667 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=0.505 $Y=1.765
+ $X2=0.505 $Y2=1.557
r119 1 3 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.505 $Y=1.765
+ $X2=0.505 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_HS__A21BOI_4%A2 3 5 7 10 12 14 17 19 21 24 26 28 29 30
+ 31 53
c86 31 0 2.25548e-19 $X=3.6 $Y=1.665
c87 5 0 3.82477e-20 $X=2.305 $Y=1.765
r88 53 54 9.87705 $w=3.66e-07 $l=7.5e-08 $layer=POLY_cond $X=3.58 $Y=1.557
+ $X2=3.655 $Y2=1.557
r89 51 53 3.95082 $w=3.66e-07 $l=3e-08 $layer=POLY_cond $X=3.55 $Y=1.557
+ $X2=3.58 $Y2=1.557
r90 51 52 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.55
+ $Y=1.515 $X2=3.55 $Y2=1.515
r91 49 52 11.1952 $w=3.48e-07 $l=3.4e-07 $layer=LI1_cond $X=3.21 $Y=1.605
+ $X2=3.55 $Y2=1.605
r92 48 51 44.776 $w=3.66e-07 $l=3.4e-07 $layer=POLY_cond $X=3.21 $Y=1.557
+ $X2=3.55 $Y2=1.557
r93 48 49 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.21
+ $Y=1.515 $X2=3.21 $Y2=1.515
r94 46 48 0.65847 $w=3.66e-07 $l=5e-09 $layer=POLY_cond $X=3.205 $Y=1.557
+ $X2=3.21 $Y2=1.557
r95 45 46 7.24317 $w=3.66e-07 $l=5.5e-08 $layer=POLY_cond $X=3.15 $Y=1.557
+ $X2=3.205 $Y2=1.557
r96 43 45 36.8743 $w=3.66e-07 $l=2.8e-07 $layer=POLY_cond $X=2.87 $Y=1.557
+ $X2=3.15 $Y2=1.557
r97 43 44 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.87
+ $Y=1.515 $X2=2.87 $Y2=1.515
r98 41 43 15.1448 $w=3.66e-07 $l=1.15e-07 $layer=POLY_cond $X=2.755 $Y=1.557
+ $X2=2.87 $Y2=1.557
r99 40 41 4.60929 $w=3.66e-07 $l=3.5e-08 $layer=POLY_cond $X=2.72 $Y=1.557
+ $X2=2.755 $Y2=1.557
r100 38 40 25.0219 $w=3.66e-07 $l=1.9e-07 $layer=POLY_cond $X=2.53 $Y=1.557
+ $X2=2.72 $Y2=1.557
r101 38 39 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.53
+ $Y=1.515 $X2=2.53 $Y2=1.515
r102 36 38 29.6311 $w=3.66e-07 $l=2.25e-07 $layer=POLY_cond $X=2.305 $Y=1.557
+ $X2=2.53 $Y2=1.557
r103 35 36 1.97541 $w=3.66e-07 $l=1.5e-08 $layer=POLY_cond $X=2.29 $Y=1.557
+ $X2=2.305 $Y2=1.557
r104 31 52 1.64635 $w=3.48e-07 $l=5e-08 $layer=LI1_cond $X=3.6 $Y=1.605 $X2=3.55
+ $Y2=1.605
r105 30 49 2.96342 $w=3.48e-07 $l=9e-08 $layer=LI1_cond $X=3.12 $Y=1.605
+ $X2=3.21 $Y2=1.605
r106 30 44 8.23174 $w=3.48e-07 $l=2.5e-07 $layer=LI1_cond $X=3.12 $Y=1.605
+ $X2=2.87 $Y2=1.605
r107 29 44 7.5732 $w=3.48e-07 $l=2.3e-07 $layer=LI1_cond $X=2.64 $Y=1.605
+ $X2=2.87 $Y2=1.605
r108 29 39 3.62196 $w=3.48e-07 $l=1.1e-07 $layer=LI1_cond $X=2.64 $Y=1.605
+ $X2=2.53 $Y2=1.605
r109 26 54 23.7042 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=3.655 $Y=1.765
+ $X2=3.655 $Y2=1.557
r110 26 28 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.655 $Y=1.765
+ $X2=3.655 $Y2=2.4
r111 22 53 23.7042 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.58 $Y=1.35
+ $X2=3.58 $Y2=1.557
r112 22 24 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=3.58 $Y=1.35
+ $X2=3.58 $Y2=0.74
r113 19 46 23.7042 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=3.205 $Y=1.765
+ $X2=3.205 $Y2=1.557
r114 19 21 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.205 $Y=1.765
+ $X2=3.205 $Y2=2.4
r115 15 45 23.7042 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.15 $Y=1.35
+ $X2=3.15 $Y2=1.557
r116 15 17 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=3.15 $Y=1.35
+ $X2=3.15 $Y2=0.74
r117 12 41 23.7042 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=2.755 $Y=1.765
+ $X2=2.755 $Y2=1.557
r118 12 14 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.755 $Y=1.765
+ $X2=2.755 $Y2=2.4
r119 8 40 23.7042 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.72 $Y=1.35
+ $X2=2.72 $Y2=1.557
r120 8 10 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.72 $Y=1.35
+ $X2=2.72 $Y2=0.74
r121 5 36 23.7042 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=2.305 $Y=1.765
+ $X2=2.305 $Y2=1.557
r122 5 7 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.305 $Y=1.765
+ $X2=2.305 $Y2=2.4
r123 1 35 23.7042 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.29 $Y=1.35
+ $X2=2.29 $Y2=1.557
r124 1 3 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.29 $Y=1.35 $X2=2.29
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HS__A21BOI_4%A_803_323# 1 2 7 9 10 11 12 14 17 19 23 25
+ 27 30 32 34 37 41 48 50 51 53 54 57 61 63
c124 63 0 1.00768e-19 $X=6.11 $Y=1.4
c125 50 0 1.93315e-19 $X=6.11 $Y=1.99
c126 48 0 1.04161e-19 $X=5.76 $Y=1.485
c127 25 0 1.60106e-19 $X=5.005 $Y=1.765
c128 11 0 1.72529e-19 $X=4.18 $Y=1.69
c129 7 0 1.47719e-20 $X=4.105 $Y=1.765
r130 67 68 4.55946 $w=3.7e-07 $l=3.5e-08 $layer=POLY_cond $X=5.42 $Y=1.542
+ $X2=5.455 $Y2=1.542
r131 64 65 1.95405 $w=3.7e-07 $l=1.5e-08 $layer=POLY_cond $X=4.99 $Y=1.542
+ $X2=5.005 $Y2=1.542
r132 59 61 4.32166 $w=2.78e-07 $l=1.05e-07 $layer=LI1_cond $X=6.675 $Y=2.16
+ $X2=6.675 $Y2=2.265
r133 55 57 28.1462 $w=2.58e-07 $l=6.35e-07 $layer=LI1_cond $X=6.53 $Y=1.15
+ $X2=6.53 $Y2=0.515
r134 53 59 7.36005 $w=1.7e-07 $l=1.77482e-07 $layer=LI1_cond $X=6.535 $Y=2.075
+ $X2=6.675 $Y2=2.16
r135 53 54 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=6.535 $Y=2.075
+ $X2=6.195 $Y2=2.075
r136 52 63 3.70735 $w=2.5e-07 $l=2.03101e-07 $layer=LI1_cond $X=6.195 $Y=1.235
+ $X2=6.11 $Y2=1.4
r137 51 55 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=6.4 $Y=1.235
+ $X2=6.53 $Y2=1.15
r138 51 52 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=6.4 $Y=1.235
+ $X2=6.195 $Y2=1.235
r139 50 54 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.11 $Y=1.99
+ $X2=6.195 $Y2=2.075
r140 49 63 2.76166 $w=1.7e-07 $l=2.5e-07 $layer=LI1_cond $X=6.11 $Y=1.65
+ $X2=6.11 $Y2=1.4
r141 49 50 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=6.11 $Y=1.65
+ $X2=6.11 $Y2=1.99
r142 48 70 11.7243 $w=3.7e-07 $l=9e-08 $layer=POLY_cond $X=5.76 $Y=1.542
+ $X2=5.85 $Y2=1.542
r143 48 68 39.7324 $w=3.7e-07 $l=3.05e-07 $layer=POLY_cond $X=5.76 $Y=1.542
+ $X2=5.455 $Y2=1.542
r144 47 48 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=5.76
+ $Y=1.485 $X2=5.76 $Y2=1.485
r145 44 67 44.2919 $w=3.7e-07 $l=3.4e-07 $layer=POLY_cond $X=5.08 $Y=1.542
+ $X2=5.42 $Y2=1.542
r146 44 65 9.77027 $w=3.7e-07 $l=7.5e-08 $layer=POLY_cond $X=5.08 $Y=1.542
+ $X2=5.005 $Y2=1.542
r147 43 47 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=5.08 $Y=1.485
+ $X2=5.76 $Y2=1.485
r148 43 44 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=5.08
+ $Y=1.485 $X2=5.08 $Y2=1.485
r149 41 63 3.70735 $w=2.5e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.025 $Y=1.485
+ $X2=6.11 $Y2=1.4
r150 41 47 9.25447 $w=3.28e-07 $l=2.65e-07 $layer=LI1_cond $X=6.025 $Y=1.485
+ $X2=5.76 $Y2=1.485
r151 39 40 34.216 $w=1.62e-07 $l=1.15e-07 $layer=POLY_cond $X=4.562 $Y=1.575
+ $X2=4.562 $Y2=1.69
r152 35 70 23.9667 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=5.85 $Y=1.32
+ $X2=5.85 $Y2=1.542
r153 35 37 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=5.85 $Y=1.32
+ $X2=5.85 $Y2=0.74
r154 32 68 23.9667 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=5.455 $Y=1.765
+ $X2=5.455 $Y2=1.542
r155 32 34 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=5.455 $Y=1.765
+ $X2=5.455 $Y2=2.4
r156 28 67 23.9667 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=5.42 $Y=1.32
+ $X2=5.42 $Y2=1.542
r157 28 30 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=5.42 $Y=1.32
+ $X2=5.42 $Y2=0.74
r158 25 65 23.9667 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=5.005 $Y=1.765
+ $X2=5.005 $Y2=1.542
r159 25 27 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=5.005 $Y=1.765
+ $X2=5.005 $Y2=2.4
r160 21 64 23.9667 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=4.99 $Y=1.32
+ $X2=4.99 $Y2=1.542
r161 21 23 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=4.99 $Y=1.32
+ $X2=4.99 $Y2=0.74
r162 20 39 4.66776 $w=1.5e-07 $l=8.3e-08 $layer=POLY_cond $X=4.645 $Y=1.575
+ $X2=4.562 $Y2=1.575
r163 19 64 27.3315 $w=3.7e-07 $l=9e-08 $layer=POLY_cond $X=4.915 $Y=1.575
+ $X2=4.99 $Y2=1.542
r164 19 20 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=4.915 $Y=1.575
+ $X2=4.645 $Y2=1.575
r165 15 39 22.6565 $w=1.62e-07 $l=7.59934e-08 $layer=POLY_cond $X=4.56 $Y=1.5
+ $X2=4.562 $Y2=1.575
r166 15 17 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=4.56 $Y=1.5
+ $X2=4.56 $Y2=0.74
r167 12 40 22.6565 $w=1.62e-07 $l=7.84219e-08 $layer=POLY_cond $X=4.555 $Y=1.765
+ $X2=4.562 $Y2=1.69
r168 12 14 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=4.555 $Y=1.765
+ $X2=4.555 $Y2=2.4
r169 10 40 4.66776 $w=1.5e-07 $l=8.2e-08 $layer=POLY_cond $X=4.48 $Y=1.69
+ $X2=4.562 $Y2=1.69
r170 10 11 153.83 $w=1.5e-07 $l=3e-07 $layer=POLY_cond $X=4.48 $Y=1.69 $X2=4.18
+ $Y2=1.69
r171 7 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.105 $Y=1.765
+ $X2=4.18 $Y2=1.69
r172 7 9 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=4.105 $Y=1.765
+ $X2=4.105 $Y2=2.4
r173 2 61 300 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=2 $X=6.5
+ $Y=2.12 $X2=6.65 $Y2=2.265
r174 1 57 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=6.355
+ $Y=0.37 $X2=6.495 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__A21BOI_4%B1_N 3 5 7 8 10 11 12 13 20
c37 20 0 1.00768e-19 $X=6.53 $Y=1.655
c38 13 0 1.04161e-19 $X=7.44 $Y=1.665
r39 20 22 41.0593 $w=4.05e-07 $l=3.45e-07 $layer=POLY_cond $X=6.53 $Y=1.767
+ $X2=6.875 $Y2=1.767
r40 18 20 12.4963 $w=4.05e-07 $l=1.05e-07 $layer=POLY_cond $X=6.425 $Y=1.767
+ $X2=6.53 $Y2=1.767
r41 12 13 16.7628 $w=3.28e-07 $l=4.8e-07 $layer=LI1_cond $X=6.96 $Y=1.655
+ $X2=7.44 $Y2=1.655
r42 11 12 16.7628 $w=3.28e-07 $l=4.8e-07 $layer=LI1_cond $X=6.48 $Y=1.655
+ $X2=6.96 $Y2=1.655
r43 11 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.53
+ $Y=1.655 $X2=6.53 $Y2=1.655
r44 8 22 26.1659 $w=1.5e-07 $l=2.78e-07 $layer=POLY_cond $X=6.875 $Y=2.045
+ $X2=6.875 $Y2=1.767
r45 8 10 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=6.875 $Y=2.045
+ $X2=6.875 $Y2=2.54
r46 5 18 26.1659 $w=1.5e-07 $l=2.78e-07 $layer=POLY_cond $X=6.425 $Y=2.045
+ $X2=6.425 $Y2=1.767
r47 5 7 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=6.425 $Y=2.045
+ $X2=6.425 $Y2=2.54
r48 1 18 17.2568 $w=4.05e-07 $l=3.41898e-07 $layer=POLY_cond $X=6.28 $Y=1.49
+ $X2=6.425 $Y2=1.767
r49 1 3 384.574 $w=1.5e-07 $l=7.5e-07 $layer=POLY_cond $X=6.28 $Y=1.49 $X2=6.28
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HS__A21BOI_4%A_31_368# 1 2 3 4 5 6 7 22 24 26 30 32 36
+ 38 42 44 46 49 50 51 54 56 60 67 69 71 74
r108 60 63 34.1617 $w=2.78e-07 $l=8.3e-07 $layer=LI1_cond $X=5.705 $Y=1.985
+ $X2=5.705 $Y2=2.815
r109 58 63 3.70428 $w=2.78e-07 $l=9e-08 $layer=LI1_cond $X=5.705 $Y=2.905
+ $X2=5.705 $Y2=2.815
r110 57 74 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=4.895 $Y=2.99
+ $X2=4.78 $Y2=2.99
r111 56 58 7.36005 $w=1.7e-07 $l=1.77482e-07 $layer=LI1_cond $X=5.565 $Y=2.99
+ $X2=5.705 $Y2=2.905
r112 56 57 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.565 $Y=2.99
+ $X2=4.895 $Y2=2.99
r113 52 74 0.280307 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.78 $Y=2.905
+ $X2=4.78 $Y2=2.99
r114 52 54 29.0616 $w=2.28e-07 $l=5.8e-07 $layer=LI1_cond $X=4.78 $Y=2.905
+ $X2=4.78 $Y2=2.325
r115 50 74 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=4.665 $Y=2.99
+ $X2=4.78 $Y2=2.99
r116 50 51 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.665 $Y=2.99
+ $X2=3.995 $Y2=2.99
r117 47 51 7.36005 $w=1.7e-07 $l=1.77482e-07 $layer=LI1_cond $X=3.855 $Y=2.905
+ $X2=3.995 $Y2=2.99
r118 47 49 3.70428 $w=2.78e-07 $l=9e-08 $layer=LI1_cond $X=3.855 $Y=2.905
+ $X2=3.855 $Y2=2.815
r119 46 73 2.78046 $w=2.8e-07 $l=8.5e-08 $layer=LI1_cond $X=3.855 $Y=2.12
+ $X2=3.855 $Y2=2.035
r120 46 49 28.6053 $w=2.78e-07 $l=6.95e-07 $layer=LI1_cond $X=3.855 $Y=2.12
+ $X2=3.855 $Y2=2.815
r121 45 71 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.145 $Y=2.035
+ $X2=2.98 $Y2=2.035
r122 44 73 4.57959 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=3.715 $Y=2.035
+ $X2=3.855 $Y2=2.035
r123 44 45 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=3.715 $Y=2.035
+ $X2=3.145 $Y2=2.035
r124 40 71 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.98 $Y=2.12
+ $X2=2.98 $Y2=2.035
r125 40 42 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=2.98 $Y=2.12
+ $X2=2.98 $Y2=2.815
r126 39 69 5.16603 $w=1.7e-07 $l=1.12916e-07 $layer=LI1_cond $X=2.165 $Y=2.035
+ $X2=2.08 $Y2=1.97
r127 38 71 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.815 $Y=2.035
+ $X2=2.98 $Y2=2.035
r128 38 39 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=2.815 $Y=2.035
+ $X2=2.165 $Y2=2.035
r129 34 69 1.34256 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=2.08 $Y=2.12
+ $X2=2.08 $Y2=1.97
r130 34 36 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=2.08 $Y=2.12
+ $X2=2.08 $Y2=2.4
r131 33 67 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.265 $Y=2.035
+ $X2=1.18 $Y2=2.035
r132 32 69 5.16603 $w=1.7e-07 $l=1.12916e-07 $layer=LI1_cond $X=1.995 $Y=2.035
+ $X2=2.08 $Y2=1.97
r133 32 33 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=1.995 $Y=2.035
+ $X2=1.265 $Y2=2.035
r134 28 67 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.18 $Y=2.12
+ $X2=1.18 $Y2=2.035
r135 28 30 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=1.18 $Y=2.12
+ $X2=1.18 $Y2=2.815
r136 27 65 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.365 $Y=2.035
+ $X2=0.24 $Y2=2.035
r137 26 67 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.095 $Y=2.035
+ $X2=1.18 $Y2=2.035
r138 26 27 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=1.095 $Y=2.035
+ $X2=0.365 $Y2=2.035
r139 22 65 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.24 $Y=2.12
+ $X2=0.24 $Y2=2.035
r140 22 24 32.0379 $w=2.48e-07 $l=6.95e-07 $layer=LI1_cond $X=0.24 $Y=2.12
+ $X2=0.24 $Y2=2.815
r141 7 63 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=5.53
+ $Y=1.84 $X2=5.68 $Y2=2.815
r142 7 60 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=5.53
+ $Y=1.84 $X2=5.68 $Y2=1.985
r143 6 54 300 $w=1.7e-07 $l=5.54955e-07 $layer=licon1_PDIFF $count=2 $X=4.63
+ $Y=1.84 $X2=4.78 $Y2=2.325
r144 5 73 400 $w=1.7e-07 $l=3.4187e-07 $layer=licon1_PDIFF $count=1 $X=3.73
+ $Y=1.84 $X2=3.88 $Y2=2.115
r145 5 49 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=3.73
+ $Y=1.84 $X2=3.88 $Y2=2.815
r146 4 71 400 $w=1.7e-07 $l=3.4187e-07 $layer=licon1_PDIFF $count=1 $X=2.83
+ $Y=1.84 $X2=2.98 $Y2=2.115
r147 4 42 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=2.83
+ $Y=1.84 $X2=2.98 $Y2=2.815
r148 3 69 600 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=1.93
+ $Y=1.84 $X2=2.08 $Y2=1.985
r149 3 36 300 $w=1.7e-07 $l=6.30555e-07 $layer=licon1_PDIFF $count=2 $X=1.93
+ $Y=1.84 $X2=2.08 $Y2=2.4
r150 2 67 400 $w=1.7e-07 $l=3.4187e-07 $layer=licon1_PDIFF $count=1 $X=1.03
+ $Y=1.84 $X2=1.18 $Y2=2.115
r151 2 30 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=1.03
+ $Y=1.84 $X2=1.18 $Y2=2.815
r152 1 65 400 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_PDIFF $count=1 $X=0.155
+ $Y=1.84 $X2=0.28 $Y2=2.115
r153 1 24 400 $w=1.7e-07 $l=1.03562e-06 $layer=licon1_PDIFF $count=1 $X=0.155
+ $Y=1.84 $X2=0.28 $Y2=2.815
.ends

.subckt PM_SKY130_FD_SC_HS__A21BOI_4%VPWR 1 2 3 4 5 6 21 25 29 33 37 41 44 45 47
+ 48 50 51 53 54 55 57 62 84 85 88 91
r110 91 92 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r111 88 89 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r112 84 85 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r113 82 85 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=7.44 $Y2=3.33
r114 81 82 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r115 79 82 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6 $Y=3.33 $X2=6.96
+ $Y2=3.33
r116 78 79 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r117 75 78 156.578 $w=1.68e-07 $l=2.4e-06 $layer=LI1_cond $X=3.6 $Y=3.33 $X2=6
+ $Y2=3.33
r118 75 76 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r119 73 76 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=3.6 $Y2=3.33
r120 72 73 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r121 70 73 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=3.12 $Y2=3.33
r122 70 92 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.68 $Y2=3.33
r123 69 70 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r124 67 91 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.795 $Y=3.33
+ $X2=1.63 $Y2=3.33
r125 67 69 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=1.795 $Y=3.33
+ $X2=2.16 $Y2=3.33
r126 66 92 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=1.68 $Y2=3.33
r127 66 89 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r128 65 66 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r129 63 88 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.895 $Y=3.33
+ $X2=0.73 $Y2=3.33
r130 63 65 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.895 $Y=3.33
+ $X2=1.2 $Y2=3.33
r131 62 91 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.465 $Y=3.33
+ $X2=1.63 $Y2=3.33
r132 62 65 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=1.465 $Y=3.33
+ $X2=1.2 $Y2=3.33
r133 60 89 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r134 59 60 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r135 57 88 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.565 $Y=3.33
+ $X2=0.73 $Y2=3.33
r136 57 59 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.565 $Y=3.33
+ $X2=0.24 $Y2=3.33
r137 55 79 0.602067 $w=4.9e-07 $l=2.16e-06 $layer=MET1_cond $X=3.84 $Y=3.33
+ $X2=6 $Y2=3.33
r138 55 76 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=3.84 $Y=3.33
+ $X2=3.6 $Y2=3.33
r139 53 81 3.58824 $w=1.68e-07 $l=5.5e-08 $layer=LI1_cond $X=7.015 $Y=3.33
+ $X2=6.96 $Y2=3.33
r140 53 54 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.015 $Y=3.33
+ $X2=7.14 $Y2=3.33
r141 52 84 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=7.265 $Y=3.33
+ $X2=7.44 $Y2=3.33
r142 52 54 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.265 $Y=3.33
+ $X2=7.14 $Y2=3.33
r143 50 78 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=6.035 $Y=3.33 $X2=6
+ $Y2=3.33
r144 50 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.035 $Y=3.33
+ $X2=6.2 $Y2=3.33
r145 49 81 38.8182 $w=1.68e-07 $l=5.95e-07 $layer=LI1_cond $X=6.365 $Y=3.33
+ $X2=6.96 $Y2=3.33
r146 49 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.365 $Y=3.33
+ $X2=6.2 $Y2=3.33
r147 47 72 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=3.345 $Y=3.33
+ $X2=3.12 $Y2=3.33
r148 47 48 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.345 $Y=3.33
+ $X2=3.43 $Y2=3.33
r149 46 75 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=3.515 $Y=3.33
+ $X2=3.6 $Y2=3.33
r150 46 48 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.515 $Y=3.33
+ $X2=3.43 $Y2=3.33
r151 44 69 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=2.365 $Y=3.33
+ $X2=2.16 $Y2=3.33
r152 44 45 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.365 $Y=3.33
+ $X2=2.49 $Y2=3.33
r153 43 72 32.9465 $w=1.68e-07 $l=5.05e-07 $layer=LI1_cond $X=2.615 $Y=3.33
+ $X2=3.12 $Y2=3.33
r154 43 45 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.615 $Y=3.33
+ $X2=2.49 $Y2=3.33
r155 39 54 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=7.14 $Y=3.245
+ $X2=7.14 $Y2=3.33
r156 39 41 45.1758 $w=2.48e-07 $l=9.8e-07 $layer=LI1_cond $X=7.14 $Y=3.245
+ $X2=7.14 $Y2=2.265
r157 35 51 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.2 $Y=3.245 $X2=6.2
+ $Y2=3.33
r158 35 37 27.938 $w=3.28e-07 $l=8e-07 $layer=LI1_cond $X=6.2 $Y=3.245 $X2=6.2
+ $Y2=2.445
r159 31 48 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.43 $Y=3.245
+ $X2=3.43 $Y2=3.33
r160 31 33 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=3.43 $Y=3.245
+ $X2=3.43 $Y2=2.455
r161 27 45 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.49 $Y=3.245
+ $X2=2.49 $Y2=3.33
r162 27 29 36.4172 $w=2.48e-07 $l=7.9e-07 $layer=LI1_cond $X=2.49 $Y=3.245
+ $X2=2.49 $Y2=2.455
r163 23 91 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.63 $Y=3.245
+ $X2=1.63 $Y2=3.33
r164 23 25 27.5888 $w=3.28e-07 $l=7.9e-07 $layer=LI1_cond $X=1.63 $Y=3.245
+ $X2=1.63 $Y2=2.455
r165 19 88 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.73 $Y=3.245
+ $X2=0.73 $Y2=3.33
r166 19 21 27.5888 $w=3.28e-07 $l=7.9e-07 $layer=LI1_cond $X=0.73 $Y=3.245
+ $X2=0.73 $Y2=2.455
r167 6 41 300 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=2 $X=6.95
+ $Y=2.12 $X2=7.1 $Y2=2.265
r168 5 37 300 $w=1.7e-07 $l=3.82426e-07 $layer=licon1_PDIFF $count=2 $X=6.075
+ $Y=2.12 $X2=6.2 $Y2=2.445
r169 4 33 300 $w=1.7e-07 $l=6.85912e-07 $layer=licon1_PDIFF $count=2 $X=3.28
+ $Y=1.84 $X2=3.43 $Y2=2.455
r170 3 29 300 $w=1.7e-07 $l=6.85912e-07 $layer=licon1_PDIFF $count=2 $X=2.38
+ $Y=1.84 $X2=2.53 $Y2=2.455
r171 2 25 300 $w=1.7e-07 $l=6.85912e-07 $layer=licon1_PDIFF $count=2 $X=1.48
+ $Y=1.84 $X2=1.63 $Y2=2.455
r172 1 21 300 $w=1.7e-07 $l=6.85912e-07 $layer=licon1_PDIFF $count=2 $X=0.58
+ $Y=1.84 $X2=0.73 $Y2=2.455
.ends

.subckt PM_SKY130_FD_SC_HS__A21BOI_4%Y 1 2 3 4 5 6 19 21 23 25 29 31 33 35 37 41
+ 43 48 56 57
c111 43 0 1.44963e-19 $X=0.825 $Y=0.855
c112 23 0 1.60106e-19 $X=4.33 $Y=1.99
c113 21 0 9.07735e-20 $X=3.965 $Y=1.175
r114 56 57 6.53256 $w=6.91e-07 $l=3.7e-07 $layer=LI1_cond $X=4.412 $Y=1.295
+ $X2=4.412 $Y2=1.665
r115 56 65 2.11867 $w=6.91e-07 $l=1.2e-07 $layer=LI1_cond $X=4.412 $Y=1.295
+ $X2=4.412 $Y2=1.175
r116 51 52 7.85757 $w=3.28e-07 $l=2.25e-07 $layer=LI1_cond $X=1.645 $Y=0.95
+ $X2=1.645 $Y2=1.175
r117 48 51 3.31764 $w=3.28e-07 $l=9.5e-08 $layer=LI1_cond $X=1.645 $Y=0.855
+ $X2=1.645 $Y2=0.95
r118 43 46 4.37928 $w=2.48e-07 $l=9.5e-08 $layer=LI1_cond $X=0.825 $Y=0.855
+ $X2=0.825 $Y2=0.95
r119 39 41 21.4354 $w=2.48e-07 $l=4.65e-07 $layer=LI1_cond $X=5.595 $Y=0.98
+ $X2=5.595 $Y2=0.515
r120 35 55 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.23 $Y=1.99 $X2=5.23
+ $Y2=1.905
r121 35 37 23.0489 $w=3.28e-07 $l=6.6e-07 $layer=LI1_cond $X=5.23 $Y=1.99
+ $X2=5.23 $Y2=2.65
r122 34 65 1.94211 $w=6.91e-07 $l=4.99984e-07 $layer=LI1_cond $X=4.86 $Y=1.065
+ $X2=4.412 $Y2=1.175
r123 33 39 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=5.47 $Y=1.065
+ $X2=5.595 $Y2=0.98
r124 33 34 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=5.47 $Y=1.065
+ $X2=4.86 $Y2=1.065
r125 32 74 1.14761 $w=6.91e-07 $l=6.5e-08 $layer=LI1_cond $X=4.412 $Y=1.905
+ $X2=4.412 $Y2=1.97
r126 32 57 4.23734 $w=6.91e-07 $l=2.4e-07 $layer=LI1_cond $X=4.412 $Y=1.905
+ $X2=4.412 $Y2=1.665
r127 31 55 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.065 $Y=1.905
+ $X2=5.23 $Y2=1.905
r128 31 32 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=5.065 $Y=1.905
+ $X2=4.745 $Y2=1.905
r129 27 34 6.74026 $w=6.91e-07 $l=1.62019e-07 $layer=LI1_cond $X=4.735 $Y=0.98
+ $X2=4.86 $Y2=1.065
r130 27 29 21.4354 $w=2.48e-07 $l=4.65e-07 $layer=LI1_cond $X=4.735 $Y=0.98
+ $X2=4.735 $Y2=0.515
r131 23 74 3.69776 $w=6.91e-07 $l=9.14549e-08 $layer=LI1_cond $X=4.33 $Y=1.99
+ $X2=4.412 $Y2=1.97
r132 23 25 23.0489 $w=3.28e-07 $l=6.6e-07 $layer=LI1_cond $X=4.33 $Y=1.99
+ $X2=4.33 $Y2=2.65
r133 22 52 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.81 $Y=1.175
+ $X2=1.645 $Y2=1.175
r134 21 65 9.23635 $w=1.7e-07 $l=4.47e-07 $layer=LI1_cond $X=3.965 $Y=1.175
+ $X2=4.412 $Y2=1.175
r135 21 22 140.594 $w=1.68e-07 $l=2.155e-06 $layer=LI1_cond $X=3.965 $Y=1.175
+ $X2=1.81 $Y2=1.175
r136 20 43 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.95 $Y=0.855
+ $X2=0.825 $Y2=0.855
r137 19 48 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.48 $Y=0.855
+ $X2=1.645 $Y2=0.855
r138 19 20 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=1.48 $Y=0.855
+ $X2=0.95 $Y2=0.855
r139 6 55 400 $w=1.7e-07 $l=2.04939e-07 $layer=licon1_PDIFF $count=1 $X=5.08
+ $Y=1.84 $X2=5.23 $Y2=1.97
r140 6 37 400 $w=1.7e-07 $l=8.81816e-07 $layer=licon1_PDIFF $count=1 $X=5.08
+ $Y=1.84 $X2=5.23 $Y2=2.65
r141 5 74 400 $w=1.7e-07 $l=2.04939e-07 $layer=licon1_PDIFF $count=1 $X=4.18
+ $Y=1.84 $X2=4.33 $Y2=1.97
r142 5 25 400 $w=1.7e-07 $l=8.81816e-07 $layer=licon1_PDIFF $count=1 $X=4.18
+ $Y=1.84 $X2=4.33 $Y2=2.65
r143 4 41 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=5.495
+ $Y=0.37 $X2=5.635 $Y2=0.515
r144 3 29 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=4.635
+ $Y=0.37 $X2=4.775 $Y2=0.515
r145 2 51 182 $w=1.7e-07 $l=6.4622e-07 $layer=licon1_NDIFF $count=1 $X=1.505
+ $Y=0.37 $X2=1.645 $Y2=0.95
r146 1 46 182 $w=1.7e-07 $l=6.4622e-07 $layer=licon1_NDIFF $count=1 $X=0.645
+ $Y=0.37 $X2=0.785 $Y2=0.95
.ends

.subckt PM_SKY130_FD_SC_HS__A21BOI_4%A_46_74# 1 2 3 4 5 18 26 27 28 31 33 38
r54 38 40 5.07075 $w=2.48e-07 $l=1.1e-07 $layer=LI1_cond $X=3.835 $Y=0.725
+ $X2=3.835 $Y2=0.835
r55 33 35 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=2.935 $Y=0.725
+ $X2=2.935 $Y2=0.835
r56 29 35 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.02 $Y=0.835
+ $X2=2.935 $Y2=0.835
r57 28 40 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.71 $Y=0.835
+ $X2=3.835 $Y2=0.835
r58 28 29 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=3.71 $Y=0.835
+ $X2=3.02 $Y2=0.835
r59 26 35 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.85 $Y=0.835
+ $X2=2.935 $Y2=0.835
r60 26 27 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=2.85 $Y=0.835
+ $X2=2.16 $Y2=0.835
r61 23 27 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.075 $Y=0.75
+ $X2=2.16 $Y2=0.835
r62 23 25 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=2.075 $Y=0.75
+ $X2=2.075 $Y2=0.725
r63 22 25 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=2.075 $Y=0.6
+ $X2=2.075 $Y2=0.725
r64 19 31 3.97509 $w=2.5e-07 $l=1.65e-07 $layer=LI1_cond $X=0.52 $Y=0.475
+ $X2=0.355 $Y2=0.475
r65 19 21 32.0379 $w=2.48e-07 $l=6.95e-07 $layer=LI1_cond $X=0.52 $Y=0.475
+ $X2=1.215 $Y2=0.475
r66 18 22 7.14316 $w=2.5e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.99 $Y=0.475
+ $X2=2.075 $Y2=0.6
r67 18 21 35.7257 $w=2.48e-07 $l=7.75e-07 $layer=LI1_cond $X=1.99 $Y=0.475
+ $X2=1.215 $Y2=0.475
r68 5 38 182 $w=1.7e-07 $l=4.19196e-07 $layer=licon1_NDIFF $count=1 $X=3.655
+ $Y=0.37 $X2=3.795 $Y2=0.725
r69 4 33 182 $w=1.7e-07 $l=4.19196e-07 $layer=licon1_NDIFF $count=1 $X=2.795
+ $Y=0.37 $X2=2.935 $Y2=0.725
r70 3 25 182 $w=1.7e-07 $l=4.19196e-07 $layer=licon1_NDIFF $count=1 $X=1.935
+ $Y=0.37 $X2=2.075 $Y2=0.725
r71 2 21 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=1.075
+ $Y=0.37 $X2=1.215 $Y2=0.515
r72 1 31 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.23
+ $Y=0.37 $X2=0.355 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__A21BOI_4%VGND 1 2 3 4 5 18 22 26 28 32 36 39 40 42
+ 43 44 45 46 61 71 72 75 78
r98 78 79 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=0 $X2=6 $Y2=0
r99 75 76 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r100 71 72 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=7.44 $Y=0 $X2=7.44
+ $Y2=0
r101 69 72 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.48 $Y=0 $X2=7.44
+ $Y2=0
r102 69 79 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=0 $X2=6
+ $Y2=0
r103 68 71 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=6.48 $Y=0 $X2=7.44
+ $Y2=0
r104 68 69 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6.48 $Y=0 $X2=6.48
+ $Y2=0
r105 66 78 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.23 $Y=0 $X2=6.065
+ $Y2=0
r106 66 68 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=6.23 $Y=0 $X2=6.48
+ $Y2=0
r107 65 79 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=6
+ $Y2=0
r108 65 76 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=5.04
+ $Y2=0
r109 64 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r110 62 75 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.29 $Y=0 $X2=5.165
+ $Y2=0
r111 62 64 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=5.29 $Y=0 $X2=5.52
+ $Y2=0
r112 61 78 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.9 $Y=0 $X2=6.065
+ $Y2=0
r113 61 64 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=5.9 $Y=0 $X2=5.52
+ $Y2=0
r114 60 76 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=5.04
+ $Y2=0
r115 59 60 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r116 56 57 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r117 54 57 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=3.12
+ $Y2=0
r118 53 54 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.16 $Y=0
+ $X2=2.16 $Y2=0
r119 50 54 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=0.24 $Y=0
+ $X2=2.16 $Y2=0
r120 49 53 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=0.24 $Y=0 $X2=2.16
+ $Y2=0
r121 49 50 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.24 $Y=0
+ $X2=0.24 $Y2=0
r122 46 60 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=3.84 $Y=0
+ $X2=4.08 $Y2=0
r123 46 57 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=3.84 $Y=0 $X2=3.12
+ $Y2=0
r124 44 59 6.52406 $w=1.68e-07 $l=1e-07 $layer=LI1_cond $X=4.18 $Y=0 $X2=4.08
+ $Y2=0
r125 44 45 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.18 $Y=0 $X2=4.305
+ $Y2=0
r126 42 56 5.21925 $w=1.68e-07 $l=8e-08 $layer=LI1_cond $X=3.2 $Y=0 $X2=3.12
+ $Y2=0
r127 42 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.2 $Y=0 $X2=3.365
+ $Y2=0
r128 41 59 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=3.53 $Y=0 $X2=4.08
+ $Y2=0
r129 41 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.53 $Y=0 $X2=3.365
+ $Y2=0
r130 39 53 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=2.34 $Y=0 $X2=2.16
+ $Y2=0
r131 39 40 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.34 $Y=0 $X2=2.505
+ $Y2=0
r132 38 56 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=2.67 $Y=0 $X2=3.12
+ $Y2=0
r133 38 40 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.67 $Y=0 $X2=2.505
+ $Y2=0
r134 34 78 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.065 $Y=0.085
+ $X2=6.065 $Y2=0
r135 34 36 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=6.065 $Y=0.085
+ $X2=6.065 $Y2=0.495
r136 30 75 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.165 $Y=0.085
+ $X2=5.165 $Y2=0
r137 30 32 25.8147 $w=2.48e-07 $l=5.6e-07 $layer=LI1_cond $X=5.165 $Y=0.085
+ $X2=5.165 $Y2=0.645
r138 29 45 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.43 $Y=0 $X2=4.305
+ $Y2=0
r139 28 75 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.04 $Y=0 $X2=5.165
+ $Y2=0
r140 28 29 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=5.04 $Y=0 $X2=4.43
+ $Y2=0
r141 24 45 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.305 $Y=0.085
+ $X2=4.305 $Y2=0
r142 24 26 29.0416 $w=2.48e-07 $l=6.3e-07 $layer=LI1_cond $X=4.305 $Y=0.085
+ $X2=4.305 $Y2=0.715
r143 20 43 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.365 $Y=0.085
+ $X2=3.365 $Y2=0
r144 20 22 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=3.365 $Y=0.085
+ $X2=3.365 $Y2=0.495
r145 16 40 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.505 $Y=0.085
+ $X2=2.505 $Y2=0
r146 16 18 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=2.505 $Y=0.085
+ $X2=2.505 $Y2=0.495
r147 5 36 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=5.925
+ $Y=0.37 $X2=6.065 $Y2=0.495
r148 4 32 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=5.065
+ $Y=0.37 $X2=5.205 $Y2=0.645
r149 3 26 182 $w=1.7e-07 $l=4.02679e-07 $layer=licon1_NDIFF $count=1 $X=4.22
+ $Y=0.37 $X2=4.345 $Y2=0.715
r150 2 22 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=3.225
+ $Y=0.37 $X2=3.365 $Y2=0.495
r151 1 18 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=2.365
+ $Y=0.37 $X2=2.505 $Y2=0.495
.ends

