* File: sky130_fd_sc_hs__ebufn_8.pxi.spice
* Created: Thu Aug 27 20:44:20 2020
* 
x_PM_SKY130_FD_SC_HS__EBUFN_8%A_84_48# N_A_84_48#_M1008_d N_A_84_48#_M1000_d
+ N_A_84_48#_M1005_g N_A_84_48#_c_218_n N_A_84_48#_M1006_g N_A_84_48#_M1009_g
+ N_A_84_48#_c_219_n N_A_84_48#_M1010_g N_A_84_48#_M1011_g N_A_84_48#_c_220_n
+ N_A_84_48#_M1013_g N_A_84_48#_M1029_g N_A_84_48#_c_221_n N_A_84_48#_M1014_g
+ N_A_84_48#_M1032_g N_A_84_48#_c_222_n N_A_84_48#_M1015_g N_A_84_48#_M1033_g
+ N_A_84_48#_c_223_n N_A_84_48#_M1017_g N_A_84_48#_c_224_n N_A_84_48#_M1019_g
+ N_A_84_48#_M1034_g N_A_84_48#_c_225_n N_A_84_48#_M1020_g N_A_84_48#_M1036_g
+ N_A_84_48#_c_329_p N_A_84_48#_c_214_n N_A_84_48#_c_226_n N_A_84_48#_c_242_p
+ N_A_84_48#_c_293_p N_A_84_48#_c_227_n N_A_84_48#_c_238_p N_A_84_48#_c_228_n
+ N_A_84_48#_c_275_p N_A_84_48#_c_215_n N_A_84_48#_c_280_p N_A_84_48#_c_229_n
+ N_A_84_48#_c_230_n N_A_84_48#_c_216_n N_A_84_48#_c_258_p N_A_84_48#_c_274_p
+ N_A_84_48#_c_217_n PM_SKY130_FD_SC_HS__EBUFN_8%A_84_48#
x_PM_SKY130_FD_SC_HS__EBUFN_8%A_833_48# N_A_833_48#_M1031_s N_A_833_48#_M1002_s
+ N_A_833_48#_c_478_n N_A_833_48#_M1001_g N_A_833_48#_c_479_n
+ N_A_833_48#_c_480_n N_A_833_48#_c_481_n N_A_833_48#_M1003_g
+ N_A_833_48#_c_482_n N_A_833_48#_c_483_n N_A_833_48#_M1004_g
+ N_A_833_48#_c_484_n N_A_833_48#_c_485_n N_A_833_48#_M1012_g
+ N_A_833_48#_c_486_n N_A_833_48#_c_487_n N_A_833_48#_M1025_g
+ N_A_833_48#_c_488_n N_A_833_48#_c_489_n N_A_833_48#_M1027_g
+ N_A_833_48#_c_490_n N_A_833_48#_c_491_n N_A_833_48#_M1035_g
+ N_A_833_48#_c_492_n N_A_833_48#_c_493_n N_A_833_48#_M1037_g
+ N_A_833_48#_c_494_n N_A_833_48#_c_495_n N_A_833_48#_c_496_n
+ N_A_833_48#_c_497_n N_A_833_48#_c_498_n N_A_833_48#_c_499_n
+ N_A_833_48#_c_500_n N_A_833_48#_c_501_n N_A_833_48#_c_502_n
+ N_A_833_48#_c_503_n N_A_833_48#_c_504_n N_A_833_48#_c_505_n
+ N_A_833_48#_c_506_n N_A_833_48#_c_507_n N_A_833_48#_c_513_n
+ N_A_833_48#_c_509_n PM_SKY130_FD_SC_HS__EBUFN_8%A_833_48#
x_PM_SKY130_FD_SC_HS__EBUFN_8%TE_B N_TE_B_c_664_n N_TE_B_M1016_g N_TE_B_c_643_n
+ N_TE_B_c_644_n N_TE_B_c_667_n N_TE_B_M1021_g N_TE_B_c_645_n N_TE_B_c_669_n
+ N_TE_B_M1022_g N_TE_B_c_646_n N_TE_B_c_671_n N_TE_B_M1023_g N_TE_B_c_647_n
+ N_TE_B_c_673_n N_TE_B_M1024_g N_TE_B_c_648_n N_TE_B_c_675_n N_TE_B_M1026_g
+ N_TE_B_c_649_n N_TE_B_c_677_n N_TE_B_M1028_g N_TE_B_c_650_n N_TE_B_c_679_n
+ N_TE_B_M1030_g N_TE_B_c_651_n N_TE_B_c_652_n N_TE_B_c_682_n N_TE_B_M1002_g
+ N_TE_B_c_653_n N_TE_B_M1031_g N_TE_B_c_654_n N_TE_B_c_655_n N_TE_B_c_656_n
+ N_TE_B_c_657_n N_TE_B_c_658_n N_TE_B_c_659_n N_TE_B_c_660_n TE_B TE_B TE_B
+ N_TE_B_c_662_n N_TE_B_c_663_n PM_SKY130_FD_SC_HS__EBUFN_8%TE_B
x_PM_SKY130_FD_SC_HS__EBUFN_8%A N_A_c_831_n N_A_M1000_g N_A_c_827_n N_A_M1008_g
+ N_A_c_832_n N_A_M1007_g N_A_c_828_n N_A_M1018_g A N_A_c_830_n
+ PM_SKY130_FD_SC_HS__EBUFN_8%A
x_PM_SKY130_FD_SC_HS__EBUFN_8%A_28_368# N_A_28_368#_M1006_d N_A_28_368#_M1010_d
+ N_A_28_368#_M1014_d N_A_28_368#_M1017_d N_A_28_368#_M1020_d
+ N_A_28_368#_M1021_d N_A_28_368#_M1023_d N_A_28_368#_M1026_d
+ N_A_28_368#_M1030_d N_A_28_368#_c_877_n N_A_28_368#_c_878_n
+ N_A_28_368#_c_879_n N_A_28_368#_c_900_n N_A_28_368#_c_880_n
+ N_A_28_368#_c_904_n N_A_28_368#_c_881_n N_A_28_368#_c_966_p
+ N_A_28_368#_c_882_n N_A_28_368#_c_910_n N_A_28_368#_c_927_n
+ N_A_28_368#_c_912_n N_A_28_368#_c_913_n N_A_28_368#_c_914_n
+ N_A_28_368#_c_915_n N_A_28_368#_c_883_n N_A_28_368#_c_884_n
+ N_A_28_368#_c_885_n N_A_28_368#_c_886_n N_A_28_368#_c_887_n
+ N_A_28_368#_c_888_n N_A_28_368#_c_889_n PM_SKY130_FD_SC_HS__EBUFN_8%A_28_368#
x_PM_SKY130_FD_SC_HS__EBUFN_8%Z N_Z_M1005_s N_Z_M1011_s N_Z_M1032_s N_Z_M1034_s
+ N_Z_M1006_s N_Z_M1013_s N_Z_M1015_s N_Z_M1019_s N_Z_c_1030_n N_Z_c_1015_n
+ N_Z_c_1022_n N_Z_c_1041_n N_Z_c_1045_n N_Z_c_1016_n N_Z_c_1023_n N_Z_c_1055_n
+ N_Z_c_1059_n N_Z_c_1024_n N_Z_c_1017_n N_Z_c_1025_n N_Z_c_1075_n N_Z_c_1077_n
+ N_Z_c_1026_n N_Z_c_1018_n N_Z_c_1027_n N_Z_c_1028_n N_Z_c_1019_n Z Z Z
+ N_Z_c_1103_n Z PM_SKY130_FD_SC_HS__EBUFN_8%Z
x_PM_SKY130_FD_SC_HS__EBUFN_8%VPWR N_VPWR_M1016_s N_VPWR_M1022_s N_VPWR_M1024_s
+ N_VPWR_M1028_s N_VPWR_M1002_d N_VPWR_M1007_s N_VPWR_c_1149_n N_VPWR_c_1150_n
+ N_VPWR_c_1151_n N_VPWR_c_1152_n N_VPWR_c_1153_n N_VPWR_c_1154_n
+ N_VPWR_c_1155_n N_VPWR_c_1156_n VPWR N_VPWR_c_1157_n N_VPWR_c_1158_n
+ N_VPWR_c_1159_n N_VPWR_c_1160_n N_VPWR_c_1161_n N_VPWR_c_1162_n
+ N_VPWR_c_1163_n N_VPWR_c_1164_n N_VPWR_c_1165_n N_VPWR_c_1166_n
+ N_VPWR_c_1148_n PM_SKY130_FD_SC_HS__EBUFN_8%VPWR
x_PM_SKY130_FD_SC_HS__EBUFN_8%A_27_74# N_A_27_74#_M1005_d N_A_27_74#_M1009_d
+ N_A_27_74#_M1029_d N_A_27_74#_M1033_d N_A_27_74#_M1036_d N_A_27_74#_M1003_d
+ N_A_27_74#_M1012_d N_A_27_74#_M1027_d N_A_27_74#_M1037_d N_A_27_74#_c_1277_n
+ N_A_27_74#_c_1278_n N_A_27_74#_c_1279_n N_A_27_74#_c_1302_n
+ N_A_27_74#_c_1280_n N_A_27_74#_c_1305_n N_A_27_74#_c_1281_n
+ N_A_27_74#_c_1309_n N_A_27_74#_c_1282_n N_A_27_74#_c_1283_n
+ N_A_27_74#_c_1284_n N_A_27_74#_c_1285_n N_A_27_74#_c_1286_n
+ N_A_27_74#_c_1287_n N_A_27_74#_c_1288_n N_A_27_74#_c_1289_n
+ N_A_27_74#_c_1290_n N_A_27_74#_c_1291_n N_A_27_74#_c_1292_n
+ N_A_27_74#_c_1293_n N_A_27_74#_c_1294_n N_A_27_74#_c_1295_n
+ N_A_27_74#_c_1296_n N_A_27_74#_c_1297_n N_A_27_74#_c_1298_n
+ PM_SKY130_FD_SC_HS__EBUFN_8%A_27_74#
x_PM_SKY130_FD_SC_HS__EBUFN_8%VGND N_VGND_M1001_s N_VGND_M1004_s N_VGND_M1025_s
+ N_VGND_M1035_s N_VGND_M1031_d N_VGND_M1018_s N_VGND_c_1442_n N_VGND_c_1443_n
+ N_VGND_c_1444_n N_VGND_c_1445_n N_VGND_c_1446_n N_VGND_c_1447_n
+ N_VGND_c_1448_n N_VGND_c_1449_n N_VGND_c_1450_n N_VGND_c_1451_n
+ N_VGND_c_1452_n N_VGND_c_1453_n N_VGND_c_1454_n VGND N_VGND_c_1455_n
+ N_VGND_c_1456_n N_VGND_c_1457_n N_VGND_c_1458_n N_VGND_c_1459_n
+ N_VGND_c_1460_n PM_SKY130_FD_SC_HS__EBUFN_8%VGND
cc_1 VNB N_A_84_48#_M1005_g 0.02824f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_2 VNB N_A_84_48#_M1009_g 0.0212213f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=0.74
cc_3 VNB N_A_84_48#_M1011_g 0.0212477f $X=-0.19 $Y=-0.245 $X2=1.38 $Y2=0.74
cc_4 VNB N_A_84_48#_M1029_g 0.0218518f $X=-0.19 $Y=-0.245 $X2=1.81 $Y2=0.74
cc_5 VNB N_A_84_48#_M1032_g 0.0227695f $X=-0.19 $Y=-0.245 $X2=2.31 $Y2=0.74
cc_6 VNB N_A_84_48#_M1033_g 0.0229504f $X=-0.19 $Y=-0.245 $X2=2.81 $Y2=0.74
cc_7 VNB N_A_84_48#_M1034_g 0.0227562f $X=-0.19 $Y=-0.245 $X2=3.325 $Y2=0.74
cc_8 VNB N_A_84_48#_M1036_g 0.022169f $X=-0.19 $Y=-0.245 $X2=3.81 $Y2=0.74
cc_9 VNB N_A_84_48#_c_214_n 0.00906377f $X=-0.19 $Y=-0.245 $X2=3.87 $Y2=1.565
cc_10 VNB N_A_84_48#_c_215_n 0.00210925f $X=-0.19 $Y=-0.245 $X2=9.845 $Y2=0.505
cc_11 VNB N_A_84_48#_c_216_n 0.0247114f $X=-0.19 $Y=-0.245 $X2=10.23 $Y2=1.72
cc_12 VNB N_A_84_48#_c_217_n 0.233364f $X=-0.19 $Y=-0.245 $X2=3.795 $Y2=1.542
cc_13 VNB N_A_833_48#_c_478_n 0.0145547f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.32
cc_14 VNB N_A_833_48#_c_479_n 0.0127756f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_833_48#_c_480_n 0.00774194f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=1.765
cc_16 VNB N_A_833_48#_c_481_n 0.0143293f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=2.4
cc_17 VNB N_A_833_48#_c_482_n 0.0109932f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=0.74
cc_18 VNB N_A_833_48#_c_483_n 0.0149279f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_833_48#_c_484_n 0.0102563f $X=-0.19 $Y=-0.245 $X2=0.96 $Y2=2.4
cc_20 VNB N_A_833_48#_c_485_n 0.0149544f $X=-0.19 $Y=-0.245 $X2=1.38 $Y2=0.74
cc_21 VNB N_A_833_48#_c_486_n 0.0109799f $X=-0.19 $Y=-0.245 $X2=1.41 $Y2=1.765
cc_22 VNB N_A_833_48#_c_487_n 0.0145943f $X=-0.19 $Y=-0.245 $X2=1.41 $Y2=2.4
cc_23 VNB N_A_833_48#_c_488_n 0.0102563f $X=-0.19 $Y=-0.245 $X2=1.81 $Y2=0.74
cc_24 VNB N_A_833_48#_c_489_n 0.0149561f $X=-0.19 $Y=-0.245 $X2=1.91 $Y2=1.765
cc_25 VNB N_A_833_48#_c_490_n 0.0109799f $X=-0.19 $Y=-0.245 $X2=2.31 $Y2=1.32
cc_26 VNB N_A_833_48#_c_491_n 0.0145943f $X=-0.19 $Y=-0.245 $X2=2.31 $Y2=0.74
cc_27 VNB N_A_833_48#_c_492_n 0.0102563f $X=-0.19 $Y=-0.245 $X2=2.36 $Y2=2.4
cc_28 VNB N_A_833_48#_c_493_n 0.0183025f $X=-0.19 $Y=-0.245 $X2=2.81 $Y2=1.32
cc_29 VNB N_A_833_48#_c_494_n 0.0292022f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_833_48#_c_495_n 0.0299788f $X=-0.19 $Y=-0.245 $X2=2.81 $Y2=2.4
cc_31 VNB N_A_833_48#_c_496_n 0.00523367f $X=-0.19 $Y=-0.245 $X2=3.31 $Y2=1.765
cc_32 VNB N_A_833_48#_c_497_n 0.00436985f $X=-0.19 $Y=-0.245 $X2=3.31 $Y2=2.4
cc_33 VNB N_A_833_48#_c_498_n 0.00436985f $X=-0.19 $Y=-0.245 $X2=3.31 $Y2=2.4
cc_34 VNB N_A_833_48#_c_499_n 0.00438315f $X=-0.19 $Y=-0.245 $X2=3.325 $Y2=1.32
cc_35 VNB N_A_833_48#_c_500_n 0.00436985f $X=-0.19 $Y=-0.245 $X2=3.325 $Y2=0.74
cc_36 VNB N_A_833_48#_c_501_n 0.00438315f $X=-0.19 $Y=-0.245 $X2=3.325 $Y2=0.74
cc_37 VNB N_A_833_48#_c_502_n 0.00436985f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_833_48#_c_503_n 0.0152858f $X=-0.19 $Y=-0.245 $X2=3.795 $Y2=1.765
cc_39 VNB N_A_833_48#_c_504_n 0.020453f $X=-0.19 $Y=-0.245 $X2=3.795 $Y2=2.4
cc_40 VNB N_A_833_48#_c_505_n 0.0111351f $X=-0.19 $Y=-0.245 $X2=3.81 $Y2=1.32
cc_41 VNB N_A_833_48#_c_506_n 0.0795427f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_833_48#_c_507_n 0.0141642f $X=-0.19 $Y=-0.245 $X2=1.14 $Y2=1.485
cc_43 VNB N_TE_B_c_643_n 0.00960637f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_TE_B_c_644_n 0.00495511f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_TE_B_c_645_n 0.00718581f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_46 VNB N_TE_B_c_646_n 0.00957048f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=1.32
cc_47 VNB N_TE_B_c_647_n 0.00720484f $X=-0.19 $Y=-0.245 $X2=0.96 $Y2=2.4
cc_48 VNB N_TE_B_c_648_n 0.0095704f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_TE_B_c_649_n 0.00720484f $X=-0.19 $Y=-0.245 $X2=1.81 $Y2=0.74
cc_50 VNB N_TE_B_c_650_n 0.0113005f $X=-0.19 $Y=-0.245 $X2=1.91 $Y2=2.4
cc_51 VNB N_TE_B_c_651_n 0.035544f $X=-0.19 $Y=-0.245 $X2=2.36 $Y2=2.4
cc_52 VNB N_TE_B_c_652_n 0.0283125f $X=-0.19 $Y=-0.245 $X2=2.81 $Y2=1.32
cc_53 VNB N_TE_B_c_653_n 0.0227572f $X=-0.19 $Y=-0.245 $X2=2.81 $Y2=1.765
cc_54 VNB N_TE_B_c_654_n 0.003679f $X=-0.19 $Y=-0.245 $X2=3.31 $Y2=1.765
cc_55 VNB N_TE_B_c_655_n 0.00367913f $X=-0.19 $Y=-0.245 $X2=3.31 $Y2=2.4
cc_56 VNB N_TE_B_c_656_n 0.00367905f $X=-0.19 $Y=-0.245 $X2=3.31 $Y2=2.4
cc_57 VNB N_TE_B_c_657_n 0.00367913f $X=-0.19 $Y=-0.245 $X2=3.325 $Y2=1.32
cc_58 VNB N_TE_B_c_658_n 0.00367913f $X=-0.19 $Y=-0.245 $X2=3.325 $Y2=0.74
cc_59 VNB N_TE_B_c_659_n 0.0036791f $X=-0.19 $Y=-0.245 $X2=3.325 $Y2=0.74
cc_60 VNB N_TE_B_c_660_n 0.00594258f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB TE_B 0.0193491f $X=-0.19 $Y=-0.245 $X2=3.795 $Y2=2.4
cc_62 VNB N_TE_B_c_662_n 0.0105317f $X=-0.19 $Y=-0.245 $X2=1.14 $Y2=1.485
cc_63 VNB N_TE_B_c_663_n 0.022361f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_A_c_827_n 0.0172452f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_A_c_828_n 0.0188503f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB A 0.0035636f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=2.4
cc_67 VNB N_A_c_830_n 0.0565653f $X=-0.19 $Y=-0.245 $X2=0.96 $Y2=2.4
cc_68 VNB N_Z_c_1015_n 0.00261517f $X=-0.19 $Y=-0.245 $X2=1.81 $Y2=0.74
cc_69 VNB N_Z_c_1016_n 0.00307912f $X=-0.19 $Y=-0.245 $X2=2.36 $Y2=2.4
cc_70 VNB N_Z_c_1017_n 0.00559895f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_Z_c_1018_n 0.00229628f $X=-0.19 $Y=-0.245 $X2=3.87 $Y2=1.565
cc_72 VNB N_Z_c_1019_n 0.00229411f $X=-0.19 $Y=-0.245 $X2=4.04 $Y2=2.135
cc_73 VNB Z 2.27624e-19 $X=-0.19 $Y=-0.245 $X2=9.805 $Y2=1.89
cc_74 VNB Z 0.00172469f $X=-0.19 $Y=-0.245 $X2=9.805 $Y2=2.22
cc_75 VNB N_VPWR_c_1148_n 0.442315f $X=-0.19 $Y=-0.245 $X2=3.655 $Y2=1.485
cc_76 VNB N_A_27_74#_c_1277_n 0.0362361f $X=-0.19 $Y=-0.245 $X2=1.81 $Y2=0.74
cc_77 VNB N_A_27_74#_c_1278_n 0.0027626f $X=-0.19 $Y=-0.245 $X2=1.91 $Y2=1.765
cc_78 VNB N_A_27_74#_c_1279_n 0.00931596f $X=-0.19 $Y=-0.245 $X2=1.91 $Y2=2.4
cc_79 VNB N_A_27_74#_c_1280_n 0.0028694f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_A_27_74#_c_1281_n 0.00280532f $X=-0.19 $Y=-0.245 $X2=2.81 $Y2=0.74
cc_81 VNB N_A_27_74#_c_1282_n 0.00488489f $X=-0.19 $Y=-0.245 $X2=3.31 $Y2=2.4
cc_82 VNB N_A_27_74#_c_1283_n 4.66026e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_83 VNB N_A_27_74#_c_1284_n 0.00627739f $X=-0.19 $Y=-0.245 $X2=3.795 $Y2=1.765
cc_84 VNB N_A_27_74#_c_1285_n 0.00583076f $X=-0.19 $Y=-0.245 $X2=3.795 $Y2=2.4
cc_85 VNB N_A_27_74#_c_1286_n 0.0023333f $X=-0.19 $Y=-0.245 $X2=3.81 $Y2=0.74
cc_86 VNB N_A_27_74#_c_1287_n 0.00528215f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_87 VNB N_A_27_74#_c_1288_n 0.00263046f $X=-0.19 $Y=-0.245 $X2=1.14 $Y2=1.485
cc_88 VNB N_A_27_74#_c_1289_n 0.00563126f $X=-0.19 $Y=-0.245 $X2=3.87 $Y2=1.565
cc_89 VNB N_A_27_74#_c_1290_n 0.00263046f $X=-0.19 $Y=-0.245 $X2=7.585 $Y2=2.135
cc_90 VNB N_A_27_74#_c_1291_n 0.00976772f $X=-0.19 $Y=-0.245 $X2=9.665 $Y2=2.305
cc_91 VNB N_A_27_74#_c_1292_n 0.00266546f $X=-0.19 $Y=-0.245 $X2=9.805 $Y2=1.985
cc_92 VNB N_A_27_74#_c_1293_n 0.00121874f $X=-0.19 $Y=-0.245 $X2=9.805 $Y2=2.39
cc_93 VNB N_A_27_74#_c_1294_n 0.00220535f $X=-0.19 $Y=-0.245 $X2=9.805 $Y2=2.815
cc_94 VNB N_A_27_74#_c_1295_n 0.00233543f $X=-0.19 $Y=-0.245 $X2=9.83 $Y2=2.815
cc_95 VNB N_A_27_74#_c_1296_n 0.0105845f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_96 VNB N_A_27_74#_c_1297_n 0.00238685f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_97 VNB N_A_27_74#_c_1298_n 0.00238685f $X=-0.19 $Y=-0.245 $X2=10.145
+ $Y2=0.925
cc_98 VNB N_VGND_c_1442_n 0.00334323f $X=-0.19 $Y=-0.245 $X2=1.38 $Y2=1.32
cc_99 VNB N_VGND_c_1443_n 0.00789915f $X=-0.19 $Y=-0.245 $X2=1.41 $Y2=1.765
cc_100 VNB N_VGND_c_1444_n 0.00582552f $X=-0.19 $Y=-0.245 $X2=1.81 $Y2=0.74
cc_101 VNB N_VGND_c_1445_n 0.00659784f $X=-0.19 $Y=-0.245 $X2=1.91 $Y2=2.4
cc_102 VNB N_VGND_c_1446_n 0.00719205f $X=-0.19 $Y=-0.245 $X2=2.31 $Y2=0.74
cc_103 VNB N_VGND_c_1447_n 0.0120978f $X=-0.19 $Y=-0.245 $X2=2.36 $Y2=1.765
cc_104 VNB N_VGND_c_1448_n 0.0189538f $X=-0.19 $Y=-0.245 $X2=2.36 $Y2=2.4
cc_105 VNB N_VGND_c_1449_n 0.0998102f $X=-0.19 $Y=-0.245 $X2=2.81 $Y2=0.74
cc_106 VNB N_VGND_c_1450_n 0.00604233f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_107 VNB N_VGND_c_1451_n 0.0172524f $X=-0.19 $Y=-0.245 $X2=2.81 $Y2=2.4
cc_108 VNB N_VGND_c_1452_n 0.00326991f $X=-0.19 $Y=-0.245 $X2=2.81 $Y2=2.4
cc_109 VNB N_VGND_c_1453_n 0.0172524f $X=-0.19 $Y=-0.245 $X2=3.31 $Y2=2.4
cc_110 VNB N_VGND_c_1454_n 0.00461913f $X=-0.19 $Y=-0.245 $X2=3.31 $Y2=2.4
cc_111 VNB N_VGND_c_1455_n 0.0172524f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_112 VNB N_VGND_c_1456_n 0.0569499f $X=-0.19 $Y=-0.245 $X2=3.955 $Y2=2.05
cc_113 VNB N_VGND_c_1457_n 0.0172141f $X=-0.19 $Y=-0.245 $X2=9.805 $Y2=1.89
cc_114 VNB N_VGND_c_1458_n 0.00461913f $X=-0.19 $Y=-0.245 $X2=9.83 $Y2=2.815
cc_115 VNB N_VGND_c_1459_n 0.00326991f $X=-0.19 $Y=-0.245 $X2=9.805 $Y2=0.505
cc_116 VNB N_VGND_c_1460_n 0.558924f $X=-0.19 $Y=-0.245 $X2=9.93 $Y2=0.925
cc_117 VPB N_A_84_48#_c_218_n 0.0181039f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=1.765
cc_118 VPB N_A_84_48#_c_219_n 0.0145458f $X=-0.19 $Y=1.66 $X2=0.96 $Y2=1.765
cc_119 VPB N_A_84_48#_c_220_n 0.0149261f $X=-0.19 $Y=1.66 $X2=1.41 $Y2=1.765
cc_120 VPB N_A_84_48#_c_221_n 0.0149468f $X=-0.19 $Y=1.66 $X2=1.91 $Y2=1.765
cc_121 VPB N_A_84_48#_c_222_n 0.0145655f $X=-0.19 $Y=1.66 $X2=2.36 $Y2=1.765
cc_122 VPB N_A_84_48#_c_223_n 0.0149469f $X=-0.19 $Y=1.66 $X2=2.81 $Y2=1.765
cc_123 VPB N_A_84_48#_c_224_n 0.0152144f $X=-0.19 $Y=1.66 $X2=3.31 $Y2=1.765
cc_124 VPB N_A_84_48#_c_225_n 0.015225f $X=-0.19 $Y=1.66 $X2=3.795 $Y2=1.765
cc_125 VPB N_A_84_48#_c_226_n 0.00229687f $X=-0.19 $Y=1.66 $X2=3.955 $Y2=2.05
cc_126 VPB N_A_84_48#_c_227_n 0.0123659f $X=-0.19 $Y=1.66 $X2=9.665 $Y2=2.305
cc_127 VPB N_A_84_48#_c_228_n 0.00243101f $X=-0.19 $Y=1.66 $X2=9.83 $Y2=2.815
cc_128 VPB N_A_84_48#_c_229_n 0.00503473f $X=-0.19 $Y=1.66 $X2=10.145 $Y2=1.805
cc_129 VPB N_A_84_48#_c_230_n 0.00205111f $X=-0.19 $Y=1.66 $X2=9.945 $Y2=1.805
cc_130 VPB N_A_84_48#_c_216_n 0.00255885f $X=-0.19 $Y=1.66 $X2=10.23 $Y2=1.72
cc_131 VPB N_A_84_48#_c_217_n 0.0552073f $X=-0.19 $Y=1.66 $X2=3.795 $Y2=1.542
cc_132 VPB N_A_833_48#_c_504_n 0.00116802f $X=-0.19 $Y=1.66 $X2=3.795 $Y2=2.4
cc_133 VPB N_A_833_48#_c_509_n 0.012324f $X=-0.19 $Y=1.66 $X2=3.87 $Y2=1.565
cc_134 VPB N_TE_B_c_664_n 0.0161921f $X=-0.19 $Y=1.66 $X2=9.705 $Y2=0.37
cc_135 VPB N_TE_B_c_643_n 0.00973153f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_136 VPB N_TE_B_c_644_n 0.00429227f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_137 VPB N_TE_B_c_667_n 0.0163477f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_138 VPB N_TE_B_c_645_n 0.00620972f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.74
cc_139 VPB N_TE_B_c_669_n 0.0163499f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=1.765
cc_140 VPB N_TE_B_c_646_n 0.00973153f $X=-0.19 $Y=1.66 $X2=0.925 $Y2=1.32
cc_141 VPB N_TE_B_c_671_n 0.0163499f $X=-0.19 $Y=1.66 $X2=0.925 $Y2=0.74
cc_142 VPB N_TE_B_c_647_n 0.00620972f $X=-0.19 $Y=1.66 $X2=0.96 $Y2=2.4
cc_143 VPB N_TE_B_c_673_n 0.0163499f $X=-0.19 $Y=1.66 $X2=1.38 $Y2=1.32
cc_144 VPB N_TE_B_c_648_n 0.00973153f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_145 VPB N_TE_B_c_675_n 0.016351f $X=-0.19 $Y=1.66 $X2=1.41 $Y2=2.4
cc_146 VPB N_TE_B_c_649_n 0.00620972f $X=-0.19 $Y=1.66 $X2=1.81 $Y2=0.74
cc_147 VPB N_TE_B_c_677_n 0.016792f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_148 VPB N_TE_B_c_650_n 0.0121704f $X=-0.19 $Y=1.66 $X2=1.91 $Y2=2.4
cc_149 VPB N_TE_B_c_679_n 0.0209085f $X=-0.19 $Y=1.66 $X2=2.31 $Y2=0.74
cc_150 VPB N_TE_B_c_651_n 0.0151939f $X=-0.19 $Y=1.66 $X2=2.36 $Y2=2.4
cc_151 VPB N_TE_B_c_652_n 0.00960941f $X=-0.19 $Y=1.66 $X2=2.81 $Y2=1.32
cc_152 VPB N_TE_B_c_682_n 0.0206913f $X=-0.19 $Y=1.66 $X2=2.81 $Y2=0.74
cc_153 VPB N_TE_B_c_654_n 0.00167153f $X=-0.19 $Y=1.66 $X2=3.31 $Y2=1.765
cc_154 VPB N_TE_B_c_655_n 0.00167153f $X=-0.19 $Y=1.66 $X2=3.31 $Y2=2.4
cc_155 VPB N_TE_B_c_656_n 0.00167153f $X=-0.19 $Y=1.66 $X2=3.31 $Y2=2.4
cc_156 VPB N_TE_B_c_657_n 0.00167153f $X=-0.19 $Y=1.66 $X2=3.325 $Y2=1.32
cc_157 VPB N_TE_B_c_658_n 0.00167153f $X=-0.19 $Y=1.66 $X2=3.325 $Y2=0.74
cc_158 VPB N_TE_B_c_659_n 0.00167153f $X=-0.19 $Y=1.66 $X2=3.325 $Y2=0.74
cc_159 VPB N_TE_B_c_660_n 0.00167153f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_160 VPB N_TE_B_c_662_n 0.00841803f $X=-0.19 $Y=1.66 $X2=1.14 $Y2=1.485
cc_161 VPB N_TE_B_c_663_n 0.00458689f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_162 VPB N_A_c_831_n 0.0159625f $X=-0.19 $Y=1.66 $X2=9.705 $Y2=0.37
cc_163 VPB N_A_c_832_n 0.0173807f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.32
cc_164 VPB N_A_c_830_n 0.0136734f $X=-0.19 $Y=1.66 $X2=0.96 $Y2=2.4
cc_165 VPB N_A_28_368#_c_877_n 0.0501935f $X=-0.19 $Y=1.66 $X2=1.81 $Y2=0.74
cc_166 VPB N_A_28_368#_c_878_n 0.0029406f $X=-0.19 $Y=1.66 $X2=1.91 $Y2=2.4
cc_167 VPB N_A_28_368#_c_879_n 0.00935849f $X=-0.19 $Y=1.66 $X2=2.31 $Y2=1.32
cc_168 VPB N_A_28_368#_c_880_n 0.00294772f $X=-0.19 $Y=1.66 $X2=2.36 $Y2=2.4
cc_169 VPB N_A_28_368#_c_881_n 0.0028338f $X=-0.19 $Y=1.66 $X2=2.81 $Y2=1.765
cc_170 VPB N_A_28_368#_c_882_n 0.0049919f $X=-0.19 $Y=1.66 $X2=3.325 $Y2=1.32
cc_171 VPB N_A_28_368#_c_883_n 0.00181992f $X=-0.19 $Y=1.66 $X2=3.87 $Y2=1.565
cc_172 VPB N_A_28_368#_c_884_n 0.00123754f $X=-0.19 $Y=1.66 $X2=3.655 $Y2=1.565
cc_173 VPB N_A_28_368#_c_885_n 0.00196551f $X=-0.19 $Y=1.66 $X2=3.955 $Y2=1.65
cc_174 VPB N_A_28_368#_c_886_n 0.00256678f $X=-0.19 $Y=1.66 $X2=9.665 $Y2=2.305
cc_175 VPB N_A_28_368#_c_887_n 0.00256678f $X=-0.19 $Y=1.66 $X2=9.805 $Y2=1.89
cc_176 VPB N_A_28_368#_c_888_n 0.00256678f $X=-0.19 $Y=1.66 $X2=9.83 $Y2=1.985
cc_177 VPB N_A_28_368#_c_889_n 0.0188798f $X=-0.19 $Y=1.66 $X2=9.83 $Y2=2.815
cc_178 VPB N_Z_c_1022_n 0.00199674f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_179 VPB N_Z_c_1023_n 0.00179576f $X=-0.19 $Y=1.66 $X2=2.81 $Y2=0.74
cc_180 VPB N_Z_c_1024_n 0.00209616f $X=-0.19 $Y=1.66 $X2=3.325 $Y2=0.74
cc_181 VPB N_Z_c_1025_n 0.00209284f $X=-0.19 $Y=1.66 $X2=3.795 $Y2=2.4
cc_182 VPB N_Z_c_1026_n 4.41918e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_183 VPB N_Z_c_1027_n 0.00193069f $X=-0.19 $Y=1.66 $X2=3.955 $Y2=1.65
cc_184 VPB N_Z_c_1028_n 0.00183525f $X=-0.19 $Y=1.66 $X2=7.585 $Y2=2.135
cc_185 VPB Z 0.00153702f $X=-0.19 $Y=1.66 $X2=9.805 $Y2=2.22
cc_186 VPB N_VPWR_c_1149_n 0.0085833f $X=-0.19 $Y=1.66 $X2=1.38 $Y2=1.32
cc_187 VPB N_VPWR_c_1150_n 0.00830446f $X=-0.19 $Y=1.66 $X2=1.41 $Y2=1.765
cc_188 VPB N_VPWR_c_1151_n 0.00900305f $X=-0.19 $Y=1.66 $X2=1.81 $Y2=0.74
cc_189 VPB N_VPWR_c_1152_n 0.0188241f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_190 VPB N_VPWR_c_1153_n 0.00804215f $X=-0.19 $Y=1.66 $X2=2.31 $Y2=1.32
cc_191 VPB N_VPWR_c_1154_n 0.00572483f $X=-0.19 $Y=1.66 $X2=2.36 $Y2=1.765
cc_192 VPB N_VPWR_c_1155_n 0.0120106f $X=-0.19 $Y=1.66 $X2=2.36 $Y2=2.4
cc_193 VPB N_VPWR_c_1156_n 0.0444341f $X=-0.19 $Y=1.66 $X2=2.81 $Y2=0.74
cc_194 VPB N_VPWR_c_1157_n 0.101629f $X=-0.19 $Y=1.66 $X2=3.31 $Y2=1.765
cc_195 VPB N_VPWR_c_1158_n 0.0186948f $X=-0.19 $Y=1.66 $X2=3.795 $Y2=2.4
cc_196 VPB N_VPWR_c_1159_n 0.0186948f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_197 VPB N_VPWR_c_1160_n 0.0417371f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_198 VPB N_VPWR_c_1161_n 0.0173363f $X=-0.19 $Y=1.66 $X2=7.755 $Y2=2.305
cc_199 VPB N_VPWR_c_1162_n 0.00631813f $X=-0.19 $Y=1.66 $X2=9.805 $Y2=2.815
cc_200 VPB N_VPWR_c_1163_n 0.00632182f $X=-0.19 $Y=1.66 $X2=9.805 $Y2=0.84
cc_201 VPB N_VPWR_c_1164_n 0.00632182f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_202 VPB N_VPWR_c_1165_n 0.00631222f $X=-0.19 $Y=1.66 $X2=10.145 $Y2=1.805
cc_203 VPB N_VPWR_c_1166_n 0.00614127f $X=-0.19 $Y=1.66 $X2=10.23 $Y2=1.72
cc_204 VPB N_VPWR_c_1148_n 0.115984f $X=-0.19 $Y=1.66 $X2=3.655 $Y2=1.485
cc_205 N_A_84_48#_c_227_n N_A_833_48#_M1002_s 0.0246237f $X=9.665 $Y=2.305 $X2=0
+ $Y2=0
cc_206 N_A_84_48#_M1036_g N_A_833_48#_c_478_n 0.00835898f $X=3.81 $Y=0.74 $X2=0
+ $Y2=0
cc_207 N_A_84_48#_c_217_n N_A_833_48#_c_480_n 0.00835898f $X=3.795 $Y=1.542
+ $X2=0 $Y2=0
cc_208 N_A_84_48#_c_227_n N_A_833_48#_c_513_n 0.00899589f $X=9.665 $Y=2.305
+ $X2=0 $Y2=0
cc_209 N_A_84_48#_c_227_n N_A_833_48#_c_509_n 0.0674273f $X=9.665 $Y=2.305 $X2=0
+ $Y2=0
cc_210 N_A_84_48#_c_238_p N_A_833_48#_c_509_n 0.00425949f $X=9.83 $Y=1.985 $X2=0
+ $Y2=0
cc_211 N_A_84_48#_c_230_n N_A_833_48#_c_509_n 0.00254884f $X=9.945 $Y=1.805
+ $X2=0 $Y2=0
cc_212 N_A_84_48#_c_225_n N_TE_B_c_664_n 0.0225535f $X=3.795 $Y=1.765 $X2=-0.19
+ $Y2=-0.245
cc_213 N_A_84_48#_c_226_n N_TE_B_c_664_n 0.00616529f $X=3.955 $Y=2.05 $X2=-0.19
+ $Y2=-0.245
cc_214 N_A_84_48#_c_242_p N_TE_B_c_664_n 0.0154121f $X=7.585 $Y=2.135 $X2=-0.19
+ $Y2=-0.245
cc_215 N_A_84_48#_c_242_p N_TE_B_c_643_n 0.00666012f $X=7.585 $Y=2.135 $X2=0
+ $Y2=0
cc_216 N_A_84_48#_c_214_n N_TE_B_c_644_n 0.00106842f $X=3.87 $Y=1.565 $X2=0
+ $Y2=0
cc_217 N_A_84_48#_c_226_n N_TE_B_c_644_n 0.00266816f $X=3.955 $Y=2.05 $X2=0
+ $Y2=0
cc_218 N_A_84_48#_c_217_n N_TE_B_c_644_n 0.00662396f $X=3.795 $Y=1.542 $X2=0
+ $Y2=0
cc_219 N_A_84_48#_c_242_p N_TE_B_c_667_n 0.012726f $X=7.585 $Y=2.135 $X2=0 $Y2=0
cc_220 N_A_84_48#_c_242_p N_TE_B_c_645_n 0.0024232f $X=7.585 $Y=2.135 $X2=0
+ $Y2=0
cc_221 N_A_84_48#_c_242_p N_TE_B_c_669_n 0.012729f $X=7.585 $Y=2.135 $X2=0 $Y2=0
cc_222 N_A_84_48#_c_242_p N_TE_B_c_646_n 0.00442441f $X=7.585 $Y=2.135 $X2=0
+ $Y2=0
cc_223 N_A_84_48#_c_242_p N_TE_B_c_671_n 0.0127271f $X=7.585 $Y=2.135 $X2=0
+ $Y2=0
cc_224 N_A_84_48#_c_242_p N_TE_B_c_647_n 0.00241357f $X=7.585 $Y=2.135 $X2=0
+ $Y2=0
cc_225 N_A_84_48#_c_242_p N_TE_B_c_673_n 0.012729f $X=7.585 $Y=2.135 $X2=0 $Y2=0
cc_226 N_A_84_48#_c_242_p N_TE_B_c_648_n 0.00442341f $X=7.585 $Y=2.135 $X2=0
+ $Y2=0
cc_227 N_A_84_48#_c_242_p N_TE_B_c_675_n 0.0126642f $X=7.585 $Y=2.135 $X2=0
+ $Y2=0
cc_228 N_A_84_48#_c_242_p N_TE_B_c_649_n 0.00241357f $X=7.585 $Y=2.135 $X2=0
+ $Y2=0
cc_229 N_A_84_48#_c_242_p N_TE_B_c_677_n 0.0131455f $X=7.585 $Y=2.135 $X2=0
+ $Y2=0
cc_230 N_A_84_48#_c_258_p N_TE_B_c_677_n 0.0036836f $X=7.67 $Y=2.135 $X2=0 $Y2=0
cc_231 N_A_84_48#_c_242_p N_TE_B_c_650_n 0.0035728f $X=7.585 $Y=2.135 $X2=0
+ $Y2=0
cc_232 N_A_84_48#_c_258_p N_TE_B_c_650_n 0.00425484f $X=7.67 $Y=2.135 $X2=0
+ $Y2=0
cc_233 N_A_84_48#_c_227_n N_TE_B_c_679_n 0.0153437f $X=9.665 $Y=2.305 $X2=0
+ $Y2=0
cc_234 N_A_84_48#_c_227_n N_TE_B_c_682_n 0.0190695f $X=9.665 $Y=2.305 $X2=0
+ $Y2=0
cc_235 N_A_84_48#_c_238_p N_TE_B_c_682_n 0.00127549f $X=9.83 $Y=1.985 $X2=0
+ $Y2=0
cc_236 N_A_84_48#_c_228_n N_TE_B_c_682_n 8.34609e-19 $X=9.83 $Y=2.815 $X2=0
+ $Y2=0
cc_237 N_A_84_48#_c_230_n N_TE_B_c_682_n 4.30703e-19 $X=9.945 $Y=1.805 $X2=0
+ $Y2=0
cc_238 N_A_84_48#_c_227_n TE_B 0.0105454f $X=9.665 $Y=2.305 $X2=0 $Y2=0
cc_239 N_A_84_48#_c_227_n N_TE_B_c_662_n 0.00128972f $X=9.665 $Y=2.305 $X2=0
+ $Y2=0
cc_240 N_A_84_48#_c_227_n N_TE_B_c_663_n 0.00127253f $X=9.665 $Y=2.305 $X2=0
+ $Y2=0
cc_241 N_A_84_48#_c_230_n N_TE_B_c_663_n 2.47064e-19 $X=9.945 $Y=1.805 $X2=0
+ $Y2=0
cc_242 N_A_84_48#_c_227_n N_A_c_831_n 0.0160358f $X=9.665 $Y=2.305 $X2=-0.19
+ $Y2=-0.245
cc_243 N_A_84_48#_c_238_p N_A_c_831_n 0.00628912f $X=9.83 $Y=1.985 $X2=-0.19
+ $Y2=-0.245
cc_244 N_A_84_48#_c_228_n N_A_c_831_n 0.00767841f $X=9.83 $Y=2.815 $X2=-0.19
+ $Y2=-0.245
cc_245 N_A_84_48#_c_230_n N_A_c_831_n 0.0032668f $X=9.945 $Y=1.805 $X2=-0.19
+ $Y2=-0.245
cc_246 N_A_84_48#_c_274_p N_A_c_831_n 2.24111e-19 $X=9.805 $Y=2.305 $X2=-0.19
+ $Y2=-0.245
cc_247 N_A_84_48#_c_275_p N_A_c_827_n 0.00208866f $X=9.805 $Y=0.84 $X2=0 $Y2=0
cc_248 N_A_84_48#_c_215_n N_A_c_827_n 0.00591333f $X=9.845 $Y=0.505 $X2=0 $Y2=0
cc_249 N_A_84_48#_c_228_n N_A_c_832_n 2.71519e-19 $X=9.83 $Y=2.815 $X2=0 $Y2=0
cc_250 N_A_84_48#_c_229_n N_A_c_832_n 0.0110436f $X=10.145 $Y=1.805 $X2=0 $Y2=0
cc_251 N_A_84_48#_c_215_n N_A_c_828_n 3.45303e-19 $X=9.845 $Y=0.505 $X2=0 $Y2=0
cc_252 N_A_84_48#_c_280_p N_A_c_828_n 0.0152487f $X=10.145 $Y=0.925 $X2=0 $Y2=0
cc_253 N_A_84_48#_c_216_n N_A_c_828_n 0.0057552f $X=10.23 $Y=1.72 $X2=0 $Y2=0
cc_254 N_A_84_48#_c_227_n A 4.25182e-19 $X=9.665 $Y=2.305 $X2=0 $Y2=0
cc_255 N_A_84_48#_c_275_p A 0.0190643f $X=9.805 $Y=0.84 $X2=0 $Y2=0
cc_256 N_A_84_48#_c_229_n A 0.00213835f $X=10.145 $Y=1.805 $X2=0 $Y2=0
cc_257 N_A_84_48#_c_230_n A 0.023783f $X=9.945 $Y=1.805 $X2=0 $Y2=0
cc_258 N_A_84_48#_c_216_n A 0.0279669f $X=10.23 $Y=1.72 $X2=0 $Y2=0
cc_259 N_A_84_48#_c_275_p N_A_c_830_n 7.03839e-19 $X=9.805 $Y=0.84 $X2=0 $Y2=0
cc_260 N_A_84_48#_c_229_n N_A_c_830_n 0.01014f $X=10.145 $Y=1.805 $X2=0 $Y2=0
cc_261 N_A_84_48#_c_230_n N_A_c_830_n 0.00299627f $X=9.945 $Y=1.805 $X2=0 $Y2=0
cc_262 N_A_84_48#_c_216_n N_A_c_830_n 0.0174888f $X=10.23 $Y=1.72 $X2=0 $Y2=0
cc_263 N_A_84_48#_c_226_n N_A_28_368#_M1020_d 0.00283534f $X=3.955 $Y=2.05 $X2=0
+ $Y2=0
cc_264 N_A_84_48#_c_242_p N_A_28_368#_M1020_d 0.00424436f $X=7.585 $Y=2.135
+ $X2=0 $Y2=0
cc_265 N_A_84_48#_c_293_p N_A_28_368#_M1020_d 0.00197336f $X=4.04 $Y=2.135 $X2=0
+ $Y2=0
cc_266 N_A_84_48#_c_242_p N_A_28_368#_M1021_d 0.00501812f $X=7.585 $Y=2.135
+ $X2=0 $Y2=0
cc_267 N_A_84_48#_c_242_p N_A_28_368#_M1023_d 0.00503421f $X=7.585 $Y=2.135
+ $X2=0 $Y2=0
cc_268 N_A_84_48#_c_242_p N_A_28_368#_M1026_d 0.00503421f $X=7.585 $Y=2.135
+ $X2=0 $Y2=0
cc_269 N_A_84_48#_c_227_n N_A_28_368#_M1030_d 0.00585261f $X=9.665 $Y=2.305
+ $X2=0 $Y2=0
cc_270 N_A_84_48#_c_218_n N_A_28_368#_c_877_n 0.00770803f $X=0.51 $Y=1.765 $X2=0
+ $Y2=0
cc_271 N_A_84_48#_c_218_n N_A_28_368#_c_878_n 0.01294f $X=0.51 $Y=1.765 $X2=0
+ $Y2=0
cc_272 N_A_84_48#_c_219_n N_A_28_368#_c_878_n 0.0128349f $X=0.96 $Y=1.765 $X2=0
+ $Y2=0
cc_273 N_A_84_48#_c_220_n N_A_28_368#_c_900_n 0.00974071f $X=1.41 $Y=1.765 $X2=0
+ $Y2=0
cc_274 N_A_84_48#_c_221_n N_A_28_368#_c_900_n 5.35939e-19 $X=1.91 $Y=1.765 $X2=0
+ $Y2=0
cc_275 N_A_84_48#_c_220_n N_A_28_368#_c_880_n 0.0111147f $X=1.41 $Y=1.765 $X2=0
+ $Y2=0
cc_276 N_A_84_48#_c_221_n N_A_28_368#_c_880_n 0.0131082f $X=1.91 $Y=1.765 $X2=0
+ $Y2=0
cc_277 N_A_84_48#_c_221_n N_A_28_368#_c_904_n 0.00553744f $X=1.91 $Y=1.765 $X2=0
+ $Y2=0
cc_278 N_A_84_48#_c_222_n N_A_28_368#_c_904_n 0.00553744f $X=2.36 $Y=1.765 $X2=0
+ $Y2=0
cc_279 N_A_84_48#_c_222_n N_A_28_368#_c_881_n 0.0128349f $X=2.36 $Y=1.765 $X2=0
+ $Y2=0
cc_280 N_A_84_48#_c_223_n N_A_28_368#_c_881_n 0.0138537f $X=2.81 $Y=1.765 $X2=0
+ $Y2=0
cc_281 N_A_84_48#_c_224_n N_A_28_368#_c_882_n 0.0132138f $X=3.31 $Y=1.765 $X2=0
+ $Y2=0
cc_282 N_A_84_48#_c_225_n N_A_28_368#_c_882_n 0.0134638f $X=3.795 $Y=1.765 $X2=0
+ $Y2=0
cc_283 N_A_84_48#_c_242_p N_A_28_368#_c_910_n 0.00822853f $X=7.585 $Y=2.135
+ $X2=0 $Y2=0
cc_284 N_A_84_48#_c_293_p N_A_28_368#_c_910_n 0.0101487f $X=4.04 $Y=2.135 $X2=0
+ $Y2=0
cc_285 N_A_84_48#_c_242_p N_A_28_368#_c_912_n 0.039006f $X=7.585 $Y=2.135 $X2=0
+ $Y2=0
cc_286 N_A_84_48#_c_242_p N_A_28_368#_c_913_n 0.039006f $X=7.585 $Y=2.135 $X2=0
+ $Y2=0
cc_287 N_A_84_48#_c_242_p N_A_28_368#_c_914_n 0.0390399f $X=7.585 $Y=2.135 $X2=0
+ $Y2=0
cc_288 N_A_84_48#_c_242_p N_A_28_368#_c_915_n 0.0136727f $X=7.585 $Y=2.135 $X2=0
+ $Y2=0
cc_289 N_A_84_48#_c_227_n N_A_28_368#_c_915_n 0.00915035f $X=9.665 $Y=2.305
+ $X2=0 $Y2=0
cc_290 N_A_84_48#_c_258_p N_A_28_368#_c_915_n 0.0124697f $X=7.67 $Y=2.135 $X2=0
+ $Y2=0
cc_291 N_A_84_48#_c_220_n N_A_28_368#_c_883_n 0.00175197f $X=1.41 $Y=1.765 $X2=0
+ $Y2=0
cc_292 N_A_84_48#_c_242_p N_A_28_368#_c_886_n 0.0171364f $X=7.585 $Y=2.135 $X2=0
+ $Y2=0
cc_293 N_A_84_48#_c_242_p N_A_28_368#_c_887_n 0.0171364f $X=7.585 $Y=2.135 $X2=0
+ $Y2=0
cc_294 N_A_84_48#_c_242_p N_A_28_368#_c_888_n 0.016984f $X=7.585 $Y=2.135 $X2=0
+ $Y2=0
cc_295 N_A_84_48#_c_227_n N_A_28_368#_c_889_n 0.0211942f $X=9.665 $Y=2.305 $X2=0
+ $Y2=0
cc_296 N_A_84_48#_c_218_n N_Z_c_1030_n 0.00932452f $X=0.51 $Y=1.765 $X2=0 $Y2=0
cc_297 N_A_84_48#_c_219_n N_Z_c_1030_n 0.00890996f $X=0.96 $Y=1.765 $X2=0 $Y2=0
cc_298 N_A_84_48#_c_220_n N_Z_c_1030_n 6.51855e-19 $X=1.41 $Y=1.765 $X2=0 $Y2=0
cc_299 N_A_84_48#_M1009_g N_Z_c_1015_n 0.0108754f $X=0.925 $Y=0.74 $X2=0 $Y2=0
cc_300 N_A_84_48#_M1011_g N_Z_c_1015_n 0.00906272f $X=1.38 $Y=0.74 $X2=0 $Y2=0
cc_301 N_A_84_48#_c_329_p N_Z_c_1015_n 0.0291873f $X=3.49 $Y=1.485 $X2=0 $Y2=0
cc_302 N_A_84_48#_c_217_n N_Z_c_1015_n 0.00280257f $X=3.795 $Y=1.542 $X2=0 $Y2=0
cc_303 N_A_84_48#_c_219_n N_Z_c_1022_n 0.0139827f $X=0.96 $Y=1.765 $X2=0 $Y2=0
cc_304 N_A_84_48#_c_220_n N_Z_c_1022_n 0.0151589f $X=1.41 $Y=1.765 $X2=0 $Y2=0
cc_305 N_A_84_48#_c_329_p N_Z_c_1022_n 0.0358513f $X=3.49 $Y=1.485 $X2=0 $Y2=0
cc_306 N_A_84_48#_c_217_n N_Z_c_1022_n 0.00850771f $X=3.795 $Y=1.542 $X2=0 $Y2=0
cc_307 N_A_84_48#_M1009_g N_Z_c_1041_n 5.43234e-19 $X=0.925 $Y=0.74 $X2=0 $Y2=0
cc_308 N_A_84_48#_M1011_g N_Z_c_1041_n 0.00600998f $X=1.38 $Y=0.74 $X2=0 $Y2=0
cc_309 N_A_84_48#_M1029_g N_Z_c_1041_n 0.00618702f $X=1.81 $Y=0.74 $X2=0 $Y2=0
cc_310 N_A_84_48#_M1032_g N_Z_c_1041_n 4.62714e-19 $X=2.31 $Y=0.74 $X2=0 $Y2=0
cc_311 N_A_84_48#_c_221_n N_Z_c_1045_n 0.00898134f $X=1.91 $Y=1.765 $X2=0 $Y2=0
cc_312 N_A_84_48#_c_222_n N_Z_c_1045_n 6.10637e-19 $X=2.36 $Y=1.765 $X2=0 $Y2=0
cc_313 N_A_84_48#_M1029_g N_Z_c_1016_n 0.00930697f $X=1.81 $Y=0.74 $X2=0 $Y2=0
cc_314 N_A_84_48#_M1032_g N_Z_c_1016_n 0.0128277f $X=2.31 $Y=0.74 $X2=0 $Y2=0
cc_315 N_A_84_48#_c_329_p N_Z_c_1016_n 0.0492574f $X=3.49 $Y=1.485 $X2=0 $Y2=0
cc_316 N_A_84_48#_c_217_n N_Z_c_1016_n 0.00387231f $X=3.795 $Y=1.542 $X2=0 $Y2=0
cc_317 N_A_84_48#_c_221_n N_Z_c_1023_n 0.0120074f $X=1.91 $Y=1.765 $X2=0 $Y2=0
cc_318 N_A_84_48#_c_222_n N_Z_c_1023_n 0.0120074f $X=2.36 $Y=1.765 $X2=0 $Y2=0
cc_319 N_A_84_48#_c_329_p N_Z_c_1023_n 0.0417603f $X=3.49 $Y=1.485 $X2=0 $Y2=0
cc_320 N_A_84_48#_c_217_n N_Z_c_1023_n 0.00740856f $X=3.795 $Y=1.542 $X2=0 $Y2=0
cc_321 N_A_84_48#_c_221_n N_Z_c_1055_n 6.10637e-19 $X=1.91 $Y=1.765 $X2=0 $Y2=0
cc_322 N_A_84_48#_c_222_n N_Z_c_1055_n 0.00898134f $X=2.36 $Y=1.765 $X2=0 $Y2=0
cc_323 N_A_84_48#_c_223_n N_Z_c_1055_n 0.00880308f $X=2.81 $Y=1.765 $X2=0 $Y2=0
cc_324 N_A_84_48#_c_224_n N_Z_c_1055_n 5.78196e-19 $X=3.31 $Y=1.765 $X2=0 $Y2=0
cc_325 N_A_84_48#_M1033_g N_Z_c_1059_n 0.00620791f $X=2.81 $Y=0.74 $X2=0 $Y2=0
cc_326 N_A_84_48#_M1034_g N_Z_c_1059_n 4.62024e-19 $X=3.325 $Y=0.74 $X2=0 $Y2=0
cc_327 N_A_84_48#_c_223_n N_Z_c_1024_n 0.0122806f $X=2.81 $Y=1.765 $X2=0 $Y2=0
cc_328 N_A_84_48#_c_224_n N_Z_c_1024_n 0.0122806f $X=3.31 $Y=1.765 $X2=0 $Y2=0
cc_329 N_A_84_48#_c_329_p N_Z_c_1024_n 0.0455181f $X=3.49 $Y=1.485 $X2=0 $Y2=0
cc_330 N_A_84_48#_c_217_n N_Z_c_1024_n 0.0086117f $X=3.795 $Y=1.542 $X2=0 $Y2=0
cc_331 N_A_84_48#_M1033_g N_Z_c_1017_n 0.00938204f $X=2.81 $Y=0.74 $X2=0 $Y2=0
cc_332 N_A_84_48#_M1034_g N_Z_c_1017_n 0.0130129f $X=3.325 $Y=0.74 $X2=0 $Y2=0
cc_333 N_A_84_48#_M1036_g N_Z_c_1017_n 0.00461775f $X=3.81 $Y=0.74 $X2=0 $Y2=0
cc_334 N_A_84_48#_c_329_p N_Z_c_1017_n 0.0678816f $X=3.49 $Y=1.485 $X2=0 $Y2=0
cc_335 N_A_84_48#_c_214_n N_Z_c_1017_n 0.0049593f $X=3.87 $Y=1.565 $X2=0 $Y2=0
cc_336 N_A_84_48#_c_217_n N_Z_c_1017_n 0.0077314f $X=3.795 $Y=1.542 $X2=0 $Y2=0
cc_337 N_A_84_48#_c_224_n N_Z_c_1025_n 6.68855e-19 $X=3.31 $Y=1.765 $X2=0 $Y2=0
cc_338 N_A_84_48#_c_329_p N_Z_c_1025_n 0.0275262f $X=3.49 $Y=1.485 $X2=0 $Y2=0
cc_339 N_A_84_48#_c_226_n N_Z_c_1025_n 0.00160357f $X=3.955 $Y=2.05 $X2=0 $Y2=0
cc_340 N_A_84_48#_c_217_n N_Z_c_1025_n 0.00802989f $X=3.795 $Y=1.542 $X2=0 $Y2=0
cc_341 N_A_84_48#_c_223_n N_Z_c_1075_n 6.54588e-19 $X=2.81 $Y=1.765 $X2=0 $Y2=0
cc_342 N_A_84_48#_c_224_n N_Z_c_1075_n 0.00893843f $X=3.31 $Y=1.765 $X2=0 $Y2=0
cc_343 N_A_84_48#_M1036_g N_Z_c_1077_n 0.00457683f $X=3.81 $Y=0.74 $X2=0 $Y2=0
cc_344 N_A_84_48#_c_218_n N_Z_c_1026_n 0.00225616f $X=0.51 $Y=1.765 $X2=0 $Y2=0
cc_345 N_A_84_48#_c_219_n N_Z_c_1026_n 8.92594e-19 $X=0.96 $Y=1.765 $X2=0 $Y2=0
cc_346 N_A_84_48#_c_217_n N_Z_c_1026_n 0.00178968f $X=3.795 $Y=1.542 $X2=0 $Y2=0
cc_347 N_A_84_48#_M1011_g N_Z_c_1018_n 0.00277555f $X=1.38 $Y=0.74 $X2=0 $Y2=0
cc_348 N_A_84_48#_M1029_g N_Z_c_1018_n 0.00277555f $X=1.81 $Y=0.74 $X2=0 $Y2=0
cc_349 N_A_84_48#_c_329_p N_Z_c_1018_n 0.0271537f $X=3.49 $Y=1.485 $X2=0 $Y2=0
cc_350 N_A_84_48#_c_217_n N_Z_c_1018_n 0.002312f $X=3.795 $Y=1.542 $X2=0 $Y2=0
cc_351 N_A_84_48#_c_221_n N_Z_c_1027_n 7.14845e-19 $X=1.91 $Y=1.765 $X2=0 $Y2=0
cc_352 N_A_84_48#_c_329_p N_Z_c_1027_n 0.0277622f $X=3.49 $Y=1.485 $X2=0 $Y2=0
cc_353 N_A_84_48#_c_217_n N_Z_c_1027_n 0.00824682f $X=3.795 $Y=1.542 $X2=0 $Y2=0
cc_354 N_A_84_48#_c_222_n N_Z_c_1028_n 6.83942e-19 $X=2.36 $Y=1.765 $X2=0 $Y2=0
cc_355 N_A_84_48#_c_223_n N_Z_c_1028_n 6.83942e-19 $X=2.81 $Y=1.765 $X2=0 $Y2=0
cc_356 N_A_84_48#_c_329_p N_Z_c_1028_n 0.0276944f $X=3.49 $Y=1.485 $X2=0 $Y2=0
cc_357 N_A_84_48#_c_217_n N_Z_c_1028_n 0.00762283f $X=3.795 $Y=1.542 $X2=0 $Y2=0
cc_358 N_A_84_48#_M1033_g N_Z_c_1019_n 0.00317348f $X=2.81 $Y=0.74 $X2=0 $Y2=0
cc_359 N_A_84_48#_c_329_p N_Z_c_1019_n 0.0272627f $X=3.49 $Y=1.485 $X2=0 $Y2=0
cc_360 N_A_84_48#_c_217_n N_Z_c_1019_n 0.0039304f $X=3.795 $Y=1.542 $X2=0 $Y2=0
cc_361 N_A_84_48#_M1005_g Z 0.00463107f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_362 N_A_84_48#_M1009_g Z 0.00294797f $X=0.925 $Y=0.74 $X2=0 $Y2=0
cc_363 N_A_84_48#_M1005_g Z 0.00883951f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_364 N_A_84_48#_c_218_n Z 0.00286344f $X=0.51 $Y=1.765 $X2=0 $Y2=0
cc_365 N_A_84_48#_M1009_g Z 0.00469957f $X=0.925 $Y=0.74 $X2=0 $Y2=0
cc_366 N_A_84_48#_c_219_n Z 0.00145091f $X=0.96 $Y=1.765 $X2=0 $Y2=0
cc_367 N_A_84_48#_c_329_p Z 0.0227592f $X=3.49 $Y=1.485 $X2=0 $Y2=0
cc_368 N_A_84_48#_c_217_n Z 0.0453979f $X=3.795 $Y=1.542 $X2=0 $Y2=0
cc_369 N_A_84_48#_M1005_g N_Z_c_1103_n 0.00480711f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_370 N_A_84_48#_M1009_g N_Z_c_1103_n 0.00588517f $X=0.925 $Y=0.74 $X2=0 $Y2=0
cc_371 N_A_84_48#_M1011_g N_Z_c_1103_n 5.35511e-19 $X=1.38 $Y=0.74 $X2=0 $Y2=0
cc_372 N_A_84_48#_c_242_p N_VPWR_M1016_s 0.00873006f $X=7.585 $Y=2.135 $X2=-0.19
+ $Y2=-0.245
cc_373 N_A_84_48#_c_242_p N_VPWR_M1022_s 0.00794746f $X=7.585 $Y=2.135 $X2=0
+ $Y2=0
cc_374 N_A_84_48#_c_242_p N_VPWR_M1024_s 0.00794599f $X=7.585 $Y=2.135 $X2=0
+ $Y2=0
cc_375 N_A_84_48#_c_242_p N_VPWR_M1028_s 0.00683659f $X=7.585 $Y=2.135 $X2=0
+ $Y2=0
cc_376 N_A_84_48#_c_258_p N_VPWR_M1028_s 0.00816719f $X=7.67 $Y=2.135 $X2=0
+ $Y2=0
cc_377 N_A_84_48#_c_227_n N_VPWR_M1002_d 0.00738851f $X=9.665 $Y=2.305 $X2=0
+ $Y2=0
cc_378 N_A_84_48#_c_229_n N_VPWR_M1007_s 0.00365985f $X=10.145 $Y=1.805 $X2=0
+ $Y2=0
cc_379 N_A_84_48#_c_227_n N_VPWR_c_1154_n 0.0202249f $X=9.665 $Y=2.305 $X2=0
+ $Y2=0
cc_380 N_A_84_48#_c_228_n N_VPWR_c_1154_n 0.0161582f $X=9.83 $Y=2.815 $X2=0
+ $Y2=0
cc_381 N_A_84_48#_c_228_n N_VPWR_c_1156_n 0.0229093f $X=9.83 $Y=2.815 $X2=0
+ $Y2=0
cc_382 N_A_84_48#_c_229_n N_VPWR_c_1156_n 0.012565f $X=10.145 $Y=1.805 $X2=0
+ $Y2=0
cc_383 N_A_84_48#_c_218_n N_VPWR_c_1157_n 0.00278271f $X=0.51 $Y=1.765 $X2=0
+ $Y2=0
cc_384 N_A_84_48#_c_219_n N_VPWR_c_1157_n 0.00278271f $X=0.96 $Y=1.765 $X2=0
+ $Y2=0
cc_385 N_A_84_48#_c_220_n N_VPWR_c_1157_n 0.00278257f $X=1.41 $Y=1.765 $X2=0
+ $Y2=0
cc_386 N_A_84_48#_c_221_n N_VPWR_c_1157_n 0.00278271f $X=1.91 $Y=1.765 $X2=0
+ $Y2=0
cc_387 N_A_84_48#_c_222_n N_VPWR_c_1157_n 0.00278271f $X=2.36 $Y=1.765 $X2=0
+ $Y2=0
cc_388 N_A_84_48#_c_223_n N_VPWR_c_1157_n 0.00278271f $X=2.81 $Y=1.765 $X2=0
+ $Y2=0
cc_389 N_A_84_48#_c_224_n N_VPWR_c_1157_n 0.00278271f $X=3.31 $Y=1.765 $X2=0
+ $Y2=0
cc_390 N_A_84_48#_c_225_n N_VPWR_c_1157_n 0.00278271f $X=3.795 $Y=1.765 $X2=0
+ $Y2=0
cc_391 N_A_84_48#_c_228_n N_VPWR_c_1161_n 0.0123628f $X=9.83 $Y=2.815 $X2=0
+ $Y2=0
cc_392 N_A_84_48#_c_218_n N_VPWR_c_1148_n 0.00357334f $X=0.51 $Y=1.765 $X2=0
+ $Y2=0
cc_393 N_A_84_48#_c_219_n N_VPWR_c_1148_n 0.00353823f $X=0.96 $Y=1.765 $X2=0
+ $Y2=0
cc_394 N_A_84_48#_c_220_n N_VPWR_c_1148_n 0.00354283f $X=1.41 $Y=1.765 $X2=0
+ $Y2=0
cc_395 N_A_84_48#_c_221_n N_VPWR_c_1148_n 0.00354284f $X=1.91 $Y=1.765 $X2=0
+ $Y2=0
cc_396 N_A_84_48#_c_222_n N_VPWR_c_1148_n 0.00353823f $X=2.36 $Y=1.765 $X2=0
+ $Y2=0
cc_397 N_A_84_48#_c_223_n N_VPWR_c_1148_n 0.00354284f $X=2.81 $Y=1.765 $X2=0
+ $Y2=0
cc_398 N_A_84_48#_c_224_n N_VPWR_c_1148_n 0.00354611f $X=3.31 $Y=1.765 $X2=0
+ $Y2=0
cc_399 N_A_84_48#_c_225_n N_VPWR_c_1148_n 0.00354367f $X=3.795 $Y=1.765 $X2=0
+ $Y2=0
cc_400 N_A_84_48#_c_228_n N_VPWR_c_1148_n 0.0101999f $X=9.83 $Y=2.815 $X2=0
+ $Y2=0
cc_401 N_A_84_48#_M1005_g N_A_27_74#_c_1277_n 0.00159289f $X=0.495 $Y=0.74 $X2=0
+ $Y2=0
cc_402 N_A_84_48#_M1005_g N_A_27_74#_c_1278_n 0.0132617f $X=0.495 $Y=0.74 $X2=0
+ $Y2=0
cc_403 N_A_84_48#_M1009_g N_A_27_74#_c_1278_n 0.0108851f $X=0.925 $Y=0.74 $X2=0
+ $Y2=0
cc_404 N_A_84_48#_M1011_g N_A_27_74#_c_1302_n 0.00394726f $X=1.38 $Y=0.74 $X2=0
+ $Y2=0
cc_405 N_A_84_48#_M1011_g N_A_27_74#_c_1280_n 0.0108851f $X=1.38 $Y=0.74 $X2=0
+ $Y2=0
cc_406 N_A_84_48#_M1029_g N_A_27_74#_c_1280_n 0.0111293f $X=1.81 $Y=0.74 $X2=0
+ $Y2=0
cc_407 N_A_84_48#_M1032_g N_A_27_74#_c_1305_n 0.0061935f $X=2.31 $Y=0.74 $X2=0
+ $Y2=0
cc_408 N_A_84_48#_M1033_g N_A_27_74#_c_1305_n 4.62714e-19 $X=2.81 $Y=0.74 $X2=0
+ $Y2=0
cc_409 N_A_84_48#_M1032_g N_A_27_74#_c_1281_n 0.00822804f $X=2.31 $Y=0.74 $X2=0
+ $Y2=0
cc_410 N_A_84_48#_M1033_g N_A_27_74#_c_1281_n 0.0115976f $X=2.81 $Y=0.74 $X2=0
+ $Y2=0
cc_411 N_A_84_48#_M1034_g N_A_27_74#_c_1309_n 0.00542481f $X=3.325 $Y=0.74 $X2=0
+ $Y2=0
cc_412 N_A_84_48#_M1036_g N_A_27_74#_c_1309_n 7.18008e-19 $X=3.81 $Y=0.74 $X2=0
+ $Y2=0
cc_413 N_A_84_48#_M1034_g N_A_27_74#_c_1282_n 0.00879688f $X=3.325 $Y=0.74 $X2=0
+ $Y2=0
cc_414 N_A_84_48#_M1036_g N_A_27_74#_c_1282_n 0.0123192f $X=3.81 $Y=0.74 $X2=0
+ $Y2=0
cc_415 N_A_84_48#_M1036_g N_A_27_74#_c_1283_n 4.60332e-19 $X=3.81 $Y=0.74 $X2=0
+ $Y2=0
cc_416 N_A_84_48#_M1036_g N_A_27_74#_c_1285_n 0.00514561f $X=3.81 $Y=0.74 $X2=0
+ $Y2=0
cc_417 N_A_84_48#_c_214_n N_A_27_74#_c_1285_n 0.00936976f $X=3.87 $Y=1.565 $X2=0
+ $Y2=0
cc_418 N_A_84_48#_c_242_p N_A_27_74#_c_1287_n 0.0140951f $X=7.585 $Y=2.135 $X2=0
+ $Y2=0
cc_419 N_A_84_48#_c_242_p N_A_27_74#_c_1289_n 0.0155632f $X=7.585 $Y=2.135 $X2=0
+ $Y2=0
cc_420 N_A_84_48#_c_242_p N_A_27_74#_c_1291_n 0.0232299f $X=7.585 $Y=2.135 $X2=0
+ $Y2=0
cc_421 N_A_84_48#_M1032_g N_A_27_74#_c_1294_n 0.00294698f $X=2.31 $Y=0.74 $X2=0
+ $Y2=0
cc_422 N_A_84_48#_M1034_g N_A_27_74#_c_1295_n 0.00270885f $X=3.325 $Y=0.74 $X2=0
+ $Y2=0
cc_423 N_A_84_48#_c_242_p N_A_27_74#_c_1296_n 0.00967233f $X=7.585 $Y=2.135
+ $X2=0 $Y2=0
cc_424 N_A_84_48#_c_242_p N_A_27_74#_c_1297_n 0.00749426f $X=7.585 $Y=2.135
+ $X2=0 $Y2=0
cc_425 N_A_84_48#_c_242_p N_A_27_74#_c_1298_n 0.00835391f $X=7.585 $Y=2.135
+ $X2=0 $Y2=0
cc_426 N_A_84_48#_c_280_p N_VGND_M1018_s 0.00916777f $X=10.145 $Y=0.925 $X2=0
+ $Y2=0
cc_427 N_A_84_48#_c_216_n N_VGND_M1018_s 0.0037774f $X=10.23 $Y=1.72 $X2=0 $Y2=0
cc_428 N_A_84_48#_c_215_n N_VGND_c_1446_n 0.0181878f $X=9.845 $Y=0.505 $X2=0
+ $Y2=0
cc_429 N_A_84_48#_c_215_n N_VGND_c_1448_n 0.0104513f $X=9.845 $Y=0.505 $X2=0
+ $Y2=0
cc_430 N_A_84_48#_c_280_p N_VGND_c_1448_n 0.00936242f $X=10.145 $Y=0.925 $X2=0
+ $Y2=0
cc_431 N_A_84_48#_M1005_g N_VGND_c_1449_n 0.00278271f $X=0.495 $Y=0.74 $X2=0
+ $Y2=0
cc_432 N_A_84_48#_M1009_g N_VGND_c_1449_n 0.00278271f $X=0.925 $Y=0.74 $X2=0
+ $Y2=0
cc_433 N_A_84_48#_M1011_g N_VGND_c_1449_n 0.00278271f $X=1.38 $Y=0.74 $X2=0
+ $Y2=0
cc_434 N_A_84_48#_M1029_g N_VGND_c_1449_n 0.00278271f $X=1.81 $Y=0.74 $X2=0
+ $Y2=0
cc_435 N_A_84_48#_M1032_g N_VGND_c_1449_n 0.00278247f $X=2.31 $Y=0.74 $X2=0
+ $Y2=0
cc_436 N_A_84_48#_M1033_g N_VGND_c_1449_n 0.00278271f $X=2.81 $Y=0.74 $X2=0
+ $Y2=0
cc_437 N_A_84_48#_M1034_g N_VGND_c_1449_n 0.00278262f $X=3.325 $Y=0.74 $X2=0
+ $Y2=0
cc_438 N_A_84_48#_M1036_g N_VGND_c_1449_n 0.00278271f $X=3.81 $Y=0.74 $X2=0
+ $Y2=0
cc_439 N_A_84_48#_c_215_n N_VGND_c_1457_n 0.0114427f $X=9.845 $Y=0.505 $X2=0
+ $Y2=0
cc_440 N_A_84_48#_M1005_g N_VGND_c_1460_n 0.00357086f $X=0.495 $Y=0.74 $X2=0
+ $Y2=0
cc_441 N_A_84_48#_M1009_g N_VGND_c_1460_n 0.00353674f $X=0.925 $Y=0.74 $X2=0
+ $Y2=0
cc_442 N_A_84_48#_M1011_g N_VGND_c_1460_n 0.00353674f $X=1.38 $Y=0.74 $X2=0
+ $Y2=0
cc_443 N_A_84_48#_M1029_g N_VGND_c_1460_n 0.00354087f $X=1.81 $Y=0.74 $X2=0
+ $Y2=0
cc_444 N_A_84_48#_M1032_g N_VGND_c_1460_n 0.00354743f $X=2.31 $Y=0.74 $X2=0
+ $Y2=0
cc_445 N_A_84_48#_M1033_g N_VGND_c_1460_n 0.00354875f $X=2.81 $Y=0.74 $X2=0
+ $Y2=0
cc_446 N_A_84_48#_M1034_g N_VGND_c_1460_n 0.0035474f $X=3.325 $Y=0.74 $X2=0
+ $Y2=0
cc_447 N_A_84_48#_M1036_g N_VGND_c_1460_n 0.0035405f $X=3.81 $Y=0.74 $X2=0 $Y2=0
cc_448 N_A_84_48#_c_215_n N_VGND_c_1460_n 0.00909435f $X=9.845 $Y=0.505 $X2=0
+ $Y2=0
cc_449 N_A_84_48#_c_280_p N_VGND_c_1460_n 0.00616274f $X=10.145 $Y=0.925 $X2=0
+ $Y2=0
cc_450 N_A_833_48#_c_479_n N_TE_B_c_643_n 0.0114525f $X=4.595 $Y=1.26 $X2=0
+ $Y2=0
cc_451 N_A_833_48#_c_480_n N_TE_B_c_644_n 0.0114525f $X=4.315 $Y=1.26 $X2=0
+ $Y2=0
cc_452 N_A_833_48#_c_482_n N_TE_B_c_645_n 0.0114525f $X=5.025 $Y=1.26 $X2=0
+ $Y2=0
cc_453 N_A_833_48#_c_484_n N_TE_B_c_646_n 0.0114525f $X=5.455 $Y=1.26 $X2=0
+ $Y2=0
cc_454 N_A_833_48#_c_486_n N_TE_B_c_647_n 0.0114525f $X=5.885 $Y=1.26 $X2=0
+ $Y2=0
cc_455 N_A_833_48#_c_488_n N_TE_B_c_648_n 0.0114525f $X=6.315 $Y=1.26 $X2=0
+ $Y2=0
cc_456 N_A_833_48#_c_490_n N_TE_B_c_649_n 0.0114525f $X=6.745 $Y=1.26 $X2=0
+ $Y2=0
cc_457 N_A_833_48#_c_513_n N_TE_B_c_677_n 0.00111159f $X=8.095 $Y=1.925 $X2=0
+ $Y2=0
cc_458 N_A_833_48#_c_492_n N_TE_B_c_650_n 0.0114525f $X=7.175 $Y=1.26 $X2=0
+ $Y2=0
cc_459 N_A_833_48#_c_504_n N_TE_B_c_679_n 0.00123064f $X=8.01 $Y=1.8 $X2=0 $Y2=0
cc_460 N_A_833_48#_c_513_n N_TE_B_c_679_n 0.012258f $X=8.095 $Y=1.925 $X2=0
+ $Y2=0
cc_461 N_A_833_48#_c_494_n N_TE_B_c_652_n 0.00317119f $X=7.72 $Y=1.26 $X2=0
+ $Y2=0
cc_462 N_A_833_48#_c_504_n N_TE_B_c_652_n 0.00462536f $X=8.01 $Y=1.8 $X2=0 $Y2=0
cc_463 N_A_833_48#_c_506_n N_TE_B_c_652_n 0.00756727f $X=8.565 $Y=0.505 $X2=0
+ $Y2=0
cc_464 N_A_833_48#_c_507_n N_TE_B_c_652_n 0.00456231f $X=8.985 $Y=0.515 $X2=0
+ $Y2=0
cc_465 N_A_833_48#_c_509_n N_TE_B_c_682_n 0.0110783f $X=8.77 $Y=1.965 $X2=0
+ $Y2=0
cc_466 N_A_833_48#_c_506_n N_TE_B_c_653_n 0.00516259f $X=8.565 $Y=0.505 $X2=0
+ $Y2=0
cc_467 N_A_833_48#_c_507_n N_TE_B_c_653_n 0.00794536f $X=8.985 $Y=0.515 $X2=0
+ $Y2=0
cc_468 N_A_833_48#_c_496_n N_TE_B_c_654_n 0.0114525f $X=4.67 $Y=1.26 $X2=0 $Y2=0
cc_469 N_A_833_48#_c_497_n N_TE_B_c_655_n 0.0114525f $X=5.1 $Y=1.26 $X2=0 $Y2=0
cc_470 N_A_833_48#_c_498_n N_TE_B_c_656_n 0.0114525f $X=5.53 $Y=1.26 $X2=0 $Y2=0
cc_471 N_A_833_48#_c_499_n N_TE_B_c_657_n 0.0114525f $X=5.96 $Y=1.26 $X2=0 $Y2=0
cc_472 N_A_833_48#_c_500_n N_TE_B_c_658_n 0.0114525f $X=6.39 $Y=1.26 $X2=0 $Y2=0
cc_473 N_A_833_48#_c_501_n N_TE_B_c_659_n 0.0114525f $X=6.82 $Y=1.26 $X2=0 $Y2=0
cc_474 N_A_833_48#_c_502_n N_TE_B_c_660_n 0.0114525f $X=7.25 $Y=1.26 $X2=0 $Y2=0
cc_475 N_A_833_48#_c_504_n N_TE_B_c_660_n 0.00777303f $X=8.01 $Y=1.8 $X2=0 $Y2=0
cc_476 N_A_833_48#_c_504_n TE_B 0.0295862f $X=8.01 $Y=1.8 $X2=0 $Y2=0
cc_477 N_A_833_48#_c_506_n TE_B 9.40747e-19 $X=8.565 $Y=0.505 $X2=0 $Y2=0
cc_478 N_A_833_48#_c_507_n TE_B 0.0751834f $X=8.985 $Y=0.515 $X2=0 $Y2=0
cc_479 N_A_833_48#_c_509_n TE_B 0.0455344f $X=8.77 $Y=1.965 $X2=0 $Y2=0
cc_480 N_A_833_48#_c_504_n N_TE_B_c_662_n 0.0129759f $X=8.01 $Y=1.8 $X2=0 $Y2=0
cc_481 N_A_833_48#_c_507_n N_TE_B_c_662_n 0.00437509f $X=8.985 $Y=0.515 $X2=0
+ $Y2=0
cc_482 N_A_833_48#_c_509_n N_TE_B_c_662_n 0.0277616f $X=8.77 $Y=1.965 $X2=0
+ $Y2=0
cc_483 N_A_833_48#_c_509_n N_A_c_831_n 7.50016e-19 $X=8.77 $Y=1.965 $X2=-0.19
+ $Y2=-0.245
cc_484 N_A_833_48#_c_513_n N_A_28_368#_M1030_d 9.20758e-19 $X=8.095 $Y=1.925
+ $X2=0 $Y2=0
cc_485 N_A_833_48#_c_509_n N_A_28_368#_M1030_d 0.00232265f $X=8.77 $Y=1.965
+ $X2=0 $Y2=0
cc_486 N_A_833_48#_c_478_n N_A_27_74#_c_1282_n 9.48753e-19 $X=4.24 $Y=1.185
+ $X2=0 $Y2=0
cc_487 N_A_833_48#_c_478_n N_A_27_74#_c_1283_n 9.29165e-19 $X=4.24 $Y=1.185
+ $X2=0 $Y2=0
cc_488 N_A_833_48#_c_478_n N_A_27_74#_c_1284_n 0.00741157f $X=4.24 $Y=1.185
+ $X2=0 $Y2=0
cc_489 N_A_833_48#_c_479_n N_A_27_74#_c_1284_n 0.00839174f $X=4.595 $Y=1.26
+ $X2=0 $Y2=0
cc_490 N_A_833_48#_c_480_n N_A_27_74#_c_1284_n 0.0049686f $X=4.315 $Y=1.26 $X2=0
+ $Y2=0
cc_491 N_A_833_48#_c_481_n N_A_27_74#_c_1284_n 0.00605219f $X=4.67 $Y=1.185
+ $X2=0 $Y2=0
cc_492 N_A_833_48#_c_496_n N_A_27_74#_c_1284_n 0.00349533f $X=4.67 $Y=1.26 $X2=0
+ $Y2=0
cc_493 N_A_833_48#_c_481_n N_A_27_74#_c_1286_n 0.00112526f $X=4.67 $Y=1.185
+ $X2=0 $Y2=0
cc_494 N_A_833_48#_c_483_n N_A_27_74#_c_1286_n 0.00943354f $X=5.1 $Y=1.185 $X2=0
+ $Y2=0
cc_495 N_A_833_48#_c_485_n N_A_27_74#_c_1286_n 3.92634e-19 $X=5.53 $Y=1.185
+ $X2=0 $Y2=0
cc_496 N_A_833_48#_c_484_n N_A_27_74#_c_1287_n 0.00945505f $X=5.455 $Y=1.26
+ $X2=0 $Y2=0
cc_497 N_A_833_48#_c_497_n N_A_27_74#_c_1287_n 0.00691356f $X=5.1 $Y=1.26 $X2=0
+ $Y2=0
cc_498 N_A_833_48#_c_498_n N_A_27_74#_c_1287_n 0.00675192f $X=5.53 $Y=1.26 $X2=0
+ $Y2=0
cc_499 N_A_833_48#_c_483_n N_A_27_74#_c_1288_n 3.93664e-19 $X=5.1 $Y=1.185 $X2=0
+ $Y2=0
cc_500 N_A_833_48#_c_485_n N_A_27_74#_c_1288_n 0.0106304f $X=5.53 $Y=1.185 $X2=0
+ $Y2=0
cc_501 N_A_833_48#_c_486_n N_A_27_74#_c_1288_n 0.00787652f $X=5.885 $Y=1.26
+ $X2=0 $Y2=0
cc_502 N_A_833_48#_c_487_n N_A_27_74#_c_1288_n 0.00126428f $X=5.96 $Y=1.185
+ $X2=0 $Y2=0
cc_503 N_A_833_48#_c_498_n N_A_27_74#_c_1288_n 0.00308673f $X=5.53 $Y=1.26 $X2=0
+ $Y2=0
cc_504 N_A_833_48#_c_486_n N_A_27_74#_c_1289_n 0.0028859f $X=5.885 $Y=1.26 $X2=0
+ $Y2=0
cc_505 N_A_833_48#_c_488_n N_A_27_74#_c_1289_n 0.00777301f $X=6.315 $Y=1.26
+ $X2=0 $Y2=0
cc_506 N_A_833_48#_c_499_n N_A_27_74#_c_1289_n 0.00743366f $X=5.96 $Y=1.26 $X2=0
+ $Y2=0
cc_507 N_A_833_48#_c_500_n N_A_27_74#_c_1289_n 0.00675192f $X=6.39 $Y=1.26 $X2=0
+ $Y2=0
cc_508 N_A_833_48#_c_487_n N_A_27_74#_c_1290_n 4.44315e-19 $X=5.96 $Y=1.185
+ $X2=0 $Y2=0
cc_509 N_A_833_48#_c_489_n N_A_27_74#_c_1290_n 0.0106978f $X=6.39 $Y=1.185 $X2=0
+ $Y2=0
cc_510 N_A_833_48#_c_490_n N_A_27_74#_c_1290_n 0.00787652f $X=6.745 $Y=1.26
+ $X2=0 $Y2=0
cc_511 N_A_833_48#_c_491_n N_A_27_74#_c_1290_n 0.00126428f $X=6.82 $Y=1.185
+ $X2=0 $Y2=0
cc_512 N_A_833_48#_c_500_n N_A_27_74#_c_1290_n 0.00333129f $X=6.39 $Y=1.26 $X2=0
+ $Y2=0
cc_513 N_A_833_48#_c_490_n N_A_27_74#_c_1291_n 0.0028859f $X=6.745 $Y=1.26 $X2=0
+ $Y2=0
cc_514 N_A_833_48#_c_492_n N_A_27_74#_c_1291_n 0.00777301f $X=7.175 $Y=1.26
+ $X2=0 $Y2=0
cc_515 N_A_833_48#_c_494_n N_A_27_74#_c_1291_n 0.00293227f $X=7.72 $Y=1.26 $X2=0
+ $Y2=0
cc_516 N_A_833_48#_c_501_n N_A_27_74#_c_1291_n 0.00743366f $X=6.82 $Y=1.26 $X2=0
+ $Y2=0
cc_517 N_A_833_48#_c_502_n N_A_27_74#_c_1291_n 0.00701045f $X=7.25 $Y=1.26 $X2=0
+ $Y2=0
cc_518 N_A_833_48#_c_504_n N_A_27_74#_c_1291_n 0.00812414f $X=8.01 $Y=1.8 $X2=0
+ $Y2=0
cc_519 N_A_833_48#_c_491_n N_A_27_74#_c_1292_n 4.44315e-19 $X=6.82 $Y=1.185
+ $X2=0 $Y2=0
cc_520 N_A_833_48#_c_493_n N_A_27_74#_c_1292_n 0.011062f $X=7.25 $Y=1.185 $X2=0
+ $Y2=0
cc_521 N_A_833_48#_c_494_n N_A_27_74#_c_1292_n 0.00763221f $X=7.72 $Y=1.26 $X2=0
+ $Y2=0
cc_522 N_A_833_48#_c_495_n N_A_27_74#_c_1292_n 0.00481512f $X=7.795 $Y=1.185
+ $X2=0 $Y2=0
cc_523 N_A_833_48#_c_502_n N_A_27_74#_c_1292_n 0.00333129f $X=7.25 $Y=1.26 $X2=0
+ $Y2=0
cc_524 N_A_833_48#_c_503_n N_A_27_74#_c_1292_n 0.00117099f $X=7.87 $Y=0.505
+ $X2=0 $Y2=0
cc_525 N_A_833_48#_c_504_n N_A_27_74#_c_1292_n 0.0123137f $X=8.01 $Y=1.8 $X2=0
+ $Y2=0
cc_526 N_A_833_48#_c_505_n N_A_27_74#_c_1292_n 0.0423085f $X=8.095 $Y=0.675
+ $X2=0 $Y2=0
cc_527 N_A_833_48#_c_481_n N_A_27_74#_c_1296_n 0.00190168f $X=4.67 $Y=1.185
+ $X2=0 $Y2=0
cc_528 N_A_833_48#_c_482_n N_A_27_74#_c_1296_n 0.00829432f $X=5.025 $Y=1.26
+ $X2=0 $Y2=0
cc_529 N_A_833_48#_c_483_n N_A_27_74#_c_1296_n 0.00128545f $X=5.1 $Y=1.185 $X2=0
+ $Y2=0
cc_530 N_A_833_48#_c_496_n N_A_27_74#_c_1296_n 0.00207909f $X=4.67 $Y=1.26 $X2=0
+ $Y2=0
cc_531 N_A_833_48#_c_497_n N_A_27_74#_c_1296_n 0.00346919f $X=5.1 $Y=1.26 $X2=0
+ $Y2=0
cc_532 N_A_833_48#_c_486_n N_A_27_74#_c_1297_n 0.00231645f $X=5.885 $Y=1.26
+ $X2=0 $Y2=0
cc_533 N_A_833_48#_c_498_n N_A_27_74#_c_1297_n 2.58532e-19 $X=5.53 $Y=1.26 $X2=0
+ $Y2=0
cc_534 N_A_833_48#_c_490_n N_A_27_74#_c_1298_n 0.00231645f $X=6.745 $Y=1.26
+ $X2=0 $Y2=0
cc_535 N_A_833_48#_c_500_n N_A_27_74#_c_1298_n 2.58532e-19 $X=6.39 $Y=1.26 $X2=0
+ $Y2=0
cc_536 N_A_833_48#_c_478_n N_VGND_c_1442_n 0.0100283f $X=4.24 $Y=1.185 $X2=0
+ $Y2=0
cc_537 N_A_833_48#_c_479_n N_VGND_c_1442_n 7.11061e-19 $X=4.595 $Y=1.26 $X2=0
+ $Y2=0
cc_538 N_A_833_48#_c_481_n N_VGND_c_1442_n 0.0108109f $X=4.67 $Y=1.185 $X2=0
+ $Y2=0
cc_539 N_A_833_48#_c_483_n N_VGND_c_1442_n 5.57989e-19 $X=5.1 $Y=1.185 $X2=0
+ $Y2=0
cc_540 N_A_833_48#_c_483_n N_VGND_c_1443_n 0.001891f $X=5.1 $Y=1.185 $X2=0 $Y2=0
cc_541 N_A_833_48#_c_484_n N_VGND_c_1443_n 0.00230361f $X=5.455 $Y=1.26 $X2=0
+ $Y2=0
cc_542 N_A_833_48#_c_485_n N_VGND_c_1443_n 0.001891f $X=5.53 $Y=1.185 $X2=0
+ $Y2=0
cc_543 N_A_833_48#_c_485_n N_VGND_c_1444_n 6.16849e-19 $X=5.53 $Y=1.185 $X2=0
+ $Y2=0
cc_544 N_A_833_48#_c_487_n N_VGND_c_1444_n 0.0128208f $X=5.96 $Y=1.185 $X2=0
+ $Y2=0
cc_545 N_A_833_48#_c_488_n N_VGND_c_1444_n 0.00230361f $X=6.315 $Y=1.26 $X2=0
+ $Y2=0
cc_546 N_A_833_48#_c_489_n N_VGND_c_1444_n 0.00198331f $X=6.39 $Y=1.185 $X2=0
+ $Y2=0
cc_547 N_A_833_48#_c_489_n N_VGND_c_1445_n 6.16849e-19 $X=6.39 $Y=1.185 $X2=0
+ $Y2=0
cc_548 N_A_833_48#_c_491_n N_VGND_c_1445_n 0.0128208f $X=6.82 $Y=1.185 $X2=0
+ $Y2=0
cc_549 N_A_833_48#_c_492_n N_VGND_c_1445_n 0.00230361f $X=7.175 $Y=1.26 $X2=0
+ $Y2=0
cc_550 N_A_833_48#_c_493_n N_VGND_c_1445_n 0.00321968f $X=7.25 $Y=1.185 $X2=0
+ $Y2=0
cc_551 N_A_833_48#_c_505_n N_VGND_c_1445_n 3.11442e-19 $X=8.095 $Y=0.675 $X2=0
+ $Y2=0
cc_552 N_A_833_48#_c_507_n N_VGND_c_1446_n 0.0278867f $X=8.985 $Y=0.515 $X2=0
+ $Y2=0
cc_553 N_A_833_48#_c_478_n N_VGND_c_1449_n 0.00383152f $X=4.24 $Y=1.185 $X2=0
+ $Y2=0
cc_554 N_A_833_48#_c_481_n N_VGND_c_1451_n 0.00383152f $X=4.67 $Y=1.185 $X2=0
+ $Y2=0
cc_555 N_A_833_48#_c_483_n N_VGND_c_1451_n 0.00434272f $X=5.1 $Y=1.185 $X2=0
+ $Y2=0
cc_556 N_A_833_48#_c_485_n N_VGND_c_1453_n 0.00434272f $X=5.53 $Y=1.185 $X2=0
+ $Y2=0
cc_557 N_A_833_48#_c_487_n N_VGND_c_1453_n 0.00383152f $X=5.96 $Y=1.185 $X2=0
+ $Y2=0
cc_558 N_A_833_48#_c_489_n N_VGND_c_1455_n 0.00434272f $X=6.39 $Y=1.185 $X2=0
+ $Y2=0
cc_559 N_A_833_48#_c_491_n N_VGND_c_1455_n 0.00383152f $X=6.82 $Y=1.185 $X2=0
+ $Y2=0
cc_560 N_A_833_48#_c_493_n N_VGND_c_1456_n 0.00434272f $X=7.25 $Y=1.185 $X2=0
+ $Y2=0
cc_561 N_A_833_48#_c_503_n N_VGND_c_1456_n 0.00215305f $X=7.87 $Y=0.505 $X2=0
+ $Y2=0
cc_562 N_A_833_48#_c_505_n N_VGND_c_1456_n 0.0158548f $X=8.095 $Y=0.675 $X2=0
+ $Y2=0
cc_563 N_A_833_48#_c_506_n N_VGND_c_1456_n 0.0129945f $X=8.565 $Y=0.505 $X2=0
+ $Y2=0
cc_564 N_A_833_48#_c_507_n N_VGND_c_1456_n 0.0467562f $X=8.985 $Y=0.515 $X2=0
+ $Y2=0
cc_565 N_A_833_48#_c_478_n N_VGND_c_1460_n 0.00757637f $X=4.24 $Y=1.185 $X2=0
+ $Y2=0
cc_566 N_A_833_48#_c_481_n N_VGND_c_1460_n 0.0075754f $X=4.67 $Y=1.185 $X2=0
+ $Y2=0
cc_567 N_A_833_48#_c_483_n N_VGND_c_1460_n 0.00820284f $X=5.1 $Y=1.185 $X2=0
+ $Y2=0
cc_568 N_A_833_48#_c_485_n N_VGND_c_1460_n 0.00820284f $X=5.53 $Y=1.185 $X2=0
+ $Y2=0
cc_569 N_A_833_48#_c_487_n N_VGND_c_1460_n 0.0075754f $X=5.96 $Y=1.185 $X2=0
+ $Y2=0
cc_570 N_A_833_48#_c_489_n N_VGND_c_1460_n 0.00820284f $X=6.39 $Y=1.185 $X2=0
+ $Y2=0
cc_571 N_A_833_48#_c_491_n N_VGND_c_1460_n 0.0075754f $X=6.82 $Y=1.185 $X2=0
+ $Y2=0
cc_572 N_A_833_48#_c_493_n N_VGND_c_1460_n 0.00825283f $X=7.25 $Y=1.185 $X2=0
+ $Y2=0
cc_573 N_A_833_48#_c_505_n N_VGND_c_1460_n 0.0134631f $X=8.095 $Y=0.675 $X2=0
+ $Y2=0
cc_574 N_A_833_48#_c_506_n N_VGND_c_1460_n 0.0193081f $X=8.565 $Y=0.505 $X2=0
+ $Y2=0
cc_575 N_A_833_48#_c_507_n N_VGND_c_1460_n 0.0385205f $X=8.985 $Y=0.515 $X2=0
+ $Y2=0
cc_576 N_TE_B_c_682_n N_A_c_831_n 0.0362093f $X=9.105 $Y=1.765 $X2=-0.19
+ $Y2=-0.245
cc_577 N_TE_B_c_653_n N_A_c_827_n 0.0133063f $X=9.2 $Y=1.22 $X2=0 $Y2=0
cc_578 TE_B N_A_c_827_n 2.95037e-19 $X=9.275 $Y=1.21 $X2=0 $Y2=0
cc_579 N_TE_B_c_653_n A 2.69981e-19 $X=9.2 $Y=1.22 $X2=0 $Y2=0
cc_580 TE_B A 0.0309922f $X=9.275 $Y=1.21 $X2=0 $Y2=0
cc_581 TE_B N_A_c_830_n 0.00304313f $X=9.275 $Y=1.21 $X2=0 $Y2=0
cc_582 N_TE_B_c_663_n N_A_c_830_n 0.028872f $X=9.11 $Y=1.385 $X2=0 $Y2=0
cc_583 N_TE_B_c_664_n N_A_28_368#_c_882_n 0.00318927f $X=4.26 $Y=1.765 $X2=0
+ $Y2=0
cc_584 N_TE_B_c_664_n N_A_28_368#_c_910_n 4.27119e-19 $X=4.26 $Y=1.765 $X2=0
+ $Y2=0
cc_585 N_TE_B_c_664_n N_A_28_368#_c_927_n 0.00497909f $X=4.26 $Y=1.765 $X2=0
+ $Y2=0
cc_586 N_TE_B_c_667_n N_A_28_368#_c_927_n 5.5844e-19 $X=4.81 $Y=1.765 $X2=0
+ $Y2=0
cc_587 N_TE_B_c_664_n N_A_28_368#_c_912_n 0.00947174f $X=4.26 $Y=1.765 $X2=0
+ $Y2=0
cc_588 N_TE_B_c_667_n N_A_28_368#_c_912_n 0.00947174f $X=4.81 $Y=1.765 $X2=0
+ $Y2=0
cc_589 N_TE_B_c_669_n N_A_28_368#_c_913_n 0.00947174f $X=5.26 $Y=1.765 $X2=0
+ $Y2=0
cc_590 N_TE_B_c_671_n N_A_28_368#_c_913_n 0.00947174f $X=5.81 $Y=1.765 $X2=0
+ $Y2=0
cc_591 N_TE_B_c_673_n N_A_28_368#_c_914_n 0.00947174f $X=6.26 $Y=1.765 $X2=0
+ $Y2=0
cc_592 N_TE_B_c_675_n N_A_28_368#_c_914_n 0.0105001f $X=6.81 $Y=1.765 $X2=0
+ $Y2=0
cc_593 N_TE_B_c_677_n N_A_28_368#_c_915_n 0.0114786f $X=7.26 $Y=1.765 $X2=0
+ $Y2=0
cc_594 N_TE_B_c_679_n N_A_28_368#_c_915_n 0.0101684f $X=7.88 $Y=1.765 $X2=0
+ $Y2=0
cc_595 N_TE_B_c_664_n N_A_28_368#_c_886_n 5.73918e-19 $X=4.26 $Y=1.765 $X2=0
+ $Y2=0
cc_596 N_TE_B_c_667_n N_A_28_368#_c_886_n 0.00650056f $X=4.81 $Y=1.765 $X2=0
+ $Y2=0
cc_597 N_TE_B_c_669_n N_A_28_368#_c_886_n 0.00650056f $X=5.26 $Y=1.765 $X2=0
+ $Y2=0
cc_598 N_TE_B_c_671_n N_A_28_368#_c_886_n 5.73918e-19 $X=5.81 $Y=1.765 $X2=0
+ $Y2=0
cc_599 N_TE_B_c_669_n N_A_28_368#_c_887_n 5.73918e-19 $X=5.26 $Y=1.765 $X2=0
+ $Y2=0
cc_600 N_TE_B_c_671_n N_A_28_368#_c_887_n 0.00650056f $X=5.81 $Y=1.765 $X2=0
+ $Y2=0
cc_601 N_TE_B_c_673_n N_A_28_368#_c_887_n 0.00650056f $X=6.26 $Y=1.765 $X2=0
+ $Y2=0
cc_602 N_TE_B_c_675_n N_A_28_368#_c_887_n 5.73918e-19 $X=6.81 $Y=1.765 $X2=0
+ $Y2=0
cc_603 N_TE_B_c_673_n N_A_28_368#_c_888_n 6.55446e-19 $X=6.26 $Y=1.765 $X2=0
+ $Y2=0
cc_604 N_TE_B_c_675_n N_A_28_368#_c_888_n 0.00702028f $X=6.81 $Y=1.765 $X2=0
+ $Y2=0
cc_605 N_TE_B_c_677_n N_A_28_368#_c_888_n 0.00910693f $X=7.26 $Y=1.765 $X2=0
+ $Y2=0
cc_606 N_TE_B_c_679_n N_A_28_368#_c_888_n 0.0015865f $X=7.88 $Y=1.765 $X2=0
+ $Y2=0
cc_607 N_TE_B_c_677_n N_A_28_368#_c_889_n 8.39036e-19 $X=7.26 $Y=1.765 $X2=0
+ $Y2=0
cc_608 N_TE_B_c_679_n N_A_28_368#_c_889_n 0.00608649f $X=7.88 $Y=1.765 $X2=0
+ $Y2=0
cc_609 N_TE_B_c_664_n N_VPWR_c_1149_n 0.00285025f $X=4.26 $Y=1.765 $X2=0 $Y2=0
cc_610 N_TE_B_c_667_n N_VPWR_c_1149_n 0.00336706f $X=4.81 $Y=1.765 $X2=0 $Y2=0
cc_611 N_TE_B_c_669_n N_VPWR_c_1150_n 0.00336706f $X=5.26 $Y=1.765 $X2=0 $Y2=0
cc_612 N_TE_B_c_671_n N_VPWR_c_1150_n 0.00336706f $X=5.81 $Y=1.765 $X2=0 $Y2=0
cc_613 N_TE_B_c_673_n N_VPWR_c_1151_n 0.00336706f $X=6.26 $Y=1.765 $X2=0 $Y2=0
cc_614 N_TE_B_c_675_n N_VPWR_c_1151_n 0.00475521f $X=6.81 $Y=1.765 $X2=0 $Y2=0
cc_615 N_TE_B_c_675_n N_VPWR_c_1152_n 0.00445602f $X=6.81 $Y=1.765 $X2=0 $Y2=0
cc_616 N_TE_B_c_677_n N_VPWR_c_1152_n 0.00320415f $X=7.26 $Y=1.765 $X2=0 $Y2=0
cc_617 N_TE_B_c_677_n N_VPWR_c_1153_n 0.00394942f $X=7.26 $Y=1.765 $X2=0 $Y2=0
cc_618 N_TE_B_c_679_n N_VPWR_c_1153_n 0.00394942f $X=7.88 $Y=1.765 $X2=0 $Y2=0
cc_619 N_TE_B_c_682_n N_VPWR_c_1154_n 0.0250504f $X=9.105 $Y=1.765 $X2=0 $Y2=0
cc_620 N_TE_B_c_664_n N_VPWR_c_1157_n 0.0044313f $X=4.26 $Y=1.765 $X2=0 $Y2=0
cc_621 N_TE_B_c_667_n N_VPWR_c_1158_n 0.00445602f $X=4.81 $Y=1.765 $X2=0 $Y2=0
cc_622 N_TE_B_c_669_n N_VPWR_c_1158_n 0.00445602f $X=5.26 $Y=1.765 $X2=0 $Y2=0
cc_623 N_TE_B_c_671_n N_VPWR_c_1159_n 0.00445602f $X=5.81 $Y=1.765 $X2=0 $Y2=0
cc_624 N_TE_B_c_673_n N_VPWR_c_1159_n 0.00445602f $X=6.26 $Y=1.765 $X2=0 $Y2=0
cc_625 N_TE_B_c_679_n N_VPWR_c_1160_n 0.00320415f $X=7.88 $Y=1.765 $X2=0 $Y2=0
cc_626 N_TE_B_c_682_n N_VPWR_c_1160_n 0.00413917f $X=9.105 $Y=1.765 $X2=0 $Y2=0
cc_627 N_TE_B_c_664_n N_VPWR_c_1148_n 0.00437782f $X=4.26 $Y=1.765 $X2=0 $Y2=0
cc_628 N_TE_B_c_667_n N_VPWR_c_1148_n 0.00437179f $X=4.81 $Y=1.765 $X2=0 $Y2=0
cc_629 N_TE_B_c_669_n N_VPWR_c_1148_n 0.00437179f $X=5.26 $Y=1.765 $X2=0 $Y2=0
cc_630 N_TE_B_c_671_n N_VPWR_c_1148_n 0.00437179f $X=5.81 $Y=1.765 $X2=0 $Y2=0
cc_631 N_TE_B_c_673_n N_VPWR_c_1148_n 0.00437179f $X=6.26 $Y=1.765 $X2=0 $Y2=0
cc_632 N_TE_B_c_675_n N_VPWR_c_1148_n 0.00437179f $X=6.81 $Y=1.765 $X2=0 $Y2=0
cc_633 N_TE_B_c_677_n N_VPWR_c_1148_n 0.00400928f $X=7.26 $Y=1.765 $X2=0 $Y2=0
cc_634 N_TE_B_c_679_n N_VPWR_c_1148_n 0.00405729f $X=7.88 $Y=1.765 $X2=0 $Y2=0
cc_635 N_TE_B_c_682_n N_VPWR_c_1148_n 0.00822528f $X=9.105 $Y=1.765 $X2=0 $Y2=0
cc_636 N_TE_B_c_644_n N_A_27_74#_c_1284_n 0.00363845f $X=4.335 $Y=1.69 $X2=0
+ $Y2=0
cc_637 N_TE_B_c_645_n N_A_27_74#_c_1287_n 0.00587659f $X=5.185 $Y=1.69 $X2=0
+ $Y2=0
cc_638 N_TE_B_c_656_n N_A_27_74#_c_1289_n 0.00689812f $X=5.81 $Y=1.69 $X2=0
+ $Y2=0
cc_639 N_TE_B_c_648_n N_A_27_74#_c_1291_n 0.00692076f $X=6.735 $Y=1.69 $X2=0
+ $Y2=0
cc_640 N_TE_B_c_659_n N_A_27_74#_c_1291_n 0.00338859f $X=7.26 $Y=1.69 $X2=0
+ $Y2=0
cc_641 N_TE_B_c_643_n N_A_27_74#_c_1296_n 0.00445864f $X=4.735 $Y=1.69 $X2=0
+ $Y2=0
cc_642 N_TE_B_c_646_n N_A_27_74#_c_1297_n 0.00347932f $X=5.735 $Y=1.69 $X2=0
+ $Y2=0
cc_643 N_TE_B_c_648_n N_A_27_74#_c_1298_n 0.00327264f $X=6.735 $Y=1.69 $X2=0
+ $Y2=0
cc_644 N_TE_B_c_653_n N_VGND_c_1446_n 0.00259633f $X=9.2 $Y=1.22 $X2=0 $Y2=0
cc_645 TE_B N_VGND_c_1446_n 0.0125437f $X=9.275 $Y=1.21 $X2=0 $Y2=0
cc_646 N_TE_B_c_653_n N_VGND_c_1456_n 0.00432935f $X=9.2 $Y=1.22 $X2=0 $Y2=0
cc_647 N_TE_B_c_653_n N_VGND_c_1460_n 0.00821561f $X=9.2 $Y=1.22 $X2=0 $Y2=0
cc_648 N_A_c_831_n N_VPWR_c_1154_n 0.00398037f $X=9.605 $Y=1.765 $X2=0 $Y2=0
cc_649 N_A_c_831_n N_VPWR_c_1156_n 6.04028e-19 $X=9.605 $Y=1.765 $X2=0 $Y2=0
cc_650 N_A_c_832_n N_VPWR_c_1156_n 0.0137742f $X=10.055 $Y=1.765 $X2=0 $Y2=0
cc_651 N_A_c_831_n N_VPWR_c_1161_n 0.00445602f $X=9.605 $Y=1.765 $X2=0 $Y2=0
cc_652 N_A_c_832_n N_VPWR_c_1161_n 0.00413917f $X=10.055 $Y=1.765 $X2=0 $Y2=0
cc_653 N_A_c_831_n N_VPWR_c_1148_n 0.00857432f $X=9.605 $Y=1.765 $X2=0 $Y2=0
cc_654 N_A_c_832_n N_VPWR_c_1148_n 0.00817726f $X=10.055 $Y=1.765 $X2=0 $Y2=0
cc_655 N_A_c_827_n N_VGND_c_1446_n 0.00144568f $X=9.63 $Y=1.22 $X2=0 $Y2=0
cc_656 N_A_c_827_n N_VGND_c_1448_n 3.97405e-19 $X=9.63 $Y=1.22 $X2=0 $Y2=0
cc_657 N_A_c_828_n N_VGND_c_1448_n 0.00805371f $X=10.06 $Y=1.22 $X2=0 $Y2=0
cc_658 N_A_c_827_n N_VGND_c_1457_n 0.00434054f $X=9.63 $Y=1.22 $X2=0 $Y2=0
cc_659 N_A_c_828_n N_VGND_c_1457_n 0.00383152f $X=10.06 $Y=1.22 $X2=0 $Y2=0
cc_660 N_A_c_827_n N_VGND_c_1460_n 0.00820221f $X=9.63 $Y=1.22 $X2=0 $Y2=0
cc_661 N_A_c_828_n N_VGND_c_1460_n 0.00383967f $X=10.06 $Y=1.22 $X2=0 $Y2=0
cc_662 N_A_28_368#_c_878_n N_Z_M1006_s 0.00197722f $X=1.085 $Y=2.99 $X2=0 $Y2=0
cc_663 N_A_28_368#_c_880_n N_Z_M1013_s 0.00250873f $X=2.05 $Y=2.99 $X2=0 $Y2=0
cc_664 N_A_28_368#_c_881_n N_Z_M1015_s 0.00197722f $X=2.92 $Y=2.99 $X2=0 $Y2=0
cc_665 N_A_28_368#_c_882_n N_Z_M1019_s 0.00234927f $X=3.87 $Y=2.99 $X2=0 $Y2=0
cc_666 N_A_28_368#_c_877_n N_Z_c_1030_n 0.0556321f $X=0.285 $Y=1.985 $X2=0 $Y2=0
cc_667 N_A_28_368#_c_878_n N_Z_c_1030_n 0.017859f $X=1.085 $Y=2.99 $X2=0 $Y2=0
cc_668 N_A_28_368#_M1010_d N_Z_c_1022_n 0.00197722f $X=1.035 $Y=1.84 $X2=0 $Y2=0
cc_669 N_A_28_368#_c_900_n N_Z_c_1022_n 0.016157f $X=1.185 $Y=2.325 $X2=0 $Y2=0
cc_670 N_A_28_368#_c_880_n N_Z_c_1045_n 0.018923f $X=2.05 $Y=2.99 $X2=0 $Y2=0
cc_671 N_A_28_368#_c_904_n N_Z_c_1045_n 0.0374537f $X=2.135 $Y=2.325 $X2=0 $Y2=0
cc_672 N_A_28_368#_M1014_d N_Z_c_1023_n 0.00247267f $X=1.985 $Y=1.84 $X2=0 $Y2=0
cc_673 N_A_28_368#_c_904_n N_Z_c_1023_n 0.0136682f $X=2.135 $Y=2.325 $X2=0 $Y2=0
cc_674 N_A_28_368#_c_904_n N_Z_c_1055_n 0.0374537f $X=2.135 $Y=2.325 $X2=0 $Y2=0
cc_675 N_A_28_368#_c_881_n N_Z_c_1055_n 0.0160777f $X=2.92 $Y=2.99 $X2=0 $Y2=0
cc_676 N_A_28_368#_M1017_d N_Z_c_1024_n 0.00250873f $X=2.885 $Y=1.84 $X2=0 $Y2=0
cc_677 N_A_28_368#_c_966_p N_Z_c_1024_n 0.0192006f $X=3.085 $Y=2.325 $X2=0 $Y2=0
cc_678 N_A_28_368#_c_882_n N_Z_c_1075_n 0.0177813f $X=3.87 $Y=2.99 $X2=0 $Y2=0
cc_679 N_A_28_368#_c_877_n N_Z_c_1026_n 0.0134523f $X=0.285 $Y=1.985 $X2=0 $Y2=0
cc_680 N_A_28_368#_c_912_n N_VPWR_M1016_s 0.00621236f $X=4.87 $Y=2.475 $X2=-0.19
+ $Y2=1.66
cc_681 N_A_28_368#_c_913_n N_VPWR_M1022_s 0.00621236f $X=5.87 $Y=2.475 $X2=0
+ $Y2=0
cc_682 N_A_28_368#_c_914_n N_VPWR_M1024_s 0.00621236f $X=6.87 $Y=2.475 $X2=0
+ $Y2=0
cc_683 N_A_28_368#_c_915_n N_VPWR_M1028_s 0.00935184f $X=7.94 $Y=2.645 $X2=0
+ $Y2=0
cc_684 N_A_28_368#_c_882_n N_VPWR_c_1149_n 0.0119239f $X=3.87 $Y=2.99 $X2=0
+ $Y2=0
cc_685 N_A_28_368#_c_912_n N_VPWR_c_1149_n 0.0226192f $X=4.87 $Y=2.475 $X2=0
+ $Y2=0
cc_686 N_A_28_368#_c_886_n N_VPWR_c_1149_n 0.0101711f $X=5.035 $Y=2.475 $X2=0
+ $Y2=0
cc_687 N_A_28_368#_c_913_n N_VPWR_c_1150_n 0.0226192f $X=5.87 $Y=2.475 $X2=0
+ $Y2=0
cc_688 N_A_28_368#_c_886_n N_VPWR_c_1150_n 0.0101711f $X=5.035 $Y=2.475 $X2=0
+ $Y2=0
cc_689 N_A_28_368#_c_887_n N_VPWR_c_1150_n 0.0101711f $X=6.035 $Y=2.475 $X2=0
+ $Y2=0
cc_690 N_A_28_368#_c_914_n N_VPWR_c_1151_n 0.0226192f $X=6.87 $Y=2.475 $X2=0
+ $Y2=0
cc_691 N_A_28_368#_c_887_n N_VPWR_c_1151_n 0.0101711f $X=6.035 $Y=2.475 $X2=0
+ $Y2=0
cc_692 N_A_28_368#_c_888_n N_VPWR_c_1151_n 0.0101711f $X=7.035 $Y=2.475 $X2=0
+ $Y2=0
cc_693 N_A_28_368#_c_915_n N_VPWR_c_1152_n 0.0032422f $X=7.94 $Y=2.645 $X2=0
+ $Y2=0
cc_694 N_A_28_368#_c_888_n N_VPWR_c_1152_n 0.0144033f $X=7.035 $Y=2.475 $X2=0
+ $Y2=0
cc_695 N_A_28_368#_c_915_n N_VPWR_c_1153_n 0.0247191f $X=7.94 $Y=2.645 $X2=0
+ $Y2=0
cc_696 N_A_28_368#_c_888_n N_VPWR_c_1153_n 0.00540816f $X=7.035 $Y=2.475 $X2=0
+ $Y2=0
cc_697 N_A_28_368#_c_889_n N_VPWR_c_1153_n 0.00540816f $X=8.105 $Y=2.645 $X2=0
+ $Y2=0
cc_698 N_A_28_368#_c_878_n N_VPWR_c_1157_n 0.0451275f $X=1.085 $Y=2.99 $X2=0
+ $Y2=0
cc_699 N_A_28_368#_c_879_n N_VPWR_c_1157_n 0.0179217f $X=0.37 $Y=2.99 $X2=0
+ $Y2=0
cc_700 N_A_28_368#_c_880_n N_VPWR_c_1157_n 0.0442078f $X=2.05 $Y=2.99 $X2=0
+ $Y2=0
cc_701 N_A_28_368#_c_881_n N_VPWR_c_1157_n 0.0441612f $X=2.92 $Y=2.99 $X2=0
+ $Y2=0
cc_702 N_A_28_368#_c_882_n N_VPWR_c_1157_n 0.0664928f $X=3.87 $Y=2.99 $X2=0
+ $Y2=0
cc_703 N_A_28_368#_c_883_n N_VPWR_c_1157_n 0.0189443f $X=1.217 $Y=2.99 $X2=0
+ $Y2=0
cc_704 N_A_28_368#_c_884_n N_VPWR_c_1157_n 0.0121867f $X=2.135 $Y=2.99 $X2=0
+ $Y2=0
cc_705 N_A_28_368#_c_885_n N_VPWR_c_1157_n 0.0193554f $X=3.055 $Y=2.99 $X2=0
+ $Y2=0
cc_706 N_A_28_368#_c_886_n N_VPWR_c_1158_n 0.0144033f $X=5.035 $Y=2.475 $X2=0
+ $Y2=0
cc_707 N_A_28_368#_c_887_n N_VPWR_c_1159_n 0.0144033f $X=6.035 $Y=2.475 $X2=0
+ $Y2=0
cc_708 N_A_28_368#_c_915_n N_VPWR_c_1160_n 0.0032422f $X=7.94 $Y=2.645 $X2=0
+ $Y2=0
cc_709 N_A_28_368#_c_889_n N_VPWR_c_1160_n 0.0140991f $X=8.105 $Y=2.645 $X2=0
+ $Y2=0
cc_710 N_A_28_368#_c_878_n N_VPWR_c_1148_n 0.0255092f $X=1.085 $Y=2.99 $X2=0
+ $Y2=0
cc_711 N_A_28_368#_c_879_n N_VPWR_c_1148_n 0.00971942f $X=0.37 $Y=2.99 $X2=0
+ $Y2=0
cc_712 N_A_28_368#_c_880_n N_VPWR_c_1148_n 0.0250141f $X=2.05 $Y=2.99 $X2=0
+ $Y2=0
cc_713 N_A_28_368#_c_881_n N_VPWR_c_1148_n 0.0249452f $X=2.92 $Y=2.99 $X2=0
+ $Y2=0
cc_714 N_A_28_368#_c_882_n N_VPWR_c_1148_n 0.0369573f $X=3.87 $Y=2.99 $X2=0
+ $Y2=0
cc_715 N_A_28_368#_c_912_n N_VPWR_c_1148_n 0.0117498f $X=4.87 $Y=2.475 $X2=0
+ $Y2=0
cc_716 N_A_28_368#_c_913_n N_VPWR_c_1148_n 0.0117498f $X=5.87 $Y=2.475 $X2=0
+ $Y2=0
cc_717 N_A_28_368#_c_914_n N_VPWR_c_1148_n 0.0117628f $X=6.87 $Y=2.475 $X2=0
+ $Y2=0
cc_718 N_A_28_368#_c_915_n N_VPWR_c_1148_n 0.0123416f $X=7.94 $Y=2.645 $X2=0
+ $Y2=0
cc_719 N_A_28_368#_c_883_n N_VPWR_c_1148_n 0.010234f $X=1.217 $Y=2.99 $X2=0
+ $Y2=0
cc_720 N_A_28_368#_c_884_n N_VPWR_c_1148_n 0.00660921f $X=2.135 $Y=2.99 $X2=0
+ $Y2=0
cc_721 N_A_28_368#_c_885_n N_VPWR_c_1148_n 0.010497f $X=3.055 $Y=2.99 $X2=0
+ $Y2=0
cc_722 N_A_28_368#_c_886_n N_VPWR_c_1148_n 0.0119211f $X=5.035 $Y=2.475 $X2=0
+ $Y2=0
cc_723 N_A_28_368#_c_887_n N_VPWR_c_1148_n 0.0119211f $X=6.035 $Y=2.475 $X2=0
+ $Y2=0
cc_724 N_A_28_368#_c_888_n N_VPWR_c_1148_n 0.0119211f $X=7.035 $Y=2.475 $X2=0
+ $Y2=0
cc_725 N_A_28_368#_c_889_n N_VPWR_c_1148_n 0.0118561f $X=8.105 $Y=2.645 $X2=0
+ $Y2=0
cc_726 N_Z_c_1015_n N_A_27_74#_M1009_d 0.00221449f $X=1.43 $Y=1.065 $X2=0 $Y2=0
cc_727 N_Z_c_1016_n N_A_27_74#_M1029_d 0.00250873f $X=2.43 $Y=1.065 $X2=0 $Y2=0
cc_728 N_Z_c_1017_n N_A_27_74#_M1033_d 0.00270388f $X=3.43 $Y=1.065 $X2=0 $Y2=0
cc_729 Z N_A_27_74#_c_1277_n 0.00676472f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_730 N_Z_M1005_s N_A_27_74#_c_1278_n 0.00176461f $X=0.57 $Y=0.37 $X2=0 $Y2=0
cc_731 N_Z_c_1015_n N_A_27_74#_c_1278_n 0.00319222f $X=1.43 $Y=1.065 $X2=0 $Y2=0
cc_732 N_Z_c_1103_n N_A_27_74#_c_1278_n 0.0159544f $X=0.71 $Y=0.76 $X2=0 $Y2=0
cc_733 N_Z_c_1015_n N_A_27_74#_c_1302_n 0.0133644f $X=1.43 $Y=1.065 $X2=0 $Y2=0
cc_734 N_Z_c_1041_n N_A_27_74#_c_1302_n 0.0137413f $X=1.595 $Y=0.76 $X2=0 $Y2=0
cc_735 N_Z_M1011_s N_A_27_74#_c_1280_n 0.00176461f $X=1.455 $Y=0.37 $X2=0 $Y2=0
cc_736 N_Z_c_1015_n N_A_27_74#_c_1280_n 0.00386975f $X=1.43 $Y=1.065 $X2=0 $Y2=0
cc_737 N_Z_c_1041_n N_A_27_74#_c_1280_n 0.0157331f $X=1.595 $Y=0.76 $X2=0 $Y2=0
cc_738 N_Z_c_1016_n N_A_27_74#_c_1280_n 0.00319222f $X=2.43 $Y=1.065 $X2=0 $Y2=0
cc_739 N_Z_c_1016_n N_A_27_74#_c_1305_n 0.0206429f $X=2.43 $Y=1.065 $X2=0 $Y2=0
cc_740 N_Z_M1032_s N_A_27_74#_c_1281_n 0.00250873f $X=2.385 $Y=0.37 $X2=0 $Y2=0
cc_741 N_Z_c_1016_n N_A_27_74#_c_1281_n 0.00319222f $X=2.43 $Y=1.065 $X2=0 $Y2=0
cc_742 N_Z_c_1059_n N_A_27_74#_c_1281_n 0.0193319f $X=2.595 $Y=0.76 $X2=0 $Y2=0
cc_743 N_Z_c_1017_n N_A_27_74#_c_1281_n 0.00319222f $X=3.43 $Y=1.065 $X2=0 $Y2=0
cc_744 N_Z_c_1017_n N_A_27_74#_c_1309_n 0.0207199f $X=3.43 $Y=1.065 $X2=0 $Y2=0
cc_745 N_Z_M1034_s N_A_27_74#_c_1282_n 0.00234927f $X=3.4 $Y=0.37 $X2=0 $Y2=0
cc_746 N_Z_c_1017_n N_A_27_74#_c_1282_n 0.00357683f $X=3.43 $Y=1.065 $X2=0 $Y2=0
cc_747 N_Z_c_1077_n N_A_27_74#_c_1282_n 0.0182078f $X=3.595 $Y=0.76 $X2=0 $Y2=0
cc_748 N_Z_c_1017_n N_A_27_74#_c_1283_n 0.00745191f $X=3.43 $Y=1.065 $X2=0 $Y2=0
cc_749 N_Z_c_1017_n N_A_27_74#_c_1285_n 8.53482e-19 $X=3.43 $Y=1.065 $X2=0 $Y2=0
cc_750 N_A_27_74#_c_1282_n N_VGND_c_1442_n 0.0112234f $X=3.94 $Y=0.34 $X2=0
+ $Y2=0
cc_751 N_A_27_74#_c_1284_n N_VGND_c_1442_n 0.0216086f $X=4.72 $Y=1.225 $X2=0
+ $Y2=0
cc_752 N_A_27_74#_c_1286_n N_VGND_c_1442_n 0.0229496f $X=4.885 $Y=0.515 $X2=0
+ $Y2=0
cc_753 N_A_27_74#_c_1286_n N_VGND_c_1443_n 0.0281649f $X=4.885 $Y=0.515 $X2=0
+ $Y2=0
cc_754 N_A_27_74#_c_1287_n N_VGND_c_1443_n 0.0135549f $X=5.58 $Y=1.385 $X2=0
+ $Y2=0
cc_755 N_A_27_74#_c_1288_n N_VGND_c_1443_n 0.0281649f $X=5.745 $Y=0.515 $X2=0
+ $Y2=0
cc_756 N_A_27_74#_c_1288_n N_VGND_c_1444_n 0.0282477f $X=5.745 $Y=0.515 $X2=0
+ $Y2=0
cc_757 N_A_27_74#_c_1289_n N_VGND_c_1444_n 0.0198685f $X=6.44 $Y=1.385 $X2=0
+ $Y2=0
cc_758 N_A_27_74#_c_1290_n N_VGND_c_1444_n 0.0282477f $X=6.605 $Y=0.515 $X2=0
+ $Y2=0
cc_759 N_A_27_74#_c_1290_n N_VGND_c_1445_n 0.0282477f $X=6.605 $Y=0.515 $X2=0
+ $Y2=0
cc_760 N_A_27_74#_c_1291_n N_VGND_c_1445_n 0.0198685f $X=7.3 $Y=1.385 $X2=0
+ $Y2=0
cc_761 N_A_27_74#_c_1292_n N_VGND_c_1445_n 0.0282477f $X=7.465 $Y=0.515 $X2=0
+ $Y2=0
cc_762 N_A_27_74#_c_1278_n N_VGND_c_1449_n 0.043517f $X=1.055 $Y=0.34 $X2=0
+ $Y2=0
cc_763 N_A_27_74#_c_1279_n N_VGND_c_1449_n 0.0179217f $X=0.365 $Y=0.34 $X2=0
+ $Y2=0
cc_764 N_A_27_74#_c_1280_n N_VGND_c_1449_n 0.0444833f $X=1.93 $Y=0.34 $X2=0
+ $Y2=0
cc_765 N_A_27_74#_c_1281_n N_VGND_c_1449_n 0.0423044f $X=2.93 $Y=0.34 $X2=0
+ $Y2=0
cc_766 N_A_27_74#_c_1282_n N_VGND_c_1449_n 0.0550916f $X=3.94 $Y=0.34 $X2=0
+ $Y2=0
cc_767 N_A_27_74#_c_1293_n N_VGND_c_1449_n 0.0120038f $X=1.14 $Y=0.34 $X2=0
+ $Y2=0
cc_768 N_A_27_74#_c_1294_n N_VGND_c_1449_n 0.0232138f $X=2.095 $Y=0.34 $X2=0
+ $Y2=0
cc_769 N_A_27_74#_c_1295_n N_VGND_c_1449_n 0.0232651f $X=3.095 $Y=0.34 $X2=0
+ $Y2=0
cc_770 N_A_27_74#_c_1286_n N_VGND_c_1451_n 0.0109942f $X=4.885 $Y=0.515 $X2=0
+ $Y2=0
cc_771 N_A_27_74#_c_1288_n N_VGND_c_1453_n 0.0109942f $X=5.745 $Y=0.515 $X2=0
+ $Y2=0
cc_772 N_A_27_74#_c_1290_n N_VGND_c_1455_n 0.0109942f $X=6.605 $Y=0.515 $X2=0
+ $Y2=0
cc_773 N_A_27_74#_c_1292_n N_VGND_c_1456_n 0.0109942f $X=7.465 $Y=0.515 $X2=0
+ $Y2=0
cc_774 N_A_27_74#_c_1278_n N_VGND_c_1460_n 0.0245693f $X=1.055 $Y=0.34 $X2=0
+ $Y2=0
cc_775 N_A_27_74#_c_1279_n N_VGND_c_1460_n 0.00971942f $X=0.365 $Y=0.34 $X2=0
+ $Y2=0
cc_776 N_A_27_74#_c_1280_n N_VGND_c_1460_n 0.0251332f $X=1.93 $Y=0.34 $X2=0
+ $Y2=0
cc_777 N_A_27_74#_c_1281_n N_VGND_c_1460_n 0.0239316f $X=2.93 $Y=0.34 $X2=0
+ $Y2=0
cc_778 N_A_27_74#_c_1282_n N_VGND_c_1460_n 0.0308486f $X=3.94 $Y=0.34 $X2=0
+ $Y2=0
cc_779 N_A_27_74#_c_1286_n N_VGND_c_1460_n 0.00904371f $X=4.885 $Y=0.515 $X2=0
+ $Y2=0
cc_780 N_A_27_74#_c_1288_n N_VGND_c_1460_n 0.00904371f $X=5.745 $Y=0.515 $X2=0
+ $Y2=0
cc_781 N_A_27_74#_c_1290_n N_VGND_c_1460_n 0.00904371f $X=6.605 $Y=0.515 $X2=0
+ $Y2=0
cc_782 N_A_27_74#_c_1292_n N_VGND_c_1460_n 0.00904371f $X=7.465 $Y=0.515 $X2=0
+ $Y2=0
cc_783 N_A_27_74#_c_1293_n N_VGND_c_1460_n 0.00657483f $X=1.14 $Y=0.34 $X2=0
+ $Y2=0
cc_784 N_A_27_74#_c_1294_n N_VGND_c_1460_n 0.0126482f $X=2.095 $Y=0.34 $X2=0
+ $Y2=0
cc_785 N_A_27_74#_c_1295_n N_VGND_c_1460_n 0.0127168f $X=3.095 $Y=0.34 $X2=0
+ $Y2=0
