* File: sky130_fd_sc_hs__o32a_4.pex.spice
* Created: Tue Sep  1 20:18:45 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HS__O32A_4%A_83_256# 1 2 3 4 14 15 17 20 22 25 26 28 31
+ 33 35 38 40 42 45 47 48 55 56 58 59 62 64 68 72 74
c173 74 0 1.29542e-19 $X=2.27 $Y=1.195
c174 64 0 6.51508e-20 $X=4.23 $Y=1.015
c175 59 0 7.30872e-20 $X=3.395 $Y=1.92
c176 40 0 7.44774e-20 $X=2.025 $Y=1.765
c177 31 0 8.40338e-20 $X=1.065 $Y=0.74
c178 25 0 1.0009e-19 $X=0.955 $Y=1.675
c179 15 0 3.73162e-20 $X=0.505 $Y=1.765
r180 86 87 58.9279 $w=3.19e-07 $l=3.9e-07 $layer=POLY_cond $X=1.635 $Y=1.522
+ $X2=2.025 $Y2=1.522
r181 85 86 27.1975 $w=3.19e-07 $l=1.8e-07 $layer=POLY_cond $X=1.455 $Y=1.522
+ $X2=1.635 $Y2=1.522
r182 78 79 7.46939 $w=2.94e-07 $l=1.8e-07 $layer=LI1_cond $X=3.395 $Y=1.015
+ $X2=3.395 $Y2=1.195
r183 70 72 4.1907 $w=3.28e-07 $l=1.2e-07 $layer=LI1_cond $X=4.395 $Y=0.93
+ $X2=4.395 $Y2=0.81
r184 66 81 4.74481 $w=1.7e-07 $l=1.96415e-07 $layer=LI1_cond $X=3.575 $Y=2.105
+ $X2=3.402 $Y2=2.055
r185 66 68 119.064 $w=1.68e-07 $l=1.825e-06 $layer=LI1_cond $X=3.575 $Y=2.105
+ $X2=5.4 $Y2=2.105
r186 65 78 3.94234 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.56 $Y=1.015
+ $X2=3.395 $Y2=1.015
r187 64 70 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.23 $Y=1.015
+ $X2=4.395 $Y2=0.93
r188 64 65 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.23 $Y=1.015
+ $X2=3.56 $Y2=1.015
r189 60 78 3.72042 $w=2.94e-07 $l=1.00995e-07 $layer=LI1_cond $X=3.43 $Y=0.93
+ $X2=3.395 $Y2=1.015
r190 60 62 5.31897 $w=2.58e-07 $l=1.2e-07 $layer=LI1_cond $X=3.43 $Y=0.93
+ $X2=3.43 $Y2=0.81
r191 59 81 3.02136 $w=3.3e-07 $l=1.38456e-07 $layer=LI1_cond $X=3.395 $Y=1.92
+ $X2=3.402 $Y2=2.055
r192 58 79 3.3163 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.395 $Y=1.28
+ $X2=3.395 $Y2=1.195
r193 58 59 22.3504 $w=3.28e-07 $l=6.4e-07 $layer=LI1_cond $X=3.395 $Y=1.28
+ $X2=3.395 $Y2=1.92
r194 57 74 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.355 $Y=1.195
+ $X2=2.27 $Y2=1.195
r195 56 79 3.94234 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.23 $Y=1.195
+ $X2=3.395 $Y2=1.195
r196 56 57 57.0856 $w=1.68e-07 $l=8.75e-07 $layer=LI1_cond $X=3.23 $Y=1.195
+ $X2=2.355 $Y2=1.195
r197 55 89 13.5987 $w=3.19e-07 $l=9e-08 $layer=POLY_cond $X=2.1 $Y=1.522
+ $X2=2.19 $Y2=1.522
r198 55 87 11.3323 $w=3.19e-07 $l=7.5e-08 $layer=POLY_cond $X=2.1 $Y=1.522
+ $X2=2.025 $Y2=1.522
r199 54 55 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=2.1
+ $Y=1.445 $X2=2.1 $Y2=1.445
r200 51 85 5.2884 $w=3.19e-07 $l=3.5e-08 $layer=POLY_cond $X=1.42 $Y=1.522
+ $X2=1.455 $Y2=1.522
r201 50 54 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=1.42 $Y=1.445
+ $X2=2.1 $Y2=1.445
r202 50 51 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.42
+ $Y=1.445 $X2=1.42 $Y2=1.445
r203 48 74 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=2.27 $Y=1.445
+ $X2=2.27 $Y2=1.195
r204 48 54 2.96841 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=2.185 $Y=1.445
+ $X2=2.1 $Y2=1.445
r205 43 89 20.418 $w=1.5e-07 $l=2.42e-07 $layer=POLY_cond $X=2.19 $Y=1.28
+ $X2=2.19 $Y2=1.522
r206 43 45 276.894 $w=1.5e-07 $l=5.4e-07 $layer=POLY_cond $X=2.19 $Y=1.28
+ $X2=2.19 $Y2=0.74
r207 40 87 20.418 $w=1.5e-07 $l=2.43e-07 $layer=POLY_cond $X=2.025 $Y=1.765
+ $X2=2.025 $Y2=1.522
r208 40 42 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.025 $Y=1.765
+ $X2=2.025 $Y2=2.4
r209 36 86 20.418 $w=1.5e-07 $l=2.42e-07 $layer=POLY_cond $X=1.635 $Y=1.28
+ $X2=1.635 $Y2=1.522
r210 36 38 276.894 $w=1.5e-07 $l=5.4e-07 $layer=POLY_cond $X=1.635 $Y=1.28
+ $X2=1.635 $Y2=0.74
r211 33 85 20.418 $w=1.5e-07 $l=2.43e-07 $layer=POLY_cond $X=1.455 $Y=1.765
+ $X2=1.455 $Y2=1.522
r212 33 35 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.455 $Y=1.765
+ $X2=1.455 $Y2=2.4
r213 29 51 53.6395 $w=3.19e-07 $l=4.60364e-07 $layer=POLY_cond $X=1.065 $Y=1.28
+ $X2=1.42 $Y2=1.522
r214 29 31 276.894 $w=1.5e-07 $l=5.4e-07 $layer=POLY_cond $X=1.065 $Y=1.28
+ $X2=1.065 $Y2=0.74
r215 26 28 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.955 $Y=1.765
+ $X2=0.955 $Y2=2.4
r216 25 26 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=0.955 $Y=1.675
+ $X2=0.955 $Y2=1.765
r217 24 29 16.6207 $w=3.19e-07 $l=1.97484e-07 $layer=POLY_cond $X=0.955 $Y=1.43
+ $X2=1.065 $Y2=1.28
r218 24 25 95.2339 $w=1.8e-07 $l=2.45e-07 $layer=POLY_cond $X=0.955 $Y=1.43
+ $X2=0.955 $Y2=1.675
r219 23 47 6.66866 $w=1.5e-07 $l=1.48e-07 $layer=POLY_cond $X=0.71 $Y=1.355
+ $X2=0.562 $Y2=1.355
r220 22 24 27.2139 $w=3.19e-07 $l=1.21861e-07 $layer=POLY_cond $X=0.865 $Y=1.355
+ $X2=0.955 $Y2=1.43
r221 22 23 79.4787 $w=1.5e-07 $l=1.55e-07 $layer=POLY_cond $X=0.865 $Y=1.355
+ $X2=0.71 $Y2=1.355
r222 18 47 18.8402 $w=1.65e-07 $l=1.05357e-07 $layer=POLY_cond $X=0.635 $Y=1.28
+ $X2=0.562 $Y2=1.355
r223 18 20 276.894 $w=1.5e-07 $l=5.4e-07 $layer=POLY_cond $X=0.635 $Y=1.28
+ $X2=0.635 $Y2=0.74
r224 15 17 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.505 $Y=1.765
+ $X2=0.505 $Y2=2.4
r225 14 15 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=0.505 $Y=1.675
+ $X2=0.505 $Y2=1.765
r226 13 47 18.8402 $w=1.65e-07 $l=9.94987e-08 $layer=POLY_cond $X=0.505 $Y=1.43
+ $X2=0.562 $Y2=1.355
r227 13 14 95.2339 $w=1.8e-07 $l=2.45e-07 $layer=POLY_cond $X=0.505 $Y=1.43
+ $X2=0.505 $Y2=1.675
r228 4 68 600 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=5.25
+ $Y=1.96 $X2=5.4 $Y2=2.105
r229 3 81 600 $w=1.7e-07 $l=2.17428e-07 $layer=licon1_PDIFF $count=1 $X=3.26
+ $Y=1.94 $X2=3.41 $Y2=2.095
r230 2 72 182 $w=1.7e-07 $l=5.3479e-07 $layer=licon1_NDIFF $count=1 $X=4.185
+ $Y=0.37 $X2=4.395 $Y2=0.81
r231 1 62 182 $w=1.7e-07 $l=5.05173e-07 $layer=licon1_NDIFF $count=1 $X=3.255
+ $Y=0.37 $X2=3.395 $Y2=0.81
.ends

.subckt PM_SKY130_FD_SC_HS__O32A_4%B1 1 3 5 6 7 8 10 11 13 15 16 18 19 20 22 23
+ 25 26 27 28 31 33 34 38 49
c148 49 0 7.44774e-20 $X=2.77 $Y=1.615
c149 34 0 6.51508e-20 $X=4.66 $Y=1.615
c150 33 0 7.47943e-20 $X=4.66 $Y=1.615
c151 11 0 7.30872e-20 $X=3.535 $Y=1.165
c152 7 0 1.29542e-19 $X=2.855 $Y=1.165
r153 38 49 4.53993 $w=3.28e-07 $l=1.3e-07 $layer=LI1_cond $X=2.64 $Y=1.615
+ $X2=2.77 $Y2=1.615
r154 38 41 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.69
+ $Y=1.615 $X2=2.69 $Y2=1.615
r155 34 45 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.66 $Y=1.615
+ $X2=4.66 $Y2=1.78
r156 33 36 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=4.66 $Y=1.615
+ $X2=4.66 $Y2=1.765
r157 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.66
+ $Y=1.615 $X2=4.66 $Y2=1.615
r158 30 31 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=5.82 $Y=1.85
+ $X2=5.82 $Y2=2.36
r159 29 36 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.825 $Y=1.765
+ $X2=4.66 $Y2=1.765
r160 28 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.735 $Y=1.765
+ $X2=5.82 $Y2=1.85
r161 28 29 59.369 $w=1.68e-07 $l=9.1e-07 $layer=LI1_cond $X=5.735 $Y=1.765
+ $X2=4.825 $Y2=1.765
r162 26 31 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.735 $Y=2.445
+ $X2=5.82 $Y2=2.36
r163 26 27 187.893 $w=1.68e-07 $l=2.88e-06 $layer=LI1_cond $X=5.735 $Y=2.445
+ $X2=2.855 $Y2=2.445
r164 25 27 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.77 $Y=2.36
+ $X2=2.855 $Y2=2.445
r165 24 49 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.77 $Y=1.78
+ $X2=2.77 $Y2=1.615
r166 24 25 37.8396 $w=1.68e-07 $l=5.8e-07 $layer=LI1_cond $X=2.77 $Y=1.78
+ $X2=2.77 $Y2=2.36
r167 22 45 633.266 $w=1.5e-07 $l=1.235e-06 $layer=POLY_cond $X=4.655 $Y=3.015
+ $X2=4.655 $Y2=1.78
r168 19 22 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.58 $Y=3.09
+ $X2=4.655 $Y2=3.015
r169 19 20 215.362 $w=1.5e-07 $l=4.2e-07 $layer=POLY_cond $X=4.58 $Y=3.09
+ $X2=4.16 $Y2=3.09
r170 16 20 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.085 $Y=3.015
+ $X2=4.16 $Y2=3.09
r171 16 18 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=4.085 $Y=3.015
+ $X2=4.085 $Y2=2.44
r172 13 15 128.533 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=3.61 $Y=1.09 $X2=3.61
+ $Y2=0.69
r173 12 23 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.255 $Y=1.165
+ $X2=3.18 $Y2=1.165
r174 11 13 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.535 $Y=1.165
+ $X2=3.61 $Y2=1.09
r175 11 12 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=3.535 $Y=1.165
+ $X2=3.255 $Y2=1.165
r176 8 23 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.18 $Y=1.09
+ $X2=3.18 $Y2=1.165
r177 8 10 128.533 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=3.18 $Y=1.09 $X2=3.18
+ $Y2=0.69
r178 6 23 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.105 $Y=1.165
+ $X2=3.18 $Y2=1.165
r179 6 7 128.191 $w=1.5e-07 $l=2.5e-07 $layer=POLY_cond $X=3.105 $Y=1.165
+ $X2=2.855 $Y2=1.165
r180 5 41 38.5363 $w=3.15e-07 $l=2.09105e-07 $layer=POLY_cond $X=2.78 $Y=1.45
+ $X2=2.68 $Y2=1.615
r181 4 7 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.78 $Y=1.24
+ $X2=2.855 $Y2=1.165
r182 4 5 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=2.78 $Y=1.24 $X2=2.78
+ $Y2=1.45
r183 1 41 51.5426 $w=3.15e-07 $l=2.89396e-07 $layer=POLY_cond $X=2.595 $Y=1.865
+ $X2=2.68 $Y2=1.615
r184 1 3 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=2.595 $Y=1.865
+ $X2=2.595 $Y2=2.44
.ends

.subckt PM_SKY130_FD_SC_HS__O32A_4%B2 1 3 4 5 6 8 9 11 13 14 16 18 22 24 27 28
r79 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.09
+ $Y=1.435 $X2=4.09 $Y2=1.435
r80 24 28 8.03218 $w=3.28e-07 $l=2.3e-07 $layer=LI1_cond $X=4.09 $Y=1.665
+ $X2=4.09 $Y2=1.435
r81 23 27 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=4.09 $Y=1.45
+ $X2=4.09 $Y2=1.435
r82 21 27 34.0979 $w=3.3e-07 $l=1.95e-07 $layer=POLY_cond $X=4.09 $Y=1.24
+ $X2=4.09 $Y2=1.435
r83 21 22 13.5877 $w=2.4e-07 $l=7.5e-08 $layer=POLY_cond $X=4.09 $Y=1.24
+ $X2=4.09 $Y2=1.165
r84 19 20 82.4064 $w=1.55e-07 $l=2.65e-07 $layer=POLY_cond $X=3.642 $Y=1.525
+ $X2=3.642 $Y2=1.79
r85 16 18 128.533 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=4.61 $Y=1.09 $X2=4.61
+ $Y2=0.69
r86 15 22 12.1617 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.255 $Y=1.165
+ $X2=4.09 $Y2=1.165
r87 14 16 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.535 $Y=1.165
+ $X2=4.61 $Y2=1.09
r88 14 15 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=4.535 $Y=1.165
+ $X2=4.255 $Y2=1.165
r89 11 22 13.5877 $w=2.4e-07 $l=8.44097e-08 $layer=POLY_cond $X=4.11 $Y=1.09
+ $X2=4.09 $Y2=1.165
r90 11 13 128.533 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=4.11 $Y=1.09 $X2=4.11
+ $Y2=0.69
r91 10 19 3.61756 $w=1.5e-07 $l=8.3e-08 $layer=POLY_cond $X=3.725 $Y=1.525
+ $X2=3.642 $Y2=1.525
r92 9 23 32.1775 $w=1.5e-07 $l=1.98997e-07 $layer=POLY_cond $X=3.925 $Y=1.525
+ $X2=4.09 $Y2=1.45
r93 9 10 102.553 $w=1.5e-07 $l=2e-07 $layer=POLY_cond $X=3.925 $Y=1.525
+ $X2=3.725 $Y2=1.525
r94 6 20 23.3226 $w=1.55e-07 $l=7.84219e-08 $layer=POLY_cond $X=3.635 $Y=1.865
+ $X2=3.642 $Y2=1.79
r95 6 8 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=3.635 $Y=1.865
+ $X2=3.635 $Y2=2.44
r96 4 20 3.61756 $w=1.5e-07 $l=8.2e-08 $layer=POLY_cond $X=3.56 $Y=1.79
+ $X2=3.642 $Y2=1.79
r97 4 5 153.83 $w=1.5e-07 $l=3e-07 $layer=POLY_cond $X=3.56 $Y=1.79 $X2=3.26
+ $Y2=1.79
r98 1 5 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.185 $Y=1.865
+ $X2=3.26 $Y2=1.79
r99 1 3 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=3.185 $Y=1.865
+ $X2=3.185 $Y2=2.44
.ends

.subckt PM_SKY130_FD_SC_HS__O32A_4%A3 3 6 7 9 12 15 19 20 21 29
c65 29 0 7.47943e-20 $X=5.66 $Y=1.345
c66 3 0 3.01827e-20 $X=5.14 $Y=0.69
r67 27 29 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=5.57 $Y=1.345 $X2=5.66
+ $Y2=1.345
r68 25 27 69.0702 $w=3.3e-07 $l=3.95e-07 $layer=POLY_cond $X=5.175 $Y=1.345
+ $X2=5.57 $Y2=1.345
r69 23 25 6.12014 $w=3.3e-07 $l=3.5e-08 $layer=POLY_cond $X=5.14 $Y=1.345
+ $X2=5.175 $Y2=1.345
r70 21 27 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.57
+ $Y=1.345 $X2=5.57 $Y2=1.345
r71 19 20 58.8086 $w=1.65e-07 $l=1.35e-07 $layer=POLY_cond $X=5.652 $Y=1.75
+ $X2=5.652 $Y2=1.885
r72 17 29 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.66 $Y=1.51
+ $X2=5.66 $Y2=1.345
r73 17 19 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=5.66 $Y=1.51
+ $X2=5.66 $Y2=1.75
r74 13 29 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.66 $Y=1.18
+ $X2=5.66 $Y2=1.345
r75 13 15 251.255 $w=1.5e-07 $l=4.9e-07 $layer=POLY_cond $X=5.66 $Y=1.18
+ $X2=5.66 $Y2=0.69
r76 12 20 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=5.645 $Y=2.46
+ $X2=5.645 $Y2=1.885
r77 7 9 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=5.175 $Y=1.885
+ $X2=5.175 $Y2=2.46
r78 6 7 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=5.175 $Y=1.795 $X2=5.175
+ $Y2=1.885
r79 5 25 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=5.175 $Y=1.51
+ $X2=5.175 $Y2=1.345
r80 5 6 110.782 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=5.175 $Y=1.51
+ $X2=5.175 $Y2=1.795
r81 1 23 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.14 $Y=1.18
+ $X2=5.14 $Y2=1.345
r82 1 3 251.255 $w=1.5e-07 $l=4.9e-07 $layer=POLY_cond $X=5.14 $Y=1.18 $X2=5.14
+ $Y2=0.69
.ends

.subckt PM_SKY130_FD_SC_HS__O32A_4%A2 1 3 4 6 7 9 10 12 15 17 18 19 20 21 29 30
+ 37 49
c93 18 0 1.50094e-19 $X=6.395 $Y=1.58
c94 7 0 1.91837e-19 $X=6.61 $Y=1.085
r95 35 37 4.15909 $w=1.98e-07 $l=7.5e-08 $layer=LI1_cond $X=6.405 $Y=1.68
+ $X2=6.48 $Y2=1.68
r96 33 49 7.53752 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=7.73 $Y=1.615
+ $X2=7.565 $Y2=1.615
r97 32 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.73
+ $Y=1.615 $X2=7.73 $Y2=1.615
r98 29 30 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.24
+ $Y=1.295 $X2=6.24 $Y2=1.295
r99 21 33 6.63528 $w=3.28e-07 $l=1.9e-07 $layer=LI1_cond $X=7.92 $Y=1.615
+ $X2=7.73 $Y2=1.615
r100 20 49 6.93182 $w=1.98e-07 $l=1.25e-07 $layer=LI1_cond $X=7.44 $Y=1.68
+ $X2=7.565 $Y2=1.68
r101 19 20 26.6182 $w=1.98e-07 $l=4.8e-07 $layer=LI1_cond $X=6.96 $Y=1.68
+ $X2=7.44 $Y2=1.68
r102 18 35 4.52169 $w=2e-07 $l=1.69926e-07 $layer=LI1_cond $X=6.24 $Y=1.69
+ $X2=6.405 $Y2=1.68
r103 18 30 9.66018 $w=3.38e-07 $l=2.85e-07 $layer=LI1_cond $X=6.24 $Y=1.58
+ $X2=6.24 $Y2=1.295
r104 18 19 26.3409 $w=1.98e-07 $l=4.75e-07 $layer=LI1_cond $X=6.485 $Y=1.68
+ $X2=6.96 $Y2=1.68
r105 18 37 0.277273 $w=1.98e-07 $l=5e-09 $layer=LI1_cond $X=6.485 $Y=1.68
+ $X2=6.48 $Y2=1.68
r106 17 29 42.4067 $w=4e-07 $l=3.05e-07 $layer=POLY_cond $X=6.205 $Y=1.6
+ $X2=6.205 $Y2=1.295
r107 15 29 8.34231 $w=4e-07 $l=6e-08 $layer=POLY_cond $X=6.205 $Y=1.235
+ $X2=6.205 $Y2=1.295
r108 15 16 131.899 $w=1.48e-07 $l=4.05e-07 $layer=POLY_cond $X=6.205 $Y=1.16
+ $X2=6.61 $Y2=1.16
r109 13 15 30.9392 $w=1.48e-07 $l=9.5e-08 $layer=POLY_cond $X=6.11 $Y=1.16
+ $X2=6.205 $Y2=1.16
r110 10 32 55.8646 $w=2.93e-07 $l=3.05205e-07 $layer=POLY_cond $X=7.655 $Y=1.885
+ $X2=7.73 $Y2=1.615
r111 10 12 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=7.655 $Y=1.885
+ $X2=7.655 $Y2=2.46
r112 7 16 2.50663 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.61 $Y=1.085
+ $X2=6.61 $Y2=1.16
r113 7 9 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=6.61 $Y=1.085
+ $X2=6.61 $Y2=0.69
r114 4 13 2.50663 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.11 $Y=1.085
+ $X2=6.11 $Y2=1.16
r115 4 6 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=6.11 $Y=1.085
+ $X2=6.11 $Y2=0.69
r116 1 17 41.1287 $w=3.34e-07 $l=3.35522e-07 $layer=POLY_cond $X=6.095 $Y=1.885
+ $X2=6.205 $Y2=1.6
r117 1 3 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=6.095 $Y=1.885
+ $X2=6.095 $Y2=2.46
.ends

.subckt PM_SKY130_FD_SC_HS__O32A_4%A1 1 3 4 5 6 8 9 11 12 14 16 18 20 21 24 25
c69 9 0 8.90518e-20 $X=7.205 $Y=1.885
c70 5 0 1.50094e-19 $X=6.81 $Y=1.81
c71 1 0 8.9584e-20 $X=6.735 $Y=1.885
r72 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.13
+ $Y=1.285 $X2=7.13 $Y2=1.285
r73 21 25 6.7557 $w=2.88e-07 $l=1.7e-07 $layer=LI1_cond $X=6.96 $Y=1.265
+ $X2=7.13 $Y2=1.265
r74 19 24 78.6876 $w=3.3e-07 $l=4.5e-07 $layer=POLY_cond $X=7.13 $Y=1.735
+ $X2=7.13 $Y2=1.285
r75 19 20 13.5877 $w=2.4e-07 $l=7.5e-08 $layer=POLY_cond $X=7.13 $Y=1.735
+ $X2=7.13 $Y2=1.81
r76 17 24 7.86876 $w=3.3e-07 $l=4.5e-08 $layer=POLY_cond $X=7.13 $Y=1.24
+ $X2=7.13 $Y2=1.285
r77 17 18 13.5877 $w=2.4e-07 $l=7.5e-08 $layer=POLY_cond $X=7.13 $Y=1.24
+ $X2=7.13 $Y2=1.165
r78 14 16 128.533 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=7.665 $Y=1.09
+ $X2=7.665 $Y2=0.69
r79 13 18 12.1617 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.295 $Y=1.165
+ $X2=7.13 $Y2=1.165
r80 12 14 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=7.59 $Y=1.165
+ $X2=7.665 $Y2=1.09
r81 12 13 151.266 $w=1.5e-07 $l=2.95e-07 $layer=POLY_cond $X=7.59 $Y=1.165
+ $X2=7.295 $Y2=1.165
r82 9 20 13.5877 $w=2.4e-07 $l=1.06066e-07 $layer=POLY_cond $X=7.205 $Y=1.885
+ $X2=7.13 $Y2=1.81
r83 9 11 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=7.205 $Y=1.885
+ $X2=7.205 $Y2=2.46
r84 6 18 13.5877 $w=2.4e-07 $l=1.21861e-07 $layer=POLY_cond $X=7.04 $Y=1.09
+ $X2=7.13 $Y2=1.165
r85 6 8 128.533 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=7.04 $Y=1.09 $X2=7.04
+ $Y2=0.69
r86 4 20 12.1617 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.965 $Y=1.81
+ $X2=7.13 $Y2=1.81
r87 4 5 79.4787 $w=1.5e-07 $l=1.55e-07 $layer=POLY_cond $X=6.965 $Y=1.81
+ $X2=6.81 $Y2=1.81
r88 1 5 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=6.735 $Y=1.885
+ $X2=6.81 $Y2=1.81
r89 1 3 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=6.735 $Y=1.885
+ $X2=6.735 $Y2=2.46
.ends

.subckt PM_SKY130_FD_SC_HS__O32A_4%VPWR 1 2 3 4 5 16 18 24 26 30 36 40 43 44 45
+ 47 59 68 69 75 78 81
r98 81 82 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r99 78 79 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r100 76 79 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.16 $Y2=3.33
r101 75 76 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r102 72 73 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r103 69 82 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=7.92 $Y=3.33
+ $X2=6.96 $Y2=3.33
r104 68 69 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r105 66 81 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.135 $Y=3.33
+ $X2=6.97 $Y2=3.33
r106 66 68 51.2139 $w=1.68e-07 $l=7.85e-07 $layer=LI1_cond $X=7.135 $Y=3.33
+ $X2=7.92 $Y2=3.33
r107 65 82 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=6.96 $Y2=3.33
r108 64 65 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r109 62 65 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=6.48 $Y2=3.33
r110 61 64 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=4.56 $Y=3.33
+ $X2=6.48 $Y2=3.33
r111 61 62 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r112 59 81 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.805 $Y=3.33
+ $X2=6.97 $Y2=3.33
r113 59 64 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=6.805 $Y=3.33
+ $X2=6.48 $Y2=3.33
r114 55 79 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=2.16 $Y2=3.33
r115 54 57 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=2.64 $Y=3.33
+ $X2=4.08 $Y2=3.33
r116 54 55 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r117 52 78 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.415 $Y=3.33
+ $X2=2.25 $Y2=3.33
r118 52 54 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=2.415 $Y=3.33
+ $X2=2.64 $Y2=3.33
r119 51 76 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r120 51 73 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r121 50 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r122 48 72 4.00981 $w=1.7e-07 $l=1.83e-07 $layer=LI1_cond $X=0.365 $Y=3.33
+ $X2=0.182 $Y2=3.33
r123 48 50 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=0.365 $Y=3.33
+ $X2=0.72 $Y2=3.33
r124 47 75 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.065 $Y=3.33
+ $X2=1.23 $Y2=3.33
r125 47 50 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.065 $Y=3.33
+ $X2=0.72 $Y2=3.33
r126 45 62 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=4.56 $Y2=3.33
r127 45 55 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=2.64 $Y2=3.33
r128 45 57 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r129 43 57 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=4.195 $Y=3.33
+ $X2=4.08 $Y2=3.33
r130 43 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.195 $Y=3.33
+ $X2=4.36 $Y2=3.33
r131 42 61 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=4.525 $Y=3.33
+ $X2=4.56 $Y2=3.33
r132 42 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.525 $Y=3.33
+ $X2=4.36 $Y2=3.33
r133 38 81 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.97 $Y=3.245
+ $X2=6.97 $Y2=3.33
r134 38 40 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=6.97 $Y=3.245
+ $X2=6.97 $Y2=2.815
r135 34 44 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.36 $Y=3.245
+ $X2=4.36 $Y2=3.33
r136 34 36 15.8897 $w=3.28e-07 $l=4.55e-07 $layer=LI1_cond $X=4.36 $Y=3.245
+ $X2=4.36 $Y2=2.79
r137 30 33 24.4458 $w=3.28e-07 $l=7e-07 $layer=LI1_cond $X=2.25 $Y=2.115
+ $X2=2.25 $Y2=2.815
r138 28 78 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.25 $Y=3.245
+ $X2=2.25 $Y2=3.33
r139 28 33 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=2.25 $Y=3.245
+ $X2=2.25 $Y2=2.815
r140 27 75 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.395 $Y=3.33
+ $X2=1.23 $Y2=3.33
r141 26 78 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.085 $Y=3.33
+ $X2=2.25 $Y2=3.33
r142 26 27 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=2.085 $Y=3.33
+ $X2=1.395 $Y2=3.33
r143 22 75 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.23 $Y=3.245
+ $X2=1.23 $Y2=3.33
r144 22 24 33.5256 $w=3.28e-07 $l=9.6e-07 $layer=LI1_cond $X=1.23 $Y=3.245
+ $X2=1.23 $Y2=2.285
r145 18 21 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=0.24 $Y=1.985
+ $X2=0.24 $Y2=2.815
r146 16 72 3.13335 $w=2.5e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.24 $Y=3.245
+ $X2=0.182 $Y2=3.33
r147 16 21 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=0.24 $Y=3.245
+ $X2=0.24 $Y2=2.815
r148 5 40 600 $w=1.7e-07 $l=9.31571e-07 $layer=licon1_PDIFF $count=1 $X=6.81
+ $Y=1.96 $X2=6.97 $Y2=2.815
r149 4 36 600 $w=1.7e-07 $l=9.44722e-07 $layer=licon1_PDIFF $count=1 $X=4.16
+ $Y=1.94 $X2=4.36 $Y2=2.79
r150 3 33 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=2.1
+ $Y=1.84 $X2=2.25 $Y2=2.815
r151 3 30 400 $w=1.7e-07 $l=3.4187e-07 $layer=licon1_PDIFF $count=1 $X=2.1
+ $Y=1.84 $X2=2.25 $Y2=2.115
r152 2 24 300 $w=1.7e-07 $l=5.35747e-07 $layer=licon1_PDIFF $count=2 $X=1.03
+ $Y=1.84 $X2=1.23 $Y2=2.285
r153 1 21 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.815
r154 1 18 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HS__O32A_4%X 1 2 3 4 13 15 16 19 25 27 29 33 39 42 45 48
+ 51
c76 27 0 3.73162e-20 $X=1.565 $Y=1.865
c77 15 0 1.0009e-19 $X=0.565 $Y=1.565
c78 13 0 8.40338e-20 $X=0.685 $Y=1.225
r79 48 51 2.9826 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.24 $Y=1.225 $X2=0.24
+ $Y2=1.31
r80 48 51 1.75372 $w=2.28e-07 $l=3.5e-08 $layer=LI1_cond $X=0.24 $Y=1.345
+ $X2=0.24 $Y2=1.31
r81 45 46 6.9845 $w=3.28e-07 $l=2e-07 $layer=LI1_cond $X=0.85 $Y=1.025 $X2=0.85
+ $Y2=1.225
r82 42 44 10.4768 $w=3.28e-07 $l=3e-07 $layer=LI1_cond $X=0.73 $Y=1.565 $X2=0.73
+ $Y2=1.865
r83 41 48 6.76434 $w=2.28e-07 $l=1.35e-07 $layer=LI1_cond $X=0.24 $Y=1.48
+ $X2=0.24 $Y2=1.345
r84 37 39 14.8421 $w=3.28e-07 $l=4.25e-07 $layer=LI1_cond $X=1.85 $Y=0.94
+ $X2=1.85 $Y2=0.515
r85 33 35 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=1.73 $Y=1.985
+ $X2=1.73 $Y2=2.815
r86 31 33 1.22229 $w=3.28e-07 $l=3.5e-08 $layer=LI1_cond $X=1.73 $Y=1.95
+ $X2=1.73 $Y2=1.985
r87 30 45 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.015 $Y=1.025
+ $X2=0.85 $Y2=1.025
r88 29 37 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.685 $Y=1.025
+ $X2=1.85 $Y2=0.94
r89 29 30 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.685 $Y=1.025
+ $X2=1.015 $Y2=1.025
r90 28 44 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.895 $Y=1.865
+ $X2=0.73 $Y2=1.865
r91 27 31 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.565 $Y=1.865
+ $X2=1.73 $Y2=1.95
r92 27 28 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.565 $Y=1.865
+ $X2=0.895 $Y2=1.865
r93 23 45 2.96841 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=0.85 $Y=0.94
+ $X2=0.85 $Y2=1.025
r94 23 25 14.8421 $w=3.28e-07 $l=4.25e-07 $layer=LI1_cond $X=0.85 $Y=0.94
+ $X2=0.85 $Y2=0.515
r95 19 21 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=0.73 $Y=1.985
+ $X2=0.73 $Y2=2.815
r96 17 44 2.96841 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=0.73 $Y=1.95
+ $X2=0.73 $Y2=1.865
r97 17 19 1.22229 $w=3.28e-07 $l=3.5e-08 $layer=LI1_cond $X=0.73 $Y=1.95
+ $X2=0.73 $Y2=1.985
r98 16 41 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=0.355 $Y=1.565
+ $X2=0.24 $Y2=1.48
r99 15 42 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.565 $Y=1.565
+ $X2=0.73 $Y2=1.565
r100 15 16 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=0.565 $Y=1.565
+ $X2=0.355 $Y2=1.565
r101 14 48 4.03528 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=0.355 $Y=1.225
+ $X2=0.24 $Y2=1.225
r102 13 46 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.685 $Y=1.225
+ $X2=0.85 $Y2=1.225
r103 13 14 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=0.685 $Y=1.225
+ $X2=0.355 $Y2=1.225
r104 4 35 400 $w=1.7e-07 $l=1.07034e-06 $layer=licon1_PDIFF $count=1 $X=1.53
+ $Y=1.84 $X2=1.73 $Y2=2.815
r105 4 33 400 $w=1.7e-07 $l=2.62678e-07 $layer=licon1_PDIFF $count=1 $X=1.53
+ $Y=1.84 $X2=1.73 $Y2=1.985
r106 3 21 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=0.58
+ $Y=1.84 $X2=0.73 $Y2=2.815
r107 3 19 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=0.58
+ $Y=1.84 $X2=0.73 $Y2=1.985
r108 2 39 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.71
+ $Y=0.37 $X2=1.85 $Y2=0.515
r109 1 25 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=0.71
+ $Y=0.37 $X2=0.85 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__O32A_4%A_534_388# 1 2 11
r18 8 11 42.995 $w=2.58e-07 $l=9.7e-07 $layer=LI1_cond $X=2.89 $Y=2.83 $X2=3.86
+ $Y2=2.83
r19 2 11 600 $w=1.7e-07 $l=9.21954e-07 $layer=licon1_PDIFF $count=1 $X=3.71
+ $Y=1.94 $X2=3.86 $Y2=2.79
r20 1 8 600 $w=1.7e-07 $l=9.48644e-07 $layer=licon1_PDIFF $count=1 $X=2.67
+ $Y=1.94 $X2=2.89 $Y2=2.785
.ends

.subckt PM_SKY130_FD_SC_HS__O32A_4%A_961_392# 1 2 3 10 17 18 19 22 26 28
c50 19 0 1.81307e-19 $X=6.245 $Y=2.475
r51 24 28 3.10218 $w=3.05e-07 $l=9.66954e-08 $layer=LI1_cond $X=7.905 $Y=2.39
+ $X2=7.88 $Y2=2.475
r52 24 26 11.3186 $w=2.78e-07 $l=2.75e-07 $layer=LI1_cond $X=7.905 $Y=2.39
+ $X2=7.905 $Y2=2.115
r53 20 28 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=7.88 $Y=2.56
+ $X2=7.88 $Y2=2.475
r54 20 22 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=7.88 $Y=2.56
+ $X2=7.88 $Y2=2.815
r55 18 28 3.51065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.715 $Y=2.475
+ $X2=7.88 $Y2=2.475
r56 18 19 95.9037 $w=1.68e-07 $l=1.47e-06 $layer=LI1_cond $X=7.715 $Y=2.475
+ $X2=6.245 $Y2=2.475
r57 16 19 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.16 $Y=2.56
+ $X2=6.245 $Y2=2.475
r58 16 17 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=6.16 $Y=2.56
+ $X2=6.16 $Y2=2.7
r59 12 15 37.866 $w=2.78e-07 $l=9.2e-07 $layer=LI1_cond $X=4.95 $Y=2.84 $X2=5.87
+ $Y2=2.84
r60 10 17 7.36005 $w=2.8e-07 $l=1.77482e-07 $layer=LI1_cond $X=6.075 $Y=2.84
+ $X2=6.16 $Y2=2.7
r61 10 15 8.43753 $w=2.78e-07 $l=2.05e-07 $layer=LI1_cond $X=6.075 $Y=2.84
+ $X2=5.87 $Y2=2.84
r62 3 26 300 $w=1.7e-07 $l=2.17428e-07 $layer=licon1_PDIFF $count=2 $X=7.73
+ $Y=1.96 $X2=7.88 $Y2=2.115
r63 3 22 600 $w=1.7e-07 $l=9.26971e-07 $layer=licon1_PDIFF $count=1 $X=7.73
+ $Y=1.96 $X2=7.88 $Y2=2.815
r64 2 15 600 $w=1.7e-07 $l=9.11921e-07 $layer=licon1_PDIFF $count=1 $X=5.72
+ $Y=1.96 $X2=5.87 $Y2=2.8
r65 1 12 600 $w=1.7e-07 $l=9.09615e-07 $layer=licon1_PDIFF $count=1 $X=4.805
+ $Y=1.96 $X2=4.95 $Y2=2.8
.ends

.subckt PM_SKY130_FD_SC_HS__O32A_4%A_1234_392# 1 2 7 13 15 16
c23 15 0 8.9584e-20 $X=7.43 $Y=2.115
c24 13 0 8.90518e-20 $X=6.675 $Y=2.095
c25 1 0 1.81307e-19 $X=6.17 $Y=1.96
r26 15 16 7.69997 $w=2.48e-07 $l=1.65e-07 $layer=LI1_cond $X=7.43 $Y=2.075
+ $X2=7.265 $Y2=2.075
r27 13 16 29.5627 $w=2.28e-07 $l=5.9e-07 $layer=LI1_cond $X=6.675 $Y=2.085
+ $X2=7.265 $Y2=2.085
r28 7 13 5.85606 $w=2.48e-07 $l=1.25e-07 $layer=LI1_cond $X=6.55 $Y=2.095
+ $X2=6.675 $Y2=2.095
r29 7 9 6.22319 $w=2.48e-07 $l=1.35e-07 $layer=LI1_cond $X=6.55 $Y=2.095
+ $X2=6.415 $Y2=2.095
r30 2 15 600 $w=1.7e-07 $l=2.17428e-07 $layer=licon1_PDIFF $count=1 $X=7.28
+ $Y=1.96 $X2=7.43 $Y2=2.115
r31 1 9 600 $w=1.7e-07 $l=3.2078e-07 $layer=licon1_PDIFF $count=1 $X=6.17
+ $Y=1.96 $X2=6.415 $Y2=2.135
.ends

.subckt PM_SKY130_FD_SC_HS__O32A_4%VGND 1 2 3 4 5 6 19 21 23 27 31 35 39 43 46
+ 47 49 50 52 53 54 69 75 76 82 85
r107 85 86 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=0 $X2=7.44
+ $Y2=0
r108 82 83 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r109 80 83 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=1.2
+ $Y2=0
r110 79 80 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r111 76 86 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=0 $X2=7.44
+ $Y2=0
r112 75 76 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=0 $X2=7.92
+ $Y2=0
r113 73 85 9.56655 $w=1.7e-07 $l=1.93e-07 $layer=LI1_cond $X=7.545 $Y=0
+ $X2=7.352 $Y2=0
r114 73 75 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=7.545 $Y=0
+ $X2=7.92 $Y2=0
r115 72 86 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=0 $X2=7.44
+ $Y2=0
r116 71 72 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.96 $Y=0 $X2=6.96
+ $Y2=0
r117 69 85 9.56655 $w=1.7e-07 $l=1.92e-07 $layer=LI1_cond $X=7.16 $Y=0 $X2=7.352
+ $Y2=0
r118 69 71 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=7.16 $Y=0 $X2=6.96
+ $Y2=0
r119 68 72 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6 $Y=0 $X2=6.96
+ $Y2=0
r120 67 68 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6 $Y=0 $X2=6 $Y2=0
r121 65 68 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=6
+ $Y2=0
r122 64 65 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r123 61 64 156.578 $w=1.68e-07 $l=2.4e-06 $layer=LI1_cond $X=2.64 $Y=0 $X2=5.04
+ $Y2=0
r124 61 62 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r125 59 62 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r126 59 83 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.2
+ $Y2=0
r127 58 59 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r128 56 82 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.515 $Y=0 $X2=1.35
+ $Y2=0
r129 56 58 42.0802 $w=1.68e-07 $l=6.45e-07 $layer=LI1_cond $X=1.515 $Y=0
+ $X2=2.16 $Y2=0
r130 54 65 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=5.04
+ $Y2=0
r131 54 62 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=4.08 $Y=0
+ $X2=2.64 $Y2=0
r132 52 67 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=6.23 $Y=0 $X2=6
+ $Y2=0
r133 52 53 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.23 $Y=0 $X2=6.395
+ $Y2=0
r134 51 71 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=6.56 $Y=0 $X2=6.96
+ $Y2=0
r135 51 53 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.56 $Y=0 $X2=6.395
+ $Y2=0
r136 49 64 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=5.23 $Y=0 $X2=5.04
+ $Y2=0
r137 49 50 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.23 $Y=0 $X2=5.395
+ $Y2=0
r138 48 67 28.7059 $w=1.68e-07 $l=4.4e-07 $layer=LI1_cond $X=5.56 $Y=0 $X2=6
+ $Y2=0
r139 48 50 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.56 $Y=0 $X2=5.395
+ $Y2=0
r140 46 58 5.21925 $w=1.68e-07 $l=8e-08 $layer=LI1_cond $X=2.24 $Y=0 $X2=2.16
+ $Y2=0
r141 46 47 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.24 $Y=0 $X2=2.405
+ $Y2=0
r142 45 61 4.56684 $w=1.68e-07 $l=7e-08 $layer=LI1_cond $X=2.57 $Y=0 $X2=2.64
+ $Y2=0
r143 45 47 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.57 $Y=0 $X2=2.405
+ $Y2=0
r144 41 85 1.35792 $w=3.85e-07 $l=8.5e-08 $layer=LI1_cond $X=7.352 $Y=0.085
+ $X2=7.352 $Y2=0
r145 41 43 12.8714 $w=3.83e-07 $l=4.3e-07 $layer=LI1_cond $X=7.352 $Y=0.085
+ $X2=7.352 $Y2=0.515
r146 37 53 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.395 $Y=0.085
+ $X2=6.395 $Y2=0
r147 37 39 15.1913 $w=3.28e-07 $l=4.35e-07 $layer=LI1_cond $X=6.395 $Y=0.085
+ $X2=6.395 $Y2=0.52
r148 33 50 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.395 $Y=0.085
+ $X2=5.395 $Y2=0
r149 33 35 15.3659 $w=3.28e-07 $l=4.4e-07 $layer=LI1_cond $X=5.395 $Y=0.085
+ $X2=5.395 $Y2=0.525
r150 29 47 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.405 $Y=0.085
+ $X2=2.405 $Y2=0
r151 29 31 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=2.405 $Y=0.085
+ $X2=2.405 $Y2=0.515
r152 25 82 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.35 $Y=0.085
+ $X2=1.35 $Y2=0
r153 25 27 16.5882 $w=3.28e-07 $l=4.75e-07 $layer=LI1_cond $X=1.35 $Y=0.085
+ $X2=1.35 $Y2=0.56
r154 24 79 4.59558 $w=1.7e-07 $l=2.58e-07 $layer=LI1_cond $X=0.515 $Y=0
+ $X2=0.257 $Y2=0
r155 23 82 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.185 $Y=0 $X2=1.35
+ $Y2=0
r156 23 24 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.185 $Y=0
+ $X2=0.515 $Y2=0
r157 19 79 3.17059 $w=3.3e-07 $l=1.28662e-07 $layer=LI1_cond $X=0.35 $Y=0.085
+ $X2=0.257 $Y2=0
r158 19 21 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=0.35 $Y=0.085
+ $X2=0.35 $Y2=0.515
r159 6 43 182 $w=1.7e-07 $l=2.98831e-07 $layer=licon1_NDIFF $count=1 $X=7.115
+ $Y=0.37 $X2=7.35 $Y2=0.515
r160 5 39 182 $w=1.7e-07 $l=2.74955e-07 $layer=licon1_NDIFF $count=1 $X=6.185
+ $Y=0.37 $X2=6.395 $Y2=0.52
r161 4 35 182 $w=1.7e-07 $l=2.45561e-07 $layer=licon1_NDIFF $count=1 $X=5.215
+ $Y=0.37 $X2=5.395 $Y2=0.525
r162 3 31 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.265
+ $Y=0.37 $X2=2.405 $Y2=0.515
r163 2 27 182 $w=1.7e-07 $l=2.89828e-07 $layer=licon1_NDIFF $count=1 $X=1.14
+ $Y=0.37 $X2=1.35 $Y2=0.56
r164 1 21 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.205
+ $Y=0.37 $X2=0.35 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__O32A_4%A_564_74# 1 2 3 4 5 6 21 23 24 27 29 32 35 39
+ 41 45 47 51 53 56 58
c99 56 0 7.70569e-20 $X=5.895 $Y=0.87
c100 45 0 1.44963e-19 $X=6.825 $Y=0.515
r101 49 51 9.25447 $w=3.28e-07 $l=2.65e-07 $layer=LI1_cond $X=7.88 $Y=0.78
+ $X2=7.88 $Y2=0.515
r102 48 58 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.99 $Y=0.865
+ $X2=6.865 $Y2=0.865
r103 47 49 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=7.715 $Y=0.865
+ $X2=7.88 $Y2=0.78
r104 47 48 47.2995 $w=1.68e-07 $l=7.25e-07 $layer=LI1_cond $X=7.715 $Y=0.865
+ $X2=6.99 $Y2=0.865
r105 43 58 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.865 $Y=0.78
+ $X2=6.865 $Y2=0.865
r106 43 45 12.2159 $w=2.48e-07 $l=2.65e-07 $layer=LI1_cond $X=6.865 $Y=0.78
+ $X2=6.865 $Y2=0.515
r107 42 56 8.61065 $w=1.7e-07 $l=1.67481e-07 $layer=LI1_cond $X=6.06 $Y=0.865
+ $X2=5.895 $Y2=0.87
r108 41 58 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.74 $Y=0.865
+ $X2=6.865 $Y2=0.865
r109 41 42 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=6.74 $Y=0.865
+ $X2=6.06 $Y2=0.865
r110 37 56 0.89609 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=5.895 $Y=0.78
+ $X2=5.895 $Y2=0.87
r111 37 39 9.25447 $w=3.28e-07 $l=2.65e-07 $layer=LI1_cond $X=5.895 $Y=0.78
+ $X2=5.895 $Y2=0.515
r112 36 55 4.91858 $w=1.7e-07 $l=1.77059e-07 $layer=LI1_cond $X=5.06 $Y=0.875
+ $X2=4.895 $Y2=0.9
r113 35 56 8.61065 $w=1.7e-07 $l=1.67481e-07 $layer=LI1_cond $X=5.73 $Y=0.875
+ $X2=5.895 $Y2=0.87
r114 35 36 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.73 $Y=0.875
+ $X2=5.06 $Y2=0.875
r115 32 55 2.8476 $w=3.3e-07 $l=1.1e-07 $layer=LI1_cond $X=4.895 $Y=0.79
+ $X2=4.895 $Y2=0.9
r116 32 34 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=4.895 $Y=0.79
+ $X2=4.895 $Y2=0.515
r117 31 34 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=4.895 $Y=0.425
+ $X2=4.895 $Y2=0.515
r118 30 53 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.06 $Y=0.34
+ $X2=3.895 $Y2=0.34
r119 29 31 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.73 $Y=0.34
+ $X2=4.895 $Y2=0.425
r120 29 30 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.73 $Y=0.34
+ $X2=4.06 $Y2=0.34
r121 25 53 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.895 $Y=0.425
+ $X2=3.895 $Y2=0.34
r122 25 27 5.93683 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=3.895 $Y=0.425
+ $X2=3.895 $Y2=0.595
r123 23 53 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.73 $Y=0.34
+ $X2=3.895 $Y2=0.34
r124 23 24 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=3.73 $Y=0.34 $X2=3.13
+ $Y2=0.34
r125 19 24 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.965 $Y=0.425
+ $X2=3.13 $Y2=0.34
r126 19 21 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=2.965 $Y=0.425
+ $X2=2.965 $Y2=0.515
r127 6 51 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=7.74
+ $Y=0.37 $X2=7.88 $Y2=0.515
r128 5 58 182 $w=1.7e-07 $l=5.60647e-07 $layer=licon1_NDIFF $count=1 $X=6.685
+ $Y=0.37 $X2=6.825 $Y2=0.865
r129 5 45 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=6.685
+ $Y=0.37 $X2=6.825 $Y2=0.515
r130 4 39 91 $w=1.7e-07 $l=2.20907e-07 $layer=licon1_NDIFF $count=2 $X=5.735
+ $Y=0.37 $X2=5.895 $Y2=0.515
r131 3 55 182 $w=1.7e-07 $l=6.11044e-07 $layer=licon1_NDIFF $count=1 $X=4.685
+ $Y=0.37 $X2=4.895 $Y2=0.885
r132 3 34 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=4.685
+ $Y=0.37 $X2=4.895 $Y2=0.515
r133 2 27 182 $w=1.7e-07 $l=3.1285e-07 $layer=licon1_NDIFF $count=1 $X=3.685
+ $Y=0.37 $X2=3.895 $Y2=0.595
r134 1 21 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=2.82
+ $Y=0.37 $X2=2.965 $Y2=0.515
.ends

