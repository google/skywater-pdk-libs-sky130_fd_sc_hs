* NGSPICE file created from sky130_fd_sc_hs__clkbuf_1.ext - technology: sky130A

.subckt sky130_fd_sc_hs__clkbuf_1 A VGND VNB VPB VPWR X
M1000 X a_27_74# VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=3.304e+11p pd=2.83e+06u as=4.48e+11p ps=3.04e+06u
M1001 X a_27_74# VGND VNB nlowvt w=420000u l=150000u
+  ad=1.19e+11p pd=1.41e+06u as=3.276e+11p ps=2.4e+06u
M1002 VGND A a_27_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.197e+11p ps=1.41e+06u
M1003 VPWR A a_27_74# VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=3.304e+11p ps=2.83e+06u
.ends

