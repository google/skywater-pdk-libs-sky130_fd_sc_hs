# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_hs__a2bb2o_2
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_hs__a2bb2o_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.800000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1_N
    ANTENNAGATEAREA  0.232500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.925000 1.180000 3.255000 2.150000 ;
    END
  END A1_N
  PIN A2_N
    ANTENNAGATEAREA  0.232500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.385000 1.180000 2.755000 1.510000 ;
    END
  END A2_N
  PIN B1
    ANTENNAGATEAREA  0.261000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105000 1.180000 0.435000 1.550000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.261000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605000 1.180000 1.315000 1.550000 ;
    END
  END B2
  PIN X
    ANTENNADIFFAREA  0.543200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.485000 0.350000 3.920000 2.150000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 4.800000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 4.800000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.800000 0.085000 ;
      RECT 0.000000  3.245000 4.800000 3.415000 ;
      RECT 0.265000  1.720000 1.415000 1.890000 ;
      RECT 0.265000  1.890000 0.515000 2.980000 ;
      RECT 0.290000  0.085000 0.620000 1.010000 ;
      RECT 0.715000  2.060000 1.045000 3.245000 ;
      RECT 1.080000  0.350000 1.480000 0.840000 ;
      RECT 1.080000  0.840000 1.655000 1.010000 ;
      RECT 1.245000  1.890000 1.415000 2.980000 ;
      RECT 1.485000  1.010000 1.655000 1.380000 ;
      RECT 1.485000  1.380000 1.755000 1.550000 ;
      RECT 1.585000  1.550000 1.755000 2.020000 ;
      RECT 1.585000  2.020000 1.945000 2.810000 ;
      RECT 1.585000  2.810000 2.920000 2.980000 ;
      RECT 1.650000  0.085000 2.520000 0.670000 ;
      RECT 1.925000  0.840000 2.870000 1.010000 ;
      RECT 1.925000  1.010000 2.175000 1.680000 ;
      RECT 1.925000  1.680000 2.580000 1.850000 ;
      RECT 2.265000  1.850000 2.580000 2.640000 ;
      RECT 2.690000  0.350000 2.870000 0.840000 ;
      RECT 2.750000  2.320000 4.470000 2.490000 ;
      RECT 2.750000  2.490000 2.920000 2.810000 ;
      RECT 3.050000  0.085000 3.315000 0.940000 ;
      RECT 3.105000  2.660000 3.495000 3.245000 ;
      RECT 4.065000  2.660000 4.395000 3.245000 ;
      RECT 4.090000  1.350000 4.470000 2.320000 ;
      RECT 4.100000  0.085000 4.350000 1.130000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
  END
END sky130_fd_sc_hs__a2bb2o_2
