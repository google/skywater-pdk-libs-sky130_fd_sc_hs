* File: sky130_fd_sc_hs__buf_1.spice
* Created: Thu Aug 27 20:34:19 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hs__buf_1.pex.spice"
.subckt sky130_fd_sc_hs__buf_1  VNB VPB A VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A	A
* VPB	VPB
* VNB	VNB
MM1002 N_VGND_M1002_d N_A_M1002_g N_A_27_164#_M1002_s VNB NLOWVT L=0.15 W=0.55
+ AD=0.129591 AS=0.24915 PD=0.997674 PS=2.37 NRD=18 NRS=0 M=1 R=3.66667
+ SA=75000.4 SB=75000.8 A=0.0825 P=1.4 MULT=1
MM1003 N_X_M1003_d N_A_27_164#_M1003_g N_VGND_M1002_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.174359 PD=2.05 PS=1.34233 NRD=0 NRS=11.34 M=1 R=4.93333
+ SA=75000.8 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1001 N_VPWR_M1001_d N_A_M1001_g N_A_27_164#_M1001_s VPB PSHORT L=0.15 W=0.84
+ AD=0.1758 AS=0.2478 PD=1.30286 PS=2.27 NRD=14.0658 NRS=2.3443 M=1 R=5.6
+ SA=75000.2 SB=75000.8 A=0.126 P=1.98 MULT=1
MM1000 N_X_M1000_d N_A_27_164#_M1000_g N_VPWR_M1001_d VPB PSHORT L=0.15 W=1.12
+ AD=0.3304 AS=0.2344 PD=2.83 PS=1.73714 NRD=1.7533 NRS=10.5395 M=1 R=7.46667
+ SA=75000.6 SB=75000.2 A=0.168 P=2.54 MULT=1
DX4_noxref VNB VPB NWDIODE A=4.278 P=8.32
*
.include "sky130_fd_sc_hs__buf_1.pxi.spice"
*
.ends
*
*
