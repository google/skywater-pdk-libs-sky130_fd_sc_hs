* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hs__einvp_1 A TE VGND VNB VPB VPWR Z
X0 VGND TE a_318_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X1 a_310_392# A Z VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=150000u
X2 a_44_549# TE VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X3 a_44_549# TE VPWR VPB sky130_fd_pr__pfet_01v8 w=420000u l=150000u
X4 VPWR a_44_549# a_310_392# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=150000u
X5 a_318_74# A Z VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
.ends
