* NGSPICE file created from sky130_fd_sc_hs__or2b_4.ext - technology: sky130A

.subckt sky130_fd_sc_hs__or2b_4 A B_N VGND VNB VPB VPWR X
M1000 X a_81_296# VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=6.72e+11p pd=5.68e+06u as=1.6394e+12p ps=1.379e+07u
M1001 VPWR a_81_296# X VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1002 X a_81_296# VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1003 VPWR a_81_296# X VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_676_48# B_N VPWR VPB pshort w=1e+06u l=150000u
+  ad=2.85e+11p pd=2.57e+06u as=0p ps=0u
M1005 a_81_296# A VGND VNB nlowvt w=640000u l=150000u
+  ad=4.672e+11p pd=4.02e+06u as=1.1509e+12p ps=1.032e+07u
M1006 a_81_296# a_676_48# a_489_392# VPB pshort w=1e+06u l=150000u
+  ad=3e+11p pd=2.6e+06u as=8.8e+11p ps=7.76e+06u
M1007 VGND a_81_296# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=4.329e+11p ps=4.13e+06u
M1008 a_81_296# a_676_48# VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_489_392# a_676_48# a_81_296# VPB pshort w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VGND A a_81_296# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_489_392# A VPWR VPB pshort w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VPWR A a_489_392# VPB pshort w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 X a_81_296# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 X a_81_296# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VGND a_81_296# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_676_48# B_N VGND VNB nlowvt w=640000u l=150000u
+  ad=6.272e+11p pd=3.24e+06u as=0p ps=0u
M1017 VGND a_676_48# a_81_296# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

