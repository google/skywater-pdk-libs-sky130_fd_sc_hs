# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_hs__a2111o_1
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_hs__a2111o_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.320000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 0.440000 0.840000 0.670000 ;
        RECT 0.510000 0.255000 0.840000 0.440000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.050000 1.500000 2.275000 1.800000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.435000 0.255000 1.795000 0.490000 ;
        RECT 1.595000 0.490000 1.795000 0.670000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.005000 0.255000 2.335000 0.490000 ;
        RECT 2.005000 0.490000 2.245000 0.670000 ;
    END
  END C1
  PIN D1
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.445000 1.500000 2.775000 1.800000 ;
    END
  END D1
  PIN X
    ANTENNADIFFAREA  0.504100 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.860000 0.370000 4.195000 2.980000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 4.320000 0.085000 ;
        RECT 1.095000  0.085000 1.265000 0.660000 ;
        RECT 1.095000  0.660000 1.425000 0.990000 ;
        RECT 2.415000  0.660000 2.675000 0.990000 ;
        RECT 2.505000  0.085000 2.675000 0.660000 ;
        RECT 3.435000  0.085000 3.685000 1.150000 ;
      LAYER mcon ;
        RECT 0.155000 -0.085000 0.325000 0.085000 ;
        RECT 0.635000 -0.085000 0.805000 0.085000 ;
        RECT 1.115000 -0.085000 1.285000 0.085000 ;
        RECT 1.595000 -0.085000 1.765000 0.085000 ;
        RECT 2.075000 -0.085000 2.245000 0.085000 ;
        RECT 2.555000 -0.085000 2.725000 0.085000 ;
        RECT 3.035000 -0.085000 3.205000 0.085000 ;
        RECT 3.515000 -0.085000 3.685000 0.085000 ;
        RECT 3.995000 -0.085000 4.165000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.245000 4.320000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 3.245000 4.320000 3.415000 ;
        RECT 0.890000 2.310000 1.100000 3.245000 ;
        RECT 3.410000 1.820000 3.660000 3.245000 ;
      LAYER mcon ;
        RECT 0.155000 3.245000 0.325000 3.415000 ;
        RECT 0.635000 3.245000 0.805000 3.415000 ;
        RECT 1.115000 3.245000 1.285000 3.415000 ;
        RECT 1.595000 3.245000 1.765000 3.415000 ;
        RECT 2.075000 3.245000 2.245000 3.415000 ;
        RECT 2.555000 3.245000 2.725000 3.415000 ;
        RECT 3.035000 3.245000 3.205000 3.415000 ;
        RECT 3.515000 3.245000 3.685000 3.415000 ;
        RECT 3.995000 3.245000 4.165000 3.415000 ;
      LAYER met1 ;
        RECT 0.000000 3.085000 4.320000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.360000 1.940000 0.690000 1.970000 ;
      RECT 0.360000 1.970000 1.630000 2.140000 ;
      RECT 0.360000 2.140000 0.690000 2.980000 ;
      RECT 0.385000 0.840000 0.715000 1.160000 ;
      RECT 0.385000 1.160000 3.115000 1.320000 ;
      RECT 0.385000 1.320000 3.690000 1.330000 ;
      RECT 0.385000 1.330000 0.715000 1.340000 ;
      RECT 1.300000 2.140000 1.630000 2.980000 ;
      RECT 1.715000 0.840000 2.045000 1.160000 ;
      RECT 2.530000 1.970000 3.115000 2.140000 ;
      RECT 2.530000 2.140000 2.860000 2.980000 ;
      RECT 2.845000 0.660000 3.115000 1.160000 ;
      RECT 2.945000 1.330000 3.690000 1.650000 ;
      RECT 2.945000 1.650000 3.115000 1.970000 ;
  END
END sky130_fd_sc_hs__a2111o_1
