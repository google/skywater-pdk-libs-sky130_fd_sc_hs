* File: sky130_fd_sc_hs__a21boi_1.spice
* Created: Tue Sep  1 19:49:16 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hs__a21boi_1.pex.spice"
.subckt sky130_fd_sc_hs__a21boi_1  VNB VPB B1_N A1 A2 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A2	A2
* A1	A1
* B1_N	B1_N
* VPB	VPB
* VNB	VNB
MM1001 N_VGND_M1001_d N_B1_N_M1001_g N_A_29_424#_M1001_s VNB NLOWVT L=0.15
+ W=0.55 AD=0.14575 AS=0.14575 PD=1.08295 PS=1.63 NRD=35.448 NRS=0 M=1 R=3.66667
+ SA=75000.2 SB=75001.8 A=0.0825 P=1.4 MULT=1
MM1005 N_Y_M1005_d N_A_29_424#_M1005_g N_VGND_M1001_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1961 PD=1.02 PS=1.45705 NRD=0 NRS=14.592 M=1 R=4.93333
+ SA=75000.7 SB=75001.1 A=0.111 P=1.78 MULT=1
MM1000 A_437_74# N_A1_M1000_g N_Y_M1005_d VNB NLOWVT L=0.15 W=0.74 AD=0.1184
+ AS=0.1036 PD=1.06 PS=1.02 NRD=17.016 NRS=0 M=1 R=4.93333 SA=75001.1 SB=75000.7
+ A=0.111 P=1.78 MULT=1
MM1007 N_VGND_M1007_d N_A2_M1007_g A_437_74# VNB NLOWVT L=0.15 W=0.74 AD=0.2109
+ AS=0.1184 PD=2.05 PS=1.06 NRD=0 NRS=17.016 M=1 R=4.93333 SA=75001.6 SB=75000.2
+ A=0.111 P=1.78 MULT=1
MM1002 N_VPWR_M1002_d N_B1_N_M1002_g N_A_29_424#_M1002_s VPB PSHORT L=0.15
+ W=0.84 AD=0.231 AS=0.231 PD=2.23 PS=2.23 NRD=2.3443 NRS=2.3443 M=1 R=5.6
+ SA=75000.2 SB=75000.2 A=0.126 P=1.98 MULT=1
MM1003 N_A_348_368#_M1003_d N_A_29_424#_M1003_g N_Y_M1003_s VPB PSHORT L=0.15
+ W=1.12 AD=0.168 AS=0.308 PD=1.42 PS=2.79 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75001.1 A=0.168 P=2.54 MULT=1
MM1006 N_VPWR_M1006_d N_A1_M1006_g N_A_348_368#_M1003_d VPB PSHORT L=0.15 W=1.12
+ AD=0.1848 AS=0.168 PD=1.45 PS=1.42 NRD=4.3931 NRS=1.7533 M=1 R=7.46667
+ SA=75000.6 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1004 N_A_348_368#_M1004_d N_A2_M1004_g N_VPWR_M1006_d VPB PSHORT L=0.15 W=1.12
+ AD=0.308 AS=0.1848 PD=2.79 PS=1.45 NRD=1.7533 NRS=4.3931 M=1 R=7.46667
+ SA=75001.1 SB=75000.2 A=0.168 P=2.54 MULT=1
DX8_noxref VNB VPB NWDIODE A=6.9564 P=11.2
*
.include "sky130_fd_sc_hs__a21boi_1.pxi.spice"
*
.ends
*
*
