* NGSPICE file created from sky130_fd_sc_hs__xor3_4.ext - technology: sky130A

.subckt sky130_fd_sc_hs__xor3_4 A B C VGND VNB VPB VPWR X
M1000 X a_1218_388# VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=6.72e+11p pd=5.68e+06u as=2.2388e+12p ps=1.511e+07u
M1001 VGND C a_1155_284# VNB nlowvt w=420000u l=150000u
+  ad=1.6131e+12p pd=1.223e+07u as=2.121e+11p ps=1.85e+06u
M1002 a_74_294# a_397_320# a_416_118# VPB pshort w=840000u l=150000u
+  ad=9.166e+11p pd=5.75e+06u as=6.8745e+11p ps=5.04e+06u
M1003 VPWR B a_397_320# VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=3.304e+11p ps=2.83e+06u
M1004 a_416_118# B a_27_118# VPB pshort w=640000u l=150000u
+  ad=0p pd=0u as=5.9475e+11p ps=5.02e+06u
M1005 VPWR a_1218_388# X VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_74_294# A VPWR VPB pshort w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VGND a_1218_388# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=4.144e+11p ps=4.08e+06u
M1008 VPWR a_74_294# a_27_118# VPB pshort w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_1218_388# a_1155_284# a_416_118# VPB pshort w=840000u l=150000u
+  ad=4.452e+11p pd=2.74e+06u as=0p ps=0u
M1010 VPWR C a_1155_284# VPB pshort w=640000u l=150000u
+  ad=0p pd=0u as=1.888e+11p ps=1.87e+06u
M1011 a_27_118# a_397_320# a_323_392# VPB pshort w=640000u l=150000u
+  ad=0p pd=0u as=5.532e+11p ps=4.72e+06u
M1012 VGND a_74_294# a_27_118# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=4.264e+11p ps=4.03e+06u
M1013 X a_1218_388# VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_323_392# B a_27_118# VNB nlowvt w=640000u l=150000u
+  ad=4.6775e+11p pd=4.06e+06u as=0p ps=0u
M1015 VPWR a_1218_388# X VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_1218_388# a_1155_284# a_323_392# VNB nlowvt w=640000u l=150000u
+  ad=3.392e+11p pd=2.34e+06u as=0p ps=0u
M1017 X a_1218_388# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 X a_1218_388# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_416_118# B a_74_294# VNB nlowvt w=640000u l=150000u
+  ad=3.899e+11p pd=3.83e+06u as=7.264e+11p ps=4.83e+06u
M1020 a_323_392# C a_1218_388# VPB pshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_416_118# C a_1218_388# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_27_118# a_397_320# a_416_118# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_323_392# B a_74_294# VPB pshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 VGND a_1218_388# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 a_74_294# A VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 VGND B a_397_320# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.072e+11p ps=2.04e+06u
M1027 a_74_294# a_397_320# a_323_392# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

