* File: sky130_fd_sc_hs__sdfrbp_1.spice
* Created: Tue Sep  1 20:22:19 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hs__sdfrbp_1.pex.spice"
.subckt sky130_fd_sc_hs__sdfrbp_1  VNB VPB SCE D SCD RESET_B CLK VPWR Q_N Q VGND
* 
* VGND	VGND
* Q	Q
* Q_N	Q_N
* VPWR	VPWR
* CLK	CLK
* RESET_B	RESET_B
* SCD	SCD
* D	D
* SCE	SCE
* VPB	VPB
* VNB	VNB
MM1040 N_VGND_M1040_d N_SCE_M1040_g N_A_27_74#_M1040_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.1197 AS=0.1197 PD=1.41 PS=1.41 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1021 noxref_26 N_A_27_74#_M1021_g N_noxref_25_M1021_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.07455 AS=0.1197 PD=0.775 PS=1.41 NRD=34.992 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75002.2 A=0.063 P=1.14 MULT=1
MM1000 N_A_413_90#_M1000_d N_D_M1000_g noxref_26 VNB NLOWVT L=0.15 W=0.42
+ AD=0.107537 AS=0.07455 PD=0.965 PS=0.775 NRD=65.712 NRS=34.992 M=1 R=2.8
+ SA=75000.7 SB=75001.7 A=0.063 P=1.14 MULT=1
MM1033 noxref_27 N_SCE_M1033_g N_A_413_90#_M1000_d VNB NLOWVT L=0.15 W=0.42
+ AD=0.0504 AS=0.107537 PD=0.66 PS=0.965 NRD=18.564 NRS=0 M=1 R=2.8 SA=75001.3
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1015 N_noxref_25_M1015_d N_SCD_M1015_g noxref_27 VNB NLOWVT L=0.15 W=0.42
+ AD=0.0858375 AS=0.0504 PD=0.855 PS=0.66 NRD=22.848 NRS=18.564 M=1 R=2.8
+ SA=75001.7 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1034 N_VGND_M1034_d N_RESET_B_M1034_g N_noxref_25_M1015_d VNB NLOWVT L=0.15
+ W=0.42 AD=0.1365 AS=0.0858375 PD=1.49 PS=0.855 NRD=11.424 NRS=8.568 M=1 R=2.8
+ SA=75002.1 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1035 N_VGND_M1035_d N_CLK_M1035_g N_A_850_74#_M1035_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.2109 PD=1.02 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1036 N_A_1023_74#_M1036_d N_A_850_74#_M1036_g N_VGND_M1035_d VNB NLOWVT L=0.15
+ W=0.74 AD=0.2109 AS=0.1036 PD=2.05 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.6 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1012 N_A_1221_97#_M1012_d N_A_850_74#_M1012_g N_A_413_90#_M1012_s VNB NLOWVT
+ L=0.15 W=0.42 AD=0.0735 AS=0.1197 PD=0.77 PS=1.41 NRD=19.992 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75004.5 A=0.063 P=1.14 MULT=1
MM1004 A_1321_97# N_A_1023_74#_M1004_g N_A_1221_97#_M1012_d VNB NLOWVT L=0.15
+ W=0.42 AD=0.0504 AS=0.0735 PD=0.66 PS=0.77 NRD=18.564 NRS=0 M=1 R=2.8
+ SA=75000.7 SB=75004 A=0.063 P=1.14 MULT=1
MM1016 A_1399_97# N_A_1369_71#_M1016_g A_1321_97# VNB NLOWVT L=0.15 W=0.42
+ AD=0.0504 AS=0.0504 PD=0.66 PS=0.66 NRD=18.564 NRS=18.564 M=1 R=2.8 SA=75001.1
+ SB=75003.6 A=0.063 P=1.14 MULT=1
MM1017 N_VGND_M1017_d N_RESET_B_M1017_g A_1399_97# VNB NLOWVT L=0.15 W=0.42
+ AD=0.190317 AS=0.0504 PD=1.25604 PS=0.66 NRD=113.748 NRS=18.564 M=1 R=2.8
+ SA=75001.5 SB=75003.2 A=0.063 P=1.14 MULT=1
MM1041 N_A_1369_71#_M1041_d N_A_1221_97#_M1041_g N_VGND_M1017_d VNB NLOWVT
+ L=0.15 W=0.64 AD=0.0896 AS=0.290008 PD=0.92 PS=1.91396 NRD=0 NRS=74.64 M=1
+ R=4.26667 SA=75001.7 SB=75002.1 A=0.096 P=1.58 MULT=1
MM1030 N_A_1747_74#_M1030_d N_A_1023_74#_M1030_g N_A_1369_71#_M1041_d VNB NLOWVT
+ L=0.15 W=0.64 AD=0.272845 AS=0.0896 PD=1.91396 PS=0.92 NRD=92.808 NRS=0 M=1
+ R=4.26667 SA=75002.2 SB=75001.7 A=0.096 P=1.58 MULT=1
MM1013 A_1966_74# N_A_850_74#_M1013_g N_A_1747_74#_M1030_d VNB NLOWVT L=0.15
+ W=0.42 AD=0.0441 AS=0.179055 PD=0.63 PS=1.25604 NRD=14.28 NRS=48.564 M=1 R=2.8
+ SA=75003.4 SB=75001.4 A=0.063 P=1.14 MULT=1
MM1005 N_VGND_M1005_d N_A_2008_48#_M1005_g A_1966_74# VNB NLOWVT L=0.15 W=0.42
+ AD=0.0588 AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75003.8
+ SB=75001 A=0.063 P=1.14 MULT=1
MM1007 A_2124_74# N_RESET_B_M1007_g N_VGND_M1005_d VNB NLOWVT L=0.15 W=0.42
+ AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75004.2
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1010 N_A_2008_48#_M1010_d N_A_1747_74#_M1010_g A_2124_74# VNB NLOWVT L=0.15
+ W=0.42 AD=0.1197 AS=0.0441 PD=1.41 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8
+ SA=75004.6 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1008 N_Q_N_M1008_d N_A_1747_74#_M1008_g N_VGND_M1008_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.2072 AS=0.3159 PD=2.04 PS=2.57 NRD=0 NRS=60.3 M=1 R=4.93333
+ SA=75000.3 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1002 N_VGND_M1002_d N_A_1747_74#_M1002_g N_A_2513_424#_M1002_s VNB NLOWVT
+ L=0.15 W=0.55 AD=0.101196 AS=0.14575 PD=0.92093 PS=1.63 NRD=13.632 NRS=0 M=1
+ R=3.66667 SA=75000.2 SB=75000.7 A=0.0825 P=1.4 MULT=1
MM1039 N_Q_M1039_d N_A_2513_424#_M1039_g N_VGND_M1002_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.136154 PD=2.05 PS=1.23907 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.6
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1027 N_VPWR_M1027_d N_SCE_M1027_g N_A_27_74#_M1027_s VPB PSHORT L=0.15 W=0.64
+ AD=0.112 AS=0.5792 PD=0.99 PS=3.09 NRD=18.4589 NRS=3.0732 M=1 R=4.26667
+ SA=75000.8 SB=75002.7 A=0.096 P=1.58 MULT=1
MM1024 A_338_464# N_SCE_M1024_g N_VPWR_M1027_d VPB PSHORT L=0.15 W=0.64
+ AD=0.0864 AS=0.112 PD=0.91 PS=0.99 NRD=24.625 NRS=3.0732 M=1 R=4.26667
+ SA=75001.3 SB=75002.2 A=0.096 P=1.58 MULT=1
MM1009 N_A_413_90#_M1009_d N_D_M1009_g A_338_464# VPB PSHORT L=0.15 W=0.64
+ AD=0.096 AS=0.0864 PD=0.94 PS=0.91 NRD=3.0732 NRS=24.625 M=1 R=4.26667
+ SA=75001.8 SB=75001.8 A=0.096 P=1.58 MULT=1
MM1014 A_512_464# N_A_27_74#_M1014_g N_A_413_90#_M1009_d VPB PSHORT L=0.15
+ W=0.64 AD=0.1248 AS=0.096 PD=1.03 PS=0.94 NRD=43.0839 NRS=3.0732 M=1 R=4.26667
+ SA=75002.2 SB=75001.3 A=0.096 P=1.58 MULT=1
MM1032 N_VPWR_M1032_d N_SCD_M1032_g A_512_464# VPB PSHORT L=0.15 W=0.64
+ AD=0.1344 AS=0.1248 PD=1.06 PS=1.03 NRD=7.683 NRS=43.0839 M=1 R=4.26667
+ SA=75002.7 SB=75000.8 A=0.096 P=1.58 MULT=1
MM1020 N_A_413_90#_M1020_d N_RESET_B_M1020_g N_VPWR_M1032_d VPB PSHORT L=0.15
+ W=0.64 AD=0.1888 AS=0.1344 PD=1.87 PS=1.06 NRD=3.0732 NRS=35.3812 M=1
+ R=4.26667 SA=75003.3 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1025 N_VPWR_M1025_d N_CLK_M1025_g N_A_850_74#_M1025_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.3304 PD=1.42 PS=2.83 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1038 N_A_1023_74#_M1038_d N_A_850_74#_M1038_g N_VPWR_M1025_d VPB PSHORT L=0.15
+ W=1.12 AD=0.3192 AS=0.168 PD=2.81 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.7 SB=75000.2 A=0.168 P=2.54 MULT=1
MM1028 N_A_1221_97#_M1028_d N_A_1023_74#_M1028_g N_A_413_90#_M1028_s VPB PSHORT
+ L=0.15 W=0.42 AD=0.063 AS=0.1197 PD=0.72 PS=1.41 NRD=4.6886 NRS=4.6886 M=1
+ R=2.8 SA=75000.2 SB=75001.6 A=0.063 P=1.14 MULT=1
MM1037 A_1328_463# N_A_850_74#_M1037_g N_A_1221_97#_M1028_d VPB PSHORT L=0.15
+ W=0.42 AD=0.0504 AS=0.063 PD=0.66 PS=0.72 NRD=30.4759 NRS=4.6886 M=1 R=2.8
+ SA=75000.7 SB=75001.2 A=0.063 P=1.14 MULT=1
MM1018 N_VPWR_M1018_d N_A_1369_71#_M1018_g A_1328_463# VPB PSHORT L=0.15 W=0.42
+ AD=0.126225 AS=0.0504 PD=1.105 PS=0.66 NRD=115.166 NRS=30.4759 M=1 R=2.8
+ SA=75001.1 SB=75000.8 A=0.063 P=1.14 MULT=1
MM1011 N_A_1221_97#_M1011_d N_RESET_B_M1011_g N_VPWR_M1018_d VPB PSHORT L=0.15
+ W=0.42 AD=0.1197 AS=0.126225 PD=1.41 PS=1.105 NRD=4.6886 NRS=115.166 M=1 R=2.8
+ SA=75001.6 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1019 N_A_1369_71#_M1019_d N_A_1221_97#_M1019_g N_VPWR_M1019_s VPB PSHORT
+ L=0.15 W=1 AD=0.15 AS=0.285 PD=1.3 PS=2.57 NRD=1.9503 NRS=1.9503 M=1 R=6.66667
+ SA=75000.2 SB=75001.5 A=0.15 P=2.3 MULT=1
MM1023 N_A_1747_74#_M1023_d N_A_850_74#_M1023_g N_A_1369_71#_M1019_d VPB PSHORT
+ L=0.15 W=1 AD=0.292148 AS=0.15 PD=2.47183 PS=1.3 NRD=23.3051 NRS=1.9503 M=1
+ R=6.66667 SA=75000.7 SB=75001.1 A=0.15 P=2.3 MULT=1
MM1001 A_1969_489# N_A_1023_74#_M1001_g N_A_1747_74#_M1023_d VPB PSHORT L=0.15
+ W=0.42 AD=0.0504 AS=0.122702 PD=0.66 PS=1.03817 NRD=30.4759 NRS=4.6886 M=1
+ R=2.8 SA=75001.1 SB=75002.4 A=0.063 P=1.14 MULT=1
MM1003 N_VPWR_M1003_d N_A_2008_48#_M1003_g A_1969_489# VPB PSHORT L=0.15 W=0.42
+ AD=0.117862 AS=0.0504 PD=1.01 PS=0.66 NRD=49.2303 NRS=30.4759 M=1 R=2.8
+ SA=75001.4 SB=75002 A=0.063 P=1.14 MULT=1
MM1026 N_A_2008_48#_M1026_d N_RESET_B_M1026_g N_VPWR_M1003_d VPB PSHORT L=0.15
+ W=0.42 AD=0.063 AS=0.117862 PD=0.72 PS=1.01 NRD=4.6886 NRS=51.5943 M=1 R=2.8
+ SA=75002.1 SB=75001.3 A=0.063 P=1.14 MULT=1
MM1031 N_VPWR_M1031_d N_A_1747_74#_M1031_g N_A_2008_48#_M1026_d VPB PSHORT
+ L=0.15 W=0.42 AD=0.121609 AS=0.063 PD=0.9 PS=0.72 NRD=75.0373 NRS=4.6886 M=1
+ R=2.8 SA=75002.5 SB=75000.9 A=0.063 P=1.14 MULT=1
MM1006 N_Q_N_M1006_d N_A_1747_74#_M1006_g N_VPWR_M1031_d VPB PSHORT L=0.15
+ W=1.12 AD=0.3304 AS=0.324291 PD=2.83 PS=2.4 NRD=1.7533 NRS=12.017 M=1
+ R=7.46667 SA=75001.4 SB=75000.2 A=0.168 P=2.54 MULT=1
MM1022 N_VPWR_M1022_d N_A_1747_74#_M1022_g N_A_2513_424#_M1022_s VPB PSHORT
+ L=0.15 W=0.84 AD=0.1662 AS=0.231 PD=1.27714 PS=2.23 NRD=10.5395 NRS=2.3443 M=1
+ R=5.6 SA=75000.2 SB=75000.7 A=0.126 P=1.98 MULT=1
MM1029 N_Q_M1029_d N_A_2513_424#_M1029_g N_VPWR_M1022_d VPB PSHORT L=0.15 W=1.12
+ AD=0.308 AS=0.2216 PD=2.79 PS=1.70286 NRD=1.7533 NRS=5.8509 M=1 R=7.46667
+ SA=75000.6 SB=75000.2 A=0.168 P=2.54 MULT=1
DX42_noxref VNB VPB NWDIODE A=26.8347 P=32.53
*
.include "sky130_fd_sc_hs__sdfrbp_1.pxi.spice"
*
.ends
*
*
