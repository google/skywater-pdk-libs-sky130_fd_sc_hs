* File: sky130_fd_sc_hs__mux4_2.spice
* Created: Thu Aug 27 20:49:43 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hs__mux4_2.pex.spice"
.subckt sky130_fd_sc_hs__mux4_2  VNB VPB S0 A1 A0 A3 A2 S1 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* S1	S1
* A2	A2
* A3	A3
* A0	A0
* A1	A1
* S0	S0
* VPB	VPB
* VNB	VNB
MM1001 N_VGND_M1001_d N_S0_M1001_g N_A_31_94#_M1001_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.172012 AS=0.1824 PD=1.18261 PS=1.85 NRD=48.276 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75005.8 A=0.096 P=1.58 MULT=1
MM1013 A_255_74# N_A1_M1013_g N_VGND_M1001_d VNB NLOWVT L=0.15 W=0.74 AD=0.0888
+ AS=0.198888 PD=0.98 PS=1.36739 NRD=10.536 NRS=0 M=1 R=4.93333 SA=75000.8
+ SB=75005.1 A=0.111 P=1.78 MULT=1
MM1010 N_A_333_74#_M1010_d N_S0_M1010_g A_255_74# VNB NLOWVT L=0.15 W=0.74
+ AD=0.2664 AS=0.0888 PD=1.46 PS=0.98 NRD=44.592 NRS=10.536 M=1 R=4.93333
+ SA=75001.2 SB=75004.7 A=0.111 P=1.78 MULT=1
MM1014 A_507_74# N_A_31_94#_M1014_g N_A_333_74#_M1010_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.2886 AS=0.2664 PD=1.52 PS=1.46 NRD=54.324 NRS=26.748 M=1 R=4.93333
+ SA=75002.1 SB=75003.8 A=0.111 P=1.78 MULT=1
MM1023 N_VGND_M1023_d N_A0_M1023_g A_507_74# VNB NLOWVT L=0.15 W=0.74 AD=0.1998
+ AS=0.2886 PD=1.28 PS=1.52 NRD=7.296 NRS=54.324 M=1 R=4.93333 SA=75003
+ SB=75002.9 A=0.111 P=1.78 MULT=1
MM1019 A_831_74# N_A3_M1019_g N_VGND_M1023_d VNB NLOWVT L=0.15 W=0.74 AD=0.0888
+ AS=0.1998 PD=0.98 PS=1.28 NRD=10.536 NRS=34.86 M=1 R=4.93333 SA=75003.7
+ SB=75002.2 A=0.111 P=1.78 MULT=1
MM1016 N_A_909_74#_M1016_d N_S0_M1016_g A_831_74# VNB NLOWVT L=0.15 W=0.74
+ AD=0.1998 AS=0.0888 PD=1.28 PS=0.98 NRD=27.564 NRS=10.536 M=1 R=4.93333
+ SA=75004.1 SB=75001.8 A=0.111 P=1.78 MULT=1
MM1005 A_1047_74# N_A_31_94#_M1005_g N_A_909_74#_M1016_d VNB NLOWVT L=0.15
+ W=0.74 AD=0.2886 AS=0.1998 PD=1.52 PS=1.28 NRD=54.324 NRS=14.592 M=1 R=4.93333
+ SA=75004.8 SB=75001.1 A=0.111 P=1.78 MULT=1
MM1011 N_VGND_M1011_d N_A2_M1011_g A_1047_74# VNB NLOWVT L=0.15 W=0.74 AD=0.2072
+ AS=0.2886 PD=2.04 PS=1.52 NRD=0 NRS=54.324 M=1 R=4.93333 SA=75005.7 SB=75000.2
+ A=0.111 P=1.78 MULT=1
MM1009 N_A_1429_74#_M1009_d N_S1_M1009_g N_A_909_74#_M1009_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.151475 AS=0.2072 PD=1.325 PS=2.04 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75000.6 A=0.111 P=1.78 MULT=1
MM1006 N_A_333_74#_M1006_d N_A_1500_94#_M1006_g N_A_1429_74#_M1009_d VNB NLOWVT
+ L=0.15 W=0.74 AD=0.2109 AS=0.151475 PD=2.05 PS=1.325 NRD=0 NRS=24.264 M=1
+ R=4.93333 SA=75000.5 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1008 N_VGND_M1008_d N_S1_M1008_g N_A_1500_94#_M1008_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.232858 AS=0.276725 PD=1.37275 PS=2.15 NRD=86.712 NRS=26.244 M=1 R=4.26667
+ SA=75000.4 SB=75001.5 A=0.096 P=1.58 MULT=1
MM1021 N_X_M1021_d N_A_1429_74#_M1021_g N_VGND_M1008_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.269242 PD=1.02 PS=1.58725 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.1
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1025 N_X_M1021_d N_A_1429_74#_M1025_g N_VGND_M1025_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.2109 PD=1.02 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.5
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1007 N_VPWR_M1007_d N_S0_M1007_g N_A_31_94#_M1007_s VPB PSHORT L=0.15 W=1
+ AD=0.225 AS=0.295 PD=1.45 PS=2.59 NRD=11.8003 NRS=1.9503 M=1 R=6.66667
+ SA=75000.2 SB=75005.7 A=0.15 P=2.3 MULT=1
MM1002 A_264_392# N_A1_M1002_g N_VPWR_M1007_d VPB PSHORT L=0.15 W=1 AD=0.45
+ AS=0.225 PD=1.9 PS=1.45 NRD=77.7953 NRS=21.67 M=1 R=6.66667 SA=75000.8
+ SB=75005.1 A=0.15 P=2.3 MULT=1
MM1000 N_A_333_74#_M1000_d N_A_31_94#_M1000_g A_264_392# VPB PSHORT L=0.15 W=1
+ AD=0.285 AS=0.45 PD=1.57 PS=1.9 NRD=29.5303 NRS=77.7953 M=1 R=6.66667
+ SA=75001.9 SB=75004 A=0.15 P=2.3 MULT=1
MM1020 A_618_392# N_S0_M1020_g N_A_333_74#_M1000_d VPB PSHORT L=0.15 W=1
+ AD=0.135 AS=0.285 PD=1.27 PS=1.57 NRD=15.7403 NRS=27.5603 M=1 R=6.66667
+ SA=75002.6 SB=75003.3 A=0.15 P=2.3 MULT=1
MM1004 N_VPWR_M1004_d N_A0_M1004_g A_618_392# VPB PSHORT L=0.15 W=1 AD=0.27
+ AS=0.135 PD=1.54 PS=1.27 NRD=25.5903 NRS=15.7403 M=1 R=6.66667 SA=75003
+ SB=75002.9 A=0.15 P=2.3 MULT=1
MM1003 A_840_392# N_A3_M1003_g N_VPWR_M1004_d VPB PSHORT L=0.15 W=1 AD=0.36
+ AS=0.27 PD=1.72 PS=1.54 NRD=60.0653 NRS=25.5903 M=1 R=6.66667 SA=75003.7
+ SB=75002.2 A=0.15 P=2.3 MULT=1
MM1015 N_A_909_74#_M1015_d N_A_31_94#_M1015_g A_840_392# VPB PSHORT L=0.15 W=1
+ AD=0.27 AS=0.36 PD=1.54 PS=1.72 NRD=25.5903 NRS=60.0653 M=1 R=6.66667
+ SA=75004.6 SB=75001.3 A=0.15 P=2.3 MULT=1
MM1022 A_1152_392# N_S0_M1022_g N_A_909_74#_M1015_d VPB PSHORT L=0.15 W=1
+ AD=0.135 AS=0.27 PD=1.27 PS=1.54 NRD=15.7403 NRS=25.5903 M=1 R=6.66667
+ SA=75005.3 SB=75000.6 A=0.15 P=2.3 MULT=1
MM1026 N_VPWR_M1026_d N_A2_M1026_g A_1152_392# VPB PSHORT L=0.15 W=1 AD=0.295
+ AS=0.135 PD=2.59 PS=1.27 NRD=1.9503 NRS=15.7403 M=1 R=6.66667 SA=75005.7
+ SB=75000.2 A=0.15 P=2.3 MULT=1
MM1012 N_A_1429_74#_M1012_d N_S1_M1012_g N_A_333_74#_M1012_s VPB PSHORT L=0.15
+ W=1 AD=0.15 AS=0.32 PD=1.3 PS=2.64 NRD=1.9503 NRS=4.9053 M=1 R=6.66667
+ SA=75000.2 SB=75000.7 A=0.15 P=2.3 MULT=1
MM1017 N_A_909_74#_M1017_d N_A_1500_94#_M1017_g N_A_1429_74#_M1012_d VPB PSHORT
+ L=0.15 W=1 AD=0.29 AS=0.15 PD=2.58 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=6.66667
+ SA=75000.7 SB=75000.2 A=0.15 P=2.3 MULT=1
MM1018 N_VPWR_M1018_d N_S1_M1018_g N_A_1500_94#_M1018_s VPB PSHORT L=0.15 W=1
+ AD=0.363113 AS=0.425 PD=1.75 PS=2.85 NRD=87.9802 NRS=28.565 M=1 R=6.66667
+ SA=75000.3 SB=75001.5 A=0.15 P=2.3 MULT=1
MM1024 N_X_M1024_d N_A_1429_74#_M1024_g N_VPWR_M1018_d VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.406687 PD=1.42 PS=1.96 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.1 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1027 N_X_M1024_d N_A_1429_74#_M1027_g N_VPWR_M1027_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.3248 PD=1.42 PS=2.82 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.6 SB=75000.2 A=0.168 P=2.54 MULT=1
DX28_noxref VNB VPB NWDIODE A=20.2119 P=25.8
c_164 VPB 0 5.38206e-20 $X=0 $Y=3.085
c_1316 A_507_74# 0 1.87351e-19 $X=2.535 $Y=0.37
*
.include "sky130_fd_sc_hs__mux4_2.pxi.spice"
*
.ends
*
*
