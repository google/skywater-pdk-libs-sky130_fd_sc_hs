* File: sky130_fd_sc_hs__dlxtp_1.spice
* Created: Thu Aug 27 20:42:59 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hs__dlxtp_1.pex.spice"
.subckt sky130_fd_sc_hs__dlxtp_1  VNB VPB D GATE VPWR Q VGND
* 
* VGND	VGND
* Q	Q
* VPWR	VPWR
* GATE	GATE
* D	D
* VPB	VPB
* VNB	VNB
MM1008 N_A_116_424#_M1008_d N_D_M1008_g N_VGND_M1008_s VNB NLOWVT L=0.15 W=0.55
+ AD=0.1815 AS=0.1705 PD=1.76 PS=1.72 NRD=9.816 NRS=5.448 M=1 R=3.66667
+ SA=75000.2 SB=75000.3 A=0.0825 P=1.4 MULT=1
MM1000 N_VGND_M1000_d N_A_116_424#_M1000_g N_A_239_85#_M1000_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.250643 AS=0.2238 PD=1.89466 PS=2.14 NRD=4.044 NRS=7.296 M=1
+ R=4.93333 SA=75000.2 SB=75001.3 A=0.111 P=1.78 MULT=1
MM1011 A_514_149# N_A_386_326#_M1011_g N_VGND_M1000_d VNB NLOWVT L=0.15 W=0.42
+ AD=0.0504 AS=0.142257 PD=0.66 PS=1.07534 NRD=18.564 NRS=125.712 M=1 R=2.8
+ SA=75001.1 SB=75001.2 A=0.063 P=1.14 MULT=1
MM1006 N_A_592_149#_M1006_d N_A_562_123#_M1006_g A_514_149# VNB NLOWVT L=0.15
+ W=0.42 AD=0.0996776 AS=0.0504 PD=0.872586 PS=0.66 NRD=24.276 NRS=18.564 M=1
+ R=2.8 SA=75001.5 SB=75000.8 A=0.063 P=1.14 MULT=1
MM1014 N_A_239_85#_M1014_d N_A_685_59#_M1014_g N_A_592_149#_M1006_d VNB NLOWVT
+ L=0.15 W=0.74 AD=0.222 AS=0.175622 PD=2.08 PS=1.53741 NRD=0.804 NRS=16.212 M=1
+ R=4.93333 SA=75001.3 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1010 N_VGND_M1010_d N_A_592_149#_M1010_g N_A_386_326#_M1010_s VNB NLOWVT
+ L=0.15 W=0.74 AD=0.19615 AS=0.2109 PD=1.41 PS=2.05 NRD=34.056 NRS=0 M=1
+ R=4.93333 SA=75000.2 SB=75000.8 A=0.111 P=1.78 MULT=1
MM1005 N_A_685_59#_M1005_d N_A_562_123#_M1005_g N_VGND_M1010_d VNB NLOWVT L=0.15
+ W=0.74 AD=0.2109 AS=0.19615 PD=2.05 PS=1.41 NRD=0 NRS=34.056 M=1 R=4.93333
+ SA=75000.8 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1015 N_VGND_M1015_d N_GATE_M1015_g N_A_562_123#_M1015_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.261625 AS=0.222 PD=1.545 PS=2.08 NRD=48.408 NRS=1.62 M=1 R=4.93333
+ SA=75000.2 SB=75000.9 A=0.111 P=1.78 MULT=1
MM1007 N_Q_M1007_d N_A_386_326#_M1007_g N_VGND_M1015_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.261625 PD=2.05 PS=1.545 NRD=0 NRS=48.408 M=1 R=4.93333
+ SA=75000.9 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1013 N_A_116_424#_M1013_d N_D_M1013_g N_VPWR_M1013_s VPB PSHORT L=0.15 W=0.84
+ AD=0.2478 AS=0.2478 PD=2.27 PS=2.27 NRD=2.3443 NRS=2.3443 M=1 R=5.6 SA=75000.2
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1012 N_VPWR_M1012_d N_A_116_424#_M1012_g N_A_229_392#_M1012_s VPB PSHORT
+ L=0.15 W=1 AD=0.272658 AS=0.295 PD=2.39437 PS=2.59 NRD=42.8672 NRS=1.9503 M=1
+ R=6.66667 SA=75000.2 SB=75000.4 A=0.15 P=2.3 MULT=1
MM1009 N_A_419_392#_M1009_d N_A_386_326#_M1009_g N_VPWR_M1012_d VPB PSHORT
+ L=0.15 W=0.42 AD=0.1239 AS=0.114517 PD=1.43 PS=1.00563 NRD=4.6886 NRS=102.085
+ M=1 R=2.8 SA=75000.7 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1003 N_A_592_149#_M1003_d N_A_562_123#_M1003_g N_A_229_392#_M1003_s VPB PSHORT
+ L=0.15 W=1 AD=0.234366 AS=0.295 PD=1.9507 PS=2.59 NRD=1.9503 NRS=1.9503 M=1
+ R=6.66667 SA=75000.2 SB=75000.5 A=0.15 P=2.3 MULT=1
MM1002 N_A_419_392#_M1002_d N_A_685_59#_M1002_g N_A_592_149#_M1003_d VPB PSHORT
+ L=0.15 W=0.42 AD=0.19295 AS=0.0984338 PD=1.83 PS=0.819296 NRD=46.886
+ NRS=84.119 M=1 R=2.8 SA=75000.8 SB=75000.3 A=0.063 P=1.14 MULT=1
MM1016 N_VPWR_M1016_d N_A_592_149#_M1016_g N_A_386_326#_M1016_s VPB PSHORT
+ L=0.15 W=1.12 AD=0.3444 AS=0.3696 PD=2.21714 PS=2.9 NRD=44.4038 NRS=5.2599 M=1
+ R=7.46667 SA=75000.3 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1017 N_A_685_59#_M1017_d N_A_562_123#_M1017_g N_VPWR_M1016_d VPB PSHORT L=0.15
+ W=0.84 AD=0.2478 AS=0.2583 PD=2.27 PS=1.66286 NRD=2.3443 NRS=59.1985 M=1 R=5.6
+ SA=75000.9 SB=75000.2 A=0.126 P=1.98 MULT=1
MM1001 N_VPWR_M1001_d N_GATE_M1001_g N_A_562_123#_M1001_s VPB PSHORT L=0.15
+ W=0.84 AD=0.198 AS=0.2478 PD=1.33286 PS=2.27 NRD=22.261 NRS=2.3443 M=1 R=5.6
+ SA=75000.2 SB=75000.8 A=0.126 P=1.98 MULT=1
MM1004 N_Q_M1004_d N_A_386_326#_M1004_g N_VPWR_M1001_d VPB PSHORT L=0.15 W=1.12
+ AD=0.3304 AS=0.264 PD=2.83 PS=1.77714 NRD=1.7533 NRS=10.5395 M=1 R=7.46667
+ SA=75000.7 SB=75000.2 A=0.168 P=2.54 MULT=1
DX18_noxref VNB VPB NWDIODE A=15.2636 P=20.15
*
.include "sky130_fd_sc_hs__dlxtp_1.pxi.spice"
*
.ends
*
*
