* File: sky130_fd_sc_hs__nand2b_2.spice
* Created: Tue Sep  1 20:09:00 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hs__nand2b_2.pex.spice"
.subckt sky130_fd_sc_hs__nand2b_2  VNB VPB A_N B VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* B	B
* A_N	A_N
* VPB	VPB
* VNB	VNB
MM1008 N_VGND_M1008_d N_A_N_M1008_g N_A_27_74#_M1008_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.16675 AS=0.1824 PD=1.81 PS=1.85 NRD=0 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75000.2 A=0.096 P=1.58 MULT=1
MM1005 N_Y_M1005_d N_A_27_74#_M1005_g N_A_242_74#_M1005_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.20635 PD=1.02 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75001.5 A=0.111 P=1.78 MULT=1
MM1009 N_Y_M1005_d N_A_27_74#_M1009_g N_A_242_74#_M1009_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.6 SB=75001.1 A=0.111 P=1.78 MULT=1
MM1000 N_VGND_M1000_d N_B_M1000_g N_A_242_74#_M1009_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.10545 AS=0.1036 PD=1.025 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.1
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1006 N_VGND_M1000_d N_B_M1006_g N_A_242_74#_M1006_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.10545 AS=0.2109 PD=1.025 PS=2.05 NRD=0.804 NRS=0 M=1 R=4.93333 SA=75001.5
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1003 N_VPWR_M1003_d N_A_N_M1003_g N_A_27_74#_M1003_s VPB PSHORT L=0.15 W=1
+ AD=0.435189 AS=0.295 PD=1.85849 PS=2.59 NRD=42.3353 NRS=1.9503 M=1 R=6.66667
+ SA=75000.2 SB=75002.6 A=0.15 P=2.3 MULT=1
MM1001 N_Y_M1001_d N_A_27_74#_M1001_g N_VPWR_M1003_d VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.487411 PD=1.42 PS=2.08151 NRD=1.7533 NRS=62.8627 M=1 R=7.46667
+ SA=75001.1 SB=75001.6 A=0.168 P=2.54 MULT=1
MM1002 N_Y_M1001_d N_A_27_74#_M1002_g N_VPWR_M1002_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.6 SB=75001.1 A=0.168 P=2.54 MULT=1
MM1004 N_Y_M1004_d N_B_M1004_g N_VPWR_M1002_s VPB PSHORT L=0.15 W=1.12 AD=0.168
+ AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667 SA=75002
+ SB=75000.7 A=0.168 P=2.54 MULT=1
MM1007 N_Y_M1004_d N_B_M1007_g N_VPWR_M1007_s VPB PSHORT L=0.15 W=1.12 AD=0.168
+ AS=0.3304 PD=1.42 PS=2.83 NRD=1.7533 NRS=1.7533 M=1 R=7.46667 SA=75002.5
+ SB=75000.2 A=0.168 P=2.54 MULT=1
DX10_noxref VNB VPB NWDIODE A=6.9564 P=11.2
c_70 VPB 0 1.91961e-19 $X=0 $Y=3.085
*
.include "sky130_fd_sc_hs__nand2b_2.pxi.spice"
*
.ends
*
*
