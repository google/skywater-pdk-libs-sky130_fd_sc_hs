* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hs__o22ai_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
X0 a_27_74# A1 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X1 a_27_74# A2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X2 VGND A1 a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X3 Y B1 a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X4 a_117_368# A1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X5 a_27_74# B2 Y VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X6 a_877_368# B1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X7 a_117_368# A2 Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X8 Y B2 a_877_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X9 Y B2 a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X10 Y B2 a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X11 a_27_74# B1 Y VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X12 Y A2 a_117_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X13 a_117_368# A1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X14 a_877_368# B1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X15 Y A2 a_117_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X16 VGND A2 a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X17 Y B2 a_877_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X18 VPWR B1 a_877_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X19 a_27_74# B2 Y VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X20 VPWR A1 a_117_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X21 a_27_74# A2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X22 a_877_368# B2 Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X23 VGND A1 a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X24 VGND A2 a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X25 VPWR A1 a_117_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X26 a_877_368# B2 Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X27 Y B1 a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X28 VPWR B1 a_877_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X29 a_117_368# A2 Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X30 a_27_74# A1 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X31 a_27_74# B1 Y VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
.ends
