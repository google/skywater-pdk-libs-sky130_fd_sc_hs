* File: sky130_fd_sc_hs__nand3b_2.pex.spice
* Created: Tue Sep  1 20:09:37 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HS__NAND3B_2%A_N 3 5 7 8 12 13
c33 5 0 1.52485e-19 $X=0.695 $Y=1.885
c34 3 0 1.99845e-19 $X=0.48 $Y=0.79
r35 13 14 35.7345 $w=2.9e-07 $l=2.15e-07 $layer=POLY_cond $X=0.48 $Y=1.667
+ $X2=0.695 $Y2=1.667
r36 11 13 15.7897 $w=2.9e-07 $l=9.5e-08 $layer=POLY_cond $X=0.385 $Y=1.667
+ $X2=0.48 $Y2=1.667
r37 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.385
+ $Y=1.615 $X2=0.385 $Y2=1.615
r38 8 12 5.06376 $w=3.28e-07 $l=1.45e-07 $layer=LI1_cond $X=0.24 $Y=1.615
+ $X2=0.385 $Y2=1.615
r39 5 14 18.1727 $w=1.5e-07 $l=2.18e-07 $layer=POLY_cond $X=0.695 $Y=1.885
+ $X2=0.695 $Y2=1.667
r40 5 7 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=0.695 $Y=1.885
+ $X2=0.695 $Y2=2.46
r41 1 13 18.1727 $w=1.5e-07 $l=2.17e-07 $layer=POLY_cond $X=0.48 $Y=1.45
+ $X2=0.48 $Y2=1.667
r42 1 3 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.48 $Y=1.45 $X2=0.48
+ $Y2=0.79
.ends

.subckt PM_SKY130_FD_SC_HS__NAND3B_2%C 1 3 4 6 7 9 10 12 13 14 21
c61 21 0 1.66669e-20 $X=1.615 $Y=1.515
r62 21 23 8.74376 $w=4.41e-07 $l=8e-08 $layer=POLY_cond $X=1.615 $Y=1.475
+ $X2=1.695 $Y2=1.475
r63 21 22 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.615
+ $Y=1.515 $X2=1.615 $Y2=1.515
r64 19 21 25.1383 $w=4.41e-07 $l=2.3e-07 $layer=POLY_cond $X=1.385 $Y=1.475
+ $X2=1.615 $Y2=1.475
r65 18 19 20.22 $w=4.41e-07 $l=1.85e-07 $layer=POLY_cond $X=1.2 $Y=1.475
+ $X2=1.385 $Y2=1.475
r66 14 22 2.14025 $w=3.48e-07 $l=6.5e-08 $layer=LI1_cond $X=1.68 $Y=1.605
+ $X2=1.615 $Y2=1.605
r67 13 22 13.6647 $w=3.48e-07 $l=4.15e-07 $layer=LI1_cond $X=1.2 $Y=1.605
+ $X2=1.615 $Y2=1.605
r68 10 23 28.2648 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=1.695 $Y=1.765
+ $X2=1.695 $Y2=1.475
r69 10 12 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.695 $Y=1.765
+ $X2=1.695 $Y2=2.4
r70 7 19 28.2648 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=1.385 $Y=1.185
+ $X2=1.385 $Y2=1.475
r71 7 9 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=1.385 $Y=1.185
+ $X2=1.385 $Y2=0.74
r72 4 18 28.2648 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=1.2 $Y=1.765 $X2=1.2
+ $Y2=1.475
r73 4 6 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.2 $Y=1.765 $X2=1.2
+ $Y2=2.4
r74 1 18 26.7778 $w=4.41e-07 $l=3.93891e-07 $layer=POLY_cond $X=0.955 $Y=1.185
+ $X2=1.2 $Y2=1.475
r75 1 3 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=0.955 $Y=1.185
+ $X2=0.955 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HS__NAND3B_2%A_27_94# 1 2 7 9 10 12 13 15 18 22 26 28 29
+ 31 32 37 39 40 47
c112 37 0 1.66669e-20 $X=0.805 $Y=2.035
c113 13 0 5.47792e-20 $X=2.645 $Y=1.765
r114 46 47 31.8971 $w=3.4e-07 $l=2.25e-07 $layer=POLY_cond $X=2.42 $Y=1.557
+ $X2=2.645 $Y2=1.557
r115 45 46 31.8971 $w=3.4e-07 $l=2.25e-07 $layer=POLY_cond $X=2.195 $Y=1.557
+ $X2=2.42 $Y2=1.557
r116 43 45 0.708824 $w=3.4e-07 $l=5e-09 $layer=POLY_cond $X=2.19 $Y=1.557
+ $X2=2.195 $Y2=1.557
r117 42 43 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.19
+ $Y=1.515 $X2=2.19 $Y2=1.515
r118 40 42 16.0154 $w=2.59e-07 $l=3.4e-07 $layer=LI1_cond $X=2.19 $Y=1.175
+ $X2=2.19 $Y2=1.515
r119 35 37 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=0.47 $Y=2.035
+ $X2=0.805 $Y2=2.035
r120 33 39 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.89 $Y=1.175
+ $X2=0.805 $Y2=1.175
r121 32 40 3.20129 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.025 $Y=1.175
+ $X2=2.19 $Y2=1.175
r122 32 33 74.0481 $w=1.68e-07 $l=1.135e-06 $layer=LI1_cond $X=2.025 $Y=1.175
+ $X2=0.89 $Y2=1.175
r123 31 37 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.805 $Y=1.95
+ $X2=0.805 $Y2=2.035
r124 30 39 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.805 $Y=1.26
+ $X2=0.805 $Y2=1.175
r125 30 31 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=0.805 $Y=1.26
+ $X2=0.805 $Y2=1.95
r126 28 39 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.72 $Y=1.175
+ $X2=0.805 $Y2=1.175
r127 28 29 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.72 $Y=1.175
+ $X2=0.35 $Y2=1.175
r128 26 35 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=0.47 $Y=2.815
+ $X2=0.47 $Y2=2.12
r129 20 29 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.225 $Y=1.09
+ $X2=0.35 $Y2=1.175
r130 20 22 21.8964 $w=2.48e-07 $l=4.75e-07 $layer=LI1_cond $X=0.225 $Y=1.09
+ $X2=0.225 $Y2=0.615
r131 16 47 29.0618 $w=3.4e-07 $l=2.05e-07 $layer=POLY_cond $X=2.85 $Y=1.557
+ $X2=2.645 $Y2=1.557
r132 16 18 271.766 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=2.85 $Y=1.4
+ $X2=2.85 $Y2=0.87
r133 13 47 21.9347 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=2.645 $Y=1.765
+ $X2=2.645 $Y2=1.557
r134 13 15 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.645 $Y=1.765
+ $X2=2.645 $Y2=2.4
r135 10 46 21.9347 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.42 $Y=1.35
+ $X2=2.42 $Y2=1.557
r136 10 12 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=2.42 $Y=1.35
+ $X2=2.42 $Y2=0.87
r137 7 45 21.9347 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=2.195 $Y=1.765
+ $X2=2.195 $Y2=1.557
r138 7 9 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.195 $Y=1.765
+ $X2=2.195 $Y2=2.4
r139 2 35 400 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_PDIFF $count=1 $X=0.325
+ $Y=1.96 $X2=0.47 $Y2=2.115
r140 2 26 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=0.325
+ $Y=1.96 $X2=0.47 $Y2=2.815
r141 1 22 91 $w=1.7e-07 $l=1.99687e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.47 $X2=0.265 $Y2=0.615
.ends

.subckt PM_SKY130_FD_SC_HS__NAND3B_2%B 1 3 4 6 7 9 10 12 13 14 15 24
c43 15 0 5.47792e-20 $X=4.08 $Y=1.665
r44 24 25 3.30137 $w=3.65e-07 $l=2.5e-08 $layer=POLY_cond $X=3.815 $Y=1.557
+ $X2=3.84 $Y2=1.557
r45 22 24 8.58356 $w=3.65e-07 $l=6.5e-08 $layer=POLY_cond $X=3.75 $Y=1.557
+ $X2=3.815 $Y2=1.557
r46 22 23 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.75
+ $Y=1.515 $X2=3.75 $Y2=1.515
r47 20 22 44.8986 $w=3.65e-07 $l=3.4e-07 $layer=POLY_cond $X=3.41 $Y=1.557
+ $X2=3.75 $Y2=1.557
r48 19 20 13.8658 $w=3.65e-07 $l=1.05e-07 $layer=POLY_cond $X=3.305 $Y=1.557
+ $X2=3.41 $Y2=1.557
r49 15 23 8.84433 $w=4.28e-07 $l=3.3e-07 $layer=LI1_cond $X=4.08 $Y=1.565
+ $X2=3.75 $Y2=1.565
r50 14 23 4.02015 $w=4.28e-07 $l=1.5e-07 $layer=LI1_cond $X=3.6 $Y=1.565
+ $X2=3.75 $Y2=1.565
r51 13 14 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=3.12 $Y=1.565
+ $X2=3.6 $Y2=1.565
r52 10 25 23.6381 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.84 $Y=1.35
+ $X2=3.84 $Y2=1.557
r53 10 12 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=3.84 $Y=1.35 $X2=3.84
+ $Y2=0.87
r54 7 24 23.6381 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=3.815 $Y=1.765
+ $X2=3.815 $Y2=1.557
r55 7 9 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.815 $Y=1.765
+ $X2=3.815 $Y2=2.4
r56 4 20 23.6381 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.41 $Y=1.35
+ $X2=3.41 $Y2=1.557
r57 4 6 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=3.41 $Y=1.35 $X2=3.41
+ $Y2=0.87
r58 1 19 23.6381 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=3.305 $Y=1.765
+ $X2=3.305 $Y2=1.557
r59 1 3 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.305 $Y=1.765
+ $X2=3.305 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_HS__NAND3B_2%VPWR 1 2 3 4 15 19 23 25 27 32 33 35 36 38
+ 39 40 52 58
r62 57 58 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r63 55 58 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.08 $Y2=3.33
r64 54 55 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r65 52 57 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=3.875 $Y=3.33
+ $X2=4.097 $Y2=3.33
r66 52 54 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=3.875 $Y=3.33
+ $X2=3.6 $Y2=3.33
r67 51 55 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.6 $Y2=3.33
r68 50 51 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r69 47 48 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r70 44 48 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.68 $Y2=3.33
r71 43 44 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r72 40 51 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r73 40 48 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.68 $Y2=3.33
r74 38 50 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=2.79 $Y=3.33 $X2=2.64
+ $Y2=3.33
r75 38 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.79 $Y=3.33
+ $X2=2.955 $Y2=3.33
r76 37 54 31.3155 $w=1.68e-07 $l=4.8e-07 $layer=LI1_cond $X=3.12 $Y=3.33 $X2=3.6
+ $Y2=3.33
r77 37 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.12 $Y=3.33
+ $X2=2.955 $Y2=3.33
r78 35 47 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=1.805 $Y=3.33
+ $X2=1.68 $Y2=3.33
r79 35 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.805 $Y=3.33
+ $X2=1.97 $Y2=3.33
r80 34 50 32.9465 $w=1.68e-07 $l=5.05e-07 $layer=LI1_cond $X=2.135 $Y=3.33
+ $X2=2.64 $Y2=3.33
r81 34 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.135 $Y=3.33
+ $X2=1.97 $Y2=3.33
r82 32 43 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=0.83 $Y=3.33
+ $X2=0.72 $Y2=3.33
r83 32 33 6.92067 $w=1.7e-07 $l=1.22e-07 $layer=LI1_cond $X=0.83 $Y=3.33
+ $X2=0.952 $Y2=3.33
r84 31 47 39.4706 $w=1.68e-07 $l=6.05e-07 $layer=LI1_cond $X=1.075 $Y=3.33
+ $X2=1.68 $Y2=3.33
r85 31 33 6.92067 $w=1.7e-07 $l=1.23e-07 $layer=LI1_cond $X=1.075 $Y=3.33
+ $X2=0.952 $Y2=3.33
r86 27 30 27.2396 $w=3.28e-07 $l=7.8e-07 $layer=LI1_cond $X=4.04 $Y=2.035
+ $X2=4.04 $Y2=2.815
r87 25 57 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=4.04 $Y=3.245
+ $X2=4.097 $Y2=3.33
r88 25 30 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=4.04 $Y=3.245
+ $X2=4.04 $Y2=2.815
r89 21 39 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.955 $Y=3.245
+ $X2=2.955 $Y2=3.33
r90 21 23 29.1603 $w=3.28e-07 $l=8.35e-07 $layer=LI1_cond $X=2.955 $Y=3.245
+ $X2=2.955 $Y2=2.41
r91 17 36 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.97 $Y=3.245
+ $X2=1.97 $Y2=3.33
r92 17 19 29.1603 $w=3.28e-07 $l=8.35e-07 $layer=LI1_cond $X=1.97 $Y=3.245
+ $X2=1.97 $Y2=2.41
r93 13 33 0.066131 $w=2.45e-07 $l=8.5e-08 $layer=LI1_cond $X=0.952 $Y=3.245
+ $X2=0.952 $Y2=3.33
r94 13 15 37.1604 $w=2.43e-07 $l=7.9e-07 $layer=LI1_cond $X=0.952 $Y=3.245
+ $X2=0.952 $Y2=2.455
r95 4 30 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=3.89
+ $Y=1.84 $X2=4.04 $Y2=2.815
r96 4 27 400 $w=1.7e-07 $l=2.59374e-07 $layer=licon1_PDIFF $count=1 $X=3.89
+ $Y=1.84 $X2=4.04 $Y2=2.035
r97 3 23 300 $w=1.7e-07 $l=6.77385e-07 $layer=licon1_PDIFF $count=2 $X=2.72
+ $Y=1.84 $X2=2.955 $Y2=2.41
r98 2 19 300 $w=1.7e-07 $l=6.62495e-07 $layer=licon1_PDIFF $count=2 $X=1.77
+ $Y=1.84 $X2=1.97 $Y2=2.41
r99 1 15 300 $w=1.7e-07 $l=5.78035e-07 $layer=licon1_PDIFF $count=2 $X=0.77
+ $Y=1.96 $X2=0.95 $Y2=2.455
.ends

.subckt PM_SKY130_FD_SC_HS__NAND3B_2%Y 1 2 3 4 13 15 17 21 23 24 25 27 37 42
c67 13 0 1.52485e-19 $X=1.447 $Y=2.12
r68 39 42 20.3249 $w=2.73e-07 $l=4.85e-07 $layer=LI1_cond $X=2.662 $Y=1.18
+ $X2=2.662 $Y2=1.665
r69 37 39 3.32251 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=2.635 $Y=1.095
+ $X2=2.635 $Y2=1.18
r70 34 42 11.9435 $w=2.73e-07 $l=2.85e-07 $layer=LI1_cond $X=2.662 $Y=1.95
+ $X2=2.662 $Y2=1.665
r71 32 34 15.7882 $w=1.68e-07 $l=2.42e-07 $layer=LI1_cond $X=2.42 $Y=2.035
+ $X2=2.662 $Y2=2.035
r72 25 41 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.53 $Y=2.12 $X2=3.53
+ $Y2=2.035
r73 25 27 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=3.53 $Y=2.12
+ $X2=3.53 $Y2=2.815
r74 24 34 9.00321 $w=1.68e-07 $l=1.38e-07 $layer=LI1_cond $X=2.8 $Y=2.035
+ $X2=2.662 $Y2=2.035
r75 23 41 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.365 $Y=2.035
+ $X2=3.53 $Y2=2.035
r76 23 24 36.861 $w=1.68e-07 $l=5.65e-07 $layer=LI1_cond $X=3.365 $Y=2.035
+ $X2=2.8 $Y2=2.035
r77 21 32 14.2903 $w=2.48e-07 $l=3.1e-07 $layer=LI1_cond $X=2.46 $Y=2.43
+ $X2=2.46 $Y2=2.12
r78 18 30 5.61466 $w=1.7e-07 $l=1.88e-07 $layer=LI1_cond $X=1.635 $Y=2.035
+ $X2=1.447 $Y2=2.035
r79 17 32 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=2.335 $Y=2.035
+ $X2=2.42 $Y2=2.035
r80 17 18 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=2.335 $Y=2.035
+ $X2=1.635 $Y2=2.035
r81 13 30 2.53854 $w=3.75e-07 $l=8.5e-08 $layer=LI1_cond $X=1.447 $Y=2.12
+ $X2=1.447 $Y2=2.035
r82 13 15 21.3586 $w=3.73e-07 $l=6.95e-07 $layer=LI1_cond $X=1.447 $Y=2.12
+ $X2=1.447 $Y2=2.815
r83 4 41 400 $w=1.7e-07 $l=2.59374e-07 $layer=licon1_PDIFF $count=1 $X=3.38
+ $Y=1.84 $X2=3.53 $Y2=2.035
r84 4 27 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=3.38
+ $Y=1.84 $X2=3.53 $Y2=2.815
r85 3 32 600 $w=1.7e-07 $l=2.59374e-07 $layer=licon1_PDIFF $count=1 $X=2.27
+ $Y=1.84 $X2=2.42 $Y2=2.035
r86 3 21 300 $w=1.7e-07 $l=6.60757e-07 $layer=licon1_PDIFF $count=2 $X=2.27
+ $Y=1.84 $X2=2.42 $Y2=2.43
r87 2 30 400 $w=1.7e-07 $l=2.66786e-07 $layer=licon1_PDIFF $count=1 $X=1.275
+ $Y=1.84 $X2=1.445 $Y2=2.035
r88 2 15 400 $w=1.7e-07 $l=1.05659e-06 $layer=licon1_PDIFF $count=1 $X=1.275
+ $Y=1.84 $X2=1.445 $Y2=2.815
r89 1 37 182 $w=1.7e-07 $l=6.61306e-07 $layer=licon1_NDIFF $count=1 $X=2.495
+ $Y=0.5 $X2=2.635 $Y2=1.095
.ends

.subckt PM_SKY130_FD_SC_HS__NAND3B_2%VGND 1 2 9 13 15 17 22 32 33 36 39
r46 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r47 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r48 32 33 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r49 29 32 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=2.16 $Y=0 $X2=4.08
+ $Y2=0
r50 27 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.765 $Y=0 $X2=1.6
+ $Y2=0
r51 27 29 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=1.765 $Y=0 $X2=2.16
+ $Y2=0
r52 26 40 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=1.68
+ $Y2=0
r53 26 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r54 25 26 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r55 23 36 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=0.82 $Y=0 $X2=0.675
+ $Y2=0
r56 23 25 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=0.82 $Y=0 $X2=1.2
+ $Y2=0
r57 22 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.435 $Y=0 $X2=1.6
+ $Y2=0
r58 22 25 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=1.435 $Y=0 $X2=1.2
+ $Y2=0
r59 20 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r60 19 20 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r61 17 36 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=0.53 $Y=0 $X2=0.675
+ $Y2=0
r62 17 19 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=0.53 $Y=0 $X2=0.24
+ $Y2=0
r63 15 33 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=2.16 $Y=0 $X2=4.08
+ $Y2=0
r64 15 40 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.68
+ $Y2=0
r65 15 29 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r66 11 39 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.6 $Y=0.085 $X2=1.6
+ $Y2=0
r67 11 13 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=1.6 $Y=0.085 $X2=1.6
+ $Y2=0.495
r68 7 36 0.489042 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=0.675 $Y=0.085
+ $X2=0.675 $Y2=0
r69 7 9 25.4332 $w=2.88e-07 $l=6.4e-07 $layer=LI1_cond $X=0.675 $Y=0.085
+ $X2=0.675 $Y2=0.725
r70 2 13 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=1.46
+ $Y=0.37 $X2=1.6 $Y2=0.495
r71 1 9 182 $w=1.7e-07 $l=3.17372e-07 $layer=licon1_NDIFF $count=1 $X=0.555
+ $Y=0.47 $X2=0.695 $Y2=0.725
.ends

.subckt PM_SKY130_FD_SC_HS__NAND3B_2%A_206_74# 1 2 7 9 17 18 20 21
c42 9 0 1.99845e-19 $X=1.17 $Y=0.495
r43 20 21 21.0706 $w=5.08e-07 $l=6.55e-07 $layer=LI1_cond $X=3.625 $Y=0.925
+ $X2=2.97 $Y2=0.925
r44 18 21 56.4332 $w=1.68e-07 $l=8.65e-07 $layer=LI1_cond $X=2.105 $Y=0.755
+ $X2=2.97 $Y2=0.755
r45 17 18 7.83661 $w=2.48e-07 $l=1.7e-07 $layer=LI1_cond $X=1.935 $Y=0.795
+ $X2=2.105 $Y2=0.795
r46 12 16 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.255 $Y=0.835
+ $X2=1.13 $Y2=0.835
r47 12 17 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.255 $Y=0.835
+ $X2=1.935 $Y2=0.835
r48 7 16 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.13 $Y=0.75 $X2=1.13
+ $Y2=0.835
r49 7 9 11.7549 $w=2.48e-07 $l=2.55e-07 $layer=LI1_cond $X=1.13 $Y=0.75 $X2=1.13
+ $Y2=0.495
r50 2 20 91 $w=1.7e-07 $l=3.17372e-07 $layer=licon1_NDIFF $count=2 $X=3.485
+ $Y=0.5 $X2=3.625 $Y2=0.755
r51 1 16 182 $w=1.7e-07 $l=5.30401e-07 $layer=licon1_NDIFF $count=1 $X=1.03
+ $Y=0.37 $X2=1.17 $Y2=0.835
r52 1 9 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=1.03
+ $Y=0.37 $X2=1.17 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_HS__NAND3B_2%A_403_54# 1 2 3 10 18
r16 16 18 6.42709 $w=2.58e-07 $l=1.45e-07 $layer=LI1_cond $X=4.09 $Y=0.5
+ $X2=4.09 $Y2=0.645
r17 12 15 64.5882 $w=1.68e-07 $l=9.9e-07 $layer=LI1_cond $X=2.14 $Y=0.415
+ $X2=3.13 $Y2=0.415
r18 10 16 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=3.96 $Y=0.415
+ $X2=4.09 $Y2=0.5
r19 10 15 54.1497 $w=1.68e-07 $l=8.3e-07 $layer=LI1_cond $X=3.96 $Y=0.415
+ $X2=3.13 $Y2=0.415
r20 3 18 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.915
+ $Y=0.5 $X2=4.055 $Y2=0.645
r21 2 15 182 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NDIFF $count=1 $X=2.925
+ $Y=0.5 $X2=3.13 $Y2=0.415
r22 1 12 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=2.015
+ $Y=0.27 $X2=2.14 $Y2=0.415
.ends

