* File: sky130_fd_sc_hs__dfbbn_1.spice
* Created: Thu Aug 27 20:37:49 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hs__dfbbn_1.pex.spice"
.subckt sky130_fd_sc_hs__dfbbn_1  VNB VPB CLK_N D SET_B RESET_B VPWR Q_N Q VGND
* 
* VGND	VGND
* Q	Q
* Q_N	Q_N
* VPWR	VPWR
* RESET_B	RESET_B
* SET_B	SET_B
* D	D
* CLK_N	CLK_N
* VPB	VPB
* VNB	VNB
MM1035 N_VGND_M1035_d N_CLK_N_M1035_g N_A_27_74#_M1035_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.2109 PD=1.02 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75000.6 A=0.111 P=1.78 MULT=1
MM1036 N_A_200_74#_M1036_d N_A_27_74#_M1036_g N_VGND_M1035_d VNB NLOWVT L=0.15
+ W=0.74 AD=0.2109 AS=0.1036 PD=2.05 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.6 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1015 N_VGND_M1015_d N_D_M1015_g N_A_311_119#_M1015_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.137937 AS=0.1197 PD=1.13 PS=1.41 NRD=78.12 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75002 A=0.063 P=1.14 MULT=1
MM1013 A_523_119# N_A_474_405#_M1013_g N_VGND_M1015_d VNB NLOWVT L=0.15 W=0.42
+ AD=0.0441 AS=0.137937 PD=0.63 PS=1.13 NRD=14.28 NRS=78.12 M=1 R=2.8 SA=75000.8
+ SB=75001.4 A=0.063 P=1.14 MULT=1
MM1004 N_A_595_119#_M1004_d N_A_27_74#_M1004_g A_523_119# VNB NLOWVT L=0.15
+ W=0.42 AD=0.0588 AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75001.2
+ SB=75001 A=0.063 P=1.14 MULT=1
MM1007 N_A_311_119#_M1007_d N_A_200_74#_M1007_g N_A_595_119#_M1004_d VNB NLOWVT
+ L=0.15 W=0.42 AD=0.40005 AS=0.0588 PD=2.58 PS=0.7 NRD=256.428 NRS=0 M=1 R=2.8
+ SA=75001.6 SB=75000.6 A=0.063 P=1.14 MULT=1
MM1020 N_A_474_405#_M1020_d N_A_595_119#_M1020_g N_A_867_119#_M1020_s VNB NLOWVT
+ L=0.15 W=0.55 AD=0.09625 AS=0.15675 PD=0.9 PS=1.67 NRD=15.264 NRS=0 M=1
+ R=3.66667 SA=75000.2 SB=75004.8 A=0.0825 P=1.4 MULT=1
MM1030 N_A_867_119#_M1030_d N_A_978_357#_M1030_g N_A_474_405#_M1020_d VNB NLOWVT
+ L=0.15 W=0.55 AD=0.09625 AS=0.09625 PD=0.9 PS=0.9 NRD=15.264 NRS=0 M=1
+ R=3.66667 SA=75000.7 SB=75004.3 A=0.0825 P=1.4 MULT=1
MM1026 N_VGND_M1026_d N_SET_B_M1026_g N_A_867_119#_M1030_d VNB NLOWVT L=0.15
+ W=0.55 AD=0.09625 AS=0.09625 PD=0.9 PS=0.9 NRD=15.264 NRS=0 M=1 R=3.66667
+ SA=75001.2 SB=75003.8 A=0.0825 P=1.4 MULT=1
MM1025 A_1254_119# N_A_474_405#_M1025_g N_VGND_M1026_d VNB NLOWVT L=0.15 W=0.55
+ AD=0.0915625 AS=0.09625 PD=0.9 PS=0.9 NRD=24.312 NRS=0 M=1 R=3.66667
+ SA=75001.7 SB=75003.3 A=0.0825 P=1.4 MULT=1
MM1027 N_A_1349_114#_M1027_d N_A_27_74#_M1027_g A_1254_119# VNB NLOWVT L=0.15
+ W=0.55 AD=0.356224 AS=0.0915625 PD=1.93918 PS=0.9 NRD=0 NRS=24.312 M=1
+ R=3.66667 SA=75002.1 SB=75002.9 A=0.0825 P=1.4 MULT=1
MM1024 A_1611_140# N_A_200_74#_M1024_g N_A_1349_114#_M1027_d VNB NLOWVT L=0.15
+ W=0.42 AD=0.0504 AS=0.272026 PD=0.66 PS=1.48082 NRD=18.564 NRS=22.848 M=1
+ R=2.8 SA=75003.5 SB=75002.2 A=0.063 P=1.14 MULT=1
MM1001 N_VGND_M1001_d N_A_1534_446#_M1001_g A_1611_140# VNB NLOWVT L=0.15 W=0.42
+ AD=0.108295 AS=0.0504 PD=0.89431 PS=0.66 NRD=57.948 NRS=18.564 M=1 R=2.8
+ SA=75003.9 SB=75001.8 A=0.063 P=1.14 MULT=1
MM1017 N_A_1818_76#_M1017_d N_SET_B_M1017_g N_VGND_M1001_d VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.190805 PD=1.02 PS=1.57569 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75002.7 SB=75001.2 A=0.111 P=1.78 MULT=1
MM1034 N_A_1534_446#_M1034_d N_A_978_357#_M1034_g N_A_1818_76#_M1017_d VNB
+ NLOWVT L=0.15 W=0.74 AD=0.1184 AS=0.1036 PD=1.06 PS=1.02 NRD=3.24 NRS=0 M=1
+ R=4.93333 SA=75003.1 SB=75000.7 A=0.111 P=1.78 MULT=1
MM1033 N_A_1818_76#_M1033_d N_A_1349_114#_M1033_g N_A_1534_446#_M1034_d VNB
+ NLOWVT L=0.15 W=0.74 AD=0.296 AS=0.1184 PD=2.52 PS=1.06 NRD=55.944 NRS=0 M=1
+ R=4.93333 SA=75003.6 SB=75000.3 A=0.111 P=1.78 MULT=1
MM1011 N_VGND_M1011_d N_RESET_B_M1011_g N_A_978_357#_M1011_s VNB NLOWVT L=0.15
+ W=0.42 AD=0.12457 AS=0.1134 PD=1.00293 PS=1.38 NRD=69.024 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75000.8 A=0.063 P=1.14 MULT=1
MM1028 N_Q_N_M1028_d N_A_1534_446#_M1028_g N_VGND_M1011_d VNB NLOWVT L=0.15
+ W=0.74 AD=0.1998 AS=0.21948 PD=2.02 PS=1.76707 NRD=0 NRS=39.168 M=1 R=4.93333
+ SA=75000.5 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1005 N_VGND_M1005_d N_A_1534_446#_M1005_g N_A_2412_410#_M1005_s VNB NLOWVT
+ L=0.15 W=0.42 AD=0.0837466 AS=0.1134 PD=0.78569 PS=1.38 NRD=18.564 NRS=0 M=1
+ R=2.8 SA=75000.2 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1012 N_Q_M1012_d N_A_2412_410#_M1012_g N_VGND_M1005_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.1998 AS=0.147553 PD=2.02 PS=1.38431 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.5
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1002 N_VPWR_M1002_d N_CLK_N_M1002_g N_A_27_74#_M1002_s VPB PSHORT L=0.15
+ W=1.12 AD=0.168 AS=0.3192 PD=1.42 PS=2.81 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1003 N_A_200_74#_M1003_d N_A_27_74#_M1003_g N_VPWR_M1002_d VPB PSHORT L=0.15
+ W=1.12 AD=0.3136 AS=0.168 PD=2.8 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.7 SB=75000.2 A=0.168 P=2.54 MULT=1
MM1029 N_VPWR_M1029_d N_D_M1029_g N_A_311_119#_M1029_s VPB PSHORT L=0.15 W=0.42
+ AD=0.0945 AS=0.17805 PD=0.87 PS=1.75 NRD=72.693 NRS=46.886 M=1 R=2.8
+ SA=75000.3 SB=75001.8 A=0.063 P=1.14 MULT=1
MM1016 A_537_503# N_A_474_405#_M1016_g N_VPWR_M1029_d VPB PSHORT L=0.15 W=0.42
+ AD=0.0567 AS=0.0945 PD=0.69 PS=0.87 NRD=37.5088 NRS=7.0329 M=1 R=2.8
+ SA=75000.9 SB=75001.2 A=0.063 P=1.14 MULT=1
MM1006 N_A_595_119#_M1006_d N_A_200_74#_M1006_g A_537_503# VPB PSHORT L=0.15
+ W=0.42 AD=0.0756 AS=0.0567 PD=0.78 PS=0.69 NRD=18.7544 NRS=37.5088 M=1 R=2.8
+ SA=75001.3 SB=75000.8 A=0.063 P=1.14 MULT=1
MM1019 N_A_311_119#_M1019_d N_A_27_74#_M1019_g N_A_595_119#_M1006_d VPB PSHORT
+ L=0.15 W=0.42 AD=0.1704 AS=0.0756 PD=1.72 PS=0.78 NRD=39.8531 NRS=18.7544 M=1
+ R=2.8 SA=75001.8 SB=75000.3 A=0.063 P=1.14 MULT=1
MM1037 A_933_424# N_A_595_119#_M1037_g N_A_474_405#_M1037_s VPB PSHORT L=0.15
+ W=0.84 AD=0.1008 AS=0.2352 PD=1.08 PS=2.24 NRD=15.2281 NRS=2.3443 M=1 R=5.6
+ SA=75000.2 SB=75001 A=0.126 P=1.98 MULT=1
MM1022 N_VPWR_M1022_d N_A_978_357#_M1022_g A_933_424# VPB PSHORT L=0.15 W=0.84
+ AD=0.126 AS=0.1008 PD=1.14 PS=1.08 NRD=2.3443 NRS=15.2281 M=1 R=5.6 SA=75000.6
+ SB=75000.7 A=0.126 P=1.98 MULT=1
MM1038 N_A_474_405#_M1038_d N_SET_B_M1038_g N_VPWR_M1022_d VPB PSHORT L=0.15
+ W=0.84 AD=0.2352 AS=0.126 PD=2.24 PS=1.14 NRD=2.3443 NRS=2.3443 M=1 R=5.6
+ SA=75001 SB=75000.2 A=0.126 P=1.98 MULT=1
MM1018 A_1297_424# N_A_474_405#_M1018_g N_VPWR_M1018_s VPB PSHORT L=0.15 W=0.84
+ AD=0.1008 AS=0.2352 PD=1.08 PS=2.24 NRD=15.2281 NRS=2.3443 M=1 R=5.6
+ SA=75000.2 SB=75001.1 A=0.126 P=1.98 MULT=1
MM1009 N_A_1349_114#_M1009_d N_A_200_74#_M1009_g A_1297_424# VPB PSHORT L=0.15
+ W=0.84 AD=0.1918 AS=0.1008 PD=1.64 PS=1.08 NRD=2.3443 NRS=15.2281 M=1 R=5.6
+ SA=75000.6 SB=75000.8 A=0.126 P=1.98 MULT=1
MM1031 A_1483_508# N_A_27_74#_M1031_g N_A_1349_114#_M1009_d VPB PSHORT L=0.15
+ W=0.42 AD=0.0567 AS=0.0959 PD=0.69 PS=0.82 NRD=37.5088 NRS=46.886 M=1 R=2.8
+ SA=75001.1 SB=75000.8 A=0.063 P=1.14 MULT=1
MM1000 N_VPWR_M1000_d N_A_1534_446#_M1000_g A_1483_508# VPB PSHORT L=0.15 W=0.42
+ AD=0.250675 AS=0.0567 PD=2.14 PS=0.69 NRD=254.15 NRS=37.5088 M=1 R=2.8
+ SA=75001.6 SB=75000.3 A=0.063 P=1.14 MULT=1
MM1039 N_VPWR_M1039_d N_SET_B_M1039_g N_A_1534_446#_M1039_s VPB PSHORT L=0.15
+ W=1 AD=0.269075 AS=0.295 PD=1.705 PS=2.59 NRD=42.158 NRS=1.9503 M=1 R=6.66667
+ SA=75000.2 SB=75001.2 A=0.15 P=2.3 MULT=1
MM1032 A_1917_392# N_A_978_357#_M1032_g N_VPWR_M1039_d VPB PSHORT L=0.15 W=1
+ AD=0.135 AS=0.269075 PD=1.27 PS=1.705 NRD=15.7403 NRS=42.158 M=1 R=6.66667
+ SA=75000.8 SB=75000.6 A=0.15 P=2.3 MULT=1
MM1014 N_A_1534_446#_M1014_d N_A_1349_114#_M1014_g A_1917_392# VPB PSHORT L=0.15
+ W=1 AD=0.28 AS=0.135 PD=2.56 PS=1.27 NRD=1.9503 NRS=15.7403 M=1 R=6.66667
+ SA=75001.3 SB=75000.2 A=0.15 P=2.3 MULT=1
MM1021 N_VPWR_M1021_d N_RESET_B_M1021_g N_A_978_357#_M1021_s VPB PSHORT L=0.15
+ W=0.64 AD=0.137018 AS=0.1792 PD=1.08727 PS=1.84 NRD=48.9545 NRS=3.0732 M=1
+ R=4.26667 SA=75000.2 SB=75000.7 A=0.096 P=1.58 MULT=1
MM1023 N_Q_N_M1023_d N_A_1534_446#_M1023_g N_VPWR_M1021_d VPB PSHORT L=0.15
+ W=1.12 AD=0.3136 AS=0.239782 PD=2.8 PS=1.90273 NRD=1.7533 NRS=1.7533 M=1
+ R=7.46667 SA=75000.5 SB=75000.2 A=0.168 P=2.54 MULT=1
MM1010 N_VPWR_M1010_d N_A_1534_446#_M1010_g N_A_2412_410#_M1010_s VPB PSHORT
+ L=0.15 W=0.84 AD=0.1692 AS=0.2394 PD=1.28143 PS=2.25 NRD=37.5088 NRS=0 M=1
+ R=5.6 SA=75000.2 SB=75000.7 A=0.126 P=1.98 MULT=1
MM1008 N_Q_M1008_d N_A_2412_410#_M1008_g N_VPWR_M1010_d VPB PSHORT L=0.15 W=1.12
+ AD=0.3192 AS=0.2256 PD=2.81 PS=1.70857 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.6 SB=75000.2 A=0.168 P=2.54 MULT=1
DX40_noxref VNB VPB NWDIODE A=25.7052 P=31.36
c_142 VNB 0 5.76555e-20 $X=0 $Y=0
c_274 VPB 0 4.72451e-19 $X=0 $Y=3.085
*
.include "sky130_fd_sc_hs__dfbbn_1.pxi.spice"
*
.ends
*
*
