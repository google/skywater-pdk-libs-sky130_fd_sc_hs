# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_hs__and4b_4
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_hs__and4b_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  7.680000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A_N
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425000 1.190000 0.835000 1.550000 ;
    END
  END A_N
  PIN B
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.845000 1.470000 7.180000 1.800000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.915000 1.350000 3.245000 1.780000 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.965000 1.470000 5.155000 1.800000 ;
    END
  END D
  PIN X
    ANTENNADIFFAREA  1.209600 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.085000 0.350000 1.470000 0.980000 ;
        RECT 1.085000 0.980000 2.540000 1.150000 ;
        RECT 1.085000 1.150000 1.315000 1.820000 ;
        RECT 1.085000 1.820000 2.405000 2.220000 ;
        RECT 2.210000 0.350000 2.540000 0.980000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 7.680000 0.085000 ;
        RECT 0.585000  0.085000 0.915000 1.020000 ;
        RECT 1.670000  0.085000 2.000000 0.810000 ;
        RECT 2.710000  0.085000 3.040000 1.130000 ;
        RECT 4.285000  0.085000 4.615000 0.620000 ;
      LAYER mcon ;
        RECT 0.155000 -0.085000 0.325000 0.085000 ;
        RECT 0.635000 -0.085000 0.805000 0.085000 ;
        RECT 1.115000 -0.085000 1.285000 0.085000 ;
        RECT 1.595000 -0.085000 1.765000 0.085000 ;
        RECT 2.075000 -0.085000 2.245000 0.085000 ;
        RECT 2.555000 -0.085000 2.725000 0.085000 ;
        RECT 3.035000 -0.085000 3.205000 0.085000 ;
        RECT 3.515000 -0.085000 3.685000 0.085000 ;
        RECT 3.995000 -0.085000 4.165000 0.085000 ;
        RECT 4.475000 -0.085000 4.645000 0.085000 ;
        RECT 4.955000 -0.085000 5.125000 0.085000 ;
        RECT 5.435000 -0.085000 5.605000 0.085000 ;
        RECT 5.915000 -0.085000 6.085000 0.085000 ;
        RECT 6.395000 -0.085000 6.565000 0.085000 ;
        RECT 6.875000 -0.085000 7.045000 0.085000 ;
        RECT 7.355000 -0.085000 7.525000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.245000 7.680000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 3.245000 7.680000 3.415000 ;
        RECT 0.650000 2.730000 1.025000 3.245000 ;
        RECT 1.595000 2.730000 1.955000 3.245000 ;
        RECT 2.635000 2.730000 2.980000 3.245000 ;
        RECT 3.720000 2.730000 4.050000 3.245000 ;
        RECT 5.180000 2.730000 5.530000 3.245000 ;
        RECT 6.100000 2.730000 6.430000 3.245000 ;
        RECT 7.000000 2.730000 7.565000 3.245000 ;
      LAYER mcon ;
        RECT 0.155000 3.245000 0.325000 3.415000 ;
        RECT 0.635000 3.245000 0.805000 3.415000 ;
        RECT 1.115000 3.245000 1.285000 3.415000 ;
        RECT 1.595000 3.245000 1.765000 3.415000 ;
        RECT 2.075000 3.245000 2.245000 3.415000 ;
        RECT 2.555000 3.245000 2.725000 3.415000 ;
        RECT 3.035000 3.245000 3.205000 3.415000 ;
        RECT 3.515000 3.245000 3.685000 3.415000 ;
        RECT 3.995000 3.245000 4.165000 3.415000 ;
        RECT 4.475000 3.245000 4.645000 3.415000 ;
        RECT 4.955000 3.245000 5.125000 3.415000 ;
        RECT 5.435000 3.245000 5.605000 3.415000 ;
        RECT 5.915000 3.245000 6.085000 3.415000 ;
        RECT 6.395000 3.245000 6.565000 3.415000 ;
        RECT 6.875000 3.245000 7.045000 3.415000 ;
        RECT 7.355000 3.245000 7.525000 3.415000 ;
      LAYER met1 ;
        RECT 0.000000 3.085000 7.680000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.085000 0.450000 0.405000 1.020000 ;
      RECT 0.085000 1.020000 0.255000 1.820000 ;
      RECT 0.085000 1.820000 0.445000 2.390000 ;
      RECT 0.085000 2.390000 7.520000 2.560000 ;
      RECT 0.085000 2.560000 0.445000 2.860000 ;
      RECT 1.485000 1.320000 2.745000 1.650000 ;
      RECT 2.575000 1.650000 2.745000 1.950000 ;
      RECT 2.575000 1.950000 3.515000 1.970000 ;
      RECT 2.575000 1.970000 6.880000 2.220000 ;
      RECT 3.300000 0.605000 3.630000 1.130000 ;
      RECT 3.300000 1.130000 5.475000 1.180000 ;
      RECT 3.460000 1.180000 5.475000 1.300000 ;
      RECT 3.810000 0.630000 4.105000 0.790000 ;
      RECT 3.810000 0.790000 5.125000 0.960000 ;
      RECT 4.795000 0.605000 5.125000 0.790000 ;
      RECT 5.305000 0.255000 7.495000 0.425000 ;
      RECT 5.305000 0.425000 5.475000 1.130000 ;
      RECT 5.650000 1.940000 6.080000 1.970000 ;
      RECT 5.655000 0.595000 6.955000 0.765000 ;
      RECT 5.655000 0.765000 5.905000 0.960000 ;
      RECT 5.910000 1.130000 6.335000 1.300000 ;
      RECT 5.910000 1.300000 6.080000 1.940000 ;
      RECT 6.080000 0.935000 6.335000 1.130000 ;
      RECT 6.250000 1.470000 6.675000 1.800000 ;
      RECT 6.505000 1.130000 7.520000 1.300000 ;
      RECT 6.505000 1.300000 6.675000 1.470000 ;
      RECT 6.625000 0.765000 6.955000 0.935000 ;
      RECT 7.165000 0.425000 7.495000 0.960000 ;
      RECT 7.350000 1.300000 7.520000 2.390000 ;
  END
END sky130_fd_sc_hs__and4b_4
