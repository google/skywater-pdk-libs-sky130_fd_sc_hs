* File: sky130_fd_sc_hs__and3_1.spice
* Created: Thu Aug 27 20:32:15 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hs__and3_1.pex.spice"
.subckt sky130_fd_sc_hs__and3_1  VNB VPB A B C VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* C	C
* B	B
* A	A
* VPB	VPB
* VNB	VNB
MM1003 A_121_136# N_A_M1003_g N_A_27_398#_M1003_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.1312 AS=0.1824 PD=1.05 PS=1.85 NRD=28.116 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75001.7 A=0.096 P=1.58 MULT=1
MM1004 A_233_136# N_B_M1004_g A_121_136# VNB NLOWVT L=0.15 W=0.64 AD=0.111
+ AS=0.1312 PD=1.045 PS=1.05 NRD=22.2 NRS=28.116 M=1 R=4.26667 SA=75000.8
+ SB=75001.1 A=0.096 P=1.58 MULT=1
MM1005 N_VGND_M1005_d N_C_M1005_g A_233_136# VNB NLOWVT L=0.15 W=0.64
+ AD=0.144093 AS=0.111 PD=1.08522 PS=1.045 NRD=15.468 NRS=22.2 M=1 R=4.26667
+ SA=75001.1 SB=75000.8 A=0.096 P=1.58 MULT=1
MM1007 N_X_M1007_d N_A_27_398#_M1007_g N_VGND_M1005_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.166607 PD=2.05 PS=1.25478 NRD=0 NRS=11.34 M=1 R=4.93333
+ SA=75001.5 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1002 N_VPWR_M1002_d N_A_M1002_g N_A_27_398#_M1002_s VPB PSHORT L=0.15 W=0.84
+ AD=0.168 AS=0.2478 PD=1.24 PS=2.27 NRD=14.0658 NRS=2.3443 M=1 R=5.6 SA=75000.2
+ SB=75002.1 A=0.126 P=1.98 MULT=1
MM1006 N_A_27_398#_M1006_d N_B_M1006_g N_VPWR_M1002_d VPB PSHORT L=0.15 W=0.84
+ AD=0.126 AS=0.168 PD=1.14 PS=1.24 NRD=2.3443 NRS=14.0658 M=1 R=5.6 SA=75000.8
+ SB=75001.5 A=0.126 P=1.98 MULT=1
MM1000 N_VPWR_M1000_d N_C_M1000_g N_A_27_398#_M1006_d VPB PSHORT L=0.15 W=0.84
+ AD=0.311336 AS=0.126 PD=1.57714 PS=1.14 NRD=9.9485 NRS=2.3443 M=1 R=5.6
+ SA=75001.2 SB=75001.1 A=0.126 P=1.98 MULT=1
MM1001 N_X_M1001_d N_A_27_398#_M1001_g N_VPWR_M1000_d VPB PSHORT L=0.15 W=1.12
+ AD=0.3304 AS=0.415114 PD=2.83 PS=2.10286 NRD=1.7533 NRS=2.6201 M=1 R=7.46667
+ SA=75001.7 SB=75000.2 A=0.168 P=2.54 MULT=1
DX8_noxref VNB VPB NWDIODE A=6.0636 P=10.24
*
.include "sky130_fd_sc_hs__and3_1.pxi.spice"
*
.ends
*
*
