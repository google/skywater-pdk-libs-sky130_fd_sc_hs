* File: sky130_fd_sc_hs__o32ai_2.pxi.spice
* Created: Thu Aug 27 21:03:53 2020
* 
x_PM_SKY130_FD_SC_HS__O32AI_2%B2 N_B2_M1017_g N_B2_c_101_n N_B2_M1007_g
+ N_B2_M1018_g N_B2_c_102_n N_B2_M1008_g B2 B2 B2 N_B2_c_100_n
+ PM_SKY130_FD_SC_HS__O32AI_2%B2
x_PM_SKY130_FD_SC_HS__O32AI_2%B1 N_B1_c_147_n N_B1_M1011_g N_B1_M1012_g
+ N_B1_c_148_n N_B1_M1013_g N_B1_M1015_g B1 N_B1_c_145_n N_B1_c_146_n
+ PM_SKY130_FD_SC_HS__O32AI_2%B1
x_PM_SKY130_FD_SC_HS__O32AI_2%A3 N_A3_M1009_g N_A3_c_202_n N_A3_M1001_g
+ N_A3_M1010_g N_A3_c_203_n N_A3_M1002_g A3 A3 N_A3_c_201_n
+ PM_SKY130_FD_SC_HS__O32AI_2%A3
x_PM_SKY130_FD_SC_HS__O32AI_2%A2 N_A2_M1016_g N_A2_c_262_n N_A2_M1004_g
+ N_A2_c_263_n N_A2_M1005_g N_A2_M1019_g A2 A2 N_A2_c_261_n
+ PM_SKY130_FD_SC_HS__O32AI_2%A2
x_PM_SKY130_FD_SC_HS__O32AI_2%A1 N_A1_M1006_g N_A1_c_315_n N_A1_M1000_g
+ N_A1_c_316_n N_A1_M1003_g N_A1_M1014_g N_A1_c_311_n A1 A1 A1 A1 N_A1_c_313_n
+ N_A1_c_314_n PM_SKY130_FD_SC_HS__O32AI_2%A1
x_PM_SKY130_FD_SC_HS__O32AI_2%A_27_368# N_A_27_368#_M1007_d N_A_27_368#_M1008_d
+ N_A_27_368#_M1013_s N_A_27_368#_c_357_n N_A_27_368#_c_358_n
+ N_A_27_368#_c_359_n N_A_27_368#_c_373_p N_A_27_368#_c_379_p
+ N_A_27_368#_c_366_n N_A_27_368#_c_360_n PM_SKY130_FD_SC_HS__O32AI_2%A_27_368#
x_PM_SKY130_FD_SC_HS__O32AI_2%Y N_Y_M1017_d N_Y_M1012_s N_Y_M1007_s N_Y_M1001_d
+ N_Y_c_401_n N_Y_c_393_n N_Y_c_394_n N_Y_c_398_n N_Y_c_424_n N_Y_c_395_n
+ N_Y_c_412_n N_Y_c_396_n Y Y N_Y_c_399_n N_Y_c_397_n
+ PM_SKY130_FD_SC_HS__O32AI_2%Y
x_PM_SKY130_FD_SC_HS__O32AI_2%VPWR N_VPWR_M1011_d N_VPWR_M1000_d N_VPWR_M1003_d
+ N_VPWR_c_485_n N_VPWR_c_486_n N_VPWR_c_487_n N_VPWR_c_488_n VPWR
+ N_VPWR_c_489_n N_VPWR_c_490_n N_VPWR_c_491_n N_VPWR_c_492_n N_VPWR_c_493_n
+ N_VPWR_c_484_n PM_SKY130_FD_SC_HS__O32AI_2%VPWR
x_PM_SKY130_FD_SC_HS__O32AI_2%A_499_368# N_A_499_368#_M1001_s
+ N_A_499_368#_M1002_s N_A_499_368#_M1005_s N_A_499_368#_c_550_n
+ N_A_499_368#_c_551_n N_A_499_368#_c_552_n N_A_499_368#_c_559_n
+ N_A_499_368#_c_553_n N_A_499_368#_c_554_n N_A_499_368#_c_555_n
+ PM_SKY130_FD_SC_HS__O32AI_2%A_499_368#
x_PM_SKY130_FD_SC_HS__O32AI_2%A_768_368# N_A_768_368#_M1004_d
+ N_A_768_368#_M1000_s N_A_768_368#_c_588_n N_A_768_368#_c_599_n
+ N_A_768_368#_c_589_n N_A_768_368#_c_592_n
+ PM_SKY130_FD_SC_HS__O32AI_2%A_768_368#
x_PM_SKY130_FD_SC_HS__O32AI_2%A_27_74# N_A_27_74#_M1017_s N_A_27_74#_M1018_s
+ N_A_27_74#_M1015_d N_A_27_74#_M1010_s N_A_27_74#_M1019_s N_A_27_74#_M1014_d
+ N_A_27_74#_c_618_n N_A_27_74#_c_619_n N_A_27_74#_c_620_n N_A_27_74#_c_635_n
+ N_A_27_74#_c_621_n N_A_27_74#_c_641_n N_A_27_74#_c_642_n N_A_27_74#_c_645_n
+ N_A_27_74#_c_646_n N_A_27_74#_c_622_n N_A_27_74#_c_623_n N_A_27_74#_c_624_n
+ N_A_27_74#_c_625_n N_A_27_74#_c_626_n N_A_27_74#_c_627_n N_A_27_74#_c_628_n
+ N_A_27_74#_c_629_n PM_SKY130_FD_SC_HS__O32AI_2%A_27_74#
x_PM_SKY130_FD_SC_HS__O32AI_2%VGND N_VGND_M1009_d N_VGND_M1016_d N_VGND_M1006_s
+ N_VGND_c_709_n N_VGND_c_710_n N_VGND_c_711_n VGND N_VGND_c_712_n
+ N_VGND_c_713_n N_VGND_c_714_n N_VGND_c_715_n N_VGND_c_716_n N_VGND_c_717_n
+ PM_SKY130_FD_SC_HS__O32AI_2%VGND
cc_1 VNB N_B2_M1017_g 0.0312487f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_2 VNB N_B2_M1018_g 0.0234839f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=0.74
cc_3 VNB B2 0.0183784f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.58
cc_4 VNB N_B2_c_100_n 0.0436067f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=1.557
cc_5 VNB N_B1_M1012_g 0.0244803f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_6 VNB N_B1_M1015_g 0.0244812f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=2.4
cc_7 VNB N_B1_c_145_n 0.0015808f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.557
cc_8 VNB N_B1_c_146_n 0.0402233f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.557
cc_9 VNB N_A3_M1009_g 0.0281248f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_10 VNB N_A3_M1010_g 0.0287756f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=0.74
cc_11 VNB A3 0.00626365f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_12 VNB N_A3_c_201_n 0.0601856f $X=-0.19 $Y=-0.245 $X2=0.835 $Y2=1.515
cc_13 VNB N_A2_M1016_g 0.0246043f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_14 VNB N_A2_M1019_g 0.0247047f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=2.4
cc_15 VNB A2 0.00438466f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_16 VNB N_A2_c_261_n 0.0352141f $X=-0.19 $Y=-0.245 $X2=0.835 $Y2=1.515
cc_17 VNB N_A1_M1006_g 0.0305737f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_18 VNB N_A1_M1014_g 0.0393239f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=2.4
cc_19 VNB N_A1_c_311_n 0.00935177f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_20 VNB A1 0.0203068f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A1_c_313_n 0.0219884f $X=-0.19 $Y=-0.245 $X2=0.835 $Y2=1.515
cc_22 VNB N_A1_c_314_n 0.0395739f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_Y_c_393_n 0.00349006f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_Y_c_394_n 0.00229732f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_Y_c_395_n 0.0091475f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=1.557
cc_26 VNB N_Y_c_396_n 0.0033895f $X=-0.19 $Y=-0.245 $X2=0.835 $Y2=1.565
cc_27 VNB N_Y_c_397_n 0.00357335f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_VPWR_c_484_n 0.263193f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_27_74#_c_618_n 0.0288468f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.557
cc_30 VNB N_A_27_74#_c_619_n 0.0026914f $X=-0.19 $Y=-0.245 $X2=0.835 $Y2=1.557
cc_31 VNB N_A_27_74#_c_620_n 0.00931596f $X=-0.19 $Y=-0.245 $X2=0.835 $Y2=1.515
cc_32 VNB N_A_27_74#_c_621_n 0.00501991f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_27_74#_c_622_n 0.00291303f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_27_74#_c_623_n 0.00565856f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_27_74#_c_624_n 0.00280814f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_27_74#_c_625_n 0.017779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_27_74#_c_626_n 0.0277086f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_27_74#_c_627_n 0.00220635f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_27_74#_c_628_n 0.00280429f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_27_74#_c_629_n 0.00725128f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_709_n 0.00582196f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=1.765
cc_42 VNB N_VGND_c_710_n 0.0181004f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_43 VNB N_VGND_c_711_n 0.00616254f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_44 VNB N_VGND_c_712_n 0.0191515f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_VGND_c_713_n 0.334788f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_VGND_c_714_n 0.060757f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_VGND_c_715_n 0.0195534f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_VGND_c_716_n 0.018682f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_VGND_c_717_n 0.0300631f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VPB N_B2_c_101_n 0.0186669f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.765
cc_51 VPB N_B2_c_102_n 0.0147903f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=1.765
cc_52 VPB B2 0.0155943f $X=-0.19 $Y=1.66 $X2=1.115 $Y2=1.58
cc_53 VPB N_B2_c_100_n 0.0231669f $X=-0.19 $Y=1.66 $X2=0.925 $Y2=1.557
cc_54 VPB N_B1_c_147_n 0.0153748f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.35
cc_55 VPB N_B1_c_148_n 0.0190439f $X=-0.19 $Y=1.66 $X2=0.925 $Y2=1.35
cc_56 VPB N_B1_c_145_n 0.00282068f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.557
cc_57 VPB N_B1_c_146_n 0.0198011f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.557
cc_58 VPB N_A3_c_202_n 0.0182852f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.765
cc_59 VPB N_A3_c_203_n 0.0147998f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=1.765
cc_60 VPB A3 0.00852759f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_61 VPB N_A3_c_201_n 0.0333645f $X=-0.19 $Y=1.66 $X2=0.835 $Y2=1.515
cc_62 VPB N_A2_c_262_n 0.0147885f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.765
cc_63 VPB N_A2_c_263_n 0.0183838f $X=-0.19 $Y=1.66 $X2=0.925 $Y2=1.35
cc_64 VPB A2 0.00762542f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_65 VPB N_A2_c_261_n 0.0198333f $X=-0.19 $Y=1.66 $X2=0.835 $Y2=1.515
cc_66 VPB N_A1_c_315_n 0.0180059f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.765
cc_67 VPB N_A1_c_316_n 0.0180207f $X=-0.19 $Y=1.66 $X2=0.925 $Y2=1.35
cc_68 VPB N_A1_c_311_n 0.0048851f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_69 VPB A1 0.0208738f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_70 VPB N_A1_c_313_n 0.0129865f $X=-0.19 $Y=1.66 $X2=0.835 $Y2=1.515
cc_71 VPB N_A1_c_314_n 0.0218282f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_72 VPB N_A_27_368#_c_357_n 0.0354954f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=1.765
cc_73 VPB N_A_27_368#_c_358_n 0.00523584f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_74 VPB N_A_27_368#_c_359_n 0.00935849f $X=-0.19 $Y=1.66 $X2=1.115 $Y2=1.58
cc_75 VPB N_A_27_368#_c_360_n 0.00909276f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=1.557
cc_76 VPB N_Y_c_398_n 0.0120361f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.557
cc_77 VPB N_Y_c_399_n 0.00161209f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_78 VPB N_Y_c_397_n 0.00115845f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_79 VPB N_VPWR_c_485_n 0.00571271f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=1.765
cc_80 VPB N_VPWR_c_486_n 0.0158037f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_81 VPB N_VPWR_c_487_n 0.0107598f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_82 VPB N_VPWR_c_488_n 0.0495498f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_83 VPB N_VPWR_c_489_n 0.037515f $X=-0.19 $Y=1.66 $X2=0.925 $Y2=1.557
cc_84 VPB N_VPWR_c_490_n 0.0760815f $X=-0.19 $Y=1.66 $X2=1.2 $Y2=1.565
cc_85 VPB N_VPWR_c_491_n 0.0197695f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_86 VPB N_VPWR_c_492_n 0.00460249f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_87 VPB N_VPWR_c_493_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_88 VPB N_VPWR_c_484_n 0.0963019f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_89 VPB N_A_499_368#_c_550_n 0.0055749f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=1.765
cc_90 VPB N_A_499_368#_c_551_n 0.0030474f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=2.4
cc_91 VPB N_A_499_368#_c_552_n 0.00455789f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_92 VPB N_A_499_368#_c_553_n 0.00693844f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.557
cc_93 VPB N_A_499_368#_c_554_n 0.00574906f $X=-0.19 $Y=1.66 $X2=0.925 $Y2=1.557
cc_94 VPB N_A_499_368#_c_555_n 0.00123754f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=1.565
cc_95 VPB N_A_768_368#_c_588_n 0.011775f $X=-0.19 $Y=1.66 $X2=0.925 $Y2=0.74
cc_96 VPB N_A_768_368#_c_589_n 0.00261637f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=2.4
cc_97 N_B2_c_102_n N_B1_c_147_n 0.0264665f $X=0.955 $Y=1.765 $X2=-0.19
+ $Y2=-0.245
cc_98 N_B2_M1018_g N_B1_M1012_g 0.0301413f $X=0.925 $Y=0.74 $X2=0 $Y2=0
cc_99 B2 N_B1_c_145_n 0.034285f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_100 N_B2_c_100_n N_B1_c_145_n 2.66807e-19 $X=0.925 $Y=1.557 $X2=0 $Y2=0
cc_101 B2 N_B1_c_146_n 0.00437097f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_102 N_B2_c_100_n N_B1_c_146_n 0.019829f $X=0.925 $Y=1.557 $X2=0 $Y2=0
cc_103 B2 N_A_27_368#_c_357_n 0.0211447f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_104 N_B2_c_100_n N_A_27_368#_c_357_n 2.09582e-19 $X=0.925 $Y=1.557 $X2=0
+ $Y2=0
cc_105 N_B2_c_101_n N_A_27_368#_c_358_n 0.0136535f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_106 N_B2_c_102_n N_A_27_368#_c_358_n 0.012504f $X=0.955 $Y=1.765 $X2=0 $Y2=0
cc_107 N_B2_M1017_g N_Y_c_401_n 0.00516364f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_108 N_B2_M1018_g N_Y_c_401_n 0.00668237f $X=0.925 $Y=0.74 $X2=0 $Y2=0
cc_109 N_B2_M1018_g N_Y_c_393_n 0.00933793f $X=0.925 $Y=0.74 $X2=0 $Y2=0
cc_110 B2 N_Y_c_393_n 0.0344043f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_111 N_B2_c_100_n N_Y_c_393_n 0.00114341f $X=0.925 $Y=1.557 $X2=0 $Y2=0
cc_112 N_B2_M1017_g N_Y_c_394_n 0.00605998f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_113 N_B2_M1018_g N_Y_c_394_n 0.00277595f $X=0.925 $Y=0.74 $X2=0 $Y2=0
cc_114 B2 N_Y_c_394_n 0.0277268f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_115 N_B2_c_100_n N_Y_c_394_n 0.00231375f $X=0.925 $Y=1.557 $X2=0 $Y2=0
cc_116 N_B2_c_102_n N_Y_c_398_n 0.0119563f $X=0.955 $Y=1.765 $X2=0 $Y2=0
cc_117 B2 N_Y_c_398_n 0.0289214f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_118 N_B2_c_101_n N_Y_c_412_n 0.00964697f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_119 N_B2_c_102_n N_Y_c_412_n 0.0089467f $X=0.955 $Y=1.765 $X2=0 $Y2=0
cc_120 B2 N_Y_c_412_n 0.0237598f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_121 N_B2_c_100_n N_Y_c_412_n 0.00144162f $X=0.925 $Y=1.557 $X2=0 $Y2=0
cc_122 N_B2_c_101_n N_VPWR_c_489_n 0.00278271f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_123 N_B2_c_102_n N_VPWR_c_489_n 0.00278271f $X=0.955 $Y=1.765 $X2=0 $Y2=0
cc_124 N_B2_c_101_n N_VPWR_c_484_n 0.00357317f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_125 N_B2_c_102_n N_VPWR_c_484_n 0.00353907f $X=0.955 $Y=1.765 $X2=0 $Y2=0
cc_126 N_B2_M1017_g N_A_27_74#_c_618_n 0.00159289f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_127 B2 N_A_27_74#_c_618_n 0.0178256f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_128 N_B2_c_100_n N_A_27_74#_c_618_n 7.71522e-19 $X=0.925 $Y=1.557 $X2=0 $Y2=0
cc_129 N_B2_M1017_g N_A_27_74#_c_619_n 0.0132764f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_130 N_B2_M1018_g N_A_27_74#_c_619_n 0.0111757f $X=0.925 $Y=0.74 $X2=0 $Y2=0
cc_131 N_B2_M1017_g N_VGND_c_713_n 0.00357086f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_132 N_B2_M1018_g N_VGND_c_713_n 0.0035414f $X=0.925 $Y=0.74 $X2=0 $Y2=0
cc_133 N_B2_M1017_g N_VGND_c_714_n 0.00278271f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_134 N_B2_M1018_g N_VGND_c_714_n 0.00278271f $X=0.925 $Y=0.74 $X2=0 $Y2=0
cc_135 N_B1_M1015_g N_A3_M1009_g 0.0178748f $X=1.925 $Y=0.74 $X2=0 $Y2=0
cc_136 N_B1_c_148_n A3 2.96095e-19 $X=1.855 $Y=1.765 $X2=0 $Y2=0
cc_137 N_B1_c_145_n A3 0.0288593f $X=1.65 $Y=1.515 $X2=0 $Y2=0
cc_138 N_B1_c_146_n A3 0.00603276f $X=1.855 $Y=1.557 $X2=0 $Y2=0
cc_139 N_B1_c_145_n N_A3_c_201_n 2.25325e-19 $X=1.65 $Y=1.515 $X2=0 $Y2=0
cc_140 N_B1_c_146_n N_A3_c_201_n 0.0226324f $X=1.855 $Y=1.557 $X2=0 $Y2=0
cc_141 N_B1_c_147_n N_A_27_368#_c_358_n 0.00125031f $X=1.405 $Y=1.765 $X2=0
+ $Y2=0
cc_142 N_B1_c_147_n N_A_27_368#_c_366_n 0.0124723f $X=1.405 $Y=1.765 $X2=0 $Y2=0
cc_143 N_B1_c_148_n N_A_27_368#_c_366_n 0.0117449f $X=1.855 $Y=1.765 $X2=0 $Y2=0
cc_144 N_B1_c_147_n N_A_27_368#_c_360_n 5.8779e-19 $X=1.405 $Y=1.765 $X2=0 $Y2=0
cc_145 N_B1_c_148_n N_A_27_368#_c_360_n 0.00765353f $X=1.855 $Y=1.765 $X2=0
+ $Y2=0
cc_146 N_B1_M1012_g N_Y_c_401_n 5.09814e-19 $X=1.425 $Y=0.74 $X2=0 $Y2=0
cc_147 N_B1_M1012_g N_Y_c_393_n 0.017016f $X=1.425 $Y=0.74 $X2=0 $Y2=0
cc_148 N_B1_c_145_n N_Y_c_393_n 0.00445816f $X=1.65 $Y=1.515 $X2=0 $Y2=0
cc_149 N_B1_c_146_n N_Y_c_393_n 0.0014099f $X=1.855 $Y=1.557 $X2=0 $Y2=0
cc_150 N_B1_c_147_n N_Y_c_398_n 0.0152274f $X=1.405 $Y=1.765 $X2=0 $Y2=0
cc_151 N_B1_c_148_n N_Y_c_398_n 0.0161939f $X=1.855 $Y=1.765 $X2=0 $Y2=0
cc_152 N_B1_c_145_n N_Y_c_398_n 0.0220806f $X=1.65 $Y=1.515 $X2=0 $Y2=0
cc_153 N_B1_c_146_n N_Y_c_398_n 0.0024691f $X=1.855 $Y=1.557 $X2=0 $Y2=0
cc_154 N_B1_M1015_g N_Y_c_424_n 0.0064205f $X=1.925 $Y=0.74 $X2=0 $Y2=0
cc_155 N_B1_M1015_g N_Y_c_395_n 0.0128778f $X=1.925 $Y=0.74 $X2=0 $Y2=0
cc_156 N_B1_c_147_n N_Y_c_412_n 7.39283e-19 $X=1.405 $Y=1.765 $X2=0 $Y2=0
cc_157 N_B1_M1015_g N_Y_c_396_n 0.00404963f $X=1.925 $Y=0.74 $X2=0 $Y2=0
cc_158 N_B1_c_145_n N_Y_c_396_n 0.0228889f $X=1.65 $Y=1.515 $X2=0 $Y2=0
cc_159 N_B1_c_146_n N_Y_c_396_n 0.00131877f $X=1.855 $Y=1.557 $X2=0 $Y2=0
cc_160 N_B1_c_147_n N_VPWR_c_485_n 0.00651069f $X=1.405 $Y=1.765 $X2=0 $Y2=0
cc_161 N_B1_c_148_n N_VPWR_c_485_n 0.00409001f $X=1.855 $Y=1.765 $X2=0 $Y2=0
cc_162 N_B1_c_147_n N_VPWR_c_489_n 0.00413917f $X=1.405 $Y=1.765 $X2=0 $Y2=0
cc_163 N_B1_c_148_n N_VPWR_c_490_n 0.00445602f $X=1.855 $Y=1.765 $X2=0 $Y2=0
cc_164 N_B1_c_147_n N_VPWR_c_484_n 0.0081781f $X=1.405 $Y=1.765 $X2=0 $Y2=0
cc_165 N_B1_c_148_n N_VPWR_c_484_n 0.00862391f $X=1.855 $Y=1.765 $X2=0 $Y2=0
cc_166 N_B1_c_148_n N_A_499_368#_c_552_n 0.00283598f $X=1.855 $Y=1.765 $X2=0
+ $Y2=0
cc_167 N_B1_M1012_g N_A_27_74#_c_635_n 0.00668986f $X=1.425 $Y=0.74 $X2=0 $Y2=0
cc_168 N_B1_M1015_g N_A_27_74#_c_635_n 5.09814e-19 $X=1.925 $Y=0.74 $X2=0 $Y2=0
cc_169 N_B1_M1012_g N_A_27_74#_c_621_n 0.00831967f $X=1.425 $Y=0.74 $X2=0 $Y2=0
cc_170 N_B1_M1015_g N_A_27_74#_c_621_n 0.011569f $X=1.925 $Y=0.74 $X2=0 $Y2=0
cc_171 N_B1_M1012_g N_A_27_74#_c_627_n 0.00288559f $X=1.425 $Y=0.74 $X2=0 $Y2=0
cc_172 N_B1_M1012_g N_VGND_c_713_n 0.00354796f $X=1.425 $Y=0.74 $X2=0 $Y2=0
cc_173 N_B1_M1015_g N_VGND_c_713_n 0.00354798f $X=1.925 $Y=0.74 $X2=0 $Y2=0
cc_174 N_B1_M1012_g N_VGND_c_714_n 0.00278247f $X=1.425 $Y=0.74 $X2=0 $Y2=0
cc_175 N_B1_M1015_g N_VGND_c_714_n 0.00278271f $X=1.925 $Y=0.74 $X2=0 $Y2=0
cc_176 N_A3_M1010_g N_A2_M1016_g 0.0150421f $X=3.255 $Y=0.74 $X2=0 $Y2=0
cc_177 N_A3_c_203_n N_A2_c_262_n 0.0119933f $X=3.315 $Y=1.765 $X2=0 $Y2=0
cc_178 N_A3_c_201_n A2 0.00520396f $X=3.255 $Y=1.557 $X2=0 $Y2=0
cc_179 N_A3_c_201_n N_A2_c_261_n 0.0257669f $X=3.255 $Y=1.557 $X2=0 $Y2=0
cc_180 N_A3_c_202_n N_Y_c_398_n 0.0188638f $X=2.865 $Y=1.765 $X2=0 $Y2=0
cc_181 A3 N_Y_c_398_n 0.0561123f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_182 N_A3_c_201_n N_Y_c_398_n 0.00215179f $X=3.255 $Y=1.557 $X2=0 $Y2=0
cc_183 N_A3_M1009_g N_Y_c_424_n 8.78205e-19 $X=2.425 $Y=0.74 $X2=0 $Y2=0
cc_184 N_A3_M1009_g N_Y_c_395_n 0.0121505f $X=2.425 $Y=0.74 $X2=0 $Y2=0
cc_185 N_A3_M1010_g N_Y_c_395_n 0.00213938f $X=3.255 $Y=0.74 $X2=0 $Y2=0
cc_186 A3 N_Y_c_395_n 0.0552068f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_187 N_A3_c_201_n N_Y_c_395_n 0.0106165f $X=3.255 $Y=1.557 $X2=0 $Y2=0
cc_188 N_A3_c_202_n Y 0.01464f $X=2.865 $Y=1.765 $X2=0 $Y2=0
cc_189 N_A3_c_203_n Y 0.00890313f $X=3.315 $Y=1.765 $X2=0 $Y2=0
cc_190 N_A3_c_202_n N_Y_c_399_n 0.00655005f $X=2.865 $Y=1.765 $X2=0 $Y2=0
cc_191 N_A3_c_203_n N_Y_c_399_n 0.00501057f $X=3.315 $Y=1.765 $X2=0 $Y2=0
cc_192 N_A3_c_201_n N_Y_c_399_n 0.00732069f $X=3.255 $Y=1.557 $X2=0 $Y2=0
cc_193 N_A3_M1009_g N_Y_c_397_n 0.00299821f $X=2.425 $Y=0.74 $X2=0 $Y2=0
cc_194 N_A3_c_202_n N_Y_c_397_n 0.00213499f $X=2.865 $Y=1.765 $X2=0 $Y2=0
cc_195 N_A3_M1010_g N_Y_c_397_n 0.00459856f $X=3.255 $Y=0.74 $X2=0 $Y2=0
cc_196 N_A3_c_203_n N_Y_c_397_n 9.81445e-19 $X=3.315 $Y=1.765 $X2=0 $Y2=0
cc_197 A3 N_Y_c_397_n 0.0331353f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_198 N_A3_c_201_n N_Y_c_397_n 0.0244276f $X=3.255 $Y=1.557 $X2=0 $Y2=0
cc_199 N_A3_c_202_n N_VPWR_c_490_n 0.00278271f $X=2.865 $Y=1.765 $X2=0 $Y2=0
cc_200 N_A3_c_203_n N_VPWR_c_490_n 0.00278271f $X=3.315 $Y=1.765 $X2=0 $Y2=0
cc_201 N_A3_c_202_n N_VPWR_c_484_n 0.00358624f $X=2.865 $Y=1.765 $X2=0 $Y2=0
cc_202 N_A3_c_203_n N_VPWR_c_484_n 0.00353907f $X=3.315 $Y=1.765 $X2=0 $Y2=0
cc_203 N_A3_c_202_n N_A_499_368#_c_551_n 0.0137046f $X=2.865 $Y=1.765 $X2=0
+ $Y2=0
cc_204 N_A3_c_203_n N_A_499_368#_c_551_n 0.0128006f $X=3.315 $Y=1.765 $X2=0
+ $Y2=0
cc_205 N_A3_M1009_g N_A_27_74#_c_621_n 0.00401363f $X=2.425 $Y=0.74 $X2=0 $Y2=0
cc_206 N_A3_M1009_g N_A_27_74#_c_641_n 0.00816247f $X=2.425 $Y=0.74 $X2=0 $Y2=0
cc_207 N_A3_M1009_g N_A_27_74#_c_642_n 0.00998617f $X=2.425 $Y=0.74 $X2=0 $Y2=0
cc_208 N_A3_M1010_g N_A_27_74#_c_642_n 0.0143601f $X=3.255 $Y=0.74 $X2=0 $Y2=0
cc_209 N_A3_c_201_n N_A_27_74#_c_642_n 9.68617e-19 $X=3.255 $Y=1.557 $X2=0 $Y2=0
cc_210 N_A3_M1009_g N_A_27_74#_c_645_n 0.00134994f $X=2.425 $Y=0.74 $X2=0 $Y2=0
cc_211 N_A3_M1010_g N_A_27_74#_c_646_n 0.00728117f $X=3.255 $Y=0.74 $X2=0 $Y2=0
cc_212 N_A3_M1010_g N_A_27_74#_c_623_n 0.00424559f $X=3.255 $Y=0.74 $X2=0 $Y2=0
cc_213 N_A3_c_201_n N_A_27_74#_c_623_n 0.00292897f $X=3.255 $Y=1.557 $X2=0 $Y2=0
cc_214 N_A3_M1010_g N_A_27_74#_c_628_n 0.0111563f $X=3.255 $Y=0.74 $X2=0 $Y2=0
cc_215 N_A3_M1010_g N_VGND_c_709_n 6.70813e-19 $X=3.255 $Y=0.74 $X2=0 $Y2=0
cc_216 N_A3_M1010_g N_VGND_c_710_n 0.00324657f $X=3.255 $Y=0.74 $X2=0 $Y2=0
cc_217 N_A3_M1009_g N_VGND_c_713_n 0.00413263f $X=2.425 $Y=0.74 $X2=0 $Y2=0
cc_218 N_A3_M1010_g N_VGND_c_713_n 0.00413208f $X=3.255 $Y=0.74 $X2=0 $Y2=0
cc_219 N_A3_M1009_g N_VGND_c_714_n 0.00321293f $X=2.425 $Y=0.74 $X2=0 $Y2=0
cc_220 N_A3_M1009_g N_VGND_c_715_n 0.00303822f $X=2.425 $Y=0.74 $X2=0 $Y2=0
cc_221 N_A3_M1010_g N_VGND_c_715_n 0.00514433f $X=3.255 $Y=0.74 $X2=0 $Y2=0
cc_222 N_A2_M1019_g N_A1_M1006_g 0.0155173f $X=4.23 $Y=0.74 $X2=0 $Y2=0
cc_223 A2 N_A1_c_311_n 2.78011e-19 $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_224 N_A2_c_261_n N_A1_c_311_n 0.0155173f $X=4.215 $Y=1.557 $X2=0 $Y2=0
cc_225 N_A2_c_263_n A1 2.85825e-19 $X=4.215 $Y=1.765 $X2=0 $Y2=0
cc_226 A2 A1 0.0285909f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_227 N_A2_c_261_n A1 0.00519513f $X=4.215 $Y=1.557 $X2=0 $Y2=0
cc_228 N_A2_c_262_n N_Y_c_399_n 7.89967e-19 $X=3.765 $Y=1.765 $X2=0 $Y2=0
cc_229 A2 N_Y_c_397_n 0.0190659f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_230 N_A2_c_261_n N_Y_c_397_n 2.34445e-19 $X=4.215 $Y=1.557 $X2=0 $Y2=0
cc_231 N_A2_c_263_n N_VPWR_c_486_n 0.00191006f $X=4.215 $Y=1.765 $X2=0 $Y2=0
cc_232 N_A2_c_262_n N_VPWR_c_490_n 0.00278271f $X=3.765 $Y=1.765 $X2=0 $Y2=0
cc_233 N_A2_c_263_n N_VPWR_c_490_n 0.00278257f $X=4.215 $Y=1.765 $X2=0 $Y2=0
cc_234 N_A2_c_262_n N_VPWR_c_484_n 0.00353907f $X=3.765 $Y=1.765 $X2=0 $Y2=0
cc_235 N_A2_c_263_n N_VPWR_c_484_n 0.00358623f $X=4.215 $Y=1.765 $X2=0 $Y2=0
cc_236 A2 N_A_499_368#_c_559_n 0.0122873f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_237 N_A2_c_262_n N_A_499_368#_c_553_n 0.0127563f $X=3.765 $Y=1.765 $X2=0
+ $Y2=0
cc_238 N_A2_c_263_n N_A_499_368#_c_553_n 0.0134708f $X=4.215 $Y=1.765 $X2=0
+ $Y2=0
cc_239 N_A2_c_262_n N_A_499_368#_c_554_n 6.14943e-19 $X=3.765 $Y=1.765 $X2=0
+ $Y2=0
cc_240 N_A2_c_263_n N_A_499_368#_c_554_n 0.00786706f $X=4.215 $Y=1.765 $X2=0
+ $Y2=0
cc_241 N_A2_c_263_n N_A_768_368#_c_588_n 0.0175073f $X=4.215 $Y=1.765 $X2=0
+ $Y2=0
cc_242 A2 N_A_768_368#_c_588_n 0.00705005f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_243 N_A2_c_262_n N_A_768_368#_c_592_n 0.00898954f $X=3.765 $Y=1.765 $X2=0
+ $Y2=0
cc_244 N_A2_c_263_n N_A_768_368#_c_592_n 0.00540976f $X=4.215 $Y=1.765 $X2=0
+ $Y2=0
cc_245 A2 N_A_768_368#_c_592_n 0.0193936f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_246 N_A2_c_261_n N_A_768_368#_c_592_n 0.00124582f $X=4.215 $Y=1.557 $X2=0
+ $Y2=0
cc_247 N_A2_M1016_g N_A_27_74#_c_622_n 0.0151193f $X=3.75 $Y=0.74 $X2=0 $Y2=0
cc_248 N_A2_M1019_g N_A_27_74#_c_622_n 0.0165847f $X=4.23 $Y=0.74 $X2=0 $Y2=0
cc_249 A2 N_A_27_74#_c_622_n 0.0423811f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_250 N_A2_c_261_n N_A_27_74#_c_622_n 0.00336308f $X=4.215 $Y=1.557 $X2=0 $Y2=0
cc_251 A2 N_A_27_74#_c_623_n 0.0135252f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_252 N_A2_M1019_g N_A_27_74#_c_624_n 4.71232e-19 $X=4.23 $Y=0.74 $X2=0 $Y2=0
cc_253 N_A2_M1016_g N_A_27_74#_c_628_n 0.00349724f $X=3.75 $Y=0.74 $X2=0 $Y2=0
cc_254 N_A2_M1019_g N_A_27_74#_c_629_n 8.63921e-19 $X=4.23 $Y=0.74 $X2=0 $Y2=0
cc_255 N_A2_M1016_g N_VGND_c_709_n 0.00955922f $X=3.75 $Y=0.74 $X2=0 $Y2=0
cc_256 N_A2_M1019_g N_VGND_c_709_n 0.00230425f $X=4.23 $Y=0.74 $X2=0 $Y2=0
cc_257 N_A2_M1016_g N_VGND_c_710_n 0.00398535f $X=3.75 $Y=0.74 $X2=0 $Y2=0
cc_258 N_A2_M1016_g N_VGND_c_713_n 0.00788205f $X=3.75 $Y=0.74 $X2=0 $Y2=0
cc_259 N_A2_M1019_g N_VGND_c_713_n 0.00908353f $X=4.23 $Y=0.74 $X2=0 $Y2=0
cc_260 N_A2_M1019_g N_VGND_c_716_n 0.00461464f $X=4.23 $Y=0.74 $X2=0 $Y2=0
cc_261 N_A1_c_315_n N_VPWR_c_486_n 0.018269f $X=5.275 $Y=1.765 $X2=0 $Y2=0
cc_262 N_A1_c_316_n N_VPWR_c_488_n 0.00831454f $X=5.73 $Y=1.765 $X2=0 $Y2=0
cc_263 A1 N_VPWR_c_488_n 0.0215956f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_264 N_A1_c_315_n N_VPWR_c_491_n 0.00445602f $X=5.275 $Y=1.765 $X2=0 $Y2=0
cc_265 N_A1_c_316_n N_VPWR_c_491_n 0.00445602f $X=5.73 $Y=1.765 $X2=0 $Y2=0
cc_266 N_A1_c_315_n N_VPWR_c_484_n 0.00861767f $X=5.275 $Y=1.765 $X2=0 $Y2=0
cc_267 N_A1_c_316_n N_VPWR_c_484_n 0.00861148f $X=5.73 $Y=1.765 $X2=0 $Y2=0
cc_268 N_A1_c_315_n N_A_768_368#_c_588_n 0.0139279f $X=5.275 $Y=1.765 $X2=0
+ $Y2=0
cc_269 N_A1_c_311_n N_A_768_368#_c_588_n 0.00303545f $X=4.76 $Y=1.515 $X2=0
+ $Y2=0
cc_270 A1 N_A_768_368#_c_588_n 0.0682409f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_271 N_A1_c_315_n N_A_768_368#_c_599_n 4.27055e-19 $X=5.275 $Y=1.765 $X2=0
+ $Y2=0
cc_272 N_A1_c_316_n N_A_768_368#_c_599_n 0.00203651f $X=5.73 $Y=1.765 $X2=0
+ $Y2=0
cc_273 A1 N_A_768_368#_c_599_n 0.0242018f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_274 N_A1_c_314_n N_A_768_368#_c_599_n 0.00148021f $X=5.73 $Y=1.557 $X2=0
+ $Y2=0
cc_275 N_A1_c_315_n N_A_768_368#_c_589_n 0.0146517f $X=5.275 $Y=1.765 $X2=0
+ $Y2=0
cc_276 N_A1_c_316_n N_A_768_368#_c_589_n 0.00980542f $X=5.73 $Y=1.765 $X2=0
+ $Y2=0
cc_277 N_A1_M1006_g N_A_27_74#_c_624_n 0.0148256f $X=4.685 $Y=0.74 $X2=0 $Y2=0
cc_278 N_A1_M1006_g N_A_27_74#_c_625_n 0.0131906f $X=4.685 $Y=0.74 $X2=0 $Y2=0
cc_279 N_A1_M1014_g N_A_27_74#_c_625_n 0.0153378f $X=5.745 $Y=0.74 $X2=0 $Y2=0
cc_280 A1 N_A_27_74#_c_625_n 0.116536f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_281 N_A1_c_313_n N_A_27_74#_c_625_n 0.0169703f $X=5.185 $Y=1.515 $X2=0 $Y2=0
cc_282 N_A1_M1014_g N_A_27_74#_c_626_n 0.0155483f $X=5.745 $Y=0.74 $X2=0 $Y2=0
cc_283 N_A1_M1006_g N_A_27_74#_c_629_n 0.0016171f $X=4.685 $Y=0.74 $X2=0 $Y2=0
cc_284 A1 N_A_27_74#_c_629_n 0.0169123f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_285 N_A1_M1014_g N_VGND_c_712_n 0.00434272f $X=5.745 $Y=0.74 $X2=0 $Y2=0
cc_286 N_A1_M1006_g N_VGND_c_713_n 0.00825362f $X=4.685 $Y=0.74 $X2=0 $Y2=0
cc_287 N_A1_M1014_g N_VGND_c_713_n 0.00828694f $X=5.745 $Y=0.74 $X2=0 $Y2=0
cc_288 N_A1_M1006_g N_VGND_c_716_n 0.00434272f $X=4.685 $Y=0.74 $X2=0 $Y2=0
cc_289 N_A1_M1006_g N_VGND_c_717_n 0.00539931f $X=4.685 $Y=0.74 $X2=0 $Y2=0
cc_290 N_A1_M1014_g N_VGND_c_717_n 0.00705014f $X=5.745 $Y=0.74 $X2=0 $Y2=0
cc_291 N_A_27_368#_c_358_n N_Y_M1007_s 0.00197722f $X=1.095 $Y=2.99 $X2=0 $Y2=0
cc_292 N_A_27_368#_M1008_d N_Y_c_398_n 0.00417966f $X=1.03 $Y=1.84 $X2=0 $Y2=0
cc_293 N_A_27_368#_M1013_s N_Y_c_398_n 0.00742599f $X=1.93 $Y=1.84 $X2=0 $Y2=0
cc_294 N_A_27_368#_c_373_p N_Y_c_398_n 0.013831f $X=1.18 $Y=2.46 $X2=0 $Y2=0
cc_295 N_A_27_368#_c_366_n N_Y_c_398_n 0.0333042f $X=1.915 $Y=2.375 $X2=0 $Y2=0
cc_296 N_A_27_368#_c_360_n N_Y_c_398_n 0.0221794f $X=2.08 $Y=2.455 $X2=0 $Y2=0
cc_297 N_A_27_368#_c_357_n N_Y_c_412_n 0.0533059f $X=0.28 $Y=2.115 $X2=0 $Y2=0
cc_298 N_A_27_368#_c_358_n N_Y_c_412_n 0.0160777f $X=1.095 $Y=2.99 $X2=0 $Y2=0
cc_299 N_A_27_368#_c_373_p N_Y_c_412_n 0.0123817f $X=1.18 $Y=2.46 $X2=0 $Y2=0
cc_300 N_A_27_368#_c_379_p N_Y_c_412_n 0.0178804f $X=1.18 $Y=2.905 $X2=0 $Y2=0
cc_301 N_A_27_368#_c_366_n N_VPWR_M1011_d 0.00404182f $X=1.915 $Y=2.375
+ $X2=-0.19 $Y2=1.66
cc_302 N_A_27_368#_c_358_n N_VPWR_c_485_n 0.0123543f $X=1.095 $Y=2.99 $X2=0
+ $Y2=0
cc_303 N_A_27_368#_c_379_p N_VPWR_c_485_n 0.0175031f $X=1.18 $Y=2.905 $X2=0
+ $Y2=0
cc_304 N_A_27_368#_c_366_n N_VPWR_c_485_n 0.0154248f $X=1.915 $Y=2.375 $X2=0
+ $Y2=0
cc_305 N_A_27_368#_c_360_n N_VPWR_c_485_n 0.0234974f $X=2.08 $Y=2.455 $X2=0
+ $Y2=0
cc_306 N_A_27_368#_c_358_n N_VPWR_c_489_n 0.0582805f $X=1.095 $Y=2.99 $X2=0
+ $Y2=0
cc_307 N_A_27_368#_c_359_n N_VPWR_c_489_n 0.0179217f $X=0.365 $Y=2.99 $X2=0
+ $Y2=0
cc_308 N_A_27_368#_c_360_n N_VPWR_c_490_n 0.0146094f $X=2.08 $Y=2.455 $X2=0
+ $Y2=0
cc_309 N_A_27_368#_c_358_n N_VPWR_c_484_n 0.0326824f $X=1.095 $Y=2.99 $X2=0
+ $Y2=0
cc_310 N_A_27_368#_c_359_n N_VPWR_c_484_n 0.00971942f $X=0.365 $Y=2.99 $X2=0
+ $Y2=0
cc_311 N_A_27_368#_c_360_n N_VPWR_c_484_n 0.0120527f $X=2.08 $Y=2.455 $X2=0
+ $Y2=0
cc_312 N_A_27_368#_c_360_n N_A_499_368#_c_550_n 0.0412428f $X=2.08 $Y=2.455
+ $X2=0 $Y2=0
cc_313 N_A_27_368#_c_360_n N_A_499_368#_c_552_n 0.00536545f $X=2.08 $Y=2.455
+ $X2=0 $Y2=0
cc_314 N_Y_c_398_n N_VPWR_M1011_d 0.00359488f $X=2.925 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_315 N_Y_c_398_n N_A_499_368#_M1001_s 0.00591542f $X=2.925 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_316 N_Y_c_398_n N_A_499_368#_c_550_n 0.0202359f $X=2.925 $Y=2.035 $X2=0 $Y2=0
cc_317 Y N_A_499_368#_c_550_n 0.0298377f $X=3.035 $Y=2.32 $X2=0 $Y2=0
cc_318 N_Y_M1001_d N_A_499_368#_c_551_n 0.00197722f $X=2.94 $Y=1.84 $X2=0 $Y2=0
cc_319 Y N_A_499_368#_c_551_n 0.0160777f $X=3.035 $Y=2.32 $X2=0 $Y2=0
cc_320 N_Y_c_399_n N_A_499_368#_c_559_n 0.0510995f $X=3.09 $Y=1.985 $X2=0 $Y2=0
cc_321 N_Y_c_393_n N_A_27_74#_M1018_s 0.0025999f $X=1.545 $Y=1.095 $X2=0 $Y2=0
cc_322 N_Y_c_395_n N_A_27_74#_M1015_d 0.00250873f $X=2.925 $Y=1.095 $X2=0 $Y2=0
cc_323 N_Y_c_394_n N_A_27_74#_c_618_n 0.00555794f $X=0.875 $Y=1.095 $X2=0 $Y2=0
cc_324 N_Y_M1017_d N_A_27_74#_c_619_n 0.00182874f $X=0.57 $Y=0.37 $X2=0 $Y2=0
cc_325 N_Y_c_401_n N_A_27_74#_c_619_n 0.0146462f $X=0.71 $Y=0.775 $X2=0 $Y2=0
cc_326 N_Y_c_393_n N_A_27_74#_c_619_n 0.00304353f $X=1.545 $Y=1.095 $X2=0 $Y2=0
cc_327 N_Y_c_393_n N_A_27_74#_c_635_n 0.0194125f $X=1.545 $Y=1.095 $X2=0 $Y2=0
cc_328 N_Y_M1012_s N_A_27_74#_c_621_n 0.0025999f $X=1.5 $Y=0.37 $X2=0 $Y2=0
cc_329 N_Y_c_393_n N_A_27_74#_c_621_n 0.00304353f $X=1.545 $Y=1.095 $X2=0 $Y2=0
cc_330 N_Y_c_424_n N_A_27_74#_c_621_n 0.0180071f $X=1.71 $Y=0.775 $X2=0 $Y2=0
cc_331 N_Y_c_395_n N_A_27_74#_c_621_n 0.00304353f $X=2.925 $Y=1.095 $X2=0 $Y2=0
cc_332 N_Y_c_395_n N_A_27_74#_c_642_n 0.0489623f $X=2.925 $Y=1.095 $X2=0 $Y2=0
cc_333 N_Y_c_395_n N_A_27_74#_c_645_n 0.0208474f $X=2.925 $Y=1.095 $X2=0 $Y2=0
cc_334 N_Y_c_395_n N_A_27_74#_c_623_n 0.0127334f $X=2.925 $Y=1.095 $X2=0 $Y2=0
cc_335 N_Y_c_395_n N_VGND_M1009_d 0.00894066f $X=2.925 $Y=1.095 $X2=-0.19
+ $Y2=-0.245
cc_336 N_VPWR_c_490_n N_A_499_368#_c_551_n 0.0460938f $X=4.835 $Y=3.33 $X2=0
+ $Y2=0
cc_337 N_VPWR_c_484_n N_A_499_368#_c_551_n 0.0260732f $X=6 $Y=3.33 $X2=0 $Y2=0
cc_338 N_VPWR_c_490_n N_A_499_368#_c_552_n 0.0179217f $X=4.835 $Y=3.33 $X2=0
+ $Y2=0
cc_339 N_VPWR_c_484_n N_A_499_368#_c_552_n 0.00971942f $X=6 $Y=3.33 $X2=0 $Y2=0
cc_340 N_VPWR_c_486_n N_A_499_368#_c_553_n 0.0121618f $X=5 $Y=2.455 $X2=0 $Y2=0
cc_341 N_VPWR_c_490_n N_A_499_368#_c_553_n 0.0645908f $X=4.835 $Y=3.33 $X2=0
+ $Y2=0
cc_342 N_VPWR_c_484_n N_A_499_368#_c_553_n 0.0358952f $X=6 $Y=3.33 $X2=0 $Y2=0
cc_343 N_VPWR_c_486_n N_A_499_368#_c_554_n 0.041429f $X=5 $Y=2.455 $X2=0 $Y2=0
cc_344 N_VPWR_c_490_n N_A_499_368#_c_555_n 0.0121867f $X=4.835 $Y=3.33 $X2=0
+ $Y2=0
cc_345 N_VPWR_c_484_n N_A_499_368#_c_555_n 0.00660921f $X=6 $Y=3.33 $X2=0 $Y2=0
cc_346 N_VPWR_M1000_d N_A_768_368#_c_588_n 0.00709867f $X=4.855 $Y=1.84 $X2=0
+ $Y2=0
cc_347 N_VPWR_c_486_n N_A_768_368#_c_588_n 0.025036f $X=5 $Y=2.455 $X2=0 $Y2=0
cc_348 N_VPWR_c_488_n N_A_768_368#_c_599_n 0.0121024f $X=5.955 $Y=2.115 $X2=0
+ $Y2=0
cc_349 N_VPWR_c_486_n N_A_768_368#_c_589_n 0.0267406f $X=5 $Y=2.455 $X2=0 $Y2=0
cc_350 N_VPWR_c_488_n N_A_768_368#_c_589_n 0.0577258f $X=5.955 $Y=2.115 $X2=0
+ $Y2=0
cc_351 N_VPWR_c_491_n N_A_768_368#_c_589_n 0.0147751f $X=5.87 $Y=3.33 $X2=0
+ $Y2=0
cc_352 N_VPWR_c_484_n N_A_768_368#_c_589_n 0.0121637f $X=6 $Y=3.33 $X2=0 $Y2=0
cc_353 N_A_499_368#_c_553_n N_A_768_368#_M1004_d 0.00222494f $X=4.275 $Y=2.99
+ $X2=-0.19 $Y2=1.66
cc_354 N_A_499_368#_M1005_s N_A_768_368#_c_588_n 0.00883045f $X=4.29 $Y=1.84
+ $X2=0 $Y2=0
cc_355 N_A_499_368#_c_554_n N_A_768_368#_c_588_n 0.0219924f $X=4.44 $Y=2.455
+ $X2=0 $Y2=0
cc_356 N_A_499_368#_c_559_n N_A_768_368#_c_592_n 0.0509595f $X=3.54 $Y=2.115
+ $X2=0 $Y2=0
cc_357 N_A_499_368#_c_553_n N_A_768_368#_c_592_n 0.0144323f $X=4.275 $Y=2.99
+ $X2=0 $Y2=0
cc_358 N_A_499_368#_c_554_n N_A_768_368#_c_592_n 0.0298377f $X=4.44 $Y=2.455
+ $X2=0 $Y2=0
cc_359 N_A_27_74#_c_642_n N_VGND_M1009_d 0.0150186f $X=3.305 $Y=0.755 $X2=-0.19
+ $Y2=-0.245
cc_360 N_A_27_74#_c_622_n N_VGND_M1016_d 0.00251619f $X=4.305 $Y=1.095 $X2=0
+ $Y2=0
cc_361 N_A_27_74#_c_625_n N_VGND_M1006_s 0.0122066f $X=5.795 $Y=1.095 $X2=0
+ $Y2=0
cc_362 N_A_27_74#_c_622_n N_VGND_c_709_n 0.0162019f $X=4.305 $Y=1.095 $X2=0
+ $Y2=0
cc_363 N_A_27_74#_c_624_n N_VGND_c_709_n 0.0169744f $X=4.47 $Y=0.515 $X2=0 $Y2=0
cc_364 N_A_27_74#_c_628_n N_VGND_c_709_n 0.0176756f $X=3.47 $Y=0.515 $X2=0 $Y2=0
cc_365 N_A_27_74#_c_642_n N_VGND_c_710_n 0.0023667f $X=3.305 $Y=0.755 $X2=0
+ $Y2=0
cc_366 N_A_27_74#_c_628_n N_VGND_c_710_n 0.0145639f $X=3.47 $Y=0.515 $X2=0 $Y2=0
cc_367 N_A_27_74#_c_626_n N_VGND_c_712_n 0.0145639f $X=5.96 $Y=0.515 $X2=0 $Y2=0
cc_368 N_A_27_74#_c_619_n N_VGND_c_713_n 0.0241933f $X=1.045 $Y=0.34 $X2=0 $Y2=0
cc_369 N_A_27_74#_c_620_n N_VGND_c_713_n 0.00971942f $X=0.365 $Y=0.34 $X2=0
+ $Y2=0
cc_370 N_A_27_74#_c_621_n N_VGND_c_713_n 0.0365966f $X=2.045 $Y=0.34 $X2=0 $Y2=0
cc_371 N_A_27_74#_c_642_n N_VGND_c_713_n 0.0111582f $X=3.305 $Y=0.755 $X2=0
+ $Y2=0
cc_372 N_A_27_74#_c_624_n N_VGND_c_713_n 0.0119984f $X=4.47 $Y=0.515 $X2=0 $Y2=0
cc_373 N_A_27_74#_c_626_n N_VGND_c_713_n 0.0119984f $X=5.96 $Y=0.515 $X2=0 $Y2=0
cc_374 N_A_27_74#_c_627_n N_VGND_c_713_n 0.0126568f $X=1.21 $Y=0.34 $X2=0 $Y2=0
cc_375 N_A_27_74#_c_628_n N_VGND_c_713_n 0.0119984f $X=3.47 $Y=0.515 $X2=0 $Y2=0
cc_376 N_A_27_74#_c_619_n N_VGND_c_714_n 0.0428729f $X=1.045 $Y=0.34 $X2=0 $Y2=0
cc_377 N_A_27_74#_c_620_n N_VGND_c_714_n 0.0179217f $X=0.365 $Y=0.34 $X2=0 $Y2=0
cc_378 N_A_27_74#_c_621_n N_VGND_c_714_n 0.0656076f $X=2.045 $Y=0.34 $X2=0 $Y2=0
cc_379 N_A_27_74#_c_642_n N_VGND_c_714_n 0.00236055f $X=3.305 $Y=0.755 $X2=0
+ $Y2=0
cc_380 N_A_27_74#_c_627_n N_VGND_c_714_n 0.0232598f $X=1.21 $Y=0.34 $X2=0 $Y2=0
cc_381 N_A_27_74#_c_621_n N_VGND_c_715_n 0.0118583f $X=2.045 $Y=0.34 $X2=0 $Y2=0
cc_382 N_A_27_74#_c_642_n N_VGND_c_715_n 0.0433812f $X=3.305 $Y=0.755 $X2=0
+ $Y2=0
cc_383 N_A_27_74#_c_628_n N_VGND_c_715_n 0.00619249f $X=3.47 $Y=0.515 $X2=0
+ $Y2=0
cc_384 N_A_27_74#_c_624_n N_VGND_c_716_n 0.0145639f $X=4.47 $Y=0.515 $X2=0 $Y2=0
cc_385 N_A_27_74#_c_624_n N_VGND_c_717_n 0.0180018f $X=4.47 $Y=0.515 $X2=0 $Y2=0
cc_386 N_A_27_74#_c_625_n N_VGND_c_717_n 0.0561308f $X=5.795 $Y=1.095 $X2=0
+ $Y2=0
cc_387 N_A_27_74#_c_626_n N_VGND_c_717_n 0.0180018f $X=5.96 $Y=0.515 $X2=0 $Y2=0
