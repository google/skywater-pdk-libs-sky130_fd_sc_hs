# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_hs__or2_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__or2_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.320000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.411000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.210000 1.350000 2.755000 1.950000 ;
        RECT 2.520000 1.950000 3.895000 2.120000 ;
        RECT 3.590000 1.450000 3.895000 1.950000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.411000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.925000 1.450000 3.255000 1.780000 ;
    END
  END B
  PIN X
    ANTENNADIFFAREA  1.149300 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 0.960000 1.700000 1.130000 ;
        RECT 0.125000 1.130000 0.355000 1.800000 ;
        RECT 0.125000 1.800000 1.795000 1.970000 ;
        RECT 0.545000 0.350000 0.795000 0.960000 ;
        RECT 0.565000 1.970000 0.895000 2.980000 ;
        RECT 1.405000 0.350000 1.700000 0.960000 ;
        RECT 1.465000 1.970000 1.795000 2.980000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 4.320000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 4.320000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.320000 0.085000 ;
      RECT 0.000000  3.245000 4.320000 3.415000 ;
      RECT 0.115000  0.085000 0.365000 0.790000 ;
      RECT 0.115000  2.140000 0.365000 3.245000 ;
      RECT 0.595000  1.300000 2.040000 1.630000 ;
      RECT 0.975000  0.085000 1.225000 0.790000 ;
      RECT 1.095000  2.140000 1.265000 3.245000 ;
      RECT 1.870000  1.010000 4.235000 1.180000 ;
      RECT 1.870000  1.180000 2.040000 1.300000 ;
      RECT 1.920000  0.085000 2.250000 0.840000 ;
      RECT 1.995000  2.120000 2.245000 3.245000 ;
      RECT 2.420000  0.350000 2.750000 1.010000 ;
      RECT 2.450000  2.290000 2.780000 2.905000 ;
      RECT 2.450000  2.905000 3.730000 3.075000 ;
      RECT 2.920000  0.085000 4.205000 0.840000 ;
      RECT 2.980000  2.290000 4.235000 2.460000 ;
      RECT 2.980000  2.460000 3.230000 2.735000 ;
      RECT 3.400000  2.630000 3.730000 2.905000 ;
      RECT 3.930000  2.630000 4.205000 3.245000 ;
      RECT 4.065000  1.180000 4.235000 2.290000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
  END
END sky130_fd_sc_hs__or2_4
END LIBRARY
