* File: sky130_fd_sc_hs__and4bb_4.spice
* Created: Thu Aug 27 20:34:05 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hs__and4bb_4.pex.spice"
.subckt sky130_fd_sc_hs__and4bb_4  VNB VPB B_N A_N C D VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* D	D
* C	C
* A_N	A_N
* B_N	B_N
* VPB	VPB
* VNB	VNB
MM1020 N_VGND_M1020_d N_B_N_M1020_g N_A_27_74#_M1020_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.0896 AS=0.1824 PD=0.92 PS=1.85 NRD=0 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75000.7 A=0.096 P=1.58 MULT=1
MM1021 N_A_200_74#_M1021_d N_A_N_M1021_g N_VGND_M1020_d VNB NLOWVT L=0.15 W=0.64
+ AD=0.1915 AS=0.0896 PD=1.99 PS=0.92 NRD=13.116 NRS=0 M=1 R=4.26667 SA=75000.6
+ SB=75000.2 A=0.096 P=1.58 MULT=1
MM1007 N_A_472_388#_M1007_d N_A_200_74#_M1007_g N_A_412_140#_M1007_s VNB NLOWVT
+ L=0.15 W=0.64 AD=0.0896 AS=0.2272 PD=0.92 PS=1.99 NRD=0 NRS=13.116 M=1
+ R=4.26667 SA=75000.3 SB=75001.5 A=0.096 P=1.58 MULT=1
MM1027 N_A_472_388#_M1007_d N_A_200_74#_M1027_g N_A_412_140#_M1027_s VNB NLOWVT
+ L=0.15 W=0.64 AD=0.0896 AS=0.0896 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.7 SB=75001.1 A=0.096 P=1.58 MULT=1
MM1000 N_A_685_140#_M1000_d N_A_27_74#_M1000_g N_A_412_140#_M1027_s VNB NLOWVT
+ L=0.15 W=0.64 AD=0.0896 AS=0.0896 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75001.1 SB=75000.6 A=0.096 P=1.58 MULT=1
MM1002 N_A_685_140#_M1000_d N_A_27_74#_M1002_g N_A_412_140#_M1002_s VNB NLOWVT
+ L=0.15 W=0.64 AD=0.0896 AS=0.1824 PD=0.92 PS=1.85 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75001.6 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1001 N_A_685_140#_M1001_d N_C_M1001_g N_A_882_137#_M1001_s VNB NLOWVT L=0.15
+ W=0.64 AD=0.0896 AS=0.2272 PD=0.92 PS=1.99 NRD=0 NRS=13.116 M=1 R=4.26667
+ SA=75000.3 SB=75000.6 A=0.096 P=1.58 MULT=1
MM1022 N_A_685_140#_M1001_d N_C_M1022_g N_A_882_137#_M1022_s VNB NLOWVT L=0.15
+ W=0.64 AD=0.0896 AS=0.1824 PD=0.92 PS=1.85 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.7 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1008 N_VGND_M1008_d N_D_M1008_g N_A_882_137#_M1008_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.1824 AS=0.0896 PD=1.85 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75002.6 A=0.096 P=1.58 MULT=1
MM1023 N_VGND_M1023_d N_D_M1023_g N_A_882_137#_M1008_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.115478 AS=0.0896 PD=1.01101 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667 SA=75000.6
+ SB=75002.1 A=0.096 P=1.58 MULT=1
MM1006 N_VGND_M1023_d N_A_472_388#_M1006_g N_X_M1006_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.133522 AS=0.1036 PD=1.16899 PS=1.02 NRD=11.34 NRS=0 M=1 R=4.93333
+ SA=75001 SB=75001.6 A=0.111 P=1.78 MULT=1
MM1009 N_VGND_M1009_d N_A_472_388#_M1009_g N_X_M1006_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1406 AS=0.1036 PD=1.12 PS=1.02 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75001.4
+ SB=75001.2 A=0.111 P=1.78 MULT=1
MM1014 N_VGND_M1009_d N_A_472_388#_M1014_g N_X_M1014_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1406 AS=0.1184 PD=1.12 PS=1.06 NRD=4.86 NRS=6.48 M=1 R=4.93333 SA=75002
+ SB=75000.7 A=0.111 P=1.78 MULT=1
MM1018 N_VGND_M1018_d N_A_472_388#_M1018_g N_X_M1014_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.2146 AS=0.1184 PD=2.06 PS=1.06 NRD=0 NRS=0 M=1 R=4.93333 SA=75002.4
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1010 N_VPWR_M1010_d N_B_N_M1010_g N_A_27_74#_M1010_s VPB PSHORT L=0.15 W=1
+ AD=0.2 AS=0.295 PD=1.4 PS=2.59 NRD=11.8003 NRS=1.9503 M=1 R=6.66667 SA=75000.2
+ SB=75000.8 A=0.15 P=2.3 MULT=1
MM1005 N_A_200_74#_M1005_d N_A_N_M1005_g N_VPWR_M1010_d VPB PSHORT L=0.15 W=1
+ AD=0.295 AS=0.2 PD=2.59 PS=1.4 NRD=1.9503 NRS=11.8003 M=1 R=6.66667 SA=75000.8
+ SB=75000.2 A=0.15 P=2.3 MULT=1
MM1004 N_A_472_388#_M1004_d N_A_200_74#_M1004_g N_VPWR_M1004_s VPB PSHORT L=0.15
+ W=1 AD=0.235 AS=0.32 PD=1.47 PS=2.64 NRD=18.715 NRS=2.9353 M=1 R=6.66667
+ SA=75000.2 SB=75006.3 A=0.15 P=2.3 MULT=1
MM1024 N_A_472_388#_M1004_d N_A_200_74#_M1024_g N_VPWR_M1024_s VPB PSHORT L=0.15
+ W=1 AD=0.235 AS=0.16 PD=1.47 PS=1.32 NRD=18.715 NRS=1.9503 M=1 R=6.66667
+ SA=75000.9 SB=75005.7 A=0.15 P=2.3 MULT=1
MM1012 N_A_472_388#_M1012_d N_A_27_74#_M1012_g N_VPWR_M1024_s VPB PSHORT L=0.15
+ W=1 AD=0.165 AS=0.16 PD=1.33 PS=1.32 NRD=7.8603 NRS=5.91 M=1 R=6.66667
+ SA=75001.3 SB=75005.2 A=0.15 P=2.3 MULT=1
MM1026 N_A_472_388#_M1012_d N_A_27_74#_M1026_g N_VPWR_M1026_s VPB PSHORT L=0.15
+ W=1 AD=0.165 AS=0.2 PD=1.33 PS=1.4 NRD=1.9503 NRS=11.8003 M=1 R=6.66667
+ SA=75001.8 SB=75004.7 A=0.15 P=2.3 MULT=1
MM1019 N_A_472_388#_M1019_d N_C_M1019_g N_VPWR_M1026_s VPB PSHORT L=0.15 W=1
+ AD=0.15 AS=0.2 PD=1.3 PS=1.4 NRD=1.9503 NRS=11.8003 M=1 R=6.66667 SA=75002.4
+ SB=75004.2 A=0.15 P=2.3 MULT=1
MM1025 N_A_472_388#_M1019_d N_C_M1025_g N_VPWR_M1025_s VPB PSHORT L=0.15 W=1
+ AD=0.15 AS=0.61 PD=1.3 PS=2.22 NRD=1.9503 NRS=11.8003 M=1 R=6.66667 SA=75002.8
+ SB=75003.7 A=0.15 P=2.3 MULT=1
MM1003 N_VPWR_M1025_s N_D_M1003_g N_A_472_388#_M1003_s VPB PSHORT L=0.15 W=1
+ AD=0.61 AS=0.18625 PD=2.22 PS=1.455 NRD=1.9503 NRS=11.8003 M=1 R=6.66667
+ SA=75004.2 SB=75002.4 A=0.15 P=2.3 MULT=1
MM1017 N_VPWR_M1017_d N_D_M1017_g N_A_472_388#_M1003_s VPB PSHORT L=0.15 W=1
+ AD=0.198302 AS=0.18625 PD=1.41981 PS=1.455 NRD=19.1878 NRS=2.9353 M=1
+ R=6.66667 SA=75004.2 SB=75002.1 A=0.15 P=2.3 MULT=1
MM1011 N_X_M1011_d N_A_472_388#_M1011_g N_VPWR_M1017_d VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.222098 PD=1.42 PS=1.59019 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75004.3 SB=75001.6 A=0.168 P=2.54 MULT=1
MM1013 N_X_M1011_d N_A_472_388#_M1013_g N_VPWR_M1013_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75004.7 SB=75001.1 A=0.168 P=2.54 MULT=1
MM1015 N_X_M1015_d N_A_472_388#_M1015_g N_VPWR_M1013_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75005.2 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1016 N_X_M1015_d N_A_472_388#_M1016_g N_VPWR_M1016_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.3304 PD=1.42 PS=2.83 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75005.6 SB=75000.2 A=0.168 P=2.54 MULT=1
DX28_noxref VNB VPB NWDIODE A=17.245 P=22.92
c_84 VNB 0 5.63592e-20 $X=0 $Y=0
*
.include "sky130_fd_sc_hs__and4bb_4.pxi.spice"
*
.ends
*
*
