* File: sky130_fd_sc_hs__nand4bb_1.pxi.spice
* Created: Tue Sep  1 20:10:25 2020
* 
x_PM_SKY130_FD_SC_HS__NAND4BB_1%A_N N_A_N_c_70_n N_A_N_c_71_n N_A_N_c_76_n
+ N_A_N_M1002_g N_A_N_M1005_g A_N N_A_N_c_73_n N_A_N_c_74_n
+ PM_SKY130_FD_SC_HS__NAND4BB_1%A_N
x_PM_SKY130_FD_SC_HS__NAND4BB_1%B_N N_B_N_c_100_n N_B_N_M1011_g N_B_N_M1003_g
+ B_N B_N PM_SKY130_FD_SC_HS__NAND4BB_1%B_N
x_PM_SKY130_FD_SC_HS__NAND4BB_1%A_27_398# N_A_27_398#_M1005_s
+ N_A_27_398#_M1002_s N_A_27_398#_c_130_n N_A_27_398#_M1008_g
+ N_A_27_398#_c_131_n N_A_27_398#_M1007_g N_A_27_398#_c_137_n
+ N_A_27_398#_c_132_n N_A_27_398#_c_133_n N_A_27_398#_c_134_n
+ N_A_27_398#_c_135_n PM_SKY130_FD_SC_HS__NAND4BB_1%A_27_398#
x_PM_SKY130_FD_SC_HS__NAND4BB_1%A_226_398# N_A_226_398#_M1003_d
+ N_A_226_398#_M1011_d N_A_226_398#_c_191_n N_A_226_398#_M1004_g
+ N_A_226_398#_c_192_n N_A_226_398#_M1001_g N_A_226_398#_c_199_n
+ N_A_226_398#_c_193_n N_A_226_398#_c_194_n N_A_226_398#_c_195_n
+ N_A_226_398#_c_201_n N_A_226_398#_c_196_n N_A_226_398#_c_197_n
+ PM_SKY130_FD_SC_HS__NAND4BB_1%A_226_398#
x_PM_SKY130_FD_SC_HS__NAND4BB_1%C N_C_c_262_n N_C_M1010_g N_C_c_263_n
+ N_C_M1000_g C C PM_SKY130_FD_SC_HS__NAND4BB_1%C
x_PM_SKY130_FD_SC_HS__NAND4BB_1%D N_D_M1006_g N_D_c_302_n N_D_M1009_g D
+ N_D_c_303_n PM_SKY130_FD_SC_HS__NAND4BB_1%D
x_PM_SKY130_FD_SC_HS__NAND4BB_1%VPWR N_VPWR_M1002_d N_VPWR_M1008_d
+ N_VPWR_M1000_d N_VPWR_c_336_n N_VPWR_c_337_n N_VPWR_c_338_n N_VPWR_c_339_n
+ N_VPWR_c_340_n N_VPWR_c_341_n N_VPWR_c_342_n VPWR N_VPWR_c_343_n
+ N_VPWR_c_344_n N_VPWR_c_335_n N_VPWR_c_346_n
+ PM_SKY130_FD_SC_HS__NAND4BB_1%VPWR
x_PM_SKY130_FD_SC_HS__NAND4BB_1%Y N_Y_M1007_s N_Y_M1008_s N_Y_M1001_d
+ N_Y_M1009_d N_Y_c_392_n N_Y_c_405_n N_Y_c_424_n N_Y_c_426_n N_Y_c_393_n
+ N_Y_c_394_n N_Y_c_396_n N_Y_c_395_n N_Y_c_398_n N_Y_c_399_n Y N_Y_c_400_n
+ N_Y_c_401_n PM_SKY130_FD_SC_HS__NAND4BB_1%Y
x_PM_SKY130_FD_SC_HS__NAND4BB_1%VGND N_VGND_M1005_d N_VGND_M1006_d
+ N_VGND_c_478_n N_VGND_c_479_n N_VGND_c_480_n VGND N_VGND_c_481_n
+ N_VGND_c_482_n N_VGND_c_483_n PM_SKY130_FD_SC_HS__NAND4BB_1%VGND
cc_1 VNB N_A_N_c_70_n 0.00666993f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.465
cc_2 VNB N_A_N_c_71_n 0.0113864f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.825
cc_3 VNB N_A_N_M1005_g 0.0158898f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=0.97
cc_4 VNB N_A_N_c_73_n 0.0211239f $X=-0.19 $Y=-0.245 $X2=0.315 $Y2=0.42
cc_5 VNB N_A_N_c_74_n 0.0537695f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=0.42
cc_6 VNB N_B_N_c_100_n 0.0181158f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.465
cc_7 VNB N_B_N_M1003_g 0.0307295f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=0.585
cc_8 VNB B_N 0.00795483f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=0.97
cc_9 VNB N_A_27_398#_c_130_n 0.0583008f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=1.375
cc_10 VNB N_A_27_398#_c_131_n 0.0213945f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.375
cc_11 VNB N_A_27_398#_c_132_n 0.0145839f $X=-0.19 $Y=-0.245 $X2=0.302 $Y2=0.42
cc_12 VNB N_A_27_398#_c_133_n 0.0221586f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_27_398#_c_134_n 0.017953f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_27_398#_c_135_n 0.00769994f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_226_398#_c_191_n 0.0184894f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=1.375
cc_16 VNB N_A_226_398#_c_192_n 0.039694f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.375
cc_17 VNB N_A_226_398#_c_193_n 0.00835289f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=0.42
cc_18 VNB N_A_226_398#_c_194_n 0.0023091f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_226_398#_c_195_n 0.00272739f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_226_398#_c_196_n 0.00733291f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_226_398#_c_197_n 0.00896425f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_C_c_262_n 0.0193704f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.465
cc_23 VNB N_C_c_263_n 0.0392521f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.41
cc_24 VNB C 0.00268364f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=1.375
cc_25 VNB N_D_M1006_g 0.0274698f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.915
cc_26 VNB N_D_c_302_n 0.0273786f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.41
cc_27 VNB N_D_c_303_n 0.00476542f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_VPWR_c_335_n 0.183584f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_Y_c_392_n 0.0206563f $X=-0.19 $Y=-0.245 $X2=0.315 $Y2=0.42
cc_30 VNB N_Y_c_393_n 0.0203676f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_Y_c_394_n 0.00111978f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_Y_c_395_n 0.0230393f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_478_n 0.0252046f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.47
cc_34 VNB N_VGND_c_479_n 0.0138117f $X=-0.19 $Y=-0.245 $X2=0.315 $Y2=0.42
cc_35 VNB N_VGND_c_480_n 0.0331513f $X=-0.19 $Y=-0.245 $X2=0.315 $Y2=0.42
cc_36 VNB N_VGND_c_481_n 0.0738552f $X=-0.19 $Y=-0.245 $X2=0.302 $Y2=0.42
cc_37 VNB N_VGND_c_482_n 0.0256348f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_483_n 0.264832f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VPB N_A_N_c_71_n 0.00979675f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.825
cc_40 VPB N_A_N_c_76_n 0.0265516f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.915
cc_41 VPB N_B_N_c_100_n 0.0452516f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.465
cc_42 VPB B_N 0.00759109f $X=-0.19 $Y=1.66 $X2=0.52 $Y2=0.97
cc_43 VPB N_A_27_398#_c_130_n 0.0303873f $X=-0.19 $Y=1.66 $X2=0.52 $Y2=1.375
cc_44 VPB N_A_27_398#_c_137_n 0.0389858f $X=-0.19 $Y=1.66 $X2=0.52 $Y2=0.42
cc_45 VPB N_A_27_398#_c_134_n 0.0149127f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_46 VPB N_A_226_398#_c_192_n 0.0239214f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.375
cc_47 VPB N_A_226_398#_c_199_n 0.0136975f $X=-0.19 $Y=1.66 $X2=0.315 $Y2=0.42
cc_48 VPB N_A_226_398#_c_195_n 0.00388136f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_49 VPB N_A_226_398#_c_201_n 0.0148222f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_50 VPB N_C_c_263_n 0.0243718f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.41
cc_51 VPB N_D_c_302_n 0.0324784f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.41
cc_52 VPB N_D_c_303_n 0.00459222f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_53 VPB N_VPWR_c_336_n 0.0238132f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_54 VPB N_VPWR_c_337_n 0.00694777f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_55 VPB N_VPWR_c_338_n 0.00900305f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_56 VPB N_VPWR_c_339_n 0.0345306f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_57 VPB N_VPWR_c_340_n 0.0078724f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_58 VPB N_VPWR_c_341_n 0.0185368f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_59 VPB N_VPWR_c_342_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_60 VPB N_VPWR_c_343_n 0.0197293f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_61 VPB N_VPWR_c_344_n 0.0216364f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_62 VPB N_VPWR_c_335_n 0.0805128f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_63 VPB N_VPWR_c_346_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_64 VPB N_Y_c_396_n 0.0419693f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_65 VPB N_Y_c_395_n 0.0129696f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_66 VPB N_Y_c_398_n 0.0101976f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_67 VPB N_Y_c_399_n 0.00786683f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_68 VPB N_Y_c_400_n 0.0111426f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_69 VPB N_Y_c_401_n 0.00289722f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_70 N_A_N_c_71_n N_B_N_c_100_n 0.0197784f $X=0.505 $Y=1.825 $X2=-0.19
+ $Y2=-0.245
cc_71 N_A_N_c_76_n N_B_N_c_100_n 0.0220088f $X=0.505 $Y=1.915 $X2=-0.19
+ $Y2=-0.245
cc_72 N_A_N_c_74_n N_B_N_M1003_g 0.02321f $X=0.52 $Y=0.42 $X2=0 $Y2=0
cc_73 N_A_N_c_71_n B_N 0.00387379f $X=0.505 $Y=1.825 $X2=0 $Y2=0
cc_74 N_A_N_c_76_n N_A_27_398#_c_137_n 0.0135766f $X=0.505 $Y=1.915 $X2=0 $Y2=0
cc_75 N_A_N_M1005_g N_A_27_398#_c_132_n 0.0154362f $X=0.52 $Y=0.97 $X2=0 $Y2=0
cc_76 N_A_N_c_73_n N_A_27_398#_c_132_n 2.7753e-19 $X=0.315 $Y=0.42 $X2=0 $Y2=0
cc_77 N_A_N_c_70_n N_A_27_398#_c_133_n 0.00111185f $X=0.505 $Y=1.465 $X2=0 $Y2=0
cc_78 N_A_N_M1005_g N_A_27_398#_c_133_n 0.00814439f $X=0.52 $Y=0.97 $X2=0 $Y2=0
cc_79 N_A_N_c_73_n N_A_27_398#_c_133_n 0.0263917f $X=0.315 $Y=0.42 $X2=0 $Y2=0
cc_80 N_A_N_c_74_n N_A_27_398#_c_133_n 0.0016705f $X=0.52 $Y=0.42 $X2=0 $Y2=0
cc_81 N_A_N_c_70_n N_A_27_398#_c_134_n 0.0151079f $X=0.505 $Y=1.465 $X2=0 $Y2=0
cc_82 N_A_N_c_76_n N_A_27_398#_c_134_n 0.00189951f $X=0.505 $Y=1.915 $X2=0 $Y2=0
cc_83 N_A_N_M1005_g N_A_27_398#_c_134_n 0.00257859f $X=0.52 $Y=0.97 $X2=0 $Y2=0
cc_84 N_A_N_c_76_n N_VPWR_c_336_n 0.00859659f $X=0.505 $Y=1.915 $X2=0 $Y2=0
cc_85 N_A_N_c_76_n N_VPWR_c_343_n 0.00475875f $X=0.505 $Y=1.915 $X2=0 $Y2=0
cc_86 N_A_N_c_76_n N_VPWR_c_335_n 0.00505379f $X=0.505 $Y=1.915 $X2=0 $Y2=0
cc_87 N_A_N_c_73_n N_VGND_c_478_n 0.0329753f $X=0.315 $Y=0.42 $X2=0 $Y2=0
cc_88 N_A_N_c_74_n N_VGND_c_478_n 0.0111733f $X=0.52 $Y=0.42 $X2=0 $Y2=0
cc_89 N_A_N_c_73_n N_VGND_c_482_n 0.0233084f $X=0.315 $Y=0.42 $X2=0 $Y2=0
cc_90 N_A_N_c_74_n N_VGND_c_482_n 0.00654921f $X=0.52 $Y=0.42 $X2=0 $Y2=0
cc_91 N_A_N_c_73_n N_VGND_c_483_n 0.0133606f $X=0.315 $Y=0.42 $X2=0 $Y2=0
cc_92 N_A_N_c_74_n N_VGND_c_483_n 0.0041842f $X=0.52 $Y=0.42 $X2=0 $Y2=0
cc_93 N_B_N_M1003_g N_A_27_398#_c_130_n 0.00760094f $X=1.1 $Y=0.925 $X2=0 $Y2=0
cc_94 B_N N_A_27_398#_c_130_n 0.00697096f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_95 N_B_N_c_100_n N_A_27_398#_c_132_n 0.00423441f $X=1.055 $Y=1.915 $X2=0
+ $Y2=0
cc_96 N_B_N_M1003_g N_A_27_398#_c_132_n 0.0161954f $X=1.1 $Y=0.925 $X2=0 $Y2=0
cc_97 B_N N_A_27_398#_c_132_n 0.0543686f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_98 N_B_N_M1003_g N_A_27_398#_c_133_n 7.96521e-19 $X=1.1 $Y=0.925 $X2=0 $Y2=0
cc_99 B_N N_A_27_398#_c_134_n 0.0178516f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_100 N_B_N_M1003_g N_A_27_398#_c_135_n 0.00116302f $X=1.1 $Y=0.925 $X2=0 $Y2=0
cc_101 B_N N_A_27_398#_c_135_n 0.00375077f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_102 N_B_N_c_100_n N_A_226_398#_c_201_n 0.0142503f $X=1.055 $Y=1.915 $X2=0
+ $Y2=0
cc_103 B_N N_A_226_398#_c_201_n 0.0173768f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_104 N_B_N_M1003_g N_A_226_398#_c_196_n 0.00452024f $X=1.1 $Y=0.925 $X2=0
+ $Y2=0
cc_105 N_B_N_c_100_n N_VPWR_c_336_n 0.0109025f $X=1.055 $Y=1.915 $X2=0 $Y2=0
cc_106 B_N N_VPWR_c_336_n 0.0286067f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_107 N_B_N_c_100_n N_VPWR_c_339_n 0.00475875f $X=1.055 $Y=1.915 $X2=0 $Y2=0
cc_108 N_B_N_c_100_n N_VPWR_c_335_n 0.00505379f $X=1.055 $Y=1.915 $X2=0 $Y2=0
cc_109 N_B_N_M1003_g N_Y_c_392_n 0.00275122f $X=1.1 $Y=0.925 $X2=0 $Y2=0
cc_110 N_B_N_c_100_n N_Y_c_398_n 0.00412288f $X=1.055 $Y=1.915 $X2=0 $Y2=0
cc_111 N_B_N_M1003_g N_VGND_c_478_n 0.00535347f $X=1.1 $Y=0.925 $X2=0 $Y2=0
cc_112 N_B_N_M1003_g N_VGND_c_481_n 0.00387193f $X=1.1 $Y=0.925 $X2=0 $Y2=0
cc_113 N_B_N_M1003_g N_VGND_c_483_n 0.00462577f $X=1.1 $Y=0.925 $X2=0 $Y2=0
cc_114 N_A_27_398#_c_132_n N_A_226_398#_M1003_d 0.00232397f $X=1.685 $Y=1.215
+ $X2=-0.19 $Y2=-0.245
cc_115 N_A_27_398#_c_131_n N_A_226_398#_c_191_n 0.0341467f $X=2.1 $Y=1.22 $X2=0
+ $Y2=0
cc_116 N_A_27_398#_c_130_n N_A_226_398#_c_192_n 0.0638771f $X=2.065 $Y=1.765
+ $X2=0 $Y2=0
cc_117 N_A_27_398#_c_135_n N_A_226_398#_c_192_n 2.21999e-19 $X=1.85 $Y=1.215
+ $X2=0 $Y2=0
cc_118 N_A_27_398#_c_130_n N_A_226_398#_c_199_n 0.0181409f $X=2.065 $Y=1.765
+ $X2=0 $Y2=0
cc_119 N_A_27_398#_c_132_n N_A_226_398#_c_199_n 0.00691896f $X=1.685 $Y=1.215
+ $X2=0 $Y2=0
cc_120 N_A_27_398#_c_135_n N_A_226_398#_c_199_n 0.0111894f $X=1.85 $Y=1.215
+ $X2=0 $Y2=0
cc_121 N_A_27_398#_c_130_n N_A_226_398#_c_193_n 0.00174052f $X=2.065 $Y=1.765
+ $X2=0 $Y2=0
cc_122 N_A_27_398#_c_131_n N_A_226_398#_c_193_n 0.0162635f $X=2.1 $Y=1.22 $X2=0
+ $Y2=0
cc_123 N_A_27_398#_c_135_n N_A_226_398#_c_193_n 0.0246367f $X=1.85 $Y=1.215
+ $X2=0 $Y2=0
cc_124 N_A_27_398#_c_131_n N_A_226_398#_c_194_n 0.00171321f $X=2.1 $Y=1.22 $X2=0
+ $Y2=0
cc_125 N_A_27_398#_c_135_n N_A_226_398#_c_194_n 0.00713039f $X=1.85 $Y=1.215
+ $X2=0 $Y2=0
cc_126 N_A_27_398#_c_130_n N_A_226_398#_c_195_n 0.00847786f $X=2.065 $Y=1.765
+ $X2=0 $Y2=0
cc_127 N_A_27_398#_c_130_n N_A_226_398#_c_201_n 0.00390716f $X=2.065 $Y=1.765
+ $X2=0 $Y2=0
cc_128 N_A_27_398#_c_132_n N_A_226_398#_c_201_n 0.00419957f $X=1.685 $Y=1.215
+ $X2=0 $Y2=0
cc_129 N_A_27_398#_c_131_n N_A_226_398#_c_196_n 0.00302206f $X=2.1 $Y=1.22 $X2=0
+ $Y2=0
cc_130 N_A_27_398#_c_132_n N_A_226_398#_c_196_n 0.0362968f $X=1.685 $Y=1.215
+ $X2=0 $Y2=0
cc_131 N_A_27_398#_c_130_n N_A_226_398#_c_197_n 0.00305474f $X=2.065 $Y=1.765
+ $X2=0 $Y2=0
cc_132 N_A_27_398#_c_135_n N_A_226_398#_c_197_n 0.0272167f $X=1.85 $Y=1.215
+ $X2=0 $Y2=0
cc_133 N_A_27_398#_c_137_n N_VPWR_c_336_n 0.0345631f $X=0.28 $Y=2.135 $X2=0
+ $Y2=0
cc_134 N_A_27_398#_c_130_n N_VPWR_c_337_n 0.00559083f $X=2.065 $Y=1.765 $X2=0
+ $Y2=0
cc_135 N_A_27_398#_c_130_n N_VPWR_c_339_n 0.00445602f $X=2.065 $Y=1.765 $X2=0
+ $Y2=0
cc_136 N_A_27_398#_c_137_n N_VPWR_c_343_n 0.00953144f $X=0.28 $Y=2.135 $X2=0
+ $Y2=0
cc_137 N_A_27_398#_c_130_n N_VPWR_c_335_n 0.00460285f $X=2.065 $Y=1.765 $X2=0
+ $Y2=0
cc_138 N_A_27_398#_c_137_n N_VPWR_c_335_n 0.0111133f $X=0.28 $Y=2.135 $X2=0
+ $Y2=0
cc_139 N_A_27_398#_c_131_n N_Y_c_392_n 0.0104202f $X=2.1 $Y=1.22 $X2=0 $Y2=0
cc_140 N_A_27_398#_c_130_n N_Y_c_405_n 0.00956746f $X=2.065 $Y=1.765 $X2=0 $Y2=0
cc_141 N_A_27_398#_c_130_n N_Y_c_398_n 0.00749136f $X=2.065 $Y=1.765 $X2=0 $Y2=0
cc_142 N_A_27_398#_c_132_n N_VGND_M1005_d 0.00380084f $X=1.685 $Y=1.215
+ $X2=-0.19 $Y2=-0.245
cc_143 N_A_27_398#_c_132_n N_VGND_c_478_n 0.0257093f $X=1.685 $Y=1.215 $X2=0
+ $Y2=0
cc_144 N_A_27_398#_c_131_n N_VGND_c_481_n 0.00291649f $X=2.1 $Y=1.22 $X2=0 $Y2=0
cc_145 N_A_27_398#_c_131_n N_VGND_c_483_n 0.0036383f $X=2.1 $Y=1.22 $X2=0 $Y2=0
cc_146 N_A_27_398#_c_133_n N_VGND_c_483_n 9.95189e-19 $X=0.47 $Y=1.07 $X2=0
+ $Y2=0
cc_147 N_A_226_398#_c_191_n N_C_c_262_n 0.0275008f $X=2.49 $Y=1.22 $X2=-0.19
+ $Y2=-0.245
cc_148 N_A_226_398#_c_192_n N_C_c_263_n 0.0522003f $X=2.655 $Y=1.765 $X2=0 $Y2=0
cc_149 N_A_226_398#_c_197_n N_C_c_263_n 0.00120656f $X=2.58 $Y=1.385 $X2=0 $Y2=0
cc_150 N_A_226_398#_c_191_n C 0.00159237f $X=2.49 $Y=1.22 $X2=0 $Y2=0
cc_151 N_A_226_398#_c_192_n C 4.19484e-19 $X=2.655 $Y=1.765 $X2=0 $Y2=0
cc_152 N_A_226_398#_c_193_n C 0.00438395f $X=2.185 $Y=0.875 $X2=0 $Y2=0
cc_153 N_A_226_398#_c_194_n C 0.00690774f $X=2.27 $Y=1.22 $X2=0 $Y2=0
cc_154 N_A_226_398#_c_197_n C 0.0195437f $X=2.58 $Y=1.385 $X2=0 $Y2=0
cc_155 N_A_226_398#_c_199_n N_VPWR_M1008_d 0.00357423f $X=2.185 $Y=2.055 $X2=0
+ $Y2=0
cc_156 N_A_226_398#_c_195_n N_VPWR_M1008_d 0.00134413f $X=2.27 $Y=1.97 $X2=0
+ $Y2=0
cc_157 N_A_226_398#_c_201_n N_VPWR_c_336_n 0.0353488f $X=1.28 $Y=2.135 $X2=0
+ $Y2=0
cc_158 N_A_226_398#_c_192_n N_VPWR_c_337_n 0.00767028f $X=2.655 $Y=1.765 $X2=0
+ $Y2=0
cc_159 N_A_226_398#_c_201_n N_VPWR_c_339_n 0.00953144f $X=1.28 $Y=2.135 $X2=0
+ $Y2=0
cc_160 N_A_226_398#_c_192_n N_VPWR_c_341_n 0.00413917f $X=2.655 $Y=1.765 $X2=0
+ $Y2=0
cc_161 N_A_226_398#_c_192_n N_VPWR_c_335_n 0.00417051f $X=2.655 $Y=1.765 $X2=0
+ $Y2=0
cc_162 N_A_226_398#_c_201_n N_VPWR_c_335_n 0.0111133f $X=1.28 $Y=2.135 $X2=0
+ $Y2=0
cc_163 N_A_226_398#_c_193_n N_Y_M1007_s 0.00433781f $X=2.185 $Y=0.875 $X2=-0.19
+ $Y2=-0.245
cc_164 N_A_226_398#_c_199_n N_Y_M1008_s 0.00683753f $X=2.185 $Y=2.055 $X2=0
+ $Y2=0
cc_165 N_A_226_398#_c_191_n N_Y_c_392_n 0.016417f $X=2.49 $Y=1.22 $X2=0 $Y2=0
cc_166 N_A_226_398#_c_192_n N_Y_c_392_n 0.00318569f $X=2.655 $Y=1.765 $X2=0
+ $Y2=0
cc_167 N_A_226_398#_c_193_n N_Y_c_392_n 0.0380801f $X=2.185 $Y=0.875 $X2=0 $Y2=0
cc_168 N_A_226_398#_c_197_n N_Y_c_392_n 0.00927084f $X=2.58 $Y=1.385 $X2=0 $Y2=0
cc_169 N_A_226_398#_c_199_n N_Y_c_405_n 0.0217794f $X=2.185 $Y=2.055 $X2=0 $Y2=0
cc_170 N_A_226_398#_c_192_n N_Y_c_398_n 7.50322e-19 $X=2.655 $Y=1.765 $X2=0
+ $Y2=0
cc_171 N_A_226_398#_c_199_n N_Y_c_398_n 0.0221264f $X=2.185 $Y=2.055 $X2=0 $Y2=0
cc_172 N_A_226_398#_c_201_n N_Y_c_398_n 0.0370729f $X=1.28 $Y=2.135 $X2=0 $Y2=0
cc_173 N_A_226_398#_c_192_n N_Y_c_400_n 0.0323345f $X=2.655 $Y=1.765 $X2=0 $Y2=0
cc_174 N_A_226_398#_c_195_n N_Y_c_400_n 0.00629661f $X=2.27 $Y=1.97 $X2=0 $Y2=0
cc_175 N_A_226_398#_c_197_n N_Y_c_400_n 0.0123502f $X=2.58 $Y=1.385 $X2=0 $Y2=0
cc_176 N_A_226_398#_c_192_n N_Y_c_401_n 0.00272481f $X=2.655 $Y=1.765 $X2=0
+ $Y2=0
cc_177 N_A_226_398#_c_196_n N_VGND_c_478_n 0.0138983f $X=1.49 $Y=0.795 $X2=0
+ $Y2=0
cc_178 N_A_226_398#_c_191_n N_VGND_c_481_n 0.00291649f $X=2.49 $Y=1.22 $X2=0
+ $Y2=0
cc_179 N_A_226_398#_c_196_n N_VGND_c_481_n 0.00651976f $X=1.49 $Y=0.795 $X2=0
+ $Y2=0
cc_180 N_A_226_398#_c_191_n N_VGND_c_483_n 0.00360083f $X=2.49 $Y=1.22 $X2=0
+ $Y2=0
cc_181 N_A_226_398#_c_193_n N_VGND_c_483_n 0.00894977f $X=2.185 $Y=0.875 $X2=0
+ $Y2=0
cc_182 N_A_226_398#_c_196_n N_VGND_c_483_n 0.00998901f $X=1.49 $Y=0.795 $X2=0
+ $Y2=0
cc_183 N_A_226_398#_c_193_n A_435_74# 0.0037689f $X=2.185 $Y=0.875 $X2=-0.19
+ $Y2=-0.245
cc_184 N_A_226_398#_c_194_n A_435_74# 0.00207986f $X=2.27 $Y=1.22 $X2=-0.19
+ $Y2=-0.245
cc_185 N_C_c_262_n N_D_M1006_g 0.0253098f $X=3.06 $Y=1.22 $X2=0 $Y2=0
cc_186 N_C_c_263_n N_D_M1006_g 0.0177788f $X=3.155 $Y=1.765 $X2=0 $Y2=0
cc_187 C N_D_M1006_g 0.00297693f $X=3.035 $Y=0.84 $X2=0 $Y2=0
cc_188 N_C_c_263_n N_D_c_302_n 0.0387693f $X=3.155 $Y=1.765 $X2=0 $Y2=0
cc_189 C N_D_c_302_n 2.21387e-19 $X=3.035 $Y=0.84 $X2=0 $Y2=0
cc_190 N_C_c_263_n N_D_c_303_n 0.00654791f $X=3.155 $Y=1.765 $X2=0 $Y2=0
cc_191 C N_D_c_303_n 0.0160735f $X=3.035 $Y=0.84 $X2=0 $Y2=0
cc_192 N_C_c_263_n N_VPWR_c_337_n 4.24137e-19 $X=3.155 $Y=1.765 $X2=0 $Y2=0
cc_193 N_C_c_263_n N_VPWR_c_338_n 0.00598632f $X=3.155 $Y=1.765 $X2=0 $Y2=0
cc_194 N_C_c_263_n N_VPWR_c_341_n 0.00445602f $X=3.155 $Y=1.765 $X2=0 $Y2=0
cc_195 N_C_c_263_n N_VPWR_c_335_n 0.00858339f $X=3.155 $Y=1.765 $X2=0 $Y2=0
cc_196 N_C_c_262_n N_Y_c_392_n 0.01594f $X=3.06 $Y=1.22 $X2=0 $Y2=0
cc_197 N_C_c_263_n N_Y_c_392_n 4.92344e-19 $X=3.155 $Y=1.765 $X2=0 $Y2=0
cc_198 C N_Y_c_392_n 0.0193446f $X=3.035 $Y=0.84 $X2=0 $Y2=0
cc_199 N_C_c_263_n N_Y_c_424_n 0.0144039f $X=3.155 $Y=1.765 $X2=0 $Y2=0
cc_200 C N_Y_c_424_n 0.00744175f $X=3.035 $Y=0.84 $X2=0 $Y2=0
cc_201 N_C_c_262_n N_Y_c_426_n 0.00381676f $X=3.06 $Y=1.22 $X2=0 $Y2=0
cc_202 C N_Y_c_426_n 0.0152478f $X=3.035 $Y=0.84 $X2=0 $Y2=0
cc_203 N_C_c_262_n N_Y_c_394_n 4.96616e-19 $X=3.06 $Y=1.22 $X2=0 $Y2=0
cc_204 C N_Y_c_394_n 0.0147075f $X=3.035 $Y=0.84 $X2=0 $Y2=0
cc_205 N_C_c_263_n N_Y_c_396_n 6.61384e-19 $X=3.155 $Y=1.765 $X2=0 $Y2=0
cc_206 N_C_c_263_n N_Y_c_400_n 0.0105243f $X=3.155 $Y=1.765 $X2=0 $Y2=0
cc_207 C N_Y_c_400_n 0.00673483f $X=3.035 $Y=0.84 $X2=0 $Y2=0
cc_208 N_C_c_263_n N_Y_c_401_n 0.00546834f $X=3.155 $Y=1.765 $X2=0 $Y2=0
cc_209 N_C_c_262_n N_VGND_c_481_n 0.00291649f $X=3.06 $Y=1.22 $X2=0 $Y2=0
cc_210 N_C_c_262_n N_VGND_c_483_n 0.00360678f $X=3.06 $Y=1.22 $X2=0 $Y2=0
cc_211 C A_627_74# 0.00402242f $X=3.035 $Y=0.84 $X2=-0.19 $Y2=-0.245
cc_212 N_D_c_302_n N_VPWR_c_338_n 0.00737447f $X=3.705 $Y=1.765 $X2=0 $Y2=0
cc_213 N_D_c_302_n N_VPWR_c_344_n 0.00445602f $X=3.705 $Y=1.765 $X2=0 $Y2=0
cc_214 N_D_c_302_n N_VPWR_c_335_n 0.00861631f $X=3.705 $Y=1.765 $X2=0 $Y2=0
cc_215 N_D_M1006_g N_Y_c_392_n 0.00950424f $X=3.63 $Y=0.74 $X2=0 $Y2=0
cc_216 N_D_c_302_n N_Y_c_424_n 0.0126927f $X=3.705 $Y=1.765 $X2=0 $Y2=0
cc_217 N_D_c_303_n N_Y_c_424_n 0.0193106f $X=3.72 $Y=1.515 $X2=0 $Y2=0
cc_218 N_D_M1006_g N_Y_c_426_n 0.0144061f $X=3.63 $Y=0.74 $X2=0 $Y2=0
cc_219 N_D_M1006_g N_Y_c_393_n 0.00742328f $X=3.63 $Y=0.74 $X2=0 $Y2=0
cc_220 N_D_c_302_n N_Y_c_393_n 0.00125438f $X=3.705 $Y=1.765 $X2=0 $Y2=0
cc_221 N_D_c_303_n N_Y_c_393_n 0.0174298f $X=3.72 $Y=1.515 $X2=0 $Y2=0
cc_222 N_D_M1006_g N_Y_c_394_n 0.0044161f $X=3.63 $Y=0.74 $X2=0 $Y2=0
cc_223 N_D_c_303_n N_Y_c_394_n 0.0144298f $X=3.72 $Y=1.515 $X2=0 $Y2=0
cc_224 N_D_c_302_n N_Y_c_396_n 0.010491f $X=3.705 $Y=1.765 $X2=0 $Y2=0
cc_225 N_D_M1006_g N_Y_c_395_n 0.00477786f $X=3.63 $Y=0.74 $X2=0 $Y2=0
cc_226 N_D_c_302_n N_Y_c_395_n 0.0126891f $X=3.705 $Y=1.765 $X2=0 $Y2=0
cc_227 N_D_c_303_n N_Y_c_395_n 0.0332222f $X=3.72 $Y=1.515 $X2=0 $Y2=0
cc_228 N_D_c_302_n N_Y_c_399_n 8.69057e-19 $X=3.705 $Y=1.765 $X2=0 $Y2=0
cc_229 N_D_c_303_n N_Y_c_399_n 0.00785128f $X=3.72 $Y=1.515 $X2=0 $Y2=0
cc_230 N_D_c_302_n N_Y_c_400_n 0.00133283f $X=3.705 $Y=1.765 $X2=0 $Y2=0
cc_231 N_D_M1006_g N_VGND_c_480_n 0.0143888f $X=3.63 $Y=0.74 $X2=0 $Y2=0
cc_232 N_D_M1006_g N_VGND_c_481_n 0.00348163f $X=3.63 $Y=0.74 $X2=0 $Y2=0
cc_233 N_D_M1006_g N_VGND_c_483_n 0.00547865f $X=3.63 $Y=0.74 $X2=0 $Y2=0
cc_234 N_VPWR_M1008_d N_Y_c_405_n 0.0122439f $X=2.14 $Y=1.84 $X2=0 $Y2=0
cc_235 N_VPWR_c_337_n N_Y_c_405_n 0.0259636f $X=2.385 $Y=2.815 $X2=0 $Y2=0
cc_236 N_VPWR_c_335_n N_Y_c_405_n 0.00598063f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_237 N_VPWR_M1000_d N_Y_c_424_n 0.0112207f $X=3.23 $Y=1.84 $X2=0 $Y2=0
cc_238 N_VPWR_c_338_n N_Y_c_424_n 0.0232685f $X=3.43 $Y=2.455 $X2=0 $Y2=0
cc_239 N_VPWR_c_338_n N_Y_c_396_n 0.0280303f $X=3.43 $Y=2.455 $X2=0 $Y2=0
cc_240 N_VPWR_c_344_n N_Y_c_396_n 0.0203945f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_241 N_VPWR_c_335_n N_Y_c_396_n 0.0168479f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_242 N_VPWR_c_337_n N_Y_c_398_n 0.0132022f $X=2.385 $Y=2.815 $X2=0 $Y2=0
cc_243 N_VPWR_c_339_n N_Y_c_398_n 0.0145781f $X=2.175 $Y=3.33 $X2=0 $Y2=0
cc_244 N_VPWR_c_335_n N_Y_c_398_n 0.0120405f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_245 N_VPWR_c_337_n N_Y_c_400_n 0.00111275f $X=2.385 $Y=2.815 $X2=0 $Y2=0
cc_246 N_VPWR_c_338_n N_Y_c_400_n 0.0272647f $X=3.43 $Y=2.455 $X2=0 $Y2=0
cc_247 N_VPWR_c_335_n N_Y_c_400_n 0.00585815f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_248 N_VPWR_c_337_n N_Y_c_401_n 0.0136383f $X=2.385 $Y=2.815 $X2=0 $Y2=0
cc_249 N_VPWR_c_341_n N_Y_c_401_n 0.0145938f $X=3.265 $Y=3.33 $X2=0 $Y2=0
cc_250 N_VPWR_c_335_n N_Y_c_401_n 0.0120466f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_251 N_Y_c_393_n N_VGND_M1006_d 0.00419683f $X=4.055 $Y=1.095 $X2=0 $Y2=0
cc_252 N_Y_c_392_n N_VGND_c_480_n 0.0222791f $X=3.485 $Y=0.485 $X2=0 $Y2=0
cc_253 N_Y_c_426_n N_VGND_c_480_n 0.0162446f $X=3.57 $Y=1.01 $X2=0 $Y2=0
cc_254 N_Y_c_393_n N_VGND_c_480_n 0.0281795f $X=4.055 $Y=1.095 $X2=0 $Y2=0
cc_255 N_Y_c_392_n N_VGND_c_481_n 0.0795465f $X=3.485 $Y=0.485 $X2=0 $Y2=0
cc_256 N_Y_c_392_n N_VGND_c_483_n 0.0668803f $X=3.485 $Y=0.485 $X2=0 $Y2=0
cc_257 N_Y_c_392_n A_435_74# 0.0013155f $X=3.485 $Y=0.485 $X2=-0.19 $Y2=-0.245
cc_258 N_Y_c_392_n A_513_74# 0.0103574f $X=3.485 $Y=0.485 $X2=-0.19 $Y2=-0.245
cc_259 N_Y_c_392_n A_627_74# 0.00894458f $X=3.485 $Y=0.485 $X2=-0.19 $Y2=-0.245
cc_260 N_Y_c_426_n A_627_74# 0.00432805f $X=3.57 $Y=1.01 $X2=-0.19 $Y2=-0.245
cc_261 N_Y_c_394_n A_627_74# 9.34031e-19 $X=3.655 $Y=1.095 $X2=-0.19 $Y2=-0.245
