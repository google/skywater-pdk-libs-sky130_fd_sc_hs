* File: sky130_fd_sc_hs__o41ai_2.pex.spice
* Created: Thu Aug 27 21:04:40 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HS__O41AI_2%B1 1 3 4 6 7 9 10 11 12 14 15 17 18 23 24 35
r61 36 37 8.5867 $w=4.21e-07 $l=7.5e-08 $layer=POLY_cond $X=0.945 $Y=1.492
+ $X2=1.02 $Y2=1.492
r62 34 36 24.0428 $w=4.21e-07 $l=2.1e-07 $layer=POLY_cond $X=0.735 $Y=1.492
+ $X2=0.945 $Y2=1.492
r63 34 35 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.735
+ $Y=1.385 $X2=0.735 $Y2=1.385
r64 32 34 27.4774 $w=4.21e-07 $l=2.4e-07 $layer=POLY_cond $X=0.495 $Y=1.492
+ $X2=0.735 $Y2=1.492
r65 31 32 16.0285 $w=4.21e-07 $l=1.4e-07 $layer=POLY_cond $X=0.355 $Y=1.492
+ $X2=0.495 $Y2=1.492
r66 27 31 0.666889 $w=4.6e-07 $l=2.72e-07 $layer=POLY_cond $X=0.355 $Y=1.22
+ $X2=0.355 $Y2=1.492
r67 24 35 0.467207 $w=3.68e-07 $l=1.5e-08 $layer=LI1_cond $X=0.72 $Y=1.365
+ $X2=0.735 $Y2=1.365
r68 24 38 8.25398 $w=3.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.72 $Y=1.365
+ $X2=0.455 $Y2=1.365
r69 23 38 3.26354 $w=3.7e-07 $l=1.83916e-07 $layer=LI1_cond $X=0.29 $Y=1.405
+ $X2=0.455 $Y2=1.365
r70 22 27 11.4858 $w=4.6e-07 $l=9.5e-08 $layer=POLY_cond $X=0.355 $Y=1.125
+ $X2=0.355 $Y2=1.22
r71 21 22 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=0.29
+ $Y=1.125 $X2=0.29 $Y2=1.125
r72 18 22 82.2141 $w=4.6e-07 $l=6.8e-07 $layer=POLY_cond $X=0.355 $Y=0.445
+ $X2=0.355 $Y2=1.125
r73 17 21 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=0.29 $Y=0.445
+ $X2=0.29 $Y2=1.125
r74 17 18 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=0.29
+ $Y=0.445 $X2=0.29 $Y2=0.445
r75 15 23 3.58194 $w=3.3e-07 $l=2.25e-07 $layer=LI1_cond $X=0.29 $Y=1.18
+ $X2=0.29 $Y2=1.405
r76 15 21 1.92074 $w=3.28e-07 $l=5.5e-08 $layer=LI1_cond $X=0.29 $Y=1.18
+ $X2=0.29 $Y2=1.125
r77 12 14 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.45 $Y=1.22 $X2=1.45
+ $Y2=0.74
r78 11 37 29.7157 $w=4.21e-07 $l=2.31482e-07 $layer=POLY_cond $X=1.095 $Y=1.295
+ $X2=1.02 $Y2=1.492
r79 10 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.375 $Y=1.295
+ $X2=1.45 $Y2=1.22
r80 10 11 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=1.375 $Y=1.295
+ $X2=1.095 $Y2=1.295
r81 7 37 27.1176 $w=1.5e-07 $l=2.72e-07 $layer=POLY_cond $X=1.02 $Y=1.22
+ $X2=1.02 $Y2=1.492
r82 7 9 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.02 $Y=1.22 $X2=1.02
+ $Y2=0.74
r83 4 36 27.1176 $w=1.5e-07 $l=2.73e-07 $layer=POLY_cond $X=0.945 $Y=1.765
+ $X2=0.945 $Y2=1.492
r84 4 6 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.945 $Y=1.765
+ $X2=0.945 $Y2=2.4
r85 1 32 27.1176 $w=1.5e-07 $l=2.73e-07 $layer=POLY_cond $X=0.495 $Y=1.765
+ $X2=0.495 $Y2=1.492
r86 1 3 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.495 $Y=1.765
+ $X2=0.495 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_HS__O41AI_2%A4 1 3 6 8 10 13 15 20 23
c57 23 0 1.5097e-19 $X=2.495 $Y=1.515
c58 13 0 1.18304e-19 $X=2.45 $Y=0.74
c59 8 0 1.06955e-19 $X=2.375 $Y=1.765
r60 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.495
+ $Y=1.515 $X2=2.495 $Y2=1.515
r61 20 22 6.2149 $w=3.49e-07 $l=4.5e-08 $layer=POLY_cond $X=2.45 $Y=1.557
+ $X2=2.495 $Y2=1.557
r62 19 20 10.3582 $w=3.49e-07 $l=7.5e-08 $layer=POLY_cond $X=2.375 $Y=1.557
+ $X2=2.45 $Y2=1.557
r63 18 19 58.6963 $w=3.49e-07 $l=4.25e-07 $layer=POLY_cond $X=1.95 $Y=1.557
+ $X2=2.375 $Y2=1.557
r64 17 18 3.45272 $w=3.49e-07 $l=2.5e-08 $layer=POLY_cond $X=1.925 $Y=1.557
+ $X2=1.95 $Y2=1.557
r65 15 23 4.93904 $w=3.48e-07 $l=1.5e-07 $layer=LI1_cond $X=2.58 $Y=1.665
+ $X2=2.58 $Y2=1.515
r66 11 20 22.56 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.45 $Y=1.35 $X2=2.45
+ $Y2=1.557
r67 11 13 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.45 $Y=1.35
+ $X2=2.45 $Y2=0.74
r68 8 19 22.56 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=2.375 $Y=1.765
+ $X2=2.375 $Y2=1.557
r69 8 10 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.375 $Y=1.765
+ $X2=2.375 $Y2=2.4
r70 4 18 22.56 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.95 $Y=1.35 $X2=1.95
+ $Y2=1.557
r71 4 6 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.95 $Y=1.35 $X2=1.95
+ $Y2=0.74
r72 1 17 22.56 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=1.925 $Y=1.765
+ $X2=1.925 $Y2=1.557
r73 1 3 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.925 $Y=1.765
+ $X2=1.925 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_HS__O41AI_2%A3 3 5 7 10 12 14 15 21 22
c48 21 0 9.6541e-21 $X=3.29 $Y=1.515
c49 5 0 1.5097e-19 $X=2.96 $Y=1.765
r50 22 23 3.96164 $w=3.65e-07 $l=3e-08 $layer=POLY_cond $X=3.38 $Y=1.557
+ $X2=3.41 $Y2=1.557
r51 20 22 11.8849 $w=3.65e-07 $l=9e-08 $layer=POLY_cond $X=3.29 $Y=1.557
+ $X2=3.38 $Y2=1.557
r52 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.29
+ $Y=1.515 $X2=3.29 $Y2=1.515
r53 18 20 43.5781 $w=3.65e-07 $l=3.3e-07 $layer=POLY_cond $X=2.96 $Y=1.557
+ $X2=3.29 $Y2=1.557
r54 17 18 1.98082 $w=3.65e-07 $l=1.5e-08 $layer=POLY_cond $X=2.945 $Y=1.557
+ $X2=2.96 $Y2=1.557
r55 15 21 4.55617 $w=4.28e-07 $l=1.7e-07 $layer=LI1_cond $X=3.12 $Y=1.565
+ $X2=3.29 $Y2=1.565
r56 12 23 23.6381 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=3.41 $Y=1.765
+ $X2=3.41 $Y2=1.557
r57 12 14 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.41 $Y=1.765
+ $X2=3.41 $Y2=2.4
r58 8 22 23.6381 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.38 $Y=1.35
+ $X2=3.38 $Y2=1.557
r59 8 10 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=3.38 $Y=1.35 $X2=3.38
+ $Y2=0.74
r60 5 18 23.6381 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=2.96 $Y=1.765
+ $X2=2.96 $Y2=1.557
r61 5 7 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.96 $Y=1.765
+ $X2=2.96 $Y2=2.4
r62 1 17 23.6381 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.945 $Y=1.35
+ $X2=2.945 $Y2=1.557
r63 1 3 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.945 $Y=1.35
+ $X2=2.945 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HS__O41AI_2%A2 3 5 7 10 12 14 16 17 18 19 25 29
c72 29 0 1.5035e-19 $X=4.925 $Y=1.565
c73 25 0 1.0309e-19 $X=5.04 $Y=1.665
c74 12 0 2.60424e-19 $X=4.755 $Y=1.65
r75 25 29 3.73456 $w=4.28e-07 $l=1.15e-07 $layer=LI1_cond $X=5.04 $Y=1.565
+ $X2=4.925 $Y2=1.565
r76 22 29 22.8742 $w=3.28e-07 $l=6.55e-07 $layer=LI1_cond $X=4.27 $Y=1.515
+ $X2=4.925 $Y2=1.515
r77 22 23 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.27
+ $Y=1.515 $X2=4.27 $Y2=1.515
r78 18 23 5.19077 $w=3.75e-07 $l=3.5e-08 $layer=POLY_cond $X=4.305 $Y=1.537
+ $X2=4.27 $Y2=1.537
r79 18 19 6.07033 $w=3.75e-07 $l=9.94987e-08 $layer=POLY_cond $X=4.305 $Y=1.537
+ $X2=4.395 $Y2=1.557
r80 17 23 52.6492 $w=3.75e-07 $l=3.55e-07 $layer=POLY_cond $X=3.915 $Y=1.537
+ $X2=4.27 $Y2=1.537
r81 14 16 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=4.845 $Y=1.765
+ $X2=4.845 $Y2=2.4
r82 13 19 6.07033 $w=1.5e-07 $l=1.30457e-07 $layer=POLY_cond $X=4.485 $Y=1.65
+ $X2=4.395 $Y2=1.557
r83 12 14 26.9307 $w=1.5e-07 $l=1.53542e-07 $layer=POLY_cond $X=4.755 $Y=1.65
+ $X2=4.845 $Y2=1.765
r84 12 13 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=4.755 $Y=1.65
+ $X2=4.485 $Y2=1.65
r85 8 19 19.3751 $w=1.5e-07 $l=2.14369e-07 $layer=POLY_cond $X=4.41 $Y=1.35
+ $X2=4.395 $Y2=1.557
r86 8 10 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=4.41 $Y=1.35 $X2=4.41
+ $Y2=0.74
r87 5 19 19.3751 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=4.395 $Y=1.765
+ $X2=4.395 $Y2=1.557
r88 5 7 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=4.395 $Y=1.765
+ $X2=4.395 $Y2=2.4
r89 1 17 33.9315 $w=3.75e-07 $l=2.21346e-07 $layer=POLY_cond $X=3.84 $Y=1.35
+ $X2=3.915 $Y2=1.537
r90 1 3 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=3.84 $Y=1.35 $X2=3.84
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HS__O41AI_2%A1 1 3 4 5 6 8 9 11 12 14 15 16 21
c53 16 0 1.36826e-19 $X=6 $Y=1.665
c54 6 0 1.0309e-19 $X=5.295 $Y=1.765
r55 23 24 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.855
+ $Y=1.515 $X2=5.855 $Y2=1.515
r56 21 23 9.96617 $w=5.32e-07 $l=1.1e-07 $layer=POLY_cond $X=5.745 $Y=1.475
+ $X2=5.855 $Y2=1.475
r57 20 21 36.6936 $w=5.32e-07 $l=4.05e-07 $layer=POLY_cond $X=5.34 $Y=1.475
+ $X2=5.745 $Y2=1.475
r58 19 20 4.07707 $w=5.32e-07 $l=4.5e-08 $layer=POLY_cond $X=5.295 $Y=1.475
+ $X2=5.34 $Y2=1.475
r59 16 24 3.88615 $w=4.28e-07 $l=1.45e-07 $layer=LI1_cond $X=6 $Y=1.565
+ $X2=5.855 $Y2=1.565
r60 15 24 8.97834 $w=4.28e-07 $l=3.35e-07 $layer=LI1_cond $X=5.52 $Y=1.565
+ $X2=5.855 $Y2=1.565
r61 12 21 32.9824 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=5.745 $Y=1.765
+ $X2=5.745 $Y2=1.475
r62 12 14 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=5.745 $Y=1.765
+ $X2=5.745 $Y2=2.4
r63 9 20 32.9824 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=5.34 $Y=1.185
+ $X2=5.34 $Y2=1.475
r64 9 11 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=5.34 $Y=1.185
+ $X2=5.34 $Y2=0.74
r65 6 19 32.9824 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=5.295 $Y=1.765
+ $X2=5.295 $Y2=1.475
r66 6 8 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=5.295 $Y=1.765
+ $X2=5.295 $Y2=2.4
r67 4 19 35.968 $w=5.32e-07 $l=2.56076e-07 $layer=POLY_cond $X=5.205 $Y=1.26
+ $X2=5.295 $Y2=1.475
r68 4 5 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=5.205 $Y=1.26
+ $X2=4.915 $Y2=1.26
r69 1 5 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.84 $Y=1.185
+ $X2=4.915 $Y2=1.26
r70 1 3 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=4.84 $Y=1.185
+ $X2=4.84 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HS__O41AI_2%VPWR 1 2 3 10 12 18 22 24 26 31 41 42 48 51
r67 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r68 48 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r69 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r70 42 52 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=3.33 $X2=5.52
+ $Y2=3.33
r71 41 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r72 39 51 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.605 $Y=3.33
+ $X2=5.52 $Y2=3.33
r73 39 41 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=5.605 $Y=3.33 $X2=6
+ $Y2=3.33
r74 38 52 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=5.52 $Y2=3.33
r75 37 38 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r76 35 49 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r77 34 37 219.209 $w=1.68e-07 $l=3.36e-06 $layer=LI1_cond $X=1.68 $Y=3.33
+ $X2=5.04 $Y2=3.33
r78 34 35 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r79 32 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.335 $Y=3.33
+ $X2=1.17 $Y2=3.33
r80 32 34 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.335 $Y=3.33
+ $X2=1.68 $Y2=3.33
r81 31 51 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.435 $Y=3.33
+ $X2=5.52 $Y2=3.33
r82 31 37 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=5.435 $Y=3.33
+ $X2=5.04 $Y2=3.33
r83 30 49 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r84 30 46 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r85 29 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r86 27 45 4.75569 $w=1.7e-07 $l=2.18e-07 $layer=LI1_cond $X=0.435 $Y=3.33
+ $X2=0.217 $Y2=3.33
r87 27 29 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.435 $Y=3.33
+ $X2=0.72 $Y2=3.33
r88 26 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.005 $Y=3.33
+ $X2=1.17 $Y2=3.33
r89 26 29 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=1.005 $Y=3.33
+ $X2=0.72 $Y2=3.33
r90 24 38 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=5.04 $Y2=3.33
r91 24 35 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=1.68 $Y2=3.33
r92 20 51 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.52 $Y=3.245
+ $X2=5.52 $Y2=3.33
r93 20 22 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=5.52 $Y=3.245
+ $X2=5.52 $Y2=2.455
r94 16 48 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.17 $Y=3.245
+ $X2=1.17 $Y2=3.33
r95 16 18 35.621 $w=3.28e-07 $l=1.02e-06 $layer=LI1_cond $X=1.17 $Y=3.245
+ $X2=1.17 $Y2=2.225
r96 12 15 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=0.27 $Y=1.985
+ $X2=0.27 $Y2=2.815
r97 10 45 3.01048 $w=3.3e-07 $l=1.08305e-07 $layer=LI1_cond $X=0.27 $Y=3.245
+ $X2=0.217 $Y2=3.33
r98 10 15 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=0.27 $Y=3.245
+ $X2=0.27 $Y2=2.815
r99 3 22 300 $w=1.7e-07 $l=6.85912e-07 $layer=licon1_PDIFF $count=2 $X=5.37
+ $Y=1.84 $X2=5.52 $Y2=2.455
r100 2 18 300 $w=1.7e-07 $l=4.53845e-07 $layer=licon1_PDIFF $count=2 $X=1.02
+ $Y=1.84 $X2=1.17 $Y2=2.225
r101 1 15 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.27 $Y2=2.815
r102 1 12 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.27 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HS__O41AI_2%Y 1 2 3 12 16 17 20 24 26 27 28
r52 28 31 9.49071 $w=3.38e-07 $l=2.8e-07 $layer=LI1_cond $X=1.68 $Y=1.72 $X2=1.4
+ $Y2=1.72
r53 27 31 6.36606 $w=2.55e-07 $l=1.65e-07 $layer=LI1_cond $X=1.235 $Y=1.72
+ $X2=1.4 $Y2=1.72
r54 26 28 12.0329 $w=3.38e-07 $l=3.55e-07 $layer=LI1_cond $X=2.035 $Y=1.72
+ $X2=1.68 $Y2=1.72
r55 22 26 7.42997 $w=3.4e-07 $l=2.14243e-07 $layer=LI1_cond $X=2.135 $Y=1.89
+ $X2=2.035 $Y2=1.72
r56 22 24 5.26818 $w=1.98e-07 $l=9.5e-08 $layer=LI1_cond $X=2.135 $Y=1.89
+ $X2=2.135 $Y2=1.985
r57 18 27 0.432806 $w=3.3e-07 $l=1.7e-07 $layer=LI1_cond $X=1.235 $Y=1.55
+ $X2=1.235 $Y2=1.72
r58 18 20 25.8427 $w=3.28e-07 $l=7.4e-07 $layer=LI1_cond $X=1.235 $Y=1.55
+ $X2=1.235 $Y2=0.81
r59 16 27 6.36606 $w=2.55e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.07 $Y=1.805
+ $X2=1.235 $Y2=1.72
r60 16 17 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=1.07 $Y=1.805
+ $X2=0.805 $Y2=1.805
r61 12 14 54.1497 $w=1.68e-07 $l=8.3e-07 $layer=LI1_cond $X=0.72 $Y=1.985
+ $X2=0.72 $Y2=2.815
r62 10 17 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.72 $Y=1.89
+ $X2=0.805 $Y2=1.805
r63 10 12 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=0.72 $Y=1.89
+ $X2=0.72 $Y2=1.985
r64 3 24 300 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=2 $X=2 $Y=1.84
+ $X2=2.15 $Y2=1.985
r65 2 14 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=0.57
+ $Y=1.84 $X2=0.72 $Y2=2.815
r66 2 12 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=0.57
+ $Y=1.84 $X2=0.72 $Y2=1.985
r67 1 20 182 $w=1.7e-07 $l=5.05173e-07 $layer=licon1_NDIFF $count=1 $X=1.095
+ $Y=0.37 $X2=1.235 $Y2=0.81
.ends

.subckt PM_SKY130_FD_SC_HS__O41AI_2%A_314_368# 1 2 3 12 14 15 16 19 20 27
r47 21 25 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.765 $Y=2.035
+ $X2=2.6 $Y2=2.035
r48 20 27 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.47 $Y=2.035
+ $X2=3.635 $Y2=2.035
r49 20 21 45.9947 $w=1.68e-07 $l=7.05e-07 $layer=LI1_cond $X=3.47 $Y=2.035
+ $X2=2.765 $Y2=2.035
r50 17 19 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=2.6 $Y=2.905 $X2=2.6
+ $Y2=2.815
r51 16 25 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.6 $Y=2.12 $X2=2.6
+ $Y2=2.035
r52 16 19 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=2.6 $Y=2.12 $X2=2.6
+ $Y2=2.815
r53 14 17 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.435 $Y=2.99
+ $X2=2.6 $Y2=2.905
r54 14 15 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=2.435 $Y=2.99
+ $X2=1.865 $Y2=2.99
r55 10 15 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.7 $Y=2.905
+ $X2=1.865 $Y2=2.99
r56 10 12 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=1.7 $Y=2.905 $X2=1.7
+ $Y2=2.225
r57 3 27 300 $w=1.7e-07 $l=3.4187e-07 $layer=licon1_PDIFF $count=2 $X=3.485
+ $Y=1.84 $X2=3.635 $Y2=2.115
r58 2 25 400 $w=1.7e-07 $l=3.4187e-07 $layer=licon1_PDIFF $count=1 $X=2.45
+ $Y=1.84 $X2=2.6 $Y2=2.115
r59 2 19 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=2.45
+ $Y=1.84 $X2=2.6 $Y2=2.815
r60 1 12 300 $w=1.7e-07 $l=4.45281e-07 $layer=licon1_PDIFF $count=2 $X=1.57
+ $Y=1.84 $X2=1.7 $Y2=2.225
.ends

.subckt PM_SKY130_FD_SC_HS__O41AI_2%A_607_368# 1 2 9 11 12 15
c25 12 0 9.73009e-20 $X=3.27 $Y=2.99
r26 13 15 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=4.62 $Y=2.905
+ $X2=4.62 $Y2=2.455
r27 11 13 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.535 $Y=2.99
+ $X2=4.62 $Y2=2.905
r28 11 12 82.5294 $w=1.68e-07 $l=1.265e-06 $layer=LI1_cond $X=4.535 $Y=2.99
+ $X2=3.27 $Y2=2.99
r29 7 12 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=3.145 $Y=2.905
+ $X2=3.27 $Y2=2.99
r30 7 9 20.744 $w=2.48e-07 $l=4.5e-07 $layer=LI1_cond $X=3.145 $Y=2.905
+ $X2=3.145 $Y2=2.455
r31 2 15 300 $w=1.7e-07 $l=6.85912e-07 $layer=licon1_PDIFF $count=2 $X=4.47
+ $Y=1.84 $X2=4.62 $Y2=2.455
r32 1 9 300 $w=1.7e-07 $l=6.85912e-07 $layer=licon1_PDIFF $count=2 $X=3.035
+ $Y=1.84 $X2=3.185 $Y2=2.455
.ends

.subckt PM_SKY130_FD_SC_HS__O41AI_2%A_807_368# 1 2 3 12 16 18 20 22 25 27
r47 20 29 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.97 $Y=2.12 $X2=5.97
+ $Y2=2.035
r48 20 22 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=5.97 $Y=2.12
+ $X2=5.97 $Y2=2.815
r49 19 27 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.235 $Y=2.035
+ $X2=5.07 $Y2=2.035
r50 18 29 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.805 $Y=2.035
+ $X2=5.97 $Y2=2.035
r51 18 19 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=5.805 $Y=2.035
+ $X2=5.235 $Y2=2.035
r52 14 27 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.07 $Y=2.12 $X2=5.07
+ $Y2=2.035
r53 14 16 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=5.07 $Y=2.12
+ $X2=5.07 $Y2=2.815
r54 13 25 4.77065 $w=1.7e-07 $l=1.88348e-07 $layer=LI1_cond $X=4.335 $Y=2.035
+ $X2=4.17 $Y2=1.985
r55 12 27 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.905 $Y=2.035
+ $X2=5.07 $Y2=2.035
r56 12 13 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=4.905 $Y=2.035
+ $X2=4.335 $Y2=2.035
r57 3 29 400 $w=1.7e-07 $l=3.4187e-07 $layer=licon1_PDIFF $count=1 $X=5.82
+ $Y=1.84 $X2=5.97 $Y2=2.115
r58 3 22 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=5.82
+ $Y=1.84 $X2=5.97 $Y2=2.815
r59 2 27 400 $w=1.7e-07 $l=3.4187e-07 $layer=licon1_PDIFF $count=1 $X=4.92
+ $Y=1.84 $X2=5.07 $Y2=2.115
r60 2 16 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=4.92
+ $Y=1.84 $X2=5.07 $Y2=2.815
r61 1 25 300 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=2 $X=4.035
+ $Y=1.84 $X2=4.17 $Y2=2.015
.ends

.subckt PM_SKY130_FD_SC_HS__O41AI_2%A_132_74# 1 2 3 4 5 6 21 23 24 28 29 30 33
+ 35 39 41 45 47 51 53 54 55
c98 47 0 1.23598e-19 $X=5.46 $Y=1.095
c99 23 0 1.18304e-19 $X=1.57 $Y=0.34
r100 49 51 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=5.625 $Y=1.01
+ $X2=5.625 $Y2=0.515
r101 48 55 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.79 $Y=1.095
+ $X2=4.625 $Y2=1.095
r102 47 49 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=5.46 $Y=1.095
+ $X2=5.625 $Y2=1.01
r103 47 48 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.46 $Y=1.095
+ $X2=4.79 $Y2=1.095
r104 43 55 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.625 $Y=1.01
+ $X2=4.625 $Y2=1.095
r105 43 45 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=4.625 $Y=1.01
+ $X2=4.625 $Y2=0.515
r106 42 54 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=3.79 $Y=1.095
+ $X2=3.65 $Y2=1.095
r107 41 55 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.46 $Y=1.095
+ $X2=4.625 $Y2=1.095
r108 41 42 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.46 $Y=1.095
+ $X2=3.79 $Y2=1.095
r109 37 54 0.375625 $w=2.8e-07 $l=8.5e-08 $layer=LI1_cond $X=3.65 $Y=1.01
+ $X2=3.65 $Y2=1.095
r110 37 39 20.3735 $w=2.78e-07 $l=4.95e-07 $layer=LI1_cond $X=3.65 $Y=1.01
+ $X2=3.65 $Y2=0.515
r111 36 53 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.83 $Y=1.095
+ $X2=2.705 $Y2=1.095
r112 35 54 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=3.51 $Y=1.095
+ $X2=3.65 $Y2=1.095
r113 35 36 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=3.51 $Y=1.095
+ $X2=2.83 $Y2=1.095
r114 31 53 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.705 $Y=1.01
+ $X2=2.705 $Y2=1.095
r115 31 33 22.8184 $w=2.48e-07 $l=4.95e-07 $layer=LI1_cond $X=2.705 $Y=1.01
+ $X2=2.705 $Y2=0.515
r116 29 53 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.58 $Y=1.095
+ $X2=2.705 $Y2=1.095
r117 29 30 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=2.58 $Y=1.095
+ $X2=1.9 $Y2=1.095
r118 26 30 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.735 $Y=1.01
+ $X2=1.9 $Y2=1.095
r119 26 28 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=1.735 $Y=1.01
+ $X2=1.735 $Y2=0.515
r120 25 28 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=1.735 $Y=0.425
+ $X2=1.735 $Y2=0.515
r121 23 25 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.57 $Y=0.34
+ $X2=1.735 $Y2=0.425
r122 23 24 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.57 $Y=0.34
+ $X2=0.89 $Y2=0.34
r123 19 24 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.765 $Y=0.425
+ $X2=0.89 $Y2=0.34
r124 19 21 3.68782 $w=2.48e-07 $l=8e-08 $layer=LI1_cond $X=0.765 $Y=0.425
+ $X2=0.765 $Y2=0.505
r125 6 51 91 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=2 $X=5.415
+ $Y=0.37 $X2=5.625 $Y2=0.515
r126 5 45 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=4.485
+ $Y=0.37 $X2=4.625 $Y2=0.515
r127 4 39 91 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_NDIFF $count=2 $X=3.455
+ $Y=0.37 $X2=3.61 $Y2=0.515
r128 3 33 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.525
+ $Y=0.37 $X2=2.665 $Y2=0.515
r129 2 28 91 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=2 $X=1.525
+ $Y=0.37 $X2=1.735 $Y2=0.515
r130 1 21 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=0.66
+ $Y=0.37 $X2=0.805 $Y2=0.505
.ends

.subckt PM_SKY130_FD_SC_HS__O41AI_2%VGND 1 2 3 4 15 19 23 25 29 31 33 41 46 53
+ 54 57 60 63 66
r77 66 67 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r78 64 67 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=5.04
+ $Y2=0
r79 63 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r80 57 58 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r81 54 67 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6 $Y=0 $X2=5.04
+ $Y2=0
r82 53 54 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6 $Y=0 $X2=6 $Y2=0
r83 51 66 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.29 $Y=0 $X2=5.125
+ $Y2=0
r84 51 53 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=5.29 $Y=0 $X2=6
+ $Y2=0
r85 50 64 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.08
+ $Y2=0
r86 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r87 47 60 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.33 $Y=0 $X2=3.165
+ $Y2=0
r88 47 49 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=3.33 $Y=0 $X2=3.6
+ $Y2=0
r89 46 63 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.96 $Y=0 $X2=4.125
+ $Y2=0
r90 46 49 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=3.96 $Y=0 $X2=3.6
+ $Y2=0
r91 45 58 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=2.16
+ $Y2=0
r92 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r93 42 57 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.4 $Y=0 $X2=2.235
+ $Y2=0
r94 42 44 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=2.4 $Y=0 $X2=2.64
+ $Y2=0
r95 41 60 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3 $Y=0 $X2=3.165
+ $Y2=0
r96 41 44 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=3 $Y=0 $X2=2.64
+ $Y2=0
r97 40 58 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r98 39 40 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r99 36 40 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=0.24 $Y=0 $X2=1.68
+ $Y2=0
r100 35 39 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=0.24 $Y=0 $X2=1.68
+ $Y2=0
r101 35 36 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r102 33 57 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.07 $Y=0 $X2=2.235
+ $Y2=0
r103 33 39 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=2.07 $Y=0 $X2=1.68
+ $Y2=0
r104 31 50 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=3.6
+ $Y2=0
r105 31 45 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=2.64
+ $Y2=0
r106 31 60 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r107 27 66 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.125 $Y=0.085
+ $X2=5.125 $Y2=0
r108 27 29 19.0328 $w=3.28e-07 $l=5.45e-07 $layer=LI1_cond $X=5.125 $Y=0.085
+ $X2=5.125 $Y2=0.63
r109 26 63 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.29 $Y=0 $X2=4.125
+ $Y2=0
r110 25 66 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.96 $Y=0 $X2=5.125
+ $Y2=0
r111 25 26 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.96 $Y=0 $X2=4.29
+ $Y2=0
r112 21 63 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.125 $Y=0.085
+ $X2=4.125 $Y2=0
r113 21 23 19.0328 $w=3.28e-07 $l=5.45e-07 $layer=LI1_cond $X=4.125 $Y=0.085
+ $X2=4.125 $Y2=0.63
r114 17 60 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.165 $Y=0.085
+ $X2=3.165 $Y2=0
r115 17 19 19.0328 $w=3.28e-07 $l=5.45e-07 $layer=LI1_cond $X=3.165 $Y=0.085
+ $X2=3.165 $Y2=0.63
r116 13 57 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.235 $Y=0.085
+ $X2=2.235 $Y2=0
r117 13 15 19.0328 $w=3.28e-07 $l=5.45e-07 $layer=LI1_cond $X=2.235 $Y=0.085
+ $X2=2.235 $Y2=0.63
r118 4 29 182 $w=1.7e-07 $l=3.49571e-07 $layer=licon1_NDIFF $count=1 $X=4.915
+ $Y=0.37 $X2=5.125 $Y2=0.63
r119 3 23 182 $w=1.7e-07 $l=3.49571e-07 $layer=licon1_NDIFF $count=1 $X=3.915
+ $Y=0.37 $X2=4.125 $Y2=0.63
r120 2 19 182 $w=1.7e-07 $l=3.245e-07 $layer=licon1_NDIFF $count=1 $X=3.02
+ $Y=0.37 $X2=3.165 $Y2=0.63
r121 1 15 182 $w=1.7e-07 $l=3.49571e-07 $layer=licon1_NDIFF $count=1 $X=2.025
+ $Y=0.37 $X2=2.235 $Y2=0.63
.ends

