* File: sky130_fd_sc_hs__a22o_1.spice
* Created: Thu Aug 27 20:26:51 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hs__a22o_1.pex.spice"
.subckt sky130_fd_sc_hs__a22o_1  VNB VPB A2 B2 B1 A1 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A1	A1
* B1	B1
* B2	B2
* A2	A2
* VPB	VPB
* VNB	VNB
MM1002 N_VGND_M1002_d N_A2_M1002_g N_A_52_123#_M1002_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.12325 AS=0.1696 PD=1.185 PS=1.81 NRD=3.744 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75001 A=0.096 P=1.58 MULT=1
MM1004 A_230_79# N_B2_M1004_g N_VGND_M1002_d VNB NLOWVT L=0.15 W=0.64 AD=0.0672
+ AS=0.12325 PD=0.85 PS=1.185 NRD=9.372 NRS=4.68 M=1 R=4.26667 SA=75000.5
+ SB=75001 A=0.096 P=1.58 MULT=1
MM1000 N_A_222_392#_M1000_d N_B1_M1000_g A_230_79# VNB NLOWVT L=0.15 W=0.64
+ AD=0.0896 AS=0.0672 PD=0.92 PS=0.85 NRD=0 NRS=9.372 M=1 R=4.26667 SA=75000.9
+ SB=75000.6 A=0.096 P=1.58 MULT=1
MM1005 N_A_52_123#_M1005_d N_A1_M1005_g N_A_222_392#_M1000_d VNB NLOWVT L=0.15
+ W=0.64 AD=0.1824 AS=0.0896 PD=1.85 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75001.3 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1008 N_X_M1008_d N_A_222_392#_M1008_g N_VGND_M1008_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1961 AS=0.1961 PD=2.01 PS=2.01 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1009 N_A_132_392#_M1009_d N_A2_M1009_g N_VPWR_M1009_s VPB PSHORT L=0.15 W=1
+ AD=0.15 AS=0.275 PD=1.3 PS=2.55 NRD=1.9503 NRS=1.9503 M=1 R=6.66667 SA=75000.2
+ SB=75002.4 A=0.15 P=2.3 MULT=1
MM1003 N_A_222_392#_M1003_d N_B2_M1003_g N_A_132_392#_M1009_d VPB PSHORT L=0.15
+ W=1 AD=0.165 AS=0.15 PD=1.33 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=6.66667
+ SA=75000.6 SB=75001.9 A=0.15 P=2.3 MULT=1
MM1006 N_A_132_392#_M1006_d N_B1_M1006_g N_A_222_392#_M1003_d VPB PSHORT L=0.15
+ W=1 AD=0.195 AS=0.165 PD=1.39 PS=1.33 NRD=12.7853 NRS=7.8603 M=1 R=6.66667
+ SA=75001.1 SB=75001.5 A=0.15 P=2.3 MULT=1
MM1001 N_VPWR_M1001_d N_A1_M1001_g N_A_132_392#_M1006_d VPB PSHORT L=0.15 W=1
+ AD=0.289151 AS=0.195 PD=1.60377 PS=1.39 NRD=30.0228 NRS=8.8453 M=1 R=6.66667
+ SA=75001.7 SB=75000.9 A=0.15 P=2.3 MULT=1
MM1007 N_X_M1007_d N_A_222_392#_M1007_g N_VPWR_M1001_d VPB PSHORT L=0.15 W=1.12
+ AD=0.308 AS=0.323849 PD=2.79 PS=1.79623 NRD=1.7533 NRS=25.9252 M=1 R=7.46667
+ SA=75002.2 SB=75000.2 A=0.168 P=2.54 MULT=1
DX10_noxref VNB VPB NWDIODE A=6.9564 P=11.2
*
.include "sky130_fd_sc_hs__a22o_1.pxi.spice"
*
.ends
*
*
