* File: sky130_fd_sc_hs__a22oi_2.pex.spice
* Created: Tue Sep  1 19:51:29 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HS__A22OI_2%A1 3 5 7 10 12 14 15 16 17 18 21 22 24 25 35
c90 22 0 2.00043e-19 $X=2.045 $Y=1.515
c91 15 0 5.96145e-20 $X=0.795 $Y=1.78
c92 10 0 1.09905e-19 $X=2.025 $Y=0.74
r93 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.605
+ $Y=1.515 $X2=0.605 $Y2=1.515
r94 25 35 2.59474 $w=3.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.795 $Y=1.605
+ $X2=0.71 $Y2=1.605
r95 25 35 1.25122 $w=3.48e-07 $l=3.8e-08 $layer=LI1_cond $X=0.672 $Y=1.605
+ $X2=0.71 $Y2=1.605
r96 25 31 2.20611 $w=3.48e-07 $l=6.7e-08 $layer=LI1_cond $X=0.672 $Y=1.605
+ $X2=0.605 $Y2=1.605
r97 24 31 12.0183 $w=3.48e-07 $l=3.65e-07 $layer=LI1_cond $X=0.24 $Y=1.605
+ $X2=0.605 $Y2=1.605
r98 22 34 39.8291 $w=3.57e-07 $l=2.95e-07 $layer=POLY_cond $X=2.045 $Y=1.557
+ $X2=2.34 $Y2=1.557
r99 22 32 2.70028 $w=3.57e-07 $l=2e-08 $layer=POLY_cond $X=2.045 $Y=1.557
+ $X2=2.025 $Y2=1.557
r100 21 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.045
+ $Y=1.515 $X2=2.045 $Y2=1.515
r101 19 21 15.1913 $w=3.28e-07 $l=4.35e-07 $layer=LI1_cond $X=2.045 $Y=1.95
+ $X2=2.045 $Y2=1.515
r102 17 19 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.88 $Y=2.035
+ $X2=2.045 $Y2=1.95
r103 17 18 65.2406 $w=1.68e-07 $l=1e-06 $layer=LI1_cond $X=1.88 $Y=2.035
+ $X2=0.88 $Y2=2.035
r104 16 18 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.795 $Y=1.95
+ $X2=0.88 $Y2=2.035
r105 15 25 5.34211 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=0.795 $Y=1.78
+ $X2=0.795 $Y2=1.605
r106 15 16 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=0.795 $Y=1.78
+ $X2=0.795 $Y2=1.95
r107 12 34 23.1043 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=2.34 $Y=1.765
+ $X2=2.34 $Y2=1.557
r108 12 14 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.34 $Y=1.765
+ $X2=2.34 $Y2=2.4
r109 8 32 23.1043 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.025 $Y=1.35
+ $X2=2.025 $Y2=1.557
r110 8 10 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.025 $Y=1.35
+ $X2=2.025 $Y2=0.74
r111 5 30 52.2586 $w=2.99e-07 $l=2.85044e-07 $layer=POLY_cond $X=0.68 $Y=1.765
+ $X2=0.605 $Y2=1.515
r112 5 7 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.68 $Y=1.765
+ $X2=0.68 $Y2=2.4
r113 1 30 38.5562 $w=2.99e-07 $l=1.92678e-07 $layer=POLY_cond $X=0.665 $Y=1.35
+ $X2=0.605 $Y2=1.515
r114 1 3 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=0.665 $Y=1.35
+ $X2=0.665 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HS__A22OI_2%A2 3 5 7 8 10 13 15 21 22
c51 5 0 5.96145e-20 $X=1.13 $Y=1.765
r52 22 23 1.91777 $w=3.77e-07 $l=1.5e-08 $layer=POLY_cond $X=1.58 $Y=1.557
+ $X2=1.595 $Y2=1.557
r53 20 22 46.6658 $w=3.77e-07 $l=3.65e-07 $layer=POLY_cond $X=1.215 $Y=1.557
+ $X2=1.58 $Y2=1.557
r54 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.215
+ $Y=1.515 $X2=1.215 $Y2=1.515
r55 18 20 10.8674 $w=3.77e-07 $l=8.5e-08 $layer=POLY_cond $X=1.13 $Y=1.557
+ $X2=1.215 $Y2=1.557
r56 17 18 4.4748 $w=3.77e-07 $l=3.5e-08 $layer=POLY_cond $X=1.095 $Y=1.557
+ $X2=1.13 $Y2=1.557
r57 15 21 4.67207 $w=3.68e-07 $l=1.5e-07 $layer=LI1_cond $X=1.235 $Y=1.665
+ $X2=1.235 $Y2=1.515
r58 11 23 24.4204 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.595 $Y=1.35
+ $X2=1.595 $Y2=1.557
r59 11 13 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.595 $Y=1.35
+ $X2=1.595 $Y2=0.74
r60 8 22 24.4204 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=1.58 $Y=1.765
+ $X2=1.58 $Y2=1.557
r61 8 10 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.58 $Y=1.765
+ $X2=1.58 $Y2=2.4
r62 5 18 24.4204 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=1.13 $Y=1.765
+ $X2=1.13 $Y2=1.557
r63 5 7 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.13 $Y=1.765
+ $X2=1.13 $Y2=2.4
r64 1 17 24.4204 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.095 $Y=1.35
+ $X2=1.095 $Y2=1.557
r65 1 3 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.095 $Y=1.35
+ $X2=1.095 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HS__A22OI_2%B1 1 3 4 6 9 11 13 14 20 30
c75 30 0 2.81767e-19 $X=3.235 $Y=1.32
r76 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.805
+ $Y=1.385 $X2=2.805 $Y2=1.385
r77 20 30 7.98002 $w=4.58e-07 $l=1.15e-07 $layer=LI1_cond $X=3.12 $Y=1.32
+ $X2=3.235 $Y2=1.32
r78 20 24 8.19054 $w=4.58e-07 $l=3.15e-07 $layer=LI1_cond $X=3.12 $Y=1.32
+ $X2=2.805 $Y2=1.32
r79 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.205
+ $Y=1.465 $X2=4.205 $Y2=1.465
r80 14 18 10.1086 $w=3.5e-07 $l=3.89076e-07 $layer=LI1_cond $X=3.905 $Y=1.175
+ $X2=4.137 $Y2=1.465
r81 14 30 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.905 $Y=1.175
+ $X2=3.235 $Y2=1.175
r82 11 19 61.4066 $w=2.86e-07 $l=3.17017e-07 $layer=POLY_cond $X=4.17 $Y=1.765
+ $X2=4.205 $Y2=1.465
r83 11 13 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=4.17 $Y=1.765
+ $X2=4.17 $Y2=2.4
r84 7 19 38.6549 $w=2.86e-07 $l=2.05122e-07 $layer=POLY_cond $X=4.115 $Y=1.3
+ $X2=4.205 $Y2=1.465
r85 7 9 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=4.115 $Y=1.3 $X2=4.115
+ $Y2=0.74
r86 4 23 77.2841 $w=2.7e-07 $l=3.87427e-07 $layer=POLY_cond $X=2.79 $Y=1.765
+ $X2=2.805 $Y2=1.385
r87 4 6 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.79 $Y=1.765
+ $X2=2.79 $Y2=2.4
r88 1 23 38.9026 $w=2.7e-07 $l=2.05122e-07 $layer=POLY_cond $X=2.715 $Y=1.22
+ $X2=2.805 $Y2=1.385
r89 1 3 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=2.715 $Y=1.22 $X2=2.715
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HS__A22OI_2%B2 3 5 7 10 12 14 15 21 22
r54 22 23 4.46296 $w=3.78e-07 $l=3.5e-08 $layer=POLY_cond $X=3.685 $Y=1.557
+ $X2=3.72 $Y2=1.557
r55 20 22 14.664 $w=3.78e-07 $l=1.15e-07 $layer=POLY_cond $X=3.57 $Y=1.557
+ $X2=3.685 $Y2=1.557
r56 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.57
+ $Y=1.515 $X2=3.57 $Y2=1.515
r57 18 20 38.254 $w=3.78e-07 $l=3e-07 $layer=POLY_cond $X=3.27 $Y=1.557 $X2=3.57
+ $Y2=1.557
r58 17 18 1.9127 $w=3.78e-07 $l=1.5e-08 $layer=POLY_cond $X=3.255 $Y=1.557
+ $X2=3.27 $Y2=1.557
r59 15 21 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=3.57 $Y=1.665
+ $X2=3.57 $Y2=1.515
r60 12 23 24.4846 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=3.72 $Y=1.765
+ $X2=3.72 $Y2=1.557
r61 12 14 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.72 $Y=1.765
+ $X2=3.72 $Y2=2.4
r62 8 22 24.4846 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.685 $Y=1.35
+ $X2=3.685 $Y2=1.557
r63 8 10 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=3.685 $Y=1.35
+ $X2=3.685 $Y2=0.74
r64 5 18 24.4846 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=3.27 $Y=1.765
+ $X2=3.27 $Y2=1.557
r65 5 7 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.27 $Y=1.765
+ $X2=3.27 $Y2=2.4
r66 1 17 24.4846 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.255 $Y=1.35
+ $X2=3.255 $Y2=1.557
r67 1 3 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=3.255 $Y=1.35
+ $X2=3.255 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HS__A22OI_2%A_66_368# 1 2 3 4 5 18 22 24 28 33 34 35 38
+ 40 44 46 48 50 53
r84 50 52 7.85757 $w=3.28e-07 $l=2.25e-07 $layer=LI1_cond $X=2.565 $Y=2.15
+ $X2=2.565 $Y2=2.375
r85 42 44 18.1597 $w=3.28e-07 $l=5.2e-07 $layer=LI1_cond $X=4.395 $Y=2.905
+ $X2=4.395 $Y2=2.385
r86 41 53 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.66 $Y=2.99
+ $X2=3.495 $Y2=2.99
r87 40 42 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.23 $Y=2.99
+ $X2=4.395 $Y2=2.905
r88 40 41 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=4.23 $Y=2.99
+ $X2=3.66 $Y2=2.99
r89 36 53 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.495 $Y=2.905
+ $X2=3.495 $Y2=2.99
r90 36 38 18.1597 $w=3.28e-07 $l=5.2e-07 $layer=LI1_cond $X=3.495 $Y=2.905
+ $X2=3.495 $Y2=2.385
r91 34 53 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.33 $Y=2.99
+ $X2=3.495 $Y2=2.99
r92 34 35 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=3.33 $Y=2.99 $X2=2.73
+ $Y2=2.99
r93 31 35 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.565 $Y=2.905
+ $X2=2.73 $Y2=2.99
r94 31 33 2.61919 $w=3.28e-07 $l=7.5e-08 $layer=LI1_cond $X=2.565 $Y=2.905
+ $X2=2.565 $Y2=2.83
r95 30 52 2.96841 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=2.565 $Y=2.46
+ $X2=2.565 $Y2=2.375
r96 30 33 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=2.565 $Y=2.46
+ $X2=2.565 $Y2=2.83
r97 29 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.52 $Y=2.375
+ $X2=1.355 $Y2=2.375
r98 28 52 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.4 $Y=2.375
+ $X2=2.565 $Y2=2.375
r99 28 29 57.4118 $w=1.68e-07 $l=8.8e-07 $layer=LI1_cond $X=2.4 $Y=2.375
+ $X2=1.52 $Y2=2.375
r100 25 46 2.76166 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.54 $Y=2.375
+ $X2=0.415 $Y2=2.375
r101 24 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.19 $Y=2.375
+ $X2=1.355 $Y2=2.375
r102 24 25 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=1.19 $Y=2.375
+ $X2=0.54 $Y2=2.375
r103 20 46 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.415 $Y=2.46
+ $X2=0.415 $Y2=2.375
r104 20 22 0.230489 $w=2.48e-07 $l=5e-09 $layer=LI1_cond $X=0.415 $Y=2.46
+ $X2=0.415 $Y2=2.465
r105 16 46 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.415 $Y=2.29
+ $X2=0.415 $Y2=2.375
r106 16 18 8.0671 $w=2.48e-07 $l=1.75e-07 $layer=LI1_cond $X=0.415 $Y=2.29
+ $X2=0.415 $Y2=2.115
r107 5 44 300 $w=1.7e-07 $l=6.15447e-07 $layer=licon1_PDIFF $count=2 $X=4.245
+ $Y=1.84 $X2=4.395 $Y2=2.385
r108 4 38 300 $w=1.7e-07 $l=6.15447e-07 $layer=licon1_PDIFF $count=2 $X=3.345
+ $Y=1.84 $X2=3.495 $Y2=2.385
r109 3 50 400 $w=1.7e-07 $l=3.77624e-07 $layer=licon1_PDIFF $count=1 $X=2.415
+ $Y=1.84 $X2=2.565 $Y2=2.15
r110 3 33 400 $w=1.7e-07 $l=1.06236e-06 $layer=licon1_PDIFF $count=1 $X=2.415
+ $Y=1.84 $X2=2.565 $Y2=2.83
r111 2 48 300 $w=1.7e-07 $l=6.05372e-07 $layer=licon1_PDIFF $count=2 $X=1.205
+ $Y=1.84 $X2=1.355 $Y2=2.375
r112 1 22 300 $w=1.7e-07 $l=6.84653e-07 $layer=licon1_PDIFF $count=2 $X=0.33
+ $Y=1.84 $X2=0.455 $Y2=2.465
r113 1 18 600 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_PDIFF $count=1 $X=0.33
+ $Y=1.84 $X2=0.455 $Y2=2.115
.ends

.subckt PM_SKY130_FD_SC_HS__A22OI_2%VPWR 1 2 9 13 16 17 18 24 30 31 34
r54 34 35 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r55 30 31 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r56 28 34 11.8214 $w=1.7e-07 $l=2.7e-07 $layer=LI1_cond $X=2.23 $Y=3.33 $X2=1.96
+ $Y2=3.33
r57 28 30 152.011 $w=1.68e-07 $l=2.33e-06 $layer=LI1_cond $X=2.23 $Y=3.33
+ $X2=4.56 $Y2=3.33
r58 27 35 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r59 26 27 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r60 24 34 11.8214 $w=1.7e-07 $l=2.7e-07 $layer=LI1_cond $X=1.69 $Y=3.33 $X2=1.96
+ $Y2=3.33
r61 24 26 0.652406 $w=1.68e-07 $l=1e-08 $layer=LI1_cond $X=1.69 $Y=3.33 $X2=1.68
+ $Y2=3.33
r62 22 27 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.68 $Y2=3.33
r63 21 22 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r64 18 31 0.602067 $w=4.9e-07 $l=2.16e-06 $layer=MET1_cond $X=2.4 $Y=3.33
+ $X2=4.56 $Y2=3.33
r65 18 35 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.4 $Y=3.33
+ $X2=2.16 $Y2=3.33
r66 16 21 1.30481 $w=1.68e-07 $l=2e-08 $layer=LI1_cond $X=0.74 $Y=3.33 $X2=0.72
+ $Y2=3.33
r67 16 17 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.74 $Y=3.33
+ $X2=0.865 $Y2=3.33
r68 15 26 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=0.99 $Y=3.33 $X2=1.68
+ $Y2=3.33
r69 15 17 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.99 $Y=3.33
+ $X2=0.865 $Y2=3.33
r70 11 34 2.26835 $w=5.4e-07 $l=8.5e-08 $layer=LI1_cond $X=1.96 $Y=3.245
+ $X2=1.96 $Y2=3.33
r71 11 13 9.74582 $w=5.38e-07 $l=4.4e-07 $layer=LI1_cond $X=1.96 $Y=3.245
+ $X2=1.96 $Y2=2.805
r72 7 17 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.865 $Y=3.245
+ $X2=0.865 $Y2=3.33
r73 7 9 20.283 $w=2.48e-07 $l=4.4e-07 $layer=LI1_cond $X=0.865 $Y=3.245
+ $X2=0.865 $Y2=2.805
r74 2 13 600 $w=1.7e-07 $l=1.10705e-06 $layer=licon1_PDIFF $count=1 $X=1.655
+ $Y=1.84 $X2=1.96 $Y2=2.805
r75 1 9 600 $w=1.7e-07 $l=1.03729e-06 $layer=licon1_PDIFF $count=1 $X=0.755
+ $Y=1.84 $X2=0.905 $Y2=2.805
.ends

.subckt PM_SKY130_FD_SC_HS__A22OI_2%Y 1 2 3 4 5 18 20 21 24 27 28 29 32 34 38 40
+ 44 47 48 54 55 56
c102 48 0 2.81812e-20 $X=3.03 $Y=1.805
r103 63 64 7.70264 $w=5.08e-07 $l=8.5e-08 $layer=LI1_cond $X=2.295 $Y=1.175
+ $X2=2.295 $Y2=1.26
r104 62 63 4.92503 $w=5.08e-07 $l=2.1e-07 $layer=LI1_cond $X=2.295 $Y=0.965
+ $X2=2.295 $Y2=1.175
r105 56 62 0.938101 $w=5.08e-07 $l=4e-08 $layer=LI1_cond $X=2.295 $Y=0.925
+ $X2=2.295 $Y2=0.965
r106 56 59 3.23794 $w=5.08e-07 $l=1.15e-07 $layer=LI1_cond $X=2.295 $Y=0.925
+ $X2=2.295 $Y2=0.81
r107 51 52 2.77273 $w=1.98e-07 $l=5e-08 $layer=LI1_cond $X=3.03 $Y=1.985
+ $X2=3.03 $Y2=2.035
r108 48 51 9.98182 $w=1.98e-07 $l=1.8e-07 $layer=LI1_cond $X=3.03 $Y=1.805
+ $X2=3.03 $Y2=1.985
r109 47 55 53.4973 $w=1.68e-07 $l=8.2e-07 $layer=LI1_cond $X=4.625 $Y=1.95
+ $X2=4.625 $Y2=1.13
r110 42 55 11.032 $w=4.63e-07 $l=2.32e-07 $layer=LI1_cond $X=4.477 $Y=0.898
+ $X2=4.477 $Y2=1.13
r111 42 44 9.85157 $w=4.63e-07 $l=3.83e-07 $layer=LI1_cond $X=4.477 $Y=0.898
+ $X2=4.477 $Y2=0.515
r112 41 54 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.03 $Y=2.035
+ $X2=3.945 $Y2=2.035
r113 40 47 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.54 $Y=2.035
+ $X2=4.625 $Y2=1.95
r114 40 41 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=4.54 $Y=2.035
+ $X2=4.03 $Y2=2.035
r115 36 54 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.945 $Y=2.12
+ $X2=3.945 $Y2=2.035
r116 36 38 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=3.945 $Y=2.12
+ $X2=3.945 $Y2=2.57
r117 35 52 1.68994 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=3.13 $Y=2.035 $X2=3.03
+ $Y2=2.035
r118 34 54 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.86 $Y=2.035
+ $X2=3.945 $Y2=2.035
r119 34 35 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=3.86 $Y=2.035
+ $X2=3.13 $Y2=2.035
r120 30 52 4.71364 $w=1.98e-07 $l=8.5e-08 $layer=LI1_cond $X=3.03 $Y=2.12
+ $X2=3.03 $Y2=2.035
r121 30 32 24.9545 $w=1.98e-07 $l=4.5e-07 $layer=LI1_cond $X=3.03 $Y=2.12
+ $X2=3.03 $Y2=2.57
r122 28 48 1.68994 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=2.93 $Y=1.805 $X2=3.03
+ $Y2=1.805
r123 28 29 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=2.93 $Y=1.805
+ $X2=2.55 $Y2=1.805
r124 27 29 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.465 $Y=1.72
+ $X2=2.55 $Y2=1.805
r125 27 64 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=2.465 $Y=1.72
+ $X2=2.465 $Y2=1.26
r126 24 59 8.39434 $w=4.03e-07 $l=2.95e-07 $layer=LI1_cond $X=2.347 $Y=0.515
+ $X2=2.347 $Y2=0.81
r127 20 63 7.28118 $w=1.7e-07 $l=2.55e-07 $layer=LI1_cond $X=2.04 $Y=1.175
+ $X2=2.295 $Y2=1.175
r128 20 21 98.1872 $w=1.68e-07 $l=1.505e-06 $layer=LI1_cond $X=2.04 $Y=1.175
+ $X2=0.535 $Y2=1.175
r129 16 21 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.41 $Y=1.09
+ $X2=0.535 $Y2=1.175
r130 16 18 26.5062 $w=2.48e-07 $l=5.75e-07 $layer=LI1_cond $X=0.41 $Y=1.09
+ $X2=0.41 $Y2=0.515
r131 5 54 600 $w=1.7e-07 $l=2.59374e-07 $layer=licon1_PDIFF $count=1 $X=3.795
+ $Y=1.84 $X2=3.945 $Y2=2.035
r132 5 38 600 $w=1.7e-07 $l=8.01499e-07 $layer=licon1_PDIFF $count=1 $X=3.795
+ $Y=1.84 $X2=3.945 $Y2=2.57
r133 4 51 600 $w=1.7e-07 $l=2.26164e-07 $layer=licon1_PDIFF $count=1 $X=2.865
+ $Y=1.84 $X2=3.03 $Y2=1.985
r134 4 32 600 $w=1.7e-07 $l=8.08301e-07 $layer=licon1_PDIFF $count=1 $X=2.865
+ $Y=1.84 $X2=3.03 $Y2=2.57
r135 3 44 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=4.19
+ $Y=0.37 $X2=4.33 $Y2=0.515
r136 2 62 182 $w=1.7e-07 $l=7.06965e-07 $layer=licon1_NDIFF $count=1 $X=2.1
+ $Y=0.37 $X2=2.345 $Y2=0.965
r137 2 24 182 $w=1.7e-07 $l=3.09112e-07 $layer=licon1_NDIFF $count=1 $X=2.1
+ $Y=0.37 $X2=2.345 $Y2=0.515
r138 1 18 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.325
+ $Y=0.37 $X2=0.45 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__A22OI_2%A_148_74# 1 2 7 9 11 16
r29 16 17 14.5817 $w=2.51e-07 $l=3e-07 $layer=LI1_cond $X=1.81 $Y=0.535 $X2=1.81
+ $Y2=0.835
r30 12 14 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.965 $Y=0.835
+ $X2=0.84 $Y2=0.835
r31 11 17 3.01842 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.645 $Y=0.835
+ $X2=1.81 $Y2=0.835
r32 11 12 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.645 $Y=0.835
+ $X2=0.965 $Y2=0.835
r33 7 14 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.84 $Y=0.75 $X2=0.84
+ $Y2=0.835
r34 7 9 11.7549 $w=2.48e-07 $l=2.55e-07 $layer=LI1_cond $X=0.84 $Y=0.75 $X2=0.84
+ $Y2=0.495
r35 2 16 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=1.67
+ $Y=0.37 $X2=1.81 $Y2=0.535
r36 1 14 182 $w=1.7e-07 $l=5.30401e-07 $layer=licon1_NDIFF $count=1 $X=0.74
+ $Y=0.37 $X2=0.88 $Y2=0.835
r37 1 9 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=0.74
+ $Y=0.37 $X2=0.88 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_HS__A22OI_2%VGND 1 2 9 13 15 17 22 32 33 36 39
r62 39 40 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r63 36 37 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r64 33 40 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=3.6
+ $Y2=0
r65 32 33 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r66 30 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.635 $Y=0 $X2=3.47
+ $Y2=0
r67 30 32 60.3476 $w=1.68e-07 $l=9.25e-07 $layer=LI1_cond $X=3.635 $Y=0 $X2=4.56
+ $Y2=0
r68 29 40 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=3.6
+ $Y2=0
r69 28 29 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r70 26 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r71 25 28 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.68 $Y=0 $X2=3.12
+ $Y2=0
r72 25 26 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r73 23 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.475 $Y=0 $X2=1.31
+ $Y2=0
r74 23 25 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=1.475 $Y=0 $X2=1.68
+ $Y2=0
r75 22 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.305 $Y=0 $X2=3.47
+ $Y2=0
r76 22 28 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=3.305 $Y=0 $X2=3.12
+ $Y2=0
r77 20 37 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=1.2
+ $Y2=0
r78 19 20 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r79 17 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.145 $Y=0 $X2=1.31
+ $Y2=0
r80 17 19 59.0428 $w=1.68e-07 $l=9.05e-07 $layer=LI1_cond $X=1.145 $Y=0 $X2=0.24
+ $Y2=0
r81 15 29 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=2.4 $Y=0 $X2=3.12
+ $Y2=0
r82 15 26 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=2.4 $Y=0 $X2=1.68
+ $Y2=0
r83 11 39 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.47 $Y=0.085
+ $X2=3.47 $Y2=0
r84 11 13 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=3.47 $Y=0.085
+ $X2=3.47 $Y2=0.495
r85 7 36 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.31 $Y=0.085 $X2=1.31
+ $Y2=0
r86 7 9 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=1.31 $Y=0.085 $X2=1.31
+ $Y2=0.495
r87 2 13 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=3.33
+ $Y=0.37 $X2=3.47 $Y2=0.495
r88 1 9 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=1.17
+ $Y=0.37 $X2=1.31 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_HS__A22OI_2%A_558_74# 1 2 7 9 11 13 15
r28 13 20 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.94 $Y=0.75 $X2=3.94
+ $Y2=0.835
r29 13 15 11.7549 $w=2.48e-07 $l=2.55e-07 $layer=LI1_cond $X=3.94 $Y=0.75
+ $X2=3.94 $Y2=0.495
r30 12 18 4.79851 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=3.135 $Y=0.835
+ $X2=2.985 $Y2=0.835
r31 11 20 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.815 $Y=0.835
+ $X2=3.94 $Y2=0.835
r32 11 12 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=3.815 $Y=0.835
+ $X2=3.135 $Y2=0.835
r33 7 18 2.71916 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.985 $Y=0.75 $X2=2.985
+ $Y2=0.835
r34 7 9 9.79577 $w=2.98e-07 $l=2.55e-07 $layer=LI1_cond $X=2.985 $Y=0.75
+ $X2=2.985 $Y2=0.495
r35 2 20 182 $w=1.7e-07 $l=5.30401e-07 $layer=licon1_NDIFF $count=1 $X=3.76
+ $Y=0.37 $X2=3.9 $Y2=0.835
r36 2 15 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=3.76
+ $Y=0.37 $X2=3.9 $Y2=0.495
r37 1 18 182 $w=1.7e-07 $l=5.60245e-07 $layer=licon1_NDIFF $count=1 $X=2.79
+ $Y=0.37 $X2=3 $Y2=0.835
r38 1 9 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=2.79
+ $Y=0.37 $X2=3 $Y2=0.495
.ends

