* File: sky130_fd_sc_hs__dlxtn_2.pxi.spice
* Created: Tue Sep  1 20:03:03 2020
* 
x_PM_SKY130_FD_SC_HS__DLXTN_2%D N_D_M1017_g N_D_c_136_n N_D_c_140_n N_D_M1008_g
+ D N_D_c_137_n N_D_c_138_n PM_SKY130_FD_SC_HS__DLXTN_2%D
x_PM_SKY130_FD_SC_HS__DLXTN_2%GATE_N N_GATE_N_M1003_g N_GATE_N_c_170_n
+ N_GATE_N_c_171_n N_GATE_N_M1004_g GATE_N N_GATE_N_c_169_n
+ PM_SKY130_FD_SC_HS__DLXTN_2%GATE_N
x_PM_SKY130_FD_SC_HS__DLXTN_2%A_232_82# N_A_232_82#_M1003_d N_A_232_82#_M1004_d
+ N_A_232_82#_c_215_n N_A_232_82#_c_216_n N_A_232_82#_c_232_n
+ N_A_232_82#_M1006_g N_A_232_82#_c_217_n N_A_232_82#_M1009_g
+ N_A_232_82#_c_218_n N_A_232_82#_M1001_g N_A_232_82#_c_219_n
+ N_A_232_82#_c_233_n N_A_232_82#_c_234_n N_A_232_82#_M1010_g
+ N_A_232_82#_c_220_n N_A_232_82#_c_221_n N_A_232_82#_c_222_n
+ N_A_232_82#_c_223_n N_A_232_82#_c_224_n N_A_232_82#_c_225_n
+ N_A_232_82#_c_235_n N_A_232_82#_c_267_p N_A_232_82#_c_236_n
+ N_A_232_82#_c_237_n N_A_232_82#_c_238_n N_A_232_82#_c_239_n
+ N_A_232_82#_c_240_n N_A_232_82#_c_226_n N_A_232_82#_c_227_n
+ N_A_232_82#_c_228_n N_A_232_82#_c_229_n N_A_232_82#_c_230_n
+ PM_SKY130_FD_SC_HS__DLXTN_2%A_232_82#
x_PM_SKY130_FD_SC_HS__DLXTN_2%A_27_120# N_A_27_120#_M1017_s N_A_27_120#_M1008_s
+ N_A_27_120#_c_383_n N_A_27_120#_c_384_n N_A_27_120#_c_394_n
+ N_A_27_120#_M1016_g N_A_27_120#_c_385_n N_A_27_120#_c_386_n
+ N_A_27_120#_M1002_g N_A_27_120#_c_395_n N_A_27_120#_c_387_n
+ N_A_27_120#_c_416_n N_A_27_120#_c_403_n N_A_27_120#_c_388_n
+ N_A_27_120#_c_389_n N_A_27_120#_c_390_n N_A_27_120#_c_391_n
+ N_A_27_120#_c_397_n N_A_27_120#_c_392_n PM_SKY130_FD_SC_HS__DLXTN_2%A_27_120#
x_PM_SKY130_FD_SC_HS__DLXTN_2%A_369_392# N_A_369_392#_M1009_s
+ N_A_369_392#_M1006_s N_A_369_392#_c_503_n N_A_369_392#_M1018_g
+ N_A_369_392#_M1015_g N_A_369_392#_c_504_n N_A_369_392#_c_513_n
+ N_A_369_392#_c_514_n N_A_369_392#_c_505_n N_A_369_392#_c_506_n
+ N_A_369_392#_c_507_n N_A_369_392#_c_508_n N_A_369_392#_c_509_n
+ N_A_369_392#_c_510_n PM_SKY130_FD_SC_HS__DLXTN_2%A_369_392#
x_PM_SKY130_FD_SC_HS__DLXTN_2%A_842_405# N_A_842_405#_M1014_d
+ N_A_842_405#_M1019_d N_A_842_405#_c_616_n N_A_842_405#_M1013_g
+ N_A_842_405#_M1005_g N_A_842_405#_M1000_g N_A_842_405#_c_618_n
+ N_A_842_405#_M1007_g N_A_842_405#_M1012_g N_A_842_405#_c_619_n
+ N_A_842_405#_M1011_g N_A_842_405#_c_610_n N_A_842_405#_c_611_n
+ N_A_842_405#_c_621_n N_A_842_405#_c_622_n N_A_842_405#_c_623_n
+ N_A_842_405#_c_624_n N_A_842_405#_c_612_n N_A_842_405#_c_613_n
+ N_A_842_405#_c_625_n N_A_842_405#_c_662_p N_A_842_405#_c_614_n
+ N_A_842_405#_c_615_n PM_SKY130_FD_SC_HS__DLXTN_2%A_842_405#
x_PM_SKY130_FD_SC_HS__DLXTN_2%A_669_392# N_A_669_392#_M1001_d
+ N_A_669_392#_M1018_d N_A_669_392#_c_705_n N_A_669_392#_M1019_g
+ N_A_669_392#_M1014_g N_A_669_392#_c_707_n N_A_669_392#_c_708_n
+ N_A_669_392#_c_719_n N_A_669_392#_c_709_n
+ PM_SKY130_FD_SC_HS__DLXTN_2%A_669_392#
x_PM_SKY130_FD_SC_HS__DLXTN_2%VPWR N_VPWR_M1008_d N_VPWR_M1006_d N_VPWR_M1013_d
+ N_VPWR_M1007_s N_VPWR_M1011_s N_VPWR_c_774_n N_VPWR_c_775_n N_VPWR_c_776_n
+ N_VPWR_c_777_n N_VPWR_c_778_n N_VPWR_c_779_n N_VPWR_c_780_n N_VPWR_c_781_n
+ N_VPWR_c_782_n VPWR N_VPWR_c_783_n N_VPWR_c_784_n N_VPWR_c_785_n
+ N_VPWR_c_786_n N_VPWR_c_787_n N_VPWR_c_773_n PM_SKY130_FD_SC_HS__DLXTN_2%VPWR
x_PM_SKY130_FD_SC_HS__DLXTN_2%Q N_Q_M1000_d N_Q_M1007_d N_Q_c_861_n N_Q_c_862_n
+ Q Q Q N_Q_c_863_n Q PM_SKY130_FD_SC_HS__DLXTN_2%Q
x_PM_SKY130_FD_SC_HS__DLXTN_2%VGND N_VGND_M1017_d N_VGND_M1009_d N_VGND_M1005_d
+ N_VGND_M1000_s N_VGND_M1012_s N_VGND_c_886_n N_VGND_c_887_n N_VGND_c_888_n
+ N_VGND_c_889_n N_VGND_c_890_n VGND N_VGND_c_891_n N_VGND_c_892_n
+ N_VGND_c_893_n N_VGND_c_894_n N_VGND_c_895_n N_VGND_c_896_n N_VGND_c_897_n
+ N_VGND_c_898_n N_VGND_c_899_n N_VGND_c_900_n PM_SKY130_FD_SC_HS__DLXTN_2%VGND
cc_1 VNB N_D_M1017_g 0.0283486f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.875
cc_2 VNB N_D_c_136_n 0.0015305f $X=-0.19 $Y=-0.245 $X2=0.655 $Y2=1.955
cc_3 VNB N_D_c_137_n 0.00404056f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.465
cc_4 VNB N_D_c_138_n 0.0694963f $X=-0.19 $Y=-0.245 $X2=0.655 $Y2=1.465
cc_5 VNB N_GATE_N_M1003_g 0.0303764f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.875
cc_6 VNB GATE_N 0.00262174f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_7 VNB N_GATE_N_c_169_n 0.0199146f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.465
cc_8 VNB N_A_232_82#_c_215_n 0.011531f $X=-0.19 $Y=-0.245 $X2=0.655 $Y2=2.045
cc_9 VNB N_A_232_82#_c_216_n 0.0168108f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_10 VNB N_A_232_82#_c_217_n 0.0183869f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.465
cc_11 VNB N_A_232_82#_c_218_n 0.0142471f $X=-0.19 $Y=-0.245 $X2=0.655 $Y2=1.465
cc_12 VNB N_A_232_82#_c_219_n 0.0167029f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.665
cc_13 VNB N_A_232_82#_c_220_n 0.00785913f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_232_82#_c_221_n 0.0137619f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_232_82#_c_222_n 0.0286494f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_232_82#_c_223_n 0.00787851f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_232_82#_c_224_n 0.00927555f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_232_82#_c_225_n 0.00410622f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_232_82#_c_226_n 0.039075f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_232_82#_c_227_n 5.48748e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_232_82#_c_228_n 0.020808f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_232_82#_c_229_n 0.00429395f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_232_82#_c_230_n 0.0275096f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_27_120#_c_383_n 0.0484154f $X=-0.19 $Y=-0.245 $X2=0.655 $Y2=2.045
cc_25 VNB N_A_27_120#_c_384_n 0.00179016f $X=-0.19 $Y=-0.245 $X2=0.655 $Y2=2.54
cc_26 VNB N_A_27_120#_c_385_n 0.0194095f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.465
cc_27 VNB N_A_27_120#_c_386_n 0.0158242f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.465
cc_28 VNB N_A_27_120#_c_387_n 0.00560545f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_27_120#_c_388_n 0.0218103f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_27_120#_c_389_n 0.00147483f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_27_120#_c_390_n 0.00304925f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_27_120#_c_391_n 0.0278554f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_27_120#_c_392_n 0.00714823f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_369_392#_c_503_n 0.0205796f $X=-0.19 $Y=-0.245 $X2=0.655 $Y2=2.045
cc_35 VNB N_A_369_392#_c_504_n 0.00241858f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_369_392#_c_505_n 0.00222566f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.665
cc_37 VNB N_A_369_392#_c_506_n 0.00974233f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_369_392#_c_507_n 0.0388791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_369_392#_c_508_n 0.00315129f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_369_392#_c_509_n 0.0080822f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_369_392#_c_510_n 0.0145211f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_842_405#_M1005_g 0.0414386f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.465
cc_43 VNB N_A_842_405#_M1000_g 0.02472f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.465
cc_44 VNB N_A_842_405#_M1012_g 0.0271225f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_A_842_405#_c_610_n 0.0597619f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_A_842_405#_c_611_n 0.0606755f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_842_405#_c_612_n 0.00795778f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_842_405#_c_613_n 0.0034055f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A_842_405#_c_614_n 0.0084286f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_A_842_405#_c_615_n 0.00202256f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_A_669_392#_c_705_n 0.0292853f $X=-0.19 $Y=-0.245 $X2=0.655 $Y2=2.045
cc_52 VNB N_A_669_392#_M1014_g 0.024451f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.465
cc_53 VNB N_A_669_392#_c_707_n 0.0399447f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.465
cc_54 VNB N_A_669_392#_c_708_n 0.00298842f $X=-0.19 $Y=-0.245 $X2=0.655
+ $Y2=1.465
cc_55 VNB N_A_669_392#_c_709_n 0.00379072f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_VPWR_c_773_n 0.302998f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_Q_c_861_n 0.00267235f $X=-0.19 $Y=-0.245 $X2=0.655 $Y2=2.54
cc_58 VNB N_Q_c_862_n 0.00227864f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.465
cc_59 VNB N_Q_c_863_n 0.00373325f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_VGND_c_886_n 0.0103486f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_VGND_c_887_n 0.0103936f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_VGND_c_888_n 0.00786656f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_VGND_c_889_n 0.0122168f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_VGND_c_890_n 0.0542709f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_VGND_c_891_n 0.0195351f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_VGND_c_892_n 0.0439744f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_VGND_c_893_n 0.0430783f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_VGND_c_894_n 0.0200091f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_VGND_c_895_n 0.0172943f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_VGND_c_896_n 0.0196327f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_VGND_c_897_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_VGND_c_898_n 0.00619583f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_VGND_c_899_n 0.0054847f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_VGND_c_900_n 0.422042f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VPB N_D_c_136_n 0.0206902f $X=-0.19 $Y=1.66 $X2=0.655 $Y2=1.955
cc_76 VPB N_D_c_140_n 0.0269575f $X=-0.19 $Y=1.66 $X2=0.655 $Y2=2.045
cc_77 VPB N_D_c_137_n 0.0123656f $X=-0.19 $Y=1.66 $X2=0.29 $Y2=1.465
cc_78 VPB N_GATE_N_c_170_n 0.0110472f $X=-0.19 $Y=1.66 $X2=0.655 $Y2=1.955
cc_79 VPB N_GATE_N_c_171_n 0.027385f $X=-0.19 $Y=1.66 $X2=0.655 $Y2=2.045
cc_80 VPB GATE_N 0.00260948f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_81 VPB N_GATE_N_c_169_n 0.0127652f $X=-0.19 $Y=1.66 $X2=0.29 $Y2=1.465
cc_82 VPB N_A_232_82#_c_216_n 0.00790287f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_83 VPB N_A_232_82#_c_232_n 0.0247527f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_84 VPB N_A_232_82#_c_233_n 0.0317657f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_85 VPB N_A_232_82#_c_234_n 0.0202606f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_86 VPB N_A_232_82#_c_235_n 0.00641792f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_87 VPB N_A_232_82#_c_236_n 0.00861901f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_88 VPB N_A_232_82#_c_237_n 8.72539e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_89 VPB N_A_232_82#_c_238_n 0.012783f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_90 VPB N_A_232_82#_c_239_n 0.0235844f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_91 VPB N_A_232_82#_c_240_n 0.00684486f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_92 VPB N_A_232_82#_c_227_n 0.00380583f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_93 VPB N_A_232_82#_c_228_n 0.0162329f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_94 VPB N_A_232_82#_c_229_n 0.00223583f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_95 VPB N_A_232_82#_c_230_n 0.0252921f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_96 VPB N_A_27_120#_c_384_n 0.00827177f $X=-0.19 $Y=1.66 $X2=0.655 $Y2=2.54
cc_97 VPB N_A_27_120#_c_394_n 0.0206811f $X=-0.19 $Y=1.66 $X2=0.655 $Y2=2.54
cc_98 VPB N_A_27_120#_c_395_n 0.0360197f $X=-0.19 $Y=1.66 $X2=0.29 $Y2=1.465
cc_99 VPB N_A_27_120#_c_387_n 0.00273869f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_100 VPB N_A_27_120#_c_397_n 0.0142359f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_101 VPB N_A_369_392#_c_503_n 0.0344759f $X=-0.19 $Y=1.66 $X2=0.655 $Y2=2.045
cc_102 VPB N_A_369_392#_c_504_n 0.00104552f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_103 VPB N_A_369_392#_c_513_n 0.0089307f $X=-0.19 $Y=1.66 $X2=0.655 $Y2=1.465
cc_104 VPB N_A_369_392#_c_514_n 0.0101851f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_105 VPB N_A_369_392#_c_508_n 0.00117638f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_106 VPB N_A_842_405#_c_616_n 0.0181711f $X=-0.19 $Y=1.66 $X2=0.655 $Y2=2.045
cc_107 VPB N_A_842_405#_M1005_g 0.0234795f $X=-0.19 $Y=1.66 $X2=0.29 $Y2=1.465
cc_108 VPB N_A_842_405#_c_618_n 0.0171142f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_109 VPB N_A_842_405#_c_619_n 0.0181803f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_110 VPB N_A_842_405#_c_611_n 0.0181745f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_111 VPB N_A_842_405#_c_621_n 0.00410771f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_112 VPB N_A_842_405#_c_622_n 0.0649433f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_113 VPB N_A_842_405#_c_623_n 0.0125822f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_114 VPB N_A_842_405#_c_624_n 0.00847633f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_115 VPB N_A_842_405#_c_625_n 0.00352309f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_116 VPB N_A_669_392#_c_705_n 0.0246656f $X=-0.19 $Y=1.66 $X2=0.655 $Y2=2.045
cc_117 VPB N_A_669_392#_c_709_n 0.00187927f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_118 VPB N_VPWR_c_774_n 0.00970163f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_119 VPB N_VPWR_c_775_n 0.014119f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_120 VPB N_VPWR_c_776_n 0.0115203f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_121 VPB N_VPWR_c_777_n 0.0106521f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_122 VPB N_VPWR_c_778_n 0.0646533f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_123 VPB N_VPWR_c_779_n 0.0239248f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_124 VPB N_VPWR_c_780_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_125 VPB N_VPWR_c_781_n 0.0218405f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_126 VPB N_VPWR_c_782_n 0.00410958f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_127 VPB N_VPWR_c_783_n 0.0345071f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_128 VPB N_VPWR_c_784_n 0.0221566f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_129 VPB N_VPWR_c_785_n 0.00660399f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_130 VPB N_VPWR_c_786_n 0.0393577f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_131 VPB N_VPWR_c_787_n 0.0265436f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_132 VPB N_VPWR_c_773_n 0.108245f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_133 VPB N_Q_c_863_n 0.00322055f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_134 N_D_M1017_g N_GATE_N_M1003_g 0.0184595f $X=0.495 $Y=0.875 $X2=0 $Y2=0
cc_135 N_D_c_138_n N_GATE_N_M1003_g 0.00663446f $X=0.655 $Y=1.465 $X2=0 $Y2=0
cc_136 N_D_c_136_n N_GATE_N_c_170_n 0.00382806f $X=0.655 $Y=1.955 $X2=0 $Y2=0
cc_137 N_D_c_140_n N_GATE_N_c_171_n 0.0266829f $X=0.655 $Y=2.045 $X2=0 $Y2=0
cc_138 N_D_c_138_n GATE_N 3.81053e-19 $X=0.655 $Y=1.465 $X2=0 $Y2=0
cc_139 N_D_c_138_n N_GATE_N_c_169_n 0.0174277f $X=0.655 $Y=1.465 $X2=0 $Y2=0
cc_140 N_D_c_140_n N_A_232_82#_c_239_n 6.85969e-19 $X=0.655 $Y=2.045 $X2=0 $Y2=0
cc_141 N_D_c_140_n N_A_27_120#_c_395_n 0.0137897f $X=0.655 $Y=2.045 $X2=0 $Y2=0
cc_142 N_D_M1017_g N_A_27_120#_c_387_n 0.00397398f $X=0.495 $Y=0.875 $X2=0 $Y2=0
cc_143 N_D_c_136_n N_A_27_120#_c_387_n 0.0129118f $X=0.655 $Y=1.955 $X2=0 $Y2=0
cc_144 N_D_c_137_n N_A_27_120#_c_387_n 0.0348574f $X=0.29 $Y=1.465 $X2=0 $Y2=0
cc_145 N_D_c_138_n N_A_27_120#_c_387_n 0.0116014f $X=0.655 $Y=1.465 $X2=0 $Y2=0
cc_146 N_D_M1017_g N_A_27_120#_c_403_n 4.90322e-19 $X=0.495 $Y=0.875 $X2=0 $Y2=0
cc_147 N_D_M1017_g N_A_27_120#_c_391_n 0.0266287f $X=0.495 $Y=0.875 $X2=0 $Y2=0
cc_148 N_D_c_137_n N_A_27_120#_c_391_n 0.024806f $X=0.29 $Y=1.465 $X2=0 $Y2=0
cc_149 N_D_c_138_n N_A_27_120#_c_391_n 0.0026784f $X=0.655 $Y=1.465 $X2=0 $Y2=0
cc_150 N_D_c_136_n N_A_27_120#_c_397_n 0.00304242f $X=0.655 $Y=1.955 $X2=0 $Y2=0
cc_151 N_D_c_140_n N_A_27_120#_c_397_n 0.0135169f $X=0.655 $Y=2.045 $X2=0 $Y2=0
cc_152 N_D_c_137_n N_A_27_120#_c_397_n 0.0155123f $X=0.29 $Y=1.465 $X2=0 $Y2=0
cc_153 N_D_c_138_n N_A_27_120#_c_397_n 0.00484569f $X=0.655 $Y=1.465 $X2=0 $Y2=0
cc_154 N_D_c_140_n N_VPWR_c_774_n 0.00737447f $X=0.655 $Y=2.045 $X2=0 $Y2=0
cc_155 N_D_c_140_n N_VPWR_c_779_n 0.00445602f $X=0.655 $Y=2.045 $X2=0 $Y2=0
cc_156 N_D_c_140_n N_VPWR_c_773_n 0.0086172f $X=0.655 $Y=2.045 $X2=0 $Y2=0
cc_157 N_D_M1017_g N_VGND_c_891_n 0.00327294f $X=0.495 $Y=0.875 $X2=0 $Y2=0
cc_158 N_D_M1017_g N_VGND_c_900_n 0.00476395f $X=0.495 $Y=0.875 $X2=0 $Y2=0
cc_159 N_GATE_N_M1003_g N_A_232_82#_c_223_n 0.00461345f $X=1.085 $Y=0.78 $X2=0
+ $Y2=0
cc_160 GATE_N N_A_232_82#_c_223_n 0.00948482f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_161 N_GATE_N_c_169_n N_A_232_82#_c_223_n 0.00100823f $X=1.15 $Y=1.615 $X2=0
+ $Y2=0
cc_162 N_GATE_N_M1003_g N_A_232_82#_c_224_n 0.00303911f $X=1.085 $Y=0.78 $X2=0
+ $Y2=0
cc_163 N_GATE_N_M1003_g N_A_232_82#_c_225_n 0.00593761f $X=1.085 $Y=0.78 $X2=0
+ $Y2=0
cc_164 GATE_N N_A_232_82#_c_225_n 0.0263887f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_165 N_GATE_N_c_169_n N_A_232_82#_c_225_n 0.00218737f $X=1.15 $Y=1.615 $X2=0
+ $Y2=0
cc_166 N_GATE_N_c_171_n N_A_232_82#_c_235_n 4.4113e-19 $X=1.205 $Y=2.045 $X2=0
+ $Y2=0
cc_167 N_GATE_N_c_171_n N_A_232_82#_c_239_n 0.0153928f $X=1.205 $Y=2.045 $X2=0
+ $Y2=0
cc_168 GATE_N N_A_232_82#_c_239_n 0.00246946f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_169 N_GATE_N_c_170_n N_A_232_82#_c_240_n 0.00903071f $X=1.205 $Y=1.955 $X2=0
+ $Y2=0
cc_170 N_GATE_N_c_171_n N_A_232_82#_c_240_n 0.00178037f $X=1.205 $Y=2.045 $X2=0
+ $Y2=0
cc_171 N_GATE_N_M1003_g N_A_232_82#_c_226_n 0.014014f $X=1.085 $Y=0.78 $X2=0
+ $Y2=0
cc_172 GATE_N N_A_232_82#_c_228_n 3.56619e-19 $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_173 N_GATE_N_c_169_n N_A_232_82#_c_228_n 0.0168587f $X=1.15 $Y=1.615 $X2=0
+ $Y2=0
cc_174 N_GATE_N_c_171_n N_A_27_120#_c_395_n 6.6422e-19 $X=1.205 $Y=2.045 $X2=0
+ $Y2=0
cc_175 N_GATE_N_M1003_g N_A_27_120#_c_387_n 0.0059942f $X=1.085 $Y=0.78 $X2=0
+ $Y2=0
cc_176 N_GATE_N_c_170_n N_A_27_120#_c_387_n 0.00308057f $X=1.205 $Y=1.955 $X2=0
+ $Y2=0
cc_177 GATE_N N_A_27_120#_c_387_n 0.0228108f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_178 N_GATE_N_c_169_n N_A_27_120#_c_387_n 0.00187493f $X=1.15 $Y=1.615 $X2=0
+ $Y2=0
cc_179 N_GATE_N_M1003_g N_A_27_120#_c_416_n 0.0164833f $X=1.085 $Y=0.78 $X2=0
+ $Y2=0
cc_180 N_GATE_N_M1003_g N_A_27_120#_c_403_n 0.00644004f $X=1.085 $Y=0.78 $X2=0
+ $Y2=0
cc_181 N_GATE_N_M1003_g N_A_27_120#_c_389_n 0.00578481f $X=1.085 $Y=0.78 $X2=0
+ $Y2=0
cc_182 N_GATE_N_M1003_g N_A_27_120#_c_391_n 0.00668497f $X=1.085 $Y=0.78 $X2=0
+ $Y2=0
cc_183 N_GATE_N_c_170_n N_A_27_120#_c_397_n 0.00212053f $X=1.205 $Y=1.955 $X2=0
+ $Y2=0
cc_184 N_GATE_N_c_171_n N_A_27_120#_c_397_n 0.00138504f $X=1.205 $Y=2.045 $X2=0
+ $Y2=0
cc_185 N_GATE_N_c_171_n N_A_369_392#_c_514_n 2.71171e-19 $X=1.205 $Y=2.045 $X2=0
+ $Y2=0
cc_186 N_GATE_N_c_171_n N_VPWR_c_774_n 0.00737447f $X=1.205 $Y=2.045 $X2=0 $Y2=0
cc_187 GATE_N N_VPWR_c_774_n 0.00338659f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_188 N_GATE_N_c_169_n N_VPWR_c_774_n 6.22093e-19 $X=1.15 $Y=1.615 $X2=0 $Y2=0
cc_189 N_GATE_N_c_171_n N_VPWR_c_783_n 0.00445602f $X=1.205 $Y=2.045 $X2=0 $Y2=0
cc_190 N_GATE_N_c_171_n N_VPWR_c_773_n 0.00862626f $X=1.205 $Y=2.045 $X2=0 $Y2=0
cc_191 N_GATE_N_M1003_g N_VGND_c_892_n 0.00382493f $X=1.085 $Y=0.78 $X2=0 $Y2=0
cc_192 N_GATE_N_M1003_g N_VGND_c_896_n 0.0029536f $X=1.085 $Y=0.78 $X2=0 $Y2=0
cc_193 N_GATE_N_M1003_g N_VGND_c_900_n 0.00479772f $X=1.085 $Y=0.78 $X2=0 $Y2=0
cc_194 N_A_232_82#_c_216_n N_A_27_120#_c_383_n 0.00952668f $X=2.215 $Y=1.795
+ $X2=0 $Y2=0
cc_195 N_A_232_82#_c_217_n N_A_27_120#_c_383_n 0.00378548f $X=2.355 $Y=1.185
+ $X2=0 $Y2=0
cc_196 N_A_232_82#_c_221_n N_A_27_120#_c_383_n 0.00491582f $X=2.355 $Y=1.26
+ $X2=0 $Y2=0
cc_197 N_A_232_82#_c_216_n N_A_27_120#_c_384_n 0.00329427f $X=2.215 $Y=1.795
+ $X2=0 $Y2=0
cc_198 N_A_232_82#_c_232_n N_A_27_120#_c_394_n 0.028046f $X=2.215 $Y=1.885 $X2=0
+ $Y2=0
cc_199 N_A_232_82#_c_235_n N_A_27_120#_c_394_n 0.0123901f $X=2.875 $Y=2.525
+ $X2=0 $Y2=0
cc_200 N_A_232_82#_c_267_p N_A_27_120#_c_394_n 0.00707689f $X=2.96 $Y=2.905
+ $X2=0 $Y2=0
cc_201 N_A_232_82#_c_237_n N_A_27_120#_c_394_n 0.00428477f $X=3.045 $Y=2.99
+ $X2=0 $Y2=0
cc_202 N_A_232_82#_c_222_n N_A_27_120#_c_385_n 0.0229627f $X=3.825 $Y=1.185
+ $X2=0 $Y2=0
cc_203 N_A_232_82#_c_217_n N_A_27_120#_c_386_n 0.00442582f $X=2.355 $Y=1.185
+ $X2=0 $Y2=0
cc_204 N_A_232_82#_c_218_n N_A_27_120#_c_386_n 0.0229627f $X=3.605 $Y=1.11 $X2=0
+ $Y2=0
cc_205 N_A_232_82#_c_239_n N_A_27_120#_c_395_n 0.0041043f $X=1.43 $Y=2.265 $X2=0
+ $Y2=0
cc_206 N_A_232_82#_c_223_n N_A_27_120#_c_387_n 0.00182037f $X=1.485 $Y=1.045
+ $X2=0 $Y2=0
cc_207 N_A_232_82#_M1003_d N_A_27_120#_c_416_n 0.00866525f $X=1.16 $Y=0.41 $X2=0
+ $Y2=0
cc_208 N_A_232_82#_c_223_n N_A_27_120#_c_416_n 0.00975585f $X=1.485 $Y=1.045
+ $X2=0 $Y2=0
cc_209 N_A_232_82#_M1003_d N_A_27_120#_c_403_n 0.0058378f $X=1.16 $Y=0.41 $X2=0
+ $Y2=0
cc_210 N_A_232_82#_M1003_d N_A_27_120#_c_388_n 0.00239893f $X=1.16 $Y=0.41 $X2=0
+ $Y2=0
cc_211 N_A_232_82#_c_217_n N_A_27_120#_c_388_n 0.0157054f $X=2.355 $Y=1.185
+ $X2=0 $Y2=0
cc_212 N_A_232_82#_c_223_n N_A_27_120#_c_388_n 0.00585336f $X=1.485 $Y=1.045
+ $X2=0 $Y2=0
cc_213 N_A_232_82#_c_224_n N_A_27_120#_c_388_n 0.0169889f $X=1.685 $Y=1.17 $X2=0
+ $Y2=0
cc_214 N_A_232_82#_c_226_n N_A_27_120#_c_388_n 0.00199179f $X=1.72 $Y=0.925
+ $X2=0 $Y2=0
cc_215 N_A_232_82#_c_217_n N_A_27_120#_c_390_n 0.00800558f $X=2.355 $Y=1.185
+ $X2=0 $Y2=0
cc_216 N_A_232_82#_c_223_n N_A_27_120#_c_391_n 0.0106332f $X=1.485 $Y=1.045
+ $X2=0 $Y2=0
cc_217 N_A_232_82#_c_239_n N_A_27_120#_c_397_n 7.413e-19 $X=1.43 $Y=2.265 $X2=0
+ $Y2=0
cc_218 N_A_232_82#_c_216_n N_A_27_120#_c_392_n 0.00202018f $X=2.215 $Y=1.795
+ $X2=0 $Y2=0
cc_219 N_A_232_82#_c_221_n N_A_27_120#_c_392_n 2.84937e-19 $X=2.355 $Y=1.26
+ $X2=0 $Y2=0
cc_220 N_A_232_82#_c_235_n N_A_369_392#_M1006_s 0.00811065f $X=2.875 $Y=2.525
+ $X2=0 $Y2=0
cc_221 N_A_232_82#_c_219_n N_A_369_392#_c_503_n 0.0174101f $X=3.825 $Y=1.485
+ $X2=0 $Y2=0
cc_222 N_A_232_82#_c_233_n N_A_369_392#_c_503_n 0.0100472f $X=3.88 $Y=2.35 $X2=0
+ $Y2=0
cc_223 N_A_232_82#_c_234_n N_A_369_392#_c_503_n 0.0104438f $X=3.88 $Y=2.44 $X2=0
+ $Y2=0
cc_224 N_A_232_82#_c_235_n N_A_369_392#_c_503_n 0.00143509f $X=2.875 $Y=2.525
+ $X2=0 $Y2=0
cc_225 N_A_232_82#_c_267_p N_A_369_392#_c_503_n 0.00443826f $X=2.96 $Y=2.905
+ $X2=0 $Y2=0
cc_226 N_A_232_82#_c_236_n N_A_369_392#_c_503_n 0.0141045f $X=4.02 $Y=2.99 $X2=0
+ $Y2=0
cc_227 N_A_232_82#_c_230_n N_A_369_392#_c_503_n 4.34343e-19 $X=4.185 $Y=1.65
+ $X2=0 $Y2=0
cc_228 N_A_232_82#_c_215_n N_A_369_392#_c_504_n 0.00462651f $X=2.125 $Y=1.26
+ $X2=0 $Y2=0
cc_229 N_A_232_82#_c_216_n N_A_369_392#_c_504_n 0.0137549f $X=2.215 $Y=1.795
+ $X2=0 $Y2=0
cc_230 N_A_232_82#_c_217_n N_A_369_392#_c_504_n 0.0094035f $X=2.355 $Y=1.185
+ $X2=0 $Y2=0
cc_231 N_A_232_82#_c_221_n N_A_369_392#_c_504_n 0.00522206f $X=2.355 $Y=1.26
+ $X2=0 $Y2=0
cc_232 N_A_232_82#_c_224_n N_A_369_392#_c_504_n 0.0326777f $X=1.685 $Y=1.17
+ $X2=0 $Y2=0
cc_233 N_A_232_82#_c_225_n N_A_369_392#_c_504_n 0.046382f $X=1.685 $Y=1.57 $X2=0
+ $Y2=0
cc_234 N_A_232_82#_c_240_n N_A_369_392#_c_504_n 0.00124535f $X=1.46 $Y=2.1 $X2=0
+ $Y2=0
cc_235 N_A_232_82#_c_226_n N_A_369_392#_c_504_n 0.00162222f $X=1.72 $Y=0.925
+ $X2=0 $Y2=0
cc_236 N_A_232_82#_c_228_n N_A_369_392#_c_504_n 0.00255297f $X=1.72 $Y=1.605
+ $X2=0 $Y2=0
cc_237 N_A_232_82#_c_221_n N_A_369_392#_c_513_n 0.00379117f $X=2.355 $Y=1.26
+ $X2=0 $Y2=0
cc_238 N_A_232_82#_c_235_n N_A_369_392#_c_513_n 0.0197139f $X=2.875 $Y=2.525
+ $X2=0 $Y2=0
cc_239 N_A_232_82#_c_215_n N_A_369_392#_c_514_n 0.00141981f $X=2.125 $Y=1.26
+ $X2=0 $Y2=0
cc_240 N_A_232_82#_c_232_n N_A_369_392#_c_514_n 0.0193539f $X=2.215 $Y=1.885
+ $X2=0 $Y2=0
cc_241 N_A_232_82#_c_235_n N_A_369_392#_c_514_n 0.0285924f $X=2.875 $Y=2.525
+ $X2=0 $Y2=0
cc_242 N_A_232_82#_c_240_n N_A_369_392#_c_514_n 0.0341527f $X=1.46 $Y=2.1 $X2=0
+ $Y2=0
cc_243 N_A_232_82#_c_227_n N_A_369_392#_c_514_n 0.00497552f $X=1.72 $Y=1.605
+ $X2=0 $Y2=0
cc_244 N_A_232_82#_c_228_n N_A_369_392#_c_514_n 4.32246e-19 $X=1.72 $Y=1.605
+ $X2=0 $Y2=0
cc_245 N_A_232_82#_c_218_n N_A_369_392#_c_506_n 0.0198684f $X=3.605 $Y=1.11
+ $X2=0 $Y2=0
cc_246 N_A_232_82#_c_222_n N_A_369_392#_c_506_n 0.0014907f $X=3.825 $Y=1.185
+ $X2=0 $Y2=0
cc_247 N_A_232_82#_c_218_n N_A_369_392#_c_507_n 0.0101699f $X=3.605 $Y=1.11
+ $X2=0 $Y2=0
cc_248 N_A_232_82#_c_219_n N_A_369_392#_c_508_n 3.61841e-19 $X=3.825 $Y=1.485
+ $X2=0 $Y2=0
cc_249 N_A_232_82#_c_233_n N_A_369_392#_c_508_n 4.6879e-19 $X=3.88 $Y=2.35 $X2=0
+ $Y2=0
cc_250 N_A_232_82#_c_218_n N_A_369_392#_c_509_n 0.00336691f $X=3.605 $Y=1.11
+ $X2=0 $Y2=0
cc_251 N_A_232_82#_c_219_n N_A_369_392#_c_509_n 0.00121983f $X=3.825 $Y=1.485
+ $X2=0 $Y2=0
cc_252 N_A_232_82#_c_218_n N_A_369_392#_c_510_n 0.0109494f $X=3.605 $Y=1.11
+ $X2=0 $Y2=0
cc_253 N_A_232_82#_c_222_n N_A_369_392#_c_510_n 0.00477162f $X=3.825 $Y=1.185
+ $X2=0 $Y2=0
cc_254 N_A_232_82#_c_230_n N_A_369_392#_c_510_n 0.00690996f $X=4.185 $Y=1.65
+ $X2=0 $Y2=0
cc_255 N_A_232_82#_c_234_n N_A_842_405#_c_616_n 0.0237787f $X=3.88 $Y=2.44 $X2=0
+ $Y2=0
cc_256 N_A_232_82#_c_236_n N_A_842_405#_c_616_n 0.00119814f $X=4.02 $Y=2.99
+ $X2=0 $Y2=0
cc_257 N_A_232_82#_c_238_n N_A_842_405#_c_616_n 0.00345868f $X=4.105 $Y=2.905
+ $X2=0 $Y2=0
cc_258 N_A_232_82#_c_233_n N_A_842_405#_M1005_g 0.00224512f $X=3.88 $Y=2.35
+ $X2=0 $Y2=0
cc_259 N_A_232_82#_c_222_n N_A_842_405#_M1005_g 0.00421996f $X=3.825 $Y=1.185
+ $X2=0 $Y2=0
cc_260 N_A_232_82#_c_238_n N_A_842_405#_M1005_g 0.00366868f $X=4.105 $Y=2.905
+ $X2=0 $Y2=0
cc_261 N_A_232_82#_c_229_n N_A_842_405#_M1005_g 0.00176725f $X=4.185 $Y=1.65
+ $X2=0 $Y2=0
cc_262 N_A_232_82#_c_230_n N_A_842_405#_M1005_g 0.0170611f $X=4.185 $Y=1.65
+ $X2=0 $Y2=0
cc_263 N_A_232_82#_c_238_n N_A_842_405#_c_621_n 0.0262086f $X=4.105 $Y=2.905
+ $X2=0 $Y2=0
cc_264 N_A_232_82#_c_233_n N_A_842_405#_c_622_n 0.0198173f $X=3.88 $Y=2.35 $X2=0
+ $Y2=0
cc_265 N_A_232_82#_c_238_n N_A_842_405#_c_622_n 0.0048616f $X=4.105 $Y=2.905
+ $X2=0 $Y2=0
cc_266 N_A_232_82#_c_229_n N_A_842_405#_c_622_n 0.00106548f $X=4.185 $Y=1.65
+ $X2=0 $Y2=0
cc_267 N_A_232_82#_c_230_n N_A_842_405#_c_622_n 0.0093115f $X=4.185 $Y=1.65
+ $X2=0 $Y2=0
cc_268 N_A_232_82#_c_236_n N_A_669_392#_M1018_d 0.00395618f $X=4.02 $Y=2.99
+ $X2=0 $Y2=0
cc_269 N_A_232_82#_c_229_n N_A_669_392#_c_707_n 0.0114859f $X=4.185 $Y=1.65
+ $X2=0 $Y2=0
cc_270 N_A_232_82#_c_230_n N_A_669_392#_c_707_n 2.9672e-19 $X=4.185 $Y=1.65
+ $X2=0 $Y2=0
cc_271 N_A_232_82#_c_218_n N_A_669_392#_c_708_n 0.00856348f $X=3.605 $Y=1.11
+ $X2=0 $Y2=0
cc_272 N_A_232_82#_c_222_n N_A_669_392#_c_708_n 0.00190905f $X=3.825 $Y=1.185
+ $X2=0 $Y2=0
cc_273 N_A_232_82#_c_229_n N_A_669_392#_c_708_n 0.0149091f $X=4.185 $Y=1.65
+ $X2=0 $Y2=0
cc_274 N_A_232_82#_c_230_n N_A_669_392#_c_708_n 0.00507885f $X=4.185 $Y=1.65
+ $X2=0 $Y2=0
cc_275 N_A_232_82#_c_233_n N_A_669_392#_c_719_n 0.0062152f $X=3.88 $Y=2.35 $X2=0
+ $Y2=0
cc_276 N_A_232_82#_c_234_n N_A_669_392#_c_719_n 0.011887f $X=3.88 $Y=2.44 $X2=0
+ $Y2=0
cc_277 N_A_232_82#_c_235_n N_A_669_392#_c_719_n 0.00974339f $X=2.875 $Y=2.525
+ $X2=0 $Y2=0
cc_278 N_A_232_82#_c_267_p N_A_669_392#_c_719_n 0.00640516f $X=2.96 $Y=2.905
+ $X2=0 $Y2=0
cc_279 N_A_232_82#_c_236_n N_A_669_392#_c_719_n 0.0302047f $X=4.02 $Y=2.99 $X2=0
+ $Y2=0
cc_280 N_A_232_82#_c_238_n N_A_669_392#_c_719_n 0.046327f $X=4.105 $Y=2.905
+ $X2=0 $Y2=0
cc_281 N_A_232_82#_c_218_n N_A_669_392#_c_709_n 6.33047e-19 $X=3.605 $Y=1.11
+ $X2=0 $Y2=0
cc_282 N_A_232_82#_c_219_n N_A_669_392#_c_709_n 0.0120805f $X=3.825 $Y=1.485
+ $X2=0 $Y2=0
cc_283 N_A_232_82#_c_233_n N_A_669_392#_c_709_n 0.00749785f $X=3.88 $Y=2.35
+ $X2=0 $Y2=0
cc_284 N_A_232_82#_c_222_n N_A_669_392#_c_709_n 0.00989251f $X=3.825 $Y=1.185
+ $X2=0 $Y2=0
cc_285 N_A_232_82#_c_229_n N_A_669_392#_c_709_n 0.046327f $X=4.185 $Y=1.65 $X2=0
+ $Y2=0
cc_286 N_A_232_82#_c_230_n N_A_669_392#_c_709_n 0.0100291f $X=4.185 $Y=1.65
+ $X2=0 $Y2=0
cc_287 N_A_232_82#_c_235_n N_VPWR_M1006_d 0.0116948f $X=2.875 $Y=2.525 $X2=0
+ $Y2=0
cc_288 N_A_232_82#_c_239_n N_VPWR_c_774_n 0.0273513f $X=1.43 $Y=2.265 $X2=0
+ $Y2=0
cc_289 N_A_232_82#_c_232_n N_VPWR_c_775_n 0.00438753f $X=2.215 $Y=1.885 $X2=0
+ $Y2=0
cc_290 N_A_232_82#_c_235_n N_VPWR_c_775_n 0.0267961f $X=2.875 $Y=2.525 $X2=0
+ $Y2=0
cc_291 N_A_232_82#_c_267_p N_VPWR_c_775_n 0.00924851f $X=2.96 $Y=2.905 $X2=0
+ $Y2=0
cc_292 N_A_232_82#_c_237_n N_VPWR_c_775_n 0.0142284f $X=3.045 $Y=2.99 $X2=0
+ $Y2=0
cc_293 N_A_232_82#_c_232_n N_VPWR_c_783_n 0.00366846f $X=2.215 $Y=1.885 $X2=0
+ $Y2=0
cc_294 N_A_232_82#_c_235_n N_VPWR_c_783_n 0.00949357f $X=2.875 $Y=2.525 $X2=0
+ $Y2=0
cc_295 N_A_232_82#_c_239_n N_VPWR_c_783_n 0.0172711f $X=1.43 $Y=2.265 $X2=0
+ $Y2=0
cc_296 N_A_232_82#_c_234_n N_VPWR_c_786_n 9.44495e-19 $X=3.88 $Y=2.44 $X2=0
+ $Y2=0
cc_297 N_A_232_82#_c_235_n N_VPWR_c_786_n 0.00197454f $X=2.875 $Y=2.525 $X2=0
+ $Y2=0
cc_298 N_A_232_82#_c_236_n N_VPWR_c_786_n 0.0744997f $X=4.02 $Y=2.99 $X2=0 $Y2=0
cc_299 N_A_232_82#_c_237_n N_VPWR_c_786_n 0.0119496f $X=3.045 $Y=2.99 $X2=0
+ $Y2=0
cc_300 N_A_232_82#_c_236_n N_VPWR_c_787_n 0.0138115f $X=4.02 $Y=2.99 $X2=0 $Y2=0
cc_301 N_A_232_82#_c_232_n N_VPWR_c_773_n 0.0049649f $X=2.215 $Y=1.885 $X2=0
+ $Y2=0
cc_302 N_A_232_82#_c_235_n N_VPWR_c_773_n 0.0241361f $X=2.875 $Y=2.525 $X2=0
+ $Y2=0
cc_303 N_A_232_82#_c_236_n N_VPWR_c_773_n 0.0425764f $X=4.02 $Y=2.99 $X2=0 $Y2=0
cc_304 N_A_232_82#_c_237_n N_VPWR_c_773_n 0.00636858f $X=3.045 $Y=2.99 $X2=0
+ $Y2=0
cc_305 N_A_232_82#_c_239_n N_VPWR_c_773_n 0.0142626f $X=1.43 $Y=2.265 $X2=0
+ $Y2=0
cc_306 N_A_232_82#_c_235_n A_585_392# 0.0029667f $X=2.875 $Y=2.525 $X2=-0.19
+ $Y2=-0.245
cc_307 N_A_232_82#_c_267_p A_585_392# 0.00320536f $X=2.96 $Y=2.905 $X2=-0.19
+ $Y2=-0.245
cc_308 N_A_232_82#_c_236_n A_585_392# 0.00351031f $X=4.02 $Y=2.99 $X2=-0.19
+ $Y2=-0.245
cc_309 N_A_232_82#_c_236_n A_791_503# 3.21886e-19 $X=4.02 $Y=2.99 $X2=-0.19
+ $Y2=-0.245
cc_310 N_A_232_82#_c_238_n A_791_503# 0.0056027f $X=4.105 $Y=2.905 $X2=-0.19
+ $Y2=-0.245
cc_311 N_A_232_82#_c_217_n N_VGND_c_886_n 0.00196494f $X=2.355 $Y=1.185 $X2=0
+ $Y2=0
cc_312 N_A_232_82#_c_218_n N_VGND_c_886_n 3.70241e-19 $X=3.605 $Y=1.11 $X2=0
+ $Y2=0
cc_313 N_A_232_82#_c_217_n N_VGND_c_892_n 0.00278271f $X=2.355 $Y=1.185 $X2=0
+ $Y2=0
cc_314 N_A_232_82#_c_218_n N_VGND_c_893_n 9.44495e-19 $X=3.605 $Y=1.11 $X2=0
+ $Y2=0
cc_315 N_A_232_82#_c_217_n N_VGND_c_900_n 0.00363426f $X=2.355 $Y=1.185 $X2=0
+ $Y2=0
cc_316 N_A_27_120#_c_388_n N_A_369_392#_M1009_s 0.00441657f $X=2.475 $Y=0.34
+ $X2=-0.19 $Y2=-0.245
cc_317 N_A_27_120#_c_383_n N_A_369_392#_c_503_n 0.0100759f $X=2.85 $Y=1.63 $X2=0
+ $Y2=0
cc_318 N_A_27_120#_c_384_n N_A_369_392#_c_503_n 0.0142064f $X=2.85 $Y=1.795
+ $X2=0 $Y2=0
cc_319 N_A_27_120#_c_394_n N_A_369_392#_c_503_n 0.0556071f $X=2.85 $Y=1.885
+ $X2=0 $Y2=0
cc_320 N_A_27_120#_c_385_n N_A_369_392#_c_503_n 0.0073783f $X=3.14 $Y=1.185
+ $X2=0 $Y2=0
cc_321 N_A_27_120#_c_392_n N_A_369_392#_c_503_n 5.53572e-19 $X=2.805 $Y=1.465
+ $X2=0 $Y2=0
cc_322 N_A_27_120#_c_383_n N_A_369_392#_c_504_n 3.44763e-19 $X=2.85 $Y=1.63
+ $X2=0 $Y2=0
cc_323 N_A_27_120#_c_384_n N_A_369_392#_c_504_n 9.53103e-19 $X=2.85 $Y=1.795
+ $X2=0 $Y2=0
cc_324 N_A_27_120#_c_388_n N_A_369_392#_c_504_n 0.0144209f $X=2.475 $Y=0.34
+ $X2=0 $Y2=0
cc_325 N_A_27_120#_c_390_n N_A_369_392#_c_504_n 0.0324263f $X=2.56 $Y=1.3 $X2=0
+ $Y2=0
cc_326 N_A_27_120#_c_392_n N_A_369_392#_c_504_n 0.0263966f $X=2.805 $Y=1.465
+ $X2=0 $Y2=0
cc_327 N_A_27_120#_c_383_n N_A_369_392#_c_513_n 0.00349359f $X=2.85 $Y=1.63
+ $X2=0 $Y2=0
cc_328 N_A_27_120#_c_394_n N_A_369_392#_c_513_n 0.0135965f $X=2.85 $Y=1.885
+ $X2=0 $Y2=0
cc_329 N_A_27_120#_c_385_n N_A_369_392#_c_513_n 0.0050599f $X=3.14 $Y=1.185
+ $X2=0 $Y2=0
cc_330 N_A_27_120#_c_392_n N_A_369_392#_c_513_n 0.0372099f $X=2.805 $Y=1.465
+ $X2=0 $Y2=0
cc_331 N_A_27_120#_c_394_n N_A_369_392#_c_514_n 0.00145506f $X=2.85 $Y=1.885
+ $X2=0 $Y2=0
cc_332 N_A_27_120#_c_386_n N_A_369_392#_c_505_n 0.00178439f $X=3.215 $Y=1.11
+ $X2=0 $Y2=0
cc_333 N_A_27_120#_c_383_n N_A_369_392#_c_508_n 2.00831e-19 $X=2.85 $Y=1.63
+ $X2=0 $Y2=0
cc_334 N_A_27_120#_c_384_n N_A_369_392#_c_508_n 0.00112116f $X=2.85 $Y=1.795
+ $X2=0 $Y2=0
cc_335 N_A_27_120#_c_385_n N_A_369_392#_c_508_n 8.35401e-19 $X=3.14 $Y=1.185
+ $X2=0 $Y2=0
cc_336 N_A_27_120#_c_392_n N_A_369_392#_c_508_n 0.0104417f $X=2.805 $Y=1.465
+ $X2=0 $Y2=0
cc_337 N_A_27_120#_c_383_n N_A_369_392#_c_509_n 0.00193199f $X=2.85 $Y=1.63
+ $X2=0 $Y2=0
cc_338 N_A_27_120#_c_386_n N_A_369_392#_c_509_n 0.0047803f $X=3.215 $Y=1.11
+ $X2=0 $Y2=0
cc_339 N_A_27_120#_c_390_n N_A_369_392#_c_509_n 0.00674121f $X=2.56 $Y=1.3 $X2=0
+ $Y2=0
cc_340 N_A_27_120#_c_392_n N_A_369_392#_c_509_n 0.00771809f $X=2.805 $Y=1.465
+ $X2=0 $Y2=0
cc_341 N_A_27_120#_c_394_n N_A_669_392#_c_719_n 0.00169621f $X=2.85 $Y=1.885
+ $X2=0 $Y2=0
cc_342 N_A_27_120#_c_395_n N_VPWR_c_774_n 0.0266809f $X=0.43 $Y=2.265 $X2=0
+ $Y2=0
cc_343 N_A_27_120#_c_397_n N_VPWR_c_774_n 0.00141767f $X=0.71 $Y=2.035 $X2=0
+ $Y2=0
cc_344 N_A_27_120#_c_394_n N_VPWR_c_775_n 0.00522314f $X=2.85 $Y=1.885 $X2=0
+ $Y2=0
cc_345 N_A_27_120#_c_395_n N_VPWR_c_779_n 0.0145938f $X=0.43 $Y=2.265 $X2=0
+ $Y2=0
cc_346 N_A_27_120#_c_394_n N_VPWR_c_786_n 0.0031609f $X=2.85 $Y=1.885 $X2=0
+ $Y2=0
cc_347 N_A_27_120#_c_394_n N_VPWR_c_773_n 0.0041189f $X=2.85 $Y=1.885 $X2=0
+ $Y2=0
cc_348 N_A_27_120#_c_395_n N_VPWR_c_773_n 0.0120466f $X=0.43 $Y=2.265 $X2=0
+ $Y2=0
cc_349 N_A_27_120#_c_387_n N_VGND_M1017_d 7.20017e-19 $X=0.71 $Y=1.95 $X2=-0.19
+ $Y2=-0.245
cc_350 N_A_27_120#_c_416_n N_VGND_M1017_d 0.00789213f $X=1.145 $Y=0.665
+ $X2=-0.19 $Y2=-0.245
cc_351 N_A_27_120#_c_391_n N_VGND_M1017_d 0.00822019f $X=0.795 $Y=0.855
+ $X2=-0.19 $Y2=-0.245
cc_352 N_A_27_120#_c_388_n N_VGND_M1009_d 6.47853e-19 $X=2.475 $Y=0.34 $X2=0
+ $Y2=0
cc_353 N_A_27_120#_c_390_n N_VGND_M1009_d 0.0113692f $X=2.56 $Y=1.3 $X2=0 $Y2=0
cc_354 N_A_27_120#_c_383_n N_VGND_c_886_n 0.0127456f $X=2.85 $Y=1.63 $X2=0 $Y2=0
cc_355 N_A_27_120#_c_386_n N_VGND_c_886_n 0.00940057f $X=3.215 $Y=1.11 $X2=0
+ $Y2=0
cc_356 N_A_27_120#_c_388_n N_VGND_c_886_n 0.0148948f $X=2.475 $Y=0.34 $X2=0
+ $Y2=0
cc_357 N_A_27_120#_c_390_n N_VGND_c_886_n 0.0481399f $X=2.56 $Y=1.3 $X2=0 $Y2=0
cc_358 N_A_27_120#_c_392_n N_VGND_c_886_n 0.00988174f $X=2.805 $Y=1.465 $X2=0
+ $Y2=0
cc_359 N_A_27_120#_c_391_n N_VGND_c_891_n 0.0110697f $X=0.795 $Y=0.855 $X2=0
+ $Y2=0
cc_360 N_A_27_120#_c_416_n N_VGND_c_892_n 0.00313112f $X=1.145 $Y=0.665 $X2=0
+ $Y2=0
cc_361 N_A_27_120#_c_388_n N_VGND_c_892_n 0.086417f $X=2.475 $Y=0.34 $X2=0 $Y2=0
cc_362 N_A_27_120#_c_389_n N_VGND_c_892_n 0.0118998f $X=1.315 $Y=0.34 $X2=0
+ $Y2=0
cc_363 N_A_27_120#_c_386_n N_VGND_c_893_n 0.00539704f $X=3.215 $Y=1.11 $X2=0
+ $Y2=0
cc_364 N_A_27_120#_c_389_n N_VGND_c_896_n 0.0120702f $X=1.315 $Y=0.34 $X2=0
+ $Y2=0
cc_365 N_A_27_120#_c_391_n N_VGND_c_896_n 0.0255806f $X=0.795 $Y=0.855 $X2=0
+ $Y2=0
cc_366 N_A_27_120#_c_386_n N_VGND_c_900_n 0.0052351f $X=3.215 $Y=1.11 $X2=0
+ $Y2=0
cc_367 N_A_27_120#_c_416_n N_VGND_c_900_n 0.00556468f $X=1.145 $Y=0.665 $X2=0
+ $Y2=0
cc_368 N_A_27_120#_c_388_n N_VGND_c_900_n 0.049532f $X=2.475 $Y=0.34 $X2=0 $Y2=0
cc_369 N_A_27_120#_c_389_n N_VGND_c_900_n 0.00655543f $X=1.315 $Y=0.34 $X2=0
+ $Y2=0
cc_370 N_A_27_120#_c_391_n N_VGND_c_900_n 0.0175471f $X=0.795 $Y=0.855 $X2=0
+ $Y2=0
cc_371 N_A_369_392#_c_507_n N_A_842_405#_M1005_g 0.0358316f $X=4.21 $Y=0.42
+ $X2=0 $Y2=0
cc_372 N_A_369_392#_c_506_n N_A_669_392#_M1001_d 0.00217732f $X=4.21 $Y=0.42
+ $X2=-0.19 $Y2=-0.245
cc_373 N_A_369_392#_c_508_n N_A_669_392#_M1018_d 0.00127066f $X=3.345 $Y=1.635
+ $X2=0 $Y2=0
cc_374 N_A_369_392#_c_506_n N_A_669_392#_c_707_n 0.00333692f $X=4.21 $Y=0.42
+ $X2=0 $Y2=0
cc_375 N_A_369_392#_c_510_n N_A_669_392#_c_707_n 0.00622744f $X=4.21 $Y=0.585
+ $X2=0 $Y2=0
cc_376 N_A_369_392#_c_506_n N_A_669_392#_c_708_n 0.032399f $X=4.21 $Y=0.42 $X2=0
+ $Y2=0
cc_377 N_A_369_392#_c_507_n N_A_669_392#_c_708_n 0.00386148f $X=4.21 $Y=0.42
+ $X2=0 $Y2=0
cc_378 N_A_369_392#_c_509_n N_A_669_392#_c_708_n 0.011037f $X=3.345 $Y=1.47
+ $X2=0 $Y2=0
cc_379 N_A_369_392#_c_510_n N_A_669_392#_c_708_n 0.0132252f $X=4.21 $Y=0.585
+ $X2=0 $Y2=0
cc_380 N_A_369_392#_c_503_n N_A_669_392#_c_719_n 0.010657f $X=3.27 $Y=1.885
+ $X2=0 $Y2=0
cc_381 N_A_369_392#_c_508_n N_A_669_392#_c_719_n 0.0106362f $X=3.345 $Y=1.635
+ $X2=0 $Y2=0
cc_382 N_A_369_392#_c_503_n N_A_669_392#_c_709_n 0.0049676f $X=3.27 $Y=1.885
+ $X2=0 $Y2=0
cc_383 N_A_369_392#_c_508_n N_A_669_392#_c_709_n 0.0382496f $X=3.345 $Y=1.635
+ $X2=0 $Y2=0
cc_384 N_A_369_392#_c_509_n N_A_669_392#_c_709_n 0.0277249f $X=3.345 $Y=1.47
+ $X2=0 $Y2=0
cc_385 N_A_369_392#_c_510_n N_A_669_392#_c_709_n 2.86089e-19 $X=4.21 $Y=0.585
+ $X2=0 $Y2=0
cc_386 N_A_369_392#_c_513_n N_VPWR_M1006_d 0.00653076f $X=3.18 $Y=1.885 $X2=0
+ $Y2=0
cc_387 N_A_369_392#_c_503_n N_VPWR_c_786_n 0.00278271f $X=3.27 $Y=1.885 $X2=0
+ $Y2=0
cc_388 N_A_369_392#_c_503_n N_VPWR_c_773_n 0.0035843f $X=3.27 $Y=1.885 $X2=0
+ $Y2=0
cc_389 N_A_369_392#_c_513_n A_585_392# 0.00464818f $X=3.18 $Y=1.885 $X2=-0.19
+ $Y2=-0.245
cc_390 N_A_369_392#_c_505_n N_VGND_c_886_n 0.0189626f $X=3.485 $Y=0.42 $X2=0
+ $Y2=0
cc_391 N_A_369_392#_c_509_n N_VGND_c_886_n 0.0183503f $X=3.345 $Y=1.47 $X2=0
+ $Y2=0
cc_392 N_A_369_392#_c_506_n N_VGND_c_887_n 0.0133466f $X=4.21 $Y=0.42 $X2=0
+ $Y2=0
cc_393 N_A_369_392#_c_507_n N_VGND_c_887_n 0.00191229f $X=4.21 $Y=0.42 $X2=0
+ $Y2=0
cc_394 N_A_369_392#_c_505_n N_VGND_c_893_n 0.0121867f $X=3.485 $Y=0.42 $X2=0
+ $Y2=0
cc_395 N_A_369_392#_c_506_n N_VGND_c_893_n 0.0589947f $X=4.21 $Y=0.42 $X2=0
+ $Y2=0
cc_396 N_A_369_392#_c_507_n N_VGND_c_893_n 0.00783549f $X=4.21 $Y=0.42 $X2=0
+ $Y2=0
cc_397 N_A_369_392#_c_505_n N_VGND_c_900_n 0.00660921f $X=3.485 $Y=0.42 $X2=0
+ $Y2=0
cc_398 N_A_369_392#_c_506_n N_VGND_c_900_n 0.0337644f $X=4.21 $Y=0.42 $X2=0
+ $Y2=0
cc_399 N_A_369_392#_c_507_n N_VGND_c_900_n 0.011167f $X=4.21 $Y=0.42 $X2=0 $Y2=0
cc_400 N_A_369_392#_c_509_n A_658_79# 0.00191955f $X=3.345 $Y=1.47 $X2=-0.19
+ $Y2=-0.245
cc_401 N_A_842_405#_M1005_g N_A_669_392#_c_705_n 0.0435149f $X=4.69 $Y=0.905
+ $X2=0 $Y2=0
cc_402 N_A_842_405#_c_610_n N_A_669_392#_c_705_n 0.0182244f $X=6.11 $Y=1.46
+ $X2=0 $Y2=0
cc_403 N_A_842_405#_c_621_n N_A_669_392#_c_705_n 0.0185734f $X=5.25 $Y=2.19
+ $X2=0 $Y2=0
cc_404 N_A_842_405#_c_623_n N_A_669_392#_c_705_n 0.00684283f $X=5.415 $Y=2.355
+ $X2=0 $Y2=0
cc_405 N_A_842_405#_c_624_n N_A_669_392#_c_705_n 0.0157975f $X=5.415 $Y=2.79
+ $X2=0 $Y2=0
cc_406 N_A_842_405#_c_625_n N_A_669_392#_c_705_n 0.00548739f $X=5.59 $Y=1.795
+ $X2=0 $Y2=0
cc_407 N_A_842_405#_c_615_n N_A_669_392#_c_705_n 0.00127754f $X=5.59 $Y=1.46
+ $X2=0 $Y2=0
cc_408 N_A_842_405#_M1005_g N_A_669_392#_M1014_g 0.0137357f $X=4.69 $Y=0.905
+ $X2=0 $Y2=0
cc_409 N_A_842_405#_c_612_n N_A_669_392#_M1014_g 0.00180139f $X=5.415 $Y=0.52
+ $X2=0 $Y2=0
cc_410 N_A_842_405#_c_613_n N_A_669_392#_M1014_g 0.00353515f $X=5.59 $Y=1.295
+ $X2=0 $Y2=0
cc_411 N_A_842_405#_M1005_g N_A_669_392#_c_707_n 0.0251514f $X=4.69 $Y=0.905
+ $X2=0 $Y2=0
cc_412 N_A_842_405#_c_610_n N_A_669_392#_c_707_n 3.60437e-19 $X=6.11 $Y=1.46
+ $X2=0 $Y2=0
cc_413 N_A_842_405#_c_621_n N_A_669_392#_c_707_n 0.00915012f $X=5.25 $Y=2.19
+ $X2=0 $Y2=0
cc_414 N_A_842_405#_c_623_n N_A_669_392#_c_707_n 0.00713557f $X=5.415 $Y=2.355
+ $X2=0 $Y2=0
cc_415 N_A_842_405#_c_613_n N_A_669_392#_c_707_n 0.0069888f $X=5.59 $Y=1.295
+ $X2=0 $Y2=0
cc_416 N_A_842_405#_c_615_n N_A_669_392#_c_707_n 0.0281337f $X=5.59 $Y=1.46
+ $X2=0 $Y2=0
cc_417 N_A_842_405#_M1005_g N_A_669_392#_c_708_n 0.00134353f $X=4.69 $Y=0.905
+ $X2=0 $Y2=0
cc_418 N_A_842_405#_c_621_n N_VPWR_M1013_d 0.00953826f $X=5.25 $Y=2.19 $X2=0
+ $Y2=0
cc_419 N_A_842_405#_c_618_n N_VPWR_c_776_n 0.0116432f $X=6.2 $Y=1.765 $X2=0
+ $Y2=0
cc_420 N_A_842_405#_c_610_n N_VPWR_c_776_n 0.00489956f $X=6.11 $Y=1.46 $X2=0
+ $Y2=0
cc_421 N_A_842_405#_c_623_n N_VPWR_c_776_n 0.0355478f $X=5.415 $Y=2.355 $X2=0
+ $Y2=0
cc_422 N_A_842_405#_c_624_n N_VPWR_c_776_n 0.0345916f $X=5.415 $Y=2.79 $X2=0
+ $Y2=0
cc_423 N_A_842_405#_c_662_p N_VPWR_c_776_n 0.0162042f $X=6.08 $Y=1.46 $X2=0
+ $Y2=0
cc_424 N_A_842_405#_c_619_n N_VPWR_c_778_n 0.0117699f $X=6.695 $Y=1.765 $X2=0
+ $Y2=0
cc_425 N_A_842_405#_c_624_n N_VPWR_c_781_n 0.0132586f $X=5.415 $Y=2.79 $X2=0
+ $Y2=0
cc_426 N_A_842_405#_c_618_n N_VPWR_c_784_n 0.00446702f $X=6.2 $Y=1.765 $X2=0
+ $Y2=0
cc_427 N_A_842_405#_c_619_n N_VPWR_c_784_n 0.00446702f $X=6.695 $Y=1.765 $X2=0
+ $Y2=0
cc_428 N_A_842_405#_c_616_n N_VPWR_c_786_n 0.00502391f $X=4.3 $Y=2.44 $X2=0
+ $Y2=0
cc_429 N_A_842_405#_c_616_n N_VPWR_c_787_n 0.00779314f $X=4.3 $Y=2.44 $X2=0
+ $Y2=0
cc_430 N_A_842_405#_c_621_n N_VPWR_c_787_n 0.0393049f $X=5.25 $Y=2.19 $X2=0
+ $Y2=0
cc_431 N_A_842_405#_c_622_n N_VPWR_c_787_n 0.00862558f $X=4.525 $Y=2.19 $X2=0
+ $Y2=0
cc_432 N_A_842_405#_c_624_n N_VPWR_c_787_n 0.0132969f $X=5.415 $Y=2.79 $X2=0
+ $Y2=0
cc_433 N_A_842_405#_c_616_n N_VPWR_c_773_n 0.00484068f $X=4.3 $Y=2.44 $X2=0
+ $Y2=0
cc_434 N_A_842_405#_c_618_n N_VPWR_c_773_n 0.0086399f $X=6.2 $Y=1.765 $X2=0
+ $Y2=0
cc_435 N_A_842_405#_c_619_n N_VPWR_c_773_n 0.00862683f $X=6.695 $Y=1.765 $X2=0
+ $Y2=0
cc_436 N_A_842_405#_c_624_n N_VPWR_c_773_n 0.0119178f $X=5.415 $Y=2.79 $X2=0
+ $Y2=0
cc_437 N_A_842_405#_M1000_g N_Q_c_861_n 5.5543e-19 $X=6.19 $Y=0.74 $X2=0 $Y2=0
cc_438 N_A_842_405#_M1012_g N_Q_c_861_n 0.00487958f $X=6.68 $Y=0.74 $X2=0 $Y2=0
cc_439 N_A_842_405#_c_611_n N_Q_c_862_n 0.00266648f $X=6.68 $Y=1.53 $X2=0 $Y2=0
cc_440 N_A_842_405#_c_618_n Q 0.0199584f $X=6.2 $Y=1.765 $X2=0 $Y2=0
cc_441 N_A_842_405#_c_619_n Q 0.0199584f $X=6.695 $Y=1.765 $X2=0 $Y2=0
cc_442 N_A_842_405#_c_611_n Q 0.00419557f $X=6.68 $Y=1.53 $X2=0 $Y2=0
cc_443 N_A_842_405#_M1000_g N_Q_c_863_n 0.00369108f $X=6.19 $Y=0.74 $X2=0 $Y2=0
cc_444 N_A_842_405#_c_618_n N_Q_c_863_n 0.00195842f $X=6.2 $Y=1.765 $X2=0 $Y2=0
cc_445 N_A_842_405#_c_619_n N_Q_c_863_n 0.00183496f $X=6.695 $Y=1.765 $X2=0
+ $Y2=0
cc_446 N_A_842_405#_c_611_n N_Q_c_863_n 0.0358515f $X=6.68 $Y=1.53 $X2=0 $Y2=0
cc_447 N_A_842_405#_c_662_p N_Q_c_863_n 0.0249855f $X=6.08 $Y=1.46 $X2=0 $Y2=0
cc_448 N_A_842_405#_M1005_g N_VGND_c_887_n 0.00480566f $X=4.69 $Y=0.905 $X2=0
+ $Y2=0
cc_449 N_A_842_405#_c_612_n N_VGND_c_887_n 0.0229496f $X=5.415 $Y=0.52 $X2=0
+ $Y2=0
cc_450 N_A_842_405#_M1000_g N_VGND_c_888_n 0.014912f $X=6.19 $Y=0.74 $X2=0 $Y2=0
cc_451 N_A_842_405#_M1012_g N_VGND_c_888_n 5.38476e-19 $X=6.68 $Y=0.74 $X2=0
+ $Y2=0
cc_452 N_A_842_405#_c_610_n N_VGND_c_888_n 0.00625479f $X=6.11 $Y=1.46 $X2=0
+ $Y2=0
cc_453 N_A_842_405#_c_612_n N_VGND_c_888_n 0.0346502f $X=5.415 $Y=0.52 $X2=0
+ $Y2=0
cc_454 N_A_842_405#_c_662_p N_VGND_c_888_n 0.0245638f $X=6.08 $Y=1.46 $X2=0
+ $Y2=0
cc_455 N_A_842_405#_c_614_n N_VGND_c_888_n 0.0138526f $X=5.502 $Y=1.125 $X2=0
+ $Y2=0
cc_456 N_A_842_405#_M1012_g N_VGND_c_890_n 0.00553267f $X=6.68 $Y=0.74 $X2=0
+ $Y2=0
cc_457 N_A_842_405#_c_611_n N_VGND_c_890_n 0.00114951f $X=6.68 $Y=1.53 $X2=0
+ $Y2=0
cc_458 N_A_842_405#_M1005_g N_VGND_c_893_n 0.00380268f $X=4.69 $Y=0.905 $X2=0
+ $Y2=0
cc_459 N_A_842_405#_c_612_n N_VGND_c_894_n 0.0108483f $X=5.415 $Y=0.52 $X2=0
+ $Y2=0
cc_460 N_A_842_405#_M1000_g N_VGND_c_895_n 0.00383152f $X=6.19 $Y=0.74 $X2=0
+ $Y2=0
cc_461 N_A_842_405#_M1012_g N_VGND_c_895_n 0.00460063f $X=6.68 $Y=0.74 $X2=0
+ $Y2=0
cc_462 N_A_842_405#_M1005_g N_VGND_c_900_n 0.0045051f $X=4.69 $Y=0.905 $X2=0
+ $Y2=0
cc_463 N_A_842_405#_M1000_g N_VGND_c_900_n 0.00758109f $X=6.19 $Y=0.74 $X2=0
+ $Y2=0
cc_464 N_A_842_405#_M1012_g N_VGND_c_900_n 0.0091141f $X=6.68 $Y=0.74 $X2=0
+ $Y2=0
cc_465 N_A_842_405#_c_612_n N_VGND_c_900_n 0.00913189f $X=5.415 $Y=0.52 $X2=0
+ $Y2=0
cc_466 N_A_669_392#_c_705_n N_VPWR_c_776_n 0.0044733f $X=5.19 $Y=1.74 $X2=0
+ $Y2=0
cc_467 N_A_669_392#_c_705_n N_VPWR_c_781_n 0.00544739f $X=5.19 $Y=1.74 $X2=0
+ $Y2=0
cc_468 N_A_669_392#_c_705_n N_VPWR_c_787_n 0.00570914f $X=5.19 $Y=1.74 $X2=0
+ $Y2=0
cc_469 N_A_669_392#_c_705_n N_VPWR_c_773_n 0.00537853f $X=5.19 $Y=1.74 $X2=0
+ $Y2=0
cc_470 N_A_669_392#_c_705_n N_VGND_c_887_n 5.31937e-19 $X=5.19 $Y=1.74 $X2=0
+ $Y2=0
cc_471 N_A_669_392#_M1014_g N_VGND_c_887_n 0.014975f $X=5.2 $Y=0.745 $X2=0 $Y2=0
cc_472 N_A_669_392#_c_707_n N_VGND_c_887_n 0.0253469f $X=4.99 $Y=1.23 $X2=0
+ $Y2=0
cc_473 N_A_669_392#_M1014_g N_VGND_c_888_n 0.0039491f $X=5.2 $Y=0.745 $X2=0
+ $Y2=0
cc_474 N_A_669_392#_M1014_g N_VGND_c_894_n 0.00379792f $X=5.2 $Y=0.745 $X2=0
+ $Y2=0
cc_475 N_A_669_392#_M1014_g N_VGND_c_900_n 0.00457201f $X=5.2 $Y=0.745 $X2=0
+ $Y2=0
cc_476 N_VPWR_c_776_n Q 0.0648992f $X=5.975 $Y=1.985 $X2=0 $Y2=0
cc_477 N_VPWR_c_778_n Q 0.0656374f $X=6.92 $Y=1.985 $X2=0 $Y2=0
cc_478 N_VPWR_c_784_n Q 0.0100771f $X=6.835 $Y=3.33 $X2=0 $Y2=0
cc_479 N_VPWR_c_773_n Q 0.0128515f $X=6.96 $Y=3.33 $X2=0 $Y2=0
cc_480 N_VPWR_c_776_n N_Q_c_863_n 0.00433555f $X=5.975 $Y=1.985 $X2=0 $Y2=0
cc_481 N_VPWR_c_778_n N_Q_c_863_n 0.00347086f $X=6.92 $Y=1.985 $X2=0 $Y2=0
cc_482 N_Q_c_861_n N_VGND_c_888_n 0.0285797f $X=6.41 $Y=0.515 $X2=0 $Y2=0
cc_483 N_Q_c_861_n N_VGND_c_890_n 0.0313502f $X=6.41 $Y=0.515 $X2=0 $Y2=0
cc_484 N_Q_c_861_n N_VGND_c_895_n 0.0117353f $X=6.41 $Y=0.515 $X2=0 $Y2=0
cc_485 N_Q_c_861_n N_VGND_c_900_n 0.00971347f $X=6.41 $Y=0.515 $X2=0 $Y2=0
