* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hs__dfbbn_1 CLK_N D RESET_B SET_B VGND VNB VPB VPWR Q Q_N
X0 VPWR a_27_74# a_200_74# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X1 a_595_119# a_200_74# a_311_119# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X2 a_1534_446# a_1349_114# a_1818_76# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X3 a_311_119# D VPWR VPB sky130_fd_pr__pfet_01v8 w=420000u l=150000u
X4 a_1349_114# a_27_74# a_1483_508# VPB sky130_fd_pr__pfet_01v8 w=420000u l=150000u
X5 VGND a_1534_446# Q_N VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X6 VPWR a_474_405# a_537_503# VPB sky130_fd_pr__pfet_01v8 w=420000u l=150000u
X7 VPWR a_1534_446# Q_N VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X8 a_1611_140# a_1534_446# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X9 a_595_119# a_27_74# a_311_119# VPB sky130_fd_pr__pfet_01v8 w=420000u l=150000u
X10 a_1483_508# a_1534_446# VPWR VPB sky130_fd_pr__pfet_01v8 w=420000u l=150000u
X11 VGND a_27_74# a_200_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X12 a_1917_392# a_1349_114# a_1534_446# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=150000u
X13 a_537_503# a_200_74# a_595_119# VPB sky130_fd_pr__pfet_01v8 w=420000u l=150000u
X14 a_978_357# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8 w=640000u l=150000u
X15 a_27_74# CLK_N VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X16 VPWR a_2412_410# Q VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X17 VPWR a_474_405# a_1297_424# VPB sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X18 a_311_119# D VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X19 a_474_405# a_978_357# a_867_119# VNB sky130_fd_pr__nfet_01v8_lvt w=550000u l=150000u
X20 a_867_119# a_595_119# a_474_405# VNB sky130_fd_pr__nfet_01v8_lvt w=550000u l=150000u
X21 VPWR a_978_357# a_1917_392# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=150000u
X22 a_1254_119# a_27_74# a_1349_114# VNB sky130_fd_pr__nfet_01v8_lvt w=550000u l=150000u
X23 VGND SET_B a_1818_76# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X24 a_978_357# RESET_B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X25 a_1297_424# a_200_74# a_1349_114# VPB sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X26 a_2412_410# a_1534_446# VPWR VPB sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X27 a_867_119# SET_B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=550000u l=150000u
X28 a_933_424# a_978_357# VPWR VPB sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X29 VGND a_2412_410# Q VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X30 VGND a_474_405# a_523_119# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X31 a_523_119# a_27_74# a_595_119# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X32 a_1534_446# SET_B VPWR VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=150000u
X33 a_1349_114# a_200_74# a_1611_140# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X34 VPWR SET_B a_474_405# VPB sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X35 a_1818_76# a_978_357# a_1534_446# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X36 a_2412_410# a_1534_446# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X37 a_27_74# CLK_N VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X38 VGND a_474_405# a_1254_119# VNB sky130_fd_pr__nfet_01v8_lvt w=550000u l=150000u
X39 a_474_405# a_595_119# a_933_424# VPB sky130_fd_pr__pfet_01v8 w=840000u l=150000u
.ends
