* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hs__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
M1000 a_527_368# A3 a_443_368# VPB pshort w=1.12e+06u l=150000u
+  ad=4.704e+11p pd=3.08e+06u as=3.024e+11p ps=2.78e+06u
M1001 VPWR A1 a_641_368# VPB pshort w=1.12e+06u l=150000u
+  ad=1.4016e+12p pd=7.2e+06u as=4.704e+11p ps=3.08e+06u
M1002 a_641_368# A2 a_527_368# VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1003 VGND A4 a_326_74# VNB nlowvt w=640000u l=150000u
+  ad=8.899e+11p pd=6.71e+06u as=6.24e+11p ps=5.79e+06u
M1004 a_326_74# B1 a_83_270# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=1.824e+11p ps=1.85e+06u
M1005 VPWR a_83_270# X VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=3.304e+11p ps=2.83e+06u
M1006 a_83_270# B1 VPWR VPB pshort w=840000u l=150000u
+  ad=4.0165e+11p pd=3.01e+06u as=0p ps=0u
M1007 VGND A2 a_326_74# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_443_368# A4 a_83_270# VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_326_74# A1 VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VGND a_83_270# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1011 a_326_74# A3 VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
