# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_hs__sdfrtp_2
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_hs__sdfrtp_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  14.40000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.565000 0.810000 2.100000 1.265000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.543200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 13.525000 0.350000 13.855000 1.410000 ;
        RECT 13.525000 1.410000 13.785000 2.980000 ;
    END
  END Q
  PIN RESET_B
    ANTENNAGATEAREA  0.411000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT  3.785000 1.830000  4.165000 2.160000 ;
        RECT  7.825000 1.795000  8.515000 2.150000 ;
        RECT 11.110000 1.920000 11.440000 2.220000 ;
      LAYER mcon ;
        RECT  3.995000 1.950000  4.165000 2.120000 ;
        RECT  8.315000 1.950000  8.485000 2.120000 ;
        RECT 11.195000 1.950000 11.365000 2.120000 ;
      LAYER met1 ;
        RECT  3.935000 1.920000  4.225000 1.965000 ;
        RECT  3.935000 1.965000 11.425000 2.105000 ;
        RECT  3.935000 2.105000  4.225000 2.150000 ;
        RECT  8.255000 1.920000  8.545000 1.965000 ;
        RECT  8.255000 2.105000  8.545000 2.150000 ;
        RECT 11.135000 1.920000 11.425000 1.965000 ;
        RECT 11.135000 2.105000 11.425000 2.150000 ;
    END
  END RESET_B
  PIN SCD
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.945000 1.480000 3.275000 2.150000 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605000 1.490000 2.705000 1.660000 ;
        RECT 0.605000 1.660000 1.795000 1.835000 ;
        RECT 2.375000 1.260000 2.705000 1.490000 ;
    END
  END SCE
  PIN CLK
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 3.965000 1.180000 4.195000 1.260000 ;
        RECT 3.965000 1.260000 4.645000 1.590000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT  0.000000 -0.085000 14.400000 0.085000 ;
        RECT  0.545000  0.085000  0.875000 0.765000 ;
        RECT  3.715000  0.085000  4.045000 0.845000 ;
        RECT  4.740000  0.085000  5.070000 0.750000 ;
        RECT  7.605000  0.085000  8.080000 0.410000 ;
        RECT 10.755000  0.085000 11.085000 0.810000 ;
        RECT 12.105000  0.085000 12.435000 0.600000 ;
        RECT 13.095000  0.085000 13.345000 1.130000 ;
        RECT 14.035000  0.085000 14.285000 1.130000 ;
      LAYER mcon ;
        RECT  0.155000 -0.085000  0.325000 0.085000 ;
        RECT  0.635000 -0.085000  0.805000 0.085000 ;
        RECT  1.115000 -0.085000  1.285000 0.085000 ;
        RECT  1.595000 -0.085000  1.765000 0.085000 ;
        RECT  2.075000 -0.085000  2.245000 0.085000 ;
        RECT  2.555000 -0.085000  2.725000 0.085000 ;
        RECT  3.035000 -0.085000  3.205000 0.085000 ;
        RECT  3.515000 -0.085000  3.685000 0.085000 ;
        RECT  3.995000 -0.085000  4.165000 0.085000 ;
        RECT  4.475000 -0.085000  4.645000 0.085000 ;
        RECT  4.955000 -0.085000  5.125000 0.085000 ;
        RECT  5.435000 -0.085000  5.605000 0.085000 ;
        RECT  5.915000 -0.085000  6.085000 0.085000 ;
        RECT  6.395000 -0.085000  6.565000 0.085000 ;
        RECT  6.875000 -0.085000  7.045000 0.085000 ;
        RECT  7.355000 -0.085000  7.525000 0.085000 ;
        RECT  7.835000 -0.085000  8.005000 0.085000 ;
        RECT  8.315000 -0.085000  8.485000 0.085000 ;
        RECT  8.795000 -0.085000  8.965000 0.085000 ;
        RECT  9.275000 -0.085000  9.445000 0.085000 ;
        RECT  9.755000 -0.085000  9.925000 0.085000 ;
        RECT 10.235000 -0.085000 10.405000 0.085000 ;
        RECT 10.715000 -0.085000 10.885000 0.085000 ;
        RECT 11.195000 -0.085000 11.365000 0.085000 ;
        RECT 11.675000 -0.085000 11.845000 0.085000 ;
        RECT 12.155000 -0.085000 12.325000 0.085000 ;
        RECT 12.635000 -0.085000 12.805000 0.085000 ;
        RECT 13.115000 -0.085000 13.285000 0.085000 ;
        RECT 13.595000 -0.085000 13.765000 0.085000 ;
        RECT 14.075000 -0.085000 14.245000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.245000 14.400000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT  0.000000 3.245000 14.400000 3.415000 ;
        RECT  0.615000 2.345000  1.565000 3.245000 ;
        RECT  3.095000 2.685000  3.425000 3.245000 ;
        RECT  4.705000 2.730000  5.035000 3.245000 ;
        RECT  7.150000 2.660000  7.485000 3.245000 ;
        RECT  8.250000 2.320000  8.580000 3.245000 ;
        RECT 10.560000 2.730000 11.240000 3.245000 ;
        RECT 11.945000 1.940000 12.275000 3.245000 ;
        RECT 13.005000 1.820000 13.335000 3.245000 ;
        RECT 13.955000 1.820000 14.285000 3.245000 ;
      LAYER mcon ;
        RECT  0.155000 3.245000  0.325000 3.415000 ;
        RECT  0.635000 3.245000  0.805000 3.415000 ;
        RECT  1.115000 3.245000  1.285000 3.415000 ;
        RECT  1.595000 3.245000  1.765000 3.415000 ;
        RECT  2.075000 3.245000  2.245000 3.415000 ;
        RECT  2.555000 3.245000  2.725000 3.415000 ;
        RECT  3.035000 3.245000  3.205000 3.415000 ;
        RECT  3.515000 3.245000  3.685000 3.415000 ;
        RECT  3.995000 3.245000  4.165000 3.415000 ;
        RECT  4.475000 3.245000  4.645000 3.415000 ;
        RECT  4.955000 3.245000  5.125000 3.415000 ;
        RECT  5.435000 3.245000  5.605000 3.415000 ;
        RECT  5.915000 3.245000  6.085000 3.415000 ;
        RECT  6.395000 3.245000  6.565000 3.415000 ;
        RECT  6.875000 3.245000  7.045000 3.415000 ;
        RECT  7.355000 3.245000  7.525000 3.415000 ;
        RECT  7.835000 3.245000  8.005000 3.415000 ;
        RECT  8.315000 3.245000  8.485000 3.415000 ;
        RECT  8.795000 3.245000  8.965000 3.415000 ;
        RECT  9.275000 3.245000  9.445000 3.415000 ;
        RECT  9.755000 3.245000  9.925000 3.415000 ;
        RECT 10.235000 3.245000 10.405000 3.415000 ;
        RECT 10.715000 3.245000 10.885000 3.415000 ;
        RECT 11.195000 3.245000 11.365000 3.415000 ;
        RECT 11.675000 3.245000 11.845000 3.415000 ;
        RECT 12.155000 3.245000 12.325000 3.415000 ;
        RECT 12.635000 3.245000 12.805000 3.415000 ;
        RECT 13.115000 3.245000 13.285000 3.415000 ;
        RECT 13.595000 3.245000 13.765000 3.415000 ;
        RECT 14.075000 3.245000 14.245000 3.415000 ;
      LAYER met1 ;
        RECT 0.000000 3.085000 14.400000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.115000 0.350000  0.365000 0.935000 ;
      RECT  0.115000 0.935000  1.140000 1.265000 ;
      RECT  0.115000 1.265000  0.285000 2.005000 ;
      RECT  0.115000 2.005000  2.705000 2.175000 ;
      RECT  0.115000 2.175000  0.445000 2.980000 ;
      RECT  1.105000 0.255000  3.545000 0.425000 ;
      RECT  1.105000 0.425000  1.435000 0.640000 ;
      RECT  2.105000 2.345000  3.995000 2.390000 ;
      RECT  2.105000 2.390000  5.995000 2.515000 ;
      RECT  2.105000 2.515000  2.435000 2.980000 ;
      RECT  2.270000 0.595000  3.045000 0.845000 ;
      RECT  2.375000 1.830000  2.705000 2.005000 ;
      RECT  2.875000 0.845000  3.045000 1.140000 ;
      RECT  2.875000 1.140000  3.615000 1.310000 ;
      RECT  3.215000 0.425000  3.545000 0.845000 ;
      RECT  3.445000 1.310000  3.615000 2.330000 ;
      RECT  3.445000 2.330000  3.995000 2.345000 ;
      RECT  3.615000 2.515000  5.995000 2.560000 ;
      RECT  3.615000 2.560000  3.995000 2.980000 ;
      RECT  4.335000 1.820000  4.985000 1.990000 ;
      RECT  4.335000 1.990000  4.585000 2.220000 ;
      RECT  4.390000 0.350000  4.560000 0.920000 ;
      RECT  4.390000 0.920000  4.985000 1.090000 ;
      RECT  4.815000 1.090000  4.985000 1.295000 ;
      RECT  4.815000 1.295000  5.305000 1.625000 ;
      RECT  4.815000 1.625000  4.985000 1.820000 ;
      RECT  5.155000 1.795000  6.190000 1.965000 ;
      RECT  5.155000 1.965000  5.485000 2.220000 ;
      RECT  5.240000 0.330000  7.210000 0.500000 ;
      RECT  5.240000 0.500000  5.645000 1.125000 ;
      RECT  5.475000 1.125000  5.645000 1.635000 ;
      RECT  5.475000 1.635000  6.190000 1.795000 ;
      RECT  5.745000 2.135000  6.530000 2.305000 ;
      RECT  5.745000 2.305000  5.995000 2.390000 ;
      RECT  5.745000 2.560000  5.995000 2.725000 ;
      RECT  5.815000 0.670000  6.145000 1.295000 ;
      RECT  5.815000 1.295000  6.530000 1.465000 ;
      RECT  6.195000 2.475000  8.020000 2.490000 ;
      RECT  6.195000 2.490000  6.870000 2.725000 ;
      RECT  6.315000 0.670000  6.645000 0.955000 ;
      RECT  6.315000 0.955000  6.870000 1.125000 ;
      RECT  6.360000 1.465000  6.530000 2.135000 ;
      RECT  6.700000 1.125000  6.870000 2.320000 ;
      RECT  6.700000 2.320000  8.020000 2.475000 ;
      RECT  7.040000 0.500000  7.210000 0.580000 ;
      RECT  7.040000 0.580000  8.420000 0.750000 ;
      RECT  7.040000 0.920000  8.920000 1.090000 ;
      RECT  7.040000 1.090000  7.315000 2.075000 ;
      RECT  7.485000 1.260000  8.420000 1.575000 ;
      RECT  7.485000 1.575000  7.655000 2.320000 ;
      RECT  7.690000 2.490000  8.020000 2.725000 ;
      RECT  8.250000 0.255000  9.260000 0.425000 ;
      RECT  8.250000 0.425000  8.420000 0.580000 ;
      RECT  8.590000 0.595000  8.920000 0.920000 ;
      RECT  8.590000 1.090000  8.920000 1.130000 ;
      RECT  8.750000 1.130000  8.920000 1.715000 ;
      RECT  8.750000 1.715000  9.115000 2.755000 ;
      RECT  9.090000 0.425000  9.260000 1.005000 ;
      RECT  9.090000 1.005000 10.050000 1.335000 ;
      RECT  9.320000 1.840000  9.600000 2.520000 ;
      RECT  9.320000 2.520000 10.390000 2.850000 ;
      RECT  9.430000 0.480000 10.390000 0.810000 ;
      RECT  9.785000 1.335000 10.050000 2.330000 ;
      RECT 10.220000 0.810000 10.390000 1.030000 ;
      RECT 10.220000 1.030000 11.190000 1.110000 ;
      RECT 10.220000 1.110000 11.890000 1.200000 ;
      RECT 10.220000 1.200000 10.390000 2.520000 ;
      RECT 10.560000 1.370000 10.850000 1.580000 ;
      RECT 10.560000 1.580000 12.230000 1.750000 ;
      RECT 10.560000 1.750000 10.850000 2.390000 ;
      RECT 10.560000 2.390000 11.740000 2.560000 ;
      RECT 11.020000 1.200000 11.890000 1.410000 ;
      RECT 11.410000 2.560000 11.740000 2.980000 ;
      RECT 11.545000 0.350000 11.875000 0.770000 ;
      RECT 11.545000 0.770000 12.230000 0.940000 ;
      RECT 12.060000 0.940000 12.230000 1.580000 ;
      RECT 12.445000 1.940000 12.775000 2.980000 ;
      RECT 12.605000 0.350000 12.865000 1.300000 ;
      RECT 12.605000 1.300000 13.355000 1.630000 ;
      RECT 12.605000 1.630000 12.775000 1.940000 ;
  END
END sky130_fd_sc_hs__sdfrtp_2
