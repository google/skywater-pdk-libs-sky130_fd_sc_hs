* File: sky130_fd_sc_hs__or2_4.pxi.spice
* Created: Thu Aug 27 21:05:14 2020
* 
x_PM_SKY130_FD_SC_HS__OR2_4%A_83_260# N_A_83_260#_M1001_d N_A_83_260#_M1009_d
+ N_A_83_260#_M1002_g N_A_83_260#_c_87_n N_A_83_260#_M1004_g N_A_83_260#_M1003_g
+ N_A_83_260#_c_88_n N_A_83_260#_M1005_g N_A_83_260#_M1012_g N_A_83_260#_c_89_n
+ N_A_83_260#_M1006_g N_A_83_260#_c_90_n N_A_83_260#_M1008_g N_A_83_260#_M1013_g
+ N_A_83_260#_c_155_p N_A_83_260#_c_80_n N_A_83_260#_c_81_n N_A_83_260#_c_82_n
+ N_A_83_260#_c_105_p N_A_83_260#_c_91_n N_A_83_260#_c_110_p N_A_83_260#_c_83_n
+ N_A_83_260#_c_84_n N_A_83_260#_c_85_n N_A_83_260#_c_86_n
+ PM_SKY130_FD_SC_HS__OR2_4%A_83_260#
x_PM_SKY130_FD_SC_HS__OR2_4%A N_A_M1001_g N_A_c_212_n N_A_M1007_g N_A_c_213_n
+ N_A_M1010_g N_A_c_234_n N_A_c_214_n A PM_SKY130_FD_SC_HS__OR2_4%A
x_PM_SKY130_FD_SC_HS__OR2_4%B N_B_c_289_n N_B_M1009_g N_B_M1000_g N_B_c_290_n
+ N_B_M1011_g B N_B_c_288_n PM_SKY130_FD_SC_HS__OR2_4%B
x_PM_SKY130_FD_SC_HS__OR2_4%VPWR N_VPWR_M1004_d N_VPWR_M1005_d N_VPWR_M1008_d
+ N_VPWR_M1010_s N_VPWR_c_333_n N_VPWR_c_334_n N_VPWR_c_335_n N_VPWR_c_336_n
+ N_VPWR_c_337_n N_VPWR_c_338_n N_VPWR_c_339_n N_VPWR_c_340_n VPWR
+ N_VPWR_c_341_n N_VPWR_c_342_n N_VPWR_c_343_n N_VPWR_c_332_n
+ PM_SKY130_FD_SC_HS__OR2_4%VPWR
x_PM_SKY130_FD_SC_HS__OR2_4%X N_X_M1002_d N_X_M1012_d N_X_M1004_s N_X_M1006_s
+ N_X_c_394_n N_X_c_395_n N_X_c_401_n N_X_c_402_n N_X_c_396_n N_X_c_403_n
+ N_X_c_397_n N_X_c_404_n N_X_c_398_n N_X_c_405_n N_X_c_399_n N_X_c_406_n X X
+ PM_SKY130_FD_SC_HS__OR2_4%X
x_PM_SKY130_FD_SC_HS__OR2_4%A_493_388# N_A_493_388#_M1007_d N_A_493_388#_M1011_s
+ N_A_493_388#_c_478_n N_A_493_388#_c_474_n N_A_493_388#_c_475_n
+ N_A_493_388#_c_476_n PM_SKY130_FD_SC_HS__OR2_4%A_493_388#
x_PM_SKY130_FD_SC_HS__OR2_4%VGND N_VGND_M1002_s N_VGND_M1003_s N_VGND_M1013_s
+ N_VGND_M1000_d N_VGND_c_506_n N_VGND_c_507_n N_VGND_c_508_n N_VGND_c_509_n
+ N_VGND_c_510_n N_VGND_c_511_n VGND N_VGND_c_512_n N_VGND_c_513_n
+ N_VGND_c_514_n N_VGND_c_515_n N_VGND_c_516_n PM_SKY130_FD_SC_HS__OR2_4%VGND
cc_1 VNB N_A_83_260#_M1002_g 0.0224607f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_2 VNB N_A_83_260#_M1003_g 0.0203442f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=0.74
cc_3 VNB N_A_83_260#_M1012_g 0.02196f $X=-0.19 $Y=-0.245 $X2=1.355 $Y2=0.74
cc_4 VNB N_A_83_260#_M1013_g 0.0216596f $X=-0.19 $Y=-0.245 $X2=1.87 $Y2=0.74
cc_5 VNB N_A_83_260#_c_80_n 0.00648005f $X=-0.19 $Y=-0.245 $X2=2.42 $Y2=1.095
cc_6 VNB N_A_83_260#_c_81_n 0.0028029f $X=-0.19 $Y=-0.245 $X2=2.585 $Y2=0.515
cc_7 VNB N_A_83_260#_c_82_n 0.0303098f $X=-0.19 $Y=-0.245 $X2=4.065 $Y2=1.095
cc_8 VNB N_A_83_260#_c_83_n 0.0298057f $X=-0.19 $Y=-0.245 $X2=4.15 $Y2=2.29
cc_9 VNB N_A_83_260#_c_84_n 0.00625835f $X=-0.19 $Y=-0.245 $X2=1.955 $Y2=1.095
cc_10 VNB N_A_83_260#_c_85_n 0.00255036f $X=-0.19 $Y=-0.245 $X2=2.585 $Y2=1.095
cc_11 VNB N_A_83_260#_c_86_n 0.102727f $X=-0.19 $Y=-0.245 $X2=1.855 $Y2=1.532
cc_12 VNB N_A_M1001_g 0.0256588f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_c_212_n 0.0234795f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_c_213_n 0.0260576f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_15 VNB N_A_c_214_n 0.00338952f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=0.74
cc_16 VNB A 0.0080355f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=1.765
cc_17 VNB N_B_M1000_g 0.0399583f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB B 0.00357747f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.765
cc_19 VNB N_B_c_288_n 0.0331402f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=0.74
cc_20 VNB N_VPWR_c_332_n 0.183584f $X=-0.19 $Y=-0.245 $X2=1.955 $Y2=1.095
cc_21 VNB N_X_c_394_n 9.41836e-19 $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_22 VNB N_X_c_395_n 0.00715794f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=1.3
cc_23 VNB N_X_c_396_n 0.00206666f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=2.4
cc_24 VNB N_X_c_397_n 0.00485313f $X=-0.19 $Y=-0.245 $X2=1.405 $Y2=2.4
cc_25 VNB N_X_c_398_n 0.0025013f $X=-0.19 $Y=-0.245 $X2=1.87 $Y2=0.74
cc_26 VNB N_X_c_399_n 0.0019324f $X=-0.19 $Y=-0.245 $X2=2.42 $Y2=1.095
cc_27 VNB X 0.0264317f $X=-0.19 $Y=-0.245 $X2=2.585 $Y2=1.01
cc_28 VNB N_VGND_c_506_n 0.010678f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_29 VNB N_VGND_c_507_n 0.0274133f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=0.74
cc_30 VNB N_VGND_c_508_n 0.00497771f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=2.4
cc_31 VNB N_VGND_c_509_n 0.00571437f $X=-0.19 $Y=-0.245 $X2=1.355 $Y2=0.74
cc_32 VNB N_VGND_c_510_n 0.0172524f $X=-0.19 $Y=-0.245 $X2=1.405 $Y2=2.4
cc_33 VNB N_VGND_c_511_n 0.00461913f $X=-0.19 $Y=-0.245 $X2=1.405 $Y2=2.4
cc_34 VNB N_VGND_c_512_n 0.0196058f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_513_n 0.0185359f $X=-0.19 $Y=-0.245 $X2=0.76 $Y2=1.465
cc_36 VNB N_VGND_c_514_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=2.585 $Y2=0.515
cc_37 VNB N_VGND_c_515_n 0.070232f $X=-0.19 $Y=-0.245 $X2=3.23 $Y2=2.375
cc_38 VNB N_VGND_c_516_n 0.248241f $X=-0.19 $Y=-0.245 $X2=1.955 $Y2=1.095
cc_39 VPB N_A_83_260#_c_87_n 0.0164089f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.765
cc_40 VPB N_A_83_260#_c_88_n 0.0152457f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=1.765
cc_41 VPB N_A_83_260#_c_89_n 0.015247f $X=-0.19 $Y=1.66 $X2=1.405 $Y2=1.765
cc_42 VPB N_A_83_260#_c_90_n 0.016349f $X=-0.19 $Y=1.66 $X2=1.855 $Y2=1.765
cc_43 VPB N_A_83_260#_c_91_n 0.00863795f $X=-0.19 $Y=1.66 $X2=4.065 $Y2=2.375
cc_44 VPB N_A_83_260#_c_83_n 0.0255824f $X=-0.19 $Y=1.66 $X2=4.15 $Y2=2.29
cc_45 VPB N_A_83_260#_c_86_n 0.0266937f $X=-0.19 $Y=1.66 $X2=1.855 $Y2=1.532
cc_46 VPB N_A_c_212_n 0.0294771f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_47 VPB N_A_c_213_n 0.0348552f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.74
cc_48 VPB N_A_c_214_n 0.00318353f $X=-0.19 $Y=1.66 $X2=0.925 $Y2=0.74
cc_49 VPB A 0.00280119f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=1.765
cc_50 VPB N_B_c_289_n 0.0139264f $X=-0.19 $Y=1.66 $X2=2.445 $Y2=0.37
cc_51 VPB N_B_c_290_n 0.0143254f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.74
cc_52 VPB B 0.00250427f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.765
cc_53 VPB N_B_c_288_n 0.0296827f $X=-0.19 $Y=1.66 $X2=0.925 $Y2=0.74
cc_54 VPB N_VPWR_c_333_n 0.0106521f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.4
cc_55 VPB N_VPWR_c_334_n 0.0428822f $X=-0.19 $Y=1.66 $X2=0.925 $Y2=0.74
cc_56 VPB N_VPWR_c_335_n 0.00799266f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=2.4
cc_57 VPB N_VPWR_c_336_n 0.00904194f $X=-0.19 $Y=1.66 $X2=1.355 $Y2=0.74
cc_58 VPB N_VPWR_c_337_n 0.011133f $X=-0.19 $Y=1.66 $X2=1.405 $Y2=1.765
cc_59 VPB N_VPWR_c_338_n 0.025299f $X=-0.19 $Y=1.66 $X2=1.405 $Y2=2.4
cc_60 VPB N_VPWR_c_339_n 0.0206041f $X=-0.19 $Y=1.66 $X2=1.855 $Y2=2.4
cc_61 VPB N_VPWR_c_340_n 0.00324402f $X=-0.19 $Y=1.66 $X2=1.87 $Y2=1.3
cc_62 VPB N_VPWR_c_341_n 0.0206041f $X=-0.19 $Y=1.66 $X2=0.76 $Y2=1.465
cc_63 VPB N_VPWR_c_342_n 0.0412895f $X=-0.19 $Y=1.66 $X2=1.78 $Y2=1.465
cc_64 VPB N_VPWR_c_343_n 0.0047828f $X=-0.19 $Y=1.66 $X2=4.065 $Y2=2.375
cc_65 VPB N_VPWR_c_332_n 0.0811823f $X=-0.19 $Y=1.66 $X2=1.955 $Y2=1.095
cc_66 VPB N_X_c_401_n 0.00102565f $X=-0.19 $Y=1.66 $X2=0.925 $Y2=0.74
cc_67 VPB N_X_c_402_n 0.00724103f $X=-0.19 $Y=1.66 $X2=0.925 $Y2=0.74
cc_68 VPB N_X_c_403_n 0.00257348f $X=-0.19 $Y=1.66 $X2=1.355 $Y2=0.74
cc_69 VPB N_X_c_404_n 0.00363002f $X=-0.19 $Y=1.66 $X2=1.855 $Y2=2.4
cc_70 VPB N_X_c_405_n 0.00257348f $X=-0.19 $Y=1.66 $X2=0.76 $Y2=1.465
cc_71 VPB N_X_c_406_n 0.00187467f $X=-0.19 $Y=1.66 $X2=2.04 $Y2=1.095
cc_72 VPB X 0.00690691f $X=-0.19 $Y=1.66 $X2=2.585 $Y2=1.01
cc_73 VPB N_A_493_388#_c_474_n 0.00467613f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.765
cc_74 VPB N_A_493_388#_c_475_n 0.00244157f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.4
cc_75 VPB N_A_493_388#_c_476_n 0.00266025f $X=-0.19 $Y=1.66 $X2=0.925 $Y2=1.3
cc_76 N_A_83_260#_M1013_g N_A_M1001_g 0.0274315f $X=1.87 $Y=0.74 $X2=0 $Y2=0
cc_77 N_A_83_260#_c_80_n N_A_M1001_g 0.0110153f $X=2.42 $Y=1.095 $X2=0 $Y2=0
cc_78 N_A_83_260#_c_81_n N_A_M1001_g 0.00943664f $X=2.585 $Y=0.515 $X2=0 $Y2=0
cc_79 N_A_83_260#_c_84_n N_A_M1001_g 0.00344278f $X=1.955 $Y=1.095 $X2=0 $Y2=0
cc_80 N_A_83_260#_c_85_n N_A_M1001_g 0.0016818f $X=2.585 $Y=1.095 $X2=0 $Y2=0
cc_81 N_A_83_260#_c_90_n N_A_c_212_n 0.0225647f $X=1.855 $Y=1.765 $X2=0 $Y2=0
cc_82 N_A_83_260#_c_80_n N_A_c_212_n 5.99205e-19 $X=2.42 $Y=1.095 $X2=0 $Y2=0
cc_83 N_A_83_260#_c_84_n N_A_c_212_n 8.67352e-19 $X=1.955 $Y=1.095 $X2=0 $Y2=0
cc_84 N_A_83_260#_c_85_n N_A_c_212_n 7.49199e-19 $X=2.585 $Y=1.095 $X2=0 $Y2=0
cc_85 N_A_83_260#_c_86_n N_A_c_212_n 0.0185112f $X=1.855 $Y=1.532 $X2=0 $Y2=0
cc_86 N_A_83_260#_c_82_n N_A_c_213_n 0.00280427f $X=4.065 $Y=1.095 $X2=0 $Y2=0
cc_87 N_A_83_260#_c_105_p N_A_c_213_n 7.20833e-19 $X=3.105 $Y=2.46 $X2=0 $Y2=0
cc_88 N_A_83_260#_c_91_n N_A_c_213_n 0.0166043f $X=4.065 $Y=2.375 $X2=0 $Y2=0
cc_89 N_A_83_260#_c_83_n N_A_c_213_n 0.0154998f $X=4.15 $Y=2.29 $X2=0 $Y2=0
cc_90 N_A_83_260#_M1009_d N_A_c_234_n 0.00375066f $X=2.915 $Y=1.94 $X2=0 $Y2=0
cc_91 N_A_83_260#_c_91_n N_A_c_234_n 0.0381755f $X=4.065 $Y=2.375 $X2=0 $Y2=0
cc_92 N_A_83_260#_c_110_p N_A_c_234_n 0.0151034f $X=3.23 $Y=2.375 $X2=0 $Y2=0
cc_93 N_A_83_260#_c_82_n N_A_c_214_n 0.0170702f $X=4.065 $Y=1.095 $X2=0 $Y2=0
cc_94 N_A_83_260#_c_83_n N_A_c_214_n 0.0375789f $X=4.15 $Y=2.29 $X2=0 $Y2=0
cc_95 N_A_83_260#_c_90_n A 0.00212985f $X=1.855 $Y=1.765 $X2=0 $Y2=0
cc_96 N_A_83_260#_c_80_n A 0.0161138f $X=2.42 $Y=1.095 $X2=0 $Y2=0
cc_97 N_A_83_260#_c_82_n A 3.8449e-19 $X=4.065 $Y=1.095 $X2=0 $Y2=0
cc_98 N_A_83_260#_c_84_n A 0.0219858f $X=1.955 $Y=1.095 $X2=0 $Y2=0
cc_99 N_A_83_260#_c_85_n A 0.0301826f $X=2.585 $Y=1.095 $X2=0 $Y2=0
cc_100 N_A_83_260#_c_86_n A 0.00266487f $X=1.855 $Y=1.532 $X2=0 $Y2=0
cc_101 N_A_83_260#_c_105_p N_B_c_289_n 0.00107601f $X=3.105 $Y=2.46 $X2=-0.19
+ $Y2=-0.245
cc_102 N_A_83_260#_c_110_p N_B_c_289_n 8.55285e-19 $X=3.23 $Y=2.375 $X2=-0.19
+ $Y2=-0.245
cc_103 N_A_83_260#_c_81_n N_B_M1000_g 4.78879e-19 $X=2.585 $Y=0.515 $X2=0 $Y2=0
cc_104 N_A_83_260#_c_82_n N_B_M1000_g 0.0200689f $X=4.065 $Y=1.095 $X2=0 $Y2=0
cc_105 N_A_83_260#_c_105_p N_B_c_290_n 0.00453488f $X=3.105 $Y=2.46 $X2=0 $Y2=0
cc_106 N_A_83_260#_c_91_n N_B_c_290_n 0.00939201f $X=4.065 $Y=2.375 $X2=0 $Y2=0
cc_107 N_A_83_260#_c_110_p N_B_c_290_n 6.68968e-19 $X=3.23 $Y=2.375 $X2=0 $Y2=0
cc_108 N_A_83_260#_c_82_n B 0.0174918f $X=4.065 $Y=1.095 $X2=0 $Y2=0
cc_109 N_A_83_260#_c_82_n N_B_c_288_n 0.00662087f $X=4.065 $Y=1.095 $X2=0 $Y2=0
cc_110 N_A_83_260#_c_91_n N_VPWR_M1010_s 0.00979801f $X=4.065 $Y=2.375 $X2=0
+ $Y2=0
cc_111 N_A_83_260#_c_83_n N_VPWR_M1010_s 0.00581094f $X=4.15 $Y=2.29 $X2=0 $Y2=0
cc_112 N_A_83_260#_c_87_n N_VPWR_c_334_n 0.00993564f $X=0.505 $Y=1.765 $X2=0
+ $Y2=0
cc_113 N_A_83_260#_c_88_n N_VPWR_c_335_n 0.00586501f $X=0.955 $Y=1.765 $X2=0
+ $Y2=0
cc_114 N_A_83_260#_c_89_n N_VPWR_c_335_n 0.00586501f $X=1.405 $Y=1.765 $X2=0
+ $Y2=0
cc_115 N_A_83_260#_c_90_n N_VPWR_c_336_n 0.00700356f $X=1.855 $Y=1.765 $X2=0
+ $Y2=0
cc_116 N_A_83_260#_c_84_n N_VPWR_c_336_n 0.00183071f $X=1.955 $Y=1.095 $X2=0
+ $Y2=0
cc_117 N_A_83_260#_c_91_n N_VPWR_c_338_n 0.0234202f $X=4.065 $Y=2.375 $X2=0
+ $Y2=0
cc_118 N_A_83_260#_c_87_n N_VPWR_c_339_n 0.00445602f $X=0.505 $Y=1.765 $X2=0
+ $Y2=0
cc_119 N_A_83_260#_c_88_n N_VPWR_c_339_n 0.00445602f $X=0.955 $Y=1.765 $X2=0
+ $Y2=0
cc_120 N_A_83_260#_c_89_n N_VPWR_c_341_n 0.00445602f $X=1.405 $Y=1.765 $X2=0
+ $Y2=0
cc_121 N_A_83_260#_c_90_n N_VPWR_c_341_n 0.00445602f $X=1.855 $Y=1.765 $X2=0
+ $Y2=0
cc_122 N_A_83_260#_c_87_n N_VPWR_c_332_n 0.00861084f $X=0.505 $Y=1.765 $X2=0
+ $Y2=0
cc_123 N_A_83_260#_c_88_n N_VPWR_c_332_n 0.00857589f $X=0.955 $Y=1.765 $X2=0
+ $Y2=0
cc_124 N_A_83_260#_c_89_n N_VPWR_c_332_n 0.00857589f $X=1.405 $Y=1.765 $X2=0
+ $Y2=0
cc_125 N_A_83_260#_c_90_n N_VPWR_c_332_n 0.00862391f $X=1.855 $Y=1.765 $X2=0
+ $Y2=0
cc_126 N_A_83_260#_M1002_g N_X_c_394_n 0.0143243f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_127 N_A_83_260#_c_87_n N_X_c_401_n 0.0152499f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_128 N_A_83_260#_c_86_n N_X_c_401_n 5.4426e-19 $X=1.855 $Y=1.532 $X2=0 $Y2=0
cc_129 N_A_83_260#_M1002_g N_X_c_396_n 0.0128625f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_130 N_A_83_260#_M1003_g N_X_c_396_n 3.97481e-19 $X=0.925 $Y=0.74 $X2=0 $Y2=0
cc_131 N_A_83_260#_c_87_n N_X_c_403_n 0.017229f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_132 N_A_83_260#_c_88_n N_X_c_403_n 0.0125029f $X=0.955 $Y=1.765 $X2=0 $Y2=0
cc_133 N_A_83_260#_c_89_n N_X_c_403_n 6.9119e-19 $X=1.405 $Y=1.765 $X2=0 $Y2=0
cc_134 N_A_83_260#_M1003_g N_X_c_397_n 0.0124434f $X=0.925 $Y=0.74 $X2=0 $Y2=0
cc_135 N_A_83_260#_M1012_g N_X_c_397_n 0.0121215f $X=1.355 $Y=0.74 $X2=0 $Y2=0
cc_136 N_A_83_260#_M1013_g N_X_c_397_n 0.00257018f $X=1.87 $Y=0.74 $X2=0 $Y2=0
cc_137 N_A_83_260#_c_155_p N_X_c_397_n 0.0695156f $X=1.87 $Y=1.465 $X2=0 $Y2=0
cc_138 N_A_83_260#_c_84_n N_X_c_397_n 0.0095065f $X=1.955 $Y=1.095 $X2=0 $Y2=0
cc_139 N_A_83_260#_c_86_n N_X_c_397_n 0.00643527f $X=1.855 $Y=1.532 $X2=0 $Y2=0
cc_140 N_A_83_260#_c_88_n N_X_c_404_n 0.0120074f $X=0.955 $Y=1.765 $X2=0 $Y2=0
cc_141 N_A_83_260#_c_89_n N_X_c_404_n 0.0129464f $X=1.405 $Y=1.765 $X2=0 $Y2=0
cc_142 N_A_83_260#_c_90_n N_X_c_404_n 0.0033951f $X=1.855 $Y=1.765 $X2=0 $Y2=0
cc_143 N_A_83_260#_c_155_p N_X_c_404_n 0.0694546f $X=1.87 $Y=1.465 $X2=0 $Y2=0
cc_144 N_A_83_260#_c_86_n N_X_c_404_n 0.0152376f $X=1.855 $Y=1.532 $X2=0 $Y2=0
cc_145 N_A_83_260#_M1003_g N_X_c_398_n 6.70758e-19 $X=0.925 $Y=0.74 $X2=0 $Y2=0
cc_146 N_A_83_260#_M1012_g N_X_c_398_n 0.00887699f $X=1.355 $Y=0.74 $X2=0 $Y2=0
cc_147 N_A_83_260#_M1013_g N_X_c_398_n 0.00731762f $X=1.87 $Y=0.74 $X2=0 $Y2=0
cc_148 N_A_83_260#_c_88_n N_X_c_405_n 6.9119e-19 $X=0.955 $Y=1.765 $X2=0 $Y2=0
cc_149 N_A_83_260#_c_89_n N_X_c_405_n 0.0125029f $X=1.405 $Y=1.765 $X2=0 $Y2=0
cc_150 N_A_83_260#_c_90_n N_X_c_405_n 0.0127172f $X=1.855 $Y=1.765 $X2=0 $Y2=0
cc_151 N_A_83_260#_M1002_g N_X_c_399_n 0.00132305f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_152 N_A_83_260#_c_155_p N_X_c_399_n 0.0168687f $X=1.87 $Y=1.465 $X2=0 $Y2=0
cc_153 N_A_83_260#_c_86_n N_X_c_399_n 0.00232957f $X=1.855 $Y=1.532 $X2=0 $Y2=0
cc_154 N_A_83_260#_c_87_n N_X_c_406_n 0.00114729f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_155 N_A_83_260#_c_88_n N_X_c_406_n 9.3899e-19 $X=0.955 $Y=1.765 $X2=0 $Y2=0
cc_156 N_A_83_260#_c_155_p N_X_c_406_n 0.0252322f $X=1.87 $Y=1.465 $X2=0 $Y2=0
cc_157 N_A_83_260#_c_86_n N_X_c_406_n 0.00805341f $X=1.855 $Y=1.532 $X2=0 $Y2=0
cc_158 N_A_83_260#_M1002_g X 0.0067245f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_159 N_A_83_260#_c_87_n X 0.00133808f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_160 N_A_83_260#_c_155_p X 0.0206535f $X=1.87 $Y=1.465 $X2=0 $Y2=0
cc_161 N_A_83_260#_c_86_n X 0.0158588f $X=1.855 $Y=1.532 $X2=0 $Y2=0
cc_162 N_A_83_260#_c_91_n N_A_493_388#_M1011_s 0.00493401f $X=4.065 $Y=2.375
+ $X2=0 $Y2=0
cc_163 N_A_83_260#_c_105_p N_A_493_388#_c_478_n 0.0184049f $X=3.105 $Y=2.46
+ $X2=0 $Y2=0
cc_164 N_A_83_260#_c_110_p N_A_493_388#_c_478_n 0.0123817f $X=3.23 $Y=2.375
+ $X2=0 $Y2=0
cc_165 N_A_83_260#_M1009_d N_A_493_388#_c_474_n 0.00222494f $X=2.915 $Y=1.94
+ $X2=0 $Y2=0
cc_166 N_A_83_260#_c_105_p N_A_493_388#_c_474_n 0.0140094f $X=3.105 $Y=2.46
+ $X2=0 $Y2=0
cc_167 N_A_83_260#_c_91_n N_A_493_388#_c_474_n 0.0041825f $X=4.065 $Y=2.375
+ $X2=0 $Y2=0
cc_168 N_A_83_260#_c_91_n N_A_493_388#_c_476_n 0.0195451f $X=4.065 $Y=2.375
+ $X2=0 $Y2=0
cc_169 N_A_83_260#_c_80_n N_VGND_M1013_s 0.0023395f $X=2.42 $Y=1.095 $X2=0 $Y2=0
cc_170 N_A_83_260#_c_84_n N_VGND_M1013_s 6.54518e-19 $X=1.955 $Y=1.095 $X2=0
+ $Y2=0
cc_171 N_A_83_260#_c_82_n N_VGND_M1000_d 0.0186685f $X=4.065 $Y=1.095 $X2=0
+ $Y2=0
cc_172 N_A_83_260#_M1002_g N_VGND_c_507_n 0.00409307f $X=0.495 $Y=0.74 $X2=0
+ $Y2=0
cc_173 N_A_83_260#_M1002_g N_VGND_c_508_n 5.05592e-19 $X=0.495 $Y=0.74 $X2=0
+ $Y2=0
cc_174 N_A_83_260#_M1003_g N_VGND_c_508_n 0.008885f $X=0.925 $Y=0.74 $X2=0 $Y2=0
cc_175 N_A_83_260#_M1012_g N_VGND_c_508_n 0.00307459f $X=1.355 $Y=0.74 $X2=0
+ $Y2=0
cc_176 N_A_83_260#_M1012_g N_VGND_c_509_n 7.0576e-19 $X=1.355 $Y=0.74 $X2=0
+ $Y2=0
cc_177 N_A_83_260#_M1013_g N_VGND_c_509_n 0.0114822f $X=1.87 $Y=0.74 $X2=0 $Y2=0
cc_178 N_A_83_260#_c_80_n N_VGND_c_509_n 0.016109f $X=2.42 $Y=1.095 $X2=0 $Y2=0
cc_179 N_A_83_260#_c_81_n N_VGND_c_509_n 0.0191765f $X=2.585 $Y=0.515 $X2=0
+ $Y2=0
cc_180 N_A_83_260#_c_84_n N_VGND_c_509_n 0.00528841f $X=1.955 $Y=1.095 $X2=0
+ $Y2=0
cc_181 N_A_83_260#_M1002_g N_VGND_c_510_n 0.00434272f $X=0.495 $Y=0.74 $X2=0
+ $Y2=0
cc_182 N_A_83_260#_M1003_g N_VGND_c_510_n 0.00383152f $X=0.925 $Y=0.74 $X2=0
+ $Y2=0
cc_183 N_A_83_260#_M1012_g N_VGND_c_512_n 0.00434272f $X=1.355 $Y=0.74 $X2=0
+ $Y2=0
cc_184 N_A_83_260#_M1013_g N_VGND_c_512_n 0.00383152f $X=1.87 $Y=0.74 $X2=0
+ $Y2=0
cc_185 N_A_83_260#_c_81_n N_VGND_c_513_n 0.0145639f $X=2.585 $Y=0.515 $X2=0
+ $Y2=0
cc_186 N_A_83_260#_c_81_n N_VGND_c_515_n 0.0214346f $X=2.585 $Y=0.515 $X2=0
+ $Y2=0
cc_187 N_A_83_260#_c_82_n N_VGND_c_515_n 0.101081f $X=4.065 $Y=1.095 $X2=0 $Y2=0
cc_188 N_A_83_260#_M1002_g N_VGND_c_516_n 0.00823942f $X=0.495 $Y=0.74 $X2=0
+ $Y2=0
cc_189 N_A_83_260#_M1003_g N_VGND_c_516_n 0.0075754f $X=0.925 $Y=0.74 $X2=0
+ $Y2=0
cc_190 N_A_83_260#_M1012_g N_VGND_c_516_n 0.00821072f $X=1.355 $Y=0.74 $X2=0
+ $Y2=0
cc_191 N_A_83_260#_M1013_g N_VGND_c_516_n 0.00758328f $X=1.87 $Y=0.74 $X2=0
+ $Y2=0
cc_192 N_A_83_260#_c_81_n N_VGND_c_516_n 0.0119984f $X=2.585 $Y=0.515 $X2=0
+ $Y2=0
cc_193 N_A_c_212_n N_B_c_289_n 0.0206787f $X=2.39 $Y=1.865 $X2=-0.19 $Y2=-0.245
cc_194 N_A_c_234_n N_B_c_289_n 0.0189467f $X=3.59 $Y=2.035 $X2=-0.19 $Y2=-0.245
cc_195 A N_B_c_289_n 0.0024151f $X=2.555 $Y=1.58 $X2=-0.19 $Y2=-0.245
cc_196 N_A_M1001_g N_B_M1000_g 0.0160308f $X=2.37 $Y=0.74 $X2=0 $Y2=0
cc_197 N_A_c_212_n N_B_M1000_g 0.0144774f $X=2.39 $Y=1.865 $X2=0 $Y2=0
cc_198 A N_B_M1000_g 0.00466058f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_199 N_A_c_213_n N_B_c_290_n 0.0351367f $X=3.79 $Y=1.865 $X2=0 $Y2=0
cc_200 N_A_c_234_n N_B_c_290_n 0.013799f $X=3.59 $Y=2.035 $X2=0 $Y2=0
cc_201 N_A_c_214_n N_B_c_290_n 0.00187813f $X=3.755 $Y=1.615 $X2=0 $Y2=0
cc_202 N_A_c_212_n B 2.24496e-19 $X=2.39 $Y=1.865 $X2=0 $Y2=0
cc_203 N_A_c_213_n B 0.00116857f $X=3.79 $Y=1.865 $X2=0 $Y2=0
cc_204 N_A_c_234_n B 0.0204896f $X=3.59 $Y=2.035 $X2=0 $Y2=0
cc_205 N_A_c_214_n B 0.0142939f $X=3.755 $Y=1.615 $X2=0 $Y2=0
cc_206 A B 0.0266673f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_207 N_A_c_212_n N_B_c_288_n 0.012021f $X=2.39 $Y=1.865 $X2=0 $Y2=0
cc_208 N_A_c_213_n N_B_c_288_n 0.0191286f $X=3.79 $Y=1.865 $X2=0 $Y2=0
cc_209 N_A_c_234_n N_B_c_288_n 0.00172007f $X=3.59 $Y=2.035 $X2=0 $Y2=0
cc_210 N_A_c_214_n N_B_c_288_n 0.00335266f $X=3.755 $Y=1.615 $X2=0 $Y2=0
cc_211 A N_B_c_288_n 0.00694941f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_212 A N_VPWR_M1008_d 0.00244786f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_213 N_A_c_212_n N_VPWR_c_336_n 0.0115626f $X=2.39 $Y=1.865 $X2=0 $Y2=0
cc_214 A N_VPWR_c_336_n 0.00303731f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_215 N_A_c_213_n N_VPWR_c_338_n 0.00401341f $X=3.79 $Y=1.865 $X2=0 $Y2=0
cc_216 N_A_c_212_n N_VPWR_c_342_n 0.0051666f $X=2.39 $Y=1.865 $X2=0 $Y2=0
cc_217 N_A_c_213_n N_VPWR_c_342_n 0.00519777f $X=3.79 $Y=1.865 $X2=0 $Y2=0
cc_218 N_A_c_212_n N_VPWR_c_332_n 0.00485508f $X=2.39 $Y=1.865 $X2=0 $Y2=0
cc_219 N_A_c_213_n N_VPWR_c_332_n 0.00489105f $X=3.79 $Y=1.865 $X2=0 $Y2=0
cc_220 N_A_c_212_n N_X_c_404_n 2.29428e-19 $X=2.39 $Y=1.865 $X2=0 $Y2=0
cc_221 A N_X_c_404_n 0.00651605f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_222 N_A_c_212_n N_X_c_405_n 8.94356e-19 $X=2.39 $Y=1.865 $X2=0 $Y2=0
cc_223 A N_A_493_388#_M1007_d 0.00205832f $X=2.555 $Y=1.58 $X2=-0.19 $Y2=-0.245
cc_224 N_A_c_234_n N_A_493_388#_M1011_s 0.00889447f $X=3.59 $Y=2.035 $X2=0 $Y2=0
cc_225 N_A_c_212_n N_A_493_388#_c_478_n 0.00680887f $X=2.39 $Y=1.865 $X2=0 $Y2=0
cc_226 N_A_c_234_n N_A_493_388#_c_478_n 0.00102433f $X=3.59 $Y=2.035 $X2=0 $Y2=0
cc_227 A N_A_493_388#_c_478_n 0.0174163f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_228 N_A_c_212_n N_A_493_388#_c_475_n 0.00353968f $X=2.39 $Y=1.865 $X2=0 $Y2=0
cc_229 N_A_c_213_n N_A_493_388#_c_476_n 0.00668659f $X=3.79 $Y=1.865 $X2=0 $Y2=0
cc_230 N_A_M1001_g N_VGND_c_509_n 0.00432719f $X=2.37 $Y=0.74 $X2=0 $Y2=0
cc_231 N_A_M1001_g N_VGND_c_513_n 0.00434272f $X=2.37 $Y=0.74 $X2=0 $Y2=0
cc_232 N_A_M1001_g N_VGND_c_515_n 4.84975e-19 $X=2.37 $Y=0.74 $X2=0 $Y2=0
cc_233 N_A_M1001_g N_VGND_c_516_n 0.00821358f $X=2.37 $Y=0.74 $X2=0 $Y2=0
cc_234 N_B_c_289_n N_VPWR_c_342_n 9.78684e-19 $X=2.84 $Y=1.865 $X2=0 $Y2=0
cc_235 N_B_c_290_n N_VPWR_c_342_n 9.59479e-19 $X=3.29 $Y=1.865 $X2=0 $Y2=0
cc_236 N_B_c_289_n N_A_493_388#_c_478_n 0.00778115f $X=2.84 $Y=1.865 $X2=0 $Y2=0
cc_237 N_B_c_290_n N_A_493_388#_c_478_n 6.70277e-19 $X=3.29 $Y=1.865 $X2=0 $Y2=0
cc_238 N_B_c_289_n N_A_493_388#_c_474_n 0.0118753f $X=2.84 $Y=1.865 $X2=0 $Y2=0
cc_239 N_B_c_290_n N_A_493_388#_c_474_n 0.0107106f $X=3.29 $Y=1.865 $X2=0 $Y2=0
cc_240 N_B_c_289_n N_A_493_388#_c_475_n 0.0020313f $X=2.84 $Y=1.865 $X2=0 $Y2=0
cc_241 N_B_c_290_n N_A_493_388#_c_476_n 4.94289e-19 $X=3.29 $Y=1.865 $X2=0 $Y2=0
cc_242 N_B_M1000_g N_VGND_c_513_n 0.00429299f $X=2.855 $Y=0.74 $X2=0 $Y2=0
cc_243 N_B_M1000_g N_VGND_c_515_n 0.0126649f $X=2.855 $Y=0.74 $X2=0 $Y2=0
cc_244 N_B_M1000_g N_VGND_c_516_n 0.00843495f $X=2.855 $Y=0.74 $X2=0 $Y2=0
cc_245 N_VPWR_M1004_d N_X_c_401_n 4.28442e-19 $X=0.135 $Y=1.84 $X2=0 $Y2=0
cc_246 N_VPWR_c_334_n N_X_c_401_n 6.9575e-19 $X=0.28 $Y=2.305 $X2=0 $Y2=0
cc_247 N_VPWR_M1004_d N_X_c_402_n 0.00326206f $X=0.135 $Y=1.84 $X2=0 $Y2=0
cc_248 N_VPWR_c_334_n N_X_c_402_n 0.0207257f $X=0.28 $Y=2.305 $X2=0 $Y2=0
cc_249 N_VPWR_c_334_n N_X_c_403_n 0.0563525f $X=0.28 $Y=2.305 $X2=0 $Y2=0
cc_250 N_VPWR_c_335_n N_X_c_403_n 0.0547423f $X=1.18 $Y=2.305 $X2=0 $Y2=0
cc_251 N_VPWR_c_339_n N_X_c_403_n 0.014552f $X=1.095 $Y=3.33 $X2=0 $Y2=0
cc_252 N_VPWR_c_332_n N_X_c_403_n 0.0119791f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_253 N_VPWR_M1005_d N_X_c_404_n 0.00247267f $X=1.03 $Y=1.84 $X2=0 $Y2=0
cc_254 N_VPWR_c_335_n N_X_c_404_n 0.0136682f $X=1.18 $Y=2.305 $X2=0 $Y2=0
cc_255 N_VPWR_c_335_n N_X_c_405_n 0.0547423f $X=1.18 $Y=2.305 $X2=0 $Y2=0
cc_256 N_VPWR_c_336_n N_X_c_405_n 0.0576935f $X=2.08 $Y=2.285 $X2=0 $Y2=0
cc_257 N_VPWR_c_341_n N_X_c_405_n 0.014552f $X=1.995 $Y=3.33 $X2=0 $Y2=0
cc_258 N_VPWR_c_332_n N_X_c_405_n 0.0119791f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_259 N_VPWR_c_336_n N_A_493_388#_c_478_n 0.0404301f $X=2.08 $Y=2.285 $X2=0
+ $Y2=0
cc_260 N_VPWR_c_342_n N_A_493_388#_c_474_n 0.0399102f $X=3.93 $Y=3.33 $X2=0
+ $Y2=0
cc_261 N_VPWR_c_332_n N_A_493_388#_c_474_n 0.0233066f $X=4.08 $Y=3.33 $X2=0
+ $Y2=0
cc_262 N_VPWR_c_336_n N_A_493_388#_c_475_n 0.012097f $X=2.08 $Y=2.285 $X2=0
+ $Y2=0
cc_263 N_VPWR_c_342_n N_A_493_388#_c_475_n 0.0236566f $X=3.93 $Y=3.33 $X2=0
+ $Y2=0
cc_264 N_VPWR_c_332_n N_A_493_388#_c_475_n 0.0128296f $X=4.08 $Y=3.33 $X2=0
+ $Y2=0
cc_265 N_VPWR_c_338_n N_A_493_388#_c_476_n 0.0302797f $X=4.025 $Y=2.795 $X2=0
+ $Y2=0
cc_266 N_VPWR_c_342_n N_A_493_388#_c_476_n 0.0227798f $X=3.93 $Y=3.33 $X2=0
+ $Y2=0
cc_267 N_VPWR_c_332_n N_A_493_388#_c_476_n 0.0126147f $X=4.08 $Y=3.33 $X2=0
+ $Y2=0
cc_268 N_X_c_395_n N_VGND_M1002_s 0.00330634f $X=0.355 $Y=1.045 $X2=-0.19
+ $Y2=-0.245
cc_269 N_X_c_397_n N_VGND_M1003_s 0.00176461f $X=1.405 $Y=1.045 $X2=0 $Y2=0
cc_270 N_X_c_394_n N_VGND_c_507_n 6.14392e-19 $X=0.545 $Y=1.045 $X2=0 $Y2=0
cc_271 N_X_c_395_n N_VGND_c_507_n 0.0207726f $X=0.355 $Y=1.045 $X2=0 $Y2=0
cc_272 N_X_c_396_n N_VGND_c_507_n 0.0158413f $X=0.71 $Y=0.515 $X2=0 $Y2=0
cc_273 N_X_c_396_n N_VGND_c_508_n 0.0158413f $X=0.71 $Y=0.515 $X2=0 $Y2=0
cc_274 N_X_c_397_n N_VGND_c_508_n 0.0153337f $X=1.405 $Y=1.045 $X2=0 $Y2=0
cc_275 N_X_c_398_n N_VGND_c_508_n 0.0162297f $X=1.59 $Y=0.515 $X2=0 $Y2=0
cc_276 N_X_c_398_n N_VGND_c_509_n 0.0309614f $X=1.59 $Y=0.515 $X2=0 $Y2=0
cc_277 N_X_c_396_n N_VGND_c_510_n 0.0109942f $X=0.71 $Y=0.515 $X2=0 $Y2=0
cc_278 N_X_c_398_n N_VGND_c_512_n 0.0130022f $X=1.59 $Y=0.515 $X2=0 $Y2=0
cc_279 N_X_c_396_n N_VGND_c_516_n 0.00904371f $X=0.71 $Y=0.515 $X2=0 $Y2=0
cc_280 N_X_c_398_n N_VGND_c_516_n 0.0107057f $X=1.59 $Y=0.515 $X2=0 $Y2=0
