# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_hs__sdfxtp_2
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_hs__sdfxtp_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  12.00000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.085000 1.190000 1.665000 1.845000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.576500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 11.055000 0.350000 11.385000 1.050000 ;
        RECT 11.105000 1.820000 11.435000 2.980000 ;
        RECT 11.215000 1.050000 11.385000 1.820000 ;
    END
  END Q
  PIN SCD
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.450000 1.435000 2.780000 2.150000 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425000 0.810000 0.835000 0.850000 ;
        RECT 0.425000 0.850000 2.205000 1.020000 ;
        RECT 0.425000 1.020000 0.835000 1.230000 ;
        RECT 1.875000 1.020000 2.205000 1.230000 ;
    END
  END SCE
  PIN CLK
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 3.290000 1.350000 3.685000 1.780000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT  0.000000 -0.085000 12.000000 0.085000 ;
        RECT  0.660000  0.085000  0.990000 0.640000 ;
        RECT  2.715000  0.085000  2.975000 0.810000 ;
        RECT  3.705000  0.085000  4.035000 0.840000 ;
        RECT  6.720000  0.085000  7.050000 0.550000 ;
        RECT  9.300000  0.085000  9.630000 0.810000 ;
        RECT 10.615000  0.085000 10.885000 1.050000 ;
        RECT 11.555000  0.085000 11.885000 1.130000 ;
      LAYER mcon ;
        RECT  0.155000 -0.085000  0.325000 0.085000 ;
        RECT  0.635000 -0.085000  0.805000 0.085000 ;
        RECT  1.115000 -0.085000  1.285000 0.085000 ;
        RECT  1.595000 -0.085000  1.765000 0.085000 ;
        RECT  2.075000 -0.085000  2.245000 0.085000 ;
        RECT  2.555000 -0.085000  2.725000 0.085000 ;
        RECT  3.035000 -0.085000  3.205000 0.085000 ;
        RECT  3.515000 -0.085000  3.685000 0.085000 ;
        RECT  3.995000 -0.085000  4.165000 0.085000 ;
        RECT  4.475000 -0.085000  4.645000 0.085000 ;
        RECT  4.955000 -0.085000  5.125000 0.085000 ;
        RECT  5.435000 -0.085000  5.605000 0.085000 ;
        RECT  5.915000 -0.085000  6.085000 0.085000 ;
        RECT  6.395000 -0.085000  6.565000 0.085000 ;
        RECT  6.875000 -0.085000  7.045000 0.085000 ;
        RECT  7.355000 -0.085000  7.525000 0.085000 ;
        RECT  7.835000 -0.085000  8.005000 0.085000 ;
        RECT  8.315000 -0.085000  8.485000 0.085000 ;
        RECT  8.795000 -0.085000  8.965000 0.085000 ;
        RECT  9.275000 -0.085000  9.445000 0.085000 ;
        RECT  9.755000 -0.085000  9.925000 0.085000 ;
        RECT 10.235000 -0.085000 10.405000 0.085000 ;
        RECT 10.715000 -0.085000 10.885000 0.085000 ;
        RECT 11.195000 -0.085000 11.365000 0.085000 ;
        RECT 11.675000 -0.085000 11.845000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.245000 12.000000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT  0.000000 3.245000 12.000000 3.415000 ;
        RECT  0.615000 2.355000  0.945000 3.245000 ;
        RECT  2.685000 2.790000  3.135000 3.245000 ;
        RECT  3.900000 2.790000  4.370000 3.245000 ;
        RECT  6.585000 2.520000  6.835000 3.245000 ;
        RECT  9.295000 2.590000  9.925000 3.245000 ;
        RECT 10.655000 1.820000 10.905000 3.245000 ;
        RECT 11.635000 1.820000 11.885000 3.245000 ;
      LAYER mcon ;
        RECT  0.155000 3.245000  0.325000 3.415000 ;
        RECT  0.635000 3.245000  0.805000 3.415000 ;
        RECT  1.115000 3.245000  1.285000 3.415000 ;
        RECT  1.595000 3.245000  1.765000 3.415000 ;
        RECT  2.075000 3.245000  2.245000 3.415000 ;
        RECT  2.555000 3.245000  2.725000 3.415000 ;
        RECT  3.035000 3.245000  3.205000 3.415000 ;
        RECT  3.515000 3.245000  3.685000 3.415000 ;
        RECT  3.995000 3.245000  4.165000 3.415000 ;
        RECT  4.475000 3.245000  4.645000 3.415000 ;
        RECT  4.955000 3.245000  5.125000 3.415000 ;
        RECT  5.435000 3.245000  5.605000 3.415000 ;
        RECT  5.915000 3.245000  6.085000 3.415000 ;
        RECT  6.395000 3.245000  6.565000 3.415000 ;
        RECT  6.875000 3.245000  7.045000 3.415000 ;
        RECT  7.355000 3.245000  7.525000 3.415000 ;
        RECT  7.835000 3.245000  8.005000 3.415000 ;
        RECT  8.315000 3.245000  8.485000 3.415000 ;
        RECT  8.795000 3.245000  8.965000 3.415000 ;
        RECT  9.275000 3.245000  9.445000 3.415000 ;
        RECT  9.755000 3.245000  9.925000 3.415000 ;
        RECT 10.235000 3.245000 10.405000 3.415000 ;
        RECT 10.715000 3.245000 10.885000 3.415000 ;
        RECT 11.195000 3.245000 11.365000 3.415000 ;
        RECT 11.675000 3.245000 11.845000 3.415000 ;
      LAYER met1 ;
        RECT 0.000000 3.085000 12.000000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.085000 0.390000  0.490000 0.640000 ;
      RECT  0.085000 0.640000  0.255000 1.470000 ;
      RECT  0.085000 1.470000  0.915000 2.015000 ;
      RECT  0.085000 2.015000  2.210000 2.185000 ;
      RECT  0.085000 2.185000  0.445000 2.925000 ;
      RECT  1.480000 0.350000  2.545000 0.680000 ;
      RECT  1.485000 2.355000  3.120000 2.450000 ;
      RECT  1.485000 2.450000  5.385000 2.620000 ;
      RECT  1.485000 2.620000  2.060000 2.945000 ;
      RECT  1.880000 1.775000  2.210000 2.015000 ;
      RECT  2.375000 0.680000  2.545000 1.095000 ;
      RECT  2.375000 1.095000  3.120000 1.265000 ;
      RECT  2.950000 1.265000  3.120000 2.355000 ;
      RECT  3.145000 0.330000  3.475000 0.920000 ;
      RECT  3.305000 0.920000  3.475000 1.010000 ;
      RECT  3.305000 1.010000  4.025000 1.180000 ;
      RECT  3.340000 1.950000  4.145000 2.280000 ;
      RECT  3.855000 1.180000  4.025000 1.300000 ;
      RECT  3.855000 1.300000  4.145000 1.950000 ;
      RECT  4.205000 0.255000  6.115000 0.425000 ;
      RECT  4.205000 0.425000  4.535000 1.130000 ;
      RECT  4.315000 1.300000  4.875000 1.470000 ;
      RECT  4.315000 1.470000  4.485000 2.450000 ;
      RECT  4.655000 1.820000  5.375000 2.280000 ;
      RECT  4.705000 0.595000  5.015000 0.940000 ;
      RECT  4.705000 0.940000  4.875000 1.300000 ;
      RECT  5.045000 1.610000  5.375000 1.820000 ;
      RECT  5.135000 2.620000  5.385000 2.980000 ;
      RECT  5.185000 0.425000  5.355000 1.610000 ;
      RECT  5.525000 0.595000  5.775000 0.940000 ;
      RECT  5.555000 0.940000  5.775000 1.630000 ;
      RECT  5.555000 1.630000  7.175000 1.800000 ;
      RECT  5.555000 1.800000  5.725000 2.520000 ;
      RECT  5.555000 2.520000  5.915000 2.980000 ;
      RECT  5.895000 1.970000  6.225000 2.130000 ;
      RECT  5.895000 2.130000  7.175000 2.300000 ;
      RECT  5.945000 0.425000  6.115000 0.720000 ;
      RECT  5.945000 0.720000  7.390000 0.890000 ;
      RECT  5.945000 0.890000  6.275000 1.360000 ;
      RECT  6.485000 1.060000  7.890000 1.230000 ;
      RECT  6.485000 1.230000  7.515000 1.390000 ;
      RECT  6.845000 1.800000  7.175000 1.960000 ;
      RECT  7.005000 2.300000  7.175000 2.905000 ;
      RECT  7.005000 2.905000  7.855000 3.075000 ;
      RECT  7.220000 0.255000  8.230000 0.425000 ;
      RECT  7.220000 0.425000  7.390000 0.720000 ;
      RECT  7.345000 1.390000  7.515000 2.610000 ;
      RECT  7.560000 0.595000  7.890000 1.060000 ;
      RECT  7.685000 1.600000  8.115000 1.930000 ;
      RECT  7.685000 1.930000  7.855000 2.905000 ;
      RECT  8.025000 2.490000  9.060000 2.660000 ;
      RECT  8.025000 2.660000  8.275000 2.920000 ;
      RECT  8.060000 0.425000  8.230000 1.030000 ;
      RECT  8.060000 1.030000  8.455000 1.360000 ;
      RECT  8.285000 1.360000  8.455000 1.990000 ;
      RECT  8.285000 1.990000  8.720000 2.320000 ;
      RECT  8.400000 0.350000  8.795000 0.640000 ;
      RECT  8.400000 0.640000  9.060000 0.810000 ;
      RECT  8.890000 0.810000  9.060000 2.075000 ;
      RECT  8.890000 2.075000 10.105000 2.245000 ;
      RECT  8.890000 2.245000  9.060000 2.490000 ;
      RECT  9.230000 1.070000 10.445000 1.220000 ;
      RECT  9.230000 1.220000 11.045000 1.240000 ;
      RECT  9.230000 1.240000  9.535000 1.905000 ;
      RECT  9.775000 1.410000 10.105000 2.075000 ;
      RECT  9.800000 0.350000 10.130000 1.070000 ;
      RECT 10.095000 2.415000 10.445000 2.920000 ;
      RECT 10.275000 1.240000 11.045000 1.550000 ;
      RECT 10.275000 1.550000 10.445000 2.415000 ;
  END
END sky130_fd_sc_hs__sdfxtp_2
