* File: sky130_fd_sc_hs__inv_4.pxi.spice
* Created: Tue Sep  1 20:07:05 2020
* 
x_PM_SKY130_FD_SC_HS__INV_4%A N_A_M1000_g N_A_c_49_n N_A_M1001_g N_A_c_50_n
+ N_A_M1002_g N_A_M1005_g N_A_c_51_n N_A_M1003_g N_A_M1006_g N_A_c_52_n
+ N_A_M1004_g N_A_M1007_g A A A A N_A_c_48_n PM_SKY130_FD_SC_HS__INV_4%A
x_PM_SKY130_FD_SC_HS__INV_4%VPWR N_VPWR_M1001_s N_VPWR_M1002_s N_VPWR_M1004_s
+ N_VPWR_c_121_n N_VPWR_c_122_n N_VPWR_c_123_n N_VPWR_c_124_n N_VPWR_c_125_n
+ N_VPWR_c_126_n VPWR N_VPWR_c_127_n N_VPWR_c_128_n N_VPWR_c_120_n
+ PM_SKY130_FD_SC_HS__INV_4%VPWR
x_PM_SKY130_FD_SC_HS__INV_4%Y N_Y_M1000_s N_Y_M1006_s N_Y_M1001_d N_Y_M1003_d
+ N_Y_c_168_n N_Y_c_164_n N_Y_c_157_n N_Y_c_158_n N_Y_c_159_n N_Y_c_184_n
+ N_Y_c_165_n N_Y_c_160_n N_Y_c_161_n N_Y_c_166_n N_Y_c_196_n N_Y_c_162_n Y
+ PM_SKY130_FD_SC_HS__INV_4%Y
x_PM_SKY130_FD_SC_HS__INV_4%VGND N_VGND_M1000_d N_VGND_M1005_d N_VGND_M1007_d
+ N_VGND_c_232_n N_VGND_c_233_n N_VGND_c_234_n N_VGND_c_235_n N_VGND_c_236_n
+ VGND N_VGND_c_237_n N_VGND_c_238_n N_VGND_c_239_n N_VGND_c_240_n
+ PM_SKY130_FD_SC_HS__INV_4%VGND
cc_1 VNB N_A_M1000_g 0.0314974f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=0.74
cc_2 VNB N_A_M1005_g 0.0238067f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=0.74
cc_3 VNB N_A_M1006_g 0.0238475f $X=-0.19 $Y=-0.245 $X2=1.475 $Y2=0.74
cc_4 VNB N_A_M1007_g 0.0261506f $X=-0.19 $Y=-0.245 $X2=1.905 $Y2=0.74
cc_5 VNB A 0.0177331f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=1.58
cc_6 VNB N_A_c_48_n 0.0763371f $X=-0.19 $Y=-0.245 $X2=1.89 $Y2=1.557
cc_7 VNB N_VPWR_c_120_n 0.103974f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=1.515
cc_8 VNB N_Y_c_157_n 0.00253214f $X=-0.19 $Y=-0.245 $X2=1.475 $Y2=0.74
cc_9 VNB N_Y_c_158_n 0.0035469f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_Y_c_159_n 0.00281969f $X=-0.19 $Y=-0.245 $X2=1.89 $Y2=1.765
cc_11 VNB N_Y_c_160_n 0.00179819f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.58
cc_12 VNB N_Y_c_161_n 0.0108018f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_Y_c_162_n 0.00127131f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=1.515
cc_14 VNB Y 0.0239872f $X=-0.19 $Y=-0.245 $X2=1.44 $Y2=1.557
cc_15 VNB N_VGND_c_232_n 0.0122168f $X=-0.19 $Y=-0.245 $X2=0.99 $Y2=2.4
cc_16 VNB N_VGND_c_233_n 0.0453501f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=0.74
cc_17 VNB N_VGND_c_234_n 0.00497255f $X=-0.19 $Y=-0.245 $X2=1.44 $Y2=2.4
cc_18 VNB N_VGND_c_235_n 0.0120272f $X=-0.19 $Y=-0.245 $X2=1.475 $Y2=1.35
cc_19 VNB N_VGND_c_236_n 0.0276369f $X=-0.19 $Y=-0.245 $X2=1.475 $Y2=0.74
cc_20 VNB N_VGND_c_237_n 0.016883f $X=-0.19 $Y=-0.245 $X2=1.89 $Y2=2.4
cc_21 VNB N_VGND_c_238_n 0.0169227f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_22 VNB N_VGND_c_239_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=1.557
cc_23 VNB N_VGND_c_240_n 0.160619f $X=-0.19 $Y=-0.245 $X2=0.99 $Y2=1.557
cc_24 VPB N_A_c_49_n 0.0179811f $X=-0.19 $Y=1.66 $X2=0.54 $Y2=1.765
cc_25 VPB N_A_c_50_n 0.0155127f $X=-0.19 $Y=1.66 $X2=0.99 $Y2=1.765
cc_26 VPB N_A_c_51_n 0.0155104f $X=-0.19 $Y=1.66 $X2=1.44 $Y2=1.765
cc_27 VPB N_A_c_52_n 0.0163707f $X=-0.19 $Y=1.66 $X2=1.89 $Y2=1.765
cc_28 VPB A 0.0196802f $X=-0.19 $Y=1.66 $X2=1.595 $Y2=1.58
cc_29 VPB N_A_c_48_n 0.0481502f $X=-0.19 $Y=1.66 $X2=1.89 $Y2=1.557
cc_30 VPB N_VPWR_c_121_n 0.0117686f $X=-0.19 $Y=1.66 $X2=0.99 $Y2=2.4
cc_31 VPB N_VPWR_c_122_n 0.0495873f $X=-0.19 $Y=1.66 $X2=0.995 $Y2=0.74
cc_32 VPB N_VPWR_c_123_n 0.0206041f $X=-0.19 $Y=1.66 $X2=1.44 $Y2=2.4
cc_33 VPB N_VPWR_c_124_n 0.00799266f $X=-0.19 $Y=1.66 $X2=1.475 $Y2=0.74
cc_34 VPB N_VPWR_c_125_n 0.0108116f $X=-0.19 $Y=1.66 $X2=1.89 $Y2=1.765
cc_35 VPB N_VPWR_c_126_n 0.0370539f $X=-0.19 $Y=1.66 $X2=1.89 $Y2=2.4
cc_36 VPB N_VPWR_c_127_n 0.0206041f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_37 VPB N_VPWR_c_128_n 0.00324402f $X=-0.19 $Y=1.66 $X2=0.525 $Y2=1.557
cc_38 VPB N_VPWR_c_120_n 0.0615795f $X=-0.19 $Y=1.66 $X2=0.615 $Y2=1.515
cc_39 VPB N_Y_c_164_n 0.00257348f $X=-0.19 $Y=1.66 $X2=1.44 $Y2=1.765
cc_40 VPB N_Y_c_165_n 0.00257348f $X=-0.19 $Y=1.66 $X2=1.905 $Y2=0.74
cc_41 VPB N_Y_c_166_n 0.00714919f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_42 VPB Y 0.0129845f $X=-0.19 $Y=1.66 $X2=1.44 $Y2=1.557
cc_43 N_A_c_49_n N_VPWR_c_122_n 0.00831454f $X=0.54 $Y=1.765 $X2=0 $Y2=0
cc_44 A N_VPWR_c_122_n 0.0219562f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_45 N_A_c_49_n N_VPWR_c_123_n 0.00445602f $X=0.54 $Y=1.765 $X2=0 $Y2=0
cc_46 N_A_c_50_n N_VPWR_c_123_n 0.00445602f $X=0.99 $Y=1.765 $X2=0 $Y2=0
cc_47 N_A_c_50_n N_VPWR_c_124_n 0.00486623f $X=0.99 $Y=1.765 $X2=0 $Y2=0
cc_48 N_A_c_51_n N_VPWR_c_124_n 0.00486623f $X=1.44 $Y=1.765 $X2=0 $Y2=0
cc_49 N_A_c_52_n N_VPWR_c_126_n 0.00714506f $X=1.89 $Y=1.765 $X2=0 $Y2=0
cc_50 N_A_c_51_n N_VPWR_c_127_n 0.00445602f $X=1.44 $Y=1.765 $X2=0 $Y2=0
cc_51 N_A_c_52_n N_VPWR_c_127_n 0.00445602f $X=1.89 $Y=1.765 $X2=0 $Y2=0
cc_52 N_A_c_49_n N_VPWR_c_120_n 0.00861194f $X=0.54 $Y=1.765 $X2=0 $Y2=0
cc_53 N_A_c_50_n N_VPWR_c_120_n 0.00857589f $X=0.99 $Y=1.765 $X2=0 $Y2=0
cc_54 N_A_c_51_n N_VPWR_c_120_n 0.00857589f $X=1.44 $Y=1.765 $X2=0 $Y2=0
cc_55 N_A_c_52_n N_VPWR_c_120_n 0.008611f $X=1.89 $Y=1.765 $X2=0 $Y2=0
cc_56 N_A_c_49_n N_Y_c_168_n 0.00203651f $X=0.54 $Y=1.765 $X2=0 $Y2=0
cc_57 N_A_c_50_n N_Y_c_168_n 4.27055e-19 $X=0.99 $Y=1.765 $X2=0 $Y2=0
cc_58 A N_Y_c_168_n 0.0237598f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_59 N_A_c_48_n N_Y_c_168_n 0.00144444f $X=1.89 $Y=1.557 $X2=0 $Y2=0
cc_60 N_A_c_49_n N_Y_c_164_n 0.00960826f $X=0.54 $Y=1.765 $X2=0 $Y2=0
cc_61 N_A_c_50_n N_Y_c_164_n 0.0103431f $X=0.99 $Y=1.765 $X2=0 $Y2=0
cc_62 N_A_c_51_n N_Y_c_164_n 6.45594e-19 $X=1.44 $Y=1.765 $X2=0 $Y2=0
cc_63 N_A_M1000_g N_Y_c_157_n 4.73925e-19 $X=0.525 $Y=0.74 $X2=0 $Y2=0
cc_64 N_A_M1005_g N_Y_c_157_n 4.39117e-19 $X=0.995 $Y=0.74 $X2=0 $Y2=0
cc_65 N_A_M1005_g N_Y_c_158_n 0.0133424f $X=0.995 $Y=0.74 $X2=0 $Y2=0
cc_66 N_A_M1006_g N_Y_c_158_n 0.0141141f $X=1.475 $Y=0.74 $X2=0 $Y2=0
cc_67 A N_Y_c_158_n 0.0555696f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_68 N_A_c_48_n N_Y_c_158_n 0.00336308f $X=1.89 $Y=1.557 $X2=0 $Y2=0
cc_69 N_A_M1000_g N_Y_c_159_n 0.00187357f $X=0.525 $Y=0.74 $X2=0 $Y2=0
cc_70 A N_Y_c_159_n 0.021475f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_71 N_A_c_48_n N_Y_c_159_n 0.00326139f $X=1.89 $Y=1.557 $X2=0 $Y2=0
cc_72 N_A_c_50_n N_Y_c_184_n 0.0120074f $X=0.99 $Y=1.765 $X2=0 $Y2=0
cc_73 N_A_c_51_n N_Y_c_184_n 0.0120074f $X=1.44 $Y=1.765 $X2=0 $Y2=0
cc_74 A N_Y_c_184_n 0.0393875f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_75 N_A_c_48_n N_Y_c_184_n 0.00131212f $X=1.89 $Y=1.557 $X2=0 $Y2=0
cc_76 N_A_c_50_n N_Y_c_165_n 6.45594e-19 $X=0.99 $Y=1.765 $X2=0 $Y2=0
cc_77 N_A_c_51_n N_Y_c_165_n 0.0103431f $X=1.44 $Y=1.765 $X2=0 $Y2=0
cc_78 N_A_c_52_n N_Y_c_165_n 0.01498f $X=1.89 $Y=1.765 $X2=0 $Y2=0
cc_79 N_A_M1006_g N_Y_c_160_n 4.06088e-19 $X=1.475 $Y=0.74 $X2=0 $Y2=0
cc_80 N_A_M1007_g N_Y_c_160_n 3.92313e-19 $X=1.905 $Y=0.74 $X2=0 $Y2=0
cc_81 N_A_M1007_g N_Y_c_161_n 0.0190067f $X=1.905 $Y=0.74 $X2=0 $Y2=0
cc_82 A N_Y_c_161_n 0.00188044f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_83 N_A_c_52_n N_Y_c_166_n 0.0173803f $X=1.89 $Y=1.765 $X2=0 $Y2=0
cc_84 N_A_c_51_n N_Y_c_196_n 4.27055e-19 $X=1.44 $Y=1.765 $X2=0 $Y2=0
cc_85 N_A_c_52_n N_Y_c_196_n 9.50925e-19 $X=1.89 $Y=1.765 $X2=0 $Y2=0
cc_86 A N_Y_c_196_n 0.0219285f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_87 N_A_c_48_n N_Y_c_196_n 0.00144162f $X=1.89 $Y=1.557 $X2=0 $Y2=0
cc_88 A N_Y_c_162_n 0.0146029f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_89 N_A_c_48_n N_Y_c_162_n 0.00232957f $X=1.89 $Y=1.557 $X2=0 $Y2=0
cc_90 N_A_c_52_n Y 0.00696961f $X=1.89 $Y=1.765 $X2=0 $Y2=0
cc_91 N_A_M1007_g Y 0.0190395f $X=1.905 $Y=0.74 $X2=0 $Y2=0
cc_92 A Y 0.0266022f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_93 N_A_M1000_g N_VGND_c_233_n 0.00551504f $X=0.525 $Y=0.74 $X2=0 $Y2=0
cc_94 A N_VGND_c_233_n 0.0239925f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_95 N_A_M1000_g N_VGND_c_234_n 4.69274e-19 $X=0.525 $Y=0.74 $X2=0 $Y2=0
cc_96 N_A_M1005_g N_VGND_c_234_n 0.0104328f $X=0.995 $Y=0.74 $X2=0 $Y2=0
cc_97 N_A_M1006_g N_VGND_c_234_n 0.00223467f $X=1.475 $Y=0.74 $X2=0 $Y2=0
cc_98 N_A_M1006_g N_VGND_c_236_n 4.78723e-19 $X=1.475 $Y=0.74 $X2=0 $Y2=0
cc_99 N_A_M1007_g N_VGND_c_236_n 0.0121476f $X=1.905 $Y=0.74 $X2=0 $Y2=0
cc_100 N_A_M1000_g N_VGND_c_237_n 0.00461464f $X=0.525 $Y=0.74 $X2=0 $Y2=0
cc_101 N_A_M1005_g N_VGND_c_237_n 0.00383152f $X=0.995 $Y=0.74 $X2=0 $Y2=0
cc_102 N_A_M1006_g N_VGND_c_238_n 0.00461464f $X=1.475 $Y=0.74 $X2=0 $Y2=0
cc_103 N_A_M1007_g N_VGND_c_238_n 0.00383152f $X=1.905 $Y=0.74 $X2=0 $Y2=0
cc_104 N_A_M1000_g N_VGND_c_240_n 0.00911356f $X=0.525 $Y=0.74 $X2=0 $Y2=0
cc_105 N_A_M1005_g N_VGND_c_240_n 0.00757927f $X=0.995 $Y=0.74 $X2=0 $Y2=0
cc_106 N_A_M1006_g N_VGND_c_240_n 0.0090814f $X=1.475 $Y=0.74 $X2=0 $Y2=0
cc_107 N_A_M1007_g N_VGND_c_240_n 0.0075754f $X=1.905 $Y=0.74 $X2=0 $Y2=0
cc_108 N_VPWR_c_122_n N_Y_c_168_n 0.0121024f $X=0.315 $Y=2.115 $X2=0 $Y2=0
cc_109 N_VPWR_c_122_n N_Y_c_164_n 0.0576605f $X=0.315 $Y=2.115 $X2=0 $Y2=0
cc_110 N_VPWR_c_123_n N_Y_c_164_n 0.014552f $X=1.13 $Y=3.33 $X2=0 $Y2=0
cc_111 N_VPWR_c_124_n N_Y_c_164_n 0.0449718f $X=1.215 $Y=2.455 $X2=0 $Y2=0
cc_112 N_VPWR_c_120_n N_Y_c_164_n 0.0119791f $X=2.16 $Y=3.33 $X2=0 $Y2=0
cc_113 N_VPWR_M1002_s N_Y_c_184_n 0.00408911f $X=1.065 $Y=1.84 $X2=0 $Y2=0
cc_114 N_VPWR_c_124_n N_Y_c_184_n 0.0136682f $X=1.215 $Y=2.455 $X2=0 $Y2=0
cc_115 N_VPWR_c_124_n N_Y_c_165_n 0.0449718f $X=1.215 $Y=2.455 $X2=0 $Y2=0
cc_116 N_VPWR_c_126_n N_Y_c_165_n 0.0462948f $X=2.115 $Y=2.455 $X2=0 $Y2=0
cc_117 N_VPWR_c_127_n N_Y_c_165_n 0.014552f $X=2.03 $Y=3.33 $X2=0 $Y2=0
cc_118 N_VPWR_c_120_n N_Y_c_165_n 0.0119791f $X=2.16 $Y=3.33 $X2=0 $Y2=0
cc_119 N_VPWR_M1004_s N_Y_c_166_n 0.00477129f $X=1.965 $Y=1.84 $X2=0 $Y2=0
cc_120 N_VPWR_c_126_n N_Y_c_166_n 0.0218009f $X=2.115 $Y=2.455 $X2=0 $Y2=0
cc_121 N_VPWR_M1004_s Y 0.00194528f $X=1.965 $Y=1.84 $X2=0 $Y2=0
cc_122 N_Y_c_158_n N_VGND_M1005_d 0.00229612f $X=1.605 $Y=1.095 $X2=0 $Y2=0
cc_123 N_Y_c_161_n N_VGND_M1007_d 0.00309016f $X=2.045 $Y=1.095 $X2=0 $Y2=0
cc_124 N_Y_c_157_n N_VGND_c_233_n 0.00154841f $X=0.78 $Y=0.515 $X2=0 $Y2=0
cc_125 N_Y_c_159_n N_VGND_c_233_n 0.00167954f $X=0.865 $Y=1.095 $X2=0 $Y2=0
cc_126 N_Y_c_157_n N_VGND_c_234_n 0.0182902f $X=0.78 $Y=0.515 $X2=0 $Y2=0
cc_127 N_Y_c_158_n N_VGND_c_234_n 0.0194017f $X=1.605 $Y=1.095 $X2=0 $Y2=0
cc_128 N_Y_c_160_n N_VGND_c_234_n 0.00121793f $X=1.69 $Y=0.515 $X2=0 $Y2=0
cc_129 N_Y_c_160_n N_VGND_c_236_n 0.0182488f $X=1.69 $Y=0.515 $X2=0 $Y2=0
cc_130 N_Y_c_161_n N_VGND_c_236_n 0.0232152f $X=2.045 $Y=1.095 $X2=0 $Y2=0
cc_131 N_Y_c_157_n N_VGND_c_237_n 0.011066f $X=0.78 $Y=0.515 $X2=0 $Y2=0
cc_132 N_Y_c_160_n N_VGND_c_238_n 0.00749631f $X=1.69 $Y=0.515 $X2=0 $Y2=0
cc_133 N_Y_c_157_n N_VGND_c_240_n 0.00915947f $X=0.78 $Y=0.515 $X2=0 $Y2=0
cc_134 N_Y_c_160_n N_VGND_c_240_n 0.0062048f $X=1.69 $Y=0.515 $X2=0 $Y2=0
