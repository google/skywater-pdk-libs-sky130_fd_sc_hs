* NGSPICE file created from sky130_fd_sc_hs__or4bb_4.ext - technology: sky130A

.subckt sky130_fd_sc_hs__or4bb_4 A B C_N D_N VGND VNB VPB VPWR X
M1000 VGND a_193_277# X VNB nlowvt w=740000u l=150000u
+  ad=2.0924e+12p pd=1.558e+07u as=6.919e+11p ps=4.83e+06u
M1001 a_1060_392# a_678_368# a_791_392# VPB pshort w=1e+06u l=150000u
+  ad=6.5e+11p pd=5.3e+06u as=8.9e+11p ps=7.78e+06u
M1002 a_791_392# a_678_368# a_1060_392# VPB pshort w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1003 VGND A a_193_277# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=1.4134e+12p ps=6.78e+06u
M1004 VGND D_N a_27_94# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=1.824e+11p ps=1.85e+06u
M1005 a_678_368# C_N VGND VNB nlowvt w=640000u l=150000u
+  ad=1.719e+11p pd=1.85e+06u as=0p ps=0u
M1006 a_678_368# C_N VPWR VPB pshort w=1e+06u l=150000u
+  ad=2.95e+11p pd=2.59e+06u as=1.65e+12p ps=1.178e+07u
M1007 a_193_277# B VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 X a_193_277# VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=9.856e+11p pd=6.24e+06u as=0p ps=0u
M1009 X a_193_277# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VPWR a_193_277# X VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_193_277# a_27_94# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VGND a_193_277# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VPWR D_N a_27_94# VPB pshort w=1e+06u l=150000u
+  ad=0p pd=0u as=2.95e+11p ps=2.59e+06u
M1014 X a_193_277# VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_1060_392# B a_1273_392# VPB pshort w=1e+06u l=150000u
+  ad=0p pd=0u as=8.9e+11p ps=7.78e+06u
M1016 a_1273_392# B a_1060_392# VPB pshort w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_1273_392# A VPWR VPB pshort w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 X a_193_277# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VPWR A a_1273_392# VPB pshort w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_193_277# a_27_94# a_791_392# VPB pshort w=1e+06u l=150000u
+  ad=3e+11p pd=2.6e+06u as=0p ps=0u
M1021 VGND a_678_368# a_193_277# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_791_392# a_27_94# a_193_277# VPB pshort w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 VPWR a_193_277# X VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

