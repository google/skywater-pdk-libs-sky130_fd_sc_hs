* File: sky130_fd_sc_hs__o2bb2ai_2.spice
* Created: Tue Sep  1 20:17:05 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hs__o2bb2ai_2.pex.spice"
.subckt sky130_fd_sc_hs__o2bb2ai_2  VNB VPB A1_N A2_N B1 B2 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* B2	B2
* B1	B1
* A2_N	A2_N
* A1_N	A1_N
* VPB	VPB
* VNB	VNB
MM1006 N_A_134_74#_M1006_d N_A1_N_M1006_g N_VGND_M1006_s VNB NLOWVT L=0.15
+ W=0.64 AD=0.0896 AS=0.2272 PD=0.92 PS=1.99 NRD=0 NRS=13.116 M=1 R=4.26667
+ SA=75000.3 SB=75001.6 A=0.096 P=1.58 MULT=1
MM1007 N_A_133_387#_M1007_d N_A2_N_M1007_g N_A_134_74#_M1006_d VNB NLOWVT L=0.15
+ W=0.64 AD=0.1136 AS=0.0896 PD=0.995 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.7 SB=75001.1 A=0.096 P=1.58 MULT=1
MM1019 N_A_133_387#_M1007_d N_A2_N_M1019_g N_A_134_74#_M1019_s VNB NLOWVT L=0.15
+ W=0.64 AD=0.1136 AS=0.0896 PD=0.995 PS=0.92 NRD=14.052 NRS=0 M=1 R=4.26667
+ SA=75001.2 SB=75000.6 A=0.096 P=1.58 MULT=1
MM1012 N_A_134_74#_M1019_s N_A1_N_M1012_g N_VGND_M1012_s VNB NLOWVT L=0.15
+ W=0.64 AD=0.0896 AS=0.1824 PD=0.92 PS=1.85 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75001.6 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1000 N_Y_M1000_d N_A_133_387#_M1000_g N_A_518_74#_M1000_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.2109 PD=1.02 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75002.5 A=0.111 P=1.78 MULT=1
MM1005 N_Y_M1000_d N_A_133_387#_M1005_g N_A_518_74#_M1005_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.1147 PD=1.02 PS=1.05 NRD=0 NRS=4.86 M=1 R=4.93333
+ SA=75000.6 SB=75002.1 A=0.111 P=1.78 MULT=1
MM1008 N_A_518_74#_M1005_s N_B1_M1008_g N_VGND_M1008_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1147 AS=0.1295 PD=1.05 PS=1.09 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75001.1
+ SB=75001.6 A=0.111 P=1.78 MULT=1
MM1002 N_VGND_M1008_s N_B2_M1002_g N_A_518_74#_M1002_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1295 AS=0.1221 PD=1.09 PS=1.07 NRD=0 NRS=4.044 M=1 R=4.93333 SA=75001.6
+ SB=75001.1 A=0.111 P=1.78 MULT=1
MM1015 N_VGND_M1015_d N_B2_M1015_g N_A_518_74#_M1002_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.10915 AS=0.1221 PD=1.035 PS=1.07 NRD=0.804 NRS=4.044 M=1 R=4.93333
+ SA=75002.1 SB=75000.7 A=0.111 P=1.78 MULT=1
MM1016 N_A_518_74#_M1016_d N_B1_M1016_g N_VGND_M1015_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.10915 PD=2.05 PS=1.035 NRD=0 NRS=1.62 M=1 R=4.93333 SA=75002.5
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1004 N_A_133_387#_M1004_d N_A1_N_M1004_g N_VPWR_M1004_s VPB PSHORT L=0.15
+ W=0.84 AD=0.126 AS=0.3801 PD=1.14 PS=2.86 NRD=0 NRS=93.2204 M=1 R=5.6
+ SA=75000.3 SB=75004.5 A=0.126 P=1.98 MULT=1
MM1003 N_A_133_387#_M1004_d N_A2_N_M1003_g N_VPWR_M1003_s VPB PSHORT L=0.15
+ W=0.84 AD=0.126 AS=0.232925 PD=1.14 PS=1.555 NRD=2.3443 NRS=52.1262 M=1 R=5.6
+ SA=75000.8 SB=75004 A=0.126 P=1.98 MULT=1
MM1009 N_A_133_387#_M1009_d N_A2_N_M1009_g N_VPWR_M1003_s VPB PSHORT L=0.15
+ W=0.84 AD=0.172312 AS=0.232925 PD=1.33 PS=1.555 NRD=4.6886 NRS=52.1262 M=1
+ R=5.6 SA=75001.4 SB=75003.4 A=0.126 P=1.98 MULT=1
MM1018 N_A_133_387#_M1009_d N_A1_N_M1018_g N_VPWR_M1018_s VPB PSHORT L=0.15
+ W=0.84 AD=0.172312 AS=0.2322 PD=1.33 PS=1.42714 NRD=22.261 NRS=58.6272 M=1
+ R=5.6 SA=75001.7 SB=75003.3 A=0.126 P=1.98 MULT=1
MM1001 N_VPWR_M1018_s N_A_133_387#_M1001_g N_Y_M1001_s VPB PSHORT L=0.15 W=1.12
+ AD=0.3096 AS=0.1764 PD=1.90286 PS=1.435 NRD=2.6201 NRS=1.7533 M=1 R=7.46667
+ SA=75001.9 SB=75002.6 A=0.168 P=2.54 MULT=1
MM1014 N_VPWR_M1014_d N_A_133_387#_M1014_g N_Y_M1001_s VPB PSHORT L=0.15 W=1.12
+ AD=0.2184 AS=0.1764 PD=1.51 PS=1.435 NRD=7.8997 NRS=4.3931 M=1 R=7.46667
+ SA=75002.3 SB=75002.1 A=0.168 P=2.54 MULT=1
MM1010 N_A_796_368#_M1010_d N_B1_M1010_g N_VPWR_M1014_d VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.2184 PD=1.42 PS=1.51 NRD=1.7533 NRS=11.426 M=1 R=7.46667
+ SA=75002.9 SB=75001.6 A=0.168 P=2.54 MULT=1
MM1011 N_Y_M1011_d N_B2_M1011_g N_A_796_368#_M1010_d VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75003.3 SB=75001.1 A=0.168 P=2.54 MULT=1
MM1013 N_Y_M1011_d N_B2_M1013_g N_A_796_368#_M1013_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75003.8 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1017 N_A_796_368#_M1013_s N_B1_M1017_g N_VPWR_M1017_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.3304 PD=1.42 PS=2.83 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75004.2 SB=75000.2 A=0.168 P=2.54 MULT=1
DX20_noxref VNB VPB NWDIODE A=11.4204 P=16
c_55 VNB 0 1.39855e-19 $X=0 $Y=0
*
.include "sky130_fd_sc_hs__o2bb2ai_2.pxi.spice"
*
.ends
*
*
