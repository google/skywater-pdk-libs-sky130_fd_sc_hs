* File: sky130_fd_sc_hs__mux2_1.pxi.spice
* Created: Tue Sep  1 20:07:35 2020
* 
x_PM_SKY130_FD_SC_HS__MUX2_1%S N_S_M1003_g N_S_c_78_n N_S_M1005_g N_S_c_79_n
+ N_S_M1000_g N_S_M1006_g N_S_c_74_n N_S_c_75_n N_S_c_76_n S N_S_c_77_n
+ PM_SKY130_FD_SC_HS__MUX2_1%S
x_PM_SKY130_FD_SC_HS__MUX2_1%A1 N_A1_M1004_g N_A1_c_129_n N_A1_M1011_g
+ N_A1_c_130_n N_A1_c_141_p N_A1_c_166_p N_A1_c_131_n N_A1_c_132_n A1 A1
+ N_A1_c_134_n N_A1_c_157_p PM_SKY130_FD_SC_HS__MUX2_1%A1
x_PM_SKY130_FD_SC_HS__MUX2_1%A0 N_A0_c_191_n N_A0_M1002_g N_A0_c_192_n
+ N_A0_M1001_g A0 PM_SKY130_FD_SC_HS__MUX2_1%A0
x_PM_SKY130_FD_SC_HS__MUX2_1%A_27_112# N_A_27_112#_M1003_s N_A_27_112#_M1005_s
+ N_A_27_112#_M1008_g N_A_27_112#_c_221_n N_A_27_112#_M1007_g
+ N_A_27_112#_c_222_n N_A_27_112#_c_223_n N_A_27_112#_c_239_n
+ N_A_27_112#_c_229_n N_A_27_112#_c_230_n N_A_27_112#_c_231_n
+ N_A_27_112#_c_224_n N_A_27_112#_c_225_n N_A_27_112#_c_233_n
+ N_A_27_112#_c_226_n PM_SKY130_FD_SC_HS__MUX2_1%A_27_112#
x_PM_SKY130_FD_SC_HS__MUX2_1%A_304_74# N_A_304_74#_M1004_d N_A_304_74#_M1002_d
+ N_A_304_74#_c_310_n N_A_304_74#_M1010_g N_A_304_74#_M1009_g
+ N_A_304_74#_c_312_n N_A_304_74#_c_406_p N_A_304_74#_c_319_n
+ N_A_304_74#_c_324_n N_A_304_74#_c_339_n N_A_304_74#_c_400_p
+ N_A_304_74#_c_346_n N_A_304_74#_c_347_n N_A_304_74#_c_313_n
+ N_A_304_74#_c_314_n N_A_304_74#_c_315_n N_A_304_74#_c_328_n
+ N_A_304_74#_c_316_n PM_SKY130_FD_SC_HS__MUX2_1%A_304_74#
x_PM_SKY130_FD_SC_HS__MUX2_1%VPWR N_VPWR_M1005_d N_VPWR_M1007_d N_VPWR_c_413_n
+ N_VPWR_c_414_n N_VPWR_c_415_n N_VPWR_c_416_n VPWR N_VPWR_c_417_n
+ N_VPWR_c_412_n N_VPWR_c_419_n PM_SKY130_FD_SC_HS__MUX2_1%VPWR
x_PM_SKY130_FD_SC_HS__MUX2_1%X N_X_M1009_d N_X_M1010_d N_X_c_457_n N_X_c_458_n X
+ X X N_X_c_461_n N_X_c_459_n X PM_SKY130_FD_SC_HS__MUX2_1%X
x_PM_SKY130_FD_SC_HS__MUX2_1%VGND N_VGND_M1003_d N_VGND_M1008_d N_VGND_c_481_n
+ N_VGND_c_482_n N_VGND_c_483_n N_VGND_c_484_n N_VGND_c_485_n N_VGND_c_486_n
+ VGND N_VGND_c_487_n N_VGND_c_488_n N_VGND_c_489_n N_VGND_c_490_n
+ PM_SKY130_FD_SC_HS__MUX2_1%VGND
cc_1 VNB N_S_M1003_g 0.0307509f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.835
cc_2 VNB N_S_M1006_g 0.0246926f $X=-0.19 $Y=-0.245 $X2=1.055 $Y2=0.74
cc_3 VNB N_S_c_74_n 0.01399f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.557
cc_4 VNB N_S_c_75_n 0.0184644f $X=-0.19 $Y=-0.245 $X2=0.95 $Y2=1.515
cc_5 VNB N_S_c_76_n 0.0111302f $X=-0.19 $Y=-0.245 $X2=1.04 $Y2=1.557
cc_6 VNB N_S_c_77_n 0.00177531f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=1.515
cc_7 VNB N_A1_c_129_n 0.0439773f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_A1_c_130_n 0.00111648f $X=-0.19 $Y=-0.245 $X2=1.04 $Y2=1.765
cc_9 VNB N_A1_c_131_n 0.0318272f $X=-0.19 $Y=-0.245 $X2=1.055 $Y2=0.74
cc_10 VNB N_A1_c_132_n 0.00427166f $X=-0.19 $Y=-0.245 $X2=0.595 $Y2=1.515
cc_11 VNB A1 0.00811709f $X=-0.19 $Y=-0.245 $X2=0.95 $Y2=1.515
cc_12 VNB N_A1_c_134_n 0.0189248f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=1.515
cc_13 VNB N_A0_c_191_n 0.037533f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.35
cc_14 VNB N_A0_c_192_n 0.0240239f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB A0 0.00774979f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.26
cc_16 VNB N_A_27_112#_M1008_g 0.0298799f $X=-0.19 $Y=-0.245 $X2=1.04 $Y2=2.34
cc_17 VNB N_A_27_112#_c_221_n 0.0303892f $X=-0.19 $Y=-0.245 $X2=1.055 $Y2=1.35
cc_18 VNB N_A_27_112#_c_222_n 0.0197085f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.557
cc_19 VNB N_A_27_112#_c_223_n 0.0250637f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_20 VNB N_A_27_112#_c_224_n 3.05599e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_27_112#_c_225_n 0.0116048f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_27_112#_c_226_n 0.00555683f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_304_74#_c_310_n 0.0370044f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.26
cc_24 VNB N_A_304_74#_M1009_g 0.0299476f $X=-0.19 $Y=-0.245 $X2=1.055 $Y2=0.74
cc_25 VNB N_A_304_74#_c_312_n 0.00662024f $X=-0.19 $Y=-0.245 $X2=0.595 $Y2=1.515
cc_26 VNB N_A_304_74#_c_313_n 0.00440116f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_304_74#_c_314_n 0.00102356f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_304_74#_c_315_n 0.00294361f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_304_74#_c_316_n 0.00564651f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_VPWR_c_412_n 0.183584f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_X_c_457_n 0.0267746f $X=-0.19 $Y=-0.245 $X2=1.04 $Y2=2.34
cc_32 VNB N_X_c_458_n 0.014426f $X=-0.19 $Y=-0.245 $X2=1.055 $Y2=0.74
cc_33 VNB N_X_c_459_n 0.0248128f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_481_n 0.0135512f $X=-0.19 $Y=-0.245 $X2=1.04 $Y2=1.765
cc_35 VNB N_VGND_c_482_n 0.00191515f $X=-0.19 $Y=-0.245 $X2=1.055 $Y2=1.35
cc_36 VNB N_VGND_c_483_n 0.00993982f $X=-0.19 $Y=-0.245 $X2=0.595 $Y2=1.515
cc_37 VNB N_VGND_c_484_n 6.638e-19 $X=-0.19 $Y=-0.245 $X2=1.04 $Y2=1.557
cc_38 VNB N_VGND_c_485_n 0.0585899f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=1.515
cc_39 VNB N_VGND_c_486_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=1.515
cc_40 VNB N_VGND_c_487_n 0.0202692f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_488_n 0.0213848f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_489_n 0.261293f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_490_n 0.00711965f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VPB N_S_c_78_n 0.0195831f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.765
cc_45 VPB N_S_c_79_n 0.017545f $X=-0.19 $Y=1.66 $X2=1.04 $Y2=1.765
cc_46 VPB N_S_c_74_n 0.00659712f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.557
cc_47 VPB N_S_c_75_n 0.0109102f $X=-0.19 $Y=1.66 $X2=0.95 $Y2=1.515
cc_48 VPB N_S_c_76_n 0.00753269f $X=-0.19 $Y=1.66 $X2=1.04 $Y2=1.557
cc_49 VPB N_S_c_77_n 0.00345632f $X=-0.19 $Y=1.66 $X2=0.67 $Y2=1.515
cc_50 VPB N_A1_c_129_n 0.024612f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_51 VPB N_A0_c_191_n 0.0264167f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.35
cc_52 VPB N_A_27_112#_c_221_n 0.0238634f $X=-0.19 $Y=1.66 $X2=1.055 $Y2=1.35
cc_53 VPB N_A_27_112#_c_223_n 0.0126863f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_54 VPB N_A_27_112#_c_229_n 0.00164517f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_55 VPB N_A_27_112#_c_230_n 0.0547494f $X=-0.19 $Y=1.66 $X2=0.67 $Y2=1.665
cc_56 VPB N_A_27_112#_c_231_n 0.00361939f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_57 VPB N_A_27_112#_c_224_n 0.00257182f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_58 VPB N_A_27_112#_c_233_n 0.0332575f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_59 VPB N_A_304_74#_c_310_n 0.029883f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.26
cc_60 VPB N_A_304_74#_c_312_n 0.00202686f $X=-0.19 $Y=1.66 $X2=0.595 $Y2=1.515
cc_61 VPB N_A_304_74#_c_319_n 0.024444f $X=-0.19 $Y=1.66 $X2=1.04 $Y2=1.557
cc_62 VPB N_VPWR_c_413_n 0.0196908f $X=-0.19 $Y=1.66 $X2=1.055 $Y2=1.35
cc_63 VPB N_VPWR_c_414_n 0.015165f $X=-0.19 $Y=1.66 $X2=0.595 $Y2=1.515
cc_64 VPB N_VPWR_c_415_n 0.0550508f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_65 VPB N_VPWR_c_416_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0.67 $Y2=1.515
cc_66 VPB N_VPWR_c_417_n 0.020838f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_67 VPB N_VPWR_c_412_n 0.0842263f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_68 VPB N_VPWR_c_419_n 0.0276744f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_69 VPB X 0.0444516f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_70 VPB N_X_c_461_n 0.017092f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_71 VPB N_X_c_459_n 0.00782691f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_72 N_S_M1006_g N_A1_c_130_n 2.24893e-19 $X=1.055 $Y=0.74 $X2=0 $Y2=0
cc_73 N_S_M1006_g N_A1_c_131_n 0.0207911f $X=1.055 $Y=0.74 $X2=0 $Y2=0
cc_74 N_S_M1006_g N_A1_c_132_n 3.74625e-19 $X=1.055 $Y=0.74 $X2=0 $Y2=0
cc_75 N_S_M1006_g N_A1_c_134_n 0.0476408f $X=1.055 $Y=0.74 $X2=0 $Y2=0
cc_76 N_S_M1003_g N_A_27_112#_c_222_n 0.00684278f $X=0.495 $Y=0.835 $X2=0 $Y2=0
cc_77 N_S_M1003_g N_A_27_112#_c_223_n 0.00602767f $X=0.495 $Y=0.835 $X2=0 $Y2=0
cc_78 N_S_c_78_n N_A_27_112#_c_223_n 0.00390035f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_79 N_S_c_74_n N_A_27_112#_c_223_n 0.0111274f $X=0.505 $Y=1.557 $X2=0 $Y2=0
cc_80 N_S_c_77_n N_A_27_112#_c_223_n 0.026603f $X=0.67 $Y=1.515 $X2=0 $Y2=0
cc_81 N_S_c_78_n N_A_27_112#_c_239_n 0.0143396f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_82 N_S_c_79_n N_A_27_112#_c_239_n 0.0175246f $X=1.04 $Y=1.765 $X2=0 $Y2=0
cc_83 N_S_c_75_n N_A_27_112#_c_239_n 0.00420822f $X=0.95 $Y=1.515 $X2=0 $Y2=0
cc_84 N_S_c_77_n N_A_27_112#_c_239_n 0.0164124f $X=0.67 $Y=1.515 $X2=0 $Y2=0
cc_85 N_S_c_79_n N_A_27_112#_c_229_n 0.0134005f $X=1.04 $Y=1.765 $X2=0 $Y2=0
cc_86 N_S_c_79_n N_A_27_112#_c_231_n 0.00153607f $X=1.04 $Y=1.765 $X2=0 $Y2=0
cc_87 N_S_M1003_g N_A_27_112#_c_225_n 0.00496391f $X=0.495 $Y=0.835 $X2=0 $Y2=0
cc_88 N_S_c_74_n N_A_27_112#_c_225_n 2.10625e-19 $X=0.505 $Y=1.557 $X2=0 $Y2=0
cc_89 N_S_c_78_n N_A_27_112#_c_233_n 0.0117673f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_90 N_S_c_79_n N_A_27_112#_c_233_n 0.00107648f $X=1.04 $Y=1.765 $X2=0 $Y2=0
cc_91 N_S_M1003_g N_A_304_74#_c_312_n 0.00123241f $X=0.495 $Y=0.835 $X2=0 $Y2=0
cc_92 N_S_M1006_g N_A_304_74#_c_312_n 0.00908273f $X=1.055 $Y=0.74 $X2=0 $Y2=0
cc_93 N_S_c_76_n N_A_304_74#_c_312_n 0.0121272f $X=1.04 $Y=1.557 $X2=0 $Y2=0
cc_94 N_S_c_77_n N_A_304_74#_c_312_n 0.0265523f $X=0.67 $Y=1.515 $X2=0 $Y2=0
cc_95 N_S_c_78_n N_A_304_74#_c_324_n 6.00232e-19 $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_96 N_S_c_79_n N_A_304_74#_c_324_n 0.00785206f $X=1.04 $Y=1.765 $X2=0 $Y2=0
cc_97 N_S_c_76_n N_A_304_74#_c_324_n 0.00214455f $X=1.04 $Y=1.557 $X2=0 $Y2=0
cc_98 N_S_c_77_n N_A_304_74#_c_324_n 0.00499246f $X=0.67 $Y=1.515 $X2=0 $Y2=0
cc_99 N_S_M1006_g N_A_304_74#_c_328_n 0.00748628f $X=1.055 $Y=0.74 $X2=0 $Y2=0
cc_100 N_S_c_78_n N_VPWR_c_413_n 0.00579539f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_101 N_S_c_79_n N_VPWR_c_413_n 0.0108017f $X=1.04 $Y=1.765 $X2=0 $Y2=0
cc_102 N_S_c_79_n N_VPWR_c_415_n 0.00443511f $X=1.04 $Y=1.765 $X2=0 $Y2=0
cc_103 N_S_c_78_n N_VPWR_c_412_n 0.00462577f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_104 N_S_c_79_n N_VPWR_c_412_n 0.00460931f $X=1.04 $Y=1.765 $X2=0 $Y2=0
cc_105 N_S_c_78_n N_VPWR_c_419_n 0.00393873f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_106 N_S_M1003_g N_VGND_c_481_n 0.00480382f $X=0.495 $Y=0.835 $X2=0 $Y2=0
cc_107 N_S_M1006_g N_VGND_c_481_n 0.006896f $X=1.055 $Y=0.74 $X2=0 $Y2=0
cc_108 N_S_M1006_g N_VGND_c_482_n 0.00352246f $X=1.055 $Y=0.74 $X2=0 $Y2=0
cc_109 N_S_c_75_n N_VGND_c_482_n 0.00133397f $X=0.95 $Y=1.515 $X2=0 $Y2=0
cc_110 N_S_c_77_n N_VGND_c_482_n 0.0147823f $X=0.67 $Y=1.515 $X2=0 $Y2=0
cc_111 N_S_M1006_g N_VGND_c_484_n 0.00308901f $X=1.055 $Y=0.74 $X2=0 $Y2=0
cc_112 N_S_c_75_n N_VGND_c_484_n 0.00145997f $X=0.95 $Y=1.515 $X2=0 $Y2=0
cc_113 N_S_M1006_g N_VGND_c_485_n 0.00383152f $X=1.055 $Y=0.74 $X2=0 $Y2=0
cc_114 N_S_M1003_g N_VGND_c_487_n 0.0043356f $X=0.495 $Y=0.835 $X2=0 $Y2=0
cc_115 N_S_M1003_g N_VGND_c_489_n 0.00487769f $X=0.495 $Y=0.835 $X2=0 $Y2=0
cc_116 N_S_M1006_g N_VGND_c_489_n 0.00384101f $X=1.055 $Y=0.74 $X2=0 $Y2=0
cc_117 N_A1_c_129_n N_A0_c_191_n 0.0477381f $X=2.545 $Y=1.765 $X2=-0.19
+ $Y2=-0.245
cc_118 N_A1_c_141_p N_A0_c_191_n 9.71665e-19 $X=2.455 $Y=0.895 $X2=-0.19
+ $Y2=-0.245
cc_119 N_A1_c_131_n N_A0_c_191_n 0.0214266f $X=1.51 $Y=1.385 $X2=-0.19
+ $Y2=-0.245
cc_120 N_A1_c_132_n N_A0_c_191_n 0.00113394f $X=1.6 $Y=1.385 $X2=-0.19
+ $Y2=-0.245
cc_121 A1 N_A0_c_191_n 3.71725e-19 $X=2.555 $Y=0.84 $X2=-0.19 $Y2=-0.245
cc_122 N_A1_c_130_n N_A0_c_192_n 0.00368858f $X=1.6 $Y=1.22 $X2=0 $Y2=0
cc_123 N_A1_c_141_p N_A0_c_192_n 0.013623f $X=2.455 $Y=0.895 $X2=0 $Y2=0
cc_124 A1 N_A0_c_192_n 0.00714134f $X=2.555 $Y=0.84 $X2=0 $Y2=0
cc_125 N_A1_c_134_n N_A0_c_192_n 0.0195334f $X=1.51 $Y=1.22 $X2=0 $Y2=0
cc_126 N_A1_c_129_n A0 0.00202561f $X=2.545 $Y=1.765 $X2=0 $Y2=0
cc_127 N_A1_c_130_n A0 0.00280644f $X=1.6 $Y=1.22 $X2=0 $Y2=0
cc_128 N_A1_c_141_p A0 0.0226197f $X=2.455 $Y=0.895 $X2=0 $Y2=0
cc_129 N_A1_c_131_n A0 4.04959e-19 $X=1.51 $Y=1.385 $X2=0 $Y2=0
cc_130 N_A1_c_132_n A0 0.0235137f $X=1.6 $Y=1.385 $X2=0 $Y2=0
cc_131 A1 A0 0.0285677f $X=2.555 $Y=0.84 $X2=0 $Y2=0
cc_132 N_A1_c_129_n N_A_27_112#_M1008_g 0.0176872f $X=2.545 $Y=1.765 $X2=0 $Y2=0
cc_133 A1 N_A_27_112#_M1008_g 0.00411883f $X=2.555 $Y=0.84 $X2=0 $Y2=0
cc_134 N_A1_c_157_p N_A_27_112#_M1008_g 0.0011484f $X=2.62 $Y=0.98 $X2=0 $Y2=0
cc_135 N_A1_c_129_n N_A_27_112#_c_221_n 0.0345836f $X=2.545 $Y=1.765 $X2=0 $Y2=0
cc_136 A1 N_A_27_112#_c_221_n 2.52902e-19 $X=2.555 $Y=0.84 $X2=0 $Y2=0
cc_137 N_A1_c_129_n N_A_27_112#_c_230_n 0.0119628f $X=2.545 $Y=1.765 $X2=0 $Y2=0
cc_138 N_A1_c_129_n N_A_27_112#_c_224_n 0.0125725f $X=2.545 $Y=1.765 $X2=0 $Y2=0
cc_139 N_A1_c_129_n N_A_27_112#_c_226_n 0.0035428f $X=2.545 $Y=1.765 $X2=0 $Y2=0
cc_140 A1 N_A_27_112#_c_226_n 0.0184934f $X=2.555 $Y=0.84 $X2=0 $Y2=0
cc_141 N_A1_c_130_n N_A_304_74#_M1004_d 0.00178335f $X=1.6 $Y=1.22 $X2=-0.19
+ $Y2=-0.245
cc_142 N_A1_c_141_p N_A_304_74#_M1004_d 0.0138145f $X=2.455 $Y=0.895 $X2=-0.19
+ $Y2=-0.245
cc_143 N_A1_c_166_p N_A_304_74#_M1004_d 0.00115008f $X=1.685 $Y=0.895 $X2=-0.19
+ $Y2=-0.245
cc_144 N_A1_c_130_n N_A_304_74#_c_312_n 0.00640423f $X=1.6 $Y=1.22 $X2=0 $Y2=0
cc_145 N_A1_c_131_n N_A_304_74#_c_312_n 9.64054e-19 $X=1.51 $Y=1.385 $X2=0 $Y2=0
cc_146 N_A1_c_132_n N_A_304_74#_c_312_n 0.0248292f $X=1.6 $Y=1.385 $X2=0 $Y2=0
cc_147 N_A1_c_134_n N_A_304_74#_c_312_n 9.75614e-19 $X=1.51 $Y=1.22 $X2=0 $Y2=0
cc_148 N_A1_c_129_n N_A_304_74#_c_319_n 0.00268326f $X=2.545 $Y=1.765 $X2=0
+ $Y2=0
cc_149 N_A1_c_131_n N_A_304_74#_c_319_n 0.00798977f $X=1.51 $Y=1.385 $X2=0 $Y2=0
cc_150 N_A1_c_132_n N_A_304_74#_c_319_n 0.0255946f $X=1.6 $Y=1.385 $X2=0 $Y2=0
cc_151 N_A1_c_129_n N_A_304_74#_c_339_n 0.00101813f $X=2.545 $Y=1.765 $X2=0
+ $Y2=0
cc_152 N_A1_c_141_p N_A_304_74#_c_339_n 0.0469474f $X=2.455 $Y=0.895 $X2=0 $Y2=0
cc_153 N_A1_c_166_p N_A_304_74#_c_339_n 0.00879433f $X=1.685 $Y=0.895 $X2=0
+ $Y2=0
cc_154 N_A1_c_131_n N_A_304_74#_c_339_n 4.1964e-19 $X=1.51 $Y=1.385 $X2=0 $Y2=0
cc_155 N_A1_c_132_n N_A_304_74#_c_339_n 0.00424542f $X=1.6 $Y=1.385 $X2=0 $Y2=0
cc_156 N_A1_c_134_n N_A_304_74#_c_339_n 0.0157207f $X=1.51 $Y=1.22 $X2=0 $Y2=0
cc_157 N_A1_c_157_p N_A_304_74#_c_339_n 0.0267499f $X=2.62 $Y=0.98 $X2=0 $Y2=0
cc_158 N_A1_c_129_n N_A_304_74#_c_346_n 0.0118341f $X=2.545 $Y=1.765 $X2=0 $Y2=0
cc_159 N_A1_c_157_p N_A_304_74#_c_347_n 0.0137943f $X=2.62 $Y=0.98 $X2=0 $Y2=0
cc_160 A1 N_A_304_74#_c_314_n 0.0145689f $X=2.555 $Y=0.84 $X2=0 $Y2=0
cc_161 N_A1_c_129_n N_VPWR_c_415_n 7.26245e-19 $X=2.545 $Y=1.765 $X2=0 $Y2=0
cc_162 N_A1_c_134_n N_VGND_c_481_n 9.47121e-19 $X=1.51 $Y=1.22 $X2=0 $Y2=0
cc_163 N_A1_c_134_n N_VGND_c_485_n 0.00296985f $X=1.51 $Y=1.22 $X2=0 $Y2=0
cc_164 N_A1_c_134_n N_VGND_c_489_n 0.00365796f $X=1.51 $Y=1.22 $X2=0 $Y2=0
cc_165 N_A1_c_141_p A_443_74# 0.00928686f $X=2.455 $Y=0.895 $X2=-0.19 $Y2=-0.245
cc_166 A1 A_443_74# 0.003907f $X=2.555 $Y=0.84 $X2=-0.19 $Y2=-0.245
cc_167 N_A1_c_157_p A_443_74# 0.00822687f $X=2.62 $Y=0.98 $X2=-0.19 $Y2=-0.245
cc_168 N_A0_c_191_n N_A_27_112#_c_239_n 0.00442776f $X=2.005 $Y=1.765 $X2=0
+ $Y2=0
cc_169 N_A0_c_191_n N_A_27_112#_c_229_n 0.0146215f $X=2.005 $Y=1.765 $X2=0 $Y2=0
cc_170 N_A0_c_191_n N_A_27_112#_c_230_n 0.012065f $X=2.005 $Y=1.765 $X2=0 $Y2=0
cc_171 N_A0_c_191_n N_A_304_74#_c_319_n 0.0209586f $X=2.005 $Y=1.765 $X2=0 $Y2=0
cc_172 A0 N_A_304_74#_c_319_n 0.0310181f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_173 N_A0_c_192_n N_A_304_74#_c_339_n 0.017902f $X=2.14 $Y=1.22 $X2=0 $Y2=0
cc_174 N_A0_c_191_n N_A_304_74#_c_346_n 0.0386202f $X=2.005 $Y=1.765 $X2=0 $Y2=0
cc_175 N_A0_c_191_n N_VPWR_c_415_n 7.26245e-19 $X=2.005 $Y=1.765 $X2=0 $Y2=0
cc_176 N_A0_c_192_n N_VGND_c_485_n 0.00296985f $X=2.14 $Y=1.22 $X2=0 $Y2=0
cc_177 N_A0_c_192_n N_VGND_c_489_n 0.00371085f $X=2.14 $Y=1.22 $X2=0 $Y2=0
cc_178 N_A_27_112#_M1008_g N_A_304_74#_c_310_n 5.37584e-19 $X=3.1 $Y=0.74 $X2=0
+ $Y2=0
cc_179 N_A_27_112#_c_221_n N_A_304_74#_c_310_n 0.0440864f $X=3.115 $Y=1.765
+ $X2=0 $Y2=0
cc_180 N_A_27_112#_c_224_n N_A_304_74#_c_310_n 0.00106764f $X=3.04 $Y=2.905
+ $X2=0 $Y2=0
cc_181 N_A_27_112#_c_226_n N_A_304_74#_c_310_n 4.74404e-19 $X=3.19 $Y=1.485
+ $X2=0 $Y2=0
cc_182 N_A_27_112#_M1008_g N_A_304_74#_M1009_g 0.0140133f $X=3.1 $Y=0.74 $X2=0
+ $Y2=0
cc_183 N_A_27_112#_c_239_n N_A_304_74#_c_319_n 0.0117605f $X=1.15 $Y=2.145 $X2=0
+ $Y2=0
cc_184 N_A_27_112#_c_224_n N_A_304_74#_c_319_n 0.00604f $X=3.04 $Y=2.905 $X2=0
+ $Y2=0
cc_185 N_A_27_112#_c_239_n N_A_304_74#_c_324_n 0.00864977f $X=1.15 $Y=2.145
+ $X2=0 $Y2=0
cc_186 N_A_27_112#_M1008_g N_A_304_74#_c_339_n 0.0110865f $X=3.1 $Y=0.74 $X2=0
+ $Y2=0
cc_187 N_A_27_112#_c_230_n N_A_304_74#_c_346_n 0.0230185f $X=2.955 $Y=2.99 $X2=0
+ $Y2=0
cc_188 N_A_27_112#_c_224_n N_A_304_74#_c_346_n 0.026447f $X=3.04 $Y=2.905 $X2=0
+ $Y2=0
cc_189 N_A_27_112#_M1008_g N_A_304_74#_c_347_n 0.0123701f $X=3.1 $Y=0.74 $X2=0
+ $Y2=0
cc_190 N_A_27_112#_M1008_g N_A_304_74#_c_313_n 0.00664159f $X=3.1 $Y=0.74 $X2=0
+ $Y2=0
cc_191 N_A_27_112#_c_221_n N_A_304_74#_c_313_n 0.00411621f $X=3.115 $Y=1.765
+ $X2=0 $Y2=0
cc_192 N_A_27_112#_c_226_n N_A_304_74#_c_313_n 0.0170649f $X=3.19 $Y=1.485 $X2=0
+ $Y2=0
cc_193 N_A_27_112#_M1008_g N_A_304_74#_c_314_n 0.00567512f $X=3.1 $Y=0.74 $X2=0
+ $Y2=0
cc_194 N_A_27_112#_c_226_n N_A_304_74#_c_314_n 0.0141748f $X=3.19 $Y=1.485 $X2=0
+ $Y2=0
cc_195 N_A_27_112#_M1008_g N_A_304_74#_c_315_n 0.00279208f $X=3.1 $Y=0.74 $X2=0
+ $Y2=0
cc_196 N_A_27_112#_M1008_g N_A_304_74#_c_316_n 3.83846e-19 $X=3.1 $Y=0.74 $X2=0
+ $Y2=0
cc_197 N_A_27_112#_c_221_n N_A_304_74#_c_316_n 0.0010311f $X=3.115 $Y=1.765
+ $X2=0 $Y2=0
cc_198 N_A_27_112#_c_226_n N_A_304_74#_c_316_n 0.0251871f $X=3.19 $Y=1.485 $X2=0
+ $Y2=0
cc_199 N_A_27_112#_c_239_n N_VPWR_M1005_d 0.00671692f $X=1.15 $Y=2.145 $X2=-0.19
+ $Y2=-0.245
cc_200 N_A_27_112#_c_239_n N_VPWR_c_413_n 0.0219335f $X=1.15 $Y=2.145 $X2=0
+ $Y2=0
cc_201 N_A_27_112#_c_229_n N_VPWR_c_413_n 0.0213191f $X=1.235 $Y=2.905 $X2=0
+ $Y2=0
cc_202 N_A_27_112#_c_231_n N_VPWR_c_413_n 0.0147692f $X=1.32 $Y=2.99 $X2=0 $Y2=0
cc_203 N_A_27_112#_c_233_n N_VPWR_c_413_n 0.0201945f $X=0.28 $Y=2.06 $X2=0 $Y2=0
cc_204 N_A_27_112#_c_221_n N_VPWR_c_414_n 0.0115271f $X=3.115 $Y=1.765 $X2=0
+ $Y2=0
cc_205 N_A_27_112#_c_230_n N_VPWR_c_414_n 0.0147425f $X=2.955 $Y=2.99 $X2=0
+ $Y2=0
cc_206 N_A_27_112#_c_224_n N_VPWR_c_414_n 0.0803764f $X=3.04 $Y=2.905 $X2=0
+ $Y2=0
cc_207 N_A_27_112#_c_226_n N_VPWR_c_414_n 0.00497567f $X=3.19 $Y=1.485 $X2=0
+ $Y2=0
cc_208 N_A_27_112#_c_221_n N_VPWR_c_415_n 0.00255182f $X=3.115 $Y=1.765 $X2=0
+ $Y2=0
cc_209 N_A_27_112#_c_230_n N_VPWR_c_415_n 0.117416f $X=2.955 $Y=2.99 $X2=0 $Y2=0
cc_210 N_A_27_112#_c_231_n N_VPWR_c_415_n 0.0121867f $X=1.32 $Y=2.99 $X2=0 $Y2=0
cc_211 N_A_27_112#_c_221_n N_VPWR_c_412_n 0.00220298f $X=3.115 $Y=1.765 $X2=0
+ $Y2=0
cc_212 N_A_27_112#_c_230_n N_VPWR_c_412_n 0.0680683f $X=2.955 $Y=2.99 $X2=0
+ $Y2=0
cc_213 N_A_27_112#_c_231_n N_VPWR_c_412_n 0.00660921f $X=1.32 $Y=2.99 $X2=0
+ $Y2=0
cc_214 N_A_27_112#_c_233_n N_VPWR_c_412_n 0.00997343f $X=0.28 $Y=2.06 $X2=0
+ $Y2=0
cc_215 N_A_27_112#_c_233_n N_VPWR_c_419_n 0.0066794f $X=0.28 $Y=2.06 $X2=0 $Y2=0
cc_216 N_A_27_112#_c_239_n A_223_368# 0.00523811f $X=1.15 $Y=2.145 $X2=-0.19
+ $Y2=-0.245
cc_217 N_A_27_112#_c_229_n A_223_368# 0.0140365f $X=1.235 $Y=2.905 $X2=-0.19
+ $Y2=-0.245
cc_218 N_A_27_112#_c_224_n A_524_368# 0.0147002f $X=3.04 $Y=2.905 $X2=-0.19
+ $Y2=-0.245
cc_219 N_A_27_112#_M1008_g N_X_c_457_n 8.05779e-19 $X=3.1 $Y=0.74 $X2=0 $Y2=0
cc_220 N_A_27_112#_c_225_n N_VGND_c_482_n 0.0112976f $X=0.28 $Y=1.13 $X2=0 $Y2=0
cc_221 N_A_27_112#_M1008_g N_VGND_c_483_n 0.00814582f $X=3.1 $Y=0.74 $X2=0 $Y2=0
cc_222 N_A_27_112#_c_222_n N_VGND_c_484_n 0.0112976f $X=0.28 $Y=0.835 $X2=0
+ $Y2=0
cc_223 N_A_27_112#_M1008_g N_VGND_c_485_n 0.00351724f $X=3.1 $Y=0.74 $X2=0 $Y2=0
cc_224 N_A_27_112#_c_222_n N_VGND_c_487_n 0.0081085f $X=0.28 $Y=0.835 $X2=0
+ $Y2=0
cc_225 N_A_27_112#_M1008_g N_VGND_c_489_n 0.0055287f $X=3.1 $Y=0.74 $X2=0 $Y2=0
cc_226 N_A_27_112#_c_222_n N_VGND_c_489_n 0.010608f $X=0.28 $Y=0.835 $X2=0 $Y2=0
cc_227 N_A_304_74#_c_310_n N_VPWR_c_414_n 0.0141871f $X=3.735 $Y=1.765 $X2=0
+ $Y2=0
cc_228 N_A_304_74#_c_313_n N_VPWR_c_414_n 0.00547729f $X=3.525 $Y=1.065 $X2=0
+ $Y2=0
cc_229 N_A_304_74#_c_316_n N_VPWR_c_414_n 0.00784726f $X=3.73 $Y=1.465 $X2=0
+ $Y2=0
cc_230 N_A_304_74#_c_310_n N_VPWR_c_417_n 0.00445602f $X=3.735 $Y=1.765 $X2=0
+ $Y2=0
cc_231 N_A_304_74#_c_310_n N_VPWR_c_412_n 0.0086545f $X=3.735 $Y=1.765 $X2=0
+ $Y2=0
cc_232 N_A_304_74#_c_319_n A_223_368# 0.0237834f $X=2.065 $Y=1.805 $X2=-0.19
+ $Y2=-0.245
cc_233 N_A_304_74#_M1009_g N_X_c_457_n 0.0105488f $X=3.815 $Y=0.74 $X2=0 $Y2=0
cc_234 N_A_304_74#_M1009_g N_X_c_458_n 0.00309954f $X=3.815 $Y=0.74 $X2=0 $Y2=0
cc_235 N_A_304_74#_c_313_n N_X_c_458_n 0.00664075f $X=3.525 $Y=1.065 $X2=0 $Y2=0
cc_236 N_A_304_74#_c_316_n N_X_c_458_n 0.00233746f $X=3.73 $Y=1.465 $X2=0 $Y2=0
cc_237 N_A_304_74#_c_310_n X 0.0107426f $X=3.735 $Y=1.765 $X2=0 $Y2=0
cc_238 N_A_304_74#_c_310_n N_X_c_461_n 0.00510184f $X=3.735 $Y=1.765 $X2=0 $Y2=0
cc_239 N_A_304_74#_c_316_n N_X_c_461_n 0.00761489f $X=3.73 $Y=1.465 $X2=0 $Y2=0
cc_240 N_A_304_74#_c_310_n N_X_c_459_n 0.00683011f $X=3.735 $Y=1.765 $X2=0 $Y2=0
cc_241 N_A_304_74#_M1009_g N_X_c_459_n 0.00252268f $X=3.815 $Y=0.74 $X2=0 $Y2=0
cc_242 N_A_304_74#_c_315_n N_X_c_459_n 0.005258f $X=3.61 $Y=1.3 $X2=0 $Y2=0
cc_243 N_A_304_74#_c_316_n N_X_c_459_n 0.0249903f $X=3.73 $Y=1.465 $X2=0 $Y2=0
cc_244 N_A_304_74#_c_313_n N_VGND_M1008_d 0.0107009f $X=3.525 $Y=1.065 $X2=0
+ $Y2=0
cc_245 N_A_304_74#_c_312_n N_VGND_c_482_n 0.00787863f $X=1.09 $Y=1.72 $X2=0
+ $Y2=0
cc_246 N_A_304_74#_c_328_n N_VGND_c_482_n 0.0126934f $X=1.26 $Y=0.935 $X2=0
+ $Y2=0
cc_247 N_A_304_74#_c_310_n N_VGND_c_483_n 2.35935e-19 $X=3.735 $Y=1.765 $X2=0
+ $Y2=0
cc_248 N_A_304_74#_M1009_g N_VGND_c_483_n 0.00795549f $X=3.815 $Y=0.74 $X2=0
+ $Y2=0
cc_249 N_A_304_74#_c_339_n N_VGND_c_483_n 0.0206009f $X=2.955 $Y=0.515 $X2=0
+ $Y2=0
cc_250 N_A_304_74#_c_347_n N_VGND_c_483_n 0.0125449f $X=3.04 $Y=0.98 $X2=0 $Y2=0
cc_251 N_A_304_74#_c_313_n N_VGND_c_483_n 0.0270533f $X=3.525 $Y=1.065 $X2=0
+ $Y2=0
cc_252 N_A_304_74#_c_339_n N_VGND_c_485_n 0.0577426f $X=2.955 $Y=0.515 $X2=0
+ $Y2=0
cc_253 N_A_304_74#_c_400_p N_VGND_c_485_n 0.0054507f $X=1.345 $Y=0.515 $X2=0
+ $Y2=0
cc_254 N_A_304_74#_M1009_g N_VGND_c_488_n 0.00434272f $X=3.815 $Y=0.74 $X2=0
+ $Y2=0
cc_255 N_A_304_74#_M1009_g N_VGND_c_489_n 0.00827137f $X=3.815 $Y=0.74 $X2=0
+ $Y2=0
cc_256 N_A_304_74#_c_339_n N_VGND_c_489_n 0.0601803f $X=2.955 $Y=0.515 $X2=0
+ $Y2=0
cc_257 N_A_304_74#_c_400_p N_VGND_c_489_n 0.00604114f $X=1.345 $Y=0.515 $X2=0
+ $Y2=0
cc_258 N_A_304_74#_c_328_n N_VGND_c_489_n 0.00496217f $X=1.26 $Y=0.935 $X2=0
+ $Y2=0
cc_259 N_A_304_74#_c_406_p A_226_74# 3.7257e-19 $X=1.26 $Y=0.85 $X2=-0.19
+ $Y2=-0.245
cc_260 N_A_304_74#_c_400_p A_226_74# 0.00162909f $X=1.345 $Y=0.515 $X2=-0.19
+ $Y2=-0.245
cc_261 N_A_304_74#_c_328_n A_226_74# 0.00520569f $X=1.26 $Y=0.935 $X2=-0.19
+ $Y2=-0.245
cc_262 N_A_304_74#_c_339_n A_443_74# 0.0266902f $X=2.955 $Y=0.515 $X2=-0.19
+ $Y2=-0.245
cc_263 N_A_304_74#_c_347_n A_443_74# 0.00824479f $X=3.04 $Y=0.98 $X2=-0.19
+ $Y2=-0.245
cc_264 N_A_304_74#_c_314_n A_443_74# 0.00144215f $X=3.125 $Y=1.065 $X2=-0.19
+ $Y2=-0.245
cc_265 N_VPWR_c_417_n X 0.0195021f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_266 N_VPWR_c_412_n X 0.0161093f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_267 N_VPWR_c_414_n N_X_c_461_n 0.0470261f $X=3.46 $Y=1.985 $X2=0 $Y2=0
cc_268 N_X_c_457_n N_VGND_c_483_n 0.0276686f $X=4.03 $Y=0.515 $X2=0 $Y2=0
cc_269 N_X_c_457_n N_VGND_c_488_n 0.0163488f $X=4.03 $Y=0.515 $X2=0 $Y2=0
cc_270 N_X_c_457_n N_VGND_c_489_n 0.0134757f $X=4.03 $Y=0.515 $X2=0 $Y2=0
