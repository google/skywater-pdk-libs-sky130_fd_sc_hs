* File: sky130_fd_sc_hs__a31o_4.spice
* Created: Tue Sep  1 19:53:01 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hs__a31o_4.pex.spice"
.subckt sky130_fd_sc_hs__a31o_4  VNB VPB B1 A1 A2 A3 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A3	A3
* A2	A2
* A1	A1
* B1	B1
* VPB	VPB
* VNB	VNB
MM1008 N_X_M1008_d N_A_83_274#_M1008_g N_VGND_M1008_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.12025 AS=0.2294 PD=1.065 PS=2.1 NRD=7.296 NRS=4.044 M=1 R=4.93333
+ SA=75000.2 SB=75001.6 A=0.111 P=1.78 MULT=1
MM1009 N_X_M1008_d N_A_83_274#_M1009_g N_VGND_M1009_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.12025 AS=0.1036 PD=1.065 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.7
+ SB=75001.1 A=0.111 P=1.78 MULT=1
MM1019 N_X_M1019_d N_A_83_274#_M1019_g N_VGND_M1009_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.11285 AS=0.1036 PD=1.045 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.1
+ SB=75000.7 A=0.111 P=1.78 MULT=1
MM1022 N_X_M1019_d N_A_83_274#_M1022_g N_VGND_M1022_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.11285 AS=0.2109 PD=1.045 PS=2.05 NRD=4.044 NRS=0 M=1 R=4.93333 SA=75001.6
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1002 N_A_83_274#_M1002_d N_B1_M1002_g N_VGND_M1002_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.1824 AS=0.112 PD=1.85 PS=0.99 NRD=0 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75001.7 A=0.096 P=1.58 MULT=1
MM1007 N_A_83_274#_M1007_d N_B1_M1007_g N_VGND_M1002_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.0896 AS=0.112 PD=0.92 PS=0.99 NRD=0 NRS=13.116 M=1 R=4.26667 SA=75000.7
+ SB=75001.2 A=0.096 P=1.58 MULT=1
MM1011 N_A_83_274#_M1007_d N_A1_M1011_g N_A_775_74#_M1011_s VNB NLOWVT L=0.15
+ W=0.64 AD=0.0896 AS=0.112 PD=0.92 PS=0.99 NRD=0 NRS=13.116 M=1 R=4.26667
+ SA=75001.1 SB=75000.8 A=0.096 P=1.58 MULT=1
MM1013 N_A_83_274#_M1013_d N_A1_M1013_g N_A_775_74#_M1011_s VNB NLOWVT L=0.15
+ W=0.64 AD=0.2272 AS=0.112 PD=1.99 PS=0.99 NRD=13.116 NRS=0 M=1 R=4.26667
+ SA=75001.6 SB=75000.3 A=0.096 P=1.58 MULT=1
MM1006 N_A_775_74#_M1006_d N_A2_M1006_g N_A_1000_74#_M1006_s VNB NLOWVT L=0.15
+ W=0.64 AD=0.0896 AS=0.1824 PD=0.92 PS=1.85 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75001.5 A=0.096 P=1.58 MULT=1
MM1018 N_A_775_74#_M1006_d N_A2_M1018_g N_A_1000_74#_M1018_s VNB NLOWVT L=0.15
+ W=0.64 AD=0.0896 AS=0.0896 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.6 SB=75001.1 A=0.096 P=1.58 MULT=1
MM1003 N_VGND_M1003_d N_A3_M1003_g N_A_1000_74#_M1018_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.0896 AS=0.0896 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667 SA=75001.1
+ SB=75000.6 A=0.096 P=1.58 MULT=1
MM1014 N_VGND_M1003_d N_A3_M1014_g N_A_1000_74#_M1014_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.0896 AS=0.1824 PD=0.92 PS=1.85 NRD=0 NRS=0 M=1 R=4.26667 SA=75001.5
+ SB=75000.2 A=0.096 P=1.58 MULT=1
MM1010 N_X_M1010_d N_A_83_274#_M1010_g N_VPWR_M1010_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.3304 PD=1.42 PS=2.83 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75001.7 A=0.168 P=2.54 MULT=1
MM1012 N_X_M1010_d N_A_83_274#_M1012_g N_VPWR_M1012_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.224 PD=1.42 PS=1.52 NRD=1.7533 NRS=10.5395 M=1 R=7.46667
+ SA=75000.7 SB=75001.3 A=0.168 P=2.54 MULT=1
MM1015 N_X_M1015_d N_A_83_274#_M1015_g N_VPWR_M1012_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.224 PD=1.42 PS=1.52 NRD=1.7533 NRS=10.5395 M=1 R=7.46667
+ SA=75001.2 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1017 N_X_M1015_d N_A_83_274#_M1017_g N_VPWR_M1017_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.3864 PD=1.42 PS=2.93 NRD=1.7533 NRS=10.5395 M=1 R=7.46667
+ SA=75001.7 SB=75000.3 A=0.168 P=2.54 MULT=1
MM1000 N_A_529_392#_M1000_d N_B1_M1000_g N_A_83_274#_M1000_s VPB PSHORT L=0.15
+ W=1 AD=0.295 AS=0.185 PD=2.59 PS=1.37 NRD=1.9503 NRS=13.7703 M=1 R=6.66667
+ SA=75000.2 SB=75003.9 A=0.15 P=2.3 MULT=1
MM1020 N_A_529_392#_M1020_d N_B1_M1020_g N_A_83_274#_M1000_s VPB PSHORT L=0.15
+ W=1 AD=0.225 AS=0.185 PD=1.45 PS=1.37 NRD=31.5003 NRS=3.9203 M=1 R=6.66667
+ SA=75000.7 SB=75003.4 A=0.15 P=2.3 MULT=1
MM1016 N_A_529_392#_M1020_d N_A1_M1016_g N_VPWR_M1016_s VPB PSHORT L=0.15 W=1
+ AD=0.225 AS=0.2 PD=1.45 PS=1.4 NRD=1.9503 NRS=11.8003 M=1 R=6.66667 SA=75001.3
+ SB=75002.8 A=0.15 P=2.3 MULT=1
MM1021 N_A_529_392#_M1021_d N_A1_M1021_g N_VPWR_M1016_s VPB PSHORT L=0.15 W=1
+ AD=0.15 AS=0.2 PD=1.3 PS=1.4 NRD=1.9503 NRS=11.8003 M=1 R=6.66667 SA=75001.9
+ SB=75002.2 A=0.15 P=2.3 MULT=1
MM1004 N_A_529_392#_M1021_d N_A2_M1004_g N_VPWR_M1004_s VPB PSHORT L=0.15 W=1
+ AD=0.15 AS=0.205 PD=1.3 PS=1.41 NRD=1.9503 NRS=11.8003 M=1 R=6.66667
+ SA=75002.3 SB=75001.8 A=0.15 P=2.3 MULT=1
MM1023 N_A_529_392#_M1023_d N_A2_M1023_g N_VPWR_M1004_s VPB PSHORT L=0.15 W=1
+ AD=0.175 AS=0.205 PD=1.35 PS=1.41 NRD=1.9503 NRS=13.7703 M=1 R=6.66667
+ SA=75002.9 SB=75001.2 A=0.15 P=2.3 MULT=1
MM1001 N_A_529_392#_M1023_d N_A3_M1001_g N_VPWR_M1001_s VPB PSHORT L=0.15 W=1
+ AD=0.175 AS=0.175 PD=1.35 PS=1.35 NRD=11.8003 NRS=1.9503 M=1 R=6.66667
+ SA=75003.4 SB=75000.7 A=0.15 P=2.3 MULT=1
MM1005 N_A_529_392#_M1005_d N_A3_M1005_g N_VPWR_M1001_s VPB PSHORT L=0.15 W=1
+ AD=0.295 AS=0.175 PD=2.59 PS=1.35 NRD=1.9503 NRS=11.8003 M=1 R=6.66667
+ SA=75003.9 SB=75000.2 A=0.15 P=2.3 MULT=1
DX24_noxref VNB VPB NWDIODE A=14.0988 P=18.88
*
.include "sky130_fd_sc_hs__a31o_4.pxi.spice"
*
.ends
*
*
