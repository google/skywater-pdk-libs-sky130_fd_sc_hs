* File: sky130_fd_sc_hs__clkdlyinv3sd1_1.spice
* Created: Tue Sep  1 19:57:59 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hs__clkdlyinv3sd1_1.pex.spice"
.subckt sky130_fd_sc_hs__clkdlyinv3sd1_1  VNB VPB A VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A	A
* VPB	VPB
* VNB	VNB
MM1003 N_VGND_M1003_d N_A_M1003_g N_A_28_74#_M1003_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.15435 AS=0.1113 PD=1.155 PS=1.37 NRD=15.708 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1004 N_A_285_392#_M1004_d N_A_28_74#_M1004_g N_VGND_M1003_d VNB NLOWVT L=0.15
+ W=0.42 AD=0.1113 AS=0.15435 PD=1.37 PS=1.155 NRD=0 NRS=114.276 M=1 R=2.8
+ SA=75001.1 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1005 N_Y_M1005_d N_A_285_392#_M1005_g N_VGND_M1005_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.1113 AS=0.1113 PD=1.37 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1000 N_VPWR_M1000_d N_A_M1000_g N_A_28_74#_M1000_s VPB PSHORT L=0.15 W=1.12
+ AD=0.389253 AS=0.3136 PD=1.9283 PS=2.8 NRD=5.2599 NRS=2.6201 M=1 R=7.46667
+ SA=75000.2 SB=75001 A=0.168 P=2.54 MULT=1
MM1002 N_A_285_392#_M1002_d N_A_28_74#_M1002_g N_VPWR_M1000_d VPB PSHORT L=0.15
+ W=1 AD=0.28 AS=0.347547 PD=2.56 PS=1.7217 NRD=2.9353 NRS=77.7953 M=1 R=6.66667
+ SA=75001.1 SB=75000.2 A=0.15 P=2.3 MULT=1
MM1001 N_Y_M1001_d N_A_285_392#_M1001_g N_VPWR_M1001_s VPB PSHORT L=0.15 W=1.12
+ AD=0.3136 AS=0.308 PD=2.8 PS=2.79 NRD=2.6201 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75000.2 A=0.168 P=2.54 MULT=1
DX6_noxref VNB VPB NWDIODE A=6.0636 P=10.24
*
.include "sky130_fd_sc_hs__clkdlyinv3sd1_1.pxi.spice"
*
.ends
*
*
