* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hs__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
X0 a_195_74# A2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X1 X a_27_368# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X2 VGND a_27_368# X VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X3 a_27_368# C1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=150000u
X4 X a_27_368# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X5 a_117_74# B1 a_195_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X6 a_27_368# C1 a_117_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X7 VGND A1 a_195_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X8 a_314_368# A1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=150000u
X9 VPWR B1 a_27_368# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=150000u
X10 VPWR a_27_368# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X11 a_27_368# A2 a_314_368# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=150000u
.ends
