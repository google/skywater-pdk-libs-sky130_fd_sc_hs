* File: sky130_fd_sc_hs__sdfbbn_2.spice
* Created: Tue Sep  1 20:22:06 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hs__sdfbbn_2.pex.spice"
.subckt sky130_fd_sc_hs__sdfbbn_2  VNB VPB SCD D SCE CLK_N SET_B RESET_B VPWR
+ Q_N Q VGND
* 
* VGND	VGND
* Q	Q
* Q_N	Q_N
* VPWR	VPWR
* RESET_B	RESET_B
* SET_B	SET_B
* CLK_N	CLK_N
* SCE	SCE
* D	D
* SCD	SCD
* VPB	VPB
* VNB	VNB
MM1004 A_119_119# N_SCD_M1004_g N_VGND_M1004_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.0504 AS=0.1197 PD=0.66 PS=1.41 NRD=18.564 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75002.5 A=0.063 P=1.14 MULT=1
MM1035 N_A_197_119#_M1035_d N_SCE_M1035_g A_119_119# VNB NLOWVT L=0.15 W=0.42
+ AD=0.1428 AS=0.0504 PD=1.1 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75000.6
+ SB=75002.1 A=0.063 P=1.14 MULT=1
MM1045 A_363_119# N_D_M1045_g N_A_197_119#_M1035_d VNB NLOWVT L=0.15 W=0.42
+ AD=0.0504 AS=0.1428 PD=0.66 PS=1.1 NRD=18.564 NRS=0 M=1 R=2.8 SA=75001.4
+ SB=75001.3 A=0.063 P=1.14 MULT=1
MM1028 N_VGND_M1028_d N_A_341_410#_M1028_g A_363_119# VNB NLOWVT L=0.15 W=0.42
+ AD=0.1113 AS=0.0504 PD=0.95 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75001.8
+ SB=75000.9 A=0.063 P=1.14 MULT=1
MM1040 N_A_341_410#_M1040_d N_SCE_M1040_g N_VGND_M1028_d VNB NLOWVT L=0.15
+ W=0.42 AD=0.1197 AS=0.1113 PD=1.41 PS=0.95 NRD=0 NRS=71.424 M=1 R=2.8
+ SA=75002.5 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1037 N_VGND_M1037_d N_CLK_N_M1037_g N_A_688_98#_M1037_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.30025 AS=0.2109 PD=1.74 PS=2.05 NRD=56.868 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75001.1 A=0.111 P=1.78 MULT=1
MM1047 N_A_868_368#_M1047_d N_A_688_98#_M1047_g N_VGND_M1037_d VNB NLOWVT L=0.15
+ W=0.74 AD=0.2109 AS=0.30025 PD=2.05 PS=1.74 NRD=0 NRS=56.868 M=1 R=4.93333
+ SA=75001.1 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1030 A_1185_125# N_A_1007_366#_M1030_g N_VGND_M1030_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.0441 AS=0.24385 PD=0.63 PS=2.14 NRD=14.28 NRS=150.168 M=1 R=2.8
+ SA=75000.3 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1016 N_A_1154_464#_M1016_d N_A_688_98#_M1016_g A_1185_125# VNB NLOWVT L=0.15
+ W=0.42 AD=0.06405 AS=0.0441 PD=0.725 PS=0.63 NRD=7.14 NRS=14.28 M=1 R=2.8
+ SA=75000.7 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1005 N_A_197_119#_M1005_d N_A_868_368#_M1005_g N_A_1154_464#_M1016_d VNB
+ NLOWVT L=0.15 W=0.42 AD=0.1491 AS=0.06405 PD=1.55 PS=0.725 NRD=19.992 NRS=0
+ M=1 R=2.8 SA=75001.1 SB=75000.3 A=0.063 P=1.14 MULT=1
MM1018 N_A_1007_366#_M1018_d N_A_1154_464#_M1018_g N_A_1473_73#_M1018_s VNB
+ NLOWVT L=0.15 W=0.55 AD=0.077 AS=0.3531 PD=0.83 PS=2.54 NRD=0 NRS=128.064 M=1
+ R=3.66667 SA=75000.4 SB=75003.2 A=0.0825 P=1.4 MULT=1
MM1021 N_A_1473_73#_M1021_d N_A_1643_257#_M1021_g N_A_1007_366#_M1018_d VNB
+ NLOWVT L=0.15 W=0.55 AD=0.125125 AS=0.077 PD=1.005 PS=0.83 NRD=26.172 NRS=0
+ M=1 R=3.66667 SA=75000.8 SB=75002.8 A=0.0825 P=1.4 MULT=1
MM1051 N_VGND_M1051_d N_SET_B_M1051_g N_A_1473_73#_M1021_d VNB NLOWVT L=0.15
+ W=0.55 AD=0.09625 AS=0.125125 PD=0.9 PS=1.005 NRD=15.264 NRS=11.988 M=1
+ R=3.66667 SA=75001.4 SB=75002.2 A=0.0825 P=1.4 MULT=1
MM1049 A_1902_125# N_A_1007_366#_M1049_g N_VGND_M1051_d VNB NLOWVT L=0.15 W=0.55
+ AD=0.108187 AS=0.09625 PD=1.09 PS=0.9 NRD=30.912 NRS=0 M=1 R=3.66667
+ SA=75001.9 SB=75001.7 A=0.0825 P=1.4 MULT=1
MM1023 N_A_1997_82#_M1023_d N_A_688_98#_M1023_g A_1902_125# VNB NLOWVT L=0.15
+ W=0.55 AD=0.280387 AS=0.108187 PD=1.87113 PS=1.09 NRD=0 NRS=30.912 M=1
+ R=3.66667 SA=75001.5 SB=75002.7 A=0.0825 P=1.4 MULT=1
MM1014 A_2247_82# N_A_868_368#_M1014_g N_A_1997_82#_M1023_d VNB NLOWVT L=0.15
+ W=0.42 AD=0.0504 AS=0.214113 PD=0.66 PS=1.42887 NRD=18.564 NRS=0 M=1 R=2.8
+ SA=75002.5 SB=75002.3 A=0.063 P=1.14 MULT=1
MM1048 N_VGND_M1048_d N_A_2216_410#_M1048_g A_2247_82# VNB NLOWVT L=0.15 W=0.42
+ AD=0.125656 AS=0.0504 PD=1.01017 PS=0.66 NRD=30 NRS=18.564 M=1 R=2.8
+ SA=75002.9 SB=75001.9 A=0.063 P=1.14 MULT=1
MM1002 N_A_2452_74#_M1002_d N_SET_B_M1002_g N_VGND_M1048_d VNB NLOWVT L=0.15
+ W=0.74 AD=0.1369 AS=0.221394 PD=1.11 PS=1.77983 NRD=0 NRS=39.588 M=1 R=4.93333
+ SA=75002.1 SB=75001.2 A=0.111 P=1.78 MULT=1
MM1041 N_A_2216_410#_M1041_d N_A_1643_257#_M1041_g N_A_2452_74#_M1002_d VNB
+ NLOWVT L=0.15 W=0.74 AD=0.1036 AS=0.1369 PD=1.02 PS=1.11 NRD=0 NRS=7.296 M=1
+ R=4.93333 SA=75002.6 SB=75000.7 A=0.111 P=1.78 MULT=1
MM1009 N_A_2452_74#_M1009_d N_A_1997_82#_M1009_g N_A_2216_410#_M1041_d VNB
+ NLOWVT L=0.15 W=0.74 AD=0.30055 AS=0.1036 PD=2.42 PS=1.02 NRD=13.776 NRS=0 M=1
+ R=4.93333 SA=75003 SB=75000.3 A=0.111 P=1.78 MULT=1
MM1007 N_VGND_M1007_d N_RESET_B_M1007_g N_A_1643_257#_M1007_s VNB NLOWVT L=0.15
+ W=0.42 AD=0.136772 AS=0.1176 PD=1.32517 PS=1.4 NRD=172.848 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75000.9 A=0.063 P=1.14 MULT=1
MM1003 N_VGND_M1007_d N_A_2216_410#_M1003_g N_Q_N_M1003_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.240978 AS=0.1036 PD=2.33483 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.5 SB=75000.7 A=0.111 P=1.78 MULT=1
MM1026 N_VGND_M1026_d N_A_2216_410#_M1026_g N_Q_N_M1003_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.2294 AS=0.1036 PD=2.1 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.9
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1022 N_VGND_M1022_d N_A_2216_410#_M1022_g N_A_3272_94#_M1022_s VNB NLOWVT
+ L=0.15 W=0.64 AD=0.150029 AS=0.1824 PD=1.10377 PS=1.85 NRD=19.212 NRS=0 M=1
+ R=4.26667 SA=75000.2 SB=75001.2 A=0.096 P=1.58 MULT=1
MM1027 N_Q_M1027_d N_A_3272_94#_M1027_g N_VGND_M1022_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.173471 PD=1.02 PS=1.27623 NRD=0 NRS=11.34 M=1 R=4.93333
+ SA=75000.7 SB=75000.6 A=0.111 P=1.78 MULT=1
MM1043 N_Q_M1027_d N_A_3272_94#_M1043_g N_VGND_M1043_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.2072 PD=1.02 PS=2.04 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.2
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1024 N_VPWR_M1024_d N_SCD_M1024_g N_A_27_464#_M1024_s VPB PSHORT L=0.15 W=0.64
+ AD=0.096 AS=0.1888 PD=0.94 PS=1.87 NRD=3.0732 NRS=3.0732 M=1 R=4.26667
+ SA=75000.2 SB=75001.5 A=0.096 P=1.58 MULT=1
MM1025 A_206_464# N_SCE_M1025_g N_VPWR_M1024_d VPB PSHORT L=0.15 W=0.64
+ AD=0.0768 AS=0.096 PD=0.88 PS=0.94 NRD=19.9955 NRS=3.0732 M=1 R=4.26667
+ SA=75000.7 SB=75001.1 A=0.096 P=1.58 MULT=1
MM1001 N_A_197_119#_M1001_d N_D_M1001_g A_206_464# VPB PSHORT L=0.15 W=0.64
+ AD=0.096 AS=0.0768 PD=0.94 PS=0.88 NRD=3.0732 NRS=19.9955 M=1 R=4.26667
+ SA=75001.1 SB=75000.7 A=0.096 P=1.58 MULT=1
MM1008 N_A_27_464#_M1008_d N_A_341_410#_M1008_g N_A_197_119#_M1001_d VPB PSHORT
+ L=0.15 W=0.64 AD=0.1888 AS=0.096 PD=1.87 PS=0.94 NRD=3.0732 NRS=3.0732 M=1
+ R=4.26667 SA=75001.5 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1032 N_A_341_410#_M1032_d N_SCE_M1032_g N_VPWR_M1032_s VPB PSHORT L=0.15
+ W=0.64 AD=0.1888 AS=0.1888 PD=1.87 PS=1.87 NRD=3.0732 NRS=3.0732 M=1 R=4.26667
+ SA=75000.2 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1012 N_VPWR_M1012_d N_CLK_N_M1012_g N_A_688_98#_M1012_s VPB PSHORT L=0.15
+ W=1.12 AD=0.168 AS=0.3304 PD=1.42 PS=2.83 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1015 N_A_868_368#_M1015_d N_A_688_98#_M1015_g N_VPWR_M1012_d VPB PSHORT L=0.15
+ W=1.12 AD=0.3304 AS=0.168 PD=2.83 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.7 SB=75000.2 A=0.168 P=2.54 MULT=1
MM1010 A_1070_464# N_A_1007_366#_M1010_g N_VPWR_M1010_s VPB PSHORT L=0.15 W=0.42
+ AD=0.0567 AS=0.1239 PD=0.69 PS=1.43 NRD=37.5088 NRS=4.6886 M=1 R=2.8
+ SA=75000.2 SB=75001.2 A=0.063 P=1.14 MULT=1
MM1017 N_A_1154_464#_M1017_d N_A_868_368#_M1017_g A_1070_464# VPB PSHORT L=0.15
+ W=0.42 AD=0.0897849 AS=0.0567 PD=0.812264 PS=0.69 NRD=44.5417 NRS=37.5088 M=1
+ R=2.8 SA=75000.6 SB=75000.8 A=0.063 P=1.14 MULT=1
MM1000 N_A_197_119#_M1000_d N_A_688_98#_M1000_g N_A_1154_464#_M1017_d VPB PSHORT
+ L=0.15 W=0.64 AD=0.2208 AS=0.136815 PD=1.97 PS=1.23774 NRD=18.4589 NRS=3.0732
+ M=1 R=4.26667 SA=75000.8 SB=75000.3 A=0.096 P=1.58 MULT=1
MM1034 A_1592_424# N_A_1154_464#_M1034_g N_A_1007_366#_M1034_s VPB PSHORT L=0.15
+ W=0.84 AD=0.1134 AS=0.7476 PD=1.11 PS=3.46 NRD=18.7544 NRS=2.3443 M=1 R=5.6
+ SA=75000.8 SB=75001.2 A=0.126 P=1.98 MULT=1
MM1044 N_VPWR_M1044_d N_A_1643_257#_M1044_g A_1592_424# VPB PSHORT L=0.15 W=0.84
+ AD=0.1638 AS=0.1134 PD=1.23 PS=1.11 NRD=2.3443 NRS=18.7544 M=1 R=5.6
+ SA=75001.2 SB=75000.8 A=0.126 P=1.98 MULT=1
MM1013 N_A_1007_366#_M1013_d N_SET_B_M1013_g N_VPWR_M1044_d VPB PSHORT L=0.15
+ W=0.84 AD=0.2478 AS=0.1638 PD=2.27 PS=1.23 NRD=2.3443 NRS=23.443 M=1 R=5.6
+ SA=75001.8 SB=75000.2 A=0.126 P=1.98 MULT=1
MM1036 A_1986_424# N_A_1007_366#_M1036_g N_VPWR_M1036_s VPB PSHORT L=0.15 W=0.84
+ AD=0.1008 AS=0.2478 PD=1.08 PS=2.27 NRD=15.2281 NRS=2.3443 M=1 R=5.6
+ SA=75000.2 SB=75001.1 A=0.126 P=1.98 MULT=1
MM1039 N_A_1997_82#_M1039_d N_A_868_368#_M1039_g A_1986_424# VPB PSHORT L=0.15
+ W=0.84 AD=0.1904 AS=0.1008 PD=1.63333 PS=1.08 NRD=2.3443 NRS=15.2281 M=1 R=5.6
+ SA=75000.6 SB=75000.7 A=0.126 P=1.98 MULT=1
MM1033 A_2171_508# N_A_688_98#_M1033_g N_A_1997_82#_M1039_d VPB PSHORT L=0.15
+ W=0.42 AD=0.0504 AS=0.0952 PD=0.66 PS=0.816667 NRD=30.4759 NRS=44.5417 M=1
+ R=2.8 SA=75001.1 SB=75000.6 A=0.063 P=1.14 MULT=1
MM1050 N_VPWR_M1050_d N_A_2216_410#_M1050_g A_2171_508# VPB PSHORT L=0.15 W=0.42
+ AD=0.1239 AS=0.0504 PD=1.43 PS=0.66 NRD=4.6886 NRS=30.4759 M=1 R=2.8
+ SA=75001.5 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1019 N_VPWR_M1019_d N_SET_B_M1019_g N_A_2216_410#_M1019_s VPB PSHORT L=0.15
+ W=1 AD=0.18 AS=0.295 PD=1.36 PS=2.59 NRD=11.8003 NRS=1.9503 M=1 R=6.66667
+ SA=75000.2 SB=75001.1 A=0.15 P=2.3 MULT=1
MM1046 A_2556_392# N_A_1643_257#_M1046_g N_VPWR_M1019_d VPB PSHORT L=0.15 W=1
+ AD=0.135 AS=0.18 PD=1.27 PS=1.36 NRD=15.7403 NRS=3.9203 M=1 R=6.66667
+ SA=75000.7 SB=75000.6 A=0.15 P=2.3 MULT=1
MM1020 N_A_2216_410#_M1020_d N_A_1997_82#_M1020_g A_2556_392# VPB PSHORT L=0.15
+ W=1 AD=0.295 AS=0.135 PD=2.59 PS=1.27 NRD=1.9503 NRS=15.7403 M=1 R=6.66667
+ SA=75001.1 SB=75000.2 A=0.15 P=2.3 MULT=1
MM1031 N_VPWR_M1031_d N_RESET_B_M1031_g N_A_1643_257#_M1031_s VPB PSHORT L=0.15
+ W=0.64 AD=0.426009 AS=0.1888 PD=1.70545 PS=1.87 NRD=202.378 NRS=3.0732 M=1
+ R=4.26667 SA=75000.2 SB=75001.8 A=0.096 P=1.58 MULT=1
MM1038 N_Q_N_M1038_d N_A_2216_410#_M1038_g N_VPWR_M1031_d VPB PSHORT L=0.15
+ W=1.12 AD=0.168 AS=0.745516 PD=1.42 PS=2.98455 NRD=1.7533 NRS=17.0011 M=1
+ R=7.46667 SA=75001.1 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1042 N_Q_N_M1038_d N_A_2216_410#_M1042_g N_VPWR_M1042_s VPB PSHORT L=0.15
+ W=1.12 AD=0.168 AS=0.3192 PD=1.42 PS=2.81 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.5 SB=75000.2 A=0.168 P=2.54 MULT=1
MM1029 N_VPWR_M1029_d N_A_2216_410#_M1029_g N_A_3272_94#_M1029_s VPB PSHORT
+ L=0.15 W=1 AD=0.192264 AS=0.29 PD=1.41038 PS=2.58 NRD=16.7253 NRS=1.9503 M=1
+ R=6.66667 SA=75000.2 SB=75001.2 A=0.15 P=2.3 MULT=1
MM1006 N_Q_M1006_d N_A_3272_94#_M1006_g N_VPWR_M1029_d VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.215336 PD=1.42 PS=1.57962 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.7 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1011 N_Q_M1006_d N_A_3272_94#_M1011_g N_VPWR_M1011_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.3304 PD=1.42 PS=2.83 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.1 SB=75000.2 A=0.168 P=2.54 MULT=1
DX52_noxref VNB VPB NWDIODE A=34.6332 P=40.96
c_195 VNB 0 3.69273e-19 $X=0 $Y=0
c_376 VPB 0 5.99464e-20 $X=0 $Y=3.085
c_2445 A_206_464# 0 2.57379e-20 $X=1.03 $Y=2.32
c_2924 A_1185_125# 0 1.91291e-19 $X=5.925 $Y=0.625
c_2968 A_1902_125# 0 7.74904e-20 $X=9.51 $Y=0.625
*
.include "sky130_fd_sc_hs__sdfbbn_2.pxi.spice"
*
.ends
*
*
