* File: sky130_fd_sc_hs__a21o_4.pex.spice
* Created: Tue Sep  1 19:49:45 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HS__A21O_4%A_91_48# 1 2 3 12 14 16 19 21 23 26 28 30 33
+ 35 37 38 45 48 50 51 54 56 60 63
c132 60 0 1.83628e-19 $X=4.055 $Y=0.76
c133 56 0 1.66816e-20 $X=3.96 $Y=1.195
c134 48 0 1.44963e-19 $X=2.525 $Y=0.615
c135 33 0 1.61246e-19 $X=1.82 $Y=0.74
r136 69 70 6.74555 $w=3.93e-07 $l=5.5e-08 $layer=POLY_cond $X=1.39 $Y=1.532
+ $X2=1.445 $Y2=1.532
r137 68 69 48.4453 $w=3.93e-07 $l=3.95e-07 $layer=POLY_cond $X=0.995 $Y=1.532
+ $X2=1.39 $Y2=1.532
r138 67 68 4.29262 $w=3.93e-07 $l=3.5e-08 $layer=POLY_cond $X=0.96 $Y=1.532
+ $X2=0.995 $Y2=1.532
r139 64 65 1.83969 $w=3.93e-07 $l=1.5e-08 $layer=POLY_cond $X=0.53 $Y=1.532
+ $X2=0.545 $Y2=1.532
r140 58 60 15.5137 $w=2.58e-07 $l=3.5e-07 $layer=LI1_cond $X=4.09 $Y=1.11
+ $X2=4.09 $Y2=0.76
r141 57 63 8.61065 $w=1.7e-07 $l=1.68953e-07 $layer=LI1_cond $X=3.255 $Y=1.195
+ $X2=3.09 $Y2=1.187
r142 56 58 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=3.96 $Y=1.195
+ $X2=4.09 $Y2=1.11
r143 56 57 45.9947 $w=1.68e-07 $l=7.05e-07 $layer=LI1_cond $X=3.96 $Y=1.195
+ $X2=3.255 $Y2=1.195
r144 52 63 0.89609 $w=3.3e-07 $l=9.3e-08 $layer=LI1_cond $X=3.09 $Y=1.28
+ $X2=3.09 $Y2=1.187
r145 52 54 29.5095 $w=3.28e-07 $l=8.45e-07 $layer=LI1_cond $X=3.09 $Y=1.28
+ $X2=3.09 $Y2=2.125
r146 50 63 8.61065 $w=1.7e-07 $l=1.68464e-07 $layer=LI1_cond $X=2.925 $Y=1.18
+ $X2=3.09 $Y2=1.187
r147 50 51 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=2.925 $Y=1.18
+ $X2=2.61 $Y2=1.18
r148 46 51 7.50571 $w=3.35e-07 $l=1.62019e-07 $layer=LI1_cond $X=2.485 $Y=1.095
+ $X2=2.61 $Y2=1.18
r149 46 48 22.1269 $w=2.48e-07 $l=4.8e-07 $layer=LI1_cond $X=2.485 $Y=1.095
+ $X2=2.485 $Y2=0.615
r150 45 72 9.19847 $w=3.93e-07 $l=7.5e-08 $layer=POLY_cond $X=1.82 $Y=1.532
+ $X2=1.895 $Y2=1.532
r151 45 70 45.9924 $w=3.93e-07 $l=3.75e-07 $layer=POLY_cond $X=1.82 $Y=1.532
+ $X2=1.445 $Y2=1.532
r152 44 45 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.82
+ $Y=1.465 $X2=1.82 $Y2=1.465
r153 41 67 19.6234 $w=3.93e-07 $l=1.6e-07 $layer=POLY_cond $X=0.8 $Y=1.532
+ $X2=0.96 $Y2=1.532
r154 41 65 31.2748 $w=3.93e-07 $l=2.55e-07 $layer=POLY_cond $X=0.8 $Y=1.532
+ $X2=0.545 $Y2=1.532
r155 40 44 35.621 $w=3.28e-07 $l=1.02e-06 $layer=LI1_cond $X=0.8 $Y=1.465
+ $X2=1.82 $Y2=1.465
r156 40 41 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.8
+ $Y=1.465 $X2=0.8 $Y2=1.465
r157 38 46 22.397 $w=3.35e-07 $l=7.78315e-07 $layer=LI1_cond $X=1.87 $Y=1.465
+ $X2=2.485 $Y2=1.095
r158 38 44 1.74613 $w=3.28e-07 $l=5e-08 $layer=LI1_cond $X=1.87 $Y=1.465
+ $X2=1.82 $Y2=1.465
r159 35 72 25.4309 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=1.895 $Y=1.765
+ $X2=1.895 $Y2=1.532
r160 35 37 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.895 $Y=1.765
+ $X2=1.895 $Y2=2.4
r161 31 45 25.4309 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=1.82 $Y=1.3
+ $X2=1.82 $Y2=1.532
r162 31 33 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=1.82 $Y=1.3
+ $X2=1.82 $Y2=0.74
r163 28 70 25.4309 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=1.445 $Y=1.765
+ $X2=1.445 $Y2=1.532
r164 28 30 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.445 $Y=1.765
+ $X2=1.445 $Y2=2.4
r165 24 69 25.4309 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=1.39 $Y=1.3
+ $X2=1.39 $Y2=1.532
r166 24 26 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=1.39 $Y=1.3
+ $X2=1.39 $Y2=0.74
r167 21 68 25.4309 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=0.995 $Y=1.765
+ $X2=0.995 $Y2=1.532
r168 21 23 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.995 $Y=1.765
+ $X2=0.995 $Y2=2.4
r169 17 67 25.4309 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=0.96 $Y=1.3
+ $X2=0.96 $Y2=1.532
r170 17 19 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=0.96 $Y=1.3
+ $X2=0.96 $Y2=0.74
r171 14 65 25.4309 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=0.545 $Y=1.765
+ $X2=0.545 $Y2=1.532
r172 14 16 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.545 $Y=1.765
+ $X2=0.545 $Y2=2.4
r173 10 64 25.4309 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=0.53 $Y=1.3
+ $X2=0.53 $Y2=1.532
r174 10 12 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=0.53 $Y=1.3
+ $X2=0.53 $Y2=0.74
r175 3 54 300 $w=1.7e-07 $l=2.2798e-07 $layer=licon1_PDIFF $count=2 $X=2.94
+ $Y=1.96 $X2=3.09 $Y2=2.125
r176 2 60 182 $w=1.7e-07 $l=4.54643e-07 $layer=licon1_NDIFF $count=1 $X=3.915
+ $Y=0.37 $X2=4.055 $Y2=0.76
r177 1 48 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.385
+ $Y=0.47 $X2=2.525 $Y2=0.615
.ends

.subckt PM_SKY130_FD_SC_HS__A21O_4%B1 3 7 9 11 12 14 15 22
c52 12 0 1.88367e-19 $X=3.315 $Y=1.885
c53 7 0 1.44963e-19 $X=2.74 $Y=0.79
r54 22 23 59.2623 $w=3.66e-07 $l=4.5e-07 $layer=POLY_cond $X=2.865 $Y=1.66
+ $X2=3.315 $Y2=1.66
r55 21 22 16.4617 $w=3.66e-07 $l=1.25e-07 $layer=POLY_cond $X=2.74 $Y=1.66
+ $X2=2.865 $Y2=1.66
r56 19 21 19.7541 $w=3.66e-07 $l=1.5e-07 $layer=POLY_cond $X=2.59 $Y=1.66
+ $X2=2.74 $Y2=1.66
r57 17 19 36.8743 $w=3.66e-07 $l=2.8e-07 $layer=POLY_cond $X=2.31 $Y=1.66
+ $X2=2.59 $Y2=1.66
r58 15 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.59
+ $Y=1.6 $X2=2.59 $Y2=1.6
r59 12 23 23.7042 $w=1.5e-07 $l=2.25e-07 $layer=POLY_cond $X=3.315 $Y=1.885
+ $X2=3.315 $Y2=1.66
r60 12 14 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=3.315 $Y=1.885
+ $X2=3.315 $Y2=2.46
r61 9 22 23.7042 $w=1.5e-07 $l=2.25e-07 $layer=POLY_cond $X=2.865 $Y=1.885
+ $X2=2.865 $Y2=1.66
r62 9 11 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=2.865 $Y=1.885
+ $X2=2.865 $Y2=2.46
r63 5 21 23.7042 $w=1.5e-07 $l=2.25e-07 $layer=POLY_cond $X=2.74 $Y=1.435
+ $X2=2.74 $Y2=1.66
r64 5 7 330.734 $w=1.5e-07 $l=6.45e-07 $layer=POLY_cond $X=2.74 $Y=1.435
+ $X2=2.74 $Y2=0.79
r65 1 17 23.7042 $w=1.5e-07 $l=2.25e-07 $layer=POLY_cond $X=2.31 $Y=1.435
+ $X2=2.31 $Y2=1.66
r66 1 3 330.734 $w=1.5e-07 $l=6.45e-07 $layer=POLY_cond $X=2.31 $Y=1.435
+ $X2=2.31 $Y2=0.79
.ends

.subckt PM_SKY130_FD_SC_HS__A21O_4%A1 1 3 6 8 10 13 15 16 23
c59 13 0 1.9142e-19 $X=4.27 $Y=0.69
r60 23 24 7.06933 $w=3.75e-07 $l=5.5e-08 $layer=POLY_cond $X=4.215 $Y=1.667
+ $X2=4.27 $Y2=1.667
r61 21 23 48.2 $w=3.75e-07 $l=3.75e-07 $layer=POLY_cond $X=3.84 $Y=1.667
+ $X2=4.215 $Y2=1.667
r62 21 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.84
+ $Y=1.615 $X2=3.84 $Y2=1.615
r63 19 21 9.64 $w=3.75e-07 $l=7.5e-08 $layer=POLY_cond $X=3.765 $Y=1.667
+ $X2=3.84 $Y2=1.667
r64 16 22 8.3814 $w=3.28e-07 $l=2.4e-07 $layer=LI1_cond $X=4.08 $Y=1.615
+ $X2=3.84 $Y2=1.615
r65 15 22 8.3814 $w=3.28e-07 $l=2.4e-07 $layer=LI1_cond $X=3.6 $Y=1.615 $X2=3.84
+ $Y2=1.615
r66 11 24 24.2915 $w=1.5e-07 $l=2.17e-07 $layer=POLY_cond $X=4.27 $Y=1.45
+ $X2=4.27 $Y2=1.667
r67 11 13 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=4.27 $Y=1.45
+ $X2=4.27 $Y2=0.69
r68 8 23 24.2915 $w=1.5e-07 $l=2.18e-07 $layer=POLY_cond $X=4.215 $Y=1.885
+ $X2=4.215 $Y2=1.667
r69 8 10 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=4.215 $Y=1.885
+ $X2=4.215 $Y2=2.46
r70 4 21 24.2915 $w=1.5e-07 $l=2.17e-07 $layer=POLY_cond $X=3.84 $Y=1.45
+ $X2=3.84 $Y2=1.667
r71 4 6 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=3.84 $Y=1.45 $X2=3.84
+ $Y2=0.69
r72 1 19 24.2915 $w=1.5e-07 $l=2.18e-07 $layer=POLY_cond $X=3.765 $Y=1.885
+ $X2=3.765 $Y2=1.667
r73 1 3 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=3.765 $Y=1.885
+ $X2=3.765 $Y2=2.46
.ends

.subckt PM_SKY130_FD_SC_HS__A21O_4%A2 2 3 5 8 11 12 14 17 19 26 28
c48 28 0 1.66816e-20 $X=5.13 $Y=1.425
c49 8 0 1.83628e-19 $X=4.7 $Y=0.69
r50 27 28 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=5.115 $Y=1.425
+ $X2=5.13 $Y2=1.425
r51 25 27 65.573 $w=3.3e-07 $l=3.75e-07 $layer=POLY_cond $X=4.74 $Y=1.425
+ $X2=5.115 $Y2=1.425
r52 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.74
+ $Y=1.425 $X2=4.74 $Y2=1.425
r53 23 25 6.99445 $w=3.3e-07 $l=4e-08 $layer=POLY_cond $X=4.7 $Y=1.425 $X2=4.74
+ $Y2=1.425
r54 21 23 6.12014 $w=3.3e-07 $l=3.5e-08 $layer=POLY_cond $X=4.665 $Y=1.425
+ $X2=4.7 $Y2=1.425
r55 19 26 6.24041 $w=4.58e-07 $l=2.4e-07 $layer=LI1_cond $X=4.675 $Y=1.665
+ $X2=4.675 $Y2=1.425
r56 15 28 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.13 $Y=1.26
+ $X2=5.13 $Y2=1.425
r57 15 17 292.277 $w=1.5e-07 $l=5.7e-07 $layer=POLY_cond $X=5.13 $Y=1.26
+ $X2=5.13 $Y2=0.69
r58 12 14 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=5.115 $Y=1.885
+ $X2=5.115 $Y2=2.46
r59 11 12 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=5.115 $Y=1.795
+ $X2=5.115 $Y2=1.885
r60 10 27 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=5.115 $Y=1.59
+ $X2=5.115 $Y2=1.425
r61 10 11 79.6855 $w=1.8e-07 $l=2.05e-07 $layer=POLY_cond $X=5.115 $Y=1.59
+ $X2=5.115 $Y2=1.795
r62 6 23 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.7 $Y=1.26 $X2=4.7
+ $Y2=1.425
r63 6 8 292.277 $w=1.5e-07 $l=5.7e-07 $layer=POLY_cond $X=4.7 $Y=1.26 $X2=4.7
+ $Y2=0.69
r64 3 5 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=4.665 $Y=1.885
+ $X2=4.665 $Y2=2.46
r65 2 3 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=4.665 $Y=1.795 $X2=4.665
+ $Y2=1.885
r66 1 21 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=4.665 $Y=1.59
+ $X2=4.665 $Y2=1.425
r67 1 2 79.6855 $w=1.8e-07 $l=2.05e-07 $layer=POLY_cond $X=4.665 $Y=1.59
+ $X2=4.665 $Y2=1.795
.ends

.subckt PM_SKY130_FD_SC_HS__A21O_4%VPWR 1 2 3 4 5 16 18 22 26 32 36 39 40 42 43
+ 44 46 51 67 68 74 77
c85 32 0 1.88367e-19 $X=3.99 $Y=2.455
r86 77 78 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r87 74 75 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r88 71 72 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r89 67 68 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r90 65 68 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=5.52 $Y2=3.33
r91 64 65 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r92 62 65 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.56 $Y2=3.33
r93 61 62 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r94 59 78 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=2.16 $Y2=3.33
r95 58 61 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=2.64 $Y=3.33 $X2=3.6
+ $Y2=3.33
r96 58 59 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r97 56 77 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.285 $Y=3.33
+ $X2=2.16 $Y2=3.33
r98 56 58 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=2.285 $Y=3.33
+ $X2=2.64 $Y2=3.33
r99 55 78 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r100 55 75 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r101 54 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r102 52 74 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.305 $Y=3.33
+ $X2=1.18 $Y2=3.33
r103 52 54 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=1.305 $Y=3.33
+ $X2=1.68 $Y2=3.33
r104 51 77 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.035 $Y=3.33
+ $X2=2.16 $Y2=3.33
r105 51 54 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=2.035 $Y=3.33
+ $X2=1.68 $Y2=3.33
r106 50 75 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r107 50 72 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r108 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r109 47 71 4.64823 $w=1.7e-07 $l=2.43e-07 $layer=LI1_cond $X=0.485 $Y=3.33
+ $X2=0.242 $Y2=3.33
r110 47 49 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=0.485 $Y=3.33
+ $X2=0.72 $Y2=3.33
r111 46 74 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.055 $Y=3.33
+ $X2=1.18 $Y2=3.33
r112 46 49 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=1.055 $Y=3.33
+ $X2=0.72 $Y2=3.33
r113 44 62 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=2.88 $Y=3.33
+ $X2=3.6 $Y2=3.33
r114 44 59 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.88 $Y=3.33
+ $X2=2.64 $Y2=3.33
r115 42 64 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=4.725 $Y=3.33
+ $X2=4.56 $Y2=3.33
r116 42 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.725 $Y=3.33
+ $X2=4.89 $Y2=3.33
r117 41 67 30.3369 $w=1.68e-07 $l=4.65e-07 $layer=LI1_cond $X=5.055 $Y=3.33
+ $X2=5.52 $Y2=3.33
r118 41 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.055 $Y=3.33
+ $X2=4.89 $Y2=3.33
r119 39 61 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=3.825 $Y=3.33
+ $X2=3.6 $Y2=3.33
r120 39 40 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.825 $Y=3.33
+ $X2=3.95 $Y2=3.33
r121 38 64 31.6417 $w=1.68e-07 $l=4.85e-07 $layer=LI1_cond $X=4.075 $Y=3.33
+ $X2=4.56 $Y2=3.33
r122 38 40 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.075 $Y=3.33
+ $X2=3.95 $Y2=3.33
r123 34 43 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.89 $Y=3.245
+ $X2=4.89 $Y2=3.33
r124 34 36 27.5888 $w=3.28e-07 $l=7.9e-07 $layer=LI1_cond $X=4.89 $Y=3.245
+ $X2=4.89 $Y2=2.455
r125 30 40 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.95 $Y=3.245
+ $X2=3.95 $Y2=3.33
r126 30 32 36.4172 $w=2.48e-07 $l=7.9e-07 $layer=LI1_cond $X=3.95 $Y=3.245
+ $X2=3.95 $Y2=2.455
r127 26 29 32.2684 $w=2.48e-07 $l=7e-07 $layer=LI1_cond $X=2.16 $Y=2.115
+ $X2=2.16 $Y2=2.815
r128 24 77 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.16 $Y=3.245
+ $X2=2.16 $Y2=3.33
r129 24 29 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=2.16 $Y=3.245
+ $X2=2.16 $Y2=2.815
r130 20 74 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.18 $Y=3.245
+ $X2=1.18 $Y2=3.33
r131 20 22 43.3319 $w=2.48e-07 $l=9.4e-07 $layer=LI1_cond $X=1.18 $Y=3.245
+ $X2=1.18 $Y2=2.305
r132 16 71 3.11795 $w=3.3e-07 $l=1.17707e-07 $layer=LI1_cond $X=0.32 $Y=3.245
+ $X2=0.242 $Y2=3.33
r133 16 18 35.621 $w=3.28e-07 $l=1.02e-06 $layer=LI1_cond $X=0.32 $Y=3.245
+ $X2=0.32 $Y2=2.225
r134 5 36 300 $w=1.7e-07 $l=5.65044e-07 $layer=licon1_PDIFF $count=2 $X=4.74
+ $Y=1.96 $X2=4.89 $Y2=2.455
r135 4 32 300 $w=1.7e-07 $l=5.65044e-07 $layer=licon1_PDIFF $count=2 $X=3.84
+ $Y=1.96 $X2=3.99 $Y2=2.455
r136 3 29 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=1.97
+ $Y=1.84 $X2=2.12 $Y2=2.815
r137 3 26 400 $w=1.7e-07 $l=3.4187e-07 $layer=licon1_PDIFF $count=1 $X=1.97
+ $Y=1.84 $X2=2.12 $Y2=2.115
r138 2 22 300 $w=1.7e-07 $l=5.34766e-07 $layer=licon1_PDIFF $count=2 $X=1.07
+ $Y=1.84 $X2=1.22 $Y2=2.305
r139 1 18 300 $w=1.7e-07 $l=4.43114e-07 $layer=licon1_PDIFF $count=2 $X=0.195
+ $Y=1.84 $X2=0.32 $Y2=2.225
.ends

.subckt PM_SKY130_FD_SC_HS__A21O_4%X 1 2 3 4 13 14 15 16 19 23 27 29 33 37 43 44
+ 45 46
c75 27 0 1.61246e-19 $X=1.44 $Y=1.045
r76 45 46 18.5393 $w=2.28e-07 $l=3.7e-07 $layer=LI1_cond $X=0.24 $Y=1.295
+ $X2=0.24 $Y2=1.665
r77 42 46 6.76434 $w=2.28e-07 $l=1.35e-07 $layer=LI1_cond $X=0.24 $Y=1.8
+ $X2=0.24 $Y2=1.665
r78 41 45 8.26753 $w=2.28e-07 $l=1.65e-07 $layer=LI1_cond $X=0.24 $Y=1.13
+ $X2=0.24 $Y2=1.295
r79 37 39 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=1.67 $Y=1.985
+ $X2=1.67 $Y2=2.815
r80 35 37 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=1.67 $Y=1.97
+ $X2=1.67 $Y2=1.985
r81 31 33 20.5135 $w=2.48e-07 $l=4.45e-07 $layer=LI1_cond $X=1.565 $Y=0.96
+ $X2=1.565 $Y2=0.515
r82 30 44 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.855 $Y=1.885
+ $X2=0.77 $Y2=1.885
r83 29 35 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.505 $Y=1.885
+ $X2=1.67 $Y2=1.97
r84 29 30 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=1.505 $Y=1.885
+ $X2=0.855 $Y2=1.885
r85 28 43 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.83 $Y=1.045
+ $X2=0.745 $Y2=1.045
r86 27 31 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.44 $Y=1.045
+ $X2=1.565 $Y2=0.96
r87 27 28 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=1.44 $Y=1.045
+ $X2=0.83 $Y2=1.045
r88 23 25 54.1497 $w=1.68e-07 $l=8.3e-07 $layer=LI1_cond $X=0.77 $Y=1.985
+ $X2=0.77 $Y2=2.815
r89 21 44 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.77 $Y=1.97 $X2=0.77
+ $Y2=1.885
r90 21 23 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=0.77 $Y=1.97
+ $X2=0.77 $Y2=1.985
r91 17 43 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.745 $Y=0.96
+ $X2=0.745 $Y2=1.045
r92 17 19 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=0.745 $Y=0.96
+ $X2=0.745 $Y2=0.515
r93 16 42 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=0.355 $Y=1.885
+ $X2=0.24 $Y2=1.8
r94 15 44 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.685 $Y=1.885
+ $X2=0.77 $Y2=1.885
r95 15 16 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=0.685 $Y=1.885
+ $X2=0.355 $Y2=1.885
r96 14 41 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=0.355 $Y=1.045
+ $X2=0.24 $Y2=1.13
r97 13 43 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.66 $Y=1.045
+ $X2=0.745 $Y2=1.045
r98 13 14 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.66 $Y=1.045
+ $X2=0.355 $Y2=1.045
r99 4 39 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=1.52
+ $Y=1.84 $X2=1.67 $Y2=2.815
r100 4 37 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=1.52
+ $Y=1.84 $X2=1.67 $Y2=1.985
r101 3 25 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=0.62
+ $Y=1.84 $X2=0.77 $Y2=2.815
r102 3 23 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=0.62
+ $Y=1.84 $X2=0.77 $Y2=1.985
r103 2 33 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.465
+ $Y=0.37 $X2=1.605 $Y2=0.515
r104 1 19 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=0.605
+ $Y=0.37 $X2=0.745 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__A21O_4%A_503_392# 1 2 3 4 15 19 20 21 24 25 29 31 33
+ 35 40
r60 33 42 2.9222 $w=2.5e-07 $l=9e-08 $layer=LI1_cond $X=5.38 $Y=2.12 $X2=5.38
+ $Y2=2.03
r61 33 35 32.0379 $w=2.48e-07 $l=6.95e-07 $layer=LI1_cond $X=5.38 $Y=2.12
+ $X2=5.38 $Y2=2.815
r62 32 40 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.525 $Y=2.035
+ $X2=4.4 $Y2=2.035
r63 31 42 4.22096 $w=1.7e-07 $l=1.27475e-07 $layer=LI1_cond $X=5.255 $Y=2.035
+ $X2=5.38 $Y2=2.03
r64 31 32 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=5.255 $Y=2.035
+ $X2=4.525 $Y2=2.035
r65 27 40 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.4 $Y=2.12
+ $X2=4.4 $Y2=2.035
r66 27 29 32.0379 $w=2.48e-07 $l=6.95e-07 $layer=LI1_cond $X=4.4 $Y=2.12 $X2=4.4
+ $Y2=2.815
r67 26 38 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.625 $Y=2.035
+ $X2=3.54 $Y2=2.035
r68 25 40 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.275 $Y=2.035
+ $X2=4.4 $Y2=2.035
r69 25 26 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=4.275 $Y=2.035
+ $X2=3.625 $Y2=2.035
r70 22 24 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=3.54 $Y=2.905 $X2=3.54
+ $Y2=2.815
r71 21 38 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.54 $Y=2.12 $X2=3.54
+ $Y2=2.035
r72 21 24 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=3.54 $Y=2.12
+ $X2=3.54 $Y2=2.815
r73 19 22 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.455 $Y=2.99
+ $X2=3.54 $Y2=2.905
r74 19 20 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=3.455 $Y=2.99
+ $X2=2.725 $Y2=2.99
r75 15 18 32.2684 $w=2.48e-07 $l=7e-07 $layer=LI1_cond $X=2.6 $Y=2.115 $X2=2.6
+ $Y2=2.815
r76 13 20 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=2.6 $Y=2.905
+ $X2=2.725 $Y2=2.99
r77 13 18 4.14879 $w=2.48e-07 $l=9e-08 $layer=LI1_cond $X=2.6 $Y=2.905 $X2=2.6
+ $Y2=2.815
r78 4 42 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=5.19
+ $Y=1.96 $X2=5.34 $Y2=2.105
r79 4 35 400 $w=1.7e-07 $l=9.26971e-07 $layer=licon1_PDIFF $count=1 $X=5.19
+ $Y=1.96 $X2=5.34 $Y2=2.815
r80 3 40 400 $w=1.7e-07 $l=2.17428e-07 $layer=licon1_PDIFF $count=1 $X=4.29
+ $Y=1.96 $X2=4.44 $Y2=2.115
r81 3 29 400 $w=1.7e-07 $l=9.26971e-07 $layer=licon1_PDIFF $count=1 $X=4.29
+ $Y=1.96 $X2=4.44 $Y2=2.815
r82 2 38 400 $w=1.7e-07 $l=2.17428e-07 $layer=licon1_PDIFF $count=1 $X=3.39
+ $Y=1.96 $X2=3.54 $Y2=2.115
r83 2 24 400 $w=1.7e-07 $l=9.26971e-07 $layer=licon1_PDIFF $count=1 $X=3.39
+ $Y=1.96 $X2=3.54 $Y2=2.815
r84 1 18 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=2.515
+ $Y=1.96 $X2=2.64 $Y2=2.815
r85 1 15 400 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_PDIFF $count=1 $X=2.515
+ $Y=1.96 $X2=2.64 $Y2=2.115
.ends

.subckt PM_SKY130_FD_SC_HS__A21O_4%VGND 1 2 3 4 5 16 18 22 26 30 34 37 38 40 41
+ 43 44 46 47 48 67 68
c87 34 0 1.9142e-19 $X=4.915 $Y=0.585
r88 71 72 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r89 67 68 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r90 65 68 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=5.52
+ $Y2=0
r91 64 65 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r92 62 65 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=3.12 $Y=0 $X2=4.56
+ $Y2=0
r93 61 64 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=3.12 $Y=0 $X2=4.56
+ $Y2=0
r94 61 62 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r95 58 59 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r96 56 59 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.64
+ $Y2=0
r97 55 56 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r98 53 56 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r99 53 72 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r100 52 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r101 50 71 4.65971 $w=1.7e-07 $l=2.4e-07 $layer=LI1_cond $X=0.48 $Y=0 $X2=0.24
+ $Y2=0
r102 50 52 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=0.48 $Y=0 $X2=0.72
+ $Y2=0
r103 48 62 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.88 $Y=0
+ $X2=3.12 $Y2=0
r104 48 59 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.88 $Y=0
+ $X2=2.64 $Y2=0
r105 46 64 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=4.75 $Y=0 $X2=4.56
+ $Y2=0
r106 46 47 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.75 $Y=0 $X2=4.915
+ $Y2=0
r107 45 67 28.7059 $w=1.68e-07 $l=4.4e-07 $layer=LI1_cond $X=5.08 $Y=0 $X2=5.52
+ $Y2=0
r108 45 47 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.08 $Y=0 $X2=4.915
+ $Y2=0
r109 44 61 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.955 $Y=0 $X2=3.12
+ $Y2=0
r110 43 58 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=2.79 $Y=0 $X2=2.64
+ $Y2=0
r111 43 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.79 $Y=0 $X2=2.955
+ $Y2=0
r112 40 55 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=1.87 $Y=0 $X2=1.68
+ $Y2=0
r113 40 41 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.87 $Y=0 $X2=1.995
+ $Y2=0
r114 39 58 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=2.12 $Y=0 $X2=2.64
+ $Y2=0
r115 39 41 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.12 $Y=0 $X2=1.995
+ $Y2=0
r116 37 52 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=1.01 $Y=0 $X2=0.72
+ $Y2=0
r117 37 38 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.01 $Y=0 $X2=1.135
+ $Y2=0
r118 36 55 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=1.26 $Y=0 $X2=1.68
+ $Y2=0
r119 36 38 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.26 $Y=0 $X2=1.135
+ $Y2=0
r120 32 47 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.915 $Y=0.085
+ $X2=4.915 $Y2=0
r121 32 34 17.4613 $w=3.28e-07 $l=5e-07 $layer=LI1_cond $X=4.915 $Y=0.085
+ $X2=4.915 $Y2=0.585
r122 28 44 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.955 $Y=0.085
+ $X2=2.955 $Y2=0
r123 28 30 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=2.955 $Y=0.085
+ $X2=2.955 $Y2=0.76
r124 24 41 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.995 $Y=0.085
+ $X2=1.995 $Y2=0
r125 24 26 28.5806 $w=2.48e-07 $l=6.2e-07 $layer=LI1_cond $X=1.995 $Y=0.085
+ $X2=1.995 $Y2=0.705
r126 20 38 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.135 $Y=0.085
+ $X2=1.135 $Y2=0
r127 20 22 24.8928 $w=2.48e-07 $l=5.4e-07 $layer=LI1_cond $X=1.135 $Y=0.085
+ $X2=1.135 $Y2=0.625
r128 16 71 3.10647 $w=3.3e-07 $l=1.16619e-07 $layer=LI1_cond $X=0.315 $Y=0.085
+ $X2=0.24 $Y2=0
r129 16 18 18.8582 $w=3.28e-07 $l=5.4e-07 $layer=LI1_cond $X=0.315 $Y=0.085
+ $X2=0.315 $Y2=0.625
r130 5 34 182 $w=1.7e-07 $l=2.7627e-07 $layer=licon1_NDIFF $count=1 $X=4.775
+ $Y=0.37 $X2=4.915 $Y2=0.585
r131 4 30 182 $w=1.7e-07 $l=3.53129e-07 $layer=licon1_NDIFF $count=1 $X=2.815
+ $Y=0.47 $X2=2.955 $Y2=0.76
r132 3 26 182 $w=1.7e-07 $l=3.98905e-07 $layer=licon1_NDIFF $count=1 $X=1.895
+ $Y=0.37 $X2=2.035 $Y2=0.705
r133 2 22 182 $w=1.7e-07 $l=3.17372e-07 $layer=licon1_NDIFF $count=1 $X=1.035
+ $Y=0.37 $X2=1.175 $Y2=0.625
r134 1 18 182 $w=1.7e-07 $l=3.19374e-07 $layer=licon1_NDIFF $count=1 $X=0.17
+ $Y=0.37 $X2=0.315 $Y2=0.625
.ends

.subckt PM_SKY130_FD_SC_HS__A21O_4%A_700_74# 1 2 3 12 14 15 20 21 24
r37 22 24 18.6696 $w=2.48e-07 $l=4.05e-07 $layer=LI1_cond $X=5.385 $Y=0.92
+ $X2=5.385 $Y2=0.515
r38 20 22 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=5.26 $Y=1.005
+ $X2=5.385 $Y2=0.92
r39 20 21 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=5.26 $Y=1.005
+ $X2=4.57 $Y2=1.005
r40 17 21 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.485 $Y=0.92
+ $X2=4.57 $Y2=1.005
r41 17 19 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=4.485 $Y=0.92
+ $X2=4.485 $Y2=0.515
r42 16 19 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=4.485 $Y=0.425
+ $X2=4.485 $Y2=0.515
r43 14 16 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.4 $Y=0.34
+ $X2=4.485 $Y2=0.425
r44 14 15 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=4.4 $Y=0.34 $X2=3.79
+ $Y2=0.34
r45 10 15 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.625 $Y=0.425
+ $X2=3.79 $Y2=0.34
r46 10 12 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=3.625 $Y=0.425
+ $X2=3.625 $Y2=0.515
r47 3 24 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=5.205
+ $Y=0.37 $X2=5.345 $Y2=0.515
r48 2 19 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=4.345
+ $Y=0.37 $X2=4.485 $Y2=0.515
r49 1 12 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=3.5
+ $Y=0.37 $X2=3.625 $Y2=0.515
.ends

