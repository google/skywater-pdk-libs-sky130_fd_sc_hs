* NGSPICE file created from sky130_fd_sc_hs__fah_1.ext - technology: sky130A

.subckt sky130_fd_sc_hs__fah_1 A B CI VGND VNB VPB VPWR COUT SUM
M1000 a_410_58# a_811_379# a_879_55# VNB nlowvt w=640000u l=150000u
+  ad=2.6395e+11p pd=2.41e+06u as=4.9405e+11p ps=5.22e+06u
M1001 a_83_21# a_811_379# a_231_132# VNB nlowvt w=640000u l=150000u
+  ad=2.375e+11p pd=2.16e+06u as=3.808e+11p ps=3.75e+06u
M1002 a_811_379# a_879_55# a_1849_374# VNB nlowvt w=640000u l=150000u
+  ad=6.528e+11p pd=3.32e+06u as=5.128e+11p ps=4.25e+06u
M1003 a_879_55# a_1023_379# a_410_58# VPB pshort w=840000u l=150000u
+  ad=4.036e+11p pd=3.01e+06u as=5.082e+11p ps=2.89e+06u
M1004 a_1023_379# a_879_55# a_1660_374# VNB nlowvt w=640000u l=150000u
+  ad=4.965e+11p pd=2.98e+06u as=5.157e+11p ps=4.37e+06u
M1005 a_231_132# a_1023_379# a_83_21# VPB pshort w=840000u l=150000u
+  ad=1.10822e+12p pd=6.61e+06u as=7.644e+11p ps=3.5e+06u
M1006 VGND a_410_58# COUT VNB nlowvt w=740000u l=150000u
+  ad=1.8144e+12p pd=1.292e+07u as=2.072e+11p ps=2.04e+06u
M1007 VPWR a_2342_48# a_1660_374# VPB pshort w=1.12e+06u l=150000u
+  ad=2.39732e+12p pd=1.594e+07u as=6.202e+11p ps=5.22e+06u
M1008 a_2342_48# A VPWR VPB pshort w=1e+06u l=150000u
+  ad=3e+11p pd=2.6e+06u as=0p ps=0u
M1009 VPWR A a_1849_374# VPB pshort w=1e+06u l=150000u
+  ad=0p pd=0u as=1.61635e+12p ps=7.38e+06u
M1010 a_231_132# CI VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_2342_48# A VGND VNB nlowvt w=640000u l=150000u
+  ad=1.824e+11p pd=1.85e+06u as=0p ps=0u
M1012 a_231_132# a_1023_379# a_410_58# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_1023_379# a_879_55# a_1849_374# VPB pshort w=840000u l=150000u
+  ad=2.52e+11p pd=2.28e+06u as=0p ps=0u
M1014 VGND A a_1849_374# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VPWR a_410_58# COUT VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=4.6765e+11p ps=3.29e+06u
M1016 a_1660_374# B a_1023_379# VPB pshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_410_58# a_811_379# a_231_132# VPB pshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_811_379# a_879_55# a_1660_374# VPB pshort w=840000u l=150000u
+  ad=2.94e+11p pd=2.38e+06u as=0p ps=0u
M1019 a_1849_374# B a_811_379# VPB pshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_644_104# a_1023_379# a_83_21# VNB nlowvt w=640000u l=150000u
+  ad=4.1745e+11p pd=3.87e+06u as=0p ps=0u
M1021 VPWR a_83_21# SUM VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=3.304e+11p ps=2.83e+06u
M1022 a_231_132# CI VPWR VPB pshort w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_83_21# a_811_379# a_644_104# VPB pshort w=840000u l=150000u
+  ad=0p pd=0u as=5.58725e+11p ps=3.27e+06u
M1024 a_644_104# a_231_132# VPWR VPB pshort w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 VGND a_2342_48# a_1660_374# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 VGND B a_879_55# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 a_1660_374# B a_811_379# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1028 a_644_104# a_231_132# VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1029 VGND a_83_21# SUM VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.072e+11p ps=2.04e+06u
M1030 a_1849_374# B a_1023_379# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1031 VPWR B a_879_55# VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

