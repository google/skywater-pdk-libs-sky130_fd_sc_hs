* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hs__dlrtp_2 D GATE RESET_B VGND VNB VPB VPWR Q
X0 VGND GATE a_235_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X1 a_568_74# a_347_98# a_646_74# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X2 VGND a_27_392# a_568_74# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X3 VPWR a_646_74# a_832_55# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X4 VGND a_832_55# Q VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X5 Q a_832_55# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X6 VPWR GATE a_235_74# VPB sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X7 a_347_98# a_235_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X8 VPWR a_27_392# a_565_392# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=150000u
X9 a_27_392# D VPWR VPB sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X10 a_832_55# a_646_74# a_1060_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X11 a_565_392# a_235_74# a_646_74# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=150000u
X12 a_784_81# a_832_55# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X13 a_646_74# a_347_98# a_756_508# VPB sky130_fd_pr__pfet_01v8 w=420000u l=150000u
X14 VPWR a_832_55# Q VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X15 Q a_832_55# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X16 a_646_74# a_235_74# a_784_81# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X17 a_832_55# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X18 a_27_392# D VGND VNB sky130_fd_pr__nfet_01v8_lvt w=550000u l=150000u
X19 a_347_98# a_235_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X20 a_756_508# a_832_55# VPWR VPB sky130_fd_pr__pfet_01v8 w=420000u l=150000u
X21 a_1060_74# RESET_B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
.ends
