* File: sky130_fd_sc_hs__dlrtn_4.pxi.spice
* Created: Tue Sep  1 20:02:15 2020
* 
x_PM_SKY130_FD_SC_HS__DLRTN_4%D N_D_M1026_g N_D_c_169_n N_D_M1006_g D
+ PM_SKY130_FD_SC_HS__DLRTN_4%D
x_PM_SKY130_FD_SC_HS__DLRTN_4%GATE_N N_GATE_N_M1004_g N_GATE_N_c_198_n
+ N_GATE_N_M1029_g GATE_N PM_SKY130_FD_SC_HS__DLRTN_4%GATE_N
x_PM_SKY130_FD_SC_HS__DLRTN_4%A_232_98# N_A_232_98#_M1004_d N_A_232_98#_M1029_d
+ N_A_232_98#_c_230_n N_A_232_98#_M1022_g N_A_232_98#_M1023_g
+ N_A_232_98#_M1020_g N_A_232_98#_c_239_n N_A_232_98#_M1013_g
+ N_A_232_98#_c_233_n N_A_232_98#_c_241_n N_A_232_98#_c_234_n
+ N_A_232_98#_c_242_n N_A_232_98#_c_243_n N_A_232_98#_c_244_n
+ N_A_232_98#_c_245_n N_A_232_98#_c_246_n N_A_232_98#_c_247_n
+ N_A_232_98#_c_248_n N_A_232_98#_c_235_n N_A_232_98#_c_236_n
+ PM_SKY130_FD_SC_HS__DLRTN_4%A_232_98#
x_PM_SKY130_FD_SC_HS__DLRTN_4%A_27_136# N_A_27_136#_M1026_s N_A_27_136#_M1006_s
+ N_A_27_136#_c_344_n N_A_27_136#_M1028_g N_A_27_136#_c_345_n
+ N_A_27_136#_c_346_n N_A_27_136#_M1021_g N_A_27_136#_c_347_n
+ N_A_27_136#_c_348_n N_A_27_136#_c_349_n N_A_27_136#_c_350_n
+ N_A_27_136#_c_351_n N_A_27_136#_c_355_n N_A_27_136#_c_352_n
+ PM_SKY130_FD_SC_HS__DLRTN_4%A_27_136#
x_PM_SKY130_FD_SC_HS__DLRTN_4%A_348_392# N_A_348_392#_M1023_s
+ N_A_348_392#_M1022_s N_A_348_392#_c_419_n N_A_348_392#_M1007_g
+ N_A_348_392#_M1011_g N_A_348_392#_c_421_n N_A_348_392#_c_428_n
+ N_A_348_392#_c_429_n N_A_348_392#_c_422_n N_A_348_392#_c_423_n
+ N_A_348_392#_c_424_n N_A_348_392#_c_425_n N_A_348_392#_c_430_n
+ PM_SKY130_FD_SC_HS__DLRTN_4%A_348_392#
x_PM_SKY130_FD_SC_HS__DLRTN_4%A_888_406# N_A_888_406#_M1015_s
+ N_A_888_406#_M1003_d N_A_888_406#_M1009_d N_A_888_406#_c_520_n
+ N_A_888_406#_M1000_g N_A_888_406#_M1019_g N_A_888_406#_c_522_n
+ N_A_888_406#_c_523_n N_A_888_406#_c_524_n N_A_888_406#_M1012_g
+ N_A_888_406#_c_507_n N_A_888_406#_M1001_g N_A_888_406#_c_525_n
+ N_A_888_406#_M1014_g N_A_888_406#_M1005_g N_A_888_406#_c_526_n
+ N_A_888_406#_M1016_g N_A_888_406#_M1018_g N_A_888_406#_c_527_n
+ N_A_888_406#_M1017_g N_A_888_406#_M1025_g N_A_888_406#_c_512_n
+ N_A_888_406#_c_529_n N_A_888_406#_c_547_p N_A_888_406#_c_513_n
+ N_A_888_406#_c_514_n N_A_888_406#_c_531_n N_A_888_406#_c_515_n
+ N_A_888_406#_c_564_p N_A_888_406#_c_532_n N_A_888_406#_c_516_n
+ N_A_888_406#_c_517_n N_A_888_406#_c_518_n N_A_888_406#_c_519_n
+ PM_SKY130_FD_SC_HS__DLRTN_4%A_888_406#
x_PM_SKY130_FD_SC_HS__DLRTN_4%A_639_392# N_A_639_392#_M1020_d
+ N_A_639_392#_M1007_d N_A_639_392#_c_702_n N_A_639_392#_c_703_n
+ N_A_639_392#_M1003_g N_A_639_392#_c_695_n N_A_639_392#_M1015_g
+ N_A_639_392#_c_704_n N_A_639_392#_c_705_n N_A_639_392#_M1008_g
+ N_A_639_392#_c_696_n N_A_639_392#_M1027_g N_A_639_392#_c_706_n
+ N_A_639_392#_c_707_n N_A_639_392#_c_708_n N_A_639_392#_c_709_n
+ N_A_639_392#_c_737_n N_A_639_392#_c_697_n N_A_639_392#_c_698_n
+ N_A_639_392#_c_699_n N_A_639_392#_c_700_n N_A_639_392#_c_701_n
+ PM_SKY130_FD_SC_HS__DLRTN_4%A_639_392#
x_PM_SKY130_FD_SC_HS__DLRTN_4%RESET_B N_RESET_B_c_813_n N_RESET_B_c_820_n
+ N_RESET_B_M1009_g N_RESET_B_c_814_n N_RESET_B_M1002_g N_RESET_B_c_815_n
+ N_RESET_B_M1024_g N_RESET_B_c_816_n N_RESET_B_c_822_n N_RESET_B_M1010_g
+ RESET_B RESET_B RESET_B N_RESET_B_c_818_n PM_SKY130_FD_SC_HS__DLRTN_4%RESET_B
x_PM_SKY130_FD_SC_HS__DLRTN_4%VPWR N_VPWR_M1006_d N_VPWR_M1022_d N_VPWR_M1000_d
+ N_VPWR_M1008_s N_VPWR_M1010_s N_VPWR_M1014_d N_VPWR_M1017_d N_VPWR_c_876_n
+ N_VPWR_c_877_n N_VPWR_c_878_n N_VPWR_c_879_n N_VPWR_c_880_n N_VPWR_c_881_n
+ N_VPWR_c_882_n N_VPWR_c_883_n N_VPWR_c_884_n N_VPWR_c_885_n N_VPWR_c_886_n
+ N_VPWR_c_887_n N_VPWR_c_888_n VPWR N_VPWR_c_889_n N_VPWR_c_890_n
+ N_VPWR_c_891_n N_VPWR_c_892_n N_VPWR_c_893_n N_VPWR_c_875_n
+ PM_SKY130_FD_SC_HS__DLRTN_4%VPWR
x_PM_SKY130_FD_SC_HS__DLRTN_4%Q N_Q_M1001_s N_Q_M1018_s N_Q_M1012_s N_Q_M1016_s
+ N_Q_c_994_n N_Q_c_989_n N_Q_c_1001_n N_Q_c_983_n N_Q_c_984_n N_Q_c_990_n
+ N_Q_c_985_n N_Q_c_991_n N_Q_c_992_n Q Q Q N_Q_c_988_n
+ PM_SKY130_FD_SC_HS__DLRTN_4%Q
x_PM_SKY130_FD_SC_HS__DLRTN_4%VGND N_VGND_M1026_d N_VGND_M1023_d N_VGND_M1019_d
+ N_VGND_M1002_s N_VGND_M1001_d N_VGND_M1005_d N_VGND_M1025_d N_VGND_c_1059_n
+ N_VGND_c_1060_n N_VGND_c_1061_n N_VGND_c_1062_n N_VGND_c_1063_n
+ N_VGND_c_1064_n N_VGND_c_1065_n N_VGND_c_1066_n N_VGND_c_1067_n
+ N_VGND_c_1068_n VGND N_VGND_c_1069_n N_VGND_c_1070_n N_VGND_c_1071_n
+ N_VGND_c_1072_n N_VGND_c_1073_n N_VGND_c_1074_n N_VGND_c_1075_n
+ N_VGND_c_1076_n N_VGND_c_1077_n N_VGND_c_1078_n N_VGND_c_1079_n
+ PM_SKY130_FD_SC_HS__DLRTN_4%VGND
x_PM_SKY130_FD_SC_HS__DLRTN_4%A_1035_74# N_A_1035_74#_M1015_d
+ N_A_1035_74#_M1027_d N_A_1035_74#_M1024_d N_A_1035_74#_c_1178_n
+ N_A_1035_74#_c_1179_n N_A_1035_74#_c_1180_n N_A_1035_74#_c_1187_n
+ N_A_1035_74#_c_1198_n N_A_1035_74#_c_1201_n N_A_1035_74#_c_1181_n
+ N_A_1035_74#_c_1182_n PM_SKY130_FD_SC_HS__DLRTN_4%A_1035_74#
cc_1 VNB N_D_M1026_g 0.0308051f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.955
cc_2 VNB N_D_c_169_n 0.0209153f $X=-0.19 $Y=-0.245 $X2=0.535 $Y2=1.895
cc_3 VNB D 0.0020826f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_4 VNB N_GATE_N_M1004_g 0.0293544f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.955
cc_5 VNB N_GATE_N_c_198_n 0.0193941f $X=-0.19 $Y=-0.245 $X2=0.535 $Y2=1.895
cc_6 VNB N_A_232_98#_c_230_n 0.0132575f $X=-0.19 $Y=-0.245 $X2=0.535 $Y2=2.39
cc_7 VNB N_A_232_98#_M1023_g 0.0274357f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.615
cc_8 VNB N_A_232_98#_M1020_g 0.0488807f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A_232_98#_c_233_n 0.0283723f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_232_98#_c_234_n 0.0101216f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_232_98#_c_235_n 0.00493468f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_232_98#_c_236_n 0.00341963f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_27_136#_c_344_n 0.0436196f $X=-0.19 $Y=-0.245 $X2=0.535 $Y2=2.39
cc_14 VNB N_A_27_136#_c_345_n 0.0319058f $X=-0.19 $Y=-0.245 $X2=0.587 $Y2=1.615
cc_15 VNB N_A_27_136#_c_346_n 0.016625f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.615
cc_16 VNB N_A_27_136#_c_347_n 0.00939626f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_27_136#_c_348_n 0.00892374f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_27_136#_c_349_n 0.0118837f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_27_136#_c_350_n 0.00172991f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_27_136#_c_351_n 0.013789f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_27_136#_c_352_n 0.0194302f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_348_392#_c_419_n 0.0176291f $X=-0.19 $Y=-0.245 $X2=0.535 $Y2=2.39
cc_23 VNB N_A_348_392#_M1011_g 0.0321721f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.615
cc_24 VNB N_A_348_392#_c_421_n 0.00310365f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.615
cc_25 VNB N_A_348_392#_c_422_n 0.00312853f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_348_392#_c_423_n 0.0216723f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_348_392#_c_424_n 0.0311398f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_348_392#_c_425_n 0.00437346f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_888_406#_M1019_g 0.064354f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.615
cc_30 VNB N_A_888_406#_c_507_n 0.0119278f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_888_406#_M1001_g 0.0237608f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_888_406#_M1005_g 0.0203648f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_888_406#_M1018_g 0.0203434f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_888_406#_M1025_g 0.0232586f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_888_406#_c_512_n 0.0125745f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_888_406#_c_513_n 0.00197983f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_888_406#_c_514_n 0.00514849f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_888_406#_c_515_n 0.0016809f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_888_406#_c_516_n 0.00244605f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_888_406#_c_517_n 0.00378547f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_888_406#_c_518_n 0.00283662f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_888_406#_c_519_n 0.100101f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_639_392#_c_695_n 0.0192663f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.615
cc_44 VNB N_A_639_392#_c_696_n 0.0163945f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_A_639_392#_c_697_n 0.0130544f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_A_639_392#_c_698_n 0.00257326f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_639_392#_c_699_n 0.0163589f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_639_392#_c_700_n 0.00339515f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A_639_392#_c_701_n 0.101808f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_RESET_B_c_813_n 0.00370409f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.955
cc_51 VNB N_RESET_B_c_814_n 0.016867f $X=-0.19 $Y=-0.245 $X2=0.535 $Y2=2.39
cc_52 VNB N_RESET_B_c_815_n 0.0211591f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_RESET_B_c_816_n 0.00392107f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.615
cc_54 VNB RESET_B 0.0270615f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_RESET_B_c_818_n 0.0651583f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_VPWR_c_875_n 0.40251f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_Q_c_983_n 0.00180794f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_Q_c_984_n 0.00165555f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_Q_c_985_n 0.0017948f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB Q 0.0171365f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB Q 0.0270077f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_Q_c_988_n 0.00306278f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_VGND_c_1059_n 0.0205322f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_VGND_c_1060_n 0.00928694f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_VGND_c_1061_n 0.00340259f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_VGND_c_1062_n 0.0187851f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_VGND_c_1063_n 0.0106146f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_VGND_c_1064_n 0.00250542f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_VGND_c_1065_n 0.012003f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_VGND_c_1066_n 0.0195864f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_VGND_c_1067_n 0.0442338f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_VGND_c_1068_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_VGND_c_1069_n 0.0197505f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_VGND_c_1070_n 0.0374084f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_VGND_c_1071_n 0.0150459f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_VGND_c_1072_n 0.0150459f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_VGND_c_1073_n 0.00631593f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_VGND_c_1074_n 0.0373356f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VNB N_VGND_c_1075_n 0.0305963f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_VGND_c_1076_n 0.00601668f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_81 VNB N_VGND_c_1077_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_82 VNB N_VGND_c_1078_n 0.00604233f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_83 VNB N_VGND_c_1079_n 0.523604f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_84 VNB N_A_1035_74#_c_1178_n 0.0057158f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.615
cc_85 VNB N_A_1035_74#_c_1179_n 0.00450979f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_86 VNB N_A_1035_74#_c_1180_n 0.00418613f $X=-0.19 $Y=-0.245 $X2=0.72
+ $Y2=1.615
cc_87 VNB N_A_1035_74#_c_1181_n 0.00179342f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_88 VNB N_A_1035_74#_c_1182_n 0.0060844f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_89 VPB N_D_c_169_n 0.0421663f $X=-0.19 $Y=1.66 $X2=0.535 $Y2=1.895
cc_90 VPB D 0.00118268f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_91 VPB N_GATE_N_c_198_n 0.0412404f $X=-0.19 $Y=1.66 $X2=0.535 $Y2=1.895
cc_92 VPB N_A_232_98#_c_230_n 0.0326318f $X=-0.19 $Y=1.66 $X2=0.535 $Y2=2.39
cc_93 VPB N_A_232_98#_M1020_g 0.025705f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_94 VPB N_A_232_98#_c_239_n 0.0182628f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_95 VPB N_A_232_98#_c_233_n 0.0188163f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_96 VPB N_A_232_98#_c_241_n 0.0189877f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_97 VPB N_A_232_98#_c_242_n 0.00652108f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_98 VPB N_A_232_98#_c_243_n 0.00569032f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_99 VPB N_A_232_98#_c_244_n 0.00752464f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_100 VPB N_A_232_98#_c_245_n 0.00562663f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_101 VPB N_A_232_98#_c_246_n 0.0441499f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_102 VPB N_A_232_98#_c_247_n 0.0108485f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_103 VPB N_A_232_98#_c_248_n 0.00381884f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_104 VPB N_A_232_98#_c_235_n 0.00748064f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_105 VPB N_A_27_136#_c_344_n 0.0346901f $X=-0.19 $Y=1.66 $X2=0.535 $Y2=2.39
cc_106 VPB N_A_27_136#_c_350_n 0.00161498f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_107 VPB N_A_27_136#_c_355_n 0.0472487f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_108 VPB N_A_27_136#_c_352_n 0.0138207f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_109 VPB N_A_348_392#_c_419_n 0.0347088f $X=-0.19 $Y=1.66 $X2=0.535 $Y2=2.39
cc_110 VPB N_A_348_392#_c_421_n 0.00315769f $X=-0.19 $Y=1.66 $X2=0.72 $Y2=1.615
cc_111 VPB N_A_348_392#_c_428_n 0.0134187f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_112 VPB N_A_348_392#_c_429_n 0.00125987f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_113 VPB N_A_348_392#_c_430_n 0.00231064f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_114 VPB N_A_888_406#_c_520_n 0.0602072f $X=-0.19 $Y=1.66 $X2=0.587 $Y2=1.615
cc_115 VPB N_A_888_406#_M1019_g 0.00498254f $X=-0.19 $Y=1.66 $X2=0.72 $Y2=1.615
cc_116 VPB N_A_888_406#_c_522_n 0.00661911f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_117 VPB N_A_888_406#_c_523_n 0.018987f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_118 VPB N_A_888_406#_c_524_n 0.0165696f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_119 VPB N_A_888_406#_c_525_n 0.0159005f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_120 VPB N_A_888_406#_c_526_n 0.0162f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_121 VPB N_A_888_406#_c_527_n 0.0180336f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_122 VPB N_A_888_406#_c_512_n 0.00607611f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_123 VPB N_A_888_406#_c_529_n 0.0124285f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_124 VPB N_A_888_406#_c_514_n 0.00473446f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_125 VPB N_A_888_406#_c_531_n 0.0072559f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_126 VPB N_A_888_406#_c_532_n 0.0026622f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_127 VPB N_A_888_406#_c_517_n 0.00856512f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_128 VPB N_A_888_406#_c_518_n 0.00126054f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_129 VPB N_A_888_406#_c_519_n 0.0204934f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_130 VPB N_A_639_392#_c_702_n 0.00893862f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_131 VPB N_A_639_392#_c_703_n 0.0211756f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_132 VPB N_A_639_392#_c_704_n 0.00753347f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_133 VPB N_A_639_392#_c_705_n 0.0207738f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_134 VPB N_A_639_392#_c_706_n 0.00185598f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_135 VPB N_A_639_392#_c_707_n 0.00335941f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_136 VPB N_A_639_392#_c_708_n 0.0295182f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_137 VPB N_A_639_392#_c_709_n 0.00146234f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_138 VPB N_A_639_392#_c_700_n 3.15148e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_139 VPB N_A_639_392#_c_701_n 0.0336549f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_140 VPB N_RESET_B_c_813_n 0.0149413f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.955
cc_141 VPB N_RESET_B_c_820_n 0.0213764f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.955
cc_142 VPB N_RESET_B_c_816_n 0.0153017f $X=-0.19 $Y=1.66 $X2=0.59 $Y2=1.615
cc_143 VPB N_RESET_B_c_822_n 0.0229917f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_144 VPB N_VPWR_c_876_n 0.0305251f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_145 VPB N_VPWR_c_877_n 0.0187933f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_146 VPB N_VPWR_c_878_n 0.010569f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_147 VPB N_VPWR_c_879_n 0.0110551f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_148 VPB N_VPWR_c_880_n 0.00526854f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_149 VPB N_VPWR_c_881_n 0.0155194f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_150 VPB N_VPWR_c_882_n 0.0408588f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_151 VPB N_VPWR_c_883_n 0.0184727f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_152 VPB N_VPWR_c_884_n 0.034657f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_153 VPB N_VPWR_c_885_n 0.0205172f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_154 VPB N_VPWR_c_886_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_155 VPB N_VPWR_c_887_n 0.0186948f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_156 VPB N_VPWR_c_888_n 0.00614127f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_157 VPB N_VPWR_c_889_n 0.0183788f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_158 VPB N_VPWR_c_890_n 0.0267333f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_159 VPB N_VPWR_c_891_n 0.0554149f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_160 VPB N_VPWR_c_892_n 0.0253974f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_161 VPB N_VPWR_c_893_n 0.00628551f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_162 VPB N_VPWR_c_875_n 0.131083f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_163 VPB N_Q_c_989_n 0.00257348f $X=-0.19 $Y=1.66 $X2=0.72 $Y2=1.615
cc_164 VPB N_Q_c_990_n 0.00326535f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_165 VPB N_Q_c_991_n 0.0142989f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_166 VPB N_Q_c_992_n 0.00251322f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_167 VPB Q 0.00747008f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_168 N_D_M1026_g N_GATE_N_M1004_g 0.0253063f $X=0.495 $Y=0.955 $X2=0 $Y2=0
cc_169 N_D_c_169_n N_GATE_N_c_198_n 0.0475112f $X=0.535 $Y=1.895 $X2=0 $Y2=0
cc_170 D N_GATE_N_c_198_n 0.00190882f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_171 N_D_c_169_n GATE_N 3.64022e-19 $X=0.535 $Y=1.895 $X2=0 $Y2=0
cc_172 D GATE_N 0.0264214f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_173 N_D_M1026_g N_A_232_98#_c_234_n 0.00111637f $X=0.495 $Y=0.955 $X2=0 $Y2=0
cc_174 N_D_M1026_g N_A_27_136#_c_347_n 0.00496207f $X=0.495 $Y=0.955 $X2=0 $Y2=0
cc_175 N_D_M1026_g N_A_27_136#_c_348_n 0.0102665f $X=0.495 $Y=0.955 $X2=0 $Y2=0
cc_176 N_D_c_169_n N_A_27_136#_c_348_n 0.0028612f $X=0.535 $Y=1.895 $X2=0 $Y2=0
cc_177 D N_A_27_136#_c_348_n 0.00871068f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_178 N_D_M1026_g N_A_27_136#_c_349_n 0.00286883f $X=0.495 $Y=0.955 $X2=0 $Y2=0
cc_179 N_D_M1026_g N_A_27_136#_c_351_n 0.00636483f $X=0.495 $Y=0.955 $X2=0 $Y2=0
cc_180 D N_A_27_136#_c_351_n 0.00131568f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_181 N_D_c_169_n N_A_27_136#_c_355_n 0.0142977f $X=0.535 $Y=1.895 $X2=0 $Y2=0
cc_182 D N_A_27_136#_c_355_n 0.00406903f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_183 N_D_M1026_g N_A_27_136#_c_352_n 0.0126381f $X=0.495 $Y=0.955 $X2=0 $Y2=0
cc_184 N_D_c_169_n N_A_27_136#_c_352_n 0.00408252f $X=0.535 $Y=1.895 $X2=0 $Y2=0
cc_185 D N_A_27_136#_c_352_n 0.0250413f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_186 N_D_c_169_n N_VPWR_c_876_n 0.0111358f $X=0.535 $Y=1.895 $X2=0 $Y2=0
cc_187 D N_VPWR_c_876_n 0.0136154f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_188 N_D_c_169_n N_VPWR_c_890_n 0.00463894f $X=0.535 $Y=1.895 $X2=0 $Y2=0
cc_189 N_D_c_169_n N_VPWR_c_875_n 0.00499434f $X=0.535 $Y=1.895 $X2=0 $Y2=0
cc_190 N_D_M1026_g N_VGND_c_1069_n 0.00301898f $X=0.495 $Y=0.955 $X2=0 $Y2=0
cc_191 N_D_M1026_g N_VGND_c_1079_n 0.00454494f $X=0.495 $Y=0.955 $X2=0 $Y2=0
cc_192 N_GATE_N_M1004_g N_A_232_98#_c_233_n 8.31894e-19 $X=1.085 $Y=0.86 $X2=0
+ $Y2=0
cc_193 N_GATE_N_c_198_n N_A_232_98#_c_233_n 0.0158557f $X=1.085 $Y=1.895 $X2=0
+ $Y2=0
cc_194 GATE_N N_A_232_98#_c_233_n 3.22315e-19 $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_195 N_GATE_N_M1004_g N_A_232_98#_c_234_n 0.00648185f $X=1.085 $Y=0.86 $X2=0
+ $Y2=0
cc_196 N_GATE_N_c_198_n N_A_232_98#_c_234_n 0.00309733f $X=1.085 $Y=1.895 $X2=0
+ $Y2=0
cc_197 GATE_N N_A_232_98#_c_234_n 0.0105236f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_198 N_GATE_N_c_198_n N_A_232_98#_c_242_n 0.00747082f $X=1.085 $Y=1.895 $X2=0
+ $Y2=0
cc_199 N_GATE_N_c_198_n N_A_232_98#_c_244_n 0.00284511f $X=1.085 $Y=1.895 $X2=0
+ $Y2=0
cc_200 N_GATE_N_c_198_n N_A_232_98#_c_247_n 0.00627857f $X=1.085 $Y=1.895 $X2=0
+ $Y2=0
cc_201 GATE_N N_A_232_98#_c_247_n 0.0120807f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_202 N_GATE_N_c_198_n N_A_232_98#_c_248_n 0.00516342f $X=1.085 $Y=1.895 $X2=0
+ $Y2=0
cc_203 N_GATE_N_c_198_n N_A_232_98#_c_235_n 0.00256913f $X=1.085 $Y=1.895 $X2=0
+ $Y2=0
cc_204 GATE_N N_A_232_98#_c_235_n 0.0262364f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_205 N_GATE_N_M1004_g N_A_232_98#_c_236_n 0.00568622f $X=1.085 $Y=0.86 $X2=0
+ $Y2=0
cc_206 N_GATE_N_M1004_g N_A_27_136#_c_347_n 0.00189038f $X=1.085 $Y=0.86 $X2=0
+ $Y2=0
cc_207 N_GATE_N_M1004_g N_A_27_136#_c_348_n 0.0160857f $X=1.085 $Y=0.86 $X2=0
+ $Y2=0
cc_208 GATE_N N_A_27_136#_c_348_n 0.00350057f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_209 N_GATE_N_M1004_g N_A_348_392#_c_425_n 3.18666e-19 $X=1.085 $Y=0.86 $X2=0
+ $Y2=0
cc_210 N_GATE_N_c_198_n N_A_348_392#_c_430_n 8.30263e-19 $X=1.085 $Y=1.895 $X2=0
+ $Y2=0
cc_211 N_GATE_N_c_198_n N_VPWR_c_876_n 0.00899622f $X=1.085 $Y=1.895 $X2=0 $Y2=0
cc_212 N_GATE_N_c_198_n N_VPWR_c_884_n 0.00463088f $X=1.085 $Y=1.895 $X2=0 $Y2=0
cc_213 N_GATE_N_c_198_n N_VPWR_c_875_n 0.00499434f $X=1.085 $Y=1.895 $X2=0 $Y2=0
cc_214 N_GATE_N_M1004_g N_VGND_c_1059_n 0.00546687f $X=1.085 $Y=0.86 $X2=0 $Y2=0
cc_215 N_GATE_N_M1004_g N_VGND_c_1074_n 0.0038134f $X=1.085 $Y=0.86 $X2=0 $Y2=0
cc_216 N_GATE_N_M1004_g N_VGND_c_1079_n 0.00508379f $X=1.085 $Y=0.86 $X2=0 $Y2=0
cc_217 N_A_232_98#_c_230_n N_A_27_136#_c_344_n 0.0347604f $X=2.11 $Y=1.885 $X2=0
+ $Y2=0
cc_218 N_A_232_98#_M1023_g N_A_27_136#_c_344_n 0.0186166f $X=2.18 $Y=0.86 $X2=0
+ $Y2=0
cc_219 N_A_232_98#_c_243_n N_A_27_136#_c_344_n 0.0135192f $X=3.87 $Y=2.685 $X2=0
+ $Y2=0
cc_220 N_A_232_98#_M1020_g N_A_27_136#_c_346_n 0.0548797f $X=3.645 $Y=0.69 $X2=0
+ $Y2=0
cc_221 N_A_232_98#_M1004_d N_A_27_136#_c_348_n 0.0113826f $X=1.16 $Y=0.49 $X2=0
+ $Y2=0
cc_222 N_A_232_98#_M1023_g N_A_27_136#_c_348_n 0.016975f $X=2.18 $Y=0.86 $X2=0
+ $Y2=0
cc_223 N_A_232_98#_c_233_n N_A_27_136#_c_348_n 0.00121652f $X=2.02 $Y=1.585
+ $X2=0 $Y2=0
cc_224 N_A_232_98#_c_234_n N_A_27_136#_c_348_n 0.0339256f $X=1.46 $Y=1.125 $X2=0
+ $Y2=0
cc_225 N_A_232_98#_c_235_n N_A_27_136#_c_348_n 0.00498546f $X=1.7 $Y=1.585 $X2=0
+ $Y2=0
cc_226 N_A_232_98#_M1023_g N_A_27_136#_c_350_n 0.0104291f $X=2.18 $Y=0.86 $X2=0
+ $Y2=0
cc_227 N_A_232_98#_c_243_n N_A_348_392#_M1022_s 0.00903093f $X=3.87 $Y=2.685
+ $X2=0 $Y2=0
cc_228 N_A_232_98#_M1020_g N_A_348_392#_c_419_n 0.0371374f $X=3.645 $Y=0.69
+ $X2=0 $Y2=0
cc_229 N_A_232_98#_c_239_n N_A_348_392#_c_419_n 0.0199787f $X=3.66 $Y=2.445
+ $X2=0 $Y2=0
cc_230 N_A_232_98#_c_243_n N_A_348_392#_c_419_n 0.0130245f $X=3.87 $Y=2.685
+ $X2=0 $Y2=0
cc_231 N_A_232_98#_M1020_g N_A_348_392#_M1011_g 0.0217567f $X=3.645 $Y=0.69
+ $X2=0 $Y2=0
cc_232 N_A_232_98#_c_230_n N_A_348_392#_c_421_n 0.0191894f $X=2.11 $Y=1.885
+ $X2=0 $Y2=0
cc_233 N_A_232_98#_M1023_g N_A_348_392#_c_421_n 0.0059554f $X=2.18 $Y=0.86 $X2=0
+ $Y2=0
cc_234 N_A_232_98#_c_248_n N_A_348_392#_c_421_n 0.00633452f $X=1.387 $Y=1.95
+ $X2=0 $Y2=0
cc_235 N_A_232_98#_c_235_n N_A_348_392#_c_421_n 0.0239603f $X=1.7 $Y=1.585 $X2=0
+ $Y2=0
cc_236 N_A_232_98#_c_236_n N_A_348_392#_c_421_n 0.00698482f $X=1.662 $Y=1.42
+ $X2=0 $Y2=0
cc_237 N_A_232_98#_c_230_n N_A_348_392#_c_428_n 0.00171935f $X=2.11 $Y=1.885
+ $X2=0 $Y2=0
cc_238 N_A_232_98#_M1020_g N_A_348_392#_c_428_n 6.59689e-19 $X=3.645 $Y=0.69
+ $X2=0 $Y2=0
cc_239 N_A_232_98#_c_243_n N_A_348_392#_c_428_n 0.0238346f $X=3.87 $Y=2.685
+ $X2=0 $Y2=0
cc_240 N_A_232_98#_M1020_g N_A_348_392#_c_429_n 0.00172231f $X=3.645 $Y=0.69
+ $X2=0 $Y2=0
cc_241 N_A_232_98#_M1020_g N_A_348_392#_c_423_n 0.0227514f $X=3.645 $Y=0.69
+ $X2=0 $Y2=0
cc_242 N_A_232_98#_M1020_g N_A_348_392#_c_424_n 0.021337f $X=3.645 $Y=0.69 $X2=0
+ $Y2=0
cc_243 N_A_232_98#_c_246_n N_A_348_392#_c_424_n 0.00489746f $X=4.035 $Y=2.195
+ $X2=0 $Y2=0
cc_244 N_A_232_98#_c_230_n N_A_348_392#_c_425_n 3.30391e-19 $X=2.11 $Y=1.885
+ $X2=0 $Y2=0
cc_245 N_A_232_98#_M1023_g N_A_348_392#_c_425_n 0.00658026f $X=2.18 $Y=0.86
+ $X2=0 $Y2=0
cc_246 N_A_232_98#_c_233_n N_A_348_392#_c_425_n 0.00528962f $X=2.02 $Y=1.585
+ $X2=0 $Y2=0
cc_247 N_A_232_98#_c_234_n N_A_348_392#_c_425_n 0.0218242f $X=1.46 $Y=1.125
+ $X2=0 $Y2=0
cc_248 N_A_232_98#_c_235_n N_A_348_392#_c_425_n 0.0049796f $X=1.7 $Y=1.585 $X2=0
+ $Y2=0
cc_249 N_A_232_98#_c_230_n N_A_348_392#_c_430_n 0.0180326f $X=2.11 $Y=1.885
+ $X2=0 $Y2=0
cc_250 N_A_232_98#_c_233_n N_A_348_392#_c_430_n 0.00505569f $X=2.02 $Y=1.585
+ $X2=0 $Y2=0
cc_251 N_A_232_98#_c_243_n N_A_348_392#_c_430_n 0.025107f $X=3.87 $Y=2.685 $X2=0
+ $Y2=0
cc_252 N_A_232_98#_c_248_n N_A_348_392#_c_430_n 0.043983f $X=1.387 $Y=1.95 $X2=0
+ $Y2=0
cc_253 N_A_232_98#_c_235_n N_A_348_392#_c_430_n 0.00527154f $X=1.7 $Y=1.585
+ $X2=0 $Y2=0
cc_254 N_A_232_98#_c_239_n N_A_888_406#_c_520_n 0.00910647f $X=3.66 $Y=2.445
+ $X2=0 $Y2=0
cc_255 N_A_232_98#_c_241_n N_A_888_406#_c_520_n 7.70197e-19 $X=3.66 $Y=2.237
+ $X2=0 $Y2=0
cc_256 N_A_232_98#_c_243_n N_A_888_406#_c_520_n 0.00251181f $X=3.87 $Y=2.685
+ $X2=0 $Y2=0
cc_257 N_A_232_98#_c_245_n N_A_888_406#_c_520_n 0.00637181f $X=4.035 $Y=2.195
+ $X2=0 $Y2=0
cc_258 N_A_232_98#_c_246_n N_A_888_406#_c_520_n 0.0185169f $X=4.035 $Y=2.195
+ $X2=0 $Y2=0
cc_259 N_A_232_98#_c_245_n N_A_888_406#_c_529_n 0.0198487f $X=4.035 $Y=2.195
+ $X2=0 $Y2=0
cc_260 N_A_232_98#_c_246_n N_A_888_406#_c_529_n 0.00136396f $X=4.035 $Y=2.195
+ $X2=0 $Y2=0
cc_261 N_A_232_98#_c_243_n N_A_639_392#_M1007_d 0.00759082f $X=3.87 $Y=2.685
+ $X2=0 $Y2=0
cc_262 N_A_232_98#_c_241_n N_A_639_392#_c_706_n 0.00819203f $X=3.66 $Y=2.237
+ $X2=0 $Y2=0
cc_263 N_A_232_98#_c_243_n N_A_639_392#_c_706_n 0.0323273f $X=3.87 $Y=2.685
+ $X2=0 $Y2=0
cc_264 N_A_232_98#_c_245_n N_A_639_392#_c_706_n 0.0135731f $X=4.035 $Y=2.195
+ $X2=0 $Y2=0
cc_265 N_A_232_98#_M1020_g N_A_639_392#_c_707_n 0.00924763f $X=3.645 $Y=0.69
+ $X2=0 $Y2=0
cc_266 N_A_232_98#_c_241_n N_A_639_392#_c_707_n 0.00734162f $X=3.66 $Y=2.237
+ $X2=0 $Y2=0
cc_267 N_A_232_98#_c_245_n N_A_639_392#_c_707_n 0.016391f $X=4.035 $Y=2.195
+ $X2=0 $Y2=0
cc_268 N_A_232_98#_M1020_g N_A_639_392#_c_708_n 0.00544814f $X=3.645 $Y=0.69
+ $X2=0 $Y2=0
cc_269 N_A_232_98#_c_241_n N_A_639_392#_c_708_n 0.00572766f $X=3.66 $Y=2.237
+ $X2=0 $Y2=0
cc_270 N_A_232_98#_c_245_n N_A_639_392#_c_708_n 0.0262124f $X=4.035 $Y=2.195
+ $X2=0 $Y2=0
cc_271 N_A_232_98#_c_246_n N_A_639_392#_c_708_n 0.0014355f $X=4.035 $Y=2.195
+ $X2=0 $Y2=0
cc_272 N_A_232_98#_M1020_g N_A_639_392#_c_709_n 0.00468408f $X=3.645 $Y=0.69
+ $X2=0 $Y2=0
cc_273 N_A_232_98#_M1020_g N_A_639_392#_c_698_n 0.00113438f $X=3.645 $Y=0.69
+ $X2=0 $Y2=0
cc_274 N_A_232_98#_c_243_n N_VPWR_M1022_d 0.0112306f $X=3.87 $Y=2.685 $X2=0
+ $Y2=0
cc_275 N_A_232_98#_c_244_n N_VPWR_c_876_n 0.0103557f $X=1.63 $Y=2.685 $X2=0
+ $Y2=0
cc_276 N_A_232_98#_c_247_n N_VPWR_c_876_n 0.0265799f $X=1.31 $Y=2.115 $X2=0
+ $Y2=0
cc_277 N_A_232_98#_c_243_n N_VPWR_c_883_n 0.0244015f $X=3.87 $Y=2.685 $X2=0
+ $Y2=0
cc_278 N_A_232_98#_c_230_n N_VPWR_c_884_n 0.00354936f $X=2.11 $Y=1.885 $X2=0
+ $Y2=0
cc_279 N_A_232_98#_c_243_n N_VPWR_c_884_n 0.0118727f $X=3.87 $Y=2.685 $X2=0
+ $Y2=0
cc_280 N_A_232_98#_c_244_n N_VPWR_c_884_n 0.0133755f $X=1.63 $Y=2.685 $X2=0
+ $Y2=0
cc_281 N_A_232_98#_c_239_n N_VPWR_c_891_n 0.00423754f $X=3.66 $Y=2.445 $X2=0
+ $Y2=0
cc_282 N_A_232_98#_c_243_n N_VPWR_c_891_n 0.0306663f $X=3.87 $Y=2.685 $X2=0
+ $Y2=0
cc_283 N_A_232_98#_c_243_n N_VPWR_c_892_n 0.00638198f $X=3.87 $Y=2.685 $X2=0
+ $Y2=0
cc_284 N_A_232_98#_c_230_n N_VPWR_c_875_n 0.0049649f $X=2.11 $Y=1.885 $X2=0
+ $Y2=0
cc_285 N_A_232_98#_c_239_n N_VPWR_c_875_n 0.00539454f $X=3.66 $Y=2.445 $X2=0
+ $Y2=0
cc_286 N_A_232_98#_c_243_n N_VPWR_c_875_n 0.0683661f $X=3.87 $Y=2.685 $X2=0
+ $Y2=0
cc_287 N_A_232_98#_c_244_n N_VPWR_c_875_n 0.0162101f $X=1.63 $Y=2.685 $X2=0
+ $Y2=0
cc_288 N_A_232_98#_c_243_n A_561_392# 0.00429882f $X=3.87 $Y=2.685 $X2=-0.19
+ $Y2=-0.245
cc_289 N_A_232_98#_c_243_n A_747_504# 0.0125198f $X=3.87 $Y=2.685 $X2=-0.19
+ $Y2=-0.245
cc_290 N_A_232_98#_c_245_n A_747_504# 0.00295795f $X=4.035 $Y=2.195 $X2=-0.19
+ $Y2=-0.245
cc_291 N_A_232_98#_M1020_g N_VGND_c_1067_n 0.00461464f $X=3.645 $Y=0.69 $X2=0
+ $Y2=0
cc_292 N_A_232_98#_M1023_g N_VGND_c_1074_n 0.0038134f $X=2.18 $Y=0.86 $X2=0
+ $Y2=0
cc_293 N_A_232_98#_M1023_g N_VGND_c_1075_n 0.0060117f $X=2.18 $Y=0.86 $X2=0
+ $Y2=0
cc_294 N_A_232_98#_M1023_g N_VGND_c_1079_n 0.00508379f $X=2.18 $Y=0.86 $X2=0
+ $Y2=0
cc_295 N_A_232_98#_M1020_g N_VGND_c_1079_n 0.00909529f $X=3.645 $Y=0.69 $X2=0
+ $Y2=0
cc_296 N_A_27_136#_c_348_n N_A_348_392#_M1023_s 0.00727646f $X=2.49 $Y=0.745
+ $X2=-0.19 $Y2=-0.245
cc_297 N_A_27_136#_c_344_n N_A_348_392#_c_419_n 0.0948126f $X=2.73 $Y=1.885
+ $X2=0 $Y2=0
cc_298 N_A_27_136#_c_345_n N_A_348_392#_c_419_n 0.0194757f $X=3.18 $Y=1.16 $X2=0
+ $Y2=0
cc_299 N_A_27_136#_c_350_n N_A_348_392#_c_419_n 6.17168e-19 $X=2.655 $Y=1.505
+ $X2=0 $Y2=0
cc_300 N_A_27_136#_c_344_n N_A_348_392#_c_421_n 0.00554509f $X=2.73 $Y=1.885
+ $X2=0 $Y2=0
cc_301 N_A_27_136#_c_350_n N_A_348_392#_c_421_n 0.0205894f $X=2.655 $Y=1.505
+ $X2=0 $Y2=0
cc_302 N_A_27_136#_c_344_n N_A_348_392#_c_428_n 0.015124f $X=2.73 $Y=1.885 $X2=0
+ $Y2=0
cc_303 N_A_27_136#_c_345_n N_A_348_392#_c_428_n 0.00421244f $X=3.18 $Y=1.16
+ $X2=0 $Y2=0
cc_304 N_A_27_136#_c_350_n N_A_348_392#_c_428_n 0.0190175f $X=2.655 $Y=1.505
+ $X2=0 $Y2=0
cc_305 N_A_27_136#_c_344_n N_A_348_392#_c_429_n 0.002713f $X=2.73 $Y=1.885 $X2=0
+ $Y2=0
cc_306 N_A_27_136#_c_350_n N_A_348_392#_c_429_n 0.00947434f $X=2.655 $Y=1.505
+ $X2=0 $Y2=0
cc_307 N_A_27_136#_c_344_n N_A_348_392#_c_422_n 0.00471724f $X=2.73 $Y=1.885
+ $X2=0 $Y2=0
cc_308 N_A_27_136#_c_345_n N_A_348_392#_c_422_n 0.0195998f $X=3.18 $Y=1.16 $X2=0
+ $Y2=0
cc_309 N_A_27_136#_c_350_n N_A_348_392#_c_422_n 0.0231983f $X=2.655 $Y=1.505
+ $X2=0 $Y2=0
cc_310 N_A_27_136#_c_348_n N_A_348_392#_c_425_n 0.0255532f $X=2.49 $Y=0.745
+ $X2=0 $Y2=0
cc_311 N_A_27_136#_c_350_n N_A_348_392#_c_425_n 0.0132245f $X=2.655 $Y=1.505
+ $X2=0 $Y2=0
cc_312 N_A_27_136#_c_344_n N_A_639_392#_c_706_n 8.12702e-19 $X=2.73 $Y=1.885
+ $X2=0 $Y2=0
cc_313 N_A_27_136#_c_355_n N_VPWR_c_876_n 0.0354172f $X=0.31 $Y=2.115 $X2=0
+ $Y2=0
cc_314 N_A_27_136#_c_344_n N_VPWR_c_883_n 0.00616653f $X=2.73 $Y=1.885 $X2=0
+ $Y2=0
cc_315 N_A_27_136#_c_355_n N_VPWR_c_890_n 0.0106954f $X=0.31 $Y=2.115 $X2=0
+ $Y2=0
cc_316 N_A_27_136#_c_344_n N_VPWR_c_891_n 0.00317855f $X=2.73 $Y=1.885 $X2=0
+ $Y2=0
cc_317 N_A_27_136#_c_344_n N_VPWR_c_875_n 0.00400204f $X=2.73 $Y=1.885 $X2=0
+ $Y2=0
cc_318 N_A_27_136#_c_355_n N_VPWR_c_875_n 0.0129659f $X=0.31 $Y=2.115 $X2=0
+ $Y2=0
cc_319 N_A_27_136#_c_348_n N_VGND_M1026_d 0.0128101f $X=2.49 $Y=0.745 $X2=-0.19
+ $Y2=-0.245
cc_320 N_A_27_136#_c_348_n N_VGND_M1023_d 0.0184416f $X=2.49 $Y=0.745 $X2=0
+ $Y2=0
cc_321 N_A_27_136#_c_350_n N_VGND_M1023_d 0.00868742f $X=2.655 $Y=1.505 $X2=0
+ $Y2=0
cc_322 N_A_27_136#_c_348_n N_VGND_c_1059_n 0.0252207f $X=2.49 $Y=0.745 $X2=0
+ $Y2=0
cc_323 N_A_27_136#_c_346_n N_VGND_c_1067_n 0.00461464f $X=3.255 $Y=1.085 $X2=0
+ $Y2=0
cc_324 N_A_27_136#_c_348_n N_VGND_c_1069_n 0.00286374f $X=2.49 $Y=0.745 $X2=0
+ $Y2=0
cc_325 N_A_27_136#_c_349_n N_VGND_c_1069_n 0.00683196f $X=0.445 $Y=0.745 $X2=0
+ $Y2=0
cc_326 N_A_27_136#_c_348_n N_VGND_c_1074_n 0.0206111f $X=2.49 $Y=0.745 $X2=0
+ $Y2=0
cc_327 N_A_27_136#_c_344_n N_VGND_c_1075_n 0.00827409f $X=2.73 $Y=1.885 $X2=0
+ $Y2=0
cc_328 N_A_27_136#_c_346_n N_VGND_c_1075_n 0.00826245f $X=3.255 $Y=1.085 $X2=0
+ $Y2=0
cc_329 N_A_27_136#_c_348_n N_VGND_c_1075_n 0.0415433f $X=2.49 $Y=0.745 $X2=0
+ $Y2=0
cc_330 N_A_27_136#_c_346_n N_VGND_c_1079_n 0.00913019f $X=3.255 $Y=1.085 $X2=0
+ $Y2=0
cc_331 N_A_27_136#_c_348_n N_VGND_c_1079_n 0.0464148f $X=2.49 $Y=0.745 $X2=0
+ $Y2=0
cc_332 N_A_27_136#_c_349_n N_VGND_c_1079_n 0.0106568f $X=0.445 $Y=0.745 $X2=0
+ $Y2=0
cc_333 N_A_348_392#_M1011_g N_A_888_406#_M1019_g 0.0429601f $X=4.12 $Y=0.58
+ $X2=0 $Y2=0
cc_334 N_A_348_392#_c_423_n N_A_888_406#_M1019_g 0.00125688f $X=4.095 $Y=1.355
+ $X2=0 $Y2=0
cc_335 N_A_348_392#_c_424_n N_A_888_406#_M1019_g 0.0196496f $X=4.095 $Y=1.355
+ $X2=0 $Y2=0
cc_336 N_A_348_392#_c_428_n N_A_639_392#_M1007_d 0.00234683f $X=3.03 $Y=2.005
+ $X2=0 $Y2=0
cc_337 N_A_348_392#_c_419_n N_A_639_392#_c_706_n 0.00386696f $X=3.12 $Y=1.885
+ $X2=0 $Y2=0
cc_338 N_A_348_392#_c_428_n N_A_639_392#_c_706_n 0.0098953f $X=3.03 $Y=2.005
+ $X2=0 $Y2=0
cc_339 N_A_348_392#_c_419_n N_A_639_392#_c_707_n 0.00318155f $X=3.12 $Y=1.885
+ $X2=0 $Y2=0
cc_340 N_A_348_392#_c_428_n N_A_639_392#_c_707_n 0.0141266f $X=3.03 $Y=2.005
+ $X2=0 $Y2=0
cc_341 N_A_348_392#_c_429_n N_A_639_392#_c_707_n 0.00467678f $X=3.195 $Y=1.61
+ $X2=0 $Y2=0
cc_342 N_A_348_392#_c_423_n N_A_639_392#_c_708_n 0.0428459f $X=4.095 $Y=1.355
+ $X2=0 $Y2=0
cc_343 N_A_348_392#_c_424_n N_A_639_392#_c_708_n 0.00393734f $X=4.095 $Y=1.355
+ $X2=0 $Y2=0
cc_344 N_A_348_392#_c_419_n N_A_639_392#_c_709_n 7.76759e-19 $X=3.12 $Y=1.885
+ $X2=0 $Y2=0
cc_345 N_A_348_392#_c_429_n N_A_639_392#_c_709_n 0.0146859f $X=3.195 $Y=1.61
+ $X2=0 $Y2=0
cc_346 N_A_348_392#_c_423_n N_A_639_392#_c_709_n 0.0139157f $X=4.095 $Y=1.355
+ $X2=0 $Y2=0
cc_347 N_A_348_392#_M1011_g N_A_639_392#_c_737_n 0.00924174f $X=4.12 $Y=0.58
+ $X2=0 $Y2=0
cc_348 N_A_348_392#_M1011_g N_A_639_392#_c_697_n 0.00848162f $X=4.12 $Y=0.58
+ $X2=0 $Y2=0
cc_349 N_A_348_392#_c_423_n N_A_639_392#_c_697_n 0.0137779f $X=4.095 $Y=1.355
+ $X2=0 $Y2=0
cc_350 N_A_348_392#_c_424_n N_A_639_392#_c_697_n 0.00145734f $X=4.095 $Y=1.355
+ $X2=0 $Y2=0
cc_351 N_A_348_392#_M1011_g N_A_639_392#_c_698_n 0.00270114f $X=4.12 $Y=0.58
+ $X2=0 $Y2=0
cc_352 N_A_348_392#_c_423_n N_A_639_392#_c_698_n 0.0282919f $X=4.095 $Y=1.355
+ $X2=0 $Y2=0
cc_353 N_A_348_392#_c_424_n N_A_639_392#_c_698_n 0.00266725f $X=4.095 $Y=1.355
+ $X2=0 $Y2=0
cc_354 N_A_348_392#_c_423_n N_A_639_392#_c_699_n 0.00454193f $X=4.095 $Y=1.355
+ $X2=0 $Y2=0
cc_355 N_A_348_392#_c_423_n N_A_639_392#_c_700_n 0.00679878f $X=4.095 $Y=1.355
+ $X2=0 $Y2=0
cc_356 N_A_348_392#_c_428_n N_VPWR_M1022_d 0.00719681f $X=3.03 $Y=2.005 $X2=0
+ $Y2=0
cc_357 N_A_348_392#_c_419_n N_VPWR_c_891_n 0.00317855f $X=3.12 $Y=1.885 $X2=0
+ $Y2=0
cc_358 N_A_348_392#_c_419_n N_VPWR_c_875_n 0.00400854f $X=3.12 $Y=1.885 $X2=0
+ $Y2=0
cc_359 N_A_348_392#_c_428_n A_561_392# 0.00230006f $X=3.03 $Y=2.005 $X2=-0.19
+ $Y2=-0.245
cc_360 N_A_348_392#_M1011_g N_VGND_c_1060_n 0.00161704f $X=4.12 $Y=0.58 $X2=0
+ $Y2=0
cc_361 N_A_348_392#_M1011_g N_VGND_c_1067_n 0.00435336f $X=4.12 $Y=0.58 $X2=0
+ $Y2=0
cc_362 N_A_348_392#_M1011_g N_VGND_c_1079_n 0.00449679f $X=4.12 $Y=0.58 $X2=0
+ $Y2=0
cc_363 N_A_888_406#_c_522_n N_A_639_392#_c_702_n 0.00218622f $X=4.56 $Y=1.825
+ $X2=0 $Y2=0
cc_364 N_A_888_406#_c_547_p N_A_639_392#_c_702_n 0.00592205f $X=5.655 $Y=2.03
+ $X2=0 $Y2=0
cc_365 N_A_888_406#_c_520_n N_A_639_392#_c_703_n 0.00475564f $X=4.53 $Y=2.445
+ $X2=0 $Y2=0
cc_366 N_A_888_406#_c_523_n N_A_639_392#_c_703_n 0.00227358f $X=4.56 $Y=2.03
+ $X2=0 $Y2=0
cc_367 N_A_888_406#_c_529_n N_A_639_392#_c_703_n 0.0239929f $X=5.49 $Y=2.195
+ $X2=0 $Y2=0
cc_368 N_A_888_406#_c_547_p N_A_639_392#_c_703_n 0.00539882f $X=5.655 $Y=2.03
+ $X2=0 $Y2=0
cc_369 N_A_888_406#_c_532_n N_A_639_392#_c_703_n 0.0184945f $X=5.655 $Y=2.245
+ $X2=0 $Y2=0
cc_370 N_A_888_406#_c_513_n N_A_639_392#_c_695_n 0.00270654f $X=5.75 $Y=0.81
+ $X2=0 $Y2=0
cc_371 N_A_888_406#_c_547_p N_A_639_392#_c_704_n 0.00465935f $X=5.655 $Y=2.03
+ $X2=0 $Y2=0
cc_372 N_A_888_406#_c_547_p N_A_639_392#_c_705_n 0.00330952f $X=5.655 $Y=2.03
+ $X2=0 $Y2=0
cc_373 N_A_888_406#_c_532_n N_A_639_392#_c_705_n 0.0126657f $X=5.655 $Y=2.245
+ $X2=0 $Y2=0
cc_374 N_A_888_406#_c_513_n N_A_639_392#_c_696_n 0.00270654f $X=5.75 $Y=0.81
+ $X2=0 $Y2=0
cc_375 N_A_888_406#_c_520_n N_A_639_392#_c_708_n 0.00343847f $X=4.53 $Y=2.445
+ $X2=0 $Y2=0
cc_376 N_A_888_406#_M1019_g N_A_639_392#_c_708_n 0.00639399f $X=4.545 $Y=0.58
+ $X2=0 $Y2=0
cc_377 N_A_888_406#_c_522_n N_A_639_392#_c_708_n 0.00540326f $X=4.56 $Y=1.825
+ $X2=0 $Y2=0
cc_378 N_A_888_406#_c_523_n N_A_639_392#_c_708_n 0.00447383f $X=4.56 $Y=2.03
+ $X2=0 $Y2=0
cc_379 N_A_888_406#_c_529_n N_A_639_392#_c_708_n 0.0634347f $X=5.49 $Y=2.195
+ $X2=0 $Y2=0
cc_380 N_A_888_406#_c_547_p N_A_639_392#_c_708_n 0.00415403f $X=5.655 $Y=2.03
+ $X2=0 $Y2=0
cc_381 N_A_888_406#_c_564_p N_A_639_392#_c_708_n 0.00582853f $X=5.662 $Y=1.705
+ $X2=0 $Y2=0
cc_382 N_A_888_406#_M1019_g N_A_639_392#_c_737_n 0.00164878f $X=4.545 $Y=0.58
+ $X2=0 $Y2=0
cc_383 N_A_888_406#_M1019_g N_A_639_392#_c_697_n 0.0153705f $X=4.545 $Y=0.58
+ $X2=0 $Y2=0
cc_384 N_A_888_406#_M1019_g N_A_639_392#_c_699_n 0.00636966f $X=4.545 $Y=0.58
+ $X2=0 $Y2=0
cc_385 N_A_888_406#_c_513_n N_A_639_392#_c_699_n 0.00674443f $X=5.75 $Y=0.81
+ $X2=0 $Y2=0
cc_386 N_A_888_406#_M1019_g N_A_639_392#_c_700_n 0.00603966f $X=4.545 $Y=0.58
+ $X2=0 $Y2=0
cc_387 N_A_888_406#_c_513_n N_A_639_392#_c_700_n 0.00989338f $X=5.75 $Y=0.81
+ $X2=0 $Y2=0
cc_388 N_A_888_406#_c_564_p N_A_639_392#_c_700_n 0.00388535f $X=5.662 $Y=1.705
+ $X2=0 $Y2=0
cc_389 N_A_888_406#_M1019_g N_A_639_392#_c_701_n 0.0267316f $X=4.545 $Y=0.58
+ $X2=0 $Y2=0
cc_390 N_A_888_406#_c_522_n N_A_639_392#_c_701_n 0.00302799f $X=4.56 $Y=1.825
+ $X2=0 $Y2=0
cc_391 N_A_888_406#_c_529_n N_A_639_392#_c_701_n 0.00690333f $X=5.49 $Y=2.195
+ $X2=0 $Y2=0
cc_392 N_A_888_406#_c_513_n N_A_639_392#_c_701_n 0.0295448f $X=5.75 $Y=0.81
+ $X2=0 $Y2=0
cc_393 N_A_888_406#_c_514_n N_A_639_392#_c_701_n 0.0183112f $X=6.49 $Y=1.705
+ $X2=0 $Y2=0
cc_394 N_A_888_406#_c_564_p N_A_639_392#_c_701_n 0.0208109f $X=5.662 $Y=1.705
+ $X2=0 $Y2=0
cc_395 N_A_888_406#_c_547_p N_RESET_B_c_813_n 7.19635e-19 $X=5.655 $Y=2.03 $X2=0
+ $Y2=0
cc_396 N_A_888_406#_c_514_n N_RESET_B_c_813_n 0.0171472f $X=6.49 $Y=1.705 $X2=0
+ $Y2=0
cc_397 N_A_888_406#_c_531_n N_RESET_B_c_813_n 0.00387749f $X=6.655 $Y=2.245
+ $X2=0 $Y2=0
cc_398 N_A_888_406#_c_531_n N_RESET_B_c_820_n 0.00592411f $X=6.655 $Y=2.245
+ $X2=0 $Y2=0
cc_399 N_A_888_406#_c_532_n N_RESET_B_c_820_n 4.44891e-19 $X=5.655 $Y=2.245
+ $X2=0 $Y2=0
cc_400 N_A_888_406#_c_524_n N_RESET_B_c_816_n 0.00755309f $X=7.485 $Y=1.765
+ $X2=0 $Y2=0
cc_401 N_A_888_406#_c_531_n N_RESET_B_c_816_n 0.00457747f $X=6.655 $Y=2.245
+ $X2=0 $Y2=0
cc_402 N_A_888_406#_c_516_n N_RESET_B_c_816_n 0.00268108f $X=6.655 $Y=1.705
+ $X2=0 $Y2=0
cc_403 N_A_888_406#_c_517_n N_RESET_B_c_816_n 0.0148205f $X=7.725 $Y=1.545 $X2=0
+ $Y2=0
cc_404 N_A_888_406#_c_524_n N_RESET_B_c_822_n 0.0191149f $X=7.485 $Y=1.765 $X2=0
+ $Y2=0
cc_405 N_A_888_406#_c_531_n N_RESET_B_c_822_n 0.00612164f $X=6.655 $Y=2.245
+ $X2=0 $Y2=0
cc_406 N_A_888_406#_M1001_g RESET_B 0.0071116f $X=7.815 $Y=0.74 $X2=0 $Y2=0
cc_407 N_A_888_406#_c_512_n RESET_B 0.00497165f $X=7.485 $Y=1.555 $X2=0 $Y2=0
cc_408 N_A_888_406#_c_513_n RESET_B 0.0106111f $X=5.75 $Y=0.81 $X2=0 $Y2=0
cc_409 N_A_888_406#_c_514_n RESET_B 0.0121777f $X=6.49 $Y=1.705 $X2=0 $Y2=0
cc_410 N_A_888_406#_c_516_n RESET_B 0.0277859f $X=6.655 $Y=1.705 $X2=0 $Y2=0
cc_411 N_A_888_406#_c_517_n RESET_B 0.056296f $X=7.725 $Y=1.545 $X2=0 $Y2=0
cc_412 N_A_888_406#_c_518_n RESET_B 0.0138646f $X=7.895 $Y=1.545 $X2=0 $Y2=0
cc_413 N_A_888_406#_c_519_n RESET_B 0.00110961f $X=8.985 $Y=1.532 $X2=0 $Y2=0
cc_414 N_A_888_406#_c_512_n N_RESET_B_c_818_n 0.0102534f $X=7.485 $Y=1.555 $X2=0
+ $Y2=0
cc_415 N_A_888_406#_c_513_n N_RESET_B_c_818_n 0.00126612f $X=5.75 $Y=0.81 $X2=0
+ $Y2=0
cc_416 N_A_888_406#_c_516_n N_RESET_B_c_818_n 0.00490094f $X=6.655 $Y=1.705
+ $X2=0 $Y2=0
cc_417 N_A_888_406#_c_529_n N_VPWR_M1000_d 0.00400885f $X=5.49 $Y=2.195 $X2=0
+ $Y2=0
cc_418 N_A_888_406#_c_532_n N_VPWR_c_877_n 0.0134657f $X=5.655 $Y=2.245 $X2=0
+ $Y2=0
cc_419 N_A_888_406#_c_514_n N_VPWR_c_878_n 0.0189103f $X=6.49 $Y=1.705 $X2=0
+ $Y2=0
cc_420 N_A_888_406#_c_531_n N_VPWR_c_878_n 0.0346007f $X=6.655 $Y=2.245 $X2=0
+ $Y2=0
cc_421 N_A_888_406#_c_532_n N_VPWR_c_878_n 0.035855f $X=5.655 $Y=2.245 $X2=0
+ $Y2=0
cc_422 N_A_888_406#_c_524_n N_VPWR_c_879_n 0.00792141f $X=7.485 $Y=1.765 $X2=0
+ $Y2=0
cc_423 N_A_888_406#_c_531_n N_VPWR_c_879_n 0.0300477f $X=6.655 $Y=2.245 $X2=0
+ $Y2=0
cc_424 N_A_888_406#_c_517_n N_VPWR_c_879_n 0.0180194f $X=7.725 $Y=1.545 $X2=0
+ $Y2=0
cc_425 N_A_888_406#_c_525_n N_VPWR_c_880_n 0.00542823f $X=7.935 $Y=1.765 $X2=0
+ $Y2=0
cc_426 N_A_888_406#_c_526_n N_VPWR_c_880_n 0.0107122f $X=8.435 $Y=1.765 $X2=0
+ $Y2=0
cc_427 N_A_888_406#_c_527_n N_VPWR_c_880_n 4.77279e-19 $X=8.985 $Y=1.765 $X2=0
+ $Y2=0
cc_428 N_A_888_406#_c_526_n N_VPWR_c_882_n 5.09864e-19 $X=8.435 $Y=1.765 $X2=0
+ $Y2=0
cc_429 N_A_888_406#_c_527_n N_VPWR_c_882_n 0.0157557f $X=8.985 $Y=1.765 $X2=0
+ $Y2=0
cc_430 N_A_888_406#_c_531_n N_VPWR_c_885_n 0.0135468f $X=6.655 $Y=2.245 $X2=0
+ $Y2=0
cc_431 N_A_888_406#_c_524_n N_VPWR_c_887_n 0.00445602f $X=7.485 $Y=1.765 $X2=0
+ $Y2=0
cc_432 N_A_888_406#_c_525_n N_VPWR_c_887_n 0.00445602f $X=7.935 $Y=1.765 $X2=0
+ $Y2=0
cc_433 N_A_888_406#_c_526_n N_VPWR_c_889_n 0.00413917f $X=8.435 $Y=1.765 $X2=0
+ $Y2=0
cc_434 N_A_888_406#_c_527_n N_VPWR_c_889_n 0.00413917f $X=8.985 $Y=1.765 $X2=0
+ $Y2=0
cc_435 N_A_888_406#_c_520_n N_VPWR_c_891_n 0.00505726f $X=4.53 $Y=2.445 $X2=0
+ $Y2=0
cc_436 N_A_888_406#_c_520_n N_VPWR_c_892_n 0.0229382f $X=4.53 $Y=2.445 $X2=0
+ $Y2=0
cc_437 N_A_888_406#_c_529_n N_VPWR_c_892_n 0.0408836f $X=5.49 $Y=2.195 $X2=0
+ $Y2=0
cc_438 N_A_888_406#_c_532_n N_VPWR_c_892_n 0.0132892f $X=5.655 $Y=2.245 $X2=0
+ $Y2=0
cc_439 N_A_888_406#_c_520_n N_VPWR_c_875_n 0.00519803f $X=4.53 $Y=2.445 $X2=0
+ $Y2=0
cc_440 N_A_888_406#_c_524_n N_VPWR_c_875_n 0.00861719f $X=7.485 $Y=1.765 $X2=0
+ $Y2=0
cc_441 N_A_888_406#_c_525_n N_VPWR_c_875_n 0.00857378f $X=7.935 $Y=1.765 $X2=0
+ $Y2=0
cc_442 N_A_888_406#_c_526_n N_VPWR_c_875_n 0.00818606f $X=8.435 $Y=1.765 $X2=0
+ $Y2=0
cc_443 N_A_888_406#_c_527_n N_VPWR_c_875_n 0.00818606f $X=8.985 $Y=1.765 $X2=0
+ $Y2=0
cc_444 N_A_888_406#_c_531_n N_VPWR_c_875_n 0.0119671f $X=6.655 $Y=2.245 $X2=0
+ $Y2=0
cc_445 N_A_888_406#_c_532_n N_VPWR_c_875_n 0.0119432f $X=5.655 $Y=2.245 $X2=0
+ $Y2=0
cc_446 N_A_888_406#_c_524_n N_Q_c_994_n 0.00320237f $X=7.485 $Y=1.765 $X2=0
+ $Y2=0
cc_447 N_A_888_406#_c_507_n N_Q_c_994_n 0.0012834f $X=7.74 $Y=1.555 $X2=0 $Y2=0
cc_448 N_A_888_406#_c_525_n N_Q_c_994_n 4.27055e-19 $X=7.935 $Y=1.765 $X2=0
+ $Y2=0
cc_449 N_A_888_406#_c_517_n N_Q_c_994_n 0.0228311f $X=7.725 $Y=1.545 $X2=0 $Y2=0
cc_450 N_A_888_406#_c_524_n N_Q_c_989_n 0.00856892f $X=7.485 $Y=1.765 $X2=0
+ $Y2=0
cc_451 N_A_888_406#_c_525_n N_Q_c_989_n 0.0101227f $X=7.935 $Y=1.765 $X2=0 $Y2=0
cc_452 N_A_888_406#_c_526_n N_Q_c_989_n 6.19463e-19 $X=8.435 $Y=1.765 $X2=0
+ $Y2=0
cc_453 N_A_888_406#_c_525_n N_Q_c_1001_n 0.0129047f $X=7.935 $Y=1.765 $X2=0
+ $Y2=0
cc_454 N_A_888_406#_c_526_n N_Q_c_1001_n 0.0150276f $X=8.435 $Y=1.765 $X2=0
+ $Y2=0
cc_455 N_A_888_406#_c_515_n N_Q_c_1001_n 0.0248579f $X=8.91 $Y=1.465 $X2=0 $Y2=0
cc_456 N_A_888_406#_c_518_n N_Q_c_1001_n 0.00144113f $X=7.895 $Y=1.545 $X2=0
+ $Y2=0
cc_457 N_A_888_406#_c_519_n N_Q_c_1001_n 0.0070359f $X=8.985 $Y=1.532 $X2=0
+ $Y2=0
cc_458 N_A_888_406#_M1001_g N_Q_c_983_n 2.84024e-19 $X=7.815 $Y=0.74 $X2=0 $Y2=0
cc_459 N_A_888_406#_M1005_g N_Q_c_983_n 2.84024e-19 $X=8.245 $Y=0.74 $X2=0 $Y2=0
cc_460 N_A_888_406#_M1001_g N_Q_c_984_n 4.35498e-19 $X=7.815 $Y=0.74 $X2=0 $Y2=0
cc_461 N_A_888_406#_c_515_n N_Q_c_984_n 0.0160251f $X=8.91 $Y=1.465 $X2=0 $Y2=0
cc_462 N_A_888_406#_c_519_n N_Q_c_984_n 0.00247261f $X=8.985 $Y=1.532 $X2=0
+ $Y2=0
cc_463 N_A_888_406#_c_526_n N_Q_c_990_n 0.00513007f $X=8.435 $Y=1.765 $X2=0
+ $Y2=0
cc_464 N_A_888_406#_c_527_n N_Q_c_990_n 0.00608252f $X=8.985 $Y=1.765 $X2=0
+ $Y2=0
cc_465 N_A_888_406#_M1018_g N_Q_c_985_n 2.84024e-19 $X=8.675 $Y=0.74 $X2=0 $Y2=0
cc_466 N_A_888_406#_M1025_g N_Q_c_985_n 2.84024e-19 $X=9.105 $Y=0.74 $X2=0 $Y2=0
cc_467 N_A_888_406#_c_527_n N_Q_c_991_n 0.0153745f $X=8.985 $Y=1.765 $X2=0 $Y2=0
cc_468 N_A_888_406#_c_515_n N_Q_c_991_n 0.0144694f $X=8.91 $Y=1.465 $X2=0 $Y2=0
cc_469 N_A_888_406#_c_519_n N_Q_c_991_n 0.00397537f $X=8.985 $Y=1.532 $X2=0
+ $Y2=0
cc_470 N_A_888_406#_c_526_n N_Q_c_992_n 0.00187133f $X=8.435 $Y=1.765 $X2=0
+ $Y2=0
cc_471 N_A_888_406#_c_527_n N_Q_c_992_n 5.64117e-19 $X=8.985 $Y=1.765 $X2=0
+ $Y2=0
cc_472 N_A_888_406#_c_515_n N_Q_c_992_n 0.0276613f $X=8.91 $Y=1.465 $X2=0 $Y2=0
cc_473 N_A_888_406#_c_519_n N_Q_c_992_n 0.00880056f $X=8.985 $Y=1.532 $X2=0
+ $Y2=0
cc_474 N_A_888_406#_M1025_g Q 0.0178501f $X=9.105 $Y=0.74 $X2=0 $Y2=0
cc_475 N_A_888_406#_c_519_n Q 0.00242112f $X=8.985 $Y=1.532 $X2=0 $Y2=0
cc_476 N_A_888_406#_c_527_n Q 0.00118721f $X=8.985 $Y=1.765 $X2=0 $Y2=0
cc_477 N_A_888_406#_M1025_g Q 0.0112629f $X=9.105 $Y=0.74 $X2=0 $Y2=0
cc_478 N_A_888_406#_c_515_n Q 0.0267934f $X=8.91 $Y=1.465 $X2=0 $Y2=0
cc_479 N_A_888_406#_c_519_n Q 0.00620365f $X=8.985 $Y=1.532 $X2=0 $Y2=0
cc_480 N_A_888_406#_M1005_g N_Q_c_988_n 0.0124418f $X=8.245 $Y=0.74 $X2=0 $Y2=0
cc_481 N_A_888_406#_M1018_g N_Q_c_988_n 0.0124434f $X=8.675 $Y=0.74 $X2=0 $Y2=0
cc_482 N_A_888_406#_c_515_n N_Q_c_988_n 0.071138f $X=8.91 $Y=1.465 $X2=0 $Y2=0
cc_483 N_A_888_406#_c_519_n N_Q_c_988_n 0.00263605f $X=8.985 $Y=1.532 $X2=0
+ $Y2=0
cc_484 N_A_888_406#_M1019_g N_VGND_c_1060_n 0.011225f $X=4.545 $Y=0.58 $X2=0
+ $Y2=0
cc_485 N_A_888_406#_M1001_g N_VGND_c_1063_n 0.0116379f $X=7.815 $Y=0.74 $X2=0
+ $Y2=0
cc_486 N_A_888_406#_M1005_g N_VGND_c_1063_n 5.21765e-19 $X=8.245 $Y=0.74 $X2=0
+ $Y2=0
cc_487 N_A_888_406#_c_512_n N_VGND_c_1063_n 0.00288892f $X=7.485 $Y=1.555 $X2=0
+ $Y2=0
cc_488 N_A_888_406#_c_517_n N_VGND_c_1063_n 0.003848f $X=7.725 $Y=1.545 $X2=0
+ $Y2=0
cc_489 N_A_888_406#_c_518_n N_VGND_c_1063_n 0.00148206f $X=7.895 $Y=1.545 $X2=0
+ $Y2=0
cc_490 N_A_888_406#_M1001_g N_VGND_c_1064_n 4.765e-19 $X=7.815 $Y=0.74 $X2=0
+ $Y2=0
cc_491 N_A_888_406#_M1005_g N_VGND_c_1064_n 0.00952924f $X=8.245 $Y=0.74 $X2=0
+ $Y2=0
cc_492 N_A_888_406#_M1018_g N_VGND_c_1064_n 0.00952924f $X=8.675 $Y=0.74 $X2=0
+ $Y2=0
cc_493 N_A_888_406#_M1025_g N_VGND_c_1064_n 4.765e-19 $X=9.105 $Y=0.74 $X2=0
+ $Y2=0
cc_494 N_A_888_406#_M1018_g N_VGND_c_1066_n 4.31235e-19 $X=8.675 $Y=0.74 $X2=0
+ $Y2=0
cc_495 N_A_888_406#_M1025_g N_VGND_c_1066_n 0.00824245f $X=9.105 $Y=0.74 $X2=0
+ $Y2=0
cc_496 N_A_888_406#_M1019_g N_VGND_c_1067_n 0.00383152f $X=4.545 $Y=0.58 $X2=0
+ $Y2=0
cc_497 N_A_888_406#_M1001_g N_VGND_c_1071_n 0.00383152f $X=7.815 $Y=0.74 $X2=0
+ $Y2=0
cc_498 N_A_888_406#_M1005_g N_VGND_c_1071_n 0.00383152f $X=8.245 $Y=0.74 $X2=0
+ $Y2=0
cc_499 N_A_888_406#_M1018_g N_VGND_c_1072_n 0.00383152f $X=8.675 $Y=0.74 $X2=0
+ $Y2=0
cc_500 N_A_888_406#_M1025_g N_VGND_c_1072_n 0.00383152f $X=9.105 $Y=0.74 $X2=0
+ $Y2=0
cc_501 N_A_888_406#_M1019_g N_VGND_c_1079_n 0.00386109f $X=4.545 $Y=0.58 $X2=0
+ $Y2=0
cc_502 N_A_888_406#_M1001_g N_VGND_c_1079_n 0.0075754f $X=7.815 $Y=0.74 $X2=0
+ $Y2=0
cc_503 N_A_888_406#_M1005_g N_VGND_c_1079_n 0.0075754f $X=8.245 $Y=0.74 $X2=0
+ $Y2=0
cc_504 N_A_888_406#_M1018_g N_VGND_c_1079_n 0.0075754f $X=8.675 $Y=0.74 $X2=0
+ $Y2=0
cc_505 N_A_888_406#_M1025_g N_VGND_c_1079_n 0.00375577f $X=9.105 $Y=0.74 $X2=0
+ $Y2=0
cc_506 N_A_888_406#_M1019_g N_A_1035_74#_c_1178_n 0.00431882f $X=4.545 $Y=0.58
+ $X2=0 $Y2=0
cc_507 N_A_888_406#_M1015_s N_A_1035_74#_c_1179_n 0.00169477f $X=5.61 $Y=0.37
+ $X2=0 $Y2=0
cc_508 N_A_888_406#_c_513_n N_A_1035_74#_c_1179_n 0.0126348f $X=5.75 $Y=0.81
+ $X2=0 $Y2=0
cc_509 N_A_888_406#_M1019_g N_A_1035_74#_c_1180_n 6.04331e-19 $X=4.545 $Y=0.58
+ $X2=0 $Y2=0
cc_510 N_A_888_406#_c_514_n N_A_1035_74#_c_1187_n 0.00658578f $X=6.49 $Y=1.705
+ $X2=0 $Y2=0
cc_511 N_A_888_406#_M1001_g N_A_1035_74#_c_1182_n 7.13159e-19 $X=7.815 $Y=0.74
+ $X2=0 $Y2=0
cc_512 N_A_639_392#_c_704_n N_RESET_B_c_813_n 0.0078189f $X=5.88 $Y=1.935 $X2=0
+ $Y2=0
cc_513 N_A_639_392#_c_705_n N_RESET_B_c_820_n 0.0271469f $X=5.88 $Y=2.025 $X2=0
+ $Y2=0
cc_514 N_A_639_392#_c_696_n N_RESET_B_c_814_n 0.00870882f $X=5.965 $Y=1.12 $X2=0
+ $Y2=0
cc_515 N_A_639_392#_c_701_n RESET_B 0.00162569f $X=5.88 $Y=1.455 $X2=0 $Y2=0
cc_516 N_A_639_392#_c_701_n N_RESET_B_c_818_n 0.0229083f $X=5.88 $Y=1.455 $X2=0
+ $Y2=0
cc_517 N_A_639_392#_c_703_n N_VPWR_c_877_n 0.00548284f $X=5.43 $Y=2.025 $X2=0
+ $Y2=0
cc_518 N_A_639_392#_c_705_n N_VPWR_c_877_n 0.00548284f $X=5.88 $Y=2.025 $X2=0
+ $Y2=0
cc_519 N_A_639_392#_c_705_n N_VPWR_c_878_n 0.00656899f $X=5.88 $Y=2.025 $X2=0
+ $Y2=0
cc_520 N_A_639_392#_c_703_n N_VPWR_c_892_n 0.0100886f $X=5.43 $Y=2.025 $X2=0
+ $Y2=0
cc_521 N_A_639_392#_c_703_n N_VPWR_c_875_n 0.00539454f $X=5.43 $Y=2.025 $X2=0
+ $Y2=0
cc_522 N_A_639_392#_c_705_n N_VPWR_c_875_n 0.00539454f $X=5.88 $Y=2.025 $X2=0
+ $Y2=0
cc_523 N_A_639_392#_c_695_n N_VGND_c_1060_n 0.00131584f $X=5.535 $Y=1.12 $X2=0
+ $Y2=0
cc_524 N_A_639_392#_c_737_n N_VGND_c_1060_n 0.00834935f $X=3.905 $Y=0.565 $X2=0
+ $Y2=0
cc_525 N_A_639_392#_c_697_n N_VGND_c_1060_n 0.0149311f $X=4.815 $Y=0.935 $X2=0
+ $Y2=0
cc_526 N_A_639_392#_c_699_n N_VGND_c_1060_n 0.00981709f $X=5.017 $Y=1.322 $X2=0
+ $Y2=0
cc_527 N_A_639_392#_c_696_n N_VGND_c_1061_n 2.42234e-19 $X=5.965 $Y=1.12 $X2=0
+ $Y2=0
cc_528 N_A_639_392#_c_737_n N_VGND_c_1067_n 0.0101443f $X=3.905 $Y=0.565 $X2=0
+ $Y2=0
cc_529 N_A_639_392#_c_695_n N_VGND_c_1070_n 0.00278247f $X=5.535 $Y=1.12 $X2=0
+ $Y2=0
cc_530 N_A_639_392#_c_696_n N_VGND_c_1070_n 0.00278247f $X=5.965 $Y=1.12 $X2=0
+ $Y2=0
cc_531 N_A_639_392#_c_695_n N_VGND_c_1079_n 0.00358425f $X=5.535 $Y=1.12 $X2=0
+ $Y2=0
cc_532 N_A_639_392#_c_696_n N_VGND_c_1079_n 0.00353524f $X=5.965 $Y=1.12 $X2=0
+ $Y2=0
cc_533 N_A_639_392#_c_737_n N_VGND_c_1079_n 0.0115712f $X=3.905 $Y=0.565 $X2=0
+ $Y2=0
cc_534 N_A_639_392#_c_697_n N_VGND_c_1079_n 0.0168958f $X=4.815 $Y=0.935 $X2=0
+ $Y2=0
cc_535 N_A_639_392#_c_699_n N_VGND_c_1079_n 0.00277523f $X=5.017 $Y=1.322 $X2=0
+ $Y2=0
cc_536 N_A_639_392#_c_695_n N_A_1035_74#_c_1178_n 0.00781452f $X=5.535 $Y=1.12
+ $X2=0 $Y2=0
cc_537 N_A_639_392#_c_696_n N_A_1035_74#_c_1178_n 6.05606e-19 $X=5.965 $Y=1.12
+ $X2=0 $Y2=0
cc_538 N_A_639_392#_c_699_n N_A_1035_74#_c_1178_n 0.0144827f $X=5.017 $Y=1.322
+ $X2=0 $Y2=0
cc_539 N_A_639_392#_c_701_n N_A_1035_74#_c_1178_n 0.0106502f $X=5.88 $Y=1.455
+ $X2=0 $Y2=0
cc_540 N_A_639_392#_c_695_n N_A_1035_74#_c_1179_n 0.0100245f $X=5.535 $Y=1.12
+ $X2=0 $Y2=0
cc_541 N_A_639_392#_c_696_n N_A_1035_74#_c_1179_n 0.0116238f $X=5.965 $Y=1.12
+ $X2=0 $Y2=0
cc_542 N_A_639_392#_c_701_n N_A_1035_74#_c_1179_n 2.49111e-19 $X=5.88 $Y=1.455
+ $X2=0 $Y2=0
cc_543 N_A_639_392#_c_695_n N_A_1035_74#_c_1180_n 0.00281658f $X=5.535 $Y=1.12
+ $X2=0 $Y2=0
cc_544 N_A_639_392#_c_696_n N_A_1035_74#_c_1187_n 0.00243926f $X=5.965 $Y=1.12
+ $X2=0 $Y2=0
cc_545 N_A_639_392#_c_695_n N_A_1035_74#_c_1198_n 5.52887e-19 $X=5.535 $Y=1.12
+ $X2=0 $Y2=0
cc_546 N_A_639_392#_c_696_n N_A_1035_74#_c_1198_n 0.00474692f $X=5.965 $Y=1.12
+ $X2=0 $Y2=0
cc_547 N_RESET_B_c_820_n N_VPWR_c_878_n 0.0153096f $X=6.38 $Y=2.025 $X2=0 $Y2=0
cc_548 N_RESET_B_c_822_n N_VPWR_c_878_n 6.98753e-19 $X=6.9 $Y=2.025 $X2=0 $Y2=0
cc_549 N_RESET_B_c_822_n N_VPWR_c_879_n 0.0119222f $X=6.9 $Y=2.025 $X2=0 $Y2=0
cc_550 N_RESET_B_c_820_n N_VPWR_c_885_n 0.00505726f $X=6.38 $Y=2.025 $X2=0 $Y2=0
cc_551 N_RESET_B_c_822_n N_VPWR_c_885_n 0.00563421f $X=6.9 $Y=2.025 $X2=0 $Y2=0
cc_552 N_RESET_B_c_820_n N_VPWR_c_875_n 0.00489105f $X=6.38 $Y=2.025 $X2=0 $Y2=0
cc_553 N_RESET_B_c_822_n N_VPWR_c_875_n 0.00539454f $X=6.9 $Y=2.025 $X2=0 $Y2=0
cc_554 N_RESET_B_c_822_n N_Q_c_994_n 5.46196e-19 $X=6.9 $Y=2.025 $X2=0 $Y2=0
cc_555 RESET_B N_Q_c_984_n 4.79428e-19 $X=7.355 $Y=1.21 $X2=0 $Y2=0
cc_556 N_RESET_B_c_814_n N_VGND_c_1061_n 0.00623004f $X=6.395 $Y=1.12 $X2=0
+ $Y2=0
cc_557 N_RESET_B_c_815_n N_VGND_c_1061_n 0.00749966f $X=6.825 $Y=1.12 $X2=0
+ $Y2=0
cc_558 N_RESET_B_c_815_n N_VGND_c_1062_n 0.00383152f $X=6.825 $Y=1.12 $X2=0
+ $Y2=0
cc_559 N_RESET_B_c_815_n N_VGND_c_1063_n 0.00252276f $X=6.825 $Y=1.12 $X2=0
+ $Y2=0
cc_560 RESET_B N_VGND_c_1063_n 0.0103498f $X=7.355 $Y=1.21 $X2=0 $Y2=0
cc_561 N_RESET_B_c_814_n N_VGND_c_1070_n 0.00383152f $X=6.395 $Y=1.12 $X2=0
+ $Y2=0
cc_562 N_RESET_B_c_814_n N_VGND_c_1079_n 0.00369368f $X=6.395 $Y=1.12 $X2=0
+ $Y2=0
cc_563 N_RESET_B_c_815_n N_VGND_c_1079_n 0.00374269f $X=6.825 $Y=1.12 $X2=0
+ $Y2=0
cc_564 N_RESET_B_c_814_n N_A_1035_74#_c_1179_n 9.48753e-19 $X=6.395 $Y=1.12
+ $X2=0 $Y2=0
cc_565 N_RESET_B_c_814_n N_A_1035_74#_c_1201_n 0.00969758f $X=6.395 $Y=1.12
+ $X2=0 $Y2=0
cc_566 N_RESET_B_c_815_n N_A_1035_74#_c_1201_n 0.00969758f $X=6.825 $Y=1.12
+ $X2=0 $Y2=0
cc_567 RESET_B N_A_1035_74#_c_1201_n 0.0397203f $X=7.355 $Y=1.21 $X2=0 $Y2=0
cc_568 N_RESET_B_c_818_n N_A_1035_74#_c_1201_n 0.0024149f $X=6.825 $Y=1.285
+ $X2=0 $Y2=0
cc_569 RESET_B N_A_1035_74#_c_1181_n 0.0216332f $X=7.355 $Y=1.21 $X2=0 $Y2=0
cc_570 N_RESET_B_c_818_n N_A_1035_74#_c_1181_n 0.00118495f $X=6.825 $Y=1.285
+ $X2=0 $Y2=0
cc_571 N_RESET_B_c_815_n N_A_1035_74#_c_1182_n 3.34329e-19 $X=6.825 $Y=1.12
+ $X2=0 $Y2=0
cc_572 N_VPWR_c_879_n N_Q_c_989_n 0.032647f $X=7.21 $Y=2.245 $X2=0 $Y2=0
cc_573 N_VPWR_c_880_n N_Q_c_989_n 0.0263057f $X=8.21 $Y=2.465 $X2=0 $Y2=0
cc_574 N_VPWR_c_887_n N_Q_c_989_n 0.014552f $X=8.045 $Y=3.33 $X2=0 $Y2=0
cc_575 N_VPWR_c_875_n N_Q_c_989_n 0.0119791f $X=9.36 $Y=3.33 $X2=0 $Y2=0
cc_576 N_VPWR_M1014_d N_Q_c_1001_n 0.00528177f $X=8.01 $Y=1.84 $X2=0 $Y2=0
cc_577 N_VPWR_c_880_n N_Q_c_1001_n 0.0202249f $X=8.21 $Y=2.465 $X2=0 $Y2=0
cc_578 N_VPWR_c_880_n N_Q_c_990_n 0.0263057f $X=8.21 $Y=2.465 $X2=0 $Y2=0
cc_579 N_VPWR_c_882_n N_Q_c_990_n 0.0323093f $X=9.21 $Y=2.305 $X2=0 $Y2=0
cc_580 N_VPWR_c_889_n N_Q_c_990_n 0.0146357f $X=9.045 $Y=3.33 $X2=0 $Y2=0
cc_581 N_VPWR_c_875_n N_Q_c_990_n 0.0121141f $X=9.36 $Y=3.33 $X2=0 $Y2=0
cc_582 N_VPWR_M1017_d N_Q_c_991_n 0.00338739f $X=9.06 $Y=1.84 $X2=0 $Y2=0
cc_583 N_VPWR_c_882_n N_Q_c_991_n 0.0230998f $X=9.21 $Y=2.305 $X2=0 $Y2=0
cc_584 N_Q_c_988_n N_VGND_M1005_d 0.00176461f $X=8.795 $Y=0.965 $X2=0 $Y2=0
cc_585 Q N_VGND_M1025_d 0.0042279f $X=9.275 $Y=0.84 $X2=0 $Y2=0
cc_586 N_Q_c_983_n N_VGND_c_1063_n 0.0224826f $X=8.03 $Y=0.525 $X2=0 $Y2=0
cc_587 N_Q_c_983_n N_VGND_c_1064_n 0.016479f $X=8.03 $Y=0.525 $X2=0 $Y2=0
cc_588 N_Q_c_985_n N_VGND_c_1064_n 0.016479f $X=8.89 $Y=0.525 $X2=0 $Y2=0
cc_589 N_Q_c_988_n N_VGND_c_1064_n 0.0170777f $X=8.795 $Y=0.965 $X2=0 $Y2=0
cc_590 N_Q_c_985_n N_VGND_c_1066_n 0.0104754f $X=8.89 $Y=0.525 $X2=0 $Y2=0
cc_591 Q N_VGND_c_1066_n 0.0216656f $X=9.275 $Y=0.84 $X2=0 $Y2=0
cc_592 N_Q_c_983_n N_VGND_c_1071_n 0.00806491f $X=8.03 $Y=0.525 $X2=0 $Y2=0
cc_593 N_Q_c_985_n N_VGND_c_1072_n 0.00781705f $X=8.89 $Y=0.525 $X2=0 $Y2=0
cc_594 N_Q_c_983_n N_VGND_c_1079_n 0.00690154f $X=8.03 $Y=0.525 $X2=0 $Y2=0
cc_595 N_Q_c_985_n N_VGND_c_1079_n 0.00680101f $X=8.89 $Y=0.525 $X2=0 $Y2=0
cc_596 Q N_VGND_c_1079_n 0.00669281f $X=9.275 $Y=0.84 $X2=0 $Y2=0
cc_597 N_VGND_c_1060_n N_A_1035_74#_c_1178_n 0.017158f $X=4.76 $Y=0.515 $X2=0
+ $Y2=0
cc_598 N_VGND_c_1061_n N_A_1035_74#_c_1179_n 0.0112234f $X=6.61 $Y=0.515 $X2=0
+ $Y2=0
cc_599 N_VGND_c_1070_n N_A_1035_74#_c_1179_n 0.0512248f $X=6.445 $Y=0 $X2=0
+ $Y2=0
cc_600 N_VGND_c_1079_n N_A_1035_74#_c_1179_n 0.0283929f $X=9.36 $Y=0 $X2=0 $Y2=0
cc_601 N_VGND_c_1060_n N_A_1035_74#_c_1180_n 0.0121616f $X=4.76 $Y=0.515 $X2=0
+ $Y2=0
cc_602 N_VGND_c_1070_n N_A_1035_74#_c_1180_n 0.0236075f $X=6.445 $Y=0 $X2=0
+ $Y2=0
cc_603 N_VGND_c_1079_n N_A_1035_74#_c_1180_n 0.0127226f $X=9.36 $Y=0 $X2=0 $Y2=0
cc_604 N_VGND_M1002_s N_A_1035_74#_c_1201_n 0.0032758f $X=6.47 $Y=0.37 $X2=0
+ $Y2=0
cc_605 N_VGND_c_1061_n N_A_1035_74#_c_1201_n 0.0166614f $X=6.61 $Y=0.515 $X2=0
+ $Y2=0
cc_606 N_VGND_c_1079_n N_A_1035_74#_c_1201_n 0.0122318f $X=9.36 $Y=0 $X2=0 $Y2=0
cc_607 N_VGND_c_1063_n N_A_1035_74#_c_1181_n 0.012877f $X=7.6 $Y=0.525 $X2=0
+ $Y2=0
cc_608 N_VGND_c_1061_n N_A_1035_74#_c_1182_n 0.00975481f $X=6.61 $Y=0.515 $X2=0
+ $Y2=0
cc_609 N_VGND_c_1062_n N_A_1035_74#_c_1182_n 0.0111768f $X=7.435 $Y=0 $X2=0
+ $Y2=0
cc_610 N_VGND_c_1063_n N_A_1035_74#_c_1182_n 0.0274502f $X=7.6 $Y=0.525 $X2=0
+ $Y2=0
cc_611 N_VGND_c_1079_n N_A_1035_74#_c_1182_n 0.00945682f $X=9.36 $Y=0 $X2=0
+ $Y2=0
