* File: sky130_fd_sc_hs__dlrtp_4.spice
* Created: Thu Aug 27 20:42:03 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hs__dlrtp_4.pex.spice"
.subckt sky130_fd_sc_hs__dlrtp_4  VNB VPB D GATE RESET_B VPWR Q VGND
* 
* VGND	VGND
* Q	Q
* VPWR	VPWR
* RESET_B	RESET_B
* GATE	GATE
* D	D
* VPB	VPB
* VNB	VNB
MM1019 N_VGND_M1019_d N_D_M1019_g N_A_27_126#_M1019_s VNB NLOWVT L=0.15 W=0.55
+ AD=0.165874 AS=0.15675 PD=1.09574 PS=1.67 NRD=29.448 NRS=0 M=1 R=3.66667
+ SA=75000.2 SB=75000.9 A=0.0825 P=1.4 MULT=1
MM1004 N_A_240_394#_M1004_d N_GATE_M1004_g N_VGND_M1019_d VNB NLOWVT L=0.15
+ W=0.74 AD=0.2109 AS=0.223176 PD=2.05 PS=1.47426 NRD=0 NRS=21.072 M=1 R=4.93333
+ SA=75000.8 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1024 N_VGND_M1024_d N_A_240_394#_M1024_g N_A_364_120#_M1024_s VNB NLOWVT
+ L=0.15 W=0.74 AD=0.160253 AS=0.2294 PD=1.43174 PS=2.1 NRD=26.196 NRS=2.424 M=1
+ R=4.93333 SA=75000.2 SB=75001 A=0.111 P=1.78 MULT=1
MM1001 A_559_74# N_A_27_126#_M1001_g N_VGND_M1024_d VNB NLOWVT L=0.15 W=0.64
+ AD=0.0816 AS=0.138597 PD=0.895 PS=1.23826 NRD=13.584 NRS=0.936 M=1 R=4.26667
+ SA=75000.6 SB=75001.3 A=0.096 P=1.58 MULT=1
MM1027 N_A_640_74#_M1027_d N_A_364_120#_M1027_g A_559_74# VNB NLOWVT L=0.15
+ W=0.64 AD=0.154264 AS=0.0816 PD=1.28604 PS=0.895 NRD=5.616 NRS=13.584 M=1
+ R=4.26667 SA=75001 SB=75000.8 A=0.096 P=1.58 MULT=1
MM1002 A_755_74# N_A_240_394#_M1002_g N_A_640_74#_M1027_d VNB NLOWVT L=0.15
+ W=0.42 AD=0.0441 AS=0.101236 PD=0.63 PS=0.843962 NRD=14.28 NRS=34.284 M=1
+ R=2.8 SA=75001.4 SB=75000.6 A=0.063 P=1.14 MULT=1
MM1026 N_VGND_M1026_d N_A_797_48#_M1026_g A_755_74# VNB NLOWVT L=0.15 W=0.42
+ AD=0.1197 AS=0.0441 PD=1.41 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75001.8
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1000 N_A_938_74#_M1000_d N_A_640_74#_M1000_g N_A_797_48#_M1000_s VNB NLOWVT
+ L=0.15 W=0.64 AD=0.1824 AS=0.0912 PD=1.85 PS=0.925 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75001.5 A=0.096 P=1.58 MULT=1
MM1006 N_A_938_74#_M1006_d N_A_640_74#_M1006_g N_A_797_48#_M1000_s VNB NLOWVT
+ L=0.15 W=0.64 AD=0.0896 AS=0.0912 PD=0.92 PS=0.925 NRD=0 NRS=0.936 M=1
+ R=4.26667 SA=75000.6 SB=75001.1 A=0.096 P=1.58 MULT=1
MM1020 N_VGND_M1020_d N_RESET_B_M1020_g N_A_938_74#_M1006_d VNB NLOWVT L=0.15
+ W=0.64 AD=0.0896 AS=0.0896 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75001.1 SB=75000.6 A=0.096 P=1.58 MULT=1
MM1028 N_VGND_M1020_d N_RESET_B_M1028_g N_A_938_74#_M1028_s VNB NLOWVT L=0.15
+ W=0.64 AD=0.0896 AS=0.1824 PD=0.92 PS=1.85 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75001.5 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1011 N_Q_M1011_d N_A_797_48#_M1011_g N_VGND_M1011_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.2109 PD=1.02 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75001.5 A=0.111 P=1.78 MULT=1
MM1015 N_Q_M1011_d N_A_797_48#_M1015_g N_VGND_M1015_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.6
+ SB=75001.1 A=0.111 P=1.78 MULT=1
MM1023 N_Q_M1023_d N_A_797_48#_M1023_g N_VGND_M1015_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.1
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1029 N_Q_M1023_d N_A_797_48#_M1029_g N_VGND_M1029_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.2109 PD=1.02 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.5
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1009 N_VPWR_M1009_d N_D_M1009_g N_A_27_126#_M1009_s VPB PSHORT L=0.15 W=0.84
+ AD=0.22785 AS=0.2478 PD=1.52 PS=2.27 NRD=50.7078 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75000.9 A=0.126 P=1.98 MULT=1
MM1007 N_A_240_394#_M1007_d N_GATE_M1007_g N_VPWR_M1009_d VPB PSHORT L=0.15
+ W=0.84 AD=0.294 AS=0.22785 PD=2.38 PS=1.52 NRD=0 NRS=50.7078 M=1 R=5.6
+ SA=75000.8 SB=75000.3 A=0.126 P=1.98 MULT=1
MM1016 N_VPWR_M1016_d N_A_240_394#_M1016_g N_A_364_120#_M1016_s VPB PSHORT
+ L=0.15 W=0.84 AD=0.173752 AS=0.2478 PD=1.2737 PS=2.27 NRD=23.443 NRS=2.3443
+ M=1 R=5.6 SA=75000.2 SB=75002.3 A=0.126 P=1.98 MULT=1
MM1018 A_562_392# N_A_27_126#_M1018_g N_VPWR_M1016_d VPB PSHORT L=0.15 W=1
+ AD=0.12 AS=0.206848 PD=1.24 PS=1.5163 NRD=12.7853 NRS=3.9203 M=1 R=6.66667
+ SA=75000.7 SB=75001.8 A=0.15 P=2.3 MULT=1
MM1008 N_A_640_74#_M1008_d N_A_240_394#_M1008_g A_562_392# VPB PSHORT L=0.15 W=1
+ AD=0.234366 AS=0.12 PD=1.9507 PS=1.24 NRD=1.9503 NRS=12.7853 M=1 R=6.66667
+ SA=75001.1 SB=75001.4 A=0.15 P=2.3 MULT=1
MM1005 A_747_508# N_A_364_120#_M1005_g N_A_640_74#_M1008_d VPB PSHORT L=0.15
+ W=0.42 AD=0.09975 AS=0.0984338 PD=0.895 PS=0.819296 NRD=85.5965 NRS=46.886 M=1
+ R=2.8 SA=75001.5 SB=75002.4 A=0.063 P=1.14 MULT=1
MM1003 N_VPWR_M1003_d N_A_797_48#_M1003_g A_747_508# VPB PSHORT L=0.15 W=0.42
+ AD=0.139533 AS=0.09975 PD=1.15667 PS=0.895 NRD=58.6272 NRS=85.5965 M=1 R=2.8
+ SA=75002.1 SB=75001.8 A=0.063 P=1.14 MULT=1
MM1017 N_A_797_48#_M1017_d N_A_640_74#_M1017_g N_VPWR_M1003_d VPB PSHORT L=0.15
+ W=0.84 AD=0.126 AS=0.279067 PD=1.14 PS=2.31333 NRD=2.3443 NRS=65.01 M=1 R=5.6
+ SA=75000.7 SB=75003.7 A=0.126 P=1.98 MULT=1
MM1025 N_A_797_48#_M1017_d N_A_640_74#_M1025_g N_VPWR_M1025_s VPB PSHORT L=0.15
+ W=0.84 AD=0.126 AS=0.147 PD=1.14 PS=1.19 NRD=2.3443 NRS=14.0658 M=1 R=5.6
+ SA=75001.1 SB=75003.3 A=0.126 P=1.98 MULT=1
MM1021 N_A_797_48#_M1021_d N_RESET_B_M1021_g N_VPWR_M1025_s VPB PSHORT L=0.15
+ W=0.84 AD=0.147 AS=0.147 PD=1.19 PS=1.19 NRD=14.0658 NRS=2.3443 M=1 R=5.6
+ SA=75001.6 SB=75002.8 A=0.126 P=1.98 MULT=1
MM1022 N_A_797_48#_M1021_d N_RESET_B_M1022_g N_VPWR_M1022_s VPB PSHORT L=0.15
+ W=0.84 AD=0.147 AS=0.174 PD=1.19 PS=1.29 NRD=2.3443 NRS=22.261 M=1 R=5.6
+ SA=75002.1 SB=75002.3 A=0.126 P=1.98 MULT=1
MM1010 N_Q_M1010_d N_A_797_48#_M1010_g N_VPWR_M1022_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.232 PD=1.42 PS=1.72 NRD=1.7533 NRS=1.7533 M=1 R=7.46667 SA=75002
+ SB=75001.7 A=0.168 P=2.54 MULT=1
MM1012 N_Q_M1010_d N_A_797_48#_M1012_g N_VPWR_M1012_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.196 PD=1.42 PS=1.47 NRD=1.7533 NRS=10.5395 M=1 R=7.46667
+ SA=75002.5 SB=75001.3 A=0.168 P=2.54 MULT=1
MM1013 N_Q_M1013_d N_A_797_48#_M1013_g N_VPWR_M1012_s VPB PSHORT L=0.15 W=1.12
+ AD=0.2072 AS=0.196 PD=1.49 PS=1.47 NRD=10.5395 NRS=1.7533 M=1 R=7.46667
+ SA=75003 SB=75000.8 A=0.168 P=2.54 MULT=1
MM1014 N_Q_M1013_d N_A_797_48#_M1014_g N_VPWR_M1014_s VPB PSHORT L=0.15 W=1.12
+ AD=0.2072 AS=0.364 PD=1.49 PS=2.89 NRD=5.2599 NRS=7.0329 M=1 R=7.46667
+ SA=75003.5 SB=75000.2 A=0.168 P=2.54 MULT=1
DX30_noxref VNB VPB NWDIODE A=17.5032 P=22.96
c_1266 A_559_74# 0 5.47968e-20 $X=2.795 $Y=0.37
*
.include "sky130_fd_sc_hs__dlrtp_4.pxi.spice"
*
.ends
*
*
