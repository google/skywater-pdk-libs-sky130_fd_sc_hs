* File: sky130_fd_sc_hs__nor4_2.pxi.spice
* Created: Thu Aug 27 20:54:48 2020
* 
x_PM_SKY130_FD_SC_HS__NOR4_2%C N_C_c_78_n N_C_c_87_n N_C_M1002_g N_C_c_79_n
+ N_C_M1008_g N_C_M1007_g N_C_c_81_n N_C_c_82_n C C N_C_c_83_n C N_C_c_85_n
+ PM_SKY130_FD_SC_HS__NOR4_2%C
x_PM_SKY130_FD_SC_HS__NOR4_2%D N_D_c_150_n N_D_c_157_n N_D_M1000_g N_D_c_151_n
+ N_D_c_152_n N_D_c_153_n N_D_c_160_n N_D_M1010_g N_D_c_154_n N_D_M1009_g D
+ N_D_c_156_n PM_SKY130_FD_SC_HS__NOR4_2%D
x_PM_SKY130_FD_SC_HS__NOR4_2%B N_B_c_211_n N_B_M1001_g N_B_M1011_g N_B_c_213_n
+ N_B_M1006_g N_B_c_219_n N_B_c_214_n B B B B N_B_c_215_n N_B_c_216_n
+ N_B_c_222_n B PM_SKY130_FD_SC_HS__NOR4_2%B
x_PM_SKY130_FD_SC_HS__NOR4_2%A N_A_c_288_n N_A_M1003_g N_A_c_285_n N_A_M1005_g
+ N_A_c_289_n N_A_M1004_g A N_A_c_287_n PM_SKY130_FD_SC_HS__NOR4_2%A
x_PM_SKY130_FD_SC_HS__NOR4_2%A_27_368# N_A_27_368#_M1002_d N_A_27_368#_M1008_d
+ N_A_27_368#_M1006_s N_A_27_368#_c_328_n N_A_27_368#_c_335_n
+ N_A_27_368#_c_329_n N_A_27_368#_c_348_n N_A_27_368#_c_330_n
+ N_A_27_368#_c_331_n N_A_27_368#_c_332_n N_A_27_368#_c_333_n
+ PM_SKY130_FD_SC_HS__NOR4_2%A_27_368#
x_PM_SKY130_FD_SC_HS__NOR4_2%A_116_368# N_A_116_368#_M1002_s
+ N_A_116_368#_M1010_d N_A_116_368#_c_387_n
+ PM_SKY130_FD_SC_HS__NOR4_2%A_116_368#
x_PM_SKY130_FD_SC_HS__NOR4_2%Y N_Y_M1009_d N_Y_M1011_d N_Y_M1000_s N_Y_c_402_n
+ N_Y_c_403_n N_Y_c_404_n N_Y_c_410_n N_Y_c_405_n N_Y_c_406_n N_Y_c_407_n
+ N_Y_c_408_n Y Y N_Y_c_412_n PM_SKY130_FD_SC_HS__NOR4_2%Y
x_PM_SKY130_FD_SC_HS__NOR4_2%A_490_368# N_A_490_368#_M1001_d
+ N_A_490_368#_M1004_s N_A_490_368#_c_488_n N_A_490_368#_c_485_n
+ N_A_490_368#_c_480_n N_A_490_368#_c_481_n
+ PM_SKY130_FD_SC_HS__NOR4_2%A_490_368#
x_PM_SKY130_FD_SC_HS__NOR4_2%VPWR N_VPWR_M1003_d N_VPWR_c_509_n VPWR
+ N_VPWR_c_510_n N_VPWR_c_511_n N_VPWR_c_508_n N_VPWR_c_513_n
+ PM_SKY130_FD_SC_HS__NOR4_2%VPWR
x_PM_SKY130_FD_SC_HS__NOR4_2%VGND N_VGND_M1009_s N_VGND_M1007_d N_VGND_M1005_d
+ N_VGND_c_555_n N_VGND_c_556_n N_VGND_c_557_n VGND N_VGND_c_558_n
+ N_VGND_c_559_n N_VGND_c_560_n N_VGND_c_561_n N_VGND_c_562_n N_VGND_c_563_n
+ N_VGND_c_564_n PM_SKY130_FD_SC_HS__NOR4_2%VGND
cc_1 VNB N_C_c_78_n 0.00985164f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.675
cc_2 VNB N_C_c_79_n 0.0277198f $X=-0.19 $Y=-0.245 $X2=1.895 $Y2=1.765
cc_3 VNB N_C_M1007_g 0.0248615f $X=-0.19 $Y=-0.245 $X2=1.93 $Y2=0.74
cc_4 VNB N_C_c_81_n 0.00272143f $X=-0.19 $Y=-0.245 $X2=0.535 $Y2=1.335
cc_5 VNB N_C_c_82_n 0.0323937f $X=-0.19 $Y=-0.245 $X2=0.535 $Y2=1.335
cc_6 VNB N_C_c_83_n 0.00590745f $X=-0.19 $Y=-0.245 $X2=1.91 $Y2=1.485
cc_7 VNB C 6.99497e-19 $X=-0.19 $Y=-0.245 $X2=1.68 $Y2=1.665
cc_8 VNB N_C_c_85_n 0.00494578f $X=-0.19 $Y=-0.245 $X2=1.565 $Y2=1.485
cc_9 VNB N_D_c_150_n 0.0378968f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.5
cc_10 VNB N_D_c_151_n 0.018773f $X=-0.19 $Y=-0.245 $X2=1.895 $Y2=2.4
cc_11 VNB N_D_c_152_n 0.0465632f $X=-0.19 $Y=-0.245 $X2=1.895 $Y2=2.4
cc_12 VNB N_D_c_153_n 0.00743291f $X=-0.19 $Y=-0.245 $X2=1.93 $Y2=1.32
cc_13 VNB N_D_c_154_n 0.016723f $X=-0.19 $Y=-0.245 $X2=1.565 $Y2=1.41
cc_14 VNB D 0.00434149f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_D_c_156_n 0.0732973f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_B_c_211_n 0.0282287f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.5
cc_17 VNB N_B_M1011_g 0.024237f $X=-0.19 $Y=-0.245 $X2=1.895 $Y2=1.765
cc_18 VNB N_B_c_213_n 0.0412845f $X=-0.19 $Y=-0.245 $X2=1.895 $Y2=2.4
cc_19 VNB N_B_c_214_n 0.00715627f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=1.41
cc_20 VNB N_B_c_215_n 0.163114f $X=-0.19 $Y=-0.245 $X2=0.535 $Y2=1.5
cc_21 VNB N_B_c_216_n 0.00361276f $X=-0.19 $Y=-0.245 $X2=1.91 $Y2=1.485
cc_22 VNB N_A_c_285_n 0.0200555f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_23 VNB A 0.021158f $X=-0.19 $Y=-0.245 $X2=1.93 $Y2=0.74
cc_24 VNB N_A_c_287_n 0.0609299f $X=-0.19 $Y=-0.245 $X2=0.562 $Y2=1.335
cc_25 VNB N_Y_c_402_n 0.0320702f $X=-0.19 $Y=-0.245 $X2=1.93 $Y2=0.74
cc_26 VNB N_Y_c_403_n 0.00804079f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_Y_c_404_n 0.00833338f $X=-0.19 $Y=-0.245 $X2=1.565 $Y2=1.41
cc_28 VNB N_Y_c_405_n 0.00280855f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_Y_c_406_n 0.00861013f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_Y_c_407_n 0.00240191f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_Y_c_408_n 0.00287885f $X=-0.19 $Y=-0.245 $X2=0.535 $Y2=1.335
cc_32 VNB N_VPWR_c_508_n 0.183584f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=1.58
cc_33 VNB N_VGND_c_555_n 0.00830622f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_556_n 0.0186948f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=1.41
cc_35 VNB N_VGND_c_557_n 0.017069f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_558_n 0.0186436f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_559_n 0.0291174f $X=-0.19 $Y=-0.245 $X2=1.68 $Y2=1.665
cc_38 VNB N_VGND_c_560_n 0.262723f $X=-0.19 $Y=-0.245 $X2=1.68 $Y2=1.7
cc_39 VNB N_VGND_c_561_n 0.0187181f $X=-0.19 $Y=-0.245 $X2=1.565 $Y2=1.485
cc_40 VNB N_VGND_c_562_n 0.0328803f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_563_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_564_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VPB N_C_c_78_n 7.07408e-19 $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.675
cc_44 VPB N_C_c_87_n 0.0254235f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.765
cc_45 VPB N_C_c_79_n 0.0235277f $X=-0.19 $Y=1.66 $X2=1.895 $Y2=1.765
cc_46 VPB C 0.00282206f $X=-0.19 $Y=1.66 $X2=1.68 $Y2=1.665
cc_47 VPB N_D_c_157_n 0.015395f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.765
cc_48 VPB N_D_c_152_n 0.00583775f $X=-0.19 $Y=1.66 $X2=1.895 $Y2=2.4
cc_49 VPB N_D_c_153_n 7.26044e-19 $X=-0.19 $Y=1.66 $X2=1.93 $Y2=1.32
cc_50 VPB N_D_c_160_n 0.0212918f $X=-0.19 $Y=1.66 $X2=1.93 $Y2=0.74
cc_51 VPB N_B_c_211_n 0.0238131f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.5
cc_52 VPB N_B_c_213_n 0.0268083f $X=-0.19 $Y=1.66 $X2=1.895 $Y2=2.4
cc_53 VPB N_B_c_219_n 0.0102383f $X=-0.19 $Y=1.66 $X2=1.93 $Y2=0.74
cc_54 VPB N_B_c_214_n 0.00113649f $X=-0.19 $Y=1.66 $X2=0.7 $Y2=1.41
cc_55 VPB N_B_c_216_n 0.00182616f $X=-0.19 $Y=1.66 $X2=1.91 $Y2=1.485
cc_56 VPB N_B_c_222_n 0.00766629f $X=-0.19 $Y=1.66 $X2=1.68 $Y2=1.7
cc_57 VPB N_A_c_288_n 0.0152808f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.5
cc_58 VPB N_A_c_289_n 0.0146527f $X=-0.19 $Y=1.66 $X2=1.895 $Y2=2.4
cc_59 VPB N_A_c_287_n 0.0124458f $X=-0.19 $Y=1.66 $X2=0.562 $Y2=1.335
cc_60 VPB N_A_27_368#_c_328_n 0.0214044f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_61 VPB N_A_27_368#_c_329_n 0.00253974f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_62 VPB N_A_27_368#_c_330_n 0.00718969f $X=-0.19 $Y=1.66 $X2=1.595 $Y2=1.95
cc_63 VPB N_A_27_368#_c_331_n 0.0306198f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_64 VPB N_A_27_368#_c_332_n 0.0184043f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_65 VPB N_A_27_368#_c_333_n 0.00419538f $X=-0.19 $Y=1.66 $X2=1.68 $Y2=1.65
cc_66 VPB N_A_116_368#_c_387_n 0.00796531f $X=-0.19 $Y=1.66 $X2=1.93 $Y2=0.74
cc_67 VPB N_Y_c_402_n 4.44592e-19 $X=-0.19 $Y=1.66 $X2=1.93 $Y2=0.74
cc_68 VPB N_Y_c_410_n 0.00926672f $X=-0.19 $Y=1.66 $X2=0.562 $Y2=1.335
cc_69 VPB Y 0.0045771f $X=-0.19 $Y=1.66 $X2=1.68 $Y2=1.65
cc_70 VPB N_Y_c_412_n 0.00432877f $X=-0.19 $Y=1.66 $X2=1.68 $Y2=2.035
cc_71 VPB N_A_490_368#_c_480_n 0.00226153f $X=-0.19 $Y=1.66 $X2=1.565 $Y2=1.41
cc_72 VPB N_A_490_368#_c_481_n 0.00371798f $X=-0.19 $Y=1.66 $X2=0.535 $Y2=1.335
cc_73 VPB N_VPWR_c_509_n 0.00396467f $X=-0.19 $Y=1.66 $X2=1.895 $Y2=1.765
cc_74 VPB N_VPWR_c_510_n 0.0801372f $X=-0.19 $Y=1.66 $X2=1.93 $Y2=0.74
cc_75 VPB N_VPWR_c_511_n 0.0302153f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_76 VPB N_VPWR_c_508_n 0.0690666f $X=-0.19 $Y=1.66 $X2=1.595 $Y2=1.58
cc_77 VPB N_VPWR_c_513_n 0.00601668f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_78 N_C_c_85_n N_D_c_150_n 0.00105479f $X=1.565 $Y=1.485 $X2=-0.19 $Y2=-0.245
cc_79 N_C_c_87_n N_D_c_157_n 0.0358376f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_80 N_C_c_81_n N_D_c_151_n 0.00113177f $X=0.535 $Y=1.335 $X2=0 $Y2=0
cc_81 N_C_c_82_n N_D_c_151_n 0.0222163f $X=0.535 $Y=1.335 $X2=0 $Y2=0
cc_82 N_C_c_78_n N_D_c_152_n 0.011803f $X=0.505 $Y=1.675 $X2=0 $Y2=0
cc_83 N_C_c_79_n N_D_c_152_n 0.0207003f $X=1.895 $Y=1.765 $X2=0 $Y2=0
cc_84 N_C_c_83_n N_D_c_152_n 0.00443665f $X=1.91 $Y=1.485 $X2=0 $Y2=0
cc_85 N_C_c_85_n N_D_c_152_n 0.0377601f $X=1.565 $Y=1.485 $X2=0 $Y2=0
cc_86 N_C_c_79_n N_D_c_153_n 0.0043173f $X=1.895 $Y=1.765 $X2=0 $Y2=0
cc_87 C N_D_c_153_n 0.00127487f $X=1.68 $Y=1.665 $X2=0 $Y2=0
cc_88 N_C_c_79_n N_D_c_160_n 0.0366793f $X=1.895 $Y=1.765 $X2=0 $Y2=0
cc_89 C N_D_c_160_n 0.00198883f $X=1.68 $Y=1.665 $X2=0 $Y2=0
cc_90 N_C_M1007_g N_D_c_154_n 0.0162664f $X=1.93 $Y=0.74 $X2=0 $Y2=0
cc_91 N_C_c_81_n N_D_c_156_n 2.88011e-19 $X=0.535 $Y=1.335 $X2=0 $Y2=0
cc_92 N_C_c_82_n N_D_c_156_n 0.0145077f $X=0.535 $Y=1.335 $X2=0 $Y2=0
cc_93 N_C_c_79_n N_B_c_211_n 0.0350736f $X=1.895 $Y=1.765 $X2=-0.19 $Y2=-0.245
cc_94 N_C_c_83_n N_B_c_211_n 4.11724e-19 $X=1.91 $Y=1.485 $X2=-0.19 $Y2=-0.245
cc_95 N_C_M1007_g N_B_M1011_g 0.0254515f $X=1.93 $Y=0.74 $X2=0 $Y2=0
cc_96 N_C_c_79_n N_B_c_214_n 7.53308e-19 $X=1.895 $Y=1.765 $X2=0 $Y2=0
cc_97 N_C_c_83_n N_B_c_214_n 0.0220044f $X=1.91 $Y=1.485 $X2=0 $Y2=0
cc_98 C N_B_c_214_n 0.00491955f $X=1.68 $Y=1.665 $X2=0 $Y2=0
cc_99 N_C_c_87_n N_A_27_368#_c_328_n 0.00590753f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_100 N_C_c_87_n N_A_27_368#_c_335_n 0.0110696f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_101 N_C_c_79_n N_A_27_368#_c_335_n 0.0128124f $X=1.895 $Y=1.765 $X2=0 $Y2=0
cc_102 N_C_c_83_n N_A_27_368#_c_335_n 0.00459743f $X=1.91 $Y=1.485 $X2=0 $Y2=0
cc_103 C N_A_27_368#_c_335_n 0.0147605f $X=1.68 $Y=1.665 $X2=0 $Y2=0
cc_104 N_C_c_87_n N_A_27_368#_c_332_n 0.00565664f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_105 N_C_c_79_n N_A_27_368#_c_333_n 0.0110562f $X=1.895 $Y=1.765 $X2=0 $Y2=0
cc_106 N_C_c_83_n N_A_27_368#_c_333_n 0.003289f $X=1.91 $Y=1.485 $X2=0 $Y2=0
cc_107 C N_A_27_368#_c_333_n 0.0104608f $X=1.68 $Y=1.665 $X2=0 $Y2=0
cc_108 C N_A_116_368#_M1010_d 0.00514296f $X=1.68 $Y=1.665 $X2=0 $Y2=0
cc_109 N_C_c_87_n N_A_116_368#_c_387_n 0.00428008f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_110 N_C_c_79_n N_A_116_368#_c_387_n 0.00382887f $X=1.895 $Y=1.765 $X2=0 $Y2=0
cc_111 N_C_c_78_n N_Y_c_402_n 0.0059715f $X=0.505 $Y=1.675 $X2=0 $Y2=0
cc_112 N_C_c_81_n N_Y_c_402_n 0.0244588f $X=0.535 $Y=1.335 $X2=0 $Y2=0
cc_113 N_C_c_82_n N_Y_c_402_n 0.00789454f $X=0.535 $Y=1.335 $X2=0 $Y2=0
cc_114 N_C_c_81_n N_Y_c_403_n 0.0206189f $X=0.535 $Y=1.335 $X2=0 $Y2=0
cc_115 N_C_c_82_n N_Y_c_403_n 0.0014919f $X=0.535 $Y=1.335 $X2=0 $Y2=0
cc_116 N_C_c_85_n N_Y_c_403_n 0.0358256f $X=1.565 $Y=1.485 $X2=0 $Y2=0
cc_117 N_C_M1007_g N_Y_c_405_n 0.00627366f $X=1.93 $Y=0.74 $X2=0 $Y2=0
cc_118 N_C_c_79_n N_Y_c_406_n 0.00156944f $X=1.895 $Y=1.765 $X2=0 $Y2=0
cc_119 N_C_M1007_g N_Y_c_406_n 0.0123739f $X=1.93 $Y=0.74 $X2=0 $Y2=0
cc_120 N_C_c_83_n N_Y_c_406_n 0.0141875f $X=1.91 $Y=1.485 $X2=0 $Y2=0
cc_121 N_C_M1007_g N_Y_c_407_n 6.22903e-19 $X=1.93 $Y=0.74 $X2=0 $Y2=0
cc_122 N_C_c_79_n N_Y_c_408_n 0.00272201f $X=1.895 $Y=1.765 $X2=0 $Y2=0
cc_123 N_C_M1007_g N_Y_c_408_n 0.00473451f $X=1.93 $Y=0.74 $X2=0 $Y2=0
cc_124 N_C_c_85_n N_Y_c_408_n 0.0282645f $X=1.565 $Y=1.485 $X2=0 $Y2=0
cc_125 C Y 0.0255283f $X=1.68 $Y=1.665 $X2=0 $Y2=0
cc_126 N_C_c_85_n Y 0.0534858f $X=1.565 $Y=1.485 $X2=0 $Y2=0
cc_127 N_C_c_78_n N_Y_c_412_n 0.00264218f $X=0.505 $Y=1.675 $X2=0 $Y2=0
cc_128 N_C_c_87_n N_Y_c_412_n 0.0118614f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_129 N_C_c_81_n N_Y_c_412_n 0.0204894f $X=0.535 $Y=1.335 $X2=0 $Y2=0
cc_130 N_C_c_82_n N_Y_c_412_n 0.00201086f $X=0.535 $Y=1.335 $X2=0 $Y2=0
cc_131 N_C_c_87_n N_VPWR_c_510_n 0.00444483f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_132 N_C_c_79_n N_VPWR_c_510_n 0.00444483f $X=1.895 $Y=1.765 $X2=0 $Y2=0
cc_133 N_C_c_87_n N_VPWR_c_508_n 0.00456474f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_134 N_C_c_79_n N_VPWR_c_508_n 0.00454867f $X=1.895 $Y=1.765 $X2=0 $Y2=0
cc_135 N_C_M1007_g N_VGND_c_555_n 0.00466065f $X=1.93 $Y=0.74 $X2=0 $Y2=0
cc_136 N_C_M1007_g N_VGND_c_558_n 0.00434272f $X=1.93 $Y=0.74 $X2=0 $Y2=0
cc_137 N_C_M1007_g N_VGND_c_560_n 0.0082177f $X=1.93 $Y=0.74 $X2=0 $Y2=0
cc_138 N_D_c_157_n N_A_27_368#_c_335_n 0.0108997f $X=0.97 $Y=1.765 $X2=0 $Y2=0
cc_139 N_D_c_160_n N_A_27_368#_c_335_n 0.01494f $X=1.445 $Y=1.765 $X2=0 $Y2=0
cc_140 N_D_c_157_n N_A_27_368#_c_332_n 9.84326e-19 $X=0.97 $Y=1.765 $X2=0 $Y2=0
cc_141 N_D_c_157_n N_A_116_368#_c_387_n 0.0128409f $X=0.97 $Y=1.765 $X2=0 $Y2=0
cc_142 N_D_c_160_n N_A_116_368#_c_387_n 0.0125604f $X=1.445 $Y=1.765 $X2=0 $Y2=0
cc_143 N_D_c_151_n N_Y_c_402_n 0.00351765f $X=0.985 $Y=1.185 $X2=0 $Y2=0
cc_144 N_D_c_150_n N_Y_c_403_n 0.0167197f $X=0.91 $Y=0.81 $X2=0 $Y2=0
cc_145 N_D_c_151_n N_Y_c_403_n 0.00870161f $X=0.985 $Y=1.185 $X2=0 $Y2=0
cc_146 N_D_c_152_n N_Y_c_403_n 0.00355636f $X=1.445 $Y=1.52 $X2=0 $Y2=0
cc_147 N_D_c_154_n N_Y_c_403_n 0.0109092f $X=1.46 $Y=1.185 $X2=0 $Y2=0
cc_148 D N_Y_c_403_n 0.012611f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_149 N_D_c_156_n N_Y_c_403_n 0.00582959f $X=0.27 $Y=0.495 $X2=0 $Y2=0
cc_150 D N_Y_c_404_n 0.0122776f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_151 N_D_c_156_n N_Y_c_404_n 0.0011793f $X=0.27 $Y=0.495 $X2=0 $Y2=0
cc_152 N_D_c_154_n N_Y_c_405_n 4.77705e-19 $X=1.46 $Y=1.185 $X2=0 $Y2=0
cc_153 N_D_c_154_n N_Y_c_408_n 0.00113886f $X=1.46 $Y=1.185 $X2=0 $Y2=0
cc_154 N_D_c_157_n Y 0.0127973f $X=0.97 $Y=1.765 $X2=0 $Y2=0
cc_155 N_D_c_152_n Y 0.00958467f $X=1.445 $Y=1.52 $X2=0 $Y2=0
cc_156 N_D_c_153_n Y 4.29608e-19 $X=1.445 $Y=1.675 $X2=0 $Y2=0
cc_157 N_D_c_160_n Y 0.0074019f $X=1.445 $Y=1.765 $X2=0 $Y2=0
cc_158 N_D_c_157_n N_VPWR_c_510_n 0.00291649f $X=0.97 $Y=1.765 $X2=0 $Y2=0
cc_159 N_D_c_160_n N_VPWR_c_510_n 0.00291649f $X=1.445 $Y=1.765 $X2=0 $Y2=0
cc_160 N_D_c_157_n N_VPWR_c_508_n 0.00359968f $X=0.97 $Y=1.765 $X2=0 $Y2=0
cc_161 N_D_c_160_n N_VPWR_c_508_n 0.00359835f $X=1.445 $Y=1.765 $X2=0 $Y2=0
cc_162 N_D_c_154_n N_VGND_c_558_n 0.00461464f $X=1.46 $Y=1.185 $X2=0 $Y2=0
cc_163 N_D_c_150_n N_VGND_c_560_n 0.00367388f $X=0.91 $Y=0.81 $X2=0 $Y2=0
cc_164 N_D_c_154_n N_VGND_c_560_n 0.00465425f $X=1.46 $Y=1.185 $X2=0 $Y2=0
cc_165 D N_VGND_c_560_n 0.0117407f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_166 N_D_c_150_n N_VGND_c_561_n 0.00272934f $X=0.91 $Y=0.81 $X2=0 $Y2=0
cc_167 D N_VGND_c_561_n 0.01419f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_168 N_D_c_156_n N_VGND_c_561_n 0.0019148f $X=0.27 $Y=0.495 $X2=0 $Y2=0
cc_169 N_D_c_150_n N_VGND_c_562_n 0.011043f $X=0.91 $Y=0.81 $X2=0 $Y2=0
cc_170 N_D_c_154_n N_VGND_c_562_n 0.00417838f $X=1.46 $Y=1.185 $X2=0 $Y2=0
cc_171 D N_VGND_c_562_n 0.0226857f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_172 N_D_c_156_n N_VGND_c_562_n 0.00626653f $X=0.27 $Y=0.495 $X2=0 $Y2=0
cc_173 N_B_c_211_n N_A_c_288_n 0.0276744f $X=2.375 $Y=1.765 $X2=-0.19 $Y2=-0.245
cc_174 N_B_c_219_n N_A_c_288_n 0.00665343f $X=3.885 $Y=1.795 $X2=-0.19
+ $Y2=-0.245
cc_175 N_B_M1011_g N_A_c_285_n 0.013405f $X=2.5 $Y=0.74 $X2=0 $Y2=0
cc_176 N_B_c_215_n N_A_c_285_n 0.00834965f $X=4.05 $Y=0.445 $X2=0 $Y2=0
cc_177 N_B_c_213_n N_A_c_289_n 0.0277412f $X=3.815 $Y=1.765 $X2=0 $Y2=0
cc_178 N_B_c_219_n N_A_c_289_n 0.00647572f $X=3.885 $Y=1.795 $X2=0 $Y2=0
cc_179 N_B_M1011_g A 3.75378e-19 $X=2.5 $Y=0.74 $X2=0 $Y2=0
cc_180 N_B_c_219_n A 0.0473225f $X=3.885 $Y=1.795 $X2=0 $Y2=0
cc_181 N_B_c_214_n A 0.00850511f $X=2.45 $Y=1.485 $X2=0 $Y2=0
cc_182 N_B_c_215_n A 0.00384508f $X=4.05 $Y=0.445 $X2=0 $Y2=0
cc_183 N_B_c_216_n A 0.0299183f $X=4.05 $Y=0.445 $X2=0 $Y2=0
cc_184 N_B_c_211_n N_A_c_287_n 0.0247101f $X=2.375 $Y=1.765 $X2=0 $Y2=0
cc_185 N_B_M1011_g N_A_c_287_n 0.00591688f $X=2.5 $Y=0.74 $X2=0 $Y2=0
cc_186 N_B_c_219_n N_A_c_287_n 0.0168603f $X=3.885 $Y=1.795 $X2=0 $Y2=0
cc_187 N_B_c_214_n N_A_c_287_n 0.00578243f $X=2.45 $Y=1.485 $X2=0 $Y2=0
cc_188 N_B_c_215_n N_A_c_287_n 0.026038f $X=4.05 $Y=0.445 $X2=0 $Y2=0
cc_189 N_B_c_216_n N_A_c_287_n 0.0010144f $X=4.05 $Y=0.445 $X2=0 $Y2=0
cc_190 N_B_c_222_n N_A_27_368#_M1006_s 0.00285517f $X=4.05 $Y=1.71 $X2=0 $Y2=0
cc_191 N_B_c_211_n N_A_27_368#_c_329_n 3.06945e-19 $X=2.375 $Y=1.765 $X2=0 $Y2=0
cc_192 N_B_c_211_n N_A_27_368#_c_348_n 0.0154029f $X=2.375 $Y=1.765 $X2=0 $Y2=0
cc_193 N_B_c_213_n N_A_27_368#_c_348_n 0.0125489f $X=3.815 $Y=1.765 $X2=0 $Y2=0
cc_194 N_B_c_219_n N_A_27_368#_c_348_n 0.0685877f $X=3.885 $Y=1.795 $X2=0 $Y2=0
cc_195 N_B_c_214_n N_A_27_368#_c_348_n 0.0152005f $X=2.45 $Y=1.485 $X2=0 $Y2=0
cc_196 N_B_c_222_n N_A_27_368#_c_348_n 3.46825e-19 $X=4.05 $Y=1.71 $X2=0 $Y2=0
cc_197 N_B_c_213_n N_A_27_368#_c_330_n 0.00117538f $X=3.815 $Y=1.765 $X2=0 $Y2=0
cc_198 N_B_c_222_n N_A_27_368#_c_330_n 0.0233324f $X=4.05 $Y=1.71 $X2=0 $Y2=0
cc_199 N_B_c_213_n N_A_27_368#_c_331_n 0.00603468f $X=3.815 $Y=1.765 $X2=0 $Y2=0
cc_200 N_B_c_214_n N_A_27_368#_c_333_n 0.00164686f $X=2.45 $Y=1.485 $X2=0 $Y2=0
cc_201 N_B_M1011_g N_Y_c_405_n 6.27466e-19 $X=2.5 $Y=0.74 $X2=0 $Y2=0
cc_202 N_B_c_211_n N_Y_c_406_n 0.0012912f $X=2.375 $Y=1.765 $X2=0 $Y2=0
cc_203 N_B_M1011_g N_Y_c_406_n 0.0129975f $X=2.5 $Y=0.74 $X2=0 $Y2=0
cc_204 N_B_c_219_n N_Y_c_406_n 0.00904733f $X=3.885 $Y=1.795 $X2=0 $Y2=0
cc_205 N_B_c_214_n N_Y_c_406_n 0.0263393f $X=2.45 $Y=1.485 $X2=0 $Y2=0
cc_206 N_B_M1011_g N_Y_c_407_n 0.00935132f $X=2.5 $Y=0.74 $X2=0 $Y2=0
cc_207 N_B_c_219_n N_A_490_368#_M1001_d 0.00167301f $X=3.885 $Y=1.795 $X2=-0.19
+ $Y2=-0.245
cc_208 N_B_c_214_n N_A_490_368#_M1001_d 0.0013013f $X=2.45 $Y=1.485 $X2=-0.19
+ $Y2=-0.245
cc_209 N_B_c_219_n N_A_490_368#_M1004_s 0.00198204f $X=3.885 $Y=1.795 $X2=0
+ $Y2=0
cc_210 N_B_c_213_n N_A_490_368#_c_485_n 0.00195471f $X=3.815 $Y=1.765 $X2=0
+ $Y2=0
cc_211 N_B_c_213_n N_A_490_368#_c_480_n 0.0056682f $X=3.815 $Y=1.765 $X2=0 $Y2=0
cc_212 N_B_c_211_n N_A_490_368#_c_481_n 7.83888e-19 $X=2.375 $Y=1.765 $X2=0
+ $Y2=0
cc_213 N_B_c_219_n N_VPWR_M1003_d 0.00198204f $X=3.885 $Y=1.795 $X2=-0.19
+ $Y2=-0.245
cc_214 N_B_c_211_n N_VPWR_c_509_n 4.76237e-19 $X=2.375 $Y=1.765 $X2=0 $Y2=0
cc_215 N_B_c_213_n N_VPWR_c_509_n 5.40305e-19 $X=3.815 $Y=1.765 $X2=0 $Y2=0
cc_216 N_B_c_211_n N_VPWR_c_510_n 0.00461464f $X=2.375 $Y=1.765 $X2=0 $Y2=0
cc_217 N_B_c_213_n N_VPWR_c_511_n 0.00445347f $X=3.815 $Y=1.765 $X2=0 $Y2=0
cc_218 N_B_c_211_n N_VPWR_c_508_n 0.00910891f $X=2.375 $Y=1.765 $X2=0 $Y2=0
cc_219 N_B_c_213_n N_VPWR_c_508_n 0.00861751f $X=3.815 $Y=1.765 $X2=0 $Y2=0
cc_220 N_B_M1011_g N_VGND_c_555_n 0.00466189f $X=2.5 $Y=0.74 $X2=0 $Y2=0
cc_221 N_B_M1011_g N_VGND_c_556_n 0.00434272f $X=2.5 $Y=0.74 $X2=0 $Y2=0
cc_222 N_B_c_215_n N_VGND_c_557_n 0.00867528f $X=4.05 $Y=0.445 $X2=0 $Y2=0
cc_223 N_B_c_216_n N_VGND_c_557_n 0.0255316f $X=4.05 $Y=0.445 $X2=0 $Y2=0
cc_224 N_B_c_215_n N_VGND_c_559_n 0.00793088f $X=4.05 $Y=0.445 $X2=0 $Y2=0
cc_225 N_B_c_216_n N_VGND_c_559_n 0.0191905f $X=4.05 $Y=0.445 $X2=0 $Y2=0
cc_226 N_B_M1011_g N_VGND_c_560_n 0.0082141f $X=2.5 $Y=0.74 $X2=0 $Y2=0
cc_227 N_B_c_215_n N_VGND_c_560_n 0.00575727f $X=4.05 $Y=0.445 $X2=0 $Y2=0
cc_228 N_B_c_216_n N_VGND_c_560_n 0.012382f $X=4.05 $Y=0.445 $X2=0 $Y2=0
cc_229 N_A_c_288_n N_A_27_368#_c_348_n 0.0111326f $X=2.915 $Y=1.765 $X2=0 $Y2=0
cc_230 N_A_c_289_n N_A_27_368#_c_348_n 0.0106815f $X=3.365 $Y=1.765 $X2=0 $Y2=0
cc_231 N_A_c_285_n N_Y_c_406_n 0.00807097f $X=2.93 $Y=1.22 $X2=0 $Y2=0
cc_232 N_A_c_287_n N_Y_c_406_n 0.0010977f $X=3.26 $Y=1.385 $X2=0 $Y2=0
cc_233 N_A_c_285_n N_Y_c_407_n 0.00786622f $X=2.93 $Y=1.22 $X2=0 $Y2=0
cc_234 N_A_c_288_n N_A_490_368#_c_488_n 0.0119611f $X=2.915 $Y=1.765 $X2=0 $Y2=0
cc_235 N_A_c_289_n N_A_490_368#_c_488_n 0.00961384f $X=3.365 $Y=1.765 $X2=0
+ $Y2=0
cc_236 N_A_c_289_n N_A_490_368#_c_480_n 0.00469694f $X=3.365 $Y=1.765 $X2=0
+ $Y2=0
cc_237 N_A_c_288_n N_A_490_368#_c_481_n 0.00269641f $X=2.915 $Y=1.765 $X2=0
+ $Y2=0
cc_238 N_A_c_288_n N_VPWR_c_509_n 0.00644223f $X=2.915 $Y=1.765 $X2=0 $Y2=0
cc_239 N_A_c_289_n N_VPWR_c_509_n 0.00647849f $X=3.365 $Y=1.765 $X2=0 $Y2=0
cc_240 N_A_c_288_n N_VPWR_c_510_n 0.00413917f $X=2.915 $Y=1.765 $X2=0 $Y2=0
cc_241 N_A_c_289_n N_VPWR_c_511_n 0.00413917f $X=3.365 $Y=1.765 $X2=0 $Y2=0
cc_242 N_A_c_288_n N_VPWR_c_508_n 0.00399473f $X=2.915 $Y=1.765 $X2=0 $Y2=0
cc_243 N_A_c_289_n N_VPWR_c_508_n 0.00398725f $X=3.365 $Y=1.765 $X2=0 $Y2=0
cc_244 N_A_c_285_n N_VGND_c_556_n 0.00434272f $X=2.93 $Y=1.22 $X2=0 $Y2=0
cc_245 N_A_c_285_n N_VGND_c_557_n 0.00279441f $X=2.93 $Y=1.22 $X2=0 $Y2=0
cc_246 A N_VGND_c_557_n 0.0248105f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_247 N_A_c_287_n N_VGND_c_557_n 0.00378955f $X=3.26 $Y=1.385 $X2=0 $Y2=0
cc_248 N_A_c_285_n N_VGND_c_560_n 0.00825157f $X=2.93 $Y=1.22 $X2=0 $Y2=0
cc_249 N_A_27_368#_c_335_n N_A_116_368#_M1002_s 0.00425462f $X=2.035 $Y=2.405
+ $X2=-0.19 $Y2=1.66
cc_250 N_A_27_368#_c_335_n N_A_116_368#_M1010_d 0.0039188f $X=2.035 $Y=2.405
+ $X2=0 $Y2=0
cc_251 N_A_27_368#_c_328_n N_A_116_368#_c_387_n 0.0226667f $X=0.28 $Y=2.495
+ $X2=0 $Y2=0
cc_252 N_A_27_368#_c_335_n N_A_116_368#_c_387_n 0.0673127f $X=2.035 $Y=2.405
+ $X2=0 $Y2=0
cc_253 N_A_27_368#_c_329_n N_A_116_368#_c_387_n 0.0226667f $X=2.12 $Y=2.815
+ $X2=0 $Y2=0
cc_254 N_A_27_368#_c_335_n N_Y_M1000_s 0.00446629f $X=2.035 $Y=2.405 $X2=0 $Y2=0
cc_255 N_A_27_368#_M1002_d N_Y_c_410_n 0.00132795f $X=0.135 $Y=1.84 $X2=0 $Y2=0
cc_256 N_A_27_368#_c_332_n N_Y_c_410_n 0.0125997f $X=0.28 $Y=2.155 $X2=0 $Y2=0
cc_257 N_A_27_368#_c_333_n N_Y_c_406_n 0.00675162f $X=2.12 $Y=1.985 $X2=0 $Y2=0
cc_258 N_A_27_368#_c_335_n Y 0.0445038f $X=2.035 $Y=2.405 $X2=0 $Y2=0
cc_259 N_A_27_368#_c_335_n N_Y_c_412_n 0.00455859f $X=2.035 $Y=2.405 $X2=0 $Y2=0
cc_260 N_A_27_368#_c_332_n N_Y_c_412_n 0.0128526f $X=0.28 $Y=2.155 $X2=0 $Y2=0
cc_261 N_A_27_368#_c_348_n N_A_490_368#_M1001_d 0.00598865f $X=3.94 $Y=2.135
+ $X2=-0.19 $Y2=1.66
cc_262 N_A_27_368#_c_348_n N_A_490_368#_M1004_s 0.00395946f $X=3.94 $Y=2.135
+ $X2=0 $Y2=0
cc_263 N_A_27_368#_c_348_n N_A_490_368#_c_488_n 0.0343548f $X=3.94 $Y=2.135
+ $X2=0 $Y2=0
cc_264 N_A_27_368#_c_348_n N_A_490_368#_c_485_n 0.0154464f $X=3.94 $Y=2.135
+ $X2=0 $Y2=0
cc_265 N_A_27_368#_c_331_n N_A_490_368#_c_480_n 0.0148001f $X=4.04 $Y=2.815
+ $X2=0 $Y2=0
cc_266 N_A_27_368#_c_329_n N_A_490_368#_c_481_n 0.00143161f $X=2.12 $Y=2.815
+ $X2=0 $Y2=0
cc_267 N_A_27_368#_c_348_n N_A_490_368#_c_481_n 0.022257f $X=3.94 $Y=2.135 $X2=0
+ $Y2=0
cc_268 N_A_27_368#_c_348_n N_VPWR_M1003_d 0.00385736f $X=3.94 $Y=2.135 $X2=-0.19
+ $Y2=1.66
cc_269 N_A_27_368#_c_328_n N_VPWR_c_510_n 0.0120294f $X=0.28 $Y=2.495 $X2=0
+ $Y2=0
cc_270 N_A_27_368#_c_329_n N_VPWR_c_510_n 0.011066f $X=2.12 $Y=2.815 $X2=0 $Y2=0
cc_271 N_A_27_368#_c_331_n N_VPWR_c_511_n 0.0117353f $X=4.04 $Y=2.815 $X2=0
+ $Y2=0
cc_272 N_A_27_368#_c_328_n N_VPWR_c_508_n 0.00926813f $X=0.28 $Y=2.495 $X2=0
+ $Y2=0
cc_273 N_A_27_368#_c_335_n N_VPWR_c_508_n 0.0108943f $X=2.035 $Y=2.405 $X2=0
+ $Y2=0
cc_274 N_A_27_368#_c_329_n N_VPWR_c_508_n 0.00915947f $X=2.12 $Y=2.815 $X2=0
+ $Y2=0
cc_275 N_A_27_368#_c_331_n N_VPWR_c_508_n 0.00971347f $X=4.04 $Y=2.815 $X2=0
+ $Y2=0
cc_276 N_A_27_368#_c_332_n N_VPWR_c_508_n 0.00286949f $X=0.28 $Y=2.155 $X2=0
+ $Y2=0
cc_277 N_A_116_368#_c_387_n N_Y_M1000_s 0.00229266f $X=1.67 $Y=2.78 $X2=0 $Y2=0
cc_278 N_A_116_368#_M1002_s Y 0.00273805f $X=0.58 $Y=1.84 $X2=0 $Y2=0
cc_279 N_A_116_368#_c_387_n N_VPWR_c_510_n 0.0525924f $X=1.67 $Y=2.78 $X2=0
+ $Y2=0
cc_280 N_A_116_368#_c_387_n N_VPWR_c_508_n 0.0441578f $X=1.67 $Y=2.78 $X2=0
+ $Y2=0
cc_281 N_Y_c_403_n N_VGND_M1009_s 0.0045742f $X=1.55 $Y=0.915 $X2=-0.19
+ $Y2=-0.245
cc_282 N_Y_c_406_n N_VGND_M1007_d 0.00368125f $X=2.55 $Y=1.065 $X2=0 $Y2=0
cc_283 N_Y_c_405_n N_VGND_c_555_n 0.0180508f $X=1.715 $Y=0.515 $X2=0 $Y2=0
cc_284 N_Y_c_406_n N_VGND_c_555_n 0.0248957f $X=2.55 $Y=1.065 $X2=0 $Y2=0
cc_285 N_Y_c_407_n N_VGND_c_555_n 0.0180508f $X=2.715 $Y=0.515 $X2=0 $Y2=0
cc_286 N_Y_c_407_n N_VGND_c_556_n 0.0144922f $X=2.715 $Y=0.515 $X2=0 $Y2=0
cc_287 N_Y_c_407_n N_VGND_c_557_n 0.0243921f $X=2.715 $Y=0.515 $X2=0 $Y2=0
cc_288 N_Y_c_405_n N_VGND_c_558_n 0.0145639f $X=1.715 $Y=0.515 $X2=0 $Y2=0
cc_289 N_Y_c_403_n N_VGND_c_560_n 0.0130998f $X=1.55 $Y=0.915 $X2=0 $Y2=0
cc_290 N_Y_c_404_n N_VGND_c_560_n 0.00111297f $X=0.255 $Y=0.915 $X2=0 $Y2=0
cc_291 N_Y_c_405_n N_VGND_c_560_n 0.0119984f $X=1.715 $Y=0.515 $X2=0 $Y2=0
cc_292 N_Y_c_407_n N_VGND_c_560_n 0.0118826f $X=2.715 $Y=0.515 $X2=0 $Y2=0
cc_293 N_Y_c_403_n N_VGND_c_562_n 0.0436524f $X=1.55 $Y=0.915 $X2=0 $Y2=0
cc_294 N_Y_c_405_n N_VGND_c_562_n 0.00167954f $X=1.715 $Y=0.515 $X2=0 $Y2=0
cc_295 N_A_490_368#_c_488_n N_VPWR_M1003_d 0.00392025f $X=3.505 $Y=2.475
+ $X2=-0.19 $Y2=1.66
cc_296 N_A_490_368#_c_488_n N_VPWR_c_509_n 0.0166996f $X=3.505 $Y=2.475 $X2=0
+ $Y2=0
cc_297 N_A_490_368#_c_480_n N_VPWR_c_509_n 0.0181628f $X=3.59 $Y=2.835 $X2=0
+ $Y2=0
cc_298 N_A_490_368#_c_481_n N_VPWR_c_509_n 0.0117536f $X=2.64 $Y=2.495 $X2=0
+ $Y2=0
cc_299 N_A_490_368#_c_481_n N_VPWR_c_510_n 0.0157837f $X=2.64 $Y=2.495 $X2=0
+ $Y2=0
cc_300 N_A_490_368#_c_480_n N_VPWR_c_511_n 0.0118914f $X=3.59 $Y=2.835 $X2=0
+ $Y2=0
cc_301 N_A_490_368#_c_488_n N_VPWR_c_508_n 0.0127927f $X=3.505 $Y=2.475 $X2=0
+ $Y2=0
cc_302 N_A_490_368#_c_480_n N_VPWR_c_508_n 0.00916858f $X=3.59 $Y=2.835 $X2=0
+ $Y2=0
cc_303 N_A_490_368#_c_481_n N_VPWR_c_508_n 0.0122146f $X=2.64 $Y=2.495 $X2=0
+ $Y2=0
