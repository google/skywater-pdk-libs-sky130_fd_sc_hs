* File: sky130_fd_sc_hs__xor3_2.pex.spice
* Created: Thu Aug 27 21:13:25 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HS__XOR3_2%A_83_289# 1 2 3 4 15 17 19 22 25 26 30 33 35
+ 36 38 41 43 44 49
c109 26 0 1.40857e-19 $X=0.745 $Y=2.005
r110 47 49 5.5876 $w=3.28e-07 $l=1.6e-07 $layer=LI1_cond $X=4.15 $Y=1.1 $X2=4.31
+ $Y2=1.1
r111 43 45 19.8947 $w=6.68e-07 $l=6.85e-07 $layer=LI1_cond $X=4.06 $Y=2.07
+ $X2=4.06 $Y2=2.755
r112 43 44 10.6117 $w=6.68e-07 $l=1.65e-07 $layer=LI1_cond $X=4.06 $Y=2.07
+ $X2=4.06 $Y2=1.905
r113 39 49 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.31 $Y=1.265
+ $X2=4.31 $Y2=1.1
r114 39 44 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=4.31 $Y=1.265
+ $X2=4.31 $Y2=1.905
r115 38 45 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=3.81 $Y=2.905
+ $X2=3.81 $Y2=2.755
r116 35 38 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.725 $Y=2.99
+ $X2=3.81 $Y2=2.905
r117 35 36 136.027 $w=1.68e-07 $l=2.085e-06 $layer=LI1_cond $X=3.725 $Y=2.99
+ $X2=1.64 $Y2=2.99
r118 31 41 3.70735 $w=2.5e-07 $l=2.3e-07 $layer=LI1_cond $X=1.54 $Y=1.92
+ $X2=1.31 $Y2=1.92
r119 31 33 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=1.54 $Y=1.92
+ $X2=1.54 $Y2=1.165
r120 28 36 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.475 $Y=2.905
+ $X2=1.64 $Y2=2.99
r121 28 30 23.2235 $w=3.28e-07 $l=6.65e-07 $layer=LI1_cond $X=1.475 $Y=2.905
+ $X2=1.475 $Y2=2.24
r122 27 41 3.70735 $w=2.5e-07 $l=2.38642e-07 $layer=LI1_cond $X=1.475 $Y=2.09
+ $X2=1.31 $Y2=1.92
r123 27 30 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=1.475 $Y=2.09
+ $X2=1.475 $Y2=2.24
r124 25 41 2.76166 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.31 $Y=2.005
+ $X2=1.31 $Y2=1.92
r125 25 26 36.861 $w=1.68e-07 $l=5.65e-07 $layer=LI1_cond $X=1.31 $Y=2.005
+ $X2=0.745 $Y2=2.005
r126 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.58
+ $Y=1.61 $X2=0.58 $Y2=1.61
r127 20 26 7.68211 $w=1.7e-07 $l=1.9799e-07 $layer=LI1_cond $X=0.585 $Y=1.92
+ $X2=0.745 $Y2=2.005
r128 20 22 11.1643 $w=3.18e-07 $l=3.1e-07 $layer=LI1_cond $X=0.585 $Y=1.92
+ $X2=0.585 $Y2=1.61
r129 17 23 52.2586 $w=2.99e-07 $l=2.85044e-07 $layer=POLY_cond $X=0.655 $Y=1.86
+ $X2=0.58 $Y2=1.61
r130 17 19 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=0.655 $Y=1.86
+ $X2=0.655 $Y2=2.435
r131 13 23 38.5562 $w=2.99e-07 $l=2.03101e-07 $layer=POLY_cond $X=0.495 $Y=1.445
+ $X2=0.58 $Y2=1.61
r132 13 15 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=0.495 $Y=1.445
+ $X2=0.495 $Y2=0.99
r133 4 43 300 $w=1.7e-07 $l=5.40463e-07 $layer=licon1_PDIFF $count=2 $X=3.35
+ $Y=1.895 $X2=3.81 $Y2=2.07
r134 3 30 300 $w=1.7e-07 $l=3.72525e-07 $layer=licon1_PDIFF $count=2 $X=1.325
+ $Y=1.935 $X2=1.475 $Y2=2.24
r135 2 47 182 $w=1.7e-07 $l=6.10635e-07 $layer=licon1_NDIFF $count=1 $X=3.84
+ $Y=0.625 $X2=4.15 $Y2=1.1
r136 1 33 182 $w=1.7e-07 $l=5.60647e-07 $layer=licon1_NDIFF $count=1 $X=1.4
+ $Y=0.67 $X2=1.54 $Y2=1.165
.ends

.subckt PM_SKY130_FD_SC_HS__XOR3_2%A 1 3 4 6 7
c34 1 0 2.38282e-19 $X=1.25 $Y=1.86
r35 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.12
+ $Y=1.585 $X2=1.12 $Y2=1.585
r36 7 11 10.1275 $w=3.28e-07 $l=2.9e-07 $layer=LI1_cond $X=1.12 $Y=1.295
+ $X2=1.12 $Y2=1.585
r37 4 10 39.1844 $w=3.78e-07 $l=2.27255e-07 $layer=POLY_cond $X=1.325 $Y=1.42
+ $X2=1.177 $Y2=1.585
r38 4 6 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=1.325 $Y=1.42
+ $X2=1.325 $Y2=0.99
r39 1 10 53.2109 $w=3.78e-07 $l=3.09354e-07 $layer=POLY_cond $X=1.25 $Y=1.86
+ $X2=1.177 $Y2=1.585
r40 1 3 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=1.25 $Y=1.86 $X2=1.25
+ $Y2=2.435
.ends

.subckt PM_SKY130_FD_SC_HS__XOR3_2%A_440_315# 1 2 8 9 11 14 16 17 18 20 21 25 30
+ 33 34 35 38 45 46
c113 46 0 7.8648e-20 $X=3.89 $Y=1.57
r114 51 52 11.4717 $w=2.23e-07 $l=2.1e-07 $layer=LI1_cond $X=4.692 $Y=0.8
+ $X2=4.692 $Y2=1.01
r115 46 54 46.6671 $w=3.65e-07 $l=1.65e-07 $layer=POLY_cond $X=3.872 $Y=1.57
+ $X2=3.872 $Y2=1.405
r116 45 46 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.89
+ $Y=1.57 $X2=3.89 $Y2=1.57
r117 42 45 3.07318 $w=2.98e-07 $l=8e-08 $layer=LI1_cond $X=3.81 $Y=1.585
+ $X2=3.89 $Y2=1.585
r118 38 40 54.1497 $w=1.68e-07 $l=8.3e-07 $layer=LI1_cond $X=4.665 $Y=1.985
+ $X2=4.665 $Y2=2.815
r119 38 52 63.6096 $w=1.68e-07 $l=9.75e-07 $layer=LI1_cond $X=4.665 $Y=1.985
+ $X2=4.665 $Y2=1.01
r120 34 51 6.14636 $w=2.23e-07 $l=1.2e-07 $layer=LI1_cond $X=4.692 $Y=0.68
+ $X2=4.692 $Y2=0.8
r121 34 35 44.6898 $w=1.68e-07 $l=6.85e-07 $layer=LI1_cond $X=4.58 $Y=0.68
+ $X2=3.895 $Y2=0.68
r122 33 42 4.061 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=3.81 $Y=1.435 $X2=3.81
+ $Y2=1.585
r123 32 35 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.81 $Y=0.765
+ $X2=3.895 $Y2=0.68
r124 32 33 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.81 $Y=0.765
+ $X2=3.81 $Y2=1.435
r125 25 54 235.872 $w=1.5e-07 $l=4.6e-07 $layer=POLY_cond $X=3.765 $Y=0.945
+ $X2=3.765 $Y2=1.405
r126 22 30 7.1379 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=3.365 $Y=1.65
+ $X2=3.275 $Y2=1.65
r127 21 46 12.6475 $w=3.65e-07 $l=8e-08 $layer=POLY_cond $X=3.872 $Y=1.65
+ $X2=3.872 $Y2=1.57
r128 21 22 166.649 $w=1.5e-07 $l=3.25e-07 $layer=POLY_cond $X=3.69 $Y=1.65
+ $X2=3.365 $Y2=1.65
r129 18 30 68.2304 $w=1.8e-07 $l=1.7e-07 $layer=POLY_cond $X=3.275 $Y=1.82
+ $X2=3.275 $Y2=1.65
r130 18 20 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=3.275 $Y=1.82
+ $X2=3.275 $Y2=2.315
r131 17 29 38.4574 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.58 $Y=1.65
+ $X2=2.505 $Y2=1.65
r132 16 30 7.1379 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=3.185 $Y=1.65
+ $X2=3.275 $Y2=1.65
r133 16 17 310.223 $w=1.5e-07 $l=6.05e-07 $layer=POLY_cond $X=3.185 $Y=1.65
+ $X2=2.58 $Y2=1.65
r134 12 29 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.505 $Y=1.575
+ $X2=2.505 $Y2=1.65
r135 12 14 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=2.505 $Y=1.575
+ $X2=2.505 $Y2=0.995
r136 9 11 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=2.29 $Y=2.02
+ $X2=2.29 $Y2=2.415
r137 8 9 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=2.29 $Y=1.93 $X2=2.29
+ $Y2=2.02
r138 7 29 110.245 $w=1.5e-07 $l=2.15e-07 $layer=POLY_cond $X=2.29 $Y=1.65
+ $X2=2.505 $Y2=1.65
r139 7 8 79.6855 $w=1.8e-07 $l=2.05e-07 $layer=POLY_cond $X=2.29 $Y=1.725
+ $X2=2.29 $Y2=1.93
r140 2 40 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=4.52
+ $Y=1.84 $X2=4.665 $Y2=2.815
r141 2 38 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=4.52
+ $Y=1.84 $X2=4.665 $Y2=1.985
r142 1 51 182 $w=1.7e-07 $l=4.929e-07 $layer=licon1_NDIFF $count=1 $X=4.585
+ $Y=0.37 $X2=4.72 $Y2=0.8
.ends

.subckt PM_SKY130_FD_SC_HS__XOR3_2%B 1 3 4 5 8 10 11 12 13 14 16 17 21 23 25 26
+ 28 29 31 33 34 36 37 38 40
c131 34 0 1.39206e-19 $X=4.935 $Y=1.22
c132 21 0 1.51563e-19 $X=3.175 $Y=0.885
c133 8 0 1.54943e-19 $X=2.005 $Y=0.885
r134 44 45 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.085
+ $Y=1.385 $X2=5.085 $Y2=1.385
r135 42 44 12.6472 $w=3.43e-07 $l=9e-08 $layer=POLY_cond $X=5.025 $Y=1.295
+ $X2=5.025 $Y2=1.385
r136 40 45 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=5.085 $Y=1.295
+ $X2=5.085 $Y2=1.385
r137 34 42 26.0611 $w=3.43e-07 $l=1.21861e-07 $layer=POLY_cond $X=4.935 $Y=1.22
+ $X2=5.025 $Y2=1.295
r138 34 36 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=4.935 $Y=1.22
+ $X2=4.935 $Y2=0.74
r139 31 44 68.9212 $w=3.43e-07 $l=4.4238e-07 $layer=POLY_cond $X=4.89 $Y=1.765
+ $X2=5.025 $Y2=1.385
r140 31 33 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=4.89 $Y=1.765
+ $X2=4.89 $Y2=2.4
r141 30 39 7.39479 $w=1.5e-07 $l=1.08e-07 $layer=POLY_cond $X=4.51 $Y=1.295
+ $X2=4.402 $Y2=1.295
r142 29 42 22.1447 $w=1.5e-07 $l=2.25e-07 $layer=POLY_cond $X=4.8 $Y=1.295
+ $X2=5.025 $Y2=1.295
r143 29 30 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=4.8 $Y=1.295
+ $X2=4.51 $Y2=1.295
r144 28 39 21.4953 $w=1.82e-07 $l=9e-08 $layer=POLY_cond $X=4.435 $Y=1.22
+ $X2=4.402 $Y2=1.295
r145 27 28 494.819 $w=1.5e-07 $l=9.65e-07 $layer=POLY_cond $X=4.435 $Y=0.255
+ $X2=4.435 $Y2=1.22
r146 25 39 61.2206 $w=1.82e-07 $l=2.40468e-07 $layer=POLY_cond $X=4.37 $Y=1.52
+ $X2=4.402 $Y2=1.295
r147 25 26 797.351 $w=1.5e-07 $l=1.555e-06 $layer=POLY_cond $X=4.37 $Y=1.52
+ $X2=4.37 $Y2=3.075
r148 24 38 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.25 $Y=0.18
+ $X2=3.175 $Y2=0.18
r149 23 27 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.36 $Y=0.18
+ $X2=4.435 $Y2=0.255
r150 23 24 569.17 $w=1.5e-07 $l=1.11e-06 $layer=POLY_cond $X=4.36 $Y=0.18
+ $X2=3.25 $Y2=0.18
r151 19 38 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.175 $Y=0.255
+ $X2=3.175 $Y2=0.18
r152 19 21 323.043 $w=1.5e-07 $l=6.3e-07 $layer=POLY_cond $X=3.175 $Y=0.255
+ $X2=3.175 $Y2=0.885
r153 18 37 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=2.83 $Y=3.15 $X2=2.74
+ $Y2=3.15
r154 17 26 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.295 $Y=3.15
+ $X2=4.37 $Y2=3.075
r155 17 18 751.202 $w=1.5e-07 $l=1.465e-06 $layer=POLY_cond $X=4.295 $Y=3.15
+ $X2=2.83 $Y2=3.15
r156 14 16 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=2.74 $Y=2.81
+ $X2=2.74 $Y2=2.415
r157 13 37 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=2.74 $Y=3.075
+ $X2=2.74 $Y2=3.15
r158 12 14 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=2.74 $Y=2.9 $X2=2.74
+ $Y2=2.81
r159 12 13 68.0242 $w=1.8e-07 $l=1.75e-07 $layer=POLY_cond $X=2.74 $Y=2.9
+ $X2=2.74 $Y2=3.075
r160 10 38 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.1 $Y=0.18
+ $X2=3.175 $Y2=0.18
r161 10 11 523.021 $w=1.5e-07 $l=1.02e-06 $layer=POLY_cond $X=3.1 $Y=0.18
+ $X2=2.08 $Y2=0.18
r162 6 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.005 $Y=0.255
+ $X2=2.08 $Y2=0.18
r163 6 8 323.043 $w=1.5e-07 $l=6.3e-07 $layer=POLY_cond $X=2.005 $Y=0.255
+ $X2=2.005 $Y2=0.885
r164 4 37 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=2.65 $Y=3.15 $X2=2.74
+ $Y2=3.15
r165 4 5 397.394 $w=1.5e-07 $l=7.75e-07 $layer=POLY_cond $X=2.65 $Y=3.15
+ $X2=1.875 $Y2=3.15
r166 1 5 26.9307 $w=1.5e-07 $l=1.79444e-07 $layer=POLY_cond $X=1.785 $Y=3.01
+ $X2=1.875 $Y2=3.15
r167 1 3 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=1.785 $Y=3.01
+ $X2=1.785 $Y2=2.515
.ends

.subckt PM_SKY130_FD_SC_HS__XOR3_2%A_1162_379# 1 2 7 9 12 15 18 21 22 23 25 27
+ 28 30 33 34
c108 30 0 2.73932e-20 $X=7.86 $Y=0.6
c109 27 0 3.42466e-19 $X=7.72 $Y=2.195
c110 15 0 1.62191e-19 $X=6.155 $Y=1.895
c111 12 0 1.40994e-19 $X=6.155 $Y=0.855
r112 37 40 3.0228 $w=3.03e-07 $l=8e-08 $layer=LI1_cond $X=7.365 $Y=2.347
+ $X2=7.445 $Y2=2.347
r113 34 49 45.2517 $w=3.8e-07 $l=1.65e-07 $layer=POLY_cond $X=6.04 $Y=1.52
+ $X2=6.04 $Y2=1.685
r114 34 48 45.2517 $w=3.8e-07 $l=1.65e-07 $layer=POLY_cond $X=6.04 $Y=1.52
+ $X2=6.04 $Y2=1.355
r115 33 36 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=6.015 $Y=1.52
+ $X2=6.015 $Y2=1.685
r116 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.015
+ $Y=1.52 $X2=6.015 $Y2=1.52
r117 28 43 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=7.9 $Y=1.52
+ $X2=7.72 $Y2=1.52
r118 28 30 38.4916 $w=2.48e-07 $l=8.35e-07 $layer=LI1_cond $X=7.9 $Y=1.435
+ $X2=7.9 $Y2=0.6
r119 27 40 10.3909 $w=3.03e-07 $l=2.75e-07 $layer=LI1_cond $X=7.72 $Y=2.347
+ $X2=7.445 $Y2=2.347
r120 26 43 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.72 $Y=1.605
+ $X2=7.72 $Y2=1.52
r121 26 27 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=7.72 $Y=1.605
+ $X2=7.72 $Y2=2.195
r122 24 37 4.15824 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=7.365 $Y=2.5
+ $X2=7.365 $Y2=2.347
r123 24 25 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=7.365 $Y=2.5
+ $X2=7.365 $Y2=2.905
r124 22 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.28 $Y=2.99
+ $X2=7.365 $Y2=2.905
r125 22 23 71.7647 $w=1.68e-07 $l=1.1e-06 $layer=LI1_cond $X=7.28 $Y=2.99
+ $X2=6.18 $Y2=2.99
r126 21 23 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.095 $Y=2.905
+ $X2=6.18 $Y2=2.99
r127 21 36 79.5936 $w=1.68e-07 $l=1.22e-06 $layer=LI1_cond $X=6.095 $Y=2.905
+ $X2=6.095 $Y2=1.685
r128 16 18 130.755 $w=1.5e-07 $l=2.55e-07 $layer=POLY_cond $X=5.9 $Y=1.97
+ $X2=6.155 $Y2=1.97
r129 15 18 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.155 $Y=1.895
+ $X2=6.155 $Y2=1.97
r130 15 49 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=6.155 $Y=1.895
+ $X2=6.155 $Y2=1.685
r131 12 48 256.383 $w=1.5e-07 $l=5e-07 $layer=POLY_cond $X=6.155 $Y=0.855
+ $X2=6.155 $Y2=1.355
r132 7 16 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.9 $Y=2.045 $X2=5.9
+ $Y2=1.97
r133 7 9 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=5.9 $Y=2.045 $X2=5.9
+ $Y2=2.54
r134 2 40 600 $w=1.7e-07 $l=5.32588e-07 $layer=licon1_PDIFF $count=1 $X=7.3
+ $Y=1.84 $X2=7.445 $Y2=2.305
r135 1 30 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=7.715
+ $Y=0.39 $X2=7.86 $Y2=0.6
.ends

.subckt PM_SKY130_FD_SC_HS__XOR3_2%C 2 3 5 6 8 9 10 12 13 15 16 17 18 20 22
c97 22 0 2.73932e-20 $X=6.96 $Y=1.295
c98 12 0 1.05114e-19 $X=7.735 $Y=1.355
c99 9 0 1.48172e-19 $X=7.66 $Y=1.43
r100 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.975
+ $Y=1.52 $X2=6.975 $Y2=1.52
r101 25 27 24.9926 $w=2.7e-07 $l=1.4e-07 $layer=POLY_cond $X=6.835 $Y=1.52
+ $X2=6.975 $Y2=1.52
r102 22 28 10.372 $w=2.48e-07 $l=2.25e-07 $layer=LI1_cond $X=7 $Y=1.295 $X2=7
+ $Y2=1.52
r103 18 20 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=8.075 $Y=0.885
+ $X2=8.075 $Y2=0.6
r104 16 18 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=8 $Y=0.96
+ $X2=8.075 $Y2=0.885
r105 16 17 97.4255 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=8 $Y=0.96 $X2=7.81
+ $Y2=0.96
r106 13 21 96.2697 $w=1.69e-07 $l=3.35e-07 $layer=POLY_cond $X=7.75 $Y=1.765
+ $X2=7.75 $Y2=1.43
r107 13 15 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=7.75 $Y=1.765
+ $X2=7.75 $Y2=2.16
r108 12 21 22.1159 $w=1.69e-07 $l=8.21584e-08 $layer=POLY_cond $X=7.735 $Y=1.355
+ $X2=7.75 $Y2=1.43
r109 11 17 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=7.735 $Y=1.035
+ $X2=7.81 $Y2=0.96
r110 11 12 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=7.735 $Y=1.035
+ $X2=7.735 $Y2=1.355
r111 10 27 38.9026 $w=2.7e-07 $l=2.05122e-07 $layer=POLY_cond $X=7.14 $Y=1.43
+ $X2=6.975 $Y2=1.52
r112 9 21 5.66465 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=7.66 $Y=1.43 $X2=7.75
+ $Y2=1.43
r113 9 10 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=7.66 $Y=1.43
+ $X2=7.14 $Y2=1.43
r114 6 25 16.5046 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.835 $Y=1.355
+ $X2=6.835 $Y2=1.52
r115 6 8 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=6.835 $Y=1.355
+ $X2=6.835 $Y2=0.925
r116 3 5 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=6.66 $Y=2.045
+ $X2=6.66 $Y2=2.54
r117 2 3 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=6.66 $Y=1.955 $X2=6.66
+ $Y2=2.045
r118 1 25 31.2407 $w=2.7e-07 $l=2.43926e-07 $layer=POLY_cond $X=6.66 $Y=1.685
+ $X2=6.835 $Y2=1.52
r119 1 2 104.952 $w=1.8e-07 $l=2.7e-07 $layer=POLY_cond $X=6.66 $Y=1.685
+ $X2=6.66 $Y2=1.955
.ends

.subckt PM_SKY130_FD_SC_HS__XOR3_2%A_1195_424# 1 2 7 9 12 14 17 20 22 24 25 26
+ 27 30 34 37 41 42 45 48 49
c112 49 0 1.49322e-19 $X=8.4 $Y=2.035
c113 37 0 1.05114e-19 $X=8.36 $Y=1.485
c114 25 0 1.94294e-19 $X=8.555 $Y=1.485
r115 48 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=2.035
+ $X2=8.4 $Y2=2.035
r116 45 55 18.4391 $w=2.48e-07 $l=4e-07 $layer=LI1_cond $X=6.475 $Y=2.035
+ $X2=6.475 $Y2=2.435
r117 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=2.035
+ $X2=6.48 $Y2=2.035
r118 42 44 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.625 $Y=2.035
+ $X2=6.48 $Y2=2.035
r119 41 48 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=8.255 $Y=2.035
+ $X2=8.4 $Y2=2.035
r120 41 42 2.01732 $w=1.4e-07 $l=1.63e-06 $layer=MET1_cond $X=8.255 $Y=2.035
+ $X2=6.625 $Y2=2.035
r121 40 49 20.3333 $w=2.08e-07 $l=3.85e-07 $layer=LI1_cond $X=8.42 $Y=1.65
+ $X2=8.42 $Y2=2.035
r122 37 40 7.28026 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=8.36 $Y=1.485
+ $X2=8.36 $Y2=1.65
r123 37 38 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.36
+ $Y=1.485 $X2=8.36 $Y2=1.485
r124 34 45 23.5098 $w=2.48e-07 $l=5.1e-07 $layer=LI1_cond $X=6.475 $Y=1.525
+ $X2=6.475 $Y2=2.035
r125 33 34 9.02376 $w=2.48e-07 $l=1.7e-07 $layer=LI1_cond $X=6.527 $Y=1.355
+ $X2=6.527 $Y2=1.525
r126 30 33 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=6.62 $Y=1.1
+ $X2=6.62 $Y2=1.355
r127 25 38 34.0979 $w=3.3e-07 $l=1.95e-07 $layer=POLY_cond $X=8.555 $Y=1.485
+ $X2=8.36 $Y2=1.485
r128 25 26 6.91837 $w=3.3e-07 $l=1.15022e-07 $layer=POLY_cond $X=8.555 $Y=1.485
+ $X2=8.645 $Y2=1.542
r129 22 24 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=9.095 $Y=1.765
+ $X2=9.095 $Y2=2.4
r130 18 27 18.8402 $w=1.65e-07 $l=7.98436e-08 $layer=POLY_cond $X=9.085 $Y=1.32
+ $X2=9.095 $Y2=1.395
r131 18 20 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=9.085 $Y=1.32
+ $X2=9.085 $Y2=0.76
r132 17 22 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=9.095 $Y=1.675
+ $X2=9.095 $Y2=1.765
r133 16 27 18.8402 $w=1.65e-07 $l=7.5e-08 $layer=POLY_cond $X=9.095 $Y=1.47
+ $X2=9.095 $Y2=1.395
r134 16 17 79.6855 $w=1.8e-07 $l=2.05e-07 $layer=POLY_cond $X=9.095 $Y=1.47
+ $X2=9.095 $Y2=1.675
r135 15 26 6.91837 $w=1.5e-07 $l=1.86652e-07 $layer=POLY_cond $X=8.735 $Y=1.395
+ $X2=8.645 $Y2=1.542
r136 14 27 6.66866 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=9.005 $Y=1.395
+ $X2=9.095 $Y2=1.395
r137 14 15 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=9.005 $Y=1.395
+ $X2=8.735 $Y2=1.395
r138 10 26 18.1359 $w=1.5e-07 $l=2.26945e-07 $layer=POLY_cond $X=8.655 $Y=1.32
+ $X2=8.645 $Y2=1.542
r139 10 12 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=8.655 $Y=1.32
+ $X2=8.655 $Y2=0.76
r140 7 26 18.1359 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=8.645 $Y=1.765
+ $X2=8.645 $Y2=1.542
r141 7 9 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=8.645 $Y=1.765
+ $X2=8.645 $Y2=2.4
r142 2 55 600 $w=1.7e-07 $l=5.97076e-07 $layer=licon1_PDIFF $count=1 $X=5.975
+ $Y=2.12 $X2=6.435 $Y2=2.435
r143 1 30 182 $w=1.7e-07 $l=7.34558e-07 $layer=licon1_NDIFF $count=1 $X=6.23
+ $Y=0.535 $X2=6.62 $Y2=1.1
.ends

.subckt PM_SKY130_FD_SC_HS__XOR3_2%A_27_134# 1 2 3 4 13 14 17 20 21 22 25 28 31
+ 33 34 36 40
r87 37 40 5.07033 $w=4.58e-07 $l=1.95e-07 $layer=LI1_cond $X=2.595 $Y=0.995
+ $X2=2.79 $Y2=0.995
r88 33 34 9.57885 $w=5.08e-07 $l=1.65e-07 $layer=LI1_cond $X=0.34 $Y=2.425
+ $X2=0.34 $Y2=2.26
r89 31 34 64.262 $w=1.68e-07 $l=9.85e-07 $layer=LI1_cond $X=0.17 $Y=1.275
+ $X2=0.17 $Y2=2.26
r90 28 36 3.70735 $w=2.5e-07 $l=1.18427e-07 $layer=LI1_cond $X=2.595 $Y=1.395
+ $X2=2.515 $Y2=1.48
r91 27 37 6.6364 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=2.595 $Y=1.225
+ $X2=2.595 $Y2=0.995
r92 27 28 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=2.595 $Y=1.225
+ $X2=2.595 $Y2=1.395
r93 23 36 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.515 $Y=1.565
+ $X2=2.515 $Y2=1.48
r94 23 25 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=2.515 $Y=1.565
+ $X2=2.515 $Y2=2.275
r95 21 36 2.76166 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.35 $Y=1.48
+ $X2=2.515 $Y2=1.48
r96 21 22 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=2.35 $Y=1.48
+ $X2=1.965 $Y2=1.48
r97 20 22 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.88 $Y=1.395
+ $X2=1.965 $Y2=1.48
r98 19 20 36.861 $w=1.68e-07 $l=5.65e-07 $layer=LI1_cond $X=1.88 $Y=0.83
+ $X2=1.88 $Y2=1.395
r99 18 30 5.39736 $w=1.7e-07 $l=1.82483e-07 $layer=LI1_cond $X=0.445 $Y=0.745
+ $X2=0.265 $Y2=0.74
r100 17 19 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.795 $Y=0.745
+ $X2=1.88 $Y2=0.83
r101 17 18 88.0749 $w=1.68e-07 $l=1.35e-06 $layer=LI1_cond $X=1.795 $Y=0.745
+ $X2=0.445 $Y2=0.745
r102 14 31 8.99121 $w=3.58e-07 $l=1.8e-07 $layer=LI1_cond $X=0.265 $Y=1.095
+ $X2=0.265 $Y2=1.275
r103 13 30 2.62574 $w=3.6e-07 $l=9e-08 $layer=LI1_cond $X=0.265 $Y=0.83
+ $X2=0.265 $Y2=0.74
r104 13 14 8.48326 $w=3.58e-07 $l=2.65e-07 $layer=LI1_cond $X=0.265 $Y=0.83
+ $X2=0.265 $Y2=1.095
r105 4 25 600 $w=1.7e-07 $l=2.43721e-07 $layer=licon1_PDIFF $count=1 $X=2.365
+ $Y=2.095 $X2=2.515 $Y2=2.275
r106 3 33 300 $w=1.7e-07 $l=5.57808e-07 $layer=licon1_PDIFF $count=2 $X=0.285
+ $Y=1.935 $X2=0.43 $Y2=2.425
r107 2 40 182 $w=1.7e-07 $l=2.96985e-07 $layer=licon1_NDIFF $count=1 $X=2.58
+ $Y=0.785 $X2=2.79 $Y2=0.995
r108 1 30 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.67 $X2=0.28 $Y2=0.815
.ends

.subckt PM_SKY130_FD_SC_HS__XOR3_2%VPWR 1 2 3 4 15 19 25 28 29 31 36 37 39 41 47
+ 54 62 68 71 75
r98 74 75 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.36 $Y=3.33
+ $X2=9.36 $Y2=3.33
r99 71 72 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=3.33 $X2=8.4
+ $Y2=3.33
r100 68 69 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r101 66 75 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=3.33
+ $X2=9.36 $Y2=3.33
r102 66 72 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=3.33
+ $X2=8.4 $Y2=3.33
r103 65 66 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r104 63 71 12.0118 $w=1.7e-07 $l=2.78e-07 $layer=LI1_cond $X=8.53 $Y=3.33
+ $X2=8.252 $Y2=3.33
r105 63 65 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=8.53 $Y=3.33
+ $X2=8.88 $Y2=3.33
r106 62 74 4.01252 $w=1.7e-07 $l=1.82e-07 $layer=LI1_cond $X=9.235 $Y=3.33
+ $X2=9.417 $Y2=3.33
r107 62 65 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=9.235 $Y=3.33
+ $X2=8.88 $Y2=3.33
r108 61 72 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=3.33
+ $X2=8.4 $Y2=3.33
r109 60 61 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r110 58 61 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=7.92 $Y2=3.33
r111 58 69 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=5.04 $Y2=3.33
r112 57 60 156.578 $w=1.68e-07 $l=2.4e-06 $layer=LI1_cond $X=5.52 $Y=3.33
+ $X2=7.92 $Y2=3.33
r113 57 58 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r114 55 68 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.2 $Y=3.33
+ $X2=5.075 $Y2=3.33
r115 55 57 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=5.2 $Y=3.33 $X2=5.52
+ $Y2=3.33
r116 54 71 12.0118 $w=1.7e-07 $l=2.77e-07 $layer=LI1_cond $X=7.975 $Y=3.33
+ $X2=8.252 $Y2=3.33
r117 54 60 3.58824 $w=1.68e-07 $l=5.5e-08 $layer=LI1_cond $X=7.975 $Y=3.33
+ $X2=7.92 $Y2=3.33
r118 52 53 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r119 50 53 0.936549 $w=4.9e-07 $l=3.36e-06 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=4.56 $Y2=3.33
r120 49 52 219.209 $w=1.68e-07 $l=3.36e-06 $layer=LI1_cond $X=1.2 $Y=3.33
+ $X2=4.56 $Y2=3.33
r121 49 50 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r122 47 68 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.95 $Y=3.33
+ $X2=5.075 $Y2=3.33
r123 47 52 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=4.95 $Y=3.33
+ $X2=4.56 $Y2=3.33
r124 45 50 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r125 44 45 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r126 41 69 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=4.8 $Y=3.33
+ $X2=5.04 $Y2=3.33
r127 41 53 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=4.8 $Y=3.33
+ $X2=4.56 $Y2=3.33
r128 39 40 9.86413 $w=5.53e-07 $l=1.65e-07 $layer=LI1_cond $X=8.252 $Y=2.485
+ $X2=8.252 $Y2=2.32
r129 36 44 2.93583 $w=1.68e-07 $l=4.5e-08 $layer=LI1_cond $X=0.765 $Y=3.33
+ $X2=0.72 $Y2=3.33
r130 36 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.765 $Y=3.33
+ $X2=0.93 $Y2=3.33
r131 35 49 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=1.095 $Y=3.33
+ $X2=1.2 $Y2=3.33
r132 35 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.095 $Y=3.33
+ $X2=0.93 $Y2=3.33
r133 31 34 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=9.36 $Y=1.985
+ $X2=9.36 $Y2=2.815
r134 29 74 3.13065 $w=2.5e-07 $l=1.09864e-07 $layer=LI1_cond $X=9.36 $Y=3.245
+ $X2=9.417 $Y2=3.33
r135 29 34 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=9.36 $Y=3.245
+ $X2=9.36 $Y2=2.815
r136 28 71 2.33542 $w=5.55e-07 $l=8.5e-08 $layer=LI1_cond $X=8.252 $Y=3.245
+ $X2=8.252 $Y2=3.33
r137 27 39 2.41371 $w=5.53e-07 $l=1.12e-07 $layer=LI1_cond $X=8.252 $Y=2.597
+ $X2=8.252 $Y2=2.485
r138 27 28 13.965 $w=5.53e-07 $l=6.48e-07 $layer=LI1_cond $X=8.252 $Y=2.597
+ $X2=8.252 $Y2=3.245
r139 25 40 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=8.06 $Y=1.985
+ $X2=8.06 $Y2=2.32
r140 19 22 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=5.075 $Y=1.985
+ $X2=5.075 $Y2=2.815
r141 17 68 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.075 $Y=3.245
+ $X2=5.075 $Y2=3.33
r142 17 22 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=5.075 $Y=3.245
+ $X2=5.075 $Y2=2.815
r143 13 37 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.93 $Y=3.245
+ $X2=0.93 $Y2=3.33
r144 13 15 28.6365 $w=3.28e-07 $l=8.2e-07 $layer=LI1_cond $X=0.93 $Y=3.245
+ $X2=0.93 $Y2=2.425
r145 4 34 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=9.17
+ $Y=1.84 $X2=9.32 $Y2=2.815
r146 4 31 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=9.17
+ $Y=1.84 $X2=9.32 $Y2=1.985
r147 3 39 200 $w=1.7e-07 $l=8.94315e-07 $layer=licon1_PDIFF $count=3 $X=7.825
+ $Y=1.84 $X2=8.42 $Y2=2.485
r148 3 25 300 $w=1.7e-07 $l=2.98831e-07 $layer=licon1_PDIFF $count=2 $X=7.825
+ $Y=1.84 $X2=8.06 $Y2=1.985
r149 2 22 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=4.965
+ $Y=1.84 $X2=5.115 $Y2=2.815
r150 2 19 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=4.965
+ $Y=1.84 $X2=5.115 $Y2=1.985
r151 1 15 300 $w=1.7e-07 $l=5.81464e-07 $layer=licon1_PDIFF $count=2 $X=0.73
+ $Y=1.935 $X2=0.93 $Y2=2.425
.ends

.subckt PM_SKY130_FD_SC_HS__XOR3_2%A_372_419# 1 2 3 4 15 17 18 22 23 24 26 27 28
+ 30 31 32 35 37 38 40 42 47
c147 22 0 7.8648e-20 $X=3.47 $Y=0.71
c148 18 0 2.51379e-19 $X=2.18 $Y=2.65
c149 15 0 1.82528e-19 $X=2.015 $Y=2.24
r150 45 47 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=7.38 $Y=1.18
+ $X2=7.52 $Y2=1.18
r151 42 47 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.52 $Y=1.095
+ $X2=7.52 $Y2=1.18
r152 41 42 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=7.52 $Y=0.425
+ $X2=7.52 $Y2=1.095
r153 39 45 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.38 $Y=1.265
+ $X2=7.38 $Y2=1.18
r154 39 40 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=7.38 $Y=1.265
+ $X2=7.38 $Y2=1.855
r155 37 40 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.295 $Y=1.94
+ $X2=7.38 $Y2=1.855
r156 37 38 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=7.295 $Y=1.94
+ $X2=7.05 $Y2=1.94
r157 33 38 7.24806 $w=1.7e-07 $l=1.70276e-07 $layer=LI1_cond $X=6.917 $Y=2.025
+ $X2=7.05 $Y2=1.94
r158 33 35 17.8302 $w=2.63e-07 $l=4.1e-07 $layer=LI1_cond $X=6.917 $Y=2.025
+ $X2=6.917 $Y2=2.435
r159 31 41 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.435 $Y=0.34
+ $X2=7.52 $Y2=0.425
r160 31 32 91.9893 $w=1.68e-07 $l=1.41e-06 $layer=LI1_cond $X=7.435 $Y=0.34
+ $X2=6.025 $Y2=0.34
r161 30 44 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.9 $Y=0.675 $X2=5.9
+ $Y2=0.76
r162 29 32 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=5.9 $Y=0.425
+ $X2=6.025 $Y2=0.34
r163 29 30 11.5244 $w=2.48e-07 $l=2.5e-07 $layer=LI1_cond $X=5.9 $Y=0.425
+ $X2=5.9 $Y2=0.675
r164 27 44 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.775 $Y=0.76
+ $X2=5.9 $Y2=0.76
r165 27 28 41.1016 $w=1.68e-07 $l=6.3e-07 $layer=LI1_cond $X=5.775 $Y=0.76
+ $X2=5.145 $Y2=0.76
r166 26 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.06 $Y=0.675
+ $X2=5.145 $Y2=0.76
r167 25 26 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=5.06 $Y=0.425
+ $X2=5.06 $Y2=0.675
r168 23 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.975 $Y=0.34
+ $X2=5.06 $Y2=0.425
r169 23 24 92.6417 $w=1.68e-07 $l=1.42e-06 $layer=LI1_cond $X=4.975 $Y=0.34
+ $X2=3.555 $Y2=0.34
r170 20 22 121.021 $w=1.68e-07 $l=1.855e-06 $layer=LI1_cond $X=3.47 $Y=2.565
+ $X2=3.47 $Y2=0.71
r171 19 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.47 $Y=0.425
+ $X2=3.555 $Y2=0.34
r172 19 22 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=3.47 $Y=0.425
+ $X2=3.47 $Y2=0.71
r173 17 20 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.385 $Y=2.65
+ $X2=3.47 $Y2=2.565
r174 17 18 78.615 $w=1.68e-07 $l=1.205e-06 $layer=LI1_cond $X=3.385 $Y=2.65
+ $X2=2.18 $Y2=2.65
r175 13 18 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.015 $Y=2.565
+ $X2=2.18 $Y2=2.65
r176 13 15 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=2.015 $Y=2.565
+ $X2=2.015 $Y2=2.24
r177 4 35 600 $w=1.7e-07 $l=3.82721e-07 $layer=licon1_PDIFF $count=1 $X=6.735
+ $Y=2.12 $X2=6.885 $Y2=2.435
r178 3 15 300 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_PDIFF $count=2 $X=1.86
+ $Y=2.095 $X2=2.015 $Y2=2.24
r179 2 44 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=5.805
+ $Y=0.535 $X2=5.94 $Y2=0.68
r180 1 22 91 $w=1.7e-07 $l=2.83373e-07 $layer=licon1_NDIFF $count=2 $X=3.25
+ $Y=0.565 $X2=3.47 $Y2=0.71
.ends

.subckt PM_SKY130_FD_SC_HS__XOR3_2%A_416_113# 1 2 3 4 15 17 18 21 27 31 32 34 36
+ 38 39 41 42 45 48 49 52 54
c125 54 0 3.01398e-19 $X=5.622 $Y=1.92
c126 42 0 1.51563e-19 $X=3.265 $Y=2.035
c127 38 0 1.40994e-19 $X=7.075 $Y=0.76
c128 15 0 1.54943e-19 $X=2.22 $Y=0.71
r129 49 54 7.48521 $w=4.33e-07 $l=1.15e-07 $layer=LI1_cond $X=5.622 $Y=2.035
+ $X2=5.622 $Y2=1.92
r130 48 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=2.035
+ $X2=5.52 $Y2=2.035
r131 45 52 8.28756 $w=3.28e-07 $l=1.6e-07 $layer=LI1_cond $X=3.05 $Y=2.035
+ $X2=3.05 $Y2=1.875
r132 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=2.035
+ $X2=3.12 $Y2=2.035
r133 42 44 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.265 $Y=2.035
+ $X2=3.12 $Y2=2.035
r134 41 48 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.375 $Y=2.035
+ $X2=5.52 $Y2=2.035
r135 41 42 2.61138 $w=1.4e-07 $l=2.11e-06 $layer=MET1_cond $X=5.375 $Y=2.035
+ $X2=3.265 $Y2=2.035
r136 38 39 9.33524 $w=3.28e-07 $l=1.9e-07 $layer=LI1_cond $X=7.075 $Y=0.76
+ $X2=6.885 $Y2=0.76
r137 36 39 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=6.365 $Y=0.68
+ $X2=6.885 $Y2=0.68
r138 33 36 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.28 $Y=0.765
+ $X2=6.365 $Y2=0.68
r139 33 34 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=6.28 $Y=0.765
+ $X2=6.28 $Y2=1.015
r140 31 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.195 $Y=1.1
+ $X2=6.28 $Y2=1.015
r141 31 32 33.5989 $w=1.68e-07 $l=5.15e-07 $layer=LI1_cond $X=6.195 $Y=1.1
+ $X2=5.68 $Y2=1.1
r142 29 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.595 $Y=1.185
+ $X2=5.68 $Y2=1.1
r143 29 54 47.9519 $w=1.68e-07 $l=7.35e-07 $layer=LI1_cond $X=5.595 $Y=1.185
+ $X2=5.595 $Y2=1.92
r144 25 49 2.70228 $w=4.33e-07 $l=1.02e-07 $layer=LI1_cond $X=5.622 $Y=2.137
+ $X2=5.622 $Y2=2.035
r145 25 27 3.3911 $w=4.33e-07 $l=1.28e-07 $layer=LI1_cond $X=5.622 $Y=2.137
+ $X2=5.622 $Y2=2.265
r146 23 52 83.508 $w=1.68e-07 $l=1.28e-06 $layer=LI1_cond $X=3.13 $Y=0.595
+ $X2=3.13 $Y2=1.875
r147 19 45 0.174613 $w=3.28e-07 $l=5e-09 $layer=LI1_cond $X=3.05 $Y=2.04
+ $X2=3.05 $Y2=2.035
r148 19 21 3.31764 $w=3.28e-07 $l=9.5e-08 $layer=LI1_cond $X=3.05 $Y=2.04
+ $X2=3.05 $Y2=2.135
r149 17 23 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.045 $Y=0.51
+ $X2=3.13 $Y2=0.595
r150 17 18 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=3.045 $Y=0.51
+ $X2=2.305 $Y2=0.51
r151 13 18 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.22 $Y=0.595
+ $X2=2.305 $Y2=0.51
r152 13 15 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=2.22 $Y=0.595
+ $X2=2.22 $Y2=0.71
r153 4 27 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=5.53
+ $Y=2.12 $X2=5.675 $Y2=2.265
r154 3 21 600 $w=1.7e-07 $l=2.54214e-07 $layer=licon1_PDIFF $count=1 $X=2.815
+ $Y=2.095 $X2=3.05 $Y2=2.135
r155 2 38 182 $w=1.7e-07 $l=2.29783e-07 $layer=licon1_NDIFF $count=1 $X=6.91
+ $Y=0.605 $X2=7.075 $Y2=0.76
r156 1 15 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.08
+ $Y=0.565 $X2=2.22 $Y2=0.71
.ends

.subckt PM_SKY130_FD_SC_HS__XOR3_2%X 1 2 7 8 9 10 11 12 13
r21 12 13 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=8.87 $Y=2.405
+ $X2=8.87 $Y2=2.775
r22 11 12 14.6675 $w=3.28e-07 $l=4.2e-07 $layer=LI1_cond $X=8.87 $Y=1.985
+ $X2=8.87 $Y2=2.405
r23 10 11 11.1752 $w=3.28e-07 $l=3.2e-07 $layer=LI1_cond $X=8.87 $Y=1.665
+ $X2=8.87 $Y2=1.985
r24 9 10 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=8.87 $Y=1.295
+ $X2=8.87 $Y2=1.665
r25 8 9 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=8.87 $Y=0.925 $X2=8.87
+ $Y2=1.295
r26 7 8 13.6198 $w=3.28e-07 $l=3.9e-07 $layer=LI1_cond $X=8.87 $Y=0.535 $X2=8.87
+ $Y2=0.925
r27 2 13 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=8.72
+ $Y=1.84 $X2=8.87 $Y2=2.815
r28 2 11 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=8.72
+ $Y=1.84 $X2=8.87 $Y2=1.985
r29 1 7 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=8.73
+ $Y=0.39 $X2=8.87 $Y2=0.535
.ends

.subckt PM_SKY130_FD_SC_HS__XOR3_2%VGND 1 2 3 4 15 19 23 25 27 34 42 47 55 58 60
+ 63 67
r81 66 67 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.36 $Y=0 $X2=9.36
+ $Y2=0
r82 63 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r83 60 61 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r84 57 58 12.4896 $w=5.73e-07 $l=2.85e-07 $layer=LI1_cond $X=0.91 $Y=0.202
+ $X2=1.195 $Y2=0.202
r85 53 57 3.95226 $w=5.73e-07 $l=1.9e-07 $layer=LI1_cond $X=0.72 $Y=0.202
+ $X2=0.91 $Y2=0.202
r86 53 55 8.53733 $w=5.73e-07 $l=9.5e-08 $layer=LI1_cond $X=0.72 $Y=0.202
+ $X2=0.625 $Y2=0.202
r87 53 54 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r88 51 67 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=0 $X2=9.36
+ $Y2=0
r89 51 64 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=0 $X2=8.4
+ $Y2=0
r90 50 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=0 $X2=8.88
+ $Y2=0
r91 48 63 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.535 $Y=0 $X2=8.37
+ $Y2=0
r92 48 50 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=8.535 $Y=0 $X2=8.88
+ $Y2=0
r93 47 66 3.98688 $w=1.7e-07 $l=1.92e-07 $layer=LI1_cond $X=9.215 $Y=0 $X2=9.407
+ $Y2=0
r94 47 50 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=9.215 $Y=0 $X2=8.88
+ $Y2=0
r95 46 64 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=0 $X2=8.4
+ $Y2=0
r96 46 61 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=7.92 $Y=0 $X2=5.52
+ $Y2=0
r97 45 46 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=7.92 $Y=0 $X2=7.92
+ $Y2=0
r98 43 60 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.565 $Y=0 $X2=5.44
+ $Y2=0
r99 43 45 153.642 $w=1.68e-07 $l=2.355e-06 $layer=LI1_cond $X=5.565 $Y=0
+ $X2=7.92 $Y2=0
r100 42 63 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.205 $Y=0 $X2=8.37
+ $Y2=0
r101 42 45 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=8.205 $Y=0
+ $X2=7.92 $Y2=0
r102 41 61 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=5.52
+ $Y2=0
r103 40 41 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=5.04 $Y=0
+ $X2=5.04 $Y2=0
r104 38 54 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r105 37 40 250.524 $w=1.68e-07 $l=3.84e-06 $layer=LI1_cond $X=1.2 $Y=0 $X2=5.04
+ $Y2=0
r106 37 58 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=1.2 $Y=0 $X2=1.195
+ $Y2=0
r107 37 38 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=1.2 $Y=0
+ $X2=1.2 $Y2=0
r108 34 60 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.315 $Y=0 $X2=5.44
+ $Y2=0
r109 34 40 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=5.315 $Y=0
+ $X2=5.04 $Y2=0
r110 32 54 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r111 31 55 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=0.24 $Y=0
+ $X2=0.625 $Y2=0
r112 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r113 27 41 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=4.8 $Y=0 $X2=5.04
+ $Y2=0
r114 27 38 1.00344 $w=4.9e-07 $l=3.6e-06 $layer=MET1_cond $X=4.8 $Y=0 $X2=1.2
+ $Y2=0
r115 23 66 3.15628 $w=2.5e-07 $l=1.13666e-07 $layer=LI1_cond $X=9.34 $Y=0.085
+ $X2=9.407 $Y2=0
r116 23 25 20.744 $w=2.48e-07 $l=4.5e-07 $layer=LI1_cond $X=9.34 $Y=0.085
+ $X2=9.34 $Y2=0.535
r117 19 21 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=8.37 $Y=0.535
+ $X2=8.37 $Y2=0.985
r118 17 63 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.37 $Y=0.085
+ $X2=8.37 $Y2=0
r119 17 19 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=8.37 $Y=0.085
+ $X2=8.37 $Y2=0.535
r120 13 60 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.44 $Y=0.085
+ $X2=5.44 $Y2=0
r121 13 15 11.7549 $w=2.48e-07 $l=2.55e-07 $layer=LI1_cond $X=5.44 $Y=0.085
+ $X2=5.44 $Y2=0.34
r122 4 25 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=9.16
+ $Y=0.39 $X2=9.3 $Y2=0.535
r123 3 21 182 $w=1.7e-07 $l=6.96366e-07 $layer=licon1_NDIFF $count=1 $X=8.15
+ $Y=0.39 $X2=8.37 $Y2=0.985
r124 3 19 182 $w=1.7e-07 $l=2.83373e-07 $layer=licon1_NDIFF $count=1 $X=8.15
+ $Y=0.39 $X2=8.37 $Y2=0.535
r125 2 15 182 $w=1.7e-07 $l=4.04722e-07 $layer=licon1_NDIFF $count=1 $X=5.01
+ $Y=0.37 $X2=5.4 $Y2=0.34
r126 1 57 182 $w=1.7e-07 $l=4.86133e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.67 $X2=0.91 $Y2=0.325
.ends

