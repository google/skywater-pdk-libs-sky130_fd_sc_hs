* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hs__a32oi_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
X0 Y A1 a_507_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X1 a_27_368# A3 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X2 a_27_74# B1 Y VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X3 a_27_368# A2 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X4 VGND B2 a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X5 Y B2 a_27_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X6 VGND A3 a_771_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X7 Y B1 a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X8 VPWR A3 a_27_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X9 a_27_368# B1 Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X10 a_771_74# A2 a_507_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X11 a_507_74# A2 a_771_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X12 a_771_74# A3 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X13 Y B1 a_27_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X14 VPWR A1 a_27_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X15 a_507_74# A1 Y VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X16 a_27_368# B2 Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X17 VPWR A2 a_27_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X18 a_27_368# A1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X19 a_27_74# B2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
.ends
