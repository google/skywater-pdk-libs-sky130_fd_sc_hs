* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hs__bufbuf_16 A VGND VNB VPB VPWR X
X0 a_27_368# A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X1 VPWR a_588_74# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X2 VPWR a_588_74# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X3 VGND a_588_74# X VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X4 VPWR a_588_74# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X5 a_203_74# a_27_368# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X6 VPWR a_588_74# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X7 VGND a_203_74# a_588_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X8 VGND a_203_74# a_588_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X9 VGND a_203_74# a_588_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X10 VPWR a_588_74# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X11 X a_588_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X12 a_588_74# a_203_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X13 X a_588_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X14 a_588_74# a_203_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X15 X a_588_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X16 VGND a_588_74# X VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X17 a_588_74# a_203_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X18 a_588_74# a_203_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X19 a_588_74# a_203_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X20 VPWR a_203_74# a_588_74# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X21 X a_588_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X22 a_27_368# A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X23 X a_588_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X24 a_588_74# a_203_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X25 VGND a_588_74# X VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X26 VPWR a_27_368# a_203_74# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X27 X a_588_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X28 X a_588_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X29 X a_588_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X30 X a_588_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X31 VGND a_588_74# X VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X32 VPWR a_588_74# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X33 VPWR a_27_368# a_203_74# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X34 X a_588_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X35 VPWR a_203_74# a_588_74# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X36 a_203_74# a_27_368# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X37 VGND a_588_74# X VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X38 VGND a_588_74# X VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X39 VGND a_588_74# X VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X40 VPWR a_588_74# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X41 VPWR a_588_74# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X42 VPWR a_203_74# a_588_74# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X43 X a_588_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X44 X a_588_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X45 VGND a_27_368# a_203_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X46 X a_588_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X47 VGND a_27_368# a_203_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X48 X a_588_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X49 VGND a_588_74# X VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X50 X a_588_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X51 X a_588_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
.ends
