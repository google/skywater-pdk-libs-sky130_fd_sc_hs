* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hs__or2b_2 A B_N VGND VNB VPB VPWR X
M1000 X a_187_48# VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=5.768e+11p pd=3.27e+06u as=8.614e+11p ps=6.09e+06u
M1001 a_470_368# A VPWR VPB pshort w=1e+06u l=150000u
+  ad=2.7e+11p pd=2.54e+06u as=0p ps=0u
M1002 VGND B_N a_27_368# VNB nlowvt w=550000u l=150000u
+  ad=9.5555e+11p pd=7.08e+06u as=1.5675e+11p ps=1.67e+06u
M1003 a_187_48# A VGND VNB nlowvt w=640000u l=150000u
+  ad=2.208e+11p pd=1.97e+06u as=0p ps=0u
M1004 a_187_48# a_27_368# a_470_368# VPB pshort w=1e+06u l=150000u
+  ad=4.15e+11p pd=2.83e+06u as=0p ps=0u
M1005 X a_187_48# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1006 VGND a_187_48# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VPWR B_N a_27_368# VPB pshort w=840000u l=150000u
+  ad=0p pd=0u as=2.478e+11p ps=2.27e+06u
M1008 VGND a_27_368# a_187_48# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VPWR a_187_48# X VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
