* File: sky130_fd_sc_hs__nand2_2.pxi.spice
* Created: Thu Aug 27 20:50:05 2020
* 
x_PM_SKY130_FD_SC_HS__NAND2_2%B N_B_M1004_g N_B_c_49_n N_B_M1001_g N_B_c_50_n
+ N_B_M1003_g N_B_M1005_g B B N_B_c_48_n PM_SKY130_FD_SC_HS__NAND2_2%B
x_PM_SKY130_FD_SC_HS__NAND2_2%A N_A_M1000_g N_A_c_89_n N_A_M1006_g N_A_c_90_n
+ N_A_M1007_g N_A_M1002_g A N_A_c_87_n N_A_c_88_n PM_SKY130_FD_SC_HS__NAND2_2%A
x_PM_SKY130_FD_SC_HS__NAND2_2%VPWR N_VPWR_M1001_d N_VPWR_M1003_d N_VPWR_M1007_s
+ N_VPWR_c_134_n N_VPWR_c_135_n N_VPWR_c_136_n N_VPWR_c_137_n N_VPWR_c_138_n
+ VPWR N_VPWR_c_139_n N_VPWR_c_140_n N_VPWR_c_141_n N_VPWR_c_133_n
+ PM_SKY130_FD_SC_HS__NAND2_2%VPWR
x_PM_SKY130_FD_SC_HS__NAND2_2%Y N_Y_M1000_d N_Y_M1001_s N_Y_M1006_d N_Y_c_180_n
+ N_Y_c_176_n N_Y_c_185_n N_Y_c_189_n N_Y_c_177_n N_Y_c_178_n N_Y_c_173_n
+ N_Y_c_174_n N_Y_c_199_n Y Y PM_SKY130_FD_SC_HS__NAND2_2%Y
x_PM_SKY130_FD_SC_HS__NAND2_2%A_27_74# N_A_27_74#_M1004_d N_A_27_74#_M1005_d
+ N_A_27_74#_M1002_s N_A_27_74#_c_224_n N_A_27_74#_c_225_n N_A_27_74#_c_226_n
+ N_A_27_74#_c_227_n N_A_27_74#_c_228_n N_A_27_74#_c_229_n
+ PM_SKY130_FD_SC_HS__NAND2_2%A_27_74#
x_PM_SKY130_FD_SC_HS__NAND2_2%VGND N_VGND_M1004_s N_VGND_c_258_n VGND
+ N_VGND_c_259_n N_VGND_c_260_n N_VGND_c_261_n N_VGND_c_262_n
+ PM_SKY130_FD_SC_HS__NAND2_2%VGND
cc_1 VNB N_B_M1004_g 0.0325972f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_2 VNB N_B_M1005_g 0.0243544f $X=-0.19 $Y=-0.245 $X2=0.975 $Y2=0.74
cc_3 VNB B 0.00631699f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.58
cc_4 VNB N_B_c_48_n 0.0453658f $X=-0.19 $Y=-0.245 $X2=0.96 $Y2=1.557
cc_5 VNB N_A_M1000_g 0.0236545f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_6 VNB N_A_M1002_g 0.0267831f $X=-0.19 $Y=-0.245 $X2=0.975 $Y2=0.74
cc_7 VNB N_A_c_87_n 0.00139482f $X=-0.19 $Y=-0.245 $X2=0.77 $Y2=1.557
cc_8 VNB N_A_c_88_n 0.0387716f $X=-0.19 $Y=-0.245 $X2=0.77 $Y2=1.515
cc_9 VNB N_VPWR_c_133_n 0.103974f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_Y_c_173_n 0.0105096f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.565
cc_11 VNB N_Y_c_174_n 0.0025404f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB Y 0.0241052f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_27_74#_c_224_n 0.0266107f $X=-0.19 $Y=-0.245 $X2=0.975 $Y2=0.74
cc_14 VNB N_A_27_74#_c_225_n 0.00790826f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_27_74#_c_226_n 0.0116953f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_16 VNB N_A_27_74#_c_227_n 0.0126678f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=1.557
cc_17 VNB N_A_27_74#_c_228_n 0.00217191f $X=-0.19 $Y=-0.245 $X2=0.77 $Y2=1.557
cc_18 VNB N_A_27_74#_c_229_n 0.0161735f $X=-0.19 $Y=-0.245 $X2=0.96 $Y2=1.557
cc_19 VNB N_VGND_c_258_n 0.00615265f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=2.4
cc_20 VNB N_VGND_c_259_n 0.0173909f $X=-0.19 $Y=-0.245 $X2=0.96 $Y2=2.4
cc_21 VNB N_VGND_c_260_n 0.0392768f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=1.557
cc_22 VNB N_VGND_c_261_n 0.163114f $X=-0.19 $Y=-0.245 $X2=0.77 $Y2=1.557
cc_23 VNB N_VGND_c_262_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0.96 $Y2=1.557
cc_24 VPB N_B_c_49_n 0.0177521f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=1.765
cc_25 VPB N_B_c_50_n 0.0151845f $X=-0.19 $Y=1.66 $X2=0.96 $Y2=1.765
cc_26 VPB B 0.00730124f $X=-0.19 $Y=1.66 $X2=1.115 $Y2=1.58
cc_27 VPB N_B_c_48_n 0.0234619f $X=-0.19 $Y=1.66 $X2=0.96 $Y2=1.557
cc_28 VPB N_A_c_89_n 0.0151869f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=1.765
cc_29 VPB N_A_c_90_n 0.0171509f $X=-0.19 $Y=1.66 $X2=0.96 $Y2=1.765
cc_30 VPB N_A_c_87_n 0.00279203f $X=-0.19 $Y=1.66 $X2=0.77 $Y2=1.557
cc_31 VPB N_A_c_88_n 0.0204862f $X=-0.19 $Y=1.66 $X2=0.77 $Y2=1.515
cc_32 VPB N_VPWR_c_134_n 0.0108116f $X=-0.19 $Y=1.66 $X2=0.96 $Y2=2.4
cc_33 VPB N_VPWR_c_135_n 0.0579743f $X=-0.19 $Y=1.66 $X2=0.975 $Y2=0.74
cc_34 VPB N_VPWR_c_136_n 0.00273118f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_35 VPB N_VPWR_c_137_n 0.012808f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=1.557
cc_36 VPB N_VPWR_c_138_n 0.035054f $X=-0.19 $Y=1.66 $X2=0.77 $Y2=1.515
cc_37 VPB N_VPWR_c_139_n 0.0185253f $X=-0.19 $Y=1.66 $X2=0.72 $Y2=1.565
cc_38 VPB N_VPWR_c_140_n 0.0167647f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_39 VPB N_VPWR_c_141_n 0.00601644f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_40 VPB N_VPWR_c_133_n 0.0597142f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_41 VPB N_Y_c_176_n 0.00216998f $X=-0.19 $Y=1.66 $X2=0.975 $Y2=0.74
cc_42 VPB N_Y_c_177_n 0.00181113f $X=-0.19 $Y=1.66 $X2=0.77 $Y2=1.515
cc_43 VPB N_Y_c_178_n 0.00793272f $X=-0.19 $Y=1.66 $X2=0.96 $Y2=1.557
cc_44 VPB Y 0.0131059f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_45 N_B_M1005_g N_A_M1000_g 0.0184614f $X=0.975 $Y=0.74 $X2=0 $Y2=0
cc_46 N_B_c_50_n N_A_c_89_n 0.0254772f $X=0.96 $Y=1.765 $X2=0 $Y2=0
cc_47 B N_A_c_87_n 0.0361808f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_48 N_B_c_48_n N_A_c_87_n 2.76228e-19 $X=0.96 $Y=1.557 $X2=0 $Y2=0
cc_49 B N_A_c_88_n 0.00423515f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_50 N_B_c_48_n N_A_c_88_n 0.0184614f $X=0.96 $Y=1.557 $X2=0 $Y2=0
cc_51 N_B_c_49_n N_VPWR_c_135_n 0.0110944f $X=0.51 $Y=1.765 $X2=0 $Y2=0
cc_52 N_B_c_49_n N_VPWR_c_136_n 5.55114e-19 $X=0.51 $Y=1.765 $X2=0 $Y2=0
cc_53 N_B_c_50_n N_VPWR_c_136_n 0.0111612f $X=0.96 $Y=1.765 $X2=0 $Y2=0
cc_54 N_B_c_49_n N_VPWR_c_139_n 0.00445602f $X=0.51 $Y=1.765 $X2=0 $Y2=0
cc_55 N_B_c_50_n N_VPWR_c_139_n 0.00413917f $X=0.96 $Y=1.765 $X2=0 $Y2=0
cc_56 N_B_c_49_n N_VPWR_c_133_n 0.008611f $X=0.51 $Y=1.765 $X2=0 $Y2=0
cc_57 N_B_c_50_n N_VPWR_c_133_n 0.00817726f $X=0.96 $Y=1.765 $X2=0 $Y2=0
cc_58 N_B_c_49_n N_Y_c_180_n 0.00256038f $X=0.51 $Y=1.765 $X2=0 $Y2=0
cc_59 B N_Y_c_180_n 0.0173447f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_60 N_B_c_48_n N_Y_c_180_n 0.0012279f $X=0.96 $Y=1.557 $X2=0 $Y2=0
cc_61 N_B_c_49_n N_Y_c_176_n 0.00955225f $X=0.51 $Y=1.765 $X2=0 $Y2=0
cc_62 N_B_c_50_n N_Y_c_176_n 0.00605728f $X=0.96 $Y=1.765 $X2=0 $Y2=0
cc_63 N_B_c_50_n N_Y_c_185_n 0.0126897f $X=0.96 $Y=1.765 $X2=0 $Y2=0
cc_64 B N_Y_c_185_n 0.0332333f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_65 N_B_M1004_g N_A_27_74#_c_224_n 0.00159319f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_66 N_B_M1004_g N_A_27_74#_c_225_n 0.018438f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_67 N_B_M1005_g N_A_27_74#_c_225_n 0.013919f $X=0.975 $Y=0.74 $X2=0 $Y2=0
cc_68 B N_A_27_74#_c_225_n 0.0533206f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_69 N_B_c_48_n N_A_27_74#_c_225_n 0.00336308f $X=0.96 $Y=1.557 $X2=0 $Y2=0
cc_70 N_B_M1005_g N_A_27_74#_c_228_n 0.00106427f $X=0.975 $Y=0.74 $X2=0 $Y2=0
cc_71 N_B_M1004_g N_VGND_c_258_n 0.0132976f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_72 N_B_M1005_g N_VGND_c_258_n 0.00192886f $X=0.975 $Y=0.74 $X2=0 $Y2=0
cc_73 N_B_M1004_g N_VGND_c_259_n 0.00383152f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_74 N_B_M1005_g N_VGND_c_260_n 0.00461464f $X=0.975 $Y=0.74 $X2=0 $Y2=0
cc_75 N_B_M1004_g N_VGND_c_261_n 0.00761198f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_76 N_B_M1005_g N_VGND_c_261_n 0.00908237f $X=0.975 $Y=0.74 $X2=0 $Y2=0
cc_77 N_A_c_89_n N_VPWR_c_136_n 0.01018f $X=1.42 $Y=1.765 $X2=0 $Y2=0
cc_78 N_A_c_90_n N_VPWR_c_136_n 5.35026e-19 $X=1.87 $Y=1.765 $X2=0 $Y2=0
cc_79 N_A_c_89_n N_VPWR_c_138_n 5.37287e-19 $X=1.42 $Y=1.765 $X2=0 $Y2=0
cc_80 N_A_c_90_n N_VPWR_c_138_n 0.0120347f $X=1.87 $Y=1.765 $X2=0 $Y2=0
cc_81 N_A_c_89_n N_VPWR_c_140_n 0.00444681f $X=1.42 $Y=1.765 $X2=0 $Y2=0
cc_82 N_A_c_90_n N_VPWR_c_140_n 0.00413917f $X=1.87 $Y=1.765 $X2=0 $Y2=0
cc_83 N_A_c_89_n N_VPWR_c_133_n 0.00877716f $X=1.42 $Y=1.765 $X2=0 $Y2=0
cc_84 N_A_c_90_n N_VPWR_c_133_n 0.00817726f $X=1.87 $Y=1.765 $X2=0 $Y2=0
cc_85 N_A_c_89_n N_Y_c_185_n 0.017247f $X=1.42 $Y=1.765 $X2=0 $Y2=0
cc_86 N_A_c_87_n N_Y_c_185_n 0.00371182f $X=1.65 $Y=1.515 $X2=0 $Y2=0
cc_87 N_A_M1000_g N_Y_c_189_n 0.00543663f $X=1.405 $Y=0.74 $X2=0 $Y2=0
cc_88 N_A_c_89_n N_Y_c_177_n 0.00564785f $X=1.42 $Y=1.765 $X2=0 $Y2=0
cc_89 N_A_c_90_n N_Y_c_177_n 0.00554978f $X=1.87 $Y=1.765 $X2=0 $Y2=0
cc_90 N_A_c_90_n N_Y_c_178_n 0.0180153f $X=1.87 $Y=1.765 $X2=0 $Y2=0
cc_91 N_A_c_87_n N_Y_c_178_n 0.00444519f $X=1.65 $Y=1.515 $X2=0 $Y2=0
cc_92 N_A_M1002_g N_Y_c_173_n 0.0177903f $X=1.885 $Y=0.74 $X2=0 $Y2=0
cc_93 N_A_c_87_n N_Y_c_173_n 0.0021829f $X=1.65 $Y=1.515 $X2=0 $Y2=0
cc_94 N_A_M1000_g N_Y_c_174_n 0.00468846f $X=1.405 $Y=0.74 $X2=0 $Y2=0
cc_95 N_A_c_87_n N_Y_c_174_n 0.0254953f $X=1.65 $Y=1.515 $X2=0 $Y2=0
cc_96 N_A_c_88_n N_Y_c_174_n 0.00116618f $X=1.87 $Y=1.557 $X2=0 $Y2=0
cc_97 N_A_c_87_n N_Y_c_199_n 0.0150976f $X=1.65 $Y=1.515 $X2=0 $Y2=0
cc_98 N_A_c_88_n N_Y_c_199_n 0.00104415f $X=1.87 $Y=1.557 $X2=0 $Y2=0
cc_99 N_A_c_90_n Y 0.00679847f $X=1.87 $Y=1.765 $X2=0 $Y2=0
cc_100 N_A_M1002_g Y 0.0182332f $X=1.885 $Y=0.74 $X2=0 $Y2=0
cc_101 N_A_c_87_n Y 0.0263485f $X=1.65 $Y=1.515 $X2=0 $Y2=0
cc_102 N_A_M1000_g N_A_27_74#_c_225_n 5.7448e-19 $X=1.405 $Y=0.74 $X2=0 $Y2=0
cc_103 N_A_M1000_g N_A_27_74#_c_227_n 0.0122924f $X=1.405 $Y=0.74 $X2=0 $Y2=0
cc_104 N_A_M1002_g N_A_27_74#_c_227_n 0.0121629f $X=1.885 $Y=0.74 $X2=0 $Y2=0
cc_105 N_A_M1000_g N_A_27_74#_c_229_n 8.69012e-19 $X=1.405 $Y=0.74 $X2=0 $Y2=0
cc_106 N_A_M1002_g N_A_27_74#_c_229_n 0.00614869f $X=1.885 $Y=0.74 $X2=0 $Y2=0
cc_107 N_A_M1000_g N_VGND_c_260_n 0.00278271f $X=1.405 $Y=0.74 $X2=0 $Y2=0
cc_108 N_A_M1002_g N_VGND_c_260_n 0.00278266f $X=1.885 $Y=0.74 $X2=0 $Y2=0
cc_109 N_A_M1000_g N_VGND_c_261_n 0.00354005f $X=1.405 $Y=0.74 $X2=0 $Y2=0
cc_110 N_A_M1002_g N_VGND_c_261_n 0.00357631f $X=1.885 $Y=0.74 $X2=0 $Y2=0
cc_111 N_VPWR_c_135_n N_Y_c_180_n 0.0121024f $X=0.285 $Y=1.985 $X2=0 $Y2=0
cc_112 N_VPWR_c_135_n N_Y_c_176_n 0.0564818f $X=0.285 $Y=1.985 $X2=0 $Y2=0
cc_113 N_VPWR_c_136_n N_Y_c_176_n 0.0462948f $X=1.185 $Y=2.455 $X2=0 $Y2=0
cc_114 N_VPWR_c_139_n N_Y_c_176_n 0.0110241f $X=1.02 $Y=3.33 $X2=0 $Y2=0
cc_115 N_VPWR_c_133_n N_Y_c_176_n 0.00909194f $X=2.16 $Y=3.33 $X2=0 $Y2=0
cc_116 N_VPWR_M1003_d N_Y_c_185_n 0.00417211f $X=1.035 $Y=1.84 $X2=0 $Y2=0
cc_117 N_VPWR_c_136_n N_Y_c_185_n 0.0172332f $X=1.185 $Y=2.455 $X2=0 $Y2=0
cc_118 N_VPWR_c_136_n N_Y_c_177_n 0.043319f $X=1.185 $Y=2.455 $X2=0 $Y2=0
cc_119 N_VPWR_c_138_n N_Y_c_177_n 0.0449718f $X=2.095 $Y=2.455 $X2=0 $Y2=0
cc_120 N_VPWR_c_140_n N_Y_c_177_n 0.00749631f $X=1.93 $Y=3.33 $X2=0 $Y2=0
cc_121 N_VPWR_c_133_n N_Y_c_177_n 0.0062048f $X=2.16 $Y=3.33 $X2=0 $Y2=0
cc_122 N_VPWR_M1007_s N_Y_c_178_n 0.00527795f $X=1.945 $Y=1.84 $X2=0 $Y2=0
cc_123 N_VPWR_c_138_n N_Y_c_178_n 0.023803f $X=2.095 $Y=2.455 $X2=0 $Y2=0
cc_124 N_VPWR_M1007_s Y 0.0019552f $X=1.945 $Y=1.84 $X2=0 $Y2=0
cc_125 N_VPWR_c_135_n N_A_27_74#_c_226_n 0.00901952f $X=0.285 $Y=1.985 $X2=0
+ $Y2=0
cc_126 N_Y_c_173_n N_A_27_74#_M1002_s 0.00341347f $X=2.045 $Y=1.095 $X2=0 $Y2=0
cc_127 N_Y_c_174_n N_A_27_74#_c_225_n 0.00997012f $X=1.785 $Y=1.095 $X2=0 $Y2=0
cc_128 N_Y_M1000_d N_A_27_74#_c_227_n 0.00229612f $X=1.48 $Y=0.37 $X2=0 $Y2=0
cc_129 N_Y_c_189_n N_A_27_74#_c_227_n 0.0179413f $X=1.62 $Y=0.86 $X2=0 $Y2=0
cc_130 N_Y_c_173_n N_A_27_74#_c_227_n 0.00352022f $X=2.045 $Y=1.095 $X2=0 $Y2=0
cc_131 N_Y_c_173_n N_A_27_74#_c_229_n 0.0230579f $X=2.045 $Y=1.095 $X2=0 $Y2=0
cc_132 N_A_27_74#_c_225_n N_VGND_M1004_s 0.00229612f $X=1.105 $Y=1.095 $X2=-0.19
+ $Y2=-0.245
cc_133 N_A_27_74#_c_224_n N_VGND_c_258_n 0.0182902f $X=0.28 $Y=0.515 $X2=0 $Y2=0
cc_134 N_A_27_74#_c_225_n N_VGND_c_258_n 0.0194017f $X=1.105 $Y=1.095 $X2=0
+ $Y2=0
cc_135 N_A_27_74#_c_228_n N_VGND_c_258_n 0.00814404f $X=1.275 $Y=0.34 $X2=0
+ $Y2=0
cc_136 N_A_27_74#_c_224_n N_VGND_c_259_n 0.011066f $X=0.28 $Y=0.515 $X2=0 $Y2=0
cc_137 N_A_27_74#_c_227_n N_VGND_c_260_n 0.066264f $X=1.955 $Y=0.34 $X2=0 $Y2=0
cc_138 N_A_27_74#_c_228_n N_VGND_c_260_n 0.0121867f $X=1.275 $Y=0.34 $X2=0 $Y2=0
cc_139 N_A_27_74#_c_224_n N_VGND_c_261_n 0.00915947f $X=0.28 $Y=0.515 $X2=0
+ $Y2=0
cc_140 N_A_27_74#_c_227_n N_VGND_c_261_n 0.0369734f $X=1.955 $Y=0.34 $X2=0 $Y2=0
cc_141 N_A_27_74#_c_228_n N_VGND_c_261_n 0.00660921f $X=1.275 $Y=0.34 $X2=0
+ $Y2=0
