* File: sky130_fd_sc_hs__dfstp_2.pex.spice
* Created: Tue Sep  1 20:00:33 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HS__DFSTP_2%D 2 4 7 9 11 12 13 17 18 21
c34 18 0 8.44909e-20 $X=0.64 $Y=1.145
r35 21 23 39.7991 $w=3.9e-07 $l=1.65e-07 $layer=POLY_cond $X=0.61 $Y=1.825
+ $X2=0.61 $Y2=1.99
r36 21 22 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=0.64
+ $Y=1.825 $X2=0.64 $Y2=1.825
r37 17 19 45.456 $w=3.9e-07 $l=1.65e-07 $layer=POLY_cond $X=0.61 $Y=1.145
+ $X2=0.61 $Y2=0.98
r38 17 18 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=0.64
+ $Y=1.145 $X2=0.64 $Y2=1.145
r39 13 22 5.5876 $w=3.28e-07 $l=1.6e-07 $layer=LI1_cond $X=0.64 $Y=1.665
+ $X2=0.64 $Y2=1.825
r40 12 13 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=0.64 $Y=1.295
+ $X2=0.64 $Y2=1.665
r41 12 18 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=0.64 $Y=1.295
+ $X2=0.64 $Y2=1.145
r42 9 11 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=0.505 $Y=2.465
+ $X2=0.505 $Y2=2.75
r43 7 19 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=0.495 $Y=0.58 $X2=0.495
+ $Y2=0.98
r44 4 9 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=0.505 $Y=2.375 $X2=0.505
+ $Y2=2.465
r45 4 23 149.653 $w=1.8e-07 $l=3.85e-07 $layer=POLY_cond $X=0.505 $Y=2.375
+ $X2=0.505 $Y2=1.99
r46 2 21 4.27811 $w=3.9e-07 $l=3e-08 $layer=POLY_cond $X=0.61 $Y=1.795 $X2=0.61
+ $Y2=1.825
r47 1 17 4.27811 $w=3.9e-07 $l=3e-08 $layer=POLY_cond $X=0.61 $Y=1.175 $X2=0.61
+ $Y2=1.145
r48 1 2 88.4142 $w=3.9e-07 $l=6.2e-07 $layer=POLY_cond $X=0.61 $Y=1.175 $X2=0.61
+ $Y2=1.795
.ends

.subckt PM_SKY130_FD_SC_HS__DFSTP_2%CLK 1 3 4 6 7
c33 4 0 1.813e-19 $X=1.515 $Y=1.715
r34 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.465
+ $Y=1.385 $X2=1.465 $Y2=1.385
r35 7 11 6.69663 $w=3.68e-07 $l=2.15e-07 $layer=LI1_cond $X=1.68 $Y=1.365
+ $X2=1.465 $Y2=1.365
r36 4 10 67.1335 $w=2.8e-07 $l=3.54119e-07 $layer=POLY_cond $X=1.515 $Y=1.715
+ $X2=1.465 $Y2=1.385
r37 4 6 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.515 $Y=1.715
+ $X2=1.515 $Y2=2.35
r38 1 10 38.7299 $w=2.8e-07 $l=1.74714e-07 $layer=POLY_cond $X=1.485 $Y=1.22
+ $X2=1.465 $Y2=1.385
r39 1 3 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.485 $Y=1.22 $X2=1.485
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HS__DFSTP_2%A_398_74# 1 2 7 8 9 11 12 14 16 20 21 23 26
+ 30 32 33 34 35 38 45 49 50 53 54 55 57 58 59 61 63 64 65 67 68 69 73 74 82
c268 74 0 1.63034e-19 $X=6.795 $Y=1.285
c269 69 0 3.40141e-19 $X=3.77 $Y=2.325
c270 59 0 4.94485e-20 $X=5.69 $Y=2.405
c271 21 0 1.55697e-19 $X=7.53 $Y=2.465
c272 14 0 1.99877e-19 $X=3.83 $Y=1.38
c273 8 0 8.44808e-20 $X=2.95 $Y=1.885
r274 77 78 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.455
+ $Y=2.215 $X2=7.455 $Y2=2.215
r275 74 82 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.795 $Y=1.285
+ $X2=6.795 $Y2=1.12
r276 73 74 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.795
+ $Y=1.285 $X2=6.795 $Y2=1.285
r277 70 73 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=6.5 $Y=1.285
+ $X2=6.795 $Y2=1.285
r278 67 77 11.5534 $w=3.29e-07 $l=2.8058e-07 $layer=LI1_cond $X=7.575 $Y=1.98
+ $X2=7.475 $Y2=2.215
r279 66 67 99.8182 $w=1.68e-07 $l=1.53e-06 $layer=LI1_cond $X=7.575 $Y=0.45
+ $X2=7.575 $Y2=1.98
r280 64 66 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.49 $Y=0.365
+ $X2=7.575 $Y2=0.45
r281 64 65 59.0428 $w=1.68e-07 $l=9.05e-07 $layer=LI1_cond $X=7.49 $Y=0.365
+ $X2=6.585 $Y2=0.365
r282 62 70 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.5 $Y=1.45 $X2=6.5
+ $Y2=1.285
r283 62 63 56.7594 $w=1.68e-07 $l=8.7e-07 $layer=LI1_cond $X=6.5 $Y=1.45 $X2=6.5
+ $Y2=2.32
r284 61 70 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.5 $Y=1.12 $X2=6.5
+ $Y2=1.285
r285 60 65 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.5 $Y=0.45
+ $X2=6.585 $Y2=0.365
r286 60 61 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=6.5 $Y=0.45 $X2=6.5
+ $Y2=1.12
r287 58 63 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.415 $Y=2.405
+ $X2=6.5 $Y2=2.32
r288 58 59 47.2995 $w=1.68e-07 $l=7.25e-07 $layer=LI1_cond $X=6.415 $Y=2.405
+ $X2=5.69 $Y2=2.405
r289 56 59 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.605 $Y=2.49
+ $X2=5.69 $Y2=2.405
r290 56 57 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=5.605 $Y=2.49
+ $X2=5.605 $Y2=2.89
r291 54 57 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.52 $Y=2.975
+ $X2=5.605 $Y2=2.89
r292 54 55 39.4706 $w=1.68e-07 $l=6.05e-07 $layer=LI1_cond $X=5.52 $Y=2.975
+ $X2=4.915 $Y2=2.975
r293 53 55 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.83 $Y=2.89
+ $X2=4.915 $Y2=2.975
r294 52 53 31.3155 $w=1.68e-07 $l=4.8e-07 $layer=LI1_cond $X=4.83 $Y=2.41
+ $X2=4.83 $Y2=2.89
r295 51 69 2.45049 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=3.915 $Y=2.325
+ $X2=3.77 $Y2=2.325
r296 50 52 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.745 $Y=2.325
+ $X2=4.83 $Y2=2.41
r297 50 51 54.1497 $w=1.68e-07 $l=8.3e-07 $layer=LI1_cond $X=4.745 $Y=2.325
+ $X2=3.915 $Y2=2.325
r298 48 69 3.98977 $w=2.3e-07 $l=1.11018e-07 $layer=LI1_cond $X=3.71 $Y=2.41
+ $X2=3.77 $Y2=2.325
r299 48 49 31.3155 $w=1.68e-07 $l=4.8e-07 $layer=LI1_cond $X=3.71 $Y=2.41
+ $X2=3.71 $Y2=2.89
r300 45 46 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.77
+ $Y=1.545 $X2=3.77 $Y2=1.545
r301 43 69 3.98977 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.77 $Y=2.24
+ $X2=3.77 $Y2=2.325
r302 43 45 27.6189 $w=2.88e-07 $l=6.95e-07 $layer=LI1_cond $X=3.77 $Y=2.24
+ $X2=3.77 $Y2=1.545
r303 41 68 62.3048 $w=1.68e-07 $l=9.55e-07 $layer=LI1_cond $X=3.03 $Y=0.425
+ $X2=3.03 $Y2=1.38
r304 38 68 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=2.95 $Y=1.545
+ $X2=2.95 $Y2=1.38
r305 38 39 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.95
+ $Y=1.545 $X2=2.95 $Y2=1.545
r306 34 49 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.625 $Y=2.975
+ $X2=3.71 $Y2=2.89
r307 34 35 88.0749 $w=1.68e-07 $l=1.35e-06 $layer=LI1_cond $X=3.625 $Y=2.975
+ $X2=2.275 $Y2=2.975
r308 32 41 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.945 $Y=0.34
+ $X2=3.03 $Y2=0.425
r309 32 33 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=2.945 $Y=0.34
+ $X2=2.215 $Y2=0.34
r310 28 35 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.19 $Y=2.89
+ $X2=2.275 $Y2=2.975
r311 28 30 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=2.19 $Y=2.89
+ $X2=2.19 $Y2=2.665
r312 24 33 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.13 $Y=0.425
+ $X2=2.215 $Y2=0.34
r313 24 26 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=2.13 $Y=0.425
+ $X2=2.13 $Y2=0.515
r314 21 78 52.2586 $w=2.99e-07 $l=2.85044e-07 $layer=POLY_cond $X=7.53 $Y=2.465
+ $X2=7.455 $Y2=2.215
r315 21 23 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=7.53 $Y=2.465
+ $X2=7.53 $Y2=2.75
r316 20 82 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=6.705 $Y=0.69
+ $X2=6.705 $Y2=1.12
r317 14 46 21.4517 $w=1.5e-07 $l=1.72337e-07 $layer=POLY_cond $X=3.83 $Y=1.38
+ $X2=3.845 $Y2=1.545
r318 14 16 410.213 $w=1.5e-07 $l=8e-07 $layer=POLY_cond $X=3.83 $Y=1.38 $X2=3.83
+ $Y2=0.58
r319 13 39 13.4654 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.115 $Y=1.545
+ $X2=2.95 $Y2=1.545
r320 12 46 10.7258 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=3.755 $Y=1.545
+ $X2=3.845 $Y2=1.545
r321 12 13 111.911 $w=3.3e-07 $l=6.4e-07 $layer=POLY_cond $X=3.755 $Y=1.545
+ $X2=3.115 $Y2=1.545
r322 9 11 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=3.005 $Y=2.205
+ $X2=3.005 $Y2=2.49
r323 8 9 60.0156 $w=2.57e-07 $l=3.4641e-07 $layer=POLY_cond $X=2.95 $Y=1.885
+ $X2=3.005 $Y2=2.205
r324 7 39 13.4654 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.95 $Y=1.71
+ $X2=2.95 $Y2=1.545
r325 7 8 30.6007 $w=3.3e-07 $l=1.75e-07 $layer=POLY_cond $X=2.95 $Y=1.71
+ $X2=2.95 $Y2=1.885
r326 2 30 600 $w=1.7e-07 $l=9.47035e-07 $layer=licon1_PDIFF $count=1 $X=2.04
+ $Y=1.79 $X2=2.19 $Y2=2.665
r327 1 26 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.99
+ $Y=0.37 $X2=2.13 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__DFSTP_2%A_767_384# 1 2 7 9 10 12 14 17 19 22 27 32
+ 33 36 40
c84 40 0 1.05311e-20 $X=4.485 $Y=1.065
c85 7 0 1.52996e-19 $X=3.925 $Y=2.205
r86 32 33 10.1743 $w=2.63e-07 $l=2e-07 $layer=LI1_cond $X=5.217 $Y=2.52
+ $X2=5.217 $Y2=2.32
r87 28 40 17.4217 $w=2.49e-07 $l=9e-08 $layer=POLY_cond $X=4.575 $Y=1.065
+ $X2=4.485 $Y2=1.065
r88 27 30 12.2584 $w=4.18e-07 $l=4.2e-07 $layer=LI1_cond $X=4.575 $Y=0.9
+ $X2=4.995 $Y2=0.9
r89 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.575
+ $Y=1.065 $X2=4.575 $Y2=1.065
r90 24 33 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=5.17 $Y=2.07
+ $X2=5.17 $Y2=2.32
r91 22 37 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=4.395 $Y=1.905
+ $X2=4.395 $Y2=1.995
r92 22 36 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.395 $Y=1.905
+ $X2=4.395 $Y2=1.74
r93 21 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.395
+ $Y=1.905 $X2=4.395 $Y2=1.905
r94 19 24 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=5.085 $Y=1.905
+ $X2=5.17 $Y2=2.07
r95 19 21 24.0965 $w=3.28e-07 $l=6.9e-07 $layer=LI1_cond $X=5.085 $Y=1.905
+ $X2=4.395 $Y2=1.905
r96 15 40 14.627 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.485 $Y=1.23
+ $X2=4.485 $Y2=1.065
r97 15 36 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=4.485 $Y=1.23
+ $X2=4.485 $Y2=1.74
r98 12 40 51.2972 $w=2.49e-07 $l=3.37565e-07 $layer=POLY_cond $X=4.22 $Y=0.9
+ $X2=4.485 $Y2=1.065
r99 12 14 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=4.22 $Y=0.9 $X2=4.22
+ $Y2=0.58
r100 11 17 7.1379 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=4.015 $Y=1.995
+ $X2=3.925 $Y2=1.995
r101 10 37 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.23 $Y=1.995
+ $X2=4.395 $Y2=1.995
r102 10 11 110.245 $w=1.5e-07 $l=2.15e-07 $layer=POLY_cond $X=4.23 $Y=1.995
+ $X2=4.015 $Y2=1.995
r103 7 17 83.7788 $w=1.8e-07 $l=2.1e-07 $layer=POLY_cond $X=3.925 $Y=2.205
+ $X2=3.925 $Y2=1.995
r104 7 9 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=3.925 $Y=2.205
+ $X2=3.925 $Y2=2.49
r105 2 32 600 $w=1.7e-07 $l=3.05941e-07 $layer=licon1_PDIFF $count=1 $X=5.115
+ $Y=2.28 $X2=5.265 $Y2=2.52
r106 1 30 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=4.85
+ $Y=0.59 $X2=4.995 $Y2=0.8
.ends

.subckt PM_SKY130_FD_SC_HS__DFSTP_2%A_612_74# 1 2 8 9 11 14 16 18 21 25 29 32 34
+ 36 38 39 41 45 47 49 54
c132 47 0 1.63034e-19 $X=6.08 $Y=1.38
c133 39 0 1.52996e-19 $X=3.285 $Y=2.26
c134 36 0 1.05311e-20 $X=5.125 $Y=1.395
c135 32 0 1.99877e-19 $X=4.17 $Y=1.4
c136 9 0 4.94485e-20 $X=5.04 $Y=2.205
r137 47 49 5.35643 $w=3.53e-07 $l=1.65e-07 $layer=LI1_cond $X=6.08 $Y=1.392
+ $X2=5.915 $Y2=1.392
r138 47 48 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.08
+ $Y=1.38 $X2=6.08 $Y2=1.38
r139 44 54 16.6118 $w=3.3e-07 $l=9.5e-08 $layer=POLY_cond $X=5.115 $Y=1.385
+ $X2=5.21 $Y2=1.385
r140 44 51 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=5.115 $Y=1.385
+ $X2=5.04 $Y2=1.385
r141 43 45 8.48848 $w=3.48e-07 $l=1.65e-07 $layer=LI1_cond $X=5.115 $Y=1.395
+ $X2=4.95 $Y2=1.395
r142 43 44 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.115
+ $Y=1.385 $X2=5.115 $Y2=1.385
r143 38 39 10.6751 $w=3.38e-07 $l=2.3e-07 $layer=LI1_cond $X=3.285 $Y=2.49
+ $X2=3.285 $Y2=2.26
r144 36 43 0.329269 $w=3.48e-07 $l=1e-08 $layer=LI1_cond $X=5.125 $Y=1.395
+ $X2=5.115 $Y2=1.395
r145 36 49 26.0123 $w=3.48e-07 $l=7.9e-07 $layer=LI1_cond $X=5.125 $Y=1.395
+ $X2=5.915 $Y2=1.395
r146 34 45 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=4.255 $Y=1.485
+ $X2=4.95 $Y2=1.485
r147 32 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.17 $Y=1.4
+ $X2=4.255 $Y2=1.485
r148 31 32 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=4.17 $Y=1.21
+ $X2=4.17 $Y2=1.4
r149 30 41 2.76166 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.615 $Y=1.125
+ $X2=3.45 $Y2=1.125
r150 29 31 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.085 $Y=1.125
+ $X2=4.17 $Y2=1.21
r151 29 30 30.6631 $w=1.68e-07 $l=4.7e-07 $layer=LI1_cond $X=4.085 $Y=1.125
+ $X2=3.615 $Y2=1.125
r152 27 41 3.70735 $w=2.5e-07 $l=1.18427e-07 $layer=LI1_cond $X=3.37 $Y=1.21
+ $X2=3.45 $Y2=1.125
r153 27 39 68.5027 $w=1.68e-07 $l=1.05e-06 $layer=LI1_cond $X=3.37 $Y=1.21
+ $X2=3.37 $Y2=2.26
r154 23 41 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.45 $Y=1.04
+ $X2=3.45 $Y2=1.125
r155 23 25 15.8897 $w=3.28e-07 $l=4.55e-07 $layer=LI1_cond $X=3.45 $Y=1.04
+ $X2=3.45 $Y2=0.585
r156 19 48 39.8702 $w=4.14e-07 $l=2.32637e-07 $layer=POLY_cond $X=6.315 $Y=1.215
+ $X2=6.152 $Y2=1.38
r157 19 21 269.202 $w=1.5e-07 $l=5.25e-07 $layer=POLY_cond $X=6.315 $Y=1.215
+ $X2=6.315 $Y2=0.69
r158 16 48 49.7663 $w=4.14e-07 $l=2.97069e-07 $layer=POLY_cond $X=6.255 $Y=1.63
+ $X2=6.152 $Y2=1.38
r159 16 18 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=6.255 $Y=1.63
+ $X2=6.255 $Y2=2.205
r160 12 54 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.21 $Y=1.22
+ $X2=5.21 $Y2=1.385
r161 12 14 215.362 $w=1.5e-07 $l=4.2e-07 $layer=POLY_cond $X=5.21 $Y=1.22
+ $X2=5.21 $Y2=0.8
r162 9 11 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=5.04 $Y=2.205
+ $X2=5.04 $Y2=2.49
r163 8 9 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=5.04 $Y=2.115 $X2=5.04
+ $Y2=2.205
r164 7 51 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=5.04 $Y=1.55
+ $X2=5.04 $Y2=1.385
r165 7 8 219.621 $w=1.8e-07 $l=5.65e-07 $layer=POLY_cond $X=5.04 $Y=1.55
+ $X2=5.04 $Y2=2.115
r166 2 38 600 $w=1.7e-07 $l=2.93428e-07 $layer=licon1_PDIFF $count=1 $X=3.08
+ $Y=2.28 $X2=3.28 $Y2=2.49
r167 1 25 182 $w=1.7e-07 $l=4.85747e-07 $layer=licon1_NDIFF $count=1 $X=3.06
+ $Y=0.37 $X2=3.45 $Y2=0.585
.ends

.subckt PM_SKY130_FD_SC_HS__DFSTP_2%SET_B 1 3 6 10 13 14 16 19 20 21 22 25 27 30
+ 31
c124 31 0 1.62395e-19 $X=8.565 $Y=1.645
c125 13 0 6.88335e-20 $X=8.49 $Y=2.375
r126 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.59
+ $Y=1.955 $X2=5.59 $Y2=1.955
r127 31 42 10.8302 $w=4.13e-07 $l=3.9e-07 $layer=LI1_cond $X=8.522 $Y=1.645
+ $X2=8.522 $Y2=2.035
r128 30 31 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=8.565
+ $Y=1.645 $X2=8.565 $Y2=1.645
r129 27 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=2.035
+ $X2=8.4 $Y2=2.035
r130 25 34 13.125 $w=3.58e-07 $l=4.1e-07 $layer=LI1_cond $X=6 $Y=1.97 $X2=5.59
+ $Y2=1.97
r131 24 25 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=2.035 $X2=6
+ $Y2=2.035
r132 22 24 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.145 $Y=2.035
+ $X2=6 $Y2=2.035
r133 21 27 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=8.255 $Y=2.035
+ $X2=8.4 $Y2=2.035
r134 21 22 2.61138 $w=1.4e-07 $l=2.11e-06 $layer=MET1_cond $X=8.255 $Y=2.035
+ $X2=6.145 $Y2=2.035
r135 19 30 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=8.565 $Y=1.985
+ $X2=8.565 $Y2=1.645
r136 19 20 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=8.565 $Y=1.985
+ $X2=8.565 $Y2=2.15
r137 18 30 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=8.565 $Y=1.48
+ $X2=8.565 $Y2=1.645
r138 14 16 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=8.49 $Y=2.465
+ $X2=8.49 $Y2=2.75
r139 13 14 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=8.49 $Y=2.375
+ $X2=8.49 $Y2=2.465
r140 13 20 87.4597 $w=1.8e-07 $l=2.25e-07 $layer=POLY_cond $X=8.49 $Y=2.375
+ $X2=8.49 $Y2=2.15
r141 10 18 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=8.475 $Y=0.8
+ $X2=8.475 $Y2=1.48
r142 4 33 38.5462 $w=3.19e-07 $l=1.76125e-07 $layer=POLY_cond $X=5.6 $Y=1.79
+ $X2=5.577 $Y2=1.955
r143 4 6 507.638 $w=1.5e-07 $l=9.9e-07 $layer=POLY_cond $X=5.6 $Y=1.79 $X2=5.6
+ $Y2=0.8
r144 1 33 51.3895 $w=3.19e-07 $l=2.90259e-07 $layer=POLY_cond $X=5.49 $Y=2.205
+ $X2=5.577 $Y2=1.955
r145 1 3 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=5.49 $Y=2.205 $X2=5.49
+ $Y2=2.49
.ends

.subckt PM_SKY130_FD_SC_HS__DFSTP_2%A_225_74# 1 2 9 11 13 15 17 18 19 20 21 24
+ 26 27 28 30 31 36 37 38 41 45 46 47 49 50 51 54 58 62 65
c194 54 0 2.99812e-20 $X=1.945 $Y=1.805
c195 31 0 1.89865e-19 $X=6.67 $Y=3.15
c196 28 0 1.36144e-19 $X=3.505 $Y=2.775
r197 62 64 17.9907 $w=4.58e-07 $l=5e-07 $layer=LI1_cond $X=1.205 $Y=0.51
+ $X2=1.205 $Y2=1.01
r198 58 59 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.11
+ $Y=1.465 $X2=2.11 $Y2=1.465
r199 56 58 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=2.11 $Y=1.72
+ $X2=2.11 $Y2=1.465
r200 54 56 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.945 $Y=1.805
+ $X2=2.11 $Y2=1.72
r201 54 65 31.9679 $w=1.68e-07 $l=4.9e-07 $layer=LI1_cond $X=1.945 $Y=1.805
+ $X2=1.455 $Y2=1.805
r202 51 53 5.57014 $w=2.98e-07 $l=1.45e-07 $layer=LI1_cond $X=1.145 $Y=1.87
+ $X2=1.29 $Y2=1.87
r203 50 65 7.90841 $w=2.98e-07 $l=1.5e-07 $layer=LI1_cond $X=1.305 $Y=1.87
+ $X2=1.455 $Y2=1.87
r204 50 53 0.576222 $w=2.98e-07 $l=1.5e-08 $layer=LI1_cond $X=1.305 $Y=1.87
+ $X2=1.29 $Y2=1.87
r205 49 51 7.51767 $w=3e-07 $l=1.8775e-07 $layer=LI1_cond $X=1.06 $Y=1.72
+ $X2=1.145 $Y2=1.87
r206 49 64 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=1.06 $Y=1.72
+ $X2=1.06 $Y2=1.01
r207 45 59 52.4584 $w=3.3e-07 $l=3e-07 $layer=POLY_cond $X=2.41 $Y=1.465
+ $X2=2.11 $Y2=1.465
r208 45 46 5.03009 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=2.41 $Y=1.465
+ $X2=2.485 $Y2=1.465
r209 44 59 9.61737 $w=3.3e-07 $l=5.5e-08 $layer=POLY_cond $X=2.055 $Y=1.465
+ $X2=2.11 $Y2=1.465
r210 39 41 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=7.37 $Y=1.66
+ $X2=7.37 $Y2=0.8
r211 37 39 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=7.295 $Y=1.735
+ $X2=7.37 $Y2=1.66
r212 37 38 228.181 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=7.295 $Y=1.735
+ $X2=6.85 $Y2=1.735
r213 34 36 294.84 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=6.76 $Y=3.035
+ $X2=6.76 $Y2=2.46
r214 33 38 26.9307 $w=1.5e-07 $l=1.89737e-07 $layer=POLY_cond $X=6.76 $Y=1.885
+ $X2=6.85 $Y2=1.735
r215 33 36 294.84 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=6.76 $Y=1.885
+ $X2=6.76 $Y2=2.46
r216 32 47 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=3.595 $Y=3.15
+ $X2=3.505 $Y2=3.15
r217 31 34 26.9307 $w=1.5e-07 $l=1.53542e-07 $layer=POLY_cond $X=6.67 $Y=3.15
+ $X2=6.76 $Y2=3.035
r218 31 32 1576.76 $w=1.5e-07 $l=3.075e-06 $layer=POLY_cond $X=6.67 $Y=3.15
+ $X2=3.595 $Y2=3.15
r219 28 30 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=3.505 $Y=2.775
+ $X2=3.505 $Y2=2.49
r220 27 47 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=3.505 $Y=3.075
+ $X2=3.505 $Y2=3.15
r221 26 28 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=3.505 $Y=2.865
+ $X2=3.505 $Y2=2.775
r222 26 27 81.629 $w=1.8e-07 $l=2.1e-07 $layer=POLY_cond $X=3.505 $Y=2.865
+ $X2=3.505 $Y2=3.075
r223 22 24 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=2.985 $Y=0.99
+ $X2=2.985 $Y2=0.58
r224 20 47 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=3.415 $Y=3.15
+ $X2=3.505 $Y2=3.15
r225 20 21 438.415 $w=1.5e-07 $l=8.55e-07 $layer=POLY_cond $X=3.415 $Y=3.15
+ $X2=2.56 $Y2=3.15
r226 18 22 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.91 $Y=1.065
+ $X2=2.985 $Y2=0.99
r227 18 19 179.468 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=2.91 $Y=1.065
+ $X2=2.56 $Y2=1.065
r228 17 21 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.485 $Y=3.075
+ $X2=2.56 $Y2=3.15
r229 16 46 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.485 $Y=1.63
+ $X2=2.485 $Y2=1.465
r230 16 17 740.947 $w=1.5e-07 $l=1.445e-06 $layer=POLY_cond $X=2.485 $Y=1.63
+ $X2=2.485 $Y2=3.075
r231 15 46 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.485 $Y=1.3
+ $X2=2.485 $Y2=1.465
r232 14 19 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.485 $Y=1.14
+ $X2=2.56 $Y2=1.065
r233 14 15 82.0426 $w=1.5e-07 $l=1.6e-07 $layer=POLY_cond $X=2.485 $Y=1.14
+ $X2=2.485 $Y2=1.3
r234 11 44 61.9504 $w=2.07e-07 $l=2.58844e-07 $layer=POLY_cond $X=1.965 $Y=1.715
+ $X2=1.947 $Y2=1.465
r235 11 13 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.965 $Y=1.715
+ $X2=1.965 $Y2=2.35
r236 7 44 42.1581 $w=2.07e-07 $l=1.80291e-07 $layer=POLY_cond $X=1.915 $Y=1.3
+ $X2=1.947 $Y2=1.465
r237 7 9 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=1.915 $Y=1.3
+ $X2=1.915 $Y2=0.74
r238 2 53 600 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=1.145
+ $Y=1.79 $X2=1.29 $Y2=1.935
r239 1 62 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.125
+ $Y=0.37 $X2=1.27 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HS__DFSTP_2%A_1566_92# 1 2 9 11 12 14 16 19 20 23 25 26
+ 29 33 35 39
c85 19 0 1.23601e-19 $X=7.995 $Y=1.285
c86 11 0 1.62395e-19 $X=7.95 $Y=2.375
r87 31 35 3.10218 $w=3.05e-07 $l=1.09087e-07 $layer=LI1_cond $X=9.765 $Y=1.24
+ $X2=9.71 $Y2=1.155
r88 31 33 69.6076 $w=2.48e-07 $l=1.51e-06 $layer=LI1_cond $X=9.765 $Y=1.24
+ $X2=9.765 $Y2=2.75
r89 27 35 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=9.71 $Y=1.07
+ $X2=9.71 $Y2=1.155
r90 27 29 8.64332 $w=3.58e-07 $l=2.7e-07 $layer=LI1_cond $X=9.71 $Y=1.07
+ $X2=9.71 $Y2=0.8
r91 25 35 3.51065 $w=1.7e-07 $l=1.8e-07 $layer=LI1_cond $X=9.53 $Y=1.155
+ $X2=9.71 $Y2=1.155
r92 25 26 90.3583 $w=1.68e-07 $l=1.385e-06 $layer=LI1_cond $X=9.53 $Y=1.155
+ $X2=8.145 $Y2=1.155
r93 23 39 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=7.995 $Y=1.965
+ $X2=7.995 $Y2=2.13
r94 22 23 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=7.995
+ $Y=1.965 $X2=7.995 $Y2=1.965
r95 20 23 118.906 $w=3.3e-07 $l=6.8e-07 $layer=POLY_cond $X=7.995 $Y=1.285
+ $X2=7.995 $Y2=1.965
r96 19 22 24.8781 $w=3.13e-07 $l=6.8e-07 $layer=LI1_cond $X=7.987 $Y=1.285
+ $X2=7.987 $Y2=1.965
r97 19 20 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=7.995
+ $Y=1.285 $X2=7.995 $Y2=1.285
r98 17 26 7.64049 $w=1.7e-07 $l=1.95944e-07 $layer=LI1_cond $X=7.987 $Y=1.24
+ $X2=8.145 $Y2=1.155
r99 17 19 1.64635 $w=3.13e-07 $l=4.5e-08 $layer=LI1_cond $X=7.987 $Y=1.24
+ $X2=7.987 $Y2=1.285
r100 16 20 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=7.995 $Y=1.12
+ $X2=7.995 $Y2=1.285
r101 12 14 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=7.95 $Y=2.465
+ $X2=7.95 $Y2=2.75
r102 11 12 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=7.95 $Y=2.375
+ $X2=7.95 $Y2=2.465
r103 11 39 95.2339 $w=1.8e-07 $l=2.45e-07 $layer=POLY_cond $X=7.95 $Y=2.375
+ $X2=7.95 $Y2=2.13
r104 9 16 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=7.905 $Y=0.8
+ $X2=7.905 $Y2=1.12
r105 2 33 600 $w=1.7e-07 $l=2.74955e-07 $layer=licon1_PDIFF $count=1 $X=9.575
+ $Y=2.54 $X2=9.725 $Y2=2.75
r106 1 29 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=9.555
+ $Y=0.59 $X2=9.695 $Y2=0.8
.ends

.subckt PM_SKY130_FD_SC_HS__DFSTP_2%A_1356_74# 1 2 3 12 14 16 17 21 23 25 27 28
+ 29 33 35 36 38 39 42 44 48 49 53 59 63 69
c158 53 0 3.20959e-20 $X=7.235 $Y=1.705
c159 39 0 6.88335e-20 $X=7.93 $Y=2.435
c160 29 0 8.20619e-20 $X=10.497 $Y=1.69
r161 61 63 6.9845 $w=3.28e-07 $l=2e-07 $layer=LI1_cond $X=7.035 $Y=0.785
+ $X2=7.235 $Y2=0.785
r162 58 59 8.41349 $w=4.28e-07 $l=1.65e-07 $layer=LI1_cond $X=7.305 $Y=2.765
+ $X2=7.47 $Y2=2.765
r163 55 58 9.64836 $w=4.28e-07 $l=3.6e-07 $layer=LI1_cond $X=6.945 $Y=2.765
+ $X2=7.305 $Y2=2.765
r164 48 49 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=9.305
+ $Y=1.78 $X2=9.305 $Y2=1.78
r165 46 48 18.8582 $w=3.28e-07 $l=5.4e-07 $layer=LI1_cond $X=9.305 $Y=2.32
+ $X2=9.305 $Y2=1.78
r166 45 69 6.19399 $w=2e-07 $l=1.39194e-07 $layer=LI1_cond $X=8.88 $Y=2.405
+ $X2=8.755 $Y2=2.435
r167 44 46 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=9.14 $Y=2.405
+ $X2=9.305 $Y2=2.32
r168 44 45 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=9.14 $Y=2.405
+ $X2=8.88 $Y2=2.405
r169 40 69 0.552779 $w=2.5e-07 $l=1.15e-07 $layer=LI1_cond $X=8.755 $Y=2.55
+ $X2=8.755 $Y2=2.435
r170 40 42 9.21954 $w=2.48e-07 $l=2e-07 $layer=LI1_cond $X=8.755 $Y=2.55
+ $X2=8.755 $Y2=2.75
r171 39 67 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=7.845 $Y=2.435
+ $X2=7.845 $Y2=2.64
r172 38 69 6.19399 $w=2e-07 $l=1.25e-07 $layer=LI1_cond $X=8.63 $Y=2.435
+ $X2=8.755 $Y2=2.435
r173 38 39 35.0744 $w=2.28e-07 $l=7e-07 $layer=LI1_cond $X=8.63 $Y=2.435
+ $X2=7.93 $Y2=2.435
r174 36 67 0.364908 $w=1.8e-07 $l=8.5e-08 $layer=LI1_cond $X=7.76 $Y=2.64
+ $X2=7.845 $Y2=2.64
r175 36 59 17.8687 $w=1.78e-07 $l=2.9e-07 $layer=LI1_cond $X=7.76 $Y=2.64
+ $X2=7.47 $Y2=2.64
r176 35 53 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.235 $Y=1.62
+ $X2=7.235 $Y2=1.705
r177 34 63 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.235 $Y=0.95
+ $X2=7.235 $Y2=0.785
r178 34 35 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=7.235 $Y=0.95
+ $X2=7.235 $Y2=1.62
r179 31 55 3.91032 $w=2.5e-07 $l=2.15e-07 $layer=LI1_cond $X=6.945 $Y=2.55
+ $X2=6.945 $Y2=2.765
r180 31 33 18.9001 $w=2.48e-07 $l=4.1e-07 $layer=LI1_cond $X=6.945 $Y=2.55
+ $X2=6.945 $Y2=2.14
r181 30 53 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=6.945 $Y=1.705
+ $X2=7.235 $Y2=1.705
r182 30 33 16.1342 $w=2.48e-07 $l=3.5e-07 $layer=LI1_cond $X=6.945 $Y=1.79
+ $X2=6.945 $Y2=2.14
r183 28 49 34.6051 $w=4.5e-07 $l=2.8e-07 $layer=POLY_cond $X=9.365 $Y=2.06
+ $X2=9.365 $Y2=1.78
r184 26 49 1.85385 $w=4.5e-07 $l=1.5e-08 $layer=POLY_cond $X=9.365 $Y=1.765
+ $X2=9.365 $Y2=1.78
r185 26 27 11.1008 $w=3e-07 $l=7.5e-08 $layer=POLY_cond $X=9.365 $Y=1.765
+ $X2=9.365 $Y2=1.69
r186 23 29 20.4101 $w=1.5e-07 $l=8.12404e-08 $layer=POLY_cond $X=10.51 $Y=1.765
+ $X2=10.497 $Y2=1.69
r187 23 25 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=10.51 $Y=1.765
+ $X2=10.51 $Y2=2.34
r188 19 29 20.4101 $w=1.5e-07 $l=8.74643e-08 $layer=POLY_cond $X=10.47 $Y=1.615
+ $X2=10.497 $Y2=1.69
r189 19 21 423.032 $w=1.5e-07 $l=8.25e-07 $layer=POLY_cond $X=10.47 $Y=1.615
+ $X2=10.47 $Y2=0.79
r190 18 27 15.4994 $w=1.5e-07 $l=2.25e-07 $layer=POLY_cond $X=9.59 $Y=1.69
+ $X2=9.365 $Y2=1.69
r191 17 29 5.30422 $w=1.5e-07 $l=1.02e-07 $layer=POLY_cond $X=10.395 $Y=1.69
+ $X2=10.497 $Y2=1.69
r192 17 18 412.777 $w=1.5e-07 $l=8.05e-07 $layer=POLY_cond $X=10.395 $Y=1.69
+ $X2=9.59 $Y2=1.69
r193 14 28 59.1545 $w=3.3e-07 $l=4.67654e-07 $layer=POLY_cond $X=9.5 $Y=2.465
+ $X2=9.365 $Y2=2.06
r194 14 16 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=9.5 $Y=2.465 $X2=9.5
+ $Y2=2.75
r195 10 27 11.1008 $w=3e-07 $l=1.47817e-07 $layer=POLY_cond $X=9.48 $Y=1.615
+ $X2=9.365 $Y2=1.69
r196 10 12 417.904 $w=1.5e-07 $l=8.15e-07 $layer=POLY_cond $X=9.48 $Y=1.615
+ $X2=9.48 $Y2=0.8
r197 3 42 600 $w=1.7e-07 $l=2.74955e-07 $layer=licon1_PDIFF $count=1 $X=8.565
+ $Y=2.54 $X2=8.715 $Y2=2.75
r198 2 58 600 $w=1.7e-07 $l=1.06437e-06 $layer=licon1_PDIFF $count=1 $X=6.835
+ $Y=1.96 $X2=7.305 $Y2=2.815
r199 2 33 300 $w=1.7e-07 $l=2.43721e-07 $layer=licon1_PDIFF $count=2 $X=6.835
+ $Y=1.96 $X2=6.985 $Y2=2.14
r200 1 61 182 $w=1.7e-07 $l=5.27304e-07 $layer=licon1_NDIFF $count=1 $X=6.78
+ $Y=0.37 $X2=7.035 $Y2=0.785
.ends

.subckt PM_SKY130_FD_SC_HS__DFSTP_2%A_2022_94# 1 2 7 9 12 16 18 20 23 27 33 36
+ 40
c68 36 0 7.76856e-20 $X=10.27 $Y=1.465
c69 7 0 1.00299e-19 $X=11.045 $Y=1.765
r70 40 41 1.84439 $w=3.92e-07 $l=1.5e-08 $layer=POLY_cond $X=11.48 $Y=1.532
+ $X2=11.495 $Y2=1.532
r71 39 40 52.8724 $w=3.92e-07 $l=4.3e-07 $layer=POLY_cond $X=11.05 $Y=1.532
+ $X2=11.48 $Y2=1.532
r72 38 39 0.614796 $w=3.92e-07 $l=5e-09 $layer=POLY_cond $X=11.045 $Y=1.532
+ $X2=11.05 $Y2=1.532
r73 34 38 8.60714 $w=3.92e-07 $l=7e-08 $layer=POLY_cond $X=10.975 $Y=1.532
+ $X2=11.045 $Y2=1.532
r74 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.975
+ $Y=1.465 $X2=10.975 $Y2=1.465
r75 31 36 1.50311 $w=3.3e-07 $l=1.8e-07 $layer=LI1_cond $X=10.45 $Y=1.465
+ $X2=10.27 $Y2=1.465
r76 31 33 18.3343 $w=3.28e-07 $l=5.25e-07 $layer=LI1_cond $X=10.45 $Y=1.465
+ $X2=10.975 $Y2=1.465
r77 27 29 22.7287 $w=3.58e-07 $l=7.1e-07 $layer=LI1_cond $X=10.27 $Y=1.985
+ $X2=10.27 $Y2=2.695
r78 25 36 4.97762 $w=3.45e-07 $l=1.65e-07 $layer=LI1_cond $X=10.27 $Y=1.63
+ $X2=10.27 $Y2=1.465
r79 25 27 11.3644 $w=3.58e-07 $l=3.55e-07 $layer=LI1_cond $X=10.27 $Y=1.63
+ $X2=10.27 $Y2=1.985
r80 21 36 4.97762 $w=3.45e-07 $l=1.72337e-07 $layer=LI1_cond $X=10.255 $Y=1.3
+ $X2=10.27 $Y2=1.465
r81 21 23 23.9219 $w=3.28e-07 $l=6.85e-07 $layer=LI1_cond $X=10.255 $Y=1.3
+ $X2=10.255 $Y2=0.615
r82 18 41 25.3688 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=11.495 $Y=1.765
+ $X2=11.495 $Y2=1.532
r83 18 20 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=11.495 $Y=1.765
+ $X2=11.495 $Y2=2.4
r84 14 40 25.3688 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=11.48 $Y=1.3
+ $X2=11.48 $Y2=1.532
r85 14 16 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=11.48 $Y=1.3
+ $X2=11.48 $Y2=0.74
r86 10 39 25.3688 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=11.05 $Y=1.3
+ $X2=11.05 $Y2=1.532
r87 10 12 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=11.05 $Y=1.3
+ $X2=11.05 $Y2=0.74
r88 7 38 25.3688 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=11.045 $Y=1.765
+ $X2=11.045 $Y2=1.532
r89 7 9 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=11.045 $Y=1.765
+ $X2=11.045 $Y2=2.4
r90 2 29 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=10.14
+ $Y=1.84 $X2=10.285 $Y2=2.695
r91 2 27 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=10.14
+ $Y=1.84 $X2=10.285 $Y2=1.985
r92 1 23 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=10.11
+ $Y=0.47 $X2=10.255 $Y2=0.615
.ends

.subckt PM_SKY130_FD_SC_HS__DFSTP_2%A_27_74# 1 2 3 4 14 17 19 21 24 26 29 30 37
c71 24 0 8.44808e-20 $X=2.53 $Y=2.06
c72 21 0 1.36144e-19 $X=2.445 $Y=2.145
r73 34 37 5.5876 $w=3.28e-07 $l=1.6e-07 $layer=LI1_cond $X=2.53 $Y=0.76 $X2=2.69
+ $Y2=0.76
r74 30 32 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=1.71 $Y=2.145
+ $X2=1.71 $Y2=2.275
r75 26 28 9.71523 $w=2.48e-07 $l=1.85e-07 $layer=LI1_cond $X=0.24 $Y=0.58
+ $X2=0.24 $Y2=0.765
r76 23 34 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.53 $Y=0.925
+ $X2=2.53 $Y2=0.76
r77 23 24 74.0481 $w=1.68e-07 $l=1.135e-06 $layer=LI1_cond $X=2.53 $Y=0.925
+ $X2=2.53 $Y2=2.06
r78 22 30 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.795 $Y=2.145
+ $X2=1.71 $Y2=2.145
r79 21 41 10.5225 $w=4e-07 $l=4.53073e-07 $layer=LI1_cond $X=2.445 $Y=2.145
+ $X2=2.695 $Y2=2.49
r80 21 24 6.71454 $w=4e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.445 $Y=2.145
+ $X2=2.53 $Y2=2.06
r81 21 22 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=2.445 $Y=2.145
+ $X2=1.795 $Y2=2.145
r82 20 29 2.11342 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.365 $Y=2.275
+ $X2=0.24 $Y2=2.275
r83 19 32 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.625 $Y=2.275
+ $X2=1.71 $Y2=2.275
r84 19 20 82.2032 $w=1.68e-07 $l=1.26e-06 $layer=LI1_cond $X=1.625 $Y=2.275
+ $X2=0.365 $Y2=2.275
r85 15 29 4.3182 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=0.24 $Y=2.36 $X2=0.24
+ $Y2=2.275
r86 15 17 17.9781 $w=2.48e-07 $l=3.9e-07 $layer=LI1_cond $X=0.24 $Y=2.36
+ $X2=0.24 $Y2=2.75
r87 14 29 4.3182 $w=2.1e-07 $l=1.03078e-07 $layer=LI1_cond $X=0.2 $Y=2.19
+ $X2=0.24 $Y2=2.275
r88 14 28 92.9679 $w=1.68e-07 $l=1.425e-06 $layer=LI1_cond $X=0.2 $Y=2.19
+ $X2=0.2 $Y2=0.765
r89 4 41 600 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_PDIFF $count=1 $X=2.635
+ $Y=2.28 $X2=2.78 $Y2=2.49
r90 3 17 600 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.54 $X2=0.28 $Y2=2.75
r91 2 37 182 $w=1.7e-07 $l=4.56782e-07 $layer=licon1_NDIFF $count=1 $X=2.545
+ $Y=0.37 $X2=2.69 $Y2=0.76
r92 1 26 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_HS__DFSTP_2%VPWR 1 2 3 4 5 6 7 8 27 31 34 37 41 45 49 53
+ 55 62 65 66 67 69 74 79 84 99 103 108 114 117 120 123 126 129 133
c149 31 0 2.99812e-20 $X=1.74 $Y=2.73
r150 132 133 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.76 $Y=3.33
+ $X2=11.76 $Y2=3.33
r151 129 130 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.8 $Y=3.33
+ $X2=10.8 $Y2=3.33
r152 126 127 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=9.36 $Y=3.33
+ $X2=9.36 $Y2=3.33
r153 120 121 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r154 117 118 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r155 114 115 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r156 112 133 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.28 $Y=3.33
+ $X2=11.76 $Y2=3.33
r157 112 130 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.28 $Y=3.33
+ $X2=10.8 $Y2=3.33
r158 111 112 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.28 $Y=3.33
+ $X2=11.28 $Y2=3.33
r159 109 129 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.985 $Y=3.33
+ $X2=10.82 $Y2=3.33
r160 109 111 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=10.985 $Y=3.33
+ $X2=11.28 $Y2=3.33
r161 108 132 4.01252 $w=1.7e-07 $l=1.82e-07 $layer=LI1_cond $X=11.635 $Y=3.33
+ $X2=11.817 $Y2=3.33
r162 108 111 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=11.635 $Y=3.33
+ $X2=11.28 $Y2=3.33
r163 107 130 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.32 $Y=3.33
+ $X2=10.8 $Y2=3.33
r164 107 127 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=10.32 $Y=3.33
+ $X2=9.36 $Y2=3.33
r165 106 107 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=10.32 $Y=3.33
+ $X2=10.32 $Y2=3.33
r166 104 126 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.44 $Y=3.33
+ $X2=9.275 $Y2=3.33
r167 104 106 57.4118 $w=1.68e-07 $l=8.8e-07 $layer=LI1_cond $X=9.44 $Y=3.33
+ $X2=10.32 $Y2=3.33
r168 103 129 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.655 $Y=3.33
+ $X2=10.82 $Y2=3.33
r169 103 106 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=10.655 $Y=3.33
+ $X2=10.32 $Y2=3.33
r170 102 127 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=3.33
+ $X2=9.36 $Y2=3.33
r171 101 102 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r172 99 126 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.11 $Y=3.33
+ $X2=9.275 $Y2=3.33
r173 99 101 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=9.11 $Y=3.33
+ $X2=8.88 $Y2=3.33
r174 98 102 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=7.92 $Y=3.33
+ $X2=8.88 $Y2=3.33
r175 97 98 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r176 95 98 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=7.92 $Y2=3.33
r177 94 97 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=6.48 $Y=3.33
+ $X2=7.92 $Y2=3.33
r178 94 95 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r179 92 123 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.11 $Y=3.33
+ $X2=5.985 $Y2=3.33
r180 92 94 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=6.11 $Y=3.33
+ $X2=6.48 $Y2=3.33
r181 90 91 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r182 88 91 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=5.52 $Y2=3.33
r183 88 121 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=4.08 $Y2=3.33
r184 87 90 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=4.56 $Y=3.33
+ $X2=5.52 $Y2=3.33
r185 87 88 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r186 85 120 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.24 $Y=3.33
+ $X2=4.155 $Y2=3.33
r187 85 87 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=4.24 $Y=3.33
+ $X2=4.56 $Y2=3.33
r188 84 123 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.86 $Y=3.33
+ $X2=5.985 $Y2=3.33
r189 84 90 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=5.86 $Y=3.33
+ $X2=5.52 $Y2=3.33
r190 83 121 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=4.08 $Y2=3.33
r191 83 118 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.68 $Y2=3.33
r192 82 83 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r193 80 117 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.905 $Y=3.33
+ $X2=1.74 $Y2=3.33
r194 80 82 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=1.905 $Y=3.33
+ $X2=2.16 $Y2=3.33
r195 79 120 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.07 $Y=3.33
+ $X2=4.155 $Y2=3.33
r196 79 82 124.61 $w=1.68e-07 $l=1.91e-06 $layer=LI1_cond $X=4.07 $Y=3.33
+ $X2=2.16 $Y2=3.33
r197 78 118 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=1.68 $Y2=3.33
r198 78 115 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r199 77 78 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r200 75 114 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.895 $Y=3.33
+ $X2=0.73 $Y2=3.33
r201 75 77 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.895 $Y=3.33
+ $X2=1.2 $Y2=3.33
r202 74 117 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.575 $Y=3.33
+ $X2=1.74 $Y2=3.33
r203 74 77 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=1.575 $Y=3.33
+ $X2=1.2 $Y2=3.33
r204 72 115 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r205 71 72 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r206 69 114 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.565 $Y=3.33
+ $X2=0.73 $Y2=3.33
r207 69 71 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.565 $Y=3.33
+ $X2=0.24 $Y2=3.33
r208 67 95 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=3.33 $X2=6.48
+ $Y2=3.33
r209 67 91 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=3.33 $X2=5.52
+ $Y2=3.33
r210 67 123 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r211 65 97 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=8.1 $Y=3.33
+ $X2=7.92 $Y2=3.33
r212 65 66 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.1 $Y=3.33
+ $X2=8.265 $Y2=3.33
r213 64 101 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=8.43 $Y=3.33
+ $X2=8.88 $Y2=3.33
r214 64 66 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.43 $Y=3.33
+ $X2=8.265 $Y2=3.33
r215 59 62 5.76222 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=4.155 $Y=2.745
+ $X2=4.32 $Y2=2.745
r216 55 58 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=11.76 $Y=1.985
+ $X2=11.76 $Y2=2.815
r217 53 132 3.13065 $w=2.5e-07 $l=1.09864e-07 $layer=LI1_cond $X=11.76 $Y=3.245
+ $X2=11.817 $Y2=3.33
r218 53 58 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=11.76 $Y=3.245
+ $X2=11.76 $Y2=2.815
r219 49 52 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=10.82 $Y=2.405
+ $X2=10.82 $Y2=2.815
r220 47 129 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=10.82 $Y=3.245
+ $X2=10.82 $Y2=3.33
r221 47 52 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=10.82 $Y=3.245
+ $X2=10.82 $Y2=2.815
r222 43 126 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.275 $Y=3.245
+ $X2=9.275 $Y2=3.33
r223 43 45 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=9.275 $Y=3.245
+ $X2=9.275 $Y2=2.78
r224 39 66 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.265 $Y=3.245
+ $X2=8.265 $Y2=3.33
r225 39 41 15.1913 $w=3.28e-07 $l=4.35e-07 $layer=LI1_cond $X=8.265 $Y=3.245
+ $X2=8.265 $Y2=2.81
r226 35 123 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.985 $Y=3.245
+ $X2=5.985 $Y2=3.33
r227 35 37 19.361 $w=2.48e-07 $l=4.2e-07 $layer=LI1_cond $X=5.985 $Y=3.245
+ $X2=5.985 $Y2=2.825
r228 34 120 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.155 $Y=3.245
+ $X2=4.155 $Y2=3.33
r229 33 59 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.155 $Y=2.91
+ $X2=4.155 $Y2=2.745
r230 33 34 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=4.155 $Y=2.91
+ $X2=4.155 $Y2=3.245
r231 29 117 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.74 $Y=3.245
+ $X2=1.74 $Y2=3.33
r232 29 31 17.9851 $w=3.28e-07 $l=5.15e-07 $layer=LI1_cond $X=1.74 $Y=3.245
+ $X2=1.74 $Y2=2.73
r233 25 114 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.73 $Y=3.245
+ $X2=0.73 $Y2=3.33
r234 25 27 17.112 $w=3.28e-07 $l=4.9e-07 $layer=LI1_cond $X=0.73 $Y=3.245
+ $X2=0.73 $Y2=2.755
r235 8 58 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=11.57
+ $Y=1.84 $X2=11.72 $Y2=2.815
r236 8 55 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=11.57
+ $Y=1.84 $X2=11.72 $Y2=1.985
r237 7 52 600 $w=1.7e-07 $l=1.08616e-06 $layer=licon1_PDIFF $count=1 $X=10.585
+ $Y=1.84 $X2=10.82 $Y2=2.815
r238 7 49 600 $w=1.7e-07 $l=6.72309e-07 $layer=licon1_PDIFF $count=1 $X=10.585
+ $Y=1.84 $X2=10.82 $Y2=2.405
r239 6 45 600 $w=1.7e-07 $l=3.03974e-07 $layer=licon1_PDIFF $count=1 $X=9.13
+ $Y=2.54 $X2=9.275 $Y2=2.78
r240 5 41 600 $w=1.7e-07 $l=3.71079e-07 $layer=licon1_PDIFF $count=1 $X=8.025
+ $Y=2.54 $X2=8.265 $Y2=2.81
r241 4 37 600 $w=1.7e-07 $l=7.10018e-07 $layer=licon1_PDIFF $count=1 $X=5.565
+ $Y=2.28 $X2=5.945 $Y2=2.825
r242 3 62 600 $w=1.7e-07 $l=6.04173e-07 $layer=licon1_PDIFF $count=1 $X=4
+ $Y=2.28 $X2=4.32 $Y2=2.745
r243 2 31 600 $w=1.7e-07 $l=1.01223e-06 $layer=licon1_PDIFF $count=1 $X=1.59
+ $Y=1.79 $X2=1.74 $Y2=2.73
r244 1 27 600 $w=1.7e-07 $l=2.80134e-07 $layer=licon1_PDIFF $count=1 $X=0.58
+ $Y=2.54 $X2=0.73 $Y2=2.755
.ends

.subckt PM_SKY130_FD_SC_HS__DFSTP_2%Q 1 2 9 13 16 17 18 19 22
c38 16 0 1.04675e-19 $X=11.38 $Y=1.82
r39 19 22 0.225187 $w=3.3e-07 $l=1.55e-07 $layer=LI1_cond $X=11.31 $Y=1.985
+ $X2=11.155 $Y2=1.985
r40 18 22 12.3975 $w=3.28e-07 $l=3.55e-07 $layer=LI1_cond $X=10.8 $Y=1.985
+ $X2=11.155 $Y2=1.985
r41 16 19 6.67463 $w=2.4e-07 $l=1.96914e-07 $layer=LI1_cond $X=11.38 $Y=1.82
+ $X2=11.31 $Y2=1.985
r42 16 17 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=11.38 $Y=1.82
+ $X2=11.38 $Y2=1.13
r43 11 19 6.67463 $w=2.4e-07 $l=1.65e-07 $layer=LI1_cond $X=11.31 $Y=2.15
+ $X2=11.31 $Y2=1.985
r44 11 13 9.29389 $w=3.08e-07 $l=2.5e-07 $layer=LI1_cond $X=11.31 $Y=2.15
+ $X2=11.31 $Y2=2.4
r45 7 17 9.06106 $w=3.63e-07 $l=1.82e-07 $layer=LI1_cond $X=11.282 $Y=0.948
+ $X2=11.282 $Y2=1.13
r46 7 9 13.6714 $w=3.63e-07 $l=4.33e-07 $layer=LI1_cond $X=11.282 $Y=0.948
+ $X2=11.282 $Y2=0.515
r47 2 19 600 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=11.12
+ $Y=1.84 $X2=11.27 $Y2=1.985
r48 2 13 300 $w=1.7e-07 $l=6.30555e-07 $layer=licon1_PDIFF $count=2 $X=11.12
+ $Y=1.84 $X2=11.27 $Y2=2.4
r49 1 9 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=11.125
+ $Y=0.37 $X2=11.265 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__DFSTP_2%VGND 1 2 3 4 5 6 7 24 26 30 34 38 42 46 48
+ 50 52 57 65 70 78 86 92 95 98 101 111 115
c110 30 0 9.68091e-20 $X=1.7 $Y=0.495
r111 114 115 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.76 $Y=0
+ $X2=11.76 $Y2=0
r112 111 112 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.8 $Y=0
+ $X2=10.8 $Y2=0
r113 98 99 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r114 95 96 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r115 93 96 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r116 92 93 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r117 90 115 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.28 $Y=0
+ $X2=11.76 $Y2=0
r118 90 112 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.28 $Y=0
+ $X2=10.8 $Y2=0
r119 89 90 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.28 $Y=0
+ $X2=11.28 $Y2=0
r120 87 111 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.93 $Y=0
+ $X2=10.765 $Y2=0
r121 87 89 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=10.93 $Y=0
+ $X2=11.28 $Y2=0
r122 86 114 4.01252 $w=1.7e-07 $l=1.82e-07 $layer=LI1_cond $X=11.635 $Y=0
+ $X2=11.817 $Y2=0
r123 86 89 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=11.635 $Y=0
+ $X2=11.28 $Y2=0
r124 85 112 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.32 $Y=0
+ $X2=10.8 $Y2=0
r125 84 85 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=10.32 $Y=0
+ $X2=10.32 $Y2=0
r126 82 85 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=9.36 $Y=0
+ $X2=10.32 $Y2=0
r127 82 106 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.36 $Y=0
+ $X2=8.88 $Y2=0
r128 81 84 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=9.36 $Y=0 $X2=10.32
+ $Y2=0
r129 81 82 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=9.36 $Y=0 $X2=9.36
+ $Y2=0
r130 78 111 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.6 $Y=0
+ $X2=10.765 $Y2=0
r131 78 84 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=10.6 $Y=0 $X2=10.32
+ $Y2=0
r132 77 106 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=0 $X2=8.88
+ $Y2=0
r133 76 77 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r134 74 77 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=6.48 $Y=0 $X2=8.4
+ $Y2=0
r135 73 76 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=6.48 $Y=0 $X2=8.4
+ $Y2=0
r136 73 74 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6.48 $Y=0
+ $X2=6.48 $Y2=0
r137 71 101 12.4999 $w=1.7e-07 $l=2.98e-07 $layer=LI1_cond $X=6.245 $Y=0
+ $X2=5.947 $Y2=0
r138 71 73 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=6.245 $Y=0
+ $X2=6.48 $Y2=0
r139 70 108 10.5284 $w=8.33e-07 $l=7.35e-07 $layer=LI1_cond $X=8.942 $Y=0
+ $X2=8.942 $Y2=0.735
r140 70 81 10.4966 $w=1.7e-07 $l=4.18e-07 $layer=LI1_cond $X=8.942 $Y=0 $X2=9.36
+ $Y2=0
r141 70 106 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=0 $X2=8.88
+ $Y2=0
r142 70 76 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=8.525 $Y=0 $X2=8.4
+ $Y2=0
r143 69 99 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=4.56
+ $Y2=0
r144 68 69 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r145 66 98 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.6 $Y=0 $X2=4.435
+ $Y2=0
r146 66 68 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=4.6 $Y=0 $X2=5.52
+ $Y2=0
r147 65 101 12.4999 $w=1.7e-07 $l=2.97e-07 $layer=LI1_cond $X=5.65 $Y=0
+ $X2=5.947 $Y2=0
r148 65 68 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=5.65 $Y=0 $X2=5.52
+ $Y2=0
r149 64 99 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=4.56
+ $Y2=0
r150 63 64 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.08 $Y=0
+ $X2=4.08 $Y2=0
r151 61 64 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=2.16 $Y=0
+ $X2=4.08 $Y2=0
r152 61 96 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.68
+ $Y2=0
r153 60 63 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=2.16 $Y=0 $X2=4.08
+ $Y2=0
r154 60 61 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.16 $Y=0
+ $X2=2.16 $Y2=0
r155 58 95 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.865 $Y=0 $X2=1.74
+ $Y2=0
r156 58 60 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=1.865 $Y=0 $X2=2.16
+ $Y2=0
r157 57 98 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.27 $Y=0 $X2=4.435
+ $Y2=0
r158 57 63 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=4.27 $Y=0 $X2=4.08
+ $Y2=0
r159 55 93 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r160 54 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r161 52 92 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.545 $Y=0 $X2=0.67
+ $Y2=0
r162 52 54 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.545 $Y=0
+ $X2=0.24 $Y2=0
r163 50 74 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=0 $X2=6.48
+ $Y2=0
r164 50 69 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=0 $X2=5.52
+ $Y2=0
r165 50 101 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=0 $X2=6 $Y2=0
r166 46 114 3.13065 $w=2.5e-07 $l=1.09864e-07 $layer=LI1_cond $X=11.76 $Y=0.085
+ $X2=11.817 $Y2=0
r167 46 48 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=11.76 $Y=0.085
+ $X2=11.76 $Y2=0.515
r168 42 44 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=10.765 $Y=0.515
+ $X2=10.765 $Y2=0.965
r169 40 111 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=10.765 $Y=0.085
+ $X2=10.765 $Y2=0
r170 40 42 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=10.765 $Y=0.085
+ $X2=10.765 $Y2=0.515
r171 36 101 2.50116 $w=5.95e-07 $l=8.5e-08 $layer=LI1_cond $X=5.947 $Y=0.085
+ $X2=5.947 $Y2=0
r172 36 38 8.64393 $w=5.93e-07 $l=4.3e-07 $layer=LI1_cond $X=5.947 $Y=0.085
+ $X2=5.947 $Y2=0.515
r173 32 98 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.435 $Y=0.085
+ $X2=4.435 $Y2=0
r174 32 34 15.5405 $w=3.28e-07 $l=4.45e-07 $layer=LI1_cond $X=4.435 $Y=0.085
+ $X2=4.435 $Y2=0.53
r175 28 95 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.74 $Y=0.085
+ $X2=1.74 $Y2=0
r176 28 30 18.9001 $w=2.48e-07 $l=4.1e-07 $layer=LI1_cond $X=1.74 $Y=0.085
+ $X2=1.74 $Y2=0.495
r177 27 92 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.795 $Y=0 $X2=0.67
+ $Y2=0
r178 26 95 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.615 $Y=0 $X2=1.74
+ $Y2=0
r179 26 27 53.4973 $w=1.68e-07 $l=8.2e-07 $layer=LI1_cond $X=1.615 $Y=0
+ $X2=0.795 $Y2=0
r180 22 92 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.67 $Y=0.085
+ $X2=0.67 $Y2=0
r181 22 24 22.8184 $w=2.48e-07 $l=4.95e-07 $layer=LI1_cond $X=0.67 $Y=0.085
+ $X2=0.67 $Y2=0.58
r182 7 48 91 $w=1.7e-07 $l=2.26164e-07 $layer=licon1_NDIFF $count=2 $X=11.555
+ $Y=0.37 $X2=11.72 $Y2=0.515
r183 6 44 182 $w=1.7e-07 $l=5.94916e-07 $layer=licon1_NDIFF $count=1 $X=10.545
+ $Y=0.47 $X2=10.765 $Y2=0.965
r184 6 42 182 $w=1.7e-07 $l=2.41454e-07 $layer=licon1_NDIFF $count=1 $X=10.545
+ $Y=0.47 $X2=10.765 $Y2=0.515
r185 5 108 91 $w=1.7e-07 $l=7.13828e-07 $layer=licon1_NDIFF $count=2 $X=8.55
+ $Y=0.59 $X2=9.195 $Y2=0.735
r186 4 38 91 $w=1.7e-07 $l=4.40908e-07 $layer=licon1_NDIFF $count=2 $X=5.675
+ $Y=0.59 $X2=6.08 $Y2=0.515
r187 3 34 182 $w=1.7e-07 $l=2.19089e-07 $layer=licon1_NDIFF $count=1 $X=4.295
+ $Y=0.37 $X2=4.435 $Y2=0.53
r188 2 30 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=1.56
+ $Y=0.37 $X2=1.7 $Y2=0.495
r189 1 24 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.37 $X2=0.71 $Y2=0.58
.ends

