* File: sky130_fd_sc_hs__dfrtp_2.pxi.spice
* Created: Tue Sep  1 20:00:03 2020
* 
x_PM_SKY130_FD_SC_HS__DFRTP_2%D N_D_c_243_n N_D_c_248_n N_D_c_249_n N_D_M1016_g
+ N_D_M1030_g D D D N_D_c_245_n N_D_c_246_n N_D_c_251_n
+ PM_SKY130_FD_SC_HS__DFRTP_2%D
x_PM_SKY130_FD_SC_HS__DFRTP_2%RESET_B N_RESET_B_M1018_g N_RESET_B_c_278_n
+ N_RESET_B_c_286_n N_RESET_B_c_287_n N_RESET_B_M1017_g N_RESET_B_c_279_n
+ N_RESET_B_M1001_g N_RESET_B_c_280_n N_RESET_B_c_289_n N_RESET_B_M1020_g
+ N_RESET_B_c_290_n N_RESET_B_M1009_g N_RESET_B_M1023_g N_RESET_B_c_282_n
+ N_RESET_B_c_292_n N_RESET_B_c_293_n N_RESET_B_c_294_n N_RESET_B_c_295_n
+ N_RESET_B_c_296_n N_RESET_B_c_297_n RESET_B N_RESET_B_c_283_n
+ N_RESET_B_c_284_n N_RESET_B_c_299_n N_RESET_B_c_300_n
+ PM_SKY130_FD_SC_HS__DFRTP_2%RESET_B
x_PM_SKY130_FD_SC_HS__DFRTP_2%CLK N_CLK_M1000_g N_CLK_c_468_n N_CLK_M1007_g CLK
+ PM_SKY130_FD_SC_HS__DFRTP_2%CLK
x_PM_SKY130_FD_SC_HS__DFRTP_2%A_490_362# N_A_490_362#_M1019_d
+ N_A_490_362#_M1012_d N_A_490_362#_c_526_n N_A_490_362#_c_527_n
+ N_A_490_362#_M1005_g N_A_490_362#_c_528_n N_A_490_362#_c_510_n
+ N_A_490_362#_M1028_g N_A_490_362#_c_512_n N_A_490_362#_M1003_g
+ N_A_490_362#_c_513_n N_A_490_362#_c_514_n N_A_490_362#_c_530_n
+ N_A_490_362#_M1026_g N_A_490_362#_c_515_n N_A_490_362#_c_516_n
+ N_A_490_362#_c_532_n N_A_490_362#_c_533_n N_A_490_362#_c_517_n
+ N_A_490_362#_c_543_n N_A_490_362#_c_518_n N_A_490_362#_c_519_n
+ N_A_490_362#_c_520_n N_A_490_362#_c_535_n N_A_490_362#_c_521_n
+ N_A_490_362#_c_522_n N_A_490_362#_c_523_n N_A_490_362#_c_524_n
+ N_A_490_362#_c_525_n N_A_490_362#_c_536_n
+ PM_SKY130_FD_SC_HS__DFRTP_2%A_490_362#
x_PM_SKY130_FD_SC_HS__DFRTP_2%A_837_359# N_A_837_359#_M1025_d
+ N_A_837_359#_M1013_d N_A_837_359#_c_708_n N_A_837_359#_M1027_g
+ N_A_837_359#_M1015_g N_A_837_359#_c_704_n N_A_837_359#_c_705_n
+ N_A_837_359#_c_734_n N_A_837_359#_c_736_n N_A_837_359#_c_711_n
+ N_A_837_359#_c_706_n N_A_837_359#_c_707_n
+ PM_SKY130_FD_SC_HS__DFRTP_2%A_837_359#
x_PM_SKY130_FD_SC_HS__DFRTP_2%A_696_457# N_A_696_457#_M1029_d
+ N_A_696_457#_M1005_d N_A_696_457#_M1020_d N_A_696_457#_M1025_g
+ N_A_696_457#_c_786_n N_A_696_457#_M1013_g N_A_696_457#_c_787_n
+ N_A_696_457#_c_788_n N_A_696_457#_c_803_n N_A_696_457#_c_795_n
+ N_A_696_457#_c_796_n N_A_696_457#_c_789_n N_A_696_457#_c_790_n
+ N_A_696_457#_c_798_n N_A_696_457#_c_791_n N_A_696_457#_c_858_n
+ PM_SKY130_FD_SC_HS__DFRTP_2%A_696_457#
x_PM_SKY130_FD_SC_HS__DFRTP_2%A_306_74# N_A_306_74#_M1000_s N_A_306_74#_M1007_s
+ N_A_306_74#_c_918_n N_A_306_74#_M1012_g N_A_306_74#_c_906_n
+ N_A_306_74#_M1019_g N_A_306_74#_c_907_n N_A_306_74#_c_919_n
+ N_A_306_74#_c_920_n N_A_306_74#_c_921_n N_A_306_74#_c_908_n
+ N_A_306_74#_M1029_g N_A_306_74#_c_922_n N_A_306_74#_c_923_n
+ N_A_306_74#_c_924_n N_A_306_74#_M1008_g N_A_306_74#_c_925_n
+ N_A_306_74#_M1021_g N_A_306_74#_c_909_n N_A_306_74#_c_928_n
+ N_A_306_74#_M1032_g N_A_306_74#_c_911_n N_A_306_74#_c_929_n
+ N_A_306_74#_c_930_n N_A_306_74#_c_931_n N_A_306_74#_c_912_n
+ N_A_306_74#_c_913_n N_A_306_74#_c_914_n N_A_306_74#_c_915_n
+ N_A_306_74#_c_916_n N_A_306_74#_c_917_n N_A_306_74#_c_934_n
+ PM_SKY130_FD_SC_HS__DFRTP_2%A_306_74#
x_PM_SKY130_FD_SC_HS__DFRTP_2%A_1525_212# N_A_1525_212#_M1024_d
+ N_A_1525_212#_M1009_d N_A_1525_212#_M1010_g N_A_1525_212#_c_1097_n
+ N_A_1525_212#_c_1098_n N_A_1525_212#_c_1099_n N_A_1525_212#_M1011_g
+ N_A_1525_212#_c_1089_n N_A_1525_212#_c_1090_n N_A_1525_212#_c_1101_n
+ N_A_1525_212#_c_1091_n N_A_1525_212#_c_1102_n N_A_1525_212#_c_1103_n
+ N_A_1525_212#_c_1104_n N_A_1525_212#_c_1092_n N_A_1525_212#_c_1093_n
+ N_A_1525_212#_c_1094_n N_A_1525_212#_c_1095_n N_A_1525_212#_c_1096_n
+ PM_SKY130_FD_SC_HS__DFRTP_2%A_1525_212#
x_PM_SKY130_FD_SC_HS__DFRTP_2%A_1271_74# N_A_1271_74#_M1003_d
+ N_A_1271_74#_M1021_d N_A_1271_74#_M1024_g N_A_1271_74#_c_1216_n
+ N_A_1271_74#_c_1217_n N_A_1271_74#_M1014_g N_A_1271_74#_c_1207_n
+ N_A_1271_74#_c_1208_n N_A_1271_74#_c_1220_n N_A_1271_74#_c_1221_n
+ N_A_1271_74#_M1002_g N_A_1271_74#_M1022_g N_A_1271_74#_c_1210_n
+ N_A_1271_74#_c_1249_n N_A_1271_74#_c_1211_n N_A_1271_74#_c_1223_n
+ N_A_1271_74#_c_1212_n N_A_1271_74#_c_1237_n N_A_1271_74#_c_1338_p
+ N_A_1271_74#_c_1224_n N_A_1271_74#_c_1213_n N_A_1271_74#_c_1214_n
+ N_A_1271_74#_c_1215_n N_A_1271_74#_c_1228_n
+ PM_SKY130_FD_SC_HS__DFRTP_2%A_1271_74#
x_PM_SKY130_FD_SC_HS__DFRTP_2%A_1921_409# N_A_1921_409#_M1022_d
+ N_A_1921_409#_M1002_d N_A_1921_409#_c_1354_n N_A_1921_409#_c_1355_n
+ N_A_1921_409#_c_1367_n N_A_1921_409#_M1004_g N_A_1921_409#_M1031_g
+ N_A_1921_409#_c_1357_n N_A_1921_409#_c_1358_n N_A_1921_409#_c_1369_n
+ N_A_1921_409#_M1006_g N_A_1921_409#_M1033_g N_A_1921_409#_c_1360_n
+ N_A_1921_409#_c_1361_n N_A_1921_409#_c_1370_n N_A_1921_409#_c_1362_n
+ N_A_1921_409#_c_1363_n N_A_1921_409#_c_1364_n N_A_1921_409#_c_1365_n
+ PM_SKY130_FD_SC_HS__DFRTP_2%A_1921_409#
x_PM_SKY130_FD_SC_HS__DFRTP_2%VPWR N_VPWR_M1016_s N_VPWR_M1017_d N_VPWR_M1007_d
+ N_VPWR_M1027_d N_VPWR_M1013_s N_VPWR_M1011_d N_VPWR_M1014_d N_VPWR_M1004_s
+ N_VPWR_M1006_s N_VPWR_c_1427_n N_VPWR_c_1428_n N_VPWR_c_1429_n N_VPWR_c_1430_n
+ N_VPWR_c_1431_n N_VPWR_c_1432_n N_VPWR_c_1433_n N_VPWR_c_1434_n
+ N_VPWR_c_1435_n N_VPWR_c_1436_n N_VPWR_c_1437_n N_VPWR_c_1438_n
+ N_VPWR_c_1439_n N_VPWR_c_1440_n VPWR N_VPWR_c_1441_n N_VPWR_c_1442_n
+ N_VPWR_c_1443_n N_VPWR_c_1444_n N_VPWR_c_1445_n N_VPWR_c_1446_n
+ N_VPWR_c_1447_n N_VPWR_c_1448_n N_VPWR_c_1449_n N_VPWR_c_1450_n
+ N_VPWR_c_1451_n N_VPWR_c_1452_n N_VPWR_c_1426_n
+ PM_SKY130_FD_SC_HS__DFRTP_2%VPWR
x_PM_SKY130_FD_SC_HS__DFRTP_2%A_30_78# N_A_30_78#_M1030_s N_A_30_78#_M1029_s
+ N_A_30_78#_M1016_d N_A_30_78#_M1005_s N_A_30_78#_c_1576_n N_A_30_78#_c_1582_n
+ N_A_30_78#_c_1583_n N_A_30_78#_c_1577_n N_A_30_78#_c_1585_n
+ N_A_30_78#_c_1578_n N_A_30_78#_c_1586_n N_A_30_78#_c_1579_n
+ N_A_30_78#_c_1580_n N_A_30_78#_c_1588_n N_A_30_78#_c_1581_n
+ PM_SKY130_FD_SC_HS__DFRTP_2%A_30_78#
x_PM_SKY130_FD_SC_HS__DFRTP_2%Q N_Q_M1031_d N_Q_M1004_d Q Q Q Q Q Q Q
+ PM_SKY130_FD_SC_HS__DFRTP_2%Q
x_PM_SKY130_FD_SC_HS__DFRTP_2%VGND N_VGND_M1018_d N_VGND_M1000_d N_VGND_M1001_d
+ N_VGND_M1010_d N_VGND_M1022_s N_VGND_M1031_s N_VGND_M1033_s N_VGND_c_1714_n
+ N_VGND_c_1715_n N_VGND_c_1716_n N_VGND_c_1717_n N_VGND_c_1718_n
+ N_VGND_c_1719_n N_VGND_c_1720_n N_VGND_c_1721_n N_VGND_c_1722_n VGND
+ N_VGND_c_1723_n N_VGND_c_1724_n N_VGND_c_1725_n N_VGND_c_1726_n
+ N_VGND_c_1727_n N_VGND_c_1728_n N_VGND_c_1729_n N_VGND_c_1730_n
+ N_VGND_c_1731_n N_VGND_c_1732_n N_VGND_c_1733_n
+ PM_SKY130_FD_SC_HS__DFRTP_2%VGND
cc_1 VNB N_D_c_243_n 0.040598f $X=-0.19 $Y=-0.245 $X2=0.402 $Y2=1.828
cc_2 VNB N_D_M1030_g 0.0286454f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=0.6
cc_3 VNB N_D_c_245_n 0.0216261f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.165
cc_4 VNB N_D_c_246_n 0.0279969f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.165
cc_5 VNB N_RESET_B_M1018_g 0.0291205f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.01
cc_6 VNB N_RESET_B_c_278_n 0.0248218f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.75
cc_7 VNB N_RESET_B_c_279_n 0.018109f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_8 VNB N_RESET_B_c_280_n 0.0106864f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_RESET_B_M1023_g 0.0519208f $X=-0.19 $Y=-0.245 $X2=0.402 $Y2=2.01
cc_10 VNB N_RESET_B_c_282_n 0.0158834f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_RESET_B_c_283_n 0.0297134f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_RESET_B_c_284_n 0.00416334f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_CLK_M1000_g 0.0270176f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.01
cc_14 VNB N_CLK_c_468_n 0.0213158f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.465
cc_15 VNB CLK 0.00455737f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=1
cc_16 VNB N_A_490_362#_c_510_n 0.0121367f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.95
cc_17 VNB N_A_490_362#_M1028_g 0.0242576f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_490_362#_c_512_n 0.0178063f $X=-0.19 $Y=-0.245 $X2=0.402 $Y2=1.165
cc_19 VNB N_A_490_362#_c_513_n 0.0205353f $X=-0.19 $Y=-0.245 $X2=0.402 $Y2=1
cc_20 VNB N_A_490_362#_c_514_n 0.010064f $X=-0.19 $Y=-0.245 $X2=0.402 $Y2=1.845
cc_21 VNB N_A_490_362#_c_515_n 0.0117162f $X=-0.19 $Y=-0.245 $X2=0.31 $Y2=1.295
cc_22 VNB N_A_490_362#_c_516_n 0.0345331f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_490_362#_c_517_n 0.00385131f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_490_362#_c_518_n 0.0145916f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_490_362#_c_519_n 0.00246106f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_490_362#_c_520_n 0.0036821f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_490_362#_c_521_n 0.00197952f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_490_362#_c_522_n 0.0141757f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_490_362#_c_523_n 0.0110381f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_490_362#_c_524_n 0.0318573f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_490_362#_c_525_n 0.00728799f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_837_359#_M1015_g 0.0304105f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_33 VNB N_A_837_359#_c_704_n 0.00259049f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_837_359#_c_705_n 0.0109483f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.165
cc_35 VNB N_A_837_359#_c_706_n 0.00239189f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_837_359#_c_707_n 0.00880031f $X=-0.19 $Y=-0.245 $X2=0.31 $Y2=1.845
cc_37 VNB N_A_696_457#_M1025_g 0.0236184f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_38 VNB N_A_696_457#_c_786_n 0.0170235f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.95
cc_39 VNB N_A_696_457#_c_787_n 0.026897f $X=-0.19 $Y=-0.245 $X2=0.402 $Y2=1.165
cc_40 VNB N_A_696_457#_c_788_n 0.00520122f $X=-0.19 $Y=-0.245 $X2=0.385
+ $Y2=1.165
cc_41 VNB N_A_696_457#_c_789_n 0.00251544f $X=-0.19 $Y=-0.245 $X2=0.402 $Y2=2.01
cc_42 VNB N_A_696_457#_c_790_n 0.00408962f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_696_457#_c_791_n 0.00300945f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_306_74#_c_906_n 0.0201899f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=0.6
cc_45 VNB N_A_306_74#_c_907_n 0.0472689f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_46 VNB N_A_306_74#_c_908_n 0.0169088f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.165
cc_47 VNB N_A_306_74#_c_909_n 0.0126064f $X=-0.19 $Y=-0.245 $X2=0.31 $Y2=2.035
cc_48 VNB N_A_306_74#_M1032_g 0.0521291f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A_306_74#_c_911_n 0.0159808f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_A_306_74#_c_912_n 0.0101157f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_A_306_74#_c_913_n 0.00770987f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_A_306_74#_c_914_n 0.00418354f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_A_306_74#_c_915_n 3.14539e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_A_306_74#_c_916_n 0.0156124f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_A_306_74#_c_917_n 0.00492726f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_A_1525_212#_M1010_g 0.0235036f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=0.6
cc_57 VNB N_A_1525_212#_c_1089_n 0.013872f $X=-0.19 $Y=-0.245 $X2=0.402
+ $Y2=1.165
cc_58 VNB N_A_1525_212#_c_1090_n 0.0150411f $X=-0.19 $Y=-0.245 $X2=0.385
+ $Y2=1.165
cc_59 VNB N_A_1525_212#_c_1091_n 0.0124228f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_A_1525_212#_c_1092_n 0.0141072f $X=-0.19 $Y=-0.245 $X2=0.31
+ $Y2=2.035
cc_61 VNB N_A_1525_212#_c_1093_n 0.00326635f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_A_1525_212#_c_1094_n 0.00415979f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_A_1525_212#_c_1095_n 0.031534f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_A_1525_212#_c_1096_n 0.00288865f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_A_1271_74#_M1024_g 0.0561848f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=0.6
cc_66 VNB N_A_1271_74#_c_1207_n 0.0155616f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_A_1271_74#_c_1208_n 0.0127478f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_A_1271_74#_M1022_g 0.0397312f $X=-0.19 $Y=-0.245 $X2=0.402 $Y2=2.01
cc_69 VNB N_A_1271_74#_c_1210_n 0.00459979f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_A_1271_74#_c_1211_n 0.00477322f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_A_1271_74#_c_1212_n 0.00415183f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_A_1271_74#_c_1213_n 0.00523477f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_A_1271_74#_c_1214_n 0.00751489f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_A_1271_74#_c_1215_n 0.00236307f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_A_1921_409#_c_1354_n 0.0140421f $X=-0.19 $Y=-0.245 $X2=0.495
+ $Y2=2.75
cc_76 VNB N_A_1921_409#_c_1355_n 0.0102109f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=0.6
cc_77 VNB N_A_1921_409#_M1031_g 0.0229651f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_A_1921_409#_c_1357_n 0.00938445f $X=-0.19 $Y=-0.245 $X2=0.402
+ $Y2=1.165
cc_79 VNB N_A_1921_409#_c_1358_n 0.0167069f $X=-0.19 $Y=-0.245 $X2=0.402 $Y2=1
cc_80 VNB N_A_1921_409#_M1033_g 0.0260342f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_81 VNB N_A_1921_409#_c_1360_n 0.00591123f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_82 VNB N_A_1921_409#_c_1361_n 0.0111562f $X=-0.19 $Y=-0.245 $X2=0.31
+ $Y2=1.665
cc_83 VNB N_A_1921_409#_c_1362_n 0.0124224f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_84 VNB N_A_1921_409#_c_1363_n 0.00109385f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_85 VNB N_A_1921_409#_c_1364_n 0.00157695f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_86 VNB N_A_1921_409#_c_1365_n 0.0465967f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_87 VNB N_VPWR_c_1426_n 0.48212f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_88 VNB N_A_30_78#_c_1576_n 0.00271393f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_89 VNB N_A_30_78#_c_1577_n 0.00538705f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.165
cc_90 VNB N_A_30_78#_c_1578_n 0.00267561f $X=-0.19 $Y=-0.245 $X2=0.402 $Y2=2.01
cc_91 VNB N_A_30_78#_c_1579_n 0.00362936f $X=-0.19 $Y=-0.245 $X2=0.31 $Y2=1.665
cc_92 VNB N_A_30_78#_c_1580_n 0.0223919f $X=-0.19 $Y=-0.245 $X2=0.31 $Y2=1.845
cc_93 VNB N_A_30_78#_c_1581_n 0.00727981f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_94 VNB Q 0.00240191f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.75
cc_95 VNB N_VGND_c_1714_n 0.016244f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.845
cc_96 VNB N_VGND_c_1715_n 0.00962093f $X=-0.19 $Y=-0.245 $X2=0.31 $Y2=1.295
cc_97 VNB N_VGND_c_1716_n 0.00612754f $X=-0.19 $Y=-0.245 $X2=0.31 $Y2=1.845
cc_98 VNB N_VGND_c_1717_n 0.0164559f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_99 VNB N_VGND_c_1718_n 0.0191664f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_100 VNB N_VGND_c_1719_n 0.0105185f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_101 VNB N_VGND_c_1720_n 0.0507342f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_102 VNB N_VGND_c_1721_n 0.0308567f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_103 VNB N_VGND_c_1722_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_104 VNB N_VGND_c_1723_n 0.0201745f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_105 VNB N_VGND_c_1724_n 0.083627f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_106 VNB N_VGND_c_1725_n 0.0578377f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_107 VNB N_VGND_c_1726_n 0.0306389f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_108 VNB N_VGND_c_1727_n 0.0209223f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_109 VNB N_VGND_c_1728_n 0.0193312f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_110 VNB N_VGND_c_1729_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_111 VNB N_VGND_c_1730_n 0.0080786f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_112 VNB N_VGND_c_1731_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_113 VNB N_VGND_c_1732_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_114 VNB N_VGND_c_1733_n 0.648176f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_115 VPB N_D_c_243_n 0.0142136f $X=-0.19 $Y=1.66 $X2=0.402 $Y2=1.828
cc_116 VPB N_D_c_248_n 0.0278558f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=2.375
cc_117 VPB N_D_c_249_n 0.0277344f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=2.465
cc_118 VPB N_D_c_246_n 0.0227717f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.165
cc_119 VPB N_D_c_251_n 0.0207699f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.845
cc_120 VPB N_RESET_B_c_278_n 0.0228603f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=2.75
cc_121 VPB N_RESET_B_c_286_n 0.0177526f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=1
cc_122 VPB N_RESET_B_c_287_n 0.0251577f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=0.6
cc_123 VPB N_RESET_B_c_280_n 0.0183715f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_124 VPB N_RESET_B_c_289_n 0.0701332f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_125 VPB N_RESET_B_c_290_n 0.0571202f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.165
cc_126 VPB N_RESET_B_M1023_g 0.0162636f $X=-0.19 $Y=1.66 $X2=0.402 $Y2=2.01
cc_127 VPB N_RESET_B_c_292_n 0.0209249f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_128 VPB N_RESET_B_c_293_n 0.00493187f $X=-0.19 $Y=1.66 $X2=0.31 $Y2=1.845
cc_129 VPB N_RESET_B_c_294_n 0.020195f $X=-0.19 $Y=1.66 $X2=0.31 $Y2=2.035
cc_130 VPB N_RESET_B_c_295_n 0.00143938f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_131 VPB N_RESET_B_c_296_n 0.00397837f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_132 VPB N_RESET_B_c_297_n 0.0019787f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_133 VPB N_RESET_B_c_284_n 9.70225e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_134 VPB N_RESET_B_c_299_n 0.0269424f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_135 VPB N_RESET_B_c_300_n 0.00930396f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_136 VPB N_CLK_c_468_n 0.0333341f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=2.465
cc_137 VPB CLK 0.00648163f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=1
cc_138 VPB N_A_490_362#_c_526_n 0.0134498f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=1
cc_139 VPB N_A_490_362#_c_527_n 0.0196842f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=0.6
cc_140 VPB N_A_490_362#_c_528_n 0.0224904f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.21
cc_141 VPB N_A_490_362#_c_510_n 0.0127361f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.95
cc_142 VPB N_A_490_362#_c_530_n 0.0194137f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.845
cc_143 VPB N_A_490_362#_c_515_n 5.88973e-19 $X=-0.19 $Y=1.66 $X2=0.31 $Y2=1.295
cc_144 VPB N_A_490_362#_c_532_n 0.00465503f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_145 VPB N_A_490_362#_c_533_n 0.00238555f $X=-0.19 $Y=1.66 $X2=0.31 $Y2=2.035
cc_146 VPB N_A_490_362#_c_520_n 0.006052f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_147 VPB N_A_490_362#_c_535_n 0.0479926f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_148 VPB N_A_490_362#_c_536_n 0.029384f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_149 VPB N_A_837_359#_c_708_n 0.0603018f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=2.75
cc_150 VPB N_A_837_359#_M1015_g 0.0134261f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.21
cc_151 VPB N_A_837_359#_c_704_n 0.00264531f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_152 VPB N_A_837_359#_c_711_n 5.83759e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_153 VPB N_A_837_359#_c_707_n 0.00377881f $X=-0.19 $Y=1.66 $X2=0.31 $Y2=1.845
cc_154 VPB N_A_696_457#_c_786_n 0.0288648f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.95
cc_155 VPB N_A_696_457#_c_787_n 0.0122975f $X=-0.19 $Y=1.66 $X2=0.402 $Y2=1.165
cc_156 VPB N_A_696_457#_c_788_n 0.00959354f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.165
cc_157 VPB N_A_696_457#_c_795_n 0.00288162f $X=-0.19 $Y=1.66 $X2=0.402 $Y2=1.845
cc_158 VPB N_A_696_457#_c_796_n 0.0112403f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.845
cc_159 VPB N_A_696_457#_c_790_n 0.00331109f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_160 VPB N_A_696_457#_c_798_n 0.00268299f $X=-0.19 $Y=1.66 $X2=0.31 $Y2=1.845
cc_161 VPB N_A_306_74#_c_918_n 0.014621f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=2.75
cc_162 VPB N_A_306_74#_c_919_n 0.0786009f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_163 VPB N_A_306_74#_c_920_n 0.0563854f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_164 VPB N_A_306_74#_c_921_n 0.0125824f $X=-0.19 $Y=1.66 $X2=0.402 $Y2=1.165
cc_165 VPB N_A_306_74#_c_922_n 0.00719725f $X=-0.19 $Y=1.66 $X2=0.402 $Y2=1.845
cc_166 VPB N_A_306_74#_c_923_n 0.0193529f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.845
cc_167 VPB N_A_306_74#_c_924_n 0.0146805f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.845
cc_168 VPB N_A_306_74#_c_925_n 0.175803f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_169 VPB N_A_306_74#_M1021_g 0.0107276f $X=-0.19 $Y=1.66 $X2=0.31 $Y2=1.845
cc_170 VPB N_A_306_74#_c_909_n 0.0397359f $X=-0.19 $Y=1.66 $X2=0.31 $Y2=2.035
cc_171 VPB N_A_306_74#_c_928_n 0.00832634f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_172 VPB N_A_306_74#_c_929_n 0.0282456f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_173 VPB N_A_306_74#_c_930_n 0.00898671f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_174 VPB N_A_306_74#_c_931_n 0.0335383f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_175 VPB N_A_306_74#_c_913_n 0.00528291f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_176 VPB N_A_306_74#_c_916_n 0.00122818f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_177 VPB N_A_306_74#_c_934_n 0.00417949f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_178 VPB N_A_1525_212#_c_1097_n 0.00452844f $X=-0.19 $Y=1.66 $X2=0.155
+ $Y2=1.58
cc_179 VPB N_A_1525_212#_c_1098_n 0.0112203f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.95
cc_180 VPB N_A_1525_212#_c_1099_n 0.0209833f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_181 VPB N_A_1525_212#_c_1089_n 0.0172903f $X=-0.19 $Y=1.66 $X2=0.402
+ $Y2=1.165
cc_182 VPB N_A_1525_212#_c_1101_n 0.0123021f $X=-0.19 $Y=1.66 $X2=0.402 $Y2=1
cc_183 VPB N_A_1525_212#_c_1102_n 0.00195592f $X=-0.19 $Y=1.66 $X2=0.31
+ $Y2=1.665
cc_184 VPB N_A_1525_212#_c_1103_n 0.00467452f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_185 VPB N_A_1525_212#_c_1104_n 0.00234171f $X=-0.19 $Y=1.66 $X2=0.31
+ $Y2=1.845
cc_186 VPB N_A_1525_212#_c_1093_n 0.00587125f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_187 VPB N_A_1271_74#_c_1216_n 0.0253818f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.21
cc_188 VPB N_A_1271_74#_c_1217_n 0.0240491f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_189 VPB N_A_1271_74#_c_1207_n 0.00814854f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_190 VPB N_A_1271_74#_c_1208_n 0.0260612f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_191 VPB N_A_1271_74#_c_1220_n 0.010774f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.165
cc_192 VPB N_A_1271_74#_c_1221_n 0.0240694f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.165
cc_193 VPB N_A_1271_74#_c_1210_n 0.00430295f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_194 VPB N_A_1271_74#_c_1223_n 0.00135315f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_195 VPB N_A_1271_74#_c_1224_n 0.0127664f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_196 VPB N_A_1271_74#_c_1213_n 0.0140489f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_197 VPB N_A_1271_74#_c_1214_n 4.13852e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_198 VPB N_A_1271_74#_c_1215_n 4.64263e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_199 VPB N_A_1271_74#_c_1228_n 0.00154868f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_200 VPB N_A_1921_409#_c_1355_n 8.65682e-19 $X=-0.19 $Y=1.66 $X2=0.51 $Y2=0.6
cc_201 VPB N_A_1921_409#_c_1367_n 0.023821f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_202 VPB N_A_1921_409#_c_1358_n 0.00111912f $X=-0.19 $Y=1.66 $X2=0.402 $Y2=1
cc_203 VPB N_A_1921_409#_c_1369_n 0.0258791f $X=-0.19 $Y=1.66 $X2=0.402
+ $Y2=1.845
cc_204 VPB N_A_1921_409#_c_1370_n 0.0117303f $X=-0.19 $Y=1.66 $X2=0.31 $Y2=2.035
cc_205 VPB N_A_1921_409#_c_1363_n 0.00710574f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_206 VPB N_VPWR_c_1427_n 0.0116916f $X=-0.19 $Y=1.66 $X2=0.31 $Y2=1.295
cc_207 VPB N_VPWR_c_1428_n 0.0302409f $X=-0.19 $Y=1.66 $X2=0.31 $Y2=1.665
cc_208 VPB N_VPWR_c_1429_n 0.00955952f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_209 VPB N_VPWR_c_1430_n 0.00426746f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_210 VPB N_VPWR_c_1431_n 0.0147915f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_211 VPB N_VPWR_c_1432_n 0.0202814f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_212 VPB N_VPWR_c_1433_n 0.0249252f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_213 VPB N_VPWR_c_1434_n 0.0152192f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_214 VPB N_VPWR_c_1435_n 0.0163857f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_215 VPB N_VPWR_c_1436_n 0.0261554f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_216 VPB N_VPWR_c_1437_n 0.0106521f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_217 VPB N_VPWR_c_1438_n 0.0638885f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_218 VPB N_VPWR_c_1439_n 0.0275707f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_219 VPB N_VPWR_c_1440_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_220 VPB N_VPWR_c_1441_n 0.0162121f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_221 VPB N_VPWR_c_1442_n 0.0206207f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_222 VPB N_VPWR_c_1443_n 0.0608968f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_223 VPB N_VPWR_c_1444_n 0.0531608f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_224 VPB N_VPWR_c_1445_n 0.0209549f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_225 VPB N_VPWR_c_1446_n 0.0188539f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_226 VPB N_VPWR_c_1447_n 0.00614127f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_227 VPB N_VPWR_c_1448_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_228 VPB N_VPWR_c_1449_n 0.00436768f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_229 VPB N_VPWR_c_1450_n 0.00436868f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_230 VPB N_VPWR_c_1451_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_231 VPB N_VPWR_c_1452_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_232 VPB N_VPWR_c_1426_n 0.119001f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_233 VPB N_A_30_78#_c_1582_n 0.00391052f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_234 VPB N_A_30_78#_c_1583_n 0.00206042f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_235 VPB N_A_30_78#_c_1577_n 0.00585658f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.165
cc_236 VPB N_A_30_78#_c_1585_n 0.0157677f $X=-0.19 $Y=1.66 $X2=0.402 $Y2=1
cc_237 VPB N_A_30_78#_c_1586_n 0.00730131f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_238 VPB N_A_30_78#_c_1579_n 0.00599832f $X=-0.19 $Y=1.66 $X2=0.31 $Y2=1.665
cc_239 VPB N_A_30_78#_c_1588_n 0.00841498f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_240 VPB Q 0.00331763f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=2.75
cc_241 N_D_M1030_g N_RESET_B_M1018_g 0.0244236f $X=0.51 $Y=0.6 $X2=0 $Y2=0
cc_242 N_D_c_246_n N_RESET_B_M1018_g 9.45409e-19 $X=0.385 $Y=1.165 $X2=0 $Y2=0
cc_243 N_D_c_243_n N_RESET_B_c_278_n 0.0244236f $X=0.402 $Y=1.828 $X2=0 $Y2=0
cc_244 N_D_c_248_n N_RESET_B_c_286_n 0.0062784f $X=0.495 $Y=2.375 $X2=0 $Y2=0
cc_245 N_D_c_249_n N_RESET_B_c_287_n 0.01449f $X=0.495 $Y=2.465 $X2=0 $Y2=0
cc_246 N_D_c_245_n N_RESET_B_c_283_n 0.0244236f $X=0.385 $Y=1.165 $X2=0 $Y2=0
cc_247 N_D_c_251_n N_RESET_B_c_299_n 0.0244236f $X=0.385 $Y=1.845 $X2=0 $Y2=0
cc_248 N_D_c_249_n N_VPWR_c_1428_n 0.0113574f $X=0.495 $Y=2.465 $X2=0 $Y2=0
cc_249 N_D_c_246_n N_VPWR_c_1428_n 0.0172326f $X=0.385 $Y=1.165 $X2=0 $Y2=0
cc_250 N_D_c_251_n N_VPWR_c_1428_n 9.92489e-19 $X=0.385 $Y=1.845 $X2=0 $Y2=0
cc_251 N_D_c_249_n N_VPWR_c_1429_n 4.09834e-19 $X=0.495 $Y=2.465 $X2=0 $Y2=0
cc_252 N_D_c_249_n N_VPWR_c_1441_n 0.00413917f $X=0.495 $Y=2.465 $X2=0 $Y2=0
cc_253 N_D_c_249_n N_VPWR_c_1426_n 0.00855638f $X=0.495 $Y=2.465 $X2=0 $Y2=0
cc_254 N_D_M1030_g N_A_30_78#_c_1576_n 0.0114706f $X=0.51 $Y=0.6 $X2=0 $Y2=0
cc_255 N_D_c_246_n N_A_30_78#_c_1576_n 0.00258996f $X=0.385 $Y=1.165 $X2=0 $Y2=0
cc_256 N_D_c_248_n N_A_30_78#_c_1582_n 0.00445133f $X=0.495 $Y=2.375 $X2=0 $Y2=0
cc_257 N_D_c_249_n N_A_30_78#_c_1582_n 0.00192676f $X=0.495 $Y=2.465 $X2=0 $Y2=0
cc_258 N_D_c_249_n N_A_30_78#_c_1583_n 0.00132898f $X=0.495 $Y=2.465 $X2=0 $Y2=0
cc_259 N_D_M1030_g N_A_30_78#_c_1577_n 0.0152471f $X=0.51 $Y=0.6 $X2=0 $Y2=0
cc_260 N_D_c_246_n N_A_30_78#_c_1577_n 0.088088f $X=0.385 $Y=1.165 $X2=0 $Y2=0
cc_261 N_D_M1030_g N_A_30_78#_c_1580_n 0.00806237f $X=0.51 $Y=0.6 $X2=0 $Y2=0
cc_262 N_D_c_245_n N_A_30_78#_c_1580_n 0.00161806f $X=0.385 $Y=1.165 $X2=0 $Y2=0
cc_263 N_D_c_246_n N_A_30_78#_c_1580_n 0.0286676f $X=0.385 $Y=1.165 $X2=0 $Y2=0
cc_264 N_D_M1030_g N_VGND_c_1721_n 0.00429844f $X=0.51 $Y=0.6 $X2=0 $Y2=0
cc_265 N_D_M1030_g N_VGND_c_1733_n 0.00539454f $X=0.51 $Y=0.6 $X2=0 $Y2=0
cc_266 N_RESET_B_c_283_n N_CLK_M1000_g 0.00270964f $X=1.12 $Y=1.305 $X2=0 $Y2=0
cc_267 N_RESET_B_c_278_n N_CLK_c_468_n 0.00555016f $X=1.055 $Y=1.92 $X2=0 $Y2=0
cc_268 N_RESET_B_c_292_n N_CLK_c_468_n 0.00422081f $X=4.895 $Y=2.035 $X2=0 $Y2=0
cc_269 N_RESET_B_c_283_n N_CLK_c_468_n 0.00646425f $X=1.12 $Y=1.305 $X2=0 $Y2=0
cc_270 N_RESET_B_c_292_n CLK 0.0118867f $X=4.895 $Y=2.035 $X2=0 $Y2=0
cc_271 N_RESET_B_c_292_n N_A_490_362#_M1012_d 0.00121208f $X=4.895 $Y=2.035
+ $X2=0 $Y2=0
cc_272 N_RESET_B_c_292_n N_A_490_362#_c_526_n 0.00396062f $X=4.895 $Y=2.035
+ $X2=0 $Y2=0
cc_273 N_RESET_B_c_292_n N_A_490_362#_c_528_n 0.00439233f $X=4.895 $Y=2.035
+ $X2=0 $Y2=0
cc_274 N_RESET_B_c_292_n N_A_490_362#_c_532_n 0.0287414f $X=4.895 $Y=2.035 $X2=0
+ $Y2=0
cc_275 N_RESET_B_c_292_n N_A_490_362#_c_533_n 0.0107516f $X=4.895 $Y=2.035 $X2=0
+ $Y2=0
cc_276 N_RESET_B_c_279_n N_A_490_362#_c_517_n 0.0123973f $X=4.79 $Y=1.185 $X2=0
+ $Y2=0
cc_277 N_RESET_B_c_279_n N_A_490_362#_c_543_n 0.00113651f $X=4.79 $Y=1.185 $X2=0
+ $Y2=0
cc_278 N_RESET_B_c_294_n N_A_490_362#_c_520_n 0.0218177f $X=7.775 $Y=2.035 $X2=0
+ $Y2=0
cc_279 N_RESET_B_c_294_n N_A_490_362#_c_535_n 0.00331406f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_280 N_RESET_B_c_279_n N_A_490_362#_c_523_n 4.35744e-19 $X=4.79 $Y=1.185 $X2=0
+ $Y2=0
cc_281 N_RESET_B_c_292_n N_A_490_362#_c_536_n 0.0038641f $X=4.895 $Y=2.035 $X2=0
+ $Y2=0
cc_282 N_RESET_B_c_294_n N_A_837_359#_M1013_d 0.00226165f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_283 N_RESET_B_c_289_n N_A_837_359#_c_708_n 0.030599f $X=4.895 $Y=2.21 $X2=0
+ $Y2=0
cc_284 N_RESET_B_c_292_n N_A_837_359#_c_708_n 0.0103415f $X=4.895 $Y=2.035 $X2=0
+ $Y2=0
cc_285 N_RESET_B_c_279_n N_A_837_359#_M1015_g 0.0419644f $X=4.79 $Y=1.185 $X2=0
+ $Y2=0
cc_286 N_RESET_B_c_280_n N_A_837_359#_M1015_g 0.0138048f $X=4.88 $Y=1.795 $X2=0
+ $Y2=0
cc_287 N_RESET_B_c_279_n N_A_837_359#_c_704_n 0.00106151f $X=4.79 $Y=1.185 $X2=0
+ $Y2=0
cc_288 N_RESET_B_c_280_n N_A_837_359#_c_704_n 4.52393e-19 $X=4.88 $Y=1.795 $X2=0
+ $Y2=0
cc_289 N_RESET_B_c_292_n N_A_837_359#_c_704_n 0.0166888f $X=4.895 $Y=2.035 $X2=0
+ $Y2=0
cc_290 N_RESET_B_c_279_n N_A_837_359#_c_705_n 0.0122236f $X=4.79 $Y=1.185 $X2=0
+ $Y2=0
cc_291 N_RESET_B_c_282_n N_A_837_359#_c_705_n 0.00269956f $X=4.88 $Y=1.26 $X2=0
+ $Y2=0
cc_292 N_RESET_B_c_294_n N_A_837_359#_c_711_n 0.0386269f $X=7.775 $Y=2.035 $X2=0
+ $Y2=0
cc_293 N_RESET_B_c_294_n N_A_696_457#_c_786_n 0.0121958f $X=7.775 $Y=2.035 $X2=0
+ $Y2=0
cc_294 N_RESET_B_c_282_n N_A_696_457#_c_787_n 0.00991362f $X=4.88 $Y=1.26 $X2=0
+ $Y2=0
cc_295 N_RESET_B_c_294_n N_A_696_457#_c_787_n 0.00341453f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_296 N_RESET_B_c_292_n N_A_696_457#_c_788_n 0.018625f $X=4.895 $Y=2.035 $X2=0
+ $Y2=0
cc_297 N_RESET_B_c_292_n N_A_696_457#_c_803_n 0.0137798f $X=4.895 $Y=2.035 $X2=0
+ $Y2=0
cc_298 N_RESET_B_c_292_n N_A_696_457#_c_795_n 0.00793203f $X=4.895 $Y=2.035
+ $X2=0 $Y2=0
cc_299 N_RESET_B_c_280_n N_A_696_457#_c_796_n 0.0102353f $X=4.88 $Y=1.795 $X2=0
+ $Y2=0
cc_300 N_RESET_B_c_289_n N_A_696_457#_c_796_n 0.00222717f $X=4.895 $Y=2.21 $X2=0
+ $Y2=0
cc_301 N_RESET_B_c_292_n N_A_696_457#_c_796_n 0.0210187f $X=4.895 $Y=2.035 $X2=0
+ $Y2=0
cc_302 N_RESET_B_c_295_n N_A_696_457#_c_796_n 0.00242233f $X=5.185 $Y=2.035
+ $X2=0 $Y2=0
cc_303 N_RESET_B_c_296_n N_A_696_457#_c_796_n 0.0245177f $X=5.04 $Y=2.035 $X2=0
+ $Y2=0
cc_304 N_RESET_B_c_282_n N_A_696_457#_c_789_n 0.00324317f $X=4.88 $Y=1.26 $X2=0
+ $Y2=0
cc_305 N_RESET_B_c_280_n N_A_696_457#_c_790_n 0.012327f $X=4.88 $Y=1.795 $X2=0
+ $Y2=0
cc_306 N_RESET_B_c_289_n N_A_696_457#_c_790_n 0.00732939f $X=4.895 $Y=2.21 $X2=0
+ $Y2=0
cc_307 N_RESET_B_c_282_n N_A_696_457#_c_790_n 0.0034188f $X=4.88 $Y=1.26 $X2=0
+ $Y2=0
cc_308 N_RESET_B_c_292_n N_A_696_457#_c_790_n 0.00355574f $X=4.895 $Y=2.035
+ $X2=0 $Y2=0
cc_309 N_RESET_B_c_294_n N_A_696_457#_c_790_n 0.0096202f $X=7.775 $Y=2.035 $X2=0
+ $Y2=0
cc_310 N_RESET_B_c_295_n N_A_696_457#_c_790_n 0.00343479f $X=5.185 $Y=2.035
+ $X2=0 $Y2=0
cc_311 N_RESET_B_c_296_n N_A_696_457#_c_790_n 0.019281f $X=5.04 $Y=2.035 $X2=0
+ $Y2=0
cc_312 N_RESET_B_c_289_n N_A_696_457#_c_798_n 0.0149971f $X=4.895 $Y=2.21 $X2=0
+ $Y2=0
cc_313 N_RESET_B_c_292_n N_A_696_457#_c_798_n 0.00433839f $X=4.895 $Y=2.035
+ $X2=0 $Y2=0
cc_314 N_RESET_B_c_294_n N_A_696_457#_c_798_n 7.0969e-19 $X=7.775 $Y=2.035 $X2=0
+ $Y2=0
cc_315 N_RESET_B_c_295_n N_A_696_457#_c_798_n 0.0087813f $X=5.185 $Y=2.035 $X2=0
+ $Y2=0
cc_316 N_RESET_B_c_296_n N_A_696_457#_c_798_n 0.0210307f $X=5.04 $Y=2.035 $X2=0
+ $Y2=0
cc_317 N_RESET_B_c_292_n N_A_306_74#_c_918_n 0.00905605f $X=4.895 $Y=2.035 $X2=0
+ $Y2=0
cc_318 N_RESET_B_c_292_n N_A_306_74#_c_919_n 0.0025035f $X=4.895 $Y=2.035 $X2=0
+ $Y2=0
cc_319 N_RESET_B_c_292_n N_A_306_74#_c_924_n 0.00257921f $X=4.895 $Y=2.035 $X2=0
+ $Y2=0
cc_320 N_RESET_B_c_289_n N_A_306_74#_c_925_n 0.00850694f $X=4.895 $Y=2.21 $X2=0
+ $Y2=0
cc_321 N_RESET_B_c_294_n N_A_306_74#_M1021_g 0.00854421f $X=7.775 $Y=2.035 $X2=0
+ $Y2=0
cc_322 N_RESET_B_c_294_n N_A_306_74#_c_909_n 0.00771224f $X=7.775 $Y=2.035 $X2=0
+ $Y2=0
cc_323 N_RESET_B_c_292_n N_A_306_74#_c_929_n 0.00211295f $X=4.895 $Y=2.035 $X2=0
+ $Y2=0
cc_324 N_RESET_B_M1018_g N_A_306_74#_c_912_n 0.0032696f $X=0.9 $Y=0.6 $X2=0
+ $Y2=0
cc_325 N_RESET_B_c_292_n N_A_306_74#_c_913_n 9.2465e-19 $X=4.895 $Y=2.035 $X2=0
+ $Y2=0
cc_326 N_RESET_B_c_283_n N_A_306_74#_c_913_n 0.00622775f $X=1.12 $Y=1.305 $X2=0
+ $Y2=0
cc_327 N_RESET_B_c_284_n N_A_306_74#_c_913_n 0.0496559f $X=1.12 $Y=1.305 $X2=0
+ $Y2=0
cc_328 N_RESET_B_c_292_n N_A_306_74#_c_915_n 0.0033665f $X=4.895 $Y=2.035 $X2=0
+ $Y2=0
cc_329 N_RESET_B_M1018_g N_A_306_74#_c_917_n 0.00281599f $X=0.9 $Y=0.6 $X2=0
+ $Y2=0
cc_330 N_RESET_B_c_284_n N_A_306_74#_c_917_n 8.33963e-19 $X=1.12 $Y=1.305 $X2=0
+ $Y2=0
cc_331 N_RESET_B_c_278_n N_A_306_74#_c_934_n 0.00281328f $X=1.055 $Y=1.92 $X2=0
+ $Y2=0
cc_332 N_RESET_B_c_292_n N_A_306_74#_c_934_n 0.0249775f $X=4.895 $Y=2.035 $X2=0
+ $Y2=0
cc_333 N_RESET_B_c_293_n N_A_306_74#_c_934_n 0.00278023f $X=1.345 $Y=2.035 $X2=0
+ $Y2=0
cc_334 N_RESET_B_c_284_n N_A_306_74#_c_934_n 0.0235472f $X=1.12 $Y=1.305 $X2=0
+ $Y2=0
cc_335 N_RESET_B_M1023_g N_A_1525_212#_M1010_g 0.0164487f $X=8.24 $Y=0.615 $X2=0
+ $Y2=0
cc_336 N_RESET_B_c_290_n N_A_1525_212#_c_1097_n 0.0164306f $X=8.235 $Y=2.39
+ $X2=0 $Y2=0
cc_337 N_RESET_B_c_294_n N_A_1525_212#_c_1097_n 4.99514e-19 $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_338 N_RESET_B_c_300_n N_A_1525_212#_c_1097_n 0.00182389f $X=8.23 $Y=2.11
+ $X2=0 $Y2=0
cc_339 N_RESET_B_c_290_n N_A_1525_212#_c_1098_n 0.00475599f $X=8.235 $Y=2.39
+ $X2=0 $Y2=0
cc_340 N_RESET_B_c_294_n N_A_1525_212#_c_1098_n 0.0054475f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_341 N_RESET_B_c_297_n N_A_1525_212#_c_1098_n 0.00136519f $X=7.92 $Y=2.035
+ $X2=0 $Y2=0
cc_342 N_RESET_B_c_300_n N_A_1525_212#_c_1098_n 0.00431246f $X=8.23 $Y=2.11
+ $X2=0 $Y2=0
cc_343 N_RESET_B_c_290_n N_A_1525_212#_c_1099_n 0.0121565f $X=8.235 $Y=2.39
+ $X2=0 $Y2=0
cc_344 N_RESET_B_c_290_n N_A_1525_212#_c_1089_n 0.00147213f $X=8.235 $Y=2.39
+ $X2=0 $Y2=0
cc_345 N_RESET_B_M1023_g N_A_1525_212#_c_1089_n 0.0193933f $X=8.24 $Y=0.615
+ $X2=0 $Y2=0
cc_346 N_RESET_B_c_294_n N_A_1525_212#_c_1089_n 0.00138661f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_347 N_RESET_B_c_297_n N_A_1525_212#_c_1089_n 8.33981e-19 $X=7.92 $Y=2.035
+ $X2=0 $Y2=0
cc_348 N_RESET_B_c_300_n N_A_1525_212#_c_1089_n 4.18149e-19 $X=8.23 $Y=2.11
+ $X2=0 $Y2=0
cc_349 N_RESET_B_M1023_g N_A_1525_212#_c_1090_n 0.013811f $X=8.24 $Y=0.615 $X2=0
+ $Y2=0
cc_350 N_RESET_B_c_290_n N_A_1525_212#_c_1101_n 0.0117959f $X=8.235 $Y=2.39
+ $X2=0 $Y2=0
cc_351 N_RESET_B_c_300_n N_A_1525_212#_c_1101_n 0.00789453f $X=8.23 $Y=2.11
+ $X2=0 $Y2=0
cc_352 N_RESET_B_M1023_g N_A_1525_212#_c_1091_n 0.00343438f $X=8.24 $Y=0.615
+ $X2=0 $Y2=0
cc_353 N_RESET_B_c_290_n N_A_1525_212#_c_1102_n 0.00297602f $X=8.235 $Y=2.39
+ $X2=0 $Y2=0
cc_354 N_RESET_B_c_290_n N_A_1525_212#_c_1104_n 8.22326e-19 $X=8.235 $Y=2.39
+ $X2=0 $Y2=0
cc_355 N_RESET_B_c_300_n N_A_1525_212#_c_1104_n 0.0092621f $X=8.23 $Y=2.11 $X2=0
+ $Y2=0
cc_356 N_RESET_B_M1023_g N_A_1525_212#_c_1094_n 0.00118187f $X=8.24 $Y=0.615
+ $X2=0 $Y2=0
cc_357 N_RESET_B_M1023_g N_A_1525_212#_c_1095_n 0.021263f $X=8.24 $Y=0.615 $X2=0
+ $Y2=0
cc_358 N_RESET_B_c_294_n N_A_1271_74#_M1021_d 0.00308066f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_359 N_RESET_B_M1023_g N_A_1271_74#_M1024_g 0.0755988f $X=8.24 $Y=0.615 $X2=0
+ $Y2=0
cc_360 N_RESET_B_c_290_n N_A_1271_74#_c_1216_n 0.00922978f $X=8.235 $Y=2.39
+ $X2=0 $Y2=0
cc_361 N_RESET_B_M1023_g N_A_1271_74#_c_1216_n 0.00125436f $X=8.24 $Y=0.615
+ $X2=0 $Y2=0
cc_362 N_RESET_B_c_300_n N_A_1271_74#_c_1216_n 0.00157069f $X=8.23 $Y=2.11 $X2=0
+ $Y2=0
cc_363 N_RESET_B_c_290_n N_A_1271_74#_c_1217_n 0.0124349f $X=8.235 $Y=2.39 $X2=0
+ $Y2=0
cc_364 N_RESET_B_M1023_g N_A_1271_74#_c_1208_n 0.0061479f $X=8.24 $Y=0.615 $X2=0
+ $Y2=0
cc_365 N_RESET_B_c_294_n N_A_1271_74#_c_1223_n 0.0172254f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_366 N_RESET_B_c_294_n N_A_1271_74#_c_1237_n 0.0184591f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_367 N_RESET_B_c_294_n N_A_1271_74#_c_1224_n 0.0225824f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_368 N_RESET_B_c_297_n N_A_1271_74#_c_1224_n 0.00231685f $X=7.92 $Y=2.035
+ $X2=0 $Y2=0
cc_369 N_RESET_B_c_300_n N_A_1271_74#_c_1224_n 0.023913f $X=8.23 $Y=2.11 $X2=0
+ $Y2=0
cc_370 N_RESET_B_c_290_n N_A_1271_74#_c_1213_n 0.00115984f $X=8.235 $Y=2.39
+ $X2=0 $Y2=0
cc_371 N_RESET_B_M1023_g N_A_1271_74#_c_1213_n 0.0108634f $X=8.24 $Y=0.615 $X2=0
+ $Y2=0
cc_372 N_RESET_B_c_294_n N_A_1271_74#_c_1213_n 0.00539223f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_373 N_RESET_B_c_297_n N_A_1271_74#_c_1213_n 0.00832147f $X=7.92 $Y=2.035
+ $X2=0 $Y2=0
cc_374 N_RESET_B_c_300_n N_A_1271_74#_c_1213_n 0.0386217f $X=8.23 $Y=2.11 $X2=0
+ $Y2=0
cc_375 N_RESET_B_c_294_n N_A_1271_74#_c_1215_n 0.00603357f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_376 N_RESET_B_M1023_g N_A_1271_74#_c_1228_n 0.00100578f $X=8.24 $Y=0.615
+ $X2=0 $Y2=0
cc_377 N_RESET_B_c_292_n N_VPWR_M1007_d 0.00537841f $X=4.895 $Y=2.035 $X2=0
+ $Y2=0
cc_378 N_RESET_B_c_287_n N_VPWR_c_1428_n 4.6593e-19 $X=0.945 $Y=2.465 $X2=0
+ $Y2=0
cc_379 N_RESET_B_c_287_n N_VPWR_c_1429_n 0.00803994f $X=0.945 $Y=2.465 $X2=0
+ $Y2=0
cc_380 N_RESET_B_c_289_n N_VPWR_c_1431_n 0.00230854f $X=4.895 $Y=2.21 $X2=0
+ $Y2=0
cc_381 N_RESET_B_c_280_n N_VPWR_c_1433_n 0.001224f $X=4.88 $Y=1.795 $X2=0 $Y2=0
cc_382 N_RESET_B_c_289_n N_VPWR_c_1433_n 0.0105924f $X=4.895 $Y=2.21 $X2=0 $Y2=0
cc_383 N_RESET_B_c_294_n N_VPWR_c_1433_n 0.0323618f $X=7.775 $Y=2.035 $X2=0
+ $Y2=0
cc_384 N_RESET_B_c_295_n N_VPWR_c_1433_n 5.54746e-19 $X=5.185 $Y=2.035 $X2=0
+ $Y2=0
cc_385 N_RESET_B_c_296_n N_VPWR_c_1433_n 0.0200056f $X=5.04 $Y=2.035 $X2=0 $Y2=0
cc_386 N_RESET_B_c_290_n N_VPWR_c_1434_n 0.0075111f $X=8.235 $Y=2.39 $X2=0 $Y2=0
cc_387 N_RESET_B_c_297_n N_VPWR_c_1434_n 0.00200394f $X=7.92 $Y=2.035 $X2=0
+ $Y2=0
cc_388 N_RESET_B_c_300_n N_VPWR_c_1434_n 0.0263442f $X=8.23 $Y=2.11 $X2=0 $Y2=0
cc_389 N_RESET_B_c_290_n N_VPWR_c_1439_n 0.00511025f $X=8.235 $Y=2.39 $X2=0
+ $Y2=0
cc_390 N_RESET_B_c_287_n N_VPWR_c_1441_n 0.00413917f $X=0.945 $Y=2.465 $X2=0
+ $Y2=0
cc_391 N_RESET_B_c_287_n N_VPWR_c_1426_n 0.00459062f $X=0.945 $Y=2.465 $X2=0
+ $Y2=0
cc_392 N_RESET_B_c_289_n N_VPWR_c_1426_n 9.49986e-19 $X=4.895 $Y=2.21 $X2=0
+ $Y2=0
cc_393 N_RESET_B_c_290_n N_VPWR_c_1426_n 0.0052212f $X=8.235 $Y=2.39 $X2=0 $Y2=0
cc_394 N_RESET_B_M1018_g N_A_30_78#_c_1576_n 0.00370091f $X=0.9 $Y=0.6 $X2=0
+ $Y2=0
cc_395 N_RESET_B_c_287_n N_A_30_78#_c_1582_n 0.00130643f $X=0.945 $Y=2.465 $X2=0
+ $Y2=0
cc_396 N_RESET_B_c_287_n N_A_30_78#_c_1583_n 2.20311e-19 $X=0.945 $Y=2.465 $X2=0
+ $Y2=0
cc_397 N_RESET_B_M1018_g N_A_30_78#_c_1577_n 0.00832998f $X=0.9 $Y=0.6 $X2=0
+ $Y2=0
cc_398 N_RESET_B_c_278_n N_A_30_78#_c_1577_n 0.011603f $X=1.055 $Y=1.92 $X2=0
+ $Y2=0
cc_399 N_RESET_B_c_286_n N_A_30_78#_c_1577_n 0.00422544f $X=0.945 $Y=2.375 $X2=0
+ $Y2=0
cc_400 N_RESET_B_c_293_n N_A_30_78#_c_1577_n 0.00138196f $X=1.345 $Y=2.035 $X2=0
+ $Y2=0
cc_401 N_RESET_B_c_283_n N_A_30_78#_c_1577_n 0.0048756f $X=1.12 $Y=1.305 $X2=0
+ $Y2=0
cc_402 N_RESET_B_c_284_n N_A_30_78#_c_1577_n 0.0697209f $X=1.12 $Y=1.305 $X2=0
+ $Y2=0
cc_403 N_RESET_B_c_299_n N_A_30_78#_c_1577_n 0.0049908f $X=1.12 $Y=1.985 $X2=0
+ $Y2=0
cc_404 N_RESET_B_c_286_n N_A_30_78#_c_1585_n 0.00991629f $X=0.945 $Y=2.375 $X2=0
+ $Y2=0
cc_405 N_RESET_B_c_287_n N_A_30_78#_c_1585_n 0.00910119f $X=0.945 $Y=2.465 $X2=0
+ $Y2=0
cc_406 N_RESET_B_c_292_n N_A_30_78#_c_1585_n 0.0343847f $X=4.895 $Y=2.035 $X2=0
+ $Y2=0
cc_407 N_RESET_B_c_293_n N_A_30_78#_c_1585_n 0.00463734f $X=1.345 $Y=2.035 $X2=0
+ $Y2=0
cc_408 N_RESET_B_c_284_n N_A_30_78#_c_1585_n 0.0184055f $X=1.12 $Y=1.305 $X2=0
+ $Y2=0
cc_409 N_RESET_B_c_299_n N_A_30_78#_c_1585_n 0.00267437f $X=1.12 $Y=1.985 $X2=0
+ $Y2=0
cc_410 N_RESET_B_c_292_n N_A_30_78#_c_1586_n 0.0179572f $X=4.895 $Y=2.035 $X2=0
+ $Y2=0
cc_411 N_RESET_B_c_292_n N_A_30_78#_c_1579_n 0.0103822f $X=4.895 $Y=2.035 $X2=0
+ $Y2=0
cc_412 N_RESET_B_M1018_g N_A_30_78#_c_1580_n 9.29579e-19 $X=0.9 $Y=0.6 $X2=0
+ $Y2=0
cc_413 N_RESET_B_c_292_n N_A_30_78#_c_1588_n 0.0132505f $X=4.895 $Y=2.035 $X2=0
+ $Y2=0
cc_414 N_RESET_B_c_292_n N_A_30_78#_c_1581_n 0.00392675f $X=4.895 $Y=2.035 $X2=0
+ $Y2=0
cc_415 N_RESET_B_M1018_g N_VGND_c_1714_n 0.0060384f $X=0.9 $Y=0.6 $X2=0 $Y2=0
cc_416 N_RESET_B_c_283_n N_VGND_c_1714_n 0.00180633f $X=1.12 $Y=1.305 $X2=0
+ $Y2=0
cc_417 N_RESET_B_c_284_n N_VGND_c_1714_n 0.0140897f $X=1.12 $Y=1.305 $X2=0 $Y2=0
cc_418 N_RESET_B_M1023_g N_VGND_c_1716_n 0.0104625f $X=8.24 $Y=0.615 $X2=0 $Y2=0
cc_419 N_RESET_B_M1018_g N_VGND_c_1721_n 0.00554804f $X=0.9 $Y=0.6 $X2=0 $Y2=0
cc_420 N_RESET_B_c_279_n N_VGND_c_1724_n 0.00296023f $X=4.79 $Y=1.185 $X2=0
+ $Y2=0
cc_421 N_RESET_B_M1023_g N_VGND_c_1726_n 0.0045897f $X=8.24 $Y=0.615 $X2=0 $Y2=0
cc_422 N_RESET_B_M1018_g N_VGND_c_1733_n 0.00539454f $X=0.9 $Y=0.6 $X2=0 $Y2=0
cc_423 N_RESET_B_c_279_n N_VGND_c_1733_n 0.00451834f $X=4.79 $Y=1.185 $X2=0
+ $Y2=0
cc_424 N_RESET_B_M1023_g N_VGND_c_1733_n 0.0044912f $X=8.24 $Y=0.615 $X2=0 $Y2=0
cc_425 CLK N_A_490_362#_c_515_n 8.33146e-19 $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_426 CLK N_A_490_362#_c_532_n 0.00810223f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_427 N_CLK_c_468_n N_A_306_74#_c_918_n 0.0412216f $X=1.925 $Y=1.735 $X2=0
+ $Y2=0
cc_428 CLK N_A_306_74#_c_918_n 4.04145e-19 $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_429 N_CLK_M1000_g N_A_306_74#_c_906_n 0.0213925f $X=1.89 $Y=0.74 $X2=0 $Y2=0
cc_430 N_CLK_M1000_g N_A_306_74#_c_911_n 0.00560421f $X=1.89 $Y=0.74 $X2=0 $Y2=0
cc_431 N_CLK_c_468_n N_A_306_74#_c_911_n 0.0213181f $X=1.925 $Y=1.735 $X2=0
+ $Y2=0
cc_432 CLK N_A_306_74#_c_911_n 0.00498195f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_433 N_CLK_c_468_n N_A_306_74#_c_929_n 0.0035155f $X=1.925 $Y=1.735 $X2=0
+ $Y2=0
cc_434 N_CLK_M1000_g N_A_306_74#_c_912_n 0.0101416f $X=1.89 $Y=0.74 $X2=0 $Y2=0
cc_435 N_CLK_M1000_g N_A_306_74#_c_913_n 0.00380568f $X=1.89 $Y=0.74 $X2=0 $Y2=0
cc_436 N_CLK_c_468_n N_A_306_74#_c_913_n 0.00515722f $X=1.925 $Y=1.735 $X2=0
+ $Y2=0
cc_437 CLK N_A_306_74#_c_913_n 0.0310013f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_438 N_CLK_M1000_g N_A_306_74#_c_914_n 0.0117933f $X=1.89 $Y=0.74 $X2=0 $Y2=0
cc_439 N_CLK_c_468_n N_A_306_74#_c_914_n 7.71729e-19 $X=1.925 $Y=1.735 $X2=0
+ $Y2=0
cc_440 CLK N_A_306_74#_c_914_n 0.0336655f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_441 N_CLK_M1000_g N_A_306_74#_c_915_n 7.82053e-19 $X=1.89 $Y=0.74 $X2=0 $Y2=0
cc_442 CLK N_A_306_74#_c_915_n 0.0184742f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_443 N_CLK_M1000_g N_A_306_74#_c_917_n 0.00151623f $X=1.89 $Y=0.74 $X2=0 $Y2=0
cc_444 N_CLK_c_468_n N_A_306_74#_c_917_n 0.00166711f $X=1.925 $Y=1.735 $X2=0
+ $Y2=0
cc_445 CLK N_A_306_74#_c_917_n 0.00370093f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_446 N_CLK_c_468_n N_A_306_74#_c_934_n 0.00728418f $X=1.925 $Y=1.735 $X2=0
+ $Y2=0
cc_447 CLK N_A_306_74#_c_934_n 0.00282549f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_448 N_CLK_c_468_n N_VPWR_c_1429_n 0.00650304f $X=1.925 $Y=1.735 $X2=0 $Y2=0
cc_449 N_CLK_c_468_n N_VPWR_c_1430_n 0.0105859f $X=1.925 $Y=1.735 $X2=0 $Y2=0
cc_450 N_CLK_c_468_n N_VPWR_c_1442_n 0.0049908f $X=1.925 $Y=1.735 $X2=0 $Y2=0
cc_451 N_CLK_c_468_n N_VPWR_c_1426_n 0.00486206f $X=1.925 $Y=1.735 $X2=0 $Y2=0
cc_452 N_CLK_c_468_n N_A_30_78#_c_1585_n 0.0155818f $X=1.925 $Y=1.735 $X2=0
+ $Y2=0
cc_453 CLK N_A_30_78#_c_1585_n 0.00451498f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_454 N_CLK_M1000_g N_VGND_c_1714_n 0.00342433f $X=1.89 $Y=0.74 $X2=0 $Y2=0
cc_455 N_CLK_M1000_g N_VGND_c_1715_n 0.00604382f $X=1.89 $Y=0.74 $X2=0 $Y2=0
cc_456 N_CLK_M1000_g N_VGND_c_1723_n 0.00434272f $X=1.89 $Y=0.74 $X2=0 $Y2=0
cc_457 N_CLK_M1000_g N_VGND_c_1733_n 0.00826311f $X=1.89 $Y=0.74 $X2=0 $Y2=0
cc_458 N_A_490_362#_c_518_n N_A_837_359#_M1025_d 0.00224297f $X=7.285 $Y=0.34
+ $X2=-0.19 $Y2=-0.245
cc_459 N_A_490_362#_c_536_n N_A_837_359#_c_708_n 0.00414301f $X=3.33 $Y=1.65
+ $X2=0 $Y2=0
cc_460 N_A_490_362#_c_510_n N_A_837_359#_M1015_g 0.00574235f $X=4.01 $Y=1.405
+ $X2=0 $Y2=0
cc_461 N_A_490_362#_M1028_g N_A_837_359#_M1015_g 0.0529896f $X=4.01 $Y=0.9 $X2=0
+ $Y2=0
cc_462 N_A_490_362#_c_517_n N_A_837_359#_M1015_g 0.00376198f $X=5.515 $Y=0.7
+ $X2=0 $Y2=0
cc_463 N_A_490_362#_c_523_n N_A_837_359#_M1015_g 0.00825047f $X=4.355 $Y=0.415
+ $X2=0 $Y2=0
cc_464 N_A_490_362#_c_510_n N_A_837_359#_c_704_n 4.1994e-19 $X=4.01 $Y=1.405
+ $X2=0 $Y2=0
cc_465 N_A_490_362#_M1028_g N_A_837_359#_c_704_n 0.00126199f $X=4.01 $Y=0.9
+ $X2=0 $Y2=0
cc_466 N_A_490_362#_c_517_n N_A_837_359#_c_705_n 0.0769509f $X=5.515 $Y=0.7
+ $X2=0 $Y2=0
cc_467 N_A_490_362#_c_518_n N_A_837_359#_c_705_n 0.00332639f $X=7.285 $Y=0.34
+ $X2=0 $Y2=0
cc_468 N_A_490_362#_c_517_n N_A_837_359#_c_734_n 3.80876e-19 $X=5.515 $Y=0.7
+ $X2=0 $Y2=0
cc_469 N_A_490_362#_c_523_n N_A_837_359#_c_734_n 0.00936402f $X=4.355 $Y=0.415
+ $X2=0 $Y2=0
cc_470 N_A_490_362#_c_518_n N_A_837_359#_c_736_n 0.0176299f $X=7.285 $Y=0.34
+ $X2=0 $Y2=0
cc_471 N_A_490_362#_c_514_n N_A_837_359#_c_711_n 0.00325656f $X=6.355 $Y=1.27
+ $X2=0 $Y2=0
cc_472 N_A_490_362#_c_512_n N_A_837_359#_c_706_n 4.62933e-19 $X=6.28 $Y=1.195
+ $X2=0 $Y2=0
cc_473 N_A_490_362#_c_512_n N_A_837_359#_c_707_n 0.00207614f $X=6.28 $Y=1.195
+ $X2=0 $Y2=0
cc_474 N_A_490_362#_c_512_n N_A_696_457#_M1025_g 0.0126968f $X=6.28 $Y=1.195
+ $X2=0 $Y2=0
cc_475 N_A_490_362#_c_518_n N_A_696_457#_M1025_g 0.0119914f $X=7.285 $Y=0.34
+ $X2=0 $Y2=0
cc_476 N_A_490_362#_c_514_n N_A_696_457#_c_786_n 0.0126968f $X=6.355 $Y=1.27
+ $X2=0 $Y2=0
cc_477 N_A_490_362#_c_526_n N_A_696_457#_c_788_n 6.06282e-19 $X=3.405 $Y=2.12
+ $X2=0 $Y2=0
cc_478 N_A_490_362#_c_510_n N_A_696_457#_c_788_n 0.0118046f $X=4.01 $Y=1.405
+ $X2=0 $Y2=0
cc_479 N_A_490_362#_M1028_g N_A_696_457#_c_788_n 0.00867235f $X=4.01 $Y=0.9
+ $X2=0 $Y2=0
cc_480 N_A_490_362#_c_527_n N_A_696_457#_c_795_n 0.00382922f $X=3.405 $Y=2.21
+ $X2=0 $Y2=0
cc_481 N_A_490_362#_c_528_n N_A_696_457#_c_795_n 0.00107261f $X=3.825 $Y=1.65
+ $X2=0 $Y2=0
cc_482 N_A_490_362#_c_528_n N_A_696_457#_c_791_n 0.00172887f $X=3.825 $Y=1.65
+ $X2=0 $Y2=0
cc_483 N_A_490_362#_c_510_n N_A_696_457#_c_791_n 0.0027075f $X=4.01 $Y=1.405
+ $X2=0 $Y2=0
cc_484 N_A_490_362#_M1028_g N_A_696_457#_c_791_n 0.00834631f $X=4.01 $Y=0.9
+ $X2=0 $Y2=0
cc_485 N_A_490_362#_c_516_n N_A_696_457#_c_791_n 0.035372f $X=4.27 $Y=0.415
+ $X2=0 $Y2=0
cc_486 N_A_490_362#_c_523_n N_A_696_457#_c_791_n 0.00147443f $X=4.355 $Y=0.415
+ $X2=0 $Y2=0
cc_487 N_A_490_362#_c_532_n N_A_306_74#_c_918_n 0.00455959f $X=3.04 $Y=1.74
+ $X2=0 $Y2=0
cc_488 N_A_490_362#_c_515_n N_A_306_74#_c_906_n 0.0057867f $X=2.955 $Y=1.575
+ $X2=0 $Y2=0
cc_489 N_A_490_362#_c_516_n N_A_306_74#_c_906_n 2.18663e-19 $X=4.27 $Y=0.415
+ $X2=0 $Y2=0
cc_490 N_A_490_362#_c_522_n N_A_306_74#_c_906_n 0.00762002f $X=2.775 $Y=0.415
+ $X2=0 $Y2=0
cc_491 N_A_490_362#_c_515_n N_A_306_74#_c_907_n 0.0133199f $X=2.955 $Y=1.575
+ $X2=0 $Y2=0
cc_492 N_A_490_362#_c_516_n N_A_306_74#_c_907_n 0.00379441f $X=4.27 $Y=0.415
+ $X2=0 $Y2=0
cc_493 N_A_490_362#_c_532_n N_A_306_74#_c_907_n 3.01079e-19 $X=3.04 $Y=1.74
+ $X2=0 $Y2=0
cc_494 N_A_490_362#_c_533_n N_A_306_74#_c_907_n 0.00480721f $X=3.33 $Y=1.74
+ $X2=0 $Y2=0
cc_495 N_A_490_362#_c_536_n N_A_306_74#_c_907_n 0.0225427f $X=3.33 $Y=1.65 $X2=0
+ $Y2=0
cc_496 N_A_490_362#_c_526_n N_A_306_74#_c_919_n 0.0100809f $X=3.405 $Y=2.12
+ $X2=0 $Y2=0
cc_497 N_A_490_362#_c_527_n N_A_306_74#_c_919_n 0.0123572f $X=3.405 $Y=2.21
+ $X2=0 $Y2=0
cc_498 N_A_490_362#_c_532_n N_A_306_74#_c_919_n 0.0172745f $X=3.04 $Y=1.74 $X2=0
+ $Y2=0
cc_499 N_A_490_362#_c_527_n N_A_306_74#_c_920_n 0.00899632f $X=3.405 $Y=2.21
+ $X2=0 $Y2=0
cc_500 N_A_490_362#_M1028_g N_A_306_74#_c_908_n 0.0184281f $X=4.01 $Y=0.9 $X2=0
+ $Y2=0
cc_501 N_A_490_362#_c_516_n N_A_306_74#_c_908_n 0.00661564f $X=4.27 $Y=0.415
+ $X2=0 $Y2=0
cc_502 N_A_490_362#_c_522_n N_A_306_74#_c_908_n 0.00456341f $X=2.775 $Y=0.415
+ $X2=0 $Y2=0
cc_503 N_A_490_362#_c_527_n N_A_306_74#_c_922_n 0.00278823f $X=3.405 $Y=2.21
+ $X2=0 $Y2=0
cc_504 N_A_490_362#_c_527_n N_A_306_74#_c_924_n 0.0102684f $X=3.405 $Y=2.21
+ $X2=0 $Y2=0
cc_505 N_A_490_362#_c_528_n N_A_306_74#_c_924_n 0.00467333f $X=3.825 $Y=1.65
+ $X2=0 $Y2=0
cc_506 N_A_490_362#_c_535_n N_A_306_74#_M1021_g 0.00727778f $X=7.12 $Y=2.14
+ $X2=0 $Y2=0
cc_507 N_A_490_362#_c_513_n N_A_306_74#_c_909_n 0.0196921f $X=6.715 $Y=1.27
+ $X2=0 $Y2=0
cc_508 N_A_490_362#_c_520_n N_A_306_74#_c_909_n 0.0166975f $X=7.12 $Y=2.14 $X2=0
+ $Y2=0
cc_509 N_A_490_362#_c_535_n N_A_306_74#_c_909_n 0.0260156f $X=7.12 $Y=2.14 $X2=0
+ $Y2=0
cc_510 N_A_490_362#_c_525_n N_A_306_74#_c_909_n 0.00239794f $X=7.37 $Y=1.18
+ $X2=0 $Y2=0
cc_511 N_A_490_362#_c_514_n N_A_306_74#_c_928_n 0.0196921f $X=6.355 $Y=1.27
+ $X2=0 $Y2=0
cc_512 N_A_490_362#_c_518_n N_A_306_74#_M1032_g 0.00912173f $X=7.285 $Y=0.34
+ $X2=0 $Y2=0
cc_513 N_A_490_362#_c_520_n N_A_306_74#_M1032_g 0.00885461f $X=7.12 $Y=2.14
+ $X2=0 $Y2=0
cc_514 N_A_490_362#_c_521_n N_A_306_74#_M1032_g 0.0230685f $X=7.37 $Y=1.015
+ $X2=0 $Y2=0
cc_515 N_A_490_362#_c_524_n N_A_306_74#_M1032_g 0.0213806f $X=6.88 $Y=1.18 $X2=0
+ $Y2=0
cc_516 N_A_490_362#_c_525_n N_A_306_74#_M1032_g 0.0123873f $X=7.37 $Y=1.18 $X2=0
+ $Y2=0
cc_517 N_A_490_362#_c_522_n N_A_306_74#_c_911_n 0.00584739f $X=2.775 $Y=0.415
+ $X2=0 $Y2=0
cc_518 N_A_490_362#_c_532_n N_A_306_74#_c_929_n 0.0181729f $X=3.04 $Y=1.74 $X2=0
+ $Y2=0
cc_519 N_A_490_362#_c_536_n N_A_306_74#_c_929_n 0.0214218f $X=3.33 $Y=1.65 $X2=0
+ $Y2=0
cc_520 N_A_490_362#_M1019_d N_A_306_74#_c_914_n 0.00261988f $X=2.535 $Y=0.37
+ $X2=0 $Y2=0
cc_521 N_A_490_362#_c_515_n N_A_306_74#_c_914_n 0.0141274f $X=2.955 $Y=1.575
+ $X2=0 $Y2=0
cc_522 N_A_490_362#_c_522_n N_A_306_74#_c_914_n 0.0112799f $X=2.775 $Y=0.415
+ $X2=0 $Y2=0
cc_523 N_A_490_362#_c_515_n N_A_306_74#_c_915_n 0.0289853f $X=2.955 $Y=1.575
+ $X2=0 $Y2=0
cc_524 N_A_490_362#_c_532_n N_A_306_74#_c_915_n 0.0137243f $X=3.04 $Y=1.74 $X2=0
+ $Y2=0
cc_525 N_A_490_362#_c_515_n N_A_306_74#_c_916_n 0.00149416f $X=2.955 $Y=1.575
+ $X2=0 $Y2=0
cc_526 N_A_490_362#_c_532_n N_A_306_74#_c_934_n 0.00600724f $X=3.04 $Y=1.74
+ $X2=0 $Y2=0
cc_527 N_A_490_362#_c_518_n N_A_1525_212#_M1010_g 0.00108131f $X=7.285 $Y=0.34
+ $X2=0 $Y2=0
cc_528 N_A_490_362#_c_521_n N_A_1525_212#_M1010_g 0.00485618f $X=7.37 $Y=1.015
+ $X2=0 $Y2=0
cc_529 N_A_490_362#_c_525_n N_A_1525_212#_M1010_g 0.00116217f $X=7.37 $Y=1.18
+ $X2=0 $Y2=0
cc_530 N_A_490_362#_c_535_n N_A_1525_212#_c_1097_n 0.0212062f $X=7.12 $Y=2.14
+ $X2=0 $Y2=0
cc_531 N_A_490_362#_c_530_n N_A_1525_212#_c_1099_n 0.0268843f $X=7.315 $Y=2.39
+ $X2=0 $Y2=0
cc_532 N_A_490_362#_c_520_n N_A_1525_212#_c_1089_n 9.8351e-19 $X=7.12 $Y=2.14
+ $X2=0 $Y2=0
cc_533 N_A_490_362#_c_520_n N_A_1525_212#_c_1094_n 0.00193736f $X=7.12 $Y=2.14
+ $X2=0 $Y2=0
cc_534 N_A_490_362#_c_525_n N_A_1525_212#_c_1094_n 0.0239506f $X=7.37 $Y=1.18
+ $X2=0 $Y2=0
cc_535 N_A_490_362#_c_525_n N_A_1525_212#_c_1095_n 0.00177987f $X=7.37 $Y=1.18
+ $X2=0 $Y2=0
cc_536 N_A_490_362#_c_518_n N_A_1271_74#_M1003_d 0.00941894f $X=7.285 $Y=0.34
+ $X2=-0.19 $Y2=-0.245
cc_537 N_A_490_362#_c_518_n N_A_1271_74#_c_1249_n 0.00860077f $X=7.285 $Y=0.34
+ $X2=0 $Y2=0
cc_538 N_A_490_362#_c_512_n N_A_1271_74#_c_1211_n 0.0041612f $X=6.28 $Y=1.195
+ $X2=0 $Y2=0
cc_539 N_A_490_362#_c_513_n N_A_1271_74#_c_1211_n 0.010955f $X=6.715 $Y=1.27
+ $X2=0 $Y2=0
cc_540 N_A_490_362#_c_520_n N_A_1271_74#_c_1211_n 0.00709969f $X=7.12 $Y=2.14
+ $X2=0 $Y2=0
cc_541 N_A_490_362#_c_524_n N_A_1271_74#_c_1211_n 0.00131723f $X=6.88 $Y=1.18
+ $X2=0 $Y2=0
cc_542 N_A_490_362#_c_525_n N_A_1271_74#_c_1211_n 0.022475f $X=7.37 $Y=1.18
+ $X2=0 $Y2=0
cc_543 N_A_490_362#_c_530_n N_A_1271_74#_c_1223_n 0.00181181f $X=7.315 $Y=2.39
+ $X2=0 $Y2=0
cc_544 N_A_490_362#_c_520_n N_A_1271_74#_c_1223_n 0.0315385f $X=7.12 $Y=2.14
+ $X2=0 $Y2=0
cc_545 N_A_490_362#_c_535_n N_A_1271_74#_c_1223_n 0.00442904f $X=7.12 $Y=2.14
+ $X2=0 $Y2=0
cc_546 N_A_490_362#_c_513_n N_A_1271_74#_c_1212_n 0.00400734f $X=6.715 $Y=1.27
+ $X2=0 $Y2=0
cc_547 N_A_490_362#_c_518_n N_A_1271_74#_c_1212_n 0.0414158f $X=7.285 $Y=0.34
+ $X2=0 $Y2=0
cc_548 N_A_490_362#_c_521_n N_A_1271_74#_c_1212_n 0.0196081f $X=7.37 $Y=1.015
+ $X2=0 $Y2=0
cc_549 N_A_490_362#_c_524_n N_A_1271_74#_c_1212_n 0.00763158f $X=6.88 $Y=1.18
+ $X2=0 $Y2=0
cc_550 N_A_490_362#_c_525_n N_A_1271_74#_c_1212_n 0.0304853f $X=7.37 $Y=1.18
+ $X2=0 $Y2=0
cc_551 N_A_490_362#_c_530_n N_A_1271_74#_c_1237_n 0.0126686f $X=7.315 $Y=2.39
+ $X2=0 $Y2=0
cc_552 N_A_490_362#_c_520_n N_A_1271_74#_c_1237_n 0.0234051f $X=7.12 $Y=2.14
+ $X2=0 $Y2=0
cc_553 N_A_490_362#_c_535_n N_A_1271_74#_c_1237_n 0.00188634f $X=7.12 $Y=2.14
+ $X2=0 $Y2=0
cc_554 N_A_490_362#_c_530_n N_A_1271_74#_c_1224_n 0.00196844f $X=7.315 $Y=2.39
+ $X2=0 $Y2=0
cc_555 N_A_490_362#_c_520_n N_A_1271_74#_c_1224_n 0.0428804f $X=7.12 $Y=2.14
+ $X2=0 $Y2=0
cc_556 N_A_490_362#_c_535_n N_A_1271_74#_c_1224_n 0.00431063f $X=7.12 $Y=2.14
+ $X2=0 $Y2=0
cc_557 N_A_490_362#_c_520_n N_A_1271_74#_c_1214_n 0.0142968f $X=7.12 $Y=2.14
+ $X2=0 $Y2=0
cc_558 N_A_490_362#_c_513_n N_A_1271_74#_c_1215_n 0.00176995f $X=6.715 $Y=1.27
+ $X2=0 $Y2=0
cc_559 N_A_490_362#_c_520_n N_A_1271_74#_c_1215_n 0.00932939f $X=7.12 $Y=2.14
+ $X2=0 $Y2=0
cc_560 N_A_490_362#_c_530_n N_VPWR_c_1434_n 0.00125875f $X=7.315 $Y=2.39 $X2=0
+ $Y2=0
cc_561 N_A_490_362#_c_530_n N_VPWR_c_1444_n 0.00391396f $X=7.315 $Y=2.39 $X2=0
+ $Y2=0
cc_562 N_A_490_362#_c_527_n N_VPWR_c_1426_n 9.49986e-19 $X=3.405 $Y=2.21 $X2=0
+ $Y2=0
cc_563 N_A_490_362#_c_530_n N_VPWR_c_1426_n 0.0052212f $X=7.315 $Y=2.39 $X2=0
+ $Y2=0
cc_564 N_A_490_362#_M1012_d N_A_30_78#_c_1585_n 0.00657073f $X=2.45 $Y=1.81
+ $X2=0 $Y2=0
cc_565 N_A_490_362#_c_532_n N_A_30_78#_c_1585_n 0.0247894f $X=3.04 $Y=1.74 $X2=0
+ $Y2=0
cc_566 N_A_490_362#_M1028_g N_A_30_78#_c_1578_n 2.83252e-19 $X=4.01 $Y=0.9 $X2=0
+ $Y2=0
cc_567 N_A_490_362#_c_516_n N_A_30_78#_c_1578_n 0.0195048f $X=4.27 $Y=0.415
+ $X2=0 $Y2=0
cc_568 N_A_490_362#_c_522_n N_A_30_78#_c_1578_n 0.0437866f $X=2.775 $Y=0.415
+ $X2=0 $Y2=0
cc_569 N_A_490_362#_c_526_n N_A_30_78#_c_1586_n 0.00410538f $X=3.405 $Y=2.12
+ $X2=0 $Y2=0
cc_570 N_A_490_362#_c_527_n N_A_30_78#_c_1586_n 0.0111572f $X=3.405 $Y=2.21
+ $X2=0 $Y2=0
cc_571 N_A_490_362#_c_528_n N_A_30_78#_c_1586_n 0.00164971f $X=3.825 $Y=1.65
+ $X2=0 $Y2=0
cc_572 N_A_490_362#_c_533_n N_A_30_78#_c_1586_n 0.0096674f $X=3.33 $Y=1.74 $X2=0
+ $Y2=0
cc_573 N_A_490_362#_c_536_n N_A_30_78#_c_1586_n 0.00109593f $X=3.33 $Y=1.65
+ $X2=0 $Y2=0
cc_574 N_A_490_362#_c_528_n N_A_30_78#_c_1579_n 0.0131253f $X=3.825 $Y=1.65
+ $X2=0 $Y2=0
cc_575 N_A_490_362#_c_510_n N_A_30_78#_c_1579_n 0.00406314f $X=4.01 $Y=1.405
+ $X2=0 $Y2=0
cc_576 N_A_490_362#_c_515_n N_A_30_78#_c_1579_n 0.00565517f $X=2.955 $Y=1.575
+ $X2=0 $Y2=0
cc_577 N_A_490_362#_c_533_n N_A_30_78#_c_1579_n 0.025441f $X=3.33 $Y=1.74 $X2=0
+ $Y2=0
cc_578 N_A_490_362#_c_536_n N_A_30_78#_c_1579_n 0.00717136f $X=3.33 $Y=1.65
+ $X2=0 $Y2=0
cc_579 N_A_490_362#_c_527_n N_A_30_78#_c_1588_n 0.00342386f $X=3.405 $Y=2.21
+ $X2=0 $Y2=0
cc_580 N_A_490_362#_c_532_n N_A_30_78#_c_1588_n 0.00323073f $X=3.04 $Y=1.74
+ $X2=0 $Y2=0
cc_581 N_A_490_362#_c_533_n N_A_30_78#_c_1588_n 0.0128199f $X=3.33 $Y=1.74 $X2=0
+ $Y2=0
cc_582 N_A_490_362#_c_536_n N_A_30_78#_c_1588_n 0.00222816f $X=3.33 $Y=1.65
+ $X2=0 $Y2=0
cc_583 N_A_490_362#_c_528_n N_A_30_78#_c_1581_n 8.36337e-19 $X=3.825 $Y=1.65
+ $X2=0 $Y2=0
cc_584 N_A_490_362#_M1028_g N_A_30_78#_c_1581_n 9.3084e-19 $X=4.01 $Y=0.9 $X2=0
+ $Y2=0
cc_585 N_A_490_362#_c_515_n N_A_30_78#_c_1581_n 0.0131356f $X=2.955 $Y=1.575
+ $X2=0 $Y2=0
cc_586 N_A_490_362#_c_533_n N_A_30_78#_c_1581_n 0.0153344f $X=3.33 $Y=1.74 $X2=0
+ $Y2=0
cc_587 N_A_490_362#_c_536_n N_A_30_78#_c_1581_n 0.00315825f $X=3.33 $Y=1.65
+ $X2=0 $Y2=0
cc_588 N_A_490_362#_c_517_n N_VGND_M1001_d 0.0203479f $X=5.515 $Y=0.7 $X2=0
+ $Y2=0
cc_589 N_A_490_362#_c_543_n N_VGND_M1001_d 0.00595426f $X=5.6 $Y=0.615 $X2=0
+ $Y2=0
cc_590 N_A_490_362#_c_519_n N_VGND_M1001_d 7.1669e-19 $X=5.685 $Y=0.34 $X2=0
+ $Y2=0
cc_591 N_A_490_362#_c_522_n N_VGND_c_1715_n 0.0209866f $X=2.775 $Y=0.415 $X2=0
+ $Y2=0
cc_592 N_A_490_362#_c_518_n N_VGND_c_1716_n 0.00865667f $X=7.285 $Y=0.34 $X2=0
+ $Y2=0
cc_593 N_A_490_362#_c_516_n N_VGND_c_1724_n 0.0538921f $X=4.27 $Y=0.415 $X2=0
+ $Y2=0
cc_594 N_A_490_362#_c_517_n N_VGND_c_1724_n 0.0408763f $X=5.515 $Y=0.7 $X2=0
+ $Y2=0
cc_595 N_A_490_362#_c_543_n N_VGND_c_1724_n 0.00152296f $X=5.6 $Y=0.615 $X2=0
+ $Y2=0
cc_596 N_A_490_362#_c_519_n N_VGND_c_1724_n 0.0151294f $X=5.685 $Y=0.34 $X2=0
+ $Y2=0
cc_597 N_A_490_362#_c_522_n N_VGND_c_1724_n 0.0251053f $X=2.775 $Y=0.415 $X2=0
+ $Y2=0
cc_598 N_A_490_362#_c_523_n N_VGND_c_1724_n 0.0124546f $X=4.355 $Y=0.415 $X2=0
+ $Y2=0
cc_599 N_A_490_362#_c_512_n N_VGND_c_1725_n 0.00278271f $X=6.28 $Y=1.195 $X2=0
+ $Y2=0
cc_600 N_A_490_362#_c_517_n N_VGND_c_1725_n 0.00309688f $X=5.515 $Y=0.7 $X2=0
+ $Y2=0
cc_601 N_A_490_362#_c_518_n N_VGND_c_1725_n 0.114324f $X=7.285 $Y=0.34 $X2=0
+ $Y2=0
cc_602 N_A_490_362#_c_519_n N_VGND_c_1725_n 0.0119604f $X=5.685 $Y=0.34 $X2=0
+ $Y2=0
cc_603 N_A_490_362#_c_512_n N_VGND_c_1733_n 0.00358928f $X=6.28 $Y=1.195 $X2=0
+ $Y2=0
cc_604 N_A_490_362#_c_516_n N_VGND_c_1733_n 0.044091f $X=4.27 $Y=0.415 $X2=0
+ $Y2=0
cc_605 N_A_490_362#_c_517_n N_VGND_c_1733_n 0.0207117f $X=5.515 $Y=0.7 $X2=0
+ $Y2=0
cc_606 N_A_490_362#_c_518_n N_VGND_c_1733_n 0.0653925f $X=7.285 $Y=0.34 $X2=0
+ $Y2=0
cc_607 N_A_490_362#_c_519_n N_VGND_c_1733_n 0.00656672f $X=5.685 $Y=0.34 $X2=0
+ $Y2=0
cc_608 N_A_490_362#_c_522_n N_VGND_c_1733_n 0.0194694f $X=2.775 $Y=0.415 $X2=0
+ $Y2=0
cc_609 N_A_490_362#_c_523_n N_VGND_c_1733_n 0.00619879f $X=4.355 $Y=0.415 $X2=0
+ $Y2=0
cc_610 N_A_490_362#_c_517_n A_895_138# 0.00134267f $X=5.515 $Y=0.7 $X2=-0.19
+ $Y2=-0.245
cc_611 N_A_837_359#_c_705_n N_A_696_457#_M1025_g 0.0124697f $X=5.855 $Y=1.04
+ $X2=0 $Y2=0
cc_612 N_A_837_359#_c_736_n N_A_696_457#_M1025_g 0.0104935f $X=6.02 $Y=0.86
+ $X2=0 $Y2=0
cc_613 N_A_837_359#_c_706_n N_A_696_457#_M1025_g 0.00268294f $X=6.02 $Y=1.042
+ $X2=0 $Y2=0
cc_614 N_A_837_359#_c_707_n N_A_696_457#_M1025_g 0.00639735f $X=6.18 $Y=1.855
+ $X2=0 $Y2=0
cc_615 N_A_837_359#_c_706_n N_A_696_457#_c_786_n 0.00463727f $X=6.02 $Y=1.042
+ $X2=0 $Y2=0
cc_616 N_A_837_359#_c_707_n N_A_696_457#_c_786_n 0.0148463f $X=6.18 $Y=1.855
+ $X2=0 $Y2=0
cc_617 N_A_837_359#_c_705_n N_A_696_457#_c_787_n 0.0091182f $X=5.855 $Y=1.04
+ $X2=0 $Y2=0
cc_618 N_A_837_359#_c_708_n N_A_696_457#_c_788_n 0.0069306f $X=4.275 $Y=2.21
+ $X2=0 $Y2=0
cc_619 N_A_837_359#_M1015_g N_A_696_457#_c_788_n 0.00213788f $X=4.4 $Y=0.9 $X2=0
+ $Y2=0
cc_620 N_A_837_359#_c_704_n N_A_696_457#_c_788_n 0.0736091f $X=4.36 $Y=1.96
+ $X2=0 $Y2=0
cc_621 N_A_837_359#_c_734_n N_A_696_457#_c_788_n 0.00118204f $X=4.445 $Y=1.04
+ $X2=0 $Y2=0
cc_622 N_A_837_359#_c_708_n N_A_696_457#_c_803_n 0.0158089f $X=4.275 $Y=2.21
+ $X2=0 $Y2=0
cc_623 N_A_837_359#_c_704_n N_A_696_457#_c_803_n 0.0065984f $X=4.36 $Y=1.96
+ $X2=0 $Y2=0
cc_624 N_A_837_359#_c_708_n N_A_696_457#_c_795_n 6.73983e-19 $X=4.275 $Y=2.21
+ $X2=0 $Y2=0
cc_625 N_A_837_359#_c_708_n N_A_696_457#_c_796_n 0.00400733f $X=4.275 $Y=2.21
+ $X2=0 $Y2=0
cc_626 N_A_837_359#_M1015_g N_A_696_457#_c_796_n 0.00140716f $X=4.4 $Y=0.9 $X2=0
+ $Y2=0
cc_627 N_A_837_359#_c_704_n N_A_696_457#_c_796_n 0.0386079f $X=4.36 $Y=1.96
+ $X2=0 $Y2=0
cc_628 N_A_837_359#_M1015_g N_A_696_457#_c_789_n 0.00201464f $X=4.4 $Y=0.9 $X2=0
+ $Y2=0
cc_629 N_A_837_359#_c_704_n N_A_696_457#_c_789_n 0.0226331f $X=4.36 $Y=1.96
+ $X2=0 $Y2=0
cc_630 N_A_837_359#_c_705_n N_A_696_457#_c_789_n 0.0137783f $X=5.855 $Y=1.04
+ $X2=0 $Y2=0
cc_631 N_A_837_359#_c_705_n N_A_696_457#_c_790_n 0.0680785f $X=5.855 $Y=1.04
+ $X2=0 $Y2=0
cc_632 N_A_837_359#_c_707_n N_A_696_457#_c_790_n 0.0134746f $X=6.18 $Y=1.855
+ $X2=0 $Y2=0
cc_633 N_A_837_359#_c_708_n N_A_696_457#_c_858_n 0.00105082f $X=4.275 $Y=2.21
+ $X2=0 $Y2=0
cc_634 N_A_837_359#_c_708_n N_A_306_74#_c_922_n 0.00284772f $X=4.275 $Y=2.21
+ $X2=0 $Y2=0
cc_635 N_A_837_359#_c_708_n N_A_306_74#_c_924_n 0.0271917f $X=4.275 $Y=2.21
+ $X2=0 $Y2=0
cc_636 N_A_837_359#_c_708_n N_A_306_74#_c_925_n 0.00850694f $X=4.275 $Y=2.21
+ $X2=0 $Y2=0
cc_637 N_A_837_359#_c_711_n N_A_306_74#_c_925_n 0.00434706f $X=6.18 $Y=2.02
+ $X2=0 $Y2=0
cc_638 N_A_837_359#_c_711_n N_A_306_74#_M1021_g 0.0106383f $X=6.18 $Y=2.02 $X2=0
+ $Y2=0
cc_639 N_A_837_359#_c_707_n N_A_306_74#_M1021_g 8.73808e-19 $X=6.18 $Y=1.855
+ $X2=0 $Y2=0
cc_640 N_A_837_359#_c_707_n N_A_306_74#_c_928_n 0.00135615f $X=6.18 $Y=1.855
+ $X2=0 $Y2=0
cc_641 N_A_837_359#_c_706_n N_A_1271_74#_c_1211_n 0.00157956f $X=6.02 $Y=1.042
+ $X2=0 $Y2=0
cc_642 N_A_837_359#_c_707_n N_A_1271_74#_c_1211_n 0.0283811f $X=6.18 $Y=1.855
+ $X2=0 $Y2=0
cc_643 N_A_837_359#_c_711_n N_A_1271_74#_c_1223_n 0.0250147f $X=6.18 $Y=2.02
+ $X2=0 $Y2=0
cc_644 N_A_837_359#_c_707_n N_A_1271_74#_c_1223_n 0.00658883f $X=6.18 $Y=1.855
+ $X2=0 $Y2=0
cc_645 N_A_837_359#_c_707_n N_A_1271_74#_c_1215_n 0.0129728f $X=6.18 $Y=1.855
+ $X2=0 $Y2=0
cc_646 N_A_837_359#_c_708_n N_VPWR_c_1431_n 0.00230854f $X=4.275 $Y=2.21 $X2=0
+ $Y2=0
cc_647 N_A_837_359#_c_705_n N_VPWR_c_1433_n 0.00367066f $X=5.855 $Y=1.04 $X2=0
+ $Y2=0
cc_648 N_A_837_359#_c_711_n N_VPWR_c_1433_n 0.0405057f $X=6.18 $Y=2.02 $X2=0
+ $Y2=0
cc_649 N_A_837_359#_c_711_n N_VPWR_c_1444_n 0.00666388f $X=6.18 $Y=2.02 $X2=0
+ $Y2=0
cc_650 N_A_837_359#_c_708_n N_VPWR_c_1426_n 9.49986e-19 $X=4.275 $Y=2.21 $X2=0
+ $Y2=0
cc_651 N_A_837_359#_c_711_n N_VPWR_c_1426_n 0.00905588f $X=6.18 $Y=2.02 $X2=0
+ $Y2=0
cc_652 N_A_837_359#_c_705_n N_VGND_M1001_d 0.0123032f $X=5.855 $Y=1.04 $X2=0
+ $Y2=0
cc_653 N_A_837_359#_M1015_g N_VGND_c_1724_n 0.00110839f $X=4.4 $Y=0.9 $X2=0
+ $Y2=0
cc_654 N_A_837_359#_M1015_g N_VGND_c_1733_n 0.0010844f $X=4.4 $Y=0.9 $X2=0 $Y2=0
cc_655 N_A_837_359#_c_705_n A_895_138# 0.00134267f $X=5.855 $Y=1.04 $X2=-0.19
+ $Y2=-0.245
cc_656 N_A_696_457#_c_788_n N_A_306_74#_c_907_n 2.17022e-19 $X=4.015 $Y=2.415
+ $X2=0 $Y2=0
cc_657 N_A_696_457#_c_795_n N_A_306_74#_c_920_n 0.0037146f $X=4.1 $Y=2.5 $X2=0
+ $Y2=0
cc_658 N_A_696_457#_c_788_n N_A_306_74#_c_908_n 0.00106324f $X=4.015 $Y=2.415
+ $X2=0 $Y2=0
cc_659 N_A_696_457#_c_791_n N_A_306_74#_c_908_n 0.00211731f $X=4.015 $Y=0.867
+ $X2=0 $Y2=0
cc_660 N_A_696_457#_c_795_n N_A_306_74#_c_922_n 4.94244e-19 $X=4.1 $Y=2.5 $X2=0
+ $Y2=0
cc_661 N_A_696_457#_c_788_n N_A_306_74#_c_924_n 0.00183744f $X=4.015 $Y=2.415
+ $X2=0 $Y2=0
cc_662 N_A_696_457#_c_795_n N_A_306_74#_c_924_n 0.0120063f $X=4.1 $Y=2.5 $X2=0
+ $Y2=0
cc_663 N_A_696_457#_c_786_n N_A_306_74#_c_925_n 0.0103562f $X=5.905 $Y=1.66
+ $X2=0 $Y2=0
cc_664 N_A_696_457#_c_803_n N_A_306_74#_c_925_n 0.00335096f $X=4.615 $Y=2.5
+ $X2=0 $Y2=0
cc_665 N_A_696_457#_c_795_n N_A_306_74#_c_925_n 0.00114785f $X=4.1 $Y=2.5 $X2=0
+ $Y2=0
cc_666 N_A_696_457#_c_798_n N_A_306_74#_c_925_n 0.00532011f $X=5.12 $Y=2.49
+ $X2=0 $Y2=0
cc_667 N_A_696_457#_c_858_n N_A_306_74#_c_925_n 0.00106642f $X=4.7 $Y=2.452
+ $X2=0 $Y2=0
cc_668 N_A_696_457#_c_786_n N_A_306_74#_M1021_g 0.0208385f $X=5.905 $Y=1.66
+ $X2=0 $Y2=0
cc_669 N_A_696_457#_c_786_n N_A_306_74#_c_928_n 0.0046962f $X=5.905 $Y=1.66
+ $X2=0 $Y2=0
cc_670 N_A_696_457#_c_803_n N_VPWR_M1027_d 0.00488949f $X=4.615 $Y=2.5 $X2=0
+ $Y2=0
cc_671 N_A_696_457#_c_796_n N_VPWR_M1027_d 4.72589e-19 $X=4.7 $Y=2.32 $X2=0
+ $Y2=0
cc_672 N_A_696_457#_c_858_n N_VPWR_M1027_d 0.00306384f $X=4.7 $Y=2.452 $X2=0
+ $Y2=0
cc_673 N_A_696_457#_c_803_n N_VPWR_c_1431_n 0.0152514f $X=4.615 $Y=2.5 $X2=0
+ $Y2=0
cc_674 N_A_696_457#_c_858_n N_VPWR_c_1431_n 0.0116304f $X=4.7 $Y=2.452 $X2=0
+ $Y2=0
cc_675 N_A_696_457#_c_798_n N_VPWR_c_1432_n 0.00636076f $X=5.12 $Y=2.49 $X2=0
+ $Y2=0
cc_676 N_A_696_457#_c_858_n N_VPWR_c_1432_n 3.55404e-19 $X=4.7 $Y=2.452 $X2=0
+ $Y2=0
cc_677 N_A_696_457#_c_786_n N_VPWR_c_1433_n 0.0144085f $X=5.905 $Y=1.66 $X2=0
+ $Y2=0
cc_678 N_A_696_457#_c_787_n N_VPWR_c_1433_n 0.00770753f $X=5.73 $Y=1.41 $X2=0
+ $Y2=0
cc_679 N_A_696_457#_c_790_n N_VPWR_c_1433_n 0.0131953f $X=5.52 $Y=1.41 $X2=0
+ $Y2=0
cc_680 N_A_696_457#_c_798_n N_VPWR_c_1433_n 0.018807f $X=5.12 $Y=2.49 $X2=0
+ $Y2=0
cc_681 N_A_696_457#_c_803_n N_VPWR_c_1443_n 0.00352361f $X=4.615 $Y=2.5 $X2=0
+ $Y2=0
cc_682 N_A_696_457#_c_795_n N_VPWR_c_1443_n 0.0105349f $X=4.1 $Y=2.5 $X2=0 $Y2=0
cc_683 N_A_696_457#_c_786_n N_VPWR_c_1426_n 8.51577e-19 $X=5.905 $Y=1.66 $X2=0
+ $Y2=0
cc_684 N_A_696_457#_c_803_n N_VPWR_c_1426_n 0.00773705f $X=4.615 $Y=2.5 $X2=0
+ $Y2=0
cc_685 N_A_696_457#_c_795_n N_VPWR_c_1426_n 0.0154763f $X=4.1 $Y=2.5 $X2=0 $Y2=0
cc_686 N_A_696_457#_c_798_n N_VPWR_c_1426_n 0.0112433f $X=5.12 $Y=2.49 $X2=0
+ $Y2=0
cc_687 N_A_696_457#_c_858_n N_VPWR_c_1426_n 0.00143814f $X=4.7 $Y=2.452 $X2=0
+ $Y2=0
cc_688 N_A_696_457#_c_788_n N_A_30_78#_c_1578_n 0.0049664f $X=4.015 $Y=2.415
+ $X2=0 $Y2=0
cc_689 N_A_696_457#_c_791_n N_A_30_78#_c_1578_n 0.014993f $X=4.015 $Y=0.867
+ $X2=0 $Y2=0
cc_690 N_A_696_457#_c_788_n N_A_30_78#_c_1586_n 0.0139725f $X=4.015 $Y=2.415
+ $X2=0 $Y2=0
cc_691 N_A_696_457#_c_795_n N_A_30_78#_c_1586_n 0.0194338f $X=4.1 $Y=2.5 $X2=0
+ $Y2=0
cc_692 N_A_696_457#_c_788_n N_A_30_78#_c_1579_n 0.0481207f $X=4.015 $Y=2.415
+ $X2=0 $Y2=0
cc_693 N_A_696_457#_c_788_n N_A_30_78#_c_1588_n 0.00310299f $X=4.015 $Y=2.415
+ $X2=0 $Y2=0
cc_694 N_A_696_457#_c_795_n N_A_30_78#_c_1588_n 0.0220686f $X=4.1 $Y=2.5 $X2=0
+ $Y2=0
cc_695 N_A_696_457#_c_788_n N_A_30_78#_c_1581_n 0.0139398f $X=4.015 $Y=2.415
+ $X2=0 $Y2=0
cc_696 N_A_696_457#_c_791_n N_A_30_78#_c_1581_n 0.00975559f $X=4.015 $Y=0.867
+ $X2=0 $Y2=0
cc_697 N_A_696_457#_c_788_n A_786_457# 0.00154981f $X=4.015 $Y=2.415 $X2=-0.19
+ $Y2=-0.245
cc_698 N_A_696_457#_c_803_n A_786_457# 0.00130488f $X=4.615 $Y=2.5 $X2=-0.19
+ $Y2=-0.245
cc_699 N_A_696_457#_c_795_n A_786_457# 0.00205983f $X=4.1 $Y=2.5 $X2=-0.19
+ $Y2=-0.245
cc_700 N_A_696_457#_M1025_g N_VGND_c_1724_n 0.0012551f $X=5.805 $Y=0.74 $X2=0
+ $Y2=0
cc_701 N_A_696_457#_M1025_g N_VGND_c_1725_n 0.00278271f $X=5.805 $Y=0.74 $X2=0
+ $Y2=0
cc_702 N_A_696_457#_M1025_g N_VGND_c_1733_n 0.00358928f $X=5.805 $Y=0.74 $X2=0
+ $Y2=0
cc_703 N_A_306_74#_M1032_g N_A_1525_212#_M1010_g 0.0390746f $X=7.33 $Y=0.615
+ $X2=0 $Y2=0
cc_704 N_A_306_74#_M1032_g N_A_1525_212#_c_1089_n 0.0184343f $X=7.33 $Y=0.615
+ $X2=0 $Y2=0
cc_705 N_A_306_74#_M1032_g N_A_1525_212#_c_1094_n 4.84439e-19 $X=7.33 $Y=0.615
+ $X2=0 $Y2=0
cc_706 N_A_306_74#_M1032_g N_A_1525_212#_c_1095_n 0.0192269f $X=7.33 $Y=0.615
+ $X2=0 $Y2=0
cc_707 N_A_306_74#_c_928_n N_A_1271_74#_c_1211_n 2.49182e-19 $X=6.485 $Y=1.66
+ $X2=0 $Y2=0
cc_708 N_A_306_74#_M1021_g N_A_1271_74#_c_1223_n 0.0101572f $X=6.41 $Y=2.31
+ $X2=0 $Y2=0
cc_709 N_A_306_74#_c_909_n N_A_1271_74#_c_1223_n 0.00688758f $X=7.255 $Y=1.66
+ $X2=0 $Y2=0
cc_710 N_A_306_74#_M1032_g N_A_1271_74#_c_1212_n 0.00513624f $X=7.33 $Y=0.615
+ $X2=0 $Y2=0
cc_711 N_A_306_74#_M1032_g N_A_1271_74#_c_1214_n 0.00152295f $X=7.33 $Y=0.615
+ $X2=0 $Y2=0
cc_712 N_A_306_74#_c_909_n N_A_1271_74#_c_1215_n 0.00544498f $X=7.255 $Y=1.66
+ $X2=0 $Y2=0
cc_713 N_A_306_74#_c_928_n N_A_1271_74#_c_1215_n 0.00457177f $X=6.485 $Y=1.66
+ $X2=0 $Y2=0
cc_714 N_A_306_74#_M1032_g N_A_1271_74#_c_1215_n 2.71569e-19 $X=7.33 $Y=0.615
+ $X2=0 $Y2=0
cc_715 N_A_306_74#_c_918_n N_VPWR_c_1430_n 0.00954209f $X=2.375 $Y=1.735 $X2=0
+ $Y2=0
cc_716 N_A_306_74#_c_919_n N_VPWR_c_1430_n 0.00503614f $X=2.88 $Y=3.075 $X2=0
+ $Y2=0
cc_717 N_A_306_74#_c_922_n N_VPWR_c_1431_n 0.00666114f $X=3.855 $Y=2.87 $X2=0
+ $Y2=0
cc_718 N_A_306_74#_c_925_n N_VPWR_c_1431_n 0.0249582f $X=6.32 $Y=3.15 $X2=0
+ $Y2=0
cc_719 N_A_306_74#_c_925_n N_VPWR_c_1432_n 0.0218115f $X=6.32 $Y=3.15 $X2=0
+ $Y2=0
cc_720 N_A_306_74#_c_925_n N_VPWR_c_1433_n 0.025868f $X=6.32 $Y=3.15 $X2=0 $Y2=0
cc_721 N_A_306_74#_M1021_g N_VPWR_c_1433_n 0.00120875f $X=6.41 $Y=2.31 $X2=0
+ $Y2=0
cc_722 N_A_306_74#_c_931_n N_VPWR_c_1433_n 0.00521396f $X=6.41 $Y=3.15 $X2=0
+ $Y2=0
cc_723 N_A_306_74#_c_918_n N_VPWR_c_1443_n 0.0049908f $X=2.375 $Y=1.735 $X2=0
+ $Y2=0
cc_724 N_A_306_74#_c_921_n N_VPWR_c_1443_n 0.04672f $X=2.955 $Y=3.15 $X2=0 $Y2=0
cc_725 N_A_306_74#_c_925_n N_VPWR_c_1444_n 0.020324f $X=6.32 $Y=3.15 $X2=0 $Y2=0
cc_726 N_A_306_74#_c_918_n N_VPWR_c_1426_n 0.00486206f $X=2.375 $Y=1.735 $X2=0
+ $Y2=0
cc_727 N_A_306_74#_c_920_n N_VPWR_c_1426_n 0.0260201f $X=3.765 $Y=3.15 $X2=0
+ $Y2=0
cc_728 N_A_306_74#_c_921_n N_VPWR_c_1426_n 0.00715677f $X=2.955 $Y=3.15 $X2=0
+ $Y2=0
cc_729 N_A_306_74#_c_925_n N_VPWR_c_1426_n 0.0546227f $X=6.32 $Y=3.15 $X2=0
+ $Y2=0
cc_730 N_A_306_74#_c_930_n N_VPWR_c_1426_n 0.0053759f $X=3.855 $Y=3.15 $X2=0
+ $Y2=0
cc_731 N_A_306_74#_c_931_n N_VPWR_c_1426_n 0.0125228f $X=6.41 $Y=3.15 $X2=0
+ $Y2=0
cc_732 N_A_306_74#_c_912_n N_A_30_78#_c_1577_n 0.0042997f $X=1.675 $Y=0.515
+ $X2=0 $Y2=0
cc_733 N_A_306_74#_c_917_n N_A_30_78#_c_1577_n 0.00486098f $X=1.647 $Y=1.065
+ $X2=0 $Y2=0
cc_734 N_A_306_74#_M1007_s N_A_30_78#_c_1585_n 0.00756572f $X=1.57 $Y=1.81 $X2=0
+ $Y2=0
cc_735 N_A_306_74#_c_918_n N_A_30_78#_c_1585_n 0.0126414f $X=2.375 $Y=1.735
+ $X2=0 $Y2=0
cc_736 N_A_306_74#_c_919_n N_A_30_78#_c_1585_n 0.013225f $X=2.88 $Y=3.075 $X2=0
+ $Y2=0
cc_737 N_A_306_74#_c_929_n N_A_30_78#_c_1585_n 0.00120812f $X=2.51 $Y=1.575
+ $X2=0 $Y2=0
cc_738 N_A_306_74#_c_934_n N_A_30_78#_c_1585_n 0.0249302f $X=1.7 $Y=1.985 $X2=0
+ $Y2=0
cc_739 N_A_306_74#_c_907_n N_A_30_78#_c_1578_n 0.00635848f $X=3.435 $Y=1.26
+ $X2=0 $Y2=0
cc_740 N_A_306_74#_c_908_n N_A_30_78#_c_1578_n 0.00853862f $X=3.51 $Y=1.185
+ $X2=0 $Y2=0
cc_741 N_A_306_74#_c_924_n N_A_30_78#_c_1586_n 7.89857e-19 $X=3.855 $Y=2.78
+ $X2=0 $Y2=0
cc_742 N_A_306_74#_c_919_n N_A_30_78#_c_1588_n 0.0120648f $X=2.88 $Y=3.075 $X2=0
+ $Y2=0
cc_743 N_A_306_74#_c_920_n N_A_30_78#_c_1588_n 0.00431186f $X=3.765 $Y=3.15
+ $X2=0 $Y2=0
cc_744 N_A_306_74#_c_907_n N_A_30_78#_c_1581_n 0.0136775f $X=3.435 $Y=1.26 $X2=0
+ $Y2=0
cc_745 N_A_306_74#_c_914_n N_VGND_M1000_d 0.00368125f $X=2.445 $Y=1.065 $X2=0
+ $Y2=0
cc_746 N_A_306_74#_c_912_n N_VGND_c_1714_n 0.0388154f $X=1.675 $Y=0.515 $X2=0
+ $Y2=0
cc_747 N_A_306_74#_c_906_n N_VGND_c_1715_n 0.00564691f $X=2.46 $Y=1.185 $X2=0
+ $Y2=0
cc_748 N_A_306_74#_c_912_n N_VGND_c_1715_n 0.0184628f $X=1.675 $Y=0.515 $X2=0
+ $Y2=0
cc_749 N_A_306_74#_c_914_n N_VGND_c_1715_n 0.0248957f $X=2.445 $Y=1.065 $X2=0
+ $Y2=0
cc_750 N_A_306_74#_M1032_g N_VGND_c_1716_n 4.38128e-19 $X=7.33 $Y=0.615 $X2=0
+ $Y2=0
cc_751 N_A_306_74#_c_912_n N_VGND_c_1723_n 0.0170181f $X=1.675 $Y=0.515 $X2=0
+ $Y2=0
cc_752 N_A_306_74#_c_906_n N_VGND_c_1724_n 0.00433834f $X=2.46 $Y=1.185 $X2=0
+ $Y2=0
cc_753 N_A_306_74#_M1032_g N_VGND_c_1725_n 9.34015e-19 $X=7.33 $Y=0.615 $X2=0
+ $Y2=0
cc_754 N_A_306_74#_c_906_n N_VGND_c_1733_n 0.00826005f $X=2.46 $Y=1.185 $X2=0
+ $Y2=0
cc_755 N_A_306_74#_c_912_n N_VGND_c_1733_n 0.0140297f $X=1.675 $Y=0.515 $X2=0
+ $Y2=0
cc_756 N_A_1525_212#_c_1090_n N_A_1271_74#_M1024_g 0.0108536f $X=8.68 $Y=1.305
+ $X2=0 $Y2=0
cc_757 N_A_1525_212#_c_1091_n N_A_1271_74#_M1024_g 0.0236543f $X=8.845 $Y=0.615
+ $X2=0 $Y2=0
cc_758 N_A_1525_212#_c_1093_n N_A_1271_74#_M1024_g 0.00397247f $X=9.29 $Y=2.105
+ $X2=0 $Y2=0
cc_759 N_A_1525_212#_c_1096_n N_A_1271_74#_M1024_g 0.00478437f $X=8.845 $Y=1.305
+ $X2=0 $Y2=0
cc_760 N_A_1525_212#_c_1102_n N_A_1271_74#_c_1216_n 7.30818e-19 $X=8.8 $Y=2.445
+ $X2=0 $Y2=0
cc_761 N_A_1525_212#_c_1103_n N_A_1271_74#_c_1216_n 0.0134689f $X=9.205 $Y=2.19
+ $X2=0 $Y2=0
cc_762 N_A_1525_212#_c_1104_n N_A_1271_74#_c_1216_n 0.00277746f $X=8.885 $Y=2.19
+ $X2=0 $Y2=0
cc_763 N_A_1525_212#_c_1101_n N_A_1271_74#_c_1217_n 0.00989487f $X=8.715 $Y=2.61
+ $X2=0 $Y2=0
cc_764 N_A_1525_212#_c_1102_n N_A_1271_74#_c_1217_n 0.00482538f $X=8.8 $Y=2.445
+ $X2=0 $Y2=0
cc_765 N_A_1525_212#_c_1103_n N_A_1271_74#_c_1207_n 0.00213341f $X=9.205 $Y=2.19
+ $X2=0 $Y2=0
cc_766 N_A_1525_212#_c_1093_n N_A_1271_74#_c_1207_n 0.0139731f $X=9.29 $Y=2.105
+ $X2=0 $Y2=0
cc_767 N_A_1525_212#_c_1104_n N_A_1271_74#_c_1208_n 0.0010617f $X=8.885 $Y=2.19
+ $X2=0 $Y2=0
cc_768 N_A_1525_212#_c_1092_n N_A_1271_74#_c_1208_n 0.00714341f $X=9.205
+ $Y=1.305 $X2=0 $Y2=0
cc_769 N_A_1525_212#_c_1093_n N_A_1271_74#_c_1208_n 0.00618579f $X=9.29 $Y=2.105
+ $X2=0 $Y2=0
cc_770 N_A_1525_212#_c_1096_n N_A_1271_74#_c_1208_n 0.00565398f $X=8.845
+ $Y=1.305 $X2=0 $Y2=0
cc_771 N_A_1525_212#_c_1093_n N_A_1271_74#_c_1220_n 0.00269774f $X=9.29 $Y=2.105
+ $X2=0 $Y2=0
cc_772 N_A_1525_212#_c_1102_n N_A_1271_74#_c_1221_n 7.46191e-19 $X=8.8 $Y=2.445
+ $X2=0 $Y2=0
cc_773 N_A_1525_212#_c_1103_n N_A_1271_74#_c_1221_n 0.00172099f $X=9.205 $Y=2.19
+ $X2=0 $Y2=0
cc_774 N_A_1525_212#_c_1093_n N_A_1271_74#_c_1221_n 0.00125184f $X=9.29 $Y=2.105
+ $X2=0 $Y2=0
cc_775 N_A_1525_212#_c_1091_n N_A_1271_74#_M1022_g 0.00350395f $X=8.845 $Y=0.615
+ $X2=0 $Y2=0
cc_776 N_A_1525_212#_c_1092_n N_A_1271_74#_M1022_g 0.00377053f $X=9.205 $Y=1.305
+ $X2=0 $Y2=0
cc_777 N_A_1525_212#_c_1093_n N_A_1271_74#_M1022_g 0.00338537f $X=9.29 $Y=2.105
+ $X2=0 $Y2=0
cc_778 N_A_1525_212#_c_1099_n N_A_1271_74#_c_1224_n 0.00151725f $X=7.735 $Y=2.39
+ $X2=0 $Y2=0
cc_779 N_A_1525_212#_c_1089_n N_A_1271_74#_c_1224_n 0.0136876f $X=7.735 $Y=1.975
+ $X2=0 $Y2=0
cc_780 N_A_1525_212#_c_1097_n N_A_1271_74#_c_1213_n 2.78684e-19 $X=7.735
+ $Y=2.065 $X2=0 $Y2=0
cc_781 N_A_1525_212#_c_1089_n N_A_1271_74#_c_1213_n 0.0105727f $X=7.735 $Y=1.975
+ $X2=0 $Y2=0
cc_782 N_A_1525_212#_c_1090_n N_A_1271_74#_c_1213_n 0.0522284f $X=8.68 $Y=1.305
+ $X2=0 $Y2=0
cc_783 N_A_1525_212#_c_1094_n N_A_1271_74#_c_1213_n 0.023491f $X=7.79 $Y=1.225
+ $X2=0 $Y2=0
cc_784 N_A_1525_212#_c_1095_n N_A_1271_74#_c_1213_n 0.00116263f $X=7.79 $Y=1.225
+ $X2=0 $Y2=0
cc_785 N_A_1525_212#_c_1096_n N_A_1271_74#_c_1213_n 0.00190438f $X=8.845
+ $Y=1.305 $X2=0 $Y2=0
cc_786 N_A_1525_212#_c_1101_n N_A_1271_74#_c_1228_n 2.74753e-19 $X=8.715 $Y=2.61
+ $X2=0 $Y2=0
cc_787 N_A_1525_212#_c_1103_n N_A_1271_74#_c_1228_n 0.00882758f $X=9.205 $Y=2.19
+ $X2=0 $Y2=0
cc_788 N_A_1525_212#_c_1104_n N_A_1271_74#_c_1228_n 0.0119175f $X=8.885 $Y=2.19
+ $X2=0 $Y2=0
cc_789 N_A_1525_212#_c_1092_n N_A_1271_74#_c_1228_n 0.00177485f $X=9.205
+ $Y=1.305 $X2=0 $Y2=0
cc_790 N_A_1525_212#_c_1093_n N_A_1271_74#_c_1228_n 0.0242588f $X=9.29 $Y=2.105
+ $X2=0 $Y2=0
cc_791 N_A_1525_212#_c_1096_n N_A_1271_74#_c_1228_n 0.0257641f $X=8.845 $Y=1.305
+ $X2=0 $Y2=0
cc_792 N_A_1525_212#_c_1103_n N_A_1921_409#_c_1370_n 0.011653f $X=9.205 $Y=2.19
+ $X2=0 $Y2=0
cc_793 N_A_1525_212#_c_1093_n N_A_1921_409#_c_1370_n 0.00461168f $X=9.29
+ $Y=2.105 $X2=0 $Y2=0
cc_794 N_A_1525_212#_c_1091_n N_A_1921_409#_c_1362_n 0.00484112f $X=8.845
+ $Y=0.615 $X2=0 $Y2=0
cc_795 N_A_1525_212#_c_1092_n N_A_1921_409#_c_1362_n 0.00459026f $X=9.205
+ $Y=1.305 $X2=0 $Y2=0
cc_796 N_A_1525_212#_c_1093_n N_A_1921_409#_c_1363_n 0.0210733f $X=9.29 $Y=2.105
+ $X2=0 $Y2=0
cc_797 N_A_1525_212#_c_1092_n N_A_1921_409#_c_1364_n 0.00528833f $X=9.205
+ $Y=1.305 $X2=0 $Y2=0
cc_798 N_A_1525_212#_c_1093_n N_A_1921_409#_c_1364_n 0.0123556f $X=9.29 $Y=2.105
+ $X2=0 $Y2=0
cc_799 N_A_1525_212#_c_1103_n N_VPWR_M1014_d 0.00763182f $X=9.205 $Y=2.19 $X2=0
+ $Y2=0
cc_800 N_A_1525_212#_c_1093_n N_VPWR_M1014_d 0.00173132f $X=9.29 $Y=2.105 $X2=0
+ $Y2=0
cc_801 N_A_1525_212#_c_1099_n N_VPWR_c_1434_n 0.0101713f $X=7.735 $Y=2.39 $X2=0
+ $Y2=0
cc_802 N_A_1525_212#_c_1101_n N_VPWR_c_1434_n 0.0142734f $X=8.715 $Y=2.61 $X2=0
+ $Y2=0
cc_803 N_A_1525_212#_c_1101_n N_VPWR_c_1435_n 0.0232957f $X=8.715 $Y=2.61 $X2=0
+ $Y2=0
cc_804 N_A_1525_212#_c_1103_n N_VPWR_c_1435_n 0.0245347f $X=9.205 $Y=2.19 $X2=0
+ $Y2=0
cc_805 N_A_1525_212#_c_1101_n N_VPWR_c_1439_n 0.01191f $X=8.715 $Y=2.61 $X2=0
+ $Y2=0
cc_806 N_A_1525_212#_c_1099_n N_VPWR_c_1444_n 0.00470366f $X=7.735 $Y=2.39 $X2=0
+ $Y2=0
cc_807 N_A_1525_212#_c_1099_n N_VPWR_c_1426_n 0.00473388f $X=7.735 $Y=2.39 $X2=0
+ $Y2=0
cc_808 N_A_1525_212#_c_1101_n N_VPWR_c_1426_n 0.0185129f $X=8.715 $Y=2.61 $X2=0
+ $Y2=0
cc_809 N_A_1525_212#_M1010_g N_VGND_c_1716_n 0.00870177f $X=7.72 $Y=0.615 $X2=0
+ $Y2=0
cc_810 N_A_1525_212#_c_1090_n N_VGND_c_1716_n 0.00751614f $X=8.68 $Y=1.305 $X2=0
+ $Y2=0
cc_811 N_A_1525_212#_c_1091_n N_VGND_c_1716_n 0.0106511f $X=8.845 $Y=0.615 $X2=0
+ $Y2=0
cc_812 N_A_1525_212#_c_1094_n N_VGND_c_1716_n 0.00718492f $X=7.79 $Y=1.225 $X2=0
+ $Y2=0
cc_813 N_A_1525_212#_c_1095_n N_VGND_c_1716_n 9.12984e-19 $X=7.79 $Y=1.225 $X2=0
+ $Y2=0
cc_814 N_A_1525_212#_c_1091_n N_VGND_c_1717_n 0.045283f $X=8.845 $Y=0.615 $X2=0
+ $Y2=0
cc_815 N_A_1525_212#_c_1092_n N_VGND_c_1717_n 0.0132803f $X=9.205 $Y=1.305 $X2=0
+ $Y2=0
cc_816 N_A_1525_212#_M1010_g N_VGND_c_1725_n 0.0045897f $X=7.72 $Y=0.615 $X2=0
+ $Y2=0
cc_817 N_A_1525_212#_c_1091_n N_VGND_c_1726_n 0.0127604f $X=8.845 $Y=0.615 $X2=0
+ $Y2=0
cc_818 N_A_1525_212#_M1010_g N_VGND_c_1733_n 0.0044912f $X=7.72 $Y=0.615 $X2=0
+ $Y2=0
cc_819 N_A_1525_212#_c_1091_n N_VGND_c_1733_n 0.011834f $X=8.845 $Y=0.615 $X2=0
+ $Y2=0
cc_820 N_A_1271_74#_c_1216_n N_A_1921_409#_c_1370_n 5.28212e-19 $X=8.945 $Y=2.3
+ $X2=0 $Y2=0
cc_821 N_A_1271_74#_c_1217_n N_A_1921_409#_c_1370_n 3.28834e-19 $X=8.945 $Y=2.39
+ $X2=0 $Y2=0
cc_822 N_A_1271_74#_c_1221_n N_A_1921_409#_c_1370_n 0.0159253f $X=9.53 $Y=1.97
+ $X2=0 $Y2=0
cc_823 N_A_1271_74#_c_1210_n N_A_1921_409#_c_1370_n 0.0016406f $X=9.562 $Y=1.63
+ $X2=0 $Y2=0
cc_824 N_A_1271_74#_M1022_g N_A_1921_409#_c_1362_n 0.0181066f $X=9.61 $Y=0.74
+ $X2=0 $Y2=0
cc_825 N_A_1271_74#_c_1220_n N_A_1921_409#_c_1363_n 0.00666991f $X=9.53 $Y=1.88
+ $X2=0 $Y2=0
cc_826 N_A_1271_74#_c_1221_n N_A_1921_409#_c_1363_n 0.00141733f $X=9.53 $Y=1.97
+ $X2=0 $Y2=0
cc_827 N_A_1271_74#_c_1210_n N_A_1921_409#_c_1363_n 0.00365747f $X=9.562 $Y=1.63
+ $X2=0 $Y2=0
cc_828 N_A_1271_74#_M1022_g N_A_1921_409#_c_1364_n 0.00613547f $X=9.61 $Y=0.74
+ $X2=0 $Y2=0
cc_829 N_A_1271_74#_c_1210_n N_A_1921_409#_c_1364_n 0.00242696f $X=9.562 $Y=1.63
+ $X2=0 $Y2=0
cc_830 N_A_1271_74#_M1022_g N_A_1921_409#_c_1365_n 0.0181431f $X=9.61 $Y=0.74
+ $X2=0 $Y2=0
cc_831 N_A_1271_74#_c_1224_n N_VPWR_c_1434_n 0.00184051f $X=7.54 $Y=2.475 $X2=0
+ $Y2=0
cc_832 N_A_1271_74#_c_1217_n N_VPWR_c_1435_n 0.0100164f $X=8.945 $Y=2.39 $X2=0
+ $Y2=0
cc_833 N_A_1271_74#_c_1221_n N_VPWR_c_1435_n 0.00627469f $X=9.53 $Y=1.97 $X2=0
+ $Y2=0
cc_834 N_A_1271_74#_c_1221_n N_VPWR_c_1436_n 0.00466121f $X=9.53 $Y=1.97 $X2=0
+ $Y2=0
cc_835 N_A_1271_74#_c_1217_n N_VPWR_c_1439_n 0.00511015f $X=8.945 $Y=2.39 $X2=0
+ $Y2=0
cc_836 N_A_1271_74#_c_1237_n N_VPWR_c_1444_n 0.0207747f $X=7.455 $Y=2.64 $X2=0
+ $Y2=0
cc_837 N_A_1271_74#_c_1338_p N_VPWR_c_1444_n 0.00391127f $X=6.685 $Y=2.64 $X2=0
+ $Y2=0
cc_838 N_A_1271_74#_c_1221_n N_VPWR_c_1445_n 0.00510653f $X=9.53 $Y=1.97 $X2=0
+ $Y2=0
cc_839 N_A_1271_74#_c_1217_n N_VPWR_c_1426_n 0.0052212f $X=8.945 $Y=2.39 $X2=0
+ $Y2=0
cc_840 N_A_1271_74#_c_1221_n N_VPWR_c_1426_n 0.0052212f $X=9.53 $Y=1.97 $X2=0
+ $Y2=0
cc_841 N_A_1271_74#_c_1237_n N_VPWR_c_1426_n 0.029938f $X=7.455 $Y=2.64 $X2=0
+ $Y2=0
cc_842 N_A_1271_74#_c_1338_p N_VPWR_c_1426_n 0.00557315f $X=6.685 $Y=2.64 $X2=0
+ $Y2=0
cc_843 N_A_1271_74#_c_1237_n A_1478_493# 0.00315877f $X=7.455 $Y=2.64 $X2=-0.19
+ $Y2=-0.245
cc_844 N_A_1271_74#_M1024_g N_VGND_c_1716_n 0.00147575f $X=8.63 $Y=0.615 $X2=0
+ $Y2=0
cc_845 N_A_1271_74#_M1024_g N_VGND_c_1717_n 0.00438924f $X=8.63 $Y=0.615 $X2=0
+ $Y2=0
cc_846 N_A_1271_74#_c_1207_n N_VGND_c_1717_n 0.00293701f $X=9.44 $Y=1.63 $X2=0
+ $Y2=0
cc_847 N_A_1271_74#_M1022_g N_VGND_c_1717_n 0.00488092f $X=9.61 $Y=0.74 $X2=0
+ $Y2=0
cc_848 N_A_1271_74#_M1022_g N_VGND_c_1718_n 0.00412165f $X=9.61 $Y=0.74 $X2=0
+ $Y2=0
cc_849 N_A_1271_74#_M1024_g N_VGND_c_1726_n 0.00527282f $X=8.63 $Y=0.615 $X2=0
+ $Y2=0
cc_850 N_A_1271_74#_M1022_g N_VGND_c_1727_n 0.00434272f $X=9.61 $Y=0.74 $X2=0
+ $Y2=0
cc_851 N_A_1271_74#_M1024_g N_VGND_c_1733_n 0.00534666f $X=8.63 $Y=0.615 $X2=0
+ $Y2=0
cc_852 N_A_1271_74#_M1022_g N_VGND_c_1733_n 0.00830282f $X=9.61 $Y=0.74 $X2=0
+ $Y2=0
cc_853 N_A_1921_409#_c_1370_n N_VPWR_c_1435_n 0.0180508f $X=9.755 $Y=2.195 $X2=0
+ $Y2=0
cc_854 N_A_1921_409#_c_1354_n N_VPWR_c_1436_n 0.00728605f $X=10.475 $Y=1.375
+ $X2=0 $Y2=0
cc_855 N_A_1921_409#_c_1367_n N_VPWR_c_1436_n 0.0053787f $X=10.565 $Y=1.765
+ $X2=0 $Y2=0
cc_856 N_A_1921_409#_c_1363_n N_VPWR_c_1436_n 0.0728323f $X=9.755 $Y=2.03 $X2=0
+ $Y2=0
cc_857 N_A_1921_409#_c_1364_n N_VPWR_c_1436_n 0.00302521f $X=10.09 $Y=1.465
+ $X2=0 $Y2=0
cc_858 N_A_1921_409#_c_1365_n N_VPWR_c_1436_n 0.00372647f $X=10.09 $Y=1.375
+ $X2=0 $Y2=0
cc_859 N_A_1921_409#_c_1369_n N_VPWR_c_1438_n 0.00835395f $X=11.015 $Y=1.765
+ $X2=0 $Y2=0
cc_860 N_A_1921_409#_c_1370_n N_VPWR_c_1445_n 0.0111926f $X=9.755 $Y=2.195 $X2=0
+ $Y2=0
cc_861 N_A_1921_409#_c_1367_n N_VPWR_c_1446_n 0.00461464f $X=10.565 $Y=1.765
+ $X2=0 $Y2=0
cc_862 N_A_1921_409#_c_1369_n N_VPWR_c_1446_n 0.00417277f $X=11.015 $Y=1.765
+ $X2=0 $Y2=0
cc_863 N_A_1921_409#_c_1367_n N_VPWR_c_1426_n 0.00912521f $X=10.565 $Y=1.765
+ $X2=0 $Y2=0
cc_864 N_A_1921_409#_c_1369_n N_VPWR_c_1426_n 0.00769367f $X=11.015 $Y=1.765
+ $X2=0 $Y2=0
cc_865 N_A_1921_409#_c_1370_n N_VPWR_c_1426_n 0.0115381f $X=9.755 $Y=2.195 $X2=0
+ $Y2=0
cc_866 N_A_1921_409#_c_1355_n Q 0.00718159f $X=10.565 $Y=1.675 $X2=0 $Y2=0
cc_867 N_A_1921_409#_c_1367_n Q 0.00700399f $X=10.565 $Y=1.765 $X2=0 $Y2=0
cc_868 N_A_1921_409#_M1031_g Q 0.0157053f $X=10.6 $Y=0.74 $X2=0 $Y2=0
cc_869 N_A_1921_409#_c_1357_n Q 0.00813241f $X=10.925 $Y=1.375 $X2=0 $Y2=0
cc_870 N_A_1921_409#_c_1358_n Q 0.0128965f $X=11.015 $Y=1.675 $X2=0 $Y2=0
cc_871 N_A_1921_409#_c_1369_n Q 0.0235958f $X=11.015 $Y=1.765 $X2=0 $Y2=0
cc_872 N_A_1921_409#_M1033_g Q 0.0192861f $X=11.03 $Y=0.74 $X2=0 $Y2=0
cc_873 N_A_1921_409#_c_1360_n Q 0.00396751f $X=10.575 $Y=1.375 $X2=0 $Y2=0
cc_874 N_A_1921_409#_c_1361_n Q 0.00693891f $X=11.015 $Y=1.375 $X2=0 $Y2=0
cc_875 N_A_1921_409#_c_1362_n Q 0.00478422f $X=9.825 $Y=0.515 $X2=0 $Y2=0
cc_876 N_A_1921_409#_c_1364_n Q 0.0113958f $X=10.09 $Y=1.465 $X2=0 $Y2=0
cc_877 N_A_1921_409#_c_1365_n Q 5.0889e-19 $X=10.09 $Y=1.375 $X2=0 $Y2=0
cc_878 N_A_1921_409#_c_1362_n N_VGND_c_1717_n 0.0258169f $X=9.825 $Y=0.515 $X2=0
+ $Y2=0
cc_879 N_A_1921_409#_M1031_g N_VGND_c_1718_n 0.00647412f $X=10.6 $Y=0.74 $X2=0
+ $Y2=0
cc_880 N_A_1921_409#_c_1362_n N_VGND_c_1718_n 0.051504f $X=9.825 $Y=0.515 $X2=0
+ $Y2=0
cc_881 N_A_1921_409#_c_1365_n N_VGND_c_1718_n 0.0102912f $X=10.09 $Y=1.375 $X2=0
+ $Y2=0
cc_882 N_A_1921_409#_M1033_g N_VGND_c_1720_n 0.00647412f $X=11.03 $Y=0.74 $X2=0
+ $Y2=0
cc_883 N_A_1921_409#_c_1362_n N_VGND_c_1727_n 0.0145639f $X=9.825 $Y=0.515 $X2=0
+ $Y2=0
cc_884 N_A_1921_409#_M1031_g N_VGND_c_1728_n 0.00434272f $X=10.6 $Y=0.74 $X2=0
+ $Y2=0
cc_885 N_A_1921_409#_M1033_g N_VGND_c_1728_n 0.00434272f $X=11.03 $Y=0.74 $X2=0
+ $Y2=0
cc_886 N_A_1921_409#_M1031_g N_VGND_c_1733_n 0.00825283f $X=10.6 $Y=0.74 $X2=0
+ $Y2=0
cc_887 N_A_1921_409#_M1033_g N_VGND_c_1733_n 0.00823925f $X=11.03 $Y=0.74 $X2=0
+ $Y2=0
cc_888 N_A_1921_409#_c_1362_n N_VGND_c_1733_n 0.0119984f $X=9.825 $Y=0.515 $X2=0
+ $Y2=0
cc_889 N_VPWR_c_1428_n N_A_30_78#_c_1582_n 0.00665174f $X=0.27 $Y=2.75 $X2=0
+ $Y2=0
cc_890 N_VPWR_c_1428_n N_A_30_78#_c_1583_n 0.0237304f $X=0.27 $Y=2.75 $X2=0
+ $Y2=0
cc_891 N_VPWR_c_1429_n N_A_30_78#_c_1583_n 0.0127399f $X=1.17 $Y=2.78 $X2=0
+ $Y2=0
cc_892 N_VPWR_c_1441_n N_A_30_78#_c_1583_n 0.00879902f $X=1.005 $Y=3.33 $X2=0
+ $Y2=0
cc_893 N_VPWR_c_1426_n N_A_30_78#_c_1583_n 0.007299f $X=11.28 $Y=3.33 $X2=0
+ $Y2=0
cc_894 N_VPWR_M1007_d N_A_30_78#_c_1585_n 0.00491303f $X=2 $Y=1.81 $X2=0 $Y2=0
cc_895 N_VPWR_c_1429_n N_A_30_78#_c_1585_n 0.0231054f $X=1.17 $Y=2.78 $X2=0
+ $Y2=0
cc_896 N_VPWR_c_1430_n N_A_30_78#_c_1585_n 0.0162642f $X=2.15 $Y=2.765 $X2=0
+ $Y2=0
cc_897 N_VPWR_c_1426_n N_A_30_78#_c_1585_n 0.0483846f $X=11.28 $Y=3.33 $X2=0
+ $Y2=0
cc_898 N_VPWR_c_1443_n N_A_30_78#_c_1588_n 0.00531752f $X=4.42 $Y=3.33 $X2=0
+ $Y2=0
cc_899 N_VPWR_c_1426_n N_A_30_78#_c_1588_n 0.00670829f $X=11.28 $Y=3.33 $X2=0
+ $Y2=0
cc_900 N_VPWR_c_1436_n Q 0.00316191f $X=10.315 $Y=1.985 $X2=0 $Y2=0
cc_901 N_VPWR_c_1438_n Q 0.0862588f $X=11.24 $Y=1.985 $X2=0 $Y2=0
cc_902 N_VPWR_c_1446_n Q 0.0145191f $X=11.155 $Y=3.33 $X2=0 $Y2=0
cc_903 N_VPWR_c_1426_n Q 0.011926f $X=11.28 $Y=3.33 $X2=0 $Y2=0
cc_904 N_A_30_78#_c_1576_n A_117_78# 0.00232882f $X=0.665 $Y=0.745 $X2=-0.19
+ $Y2=-0.245
cc_905 N_A_30_78#_c_1576_n N_VGND_c_1714_n 0.00655394f $X=0.665 $Y=0.745 $X2=0
+ $Y2=0
cc_906 N_A_30_78#_c_1580_n N_VGND_c_1714_n 0.00436551f $X=0.295 $Y=0.6 $X2=0
+ $Y2=0
cc_907 N_A_30_78#_c_1576_n N_VGND_c_1721_n 0.00539861f $X=0.665 $Y=0.745 $X2=0
+ $Y2=0
cc_908 N_A_30_78#_c_1580_n N_VGND_c_1721_n 0.0131067f $X=0.295 $Y=0.6 $X2=0
+ $Y2=0
cc_909 N_A_30_78#_c_1576_n N_VGND_c_1733_n 0.0106557f $X=0.665 $Y=0.745 $X2=0
+ $Y2=0
cc_910 N_A_30_78#_c_1580_n N_VGND_c_1733_n 0.0117869f $X=0.295 $Y=0.6 $X2=0
+ $Y2=0
cc_911 Q N_VGND_c_1718_n 0.0294122f $X=10.715 $Y=0.47 $X2=0 $Y2=0
cc_912 Q N_VGND_c_1720_n 0.0294122f $X=10.715 $Y=0.47 $X2=0 $Y2=0
cc_913 Q N_VGND_c_1728_n 0.0144922f $X=10.715 $Y=0.47 $X2=0 $Y2=0
cc_914 Q N_VGND_c_1733_n 0.0118826f $X=10.715 $Y=0.47 $X2=0 $Y2=0
