* File: sky130_fd_sc_hs__sdfstp_2.pex.spice
* Created: Tue Sep  1 20:23:17 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HS__SDFSTP_2%SCE 2 5 7 9 10 12 15 20 21 23 24 28 32
r76 32 34 45.456 $w=3.9e-07 $l=1.65e-07 $layer=POLY_cond $X=0.61 $Y=1.635
+ $X2=0.61 $Y2=1.47
r77 28 32 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.64
+ $Y=1.635 $X2=0.64 $Y2=1.635
r78 24 36 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.96 $Y=1.415
+ $X2=1.96 $Y2=1.25
r79 23 26 3.68782 $w=2.48e-07 $l=8e-08 $layer=LI1_cond $X=1.92 $Y=1.415 $X2=1.92
+ $Y2=1.495
r80 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.96
+ $Y=1.415 $X2=1.96 $Y2=1.415
r81 21 28 9.23067 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.805 $Y=1.495
+ $X2=0.72 $Y2=1.58
r82 20 26 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.795 $Y=1.495
+ $X2=1.92 $Y2=1.495
r83 20 21 64.5882 $w=1.68e-07 $l=9.9e-07 $layer=LI1_cond $X=1.795 $Y=1.495
+ $X2=0.805 $Y2=1.495
r84 15 36 343.553 $w=1.5e-07 $l=6.7e-07 $layer=POLY_cond $X=1.94 $Y=0.58
+ $X2=1.94 $Y2=1.25
r85 10 19 10.701 $w=1.5e-07 $l=1.28e-07 $layer=POLY_cond $X=0.955 $Y=2.245
+ $X2=0.955 $Y2=2.117
r86 10 12 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=0.955 $Y=2.245
+ $X2=0.955 $Y2=2.64
r87 7 17 10.701 $w=1.5e-07 $l=1.28e-07 $layer=POLY_cond $X=0.505 $Y=2.245
+ $X2=0.505 $Y2=2.117
r88 7 9 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=0.505 $Y=2.245
+ $X2=0.505 $Y2=2.64
r89 5 34 456.362 $w=1.5e-07 $l=8.9e-07 $layer=POLY_cond $X=0.495 $Y=0.58
+ $X2=0.495 $Y2=1.47
r90 2 19 79.1857 $w=2.1e-07 $l=3.45e-07 $layer=POLY_cond $X=0.61 $Y=2.117
+ $X2=0.955 $Y2=2.117
r91 2 17 24.1 $w=2.1e-07 $l=1.05e-07 $layer=POLY_cond $X=0.61 $Y=2.117 $X2=0.505
+ $Y2=2.117
r92 1 32 4.27811 $w=3.9e-07 $l=3e-08 $layer=POLY_cond $X=0.61 $Y=1.665 $X2=0.61
+ $Y2=1.635
r93 1 2 46.3462 $w=3.9e-07 $l=3.25e-07 $layer=POLY_cond $X=0.61 $Y=1.665
+ $X2=0.61 $Y2=1.99
.ends

.subckt PM_SKY130_FD_SC_HS__SDFSTP_2%A_27_74# 1 2 9 10 12 15 18 21 25 26 30 33
+ 35 37
c73 30 0 7.10762e-20 $X=1.96 $Y=1.995
c74 26 0 1.86174e-19 $X=1.06 $Y=1.065
c75 21 0 1.64533e-19 $X=1.795 $Y=2.405
r76 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.96
+ $Y=1.995 $X2=1.96 $Y2=1.995
r77 28 30 14.9818 $w=2.48e-07 $l=3.25e-07 $layer=LI1_cond $X=1.92 $Y=2.32
+ $X2=1.92 $Y2=1.995
r78 26 37 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.06 $Y=1.065
+ $X2=1.06 $Y2=0.9
r79 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.06
+ $Y=1.065 $X2=1.06 $Y2=1.065
r80 23 33 0.364692 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=0.445 $Y=1.065
+ $X2=0.28 $Y2=1.065
r81 23 25 21.4773 $w=3.28e-07 $l=6.15e-07 $layer=LI1_cond $X=0.445 $Y=1.065
+ $X2=1.06 $Y2=1.065
r82 22 35 2.11342 $w=1.7e-07 $l=1.27475e-07 $layer=LI1_cond $X=0.365 $Y=2.405
+ $X2=0.24 $Y2=2.4
r83 21 28 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.795 $Y=2.405
+ $X2=1.92 $Y2=2.32
r84 21 22 93.2941 $w=1.68e-07 $l=1.43e-06 $layer=LI1_cond $X=1.795 $Y=2.405
+ $X2=0.365 $Y2=2.405
r85 18 35 4.3182 $w=2.1e-07 $l=1.08167e-07 $layer=LI1_cond $X=0.2 $Y=2.31
+ $X2=0.24 $Y2=2.4
r86 17 33 6.46576 $w=2.5e-07 $l=2.0106e-07 $layer=LI1_cond $X=0.2 $Y=1.23
+ $X2=0.28 $Y2=1.065
r87 17 18 70.4599 $w=1.68e-07 $l=1.08e-06 $layer=LI1_cond $X=0.2 $Y=1.23 $X2=0.2
+ $Y2=2.31
r88 13 33 6.46576 $w=2.5e-07 $l=1.65e-07 $layer=LI1_cond $X=0.28 $Y=0.9 $X2=0.28
+ $Y2=1.065
r89 13 15 11.1752 $w=3.28e-07 $l=3.2e-07 $layer=LI1_cond $X=0.28 $Y=0.9 $X2=0.28
+ $Y2=0.58
r90 10 31 52.2586 $w=2.99e-07 $l=2.7157e-07 $layer=POLY_cond $X=2.005 $Y=2.245
+ $X2=1.96 $Y2=1.995
r91 10 12 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=2.005 $Y=2.245
+ $X2=2.005 $Y2=2.64
r92 9 37 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.12 $Y=0.58 $X2=1.12
+ $Y2=0.9
r93 2 35 300 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=2.32 $X2=0.28 $Y2=2.475
r94 1 15 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_HS__SDFSTP_2%D 1 3 6 8 12
c37 1 0 4.46515e-20 $X=1.375 $Y=2.245
r38 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.42
+ $Y=1.985 $X2=1.42 $Y2=1.985
r39 8 12 7.68295 $w=3.28e-07 $l=2.2e-07 $layer=LI1_cond $X=1.2 $Y=1.985 $X2=1.42
+ $Y2=1.985
r40 4 11 38.5718 $w=2.96e-07 $l=2.05122e-07 $layer=POLY_cond $X=1.51 $Y=1.82
+ $X2=1.42 $Y2=1.985
r41 4 6 635.83 $w=1.5e-07 $l=1.24e-06 $layer=POLY_cond $X=1.51 $Y=1.82 $X2=1.51
+ $Y2=0.58
r42 1 11 54.0414 $w=2.96e-07 $l=2.81603e-07 $layer=POLY_cond $X=1.375 $Y=2.245
+ $X2=1.42 $Y2=1.985
r43 1 3 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=1.375 $Y=2.245
+ $X2=1.375 $Y2=2.64
.ends

.subckt PM_SKY130_FD_SC_HS__SDFSTP_2%SCD 3 6 7 9 10 11 12 17
c41 10 0 6.51157e-20 $X=2.64 $Y=1.295
c42 7 0 2.35609e-19 $X=2.425 $Y=2.245
r43 17 19 46.3954 $w=4.95e-07 $l=1.65e-07 $layer=POLY_cond $X=2.582 $Y=1.305
+ $X2=2.582 $Y2=1.14
r44 12 21 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=2.665
+ $Y=1.985 $X2=2.665 $Y2=1.985
r45 11 12 16.3903 $w=2.23e-07 $l=3.2e-07 $layer=LI1_cond $X=2.667 $Y=1.665
+ $X2=2.667 $Y2=1.985
r46 10 11 18.9513 $w=2.23e-07 $l=3.7e-07 $layer=LI1_cond $X=2.667 $Y=1.295
+ $X2=2.667 $Y2=1.665
r47 10 17 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=2.665
+ $Y=1.305 $X2=2.665 $Y2=1.305
r48 7 21 50.9758 $w=4.07e-07 $l=3.29272e-07 $layer=POLY_cond $X=2.425 $Y=2.245
+ $X2=2.582 $Y2=1.985
r49 7 9 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=2.425 $Y=2.245
+ $X2=2.425 $Y2=2.64
r50 6 21 9.65061 $w=4.95e-07 $l=8.2e-08 $layer=POLY_cond $X=2.582 $Y=1.903
+ $X2=2.582 $Y2=1.985
r51 5 17 8.86311 $w=4.95e-07 $l=8.2e-08 $layer=POLY_cond $X=2.582 $Y=1.387
+ $X2=2.582 $Y2=1.305
r52 5 6 55.7728 $w=4.95e-07 $l=5.16e-07 $layer=POLY_cond $X=2.582 $Y=1.387
+ $X2=2.582 $Y2=1.903
r53 3 19 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=2.41 $Y=0.58 $X2=2.41
+ $Y2=1.14
.ends

.subckt PM_SKY130_FD_SC_HS__SDFSTP_2%CLK 1 3 4 6 7
c35 4 0 6.51157e-20 $X=3.485 $Y=1.765
r36 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.42
+ $Y=1.385 $X2=3.42 $Y2=1.385
r37 7 11 5.60648 $w=3.68e-07 $l=1.8e-07 $layer=LI1_cond $X=3.6 $Y=1.365 $X2=3.42
+ $Y2=1.365
r38 4 10 77.2841 $w=2.7e-07 $l=4.11218e-07 $layer=POLY_cond $X=3.485 $Y=1.765
+ $X2=3.42 $Y2=1.385
r39 4 6 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.485 $Y=1.765
+ $X2=3.485 $Y2=2.4
r40 1 10 38.9026 $w=2.7e-07 $l=1.74714e-07 $layer=POLY_cond $X=3.4 $Y=1.22
+ $X2=3.42 $Y2=1.385
r41 1 3 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=3.4 $Y=1.22 $X2=3.4
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HS__SDFSTP_2%A_795_74# 1 2 8 9 11 12 14 18 22 23 24 26
+ 27 29 31 33 34 36 38 41 45 47 48 49 50 53 57 58 59 60 63 64 65 67 69 70 74 77
+ 78 82 88 89 97 98 99 103
c296 77 0 3.7885e-19 $X=10.555 $Y=1.97
c297 70 0 1.11484e-19 $X=10 $Y=1.64
c298 67 0 1.15295e-19 $X=7.28 $Y=2.905
c299 29 0 3.01101e-20 $X=10.13 $Y=1.085
c300 12 0 1.3233e-19 $X=5.4 $Y=1.655
c301 9 0 4.69178e-20 $X=4.975 $Y=2.21
r302 98 99 24.9528 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=5.565 $Y=1.655
+ $X2=5.565 $Y2=1.58
r303 96 97 33.0969 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=4.975 $Y=1.565
+ $X2=5.065 $Y2=1.565
r304 88 89 8.63679 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=8.255 $Y=1.685
+ $X2=8.425 $Y2=1.685
r305 86 98 39.3438 $w=3.3e-07 $l=2.25e-07 $layer=POLY_cond $X=5.565 $Y=1.88
+ $X2=5.565 $Y2=1.655
r306 85 87 16.0091 $w=2.21e-07 $l=2.9e-07 $layer=LI1_cond $X=5.602 $Y=1.88
+ $X2=5.602 $Y2=2.17
r307 85 86 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.565
+ $Y=1.88 $X2=5.565 $Y2=1.88
r308 78 107 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=10.555 $Y=1.97
+ $X2=10.555 $Y2=2.135
r309 77 78 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.555
+ $Y=1.97 $X2=10.555 $Y2=1.97
r310 75 77 13.4452 $w=3.28e-07 $l=3.85e-07 $layer=LI1_cond $X=10.17 $Y=1.97
+ $X2=10.555 $Y2=1.97
r311 74 103 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=8.975 $Y=1.64
+ $X2=8.975 $Y2=1.475
r312 73 89 19.2074 $w=3.28e-07 $l=5.5e-07 $layer=LI1_cond $X=8.975 $Y=1.64
+ $X2=8.425 $Y2=1.64
r313 73 74 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.975
+ $Y=1.64 $X2=8.975 $Y2=1.64
r314 70 75 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=10.085 $Y=1.64
+ $X2=10.085 $Y2=1.97
r315 70 73 35.7956 $w=3.28e-07 $l=1.025e-06 $layer=LI1_cond $X=10 $Y=1.64
+ $X2=8.975 $Y2=1.64
r316 69 88 58.0642 $w=1.68e-07 $l=8.9e-07 $layer=LI1_cond $X=7.365 $Y=1.81
+ $X2=8.255 $Y2=1.81
r317 66 69 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.28 $Y=1.895
+ $X2=7.365 $Y2=1.81
r318 66 67 65.8931 $w=1.68e-07 $l=1.01e-06 $layer=LI1_cond $X=7.28 $Y=1.895
+ $X2=7.28 $Y2=2.905
r319 64 67 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.195 $Y=2.99
+ $X2=7.28 $Y2=2.905
r320 64 65 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=7.195 $Y=2.99
+ $X2=6.685 $Y2=2.99
r321 63 65 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.6 $Y=2.905
+ $X2=6.685 $Y2=2.99
r322 62 63 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=6.6 $Y=2.255
+ $X2=6.6 $Y2=2.905
r323 61 87 2.27611 $w=1.7e-07 $l=1.28e-07 $layer=LI1_cond $X=5.73 $Y=2.17
+ $X2=5.602 $Y2=2.17
r324 60 62 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.515 $Y=2.17
+ $X2=6.6 $Y2=2.255
r325 60 61 51.2139 $w=1.68e-07 $l=7.85e-07 $layer=LI1_cond $X=6.515 $Y=2.17
+ $X2=5.73 $Y2=2.17
r326 58 87 5.3732 $w=2.21e-07 $l=1.04307e-07 $layer=LI1_cond $X=5.645 $Y=2.255
+ $X2=5.602 $Y2=2.17
r327 58 59 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=5.645 $Y=2.255
+ $X2=5.645 $Y2=2.895
r328 57 82 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.085 $Y=1.015
+ $X2=5.085 $Y2=1.1
r329 56 57 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=5.085 $Y=0.425
+ $X2=5.085 $Y2=1.015
r330 54 96 17.4861 $w=3.3e-07 $l=1e-07 $layer=POLY_cond $X=4.875 $Y=1.565
+ $X2=4.975 $Y2=1.565
r331 53 54 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.875
+ $Y=1.565 $X2=4.875 $Y2=1.565
r332 51 82 14.5487 $w=1.68e-07 $l=2.23e-07 $layer=LI1_cond $X=4.862 $Y=1.1
+ $X2=5.085 $Y2=1.1
r333 51 53 20.5588 $w=2.03e-07 $l=3.8e-07 $layer=LI1_cond $X=4.862 $Y=1.185
+ $X2=4.862 $Y2=1.565
r334 49 59 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.56 $Y=2.98
+ $X2=5.645 $Y2=2.895
r335 49 50 80.5722 $w=1.68e-07 $l=1.235e-06 $layer=LI1_cond $X=5.56 $Y=2.98
+ $X2=4.325 $Y2=2.98
r336 47 56 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5 $Y=0.34
+ $X2=5.085 $Y2=0.425
r337 47 48 52.1925 $w=1.68e-07 $l=8e-07 $layer=LI1_cond $X=5 $Y=0.34 $X2=4.2
+ $Y2=0.34
r338 43 50 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=4.2 $Y=2.895
+ $X2=4.325 $Y2=2.98
r339 43 45 5.30124 $w=2.48e-07 $l=1.15e-07 $layer=LI1_cond $X=4.2 $Y=2.895
+ $X2=4.2 $Y2=2.78
r340 39 48 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.115 $Y=0.425
+ $X2=4.2 $Y2=0.34
r341 39 41 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=4.115 $Y=0.425
+ $X2=4.115 $Y2=0.515
r342 34 36 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=10.63 $Y=2.465
+ $X2=10.63 $Y2=2.75
r343 33 34 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=10.63 $Y=2.375
+ $X2=10.63 $Y2=2.465
r344 33 107 93.2903 $w=1.8e-07 $l=2.4e-07 $layer=POLY_cond $X=10.63 $Y=2.375
+ $X2=10.63 $Y2=2.135
r345 29 31 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=10.13 $Y=1.085
+ $X2=10.13 $Y2=0.69
r346 28 38 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=9.775 $Y=1.16
+ $X2=9.7 $Y2=1.16
r347 27 29 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=10.055 $Y=1.16
+ $X2=10.13 $Y2=1.085
r348 27 28 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=10.055 $Y=1.16
+ $X2=9.775 $Y2=1.16
r349 24 38 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=9.7 $Y=1.085
+ $X2=9.7 $Y2=1.16
r350 24 26 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=9.7 $Y=1.085
+ $X2=9.7 $Y2=0.69
r351 22 38 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=9.625 $Y=1.16
+ $X2=9.7 $Y2=1.16
r352 22 23 248.691 $w=1.5e-07 $l=4.85e-07 $layer=POLY_cond $X=9.625 $Y=1.16
+ $X2=9.14 $Y2=1.16
r353 20 23 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=9.065 $Y=1.235
+ $X2=9.14 $Y2=1.16
r354 20 103 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=9.065 $Y=1.235
+ $X2=9.065 $Y2=1.475
r355 18 37 330.734 $w=1.5e-07 $l=6.45e-07 $layer=POLY_cond $X=5.64 $Y=0.615
+ $X2=5.64 $Y2=1.26
r356 14 37 37.1337 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=5.625 $Y=1.35
+ $X2=5.625 $Y2=1.26
r357 14 99 89.4032 $w=1.8e-07 $l=2.3e-07 $layer=POLY_cond $X=5.625 $Y=1.35
+ $X2=5.625 $Y2=1.58
r358 12 98 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.4 $Y=1.655
+ $X2=5.565 $Y2=1.655
r359 12 97 171.777 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=5.4 $Y=1.655
+ $X2=5.065 $Y2=1.655
r360 9 11 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=4.975 $Y=2.21
+ $X2=4.975 $Y2=2.495
r361 8 9 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=4.975 $Y=2.12 $X2=4.975
+ $Y2=2.21
r362 7 96 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=4.975 $Y=1.73
+ $X2=4.975 $Y2=1.565
r363 7 8 151.597 $w=1.8e-07 $l=3.9e-07 $layer=POLY_cond $X=4.975 $Y=1.73
+ $X2=4.975 $Y2=2.12
r364 2 45 600 $w=1.7e-07 $l=1.01223e-06 $layer=licon1_PDIFF $count=1 $X=4.01
+ $Y=1.84 $X2=4.16 $Y2=2.78
r365 1 41 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.975
+ $Y=0.37 $X2=4.115 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__SDFSTP_2%A_1185_55# 1 2 7 9 11 12 14 15 19 22 24 25
+ 28 32 34 36 41
c101 34 0 1.75838e-19 $X=6.27 $Y=1.815
c102 12 0 6.64302e-20 $X=6.03 $Y=2.24
c103 7 0 5.96633e-20 $X=6 $Y=0.935
r104 36 38 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=6.855 $Y=0.525
+ $X2=6.855 $Y2=0.615
r105 32 42 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.105 $Y=1.815
+ $X2=6.105 $Y2=1.98
r106 32 41 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.105 $Y=1.815
+ $X2=6.105 $Y2=1.65
r107 31 34 9.43135 $w=1.98e-07 $l=1.65e-07 $layer=LI1_cond $X=6.105 $Y=1.815
+ $X2=6.27 $Y2=1.815
r108 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.105
+ $Y=1.815 $X2=6.105 $Y2=1.815
r109 26 28 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=6.94 $Y=1.915
+ $X2=6.94 $Y2=2.515
r110 24 38 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.69 $Y=0.615
+ $X2=6.855 $Y2=0.615
r111 24 25 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=6.69 $Y=0.615
+ $X2=6.31 $Y2=0.615
r112 22 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.855 $Y=1.83
+ $X2=6.94 $Y2=1.915
r113 22 34 38.1658 $w=1.68e-07 $l=5.85e-07 $layer=LI1_cond $X=6.855 $Y=1.83
+ $X2=6.27 $Y2=1.83
r114 19 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.145
+ $Y=1.1 $X2=6.145 $Y2=1.1
r115 17 25 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=6.145 $Y=0.7
+ $X2=6.31 $Y2=0.615
r116 17 19 13.969 $w=3.28e-07 $l=4e-07 $layer=LI1_cond $X=6.145 $Y=0.7 $X2=6.145
+ $Y2=1.1
r117 15 20 38.8445 $w=3.55e-07 $l=1.93533e-07 $layer=POLY_cond $X=6.055 $Y=1.265
+ $X2=6.117 $Y2=1.1
r118 15 41 197.415 $w=1.5e-07 $l=3.85e-07 $layer=POLY_cond $X=6.055 $Y=1.265
+ $X2=6.055 $Y2=1.65
r119 12 14 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=6.03 $Y=2.24
+ $X2=6.03 $Y2=2.525
r120 11 12 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=6.03 $Y=2.15 $X2=6.03
+ $Y2=2.24
r121 11 42 66.0806 $w=1.8e-07 $l=1.7e-07 $layer=POLY_cond $X=6.03 $Y=2.15
+ $X2=6.03 $Y2=1.98
r122 7 20 38.8445 $w=3.55e-07 $l=2.15708e-07 $layer=POLY_cond $X=6 $Y=0.935
+ $X2=6.117 $Y2=1.1
r123 7 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=6 $Y=0.935 $X2=6
+ $Y2=0.615
r124 2 28 600 $w=1.7e-07 $l=2.64575e-07 $layer=licon1_PDIFF $count=1 $X=6.79
+ $Y=2.315 $X2=6.94 $Y2=2.515
r125 1 36 182 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_NDIFF $count=1 $X=6.71
+ $Y=0.37 $X2=6.855 $Y2=0.525
.ends

.subckt PM_SKY130_FD_SC_HS__SDFSTP_2%A_991_81# 1 2 7 8 9 11 12 14 16 17 19 20 22
+ 24 25 27 28 30 34 37 39 45 47 48 52 53 54 55 58 63 65 71
c195 58 0 6.64302e-20 $X=5.24 $Y=2.265
c196 55 0 5.96633e-20 $X=6.88 $Y=0.955
c197 45 0 2.09475e-20 $X=5.425 $Y=0.615
c198 37 0 1.3233e-19 $X=5.24 $Y=2.39
c199 34 0 2.52187e-20 $X=7.07 $Y=0.94
c200 8 0 2.91132e-19 $X=6.715 $Y=2.15
r201 70 71 24.0272 $w=3.31e-07 $l=1.65e-07 $layer=POLY_cond $X=8.13 $Y=1.32
+ $X2=8.295 $Y2=1.32
r202 64 70 30.5801 $w=3.31e-07 $l=2.1e-07 $layer=POLY_cond $X=7.92 $Y=1.32
+ $X2=8.13 $Y2=1.32
r203 64 68 10.9215 $w=3.31e-07 $l=7.5e-08 $layer=POLY_cond $X=7.92 $Y=1.32
+ $X2=7.845 $Y2=1.32
r204 63 65 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=7.92 $Y=1.39
+ $X2=7.92 $Y2=1.225
r205 63 64 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.92
+ $Y=1.39 $X2=7.92 $Y2=1.39
r206 56 65 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=7.84 $Y=1.04
+ $X2=7.84 $Y2=1.225
r207 54 56 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.755 $Y=0.955
+ $X2=7.84 $Y2=1.04
r208 54 55 57.0856 $w=1.68e-07 $l=8.75e-07 $layer=LI1_cond $X=7.755 $Y=0.955
+ $X2=6.88 $Y2=0.955
r209 52 53 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.715
+ $Y=1.065 $X2=6.715 $Y2=1.065
r210 50 52 10.826 $w=3.28e-07 $l=3.1e-07 $layer=LI1_cond $X=6.715 $Y=1.375
+ $X2=6.715 $Y2=1.065
r211 49 55 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=6.715 $Y=1.04
+ $X2=6.88 $Y2=0.955
r212 49 52 0.873063 $w=3.28e-07 $l=2.5e-08 $layer=LI1_cond $X=6.715 $Y=1.04
+ $X2=6.715 $Y2=1.065
r213 47 50 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=6.55 $Y=1.46
+ $X2=6.715 $Y2=1.375
r214 47 48 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=6.55 $Y=1.46
+ $X2=5.59 $Y2=1.46
r215 43 48 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=5.465 $Y=1.46
+ $X2=5.59 $Y2=1.46
r216 43 59 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=5.465 $Y=1.46
+ $X2=5.22 $Y2=1.46
r217 43 45 35.0343 $w=2.48e-07 $l=7.6e-07 $layer=LI1_cond $X=5.465 $Y=1.375
+ $X2=5.465 $Y2=0.615
r218 41 59 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.22 $Y=1.545
+ $X2=5.22 $Y2=1.46
r219 41 58 46.9733 $w=1.68e-07 $l=7.2e-07 $layer=LI1_cond $X=5.22 $Y=1.545
+ $X2=5.22 $Y2=2.265
r220 37 58 6.55365 $w=2.48e-07 $l=1.25e-07 $layer=LI1_cond $X=5.24 $Y=2.39
+ $X2=5.24 $Y2=2.265
r221 37 39 4.84026 $w=2.48e-07 $l=1.05e-07 $layer=LI1_cond $X=5.24 $Y=2.39
+ $X2=5.24 $Y2=2.495
r222 36 53 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=6.715 $Y=1.405
+ $X2=6.715 $Y2=1.065
r223 32 53 8.74306 $w=3.3e-07 $l=5e-08 $layer=POLY_cond $X=6.715 $Y=1.015
+ $X2=6.715 $Y2=1.065
r224 32 34 182.032 $w=1.5e-07 $l=3.55e-07 $layer=POLY_cond $X=6.715 $Y=0.94
+ $X2=7.07 $Y2=0.94
r225 28 71 38.5891 $w=3.31e-07 $l=3.64005e-07 $layer=POLY_cond $X=8.56 $Y=1.085
+ $X2=8.295 $Y2=1.32
r226 28 30 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=8.56 $Y=1.085
+ $X2=8.56 $Y2=0.69
r227 25 27 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=8.295 $Y=1.82
+ $X2=8.295 $Y2=2.315
r228 24 25 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=8.295 $Y=1.73
+ $X2=8.295 $Y2=1.82
r229 23 71 17.0024 $w=1.8e-07 $l=2.35e-07 $layer=POLY_cond $X=8.295 $Y=1.555
+ $X2=8.295 $Y2=1.32
r230 23 24 68.0242 $w=1.8e-07 $l=1.75e-07 $layer=POLY_cond $X=8.295 $Y=1.555
+ $X2=8.295 $Y2=1.73
r231 20 70 21.295 $w=1.5e-07 $l=2.35e-07 $layer=POLY_cond $X=8.13 $Y=1.085
+ $X2=8.13 $Y2=1.32
r232 20 22 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=8.13 $Y=1.085
+ $X2=8.13 $Y2=0.69
r233 17 19 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=7.845 $Y=1.82
+ $X2=7.845 $Y2=2.315
r234 16 17 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=7.845 $Y=1.73
+ $X2=7.845 $Y2=1.82
r235 15 68 17.0024 $w=1.8e-07 $l=2.35e-07 $layer=POLY_cond $X=7.845 $Y=1.555
+ $X2=7.845 $Y2=1.32
r236 15 16 68.0242 $w=1.8e-07 $l=1.75e-07 $layer=POLY_cond $X=7.845 $Y=1.555
+ $X2=7.845 $Y2=1.73
r237 12 34 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.07 $Y=0.865
+ $X2=7.07 $Y2=0.94
r238 12 14 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=7.07 $Y=0.865
+ $X2=7.07 $Y2=0.58
r239 9 11 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=6.715 $Y=2.24
+ $X2=6.715 $Y2=2.525
r240 8 9 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=6.715 $Y=2.15 $X2=6.715
+ $Y2=2.24
r241 7 36 34.7712 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.715 $Y=1.57
+ $X2=6.715 $Y2=1.405
r242 7 8 225.452 $w=1.8e-07 $l=5.8e-07 $layer=POLY_cond $X=6.715 $Y=1.57
+ $X2=6.715 $Y2=2.15
r243 2 39 600 $w=1.7e-07 $l=2.74955e-07 $layer=licon1_PDIFF $count=1 $X=5.05
+ $Y=2.285 $X2=5.2 $Y2=2.495
r244 1 45 182 $w=1.7e-07 $l=5.65332e-07 $layer=licon1_NDIFF $count=1 $X=4.955
+ $Y=0.405 $X2=5.425 $Y2=0.615
.ends

.subckt PM_SKY130_FD_SC_HS__SDFSTP_2%SET_B 2 3 5 8 11 12 14 17 19 20 23 25 32 35
+ 43
c143 25 0 5.34496e-20 $X=11.76 $Y=1.295
c144 17 0 7.44554e-20 $X=11.59 $Y=0.58
c145 12 0 5.57434e-20 $X=11.47 $Y=2.465
c146 11 0 3.15842e-21 $X=11.47 $Y=2.375
c147 8 0 1.09822e-19 $X=7.46 $Y=0.58
r148 36 43 9.11234 $w=4.28e-07 $l=3.4e-07 $layer=LI1_cond $X=11.66 $Y=1.635
+ $X2=11.66 $Y2=1.295
r149 35 38 39.8861 $w=3.95e-07 $l=1.65e-07 $layer=POLY_cond $X=11.577 $Y=1.635
+ $X2=11.577 $Y2=1.8
r150 35 37 45.5639 $w=3.95e-07 $l=1.65e-07 $layer=POLY_cond $X=11.577 $Y=1.635
+ $X2=11.577 $Y2=1.47
r151 35 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=11.61
+ $Y=1.635 $X2=11.61 $Y2=1.635
r152 30 32 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=7.37 $Y=1.39 $X2=7.46
+ $Y2=1.39
r153 27 30 27.9778 $w=3.3e-07 $l=1.6e-07 $layer=POLY_cond $X=7.21 $Y=1.39
+ $X2=7.37 $Y2=1.39
r154 25 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.76 $Y=1.295
+ $X2=11.76 $Y2=1.295
r155 23 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.37
+ $Y=1.39 $X2=7.37 $Y2=1.39
r156 22 23 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=1.295
+ $X2=7.44 $Y2=1.295
r157 20 22 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=7.585 $Y=1.295
+ $X2=7.44 $Y2=1.295
r158 19 25 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=11.615 $Y=1.295
+ $X2=11.76 $Y2=1.295
r159 19 20 4.98761 $w=1.4e-07 $l=4.03e-06 $layer=MET1_cond $X=11.615 $Y=1.295
+ $X2=7.585 $Y2=1.295
r160 17 37 456.362 $w=1.5e-07 $l=8.9e-07 $layer=POLY_cond $X=11.59 $Y=0.58
+ $X2=11.59 $Y2=1.47
r161 12 14 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=11.47 $Y=2.465
+ $X2=11.47 $Y2=2.75
r162 11 12 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=11.47 $Y=2.375
+ $X2=11.47 $Y2=2.465
r163 11 38 223.508 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=11.47 $Y=2.375
+ $X2=11.47 $Y2=1.8
r164 6 32 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.46 $Y=1.225
+ $X2=7.46 $Y2=1.39
r165 6 8 330.734 $w=1.5e-07 $l=6.45e-07 $layer=POLY_cond $X=7.46 $Y=1.225
+ $X2=7.46 $Y2=0.58
r166 3 5 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=7.21 $Y=2.24 $X2=7.21
+ $Y2=2.525
r167 2 3 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=7.21 $Y=2.15 $X2=7.21
+ $Y2=2.24
r168 1 27 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=7.21 $Y=1.555
+ $X2=7.21 $Y2=1.39
r169 1 2 231.282 $w=1.8e-07 $l=5.95e-07 $layer=POLY_cond $X=7.21 $Y=1.555
+ $X2=7.21 $Y2=2.15
.ends

.subckt PM_SKY130_FD_SC_HS__SDFSTP_2%A_608_74# 1 2 9 11 13 15 16 19 20 21 22 23
+ 26 28 30 31 34 35 38 39 40 41 43 45 48 50 51 52 54 57 60 61 62 67 70
c207 54 0 1.37364e-19 $X=9.44 $Y=3.13
c208 35 0 2.15509e-19 $X=9.44 $Y=2.045
c209 20 0 2.09475e-20 $X=4.805 $Y=1.115
r210 71 72 4.79261 $w=3.52e-07 $l=3.5e-08 $layer=POLY_cond $X=3.9 $Y=1.557
+ $X2=3.935 $Y2=1.557
r211 68 72 15.7472 $w=3.52e-07 $l=1.15e-07 $layer=POLY_cond $X=4.05 $Y=1.557
+ $X2=3.935 $Y2=1.557
r212 67 68 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.05
+ $Y=1.515 $X2=4.05 $Y2=1.515
r213 65 67 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=4.05 $Y=1.82
+ $X2=4.05 $Y2=1.515
r214 62 64 5.9927 $w=2.48e-07 $l=1.3e-07 $layer=LI1_cond $X=3.13 $Y=1.945
+ $X2=3.26 $Y2=1.945
r215 61 65 6.98653 $w=2.5e-07 $l=2.18746e-07 $layer=LI1_cond $X=3.885 $Y=1.945
+ $X2=4.05 $Y2=1.82
r216 61 64 28.8111 $w=2.48e-07 $l=6.25e-07 $layer=LI1_cond $X=3.885 $Y=1.945
+ $X2=3.26 $Y2=1.945
r217 60 62 7.14316 $w=2.5e-07 $l=1.62019e-07 $layer=LI1_cond $X=3.045 $Y=1.82
+ $X2=3.13 $Y2=1.945
r218 60 70 52.8449 $w=1.68e-07 $l=8.1e-07 $layer=LI1_cond $X=3.045 $Y=1.82
+ $X2=3.045 $Y2=1.01
r219 55 70 9.49412 $w=3.88e-07 $l=1.95e-07 $layer=LI1_cond $X=3.155 $Y=0.815
+ $X2=3.155 $Y2=1.01
r220 55 57 8.86495 $w=3.88e-07 $l=3e-07 $layer=LI1_cond $X=3.155 $Y=0.815
+ $X2=3.155 $Y2=0.515
r221 50 51 58.3064 $w=1.8e-07 $l=1.5e-07 $layer=POLY_cond $X=4.44 $Y=1.97
+ $X2=4.44 $Y2=2.12
r222 46 48 443.543 $w=1.5e-07 $l=8.65e-07 $layer=POLY_cond $X=10.63 $Y=1.445
+ $X2=10.63 $Y2=0.58
r223 43 45 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=9.89 $Y=3.035
+ $X2=9.89 $Y2=2.54
r224 42 54 20.4101 $w=1.5e-07 $l=9.94987e-08 $layer=POLY_cond $X=9.53 $Y=3.15
+ $X2=9.44 $Y2=3.13
r225 41 43 26.9307 $w=1.5e-07 $l=1.53542e-07 $layer=POLY_cond $X=9.8 $Y=3.15
+ $X2=9.89 $Y2=3.035
r226 41 42 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=9.8 $Y=3.15
+ $X2=9.53 $Y2=3.15
r227 39 46 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=10.555 $Y=1.52
+ $X2=10.63 $Y2=1.445
r228 39 40 525.585 $w=1.5e-07 $l=1.025e-06 $layer=POLY_cond $X=10.555 $Y=1.52
+ $X2=9.53 $Y2=1.52
r229 36 54 5.30422 $w=1.5e-07 $l=9.5e-08 $layer=POLY_cond $X=9.44 $Y=3.035
+ $X2=9.44 $Y2=3.13
r230 36 38 253.819 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=9.44 $Y=3.035
+ $X2=9.44 $Y2=2.54
r231 35 38 253.819 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=9.44 $Y=2.045
+ $X2=9.44 $Y2=2.54
r232 34 35 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=9.44 $Y=1.955
+ $X2=9.44 $Y2=2.045
r233 33 40 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=9.44 $Y=1.595
+ $X2=9.53 $Y2=1.52
r234 33 34 139.935 $w=1.8e-07 $l=3.6e-07 $layer=POLY_cond $X=9.44 $Y=1.595
+ $X2=9.44 $Y2=1.955
r235 32 52 7.1379 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=5.6 $Y=3.15 $X2=5.51
+ $Y2=3.15
r236 31 54 20.4101 $w=1.5e-07 $l=9.94987e-08 $layer=POLY_cond $X=9.35 $Y=3.15
+ $X2=9.44 $Y2=3.13
r237 31 32 1922.87 $w=1.5e-07 $l=3.75e-06 $layer=POLY_cond $X=9.35 $Y=3.15
+ $X2=5.6 $Y2=3.15
r238 28 52 95.4401 $w=1.8e-07 $l=2.4e-07 $layer=POLY_cond $X=5.51 $Y=2.91
+ $X2=5.51 $Y2=3.15
r239 28 30 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=5.51 $Y=2.91
+ $X2=5.51 $Y2=2.625
r240 24 26 217.926 $w=1.5e-07 $l=4.25e-07 $layer=POLY_cond $X=4.88 $Y=1.04
+ $X2=4.88 $Y2=0.615
r241 22 52 7.1379 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=5.42 $Y=3.15 $X2=5.51
+ $Y2=3.15
r242 22 23 456.362 $w=1.5e-07 $l=8.9e-07 $layer=POLY_cond $X=5.42 $Y=3.15
+ $X2=4.53 $Y2=3.15
r243 20 24 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.805 $Y=1.115
+ $X2=4.88 $Y2=1.04
r244 20 21 156.394 $w=1.5e-07 $l=3.05e-07 $layer=POLY_cond $X=4.805 $Y=1.115
+ $X2=4.5 $Y2=1.115
r245 19 23 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.455 $Y=3.075
+ $X2=4.53 $Y2=3.15
r246 19 51 489.691 $w=1.5e-07 $l=9.55e-07 $layer=POLY_cond $X=4.455 $Y=3.075
+ $X2=4.455 $Y2=2.12
r247 16 68 51.3494 $w=3.52e-07 $l=3.75e-07 $layer=POLY_cond $X=4.425 $Y=1.557
+ $X2=4.05 $Y2=1.557
r248 16 50 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=4.425 $Y=1.68
+ $X2=4.425 $Y2=1.97
r249 15 16 22.7654 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.425 $Y=1.35
+ $X2=4.425 $Y2=1.557
r250 14 21 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.425 $Y=1.19
+ $X2=4.5 $Y2=1.115
r251 14 15 82.0426 $w=1.5e-07 $l=1.6e-07 $layer=POLY_cond $X=4.425 $Y=1.19
+ $X2=4.425 $Y2=1.35
r252 11 72 22.7654 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=3.935 $Y=1.765
+ $X2=3.935 $Y2=1.557
r253 11 13 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.935 $Y=1.765
+ $X2=3.935 $Y2=2.4
r254 7 71 22.7654 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.9 $Y=1.35 $X2=3.9
+ $Y2=1.557
r255 7 9 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=3.9 $Y=1.35 $X2=3.9
+ $Y2=0.74
r256 2 64 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=3.125
+ $Y=1.84 $X2=3.26 $Y2=1.985
r257 1 57 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=3.04
+ $Y=0.37 $X2=3.185 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__SDFSTP_2%A_2186_367# 1 2 7 8 11 12 14 17 18 22 24 25
+ 28 31 32 36 38 40
c111 36 0 6.56335e-20 $X=11.11 $Y=1.065
c112 25 0 5.57434e-20 $X=12.31 $Y=2.395
c113 17 0 3.1683e-20 $X=11.02 $Y=1.835
c114 8 0 1.88308e-19 $X=11.02 $Y=2.375
c115 7 0 1.557e-19 $X=11.02 $Y=1.925
r116 36 41 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=11.11 $Y=1.065
+ $X2=11.11 $Y2=1.23
r117 36 40 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=11.11 $Y=1.065
+ $X2=11.11 $Y2=0.9
r118 35 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=11.11
+ $Y=1.065 $X2=11.11 $Y2=1.065
r119 32 35 6.63528 $w=3.28e-07 $l=1.9e-07 $layer=LI1_cond $X=11.11 $Y=0.875
+ $X2=11.11 $Y2=1.065
r120 30 38 3.87901 $w=2.37e-07 $l=1.14039e-07 $layer=LI1_cond $X=12.72 $Y=0.96
+ $X2=12.652 $Y2=0.875
r121 30 31 88.0749 $w=1.68e-07 $l=1.35e-06 $layer=LI1_cond $X=12.72 $Y=0.96
+ $X2=12.72 $Y2=2.31
r122 26 38 3.87901 $w=2.37e-07 $l=8.5e-08 $layer=LI1_cond $X=12.652 $Y=0.79
+ $X2=12.652 $Y2=0.875
r123 26 28 7.93485 $w=3.03e-07 $l=2.1e-07 $layer=LI1_cond $X=12.652 $Y=0.79
+ $X2=12.652 $Y2=0.58
r124 24 31 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=12.635 $Y=2.395
+ $X2=12.72 $Y2=2.31
r125 24 25 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=12.635 $Y=2.395
+ $X2=12.31 $Y2=2.395
r126 20 25 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=12.185 $Y=2.48
+ $X2=12.31 $Y2=2.395
r127 20 22 12.4464 $w=2.48e-07 $l=2.7e-07 $layer=LI1_cond $X=12.185 $Y=2.48
+ $X2=12.185 $Y2=2.75
r128 19 32 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.275 $Y=0.875
+ $X2=11.11 $Y2=0.875
r129 18 38 2.57001 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=12.5 $Y=0.875
+ $X2=12.652 $Y2=0.875
r130 18 19 79.9198 $w=1.68e-07 $l=1.225e-06 $layer=LI1_cond $X=12.5 $Y=0.875
+ $X2=11.275 $Y2=0.875
r131 17 41 310.223 $w=1.5e-07 $l=6.05e-07 $layer=POLY_cond $X=11.035 $Y=1.835
+ $X2=11.035 $Y2=1.23
r132 12 14 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=11.02 $Y=2.465
+ $X2=11.02 $Y2=2.75
r133 11 40 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=11.02 $Y=0.58
+ $X2=11.02 $Y2=0.9
r134 8 12 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=11.02 $Y=2.375
+ $X2=11.02 $Y2=2.465
r135 7 17 37.1337 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=11.02 $Y=1.925
+ $X2=11.02 $Y2=1.835
r136 7 8 174.919 $w=1.8e-07 $l=4.5e-07 $layer=POLY_cond $X=11.02 $Y=1.925
+ $X2=11.02 $Y2=2.375
r137 2 22 600 $w=1.7e-07 $l=2.67208e-07 $layer=licon1_PDIFF $count=1 $X=12.095
+ $Y=2.54 $X2=12.225 $Y2=2.75
r138 1 28 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=12.5
+ $Y=0.37 $X2=12.64 $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_HS__SDFSTP_2%A_1804_424# 1 2 3 4 5 18 21 22 24 25 27 29
+ 31 32 34 37 38 41 43 44 45 50 54 56 58 59 60 62 65 67 69 71 72 74 79 81 83 86
c205 59 0 1.93538e-19 $X=10.89 $Y=1.485
c206 38 0 5.67555e-20 $X=13.43 $Y=1.365
r207 86 87 66.7385 $w=3.75e-07 $l=4.5e-07 $layer=POLY_cond $X=12.322 $Y=1.975
+ $X2=12.322 $Y2=1.525
r208 85 86 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=12.3
+ $Y=1.975 $X2=12.3 $Y2=1.975
r209 82 83 9.54788 $w=5.03e-07 $l=1.65e-07 $layer=LI1_cond $X=11.695 $Y=2.222
+ $X2=11.86 $Y2=2.222
r210 74 77 6.63528 $w=3.28e-07 $l=1.9e-07 $layer=LI1_cond $X=9.415 $Y=0.34
+ $X2=9.415 $Y2=0.53
r211 72 87 23.988 $w=2.62e-07 $l=1.98e-07 $layer=POLY_cond $X=12.322 $Y=1.327
+ $X2=12.322 $Y2=1.525
r212 71 72 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=12.3
+ $Y=1.295 $X2=12.3 $Y2=1.295
r213 69 85 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=12.3 $Y=1.97 $X2=12.3
+ $Y2=2.055
r214 69 71 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=12.3 $Y=1.97
+ $X2=12.3 $Y2=1.295
r215 67 85 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12.135 $Y=2.055
+ $X2=12.3 $Y2=2.055
r216 67 83 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=12.135 $Y=2.055
+ $X2=11.86 $Y2=2.055
r217 63 82 3.22715 $w=3.3e-07 $l=2.53e-07 $layer=LI1_cond $X=11.695 $Y=2.475
+ $X2=11.695 $Y2=2.222
r218 63 65 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=11.695 $Y=2.475
+ $X2=11.695 $Y2=2.75
r219 62 82 17.053 $w=5.03e-07 $l=7.2e-07 $layer=LI1_cond $X=10.975 $Y=2.222
+ $X2=11.695 $Y2=2.222
r220 62 81 7.65311 $w=5.03e-07 $l=8.5e-08 $layer=LI1_cond $X=10.975 $Y=2.222
+ $X2=10.89 $Y2=2.222
r221 61 62 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=10.975 $Y=1.57
+ $X2=10.975 $Y2=1.97
r222 59 61 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=10.89 $Y=1.485
+ $X2=10.975 $Y2=1.57
r223 59 60 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=10.89 $Y=1.485
+ $X2=10.58 $Y2=1.485
r224 58 81 29.6845 $w=1.68e-07 $l=4.55e-07 $layer=LI1_cond $X=10.435 $Y=2.39
+ $X2=10.89 $Y2=2.39
r225 56 60 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=10.495 $Y=1.4
+ $X2=10.58 $Y2=1.485
r226 56 79 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=10.495 $Y=1.4
+ $X2=10.495 $Y2=0.81
r227 52 79 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=10.415 $Y=0.645
+ $X2=10.415 $Y2=0.81
r228 52 54 2.26996 $w=3.28e-07 $l=6.5e-08 $layer=LI1_cond $X=10.415 $Y=0.645
+ $X2=10.415 $Y2=0.58
r229 51 54 5.41299 $w=3.28e-07 $l=1.55e-07 $layer=LI1_cond $X=10.415 $Y=0.425
+ $X2=10.415 $Y2=0.58
r230 48 50 5.5876 $w=3.28e-07 $l=1.6e-07 $layer=LI1_cond $X=10.27 $Y=2.905
+ $X2=10.27 $Y2=2.745
r231 47 58 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=10.27 $Y=2.475
+ $X2=10.435 $Y2=2.39
r232 47 50 9.42908 $w=3.28e-07 $l=2.7e-07 $layer=LI1_cond $X=10.27 $Y=2.475
+ $X2=10.27 $Y2=2.745
r233 46 74 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.58 $Y=0.34
+ $X2=9.415 $Y2=0.34
r234 45 51 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=10.25 $Y=0.34
+ $X2=10.415 $Y2=0.425
r235 45 46 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=10.25 $Y=0.34
+ $X2=9.58 $Y2=0.34
r236 43 48 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=10.105 $Y=2.99
+ $X2=10.27 $Y2=2.905
r237 43 44 50.5615 $w=1.68e-07 $l=7.75e-07 $layer=LI1_cond $X=10.105 $Y=2.99
+ $X2=9.33 $Y2=2.99
r238 39 44 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=9.165 $Y=2.905
+ $X2=9.33 $Y2=2.99
r239 39 41 17.6359 $w=3.28e-07 $l=5.05e-07 $layer=LI1_cond $X=9.165 $Y=2.905
+ $X2=9.165 $Y2=2.4
r240 36 86 2.22462 $w=3.75e-07 $l=1.5e-08 $layer=POLY_cond $X=12.322 $Y=1.99
+ $X2=12.322 $Y2=1.975
r241 36 37 37.3423 $w=3.75e-07 $l=1.5e-07 $layer=POLY_cond $X=12.337 $Y=1.99
+ $X2=12.337 $Y2=2.14
r242 32 34 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=13.43 $Y=1.885
+ $X2=13.43 $Y2=2.46
r243 31 32 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=13.43 $Y=1.795
+ $X2=13.43 $Y2=1.885
r244 30 38 33.9972 $w=1.65e-07 $l=1.6e-07 $layer=POLY_cond $X=13.43 $Y=1.525
+ $X2=13.43 $Y2=1.365
r245 30 31 104.952 $w=1.8e-07 $l=2.7e-07 $layer=POLY_cond $X=13.43 $Y=1.525
+ $X2=13.43 $Y2=1.795
r246 27 38 33.9972 $w=1.65e-07 $l=1.67332e-07 $layer=POLY_cond $X=13.415
+ $Y=1.205 $X2=13.43 $Y2=1.365
r247 27 29 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=13.415 $Y=1.205
+ $X2=13.415 $Y2=0.81
r248 26 72 2.52859 $w=3.2e-07 $l=2.06126e-07 $layer=POLY_cond $X=12.51 $Y=1.365
+ $X2=12.322 $Y2=1.327
r249 25 38 3.5291 $w=3.2e-07 $l=9e-08 $layer=POLY_cond $X=13.34 $Y=1.365
+ $X2=13.43 $Y2=1.365
r250 25 26 149.67 $w=3.2e-07 $l=8.3e-07 $layer=POLY_cond $X=13.34 $Y=1.365
+ $X2=12.51 $Y2=1.365
r251 22 24 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=12.45 $Y=2.465
+ $X2=12.45 $Y2=2.75
r252 21 22 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=12.45 $Y=2.375
+ $X2=12.45 $Y2=2.465
r253 21 37 91.3468 $w=1.8e-07 $l=2.35e-07 $layer=POLY_cond $X=12.45 $Y=2.375
+ $X2=12.45 $Y2=2.14
r254 16 72 23.988 $w=2.62e-07 $l=2.43105e-07 $layer=POLY_cond $X=12.425 $Y=1.13
+ $X2=12.322 $Y2=1.327
r255 16 18 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=12.425 $Y=1.13
+ $X2=12.425 $Y2=0.58
r256 5 65 600 $w=1.7e-07 $l=2.74955e-07 $layer=licon1_PDIFF $count=1 $X=11.545
+ $Y=2.54 $X2=11.695 $Y2=2.75
r257 4 50 600 $w=1.7e-07 $l=7.62398e-07 $layer=licon1_PDIFF $count=1 $X=9.965
+ $Y=2.12 $X2=10.27 $Y2=2.745
r258 3 41 300 $w=1.7e-07 $l=3.44964e-07 $layer=licon1_PDIFF $count=2 $X=9.02
+ $Y=2.12 $X2=9.165 $Y2=2.4
r259 2 54 182 $w=1.7e-07 $l=2.96985e-07 $layer=licon1_NDIFF $count=1 $X=10.205
+ $Y=0.37 $X2=10.415 $Y2=0.58
r260 1 77 182 $w=1.7e-07 $l=2.20907e-07 $layer=licon1_NDIFF $count=1 $X=9.27
+ $Y=0.37 $X2=9.415 $Y2=0.53
.ends

.subckt PM_SKY130_FD_SC_HS__SDFSTP_2%A_2611_98# 1 2 7 9 12 14 16 17 19 22 26 32
+ 35 39
c80 26 0 7.29682e-20 $X=13.205 $Y=2.105
r81 39 40 1.75061 $w=4.13e-07 $l=1.5e-08 $layer=POLY_cond $X=14.37 $Y=1.485
+ $X2=14.385 $Y2=1.485
r82 33 37 4.66828 $w=4.13e-07 $l=4e-08 $layer=POLY_cond $X=13.895 $Y=1.485
+ $X2=13.935 $Y2=1.485
r83 32 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=13.895
+ $Y=1.485 $X2=13.895 $Y2=1.485
r84 30 35 1.36975 $w=3.3e-07 $l=1.68e-07 $layer=LI1_cond $X=13.37 $Y=1.485
+ $X2=13.202 $Y2=1.485
r85 30 32 18.3343 $w=3.28e-07 $l=5.25e-07 $layer=LI1_cond $X=13.37 $Y=1.485
+ $X2=13.895 $Y2=1.485
r86 26 28 24.4249 $w=3.33e-07 $l=7.1e-07 $layer=LI1_cond $X=13.202 $Y=2.105
+ $X2=13.202 $Y2=2.815
r87 24 35 5.13366 $w=3.32e-07 $l=1.65e-07 $layer=LI1_cond $X=13.202 $Y=1.65
+ $X2=13.202 $Y2=1.485
r88 24 26 15.6526 $w=3.33e-07 $l=4.55e-07 $layer=LI1_cond $X=13.202 $Y=1.65
+ $X2=13.202 $Y2=2.105
r89 20 35 5.13366 $w=3.32e-07 $l=1.65997e-07 $layer=LI1_cond $X=13.2 $Y=1.32
+ $X2=13.202 $Y2=1.485
r90 20 22 23.9219 $w=3.28e-07 $l=6.85e-07 $layer=LI1_cond $X=13.2 $Y=1.32
+ $X2=13.2 $Y2=0.635
r91 17 40 26.6457 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=14.385 $Y=1.765
+ $X2=14.385 $Y2=1.485
r92 17 19 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=14.385 $Y=1.765
+ $X2=14.385 $Y2=2.4
r93 14 39 26.6457 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=14.37 $Y=1.205
+ $X2=14.37 $Y2=1.485
r94 14 16 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=14.37 $Y=1.205
+ $X2=14.37 $Y2=0.76
r95 10 39 50.184 $w=4.13e-07 $l=4.3e-07 $layer=POLY_cond $X=13.94 $Y=1.485
+ $X2=14.37 $Y2=1.485
r96 10 37 0.583535 $w=4.13e-07 $l=5e-09 $layer=POLY_cond $X=13.94 $Y=1.485
+ $X2=13.935 $Y2=1.485
r97 10 12 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=13.94 $Y=1.32
+ $X2=13.94 $Y2=0.76
r98 7 37 26.6457 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=13.935 $Y=1.765
+ $X2=13.935 $Y2=1.485
r99 7 9 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=13.935 $Y=1.765
+ $X2=13.935 $Y2=2.4
r100 2 28 400 $w=1.7e-07 $l=9.17701e-07 $layer=licon1_PDIFF $count=1 $X=13.075
+ $Y=1.96 $X2=13.205 $Y2=2.815
r101 2 26 400 $w=1.7e-07 $l=1.99687e-07 $layer=licon1_PDIFF $count=1 $X=13.075
+ $Y=1.96 $X2=13.205 $Y2=2.105
r102 1 22 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=13.055
+ $Y=0.49 $X2=13.2 $Y2=0.635
.ends

.subckt PM_SKY130_FD_SC_HS__SDFSTP_2%VPWR 1 2 3 4 5 6 7 8 9 10 33 37 39 43 47 51
+ 55 59 63 67 71 73 76 77 79 80 82 83 84 86 91 112 119 124 129 135 138 141 144
+ 147 150 154
c186 55 0 1.72142e-19 $X=8.52 $Y=2.58
r187 153 154 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=14.64 $Y=3.33
+ $X2=14.64 $Y2=3.33
r188 150 151 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.68 $Y=3.33
+ $X2=13.68 $Y2=3.33
r189 147 148 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.72 $Y=3.33
+ $X2=12.72 $Y2=3.33
r190 144 145 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=11.28 $Y=3.33
+ $X2=11.28 $Y2=3.33
r191 141 142 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r192 139 142 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.6 $Y2=3.33
r193 138 139 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r194 135 136 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r195 133 154 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=14.16 $Y=3.33
+ $X2=14.64 $Y2=3.33
r196 133 151 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=14.16 $Y=3.33
+ $X2=13.68 $Y2=3.33
r197 132 133 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=14.16 $Y=3.33
+ $X2=14.16 $Y2=3.33
r198 130 150 7.75133 $w=1.7e-07 $l=1.43e-07 $layer=LI1_cond $X=13.825 $Y=3.33
+ $X2=13.682 $Y2=3.33
r199 130 132 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=13.825 $Y=3.33
+ $X2=14.16 $Y2=3.33
r200 129 153 4.76062 $w=1.7e-07 $l=2.17e-07 $layer=LI1_cond $X=14.445 $Y=3.33
+ $X2=14.662 $Y2=3.33
r201 129 132 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=14.445 $Y=3.33
+ $X2=14.16 $Y2=3.33
r202 128 151 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=13.2 $Y=3.33
+ $X2=13.68 $Y2=3.33
r203 128 148 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=13.2 $Y=3.33
+ $X2=12.72 $Y2=3.33
r204 127 128 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.2 $Y=3.33
+ $X2=13.2 $Y2=3.33
r205 125 147 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12.84 $Y=3.33
+ $X2=12.675 $Y2=3.33
r206 125 127 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=12.84 $Y=3.33
+ $X2=13.2 $Y2=3.33
r207 124 150 7.75133 $w=1.7e-07 $l=1.42e-07 $layer=LI1_cond $X=13.54 $Y=3.33
+ $X2=13.682 $Y2=3.33
r208 124 127 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=13.54 $Y=3.33
+ $X2=13.2 $Y2=3.33
r209 123 148 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.24 $Y=3.33
+ $X2=12.72 $Y2=3.33
r210 123 145 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=12.24 $Y=3.33
+ $X2=11.28 $Y2=3.33
r211 122 123 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=12.24 $Y=3.33
+ $X2=12.24 $Y2=3.33
r212 120 144 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=11.33 $Y=3.33
+ $X2=11.205 $Y2=3.33
r213 120 122 59.369 $w=1.68e-07 $l=9.1e-07 $layer=LI1_cond $X=11.33 $Y=3.33
+ $X2=12.24 $Y2=3.33
r214 119 147 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12.51 $Y=3.33
+ $X2=12.675 $Y2=3.33
r215 119 122 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=12.51 $Y=3.33
+ $X2=12.24 $Y2=3.33
r216 118 145 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.8 $Y=3.33
+ $X2=11.28 $Y2=3.33
r217 117 118 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=10.8 $Y=3.33
+ $X2=10.8 $Y2=3.33
r218 115 118 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=8.88 $Y=3.33
+ $X2=10.8 $Y2=3.33
r219 114 117 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=8.88 $Y=3.33
+ $X2=10.8 $Y2=3.33
r220 114 115 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r221 112 144 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=11.08 $Y=3.33
+ $X2=11.205 $Y2=3.33
r222 112 117 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=11.08 $Y=3.33
+ $X2=10.8 $Y2=3.33
r223 111 115 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=3.33
+ $X2=8.88 $Y2=3.33
r224 110 111 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.4 $Y=3.33
+ $X2=8.4 $Y2=3.33
r225 104 107 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=6.48 $Y=3.33
+ $X2=7.44 $Y2=3.33
r226 104 105 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r227 102 105 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=3.33
+ $X2=6.48 $Y2=3.33
r228 101 102 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r229 99 102 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=6 $Y2=3.33
r230 99 142 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=3.6 $Y2=3.33
r231 98 101 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=4.08 $Y=3.33
+ $X2=6 $Y2=3.33
r232 98 99 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r233 96 141 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.875 $Y=3.33
+ $X2=3.71 $Y2=3.33
r234 96 98 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=3.875 $Y=3.33
+ $X2=4.08 $Y2=3.33
r235 95 139 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.64 $Y2=3.33
r236 95 136 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r237 94 95 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r238 92 135 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.895 $Y=3.33
+ $X2=0.73 $Y2=3.33
r239 92 94 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.895 $Y=3.33
+ $X2=1.2 $Y2=3.33
r240 91 138 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.56 $Y=3.33
+ $X2=2.725 $Y2=3.33
r241 91 94 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=2.56 $Y=3.33
+ $X2=1.2 $Y2=3.33
r242 89 136 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r243 88 89 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r244 86 135 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.565 $Y=3.33
+ $X2=0.73 $Y2=3.33
r245 86 88 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.565 $Y=3.33
+ $X2=0.24 $Y2=3.33
r246 84 111 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=8.4 $Y2=3.33
r247 84 105 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=6.48 $Y2=3.33
r248 84 107 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r249 82 110 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=8.435 $Y=3.33
+ $X2=8.4 $Y2=3.33
r250 82 83 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.435 $Y=3.33
+ $X2=8.56 $Y2=3.33
r251 81 114 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=8.685 $Y=3.33
+ $X2=8.88 $Y2=3.33
r252 81 83 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.685 $Y=3.33
+ $X2=8.56 $Y2=3.33
r253 79 107 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=7.535 $Y=3.33
+ $X2=7.44 $Y2=3.33
r254 79 80 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.535 $Y=3.33
+ $X2=7.62 $Y2=3.33
r255 78 110 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=7.705 $Y=3.33
+ $X2=8.4 $Y2=3.33
r256 78 80 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.705 $Y=3.33
+ $X2=7.62 $Y2=3.33
r257 76 101 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=6.095 $Y=3.33
+ $X2=6 $Y2=3.33
r258 76 77 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.095 $Y=3.33
+ $X2=6.22 $Y2=3.33
r259 75 104 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=6.345 $Y=3.33
+ $X2=6.48 $Y2=3.33
r260 75 77 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.345 $Y=3.33
+ $X2=6.22 $Y2=3.33
r261 71 153 3.00555 $w=3.3e-07 $l=1.07912e-07 $layer=LI1_cond $X=14.61 $Y=3.245
+ $X2=14.662 $Y2=3.33
r262 71 73 29.3349 $w=3.28e-07 $l=8.4e-07 $layer=LI1_cond $X=14.61 $Y=3.245
+ $X2=14.61 $Y2=2.405
r263 67 70 29.5187 $w=2.83e-07 $l=7.3e-07 $layer=LI1_cond $X=13.682 $Y=2.085
+ $X2=13.682 $Y2=2.815
r264 65 150 0.432977 $w=2.85e-07 $l=8.5e-08 $layer=LI1_cond $X=13.682 $Y=3.245
+ $X2=13.682 $Y2=3.33
r265 65 70 17.3877 $w=2.83e-07 $l=4.3e-07 $layer=LI1_cond $X=13.682 $Y=3.245
+ $X2=13.682 $Y2=2.815
r266 61 147 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=12.675 $Y=3.245
+ $X2=12.675 $Y2=3.33
r267 61 63 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=12.675 $Y=3.245
+ $X2=12.675 $Y2=2.815
r268 57 144 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=11.205 $Y=3.245
+ $X2=11.205 $Y2=3.33
r269 57 59 20.0525 $w=2.48e-07 $l=4.35e-07 $layer=LI1_cond $X=11.205 $Y=3.245
+ $X2=11.205 $Y2=2.81
r270 53 83 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=8.56 $Y=3.245
+ $X2=8.56 $Y2=3.33
r271 53 55 30.655 $w=2.48e-07 $l=6.65e-07 $layer=LI1_cond $X=8.56 $Y=3.245
+ $X2=8.56 $Y2=2.58
r272 49 80 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.62 $Y=3.245
+ $X2=7.62 $Y2=3.33
r273 49 51 66.2193 $w=1.68e-07 $l=1.015e-06 $layer=LI1_cond $X=7.62 $Y=3.245
+ $X2=7.62 $Y2=2.23
r274 45 77 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.22 $Y=3.245
+ $X2=6.22 $Y2=3.33
r275 45 47 30.194 $w=2.48e-07 $l=6.55e-07 $layer=LI1_cond $X=6.22 $Y=3.245
+ $X2=6.22 $Y2=2.59
r276 41 141 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.71 $Y=3.245
+ $X2=3.71 $Y2=3.33
r277 41 43 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=3.71 $Y=3.245
+ $X2=3.71 $Y2=2.78
r278 40 138 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.89 $Y=3.33
+ $X2=2.725 $Y2=3.33
r279 39 141 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.545 $Y=3.33
+ $X2=3.71 $Y2=3.33
r280 39 40 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=3.545 $Y=3.33
+ $X2=2.89 $Y2=3.33
r281 35 138 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.725 $Y=3.245
+ $X2=2.725 $Y2=3.33
r282 35 37 8.73063 $w=3.28e-07 $l=2.5e-07 $layer=LI1_cond $X=2.725 $Y=3.245
+ $X2=2.725 $Y2=2.995
r283 31 135 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.73 $Y=3.245
+ $X2=0.73 $Y2=3.33
r284 31 33 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=0.73 $Y=3.245
+ $X2=0.73 $Y2=2.78
r285 10 73 300 $w=1.7e-07 $l=6.3559e-07 $layer=licon1_PDIFF $count=2 $X=14.46
+ $Y=1.84 $X2=14.61 $Y2=2.405
r286 9 70 400 $w=1.7e-07 $l=9.4975e-07 $layer=licon1_PDIFF $count=1 $X=13.505
+ $Y=1.96 $X2=13.705 $Y2=2.815
r287 9 67 400 $w=1.7e-07 $l=2.54951e-07 $layer=licon1_PDIFF $count=1 $X=13.505
+ $Y=1.96 $X2=13.705 $Y2=2.085
r288 8 63 600 $w=1.7e-07 $l=3.4187e-07 $layer=licon1_PDIFF $count=1 $X=12.525
+ $Y=2.54 $X2=12.675 $Y2=2.815
r289 7 59 600 $w=1.7e-07 $l=3.36749e-07 $layer=licon1_PDIFF $count=1 $X=11.095
+ $Y=2.54 $X2=11.245 $Y2=2.81
r290 6 55 600 $w=1.7e-07 $l=7.5629e-07 $layer=licon1_PDIFF $count=1 $X=8.37
+ $Y=1.895 $X2=8.52 $Y2=2.58
r291 5 51 300 $w=1.7e-07 $l=3.751e-07 $layer=licon1_PDIFF $count=2 $X=7.285
+ $Y=2.315 $X2=7.62 $Y2=2.23
r292 4 47 600 $w=1.7e-07 $l=3.43875e-07 $layer=licon1_PDIFF $count=1 $X=6.105
+ $Y=2.315 $X2=6.26 $Y2=2.59
r293 3 43 600 $w=1.7e-07 $l=1.01223e-06 $layer=licon1_PDIFF $count=1 $X=3.56
+ $Y=1.84 $X2=3.71 $Y2=2.78
r294 2 37 600 $w=1.7e-07 $l=7.79423e-07 $layer=licon1_PDIFF $count=1 $X=2.5
+ $Y=2.32 $X2=2.725 $Y2=2.995
r295 1 33 600 $w=1.7e-07 $l=5.29717e-07 $layer=licon1_PDIFF $count=1 $X=0.58
+ $Y=2.32 $X2=0.73 $Y2=2.78
.ends

.subckt PM_SKY130_FD_SC_HS__SDFSTP_2%A_290_464# 1 2 3 4 13 19 21 22 24 25 27 32
+ 33 36 43 45 46 47
c130 27 0 4.69178e-20 $X=4.585 $Y=2.325
c131 24 0 4.46515e-20 $X=2.3 $Y=2.49
c132 22 0 1.77325e-19 $X=1.89 $Y=0.995
c133 19 0 8.84878e-21 $X=1.725 $Y=0.58
r134 47 49 5.93683 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=4.75 $Y=2.325
+ $X2=4.75 $Y2=2.495
r135 45 46 8.63679 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=4.667 $Y=1.9
+ $X2=4.667 $Y2=2.07
r136 40 43 7.37564 $w=2.48e-07 $l=1.6e-07 $layer=LI1_cond $X=4.505 $Y=0.72
+ $X2=4.665 $Y2=0.72
r137 36 38 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=3.035 $Y=2.325
+ $X2=3.035 $Y2=2.575
r138 32 47 2.96841 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=4.75 $Y=2.24
+ $X2=4.75 $Y2=2.325
r139 32 46 5.93683 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=4.75 $Y=2.24
+ $X2=4.75 $Y2=2.07
r140 29 40 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.505 $Y=0.845
+ $X2=4.505 $Y2=0.72
r141 29 45 68.8289 $w=1.68e-07 $l=1.055e-06 $layer=LI1_cond $X=4.505 $Y=0.845
+ $X2=4.505 $Y2=1.9
r142 28 36 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.12 $Y=2.325
+ $X2=3.035 $Y2=2.325
r143 27 47 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.585 $Y=2.325
+ $X2=4.75 $Y2=2.325
r144 27 28 95.5775 $w=1.68e-07 $l=1.465e-06 $layer=LI1_cond $X=4.585 $Y=2.325
+ $X2=3.12 $Y2=2.325
r145 26 33 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.385 $Y=2.575
+ $X2=2.3 $Y2=2.575
r146 25 38 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.95 $Y=2.575
+ $X2=3.035 $Y2=2.575
r147 25 26 36.861 $w=1.68e-07 $l=5.65e-07 $layer=LI1_cond $X=2.95 $Y=2.575
+ $X2=2.385 $Y2=2.575
r148 24 33 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=2.3 $Y=2.49 $X2=2.3
+ $Y2=2.575
r149 23 24 91.9893 $w=1.68e-07 $l=1.41e-06 $layer=LI1_cond $X=2.3 $Y=1.08
+ $X2=2.3 $Y2=2.49
r150 21 23 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.215 $Y=0.995
+ $X2=2.3 $Y2=1.08
r151 21 22 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=2.215 $Y=0.995
+ $X2=1.89 $Y2=0.995
r152 17 22 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.725 $Y=0.91
+ $X2=1.89 $Y2=0.995
r153 17 19 11.5244 $w=3.28e-07 $l=3.3e-07 $layer=LI1_cond $X=1.725 $Y=0.91
+ $X2=1.725 $Y2=0.58
r154 13 33 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=2.3 $Y=2.785
+ $X2=2.3 $Y2=2.575
r155 13 15 24.2013 $w=2.48e-07 $l=5.25e-07 $layer=LI1_cond $X=2.215 $Y=2.785
+ $X2=1.69 $Y2=2.785
r156 4 49 600 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_PDIFF $count=1 $X=4.605
+ $Y=2.285 $X2=4.75 $Y2=2.495
r157 3 15 600 $w=1.7e-07 $l=5.31625e-07 $layer=licon1_PDIFF $count=1 $X=1.45
+ $Y=2.32 $X2=1.69 $Y2=2.745
r158 2 43 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=4.525
+ $Y=0.405 $X2=4.665 $Y2=0.68
r159 1 19 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.585
+ $Y=0.37 $X2=1.725 $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_HS__SDFSTP_2%A_1584_379# 1 2 9 11 15 18 19
c35 19 0 1.38803e-19 $X=8.68 $Y=2.06
r36 19 21 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=8.68 $Y=2.06 $X2=8.68
+ $Y2=2.15
r37 13 15 4.1907 $w=3.28e-07 $l=1.2e-07 $layer=LI1_cond $X=9.665 $Y=2.145
+ $X2=9.665 $Y2=2.265
r38 12 19 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.765 $Y=2.06
+ $X2=8.68 $Y2=2.06
r39 11 13 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=9.5 $Y=2.06
+ $X2=9.665 $Y2=2.145
r40 11 12 47.9519 $w=1.68e-07 $l=7.35e-07 $layer=LI1_cond $X=9.5 $Y=2.06
+ $X2=8.765 $Y2=2.06
r41 10 18 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.235 $Y=2.15
+ $X2=8.07 $Y2=2.15
r42 9 21 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.595 $Y=2.15
+ $X2=8.68 $Y2=2.15
r43 9 10 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=8.595 $Y=2.15
+ $X2=8.235 $Y2=2.15
r44 2 15 300 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=2 $X=9.515
+ $Y=2.12 $X2=9.665 $Y2=2.265
r45 1 18 300 $w=1.7e-07 $l=4.03082e-07 $layer=licon1_PDIFF $count=2 $X=7.92
+ $Y=1.895 $X2=8.07 $Y2=2.23
.ends

.subckt PM_SKY130_FD_SC_HS__SDFSTP_2%Q 1 2 9 13 17 19 20 21 22
c41 20 0 5.67555e-20 $X=14.465 $Y=1.49
r42 28 31 0.873063 $w=3.28e-07 $l=2.5e-08 $layer=LI1_cond $X=14.135 $Y=1.985
+ $X2=14.16 $Y2=1.985
r43 25 31 13.2706 $w=3.28e-07 $l=3.8e-07 $layer=LI1_cond $X=14.54 $Y=1.985
+ $X2=14.16 $Y2=1.985
r44 22 25 3.49225 $w=3.28e-07 $l=1e-07 $layer=LI1_cond $X=14.64 $Y=1.985
+ $X2=14.54 $Y2=1.985
r45 21 25 4.15415 $w=4.28e-07 $l=1.55e-07 $layer=LI1_cond $X=14.54 $Y=1.665
+ $X2=14.54 $Y2=1.82
r46 20 21 4.69018 $w=4.28e-07 $l=1.75e-07 $layer=LI1_cond $X=14.54 $Y=1.49
+ $X2=14.54 $Y2=1.665
r47 19 20 8.9189 $w=4.28e-07 $l=1.7e-07 $layer=LI1_cond $X=14.465 $Y=1.32
+ $X2=14.465 $Y2=1.49
r48 17 19 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=14.26 $Y=1.15
+ $X2=14.26 $Y2=1.32
r49 11 28 1.70047 $w=2.8e-07 $l=1.65e-07 $layer=LI1_cond $X=14.135 $Y=2.15
+ $X2=14.135 $Y2=1.985
r50 11 13 10.7013 $w=2.78e-07 $l=2.6e-07 $layer=LI1_cond $X=14.135 $Y=2.15
+ $X2=14.135 $Y2=2.41
r51 7 17 8.88861 $w=3.53e-07 $l=1.77e-07 $layer=LI1_cond $X=14.167 $Y=0.973
+ $X2=14.167 $Y2=1.15
r52 7 9 14.2189 $w=3.53e-07 $l=4.38e-07 $layer=LI1_cond $X=14.167 $Y=0.973
+ $X2=14.167 $Y2=0.535
r53 2 31 600 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=14.01
+ $Y=1.84 $X2=14.16 $Y2=1.985
r54 2 13 300 $w=1.7e-07 $l=6.40625e-07 $layer=licon1_PDIFF $count=2 $X=14.01
+ $Y=1.84 $X2=14.16 $Y2=2.41
r55 1 9 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=14.015
+ $Y=0.39 $X2=14.155 $Y2=0.535
.ends

.subckt PM_SKY130_FD_SC_HS__SDFSTP_2%VGND 1 2 3 4 5 6 7 8 9 30 34 36 40 44 48 52
+ 54 56 58 59 65 67 72 87 94 107 112 118 121 124 127 130 135 141 143 147
c162 147 0 2.52187e-20 $X=14.64 $Y=0
r163 146 147 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=14.64 $Y=0
+ $X2=14.64 $Y2=0
r164 143 144 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.68 $Y=0
+ $X2=13.68 $Y2=0
r165 139 141 9.39905 $w=6.83e-07 $l=9e-08 $layer=LI1_cond $X=12.24 $Y=0.257
+ $X2=12.33 $Y2=0.257
r166 139 140 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.24 $Y=0
+ $X2=12.24 $Y2=0
r167 137 139 1.30957 $w=6.83e-07 $l=7.5e-08 $layer=LI1_cond $X=12.165 $Y=0.257
+ $X2=12.24 $Y2=0.257
r168 134 140 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.76 $Y=0
+ $X2=12.24 $Y2=0
r169 133 137 7.0717 $w=6.83e-07 $l=4.05e-07 $layer=LI1_cond $X=11.76 $Y=0.257
+ $X2=12.165 $Y2=0.257
r170 133 135 9.92288 $w=6.83e-07 $l=1.2e-07 $layer=LI1_cond $X=11.76 $Y=0.257
+ $X2=11.64 $Y2=0.257
r171 133 134 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.76 $Y=0
+ $X2=11.76 $Y2=0
r172 130 131 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=0
+ $X2=8.88 $Y2=0
r173 127 128 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=0
+ $X2=7.92 $Y2=0
r174 124 125 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r175 122 125 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=0
+ $X2=3.6 $Y2=0
r176 121 122 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0
+ $X2=2.64 $Y2=0
r177 118 119 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0
+ $X2=0.72 $Y2=0
r178 116 147 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=14.16 $Y=0
+ $X2=14.64 $Y2=0
r179 116 144 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=14.16 $Y=0
+ $X2=13.68 $Y2=0
r180 115 116 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=14.16 $Y=0
+ $X2=14.16 $Y2=0
r181 113 143 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=13.805 $Y=0
+ $X2=13.68 $Y2=0
r182 113 115 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=13.805 $Y=0
+ $X2=14.16 $Y2=0
r183 112 146 4.01252 $w=1.7e-07 $l=1.82e-07 $layer=LI1_cond $X=14.515 $Y=0
+ $X2=14.697 $Y2=0
r184 112 115 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=14.515 $Y=0
+ $X2=14.16 $Y2=0
r185 111 144 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=13.2 $Y=0
+ $X2=13.68 $Y2=0
r186 111 140 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=13.2 $Y=0
+ $X2=12.24 $Y2=0
r187 110 141 56.7594 $w=1.68e-07 $l=8.7e-07 $layer=LI1_cond $X=13.2 $Y=0
+ $X2=12.33 $Y2=0
r188 110 111 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=13.2 $Y=0
+ $X2=13.2 $Y2=0
r189 107 143 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=13.555 $Y=0
+ $X2=13.68 $Y2=0
r190 107 110 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=13.555 $Y=0
+ $X2=13.2 $Y2=0
r191 106 134 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.28 $Y=0
+ $X2=11.76 $Y2=0
r192 105 135 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=11.28 $Y=0
+ $X2=11.64 $Y2=0
r193 105 106 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=11.28 $Y=0
+ $X2=11.28 $Y2=0
r194 103 106 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=9.36 $Y=0
+ $X2=11.28 $Y2=0
r195 103 131 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.36 $Y=0
+ $X2=8.88 $Y2=0
r196 102 105 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=9.36 $Y=0
+ $X2=11.28 $Y2=0
r197 102 103 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=9.36 $Y=0
+ $X2=9.36 $Y2=0
r198 100 130 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.02 $Y=0
+ $X2=8.855 $Y2=0
r199 100 102 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=9.02 $Y=0
+ $X2=9.36 $Y2=0
r200 98 131 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=0 $X2=8.88
+ $Y2=0
r201 98 128 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=0 $X2=7.92
+ $Y2=0
r202 97 98 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r203 95 127 11.2921 $w=1.7e-07 $l=2.5e-07 $layer=LI1_cond $X=8.01 $Y=0 $X2=7.76
+ $Y2=0
r204 95 97 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=8.01 $Y=0 $X2=8.4
+ $Y2=0
r205 94 130 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.69 $Y=0
+ $X2=8.855 $Y2=0
r206 94 97 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=8.69 $Y=0 $X2=8.4
+ $Y2=0
r207 89 92 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=6.48 $Y=0 $X2=7.44
+ $Y2=0
r208 89 90 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6.48 $Y=0 $X2=6.48
+ $Y2=0
r209 87 127 11.2921 $w=1.7e-07 $l=2.5e-07 $layer=LI1_cond $X=7.51 $Y=0 $X2=7.76
+ $Y2=0
r210 87 92 4.56684 $w=1.68e-07 $l=7e-08 $layer=LI1_cond $X=7.51 $Y=0 $X2=7.44
+ $Y2=0
r211 86 90 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=0 $X2=6.48
+ $Y2=0
r212 85 86 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6 $Y=0 $X2=6
+ $Y2=0
r213 83 86 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=4.08 $Y=0 $X2=6
+ $Y2=0
r214 83 125 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=3.6
+ $Y2=0
r215 82 85 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=4.08 $Y=0 $X2=6
+ $Y2=0
r216 82 83 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.08 $Y=0
+ $X2=4.08 $Y2=0
r217 80 124 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.85 $Y=0
+ $X2=3.685 $Y2=0
r218 80 82 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=3.85 $Y=0 $X2=4.08
+ $Y2=0
r219 79 122 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0
+ $X2=2.64 $Y2=0
r220 78 79 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r221 76 79 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r222 76 119 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r223 75 78 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r224 75 76 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r225 73 118 10.6558 $w=1.7e-07 $l=2.28e-07 $layer=LI1_cond $X=1.07 $Y=0
+ $X2=0.842 $Y2=0
r226 73 75 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=1.07 $Y=0 $X2=1.2
+ $Y2=0
r227 72 121 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.46 $Y=0
+ $X2=2.625 $Y2=0
r228 72 78 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=2.46 $Y=0 $X2=2.16
+ $Y2=0
r229 70 119 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0
+ $X2=0.72 $Y2=0
r230 69 70 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r231 67 118 10.6558 $w=1.7e-07 $l=2.27e-07 $layer=LI1_cond $X=0.615 $Y=0
+ $X2=0.842 $Y2=0
r232 67 69 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=0.615 $Y=0
+ $X2=0.24 $Y2=0
r233 65 128 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=0
+ $X2=7.92 $Y2=0
r234 65 90 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=7.44 $Y=0 $X2=6.48
+ $Y2=0
r235 65 92 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=7.44 $Y=0 $X2=7.44
+ $Y2=0
r236 61 89 1.30481 $w=1.68e-07 $l=2e-08 $layer=LI1_cond $X=6.46 $Y=0 $X2=6.48
+ $Y2=0
r237 59 85 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=6.13 $Y=0 $X2=6
+ $Y2=0
r238 58 63 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=6.295 $Y=0
+ $X2=6.295 $Y2=0.275
r239 58 61 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.295 $Y=0 $X2=6.46
+ $Y2=0
r240 58 59 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.295 $Y=0 $X2=6.13
+ $Y2=0
r241 54 146 3.13065 $w=2.5e-07 $l=1.09864e-07 $layer=LI1_cond $X=14.64 $Y=0.085
+ $X2=14.697 $Y2=0
r242 54 56 20.283 $w=2.48e-07 $l=4.4e-07 $layer=LI1_cond $X=14.64 $Y=0.085
+ $X2=14.64 $Y2=0.525
r243 50 143 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=13.68 $Y=0.085
+ $X2=13.68 $Y2=0
r244 50 52 20.744 $w=2.48e-07 $l=4.5e-07 $layer=LI1_cond $X=13.68 $Y=0.085
+ $X2=13.68 $Y2=0.535
r245 46 130 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.855 $Y=0.085
+ $X2=8.855 $Y2=0
r246 46 48 15.5405 $w=3.28e-07 $l=4.45e-07 $layer=LI1_cond $X=8.855 $Y=0.085
+ $X2=8.855 $Y2=0.53
r247 42 127 2.07448 $w=5e-07 $l=8.5e-08 $layer=LI1_cond $X=7.76 $Y=0.085
+ $X2=7.76 $Y2=0
r248 42 44 10.2863 $w=4.98e-07 $l=4.3e-07 $layer=LI1_cond $X=7.76 $Y=0.085
+ $X2=7.76 $Y2=0.515
r249 38 124 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.685 $Y=0.085
+ $X2=3.685 $Y2=0
r250 38 40 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=3.685 $Y=0.085
+ $X2=3.685 $Y2=0.515
r251 37 121 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.79 $Y=0
+ $X2=2.625 $Y2=0
r252 36 124 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.52 $Y=0
+ $X2=3.685 $Y2=0
r253 36 37 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=3.52 $Y=0 $X2=2.79
+ $Y2=0
r254 32 121 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.625 $Y=0.085
+ $X2=2.625 $Y2=0
r255 32 34 16.0644 $w=3.28e-07 $l=4.6e-07 $layer=LI1_cond $X=2.625 $Y=0.085
+ $X2=2.625 $Y2=0.545
r256 28 118 1.82608 $w=4.55e-07 $l=8.5e-08 $layer=LI1_cond $X=0.842 $Y=0.085
+ $X2=0.842 $Y2=0
r257 28 30 11.3036 $w=4.53e-07 $l=4.3e-07 $layer=LI1_cond $X=0.842 $Y=0.085
+ $X2=0.842 $Y2=0.515
r258 9 56 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=14.445
+ $Y=0.39 $X2=14.6 $Y2=0.525
r259 8 52 91 $w=1.7e-07 $l=2.51496e-07 $layer=licon1_NDIFF $count=2 $X=13.49
+ $Y=0.49 $X2=13.72 $Y2=0.535
r260 7 137 91 $w=1.7e-07 $l=5.67891e-07 $layer=licon1_NDIFF $count=2 $X=11.665
+ $Y=0.37 $X2=12.165 $Y2=0.515
r261 6 48 182 $w=1.7e-07 $l=2.89137e-07 $layer=licon1_NDIFF $count=1 $X=8.635
+ $Y=0.37 $X2=8.855 $Y2=0.53
r262 5 44 182 $w=1.7e-07 $l=2.88531e-07 $layer=licon1_NDIFF $count=1 $X=7.535
+ $Y=0.37 $X2=7.76 $Y2=0.515
r263 4 63 182 $w=1.7e-07 $l=2.77489e-07 $layer=licon1_NDIFF $count=1 $X=6.075
+ $Y=0.405 $X2=6.295 $Y2=0.275
r264 3 40 91 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=2 $X=3.475
+ $Y=0.37 $X2=3.685 $Y2=0.515
r265 2 34 182 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_NDIFF $count=1 $X=2.485
+ $Y=0.37 $X2=2.625 $Y2=0.545
r266 1 30 182 $w=1.7e-07 $l=3.34739e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.37 $X2=0.84 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__SDFSTP_2%A_1641_74# 1 2 9 11 12 14
c42 12 0 1.09822e-19 $X=8.51 $Y=0.97
c43 11 0 3.01101e-20 $X=9.75 $Y=0.97
r44 14 16 5.5876 $w=3.28e-07 $l=1.6e-07 $layer=LI1_cond $X=9.915 $Y=0.81
+ $X2=9.915 $Y2=0.97
r45 11 16 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.75 $Y=0.97
+ $X2=9.915 $Y2=0.97
r46 11 12 80.8984 $w=1.68e-07 $l=1.24e-06 $layer=LI1_cond $X=9.75 $Y=0.97
+ $X2=8.51 $Y2=0.97
r47 7 12 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=8.345 $Y=0.885
+ $X2=8.51 $Y2=0.97
r48 7 9 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=8.345 $Y=0.885
+ $X2=8.345 $Y2=0.515
r49 2 14 182 $w=1.7e-07 $l=5.05173e-07 $layer=licon1_NDIFF $count=1 $X=9.775
+ $Y=0.37 $X2=9.915 $Y2=0.81
r50 1 9 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=8.205
+ $Y=0.37 $X2=8.345 $Y2=0.515
.ends

