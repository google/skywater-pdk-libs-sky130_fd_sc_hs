* File: sky130_fd_sc_hs__o32ai_1.spice
* Created: Thu Aug 27 21:03:42 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hs__o32ai_1.pex.spice"
.subckt sky130_fd_sc_hs__o32ai_1  VNB VPB B1 B2 A3 A2 A1 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A1	A1
* A2	A2
* A3	A3
* B2	B2
* B1	B1
* VPB	VPB
* VNB	VNB
MM1008 N_Y_M1008_d N_B1_M1008_g N_A_27_74#_M1008_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.21645 AS=0.2109 PD=1.325 PS=2.05 NRD=30 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75002.5 A=0.111 P=1.78 MULT=1
MM1006 N_A_27_74#_M1006_d N_B2_M1006_g N_Y_M1008_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.1295 AS=0.21645 PD=1.09 PS=1.325 NRD=11.34 NRS=19.452 M=1 R=4.93333
+ SA=75000.9 SB=75001.7 A=0.111 P=1.78 MULT=1
MM1003 N_VGND_M1003_d N_A3_M1003_g N_A_27_74#_M1006_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.1665 AS=0.1295 PD=1.19 PS=1.09 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75001.4
+ SB=75001.2 A=0.111 P=1.78 MULT=1
MM1007 N_A_27_74#_M1007_d N_A2_M1007_g N_VGND_M1003_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1665 PD=1.02 PS=1.19 NRD=0 NRS=16.212 M=1 R=4.93333 SA=75002
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1004 N_VGND_M1004_d N_A1_M1004_g N_A_27_74#_M1007_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.1036 PD=2.05 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75002.5
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1000 A_128_368# N_B1_M1000_g N_VPWR_M1000_s VPB PSHORT L=0.15 W=1.12 AD=0.1512
+ AS=0.3752 PD=1.39 PS=2.91 NRD=14.0658 NRS=8.7862 M=1 R=7.46667 SA=75000.3
+ SB=75002.4 A=0.168 P=2.54 MULT=1
MM1005 N_Y_M1005_d N_B2_M1005_g A_128_368# VPB PSHORT L=0.15 W=1.12 AD=0.28
+ AS=0.1512 PD=1.62 PS=1.39 NRD=1.7533 NRS=14.0658 M=1 R=7.46667 SA=75000.7
+ SB=75002 A=0.168 P=2.54 MULT=1
MM1001 A_342_368# N_A3_M1001_g N_Y_M1005_d VPB PSHORT L=0.15 W=1.12 AD=0.2352
+ AS=0.28 PD=1.54 PS=1.62 NRD=27.2451 NRS=36.9178 M=1 R=7.46667 SA=75001.3
+ SB=75001.4 A=0.168 P=2.54 MULT=1
MM1009 A_456_368# N_A2_M1009_g A_342_368# VPB PSHORT L=0.15 W=1.12 AD=0.2352
+ AS=0.2352 PD=1.54 PS=1.54 NRD=27.2451 NRS=27.2451 M=1 R=7.46667 SA=75001.9
+ SB=75000.8 A=0.168 P=2.54 MULT=1
MM1002 N_VPWR_M1002_d N_A1_M1002_g A_456_368# VPB PSHORT L=0.15 W=1.12 AD=0.3304
+ AS=0.2352 PD=2.83 PS=1.54 NRD=1.7533 NRS=27.2451 M=1 R=7.46667 SA=75002.5
+ SB=75000.2 A=0.168 P=2.54 MULT=1
DX10_noxref VNB VPB NWDIODE A=6.9564 P=11.2
*
.include "sky130_fd_sc_hs__o32ai_1.pxi.spice"
*
.ends
*
*
