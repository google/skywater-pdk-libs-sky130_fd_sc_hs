* File: sky130_fd_sc_hs__clkbuf_16.pex.spice
* Created: Thu Aug 27 20:35:22 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HS__CLKBUF_16%A 3 5 7 10 12 14 17 19 21 24 26 28 29 30
+ 31 32 49
c88 26 0 1.47033e-19 $X=1.86 $Y=1.765
r89 49 50 7.16487 $w=3.7e-07 $l=5.5e-08 $layer=POLY_cond $X=1.805 $Y=1.557
+ $X2=1.86 $Y2=1.557
r90 47 49 26.0541 $w=3.7e-07 $l=2e-07 $layer=POLY_cond $X=1.605 $Y=1.557
+ $X2=1.805 $Y2=1.557
r91 47 48 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.605
+ $Y=1.515 $X2=1.605 $Y2=1.515
r92 45 47 25.4027 $w=3.7e-07 $l=1.95e-07 $layer=POLY_cond $X=1.41 $Y=1.557
+ $X2=1.605 $Y2=1.557
r93 44 45 4.55946 $w=3.7e-07 $l=3.5e-08 $layer=POLY_cond $X=1.375 $Y=1.557
+ $X2=1.41 $Y2=1.557
r94 43 44 54.0622 $w=3.7e-07 $l=4.15e-07 $layer=POLY_cond $X=0.96 $Y=1.557
+ $X2=1.375 $Y2=1.557
r95 42 43 4.55946 $w=3.7e-07 $l=3.5e-08 $layer=POLY_cond $X=0.925 $Y=1.557
+ $X2=0.96 $Y2=1.557
r96 40 42 44.2919 $w=3.7e-07 $l=3.4e-07 $layer=POLY_cond $X=0.585 $Y=1.557
+ $X2=0.925 $Y2=1.557
r97 40 41 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.585
+ $Y=1.515 $X2=0.585 $Y2=1.515
r98 38 40 9.77027 $w=3.7e-07 $l=7.5e-08 $layer=POLY_cond $X=0.51 $Y=1.557
+ $X2=0.585 $Y2=1.557
r99 37 38 1.95405 $w=3.7e-07 $l=1.5e-08 $layer=POLY_cond $X=0.495 $Y=1.557
+ $X2=0.51 $Y2=1.557
r100 32 48 2.01008 $w=4.28e-07 $l=7.5e-08 $layer=LI1_cond $X=1.68 $Y=1.565
+ $X2=1.605 $Y2=1.565
r101 31 48 10.8544 $w=4.28e-07 $l=4.05e-07 $layer=LI1_cond $X=1.2 $Y=1.565
+ $X2=1.605 $Y2=1.565
r102 30 31 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=0.72 $Y=1.565
+ $X2=1.2 $Y2=1.565
r103 30 41 3.61813 $w=4.28e-07 $l=1.35e-07 $layer=LI1_cond $X=0.72 $Y=1.565
+ $X2=0.585 $Y2=1.565
r104 29 41 9.24634 $w=4.28e-07 $l=3.45e-07 $layer=LI1_cond $X=0.24 $Y=1.565
+ $X2=0.585 $Y2=1.565
r105 26 50 23.9667 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=1.86 $Y=1.765
+ $X2=1.86 $Y2=1.557
r106 26 28 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.86 $Y=1.765
+ $X2=1.86 $Y2=2.4
r107 22 49 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.805 $Y=1.35
+ $X2=1.805 $Y2=1.557
r108 22 24 394.83 $w=1.5e-07 $l=7.7e-07 $layer=POLY_cond $X=1.805 $Y=1.35
+ $X2=1.805 $Y2=0.58
r109 19 45 23.9667 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=1.41 $Y=1.765
+ $X2=1.41 $Y2=1.557
r110 19 21 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.41 $Y=1.765
+ $X2=1.41 $Y2=2.4
r111 15 44 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.375 $Y=1.35
+ $X2=1.375 $Y2=1.557
r112 15 17 394.83 $w=1.5e-07 $l=7.7e-07 $layer=POLY_cond $X=1.375 $Y=1.35
+ $X2=1.375 $Y2=0.58
r113 12 43 23.9667 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=0.96 $Y=1.765
+ $X2=0.96 $Y2=1.557
r114 12 14 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.96 $Y=1.765
+ $X2=0.96 $Y2=2.4
r115 8 42 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.925 $Y=1.35
+ $X2=0.925 $Y2=1.557
r116 8 10 394.83 $w=1.5e-07 $l=7.7e-07 $layer=POLY_cond $X=0.925 $Y=1.35
+ $X2=0.925 $Y2=0.58
r117 5 38 23.9667 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=0.51 $Y=1.765
+ $X2=0.51 $Y2=1.557
r118 5 7 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.51 $Y=1.765
+ $X2=0.51 $Y2=2.4
r119 1 37 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.495 $Y=1.35
+ $X2=0.495 $Y2=1.557
r120 1 3 394.83 $w=1.5e-07 $l=7.7e-07 $layer=POLY_cond $X=0.495 $Y=1.35
+ $X2=0.495 $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_HS__CLKBUF_16%A_114_74# 1 2 3 4 15 18 19 21 24 27 28 30
+ 33 36 37 39 42 45 46 48 51 54 55 57 60 63 64 66 69 72 73 75 78 81 82 84 87 90
+ 91 93 96 99 100 102 104 107 109 111 114 117 118 120 122 123 125 128 131 132
+ 134 137 140 141 143 146 149 150 152 155 159 161 163 165 166 167 171 175 177
+ 179 180 183 186 194 197 200 203 206 209 211 212 267
c470 267 0 1.81624e-20 $X=9.105 $Y=1.355
c471 132 0 1.75614e-19 $X=8.17 $Y=1.765
r472 266 267 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=9.09 $Y=1.355
+ $X2=9.105 $Y2=1.355
r473 265 266 72.5674 $w=3.3e-07 $l=4.15e-07 $layer=POLY_cond $X=8.675 $Y=1.355
+ $X2=9.09 $Y2=1.355
r474 264 265 6.12014 $w=3.3e-07 $l=3.5e-08 $layer=POLY_cond $X=8.64 $Y=1.355
+ $X2=8.675 $Y2=1.355
r475 262 264 43.7153 $w=3.3e-07 $l=2.5e-07 $layer=POLY_cond $X=8.39 $Y=1.355
+ $X2=8.64 $Y2=1.355
r476 260 262 37.5952 $w=3.3e-07 $l=2.15e-07 $layer=POLY_cond $X=8.175 $Y=1.355
+ $X2=8.39 $Y2=1.355
r477 259 260 0.874306 $w=3.3e-07 $l=5e-09 $layer=POLY_cond $X=8.17 $Y=1.355
+ $X2=8.175 $Y2=1.355
r478 258 259 74.316 $w=3.3e-07 $l=4.25e-07 $layer=POLY_cond $X=7.745 $Y=1.355
+ $X2=8.17 $Y2=1.355
r479 257 258 4.37153 $w=3.3e-07 $l=2.5e-08 $layer=POLY_cond $X=7.72 $Y=1.355
+ $X2=7.745 $Y2=1.355
r480 255 257 45.4639 $w=3.3e-07 $l=2.6e-07 $layer=POLY_cond $X=7.46 $Y=1.355
+ $X2=7.72 $Y2=1.355
r481 253 255 33.2236 $w=3.3e-07 $l=1.9e-07 $layer=POLY_cond $X=7.27 $Y=1.355
+ $X2=7.46 $Y2=1.355
r482 252 253 4.37153 $w=3.3e-07 $l=2.5e-08 $layer=POLY_cond $X=7.245 $Y=1.355
+ $X2=7.27 $Y2=1.355
r483 251 252 74.316 $w=3.3e-07 $l=4.25e-07 $layer=POLY_cond $X=6.82 $Y=1.355
+ $X2=7.245 $Y2=1.355
r484 250 251 0.874306 $w=3.3e-07 $l=5e-09 $layer=POLY_cond $X=6.815 $Y=1.355
+ $X2=6.82 $Y2=1.355
r485 248 250 49.8355 $w=3.3e-07 $l=2.85e-07 $layer=POLY_cond $X=6.53 $Y=1.355
+ $X2=6.815 $Y2=1.355
r486 246 248 27.9778 $w=3.3e-07 $l=1.6e-07 $layer=POLY_cond $X=6.37 $Y=1.355
+ $X2=6.53 $Y2=1.355
r487 245 246 9.61737 $w=3.3e-07 $l=5.5e-08 $layer=POLY_cond $X=6.315 $Y=1.355
+ $X2=6.37 $Y2=1.355
r488 244 245 69.0702 $w=3.3e-07 $l=3.95e-07 $layer=POLY_cond $X=5.92 $Y=1.355
+ $X2=6.315 $Y2=1.355
r489 243 244 6.12014 $w=3.3e-07 $l=3.5e-08 $layer=POLY_cond $X=5.885 $Y=1.355
+ $X2=5.92 $Y2=1.355
r490 241 243 51.5841 $w=3.3e-07 $l=2.95e-07 $layer=POLY_cond $X=5.59 $Y=1.355
+ $X2=5.885 $Y2=1.355
r491 239 241 20.9834 $w=3.3e-07 $l=1.2e-07 $layer=POLY_cond $X=5.47 $Y=1.355
+ $X2=5.59 $Y2=1.355
r492 238 239 14.8632 $w=3.3e-07 $l=8.5e-08 $layer=POLY_cond $X=5.385 $Y=1.355
+ $X2=5.47 $Y2=1.355
r493 237 238 63.8244 $w=3.3e-07 $l=3.65e-07 $layer=POLY_cond $X=5.02 $Y=1.355
+ $X2=5.385 $Y2=1.355
r494 236 237 11.366 $w=3.3e-07 $l=6.5e-08 $layer=POLY_cond $X=4.955 $Y=1.355
+ $X2=5.02 $Y2=1.355
r495 234 236 48.9612 $w=3.3e-07 $l=2.8e-07 $layer=POLY_cond $X=4.675 $Y=1.355
+ $X2=4.955 $Y2=1.355
r496 232 234 18.3604 $w=3.3e-07 $l=1.05e-07 $layer=POLY_cond $X=4.57 $Y=1.355
+ $X2=4.675 $Y2=1.355
r497 231 232 20.109 $w=3.3e-07 $l=1.15e-07 $layer=POLY_cond $X=4.455 $Y=1.355
+ $X2=4.57 $Y2=1.355
r498 230 231 58.5785 $w=3.3e-07 $l=3.35e-07 $layer=POLY_cond $X=4.12 $Y=1.355
+ $X2=4.455 $Y2=1.355
r499 229 230 16.6118 $w=3.3e-07 $l=9.5e-08 $layer=POLY_cond $X=4.025 $Y=1.355
+ $X2=4.12 $Y2=1.355
r500 227 229 33.2236 $w=3.3e-07 $l=1.9e-07 $layer=POLY_cond $X=3.835 $Y=1.355
+ $X2=4.025 $Y2=1.355
r501 225 227 28.8521 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.67 $Y=1.355
+ $X2=3.835 $Y2=1.355
r502 224 225 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=3.595 $Y=1.355
+ $X2=3.67 $Y2=1.355
r503 223 224 65.573 $w=3.3e-07 $l=3.75e-07 $layer=POLY_cond $X=3.22 $Y=1.355
+ $X2=3.595 $Y2=1.355
r504 222 223 9.61737 $w=3.3e-07 $l=5.5e-08 $layer=POLY_cond $X=3.165 $Y=1.355
+ $X2=3.22 $Y2=1.355
r505 220 222 33.2236 $w=3.3e-07 $l=1.9e-07 $layer=POLY_cond $X=2.975 $Y=1.355
+ $X2=3.165 $Y2=1.355
r506 218 220 35.8466 $w=3.3e-07 $l=2.05e-07 $layer=POLY_cond $X=2.77 $Y=1.355
+ $X2=2.975 $Y2=1.355
r507 217 218 6.12014 $w=3.3e-07 $l=3.5e-08 $layer=POLY_cond $X=2.735 $Y=1.355
+ $X2=2.77 $Y2=1.355
r508 216 217 72.5674 $w=3.3e-07 $l=4.15e-07 $layer=POLY_cond $X=2.32 $Y=1.355
+ $X2=2.735 $Y2=1.355
r509 214 216 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=2.305 $Y=1.355
+ $X2=2.32 $Y2=1.355
r510 212 262 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.39
+ $Y=1.355 $X2=8.39 $Y2=1.355
r511 211 212 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.39 $Y=1.295
+ $X2=8.39 $Y2=1.295
r512 209 255 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.46
+ $Y=1.355 $X2=7.46 $Y2=1.355
r513 208 211 0.596692 $w=2.3e-07 $l=9.3e-07 $layer=MET1_cond $X=7.46 $Y=1.295
+ $X2=8.39 $Y2=1.295
r514 208 209 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.46 $Y=1.295
+ $X2=7.46 $Y2=1.295
r515 206 248 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.53
+ $Y=1.355 $X2=6.53 $Y2=1.355
r516 205 208 0.596692 $w=2.3e-07 $l=9.3e-07 $layer=MET1_cond $X=6.53 $Y=1.295
+ $X2=7.46 $Y2=1.295
r517 205 206 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.53 $Y=1.295
+ $X2=6.53 $Y2=1.295
r518 203 241 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.59
+ $Y=1.355 $X2=5.59 $Y2=1.355
r519 202 205 0.603108 $w=2.3e-07 $l=9.4e-07 $layer=MET1_cond $X=5.59 $Y=1.295
+ $X2=6.53 $Y2=1.295
r520 202 203 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.59 $Y=1.295
+ $X2=5.59 $Y2=1.295
r521 200 234 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.675
+ $Y=1.355 $X2=4.675 $Y2=1.355
r522 199 202 0.587068 $w=2.3e-07 $l=9.15e-07 $layer=MET1_cond $X=4.675 $Y=1.295
+ $X2=5.59 $Y2=1.295
r523 199 200 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.675 $Y=1.295
+ $X2=4.675 $Y2=1.295
r524 197 227 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.835
+ $Y=1.355 $X2=3.835 $Y2=1.355
r525 196 199 0.538948 $w=2.3e-07 $l=8.4e-07 $layer=MET1_cond $X=3.835 $Y=1.295
+ $X2=4.675 $Y2=1.295
r526 196 197 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.835 $Y=1.295
+ $X2=3.835 $Y2=1.295
r527 194 220 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.975
+ $Y=1.355 $X2=2.975 $Y2=1.355
r528 193 196 0.55178 $w=2.3e-07 $l=8.6e-07 $layer=MET1_cond $X=2.975 $Y=1.295
+ $X2=3.835 $Y2=1.295
r529 193 194 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.975 $Y=1.295
+ $X2=2.975 $Y2=1.295
r530 190 290 13.3619 $w=2.1e-07 $l=2.3e-07 $layer=LI1_cond $X=2.087 $Y=1.295
+ $X2=2.087 $Y2=1.065
r531 189 193 0.564612 $w=2.3e-07 $l=8.8e-07 $layer=MET1_cond $X=2.095 $Y=1.295
+ $X2=2.975 $Y2=1.295
r532 189 190 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.095 $Y=1.295
+ $X2=2.095 $Y2=1.295
r533 185 186 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=1.635 $Y=2.035
+ $X2=2.05 $Y2=2.035
r534 180 186 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.05 $Y=1.95
+ $X2=2.05 $Y2=2.035
r535 179 190 7.15932 $w=2.1e-07 $l=1.32212e-07 $layer=LI1_cond $X=2.05 $Y=1.41
+ $X2=2.087 $Y2=1.295
r536 179 180 35.2299 $w=1.68e-07 $l=5.4e-07 $layer=LI1_cond $X=2.05 $Y=1.41
+ $X2=2.05 $Y2=1.95
r537 178 183 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.675 $Y=1.065
+ $X2=1.55 $Y2=1.065
r538 177 290 1.9771 $w=1.7e-07 $l=1.22e-07 $layer=LI1_cond $X=1.965 $Y=1.065
+ $X2=2.087 $Y2=1.065
r539 177 178 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=1.965 $Y=1.065
+ $X2=1.675 $Y2=1.065
r540 175 185 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=1.635 $Y=2.815
+ $X2=1.635 $Y2=2.12
r541 169 183 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.55 $Y=0.98
+ $X2=1.55 $Y2=1.065
r542 169 171 18.4391 $w=2.48e-07 $l=4e-07 $layer=LI1_cond $X=1.55 $Y=0.98
+ $X2=1.55 $Y2=0.58
r543 168 182 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.9 $Y=2.035
+ $X2=0.735 $Y2=2.035
r544 167 185 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=1.47 $Y=2.035
+ $X2=1.635 $Y2=2.035
r545 167 168 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=1.47 $Y=2.035
+ $X2=0.9 $Y2=2.035
r546 165 183 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.425 $Y=1.065
+ $X2=1.55 $Y2=1.065
r547 165 166 41.1016 $w=1.68e-07 $l=6.3e-07 $layer=LI1_cond $X=1.425 $Y=1.065
+ $X2=0.795 $Y2=1.065
r548 161 182 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.735 $Y=2.12
+ $X2=0.735 $Y2=2.035
r549 161 163 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=0.735 $Y=2.12
+ $X2=0.735 $Y2=2.815
r550 157 166 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.67 $Y=0.98
+ $X2=0.795 $Y2=1.065
r551 157 159 18.4391 $w=2.48e-07 $l=4e-07 $layer=LI1_cond $X=0.67 $Y=0.98
+ $X2=0.67 $Y2=0.58
r552 153 267 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.105 $Y=1.19
+ $X2=9.105 $Y2=1.355
r553 153 155 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=9.105 $Y=1.19
+ $X2=9.105 $Y2=0.58
r554 150 152 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=9.09 $Y=1.765
+ $X2=9.09 $Y2=2.4
r555 149 150 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=9.09 $Y=1.675
+ $X2=9.09 $Y2=1.765
r556 148 266 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=9.09 $Y=1.52
+ $X2=9.09 $Y2=1.355
r557 148 149 60.25 $w=1.8e-07 $l=1.55e-07 $layer=POLY_cond $X=9.09 $Y=1.52
+ $X2=9.09 $Y2=1.675
r558 144 265 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.675 $Y=1.19
+ $X2=8.675 $Y2=1.355
r559 144 146 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=8.675 $Y=1.19
+ $X2=8.675 $Y2=0.58
r560 141 143 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=8.64 $Y=1.765
+ $X2=8.64 $Y2=2.4
r561 140 141 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=8.64 $Y=1.675
+ $X2=8.64 $Y2=1.765
r562 139 264 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=8.64 $Y=1.52
+ $X2=8.64 $Y2=1.355
r563 139 140 60.25 $w=1.8e-07 $l=1.55e-07 $layer=POLY_cond $X=8.64 $Y=1.52
+ $X2=8.64 $Y2=1.675
r564 135 260 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.175 $Y=1.19
+ $X2=8.175 $Y2=1.355
r565 135 137 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=8.175 $Y=1.19
+ $X2=8.175 $Y2=0.58
r566 132 134 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=8.17 $Y=1.765
+ $X2=8.17 $Y2=2.4
r567 131 132 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=8.17 $Y=1.675
+ $X2=8.17 $Y2=1.765
r568 130 259 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=8.17 $Y=1.52
+ $X2=8.17 $Y2=1.355
r569 130 131 60.25 $w=1.8e-07 $l=1.55e-07 $layer=POLY_cond $X=8.17 $Y=1.52
+ $X2=8.17 $Y2=1.675
r570 126 258 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.745 $Y=1.19
+ $X2=7.745 $Y2=1.355
r571 126 128 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=7.745 $Y=1.19
+ $X2=7.745 $Y2=0.58
r572 123 125 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=7.72 $Y=1.765
+ $X2=7.72 $Y2=2.4
r573 122 123 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=7.72 $Y=1.675
+ $X2=7.72 $Y2=1.765
r574 121 257 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=7.72 $Y=1.52
+ $X2=7.72 $Y2=1.355
r575 121 122 60.25 $w=1.8e-07 $l=1.55e-07 $layer=POLY_cond $X=7.72 $Y=1.52
+ $X2=7.72 $Y2=1.675
r576 118 120 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=7.27 $Y=1.765
+ $X2=7.27 $Y2=2.4
r577 117 118 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=7.27 $Y=1.675
+ $X2=7.27 $Y2=1.765
r578 116 253 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=7.27 $Y=1.52
+ $X2=7.27 $Y2=1.355
r579 116 117 60.25 $w=1.8e-07 $l=1.55e-07 $layer=POLY_cond $X=7.27 $Y=1.52
+ $X2=7.27 $Y2=1.675
r580 112 252 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.245 $Y=1.19
+ $X2=7.245 $Y2=1.355
r581 112 114 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=7.245 $Y=1.19
+ $X2=7.245 $Y2=0.58
r582 109 111 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=6.82 $Y=1.765
+ $X2=6.82 $Y2=2.4
r583 105 250 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.815 $Y=1.19
+ $X2=6.815 $Y2=1.355
r584 105 107 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=6.815 $Y=1.19
+ $X2=6.815 $Y2=0.58
r585 104 109 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=6.82 $Y=1.675
+ $X2=6.82 $Y2=1.765
r586 103 251 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=6.82 $Y=1.52
+ $X2=6.82 $Y2=1.355
r587 103 104 60.25 $w=1.8e-07 $l=1.55e-07 $layer=POLY_cond $X=6.82 $Y=1.52
+ $X2=6.82 $Y2=1.675
r588 100 102 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=6.37 $Y=1.765
+ $X2=6.37 $Y2=2.4
r589 99 100 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=6.37 $Y=1.675
+ $X2=6.37 $Y2=1.765
r590 98 246 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=6.37 $Y=1.52
+ $X2=6.37 $Y2=1.355
r591 98 99 60.25 $w=1.8e-07 $l=1.55e-07 $layer=POLY_cond $X=6.37 $Y=1.52
+ $X2=6.37 $Y2=1.675
r592 94 245 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.315 $Y=1.19
+ $X2=6.315 $Y2=1.355
r593 94 96 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=6.315 $Y=1.19
+ $X2=6.315 $Y2=0.58
r594 91 93 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=5.92 $Y=1.765
+ $X2=5.92 $Y2=2.4
r595 90 91 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=5.92 $Y=1.675
+ $X2=5.92 $Y2=1.765
r596 89 244 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=5.92 $Y=1.52
+ $X2=5.92 $Y2=1.355
r597 89 90 60.25 $w=1.8e-07 $l=1.55e-07 $layer=POLY_cond $X=5.92 $Y=1.52
+ $X2=5.92 $Y2=1.675
r598 85 243 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.885 $Y=1.19
+ $X2=5.885 $Y2=1.355
r599 85 87 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=5.885 $Y=1.19
+ $X2=5.885 $Y2=0.58
r600 82 84 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=5.47 $Y=1.765
+ $X2=5.47 $Y2=2.4
r601 81 82 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=5.47 $Y=1.675
+ $X2=5.47 $Y2=1.765
r602 80 239 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=5.47 $Y=1.52
+ $X2=5.47 $Y2=1.355
r603 80 81 60.25 $w=1.8e-07 $l=1.55e-07 $layer=POLY_cond $X=5.47 $Y=1.52
+ $X2=5.47 $Y2=1.675
r604 76 238 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.385 $Y=1.19
+ $X2=5.385 $Y2=1.355
r605 76 78 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=5.385 $Y=1.19
+ $X2=5.385 $Y2=0.58
r606 73 75 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=5.02 $Y=1.765
+ $X2=5.02 $Y2=2.4
r607 72 73 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=5.02 $Y=1.675
+ $X2=5.02 $Y2=1.765
r608 71 237 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=5.02 $Y=1.52
+ $X2=5.02 $Y2=1.355
r609 71 72 60.25 $w=1.8e-07 $l=1.55e-07 $layer=POLY_cond $X=5.02 $Y=1.52
+ $X2=5.02 $Y2=1.675
r610 67 236 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.955 $Y=1.19
+ $X2=4.955 $Y2=1.355
r611 67 69 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=4.955 $Y=1.19
+ $X2=4.955 $Y2=0.58
r612 64 66 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=4.57 $Y=1.765
+ $X2=4.57 $Y2=2.4
r613 63 64 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=4.57 $Y=1.675
+ $X2=4.57 $Y2=1.765
r614 62 232 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=4.57 $Y=1.52
+ $X2=4.57 $Y2=1.355
r615 62 63 60.25 $w=1.8e-07 $l=1.55e-07 $layer=POLY_cond $X=4.57 $Y=1.52
+ $X2=4.57 $Y2=1.675
r616 58 231 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.455 $Y=1.19
+ $X2=4.455 $Y2=1.355
r617 58 60 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=4.455 $Y=1.19
+ $X2=4.455 $Y2=0.58
r618 55 57 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=4.12 $Y=1.765
+ $X2=4.12 $Y2=2.4
r619 54 55 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=4.12 $Y=1.675
+ $X2=4.12 $Y2=1.765
r620 53 230 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=4.12 $Y=1.52
+ $X2=4.12 $Y2=1.355
r621 53 54 60.25 $w=1.8e-07 $l=1.55e-07 $layer=POLY_cond $X=4.12 $Y=1.52
+ $X2=4.12 $Y2=1.675
r622 49 229 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.025 $Y=1.19
+ $X2=4.025 $Y2=1.355
r623 49 51 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=4.025 $Y=1.19
+ $X2=4.025 $Y2=0.58
r624 46 48 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.67 $Y=1.765
+ $X2=3.67 $Y2=2.4
r625 45 46 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=3.67 $Y=1.675
+ $X2=3.67 $Y2=1.765
r626 44 225 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=3.67 $Y=1.52
+ $X2=3.67 $Y2=1.355
r627 44 45 60.25 $w=1.8e-07 $l=1.55e-07 $layer=POLY_cond $X=3.67 $Y=1.52
+ $X2=3.67 $Y2=1.675
r628 40 224 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.595 $Y=1.19
+ $X2=3.595 $Y2=1.355
r629 40 42 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=3.595 $Y=1.19
+ $X2=3.595 $Y2=0.58
r630 37 39 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.22 $Y=1.765
+ $X2=3.22 $Y2=2.4
r631 36 37 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=3.22 $Y=1.675
+ $X2=3.22 $Y2=1.765
r632 35 223 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=3.22 $Y=1.52
+ $X2=3.22 $Y2=1.355
r633 35 36 60.25 $w=1.8e-07 $l=1.55e-07 $layer=POLY_cond $X=3.22 $Y=1.52
+ $X2=3.22 $Y2=1.675
r634 31 222 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.165 $Y=1.19
+ $X2=3.165 $Y2=1.355
r635 31 33 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=3.165 $Y=1.19
+ $X2=3.165 $Y2=0.58
r636 28 30 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.77 $Y=1.765
+ $X2=2.77 $Y2=2.4
r637 27 28 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=2.77 $Y=1.675
+ $X2=2.77 $Y2=1.765
r638 26 218 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=2.77 $Y=1.52
+ $X2=2.77 $Y2=1.355
r639 26 27 60.25 $w=1.8e-07 $l=1.55e-07 $layer=POLY_cond $X=2.77 $Y=1.52
+ $X2=2.77 $Y2=1.675
r640 22 217 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.735 $Y=1.19
+ $X2=2.735 $Y2=1.355
r641 22 24 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.735 $Y=1.19
+ $X2=2.735 $Y2=0.58
r642 19 21 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.32 $Y=1.765
+ $X2=2.32 $Y2=2.4
r643 18 19 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=2.32 $Y=1.675
+ $X2=2.32 $Y2=1.765
r644 17 216 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=2.32 $Y=1.52
+ $X2=2.32 $Y2=1.355
r645 17 18 60.25 $w=1.8e-07 $l=1.55e-07 $layer=POLY_cond $X=2.32 $Y=1.52
+ $X2=2.32 $Y2=1.675
r646 13 214 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.305 $Y=1.19
+ $X2=2.305 $Y2=1.355
r647 13 15 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.305 $Y=1.19
+ $X2=2.305 $Y2=0.58
r648 4 185 400 $w=1.7e-07 $l=3.4187e-07 $layer=licon1_PDIFF $count=1 $X=1.485
+ $Y=1.84 $X2=1.635 $Y2=2.115
r649 4 175 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=1.485
+ $Y=1.84 $X2=1.635 $Y2=2.815
r650 3 182 400 $w=1.7e-07 $l=3.4187e-07 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=1.84 $X2=0.735 $Y2=2.115
r651 3 163 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=1.84 $X2=0.735 $Y2=2.815
r652 2 171 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.45
+ $Y=0.37 $X2=1.59 $Y2=0.58
r653 1 159 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.37 $X2=0.71 $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_HS__CLKBUF_16%VPWR 1 2 3 4 5 6 7 8 9 10 11 34 36 42 46
+ 50 56 62 68 72 76 82 88 92 94 99 100 102 103 105 106 108 109 110 111 112 118
+ 135 140 145 154 157 160 163 167
r192 166 167 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.36 $Y=3.33
+ $X2=9.36 $Y2=3.33
r193 163 164 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=3.33
+ $X2=8.4 $Y2=3.33
r194 160 161 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r195 157 158 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r196 154 155 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r197 151 152 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r198 149 167 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=3.33
+ $X2=9.36 $Y2=3.33
r199 149 164 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=3.33
+ $X2=8.4 $Y2=3.33
r200 148 149 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r201 146 163 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.56 $Y=3.33
+ $X2=8.395 $Y2=3.33
r202 146 148 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=8.56 $Y=3.33
+ $X2=8.88 $Y2=3.33
r203 145 166 4.72267 $w=1.7e-07 $l=2.25e-07 $layer=LI1_cond $X=9.15 $Y=3.33
+ $X2=9.375 $Y2=3.33
r204 145 148 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=9.15 $Y=3.33
+ $X2=8.88 $Y2=3.33
r205 144 164 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=3.33
+ $X2=8.4 $Y2=3.33
r206 144 161 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=3.33
+ $X2=7.44 $Y2=3.33
r207 143 144 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r208 141 160 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.66 $Y=3.33
+ $X2=7.495 $Y2=3.33
r209 141 143 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=7.66 $Y=3.33
+ $X2=7.92 $Y2=3.33
r210 140 163 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.23 $Y=3.33
+ $X2=8.395 $Y2=3.33
r211 140 143 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=8.23 $Y=3.33
+ $X2=7.92 $Y2=3.33
r212 139 161 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=7.44 $Y2=3.33
r213 139 158 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=6.48 $Y2=3.33
r214 138 139 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r215 136 157 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.76 $Y=3.33
+ $X2=6.595 $Y2=3.33
r216 136 138 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=6.76 $Y=3.33
+ $X2=6.96 $Y2=3.33
r217 135 160 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.33 $Y=3.33
+ $X2=7.495 $Y2=3.33
r218 135 138 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=7.33 $Y=3.33
+ $X2=6.96 $Y2=3.33
r219 134 158 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=6.48 $Y2=3.33
r220 133 134 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r221 130 131 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r222 128 131 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.56 $Y2=3.33
r223 127 128 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r224 125 128 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.6 $Y2=3.33
r225 125 155 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=2.16 $Y2=3.33
r226 124 125 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r227 122 154 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.25 $Y=3.33
+ $X2=2.125 $Y2=3.33
r228 122 124 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=2.25 $Y=3.33
+ $X2=2.64 $Y2=3.33
r229 121 155 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r230 120 121 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r231 118 154 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2 $Y=3.33
+ $X2=2.125 $Y2=3.33
r232 118 120 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=2 $Y=3.33 $X2=1.68
+ $Y2=3.33
r233 117 121 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.68 $Y2=3.33
r234 117 152 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r235 116 117 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r236 114 151 4.0045 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=0.37 $Y=3.33
+ $X2=0.185 $Y2=3.33
r237 114 116 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=0.37 $Y=3.33
+ $X2=0.72 $Y2=3.33
r238 112 134 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=4.8 $Y=3.33
+ $X2=5.52 $Y2=3.33
r239 112 131 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=4.8 $Y=3.33
+ $X2=4.56 $Y2=3.33
r240 110 133 0.652406 $w=1.68e-07 $l=1e-08 $layer=LI1_cond $X=5.53 $Y=3.33
+ $X2=5.52 $Y2=3.33
r241 110 111 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.53 $Y=3.33
+ $X2=5.695 $Y2=3.33
r242 108 130 4.56684 $w=1.68e-07 $l=7e-08 $layer=LI1_cond $X=4.63 $Y=3.33
+ $X2=4.56 $Y2=3.33
r243 108 109 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.63 $Y=3.33
+ $X2=4.795 $Y2=3.33
r244 107 133 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=4.96 $Y=3.33
+ $X2=5.52 $Y2=3.33
r245 107 109 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.96 $Y=3.33
+ $X2=4.795 $Y2=3.33
r246 105 127 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=3.73 $Y=3.33
+ $X2=3.6 $Y2=3.33
r247 105 106 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.73 $Y=3.33
+ $X2=3.895 $Y2=3.33
r248 104 130 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=4.06 $Y=3.33
+ $X2=4.56 $Y2=3.33
r249 104 106 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.06 $Y=3.33
+ $X2=3.895 $Y2=3.33
r250 102 124 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=2.83 $Y=3.33
+ $X2=2.64 $Y2=3.33
r251 102 103 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.83 $Y=3.33
+ $X2=2.995 $Y2=3.33
r252 101 127 28.7059 $w=1.68e-07 $l=4.4e-07 $layer=LI1_cond $X=3.16 $Y=3.33
+ $X2=3.6 $Y2=3.33
r253 101 103 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.16 $Y=3.33
+ $X2=2.995 $Y2=3.33
r254 99 116 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=1.1 $Y=3.33
+ $X2=0.72 $Y2=3.33
r255 99 100 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.1 $Y=3.33
+ $X2=1.185 $Y2=3.33
r256 98 120 26.7487 $w=1.68e-07 $l=4.1e-07 $layer=LI1_cond $X=1.27 $Y=3.33
+ $X2=1.68 $Y2=3.33
r257 98 100 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.27 $Y=3.33
+ $X2=1.185 $Y2=3.33
r258 94 97 24.4458 $w=3.28e-07 $l=7e-07 $layer=LI1_cond $X=9.315 $Y=2.115
+ $X2=9.315 $Y2=2.815
r259 92 166 3.0435 $w=3.3e-07 $l=1.11018e-07 $layer=LI1_cond $X=9.315 $Y=3.245
+ $X2=9.375 $Y2=3.33
r260 92 97 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=9.315 $Y=3.245
+ $X2=9.315 $Y2=2.815
r261 88 91 24.4458 $w=3.28e-07 $l=7e-07 $layer=LI1_cond $X=8.395 $Y=2.115
+ $X2=8.395 $Y2=2.815
r262 86 163 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.395 $Y=3.245
+ $X2=8.395 $Y2=3.33
r263 86 91 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=8.395 $Y=3.245
+ $X2=8.395 $Y2=2.815
r264 82 85 24.4458 $w=3.28e-07 $l=7e-07 $layer=LI1_cond $X=7.495 $Y=2.115
+ $X2=7.495 $Y2=2.815
r265 80 160 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.495 $Y=3.245
+ $X2=7.495 $Y2=3.33
r266 80 85 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=7.495 $Y=3.245
+ $X2=7.495 $Y2=2.815
r267 76 79 24.4458 $w=3.28e-07 $l=7e-07 $layer=LI1_cond $X=6.595 $Y=2.115
+ $X2=6.595 $Y2=2.815
r268 74 157 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.595 $Y=3.245
+ $X2=6.595 $Y2=3.33
r269 74 79 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=6.595 $Y=3.245
+ $X2=6.595 $Y2=2.815
r270 73 111 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.86 $Y=3.33
+ $X2=5.695 $Y2=3.33
r271 72 157 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.43 $Y=3.33
+ $X2=6.595 $Y2=3.33
r272 72 73 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=6.43 $Y=3.33
+ $X2=5.86 $Y2=3.33
r273 68 71 24.4458 $w=3.28e-07 $l=7e-07 $layer=LI1_cond $X=5.695 $Y=2.115
+ $X2=5.695 $Y2=2.815
r274 66 111 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.695 $Y=3.245
+ $X2=5.695 $Y2=3.33
r275 66 71 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=5.695 $Y=3.245
+ $X2=5.695 $Y2=2.815
r276 62 65 24.4458 $w=3.28e-07 $l=7e-07 $layer=LI1_cond $X=4.795 $Y=2.115
+ $X2=4.795 $Y2=2.815
r277 60 109 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.795 $Y=3.245
+ $X2=4.795 $Y2=3.33
r278 60 65 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=4.795 $Y=3.245
+ $X2=4.795 $Y2=2.815
r279 56 59 24.4458 $w=3.28e-07 $l=7e-07 $layer=LI1_cond $X=3.895 $Y=2.115
+ $X2=3.895 $Y2=2.815
r280 54 106 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.895 $Y=3.245
+ $X2=3.895 $Y2=3.33
r281 54 59 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=3.895 $Y=3.245
+ $X2=3.895 $Y2=2.815
r282 50 53 24.4458 $w=3.28e-07 $l=7e-07 $layer=LI1_cond $X=2.995 $Y=2.115
+ $X2=2.995 $Y2=2.815
r283 48 103 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.995 $Y=3.245
+ $X2=2.995 $Y2=3.33
r284 48 53 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=2.995 $Y=3.245
+ $X2=2.995 $Y2=2.815
r285 44 154 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.125 $Y=3.245
+ $X2=2.125 $Y2=3.33
r286 44 46 36.4172 $w=2.48e-07 $l=7.9e-07 $layer=LI1_cond $X=2.125 $Y=3.245
+ $X2=2.125 $Y2=2.455
r287 40 100 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.185 $Y=3.245
+ $X2=1.185 $Y2=3.33
r288 40 42 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=1.185 $Y=3.245
+ $X2=1.185 $Y2=2.455
r289 36 39 32.2684 $w=2.48e-07 $l=7e-07 $layer=LI1_cond $X=0.245 $Y=2.115
+ $X2=0.245 $Y2=2.815
r290 34 151 3.13866 $w=2.5e-07 $l=1.11018e-07 $layer=LI1_cond $X=0.245 $Y=3.245
+ $X2=0.185 $Y2=3.33
r291 34 39 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=0.245 $Y=3.245
+ $X2=0.245 $Y2=2.815
r292 11 97 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=9.165
+ $Y=1.84 $X2=9.315 $Y2=2.815
r293 11 94 400 $w=1.7e-07 $l=3.4187e-07 $layer=licon1_PDIFF $count=1 $X=9.165
+ $Y=1.84 $X2=9.315 $Y2=2.115
r294 10 91 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=8.245
+ $Y=1.84 $X2=8.395 $Y2=2.815
r295 10 88 400 $w=1.7e-07 $l=3.4187e-07 $layer=licon1_PDIFF $count=1 $X=8.245
+ $Y=1.84 $X2=8.395 $Y2=2.115
r296 9 85 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=7.345
+ $Y=1.84 $X2=7.495 $Y2=2.815
r297 9 82 400 $w=1.7e-07 $l=3.4187e-07 $layer=licon1_PDIFF $count=1 $X=7.345
+ $Y=1.84 $X2=7.495 $Y2=2.115
r298 8 79 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=6.445
+ $Y=1.84 $X2=6.595 $Y2=2.815
r299 8 76 400 $w=1.7e-07 $l=3.4187e-07 $layer=licon1_PDIFF $count=1 $X=6.445
+ $Y=1.84 $X2=6.595 $Y2=2.115
r300 7 71 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=5.545
+ $Y=1.84 $X2=5.695 $Y2=2.815
r301 7 68 400 $w=1.7e-07 $l=3.4187e-07 $layer=licon1_PDIFF $count=1 $X=5.545
+ $Y=1.84 $X2=5.695 $Y2=2.115
r302 6 65 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=4.645
+ $Y=1.84 $X2=4.795 $Y2=2.815
r303 6 62 400 $w=1.7e-07 $l=3.4187e-07 $layer=licon1_PDIFF $count=1 $X=4.645
+ $Y=1.84 $X2=4.795 $Y2=2.115
r304 5 59 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=3.745
+ $Y=1.84 $X2=3.895 $Y2=2.815
r305 5 56 400 $w=1.7e-07 $l=3.4187e-07 $layer=licon1_PDIFF $count=1 $X=3.745
+ $Y=1.84 $X2=3.895 $Y2=2.115
r306 4 53 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=2.845
+ $Y=1.84 $X2=2.995 $Y2=2.815
r307 4 50 400 $w=1.7e-07 $l=3.4187e-07 $layer=licon1_PDIFF $count=1 $X=2.845
+ $Y=1.84 $X2=2.995 $Y2=2.115
r308 3 46 300 $w=1.7e-07 $l=6.85912e-07 $layer=licon1_PDIFF $count=2 $X=1.935
+ $Y=1.84 $X2=2.085 $Y2=2.455
r309 2 42 300 $w=1.7e-07 $l=6.85912e-07 $layer=licon1_PDIFF $count=2 $X=1.035
+ $Y=1.84 $X2=1.185 $Y2=2.455
r310 1 39 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=0.14
+ $Y=1.84 $X2=0.285 $Y2=2.815
r311 1 36 400 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_PDIFF $count=1 $X=0.14
+ $Y=1.84 $X2=0.285 $Y2=2.115
.ends

.subckt PM_SKY130_FD_SC_HS__CLKBUF_16%X 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16
+ 51 55 59 65 69 73 77 79 81 85 87 91 92 95 98 101 104 106 109 116 123 130 137
+ 144 151 153 161
c266 153 0 1.65196e-19 $X=8.865 $Y=2.035
c267 79 0 1.75614e-19 $X=8.85 $Y=1.705
r268 158 161 6.04804 $w=2.68e-07 $l=1.35e-07 $layer=LI1_cond $X=2.525 $Y=1.985
+ $X2=2.525 $Y2=2.12
r269 158 160 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.545 $Y=2.035
+ $X2=2.545 $Y2=2.035
r270 151 155 43.4785 $w=2.18e-07 $l=8.3e-07 $layer=LI1_cond $X=8.86 $Y=1.985
+ $X2=8.86 $Y2=2.815
r271 151 153 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.865 $Y=2.035
+ $X2=8.865 $Y2=2.035
r272 146 153 0.590276 $w=2.3e-07 $l=9.2e-07 $layer=MET1_cond $X=7.945 $Y=2.035
+ $X2=8.865 $Y2=2.035
r273 144 148 43.8355 $w=2.08e-07 $l=8.3e-07 $layer=LI1_cond $X=7.945 $Y=1.985
+ $X2=7.945 $Y2=2.815
r274 144 146 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.945 $Y=2.035
+ $X2=7.945 $Y2=2.035
r275 139 146 0.577444 $w=2.3e-07 $l=9e-07 $layer=MET1_cond $X=7.045 $Y=2.035
+ $X2=7.945 $Y2=2.035
r276 137 141 44.9047 $w=2.03e-07 $l=8.3e-07 $layer=LI1_cond $X=7.047 $Y=1.985
+ $X2=7.047 $Y2=2.815
r277 137 139 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.045 $Y=2.035
+ $X2=7.045 $Y2=2.035
r278 132 139 0.577444 $w=2.3e-07 $l=9e-07 $layer=MET1_cond $X=6.145 $Y=2.035
+ $X2=7.045 $Y2=2.035
r279 130 134 44.9047 $w=2.03e-07 $l=8.3e-07 $layer=LI1_cond $X=6.142 $Y=1.985
+ $X2=6.142 $Y2=2.815
r280 130 132 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.145 $Y=2.035
+ $X2=6.145 $Y2=2.035
r281 123 127 43.8355 $w=2.08e-07 $l=8.3e-07 $layer=LI1_cond $X=5.245 $Y=1.985
+ $X2=5.245 $Y2=2.815
r282 123 125 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.245 $Y=2.035
+ $X2=5.245 $Y2=2.035
r283 118 125 0.587068 $w=2.3e-07 $l=9.15e-07 $layer=MET1_cond $X=4.33 $Y=2.035
+ $X2=5.245 $Y2=2.035
r284 116 120 46.0273 $w=1.98e-07 $l=8.3e-07 $layer=LI1_cond $X=4.33 $Y=1.985
+ $X2=4.33 $Y2=2.815
r285 116 118 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.33 $Y=2.035
+ $X2=4.33 $Y2=2.035
r286 111 118 0.56782 $w=2.3e-07 $l=8.85e-07 $layer=MET1_cond $X=3.445 $Y=2.035
+ $X2=4.33 $Y2=2.035
r287 111 160 0.577444 $w=2.3e-07 $l=9e-07 $layer=MET1_cond $X=3.445 $Y=2.035
+ $X2=2.545 $Y2=2.035
r288 109 113 44.9047 $w=2.03e-07 $l=8.3e-07 $layer=LI1_cond $X=3.442 $Y=1.985
+ $X2=3.442 $Y2=2.815
r289 109 111 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.445 $Y=2.035
+ $X2=3.445 $Y2=2.035
r290 106 132 0.25985 $w=2.3e-07 $l=4.05e-07 $layer=MET1_cond $X=5.74 $Y=2.035
+ $X2=6.145 $Y2=2.035
r291 106 125 0.317594 $w=2.3e-07 $l=4.95e-07 $layer=MET1_cond $X=5.74 $Y=2.035
+ $X2=5.245 $Y2=2.035
r292 105 151 6.54797 $w=2.18e-07 $l=1.25e-07 $layer=LI1_cond $X=8.86 $Y=1.86
+ $X2=8.86 $Y2=1.985
r293 104 144 6.60173 $w=2.08e-07 $l=1.25e-07 $layer=LI1_cond $X=7.945 $Y=1.86
+ $X2=7.945 $Y2=1.985
r294 103 104 8.16535 $w=2.48e-07 $l=1.7e-07 $layer=LI1_cond $X=7.922 $Y=1.69
+ $X2=7.922 $Y2=1.86
r295 101 137 6.76275 $w=2.03e-07 $l=1.25e-07 $layer=LI1_cond $X=7.047 $Y=1.86
+ $X2=7.047 $Y2=1.985
r296 100 101 8.24408 $w=2.48e-07 $l=1.7e-07 $layer=LI1_cond $X=7.007 $Y=1.69
+ $X2=7.007 $Y2=1.86
r297 98 130 6.76275 $w=2.03e-07 $l=1.25e-07 $layer=LI1_cond $X=6.142 $Y=1.86
+ $X2=6.142 $Y2=1.985
r298 97 98 8.24408 $w=2.48e-07 $l=1.7e-07 $layer=LI1_cond $X=6.09 $Y=1.69
+ $X2=6.09 $Y2=1.86
r299 95 123 6.60173 $w=2.08e-07 $l=1.25e-07 $layer=LI1_cond $X=5.245 $Y=1.86
+ $X2=5.245 $Y2=1.985
r300 94 95 8.62714 $w=2.28e-07 $l=1.7e-07 $layer=LI1_cond $X=5.187 $Y=1.69
+ $X2=5.187 $Y2=1.86
r301 92 116 6.93182 $w=1.98e-07 $l=1.25e-07 $layer=LI1_cond $X=4.33 $Y=1.86
+ $X2=4.33 $Y2=1.985
r302 91 92 9.70862 $w=1.98e-07 $l=1.7e-07 $layer=LI1_cond $X=4.3 $Y=1.69 $X2=4.3
+ $Y2=1.86
r303 89 91 61.6524 $w=1.68e-07 $l=9.45e-07 $layer=LI1_cond $X=4.255 $Y=0.745
+ $X2=4.255 $Y2=1.69
r304 87 89 8.65224 $w=2.63e-07 $l=1.65e-07 $layer=LI1_cond $X=4.207 $Y=0.58
+ $X2=4.207 $Y2=0.745
r305 85 109 6.76275 $w=2.03e-07 $l=1.25e-07 $layer=LI1_cond $X=3.442 $Y=1.86
+ $X2=3.442 $Y2=1.985
r306 84 85 8.82084 $w=2.23e-07 $l=1.7e-07 $layer=LI1_cond $X=3.41 $Y=1.69
+ $X2=3.41 $Y2=1.86
r307 79 105 7.59438 $w=2.49e-07 $l=1.59922e-07 $layer=LI1_cond $X=8.85 $Y=1.705
+ $X2=8.86 $Y2=1.86
r308 79 81 51.8599 $w=2.48e-07 $l=1.125e-06 $layer=LI1_cond $X=8.85 $Y=1.705
+ $X2=8.85 $Y2=0.58
r309 77 103 51.1685 $w=2.48e-07 $l=1.11e-06 $layer=LI1_cond $X=7.92 $Y=0.58
+ $X2=7.92 $Y2=1.69
r310 73 100 51.1685 $w=2.48e-07 $l=1.11e-06 $layer=LI1_cond $X=6.99 $Y=0.58
+ $X2=6.99 $Y2=1.69
r311 69 97 51.1685 $w=2.48e-07 $l=1.11e-06 $layer=LI1_cond $X=6.06 $Y=0.58
+ $X2=6.06 $Y2=1.69
r312 65 94 55.6179 $w=2.28e-07 $l=1.11e-06 $layer=LI1_cond $X=5.14 $Y=0.58
+ $X2=5.14 $Y2=1.69
r313 59 84 56.8539 $w=2.23e-07 $l=1.11e-06 $layer=LI1_cond $X=3.387 $Y=0.58
+ $X2=3.387 $Y2=1.69
r314 55 161 14.0297 $w=2.28e-07 $l=2.8e-07 $layer=LI1_cond $X=2.545 $Y=2.4
+ $X2=2.545 $Y2=2.12
r315 51 158 59.9697 $w=2.68e-07 $l=1.405e-06 $layer=LI1_cond $X=2.525 $Y=0.58
+ $X2=2.525 $Y2=1.985
r316 16 155 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=8.715
+ $Y=1.84 $X2=8.865 $Y2=2.815
r317 16 151 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=8.715
+ $Y=1.84 $X2=8.865 $Y2=1.985
r318 15 148 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=7.795
+ $Y=1.84 $X2=7.945 $Y2=2.815
r319 15 144 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=7.795
+ $Y=1.84 $X2=7.945 $Y2=1.985
r320 14 141 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=6.895
+ $Y=1.84 $X2=7.045 $Y2=2.815
r321 14 137 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=6.895
+ $Y=1.84 $X2=7.045 $Y2=1.985
r322 13 134 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=5.995
+ $Y=1.84 $X2=6.145 $Y2=2.815
r323 13 130 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=5.995
+ $Y=1.84 $X2=6.145 $Y2=1.985
r324 12 127 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=5.095
+ $Y=1.84 $X2=5.245 $Y2=2.815
r325 12 123 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=5.095
+ $Y=1.84 $X2=5.245 $Y2=1.985
r326 11 120 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=4.195
+ $Y=1.84 $X2=4.345 $Y2=2.815
r327 11 116 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=4.195
+ $Y=1.84 $X2=4.345 $Y2=1.985
r328 10 113 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=3.295
+ $Y=1.84 $X2=3.445 $Y2=2.815
r329 10 109 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=3.295
+ $Y=1.84 $X2=3.445 $Y2=1.985
r330 9 158 600 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=2.395
+ $Y=1.84 $X2=2.545 $Y2=1.985
r331 9 55 300 $w=1.7e-07 $l=6.30555e-07 $layer=licon1_PDIFF $count=2 $X=2.395
+ $Y=1.84 $X2=2.545 $Y2=2.4
r332 8 81 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=8.75
+ $Y=0.37 $X2=8.89 $Y2=0.58
r333 7 77 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=7.82
+ $Y=0.37 $X2=7.96 $Y2=0.58
r334 6 73 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=6.89
+ $Y=0.37 $X2=7.03 $Y2=0.58
r335 5 69 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=5.96
+ $Y=0.37 $X2=6.1 $Y2=0.58
r336 4 65 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=5.03
+ $Y=0.37 $X2=5.17 $Y2=0.58
r337 3 87 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=4.1
+ $Y=0.37 $X2=4.24 $Y2=0.58
r338 2 59 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=3.24
+ $Y=0.37 $X2=3.38 $Y2=0.58
r339 1 51 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.38
+ $Y=0.37 $X2=2.52 $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_HS__CLKBUF_16%VGND 1 2 3 4 5 6 7 8 9 10 11 34 36 40 44
+ 48 52 54 58 62 66 70 74 76 78 81 82 84 85 87 88 89 90 91 106 111 116 121 126
+ 135 138 141 144 147 151
r167 150 151 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.36 $Y=0
+ $X2=9.36 $Y2=0
r168 147 148 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r169 144 145 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=0
+ $X2=7.44 $Y2=0
r170 141 142 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=0
+ $X2=6.48 $Y2=0
r171 138 139 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=0
+ $X2=5.52 $Y2=0
r172 135 136 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=0
+ $X2=4.56 $Y2=0
r173 132 133 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0
+ $X2=0.24 $Y2=0
r174 130 151 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=0
+ $X2=9.36 $Y2=0
r175 130 148 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=0
+ $X2=8.4 $Y2=0
r176 129 130 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=0
+ $X2=8.88 $Y2=0
r177 127 147 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.555 $Y=0
+ $X2=8.39 $Y2=0
r178 127 129 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=8.555 $Y=0
+ $X2=8.88 $Y2=0
r179 126 150 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=9.155 $Y=0
+ $X2=9.377 $Y2=0
r180 126 129 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=9.155 $Y=0
+ $X2=8.88 $Y2=0
r181 125 148 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=0
+ $X2=8.4 $Y2=0
r182 125 145 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=0
+ $X2=7.44 $Y2=0
r183 124 125 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=0
+ $X2=7.92 $Y2=0
r184 122 144 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.625 $Y=0
+ $X2=7.46 $Y2=0
r185 122 124 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=7.625 $Y=0
+ $X2=7.92 $Y2=0
r186 121 147 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.225 $Y=0
+ $X2=8.39 $Y2=0
r187 121 124 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=8.225 $Y=0
+ $X2=7.92 $Y2=0
r188 120 145 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=0
+ $X2=7.44 $Y2=0
r189 120 142 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=0
+ $X2=6.48 $Y2=0
r190 119 120 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=0
+ $X2=6.96 $Y2=0
r191 117 141 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.695 $Y=0
+ $X2=6.53 $Y2=0
r192 117 119 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=6.695 $Y=0
+ $X2=6.96 $Y2=0
r193 116 144 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.295 $Y=0
+ $X2=7.46 $Y2=0
r194 116 119 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=7.295 $Y=0
+ $X2=6.96 $Y2=0
r195 115 142 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=0 $X2=6.48
+ $Y2=0
r196 115 139 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=0 $X2=5.52
+ $Y2=0
r197 114 115 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=0 $X2=6
+ $Y2=0
r198 112 138 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.765 $Y=0
+ $X2=5.6 $Y2=0
r199 112 114 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=5.765 $Y=0 $X2=6
+ $Y2=0
r200 111 141 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.365 $Y=0
+ $X2=6.53 $Y2=0
r201 111 114 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=6.365 $Y=0 $X2=6
+ $Y2=0
r202 110 139 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=0
+ $X2=5.52 $Y2=0
r203 109 110 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=0
+ $X2=5.04 $Y2=0
r204 107 135 8.5188 $w=1.7e-07 $l=1.63e-07 $layer=LI1_cond $X=4.835 $Y=0
+ $X2=4.672 $Y2=0
r205 107 109 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=4.835 $Y=0
+ $X2=5.04 $Y2=0
r206 106 138 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.435 $Y=0
+ $X2=5.6 $Y2=0
r207 106 109 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=5.435 $Y=0
+ $X2=5.04 $Y2=0
r208 105 136 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=0
+ $X2=4.56 $Y2=0
r209 104 105 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r210 102 105 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=0
+ $X2=3.6 $Y2=0
r211 101 102 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0
+ $X2=2.64 $Y2=0
r212 99 102 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0
+ $X2=2.64 $Y2=0
r213 98 99 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r214 96 99 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r215 96 133 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0
+ $X2=0.24 $Y2=0
r216 95 96 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r217 93 132 4.00981 $w=1.7e-07 $l=1.83e-07 $layer=LI1_cond $X=0.365 $Y=0
+ $X2=0.182 $Y2=0
r218 93 95 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=0.365 $Y=0
+ $X2=0.72 $Y2=0
r219 91 110 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=4.8 $Y=0
+ $X2=5.04 $Y2=0
r220 91 136 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=4.8 $Y=0
+ $X2=4.56 $Y2=0
r221 89 104 4.56684 $w=1.68e-07 $l=7e-08 $layer=LI1_cond $X=3.67 $Y=0 $X2=3.6
+ $Y2=0
r222 89 90 6.47928 $w=1.7e-07 $l=1.12e-07 $layer=LI1_cond $X=3.67 $Y=0 $X2=3.782
+ $Y2=0
r223 87 101 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=2.865 $Y=0
+ $X2=2.64 $Y2=0
r224 87 88 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.865 $Y=0 $X2=2.95
+ $Y2=0
r225 86 104 36.861 $w=1.68e-07 $l=5.65e-07 $layer=LI1_cond $X=3.035 $Y=0 $X2=3.6
+ $Y2=0
r226 86 88 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.035 $Y=0 $X2=2.95
+ $Y2=0
r227 84 98 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=1.855 $Y=0
+ $X2=1.68 $Y2=0
r228 84 85 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.855 $Y=0 $X2=2.02
+ $Y2=0
r229 83 101 29.6845 $w=1.68e-07 $l=4.55e-07 $layer=LI1_cond $X=2.185 $Y=0
+ $X2=2.64 $Y2=0
r230 83 85 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.185 $Y=0 $X2=2.02
+ $Y2=0
r231 81 95 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.975 $Y=0
+ $X2=0.72 $Y2=0
r232 81 82 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.975 $Y=0 $X2=1.1
+ $Y2=0
r233 80 98 29.6845 $w=1.68e-07 $l=4.55e-07 $layer=LI1_cond $X=1.225 $Y=0
+ $X2=1.68 $Y2=0
r234 80 82 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.225 $Y=0 $X2=1.1
+ $Y2=0
r235 76 150 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=9.32 $Y=0.085
+ $X2=9.377 $Y2=0
r236 76 78 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=9.32 $Y=0.085
+ $X2=9.32 $Y2=0.58
r237 72 147 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.39 $Y=0.085
+ $X2=8.39 $Y2=0
r238 72 74 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=8.39 $Y=0.085
+ $X2=8.39 $Y2=0.515
r239 68 144 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.46 $Y=0.085
+ $X2=7.46 $Y2=0
r240 68 70 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=7.46 $Y=0.085
+ $X2=7.46 $Y2=0.515
r241 64 141 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.53 $Y=0.085
+ $X2=6.53 $Y2=0
r242 64 66 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=6.53 $Y=0.085
+ $X2=6.53 $Y2=0.515
r243 60 138 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.6 $Y=0.085
+ $X2=5.6 $Y2=0
r244 60 62 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=5.6 $Y=0.085
+ $X2=5.6 $Y2=0.515
r245 56 135 0.848899 $w=3.25e-07 $l=8.5e-08 $layer=LI1_cond $X=4.672 $Y=0.085
+ $X2=4.672 $Y2=0
r246 56 58 17.3753 $w=3.23e-07 $l=4.9e-07 $layer=LI1_cond $X=4.672 $Y=0.085
+ $X2=4.672 $Y2=0.575
r247 55 90 6.47928 $w=1.7e-07 $l=1.13e-07 $layer=LI1_cond $X=3.895 $Y=0
+ $X2=3.782 $Y2=0
r248 54 135 8.5188 $w=1.7e-07 $l=1.62e-07 $layer=LI1_cond $X=4.51 $Y=0 $X2=4.672
+ $Y2=0
r249 54 55 40.123 $w=1.68e-07 $l=6.15e-07 $layer=LI1_cond $X=4.51 $Y=0 $X2=3.895
+ $Y2=0
r250 50 90 0.355529 $w=2.25e-07 $l=8.5e-08 $layer=LI1_cond $X=3.782 $Y=0.085
+ $X2=3.782 $Y2=0
r251 50 52 24.3294 $w=2.23e-07 $l=4.75e-07 $layer=LI1_cond $X=3.782 $Y=0.085
+ $X2=3.782 $Y2=0.56
r252 46 88 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.95 $Y=0.085
+ $X2=2.95 $Y2=0
r253 46 48 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=2.95 $Y=0.085
+ $X2=2.95 $Y2=0.515
r254 42 85 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.02 $Y=0.085
+ $X2=2.02 $Y2=0
r255 42 44 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=2.02 $Y=0.085
+ $X2=2.02 $Y2=0.58
r256 38 82 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.1 $Y=0.085
+ $X2=1.1 $Y2=0
r257 38 40 22.8184 $w=2.48e-07 $l=4.95e-07 $layer=LI1_cond $X=1.1 $Y=0.085
+ $X2=1.1 $Y2=0.58
r258 34 132 3.13335 $w=2.5e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.24 $Y=0.085
+ $X2=0.182 $Y2=0
r259 34 36 22.8184 $w=2.48e-07 $l=4.95e-07 $layer=LI1_cond $X=0.24 $Y=0.085
+ $X2=0.24 $Y2=0.58
r260 11 78 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=9.18
+ $Y=0.37 $X2=9.32 $Y2=0.58
r261 10 74 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=8.25
+ $Y=0.37 $X2=8.39 $Y2=0.515
r262 9 70 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=7.32
+ $Y=0.37 $X2=7.46 $Y2=0.515
r263 8 66 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=6.39
+ $Y=0.37 $X2=6.53 $Y2=0.515
r264 7 62 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=5.46
+ $Y=0.37 $X2=5.6 $Y2=0.515
r265 6 58 182 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_NDIFF $count=1 $X=4.53
+ $Y=0.37 $X2=4.67 $Y2=0.575
r266 5 52 182 $w=1.7e-07 $l=2.504e-07 $layer=licon1_NDIFF $count=1 $X=3.67
+ $Y=0.37 $X2=3.81 $Y2=0.56
r267 4 48 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=2.81
+ $Y=0.37 $X2=2.95 $Y2=0.515
r268 3 44 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.88
+ $Y=0.37 $X2=2.02 $Y2=0.58
r269 2 40 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1
+ $Y=0.37 $X2=1.14 $Y2=0.58
r270 1 36 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.58
.ends

