* NGSPICE file created from sky130_fd_sc_hs__a2111o_2.ext - technology: sky130A

.subckt sky130_fd_sc_hs__a2111o_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
M1000 a_522_368# C1 a_444_368# VPB pshort w=1.12e+06u l=150000u
+  ad=4.368e+11p pd=3.02e+06u as=2.688e+11p ps=2.72e+06u
M1001 a_444_368# D1 a_91_244# VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=3.08e+11p ps=2.79e+06u
M1002 a_630_368# B1 a_522_368# VPB pshort w=1.12e+06u l=150000u
+  ad=7.448e+11p pd=5.81e+06u as=0p ps=0u
M1003 VPWR A2 a_630_368# VPB pshort w=1.12e+06u l=150000u
+  ad=1.0528e+12p pd=8.6e+06u as=0p ps=0u
M1004 a_91_244# C1 VGND VNB nlowvt w=740000u l=150000u
+  ad=5.994e+11p pd=6.06e+06u as=1.0508e+12p ps=8.76e+06u
M1005 VGND a_91_244# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.072e+11p ps=2.04e+06u
M1006 X a_91_244# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_771_74# A2 VGND VNB nlowvt w=740000u l=150000u
+  ad=1.554e+11p pd=1.9e+06u as=0p ps=0u
M1008 a_91_244# A1 a_771_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VGND B1 a_91_244# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VGND D1 a_91_244# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 X a_91_244# VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=3.36e+11p pd=2.84e+06u as=0p ps=0u
M1012 VPWR a_91_244# X VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_630_368# A1 VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

