* File: sky130_fd_sc_hs__o21a_2.pxi.spice
* Created: Tue Sep  1 20:14:18 2020
* 
x_PM_SKY130_FD_SC_HS__O21A_2%A1 N_A1_c_59_n N_A1_M1006_g N_A1_c_60_n
+ N_A1_M1001_g N_A1_c_61_n A1 A1 PM_SKY130_FD_SC_HS__O21A_2%A1
x_PM_SKY130_FD_SC_HS__O21A_2%A2 N_A2_c_82_n N_A2_M1004_g N_A2_c_83_n
+ N_A2_M1002_g A2 PM_SKY130_FD_SC_HS__O21A_2%A2
x_PM_SKY130_FD_SC_HS__O21A_2%B1 N_B1_c_109_n N_B1_M1003_g N_B1_c_110_n
+ N_B1_M1009_g B1 N_B1_c_111_n PM_SKY130_FD_SC_HS__O21A_2%B1
x_PM_SKY130_FD_SC_HS__O21A_2%A_244_368# N_A_244_368#_M1009_d
+ N_A_244_368#_M1004_d N_A_244_368#_c_154_n N_A_244_368#_M1005_g
+ N_A_244_368#_c_155_n N_A_244_368#_M1007_g N_A_244_368#_c_145_n
+ N_A_244_368#_M1000_g N_A_244_368#_c_146_n N_A_244_368#_c_147_n
+ N_A_244_368#_c_148_n N_A_244_368#_M1008_g N_A_244_368#_c_157_n
+ N_A_244_368#_c_158_n N_A_244_368#_c_159_n N_A_244_368#_c_149_n
+ N_A_244_368#_c_150_n N_A_244_368#_c_151_n N_A_244_368#_c_152_n
+ N_A_244_368#_c_153_n PM_SKY130_FD_SC_HS__O21A_2%A_244_368#
x_PM_SKY130_FD_SC_HS__O21A_2%VPWR N_VPWR_M1001_s N_VPWR_M1003_d N_VPWR_M1007_s
+ N_VPWR_c_220_n N_VPWR_c_221_n N_VPWR_c_222_n N_VPWR_c_223_n N_VPWR_c_224_n
+ VPWR N_VPWR_c_225_n N_VPWR_c_226_n N_VPWR_c_227_n N_VPWR_c_219_n
+ N_VPWR_c_229_n N_VPWR_c_230_n PM_SKY130_FD_SC_HS__O21A_2%VPWR
x_PM_SKY130_FD_SC_HS__O21A_2%X N_X_M1000_d N_X_M1005_d N_X_c_262_n X X X X
+ N_X_c_264_n X PM_SKY130_FD_SC_HS__O21A_2%X
x_PM_SKY130_FD_SC_HS__O21A_2%A_54_74# N_A_54_74#_M1006_s N_A_54_74#_M1002_d
+ N_A_54_74#_c_291_n N_A_54_74#_c_292_n N_A_54_74#_c_297_n N_A_54_74#_c_303_n
+ N_A_54_74#_c_293_n PM_SKY130_FD_SC_HS__O21A_2%A_54_74#
x_PM_SKY130_FD_SC_HS__O21A_2%VGND N_VGND_M1006_d N_VGND_M1000_s N_VGND_M1008_s
+ N_VGND_c_317_n N_VGND_c_318_n N_VGND_c_319_n N_VGND_c_320_n VGND
+ N_VGND_c_321_n N_VGND_c_322_n N_VGND_c_323_n N_VGND_c_324_n N_VGND_c_325_n
+ N_VGND_c_326_n PM_SKY130_FD_SC_HS__O21A_2%VGND
cc_1 VNB N_A1_c_59_n 0.0234618f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=1.22
cc_2 VNB N_A1_c_60_n 0.020755f $X=-0.19 $Y=-0.245 $X2=0.725 $Y2=1.765
cc_3 VNB N_A1_c_61_n 0.0616222f $X=-0.19 $Y=-0.245 $X2=0.625 $Y2=1.385
cc_4 VNB A1 0.0278098f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_5 VNB N_A2_c_82_n 0.0394941f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=1.22
cc_6 VNB N_A2_c_83_n 0.0194558f $X=-0.19 $Y=-0.245 $X2=0.725 $Y2=1.765
cc_7 VNB A2 0.00587703f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.385
cc_8 VNB N_B1_c_109_n 0.0371505f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=1.22
cc_9 VNB N_B1_c_110_n 0.0199025f $X=-0.19 $Y=-0.245 $X2=0.725 $Y2=1.765
cc_10 VNB N_B1_c_111_n 0.00895346f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_244_368#_c_145_n 0.0184836f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.385
cc_12 VNB N_A_244_368#_c_146_n 0.0335612f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_244_368#_c_147_n 0.0688155f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.365
cc_14 VNB N_A_244_368#_c_148_n 0.0199304f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_244_368#_c_149_n 0.00868066f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_244_368#_c_150_n 0.0039379f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_244_368#_c_151_n 0.00271468f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_244_368#_c_152_n 0.00201793f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_244_368#_c_153_n 0.00452572f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_VPWR_c_219_n 0.163682f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB X 0.0162439f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.385
cc_22 VNB N_A_54_74#_c_291_n 0.0071683f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.385
cc_23 VNB N_A_54_74#_c_292_n 0.0222165f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_24 VNB N_A_54_74#_c_293_n 0.00286839f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.385
cc_25 VNB N_VGND_c_317_n 0.00811421f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_VGND_c_318_n 0.0160569f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_VGND_c_319_n 0.010678f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_320_n 0.0505973f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.365
cc_29 VNB N_VGND_c_321_n 0.0232388f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_322_n 0.0333734f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_323_n 0.019013f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_324_n 0.00911377f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_325_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_326_n 0.238533f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VPB N_A1_c_60_n 0.0280881f $X=-0.19 $Y=1.66 $X2=0.725 $Y2=1.765
cc_36 VPB N_A2_c_82_n 0.0240012f $X=-0.19 $Y=1.66 $X2=0.7 $Y2=1.22
cc_37 VPB N_B1_c_109_n 0.0242645f $X=-0.19 $Y=1.66 $X2=0.7 $Y2=1.22
cc_38 VPB N_A_244_368#_c_154_n 0.0164449f $X=-0.19 $Y=1.66 $X2=0.72 $Y2=1.385
cc_39 VPB N_A_244_368#_c_155_n 0.0165253f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.21
cc_40 VPB N_A_244_368#_c_147_n 0.0145303f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=1.365
cc_41 VPB N_A_244_368#_c_157_n 0.00357711f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_42 VPB N_A_244_368#_c_158_n 0.00862872f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_43 VPB N_A_244_368#_c_159_n 0.0100753f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_44 VPB N_A_244_368#_c_151_n 0.00119878f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_45 VPB N_VPWR_c_220_n 0.0613622f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_46 VPB N_VPWR_c_221_n 0.012312f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_47 VPB N_VPWR_c_222_n 0.0469052f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_48 VPB N_VPWR_c_223_n 0.0128037f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_49 VPB N_VPWR_c_224_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_50 VPB N_VPWR_c_225_n 0.0392809f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_51 VPB N_VPWR_c_226_n 0.0186948f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_52 VPB N_VPWR_c_227_n 0.0194863f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_53 VPB N_VPWR_c_219_n 0.110451f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_54 VPB N_VPWR_c_229_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_55 VPB N_VPWR_c_230_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_56 VPB N_X_c_262_n 0.00257348f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.21
cc_57 VPB X 0.00412425f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=1.385
cc_58 VPB N_X_c_264_n 0.0116776f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_59 N_A1_c_60_n N_A2_c_82_n 0.0816953f $X=0.725 $Y=1.765 $X2=-0.19 $Y2=-0.245
cc_60 A1 N_A2_c_82_n 0.00227871f $X=0.635 $Y=1.21 $X2=-0.19 $Y2=-0.245
cc_61 N_A1_c_59_n N_A2_c_83_n 0.0226983f $X=0.7 $Y=1.22 $X2=0 $Y2=0
cc_62 N_A1_c_60_n A2 3.8796e-19 $X=0.725 $Y=1.765 $X2=0 $Y2=0
cc_63 A1 A2 0.0257541f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_64 N_A1_c_60_n N_VPWR_c_220_n 0.0254152f $X=0.725 $Y=1.765 $X2=0 $Y2=0
cc_65 N_A1_c_61_n N_VPWR_c_220_n 0.00660418f $X=0.625 $Y=1.385 $X2=0 $Y2=0
cc_66 A1 N_VPWR_c_220_n 0.0196555f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_67 N_A1_c_60_n N_VPWR_c_225_n 0.00443511f $X=0.725 $Y=1.765 $X2=0 $Y2=0
cc_68 N_A1_c_60_n N_VPWR_c_219_n 0.00460931f $X=0.725 $Y=1.765 $X2=0 $Y2=0
cc_69 N_A1_c_61_n N_A_54_74#_c_291_n 0.00229997f $X=0.625 $Y=1.385 $X2=0 $Y2=0
cc_70 A1 N_A_54_74#_c_291_n 0.0283136f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_71 N_A1_c_59_n N_A_54_74#_c_292_n 0.00977947f $X=0.7 $Y=1.22 $X2=0 $Y2=0
cc_72 N_A1_c_59_n N_A_54_74#_c_297_n 0.0140987f $X=0.7 $Y=1.22 $X2=0 $Y2=0
cc_73 A1 N_A_54_74#_c_297_n 0.0153682f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_74 N_A1_c_59_n N_VGND_c_317_n 0.0138709f $X=0.7 $Y=1.22 $X2=0 $Y2=0
cc_75 N_A1_c_59_n N_VGND_c_321_n 0.00383152f $X=0.7 $Y=1.22 $X2=0 $Y2=0
cc_76 N_A1_c_59_n N_VGND_c_326_n 0.00388149f $X=0.7 $Y=1.22 $X2=0 $Y2=0
cc_77 N_A2_c_82_n N_B1_c_109_n 0.0407612f $X=1.145 $Y=1.765 $X2=-0.19 $Y2=-0.245
cc_78 A2 N_B1_c_109_n 3.71725e-19 $X=1.115 $Y=1.21 $X2=-0.19 $Y2=-0.245
cc_79 N_A2_c_83_n N_B1_c_110_n 0.0103208f $X=1.31 $Y=1.22 $X2=0 $Y2=0
cc_80 N_A2_c_83_n N_B1_c_111_n 0.00227475f $X=1.31 $Y=1.22 $X2=0 $Y2=0
cc_81 A2 N_B1_c_111_n 0.0283697f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_82 N_A2_c_82_n N_A_244_368#_c_157_n 0.0141861f $X=1.145 $Y=1.765 $X2=0 $Y2=0
cc_83 N_A2_c_82_n N_A_244_368#_c_159_n 0.00476672f $X=1.145 $Y=1.765 $X2=0 $Y2=0
cc_84 A2 N_A_244_368#_c_159_n 0.00503923f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_85 N_A2_c_82_n N_VPWR_c_220_n 0.00367695f $X=1.145 $Y=1.765 $X2=0 $Y2=0
cc_86 N_A2_c_82_n N_VPWR_c_225_n 0.0049405f $X=1.145 $Y=1.765 $X2=0 $Y2=0
cc_87 N_A2_c_82_n N_VPWR_c_219_n 0.00508379f $X=1.145 $Y=1.765 $X2=0 $Y2=0
cc_88 N_A2_c_82_n N_A_54_74#_c_297_n 9.99496e-19 $X=1.145 $Y=1.765 $X2=0 $Y2=0
cc_89 N_A2_c_83_n N_A_54_74#_c_297_n 0.0106434f $X=1.31 $Y=1.22 $X2=0 $Y2=0
cc_90 A2 N_A_54_74#_c_297_n 0.0228656f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_91 N_A2_c_83_n N_A_54_74#_c_293_n 4.10343e-19 $X=1.31 $Y=1.22 $X2=0 $Y2=0
cc_92 N_A2_c_83_n N_VGND_c_317_n 0.00532072f $X=1.31 $Y=1.22 $X2=0 $Y2=0
cc_93 N_A2_c_83_n N_VGND_c_322_n 0.00460063f $X=1.31 $Y=1.22 $X2=0 $Y2=0
cc_94 N_A2_c_83_n N_VGND_c_326_n 0.00464404f $X=1.31 $Y=1.22 $X2=0 $Y2=0
cc_95 N_B1_c_109_n N_A_244_368#_c_154_n 0.0167757f $X=1.715 $Y=1.765 $X2=0 $Y2=0
cc_96 N_B1_c_109_n N_A_244_368#_c_147_n 0.0141471f $X=1.715 $Y=1.765 $X2=0 $Y2=0
cc_97 N_B1_c_111_n N_A_244_368#_c_147_n 3.0788e-19 $X=1.79 $Y=1.385 $X2=0 $Y2=0
cc_98 N_B1_c_109_n N_A_244_368#_c_157_n 0.0145853f $X=1.715 $Y=1.765 $X2=0 $Y2=0
cc_99 N_B1_c_109_n N_A_244_368#_c_158_n 0.0168786f $X=1.715 $Y=1.765 $X2=0 $Y2=0
cc_100 N_B1_c_111_n N_A_244_368#_c_158_n 0.0221503f $X=1.79 $Y=1.385 $X2=0 $Y2=0
cc_101 N_B1_c_109_n N_A_244_368#_c_159_n 0.00266381f $X=1.715 $Y=1.765 $X2=0
+ $Y2=0
cc_102 N_B1_c_111_n N_A_244_368#_c_159_n 0.00776619f $X=1.79 $Y=1.385 $X2=0
+ $Y2=0
cc_103 N_B1_c_110_n N_A_244_368#_c_149_n 6.80643e-19 $X=1.785 $Y=1.22 $X2=0
+ $Y2=0
cc_104 N_B1_c_110_n N_A_244_368#_c_150_n 0.00502808f $X=1.785 $Y=1.22 $X2=0
+ $Y2=0
cc_105 N_B1_c_111_n N_A_244_368#_c_150_n 0.00314775f $X=1.79 $Y=1.385 $X2=0
+ $Y2=0
cc_106 N_B1_c_109_n N_A_244_368#_c_151_n 0.00325044f $X=1.715 $Y=1.765 $X2=0
+ $Y2=0
cc_107 N_B1_c_109_n N_A_244_368#_c_152_n 3.15972e-19 $X=1.715 $Y=1.765 $X2=0
+ $Y2=0
cc_108 N_B1_c_111_n N_A_244_368#_c_152_n 0.00378611f $X=1.79 $Y=1.385 $X2=0
+ $Y2=0
cc_109 N_B1_c_109_n N_A_244_368#_c_153_n 0.00131824f $X=1.715 $Y=1.765 $X2=0
+ $Y2=0
cc_110 N_B1_c_111_n N_A_244_368#_c_153_n 0.0275093f $X=1.79 $Y=1.385 $X2=0 $Y2=0
cc_111 N_B1_c_109_n N_VPWR_c_221_n 0.0109634f $X=1.715 $Y=1.765 $X2=0 $Y2=0
cc_112 N_B1_c_109_n N_VPWR_c_225_n 0.00481995f $X=1.715 $Y=1.765 $X2=0 $Y2=0
cc_113 N_B1_c_109_n N_VPWR_c_219_n 0.00508379f $X=1.715 $Y=1.765 $X2=0 $Y2=0
cc_114 N_B1_c_109_n N_X_c_262_n 8.49317e-19 $X=1.715 $Y=1.765 $X2=0 $Y2=0
cc_115 N_B1_c_109_n N_A_54_74#_c_303_n 4.36459e-19 $X=1.715 $Y=1.765 $X2=0 $Y2=0
cc_116 N_B1_c_110_n N_A_54_74#_c_303_n 0.00215143f $X=1.785 $Y=1.22 $X2=0 $Y2=0
cc_117 N_B1_c_111_n N_A_54_74#_c_303_n 0.012077f $X=1.79 $Y=1.385 $X2=0 $Y2=0
cc_118 N_B1_c_110_n N_A_54_74#_c_293_n 0.00622341f $X=1.785 $Y=1.22 $X2=0 $Y2=0
cc_119 N_B1_c_110_n N_VGND_c_318_n 0.00313679f $X=1.785 $Y=1.22 $X2=0 $Y2=0
cc_120 N_B1_c_110_n N_VGND_c_322_n 0.00434054f $X=1.785 $Y=1.22 $X2=0 $Y2=0
cc_121 N_B1_c_110_n N_VGND_c_326_n 0.0082661f $X=1.785 $Y=1.22 $X2=0 $Y2=0
cc_122 N_A_244_368#_c_158_n N_VPWR_M1003_d 0.00859937f $X=2.125 $Y=1.805 $X2=0
+ $Y2=0
cc_123 N_A_244_368#_c_157_n N_VPWR_c_220_n 0.0255995f $X=1.49 $Y=1.985 $X2=0
+ $Y2=0
cc_124 N_A_244_368#_c_159_n N_VPWR_c_220_n 0.00199817f $X=1.655 $Y=1.805 $X2=0
+ $Y2=0
cc_125 N_A_244_368#_c_154_n N_VPWR_c_221_n 0.0104597f $X=2.405 $Y=1.765 $X2=0
+ $Y2=0
cc_126 N_A_244_368#_c_157_n N_VPWR_c_221_n 0.0391828f $X=1.49 $Y=1.985 $X2=0
+ $Y2=0
cc_127 N_A_244_368#_c_158_n N_VPWR_c_221_n 0.0255961f $X=2.125 $Y=1.805 $X2=0
+ $Y2=0
cc_128 N_A_244_368#_c_155_n N_VPWR_c_222_n 0.0213847f $X=2.855 $Y=1.765 $X2=0
+ $Y2=0
cc_129 N_A_244_368#_c_157_n N_VPWR_c_225_n 0.0097982f $X=1.49 $Y=1.985 $X2=0
+ $Y2=0
cc_130 N_A_244_368#_c_154_n N_VPWR_c_226_n 0.00445602f $X=2.405 $Y=1.765 $X2=0
+ $Y2=0
cc_131 N_A_244_368#_c_155_n N_VPWR_c_226_n 0.00445602f $X=2.855 $Y=1.765 $X2=0
+ $Y2=0
cc_132 N_A_244_368#_c_154_n N_VPWR_c_219_n 0.00861719f $X=2.405 $Y=1.765 $X2=0
+ $Y2=0
cc_133 N_A_244_368#_c_155_n N_VPWR_c_219_n 0.00861719f $X=2.855 $Y=1.765 $X2=0
+ $Y2=0
cc_134 N_A_244_368#_c_157_n N_VPWR_c_219_n 0.0111907f $X=1.49 $Y=1.985 $X2=0
+ $Y2=0
cc_135 N_A_244_368#_c_154_n N_X_c_262_n 0.0137147f $X=2.405 $Y=1.765 $X2=0 $Y2=0
cc_136 N_A_244_368#_c_155_n N_X_c_262_n 0.0174943f $X=2.855 $Y=1.765 $X2=0 $Y2=0
cc_137 N_A_244_368#_c_145_n X 0.0137211f $X=2.915 $Y=1.22 $X2=0 $Y2=0
cc_138 N_A_244_368#_c_146_n X 0.0191488f $X=3.27 $Y=1.295 $X2=0 $Y2=0
cc_139 N_A_244_368#_c_147_n X 0.0155597f $X=2.99 $Y=1.295 $X2=0 $Y2=0
cc_140 N_A_244_368#_c_148_n X 0.0148558f $X=3.345 $Y=1.22 $X2=0 $Y2=0
cc_141 N_A_244_368#_c_150_n X 0.00446539f $X=2.21 $Y=1.22 $X2=0 $Y2=0
cc_142 N_A_244_368#_c_151_n X 0.00504242f $X=2.21 $Y=1.72 $X2=0 $Y2=0
cc_143 N_A_244_368#_c_153_n X 0.0161585f $X=2.48 $Y=1.385 $X2=0 $Y2=0
cc_144 N_A_244_368#_c_154_n N_X_c_264_n 0.00217371f $X=2.405 $Y=1.765 $X2=0
+ $Y2=0
cc_145 N_A_244_368#_c_155_n N_X_c_264_n 0.0113027f $X=2.855 $Y=1.765 $X2=0 $Y2=0
cc_146 N_A_244_368#_c_147_n N_X_c_264_n 0.0156994f $X=2.99 $Y=1.295 $X2=0 $Y2=0
cc_147 N_A_244_368#_c_158_n N_X_c_264_n 0.0125926f $X=2.125 $Y=1.805 $X2=0 $Y2=0
cc_148 N_A_244_368#_c_153_n N_X_c_264_n 0.0134173f $X=2.48 $Y=1.385 $X2=0 $Y2=0
cc_149 N_A_244_368#_c_149_n N_A_54_74#_c_293_n 0.0199611f $X=2 $Y=0.505 $X2=0
+ $Y2=0
cc_150 N_A_244_368#_c_145_n N_VGND_c_318_n 0.0182605f $X=2.915 $Y=1.22 $X2=0
+ $Y2=0
cc_151 N_A_244_368#_c_147_n N_VGND_c_318_n 0.00945103f $X=2.99 $Y=1.295 $X2=0
+ $Y2=0
cc_152 N_A_244_368#_c_149_n N_VGND_c_318_n 0.0595951f $X=2 $Y=0.505 $X2=0 $Y2=0
cc_153 N_A_244_368#_c_153_n N_VGND_c_318_n 0.0148152f $X=2.48 $Y=1.385 $X2=0
+ $Y2=0
cc_154 N_A_244_368#_c_148_n N_VGND_c_320_n 0.00647412f $X=3.345 $Y=1.22 $X2=0
+ $Y2=0
cc_155 N_A_244_368#_c_149_n N_VGND_c_322_n 0.0180247f $X=2 $Y=0.505 $X2=0 $Y2=0
cc_156 N_A_244_368#_c_145_n N_VGND_c_323_n 0.00434272f $X=2.915 $Y=1.22 $X2=0
+ $Y2=0
cc_157 N_A_244_368#_c_148_n N_VGND_c_323_n 0.00434272f $X=3.345 $Y=1.22 $X2=0
+ $Y2=0
cc_158 N_A_244_368#_c_145_n N_VGND_c_326_n 0.00825059f $X=2.915 $Y=1.22 $X2=0
+ $Y2=0
cc_159 N_A_244_368#_c_148_n N_VGND_c_326_n 0.00823942f $X=3.345 $Y=1.22 $X2=0
+ $Y2=0
cc_160 N_A_244_368#_c_149_n N_VGND_c_326_n 0.0144116f $X=2 $Y=0.505 $X2=0 $Y2=0
cc_161 N_VPWR_c_221_n N_X_c_262_n 0.0353111f $X=2.13 $Y=2.145 $X2=0 $Y2=0
cc_162 N_VPWR_c_222_n N_X_c_262_n 0.0353111f $X=3.13 $Y=2.225 $X2=0 $Y2=0
cc_163 N_VPWR_c_226_n N_X_c_262_n 0.014552f $X=2.965 $Y=3.33 $X2=0 $Y2=0
cc_164 N_VPWR_c_219_n N_X_c_262_n 0.0119791f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_165 N_VPWR_M1007_s N_X_c_264_n 0.00346832f $X=2.93 $Y=1.84 $X2=0 $Y2=0
cc_166 N_VPWR_c_222_n N_X_c_264_n 0.025036f $X=3.13 $Y=2.225 $X2=0 $Y2=0
cc_167 X N_VGND_c_318_n 0.0270562f $X=3.035 $Y=0.47 $X2=0 $Y2=0
cc_168 N_X_c_264_n N_VGND_c_318_n 0.00421771f $X=3.13 $Y=1.72 $X2=0 $Y2=0
cc_169 X N_VGND_c_320_n 0.0294122f $X=3.035 $Y=0.47 $X2=0 $Y2=0
cc_170 X N_VGND_c_323_n 0.0144922f $X=3.035 $Y=0.47 $X2=0 $Y2=0
cc_171 X N_VGND_c_326_n 0.0118826f $X=3.035 $Y=0.47 $X2=0 $Y2=0
cc_172 N_A_54_74#_c_297_n N_VGND_M1006_d 0.0146092f $X=1.405 $Y=0.925 $X2=-0.19
+ $Y2=-0.245
cc_173 N_A_54_74#_c_292_n N_VGND_c_317_n 0.0115542f $X=0.415 $Y=0.505 $X2=0
+ $Y2=0
cc_174 N_A_54_74#_c_297_n N_VGND_c_317_n 0.0219781f $X=1.405 $Y=0.925 $X2=0
+ $Y2=0
cc_175 N_A_54_74#_c_293_n N_VGND_c_317_n 0.00248533f $X=1.57 $Y=0.505 $X2=0
+ $Y2=0
cc_176 N_A_54_74#_c_292_n N_VGND_c_321_n 0.0152302f $X=0.415 $Y=0.505 $X2=0
+ $Y2=0
cc_177 N_A_54_74#_c_293_n N_VGND_c_322_n 0.0151574f $X=1.57 $Y=0.505 $X2=0 $Y2=0
cc_178 N_A_54_74#_c_292_n N_VGND_c_326_n 0.0121804f $X=0.415 $Y=0.505 $X2=0
+ $Y2=0
cc_179 N_A_54_74#_c_297_n N_VGND_c_326_n 0.0115606f $X=1.405 $Y=0.925 $X2=0
+ $Y2=0
cc_180 N_A_54_74#_c_293_n N_VGND_c_326_n 0.0120652f $X=1.57 $Y=0.505 $X2=0 $Y2=0
