* File: sky130_fd_sc_hs__sedfxtp_4.pxi.spice
* Created: Tue Sep  1 20:24:46 2020
* 
x_PM_SKY130_FD_SC_HS__SEDFXTP_4%D N_D_c_351_n N_D_c_352_n N_D_M1018_g
+ N_D_M1002_g D D N_D_c_348_n N_D_c_349_n N_D_c_350_n N_D_c_355_n
+ PM_SKY130_FD_SC_HS__SEDFXTP_4%D
x_PM_SKY130_FD_SC_HS__SEDFXTP_4%A_177_290# N_A_177_290#_M1008_s
+ N_A_177_290#_M1001_s N_A_177_290#_c_397_n N_A_177_290#_M1037_g
+ N_A_177_290#_M1038_g N_A_177_290#_c_398_n N_A_177_290#_c_390_n
+ N_A_177_290#_c_391_n N_A_177_290#_c_392_n N_A_177_290#_c_393_n
+ N_A_177_290#_c_400_n N_A_177_290#_c_401_n N_A_177_290#_c_394_n
+ N_A_177_290#_c_402_n N_A_177_290#_c_403_n N_A_177_290#_c_395_n
+ N_A_177_290#_c_396_n PM_SKY130_FD_SC_HS__SEDFXTP_4%A_177_290#
x_PM_SKY130_FD_SC_HS__SEDFXTP_4%DE N_DE_M1034_g N_DE_c_498_n N_DE_c_499_n
+ N_DE_c_500_n N_DE_c_506_n N_DE_c_507_n N_DE_c_501_n N_DE_M1008_g N_DE_c_508_n
+ N_DE_M1001_g N_DE_c_509_n N_DE_c_510_n N_DE_M1030_g N_DE_c_502_n N_DE_c_511_n
+ DE N_DE_c_503_n N_DE_c_512_n N_DE_c_504_n PM_SKY130_FD_SC_HS__SEDFXTP_4%DE
x_PM_SKY130_FD_SC_HS__SEDFXTP_4%A_545_87# N_A_545_87#_M1021_d
+ N_A_545_87#_M1020_d N_A_545_87#_M1023_g N_A_545_87#_c_601_n
+ N_A_545_87#_c_602_n N_A_545_87#_M1015_g N_A_545_87#_c_591_n
+ N_A_545_87#_M1017_g N_A_545_87#_c_592_n N_A_545_87#_c_593_n
+ N_A_545_87#_c_603_n N_A_545_87#_M1035_g N_A_545_87#_c_594_n
+ N_A_545_87#_c_605_n N_A_545_87#_c_606_n N_A_545_87#_c_595_n
+ N_A_545_87#_c_607_n N_A_545_87#_c_608_n N_A_545_87#_c_596_n
+ N_A_545_87#_c_609_n N_A_545_87#_c_610_n N_A_545_87#_c_597_n
+ N_A_545_87#_c_598_n N_A_545_87#_c_613_n N_A_545_87#_c_614_n
+ N_A_545_87#_c_599_n N_A_545_87#_c_600_n
+ PM_SKY130_FD_SC_HS__SEDFXTP_4%A_545_87#
x_PM_SKY130_FD_SC_HS__SEDFXTP_4%A_631_87# N_A_631_87#_M1045_s
+ N_A_631_87#_M1044_s N_A_631_87#_c_831_n N_A_631_87#_M1024_g
+ N_A_631_87#_c_832_n N_A_631_87#_c_833_n N_A_631_87#_c_842_n
+ N_A_631_87#_M1000_g N_A_631_87#_c_834_n N_A_631_87#_c_843_n
+ N_A_631_87#_c_835_n N_A_631_87#_c_836_n N_A_631_87#_c_837_n
+ N_A_631_87#_c_838_n N_A_631_87#_c_846_n N_A_631_87#_c_847_n
+ N_A_631_87#_c_839_n N_A_631_87#_c_840_n N_A_631_87#_c_841_n
+ N_A_631_87#_c_849_n N_A_631_87#_c_850_n
+ PM_SKY130_FD_SC_HS__SEDFXTP_4%A_631_87#
x_PM_SKY130_FD_SC_HS__SEDFXTP_4%SCD N_SCD_M1011_g N_SCD_c_949_n N_SCD_c_950_n
+ N_SCD_M1033_g SCD N_SCD_c_948_n PM_SKY130_FD_SC_HS__SEDFXTP_4%SCD
x_PM_SKY130_FD_SC_HS__SEDFXTP_4%SCE N_SCE_c_999_n N_SCE_M1019_g N_SCE_c_1000_n
+ N_SCE_c_1001_n N_SCE_c_992_n N_SCE_c_1003_n N_SCE_M1044_g N_SCE_M1045_g
+ N_SCE_c_994_n N_SCE_c_995_n N_SCE_M1003_g SCE N_SCE_c_998_n
+ PM_SKY130_FD_SC_HS__SEDFXTP_4%SCE
x_PM_SKY130_FD_SC_HS__SEDFXTP_4%CLK N_CLK_c_1080_n N_CLK_M1026_g N_CLK_c_1081_n
+ N_CLK_M1025_g CLK PM_SKY130_FD_SC_HS__SEDFXTP_4%CLK
x_PM_SKY130_FD_SC_HS__SEDFXTP_4%A_1510_74# N_A_1510_74#_M1013_d
+ N_A_1510_74#_M1029_d N_A_1510_74#_c_1140_n N_A_1510_74#_M1005_g
+ N_A_1510_74#_c_1115_n N_A_1510_74#_M1036_g N_A_1510_74#_M1031_g
+ N_A_1510_74#_c_1117_n N_A_1510_74#_c_1142_n N_A_1510_74#_M1014_g
+ N_A_1510_74#_c_1118_n N_A_1510_74#_c_1119_n N_A_1510_74#_c_1120_n
+ N_A_1510_74#_c_1143_n N_A_1510_74#_c_1121_n N_A_1510_74#_c_1122_n
+ N_A_1510_74#_c_1123_n N_A_1510_74#_c_1124_n N_A_1510_74#_c_1221_p
+ N_A_1510_74#_c_1125_n N_A_1510_74#_c_1126_n N_A_1510_74#_c_1127_n
+ N_A_1510_74#_c_1128_n N_A_1510_74#_c_1129_n N_A_1510_74#_c_1130_n
+ N_A_1510_74#_c_1131_n N_A_1510_74#_c_1132_n N_A_1510_74#_c_1133_n
+ N_A_1510_74#_c_1134_n N_A_1510_74#_c_1147_n N_A_1510_74#_c_1148_n
+ N_A_1510_74#_c_1135_n N_A_1510_74#_c_1136_n N_A_1510_74#_c_1137_n
+ N_A_1510_74#_c_1138_n N_A_1510_74#_c_1139_n
+ PM_SKY130_FD_SC_HS__SEDFXTP_4%A_1510_74#
x_PM_SKY130_FD_SC_HS__SEDFXTP_4%A_1313_74# N_A_1313_74#_M1026_d
+ N_A_1313_74#_M1025_d N_A_1313_74#_M1013_g N_A_1313_74#_c_1343_n
+ N_A_1313_74#_c_1358_n N_A_1313_74#_M1029_g N_A_1313_74#_c_1344_n
+ N_A_1313_74#_M1040_g N_A_1313_74#_c_1346_n N_A_1313_74#_c_1361_n
+ N_A_1313_74#_c_1362_n N_A_1313_74#_M1010_g N_A_1313_74#_c_1347_n
+ N_A_1313_74#_M1006_g N_A_1313_74#_M1016_g N_A_1313_74#_c_1349_n
+ N_A_1313_74#_c_1350_n N_A_1313_74#_c_1351_n N_A_1313_74#_c_1366_n
+ N_A_1313_74#_c_1352_n N_A_1313_74#_c_1353_n N_A_1313_74#_c_1354_n
+ N_A_1313_74#_c_1368_n N_A_1313_74#_c_1369_n N_A_1313_74#_c_1370_n
+ N_A_1313_74#_c_1355_n N_A_1313_74#_c_1356_n
+ PM_SKY130_FD_SC_HS__SEDFXTP_4%A_1313_74#
x_PM_SKY130_FD_SC_HS__SEDFXTP_4%A_1943_53# N_A_1943_53#_M1046_d
+ N_A_1943_53#_M1043_d N_A_1943_53#_M1032_g N_A_1943_53#_c_1534_n
+ N_A_1943_53#_c_1546_n N_A_1943_53#_M1007_g N_A_1943_53#_c_1535_n
+ N_A_1943_53#_c_1548_n N_A_1943_53#_M1027_g N_A_1943_53#_c_1536_n
+ N_A_1943_53#_M1047_g N_A_1943_53#_c_1537_n N_A_1943_53#_c_1549_n
+ N_A_1943_53#_c_1538_n N_A_1943_53#_c_1539_n N_A_1943_53#_c_1540_n
+ N_A_1943_53#_c_1541_n N_A_1943_53#_c_1542_n N_A_1943_53#_c_1543_n
+ N_A_1943_53#_c_1544_n PM_SKY130_FD_SC_HS__SEDFXTP_4%A_1943_53#
x_PM_SKY130_FD_SC_HS__SEDFXTP_4%A_1756_97# N_A_1756_97#_M1040_d
+ N_A_1756_97#_M1005_d N_A_1756_97#_c_1639_n N_A_1756_97#_M1043_g
+ N_A_1756_97#_M1046_g N_A_1756_97#_c_1641_n N_A_1756_97#_c_1645_n
+ N_A_1756_97#_c_1646_n N_A_1756_97#_c_1647_n N_A_1756_97#_c_1642_n
+ N_A_1756_97#_c_1643_n PM_SKY130_FD_SC_HS__SEDFXTP_4%A_1756_97#
x_PM_SKY130_FD_SC_HS__SEDFXTP_4%A_2403_74# N_A_2403_74#_M1031_d
+ N_A_2403_74#_M1006_d N_A_2403_74#_c_1727_n N_A_2403_74#_M1021_g
+ N_A_2403_74#_c_1741_n N_A_2403_74#_c_1742_n N_A_2403_74#_M1020_g
+ N_A_2403_74#_c_1729_n N_A_2403_74#_c_1730_n N_A_2403_74#_M1022_g
+ N_A_2403_74#_c_1744_n N_A_2403_74#_M1004_g N_A_2403_74#_c_1731_n
+ N_A_2403_74#_M1039_g N_A_2403_74#_c_1745_n N_A_2403_74#_M1009_g
+ N_A_2403_74#_c_1746_n N_A_2403_74#_M1012_g N_A_2403_74#_c_1732_n
+ N_A_2403_74#_M1041_g N_A_2403_74#_c_1747_n N_A_2403_74#_M1028_g
+ N_A_2403_74#_c_1733_n N_A_2403_74#_M1042_g N_A_2403_74#_c_1734_n
+ N_A_2403_74#_c_1735_n N_A_2403_74#_c_1736_n N_A_2403_74#_c_1737_n
+ N_A_2403_74#_c_1749_n N_A_2403_74#_c_1750_n N_A_2403_74#_c_1751_n
+ N_A_2403_74#_c_1752_n N_A_2403_74#_c_1738_n N_A_2403_74#_c_1739_n
+ N_A_2403_74#_c_1740_n PM_SKY130_FD_SC_HS__SEDFXTP_4%A_2403_74#
x_PM_SKY130_FD_SC_HS__SEDFXTP_4%A_37_464# N_A_37_464#_M1002_s
+ N_A_37_464#_M1023_d N_A_37_464#_M1018_s N_A_37_464#_M1015_d
+ N_A_37_464#_c_1912_n N_A_37_464#_c_1918_n N_A_37_464#_c_1919_n
+ N_A_37_464#_c_1920_n N_A_37_464#_c_1921_n N_A_37_464#_c_1922_n
+ N_A_37_464#_c_1954_n N_A_37_464#_c_1923_n N_A_37_464#_c_1924_n
+ N_A_37_464#_c_1913_n N_A_37_464#_c_1925_n N_A_37_464#_c_1914_n
+ N_A_37_464#_c_1915_n N_A_37_464#_c_1927_n N_A_37_464#_c_1916_n
+ N_A_37_464#_c_1928_n PM_SKY130_FD_SC_HS__SEDFXTP_4%A_37_464#
x_PM_SKY130_FD_SC_HS__SEDFXTP_4%VPWR N_VPWR_M1037_d N_VPWR_M1001_d
+ N_VPWR_M1044_d N_VPWR_M1025_s N_VPWR_M1029_s N_VPWR_M1007_d N_VPWR_M1027_s
+ N_VPWR_M1035_d N_VPWR_M1004_d N_VPWR_M1009_d N_VPWR_M1028_d N_VPWR_c_2038_n
+ N_VPWR_c_2039_n N_VPWR_c_2040_n N_VPWR_c_2041_n N_VPWR_c_2042_n
+ N_VPWR_c_2043_n N_VPWR_c_2044_n N_VPWR_c_2045_n N_VPWR_c_2046_n
+ N_VPWR_c_2047_n N_VPWR_c_2048_n N_VPWR_c_2049_n N_VPWR_c_2050_n
+ N_VPWR_c_2051_n N_VPWR_c_2052_n VPWR N_VPWR_c_2053_n N_VPWR_c_2054_n
+ N_VPWR_c_2055_n N_VPWR_c_2056_n N_VPWR_c_2057_n N_VPWR_c_2058_n
+ N_VPWR_c_2059_n N_VPWR_c_2060_n N_VPWR_c_2061_n N_VPWR_c_2062_n
+ N_VPWR_c_2063_n N_VPWR_c_2064_n N_VPWR_c_2065_n N_VPWR_c_2066_n
+ N_VPWR_c_2067_n N_VPWR_c_2068_n N_VPWR_c_2069_n N_VPWR_c_2070_n
+ N_VPWR_c_2037_n PM_SKY130_FD_SC_HS__SEDFXTP_4%VPWR
x_PM_SKY130_FD_SC_HS__SEDFXTP_4%A_661_113# N_A_661_113#_M1024_d
+ N_A_661_113#_M1003_d N_A_661_113#_M1040_s N_A_661_113#_M1019_d
+ N_A_661_113#_M1000_d N_A_661_113#_M1005_s N_A_661_113#_c_2241_n
+ N_A_661_113#_c_2309_n N_A_661_113#_c_2242_n N_A_661_113#_c_2253_n
+ N_A_661_113#_c_2269_n N_A_661_113#_c_2243_n N_A_661_113#_c_2233_n
+ N_A_661_113#_c_2234_n N_A_661_113#_c_2245_n N_A_661_113#_c_2246_n
+ N_A_661_113#_c_2235_n N_A_661_113#_c_2236_n N_A_661_113#_c_2247_n
+ N_A_661_113#_c_2237_n N_A_661_113#_c_2238_n N_A_661_113#_c_2239_n
+ N_A_661_113#_c_2240_n N_A_661_113#_c_2249_n N_A_661_113#_c_2250_n
+ N_A_661_113#_c_2251_n N_A_661_113#_c_2398_n
+ PM_SKY130_FD_SC_HS__SEDFXTP_4%A_661_113#
x_PM_SKY130_FD_SC_HS__SEDFXTP_4%Q N_Q_M1022_d N_Q_M1041_d N_Q_M1004_s
+ N_Q_M1012_s N_Q_c_2418_n N_Q_c_2415_n N_Q_c_2419_n N_Q_c_2416_n Q
+ PM_SKY130_FD_SC_HS__SEDFXTP_4%Q
x_PM_SKY130_FD_SC_HS__SEDFXTP_4%VGND N_VGND_M1034_d N_VGND_M1008_d
+ N_VGND_M1045_d N_VGND_M1026_s N_VGND_M1013_s N_VGND_M1032_d N_VGND_M1047_s
+ N_VGND_M1017_d N_VGND_M1022_s N_VGND_M1039_s N_VGND_M1042_s N_VGND_c_2467_n
+ N_VGND_c_2468_n N_VGND_c_2469_n N_VGND_c_2470_n N_VGND_c_2471_n
+ N_VGND_c_2472_n N_VGND_c_2473_n N_VGND_c_2474_n N_VGND_c_2475_n
+ N_VGND_c_2476_n N_VGND_c_2477_n N_VGND_c_2478_n N_VGND_c_2479_n
+ N_VGND_c_2480_n N_VGND_c_2481_n N_VGND_c_2482_n VGND N_VGND_c_2483_n
+ N_VGND_c_2484_n N_VGND_c_2485_n N_VGND_c_2486_n N_VGND_c_2487_n
+ N_VGND_c_2488_n N_VGND_c_2489_n N_VGND_c_2490_n N_VGND_c_2491_n
+ N_VGND_c_2492_n N_VGND_c_2493_n N_VGND_c_2494_n N_VGND_c_2495_n
+ N_VGND_c_2496_n N_VGND_c_2497_n N_VGND_c_2498_n N_VGND_c_2499_n
+ PM_SKY130_FD_SC_HS__SEDFXTP_4%VGND
cc_1 VNB N_D_M1002_g 0.0257827f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=0.58
cc_2 VNB N_D_c_348_n 0.0164802f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=1.145
cc_3 VNB N_D_c_349_n 0.0118303f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=1.145
cc_4 VNB N_D_c_350_n 0.0396651f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=1.825
cc_5 VNB N_A_177_290#_M1038_g 0.0403695f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_6 VNB N_A_177_290#_c_390_n 0.00361826f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=1.145
cc_7 VNB N_A_177_290#_c_391_n 0.0238207f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=1.145
cc_8 VNB N_A_177_290#_c_392_n 0.00900198f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=1.825
cc_9 VNB N_A_177_290#_c_393_n 0.0024367f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=1.825
cc_10 VNB N_A_177_290#_c_394_n 0.00790857f $X=-0.19 $Y=-0.245 $X2=0.625
+ $Y2=1.295
cc_11 VNB N_A_177_290#_c_395_n 0.00328079f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_177_290#_c_396_n 0.0184501f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_DE_M1034_g 0.0296548f $X=-0.19 $Y=-0.245 $X2=0.555 $Y2=2.245
cc_14 VNB N_DE_c_498_n 0.0311116f $X=-0.19 $Y=-0.245 $X2=0.555 $Y2=2.64
cc_15 VNB N_DE_c_499_n 0.00739824f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=0.98
cc_16 VNB N_DE_c_500_n 3.94837e-19 $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=1.145
cc_17 VNB N_DE_c_501_n 0.0158293f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_18 VNB N_DE_c_502_n 0.0297232f $X=-0.19 $Y=-0.245 $X2=0.625 $Y2=1.145
cc_19 VNB N_DE_c_503_n 0.0232037f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_DE_c_504_n 0.0163775f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_545_87#_M1023_g 0.0405741f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_545_87#_c_591_n 0.0186115f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=1.825
cc_23 VNB N_A_545_87#_c_592_n 0.039284f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=1.145
cc_24 VNB N_A_545_87#_c_593_n 0.00644191f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=1.825
cc_25 VNB N_A_545_87#_c_594_n 0.0294864f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_545_87#_c_595_n 0.0109324f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_545_87#_c_596_n 0.0129179f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_545_87#_c_597_n 0.0623893f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_545_87#_c_598_n 0.00229751f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_545_87#_c_599_n 0.0076271f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_545_87#_c_600_n 0.0226673f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_631_87#_c_831_n 0.016594f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=0.58
cc_33 VNB N_A_631_87#_c_832_n 0.039446f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=1.145
cc_34 VNB N_A_631_87#_c_833_n 0.0071047f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=0.98
cc_35 VNB N_A_631_87#_c_834_n 0.00763236f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=1.145
cc_36 VNB N_A_631_87#_c_835_n 0.00555818f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=1.825
cc_37 VNB N_A_631_87#_c_836_n 0.0777051f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=1.825
cc_38 VNB N_A_631_87#_c_837_n 0.00586902f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_631_87#_c_838_n 0.0316144f $X=-0.19 $Y=-0.245 $X2=0.625 $Y2=1.665
cc_40 VNB N_A_631_87#_c_839_n 0.0026099f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_631_87#_c_840_n 0.0279495f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_631_87#_c_841_n 0.00583512f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_SCD_M1011_g 0.028991f $X=-0.19 $Y=-0.245 $X2=0.555 $Y2=2.245
cc_44 VNB SCD 0.0143176f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=1.145
cc_45 VNB N_SCD_c_948_n 0.020908f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_46 VNB N_SCE_c_992_n 0.00813877f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=0.58
cc_47 VNB N_SCE_M1045_g 0.0292433f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_SCE_c_994_n 0.0563111f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=1.825
cc_49 VNB N_SCE_c_995_n 0.0126405f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=1.145
cc_50 VNB N_SCE_M1003_g 0.0390656f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=1.825
cc_51 VNB SCE 0.00220979f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=1.825
cc_52 VNB N_SCE_c_998_n 0.0323386f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_CLK_c_1080_n 0.021307f $X=-0.19 $Y=-0.245 $X2=0.555 $Y2=1.99
cc_54 VNB N_CLK_c_1081_n 0.0439821f $X=-0.19 $Y=-0.245 $X2=0.555 $Y2=2.64
cc_55 VNB CLK 0.0118416f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=0.58
cc_56 VNB N_A_1510_74#_c_1115_n 0.0178999f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=1.145
cc_57 VNB N_A_1510_74#_M1031_g 0.035059f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_A_1510_74#_c_1117_n 0.00362656f $X=-0.19 $Y=-0.245 $X2=0.51
+ $Y2=1.145
cc_59 VNB N_A_1510_74#_c_1118_n 0.0111034f $X=-0.19 $Y=-0.245 $X2=0.625
+ $Y2=1.145
cc_60 VNB N_A_1510_74#_c_1119_n 0.0239053f $X=-0.19 $Y=-0.245 $X2=0.625
+ $Y2=1.295
cc_61 VNB N_A_1510_74#_c_1120_n 0.00362036f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_A_1510_74#_c_1121_n 0.00727581f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_A_1510_74#_c_1122_n 0.00977192f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_A_1510_74#_c_1123_n 4.71639e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_A_1510_74#_c_1124_n 0.0122213f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_A_1510_74#_c_1125_n 0.0120634f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_A_1510_74#_c_1126_n 0.00223246f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_A_1510_74#_c_1127_n 0.00973757f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_A_1510_74#_c_1128_n 0.00548977f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_A_1510_74#_c_1129_n 0.00370687f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_A_1510_74#_c_1130_n 0.00285285f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_A_1510_74#_c_1131_n 7.17725e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_A_1510_74#_c_1132_n 0.0173419f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_A_1510_74#_c_1133_n 0.011428f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_A_1510_74#_c_1134_n 0.00123754f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_A_1510_74#_c_1135_n 0.0029202f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_A_1510_74#_c_1136_n 0.0382543f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_A_1510_74#_c_1137_n 0.0015589f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VNB N_A_1510_74#_c_1138_n 0.00361396f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_A_1510_74#_c_1139_n 0.0309263f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_81 VNB N_A_1313_74#_M1013_g 0.0477158f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_82 VNB N_A_1313_74#_c_1343_n 0.0102894f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=0.98
cc_83 VNB N_A_1313_74#_c_1344_n 0.0168013f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=1.825
cc_84 VNB N_A_1313_74#_M1040_g 0.0593878f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=1.825
cc_85 VNB N_A_1313_74#_c_1346_n 0.0197045f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=1.825
cc_86 VNB N_A_1313_74#_c_1347_n 0.0156746f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_87 VNB N_A_1313_74#_M1016_g 0.0508999f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_88 VNB N_A_1313_74#_c_1349_n 0.00496867f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_89 VNB N_A_1313_74#_c_1350_n 7.16371e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_90 VNB N_A_1313_74#_c_1351_n 0.00811038f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_91 VNB N_A_1313_74#_c_1352_n 0.00802109f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_92 VNB N_A_1313_74#_c_1353_n 3.70884e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_93 VNB N_A_1313_74#_c_1354_n 0.00455076f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_94 VNB N_A_1313_74#_c_1355_n 0.00283324f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_95 VNB N_A_1313_74#_c_1356_n 0.00926081f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_96 VNB N_A_1943_53#_M1032_g 0.0303996f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_97 VNB N_A_1943_53#_c_1534_n 0.0133486f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_98 VNB N_A_1943_53#_c_1535_n 0.00784676f $X=-0.19 $Y=-0.245 $X2=0.51
+ $Y2=1.145
cc_99 VNB N_A_1943_53#_c_1536_n 0.0200998f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=1.825
cc_100 VNB N_A_1943_53#_c_1537_n 0.00793133f $X=-0.19 $Y=-0.245 $X2=0.625
+ $Y2=1.145
cc_101 VNB N_A_1943_53#_c_1538_n 0.00534086f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_102 VNB N_A_1943_53#_c_1539_n 0.0029595f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_103 VNB N_A_1943_53#_c_1540_n 0.0120372f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_104 VNB N_A_1943_53#_c_1541_n 0.00726422f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_105 VNB N_A_1943_53#_c_1542_n 0.0353896f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_106 VNB N_A_1943_53#_c_1543_n 0.00672473f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_107 VNB N_A_1943_53#_c_1544_n 0.0555109f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_108 VNB N_A_1756_97#_c_1639_n 0.0170806f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=0.58
cc_109 VNB N_A_1756_97#_M1046_g 0.0405995f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_110 VNB N_A_1756_97#_c_1641_n 0.0210446f $X=-0.19 $Y=-0.245 $X2=0.51
+ $Y2=1.825
cc_111 VNB N_A_1756_97#_c_1642_n 0.00177868f $X=-0.19 $Y=-0.245 $X2=0.625
+ $Y2=1.825
cc_112 VNB N_A_1756_97#_c_1643_n 0.00410966f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_113 VNB N_A_2403_74#_c_1727_n 0.0173241f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=0.58
cc_114 VNB N_A_2403_74#_M1021_g 0.0269829f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=0.98
cc_115 VNB N_A_2403_74#_c_1729_n 0.0423887f $X=-0.19 $Y=-0.245 $X2=0.51
+ $Y2=1.145
cc_116 VNB N_A_2403_74#_c_1730_n 0.0169461f $X=-0.19 $Y=-0.245 $X2=0.51
+ $Y2=1.825
cc_117 VNB N_A_2403_74#_c_1731_n 0.0145959f $X=-0.19 $Y=-0.245 $X2=0.625
+ $Y2=1.295
cc_118 VNB N_A_2403_74#_c_1732_n 0.0142433f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_119 VNB N_A_2403_74#_c_1733_n 0.0168044f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_120 VNB N_A_2403_74#_c_1734_n 0.0612794f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_121 VNB N_A_2403_74#_c_1735_n 0.00286116f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_122 VNB N_A_2403_74#_c_1736_n 0.0225925f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_123 VNB N_A_2403_74#_c_1737_n 0.0025106f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_124 VNB N_A_2403_74#_c_1738_n 0.010486f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_125 VNB N_A_2403_74#_c_1739_n 0.0183869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_126 VNB N_A_2403_74#_c_1740_n 0.0129102f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_127 VNB N_A_37_464#_c_1912_n 0.040423f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_128 VNB N_A_37_464#_c_1913_n 0.00382492f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_129 VNB N_A_37_464#_c_1914_n 0.00686236f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_130 VNB N_A_37_464#_c_1915_n 0.030233f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_131 VNB N_A_37_464#_c_1916_n 0.00440078f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_132 VNB N_VPWR_c_2037_n 0.701046f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_133 VNB N_A_661_113#_c_2233_n 0.00969603f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_134 VNB N_A_661_113#_c_2234_n 0.00995999f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_135 VNB N_A_661_113#_c_2235_n 0.00711123f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_136 VNB N_A_661_113#_c_2236_n 0.00411745f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_137 VNB N_A_661_113#_c_2237_n 0.017599f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_138 VNB N_A_661_113#_c_2238_n 0.00447938f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_139 VNB N_A_661_113#_c_2239_n 0.00896457f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_140 VNB N_A_661_113#_c_2240_n 0.0172427f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_141 VNB N_Q_c_2415_n 0.00282627f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=1.145
cc_142 VNB N_Q_c_2416_n 0.00251582f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_143 VNB Q 0.0262057f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_144 VNB N_VGND_c_2467_n 0.0134335f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_145 VNB N_VGND_c_2468_n 0.0194143f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_146 VNB N_VGND_c_2469_n 0.00335587f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_147 VNB N_VGND_c_2470_n 0.0157372f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_148 VNB N_VGND_c_2471_n 0.00980185f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_149 VNB N_VGND_c_2472_n 0.00636294f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_150 VNB N_VGND_c_2473_n 0.00590394f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_151 VNB N_VGND_c_2474_n 0.0201354f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_152 VNB N_VGND_c_2475_n 0.0219434f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_153 VNB N_VGND_c_2476_n 0.0129417f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_154 VNB N_VGND_c_2477_n 0.0117383f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_155 VNB N_VGND_c_2478_n 0.0364019f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_156 VNB N_VGND_c_2479_n 0.029639f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_157 VNB N_VGND_c_2480_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_158 VNB N_VGND_c_2481_n 0.0207632f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_159 VNB N_VGND_c_2482_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_160 VNB N_VGND_c_2483_n 0.031383f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_161 VNB N_VGND_c_2484_n 0.0196191f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_162 VNB N_VGND_c_2485_n 0.0674297f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_163 VNB N_VGND_c_2486_n 0.058775f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_164 VNB N_VGND_c_2487_n 0.0298174f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_165 VNB N_VGND_c_2488_n 0.0177484f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_166 VNB N_VGND_c_2489_n 0.0162614f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_167 VNB N_VGND_c_2490_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_168 VNB N_VGND_c_2491_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_169 VNB N_VGND_c_2492_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_170 VNB N_VGND_c_2493_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_171 VNB N_VGND_c_2494_n 0.00461913f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_172 VNB N_VGND_c_2495_n 0.0392213f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_173 VNB N_VGND_c_2496_n 0.0320452f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_174 VNB N_VGND_c_2497_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_175 VNB N_VGND_c_2498_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_176 VNB N_VGND_c_2499_n 0.914074f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_177 VPB N_D_c_351_n 0.00978105f $X=-0.19 $Y=1.66 $X2=0.555 $Y2=2.155
cc_178 VPB N_D_c_352_n 0.0256033f $X=-0.19 $Y=1.66 $X2=0.555 $Y2=2.245
cc_179 VPB N_D_c_349_n 0.00449143f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=1.145
cc_180 VPB N_D_c_350_n 0.0112314f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=1.825
cc_181 VPB N_D_c_355_n 0.0155819f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=1.99
cc_182 VPB N_A_177_290#_c_397_n 0.0184392f $X=-0.19 $Y=1.66 $X2=0.6 $Y2=0.58
cc_183 VPB N_A_177_290#_c_398_n 0.0346249f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_184 VPB N_A_177_290#_c_391_n 0.0205394f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=1.145
cc_185 VPB N_A_177_290#_c_400_n 0.0129756f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=1.825
cc_186 VPB N_A_177_290#_c_401_n 0.00243214f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=1.99
cc_187 VPB N_A_177_290#_c_402_n 0.00254697f $X=-0.19 $Y=1.66 $X2=0.625 $Y2=1.825
cc_188 VPB N_A_177_290#_c_403_n 0.0139428f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_189 VPB N_A_177_290#_c_395_n 0.00517521f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_190 VPB N_A_177_290#_c_396_n 0.0208831f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_191 VPB N_DE_c_500_n 0.0237135f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=1.145
cc_192 VPB N_DE_c_506_n 0.0140005f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=0.98
cc_193 VPB N_DE_c_507_n 0.0118045f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.21
cc_194 VPB N_DE_c_508_n 0.0183363f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=1.825
cc_195 VPB N_DE_c_509_n 0.0349677f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=1.145
cc_196 VPB N_DE_c_510_n 0.0161255f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=1.825
cc_197 VPB N_DE_c_511_n 0.00488727f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_198 VPB N_DE_c_512_n 0.00321719f $X=-0.19 $Y=1.66 $X2=0.625 $Y2=1.825
cc_199 VPB N_A_545_87#_c_601_n 0.0252398f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.21
cc_200 VPB N_A_545_87#_c_602_n 0.0212328f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_201 VPB N_A_545_87#_c_603_n 0.0545994f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=1.825
cc_202 VPB N_A_545_87#_c_594_n 0.0192049f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_203 VPB N_A_545_87#_c_605_n 0.00534374f $X=-0.19 $Y=1.66 $X2=0.625 $Y2=1.295
cc_204 VPB N_A_545_87#_c_606_n 0.00883806f $X=-0.19 $Y=1.66 $X2=0.625 $Y2=1.825
cc_205 VPB N_A_545_87#_c_607_n 0.00845542f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_206 VPB N_A_545_87#_c_608_n 0.00288991f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_207 VPB N_A_545_87#_c_609_n 0.0030155f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_208 VPB N_A_545_87#_c_610_n 4.54166e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_209 VPB N_A_545_87#_c_597_n 0.0504699f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_210 VPB N_A_545_87#_c_598_n 0.00132032f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_211 VPB N_A_545_87#_c_613_n 0.00520352f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_212 VPB N_A_545_87#_c_614_n 0.00577276f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_213 VPB N_A_545_87#_c_599_n 0.0024967f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_214 VPB N_A_545_87#_c_600_n 0.0272242f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_215 VPB N_A_631_87#_c_842_n 0.0161815f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.21
cc_216 VPB N_A_631_87#_c_843_n 0.0241322f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=1.145
cc_217 VPB N_A_631_87#_c_837_n 0.0028825f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_218 VPB N_A_631_87#_c_838_n 0.0326079f $X=-0.19 $Y=1.66 $X2=0.625 $Y2=1.665
cc_219 VPB N_A_631_87#_c_846_n 0.00466068f $X=-0.19 $Y=1.66 $X2=0.625 $Y2=1.825
cc_220 VPB N_A_631_87#_c_847_n 0.019831f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_221 VPB N_A_631_87#_c_840_n 0.0201771f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_222 VPB N_A_631_87#_c_849_n 0.00579469f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_223 VPB N_A_631_87#_c_850_n 0.00833556f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_224 VPB N_SCD_c_949_n 0.0204058f $X=-0.19 $Y=1.66 $X2=0.6 $Y2=0.98
cc_225 VPB N_SCD_c_950_n 0.0215738f $X=-0.19 $Y=1.66 $X2=0.6 $Y2=0.58
cc_226 VPB SCD 0.00327296f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=1.145
cc_227 VPB N_SCD_c_948_n 0.00959317f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_228 VPB N_SCE_c_999_n 0.0185503f $X=-0.19 $Y=1.66 $X2=0.555 $Y2=1.99
cc_229 VPB N_SCE_c_1000_n 0.0805259f $X=-0.19 $Y=1.66 $X2=0.555 $Y2=2.64
cc_230 VPB N_SCE_c_1001_n 0.0132883f $X=-0.19 $Y=1.66 $X2=0.555 $Y2=2.64
cc_231 VPB N_SCE_c_992_n 0.0278804f $X=-0.19 $Y=1.66 $X2=0.6 $Y2=0.58
cc_232 VPB N_SCE_c_1003_n 0.00745008f $X=-0.19 $Y=1.66 $X2=0.6 $Y2=0.58
cc_233 VPB N_SCE_M1044_g 0.00949617f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=0.98
cc_234 VPB N_CLK_c_1081_n 0.0282303f $X=-0.19 $Y=1.66 $X2=0.555 $Y2=2.64
cc_235 VPB N_A_1510_74#_c_1140_n 0.0192339f $X=-0.19 $Y=1.66 $X2=0.6 $Y2=0.58
cc_236 VPB N_A_1510_74#_c_1117_n 0.0371508f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=1.145
cc_237 VPB N_A_1510_74#_c_1142_n 0.0218221f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=1.145
cc_238 VPB N_A_1510_74#_c_1143_n 0.00367481f $X=-0.19 $Y=1.66 $X2=0.625
+ $Y2=1.665
cc_239 VPB N_A_1510_74#_c_1121_n 0.0010342f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_240 VPB N_A_1510_74#_c_1131_n 0.00434787f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_241 VPB N_A_1510_74#_c_1132_n 0.018478f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_242 VPB N_A_1510_74#_c_1147_n 0.00744032f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_243 VPB N_A_1510_74#_c_1148_n 0.0566084f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_244 VPB N_A_1313_74#_c_1343_n 0.00979014f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=0.98
cc_245 VPB N_A_1313_74#_c_1358_n 0.0209485f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_246 VPB N_A_1313_74#_c_1344_n 0.0149626f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=1.825
cc_247 VPB N_A_1313_74#_c_1346_n 0.0172962f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=1.825
cc_248 VPB N_A_1313_74#_c_1361_n 0.0140471f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_249 VPB N_A_1313_74#_c_1362_n 0.056139f $X=-0.19 $Y=1.66 $X2=0.625 $Y2=1.295
cc_250 VPB N_A_1313_74#_c_1347_n 0.0406928f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_251 VPB N_A_1313_74#_c_1349_n 0.00167153f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_252 VPB N_A_1313_74#_c_1350_n 0.00416248f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_253 VPB N_A_1313_74#_c_1366_n 0.0060269f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_254 VPB N_A_1313_74#_c_1354_n 0.00267709f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_255 VPB N_A_1313_74#_c_1368_n 0.0140375f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_256 VPB N_A_1313_74#_c_1369_n 0.00283904f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_257 VPB N_A_1313_74#_c_1370_n 0.00864504f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_258 VPB N_A_1313_74#_c_1355_n 0.00182932f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_259 VPB N_A_1313_74#_c_1356_n 0.0466322f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_260 VPB N_A_1943_53#_c_1534_n 0.0410992f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.21
cc_261 VPB N_A_1943_53#_c_1546_n 0.0223908f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_262 VPB N_A_1943_53#_c_1535_n 0.00805235f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=1.145
cc_263 VPB N_A_1943_53#_c_1548_n 0.0301981f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=1.145
cc_264 VPB N_A_1943_53#_c_1549_n 0.00854378f $X=-0.19 $Y=1.66 $X2=0.625
+ $Y2=1.295
cc_265 VPB N_A_1943_53#_c_1539_n 0.00782072f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_266 VPB N_A_1756_97#_c_1639_n 0.0403098f $X=-0.19 $Y=1.66 $X2=0.6 $Y2=0.58
cc_267 VPB N_A_1756_97#_c_1645_n 0.00266461f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=1.825
cc_268 VPB N_A_1756_97#_c_1646_n 0.00723895f $X=-0.19 $Y=1.66 $X2=0.625
+ $Y2=1.295
cc_269 VPB N_A_1756_97#_c_1647_n 0.00923878f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_270 VPB N_A_1756_97#_c_1642_n 8.57241e-19 $X=-0.19 $Y=1.66 $X2=0.625
+ $Y2=1.825
cc_271 VPB N_A_1756_97#_c_1643_n 0.0115657f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_272 VPB N_A_2403_74#_c_1741_n 0.0106555f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_273 VPB N_A_2403_74#_c_1742_n 0.025635f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_274 VPB N_A_2403_74#_c_1729_n 0.0250854f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=1.145
cc_275 VPB N_A_2403_74#_c_1744_n 0.0175624f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=1.99
cc_276 VPB N_A_2403_74#_c_1745_n 0.0144283f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_277 VPB N_A_2403_74#_c_1746_n 0.0144424f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_278 VPB N_A_2403_74#_c_1747_n 0.0173786f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_279 VPB N_A_2403_74#_c_1734_n 0.048571f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_280 VPB N_A_2403_74#_c_1749_n 0.0029852f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_281 VPB N_A_2403_74#_c_1750_n 0.0104253f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_282 VPB N_A_2403_74#_c_1751_n 0.00470338f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_283 VPB N_A_2403_74#_c_1752_n 0.00541123f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_284 VPB N_A_2403_74#_c_1738_n 0.00121564f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_285 VPB N_A_2403_74#_c_1740_n 0.0289213f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_286 VPB N_A_37_464#_c_1912_n 0.0302506f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_287 VPB N_A_37_464#_c_1918_n 0.0252204f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=1.145
cc_288 VPB N_A_37_464#_c_1919_n 0.015179f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=1.145
cc_289 VPB N_A_37_464#_c_1920_n 0.00998336f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=1.825
cc_290 VPB N_A_37_464#_c_1921_n 0.00857095f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=1.99
cc_291 VPB N_A_37_464#_c_1922_n 0.00349119f $X=-0.19 $Y=1.66 $X2=0.625 $Y2=1.145
cc_292 VPB N_A_37_464#_c_1923_n 0.00548383f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_293 VPB N_A_37_464#_c_1924_n 8.46064e-19 $X=-0.19 $Y=1.66 $X2=0.625 $Y2=1.665
cc_294 VPB N_A_37_464#_c_1925_n 0.00216571f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_295 VPB N_A_37_464#_c_1914_n 0.0126751f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_296 VPB N_A_37_464#_c_1927_n 0.0127953f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_297 VPB N_A_37_464#_c_1928_n 0.00125429f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_298 VPB N_VPWR_c_2038_n 0.00600898f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_299 VPB N_VPWR_c_2039_n 0.00554607f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_300 VPB N_VPWR_c_2040_n 0.00745483f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_301 VPB N_VPWR_c_2041_n 0.0125325f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_302 VPB N_VPWR_c_2042_n 0.021494f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_303 VPB N_VPWR_c_2043_n 0.0115519f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_304 VPB N_VPWR_c_2044_n 0.0140087f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_305 VPB N_VPWR_c_2045_n 0.00880467f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_306 VPB N_VPWR_c_2046_n 0.019175f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_307 VPB N_VPWR_c_2047_n 0.0153587f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_308 VPB N_VPWR_c_2048_n 0.00261791f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_309 VPB N_VPWR_c_2049_n 0.0116916f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_310 VPB N_VPWR_c_2050_n 0.0348277f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_311 VPB N_VPWR_c_2051_n 0.0558311f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_312 VPB N_VPWR_c_2052_n 0.00614151f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_313 VPB N_VPWR_c_2053_n 0.0317338f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_314 VPB N_VPWR_c_2054_n 0.0296515f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_315 VPB N_VPWR_c_2055_n 0.0581188f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_316 VPB N_VPWR_c_2056_n 0.0306855f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_317 VPB N_VPWR_c_2057_n 0.0323948f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_318 VPB N_VPWR_c_2058_n 0.0223709f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_319 VPB N_VPWR_c_2059_n 0.0602391f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_320 VPB N_VPWR_c_2060_n 0.0160559f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_321 VPB N_VPWR_c_2061_n 0.0160949f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_322 VPB N_VPWR_c_2062_n 0.00460249f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_323 VPB N_VPWR_c_2063_n 0.00463855f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_324 VPB N_VPWR_c_2064_n 0.0047828f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_325 VPB N_VPWR_c_2065_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_326 VPB N_VPWR_c_2066_n 0.00614127f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_327 VPB N_VPWR_c_2067_n 0.00614151f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_328 VPB N_VPWR_c_2068_n 0.0101806f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_329 VPB N_VPWR_c_2069_n 0.00614127f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_330 VPB N_VPWR_c_2070_n 0.00601644f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_331 VPB N_VPWR_c_2037_n 0.20662f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_332 VPB N_A_661_113#_c_2241_n 0.0020929f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=1.825
cc_333 VPB N_A_661_113#_c_2242_n 0.00773134f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_334 VPB N_A_661_113#_c_2243_n 0.00104828f $X=-0.19 $Y=1.66 $X2=0.625
+ $Y2=1.825
cc_335 VPB N_A_661_113#_c_2234_n 0.0149909f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_336 VPB N_A_661_113#_c_2245_n 0.0235482f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_337 VPB N_A_661_113#_c_2246_n 0.00111442f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_338 VPB N_A_661_113#_c_2247_n 0.0152091f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_339 VPB N_A_661_113#_c_2239_n 0.00997354f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_340 VPB N_A_661_113#_c_2249_n 0.00798999f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_341 VPB N_A_661_113#_c_2250_n 0.00520801f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_342 VPB N_A_661_113#_c_2251_n 0.00866973f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_343 VPB N_Q_c_2418_n 0.00224686f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_344 VPB N_Q_c_2419_n 0.00220489f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=1.99
cc_345 VPB Q 0.0229398f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_346 N_D_c_352_n N_A_177_290#_c_397_n 0.0383469f $X=0.555 $Y=2.245 $X2=0 $Y2=0
cc_347 N_D_c_351_n N_A_177_290#_c_398_n 0.0143836f $X=0.555 $Y=2.155 $X2=0 $Y2=0
cc_348 N_D_c_355_n N_A_177_290#_c_398_n 0.0169938f $X=0.51 $Y=1.99 $X2=0 $Y2=0
cc_349 N_D_c_349_n N_A_177_290#_c_390_n 0.0651656f $X=0.51 $Y=1.145 $X2=0 $Y2=0
cc_350 N_D_c_350_n N_A_177_290#_c_390_n 0.00168519f $X=0.51 $Y=1.825 $X2=0 $Y2=0
cc_351 N_D_c_349_n N_A_177_290#_c_391_n 0.00402407f $X=0.51 $Y=1.145 $X2=0 $Y2=0
cc_352 N_D_c_350_n N_A_177_290#_c_391_n 0.0169938f $X=0.51 $Y=1.825 $X2=0 $Y2=0
cc_353 N_D_c_349_n N_A_177_290#_c_393_n 0.0144317f $X=0.51 $Y=1.145 $X2=0 $Y2=0
cc_354 N_D_c_351_n N_A_177_290#_c_401_n 6.66707e-19 $X=0.555 $Y=2.155 $X2=0
+ $Y2=0
cc_355 N_D_c_349_n N_A_177_290#_c_401_n 0.0034055f $X=0.51 $Y=1.145 $X2=0 $Y2=0
cc_356 N_D_M1002_g N_DE_M1034_g 0.0249061f $X=0.6 $Y=0.58 $X2=0 $Y2=0
cc_357 N_D_c_349_n N_DE_M1034_g 0.00172189f $X=0.51 $Y=1.145 $X2=0 $Y2=0
cc_358 N_D_c_348_n N_DE_c_499_n 0.0249061f $X=0.51 $Y=1.145 $X2=0 $Y2=0
cc_359 N_D_c_351_n N_A_37_464#_c_1912_n 0.00850381f $X=0.555 $Y=2.155 $X2=0
+ $Y2=0
cc_360 N_D_c_352_n N_A_37_464#_c_1912_n 0.00141989f $X=0.555 $Y=2.245 $X2=0
+ $Y2=0
cc_361 N_D_M1002_g N_A_37_464#_c_1912_n 0.00521378f $X=0.6 $Y=0.58 $X2=0 $Y2=0
cc_362 N_D_c_348_n N_A_37_464#_c_1912_n 0.0248496f $X=0.51 $Y=1.145 $X2=0 $Y2=0
cc_363 N_D_c_349_n N_A_37_464#_c_1912_n 0.0769553f $X=0.51 $Y=1.145 $X2=0 $Y2=0
cc_364 N_D_c_352_n N_A_37_464#_c_1918_n 0.0094621f $X=0.555 $Y=2.245 $X2=0 $Y2=0
cc_365 N_D_c_352_n N_A_37_464#_c_1919_n 0.0127112f $X=0.555 $Y=2.245 $X2=0 $Y2=0
cc_366 N_D_c_349_n N_A_37_464#_c_1919_n 0.0173118f $X=0.51 $Y=1.145 $X2=0 $Y2=0
cc_367 N_D_M1002_g N_A_37_464#_c_1915_n 0.0100933f $X=0.6 $Y=0.58 $X2=0 $Y2=0
cc_368 N_D_c_348_n N_A_37_464#_c_1915_n 0.00447722f $X=0.51 $Y=1.145 $X2=0 $Y2=0
cc_369 N_D_c_349_n N_A_37_464#_c_1915_n 0.0105828f $X=0.51 $Y=1.145 $X2=0 $Y2=0
cc_370 N_D_c_352_n N_A_37_464#_c_1927_n 0.00163791f $X=0.555 $Y=2.245 $X2=0
+ $Y2=0
cc_371 N_D_c_349_n N_A_37_464#_c_1927_n 0.0039504f $X=0.51 $Y=1.145 $X2=0 $Y2=0
cc_372 N_D_c_355_n N_A_37_464#_c_1927_n 0.00367821f $X=0.51 $Y=1.99 $X2=0 $Y2=0
cc_373 N_D_c_352_n N_VPWR_c_2038_n 0.001556f $X=0.555 $Y=2.245 $X2=0 $Y2=0
cc_374 N_D_c_352_n N_VPWR_c_2053_n 0.00445602f $X=0.555 $Y=2.245 $X2=0 $Y2=0
cc_375 N_D_c_352_n N_VPWR_c_2037_n 0.00861806f $X=0.555 $Y=2.245 $X2=0 $Y2=0
cc_376 N_D_M1002_g N_VGND_c_2467_n 0.00184547f $X=0.6 $Y=0.58 $X2=0 $Y2=0
cc_377 N_D_M1002_g N_VGND_c_2483_n 0.00432935f $X=0.6 $Y=0.58 $X2=0 $Y2=0
cc_378 N_D_M1002_g N_VGND_c_2499_n 0.00821127f $X=0.6 $Y=0.58 $X2=0 $Y2=0
cc_379 N_A_177_290#_c_393_n N_DE_M1034_g 0.00568157f $X=1.325 $Y=1.065 $X2=0
+ $Y2=0
cc_380 N_A_177_290#_c_394_n N_DE_M1034_g 0.00465695f $X=1.765 $Y=0.775 $X2=0
+ $Y2=0
cc_381 N_A_177_290#_c_390_n N_DE_c_498_n 0.00689963f $X=1.16 $Y=1.615 $X2=0
+ $Y2=0
cc_382 N_A_177_290#_c_392_n N_DE_c_498_n 0.012769f $X=1.6 $Y=1.065 $X2=0 $Y2=0
cc_383 N_A_177_290#_c_393_n N_DE_c_498_n 0.00487554f $X=1.325 $Y=1.065 $X2=0
+ $Y2=0
cc_384 N_A_177_290#_c_390_n N_DE_c_499_n 0.00149654f $X=1.16 $Y=1.615 $X2=0
+ $Y2=0
cc_385 N_A_177_290#_c_391_n N_DE_c_499_n 0.0241421f $X=1.16 $Y=1.615 $X2=0 $Y2=0
cc_386 N_A_177_290#_c_393_n N_DE_c_499_n 0.0011888f $X=1.325 $Y=1.065 $X2=0
+ $Y2=0
cc_387 N_A_177_290#_c_390_n N_DE_c_500_n 0.00113204f $X=1.16 $Y=1.615 $X2=0
+ $Y2=0
cc_388 N_A_177_290#_c_391_n N_DE_c_500_n 0.00797738f $X=1.16 $Y=1.615 $X2=0
+ $Y2=0
cc_389 N_A_177_290#_c_400_n N_DE_c_500_n 0.00486542f $X=1.795 $Y=2.035 $X2=0
+ $Y2=0
cc_390 N_A_177_290#_c_403_n N_DE_c_500_n 0.00420828f $X=2.24 $Y=1.95 $X2=0 $Y2=0
cc_391 N_A_177_290#_c_395_n N_DE_c_500_n 0.00375194f $X=2.24 $Y=1.685 $X2=0
+ $Y2=0
cc_392 N_A_177_290#_c_396_n N_DE_c_500_n 0.0109698f $X=2.41 $Y=1.685 $X2=0 $Y2=0
cc_393 N_A_177_290#_c_402_n N_DE_c_506_n 0.0100315f $X=1.88 $Y=2.515 $X2=0 $Y2=0
cc_394 N_A_177_290#_c_403_n N_DE_c_506_n 0.00650102f $X=2.24 $Y=1.95 $X2=0 $Y2=0
cc_395 N_A_177_290#_c_398_n N_DE_c_507_n 0.0113421f $X=1.105 $Y=1.9 $X2=0 $Y2=0
cc_396 N_A_177_290#_c_400_n N_DE_c_507_n 0.00486672f $X=1.795 $Y=2.035 $X2=0
+ $Y2=0
cc_397 N_A_177_290#_c_402_n N_DE_c_507_n 0.00599009f $X=1.88 $Y=2.515 $X2=0
+ $Y2=0
cc_398 N_A_177_290#_c_403_n N_DE_c_507_n 2.32181e-19 $X=2.24 $Y=1.95 $X2=0 $Y2=0
cc_399 N_A_177_290#_M1038_g N_DE_c_501_n 0.0188666f $X=2.41 $Y=0.775 $X2=0 $Y2=0
cc_400 N_A_177_290#_c_392_n N_DE_c_501_n 0.00310065f $X=1.6 $Y=1.065 $X2=0 $Y2=0
cc_401 N_A_177_290#_c_394_n N_DE_c_501_n 9.22767e-19 $X=1.765 $Y=0.775 $X2=0
+ $Y2=0
cc_402 N_A_177_290#_c_402_n N_DE_c_508_n 0.00415054f $X=1.88 $Y=2.515 $X2=0
+ $Y2=0
cc_403 N_A_177_290#_c_403_n N_DE_c_509_n 0.00505749f $X=2.24 $Y=1.95 $X2=0 $Y2=0
cc_404 N_A_177_290#_c_392_n N_DE_c_502_n 0.0146667f $X=1.6 $Y=1.065 $X2=0 $Y2=0
cc_405 N_A_177_290#_c_403_n N_DE_c_511_n 0.00708655f $X=2.24 $Y=1.95 $X2=0 $Y2=0
cc_406 N_A_177_290#_c_395_n N_DE_c_511_n 2.41872e-19 $X=2.24 $Y=1.685 $X2=0
+ $Y2=0
cc_407 N_A_177_290#_c_396_n N_DE_c_511_n 0.0231424f $X=2.41 $Y=1.685 $X2=0 $Y2=0
cc_408 N_A_177_290#_M1038_g N_DE_c_503_n 0.0092673f $X=2.41 $Y=0.775 $X2=0 $Y2=0
cc_409 N_A_177_290#_c_390_n N_DE_c_503_n 0.00782514f $X=1.16 $Y=1.615 $X2=0
+ $Y2=0
cc_410 N_A_177_290#_c_391_n N_DE_c_503_n 0.0124286f $X=1.16 $Y=1.615 $X2=0 $Y2=0
cc_411 N_A_177_290#_M1038_g N_DE_c_512_n 0.0010882f $X=2.41 $Y=0.775 $X2=0 $Y2=0
cc_412 N_A_177_290#_c_390_n N_DE_c_512_n 0.0302117f $X=1.16 $Y=1.615 $X2=0 $Y2=0
cc_413 N_A_177_290#_c_391_n N_DE_c_512_n 0.0017489f $X=1.16 $Y=1.615 $X2=0 $Y2=0
cc_414 N_A_177_290#_c_392_n N_DE_c_512_n 0.0250522f $X=1.6 $Y=1.065 $X2=0 $Y2=0
cc_415 N_A_177_290#_c_400_n N_DE_c_512_n 0.0255862f $X=1.795 $Y=2.035 $X2=0
+ $Y2=0
cc_416 N_A_177_290#_c_395_n N_DE_c_512_n 0.0145882f $X=2.24 $Y=1.685 $X2=0 $Y2=0
cc_417 N_A_177_290#_c_396_n N_DE_c_512_n 0.00136208f $X=2.41 $Y=1.685 $X2=0
+ $Y2=0
cc_418 N_A_177_290#_c_400_n N_DE_c_504_n 7.51173e-19 $X=1.795 $Y=2.035 $X2=0
+ $Y2=0
cc_419 N_A_177_290#_c_395_n N_DE_c_504_n 4.2711e-19 $X=2.24 $Y=1.685 $X2=0 $Y2=0
cc_420 N_A_177_290#_c_396_n N_DE_c_504_n 0.00811139f $X=2.41 $Y=1.685 $X2=0
+ $Y2=0
cc_421 N_A_177_290#_M1038_g N_A_545_87#_M1023_g 0.0369968f $X=2.41 $Y=0.775
+ $X2=0 $Y2=0
cc_422 N_A_177_290#_c_395_n N_A_545_87#_c_598_n 0.0074941f $X=2.24 $Y=1.685
+ $X2=0 $Y2=0
cc_423 N_A_177_290#_c_396_n N_A_545_87#_c_598_n 0.00471443f $X=2.41 $Y=1.685
+ $X2=0 $Y2=0
cc_424 N_A_177_290#_c_395_n N_A_545_87#_c_599_n 0.0230196f $X=2.24 $Y=1.685
+ $X2=0 $Y2=0
cc_425 N_A_177_290#_c_396_n N_A_545_87#_c_599_n 0.00251924f $X=2.41 $Y=1.685
+ $X2=0 $Y2=0
cc_426 N_A_177_290#_c_395_n N_A_545_87#_c_600_n 2.47097e-19 $X=2.24 $Y=1.685
+ $X2=0 $Y2=0
cc_427 N_A_177_290#_c_396_n N_A_545_87#_c_600_n 0.0369968f $X=2.41 $Y=1.685
+ $X2=0 $Y2=0
cc_428 N_A_177_290#_c_397_n N_A_37_464#_c_1918_n 0.00182013f $X=0.975 $Y=2.245
+ $X2=0 $Y2=0
cc_429 N_A_177_290#_c_397_n N_A_37_464#_c_1919_n 0.0190988f $X=0.975 $Y=2.245
+ $X2=0 $Y2=0
cc_430 N_A_177_290#_c_398_n N_A_37_464#_c_1919_n 0.00298207f $X=1.105 $Y=1.9
+ $X2=0 $Y2=0
cc_431 N_A_177_290#_c_400_n N_A_37_464#_c_1919_n 0.0240721f $X=1.795 $Y=2.035
+ $X2=0 $Y2=0
cc_432 N_A_177_290#_c_401_n N_A_37_464#_c_1919_n 0.0260821f $X=1.325 $Y=2.035
+ $X2=0 $Y2=0
cc_433 N_A_177_290#_c_402_n N_A_37_464#_c_1919_n 0.0141649f $X=1.88 $Y=2.515
+ $X2=0 $Y2=0
cc_434 N_A_177_290#_c_397_n N_A_37_464#_c_1920_n 0.00426176f $X=0.975 $Y=2.245
+ $X2=0 $Y2=0
cc_435 N_A_177_290#_c_402_n N_A_37_464#_c_1920_n 0.0203028f $X=1.88 $Y=2.515
+ $X2=0 $Y2=0
cc_436 N_A_177_290#_M1001_s N_A_37_464#_c_1921_n 0.00320543f $X=1.735 $Y=2.315
+ $X2=0 $Y2=0
cc_437 N_A_177_290#_c_402_n N_A_37_464#_c_1921_n 0.0126885f $X=1.88 $Y=2.515
+ $X2=0 $Y2=0
cc_438 N_A_177_290#_c_397_n N_A_37_464#_c_1922_n 6.5162e-19 $X=0.975 $Y=2.245
+ $X2=0 $Y2=0
cc_439 N_A_177_290#_c_402_n N_A_37_464#_c_1954_n 0.0192722f $X=1.88 $Y=2.515
+ $X2=0 $Y2=0
cc_440 N_A_177_290#_c_403_n N_A_37_464#_c_1923_n 0.00425322f $X=2.24 $Y=1.95
+ $X2=0 $Y2=0
cc_441 N_A_177_290#_c_402_n N_A_37_464#_c_1924_n 0.0133944f $X=1.88 $Y=2.515
+ $X2=0 $Y2=0
cc_442 N_A_177_290#_c_403_n N_A_37_464#_c_1924_n 0.0134805f $X=2.24 $Y=1.95
+ $X2=0 $Y2=0
cc_443 N_A_177_290#_M1038_g N_A_37_464#_c_1913_n 0.00214472f $X=2.41 $Y=0.775
+ $X2=0 $Y2=0
cc_444 N_A_177_290#_M1038_g N_A_37_464#_c_1916_n 8.26272e-19 $X=2.41 $Y=0.775
+ $X2=0 $Y2=0
cc_445 N_A_177_290#_c_397_n N_VPWR_c_2038_n 0.0107235f $X=0.975 $Y=2.245 $X2=0
+ $Y2=0
cc_446 N_A_177_290#_c_397_n N_VPWR_c_2053_n 0.00413917f $X=0.975 $Y=2.245 $X2=0
+ $Y2=0
cc_447 N_A_177_290#_c_397_n N_VPWR_c_2037_n 0.00817532f $X=0.975 $Y=2.245 $X2=0
+ $Y2=0
cc_448 N_A_177_290#_c_392_n N_VGND_c_2467_n 0.00367796f $X=1.6 $Y=1.065 $X2=0
+ $Y2=0
cc_449 N_A_177_290#_c_393_n N_VGND_c_2467_n 0.0263911f $X=1.325 $Y=1.065 $X2=0
+ $Y2=0
cc_450 N_A_177_290#_c_394_n N_VGND_c_2467_n 0.0174982f $X=1.765 $Y=0.775 $X2=0
+ $Y2=0
cc_451 N_A_177_290#_M1038_g N_VGND_c_2468_n 0.0128771f $X=2.41 $Y=0.775 $X2=0
+ $Y2=0
cc_452 N_A_177_290#_c_392_n N_VGND_c_2468_n 0.00175056f $X=1.6 $Y=1.065 $X2=0
+ $Y2=0
cc_453 N_A_177_290#_c_394_n N_VGND_c_2468_n 0.0163189f $X=1.765 $Y=0.775 $X2=0
+ $Y2=0
cc_454 N_A_177_290#_c_395_n N_VGND_c_2468_n 0.00899549f $X=2.24 $Y=1.685 $X2=0
+ $Y2=0
cc_455 N_A_177_290#_c_396_n N_VGND_c_2468_n 0.00272206f $X=2.41 $Y=1.685 $X2=0
+ $Y2=0
cc_456 N_A_177_290#_c_394_n N_VGND_c_2484_n 0.00607888f $X=1.765 $Y=0.775 $X2=0
+ $Y2=0
cc_457 N_A_177_290#_M1038_g N_VGND_c_2485_n 0.00372658f $X=2.41 $Y=0.775 $X2=0
+ $Y2=0
cc_458 N_A_177_290#_M1038_g N_VGND_c_2499_n 0.00408518f $X=2.41 $Y=0.775 $X2=0
+ $Y2=0
cc_459 N_A_177_290#_c_394_n N_VGND_c_2499_n 0.00799492f $X=1.765 $Y=0.775 $X2=0
+ $Y2=0
cc_460 N_DE_c_509_n N_A_545_87#_c_601_n 0.0106312f $X=2.71 $Y=2.165 $X2=0 $Y2=0
cc_461 N_DE_c_510_n N_A_545_87#_c_602_n 0.0437219f $X=2.785 $Y=2.24 $X2=0 $Y2=0
cc_462 N_DE_c_509_n N_A_545_87#_c_598_n 8.44289e-19 $X=2.71 $Y=2.165 $X2=0 $Y2=0
cc_463 N_DE_c_509_n N_A_545_87#_c_599_n 0.00534454f $X=2.71 $Y=2.165 $X2=0 $Y2=0
cc_464 N_DE_c_509_n N_A_545_87#_c_600_n 0.0090241f $X=2.71 $Y=2.165 $X2=0 $Y2=0
cc_465 N_DE_c_508_n N_A_37_464#_c_1920_n 0.00326422f $X=2.105 $Y=2.24 $X2=0
+ $Y2=0
cc_466 N_DE_c_506_n N_A_37_464#_c_1921_n 7.52982e-19 $X=2.03 $Y=2.165 $X2=0
+ $Y2=0
cc_467 N_DE_c_507_n N_A_37_464#_c_1921_n 0.00321107f $X=1.835 $Y=2.165 $X2=0
+ $Y2=0
cc_468 N_DE_c_508_n N_A_37_464#_c_1921_n 0.0134964f $X=2.105 $Y=2.24 $X2=0 $Y2=0
cc_469 N_DE_c_510_n N_A_37_464#_c_1921_n 4.28313e-19 $X=2.785 $Y=2.24 $X2=0
+ $Y2=0
cc_470 N_DE_c_508_n N_A_37_464#_c_1954_n 0.0118088f $X=2.105 $Y=2.24 $X2=0 $Y2=0
cc_471 N_DE_c_510_n N_A_37_464#_c_1954_n 0.00283455f $X=2.785 $Y=2.24 $X2=0
+ $Y2=0
cc_472 N_DE_c_509_n N_A_37_464#_c_1923_n 0.0105252f $X=2.71 $Y=2.165 $X2=0 $Y2=0
cc_473 N_DE_c_510_n N_A_37_464#_c_1923_n 0.0154946f $X=2.785 $Y=2.24 $X2=0 $Y2=0
cc_474 N_DE_c_508_n N_A_37_464#_c_1924_n 0.00584584f $X=2.105 $Y=2.24 $X2=0
+ $Y2=0
cc_475 N_DE_c_509_n N_A_37_464#_c_1924_n 8.1141e-19 $X=2.71 $Y=2.165 $X2=0 $Y2=0
cc_476 N_DE_c_510_n N_A_37_464#_c_1925_n 0.00179485f $X=2.785 $Y=2.24 $X2=0
+ $Y2=0
cc_477 N_DE_M1034_g N_A_37_464#_c_1915_n 0.00132346f $X=0.99 $Y=0.58 $X2=0 $Y2=0
cc_478 N_DE_c_508_n N_VPWR_c_2039_n 0.00153478f $X=2.105 $Y=2.24 $X2=0 $Y2=0
cc_479 N_DE_c_510_n N_VPWR_c_2039_n 0.00967911f $X=2.785 $Y=2.24 $X2=0 $Y2=0
cc_480 N_DE_c_508_n N_VPWR_c_2054_n 0.00275664f $X=2.105 $Y=2.24 $X2=0 $Y2=0
cc_481 N_DE_c_510_n N_VPWR_c_2055_n 0.00410286f $X=2.785 $Y=2.24 $X2=0 $Y2=0
cc_482 N_DE_c_508_n N_VPWR_c_2037_n 0.00544287f $X=2.105 $Y=2.24 $X2=0 $Y2=0
cc_483 N_DE_c_510_n N_VPWR_c_2037_n 0.00493487f $X=2.785 $Y=2.24 $X2=0 $Y2=0
cc_484 N_DE_M1034_g N_VGND_c_2467_n 0.0140397f $X=0.99 $Y=0.58 $X2=0 $Y2=0
cc_485 N_DE_c_498_n N_VGND_c_2467_n 0.00140666f $X=1.535 $Y=1.135 $X2=0 $Y2=0
cc_486 N_DE_c_501_n N_VGND_c_2467_n 0.00221288f $X=1.98 $Y=1.06 $X2=0 $Y2=0
cc_487 N_DE_c_501_n N_VGND_c_2468_n 0.0112174f $X=1.98 $Y=1.06 $X2=0 $Y2=0
cc_488 N_DE_M1034_g N_VGND_c_2483_n 0.00383152f $X=0.99 $Y=0.58 $X2=0 $Y2=0
cc_489 N_DE_c_501_n N_VGND_c_2484_n 0.00372658f $X=1.98 $Y=1.06 $X2=0 $Y2=0
cc_490 N_DE_M1034_g N_VGND_c_2499_n 0.0075725f $X=0.99 $Y=0.58 $X2=0 $Y2=0
cc_491 N_DE_c_501_n N_VGND_c_2499_n 0.00408518f $X=1.98 $Y=1.06 $X2=0 $Y2=0
cc_492 N_A_545_87#_M1023_g N_A_631_87#_c_831_n 0.0180128f $X=2.8 $Y=0.775 $X2=0
+ $Y2=0
cc_493 N_A_545_87#_c_597_n N_A_631_87#_c_832_n 0.00541449f $X=14.495 $Y=1.665
+ $X2=0 $Y2=0
cc_494 N_A_545_87#_c_600_n N_A_631_87#_c_833_n 0.00439178f $X=3.175 $Y=1.685
+ $X2=0 $Y2=0
cc_495 N_A_545_87#_c_597_n N_A_631_87#_c_837_n 0.0247491f $X=14.495 $Y=1.665
+ $X2=0 $Y2=0
cc_496 N_A_545_87#_c_597_n N_A_631_87#_c_838_n 0.00741108f $X=14.495 $Y=1.665
+ $X2=0 $Y2=0
cc_497 N_A_545_87#_c_600_n N_A_631_87#_c_838_n 0.00544411f $X=3.175 $Y=1.685
+ $X2=0 $Y2=0
cc_498 N_A_545_87#_c_597_n N_A_631_87#_c_847_n 0.0362481f $X=14.495 $Y=1.665
+ $X2=0 $Y2=0
cc_499 N_A_545_87#_c_597_n N_A_631_87#_c_839_n 0.0160887f $X=14.495 $Y=1.665
+ $X2=0 $Y2=0
cc_500 N_A_545_87#_c_597_n N_A_631_87#_c_840_n 0.00341536f $X=14.495 $Y=1.665
+ $X2=0 $Y2=0
cc_501 N_A_545_87#_c_597_n N_A_631_87#_c_841_n 0.00653743f $X=14.495 $Y=1.665
+ $X2=0 $Y2=0
cc_502 N_A_545_87#_c_597_n N_A_631_87#_c_850_n 7.90379e-19 $X=14.495 $Y=1.665
+ $X2=0 $Y2=0
cc_503 N_A_545_87#_c_597_n SCD 0.0332863f $X=14.495 $Y=1.665 $X2=0 $Y2=0
cc_504 N_A_545_87#_c_597_n N_SCD_c_948_n 6.94548e-19 $X=14.495 $Y=1.665 $X2=0
+ $Y2=0
cc_505 N_A_545_87#_c_602_n N_SCE_c_999_n 0.0074134f $X=3.175 $Y=2.24 $X2=-0.19
+ $Y2=-0.245
cc_506 N_A_545_87#_c_597_n N_SCE_c_999_n 0.00250527f $X=14.495 $Y=1.665
+ $X2=-0.19 $Y2=-0.245
cc_507 N_A_545_87#_c_602_n N_SCE_c_1001_n 0.00288121f $X=3.175 $Y=2.24 $X2=0
+ $Y2=0
cc_508 N_A_545_87#_c_597_n N_SCE_c_992_n 0.0060229f $X=14.495 $Y=1.665 $X2=0
+ $Y2=0
cc_509 N_A_545_87#_c_597_n N_SCE_M1003_g 0.0030065f $X=14.495 $Y=1.665 $X2=0
+ $Y2=0
cc_510 N_A_545_87#_c_597_n SCE 0.0100898f $X=14.495 $Y=1.665 $X2=0 $Y2=0
cc_511 N_A_545_87#_c_597_n N_SCE_c_998_n 0.00432538f $X=14.495 $Y=1.665 $X2=0
+ $Y2=0
cc_512 N_A_545_87#_c_597_n N_CLK_c_1081_n 0.0120231f $X=14.495 $Y=1.665 $X2=0
+ $Y2=0
cc_513 N_A_545_87#_c_597_n CLK 0.0239464f $X=14.495 $Y=1.665 $X2=0 $Y2=0
cc_514 N_A_545_87#_c_603_n N_A_1510_74#_c_1117_n 0.020204f $X=13.275 $Y=2.465
+ $X2=0 $Y2=0
cc_515 N_A_545_87#_c_594_n N_A_1510_74#_c_1117_n 0.0141746f $X=13.41 $Y=2.05
+ $X2=0 $Y2=0
cc_516 N_A_545_87#_c_608_n N_A_1510_74#_c_1117_n 8.21089e-19 $X=13.485 $Y=2.222
+ $X2=0 $Y2=0
cc_517 N_A_545_87#_c_597_n N_A_1510_74#_c_1117_n 0.00571827f $X=14.495 $Y=1.665
+ $X2=0 $Y2=0
cc_518 N_A_545_87#_c_603_n N_A_1510_74#_c_1142_n 0.032062f $X=13.275 $Y=2.465
+ $X2=0 $Y2=0
cc_519 N_A_545_87#_c_597_n N_A_1510_74#_c_1118_n 0.00543427f $X=14.495 $Y=1.665
+ $X2=0 $Y2=0
cc_520 N_A_545_87#_c_597_n N_A_1510_74#_c_1143_n 0.0148651f $X=14.495 $Y=1.665
+ $X2=0 $Y2=0
cc_521 N_A_545_87#_c_597_n N_A_1510_74#_c_1121_n 0.0201438f $X=14.495 $Y=1.665
+ $X2=0 $Y2=0
cc_522 N_A_545_87#_c_597_n N_A_1510_74#_c_1124_n 0.00493977f $X=14.495 $Y=1.665
+ $X2=0 $Y2=0
cc_523 N_A_545_87#_c_597_n N_A_1510_74#_c_1128_n 0.00657297f $X=14.495 $Y=1.665
+ $X2=0 $Y2=0
cc_524 N_A_545_87#_c_597_n N_A_1510_74#_c_1131_n 0.0345923f $X=14.495 $Y=1.665
+ $X2=0 $Y2=0
cc_525 N_A_545_87#_c_597_n N_A_1510_74#_c_1132_n 0.0041349f $X=14.495 $Y=1.665
+ $X2=0 $Y2=0
cc_526 N_A_545_87#_c_593_n N_A_1510_74#_c_1133_n 2.40283e-19 $X=12.88 $Y=0.94
+ $X2=0 $Y2=0
cc_527 N_A_545_87#_c_597_n N_A_1510_74#_c_1133_n 0.0153966f $X=14.495 $Y=1.665
+ $X2=0 $Y2=0
cc_528 N_A_545_87#_c_597_n N_A_1510_74#_c_1147_n 0.00675777f $X=14.495 $Y=1.665
+ $X2=0 $Y2=0
cc_529 N_A_545_87#_c_597_n N_A_1510_74#_c_1135_n 0.00778786f $X=14.495 $Y=1.665
+ $X2=0 $Y2=0
cc_530 N_A_545_87#_c_597_n N_A_1510_74#_c_1136_n 4.85293e-19 $X=14.495 $Y=1.665
+ $X2=0 $Y2=0
cc_531 N_A_545_87#_c_593_n N_A_1510_74#_c_1138_n 0.0011337f $X=12.88 $Y=0.94
+ $X2=0 $Y2=0
cc_532 N_A_545_87#_c_594_n N_A_1510_74#_c_1138_n 7.75578e-19 $X=13.41 $Y=2.05
+ $X2=0 $Y2=0
cc_533 N_A_545_87#_c_597_n N_A_1510_74#_c_1138_n 0.00932399f $X=14.495 $Y=1.665
+ $X2=0 $Y2=0
cc_534 N_A_545_87#_c_593_n N_A_1510_74#_c_1139_n 0.0181563f $X=12.88 $Y=0.94
+ $X2=0 $Y2=0
cc_535 N_A_545_87#_c_594_n N_A_1510_74#_c_1139_n 0.0173139f $X=13.41 $Y=2.05
+ $X2=0 $Y2=0
cc_536 N_A_545_87#_c_597_n N_A_1313_74#_M1013_g 0.00592482f $X=14.495 $Y=1.665
+ $X2=0 $Y2=0
cc_537 N_A_545_87#_c_597_n N_A_1313_74#_c_1343_n 0.00385573f $X=14.495 $Y=1.665
+ $X2=0 $Y2=0
cc_538 N_A_545_87#_c_597_n N_A_1313_74#_c_1344_n 0.00449609f $X=14.495 $Y=1.665
+ $X2=0 $Y2=0
cc_539 N_A_545_87#_c_597_n N_A_1313_74#_M1040_g 0.00507242f $X=14.495 $Y=1.665
+ $X2=0 $Y2=0
cc_540 N_A_545_87#_c_597_n N_A_1313_74#_c_1346_n 0.00251542f $X=14.495 $Y=1.665
+ $X2=0 $Y2=0
cc_541 N_A_545_87#_c_597_n N_A_1313_74#_c_1347_n 6.94548e-19 $X=14.495 $Y=1.665
+ $X2=0 $Y2=0
cc_542 N_A_545_87#_c_591_n N_A_1313_74#_M1016_g 0.04003f $X=12.805 $Y=0.865
+ $X2=0 $Y2=0
cc_543 N_A_545_87#_c_597_n N_A_1313_74#_c_1349_n 0.002118f $X=14.495 $Y=1.665
+ $X2=0 $Y2=0
cc_544 N_A_545_87#_c_597_n N_A_1313_74#_c_1350_n 9.81771e-19 $X=14.495 $Y=1.665
+ $X2=0 $Y2=0
cc_545 N_A_545_87#_c_597_n N_A_1313_74#_c_1366_n 0.0200713f $X=14.495 $Y=1.665
+ $X2=0 $Y2=0
cc_546 N_A_545_87#_c_597_n N_A_1313_74#_c_1352_n 0.00549588f $X=14.495 $Y=1.665
+ $X2=0 $Y2=0
cc_547 N_A_545_87#_c_597_n N_A_1313_74#_c_1354_n 0.0245154f $X=14.495 $Y=1.665
+ $X2=0 $Y2=0
cc_548 N_A_545_87#_c_597_n N_A_1313_74#_c_1369_n 0.0030857f $X=14.495 $Y=1.665
+ $X2=0 $Y2=0
cc_549 N_A_545_87#_c_597_n N_A_1313_74#_c_1370_n 0.00240344f $X=14.495 $Y=1.665
+ $X2=0 $Y2=0
cc_550 N_A_545_87#_c_597_n N_A_1313_74#_c_1355_n 0.0267747f $X=14.495 $Y=1.665
+ $X2=0 $Y2=0
cc_551 N_A_545_87#_c_597_n N_A_1313_74#_c_1356_n 0.00390688f $X=14.495 $Y=1.665
+ $X2=0 $Y2=0
cc_552 N_A_545_87#_c_597_n N_A_1943_53#_c_1534_n 0.00219985f $X=14.495 $Y=1.665
+ $X2=0 $Y2=0
cc_553 N_A_545_87#_c_597_n N_A_1943_53#_c_1535_n 0.0120698f $X=14.495 $Y=1.665
+ $X2=0 $Y2=0
cc_554 N_A_545_87#_c_597_n N_A_1943_53#_c_1537_n 0.00782264f $X=14.495 $Y=1.665
+ $X2=0 $Y2=0
cc_555 N_A_545_87#_c_597_n N_A_1943_53#_c_1549_n 0.00570645f $X=14.495 $Y=1.665
+ $X2=0 $Y2=0
cc_556 N_A_545_87#_c_597_n N_A_1943_53#_c_1539_n 0.0251769f $X=14.495 $Y=1.665
+ $X2=0 $Y2=0
cc_557 N_A_545_87#_c_597_n N_A_1943_53#_c_1540_n 0.00488667f $X=14.495 $Y=1.665
+ $X2=0 $Y2=0
cc_558 N_A_545_87#_c_597_n N_A_1943_53#_c_1541_n 0.0277714f $X=14.495 $Y=1.665
+ $X2=0 $Y2=0
cc_559 N_A_545_87#_c_597_n N_A_1943_53#_c_1542_n 0.00410529f $X=14.495 $Y=1.665
+ $X2=0 $Y2=0
cc_560 N_A_545_87#_c_597_n N_A_1943_53#_c_1543_n 0.0075983f $X=14.495 $Y=1.665
+ $X2=0 $Y2=0
cc_561 N_A_545_87#_c_597_n N_A_1943_53#_c_1544_n 0.00838974f $X=14.495 $Y=1.665
+ $X2=0 $Y2=0
cc_562 N_A_545_87#_c_597_n N_A_1756_97#_c_1639_n 0.00189408f $X=14.495 $Y=1.665
+ $X2=0 $Y2=0
cc_563 N_A_545_87#_c_597_n N_A_1756_97#_c_1641_n 0.0110565f $X=14.495 $Y=1.665
+ $X2=0 $Y2=0
cc_564 N_A_545_87#_c_597_n N_A_1756_97#_c_1645_n 0.0126357f $X=14.495 $Y=1.665
+ $X2=0 $Y2=0
cc_565 N_A_545_87#_c_597_n N_A_1756_97#_c_1647_n 0.00152612f $X=14.495 $Y=1.665
+ $X2=0 $Y2=0
cc_566 N_A_545_87#_c_597_n N_A_1756_97#_c_1642_n 0.0219629f $X=14.495 $Y=1.665
+ $X2=0 $Y2=0
cc_567 N_A_545_87#_c_597_n N_A_1756_97#_c_1643_n 0.0554309f $X=14.495 $Y=1.665
+ $X2=0 $Y2=0
cc_568 N_A_545_87#_c_594_n N_A_2403_74#_c_1727_n 0.0275433f $X=13.41 $Y=2.05
+ $X2=0 $Y2=0
cc_569 N_A_545_87#_c_592_n N_A_2403_74#_M1021_g 0.00417986f $X=13.335 $Y=0.94
+ $X2=0 $Y2=0
cc_570 N_A_545_87#_c_595_n N_A_2403_74#_M1021_g 0.00563211f $X=14.31 $Y=1.55
+ $X2=0 $Y2=0
cc_571 N_A_545_87#_c_596_n N_A_2403_74#_M1021_g 0.0113373f $X=14.17 $Y=0.58
+ $X2=0 $Y2=0
cc_572 N_A_545_87#_c_594_n N_A_2403_74#_c_1741_n 0.00391262f $X=13.41 $Y=2.05
+ $X2=0 $Y2=0
cc_573 N_A_545_87#_c_608_n N_A_2403_74#_c_1741_n 4.87494e-19 $X=13.485 $Y=2.222
+ $X2=0 $Y2=0
cc_574 N_A_545_87#_c_603_n N_A_2403_74#_c_1742_n 0.0196904f $X=13.275 $Y=2.465
+ $X2=0 $Y2=0
cc_575 N_A_545_87#_c_605_n N_A_2403_74#_c_1742_n 0.0131432f $X=14.045 $Y=2.265
+ $X2=0 $Y2=0
cc_576 N_A_545_87#_c_606_n N_A_2403_74#_c_1742_n 0.0102172f $X=14.21 $Y=2.465
+ $X2=0 $Y2=0
cc_577 N_A_545_87#_c_609_n N_A_2403_74#_c_1742_n 0.00416765f $X=14.22 $Y=2.265
+ $X2=0 $Y2=0
cc_578 N_A_545_87#_c_595_n N_A_2403_74#_c_1729_n 0.0154738f $X=14.31 $Y=1.55
+ $X2=0 $Y2=0
cc_579 N_A_545_87#_c_596_n N_A_2403_74#_c_1729_n 0.00161436f $X=14.17 $Y=0.58
+ $X2=0 $Y2=0
cc_580 N_A_545_87#_c_609_n N_A_2403_74#_c_1729_n 0.00386993f $X=14.22 $Y=2.265
+ $X2=0 $Y2=0
cc_581 N_A_545_87#_c_610_n N_A_2403_74#_c_1729_n 0.00751453f $X=14.31 $Y=1.665
+ $X2=0 $Y2=0
cc_582 N_A_545_87#_c_597_n N_A_2403_74#_c_1729_n 0.00714857f $X=14.495 $Y=1.665
+ $X2=0 $Y2=0
cc_583 N_A_545_87#_c_613_n N_A_2403_74#_c_1729_n 0.00647787f $X=14.64 $Y=1.665
+ $X2=0 $Y2=0
cc_584 N_A_545_87#_c_614_n N_A_2403_74#_c_1729_n 0.0187409f $X=14.64 $Y=1.665
+ $X2=0 $Y2=0
cc_585 N_A_545_87#_c_595_n N_A_2403_74#_c_1730_n 0.00135428f $X=14.31 $Y=1.55
+ $X2=0 $Y2=0
cc_586 N_A_545_87#_c_596_n N_A_2403_74#_c_1730_n 0.00171167f $X=14.17 $Y=0.58
+ $X2=0 $Y2=0
cc_587 N_A_545_87#_c_606_n N_A_2403_74#_c_1744_n 9.56764e-19 $X=14.21 $Y=2.465
+ $X2=0 $Y2=0
cc_588 N_A_545_87#_c_607_n N_A_2403_74#_c_1744_n 0.00175174f $X=14.31 $Y=2.18
+ $X2=0 $Y2=0
cc_589 N_A_545_87#_c_609_n N_A_2403_74#_c_1744_n 3.36721e-19 $X=14.22 $Y=2.265
+ $X2=0 $Y2=0
cc_590 N_A_545_87#_c_613_n N_A_2403_74#_c_1744_n 3.62444e-19 $X=14.64 $Y=1.665
+ $X2=0 $Y2=0
cc_591 N_A_545_87#_c_614_n N_A_2403_74#_c_1744_n 2.99261e-19 $X=14.64 $Y=1.665
+ $X2=0 $Y2=0
cc_592 N_A_545_87#_c_613_n N_A_2403_74#_c_1734_n 0.00243858f $X=14.64 $Y=1.665
+ $X2=0 $Y2=0
cc_593 N_A_545_87#_c_614_n N_A_2403_74#_c_1734_n 0.00203152f $X=14.64 $Y=1.665
+ $X2=0 $Y2=0
cc_594 N_A_545_87#_c_591_n N_A_2403_74#_c_1735_n 0.00177547f $X=12.805 $Y=0.865
+ $X2=0 $Y2=0
cc_595 N_A_545_87#_c_591_n N_A_2403_74#_c_1736_n 0.00387158f $X=12.805 $Y=0.865
+ $X2=0 $Y2=0
cc_596 N_A_545_87#_c_592_n N_A_2403_74#_c_1736_n 0.0231504f $X=13.335 $Y=0.94
+ $X2=0 $Y2=0
cc_597 N_A_545_87#_c_593_n N_A_2403_74#_c_1736_n 0.00439386f $X=12.88 $Y=0.94
+ $X2=0 $Y2=0
cc_598 N_A_545_87#_c_595_n N_A_2403_74#_c_1736_n 0.00315267f $X=14.31 $Y=1.55
+ $X2=0 $Y2=0
cc_599 N_A_545_87#_c_596_n N_A_2403_74#_c_1736_n 0.00413501f $X=14.17 $Y=0.58
+ $X2=0 $Y2=0
cc_600 N_A_545_87#_c_597_n N_A_2403_74#_c_1736_n 0.00608858f $X=14.495 $Y=1.665
+ $X2=0 $Y2=0
cc_601 N_A_545_87#_c_603_n N_A_2403_74#_c_1749_n 0.00312272f $X=13.275 $Y=2.465
+ $X2=0 $Y2=0
cc_602 N_A_545_87#_c_608_n N_A_2403_74#_c_1749_n 0.0119401f $X=13.485 $Y=2.222
+ $X2=0 $Y2=0
cc_603 N_A_545_87#_c_603_n N_A_2403_74#_c_1750_n 0.00288406f $X=13.275 $Y=2.465
+ $X2=0 $Y2=0
cc_604 N_A_545_87#_c_608_n N_A_2403_74#_c_1750_n 0.00761573f $X=13.485 $Y=2.222
+ $X2=0 $Y2=0
cc_605 N_A_545_87#_c_597_n N_A_2403_74#_c_1750_n 0.0147772f $X=14.495 $Y=1.665
+ $X2=0 $Y2=0
cc_606 N_A_545_87#_c_603_n N_A_2403_74#_c_1751_n 3.41912e-19 $X=13.275 $Y=2.465
+ $X2=0 $Y2=0
cc_607 N_A_545_87#_c_594_n N_A_2403_74#_c_1751_n 6.56155e-19 $X=13.41 $Y=2.05
+ $X2=0 $Y2=0
cc_608 N_A_545_87#_c_608_n N_A_2403_74#_c_1751_n 0.0024169f $X=13.485 $Y=2.222
+ $X2=0 $Y2=0
cc_609 N_A_545_87#_c_597_n N_A_2403_74#_c_1751_n 0.0112472f $X=14.495 $Y=1.665
+ $X2=0 $Y2=0
cc_610 N_A_545_87#_c_603_n N_A_2403_74#_c_1752_n 0.00200844f $X=13.275 $Y=2.465
+ $X2=0 $Y2=0
cc_611 N_A_545_87#_c_594_n N_A_2403_74#_c_1752_n 0.00928497f $X=13.41 $Y=2.05
+ $X2=0 $Y2=0
cc_612 N_A_545_87#_c_605_n N_A_2403_74#_c_1752_n 0.0356642f $X=14.045 $Y=2.265
+ $X2=0 $Y2=0
cc_613 N_A_545_87#_c_607_n N_A_2403_74#_c_1752_n 0.0164589f $X=14.31 $Y=2.18
+ $X2=0 $Y2=0
cc_614 N_A_545_87#_c_608_n N_A_2403_74#_c_1752_n 0.0166089f $X=13.485 $Y=2.222
+ $X2=0 $Y2=0
cc_615 N_A_545_87#_c_609_n N_A_2403_74#_c_1752_n 7.31419e-19 $X=14.22 $Y=2.265
+ $X2=0 $Y2=0
cc_616 N_A_545_87#_c_610_n N_A_2403_74#_c_1752_n 0.00210074f $X=14.31 $Y=1.665
+ $X2=0 $Y2=0
cc_617 N_A_545_87#_c_594_n N_A_2403_74#_c_1738_n 0.02408f $X=13.41 $Y=2.05 $X2=0
+ $Y2=0
cc_618 N_A_545_87#_c_595_n N_A_2403_74#_c_1738_n 0.0414257f $X=14.31 $Y=1.55
+ $X2=0 $Y2=0
cc_619 N_A_545_87#_c_610_n N_A_2403_74#_c_1738_n 0.0146426f $X=14.31 $Y=1.665
+ $X2=0 $Y2=0
cc_620 N_A_545_87#_c_597_n N_A_2403_74#_c_1738_n 0.0712682f $X=14.495 $Y=1.665
+ $X2=0 $Y2=0
cc_621 N_A_545_87#_c_613_n N_A_2403_74#_c_1738_n 2.75883e-19 $X=14.64 $Y=1.665
+ $X2=0 $Y2=0
cc_622 N_A_545_87#_c_592_n N_A_2403_74#_c_1739_n 0.0275433f $X=13.335 $Y=0.94
+ $X2=0 $Y2=0
cc_623 N_A_545_87#_c_595_n N_A_2403_74#_c_1739_n 0.00959895f $X=14.31 $Y=1.55
+ $X2=0 $Y2=0
cc_624 N_A_545_87#_c_596_n N_A_2403_74#_c_1739_n 0.00110885f $X=14.17 $Y=0.58
+ $X2=0 $Y2=0
cc_625 N_A_545_87#_c_605_n N_A_2403_74#_c_1740_n 0.00115499f $X=14.045 $Y=2.265
+ $X2=0 $Y2=0
cc_626 N_A_545_87#_c_607_n N_A_2403_74#_c_1740_n 0.0116068f $X=14.31 $Y=2.18
+ $X2=0 $Y2=0
cc_627 N_A_545_87#_c_610_n N_A_2403_74#_c_1740_n 0.00204394f $X=14.31 $Y=1.665
+ $X2=0 $Y2=0
cc_628 N_A_545_87#_c_597_n N_A_2403_74#_c_1740_n 0.00191903f $X=14.495 $Y=1.665
+ $X2=0 $Y2=0
cc_629 N_A_545_87#_c_602_n N_A_37_464#_c_1923_n 0.0133663f $X=3.175 $Y=2.24
+ $X2=0 $Y2=0
cc_630 N_A_545_87#_c_597_n N_A_37_464#_c_1923_n 0.00606879f $X=14.495 $Y=1.665
+ $X2=0 $Y2=0
cc_631 N_A_545_87#_c_598_n N_A_37_464#_c_1923_n 0.00281723f $X=2.785 $Y=1.665
+ $X2=0 $Y2=0
cc_632 N_A_545_87#_c_599_n N_A_37_464#_c_1923_n 0.0161246f $X=2.89 $Y=1.685
+ $X2=0 $Y2=0
cc_633 N_A_545_87#_c_600_n N_A_37_464#_c_1923_n 0.00461297f $X=3.175 $Y=1.685
+ $X2=0 $Y2=0
cc_634 N_A_545_87#_M1023_g N_A_37_464#_c_1913_n 0.0139537f $X=2.8 $Y=0.775 $X2=0
+ $Y2=0
cc_635 N_A_545_87#_c_602_n N_A_37_464#_c_1925_n 0.00870642f $X=3.175 $Y=2.24
+ $X2=0 $Y2=0
cc_636 N_A_545_87#_M1023_g N_A_37_464#_c_1914_n 0.004494f $X=2.8 $Y=0.775 $X2=0
+ $Y2=0
cc_637 N_A_545_87#_c_602_n N_A_37_464#_c_1914_n 0.00116727f $X=3.175 $Y=2.24
+ $X2=0 $Y2=0
cc_638 N_A_545_87#_c_597_n N_A_37_464#_c_1914_n 0.0171244f $X=14.495 $Y=1.665
+ $X2=0 $Y2=0
cc_639 N_A_545_87#_c_598_n N_A_37_464#_c_1914_n 3.93276e-19 $X=2.785 $Y=1.665
+ $X2=0 $Y2=0
cc_640 N_A_545_87#_c_599_n N_A_37_464#_c_1914_n 0.0163889f $X=2.89 $Y=1.685
+ $X2=0 $Y2=0
cc_641 N_A_545_87#_c_600_n N_A_37_464#_c_1914_n 0.0182371f $X=3.175 $Y=1.685
+ $X2=0 $Y2=0
cc_642 N_A_545_87#_M1023_g N_A_37_464#_c_1916_n 0.00714755f $X=2.8 $Y=0.775
+ $X2=0 $Y2=0
cc_643 N_A_545_87#_c_597_n N_A_37_464#_c_1916_n 0.012122f $X=14.495 $Y=1.665
+ $X2=0 $Y2=0
cc_644 N_A_545_87#_c_599_n N_A_37_464#_c_1916_n 0.0137413f $X=2.89 $Y=1.685
+ $X2=0 $Y2=0
cc_645 N_A_545_87#_c_600_n N_A_37_464#_c_1916_n 0.0105002f $X=3.175 $Y=1.685
+ $X2=0 $Y2=0
cc_646 N_A_545_87#_c_602_n N_A_37_464#_c_1928_n 0.00166465f $X=3.175 $Y=2.24
+ $X2=0 $Y2=0
cc_647 N_A_545_87#_c_597_n N_A_37_464#_c_1928_n 0.00276825f $X=14.495 $Y=1.665
+ $X2=0 $Y2=0
cc_648 N_A_545_87#_c_605_n N_VPWR_M1035_d 0.00295338f $X=14.045 $Y=2.265 $X2=0
+ $Y2=0
cc_649 N_A_545_87#_c_602_n N_VPWR_c_2039_n 0.00150486f $X=3.175 $Y=2.24 $X2=0
+ $Y2=0
cc_650 N_A_545_87#_c_603_n N_VPWR_c_2045_n 0.0184894f $X=13.275 $Y=2.465 $X2=0
+ $Y2=0
cc_651 N_A_545_87#_c_606_n N_VPWR_c_2045_n 0.013346f $X=14.21 $Y=2.465 $X2=0
+ $Y2=0
cc_652 N_A_545_87#_c_608_n N_VPWR_c_2045_n 0.0259876f $X=13.485 $Y=2.222 $X2=0
+ $Y2=0
cc_653 N_A_545_87#_c_606_n N_VPWR_c_2046_n 0.0154862f $X=14.21 $Y=2.465 $X2=0
+ $Y2=0
cc_654 N_A_545_87#_c_606_n N_VPWR_c_2047_n 0.0526516f $X=14.21 $Y=2.465 $X2=0
+ $Y2=0
cc_655 N_A_545_87#_c_607_n N_VPWR_c_2047_n 0.0181977f $X=14.31 $Y=2.18 $X2=0
+ $Y2=0
cc_656 N_A_545_87#_c_609_n N_VPWR_c_2047_n 0.0150382f $X=14.22 $Y=2.265 $X2=0
+ $Y2=0
cc_657 N_A_545_87#_c_613_n N_VPWR_c_2047_n 0.00645519f $X=14.64 $Y=1.665 $X2=0
+ $Y2=0
cc_658 N_A_545_87#_c_614_n N_VPWR_c_2047_n 0.0137154f $X=14.64 $Y=1.665 $X2=0
+ $Y2=0
cc_659 N_A_545_87#_c_602_n N_VPWR_c_2055_n 0.0044174f $X=3.175 $Y=2.24 $X2=0
+ $Y2=0
cc_660 N_A_545_87#_c_603_n N_VPWR_c_2059_n 0.00413917f $X=13.275 $Y=2.465 $X2=0
+ $Y2=0
cc_661 N_A_545_87#_c_602_n N_VPWR_c_2037_n 0.00544287f $X=3.175 $Y=2.24 $X2=0
+ $Y2=0
cc_662 N_A_545_87#_c_603_n N_VPWR_c_2037_n 0.00852225f $X=13.275 $Y=2.465 $X2=0
+ $Y2=0
cc_663 N_A_545_87#_c_606_n N_VPWR_c_2037_n 0.0127853f $X=14.21 $Y=2.465 $X2=0
+ $Y2=0
cc_664 N_A_545_87#_c_597_n N_A_661_113#_c_2241_n 0.00390489f $X=14.495 $Y=1.665
+ $X2=0 $Y2=0
cc_665 N_A_545_87#_c_602_n N_A_661_113#_c_2253_n 5.18926e-19 $X=3.175 $Y=2.24
+ $X2=0 $Y2=0
cc_666 N_A_545_87#_c_597_n N_A_661_113#_c_2234_n 0.0143992f $X=14.495 $Y=1.665
+ $X2=0 $Y2=0
cc_667 N_A_545_87#_c_597_n N_A_661_113#_c_2245_n 0.0221561f $X=14.495 $Y=1.665
+ $X2=0 $Y2=0
cc_668 N_A_545_87#_c_597_n N_A_661_113#_c_2246_n 0.0136971f $X=14.495 $Y=1.665
+ $X2=0 $Y2=0
cc_669 N_A_545_87#_c_597_n N_A_661_113#_c_2235_n 0.0282403f $X=14.495 $Y=1.665
+ $X2=0 $Y2=0
cc_670 N_A_545_87#_c_597_n N_A_661_113#_c_2236_n 0.00557308f $X=14.495 $Y=1.665
+ $X2=0 $Y2=0
cc_671 N_A_545_87#_c_597_n N_A_661_113#_c_2247_n 0.00423412f $X=14.495 $Y=1.665
+ $X2=0 $Y2=0
cc_672 N_A_545_87#_c_597_n N_A_661_113#_c_2238_n 0.00594784f $X=14.495 $Y=1.665
+ $X2=0 $Y2=0
cc_673 N_A_545_87#_c_597_n N_A_661_113#_c_2239_n 0.0169423f $X=14.495 $Y=1.665
+ $X2=0 $Y2=0
cc_674 N_A_545_87#_c_597_n N_A_661_113#_c_2240_n 0.00894617f $X=14.495 $Y=1.665
+ $X2=0 $Y2=0
cc_675 N_A_545_87#_c_597_n N_A_661_113#_c_2250_n 0.00101595f $X=14.495 $Y=1.665
+ $X2=0 $Y2=0
cc_676 N_A_545_87#_c_597_n N_A_661_113#_c_2251_n 0.00600127f $X=14.495 $Y=1.665
+ $X2=0 $Y2=0
cc_677 N_A_545_87#_c_607_n Q 0.00220553f $X=14.31 $Y=2.18 $X2=0 $Y2=0
cc_678 N_A_545_87#_c_613_n Q 0.00608382f $X=14.64 $Y=1.665 $X2=0 $Y2=0
cc_679 N_A_545_87#_c_614_n Q 0.00604625f $X=14.64 $Y=1.665 $X2=0 $Y2=0
cc_680 N_A_545_87#_M1023_g N_VGND_c_2468_n 0.0018473f $X=2.8 $Y=0.775 $X2=0
+ $Y2=0
cc_681 N_A_545_87#_c_597_n N_VGND_c_2469_n 0.00662369f $X=14.495 $Y=1.665 $X2=0
+ $Y2=0
cc_682 N_A_545_87#_c_596_n N_VGND_c_2474_n 0.0169737f $X=14.17 $Y=0.58 $X2=0
+ $Y2=0
cc_683 N_A_545_87#_c_596_n N_VGND_c_2475_n 0.0807764f $X=14.17 $Y=0.58 $X2=0
+ $Y2=0
cc_684 N_A_545_87#_c_613_n N_VGND_c_2475_n 0.00547886f $X=14.64 $Y=1.665 $X2=0
+ $Y2=0
cc_685 N_A_545_87#_c_614_n N_VGND_c_2475_n 0.0106518f $X=14.64 $Y=1.665 $X2=0
+ $Y2=0
cc_686 N_A_545_87#_M1023_g N_VGND_c_2485_n 0.00430863f $X=2.8 $Y=0.775 $X2=0
+ $Y2=0
cc_687 N_A_545_87#_c_591_n N_VGND_c_2495_n 0.00383152f $X=12.805 $Y=0.865 $X2=0
+ $Y2=0
cc_688 N_A_545_87#_c_591_n N_VGND_c_2496_n 0.0115585f $X=12.805 $Y=0.865 $X2=0
+ $Y2=0
cc_689 N_A_545_87#_c_592_n N_VGND_c_2496_n 0.00552448f $X=13.335 $Y=0.94 $X2=0
+ $Y2=0
cc_690 N_A_545_87#_c_596_n N_VGND_c_2496_n 0.0136104f $X=14.17 $Y=0.58 $X2=0
+ $Y2=0
cc_691 N_A_545_87#_M1023_g N_VGND_c_2499_n 0.00486331f $X=2.8 $Y=0.775 $X2=0
+ $Y2=0
cc_692 N_A_545_87#_c_591_n N_VGND_c_2499_n 0.00384101f $X=12.805 $Y=0.865 $X2=0
+ $Y2=0
cc_693 N_A_545_87#_c_596_n N_VGND_c_2499_n 0.0141105f $X=14.17 $Y=0.58 $X2=0
+ $Y2=0
cc_694 N_A_631_87#_c_843_n N_SCD_c_949_n 0.0255091f $X=5.745 $Y=1.92 $X2=0 $Y2=0
cc_695 N_A_631_87#_c_847_n N_SCD_c_949_n 0.01197f $X=5.58 $Y=2 $X2=0 $Y2=0
cc_696 N_A_631_87#_c_842_n N_SCD_c_950_n 0.0438474f $X=5.67 $Y=2.2 $X2=0 $Y2=0
cc_697 N_A_631_87#_c_847_n SCD 0.0294802f $X=5.58 $Y=2 $X2=0 $Y2=0
cc_698 N_A_631_87#_c_839_n SCD 0.0193335f $X=5.745 $Y=1.58 $X2=0 $Y2=0
cc_699 N_A_631_87#_c_840_n SCD 0.00113695f $X=5.745 $Y=1.58 $X2=0 $Y2=0
cc_700 N_A_631_87#_c_847_n N_SCD_c_948_n 0.00104612f $X=5.58 $Y=2 $X2=0 $Y2=0
cc_701 N_A_631_87#_c_839_n N_SCD_c_948_n 0.00227836f $X=5.745 $Y=1.58 $X2=0
+ $Y2=0
cc_702 N_A_631_87#_c_840_n N_SCD_c_948_n 0.0255091f $X=5.745 $Y=1.58 $X2=0 $Y2=0
cc_703 N_A_631_87#_c_846_n N_SCE_c_999_n 3.50071e-19 $X=4.19 $Y=2.255 $X2=-0.19
+ $Y2=-0.245
cc_704 N_A_631_87#_c_850_n N_SCE_c_999_n 0.00100796f $X=4.375 $Y=2.495 $X2=-0.19
+ $Y2=-0.245
cc_705 N_A_631_87#_c_850_n N_SCE_c_1000_n 0.00201936f $X=4.375 $Y=2.495 $X2=0
+ $Y2=0
cc_706 N_A_631_87#_c_837_n N_SCE_c_992_n 0.0076784f $X=4.08 $Y=1.78 $X2=0 $Y2=0
cc_707 N_A_631_87#_c_838_n N_SCE_c_992_n 0.020518f $X=4.08 $Y=1.78 $X2=0 $Y2=0
cc_708 N_A_631_87#_c_846_n N_SCE_c_992_n 0.00371596f $X=4.19 $Y=2.255 $X2=0
+ $Y2=0
cc_709 N_A_631_87#_c_847_n N_SCE_c_992_n 0.0189076f $X=5.58 $Y=2 $X2=0 $Y2=0
cc_710 N_A_631_87#_c_846_n N_SCE_M1044_g 0.00171259f $X=4.19 $Y=2.255 $X2=0
+ $Y2=0
cc_711 N_A_631_87#_c_850_n N_SCE_M1044_g 0.00320341f $X=4.375 $Y=2.495 $X2=0
+ $Y2=0
cc_712 N_A_631_87#_c_835_n N_SCE_M1045_g 0.00263665f $X=4.08 $Y=0.42 $X2=0 $Y2=0
cc_713 N_A_631_87#_c_836_n N_SCE_M1045_g 0.0198324f $X=4.08 $Y=0.42 $X2=0 $Y2=0
cc_714 N_A_631_87#_c_837_n N_SCE_M1045_g 0.0032212f $X=4.08 $Y=1.78 $X2=0 $Y2=0
cc_715 N_A_631_87#_c_841_n N_SCE_M1045_g 2.28678e-19 $X=4.5 $Y=0.805 $X2=0 $Y2=0
cc_716 N_A_631_87#_c_834_n SCE 0.00100831f $X=4.08 $Y=1.135 $X2=0 $Y2=0
cc_717 N_A_631_87#_c_837_n SCE 0.027154f $X=4.08 $Y=1.78 $X2=0 $Y2=0
cc_718 N_A_631_87#_c_847_n SCE 0.00626904f $X=5.58 $Y=2 $X2=0 $Y2=0
cc_719 N_A_631_87#_c_841_n SCE 0.0107055f $X=4.5 $Y=0.805 $X2=0 $Y2=0
cc_720 N_A_631_87#_c_834_n N_SCE_c_998_n 0.0213991f $X=4.08 $Y=1.135 $X2=0 $Y2=0
cc_721 N_A_631_87#_c_837_n N_SCE_c_998_n 0.00101987f $X=4.08 $Y=1.78 $X2=0 $Y2=0
cc_722 N_A_631_87#_c_847_n N_SCE_c_998_n 0.00328462f $X=5.58 $Y=2 $X2=0 $Y2=0
cc_723 N_A_631_87#_c_841_n N_SCE_c_998_n 0.00326781f $X=4.5 $Y=0.805 $X2=0 $Y2=0
cc_724 N_A_631_87#_c_840_n N_CLK_c_1081_n 0.00882105f $X=5.745 $Y=1.58 $X2=0
+ $Y2=0
cc_725 N_A_631_87#_c_831_n N_A_37_464#_c_1913_n 0.0119582f $X=3.23 $Y=1.06 $X2=0
+ $Y2=0
cc_726 N_A_631_87#_c_833_n N_A_37_464#_c_1913_n 0.00456059f $X=3.305 $Y=1.135
+ $X2=0 $Y2=0
cc_727 N_A_631_87#_c_832_n N_A_37_464#_c_1914_n 9.40513e-19 $X=3.915 $Y=1.135
+ $X2=0 $Y2=0
cc_728 N_A_631_87#_c_832_n N_A_37_464#_c_1916_n 0.00739581f $X=3.915 $Y=1.135
+ $X2=0 $Y2=0
cc_729 N_A_631_87#_c_833_n N_A_37_464#_c_1916_n 0.00806291f $X=3.305 $Y=1.135
+ $X2=0 $Y2=0
cc_730 N_A_631_87#_c_842_n N_VPWR_c_2040_n 0.00149083f $X=5.67 $Y=2.2 $X2=0
+ $Y2=0
cc_731 N_A_631_87#_c_842_n N_VPWR_c_2041_n 0.00329869f $X=5.67 $Y=2.2 $X2=0
+ $Y2=0
cc_732 N_A_631_87#_c_842_n N_VPWR_c_2056_n 0.00530811f $X=5.67 $Y=2.2 $X2=0
+ $Y2=0
cc_733 N_A_631_87#_c_842_n N_VPWR_c_2037_n 0.005315f $X=5.67 $Y=2.2 $X2=0 $Y2=0
cc_734 N_A_631_87#_c_838_n N_A_661_113#_c_2241_n 7.59117e-19 $X=4.08 $Y=1.78
+ $X2=0 $Y2=0
cc_735 N_A_631_87#_c_850_n N_A_661_113#_c_2241_n 0.0358182f $X=4.375 $Y=2.495
+ $X2=0 $Y2=0
cc_736 N_A_631_87#_M1044_s N_A_661_113#_c_2242_n 0.00259631f $X=4.245 $Y=2.275
+ $X2=0 $Y2=0
cc_737 N_A_631_87#_c_850_n N_A_661_113#_c_2242_n 0.0265612f $X=4.375 $Y=2.495
+ $X2=0 $Y2=0
cc_738 N_A_631_87#_c_850_n N_A_661_113#_c_2269_n 0.0230808f $X=4.375 $Y=2.495
+ $X2=0 $Y2=0
cc_739 N_A_631_87#_c_847_n N_A_661_113#_c_2243_n 0.0134263f $X=5.58 $Y=2 $X2=0
+ $Y2=0
cc_740 N_A_631_87#_c_850_n N_A_661_113#_c_2243_n 0.0140999f $X=4.375 $Y=2.495
+ $X2=0 $Y2=0
cc_741 N_A_631_87#_c_842_n N_A_661_113#_c_2234_n 0.00165009f $X=5.67 $Y=2.2
+ $X2=0 $Y2=0
cc_742 N_A_631_87#_c_843_n N_A_661_113#_c_2234_n 0.00361138f $X=5.745 $Y=1.92
+ $X2=0 $Y2=0
cc_743 N_A_631_87#_c_847_n N_A_661_113#_c_2234_n 0.0135427f $X=5.58 $Y=2 $X2=0
+ $Y2=0
cc_744 N_A_631_87#_c_839_n N_A_661_113#_c_2234_n 0.0361817f $X=5.745 $Y=1.58
+ $X2=0 $Y2=0
cc_745 N_A_631_87#_c_840_n N_A_661_113#_c_2234_n 0.00703953f $X=5.745 $Y=1.58
+ $X2=0 $Y2=0
cc_746 N_A_631_87#_c_831_n N_A_661_113#_c_2238_n 0.00274432f $X=3.23 $Y=1.06
+ $X2=0 $Y2=0
cc_747 N_A_631_87#_c_832_n N_A_661_113#_c_2238_n 0.0107113f $X=3.915 $Y=1.135
+ $X2=0 $Y2=0
cc_748 N_A_631_87#_c_836_n N_A_661_113#_c_2238_n 0.00400614f $X=4.08 $Y=0.42
+ $X2=0 $Y2=0
cc_749 N_A_631_87#_c_841_n N_A_661_113#_c_2238_n 0.0281364f $X=4.5 $Y=0.805
+ $X2=0 $Y2=0
cc_750 N_A_631_87#_c_831_n N_A_661_113#_c_2239_n 4.67525e-19 $X=3.23 $Y=1.06
+ $X2=0 $Y2=0
cc_751 N_A_631_87#_c_832_n N_A_661_113#_c_2239_n 0.0142405f $X=3.915 $Y=1.135
+ $X2=0 $Y2=0
cc_752 N_A_631_87#_c_836_n N_A_661_113#_c_2239_n 7.07121e-19 $X=4.08 $Y=0.42
+ $X2=0 $Y2=0
cc_753 N_A_631_87#_c_837_n N_A_661_113#_c_2239_n 0.0656047f $X=4.08 $Y=1.78
+ $X2=0 $Y2=0
cc_754 N_A_631_87#_c_838_n N_A_661_113#_c_2239_n 0.0123483f $X=4.08 $Y=1.78
+ $X2=0 $Y2=0
cc_755 N_A_631_87#_c_846_n N_A_661_113#_c_2239_n 0.00902514f $X=4.19 $Y=2.255
+ $X2=0 $Y2=0
cc_756 N_A_631_87#_c_849_n N_A_661_113#_c_2239_n 0.0142217f $X=4.135 $Y=2 $X2=0
+ $Y2=0
cc_757 N_A_631_87#_c_850_n N_A_661_113#_c_2239_n 0.00217874f $X=4.375 $Y=2.495
+ $X2=0 $Y2=0
cc_758 N_A_631_87#_c_847_n N_A_661_113#_c_2240_n 2.73581e-19 $X=5.58 $Y=2 $X2=0
+ $Y2=0
cc_759 N_A_631_87#_c_839_n N_A_661_113#_c_2240_n 0.0209662f $X=5.745 $Y=1.58
+ $X2=0 $Y2=0
cc_760 N_A_631_87#_c_840_n N_A_661_113#_c_2240_n 0.00403118f $X=5.745 $Y=1.58
+ $X2=0 $Y2=0
cc_761 N_A_631_87#_c_842_n N_A_661_113#_c_2249_n 0.0076275f $X=5.67 $Y=2.2 $X2=0
+ $Y2=0
cc_762 N_A_631_87#_c_842_n N_A_661_113#_c_2250_n 0.011357f $X=5.67 $Y=2.2 $X2=0
+ $Y2=0
cc_763 N_A_631_87#_c_843_n N_A_661_113#_c_2250_n 4.52395e-19 $X=5.745 $Y=1.92
+ $X2=0 $Y2=0
cc_764 N_A_631_87#_c_847_n N_A_661_113#_c_2250_n 0.0769068f $X=5.58 $Y=2 $X2=0
+ $Y2=0
cc_765 N_A_631_87#_c_842_n N_A_661_113#_c_2251_n 0.00236127f $X=5.67 $Y=2.2
+ $X2=0 $Y2=0
cc_766 N_A_631_87#_c_843_n N_A_661_113#_c_2251_n 0.0033091f $X=5.745 $Y=1.92
+ $X2=0 $Y2=0
cc_767 N_A_631_87#_c_835_n N_VGND_c_2469_n 0.0123486f $X=4.08 $Y=0.42 $X2=0
+ $Y2=0
cc_768 N_A_631_87#_c_836_n N_VGND_c_2469_n 6.24286e-19 $X=4.08 $Y=0.42 $X2=0
+ $Y2=0
cc_769 N_A_631_87#_c_841_n N_VGND_c_2469_n 0.0152974f $X=4.5 $Y=0.805 $X2=0
+ $Y2=0
cc_770 N_A_631_87#_c_831_n N_VGND_c_2485_n 0.00430863f $X=3.23 $Y=1.06 $X2=0
+ $Y2=0
cc_771 N_A_631_87#_c_835_n N_VGND_c_2485_n 0.0181716f $X=4.08 $Y=0.42 $X2=0
+ $Y2=0
cc_772 N_A_631_87#_c_836_n N_VGND_c_2485_n 0.00466976f $X=4.08 $Y=0.42 $X2=0
+ $Y2=0
cc_773 N_A_631_87#_c_841_n N_VGND_c_2485_n 0.00645779f $X=4.5 $Y=0.805 $X2=0
+ $Y2=0
cc_774 N_A_631_87#_c_831_n N_VGND_c_2499_n 0.00486331f $X=3.23 $Y=1.06 $X2=0
+ $Y2=0
cc_775 N_A_631_87#_c_835_n N_VGND_c_2499_n 0.0104851f $X=4.08 $Y=0.42 $X2=0
+ $Y2=0
cc_776 N_A_631_87#_c_836_n N_VGND_c_2499_n 0.00292172f $X=4.08 $Y=0.42 $X2=0
+ $Y2=0
cc_777 N_A_631_87#_c_841_n N_VGND_c_2499_n 0.00945185f $X=4.5 $Y=0.805 $X2=0
+ $Y2=0
cc_778 N_SCD_c_950_n N_SCE_c_1000_n 0.00100522f $X=5.28 $Y=2.2 $X2=0 $Y2=0
cc_779 N_SCD_c_949_n N_SCE_c_992_n 0.00601231f $X=5.28 $Y=2.11 $X2=0 $Y2=0
cc_780 SCD N_SCE_c_992_n 0.00432722f $X=4.955 $Y=1.21 $X2=0 $Y2=0
cc_781 N_SCD_c_948_n N_SCE_c_992_n 0.00806113f $X=5.205 $Y=1.58 $X2=0 $Y2=0
cc_782 N_SCD_c_950_n N_SCE_c_1003_n 0.00601231f $X=5.28 $Y=2.2 $X2=0 $Y2=0
cc_783 N_SCD_c_950_n N_SCE_M1044_g 0.0111767f $X=5.28 $Y=2.2 $X2=0 $Y2=0
cc_784 N_SCD_M1011_g N_SCE_M1045_g 0.0249668f $X=5.145 $Y=0.835 $X2=0 $Y2=0
cc_785 N_SCD_M1011_g N_SCE_c_994_n 0.00894529f $X=5.145 $Y=0.835 $X2=0 $Y2=0
cc_786 N_SCD_M1011_g N_SCE_M1003_g 0.0397856f $X=5.145 $Y=0.835 $X2=0 $Y2=0
cc_787 N_SCD_M1011_g SCE 2.44439e-19 $X=5.145 $Y=0.835 $X2=0 $Y2=0
cc_788 SCD SCE 0.0266241f $X=4.955 $Y=1.21 $X2=0 $Y2=0
cc_789 SCD N_SCE_c_998_n 0.00222986f $X=4.955 $Y=1.21 $X2=0 $Y2=0
cc_790 N_SCD_c_948_n N_SCE_c_998_n 0.00474864f $X=5.205 $Y=1.58 $X2=0 $Y2=0
cc_791 N_SCD_c_950_n N_VPWR_c_2040_n 0.00959399f $X=5.28 $Y=2.2 $X2=0 $Y2=0
cc_792 N_SCD_c_950_n N_VPWR_c_2056_n 0.00489294f $X=5.28 $Y=2.2 $X2=0 $Y2=0
cc_793 N_SCD_c_950_n N_VPWR_c_2037_n 0.00481893f $X=5.28 $Y=2.2 $X2=0 $Y2=0
cc_794 N_SCD_c_950_n N_A_661_113#_c_2242_n 3.76568e-19 $X=5.28 $Y=2.2 $X2=0
+ $Y2=0
cc_795 N_SCD_c_950_n N_A_661_113#_c_2269_n 0.00283455f $X=5.28 $Y=2.2 $X2=0
+ $Y2=0
cc_796 N_SCD_M1011_g N_A_661_113#_c_2233_n 0.00142836f $X=5.145 $Y=0.835 $X2=0
+ $Y2=0
cc_797 SCD N_A_661_113#_c_2234_n 0.00532608f $X=4.955 $Y=1.21 $X2=0 $Y2=0
cc_798 N_SCD_M1011_g N_A_661_113#_c_2240_n 0.00101742f $X=5.145 $Y=0.835 $X2=0
+ $Y2=0
cc_799 SCD N_A_661_113#_c_2240_n 0.0053986f $X=4.955 $Y=1.21 $X2=0 $Y2=0
cc_800 N_SCD_c_950_n N_A_661_113#_c_2249_n 0.00138942f $X=5.28 $Y=2.2 $X2=0
+ $Y2=0
cc_801 N_SCD_c_950_n N_A_661_113#_c_2250_n 0.0160628f $X=5.28 $Y=2.2 $X2=0 $Y2=0
cc_802 N_SCD_c_950_n N_A_661_113#_c_2251_n 3.80333e-19 $X=5.28 $Y=2.2 $X2=0
+ $Y2=0
cc_803 N_SCD_M1011_g N_VGND_c_2469_n 0.0105685f $X=5.145 $Y=0.835 $X2=0 $Y2=0
cc_804 SCD N_VGND_c_2469_n 0.00958749f $X=4.955 $Y=1.21 $X2=0 $Y2=0
cc_805 N_SCD_M1011_g N_VGND_c_2499_n 7.97988e-19 $X=5.145 $Y=0.835 $X2=0 $Y2=0
cc_806 N_SCE_c_999_n N_A_37_464#_c_1925_n 0.00161473f $X=3.625 $Y=3.03 $X2=0
+ $Y2=0
cc_807 N_SCE_c_999_n N_A_37_464#_c_1914_n 7.32247e-19 $X=3.625 $Y=3.03 $X2=0
+ $Y2=0
cc_808 N_SCE_c_999_n N_A_37_464#_c_1928_n 7.52181e-19 $X=3.625 $Y=3.03 $X2=0
+ $Y2=0
cc_809 N_SCE_c_1000_n N_VPWR_c_2040_n 0.00310923f $X=4.51 $Y=3.105 $X2=0 $Y2=0
cc_810 N_SCE_M1044_g N_VPWR_c_2040_n 0.00117443f $X=4.6 $Y=2.595 $X2=0 $Y2=0
cc_811 N_SCE_c_1001_n N_VPWR_c_2055_n 0.0240584f $X=3.7 $Y=3.105 $X2=0 $Y2=0
cc_812 N_SCE_c_1000_n N_VPWR_c_2037_n 0.0252128f $X=4.51 $Y=3.105 $X2=0 $Y2=0
cc_813 N_SCE_c_1001_n N_VPWR_c_2037_n 0.0100661f $X=3.7 $Y=3.105 $X2=0 $Y2=0
cc_814 N_SCE_c_999_n N_A_661_113#_c_2241_n 0.00196983f $X=3.625 $Y=3.03 $X2=0
+ $Y2=0
cc_815 N_SCE_M1044_g N_A_661_113#_c_2241_n 0.00450557f $X=4.6 $Y=2.595 $X2=0
+ $Y2=0
cc_816 N_SCE_c_999_n N_A_661_113#_c_2309_n 0.00538071f $X=3.625 $Y=3.03 $X2=0
+ $Y2=0
cc_817 N_SCE_c_1000_n N_A_661_113#_c_2242_n 0.0217336f $X=4.51 $Y=3.105 $X2=0
+ $Y2=0
cc_818 N_SCE_M1044_g N_A_661_113#_c_2242_n 0.00872278f $X=4.6 $Y=2.595 $X2=0
+ $Y2=0
cc_819 N_SCE_c_999_n N_A_661_113#_c_2253_n 0.00373701f $X=3.625 $Y=3.03 $X2=0
+ $Y2=0
cc_820 N_SCE_c_1000_n N_A_661_113#_c_2253_n 0.00837949f $X=4.51 $Y=3.105 $X2=0
+ $Y2=0
cc_821 N_SCE_c_1001_n N_A_661_113#_c_2253_n 0.0013142f $X=3.7 $Y=3.105 $X2=0
+ $Y2=0
cc_822 N_SCE_M1044_g N_A_661_113#_c_2269_n 0.0162802f $X=4.6 $Y=2.595 $X2=0
+ $Y2=0
cc_823 N_SCE_c_1003_n N_A_661_113#_c_2243_n 4.69291e-19 $X=4.6 $Y=2.2 $X2=0
+ $Y2=0
cc_824 N_SCE_M1044_g N_A_661_113#_c_2243_n 0.00578626f $X=4.6 $Y=2.595 $X2=0
+ $Y2=0
cc_825 N_SCE_M1003_g N_A_661_113#_c_2233_n 0.00979553f $X=5.505 $Y=0.835 $X2=0
+ $Y2=0
cc_826 N_SCE_c_999_n N_A_661_113#_c_2239_n 0.00415211f $X=3.625 $Y=3.03 $X2=0
+ $Y2=0
cc_827 N_SCE_c_992_n N_A_661_113#_c_2239_n 5.38464e-19 $X=4.6 $Y=2.11 $X2=0
+ $Y2=0
cc_828 N_SCE_M1003_g N_A_661_113#_c_2240_n 0.00463009f $X=5.505 $Y=0.835 $X2=0
+ $Y2=0
cc_829 N_SCE_M1045_g N_VGND_c_2469_n 0.01623f $X=4.715 $Y=0.835 $X2=0 $Y2=0
cc_830 N_SCE_c_994_n N_VGND_c_2469_n 0.0182613f $X=5.43 $Y=0.18 $X2=0 $Y2=0
cc_831 N_SCE_c_995_n N_VGND_c_2469_n 0.00388727f $X=4.79 $Y=0.18 $X2=0 $Y2=0
cc_832 N_SCE_M1003_g N_VGND_c_2469_n 0.00691201f $X=5.505 $Y=0.835 $X2=0 $Y2=0
cc_833 SCE N_VGND_c_2469_n 0.00147588f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_834 N_SCE_c_994_n N_VGND_c_2470_n 0.01117f $X=5.43 $Y=0.18 $X2=0 $Y2=0
cc_835 N_SCE_M1003_g N_VGND_c_2470_n 5.60011e-19 $X=5.505 $Y=0.835 $X2=0 $Y2=0
cc_836 N_SCE_c_994_n N_VGND_c_2479_n 0.0177114f $X=5.43 $Y=0.18 $X2=0 $Y2=0
cc_837 N_SCE_c_995_n N_VGND_c_2485_n 0.00486043f $X=4.79 $Y=0.18 $X2=0 $Y2=0
cc_838 N_SCE_c_994_n N_VGND_c_2499_n 0.0266988f $X=5.43 $Y=0.18 $X2=0 $Y2=0
cc_839 N_SCE_c_995_n N_VGND_c_2499_n 0.00983503f $X=4.79 $Y=0.18 $X2=0 $Y2=0
cc_840 N_CLK_c_1081_n N_A_1313_74#_M1013_g 0.00452821f $X=6.65 $Y=1.73 $X2=0
+ $Y2=0
cc_841 CLK N_A_1313_74#_M1013_g 0.00132157f $X=6.875 $Y=1.21 $X2=0 $Y2=0
cc_842 N_CLK_c_1080_n N_A_1313_74#_c_1351_n 0.00636314f $X=6.49 $Y=1.22 $X2=0
+ $Y2=0
cc_843 N_CLK_c_1081_n N_A_1313_74#_c_1366_n 0.00814396f $X=6.65 $Y=1.73 $X2=0
+ $Y2=0
cc_844 CLK N_A_1313_74#_c_1366_n 0.0162653f $X=6.875 $Y=1.21 $X2=0 $Y2=0
cc_845 CLK N_A_1313_74#_c_1352_n 0.0159681f $X=6.875 $Y=1.21 $X2=0 $Y2=0
cc_846 N_CLK_c_1080_n N_A_1313_74#_c_1353_n 0.0033074f $X=6.49 $Y=1.22 $X2=0
+ $Y2=0
cc_847 N_CLK_c_1081_n N_A_1313_74#_c_1353_n 0.00109995f $X=6.65 $Y=1.73 $X2=0
+ $Y2=0
cc_848 CLK N_A_1313_74#_c_1353_n 0.0254473f $X=6.875 $Y=1.21 $X2=0 $Y2=0
cc_849 N_CLK_c_1080_n N_A_1313_74#_c_1354_n 0.0025538f $X=6.49 $Y=1.22 $X2=0
+ $Y2=0
cc_850 N_CLK_c_1081_n N_A_1313_74#_c_1354_n 0.00259477f $X=6.65 $Y=1.73 $X2=0
+ $Y2=0
cc_851 CLK N_A_1313_74#_c_1354_n 0.0308424f $X=6.875 $Y=1.21 $X2=0 $Y2=0
cc_852 N_CLK_c_1081_n N_A_1313_74#_c_1356_n 0.00979722f $X=6.65 $Y=1.73 $X2=0
+ $Y2=0
cc_853 N_CLK_c_1081_n N_VPWR_c_2041_n 0.0192789f $X=6.65 $Y=1.73 $X2=0 $Y2=0
cc_854 N_CLK_c_1081_n N_VPWR_c_2057_n 0.00495793f $X=6.65 $Y=1.73 $X2=0 $Y2=0
cc_855 N_CLK_c_1081_n N_VPWR_c_2037_n 0.00484764f $X=6.65 $Y=1.73 $X2=0 $Y2=0
cc_856 N_CLK_c_1080_n N_A_661_113#_c_2233_n 0.00384909f $X=6.49 $Y=1.22 $X2=0
+ $Y2=0
cc_857 N_CLK_c_1081_n N_A_661_113#_c_2234_n 0.0151779f $X=6.65 $Y=1.73 $X2=0
+ $Y2=0
cc_858 CLK N_A_661_113#_c_2234_n 0.0177648f $X=6.875 $Y=1.21 $X2=0 $Y2=0
cc_859 N_CLK_c_1081_n N_A_661_113#_c_2245_n 0.0172018f $X=6.65 $Y=1.73 $X2=0
+ $Y2=0
cc_860 N_CLK_c_1080_n N_A_661_113#_c_2240_n 0.00537533f $X=6.49 $Y=1.22 $X2=0
+ $Y2=0
cc_861 CLK N_A_661_113#_c_2240_n 0.00406505f $X=6.875 $Y=1.21 $X2=0 $Y2=0
cc_862 N_CLK_c_1081_n N_A_661_113#_c_2249_n 0.00364957f $X=6.65 $Y=1.73 $X2=0
+ $Y2=0
cc_863 N_CLK_c_1081_n N_A_661_113#_c_2251_n 0.00261254f $X=6.65 $Y=1.73 $X2=0
+ $Y2=0
cc_864 N_CLK_c_1080_n N_VGND_c_2470_n 0.0076584f $X=6.49 $Y=1.22 $X2=0 $Y2=0
cc_865 N_CLK_c_1080_n N_VGND_c_2471_n 0.00334136f $X=6.49 $Y=1.22 $X2=0 $Y2=0
cc_866 N_CLK_c_1080_n N_VGND_c_2481_n 0.00434272f $X=6.49 $Y=1.22 $X2=0 $Y2=0
cc_867 N_CLK_c_1080_n N_VGND_c_2499_n 0.00830282f $X=6.49 $Y=1.22 $X2=0 $Y2=0
cc_868 N_A_1510_74#_c_1118_n N_A_1313_74#_M1013_g 0.00159626f $X=7.69 $Y=0.515
+ $X2=0 $Y2=0
cc_869 N_A_1510_74#_c_1120_n N_A_1313_74#_M1013_g 0.00266901f $X=7.855 $Y=0.34
+ $X2=0 $Y2=0
cc_870 N_A_1510_74#_c_1118_n N_A_1313_74#_c_1343_n 0.00277021f $X=7.69 $Y=0.515
+ $X2=0 $Y2=0
cc_871 N_A_1510_74#_c_1143_n N_A_1313_74#_c_1358_n 0.00413487f $X=8.495 $Y=1.992
+ $X2=0 $Y2=0
cc_872 N_A_1510_74#_c_1121_n N_A_1313_74#_c_1358_n 9.29699e-19 $X=8.58 $Y=1.82
+ $X2=0 $Y2=0
cc_873 N_A_1510_74#_c_1147_n N_A_1313_74#_c_1358_n 0.00131308f $X=8.58 $Y=2.077
+ $X2=0 $Y2=0
cc_874 N_A_1510_74#_c_1148_n N_A_1313_74#_c_1358_n 0.00570117f $X=8.675 $Y=2.17
+ $X2=0 $Y2=0
cc_875 N_A_1510_74#_c_1143_n N_A_1313_74#_c_1344_n 0.0107509f $X=8.495 $Y=1.992
+ $X2=0 $Y2=0
cc_876 N_A_1510_74#_c_1121_n N_A_1313_74#_c_1344_n 0.00722536f $X=8.58 $Y=1.82
+ $X2=0 $Y2=0
cc_877 N_A_1510_74#_c_1148_n N_A_1313_74#_c_1344_n 0.0180858f $X=8.675 $Y=2.17
+ $X2=0 $Y2=0
cc_878 N_A_1510_74#_c_1115_n N_A_1313_74#_M1040_g 0.0197489f $X=9.215 $Y=0.925
+ $X2=0 $Y2=0
cc_879 N_A_1510_74#_c_1121_n N_A_1313_74#_M1040_g 0.0345945f $X=8.58 $Y=1.82
+ $X2=0 $Y2=0
cc_880 N_A_1510_74#_c_1122_n N_A_1313_74#_M1040_g 0.00861265f $X=9.175 $Y=0.34
+ $X2=0 $Y2=0
cc_881 N_A_1510_74#_c_1123_n N_A_1313_74#_M1040_g 7.08973e-19 $X=9.34 $Y=0.86
+ $X2=0 $Y2=0
cc_882 N_A_1510_74#_c_1134_n N_A_1313_74#_M1040_g 0.00248552f $X=8.58 $Y=0.34
+ $X2=0 $Y2=0
cc_883 N_A_1510_74#_c_1148_n N_A_1313_74#_c_1346_n 0.00575555f $X=8.675 $Y=2.17
+ $X2=0 $Y2=0
cc_884 N_A_1510_74#_c_1135_n N_A_1313_74#_c_1346_n 7.59768e-19 $X=9.34 $Y=0.945
+ $X2=0 $Y2=0
cc_885 N_A_1510_74#_c_1136_n N_A_1313_74#_c_1346_n 0.0101403f $X=9.34 $Y=1.09
+ $X2=0 $Y2=0
cc_886 N_A_1510_74#_c_1140_n N_A_1313_74#_c_1362_n 0.0101282f $X=8.97 $Y=2.465
+ $X2=0 $Y2=0
cc_887 N_A_1510_74#_c_1148_n N_A_1313_74#_c_1362_n 0.0186322f $X=8.675 $Y=2.17
+ $X2=0 $Y2=0
cc_888 N_A_1510_74#_c_1117_n N_A_1313_74#_c_1347_n 0.0202897f $X=12.855 $Y=2.375
+ $X2=0 $Y2=0
cc_889 N_A_1510_74#_c_1142_n N_A_1313_74#_c_1347_n 0.0126385f $X=12.855 $Y=2.465
+ $X2=0 $Y2=0
cc_890 N_A_1510_74#_c_1131_n N_A_1313_74#_c_1347_n 6.96576e-19 $X=11.85 $Y=1.635
+ $X2=0 $Y2=0
cc_891 N_A_1510_74#_c_1132_n N_A_1313_74#_c_1347_n 0.0216845f $X=11.85 $Y=1.635
+ $X2=0 $Y2=0
cc_892 N_A_1510_74#_c_1133_n N_A_1313_74#_c_1347_n 0.00464354f $X=12.765
+ $Y=1.275 $X2=0 $Y2=0
cc_893 N_A_1510_74#_c_1138_n N_A_1313_74#_c_1347_n 5.03473e-19 $X=12.93 $Y=1.275
+ $X2=0 $Y2=0
cc_894 N_A_1510_74#_c_1139_n N_A_1313_74#_c_1347_n 0.02153f $X=12.93 $Y=1.42
+ $X2=0 $Y2=0
cc_895 N_A_1510_74#_M1031_g N_A_1313_74#_M1016_g 0.0312272f $X=11.94 $Y=0.69
+ $X2=0 $Y2=0
cc_896 N_A_1510_74#_c_1131_n N_A_1313_74#_M1016_g 5.85904e-19 $X=11.85 $Y=1.635
+ $X2=0 $Y2=0
cc_897 N_A_1510_74#_c_1133_n N_A_1313_74#_M1016_g 0.0110881f $X=12.765 $Y=1.275
+ $X2=0 $Y2=0
cc_898 N_A_1510_74#_c_1138_n N_A_1313_74#_M1016_g 0.001f $X=12.93 $Y=1.275 $X2=0
+ $Y2=0
cc_899 N_A_1510_74#_c_1139_n N_A_1313_74#_M1016_g 0.0101758f $X=12.93 $Y=1.42
+ $X2=0 $Y2=0
cc_900 N_A_1510_74#_c_1121_n N_A_1313_74#_c_1350_n 0.00213866f $X=8.58 $Y=1.82
+ $X2=0 $Y2=0
cc_901 N_A_1510_74#_c_1147_n N_A_1313_74#_c_1350_n 0.00370702f $X=8.58 $Y=2.077
+ $X2=0 $Y2=0
cc_902 N_A_1510_74#_c_1118_n N_A_1313_74#_c_1354_n 0.00438992f $X=7.69 $Y=0.515
+ $X2=0 $Y2=0
cc_903 N_A_1510_74#_c_1131_n N_A_1313_74#_c_1368_n 0.00785016f $X=11.85 $Y=1.635
+ $X2=0 $Y2=0
cc_904 N_A_1510_74#_c_1132_n N_A_1313_74#_c_1368_n 0.00300142f $X=11.85 $Y=1.635
+ $X2=0 $Y2=0
cc_905 N_A_1510_74#_c_1117_n N_A_1313_74#_c_1369_n 4.93293e-19 $X=12.855
+ $Y=2.375 $X2=0 $Y2=0
cc_906 N_A_1510_74#_c_1131_n N_A_1313_74#_c_1369_n 0.00333066f $X=11.85 $Y=1.635
+ $X2=0 $Y2=0
cc_907 N_A_1510_74#_c_1132_n N_A_1313_74#_c_1369_n 2.67802e-19 $X=11.85 $Y=1.635
+ $X2=0 $Y2=0
cc_908 N_A_1510_74#_c_1131_n N_A_1313_74#_c_1355_n 0.016352f $X=11.85 $Y=1.635
+ $X2=0 $Y2=0
cc_909 N_A_1510_74#_c_1132_n N_A_1313_74#_c_1355_n 0.00123323f $X=11.85 $Y=1.635
+ $X2=0 $Y2=0
cc_910 N_A_1510_74#_c_1133_n N_A_1313_74#_c_1355_n 0.0286707f $X=12.765 $Y=1.275
+ $X2=0 $Y2=0
cc_911 N_A_1510_74#_c_1138_n N_A_1313_74#_c_1355_n 0.00350748f $X=12.93 $Y=1.275
+ $X2=0 $Y2=0
cc_912 N_A_1510_74#_c_1139_n N_A_1313_74#_c_1355_n 0.00194604f $X=12.93 $Y=1.42
+ $X2=0 $Y2=0
cc_913 N_A_1510_74#_c_1125_n N_A_1943_53#_M1046_d 0.00427127f $X=10.94 $Y=0.34
+ $X2=-0.19 $Y2=-0.245
cc_914 N_A_1510_74#_c_1115_n N_A_1943_53#_M1032_g 0.0150403f $X=9.215 $Y=0.925
+ $X2=0 $Y2=0
cc_915 N_A_1510_74#_c_1122_n N_A_1943_53#_M1032_g 0.00154688f $X=9.175 $Y=0.34
+ $X2=0 $Y2=0
cc_916 N_A_1510_74#_c_1123_n N_A_1943_53#_M1032_g 0.00637996f $X=9.34 $Y=0.86
+ $X2=0 $Y2=0
cc_917 N_A_1510_74#_c_1124_n N_A_1943_53#_M1032_g 0.0124305f $X=10.26 $Y=0.945
+ $X2=0 $Y2=0
cc_918 N_A_1510_74#_c_1221_p N_A_1943_53#_M1032_g 0.00284853f $X=10.345 $Y=0.86
+ $X2=0 $Y2=0
cc_919 N_A_1510_74#_c_1126_n N_A_1943_53#_M1032_g 4.25169e-19 $X=10.43 $Y=0.34
+ $X2=0 $Y2=0
cc_920 N_A_1510_74#_c_1135_n N_A_1943_53#_M1032_g 0.00131332f $X=9.34 $Y=0.945
+ $X2=0 $Y2=0
cc_921 N_A_1510_74#_c_1136_n N_A_1943_53#_M1032_g 0.0214344f $X=9.34 $Y=1.09
+ $X2=0 $Y2=0
cc_922 N_A_1510_74#_M1031_g N_A_1943_53#_c_1536_n 0.0596831f $X=11.94 $Y=0.69
+ $X2=0 $Y2=0
cc_923 N_A_1510_74#_c_1125_n N_A_1943_53#_c_1536_n 6.63977e-19 $X=10.94 $Y=0.34
+ $X2=0 $Y2=0
cc_924 N_A_1510_74#_c_1127_n N_A_1943_53#_c_1536_n 0.00423957f $X=11.025 $Y=0.86
+ $X2=0 $Y2=0
cc_925 N_A_1510_74#_c_1128_n N_A_1943_53#_c_1536_n 0.0138048f $X=11.685 $Y=0.945
+ $X2=0 $Y2=0
cc_926 N_A_1510_74#_c_1130_n N_A_1943_53#_c_1536_n 0.00382611f $X=11.77 $Y=1.19
+ $X2=0 $Y2=0
cc_927 N_A_1510_74#_c_1124_n N_A_1943_53#_c_1537_n 0.0109975f $X=10.26 $Y=0.945
+ $X2=0 $Y2=0
cc_928 N_A_1510_74#_c_1125_n N_A_1943_53#_c_1538_n 0.0127109f $X=10.94 $Y=0.34
+ $X2=0 $Y2=0
cc_929 N_A_1510_74#_c_1127_n N_A_1943_53#_c_1538_n 0.0195631f $X=11.025 $Y=0.86
+ $X2=0 $Y2=0
cc_930 N_A_1510_74#_c_1129_n N_A_1943_53#_c_1538_n 0.0141315f $X=11.11 $Y=0.945
+ $X2=0 $Y2=0
cc_931 N_A_1510_74#_M1031_g N_A_1943_53#_c_1541_n 2.51383e-19 $X=11.94 $Y=0.69
+ $X2=0 $Y2=0
cc_932 N_A_1510_74#_c_1128_n N_A_1943_53#_c_1541_n 0.0267734f $X=11.685 $Y=0.945
+ $X2=0 $Y2=0
cc_933 N_A_1510_74#_c_1129_n N_A_1943_53#_c_1541_n 0.0146025f $X=11.11 $Y=0.945
+ $X2=0 $Y2=0
cc_934 N_A_1510_74#_c_1131_n N_A_1943_53#_c_1541_n 0.0116825f $X=11.85 $Y=1.635
+ $X2=0 $Y2=0
cc_935 N_A_1510_74#_c_1132_n N_A_1943_53#_c_1541_n 2.05067e-19 $X=11.85 $Y=1.635
+ $X2=0 $Y2=0
cc_936 N_A_1510_74#_c_1137_n N_A_1943_53#_c_1541_n 0.0120804f $X=11.82 $Y=1.275
+ $X2=0 $Y2=0
cc_937 N_A_1510_74#_c_1124_n N_A_1943_53#_c_1542_n 0.00480056f $X=10.26 $Y=0.945
+ $X2=0 $Y2=0
cc_938 N_A_1510_74#_c_1124_n N_A_1943_53#_c_1543_n 0.038229f $X=10.26 $Y=0.945
+ $X2=0 $Y2=0
cc_939 N_A_1510_74#_c_1135_n N_A_1943_53#_c_1543_n 0.00363676f $X=9.34 $Y=0.945
+ $X2=0 $Y2=0
cc_940 N_A_1510_74#_M1031_g N_A_1943_53#_c_1544_n 0.00604034f $X=11.94 $Y=0.69
+ $X2=0 $Y2=0
cc_941 N_A_1510_74#_c_1128_n N_A_1943_53#_c_1544_n 0.010336f $X=11.685 $Y=0.945
+ $X2=0 $Y2=0
cc_942 N_A_1510_74#_c_1131_n N_A_1943_53#_c_1544_n 0.00288564f $X=11.85 $Y=1.635
+ $X2=0 $Y2=0
cc_943 N_A_1510_74#_c_1132_n N_A_1943_53#_c_1544_n 0.0220039f $X=11.85 $Y=1.635
+ $X2=0 $Y2=0
cc_944 N_A_1510_74#_c_1137_n N_A_1943_53#_c_1544_n 0.00136894f $X=11.82 $Y=1.275
+ $X2=0 $Y2=0
cc_945 N_A_1510_74#_c_1122_n N_A_1756_97#_M1040_d 0.00422613f $X=9.175 $Y=0.34
+ $X2=-0.19 $Y2=-0.245
cc_946 N_A_1510_74#_c_1124_n N_A_1756_97#_M1046_g 0.00554f $X=10.26 $Y=0.945
+ $X2=0 $Y2=0
cc_947 N_A_1510_74#_c_1221_p N_A_1756_97#_M1046_g 0.0113905f $X=10.345 $Y=0.86
+ $X2=0 $Y2=0
cc_948 N_A_1510_74#_c_1125_n N_A_1756_97#_M1046_g 0.0120035f $X=10.94 $Y=0.34
+ $X2=0 $Y2=0
cc_949 N_A_1510_74#_c_1126_n N_A_1756_97#_M1046_g 0.00287637f $X=10.43 $Y=0.34
+ $X2=0 $Y2=0
cc_950 N_A_1510_74#_c_1127_n N_A_1756_97#_M1046_g 0.00329118f $X=11.025 $Y=0.86
+ $X2=0 $Y2=0
cc_951 N_A_1510_74#_c_1115_n N_A_1756_97#_c_1641_n 0.00482329f $X=9.215 $Y=0.925
+ $X2=0 $Y2=0
cc_952 N_A_1510_74#_c_1121_n N_A_1756_97#_c_1641_n 0.0621438f $X=8.58 $Y=1.82
+ $X2=0 $Y2=0
cc_953 N_A_1510_74#_c_1122_n N_A_1756_97#_c_1641_n 0.0128192f $X=9.175 $Y=0.34
+ $X2=0 $Y2=0
cc_954 N_A_1510_74#_c_1123_n N_A_1756_97#_c_1641_n 0.049118f $X=9.34 $Y=0.86
+ $X2=0 $Y2=0
cc_955 N_A_1510_74#_c_1121_n N_A_1756_97#_c_1645_n 0.0119898f $X=8.58 $Y=1.82
+ $X2=0 $Y2=0
cc_956 N_A_1510_74#_c_1148_n N_A_1756_97#_c_1645_n 0.00303355f $X=8.675 $Y=2.17
+ $X2=0 $Y2=0
cc_957 N_A_1510_74#_c_1136_n N_A_1756_97#_c_1645_n 3.64767e-19 $X=9.34 $Y=1.09
+ $X2=0 $Y2=0
cc_958 N_A_1510_74#_c_1140_n N_A_1756_97#_c_1646_n 0.00681887f $X=8.97 $Y=2.465
+ $X2=0 $Y2=0
cc_959 N_A_1510_74#_c_1140_n N_A_1756_97#_c_1647_n 0.00148452f $X=8.97 $Y=2.465
+ $X2=0 $Y2=0
cc_960 N_A_1510_74#_c_1121_n N_A_1756_97#_c_1647_n 9.18312e-19 $X=8.58 $Y=1.82
+ $X2=0 $Y2=0
cc_961 N_A_1510_74#_c_1147_n N_A_1756_97#_c_1647_n 0.03506f $X=8.58 $Y=2.077
+ $X2=0 $Y2=0
cc_962 N_A_1510_74#_c_1148_n N_A_1756_97#_c_1647_n 0.0103718f $X=8.675 $Y=2.17
+ $X2=0 $Y2=0
cc_963 N_A_1510_74#_c_1124_n N_A_1756_97#_c_1643_n 0.00365265f $X=10.26 $Y=0.945
+ $X2=0 $Y2=0
cc_964 N_A_1510_74#_c_1135_n N_A_1756_97#_c_1643_n 0.00889803f $X=9.34 $Y=0.945
+ $X2=0 $Y2=0
cc_965 N_A_1510_74#_c_1136_n N_A_1756_97#_c_1643_n 8.95132e-19 $X=9.34 $Y=1.09
+ $X2=0 $Y2=0
cc_966 N_A_1510_74#_M1031_g N_A_2403_74#_c_1735_n 7.35604e-19 $X=11.94 $Y=0.69
+ $X2=0 $Y2=0
cc_967 N_A_1510_74#_c_1133_n N_A_2403_74#_c_1736_n 0.028365f $X=12.765 $Y=1.275
+ $X2=0 $Y2=0
cc_968 N_A_1510_74#_c_1138_n N_A_2403_74#_c_1736_n 0.02584f $X=12.93 $Y=1.275
+ $X2=0 $Y2=0
cc_969 N_A_1510_74#_c_1139_n N_A_2403_74#_c_1736_n 8.40831e-19 $X=12.93 $Y=1.42
+ $X2=0 $Y2=0
cc_970 N_A_1510_74#_M1031_g N_A_2403_74#_c_1737_n 9.17078e-19 $X=11.94 $Y=0.69
+ $X2=0 $Y2=0
cc_971 N_A_1510_74#_c_1128_n N_A_2403_74#_c_1737_n 8.0891e-19 $X=11.685 $Y=0.945
+ $X2=0 $Y2=0
cc_972 N_A_1510_74#_c_1133_n N_A_2403_74#_c_1737_n 0.0268237f $X=12.765 $Y=1.275
+ $X2=0 $Y2=0
cc_973 N_A_1510_74#_c_1117_n N_A_2403_74#_c_1749_n 0.00754943f $X=12.855
+ $Y=2.375 $X2=0 $Y2=0
cc_974 N_A_1510_74#_c_1142_n N_A_2403_74#_c_1749_n 0.018329f $X=12.855 $Y=2.465
+ $X2=0 $Y2=0
cc_975 N_A_1510_74#_c_1117_n N_A_2403_74#_c_1750_n 0.00607654f $X=12.855
+ $Y=2.375 $X2=0 $Y2=0
cc_976 N_A_1510_74#_c_1138_n N_A_2403_74#_c_1750_n 0.0116579f $X=12.93 $Y=1.275
+ $X2=0 $Y2=0
cc_977 N_A_1510_74#_c_1139_n N_A_2403_74#_c_1750_n 0.00105037f $X=12.93 $Y=1.42
+ $X2=0 $Y2=0
cc_978 N_A_1510_74#_c_1117_n N_A_2403_74#_c_1751_n 0.0128966f $X=12.855 $Y=2.375
+ $X2=0 $Y2=0
cc_979 N_A_1510_74#_c_1133_n N_A_2403_74#_c_1751_n 0.00352142f $X=12.765
+ $Y=1.275 $X2=0 $Y2=0
cc_980 N_A_1510_74#_c_1138_n N_A_2403_74#_c_1751_n 0.00816138f $X=12.93 $Y=1.275
+ $X2=0 $Y2=0
cc_981 N_A_1510_74#_c_1117_n N_A_2403_74#_c_1738_n 0.00280042f $X=12.855
+ $Y=2.375 $X2=0 $Y2=0
cc_982 N_A_1510_74#_c_1138_n N_A_2403_74#_c_1738_n 0.0334325f $X=12.93 $Y=1.275
+ $X2=0 $Y2=0
cc_983 N_A_1510_74#_c_1139_n N_A_2403_74#_c_1738_n 0.00215716f $X=12.93 $Y=1.42
+ $X2=0 $Y2=0
cc_984 N_A_1510_74#_c_1142_n N_VPWR_c_2045_n 0.00144848f $X=12.855 $Y=2.465
+ $X2=0 $Y2=0
cc_985 N_A_1510_74#_c_1140_n N_VPWR_c_2051_n 0.00411612f $X=8.97 $Y=2.465 $X2=0
+ $Y2=0
cc_986 N_A_1510_74#_c_1142_n N_VPWR_c_2059_n 0.00332301f $X=12.855 $Y=2.465
+ $X2=0 $Y2=0
cc_987 N_A_1510_74#_c_1140_n N_VPWR_c_2037_n 0.00753176f $X=8.97 $Y=2.465 $X2=0
+ $Y2=0
cc_988 N_A_1510_74#_c_1142_n N_VPWR_c_2037_n 0.00529713f $X=12.855 $Y=2.465
+ $X2=0 $Y2=0
cc_989 N_A_1510_74#_c_1148_n N_VPWR_c_2037_n 3.2759e-19 $X=8.675 $Y=2.17 $X2=0
+ $Y2=0
cc_990 N_A_1510_74#_c_1121_n N_A_661_113#_M1040_s 0.00544605f $X=8.58 $Y=1.82
+ $X2=0 $Y2=0
cc_991 N_A_1510_74#_c_1143_n N_A_661_113#_c_2246_n 0.0149994f $X=8.495 $Y=1.992
+ $X2=0 $Y2=0
cc_992 N_A_1510_74#_c_1121_n N_A_661_113#_c_2246_n 0.00327926f $X=8.58 $Y=1.82
+ $X2=0 $Y2=0
cc_993 N_A_1510_74#_c_1143_n N_A_661_113#_c_2235_n 0.0174322f $X=8.495 $Y=1.992
+ $X2=0 $Y2=0
cc_994 N_A_1510_74#_c_1121_n N_A_661_113#_c_2235_n 0.0133653f $X=8.58 $Y=1.82
+ $X2=0 $Y2=0
cc_995 N_A_1510_74#_c_1118_n N_A_661_113#_c_2236_n 0.00648607f $X=7.69 $Y=0.515
+ $X2=0 $Y2=0
cc_996 N_A_1510_74#_M1029_d N_A_661_113#_c_2247_n 0.0153668f $X=8.075 $Y=1.84
+ $X2=0 $Y2=0
cc_997 N_A_1510_74#_c_1140_n N_A_661_113#_c_2247_n 0.00401873f $X=8.97 $Y=2.465
+ $X2=0 $Y2=0
cc_998 N_A_1510_74#_c_1143_n N_A_661_113#_c_2247_n 0.02575f $X=8.495 $Y=1.992
+ $X2=0 $Y2=0
cc_999 N_A_1510_74#_c_1147_n N_A_661_113#_c_2247_n 0.0284119f $X=8.58 $Y=2.077
+ $X2=0 $Y2=0
cc_1000 N_A_1510_74#_c_1148_n N_A_661_113#_c_2247_n 0.00465406f $X=8.675 $Y=2.17
+ $X2=0 $Y2=0
cc_1001 N_A_1510_74#_c_1118_n N_A_661_113#_c_2237_n 0.0356656f $X=7.69 $Y=0.515
+ $X2=0 $Y2=0
cc_1002 N_A_1510_74#_c_1119_n N_A_661_113#_c_2237_n 0.0192437f $X=8.495 $Y=0.34
+ $X2=0 $Y2=0
cc_1003 N_A_1510_74#_c_1121_n N_A_661_113#_c_2237_n 0.0677461f $X=8.58 $Y=1.82
+ $X2=0 $Y2=0
cc_1004 N_A_1510_74#_c_1124_n N_VGND_M1032_d 0.00485076f $X=10.26 $Y=0.945 $X2=0
+ $Y2=0
cc_1005 N_A_1510_74#_c_1221_p N_VGND_M1032_d 0.0047792f $X=10.345 $Y=0.86 $X2=0
+ $Y2=0
cc_1006 N_A_1510_74#_c_1126_n N_VGND_M1032_d 2.8512e-19 $X=10.43 $Y=0.34 $X2=0
+ $Y2=0
cc_1007 N_A_1510_74#_c_1128_n N_VGND_M1047_s 0.00386678f $X=11.685 $Y=0.945
+ $X2=0 $Y2=0
cc_1008 N_A_1510_74#_c_1120_n N_VGND_c_2471_n 0.0112234f $X=7.855 $Y=0.34 $X2=0
+ $Y2=0
cc_1009 N_A_1510_74#_c_1115_n N_VGND_c_2472_n 3.55414e-19 $X=9.215 $Y=0.925
+ $X2=0 $Y2=0
cc_1010 N_A_1510_74#_c_1122_n N_VGND_c_2472_n 0.00848359f $X=9.175 $Y=0.34 $X2=0
+ $Y2=0
cc_1011 N_A_1510_74#_c_1123_n N_VGND_c_2472_n 0.0119616f $X=9.34 $Y=0.86 $X2=0
+ $Y2=0
cc_1012 N_A_1510_74#_c_1124_n N_VGND_c_2472_n 0.01733f $X=10.26 $Y=0.945 $X2=0
+ $Y2=0
cc_1013 N_A_1510_74#_c_1221_p N_VGND_c_2472_n 0.0197837f $X=10.345 $Y=0.86 $X2=0
+ $Y2=0
cc_1014 N_A_1510_74#_c_1126_n N_VGND_c_2472_n 0.0146484f $X=10.43 $Y=0.34 $X2=0
+ $Y2=0
cc_1015 N_A_1510_74#_M1031_g N_VGND_c_2473_n 0.00152129f $X=11.94 $Y=0.69 $X2=0
+ $Y2=0
cc_1016 N_A_1510_74#_c_1125_n N_VGND_c_2473_n 0.0146661f $X=10.94 $Y=0.34 $X2=0
+ $Y2=0
cc_1017 N_A_1510_74#_c_1127_n N_VGND_c_2473_n 0.0201354f $X=11.025 $Y=0.86 $X2=0
+ $Y2=0
cc_1018 N_A_1510_74#_c_1128_n N_VGND_c_2473_n 0.0150603f $X=11.685 $Y=0.945
+ $X2=0 $Y2=0
cc_1019 N_A_1510_74#_c_1115_n N_VGND_c_2486_n 9.62735e-19 $X=9.215 $Y=0.925
+ $X2=0 $Y2=0
cc_1020 N_A_1510_74#_c_1119_n N_VGND_c_2486_n 0.0411694f $X=8.495 $Y=0.34 $X2=0
+ $Y2=0
cc_1021 N_A_1510_74#_c_1120_n N_VGND_c_2486_n 0.0179217f $X=7.855 $Y=0.34 $X2=0
+ $Y2=0
cc_1022 N_A_1510_74#_c_1122_n N_VGND_c_2486_n 0.0564517f $X=9.175 $Y=0.34 $X2=0
+ $Y2=0
cc_1023 N_A_1510_74#_c_1134_n N_VGND_c_2486_n 0.0121867f $X=8.58 $Y=0.34 $X2=0
+ $Y2=0
cc_1024 N_A_1510_74#_c_1125_n N_VGND_c_2487_n 0.0449818f $X=10.94 $Y=0.34 $X2=0
+ $Y2=0
cc_1025 N_A_1510_74#_c_1126_n N_VGND_c_2487_n 0.0121867f $X=10.43 $Y=0.34 $X2=0
+ $Y2=0
cc_1026 N_A_1510_74#_M1031_g N_VGND_c_2495_n 0.00461464f $X=11.94 $Y=0.69 $X2=0
+ $Y2=0
cc_1027 N_A_1510_74#_M1031_g N_VGND_c_2499_n 0.0090922f $X=11.94 $Y=0.69 $X2=0
+ $Y2=0
cc_1028 N_A_1510_74#_c_1119_n N_VGND_c_2499_n 0.0240545f $X=8.495 $Y=0.34 $X2=0
+ $Y2=0
cc_1029 N_A_1510_74#_c_1120_n N_VGND_c_2499_n 0.00971942f $X=7.855 $Y=0.34 $X2=0
+ $Y2=0
cc_1030 N_A_1510_74#_c_1122_n N_VGND_c_2499_n 0.0319965f $X=9.175 $Y=0.34 $X2=0
+ $Y2=0
cc_1031 N_A_1510_74#_c_1124_n N_VGND_c_2499_n 0.017544f $X=10.26 $Y=0.945 $X2=0
+ $Y2=0
cc_1032 N_A_1510_74#_c_1125_n N_VGND_c_2499_n 0.025776f $X=10.94 $Y=0.34 $X2=0
+ $Y2=0
cc_1033 N_A_1510_74#_c_1126_n N_VGND_c_2499_n 0.00660921f $X=10.43 $Y=0.34 $X2=0
+ $Y2=0
cc_1034 N_A_1510_74#_c_1128_n N_VGND_c_2499_n 0.0175282f $X=11.685 $Y=0.945
+ $X2=0 $Y2=0
cc_1035 N_A_1510_74#_c_1134_n N_VGND_c_2499_n 0.00660921f $X=8.58 $Y=0.34 $X2=0
+ $Y2=0
cc_1036 N_A_1510_74#_c_1122_n A_1858_79# 4.09921e-19 $X=9.175 $Y=0.34 $X2=-0.19
+ $Y2=-0.245
cc_1037 N_A_1510_74#_c_1123_n A_1858_79# 0.00524566f $X=9.34 $Y=0.86 $X2=-0.19
+ $Y2=-0.245
cc_1038 N_A_1510_74#_c_1128_n A_2331_74# 0.00231857f $X=11.685 $Y=0.945
+ $X2=-0.19 $Y2=-0.245
cc_1039 N_A_1313_74#_c_1368_n N_A_1943_53#_M1043_d 0.00728602f $X=12.125
+ $Y=2.475 $X2=0 $Y2=0
cc_1040 N_A_1313_74#_c_1346_n N_A_1943_53#_c_1534_n 0.0121937f $X=9.27 $Y=1.69
+ $X2=0 $Y2=0
cc_1041 N_A_1313_74#_c_1362_n N_A_1943_53#_c_1534_n 0.0243178f $X=9.42 $Y=2.465
+ $X2=0 $Y2=0
cc_1042 N_A_1313_74#_c_1370_n N_A_1943_53#_c_1534_n 0.00963636f $X=9.435
+ $Y=2.165 $X2=0 $Y2=0
cc_1043 N_A_1313_74#_c_1362_n N_A_1943_53#_c_1546_n 0.0221968f $X=9.42 $Y=2.465
+ $X2=0 $Y2=0
cc_1044 N_A_1313_74#_c_1368_n N_A_1943_53#_c_1546_n 0.0152453f $X=12.125
+ $Y=2.475 $X2=0 $Y2=0
cc_1045 N_A_1313_74#_c_1368_n N_A_1943_53#_c_1548_n 0.0202137f $X=12.125
+ $Y=2.475 $X2=0 $Y2=0
cc_1046 N_A_1313_74#_c_1369_n N_A_1943_53#_c_1548_n 0.0121681f $X=12.21 $Y=2.39
+ $X2=0 $Y2=0
cc_1047 N_A_1313_74#_c_1368_n N_A_1943_53#_c_1549_n 0.0308108f $X=12.125
+ $Y=2.475 $X2=0 $Y2=0
cc_1048 N_A_1313_74#_c_1368_n N_A_1756_97#_c_1639_n 0.0168265f $X=12.125
+ $Y=2.475 $X2=0 $Y2=0
cc_1049 N_A_1313_74#_M1040_g N_A_1756_97#_c_1641_n 0.0106185f $X=8.705 $Y=0.695
+ $X2=0 $Y2=0
cc_1050 N_A_1313_74#_c_1346_n N_A_1756_97#_c_1641_n 0.00473461f $X=9.27 $Y=1.69
+ $X2=0 $Y2=0
cc_1051 N_A_1313_74#_c_1346_n N_A_1756_97#_c_1645_n 0.0113733f $X=9.27 $Y=1.69
+ $X2=0 $Y2=0
cc_1052 N_A_1313_74#_c_1362_n N_A_1756_97#_c_1646_n 0.0126416f $X=9.42 $Y=2.465
+ $X2=0 $Y2=0
cc_1053 N_A_1313_74#_c_1370_n N_A_1756_97#_c_1646_n 0.00378639f $X=9.435
+ $Y=2.165 $X2=0 $Y2=0
cc_1054 N_A_1313_74#_c_1346_n N_A_1756_97#_c_1647_n 0.00143134f $X=9.27 $Y=1.69
+ $X2=0 $Y2=0
cc_1055 N_A_1313_74#_c_1361_n N_A_1756_97#_c_1647_n 0.0100195f $X=9.345 $Y=2
+ $X2=0 $Y2=0
cc_1056 N_A_1313_74#_c_1362_n N_A_1756_97#_c_1647_n 0.00147297f $X=9.42 $Y=2.465
+ $X2=0 $Y2=0
cc_1057 N_A_1313_74#_c_1370_n N_A_1756_97#_c_1647_n 0.0342485f $X=9.435 $Y=2.165
+ $X2=0 $Y2=0
cc_1058 N_A_1313_74#_c_1346_n N_A_1756_97#_c_1643_n 0.0066017f $X=9.27 $Y=1.69
+ $X2=0 $Y2=0
cc_1059 N_A_1313_74#_c_1361_n N_A_1756_97#_c_1643_n 0.00582153f $X=9.345 $Y=2
+ $X2=0 $Y2=0
cc_1060 N_A_1313_74#_c_1362_n N_A_1756_97#_c_1643_n 0.0012185f $X=9.42 $Y=2.465
+ $X2=0 $Y2=0
cc_1061 N_A_1313_74#_c_1368_n N_A_1756_97#_c_1643_n 0.0208427f $X=12.125
+ $Y=2.475 $X2=0 $Y2=0
cc_1062 N_A_1313_74#_c_1370_n N_A_1756_97#_c_1643_n 0.0221092f $X=9.435 $Y=2.165
+ $X2=0 $Y2=0
cc_1063 N_A_1313_74#_M1016_g N_A_2403_74#_c_1735_n 0.00995617f $X=12.415 $Y=0.58
+ $X2=0 $Y2=0
cc_1064 N_A_1313_74#_M1016_g N_A_2403_74#_c_1736_n 0.00821531f $X=12.415 $Y=0.58
+ $X2=0 $Y2=0
cc_1065 N_A_1313_74#_M1016_g N_A_2403_74#_c_1737_n 0.00270117f $X=12.415 $Y=0.58
+ $X2=0 $Y2=0
cc_1066 N_A_1313_74#_c_1347_n N_A_2403_74#_c_1749_n 0.0048907f $X=12.345
+ $Y=1.885 $X2=0 $Y2=0
cc_1067 N_A_1313_74#_c_1347_n N_A_2403_74#_c_1751_n 0.00508401f $X=12.345
+ $Y=1.885 $X2=0 $Y2=0
cc_1068 N_A_1313_74#_c_1369_n N_A_2403_74#_c_1751_n 0.0156644f $X=12.21 $Y=2.39
+ $X2=0 $Y2=0
cc_1069 N_A_1313_74#_c_1355_n N_A_2403_74#_c_1751_n 0.00663964f $X=12.39
+ $Y=1.635 $X2=0 $Y2=0
cc_1070 N_A_1313_74#_c_1368_n N_VPWR_M1007_d 0.00663907f $X=12.125 $Y=2.475
+ $X2=0 $Y2=0
cc_1071 N_A_1313_74#_c_1368_n N_VPWR_M1027_s 0.011473f $X=12.125 $Y=2.475 $X2=0
+ $Y2=0
cc_1072 N_A_1313_74#_c_1358_n N_VPWR_c_2042_n 0.0110684f $X=8 $Y=1.765 $X2=0
+ $Y2=0
cc_1073 N_A_1313_74#_c_1362_n N_VPWR_c_2043_n 0.00127908f $X=9.42 $Y=2.465 $X2=0
+ $Y2=0
cc_1074 N_A_1313_74#_c_1368_n N_VPWR_c_2043_n 0.0208457f $X=12.125 $Y=2.475
+ $X2=0 $Y2=0
cc_1075 N_A_1313_74#_c_1368_n N_VPWR_c_2044_n 0.021438f $X=12.125 $Y=2.475 $X2=0
+ $Y2=0
cc_1076 N_A_1313_74#_c_1358_n N_VPWR_c_2051_n 0.00413917f $X=8 $Y=1.765 $X2=0
+ $Y2=0
cc_1077 N_A_1313_74#_c_1362_n N_VPWR_c_2051_n 0.00445602f $X=9.42 $Y=2.465 $X2=0
+ $Y2=0
cc_1078 N_A_1313_74#_c_1347_n N_VPWR_c_2059_n 0.00461464f $X=12.345 $Y=1.885
+ $X2=0 $Y2=0
cc_1079 N_A_1313_74#_c_1358_n N_VPWR_c_2037_n 0.00415915f $X=8 $Y=1.765 $X2=0
+ $Y2=0
cc_1080 N_A_1313_74#_c_1362_n N_VPWR_c_2037_n 0.00894079f $X=9.42 $Y=2.465 $X2=0
+ $Y2=0
cc_1081 N_A_1313_74#_c_1347_n N_VPWR_c_2037_n 0.00838031f $X=12.345 $Y=1.885
+ $X2=0 $Y2=0
cc_1082 N_A_1313_74#_c_1368_n N_VPWR_c_2037_n 0.0717358f $X=12.125 $Y=2.475
+ $X2=0 $Y2=0
cc_1083 N_A_1313_74#_c_1370_n N_VPWR_c_2037_n 0.00699572f $X=9.435 $Y=2.165
+ $X2=0 $Y2=0
cc_1084 N_A_1313_74#_c_1353_n N_A_661_113#_c_2233_n 0.0031353f $X=6.87 $Y=0.925
+ $X2=0 $Y2=0
cc_1085 N_A_1313_74#_c_1366_n N_A_661_113#_c_2234_n 0.0131194f $X=7.245 $Y=1.975
+ $X2=0 $Y2=0
cc_1086 N_A_1313_74#_M1025_d N_A_661_113#_c_2245_n 0.00750239f $X=6.725 $Y=1.805
+ $X2=0 $Y2=0
cc_1087 N_A_1313_74#_c_1343_n N_A_661_113#_c_2245_n 0.0017945f $X=7.925 $Y=1.69
+ $X2=0 $Y2=0
cc_1088 N_A_1313_74#_c_1366_n N_A_661_113#_c_2245_n 0.0366312f $X=7.245 $Y=1.975
+ $X2=0 $Y2=0
cc_1089 N_A_1313_74#_c_1354_n N_A_661_113#_c_2245_n 0.0199529f $X=7.33 $Y=1.785
+ $X2=0 $Y2=0
cc_1090 N_A_1313_74#_c_1356_n N_A_661_113#_c_2245_n 0.00438727f $X=7.355 $Y=1.69
+ $X2=0 $Y2=0
cc_1091 N_A_1313_74#_c_1343_n N_A_661_113#_c_2246_n 0.00864063f $X=7.925 $Y=1.69
+ $X2=0 $Y2=0
cc_1092 N_A_1313_74#_c_1358_n N_A_661_113#_c_2246_n 0.00681616f $X=8 $Y=1.765
+ $X2=0 $Y2=0
cc_1093 N_A_1313_74#_c_1354_n N_A_661_113#_c_2246_n 0.0289113f $X=7.33 $Y=1.785
+ $X2=0 $Y2=0
cc_1094 N_A_1313_74#_c_1356_n N_A_661_113#_c_2246_n 0.0029034f $X=7.355 $Y=1.69
+ $X2=0 $Y2=0
cc_1095 N_A_1313_74#_c_1343_n N_A_661_113#_c_2235_n 0.00146076f $X=7.925 $Y=1.69
+ $X2=0 $Y2=0
cc_1096 N_A_1313_74#_c_1344_n N_A_661_113#_c_2235_n 0.00852537f $X=8.63 $Y=1.69
+ $X2=0 $Y2=0
cc_1097 N_A_1313_74#_M1040_g N_A_661_113#_c_2235_n 7.47252e-19 $X=8.705 $Y=0.695
+ $X2=0 $Y2=0
cc_1098 N_A_1313_74#_c_1349_n N_A_661_113#_c_2235_n 0.00636466f $X=8 $Y=1.69
+ $X2=0 $Y2=0
cc_1099 N_A_1313_74#_M1013_g N_A_661_113#_c_2236_n 0.0028423f $X=7.475 $Y=0.74
+ $X2=0 $Y2=0
cc_1100 N_A_1313_74#_c_1343_n N_A_661_113#_c_2236_n 0.00390297f $X=7.925 $Y=1.69
+ $X2=0 $Y2=0
cc_1101 N_A_1313_74#_c_1354_n N_A_661_113#_c_2236_n 0.0078668f $X=7.33 $Y=1.785
+ $X2=0 $Y2=0
cc_1102 N_A_1313_74#_c_1358_n N_A_661_113#_c_2247_n 0.0311109f $X=8 $Y=1.765
+ $X2=0 $Y2=0
cc_1103 N_A_1313_74#_M1013_g N_A_661_113#_c_2237_n 0.00639263f $X=7.475 $Y=0.74
+ $X2=0 $Y2=0
cc_1104 N_A_1313_74#_M1040_g N_A_661_113#_c_2237_n 0.00466103f $X=8.705 $Y=0.695
+ $X2=0 $Y2=0
cc_1105 N_A_1313_74#_c_1354_n N_A_661_113#_c_2237_n 0.00921645f $X=7.33 $Y=1.785
+ $X2=0 $Y2=0
cc_1106 N_A_1313_74#_c_1368_n A_1899_508# 0.00126545f $X=12.125 $Y=2.475
+ $X2=-0.19 $Y2=-0.245
cc_1107 N_A_1313_74#_c_1370_n A_1899_508# 0.00331222f $X=9.435 $Y=2.165
+ $X2=-0.19 $Y2=-0.245
cc_1108 N_A_1313_74#_c_1368_n A_2292_392# 0.0337585f $X=12.125 $Y=2.475
+ $X2=-0.19 $Y2=-0.245
cc_1109 N_A_1313_74#_c_1369_n A_2292_392# 0.00757088f $X=12.21 $Y=2.39 $X2=-0.19
+ $Y2=-0.245
cc_1110 N_A_1313_74#_c_1352_n N_VGND_M1013_s 0.00503458f $X=7.245 $Y=0.925 $X2=0
+ $Y2=0
cc_1111 N_A_1313_74#_c_1354_n N_VGND_M1013_s 0.00176713f $X=7.33 $Y=1.785 $X2=0
+ $Y2=0
cc_1112 N_A_1313_74#_c_1351_n N_VGND_c_2470_n 0.0182544f $X=6.705 $Y=0.515 $X2=0
+ $Y2=0
cc_1113 N_A_1313_74#_M1013_g N_VGND_c_2471_n 0.0088425f $X=7.475 $Y=0.74 $X2=0
+ $Y2=0
cc_1114 N_A_1313_74#_c_1351_n N_VGND_c_2471_n 0.0219045f $X=6.705 $Y=0.515 $X2=0
+ $Y2=0
cc_1115 N_A_1313_74#_c_1352_n N_VGND_c_2471_n 0.0216996f $X=7.245 $Y=0.925 $X2=0
+ $Y2=0
cc_1116 N_A_1313_74#_c_1351_n N_VGND_c_2481_n 0.0145323f $X=6.705 $Y=0.515 $X2=0
+ $Y2=0
cc_1117 N_A_1313_74#_M1013_g N_VGND_c_2486_n 0.00383152f $X=7.475 $Y=0.74 $X2=0
+ $Y2=0
cc_1118 N_A_1313_74#_M1040_g N_VGND_c_2486_n 7.53287e-19 $X=8.705 $Y=0.695 $X2=0
+ $Y2=0
cc_1119 N_A_1313_74#_M1016_g N_VGND_c_2495_n 0.00434272f $X=12.415 $Y=0.58 $X2=0
+ $Y2=0
cc_1120 N_A_1313_74#_M1016_g N_VGND_c_2496_n 0.00148617f $X=12.415 $Y=0.58 $X2=0
+ $Y2=0
cc_1121 N_A_1313_74#_M1013_g N_VGND_c_2499_n 0.00762539f $X=7.475 $Y=0.74 $X2=0
+ $Y2=0
cc_1122 N_A_1313_74#_M1016_g N_VGND_c_2499_n 0.00448332f $X=12.415 $Y=0.58 $X2=0
+ $Y2=0
cc_1123 N_A_1313_74#_c_1351_n N_VGND_c_2499_n 0.0119861f $X=6.705 $Y=0.515 $X2=0
+ $Y2=0
cc_1124 N_A_1313_74#_c_1352_n N_VGND_c_2499_n 0.00888394f $X=7.245 $Y=0.925
+ $X2=0 $Y2=0
cc_1125 N_A_1943_53#_c_1534_n N_A_1756_97#_c_1639_n 0.040416f $X=9.9 $Y=2.375
+ $X2=0 $Y2=0
cc_1126 N_A_1943_53#_c_1546_n N_A_1756_97#_c_1639_n 0.0103066f $X=9.9 $Y=2.465
+ $X2=0 $Y2=0
cc_1127 N_A_1943_53#_c_1535_n N_A_1756_97#_c_1639_n 0.00312006f $X=11.385
+ $Y=1.795 $X2=0 $Y2=0
cc_1128 N_A_1943_53#_c_1537_n N_A_1756_97#_c_1639_n 0.00452842f $X=10.6 $Y=1.285
+ $X2=0 $Y2=0
cc_1129 N_A_1943_53#_c_1549_n N_A_1756_97#_c_1639_n 0.00804707f $X=10.755
+ $Y=2.095 $X2=0 $Y2=0
cc_1130 N_A_1943_53#_c_1539_n N_A_1756_97#_c_1639_n 0.00656693f $X=10.84 $Y=1.97
+ $X2=0 $Y2=0
cc_1131 N_A_1943_53#_c_1540_n N_A_1756_97#_c_1639_n 0.00125647f $X=10.925
+ $Y=1.365 $X2=0 $Y2=0
cc_1132 N_A_1943_53#_c_1544_n N_A_1756_97#_c_1639_n 6.01846e-19 $X=11.385
+ $Y=1.32 $X2=0 $Y2=0
cc_1133 N_A_1943_53#_M1032_g N_A_1756_97#_M1046_g 0.0137291f $X=9.79 $Y=0.605
+ $X2=0 $Y2=0
cc_1134 N_A_1943_53#_c_1534_n N_A_1756_97#_M1046_g 3.31869e-19 $X=9.9 $Y=2.375
+ $X2=0 $Y2=0
cc_1135 N_A_1943_53#_c_1537_n N_A_1756_97#_M1046_g 0.0155121f $X=10.6 $Y=1.285
+ $X2=0 $Y2=0
cc_1136 N_A_1943_53#_c_1538_n N_A_1756_97#_M1046_g 0.0063093f $X=10.685 $Y=0.825
+ $X2=0 $Y2=0
cc_1137 N_A_1943_53#_c_1540_n N_A_1756_97#_M1046_g 0.00348498f $X=10.925
+ $Y=1.365 $X2=0 $Y2=0
cc_1138 N_A_1943_53#_c_1542_n N_A_1756_97#_M1046_g 0.0121102f $X=9.88 $Y=1.315
+ $X2=0 $Y2=0
cc_1139 N_A_1943_53#_c_1543_n N_A_1756_97#_M1046_g 2.02651e-19 $X=10.045
+ $Y=1.302 $X2=0 $Y2=0
cc_1140 N_A_1943_53#_c_1544_n N_A_1756_97#_M1046_g 0.00500556f $X=11.385 $Y=1.32
+ $X2=0 $Y2=0
cc_1141 N_A_1943_53#_c_1546_n N_A_1756_97#_c_1646_n 0.00157645f $X=9.9 $Y=2.465
+ $X2=0 $Y2=0
cc_1142 N_A_1943_53#_c_1534_n N_A_1756_97#_c_1642_n 7.04905e-19 $X=9.9 $Y=2.375
+ $X2=0 $Y2=0
cc_1143 N_A_1943_53#_c_1537_n N_A_1756_97#_c_1642_n 0.0218067f $X=10.6 $Y=1.285
+ $X2=0 $Y2=0
cc_1144 N_A_1943_53#_c_1549_n N_A_1756_97#_c_1642_n 0.00760086f $X=10.755
+ $Y=2.095 $X2=0 $Y2=0
cc_1145 N_A_1943_53#_c_1539_n N_A_1756_97#_c_1642_n 0.0187791f $X=10.84 $Y=1.97
+ $X2=0 $Y2=0
cc_1146 N_A_1943_53#_c_1534_n N_A_1756_97#_c_1643_n 0.0139188f $X=9.9 $Y=2.375
+ $X2=0 $Y2=0
cc_1147 N_A_1943_53#_c_1537_n N_A_1756_97#_c_1643_n 0.00890429f $X=10.6 $Y=1.285
+ $X2=0 $Y2=0
cc_1148 N_A_1943_53#_c_1542_n N_A_1756_97#_c_1643_n 0.00383582f $X=9.88 $Y=1.315
+ $X2=0 $Y2=0
cc_1149 N_A_1943_53#_c_1543_n N_A_1756_97#_c_1643_n 0.0149674f $X=10.045
+ $Y=1.302 $X2=0 $Y2=0
cc_1150 N_A_1943_53#_c_1546_n N_VPWR_c_2043_n 0.00966968f $X=9.9 $Y=2.465 $X2=0
+ $Y2=0
cc_1151 N_A_1943_53#_c_1548_n N_VPWR_c_2044_n 0.0183124f $X=11.385 $Y=1.885
+ $X2=0 $Y2=0
cc_1152 N_A_1943_53#_c_1546_n N_VPWR_c_2051_n 0.00413917f $X=9.9 $Y=2.465 $X2=0
+ $Y2=0
cc_1153 N_A_1943_53#_c_1548_n N_VPWR_c_2059_n 0.00413917f $X=11.385 $Y=1.885
+ $X2=0 $Y2=0
cc_1154 N_A_1943_53#_c_1546_n N_VPWR_c_2037_n 0.00398988f $X=9.9 $Y=2.465 $X2=0
+ $Y2=0
cc_1155 N_A_1943_53#_c_1548_n N_VPWR_c_2037_n 0.00403443f $X=11.385 $Y=1.885
+ $X2=0 $Y2=0
cc_1156 N_A_1943_53#_M1032_g N_VGND_c_2472_n 0.00862979f $X=9.79 $Y=0.605 $X2=0
+ $Y2=0
cc_1157 N_A_1943_53#_c_1536_n N_VGND_c_2473_n 0.0108108f $X=11.58 $Y=1.11 $X2=0
+ $Y2=0
cc_1158 N_A_1943_53#_M1032_g N_VGND_c_2486_n 0.00465077f $X=9.79 $Y=0.605 $X2=0
+ $Y2=0
cc_1159 N_A_1943_53#_c_1536_n N_VGND_c_2495_n 0.00383152f $X=11.58 $Y=1.11 $X2=0
+ $Y2=0
cc_1160 N_A_1943_53#_M1032_g N_VGND_c_2499_n 0.00451796f $X=9.79 $Y=0.605 $X2=0
+ $Y2=0
cc_1161 N_A_1943_53#_c_1536_n N_VGND_c_2499_n 0.00387546f $X=11.58 $Y=1.11 $X2=0
+ $Y2=0
cc_1162 N_A_1756_97#_c_1639_n N_VPWR_c_2043_n 0.00419996f $X=10.415 $Y=1.915
+ $X2=0 $Y2=0
cc_1163 N_A_1756_97#_c_1646_n N_VPWR_c_2043_n 0.00665231f $X=9.195 $Y=2.75 $X2=0
+ $Y2=0
cc_1164 N_A_1756_97#_c_1639_n N_VPWR_c_2044_n 0.00600586f $X=10.415 $Y=1.915
+ $X2=0 $Y2=0
cc_1165 N_A_1756_97#_c_1646_n N_VPWR_c_2051_n 0.015569f $X=9.195 $Y=2.75 $X2=0
+ $Y2=0
cc_1166 N_A_1756_97#_c_1639_n N_VPWR_c_2058_n 0.00487664f $X=10.415 $Y=1.915
+ $X2=0 $Y2=0
cc_1167 N_A_1756_97#_c_1639_n N_VPWR_c_2037_n 0.00505379f $X=10.415 $Y=1.915
+ $X2=0 $Y2=0
cc_1168 N_A_1756_97#_c_1646_n N_VPWR_c_2037_n 0.0128526f $X=9.195 $Y=2.75 $X2=0
+ $Y2=0
cc_1169 N_A_1756_97#_c_1647_n N_A_661_113#_c_2247_n 0.0439389f $X=9.18 $Y=2.52
+ $X2=0 $Y2=0
cc_1170 N_A_1756_97#_M1046_g N_VGND_c_2472_n 0.00123511f $X=10.47 $Y=0.715 $X2=0
+ $Y2=0
cc_1171 N_A_1756_97#_M1046_g N_VGND_c_2487_n 9.63466e-19 $X=10.47 $Y=0.715 $X2=0
+ $Y2=0
cc_1172 N_A_2403_74#_c_1742_n N_VPWR_c_2045_n 0.00634677f $X=13.985 $Y=2.245
+ $X2=0 $Y2=0
cc_1173 N_A_2403_74#_c_1749_n N_VPWR_c_2045_n 0.0121541f $X=12.63 $Y=2.75 $X2=0
+ $Y2=0
cc_1174 N_A_2403_74#_c_1742_n N_VPWR_c_2046_n 0.00445602f $X=13.985 $Y=2.245
+ $X2=0 $Y2=0
cc_1175 N_A_2403_74#_c_1742_n N_VPWR_c_2047_n 0.00429291f $X=13.985 $Y=2.245
+ $X2=0 $Y2=0
cc_1176 N_A_2403_74#_c_1729_n N_VPWR_c_2047_n 0.00378253f $X=14.865 $Y=1.537
+ $X2=0 $Y2=0
cc_1177 N_A_2403_74#_c_1744_n N_VPWR_c_2047_n 0.0153471f $X=14.955 $Y=1.765
+ $X2=0 $Y2=0
cc_1178 N_A_2403_74#_c_1745_n N_VPWR_c_2047_n 5.43055e-19 $X=15.405 $Y=1.765
+ $X2=0 $Y2=0
cc_1179 N_A_2403_74#_c_1744_n N_VPWR_c_2048_n 5.08113e-19 $X=14.955 $Y=1.765
+ $X2=0 $Y2=0
cc_1180 N_A_2403_74#_c_1745_n N_VPWR_c_2048_n 0.01067f $X=15.405 $Y=1.765 $X2=0
+ $Y2=0
cc_1181 N_A_2403_74#_c_1746_n N_VPWR_c_2048_n 0.0105935f $X=15.855 $Y=1.765
+ $X2=0 $Y2=0
cc_1182 N_A_2403_74#_c_1747_n N_VPWR_c_2048_n 5.03387e-19 $X=16.305 $Y=1.765
+ $X2=0 $Y2=0
cc_1183 N_A_2403_74#_c_1734_n N_VPWR_c_2048_n 7.29495e-19 $X=16.305 $Y=1.58
+ $X2=0 $Y2=0
cc_1184 N_A_2403_74#_c_1746_n N_VPWR_c_2050_n 5.08113e-19 $X=15.855 $Y=1.765
+ $X2=0 $Y2=0
cc_1185 N_A_2403_74#_c_1747_n N_VPWR_c_2050_n 0.0118145f $X=16.305 $Y=1.765
+ $X2=0 $Y2=0
cc_1186 N_A_2403_74#_c_1749_n N_VPWR_c_2059_n 0.018757f $X=12.63 $Y=2.75 $X2=0
+ $Y2=0
cc_1187 N_A_2403_74#_c_1744_n N_VPWR_c_2060_n 0.00413917f $X=14.955 $Y=1.765
+ $X2=0 $Y2=0
cc_1188 N_A_2403_74#_c_1745_n N_VPWR_c_2060_n 0.00413917f $X=15.405 $Y=1.765
+ $X2=0 $Y2=0
cc_1189 N_A_2403_74#_c_1746_n N_VPWR_c_2061_n 0.00413917f $X=15.855 $Y=1.765
+ $X2=0 $Y2=0
cc_1190 N_A_2403_74#_c_1747_n N_VPWR_c_2061_n 0.00413917f $X=16.305 $Y=1.765
+ $X2=0 $Y2=0
cc_1191 N_A_2403_74#_c_1742_n N_VPWR_c_2037_n 0.00863669f $X=13.985 $Y=2.245
+ $X2=0 $Y2=0
cc_1192 N_A_2403_74#_c_1744_n N_VPWR_c_2037_n 0.00817726f $X=14.955 $Y=1.765
+ $X2=0 $Y2=0
cc_1193 N_A_2403_74#_c_1745_n N_VPWR_c_2037_n 0.00817726f $X=15.405 $Y=1.765
+ $X2=0 $Y2=0
cc_1194 N_A_2403_74#_c_1746_n N_VPWR_c_2037_n 0.00817726f $X=15.855 $Y=1.765
+ $X2=0 $Y2=0
cc_1195 N_A_2403_74#_c_1747_n N_VPWR_c_2037_n 0.00817726f $X=16.305 $Y=1.765
+ $X2=0 $Y2=0
cc_1196 N_A_2403_74#_c_1749_n N_VPWR_c_2037_n 0.0152576f $X=12.63 $Y=2.75 $X2=0
+ $Y2=0
cc_1197 N_A_2403_74#_c_1744_n N_Q_c_2418_n 4.77902e-19 $X=14.955 $Y=1.765 $X2=0
+ $Y2=0
cc_1198 N_A_2403_74#_c_1745_n N_Q_c_2418_n 4.71103e-19 $X=15.405 $Y=1.765 $X2=0
+ $Y2=0
cc_1199 N_A_2403_74#_c_1730_n N_Q_c_2415_n 3.97481e-19 $X=14.945 $Y=1.395 $X2=0
+ $Y2=0
cc_1200 N_A_2403_74#_c_1731_n N_Q_c_2415_n 0.00813388f $X=15.375 $Y=1.395 $X2=0
+ $Y2=0
cc_1201 N_A_2403_74#_c_1732_n N_Q_c_2415_n 5.93572e-19 $X=15.875 $Y=1.395 $X2=0
+ $Y2=0
cc_1202 N_A_2403_74#_c_1746_n N_Q_c_2419_n 4.74176e-19 $X=15.855 $Y=1.765 $X2=0
+ $Y2=0
cc_1203 N_A_2403_74#_c_1747_n N_Q_c_2419_n 4.70785e-19 $X=16.305 $Y=1.765 $X2=0
+ $Y2=0
cc_1204 N_A_2403_74#_c_1732_n N_Q_c_2416_n 2.36759e-19 $X=15.875 $Y=1.395 $X2=0
+ $Y2=0
cc_1205 N_A_2403_74#_c_1733_n N_Q_c_2416_n 2.36759e-19 $X=16.32 $Y=1.395 $X2=0
+ $Y2=0
cc_1206 N_A_2403_74#_c_1730_n Q 0.00171856f $X=14.945 $Y=1.395 $X2=0 $Y2=0
cc_1207 N_A_2403_74#_c_1744_n Q 0.00167228f $X=14.955 $Y=1.765 $X2=0 $Y2=0
cc_1208 N_A_2403_74#_c_1731_n Q 0.0129525f $X=15.375 $Y=1.395 $X2=0 $Y2=0
cc_1209 N_A_2403_74#_c_1745_n Q 0.0179427f $X=15.405 $Y=1.765 $X2=0 $Y2=0
cc_1210 N_A_2403_74#_c_1746_n Q 0.0178583f $X=15.855 $Y=1.765 $X2=0 $Y2=0
cc_1211 N_A_2403_74#_c_1732_n Q 0.015929f $X=15.875 $Y=1.395 $X2=0 $Y2=0
cc_1212 N_A_2403_74#_c_1747_n Q 0.0212283f $X=16.305 $Y=1.765 $X2=0 $Y2=0
cc_1213 N_A_2403_74#_c_1733_n Q 0.0177773f $X=16.32 $Y=1.395 $X2=0 $Y2=0
cc_1214 N_A_2403_74#_c_1734_n Q 0.0918412f $X=16.305 $Y=1.58 $X2=0 $Y2=0
cc_1215 N_A_2403_74#_c_1735_n N_VGND_c_2473_n 0.00539463f $X=12.2 $Y=0.58 $X2=0
+ $Y2=0
cc_1216 N_A_2403_74#_M1021_g N_VGND_c_2474_n 0.00434272f $X=13.955 $Y=0.58 $X2=0
+ $Y2=0
cc_1217 N_A_2403_74#_M1021_g N_VGND_c_2475_n 0.00348962f $X=13.955 $Y=0.58 $X2=0
+ $Y2=0
cc_1218 N_A_2403_74#_c_1729_n N_VGND_c_2475_n 0.00592208f $X=14.865 $Y=1.537
+ $X2=0 $Y2=0
cc_1219 N_A_2403_74#_c_1730_n N_VGND_c_2475_n 0.0155123f $X=14.945 $Y=1.395
+ $X2=0 $Y2=0
cc_1220 N_A_2403_74#_c_1731_n N_VGND_c_2475_n 6.10916e-19 $X=15.375 $Y=1.395
+ $X2=0 $Y2=0
cc_1221 N_A_2403_74#_c_1731_n N_VGND_c_2476_n 0.00357456f $X=15.375 $Y=1.395
+ $X2=0 $Y2=0
cc_1222 N_A_2403_74#_c_1732_n N_VGND_c_2476_n 0.00815698f $X=15.875 $Y=1.395
+ $X2=0 $Y2=0
cc_1223 N_A_2403_74#_c_1733_n N_VGND_c_2476_n 4.66019e-19 $X=16.32 $Y=1.395
+ $X2=0 $Y2=0
cc_1224 N_A_2403_74#_c_1734_n N_VGND_c_2476_n 6.99498e-19 $X=16.305 $Y=1.58
+ $X2=0 $Y2=0
cc_1225 N_A_2403_74#_c_1732_n N_VGND_c_2478_n 4.66019e-19 $X=15.875 $Y=1.395
+ $X2=0 $Y2=0
cc_1226 N_A_2403_74#_c_1733_n N_VGND_c_2478_n 0.00921274f $X=16.32 $Y=1.395
+ $X2=0 $Y2=0
cc_1227 N_A_2403_74#_c_1730_n N_VGND_c_2488_n 0.00365567f $X=14.945 $Y=1.395
+ $X2=0 $Y2=0
cc_1228 N_A_2403_74#_c_1731_n N_VGND_c_2488_n 0.00422883f $X=15.375 $Y=1.395
+ $X2=0 $Y2=0
cc_1229 N_A_2403_74#_c_1732_n N_VGND_c_2489_n 0.00365567f $X=15.875 $Y=1.395
+ $X2=0 $Y2=0
cc_1230 N_A_2403_74#_c_1733_n N_VGND_c_2489_n 0.00365567f $X=16.32 $Y=1.395
+ $X2=0 $Y2=0
cc_1231 N_A_2403_74#_c_1735_n N_VGND_c_2495_n 0.0145482f $X=12.2 $Y=0.58 $X2=0
+ $Y2=0
cc_1232 N_A_2403_74#_M1021_g N_VGND_c_2496_n 0.0115871f $X=13.955 $Y=0.58 $X2=0
+ $Y2=0
cc_1233 N_A_2403_74#_c_1735_n N_VGND_c_2496_n 0.0110541f $X=12.2 $Y=0.58 $X2=0
+ $Y2=0
cc_1234 N_A_2403_74#_c_1736_n N_VGND_c_2496_n 0.068269f $X=13.265 $Y=0.935 $X2=0
+ $Y2=0
cc_1235 N_A_2403_74#_c_1739_n N_VGND_c_2496_n 7.56504e-19 $X=13.89 $Y=1.145
+ $X2=0 $Y2=0
cc_1236 N_A_2403_74#_M1021_g N_VGND_c_2499_n 0.00830035f $X=13.955 $Y=0.58 $X2=0
+ $Y2=0
cc_1237 N_A_2403_74#_c_1730_n N_VGND_c_2499_n 0.00404919f $X=14.945 $Y=1.395
+ $X2=0 $Y2=0
cc_1238 N_A_2403_74#_c_1731_n N_VGND_c_2499_n 0.00482046f $X=15.375 $Y=1.395
+ $X2=0 $Y2=0
cc_1239 N_A_2403_74#_c_1732_n N_VGND_c_2499_n 0.00404919f $X=15.875 $Y=1.395
+ $X2=0 $Y2=0
cc_1240 N_A_2403_74#_c_1733_n N_VGND_c_2499_n 0.00404919f $X=16.32 $Y=1.395
+ $X2=0 $Y2=0
cc_1241 N_A_2403_74#_c_1735_n N_VGND_c_2499_n 0.0119922f $X=12.2 $Y=0.58 $X2=0
+ $Y2=0
cc_1242 N_A_2403_74#_c_1736_n N_VGND_c_2499_n 0.0168873f $X=13.265 $Y=0.935
+ $X2=0 $Y2=0
cc_1243 N_A_37_464#_c_1919_n A_126_464# 0.00595227f $X=1.455 $Y=2.375 $X2=-0.19
+ $Y2=-0.245
cc_1244 N_A_37_464#_c_1919_n N_VPWR_M1037_d 0.00509381f $X=1.455 $Y=2.375
+ $X2=-0.19 $Y2=-0.245
cc_1245 N_A_37_464#_c_1921_n N_VPWR_M1001_d 4.76982e-19 $X=2.135 $Y=2.99 $X2=0
+ $Y2=0
cc_1246 N_A_37_464#_c_1954_n N_VPWR_M1001_d 0.00490162f $X=2.22 $Y=2.905 $X2=0
+ $Y2=0
cc_1247 N_A_37_464#_c_1923_n N_VPWR_M1001_d 0.00972296f $X=3.235 $Y=2.375 $X2=0
+ $Y2=0
cc_1248 N_A_37_464#_c_1918_n N_VPWR_c_2038_n 0.010138f $X=0.33 $Y=2.465 $X2=0
+ $Y2=0
cc_1249 N_A_37_464#_c_1919_n N_VPWR_c_2038_n 0.0154248f $X=1.455 $Y=2.375 $X2=0
+ $Y2=0
cc_1250 N_A_37_464#_c_1920_n N_VPWR_c_2038_n 0.0208967f $X=1.54 $Y=2.905 $X2=0
+ $Y2=0
cc_1251 N_A_37_464#_c_1922_n N_VPWR_c_2038_n 0.0146662f $X=1.625 $Y=2.99 $X2=0
+ $Y2=0
cc_1252 N_A_37_464#_c_1921_n N_VPWR_c_2039_n 0.0145842f $X=2.135 $Y=2.99 $X2=0
+ $Y2=0
cc_1253 N_A_37_464#_c_1954_n N_VPWR_c_2039_n 0.0205316f $X=2.22 $Y=2.905 $X2=0
+ $Y2=0
cc_1254 N_A_37_464#_c_1923_n N_VPWR_c_2039_n 0.0154248f $X=3.235 $Y=2.375 $X2=0
+ $Y2=0
cc_1255 N_A_37_464#_c_1925_n N_VPWR_c_2039_n 0.0101141f $X=3.4 $Y=2.46 $X2=0
+ $Y2=0
cc_1256 N_A_37_464#_c_1918_n N_VPWR_c_2053_n 0.0181748f $X=0.33 $Y=2.465 $X2=0
+ $Y2=0
cc_1257 N_A_37_464#_c_1921_n N_VPWR_c_2054_n 0.0445209f $X=2.135 $Y=2.99 $X2=0
+ $Y2=0
cc_1258 N_A_37_464#_c_1922_n N_VPWR_c_2054_n 0.0121867f $X=1.625 $Y=2.99 $X2=0
+ $Y2=0
cc_1259 N_A_37_464#_c_1925_n N_VPWR_c_2055_n 0.0108086f $X=3.4 $Y=2.46 $X2=0
+ $Y2=0
cc_1260 N_A_37_464#_c_1918_n N_VPWR_c_2037_n 0.0150057f $X=0.33 $Y=2.465 $X2=0
+ $Y2=0
cc_1261 N_A_37_464#_c_1921_n N_VPWR_c_2037_n 0.0250929f $X=2.135 $Y=2.99 $X2=0
+ $Y2=0
cc_1262 N_A_37_464#_c_1922_n N_VPWR_c_2037_n 0.00660921f $X=1.625 $Y=2.99 $X2=0
+ $Y2=0
cc_1263 N_A_37_464#_c_1925_n N_VPWR_c_2037_n 0.00906495f $X=3.4 $Y=2.46 $X2=0
+ $Y2=0
cc_1264 N_A_37_464#_c_1923_n A_572_463# 0.0048076f $X=3.235 $Y=2.375 $X2=-0.19
+ $Y2=-0.245
cc_1265 N_A_37_464#_c_1925_n N_A_661_113#_c_2309_n 0.033328f $X=3.4 $Y=2.46
+ $X2=0 $Y2=0
cc_1266 N_A_37_464#_c_1925_n N_A_661_113#_c_2253_n 0.00568204f $X=3.4 $Y=2.46
+ $X2=0 $Y2=0
cc_1267 N_A_37_464#_c_1913_n N_A_661_113#_c_2238_n 0.0131609f $X=3.015 $Y=0.775
+ $X2=0 $Y2=0
cc_1268 N_A_37_464#_c_1916_n N_A_661_113#_c_2238_n 0.00990851f $X=3.4 $Y=1.26
+ $X2=0 $Y2=0
cc_1269 N_A_37_464#_c_1913_n N_A_661_113#_c_2239_n 0.00545722f $X=3.015 $Y=0.775
+ $X2=0 $Y2=0
cc_1270 N_A_37_464#_c_1914_n N_A_661_113#_c_2239_n 0.0700563f $X=3.4 $Y=2.29
+ $X2=0 $Y2=0
cc_1271 N_A_37_464#_c_1916_n N_A_661_113#_c_2239_n 0.0138286f $X=3.4 $Y=1.26
+ $X2=0 $Y2=0
cc_1272 N_A_37_464#_c_1928_n N_A_661_113#_c_2239_n 0.0138383f $X=3.36 $Y=2.375
+ $X2=0 $Y2=0
cc_1273 N_A_37_464#_c_1915_n N_VGND_c_2467_n 0.015258f $X=0.385 $Y=0.575 $X2=0
+ $Y2=0
cc_1274 N_A_37_464#_c_1913_n N_VGND_c_2468_n 0.0145731f $X=3.015 $Y=0.775 $X2=0
+ $Y2=0
cc_1275 N_A_37_464#_c_1915_n N_VGND_c_2483_n 0.0208797f $X=0.385 $Y=0.575 $X2=0
+ $Y2=0
cc_1276 N_A_37_464#_c_1913_n N_VGND_c_2485_n 0.00794834f $X=3.015 $Y=0.775 $X2=0
+ $Y2=0
cc_1277 N_A_37_464#_c_1913_n N_VGND_c_2499_n 0.0105391f $X=3.015 $Y=0.775 $X2=0
+ $Y2=0
cc_1278 N_A_37_464#_c_1915_n N_VGND_c_2499_n 0.0169374f $X=0.385 $Y=0.575 $X2=0
+ $Y2=0
cc_1279 N_VPWR_c_2040_n N_A_661_113#_c_2242_n 0.0147124f $X=5.055 $Y=2.765 $X2=0
+ $Y2=0
cc_1280 N_VPWR_c_2055_n N_A_661_113#_c_2242_n 0.0546448f $X=4.97 $Y=3.33 $X2=0
+ $Y2=0
cc_1281 N_VPWR_c_2037_n N_A_661_113#_c_2242_n 0.0292625f $X=16.56 $Y=3.33 $X2=0
+ $Y2=0
cc_1282 N_VPWR_c_2055_n N_A_661_113#_c_2253_n 0.0190556f $X=4.97 $Y=3.33 $X2=0
+ $Y2=0
cc_1283 N_VPWR_c_2037_n N_A_661_113#_c_2253_n 0.00957028f $X=16.56 $Y=3.33 $X2=0
+ $Y2=0
cc_1284 N_VPWR_M1044_d N_A_661_113#_c_2269_n 0.00522241f $X=4.675 $Y=2.275 $X2=0
+ $Y2=0
cc_1285 N_VPWR_c_2040_n N_A_661_113#_c_2269_n 0.0231493f $X=5.055 $Y=2.765 $X2=0
+ $Y2=0
cc_1286 N_VPWR_M1025_s N_A_661_113#_c_2245_n 0.007768f $X=6.295 $Y=1.805 $X2=0
+ $Y2=0
cc_1287 N_VPWR_M1029_s N_A_661_113#_c_2245_n 0.00196153f $X=7.65 $Y=1.84 $X2=0
+ $Y2=0
cc_1288 N_VPWR_c_2041_n N_A_661_113#_c_2245_n 0.0215269f $X=6.425 $Y=2.77 $X2=0
+ $Y2=0
cc_1289 N_VPWR_c_2042_n N_A_661_113#_c_2245_n 0.00874606f $X=7.775 $Y=2.785
+ $X2=0 $Y2=0
cc_1290 N_VPWR_c_2037_n N_A_661_113#_c_2245_n 0.0367495f $X=16.56 $Y=3.33 $X2=0
+ $Y2=0
cc_1291 N_VPWR_M1029_s N_A_661_113#_c_2246_n 0.0115959f $X=7.65 $Y=1.84 $X2=0
+ $Y2=0
cc_1292 N_VPWR_c_2042_n N_A_661_113#_c_2247_n 0.0220369f $X=7.775 $Y=2.785 $X2=0
+ $Y2=0
cc_1293 N_VPWR_c_2051_n N_A_661_113#_c_2247_n 0.0295144f $X=9.96 $Y=3.33 $X2=0
+ $Y2=0
cc_1294 N_VPWR_c_2037_n N_A_661_113#_c_2247_n 0.0314214f $X=16.56 $Y=3.33 $X2=0
+ $Y2=0
cc_1295 N_VPWR_c_2040_n N_A_661_113#_c_2249_n 0.0101841f $X=5.055 $Y=2.765 $X2=0
+ $Y2=0
cc_1296 N_VPWR_c_2041_n N_A_661_113#_c_2249_n 0.0193156f $X=6.425 $Y=2.77 $X2=0
+ $Y2=0
cc_1297 N_VPWR_c_2056_n N_A_661_113#_c_2249_n 0.0119549f $X=6.26 $Y=3.33 $X2=0
+ $Y2=0
cc_1298 N_VPWR_c_2037_n N_A_661_113#_c_2249_n 0.011576f $X=16.56 $Y=3.33 $X2=0
+ $Y2=0
cc_1299 N_VPWR_M1044_d N_A_661_113#_c_2250_n 0.00977001f $X=4.675 $Y=2.275 $X2=0
+ $Y2=0
cc_1300 N_VPWR_c_2040_n N_A_661_113#_c_2250_n 0.0154248f $X=5.055 $Y=2.765 $X2=0
+ $Y2=0
cc_1301 N_VPWR_c_2037_n N_A_661_113#_c_2251_n 0.00725008f $X=16.56 $Y=3.33 $X2=0
+ $Y2=0
cc_1302 N_VPWR_M1029_s N_A_661_113#_c_2398_n 0.00183801f $X=7.65 $Y=1.84 $X2=0
+ $Y2=0
cc_1303 N_VPWR_c_2042_n N_A_661_113#_c_2398_n 0.0129606f $X=7.775 $Y=2.785 $X2=0
+ $Y2=0
cc_1304 N_VPWR_c_2037_n N_A_661_113#_c_2398_n 6.28937e-19 $X=16.56 $Y=3.33 $X2=0
+ $Y2=0
cc_1305 N_VPWR_c_2047_n N_Q_c_2418_n 0.031887f $X=14.73 $Y=2.035 $X2=0 $Y2=0
cc_1306 N_VPWR_c_2048_n N_Q_c_2418_n 0.0243693f $X=15.63 $Y=2.405 $X2=0 $Y2=0
cc_1307 N_VPWR_c_2060_n N_Q_c_2418_n 0.00972736f $X=15.465 $Y=3.33 $X2=0 $Y2=0
cc_1308 N_VPWR_c_2037_n N_Q_c_2418_n 0.00805147f $X=16.56 $Y=3.33 $X2=0 $Y2=0
cc_1309 N_VPWR_c_2048_n N_Q_c_2419_n 0.0249212f $X=15.63 $Y=2.405 $X2=0 $Y2=0
cc_1310 N_VPWR_c_2050_n N_Q_c_2419_n 0.0243668f $X=16.53 $Y=2.405 $X2=0 $Y2=0
cc_1311 N_VPWR_c_2061_n N_Q_c_2419_n 0.00950426f $X=16.365 $Y=3.33 $X2=0 $Y2=0
cc_1312 N_VPWR_c_2037_n N_Q_c_2419_n 0.0078668f $X=16.56 $Y=3.33 $X2=0 $Y2=0
cc_1313 N_VPWR_M1009_d Q 0.00205832f $X=15.48 $Y=1.84 $X2=0 $Y2=0
cc_1314 N_VPWR_M1028_d Q 0.00423758f $X=16.38 $Y=1.84 $X2=0 $Y2=0
cc_1315 N_VPWR_c_2048_n Q 0.0190557f $X=15.63 $Y=2.405 $X2=0 $Y2=0
cc_1316 N_VPWR_c_2050_n Q 0.0226366f $X=16.53 $Y=2.405 $X2=0 $Y2=0
cc_1317 N_VPWR_c_2047_n N_VGND_c_2475_n 0.00323216f $X=14.73 $Y=2.035 $X2=0
+ $Y2=0
cc_1318 N_A_661_113#_c_2250_n A_1071_455# 0.0048076f $X=5.73 $Y=2.38 $X2=-0.19
+ $Y2=-0.245
cc_1319 N_A_661_113#_c_2240_n N_VGND_M1026_s 0.00135398f $X=6.115 $Y=1.16 $X2=0
+ $Y2=0
cc_1320 N_A_661_113#_c_2233_n N_VGND_c_2469_n 0.0135502f $X=5.72 $Y=0.835 $X2=0
+ $Y2=0
cc_1321 N_A_661_113#_c_2233_n N_VGND_c_2470_n 0.0201128f $X=5.72 $Y=0.835 $X2=0
+ $Y2=0
cc_1322 N_A_661_113#_c_2240_n N_VGND_c_2470_n 0.00729985f $X=6.115 $Y=1.16 $X2=0
+ $Y2=0
cc_1323 N_A_661_113#_c_2233_n N_VGND_c_2479_n 0.00683013f $X=5.72 $Y=0.835 $X2=0
+ $Y2=0
cc_1324 N_A_661_113#_c_2238_n N_VGND_c_2485_n 0.00788726f $X=3.74 $Y=0.84 $X2=0
+ $Y2=0
cc_1325 N_A_661_113#_c_2233_n N_VGND_c_2499_n 0.00988536f $X=5.72 $Y=0.835 $X2=0
+ $Y2=0
cc_1326 N_A_661_113#_c_2238_n N_VGND_c_2499_n 0.0135252f $X=3.74 $Y=0.84 $X2=0
+ $Y2=0
cc_1327 Q N_VGND_M1039_s 0.00261163f $X=16.475 $Y=1.21 $X2=0 $Y2=0
cc_1328 Q N_VGND_M1042_s 0.00350286f $X=16.475 $Y=1.21 $X2=0 $Y2=0
cc_1329 N_Q_c_2415_n N_VGND_c_2475_n 0.0197239f $X=15.16 $Y=0.725 $X2=0 $Y2=0
cc_1330 Q N_VGND_c_2475_n 0.00985092f $X=16.475 $Y=1.21 $X2=0 $Y2=0
cc_1331 N_Q_c_2415_n N_VGND_c_2476_n 0.0137359f $X=15.16 $Y=0.725 $X2=0 $Y2=0
cc_1332 N_Q_c_2416_n N_VGND_c_2476_n 0.0131001f $X=16.095 $Y=0.74 $X2=0 $Y2=0
cc_1333 Q N_VGND_c_2476_n 0.0232675f $X=16.475 $Y=1.21 $X2=0 $Y2=0
cc_1334 N_Q_c_2416_n N_VGND_c_2478_n 0.0131001f $X=16.095 $Y=0.74 $X2=0 $Y2=0
cc_1335 Q N_VGND_c_2478_n 0.0221307f $X=16.475 $Y=1.21 $X2=0 $Y2=0
cc_1336 N_Q_c_2415_n N_VGND_c_2488_n 0.00586114f $X=15.16 $Y=0.725 $X2=0 $Y2=0
cc_1337 N_Q_c_2416_n N_VGND_c_2489_n 0.00468116f $X=16.095 $Y=0.74 $X2=0 $Y2=0
cc_1338 N_Q_c_2415_n N_VGND_c_2499_n 0.00792225f $X=15.16 $Y=0.725 $X2=0 $Y2=0
cc_1339 N_Q_c_2416_n N_VGND_c_2499_n 0.0064368f $X=16.095 $Y=0.74 $X2=0 $Y2=0
