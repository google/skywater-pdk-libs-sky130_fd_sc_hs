* File: sky130_fd_sc_hs__sdfrbp_1.pxi.spice
* Created: Tue Sep  1 20:22:19 2020
* 
x_PM_SKY130_FD_SC_HS__SDFRBP_1%A_27_74# N_A_27_74#_M1040_s N_A_27_74#_M1027_s
+ N_A_27_74#_c_288_n N_A_27_74#_M1021_g N_A_27_74#_c_294_n N_A_27_74#_M1014_g
+ N_A_27_74#_c_289_n N_A_27_74#_c_290_n N_A_27_74#_c_291_n N_A_27_74#_c_292_n
+ N_A_27_74#_c_296_n N_A_27_74#_c_293_n N_A_27_74#_c_297_n N_A_27_74#_c_298_n
+ PM_SKY130_FD_SC_HS__SDFRBP_1%A_27_74#
x_PM_SKY130_FD_SC_HS__SDFRBP_1%SCE N_SCE_M1040_g N_SCE_c_378_n N_SCE_c_379_n
+ N_SCE_M1027_g N_SCE_c_380_n N_SCE_c_381_n N_SCE_M1024_g N_SCE_M1033_g
+ N_SCE_c_370_n N_SCE_c_371_n N_SCE_c_372_n N_SCE_c_373_n SCE SCE SCE
+ N_SCE_c_374_n N_SCE_c_375_n N_SCE_c_376_n SCE N_SCE_c_377_n
+ PM_SKY130_FD_SC_HS__SDFRBP_1%SCE
x_PM_SKY130_FD_SC_HS__SDFRBP_1%D N_D_M1000_g N_D_c_457_n N_D_c_462_n N_D_M1009_g
+ D N_D_c_458_n N_D_c_459_n N_D_c_460_n PM_SKY130_FD_SC_HS__SDFRBP_1%D
x_PM_SKY130_FD_SC_HS__SDFRBP_1%SCD N_SCD_c_505_n N_SCD_M1032_g N_SCD_M1015_g
+ N_SCD_c_502_n SCD SCD N_SCD_c_504_n PM_SKY130_FD_SC_HS__SDFRBP_1%SCD
x_PM_SKY130_FD_SC_HS__SDFRBP_1%RESET_B N_RESET_B_M1034_g N_RESET_B_c_553_n
+ N_RESET_B_M1020_g N_RESET_B_M1017_g N_RESET_B_c_554_n N_RESET_B_M1011_g
+ N_RESET_B_c_547_n N_RESET_B_M1007_g N_RESET_B_M1026_g N_RESET_B_c_549_n
+ N_RESET_B_c_550_n N_RESET_B_c_556_n N_RESET_B_c_557_n N_RESET_B_c_558_n
+ N_RESET_B_c_559_n N_RESET_B_c_560_n N_RESET_B_c_561_n RESET_B
+ N_RESET_B_c_563_n N_RESET_B_c_564_n N_RESET_B_c_565_n N_RESET_B_c_566_n
+ N_RESET_B_c_567_n N_RESET_B_c_568_n N_RESET_B_c_551_n
+ PM_SKY130_FD_SC_HS__SDFRBP_1%RESET_B
x_PM_SKY130_FD_SC_HS__SDFRBP_1%CLK N_CLK_c_765_n N_CLK_M1035_g N_CLK_c_766_n
+ N_CLK_M1025_g N_CLK_c_767_n CLK N_CLK_c_768_n PM_SKY130_FD_SC_HS__SDFRBP_1%CLK
x_PM_SKY130_FD_SC_HS__SDFRBP_1%A_1023_74# N_A_1023_74#_M1036_d
+ N_A_1023_74#_M1038_d N_A_1023_74#_c_833_n N_A_1023_74#_c_834_n
+ N_A_1023_74#_M1028_g N_A_1023_74#_c_813_n N_A_1023_74#_M1004_g
+ N_A_1023_74#_c_815_n N_A_1023_74#_M1030_g N_A_1023_74#_c_816_n
+ N_A_1023_74#_c_817_n N_A_1023_74#_c_836_n N_A_1023_74#_M1001_g
+ N_A_1023_74#_c_818_n N_A_1023_74#_c_819_n N_A_1023_74#_c_820_n
+ N_A_1023_74#_c_821_n N_A_1023_74#_c_822_n N_A_1023_74#_c_823_n
+ N_A_1023_74#_c_824_n N_A_1023_74#_c_848_n N_A_1023_74#_c_863_p
+ N_A_1023_74#_c_850_n N_A_1023_74#_c_825_n N_A_1023_74#_c_826_n
+ N_A_1023_74#_c_944_p N_A_1023_74#_c_827_n N_A_1023_74#_c_839_n
+ N_A_1023_74#_c_828_n N_A_1023_74#_c_829_n N_A_1023_74#_c_830_n
+ N_A_1023_74#_c_831_n N_A_1023_74#_c_832_n
+ PM_SKY130_FD_SC_HS__SDFRBP_1%A_1023_74#
x_PM_SKY130_FD_SC_HS__SDFRBP_1%A_1369_71# N_A_1369_71#_M1041_d
+ N_A_1369_71#_M1019_d N_A_1369_71#_M1016_g N_A_1369_71#_c_1031_n
+ N_A_1369_71#_c_1032_n N_A_1369_71#_M1018_g N_A_1369_71#_c_1023_n
+ N_A_1369_71#_c_1024_n N_A_1369_71#_c_1025_n N_A_1369_71#_c_1026_n
+ N_A_1369_71#_c_1068_n N_A_1369_71#_c_1027_n N_A_1369_71#_c_1028_n
+ N_A_1369_71#_c_1029_n N_A_1369_71#_c_1030_n
+ PM_SKY130_FD_SC_HS__SDFRBP_1%A_1369_71#
x_PM_SKY130_FD_SC_HS__SDFRBP_1%A_1221_97# N_A_1221_97#_M1012_d
+ N_A_1221_97#_M1028_d N_A_1221_97#_M1011_d N_A_1221_97#_M1041_g
+ N_A_1221_97#_c_1137_n N_A_1221_97#_M1019_g N_A_1221_97#_c_1131_n
+ N_A_1221_97#_c_1138_n N_A_1221_97#_c_1132_n N_A_1221_97#_c_1148_n
+ N_A_1221_97#_c_1133_n N_A_1221_97#_c_1134_n N_A_1221_97#_c_1135_n
+ N_A_1221_97#_c_1141_n N_A_1221_97#_c_1136_n
+ PM_SKY130_FD_SC_HS__SDFRBP_1%A_1221_97#
x_PM_SKY130_FD_SC_HS__SDFRBP_1%A_850_74# N_A_850_74#_M1035_s N_A_850_74#_M1025_s
+ N_A_850_74#_c_1245_n N_A_850_74#_M1036_g N_A_850_74#_c_1246_n
+ N_A_850_74#_M1038_g N_A_850_74#_c_1247_n N_A_850_74#_c_1248_n
+ N_A_850_74#_c_1249_n N_A_850_74#_c_1262_n N_A_850_74#_c_1263_n
+ N_A_850_74#_M1012_g N_A_850_74#_c_1264_n N_A_850_74#_c_1265_n
+ N_A_850_74#_c_1266_n N_A_850_74#_M1037_g N_A_850_74#_c_1267_n
+ N_A_850_74#_c_1268_n N_A_850_74#_c_1269_n N_A_850_74#_M1023_g
+ N_A_850_74#_c_1251_n N_A_850_74#_c_1252_n N_A_850_74#_M1013_g
+ N_A_850_74#_c_1254_n N_A_850_74#_c_1273_n N_A_850_74#_c_1255_n
+ N_A_850_74#_c_1256_n N_A_850_74#_c_1299_n N_A_850_74#_c_1274_n
+ N_A_850_74#_c_1257_n N_A_850_74#_c_1258_n N_A_850_74#_c_1276_n
+ N_A_850_74#_c_1259_n PM_SKY130_FD_SC_HS__SDFRBP_1%A_850_74#
x_PM_SKY130_FD_SC_HS__SDFRBP_1%A_2008_48# N_A_2008_48#_M1010_d
+ N_A_2008_48#_M1026_d N_A_2008_48#_M1005_g N_A_2008_48#_c_1438_n
+ N_A_2008_48#_c_1445_n N_A_2008_48#_c_1446_n N_A_2008_48#_M1003_g
+ N_A_2008_48#_c_1439_n N_A_2008_48#_c_1448_n N_A_2008_48#_c_1449_n
+ N_A_2008_48#_c_1450_n N_A_2008_48#_c_1451_n N_A_2008_48#_c_1440_n
+ N_A_2008_48#_c_1452_n N_A_2008_48#_c_1441_n N_A_2008_48#_c_1442_n
+ N_A_2008_48#_c_1454_n N_A_2008_48#_c_1443_n
+ PM_SKY130_FD_SC_HS__SDFRBP_1%A_2008_48#
x_PM_SKY130_FD_SC_HS__SDFRBP_1%A_1747_74# N_A_1747_74#_M1030_d
+ N_A_1747_74#_M1023_d N_A_1747_74#_c_1573_n N_A_1747_74#_M1010_g
+ N_A_1747_74#_c_1574_n N_A_1747_74#_c_1575_n N_A_1747_74#_c_1585_n
+ N_A_1747_74#_M1031_g N_A_1747_74#_c_1586_n N_A_1747_74#_c_1587_n
+ N_A_1747_74#_M1006_g N_A_1747_74#_c_1576_n N_A_1747_74#_M1008_g
+ N_A_1747_74#_c_1577_n N_A_1747_74#_c_1578_n N_A_1747_74#_c_1590_n
+ N_A_1747_74#_c_1591_n N_A_1747_74#_M1022_g N_A_1747_74#_M1002_g
+ N_A_1747_74#_c_1592_n N_A_1747_74#_c_1580_n N_A_1747_74#_c_1609_n
+ N_A_1747_74#_c_1627_n N_A_1747_74#_c_1594_n N_A_1747_74#_c_1595_n
+ N_A_1747_74#_c_1581_n N_A_1747_74#_c_1582_n N_A_1747_74#_c_1583_n
+ N_A_1747_74#_c_1584_n PM_SKY130_FD_SC_HS__SDFRBP_1%A_1747_74#
x_PM_SKY130_FD_SC_HS__SDFRBP_1%A_2513_424# N_A_2513_424#_M1002_s
+ N_A_2513_424#_M1022_s N_A_2513_424#_M1039_g N_A_2513_424#_c_1754_n
+ N_A_2513_424#_M1029_g N_A_2513_424#_c_1755_n N_A_2513_424#_c_1759_n
+ N_A_2513_424#_c_1756_n N_A_2513_424#_c_1757_n
+ PM_SKY130_FD_SC_HS__SDFRBP_1%A_2513_424#
x_PM_SKY130_FD_SC_HS__SDFRBP_1%VPWR N_VPWR_M1027_d N_VPWR_M1032_d N_VPWR_M1025_d
+ N_VPWR_M1018_d N_VPWR_M1019_s N_VPWR_M1003_d N_VPWR_M1031_d N_VPWR_M1022_d
+ N_VPWR_c_1804_n N_VPWR_c_1805_n N_VPWR_c_1806_n N_VPWR_c_1807_n
+ N_VPWR_c_1808_n N_VPWR_c_1809_n N_VPWR_c_1810_n N_VPWR_c_1923_n
+ N_VPWR_c_1811_n N_VPWR_c_1812_n N_VPWR_c_1813_n N_VPWR_c_1814_n
+ N_VPWR_c_1815_n N_VPWR_c_1816_n N_VPWR_c_1817_n N_VPWR_c_1818_n VPWR
+ N_VPWR_c_1819_n N_VPWR_c_1820_n N_VPWR_c_1821_n N_VPWR_c_1822_n
+ N_VPWR_c_1823_n N_VPWR_c_1824_n N_VPWR_c_1803_n N_VPWR_c_1826_n
+ N_VPWR_c_1827_n N_VPWR_c_1828_n N_VPWR_c_1829_n N_VPWR_c_1830_n
+ PM_SKY130_FD_SC_HS__SDFRBP_1%VPWR
x_PM_SKY130_FD_SC_HS__SDFRBP_1%A_413_90# N_A_413_90#_M1000_d N_A_413_90#_M1012_s
+ N_A_413_90#_M1009_d N_A_413_90#_M1020_d N_A_413_90#_M1028_s
+ N_A_413_90#_c_1985_n N_A_413_90#_c_1986_n N_A_413_90#_c_1994_n
+ N_A_413_90#_c_1995_n N_A_413_90#_c_1987_n N_A_413_90#_c_1996_n
+ N_A_413_90#_c_1988_n N_A_413_90#_c_1989_n N_A_413_90#_c_1990_n
+ N_A_413_90#_c_1998_n N_A_413_90#_c_1991_n N_A_413_90#_c_2004_n
+ N_A_413_90#_c_1999_n N_A_413_90#_c_1992_n N_A_413_90#_c_2000_n
+ PM_SKY130_FD_SC_HS__SDFRBP_1%A_413_90#
x_PM_SKY130_FD_SC_HS__SDFRBP_1%Q_N N_Q_N_M1008_d N_Q_N_M1006_d Q_N Q_N Q_N Q_N
+ Q_N Q_N Q_N PM_SKY130_FD_SC_HS__SDFRBP_1%Q_N
x_PM_SKY130_FD_SC_HS__SDFRBP_1%Q N_Q_M1039_d N_Q_M1029_d Q Q Q Q Q Q Q
+ N_Q_c_2156_n PM_SKY130_FD_SC_HS__SDFRBP_1%Q
x_PM_SKY130_FD_SC_HS__SDFRBP_1%VGND N_VGND_M1040_d N_VGND_M1034_d N_VGND_M1035_d
+ N_VGND_M1017_d N_VGND_M1005_d N_VGND_M1008_s N_VGND_M1002_d N_VGND_c_2174_n
+ N_VGND_c_2175_n N_VGND_c_2176_n N_VGND_c_2177_n N_VGND_c_2178_n
+ N_VGND_c_2179_n N_VGND_c_2180_n N_VGND_c_2181_n N_VGND_c_2182_n
+ N_VGND_c_2183_n N_VGND_c_2184_n VGND N_VGND_c_2185_n N_VGND_c_2186_n
+ N_VGND_c_2187_n N_VGND_c_2188_n N_VGND_c_2189_n N_VGND_c_2190_n
+ N_VGND_c_2191_n N_VGND_c_2192_n N_VGND_c_2193_n N_VGND_c_2194_n
+ N_VGND_c_2195_n PM_SKY130_FD_SC_HS__SDFRBP_1%VGND
x_PM_SKY130_FD_SC_HS__SDFRBP_1%noxref_25 N_noxref_25_M1021_s N_noxref_25_M1015_d
+ N_noxref_25_c_2313_n N_noxref_25_c_2314_n N_noxref_25_c_2315_n
+ N_noxref_25_c_2316_n PM_SKY130_FD_SC_HS__SDFRBP_1%noxref_25
cc_1 VNB N_A_27_74#_c_288_n 0.0213036f $X=-0.19 $Y=-0.245 $X2=1.485 $Y2=0.98
cc_2 VNB N_A_27_74#_c_289_n 0.0280153f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=0.58
cc_3 VNB N_A_27_74#_c_290_n 0.0167958f $X=-0.19 $Y=-0.245 $X2=0.2 $Y2=2.05
cc_4 VNB N_A_27_74#_c_291_n 0.0201543f $X=-0.19 $Y=-0.245 $X2=1.23 $Y2=1.145
cc_5 VNB N_A_27_74#_c_292_n 0.0460387f $X=-0.19 $Y=-0.245 $X2=1.23 $Y2=1.145
cc_6 VNB N_A_27_74#_c_293_n 0.018224f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.145
cc_7 VNB N_SCE_M1040_g 0.0718805f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_SCE_M1033_g 0.0299239f $X=-0.19 $Y=-0.245 $X2=0.2 $Y2=1.31
cc_9 VNB N_SCE_c_370_n 0.00457743f $X=-0.19 $Y=-0.245 $X2=0.365 $Y2=1.145
cc_10 VNB N_SCE_c_371_n 0.012877f $X=-0.19 $Y=-0.245 $X2=1.23 $Y2=1.145
cc_11 VNB N_SCE_c_372_n 0.00226615f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_SCE_c_373_n 0.0323948f $X=-0.19 $Y=-0.245 $X2=2.365 $Y2=2.135
cc_13 VNB N_SCE_c_374_n 0.0181262f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_SCE_c_375_n 0.0212614f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_SCE_c_376_n 0.00943038f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_SCE_c_377_n 0.001771f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_D_c_457_n 0.0248832f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_D_c_458_n 0.0352988f $X=-0.19 $Y=-0.245 $X2=2.485 $Y2=2.64
cc_19 VNB N_D_c_459_n 0.0056581f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=0.98
cc_20 VNB N_D_c_460_n 0.0173597f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=0.58
cc_21 VNB N_SCD_M1015_g 0.0388904f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_SCD_c_502_n 0.00416515f $X=-0.19 $Y=-0.245 $X2=2.485 $Y2=2.245
cc_23 VNB SCD 0.00223563f $X=-0.19 $Y=-0.245 $X2=2.485 $Y2=2.64
cc_24 VNB N_SCD_c_504_n 0.0166407f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_RESET_B_M1034_g 0.0627625f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_RESET_B_M1017_g 0.0217161f $X=-0.19 $Y=-0.245 $X2=2.485 $Y2=2.245
cc_27 VNB N_RESET_B_c_547_n 0.0213998f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_RESET_B_M1007_g 0.0341606f $X=-0.19 $Y=-0.245 $X2=0.365 $Y2=1.145
cc_29 VNB N_RESET_B_c_549_n 0.0315124f $X=-0.19 $Y=-0.245 $X2=0.89 $Y2=2.465
cc_30 VNB N_RESET_B_c_550_n 0.0234009f $X=-0.19 $Y=-0.245 $X2=2.53 $Y2=2.135
cc_31 VNB N_RESET_B_c_551_n 0.0158526f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_CLK_c_765_n 0.0205826f $X=-0.19 $Y=-0.245 $X2=0.135 $Y2=0.37
cc_33 VNB N_CLK_c_766_n 0.0218565f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_CLK_c_767_n 0.0558522f $X=-0.19 $Y=-0.245 $X2=1.485 $Y2=0.66
cc_35 VNB N_CLK_c_768_n 0.0152334f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=0.98
cc_36 VNB N_A_1023_74#_c_813_n 0.00999582f $X=-0.19 $Y=-0.245 $X2=2.485 $Y2=2.64
cc_37 VNB N_A_1023_74#_M1004_g 0.0473872f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_1023_74#_c_815_n 0.0165132f $X=-0.19 $Y=-0.245 $X2=0.2 $Y2=2.05
cc_39 VNB N_A_1023_74#_c_816_n 0.0213887f $X=-0.19 $Y=-0.245 $X2=1.23 $Y2=1.145
cc_40 VNB N_A_1023_74#_c_817_n 0.007535f $X=-0.19 $Y=-0.245 $X2=1.23 $Y2=1.145
cc_41 VNB N_A_1023_74#_c_818_n 0.00602149f $X=-0.19 $Y=-0.245 $X2=0.89 $Y2=2.512
cc_42 VNB N_A_1023_74#_c_819_n 0.029262f $X=-0.19 $Y=-0.245 $X2=0.89 $Y2=2.465
cc_43 VNB N_A_1023_74#_c_820_n 0.00359674f $X=-0.19 $Y=-0.245 $X2=1.055
+ $Y2=2.512
cc_44 VNB N_A_1023_74#_c_821_n 0.00279565f $X=-0.19 $Y=-0.245 $X2=2.53 $Y2=1.995
cc_45 VNB N_A_1023_74#_c_822_n 4.16166e-19 $X=-0.19 $Y=-0.245 $X2=2.53 $Y2=1.995
cc_46 VNB N_A_1023_74#_c_823_n 0.00204418f $X=-0.19 $Y=-0.245 $X2=2.53 $Y2=2.135
cc_47 VNB N_A_1023_74#_c_824_n 0.00104961f $X=-0.19 $Y=-0.245 $X2=2.53 $Y2=1.995
cc_48 VNB N_A_1023_74#_c_825_n 0.00867477f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A_1023_74#_c_826_n 0.00243212f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_A_1023_74#_c_827_n 0.00269633f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_A_1023_74#_c_828_n 0.00688208f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_A_1023_74#_c_829_n 0.00830295f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_A_1023_74#_c_830_n 0.0326227f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_A_1023_74#_c_831_n 0.00544115f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_A_1023_74#_c_832_n 0.0100685f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_A_1369_71#_M1016_g 0.0382884f $X=-0.19 $Y=-0.245 $X2=1.485 $Y2=0.66
cc_57 VNB N_A_1369_71#_c_1023_n 0.00474911f $X=-0.19 $Y=-0.245 $X2=0.2 $Y2=2.05
cc_58 VNB N_A_1369_71#_c_1024_n 0.0257402f $X=-0.19 $Y=-0.245 $X2=0.365
+ $Y2=1.145
cc_59 VNB N_A_1369_71#_c_1025_n 0.00892994f $X=-0.19 $Y=-0.245 $X2=1.23
+ $Y2=1.145
cc_60 VNB N_A_1369_71#_c_1026_n 0.00332197f $X=-0.19 $Y=-0.245 $X2=1.23
+ $Y2=1.145
cc_61 VNB N_A_1369_71#_c_1027_n 0.00177944f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_A_1369_71#_c_1028_n 0.00845443f $X=-0.19 $Y=-0.245 $X2=0.89
+ $Y2=2.512
cc_63 VNB N_A_1369_71#_c_1029_n 0.00273128f $X=-0.19 $Y=-0.245 $X2=1.055
+ $Y2=2.512
cc_64 VNB N_A_1369_71#_c_1030_n 0.00145912f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_A_1221_97#_M1041_g 0.0262153f $X=-0.19 $Y=-0.245 $X2=2.485 $Y2=2.64
cc_66 VNB N_A_1221_97#_c_1131_n 0.00511822f $X=-0.19 $Y=-0.245 $X2=0.2 $Y2=1.31
cc_67 VNB N_A_1221_97#_c_1132_n 0.012253f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.145
cc_68 VNB N_A_1221_97#_c_1133_n 5.52581e-19 $X=-0.19 $Y=-0.245 $X2=0.89
+ $Y2=2.465
cc_69 VNB N_A_1221_97#_c_1134_n 0.00251373f $X=-0.19 $Y=-0.245 $X2=1.055
+ $Y2=2.512
cc_70 VNB N_A_1221_97#_c_1135_n 0.00399797f $X=-0.19 $Y=-0.245 $X2=2.53
+ $Y2=1.995
cc_71 VNB N_A_1221_97#_c_1136_n 0.0423512f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_A_850_74#_c_1245_n 0.0156779f $X=-0.19 $Y=-0.245 $X2=1.485 $Y2=0.98
cc_73 VNB N_A_850_74#_c_1246_n 0.0323814f $X=-0.19 $Y=-0.245 $X2=2.485 $Y2=2.245
cc_74 VNB N_A_850_74#_c_1247_n 0.0111162f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=0.98
cc_75 VNB N_A_850_74#_c_1248_n 0.0136262f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_A_850_74#_c_1249_n 0.0233578f $X=-0.19 $Y=-0.245 $X2=0.2 $Y2=1.31
cc_77 VNB N_A_850_74#_M1012_g 0.0303219f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_A_850_74#_c_1251_n 0.0216126f $X=-0.19 $Y=-0.245 $X2=1.23 $Y2=1.145
cc_79 VNB N_A_850_74#_c_1252_n 0.00443907f $X=-0.19 $Y=-0.245 $X2=1.485 $Y2=0.98
cc_80 VNB N_A_850_74#_M1013_g 0.0521391f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_81 VNB N_A_850_74#_c_1254_n 0.00756215f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_82 VNB N_A_850_74#_c_1255_n 0.0026699f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_83 VNB N_A_850_74#_c_1256_n 0.00733274f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_84 VNB N_A_850_74#_c_1257_n 0.00179234f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_85 VNB N_A_850_74#_c_1258_n 5.99108e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_86 VNB N_A_850_74#_c_1259_n 0.0031096f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_87 VNB N_A_2008_48#_M1005_g 0.0424527f $X=-0.19 $Y=-0.245 $X2=1.485 $Y2=0.66
cc_88 VNB N_A_2008_48#_c_1438_n 0.0184816f $X=-0.19 $Y=-0.245 $X2=2.485 $Y2=2.64
cc_89 VNB N_A_2008_48#_c_1439_n 0.00245359f $X=-0.19 $Y=-0.245 $X2=0.2 $Y2=2.05
cc_90 VNB N_A_2008_48#_c_1440_n 0.00907094f $X=-0.19 $Y=-0.245 $X2=0.89
+ $Y2=2.512
cc_91 VNB N_A_2008_48#_c_1441_n 6.5078e-19 $X=-0.19 $Y=-0.245 $X2=2.53 $Y2=1.995
cc_92 VNB N_A_2008_48#_c_1442_n 0.00160142f $X=-0.19 $Y=-0.245 $X2=2.53
+ $Y2=1.995
cc_93 VNB N_A_2008_48#_c_1443_n 0.00658078f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_94 VNB N_A_1747_74#_c_1573_n 0.0180751f $X=-0.19 $Y=-0.245 $X2=1.485 $Y2=0.98
cc_95 VNB N_A_1747_74#_c_1574_n 0.031848f $X=-0.19 $Y=-0.245 $X2=2.485 $Y2=2.245
cc_96 VNB N_A_1747_74#_c_1575_n 0.0157622f $X=-0.19 $Y=-0.245 $X2=2.485 $Y2=2.64
cc_97 VNB N_A_1747_74#_c_1576_n 0.0240396f $X=-0.19 $Y=-0.245 $X2=1.23 $Y2=1.145
cc_98 VNB N_A_1747_74#_c_1577_n 0.0485723f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_99 VNB N_A_1747_74#_c_1578_n 0.0663668f $X=-0.19 $Y=-0.245 $X2=2.365
+ $Y2=2.135
cc_100 VNB N_A_1747_74#_M1002_g 0.0405544f $X=-0.19 $Y=-0.245 $X2=2.53 $Y2=1.995
cc_101 VNB N_A_1747_74#_c_1580_n 0.00927852f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_102 VNB N_A_1747_74#_c_1581_n 0.00249714f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_103 VNB N_A_1747_74#_c_1582_n 0.00130137f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_104 VNB N_A_1747_74#_c_1583_n 0.0147798f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_105 VNB N_A_1747_74#_c_1584_n 0.020816f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_106 VNB N_A_2513_424#_M1039_g 0.0280908f $X=-0.19 $Y=-0.245 $X2=1.485
+ $Y2=0.66
cc_107 VNB N_A_2513_424#_c_1754_n 0.0352088f $X=-0.19 $Y=-0.245 $X2=2.485
+ $Y2=2.64
cc_108 VNB N_A_2513_424#_c_1755_n 0.0126466f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_109 VNB N_A_2513_424#_c_1756_n 0.00835153f $X=-0.19 $Y=-0.245 $X2=2.365
+ $Y2=2.135
cc_110 VNB N_A_2513_424#_c_1757_n 4.48326e-19 $X=-0.19 $Y=-0.245 $X2=0.2
+ $Y2=2.512
cc_111 VNB N_VPWR_c_1803_n 0.581632f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_112 VNB N_A_413_90#_c_1985_n 0.0226398f $X=-0.19 $Y=-0.245 $X2=1.23 $Y2=1.145
cc_113 VNB N_A_413_90#_c_1986_n 0.00517566f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_114 VNB N_A_413_90#_c_1987_n 0.00165194f $X=-0.19 $Y=-0.245 $X2=0.89
+ $Y2=2.512
cc_115 VNB N_A_413_90#_c_1988_n 0.0058676f $X=-0.19 $Y=-0.245 $X2=2.53 $Y2=1.995
cc_116 VNB N_A_413_90#_c_1989_n 7.33295e-19 $X=-0.19 $Y=-0.245 $X2=2.53
+ $Y2=1.995
cc_117 VNB N_A_413_90#_c_1990_n 0.00598059f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_118 VNB N_A_413_90#_c_1991_n 0.00483383f $X=-0.19 $Y=-0.245 $X2=1.485
+ $Y2=0.98
cc_119 VNB N_A_413_90#_c_1992_n 0.00211107f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_120 VNB Q_N 0.0123064f $X=-0.19 $Y=-0.245 $X2=1.485 $Y2=0.98
cc_121 VNB Q 0.0267037f $X=-0.19 $Y=-0.245 $X2=1.485 $Y2=0.66
cc_122 VNB Q 0.0127641f $X=-0.19 $Y=-0.245 $X2=2.485 $Y2=2.245
cc_123 VNB N_Q_c_2156_n 0.0251085f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_124 VNB N_VGND_c_2174_n 0.0135998f $X=-0.19 $Y=-0.245 $X2=2.365 $Y2=2.135
cc_125 VNB N_VGND_c_2175_n 0.014263f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_126 VNB N_VGND_c_2176_n 0.00340259f $X=-0.19 $Y=-0.245 $X2=2.53 $Y2=1.995
cc_127 VNB N_VGND_c_2177_n 0.00865424f $X=-0.19 $Y=-0.245 $X2=2.53 $Y2=2.135
cc_128 VNB N_VGND_c_2178_n 0.00396467f $X=-0.19 $Y=-0.245 $X2=2.53 $Y2=1.995
cc_129 VNB N_VGND_c_2179_n 0.0363017f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_130 VNB N_VGND_c_2180_n 0.0097163f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_131 VNB N_VGND_c_2181_n 0.0663868f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_132 VNB N_VGND_c_2182_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_133 VNB N_VGND_c_2183_n 0.0188435f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_134 VNB N_VGND_c_2184_n 0.00604233f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_135 VNB N_VGND_c_2185_n 0.0173909f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_136 VNB N_VGND_c_2186_n 0.0575933f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_137 VNB N_VGND_c_2187_n 0.0609299f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_138 VNB N_VGND_c_2188_n 0.0284194f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_139 VNB N_VGND_c_2189_n 0.0193554f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_140 VNB N_VGND_c_2190_n 0.765774f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_141 VNB N_VGND_c_2191_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_142 VNB N_VGND_c_2192_n 0.00631189f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_143 VNB N_VGND_c_2193_n 0.00604233f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_144 VNB N_VGND_c_2194_n 0.0153005f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_145 VNB N_VGND_c_2195_n 0.00326991f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_146 VNB N_noxref_25_c_2313_n 0.00380385f $X=-0.19 $Y=-0.245 $X2=1.485
+ $Y2=0.66
cc_147 VNB N_noxref_25_c_2314_n 0.0318599f $X=-0.19 $Y=-0.245 $X2=2.485 $Y2=2.64
cc_148 VNB N_noxref_25_c_2315_n 0.00398497f $X=-0.19 $Y=-0.245 $X2=2.485
+ $Y2=2.64
cc_149 VNB N_noxref_25_c_2316_n 0.00603433f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=0.98
cc_150 VPB N_A_27_74#_c_294_n 0.0531412f $X=-0.19 $Y=1.66 $X2=2.485 $Y2=2.245
cc_151 VPB N_A_27_74#_c_290_n 0.0237442f $X=-0.19 $Y=1.66 $X2=0.2 $Y2=2.05
cc_152 VPB N_A_27_74#_c_296_n 0.022353f $X=-0.19 $Y=1.66 $X2=2.365 $Y2=2.135
cc_153 VPB N_A_27_74#_c_297_n 0.064305f $X=-0.19 $Y=1.66 $X2=1.055 $Y2=2.512
cc_154 VPB N_A_27_74#_c_298_n 0.00429588f $X=-0.19 $Y=1.66 $X2=2.53 $Y2=1.995
cc_155 VPB N_SCE_c_378_n 0.021095f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_156 VPB N_SCE_c_379_n 0.0272472f $X=-0.19 $Y=1.66 $X2=1.485 $Y2=0.98
cc_157 VPB N_SCE_c_380_n 0.0141937f $X=-0.19 $Y=1.66 $X2=2.485 $Y2=2.64
cc_158 VPB N_SCE_c_381_n 0.0211524f $X=-0.19 $Y=1.66 $X2=2.485 $Y2=2.64
cc_159 VPB N_SCE_c_370_n 0.0130807f $X=-0.19 $Y=1.66 $X2=0.365 $Y2=1.145
cc_160 VPB N_SCE_c_372_n 0.00295534f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_161 VPB N_SCE_c_374_n 0.0215244f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_162 VPB N_SCE_c_375_n 0.0217946f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_163 VPB N_SCE_c_377_n 0.00321268f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_164 VPB N_D_c_457_n 0.0307331f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_165 VPB N_D_c_462_n 0.0213891f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_166 VPB N_SCD_c_505_n 0.0170207f $X=-0.19 $Y=1.66 $X2=0.135 $Y2=0.37
cc_167 VPB N_SCD_c_502_n 0.0505553f $X=-0.19 $Y=1.66 $X2=2.485 $Y2=2.245
cc_168 VPB SCD 0.00183951f $X=-0.19 $Y=1.66 $X2=2.485 $Y2=2.64
cc_169 VPB N_RESET_B_M1034_g 0.0115735f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_170 VPB N_RESET_B_c_553_n 0.0213877f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_171 VPB N_RESET_B_c_554_n 0.0386858f $X=-0.19 $Y=1.66 $X2=2.485 $Y2=2.64
cc_172 VPB N_RESET_B_c_547_n 0.0119976f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_173 VPB N_RESET_B_c_556_n 0.0117494f $X=-0.19 $Y=1.66 $X2=1.23 $Y2=1.145
cc_174 VPB N_RESET_B_c_557_n 0.0274905f $X=-0.19 $Y=1.66 $X2=1.485 $Y2=0.98
cc_175 VPB N_RESET_B_c_558_n 0.0206649f $X=-0.19 $Y=1.66 $X2=2.53 $Y2=1.995
cc_176 VPB N_RESET_B_c_559_n 0.00331698f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_177 VPB N_RESET_B_c_560_n 0.0138334f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_178 VPB N_RESET_B_c_561_n 0.00662848f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_179 VPB RESET_B 0.00207862f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_180 VPB N_RESET_B_c_563_n 0.0371391f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_181 VPB N_RESET_B_c_564_n 0.00183211f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_182 VPB N_RESET_B_c_565_n 0.0709137f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_183 VPB N_RESET_B_c_566_n 0.00202094f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_184 VPB N_RESET_B_c_567_n 0.0307002f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_185 VPB N_RESET_B_c_568_n 0.0048181f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_186 VPB N_RESET_B_c_551_n 0.00104493f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_187 VPB N_CLK_c_766_n 0.0282017f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_188 VPB N_A_1023_74#_c_833_n 0.0149784f $X=-0.19 $Y=1.66 $X2=1.485 $Y2=0.66
cc_189 VPB N_A_1023_74#_c_834_n 0.019571f $X=-0.19 $Y=1.66 $X2=1.485 $Y2=0.66
cc_190 VPB N_A_1023_74#_c_813_n 0.0151986f $X=-0.19 $Y=1.66 $X2=2.485 $Y2=2.64
cc_191 VPB N_A_1023_74#_c_836_n 0.0616091f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_192 VPB N_A_1023_74#_c_822_n 0.00517344f $X=-0.19 $Y=1.66 $X2=2.53 $Y2=1.995
cc_193 VPB N_A_1023_74#_c_823_n 0.00184525f $X=-0.19 $Y=1.66 $X2=2.53 $Y2=2.135
cc_194 VPB N_A_1023_74#_c_839_n 0.00535343f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_195 VPB N_A_1023_74#_c_832_n 0.0208444f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_196 VPB N_A_1369_71#_c_1031_n 0.0269225f $X=-0.19 $Y=1.66 $X2=2.485 $Y2=2.64
cc_197 VPB N_A_1369_71#_c_1032_n 0.0207894f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=0.98
cc_198 VPB N_A_1369_71#_c_1023_n 0.00226924f $X=-0.19 $Y=1.66 $X2=0.2 $Y2=2.05
cc_199 VPB N_A_1369_71#_c_1024_n 0.0182294f $X=-0.19 $Y=1.66 $X2=0.365 $Y2=1.145
cc_200 VPB N_A_1369_71#_c_1029_n 0.00432622f $X=-0.19 $Y=1.66 $X2=1.055
+ $Y2=2.512
cc_201 VPB N_A_1221_97#_c_1137_n 0.0164664f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=0.58
cc_202 VPB N_A_1221_97#_c_1138_n 0.00309276f $X=-0.19 $Y=1.66 $X2=1.23 $Y2=1.145
cc_203 VPB N_A_1221_97#_c_1132_n 0.0122061f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=1.145
cc_204 VPB N_A_1221_97#_c_1133_n 0.0127694f $X=-0.19 $Y=1.66 $X2=0.89 $Y2=2.465
cc_205 VPB N_A_1221_97#_c_1141_n 0.00178603f $X=-0.19 $Y=1.66 $X2=2.53 $Y2=2.135
cc_206 VPB N_A_1221_97#_c_1136_n 0.023248f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_207 VPB N_A_850_74#_c_1246_n 0.0214835f $X=-0.19 $Y=1.66 $X2=2.485 $Y2=2.245
cc_208 VPB N_A_850_74#_c_1248_n 0.0767109f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_209 VPB N_A_850_74#_c_1262_n 0.0548537f $X=-0.19 $Y=1.66 $X2=0.365 $Y2=1.145
cc_210 VPB N_A_850_74#_c_1263_n 0.0125836f $X=-0.19 $Y=1.66 $X2=1.23 $Y2=1.145
cc_211 VPB N_A_850_74#_c_1264_n 0.00707451f $X=-0.19 $Y=1.66 $X2=1.055 $Y2=2.135
cc_212 VPB N_A_850_74#_c_1265_n 0.0163525f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=1.145
cc_213 VPB N_A_850_74#_c_1266_n 0.0144828f $X=-0.19 $Y=1.66 $X2=0.2 $Y2=2.512
cc_214 VPB N_A_850_74#_c_1267_n 0.181289f $X=-0.19 $Y=1.66 $X2=0.89 $Y2=2.465
cc_215 VPB N_A_850_74#_c_1268_n 0.00753678f $X=-0.19 $Y=1.66 $X2=2.53 $Y2=1.995
cc_216 VPB N_A_850_74#_c_1269_n 0.0145726f $X=-0.19 $Y=1.66 $X2=2.53 $Y2=1.995
cc_217 VPB N_A_850_74#_M1023_g 0.00889026f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_218 VPB N_A_850_74#_c_1251_n 0.0212414f $X=-0.19 $Y=1.66 $X2=1.23 $Y2=1.145
cc_219 VPB N_A_850_74#_c_1252_n 0.00362133f $X=-0.19 $Y=1.66 $X2=1.485 $Y2=0.98
cc_220 VPB N_A_850_74#_c_1273_n 0.0089864f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_221 VPB N_A_850_74#_c_1274_n 0.00298529f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_222 VPB N_A_850_74#_c_1258_n 0.00276522f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_223 VPB N_A_850_74#_c_1276_n 0.00202514f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_224 VPB N_A_2008_48#_c_1438_n 0.0363084f $X=-0.19 $Y=1.66 $X2=2.485 $Y2=2.64
cc_225 VPB N_A_2008_48#_c_1445_n 0.0157644f $X=-0.19 $Y=1.66 $X2=2.485 $Y2=2.64
cc_226 VPB N_A_2008_48#_c_1446_n 0.0216925f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=0.98
cc_227 VPB N_A_2008_48#_c_1439_n 0.00554437f $X=-0.19 $Y=1.66 $X2=0.2 $Y2=2.05
cc_228 VPB N_A_2008_48#_c_1448_n 0.00200572f $X=-0.19 $Y=1.66 $X2=1.23 $Y2=1.145
cc_229 VPB N_A_2008_48#_c_1449_n 0.00188008f $X=-0.19 $Y=1.66 $X2=1.23 $Y2=1.145
cc_230 VPB N_A_2008_48#_c_1450_n 0.0030033f $X=-0.19 $Y=1.66 $X2=1.055 $Y2=2.135
cc_231 VPB N_A_2008_48#_c_1451_n 0.00272239f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_232 VPB N_A_2008_48#_c_1452_n 0.00910875f $X=-0.19 $Y=1.66 $X2=1.055
+ $Y2=2.512
cc_233 VPB N_A_2008_48#_c_1441_n 0.00102188f $X=-0.19 $Y=1.66 $X2=2.53 $Y2=1.995
cc_234 VPB N_A_2008_48#_c_1454_n 0.00510966f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_235 VPB N_A_1747_74#_c_1585_n 0.0156363f $X=-0.19 $Y=1.66 $X2=2.485 $Y2=2.64
cc_236 VPB N_A_1747_74#_c_1586_n 0.0266893f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_237 VPB N_A_1747_74#_c_1587_n 0.0200685f $X=-0.19 $Y=1.66 $X2=0.2 $Y2=1.31
cc_238 VPB N_A_1747_74#_c_1577_n 0.0295508f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_239 VPB N_A_1747_74#_c_1578_n 0.0208636f $X=-0.19 $Y=1.66 $X2=2.365 $Y2=2.135
cc_240 VPB N_A_1747_74#_c_1590_n 0.0185739f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=1.145
cc_241 VPB N_A_1747_74#_c_1591_n 0.0280061f $X=-0.19 $Y=1.66 $X2=0.2 $Y2=2.512
cc_242 VPB N_A_1747_74#_c_1592_n 0.0189178f $X=-0.19 $Y=1.66 $X2=2.53 $Y2=1.995
cc_243 VPB N_A_1747_74#_c_1580_n 0.00103641f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_244 VPB N_A_1747_74#_c_1594_n 0.00533426f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_245 VPB N_A_1747_74#_c_1595_n 0.00295698f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_246 VPB N_A_1747_74#_c_1582_n 0.00536747f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_247 VPB N_A_2513_424#_c_1754_n 0.0293072f $X=-0.19 $Y=1.66 $X2=2.485 $Y2=2.64
cc_248 VPB N_A_2513_424#_c_1759_n 0.00679439f $X=-0.19 $Y=1.66 $X2=1.23
+ $Y2=1.145
cc_249 VPB N_VPWR_c_1804_n 0.00653637f $X=-0.19 $Y=1.66 $X2=0.2 $Y2=2.512
cc_250 VPB N_VPWR_c_1805_n 0.00677641f $X=-0.19 $Y=1.66 $X2=1.055 $Y2=2.512
cc_251 VPB N_VPWR_c_1806_n 0.00486025f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_252 VPB N_VPWR_c_1807_n 0.0138299f $X=-0.19 $Y=1.66 $X2=1.485 $Y2=0.98
cc_253 VPB N_VPWR_c_1808_n 0.015124f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_254 VPB N_VPWR_c_1809_n 0.0169757f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_255 VPB N_VPWR_c_1810_n 0.0142672f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_256 VPB N_VPWR_c_1811_n 0.0141486f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_257 VPB N_VPWR_c_1812_n 0.0338628f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_258 VPB N_VPWR_c_1813_n 0.00614127f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_259 VPB N_VPWR_c_1814_n 0.0370161f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_260 VPB N_VPWR_c_1815_n 0.00626055f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_261 VPB N_VPWR_c_1816_n 0.0596332f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_262 VPB N_VPWR_c_1817_n 0.00436868f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_263 VPB N_VPWR_c_1818_n 5.16032e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_264 VPB N_VPWR_c_1819_n 0.0456433f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_265 VPB N_VPWR_c_1820_n 0.0221228f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_266 VPB N_VPWR_c_1821_n 0.0505955f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_267 VPB N_VPWR_c_1822_n 0.020722f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_268 VPB N_VPWR_c_1823_n 0.0343043f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_269 VPB N_VPWR_c_1824_n 0.0189057f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_270 VPB N_VPWR_c_1803_n 0.140667f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_271 VPB N_VPWR_c_1826_n 0.00671858f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_272 VPB N_VPWR_c_1827_n 0.00330333f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_273 VPB N_VPWR_c_1828_n 0.0066101f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_274 VPB N_VPWR_c_1829_n 0.00853483f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_275 VPB N_VPWR_c_1830_n 0.00535984f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_276 VPB N_A_413_90#_c_1986_n 0.00490368f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_277 VPB N_A_413_90#_c_1994_n 0.00979095f $X=-0.19 $Y=1.66 $X2=2.365 $Y2=2.135
cc_278 VPB N_A_413_90#_c_1995_n 0.0120995f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=1.145
cc_279 VPB N_A_413_90#_c_1996_n 0.007415f $X=-0.19 $Y=1.66 $X2=0.89 $Y2=2.465
cc_280 VPB N_A_413_90#_c_1990_n 0.00541415f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_281 VPB N_A_413_90#_c_1998_n 0.00248229f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_282 VPB N_A_413_90#_c_1999_n 0.00142001f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_283 VPB N_A_413_90#_c_2000_n 0.00949635f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_284 VPB Q_N 0.0164214f $X=-0.19 $Y=1.66 $X2=1.485 $Y2=0.98
cc_285 VPB Q 0.0100975f $X=-0.19 $Y=1.66 $X2=2.485 $Y2=2.64
cc_286 VPB Q 0.0417421f $X=-0.19 $Y=1.66 $X2=2.53 $Y2=1.995
cc_287 VPB N_Q_c_2156_n 0.00779891f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_288 N_A_27_74#_c_289_n N_SCE_M1040_g 0.00834942f $X=0.28 $Y=0.58 $X2=0 $Y2=0
cc_289 N_A_27_74#_c_290_n N_SCE_M1040_g 0.017345f $X=0.2 $Y=2.05 $X2=0 $Y2=0
cc_290 N_A_27_74#_c_291_n N_SCE_M1040_g 0.0301676f $X=1.23 $Y=1.145 $X2=0 $Y2=0
cc_291 N_A_27_74#_c_292_n N_SCE_M1040_g 0.00651386f $X=1.23 $Y=1.145 $X2=0 $Y2=0
cc_292 N_A_27_74#_c_296_n N_SCE_c_378_n 0.00485819f $X=2.365 $Y=2.135 $X2=0
+ $Y2=0
cc_293 N_A_27_74#_c_297_n N_SCE_c_378_n 0.00322075f $X=1.055 $Y=2.512 $X2=0
+ $Y2=0
cc_294 N_A_27_74#_c_296_n N_SCE_c_379_n 0.00822995f $X=2.365 $Y=2.135 $X2=0
+ $Y2=0
cc_295 N_A_27_74#_c_297_n N_SCE_c_379_n 0.014007f $X=1.055 $Y=2.512 $X2=0 $Y2=0
cc_296 N_A_27_74#_c_296_n N_SCE_c_380_n 0.00663467f $X=2.365 $Y=2.135 $X2=0
+ $Y2=0
cc_297 N_A_27_74#_c_296_n N_SCE_c_381_n 0.00943326f $X=2.365 $Y=2.135 $X2=0
+ $Y2=0
cc_298 N_A_27_74#_c_297_n N_SCE_c_381_n 7.55381e-19 $X=1.055 $Y=2.512 $X2=0
+ $Y2=0
cc_299 N_A_27_74#_c_297_n N_SCE_c_370_n 0.0185427f $X=1.055 $Y=2.512 $X2=0 $Y2=0
cc_300 N_A_27_74#_c_294_n N_SCE_c_371_n 2.04435e-19 $X=2.485 $Y=2.245 $X2=0
+ $Y2=0
cc_301 N_A_27_74#_c_296_n N_SCE_c_371_n 0.0227799f $X=2.365 $Y=2.135 $X2=0 $Y2=0
cc_302 N_A_27_74#_c_298_n N_SCE_c_371_n 0.00221846f $X=2.53 $Y=1.995 $X2=0 $Y2=0
cc_303 N_A_27_74#_c_294_n N_SCE_c_372_n 0.00103776f $X=2.485 $Y=2.245 $X2=0
+ $Y2=0
cc_304 N_A_27_74#_c_298_n N_SCE_c_372_n 0.0244747f $X=2.53 $Y=1.995 $X2=0 $Y2=0
cc_305 N_A_27_74#_c_294_n N_SCE_c_373_n 0.0165737f $X=2.485 $Y=2.245 $X2=0 $Y2=0
cc_306 N_A_27_74#_c_298_n N_SCE_c_373_n 3.27431e-19 $X=2.53 $Y=1.995 $X2=0 $Y2=0
cc_307 N_A_27_74#_c_291_n N_SCE_c_374_n 0.00418014f $X=1.23 $Y=1.145 $X2=0 $Y2=0
cc_308 N_A_27_74#_c_291_n N_SCE_c_375_n 3.70862e-19 $X=1.23 $Y=1.145 $X2=0 $Y2=0
cc_309 N_A_27_74#_c_292_n N_SCE_c_375_n 0.0219042f $X=1.23 $Y=1.145 $X2=0 $Y2=0
cc_310 N_A_27_74#_c_296_n N_SCE_c_375_n 0.00313888f $X=2.365 $Y=2.135 $X2=0
+ $Y2=0
cc_311 N_A_27_74#_c_290_n N_SCE_c_376_n 0.0195247f $X=0.2 $Y=2.05 $X2=0 $Y2=0
cc_312 N_A_27_74#_c_291_n N_SCE_c_376_n 0.0626128f $X=1.23 $Y=1.145 $X2=0 $Y2=0
cc_313 N_A_27_74#_c_292_n N_SCE_c_376_n 0.00563186f $X=1.23 $Y=1.145 $X2=0 $Y2=0
cc_314 N_A_27_74#_c_297_n N_SCE_c_376_n 0.0467278f $X=1.055 $Y=2.512 $X2=0 $Y2=0
cc_315 N_A_27_74#_c_296_n N_SCE_c_377_n 0.0467278f $X=2.365 $Y=2.135 $X2=0 $Y2=0
cc_316 N_A_27_74#_c_298_n N_SCE_c_377_n 0.00165158f $X=2.53 $Y=1.995 $X2=0 $Y2=0
cc_317 N_A_27_74#_c_294_n N_D_c_457_n 0.0182683f $X=2.485 $Y=2.245 $X2=0 $Y2=0
cc_318 N_A_27_74#_c_296_n N_D_c_457_n 0.00773295f $X=2.365 $Y=2.135 $X2=0 $Y2=0
cc_319 N_A_27_74#_c_298_n N_D_c_457_n 0.00139926f $X=2.53 $Y=1.995 $X2=0 $Y2=0
cc_320 N_A_27_74#_c_294_n N_D_c_462_n 0.0136568f $X=2.485 $Y=2.245 $X2=0 $Y2=0
cc_321 N_A_27_74#_c_296_n N_D_c_462_n 0.00913859f $X=2.365 $Y=2.135 $X2=0 $Y2=0
cc_322 N_A_27_74#_c_291_n N_D_c_458_n 2.658e-19 $X=1.23 $Y=1.145 $X2=0 $Y2=0
cc_323 N_A_27_74#_c_292_n N_D_c_458_n 0.0150607f $X=1.23 $Y=1.145 $X2=0 $Y2=0
cc_324 N_A_27_74#_c_288_n N_D_c_459_n 0.00525376f $X=1.485 $Y=0.98 $X2=0 $Y2=0
cc_325 N_A_27_74#_c_291_n N_D_c_459_n 0.0286966f $X=1.23 $Y=1.145 $X2=0 $Y2=0
cc_326 N_A_27_74#_c_292_n N_D_c_459_n 7.30413e-19 $X=1.23 $Y=1.145 $X2=0 $Y2=0
cc_327 N_A_27_74#_c_288_n N_D_c_460_n 0.0223399f $X=1.485 $Y=0.98 $X2=0 $Y2=0
cc_328 N_A_27_74#_c_294_n N_SCD_c_505_n 0.0262181f $X=2.485 $Y=2.245 $X2=-0.19
+ $Y2=-0.245
cc_329 N_A_27_74#_c_294_n N_SCD_c_502_n 0.0198258f $X=2.485 $Y=2.245 $X2=0 $Y2=0
cc_330 N_A_27_74#_c_298_n N_SCD_c_502_n 0.00257757f $X=2.53 $Y=1.995 $X2=0 $Y2=0
cc_331 N_A_27_74#_c_294_n SCD 0.00117743f $X=2.485 $Y=2.245 $X2=0 $Y2=0
cc_332 N_A_27_74#_c_298_n SCD 0.0182021f $X=2.53 $Y=1.995 $X2=0 $Y2=0
cc_333 N_A_27_74#_c_296_n N_VPWR_c_1804_n 0.0234317f $X=2.365 $Y=2.135 $X2=0
+ $Y2=0
cc_334 N_A_27_74#_c_297_n N_VPWR_c_1804_n 0.0251436f $X=1.055 $Y=2.512 $X2=0
+ $Y2=0
cc_335 N_A_27_74#_c_294_n N_VPWR_c_1805_n 0.00124919f $X=2.485 $Y=2.245 $X2=0
+ $Y2=0
cc_336 N_A_27_74#_c_297_n N_VPWR_c_1812_n 0.0408917f $X=1.055 $Y=2.512 $X2=0
+ $Y2=0
cc_337 N_A_27_74#_c_294_n N_VPWR_c_1819_n 0.00445347f $X=2.485 $Y=2.245 $X2=0
+ $Y2=0
cc_338 N_A_27_74#_c_294_n N_VPWR_c_1803_n 0.0043847f $X=2.485 $Y=2.245 $X2=0
+ $Y2=0
cc_339 N_A_27_74#_c_297_n N_VPWR_c_1803_n 0.0345127f $X=1.055 $Y=2.512 $X2=0
+ $Y2=0
cc_340 N_A_27_74#_c_294_n N_A_413_90#_c_1998_n 0.00949185f $X=2.485 $Y=2.245
+ $X2=0 $Y2=0
cc_341 N_A_27_74#_c_296_n N_A_413_90#_c_1998_n 0.0188908f $X=2.365 $Y=2.135
+ $X2=0 $Y2=0
cc_342 N_A_27_74#_c_298_n N_A_413_90#_c_1998_n 0.00299996f $X=2.53 $Y=1.995
+ $X2=0 $Y2=0
cc_343 N_A_27_74#_c_294_n N_A_413_90#_c_2004_n 0.00998537f $X=2.485 $Y=2.245
+ $X2=0 $Y2=0
cc_344 N_A_27_74#_c_298_n N_A_413_90#_c_2004_n 0.018284f $X=2.53 $Y=1.995 $X2=0
+ $Y2=0
cc_345 N_A_27_74#_c_288_n N_VGND_c_2174_n 0.00108896f $X=1.485 $Y=0.98 $X2=0
+ $Y2=0
cc_346 N_A_27_74#_c_289_n N_VGND_c_2174_n 0.0179429f $X=0.28 $Y=0.58 $X2=0 $Y2=0
cc_347 N_A_27_74#_c_291_n N_VGND_c_2174_n 0.0288081f $X=1.23 $Y=1.145 $X2=0
+ $Y2=0
cc_348 N_A_27_74#_c_288_n N_VGND_c_2181_n 8.05596e-19 $X=1.485 $Y=0.98 $X2=0
+ $Y2=0
cc_349 N_A_27_74#_c_289_n N_VGND_c_2185_n 0.011066f $X=0.28 $Y=0.58 $X2=0 $Y2=0
cc_350 N_A_27_74#_c_289_n N_VGND_c_2190_n 0.00915947f $X=0.28 $Y=0.58 $X2=0
+ $Y2=0
cc_351 N_A_27_74#_c_288_n N_noxref_25_c_2313_n 9.72985e-19 $X=1.485 $Y=0.98
+ $X2=0 $Y2=0
cc_352 N_A_27_74#_c_291_n N_noxref_25_c_2313_n 0.0201381f $X=1.23 $Y=1.145 $X2=0
+ $Y2=0
cc_353 N_A_27_74#_c_292_n N_noxref_25_c_2313_n 0.00573089f $X=1.23 $Y=1.145
+ $X2=0 $Y2=0
cc_354 N_A_27_74#_c_288_n N_noxref_25_c_2314_n 0.0139744f $X=1.485 $Y=0.98 $X2=0
+ $Y2=0
cc_355 N_A_27_74#_c_291_n N_noxref_25_c_2314_n 0.00121356f $X=1.23 $Y=1.145
+ $X2=0 $Y2=0
cc_356 N_A_27_74#_c_292_n N_noxref_25_c_2314_n 0.00100866f $X=1.23 $Y=1.145
+ $X2=0 $Y2=0
cc_357 N_SCE_c_371_n N_D_c_457_n 0.0149823f $X=2.395 $Y=1.575 $X2=0 $Y2=0
cc_358 N_SCE_c_372_n N_D_c_457_n 3.21106e-19 $X=2.56 $Y=1.425 $X2=0 $Y2=0
cc_359 N_SCE_c_375_n N_D_c_457_n 0.0188435f $X=1.615 $Y=1.715 $X2=0 $Y2=0
cc_360 N_SCE_c_377_n N_D_c_457_n 0.00533998f $X=1.795 $Y=1.685 $X2=0 $Y2=0
cc_361 N_SCE_c_380_n N_D_c_462_n 0.0188435f $X=1.615 $Y=2.155 $X2=0 $Y2=0
cc_362 N_SCE_c_381_n N_D_c_462_n 0.0377129f $X=1.615 $Y=2.245 $X2=0 $Y2=0
cc_363 N_SCE_M1033_g N_D_c_458_n 0.00739628f $X=2.65 $Y=0.695 $X2=0 $Y2=0
cc_364 N_SCE_c_372_n N_D_c_458_n 0.00136148f $X=2.56 $Y=1.425 $X2=0 $Y2=0
cc_365 N_SCE_c_373_n N_D_c_458_n 0.0159923f $X=2.56 $Y=1.425 $X2=0 $Y2=0
cc_366 N_SCE_c_377_n N_D_c_458_n 0.00402499f $X=1.795 $Y=1.685 $X2=0 $Y2=0
cc_367 N_SCE_M1033_g N_D_c_459_n 0.00121036f $X=2.65 $Y=0.695 $X2=0 $Y2=0
cc_368 N_SCE_c_372_n N_D_c_459_n 0.00246473f $X=2.56 $Y=1.425 $X2=0 $Y2=0
cc_369 N_SCE_c_375_n N_D_c_459_n 9.21412e-19 $X=1.615 $Y=1.715 $X2=0 $Y2=0
cc_370 N_SCE_c_376_n N_D_c_459_n 0.0411265f $X=1.6 $Y=1.685 $X2=0 $Y2=0
cc_371 N_SCE_M1033_g N_D_c_460_n 0.0097239f $X=2.65 $Y=0.695 $X2=0 $Y2=0
cc_372 N_SCE_M1033_g N_SCD_M1015_g 0.0589665f $X=2.65 $Y=0.695 $X2=0 $Y2=0
cc_373 N_SCE_c_372_n N_SCD_M1015_g 0.00116379f $X=2.56 $Y=1.425 $X2=0 $Y2=0
cc_374 N_SCE_c_372_n SCD 0.0142044f $X=2.56 $Y=1.425 $X2=0 $Y2=0
cc_375 N_SCE_c_373_n SCD 5.22436e-19 $X=2.56 $Y=1.425 $X2=0 $Y2=0
cc_376 N_SCE_c_372_n N_SCD_c_504_n 0.00206001f $X=2.56 $Y=1.425 $X2=0 $Y2=0
cc_377 N_SCE_c_373_n N_SCD_c_504_n 0.00914109f $X=2.56 $Y=1.425 $X2=0 $Y2=0
cc_378 N_SCE_c_379_n N_VPWR_c_1804_n 0.00645742f $X=1.115 $Y=2.245 $X2=0 $Y2=0
cc_379 N_SCE_c_381_n N_VPWR_c_1804_n 0.0139313f $X=1.615 $Y=2.245 $X2=0 $Y2=0
cc_380 N_SCE_c_379_n N_VPWR_c_1812_n 0.0044455f $X=1.115 $Y=2.245 $X2=0 $Y2=0
cc_381 N_SCE_c_381_n N_VPWR_c_1819_n 0.00413917f $X=1.615 $Y=2.245 $X2=0 $Y2=0
cc_382 N_SCE_c_379_n N_VPWR_c_1803_n 0.00858576f $X=1.115 $Y=2.245 $X2=0 $Y2=0
cc_383 N_SCE_c_381_n N_VPWR_c_1803_n 0.00817532f $X=1.615 $Y=2.245 $X2=0 $Y2=0
cc_384 N_SCE_M1033_g N_A_413_90#_c_1985_n 0.00897206f $X=2.65 $Y=0.695 $X2=0
+ $Y2=0
cc_385 N_SCE_c_372_n N_A_413_90#_c_1985_n 0.00904054f $X=2.56 $Y=1.425 $X2=0
+ $Y2=0
cc_386 N_SCE_c_381_n N_A_413_90#_c_1998_n 0.00175747f $X=1.615 $Y=2.245 $X2=0
+ $Y2=0
cc_387 N_SCE_M1033_g N_A_413_90#_c_1991_n 0.00996051f $X=2.65 $Y=0.695 $X2=0
+ $Y2=0
cc_388 N_SCE_c_371_n N_A_413_90#_c_1991_n 0.00563615f $X=2.395 $Y=1.575 $X2=0
+ $Y2=0
cc_389 N_SCE_c_372_n N_A_413_90#_c_1991_n 0.016885f $X=2.56 $Y=1.425 $X2=0 $Y2=0
cc_390 N_SCE_c_373_n N_A_413_90#_c_1991_n 0.0013723f $X=2.56 $Y=1.425 $X2=0
+ $Y2=0
cc_391 N_SCE_M1040_g N_VGND_c_2174_n 0.0141679f $X=0.495 $Y=0.58 $X2=0 $Y2=0
cc_392 N_SCE_M1033_g N_VGND_c_2181_n 7.35405e-19 $X=2.65 $Y=0.695 $X2=0 $Y2=0
cc_393 N_SCE_M1040_g N_VGND_c_2185_n 0.00383152f $X=0.495 $Y=0.58 $X2=0 $Y2=0
cc_394 N_SCE_M1040_g N_VGND_c_2190_n 0.00761198f $X=0.495 $Y=0.58 $X2=0 $Y2=0
cc_395 N_SCE_M1040_g N_noxref_25_c_2313_n 7.01965e-19 $X=0.495 $Y=0.58 $X2=0
+ $Y2=0
cc_396 N_SCE_M1033_g N_noxref_25_c_2314_n 0.00874184f $X=2.65 $Y=0.695 $X2=0
+ $Y2=0
cc_397 N_SCE_M1040_g N_noxref_25_c_2315_n 6.37214e-19 $X=0.495 $Y=0.58 $X2=0
+ $Y2=0
cc_398 N_D_c_462_n N_VPWR_c_1804_n 0.00220672f $X=2.035 $Y=2.245 $X2=0 $Y2=0
cc_399 N_D_c_462_n N_VPWR_c_1819_n 0.00445347f $X=2.035 $Y=2.245 $X2=0 $Y2=0
cc_400 N_D_c_462_n N_VPWR_c_1803_n 0.00858062f $X=2.035 $Y=2.245 $X2=0 $Y2=0
cc_401 N_D_c_462_n N_A_413_90#_c_1998_n 0.0110864f $X=2.035 $Y=2.245 $X2=0 $Y2=0
cc_402 N_D_c_458_n N_A_413_90#_c_1991_n 0.00100119f $X=1.935 $Y=1.145 $X2=0
+ $Y2=0
cc_403 N_D_c_459_n N_A_413_90#_c_1991_n 0.0209433f $X=1.935 $Y=1.145 $X2=0 $Y2=0
cc_404 N_D_c_460_n N_A_413_90#_c_1991_n 0.00597193f $X=1.947 $Y=0.98 $X2=0 $Y2=0
cc_405 N_D_c_460_n N_VGND_c_2181_n 8.05596e-19 $X=1.947 $Y=0.98 $X2=0 $Y2=0
cc_406 N_D_c_458_n N_noxref_25_c_2314_n 0.0014811f $X=1.935 $Y=1.145 $X2=0 $Y2=0
cc_407 N_D_c_459_n N_noxref_25_c_2314_n 0.0171941f $X=1.935 $Y=1.145 $X2=0 $Y2=0
cc_408 N_D_c_460_n N_noxref_25_c_2314_n 0.0105212f $X=1.947 $Y=0.98 $X2=0 $Y2=0
cc_409 N_D_c_459_n noxref_26 0.00381079f $X=1.935 $Y=1.145 $X2=-0.19 $Y2=-0.245
cc_410 N_SCD_M1015_g N_RESET_B_M1034_g 0.0253875f $X=3.04 $Y=0.695 $X2=0 $Y2=0
cc_411 SCD N_RESET_B_M1034_g 7.5908e-19 $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_412 N_SCD_c_504_n N_RESET_B_M1034_g 0.0176254f $X=3.1 $Y=1.605 $X2=0 $Y2=0
cc_413 N_SCD_c_505_n N_RESET_B_c_553_n 0.0166903f $X=3.025 $Y=2.245 $X2=0 $Y2=0
cc_414 N_SCD_c_502_n N_RESET_B_c_565_n 0.0213431f $X=3.1 $Y=1.945 $X2=0 $Y2=0
cc_415 N_SCD_c_505_n N_VPWR_c_1805_n 0.00926326f $X=3.025 $Y=2.245 $X2=0 $Y2=0
cc_416 N_SCD_c_505_n N_VPWR_c_1819_n 0.00413917f $X=3.025 $Y=2.245 $X2=0 $Y2=0
cc_417 N_SCD_c_505_n N_VPWR_c_1803_n 0.00399473f $X=3.025 $Y=2.245 $X2=0 $Y2=0
cc_418 N_SCD_M1015_g N_A_413_90#_c_1985_n 0.0133448f $X=3.04 $Y=0.695 $X2=0
+ $Y2=0
cc_419 SCD N_A_413_90#_c_1985_n 0.0147015f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_420 N_SCD_c_504_n N_A_413_90#_c_1985_n 0.00106413f $X=3.1 $Y=1.605 $X2=0
+ $Y2=0
cc_421 N_SCD_c_505_n N_A_413_90#_c_1986_n 0.00133463f $X=3.025 $Y=2.245 $X2=0
+ $Y2=0
cc_422 N_SCD_M1015_g N_A_413_90#_c_1986_n 0.00626156f $X=3.04 $Y=0.695 $X2=0
+ $Y2=0
cc_423 N_SCD_c_502_n N_A_413_90#_c_1986_n 0.00181592f $X=3.1 $Y=1.945 $X2=0
+ $Y2=0
cc_424 SCD N_A_413_90#_c_1986_n 0.051206f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_425 N_SCD_c_504_n N_A_413_90#_c_1986_n 0.00379786f $X=3.1 $Y=1.605 $X2=0
+ $Y2=0
cc_426 N_SCD_c_505_n N_A_413_90#_c_1994_n 6.08409e-19 $X=3.025 $Y=2.245 $X2=0
+ $Y2=0
cc_427 N_SCD_c_505_n N_A_413_90#_c_1998_n 0.00160234f $X=3.025 $Y=2.245 $X2=0
+ $Y2=0
cc_428 N_SCD_M1015_g N_A_413_90#_c_1991_n 0.00137758f $X=3.04 $Y=0.695 $X2=0
+ $Y2=0
cc_429 N_SCD_c_505_n N_A_413_90#_c_2004_n 0.0131275f $X=3.025 $Y=2.245 $X2=0
+ $Y2=0
cc_430 N_SCD_c_502_n N_A_413_90#_c_2004_n 7.80289e-19 $X=3.1 $Y=1.945 $X2=0
+ $Y2=0
cc_431 SCD N_A_413_90#_c_2004_n 0.0181419f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_432 N_SCD_c_505_n N_A_413_90#_c_1999_n 0.00158693f $X=3.025 $Y=2.245 $X2=0
+ $Y2=0
cc_433 N_SCD_M1015_g N_VGND_c_2181_n 7.35405e-19 $X=3.04 $Y=0.695 $X2=0 $Y2=0
cc_434 N_SCD_M1015_g N_noxref_25_c_2314_n 0.00828992f $X=3.04 $Y=0.695 $X2=0
+ $Y2=0
cc_435 N_SCD_M1015_g N_noxref_25_c_2316_n 0.00337997f $X=3.04 $Y=0.695 $X2=0
+ $Y2=0
cc_436 N_RESET_B_c_558_n N_CLK_c_766_n 0.002278f $X=7.775 $Y=2.035 $X2=0 $Y2=0
cc_437 N_RESET_B_M1034_g N_CLK_c_767_n 0.0116585f $X=3.58 $Y=0.65 $X2=0 $Y2=0
cc_438 N_RESET_B_c_558_n N_CLK_c_767_n 0.00231089f $X=7.775 $Y=2.035 $X2=0 $Y2=0
cc_439 N_RESET_B_c_559_n N_CLK_c_767_n 0.0013801f $X=4.225 $Y=2.035 $X2=0 $Y2=0
cc_440 N_RESET_B_c_565_n N_CLK_c_767_n 0.006271f $X=3.595 $Y=2.032 $X2=0 $Y2=0
cc_441 N_RESET_B_c_566_n N_CLK_c_767_n 0.00160713f $X=3.95 $Y=1.985 $X2=0 $Y2=0
cc_442 N_RESET_B_M1034_g N_CLK_c_768_n 0.00315336f $X=3.58 $Y=0.65 $X2=0 $Y2=0
cc_443 N_RESET_B_c_558_n N_CLK_c_768_n 0.00546318f $X=7.775 $Y=2.035 $X2=0 $Y2=0
cc_444 N_RESET_B_c_559_n N_CLK_c_768_n 0.00346896f $X=4.225 $Y=2.035 $X2=0 $Y2=0
cc_445 N_RESET_B_c_565_n N_CLK_c_768_n 7.52322e-19 $X=3.595 $Y=2.032 $X2=0 $Y2=0
cc_446 N_RESET_B_c_566_n N_CLK_c_768_n 0.00939458f $X=3.95 $Y=1.985 $X2=0 $Y2=0
cc_447 N_RESET_B_c_558_n N_A_1023_74#_c_833_n 0.00468421f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_448 N_RESET_B_c_558_n N_A_1023_74#_c_813_n 0.00384754f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_449 N_RESET_B_c_560_n N_A_1023_74#_c_836_n 0.0053373f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_450 N_RESET_B_M1017_g N_A_1023_74#_c_819_n 6.5419e-19 $X=7.31 $Y=0.695 $X2=0
+ $Y2=0
cc_451 N_RESET_B_c_558_n N_A_1023_74#_c_822_n 0.0359131f $X=7.775 $Y=2.035 $X2=0
+ $Y2=0
cc_452 N_RESET_B_c_558_n N_A_1023_74#_c_823_n 0.0158048f $X=7.775 $Y=2.035 $X2=0
+ $Y2=0
cc_453 N_RESET_B_M1017_g N_A_1023_74#_c_824_n 0.00177674f $X=7.31 $Y=0.695 $X2=0
+ $Y2=0
cc_454 N_RESET_B_M1017_g N_A_1023_74#_c_848_n 0.0125562f $X=7.31 $Y=0.695 $X2=0
+ $Y2=0
cc_455 N_RESET_B_c_549_n N_A_1023_74#_c_848_n 0.0013918f $X=7.605 $Y=1.145 $X2=0
+ $Y2=0
cc_456 N_RESET_B_M1017_g N_A_1023_74#_c_850_n 0.00387243f $X=7.31 $Y=0.695 $X2=0
+ $Y2=0
cc_457 N_RESET_B_c_560_n N_A_1023_74#_c_839_n 0.0136948f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_458 N_RESET_B_c_560_n N_A_1023_74#_c_831_n 0.0078678f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_459 N_RESET_B_c_558_n N_A_1023_74#_c_832_n 0.0038641f $X=7.775 $Y=2.035 $X2=0
+ $Y2=0
cc_460 N_RESET_B_c_560_n N_A_1369_71#_M1019_d 0.00328043f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_461 N_RESET_B_M1017_g N_A_1369_71#_M1016_g 0.0419455f $X=7.31 $Y=0.695 $X2=0
+ $Y2=0
cc_462 N_RESET_B_c_547_n N_A_1369_71#_M1016_g 0.00304499f $X=7.605 $Y=1.82 $X2=0
+ $Y2=0
cc_463 N_RESET_B_c_554_n N_A_1369_71#_c_1031_n 0.00631034f $X=7.555 $Y=2.24
+ $X2=0 $Y2=0
cc_464 N_RESET_B_c_547_n N_A_1369_71#_c_1031_n 0.0047841f $X=7.605 $Y=1.82 $X2=0
+ $Y2=0
cc_465 N_RESET_B_c_558_n N_A_1369_71#_c_1031_n 0.0115086f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_466 N_RESET_B_c_554_n N_A_1369_71#_c_1032_n 0.0131242f $X=7.555 $Y=2.24 $X2=0
+ $Y2=0
cc_467 N_RESET_B_c_547_n N_A_1369_71#_c_1023_n 0.00189704f $X=7.605 $Y=1.82
+ $X2=0 $Y2=0
cc_468 N_RESET_B_c_549_n N_A_1369_71#_c_1023_n 0.0031348f $X=7.605 $Y=1.145
+ $X2=0 $Y2=0
cc_469 N_RESET_B_c_558_n N_A_1369_71#_c_1023_n 0.00650511f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_470 N_RESET_B_c_547_n N_A_1369_71#_c_1024_n 0.0175446f $X=7.605 $Y=1.82 $X2=0
+ $Y2=0
cc_471 N_RESET_B_c_549_n N_A_1369_71#_c_1024_n 0.0040469f $X=7.605 $Y=1.145
+ $X2=0 $Y2=0
cc_472 N_RESET_B_c_558_n N_A_1369_71#_c_1024_n 0.00186974f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_473 N_RESET_B_M1017_g N_A_1369_71#_c_1025_n 0.00710957f $X=7.31 $Y=0.695
+ $X2=0 $Y2=0
cc_474 N_RESET_B_c_549_n N_A_1369_71#_c_1025_n 0.015222f $X=7.605 $Y=1.145 $X2=0
+ $Y2=0
cc_475 N_RESET_B_M1017_g N_A_1369_71#_c_1026_n 0.00106261f $X=7.31 $Y=0.695
+ $X2=0 $Y2=0
cc_476 N_RESET_B_c_549_n N_A_1369_71#_c_1026_n 2.71646e-19 $X=7.605 $Y=1.145
+ $X2=0 $Y2=0
cc_477 N_RESET_B_c_560_n N_A_1369_71#_c_1028_n 0.00664109f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_478 N_RESET_B_c_560_n N_A_1369_71#_c_1029_n 0.0247803f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_479 N_RESET_B_c_549_n N_A_1221_97#_M1041_g 0.00544172f $X=7.605 $Y=1.145
+ $X2=0 $Y2=0
cc_480 N_RESET_B_c_560_n N_A_1221_97#_c_1137_n 0.00728194f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_481 N_RESET_B_M1017_g N_A_1221_97#_c_1131_n 8.68322e-19 $X=7.31 $Y=0.695
+ $X2=0 $Y2=0
cc_482 N_RESET_B_c_558_n N_A_1221_97#_c_1138_n 0.00858152f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_483 N_RESET_B_c_558_n N_A_1221_97#_c_1132_n 0.025309f $X=7.775 $Y=2.035 $X2=0
+ $Y2=0
cc_484 N_RESET_B_c_558_n N_A_1221_97#_c_1148_n 0.0199315f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_485 N_RESET_B_c_554_n N_A_1221_97#_c_1133_n 0.037162f $X=7.555 $Y=2.24 $X2=0
+ $Y2=0
cc_486 N_RESET_B_c_547_n N_A_1221_97#_c_1133_n 0.0102695f $X=7.605 $Y=1.82 $X2=0
+ $Y2=0
cc_487 N_RESET_B_c_558_n N_A_1221_97#_c_1133_n 0.0312198f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_488 N_RESET_B_c_561_n N_A_1221_97#_c_1133_n 0.00470341f $X=8.065 $Y=2.035
+ $X2=0 $Y2=0
cc_489 N_RESET_B_c_564_n N_A_1221_97#_c_1133_n 0.0355881f $X=7.86 $Y=1.985 $X2=0
+ $Y2=0
cc_490 N_RESET_B_c_547_n N_A_1221_97#_c_1134_n 0.00423725f $X=7.605 $Y=1.82
+ $X2=0 $Y2=0
cc_491 N_RESET_B_c_549_n N_A_1221_97#_c_1134_n 0.00287951f $X=7.605 $Y=1.145
+ $X2=0 $Y2=0
cc_492 N_RESET_B_c_547_n N_A_1221_97#_c_1135_n 0.00921867f $X=7.605 $Y=1.82
+ $X2=0 $Y2=0
cc_493 N_RESET_B_c_558_n N_A_1221_97#_c_1135_n 0.00551265f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_494 N_RESET_B_c_560_n N_A_1221_97#_c_1135_n 0.00588285f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_495 N_RESET_B_c_561_n N_A_1221_97#_c_1135_n 0.0026603f $X=8.065 $Y=2.035
+ $X2=0 $Y2=0
cc_496 N_RESET_B_c_563_n N_A_1221_97#_c_1135_n 0.00668769f $X=7.86 $Y=1.985
+ $X2=0 $Y2=0
cc_497 N_RESET_B_c_564_n N_A_1221_97#_c_1135_n 0.0134428f $X=7.86 $Y=1.985 $X2=0
+ $Y2=0
cc_498 N_RESET_B_c_547_n N_A_1221_97#_c_1136_n 0.0179208f $X=7.605 $Y=1.82 $X2=0
+ $Y2=0
cc_499 N_RESET_B_c_560_n N_A_1221_97#_c_1136_n 0.00424919f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_500 N_RESET_B_c_561_n N_A_1221_97#_c_1136_n 7.15345e-19 $X=8.065 $Y=2.035
+ $X2=0 $Y2=0
cc_501 N_RESET_B_c_563_n N_A_1221_97#_c_1136_n 0.00483051f $X=7.86 $Y=1.985
+ $X2=0 $Y2=0
cc_502 N_RESET_B_c_564_n N_A_1221_97#_c_1136_n 5.47888e-19 $X=7.86 $Y=1.985
+ $X2=0 $Y2=0
cc_503 N_RESET_B_c_558_n N_A_850_74#_M1025_s 0.00117465f $X=7.775 $Y=2.035 $X2=0
+ $Y2=0
cc_504 N_RESET_B_c_558_n N_A_850_74#_c_1246_n 0.0046943f $X=7.775 $Y=2.035 $X2=0
+ $Y2=0
cc_505 N_RESET_B_c_558_n N_A_850_74#_c_1248_n 0.00212115f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_506 N_RESET_B_c_558_n N_A_850_74#_c_1266_n 0.00273429f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_507 N_RESET_B_c_554_n N_A_850_74#_c_1267_n 0.0100134f $X=7.555 $Y=2.24 $X2=0
+ $Y2=0
cc_508 N_RESET_B_c_560_n N_A_850_74#_M1023_g 0.0105606f $X=10.655 $Y=2.035 $X2=0
+ $Y2=0
cc_509 N_RESET_B_c_560_n N_A_850_74#_c_1251_n 0.00463969f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_510 N_RESET_B_M1034_g N_A_850_74#_c_1255_n 0.00357469f $X=3.58 $Y=0.65 $X2=0
+ $Y2=0
cc_511 N_RESET_B_M1034_g N_A_850_74#_c_1256_n 0.0023811f $X=3.58 $Y=0.65 $X2=0
+ $Y2=0
cc_512 N_RESET_B_c_558_n N_A_850_74#_c_1274_n 0.0150045f $X=7.775 $Y=2.035 $X2=0
+ $Y2=0
cc_513 N_RESET_B_M1034_g N_A_850_74#_c_1276_n 4.14135e-19 $X=3.58 $Y=0.65 $X2=0
+ $Y2=0
cc_514 N_RESET_B_c_558_n N_A_850_74#_c_1276_n 0.0148387f $X=7.775 $Y=2.035 $X2=0
+ $Y2=0
cc_515 N_RESET_B_c_559_n N_A_850_74#_c_1276_n 0.00279861f $X=4.225 $Y=2.035
+ $X2=0 $Y2=0
cc_516 N_RESET_B_c_565_n N_A_850_74#_c_1276_n 0.00168423f $X=3.595 $Y=2.032
+ $X2=0 $Y2=0
cc_517 N_RESET_B_c_566_n N_A_850_74#_c_1276_n 0.0240051f $X=3.95 $Y=1.985 $X2=0
+ $Y2=0
cc_518 N_RESET_B_c_558_n N_A_850_74#_c_1259_n 0.00708562f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_519 N_RESET_B_M1007_g N_A_2008_48#_M1005_g 0.0358144f $X=10.545 $Y=0.58 $X2=0
+ $Y2=0
cc_520 N_RESET_B_c_551_n N_A_2008_48#_M1005_g 0.00188557f $X=10.9 $Y=1.68 $X2=0
+ $Y2=0
cc_521 N_RESET_B_c_550_n N_A_2008_48#_c_1438_n 0.0030428f $X=10.81 $Y=1.335
+ $X2=0 $Y2=0
cc_522 N_RESET_B_c_560_n N_A_2008_48#_c_1438_n 0.00247648f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_523 RESET_B N_A_2008_48#_c_1438_n 7.14482e-19 $X=10.715 $Y=1.95 $X2=0 $Y2=0
cc_524 N_RESET_B_c_568_n N_A_2008_48#_c_1438_n 0.00169359f $X=10.9 $Y=1.845
+ $X2=0 $Y2=0
cc_525 N_RESET_B_c_551_n N_A_2008_48#_c_1438_n 0.0249721f $X=10.9 $Y=1.68 $X2=0
+ $Y2=0
cc_526 N_RESET_B_c_556_n N_A_2008_48#_c_1445_n 0.00373821f $X=10.81 $Y=2.22
+ $X2=0 $Y2=0
cc_527 N_RESET_B_c_557_n N_A_2008_48#_c_1445_n 0.00276573f $X=10.81 $Y=2.37
+ $X2=0 $Y2=0
cc_528 N_RESET_B_c_560_n N_A_2008_48#_c_1445_n 0.00755701f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_529 N_RESET_B_c_567_n N_A_2008_48#_c_1445_n 6.88508e-19 $X=10.9 $Y=1.845
+ $X2=0 $Y2=0
cc_530 N_RESET_B_c_557_n N_A_2008_48#_c_1446_n 0.0107901f $X=10.81 $Y=2.37 $X2=0
+ $Y2=0
cc_531 N_RESET_B_c_556_n N_A_2008_48#_c_1439_n 0.00199769f $X=10.81 $Y=2.22
+ $X2=0 $Y2=0
cc_532 N_RESET_B_c_557_n N_A_2008_48#_c_1439_n 0.00241136f $X=10.81 $Y=2.37
+ $X2=0 $Y2=0
cc_533 N_RESET_B_c_560_n N_A_2008_48#_c_1439_n 0.0174665f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_534 RESET_B N_A_2008_48#_c_1439_n 0.00269473f $X=10.715 $Y=1.95 $X2=0 $Y2=0
cc_535 N_RESET_B_c_567_n N_A_2008_48#_c_1439_n 4.38169e-19 $X=10.9 $Y=1.845
+ $X2=0 $Y2=0
cc_536 N_RESET_B_c_568_n N_A_2008_48#_c_1439_n 0.0344591f $X=10.9 $Y=1.845 $X2=0
+ $Y2=0
cc_537 N_RESET_B_c_551_n N_A_2008_48#_c_1439_n 2.34208e-19 $X=10.9 $Y=1.68 $X2=0
+ $Y2=0
cc_538 N_RESET_B_c_557_n N_A_2008_48#_c_1448_n 0.00976826f $X=10.81 $Y=2.37
+ $X2=0 $Y2=0
cc_539 N_RESET_B_c_560_n N_A_2008_48#_c_1448_n 0.00560031f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_540 RESET_B N_A_2008_48#_c_1448_n 0.00309934f $X=10.715 $Y=1.95 $X2=0 $Y2=0
cc_541 N_RESET_B_c_568_n N_A_2008_48#_c_1448_n 0.00989058f $X=10.9 $Y=1.845
+ $X2=0 $Y2=0
cc_542 N_RESET_B_c_557_n N_A_2008_48#_c_1450_n 0.00646344f $X=10.81 $Y=2.37
+ $X2=0 $Y2=0
cc_543 N_RESET_B_c_556_n N_A_2008_48#_c_1451_n 0.0015825f $X=10.81 $Y=2.22 $X2=0
+ $Y2=0
cc_544 N_RESET_B_c_557_n N_A_2008_48#_c_1451_n 5.62382e-19 $X=10.81 $Y=2.37
+ $X2=0 $Y2=0
cc_545 RESET_B N_A_2008_48#_c_1451_n 0.00125949f $X=10.715 $Y=1.95 $X2=0 $Y2=0
cc_546 N_RESET_B_c_567_n N_A_2008_48#_c_1451_n 0.00110518f $X=10.9 $Y=1.845
+ $X2=0 $Y2=0
cc_547 N_RESET_B_c_568_n N_A_2008_48#_c_1451_n 0.0258608f $X=10.9 $Y=1.845 $X2=0
+ $Y2=0
cc_548 N_RESET_B_c_567_n N_A_2008_48#_c_1441_n 8.24141e-19 $X=10.9 $Y=1.845
+ $X2=0 $Y2=0
cc_549 N_RESET_B_c_568_n N_A_2008_48#_c_1441_n 0.00968802f $X=10.9 $Y=1.845
+ $X2=0 $Y2=0
cc_550 N_RESET_B_c_551_n N_A_2008_48#_c_1441_n 0.00111902f $X=10.9 $Y=1.68 $X2=0
+ $Y2=0
cc_551 N_RESET_B_c_557_n N_A_2008_48#_c_1454_n 0.00389165f $X=10.81 $Y=2.37
+ $X2=0 $Y2=0
cc_552 RESET_B N_A_2008_48#_c_1454_n 7.29139e-19 $X=10.715 $Y=1.95 $X2=0 $Y2=0
cc_553 N_RESET_B_c_567_n N_A_2008_48#_c_1454_n 8.21335e-19 $X=10.9 $Y=1.845
+ $X2=0 $Y2=0
cc_554 N_RESET_B_c_568_n N_A_2008_48#_c_1454_n 0.0169044f $X=10.9 $Y=1.845 $X2=0
+ $Y2=0
cc_555 N_RESET_B_M1007_g N_A_2008_48#_c_1443_n 0.00108873f $X=10.545 $Y=0.58
+ $X2=0 $Y2=0
cc_556 N_RESET_B_c_560_n N_A_1747_74#_M1023_d 0.00220193f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_557 N_RESET_B_M1007_g N_A_1747_74#_c_1573_n 0.0481778f $X=10.545 $Y=0.58
+ $X2=0 $Y2=0
cc_558 N_RESET_B_c_550_n N_A_1747_74#_c_1574_n 0.00304958f $X=10.81 $Y=1.335
+ $X2=0 $Y2=0
cc_559 N_RESET_B_c_567_n N_A_1747_74#_c_1574_n 0.00202705f $X=10.9 $Y=1.845
+ $X2=0 $Y2=0
cc_560 N_RESET_B_M1007_g N_A_1747_74#_c_1575_n 0.00503338f $X=10.545 $Y=0.58
+ $X2=0 $Y2=0
cc_561 N_RESET_B_c_557_n N_A_1747_74#_c_1585_n 0.00937718f $X=10.81 $Y=2.37
+ $X2=0 $Y2=0
cc_562 N_RESET_B_c_556_n N_A_1747_74#_c_1586_n 0.00655145f $X=10.81 $Y=2.22
+ $X2=0 $Y2=0
cc_563 N_RESET_B_c_568_n N_A_1747_74#_c_1586_n 8.64724e-19 $X=10.9 $Y=1.845
+ $X2=0 $Y2=0
cc_564 N_RESET_B_c_550_n N_A_1747_74#_c_1578_n 0.0113835f $X=10.81 $Y=1.335
+ $X2=0 $Y2=0
cc_565 N_RESET_B_c_567_n N_A_1747_74#_c_1578_n 0.0205072f $X=10.9 $Y=1.845 $X2=0
+ $Y2=0
cc_566 N_RESET_B_c_551_n N_A_1747_74#_c_1578_n 0.00965718f $X=10.9 $Y=1.68 $X2=0
+ $Y2=0
cc_567 N_RESET_B_c_557_n N_A_1747_74#_c_1592_n 0.00814266f $X=10.81 $Y=2.37
+ $X2=0 $Y2=0
cc_568 N_RESET_B_c_560_n N_A_1747_74#_c_1609_n 0.0211312f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_569 N_RESET_B_c_557_n N_A_1747_74#_c_1594_n 7.86001e-19 $X=10.81 $Y=2.37
+ $X2=0 $Y2=0
cc_570 N_RESET_B_c_560_n N_A_1747_74#_c_1594_n 0.0154438f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_571 N_RESET_B_c_560_n N_A_1747_74#_c_1582_n 0.0224891f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_572 N_RESET_B_c_551_n N_A_1747_74#_c_1582_n 9.47605e-19 $X=10.9 $Y=1.68 $X2=0
+ $Y2=0
cc_573 N_RESET_B_M1007_g N_A_1747_74#_c_1584_n 0.0173454f $X=10.545 $Y=0.58
+ $X2=0 $Y2=0
cc_574 N_RESET_B_c_550_n N_A_1747_74#_c_1584_n 0.0168092f $X=10.81 $Y=1.335
+ $X2=0 $Y2=0
cc_575 N_RESET_B_c_560_n N_A_1747_74#_c_1584_n 0.0108974f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_576 RESET_B N_A_1747_74#_c_1584_n 0.00277891f $X=10.715 $Y=1.95 $X2=0 $Y2=0
cc_577 N_RESET_B_c_567_n N_A_1747_74#_c_1584_n 0.00194273f $X=10.9 $Y=1.845
+ $X2=0 $Y2=0
cc_578 N_RESET_B_c_568_n N_A_1747_74#_c_1584_n 0.0211796f $X=10.9 $Y=1.845 $X2=0
+ $Y2=0
cc_579 N_RESET_B_c_551_n N_A_1747_74#_c_1584_n 0.00355179f $X=10.9 $Y=1.68 $X2=0
+ $Y2=0
cc_580 N_RESET_B_c_558_n N_VPWR_M1025_d 0.00290995f $X=7.775 $Y=2.035 $X2=0
+ $Y2=0
cc_581 N_RESET_B_c_560_n N_VPWR_M1019_s 0.00248619f $X=10.655 $Y=2.035 $X2=0
+ $Y2=0
cc_582 N_RESET_B_c_553_n N_VPWR_c_1805_n 0.00494016f $X=3.595 $Y=2.245 $X2=0
+ $Y2=0
cc_583 N_RESET_B_c_554_n N_VPWR_c_1807_n 0.00412651f $X=7.555 $Y=2.24 $X2=0
+ $Y2=0
cc_584 N_RESET_B_c_558_n N_VPWR_c_1807_n 6.86441e-19 $X=7.775 $Y=2.035 $X2=0
+ $Y2=0
cc_585 N_RESET_B_c_554_n N_VPWR_c_1808_n 0.00588806f $X=7.555 $Y=2.24 $X2=0
+ $Y2=0
cc_586 N_RESET_B_c_547_n N_VPWR_c_1808_n 0.00159571f $X=7.605 $Y=1.82 $X2=0
+ $Y2=0
cc_587 N_RESET_B_c_560_n N_VPWR_c_1808_n 0.025533f $X=10.655 $Y=2.035 $X2=0
+ $Y2=0
cc_588 N_RESET_B_c_561_n N_VPWR_c_1808_n 0.00264729f $X=8.065 $Y=2.035 $X2=0
+ $Y2=0
cc_589 N_RESET_B_c_563_n N_VPWR_c_1808_n 0.00114271f $X=7.86 $Y=1.985 $X2=0
+ $Y2=0
cc_590 N_RESET_B_c_564_n N_VPWR_c_1808_n 0.0204823f $X=7.86 $Y=1.985 $X2=0 $Y2=0
cc_591 N_RESET_B_c_557_n N_VPWR_c_1809_n 0.00552432f $X=10.81 $Y=2.37 $X2=0
+ $Y2=0
cc_592 N_RESET_B_c_560_n N_VPWR_c_1809_n 0.00114209f $X=10.655 $Y=2.035 $X2=0
+ $Y2=0
cc_593 N_RESET_B_c_553_n N_VPWR_c_1814_n 0.00399297f $X=3.595 $Y=2.245 $X2=0
+ $Y2=0
cc_594 N_RESET_B_c_557_n N_VPWR_c_1822_n 0.00497687f $X=10.81 $Y=2.37 $X2=0
+ $Y2=0
cc_595 N_RESET_B_c_553_n N_VPWR_c_1803_n 0.0042041f $X=3.595 $Y=2.245 $X2=0
+ $Y2=0
cc_596 N_RESET_B_c_554_n N_VPWR_c_1803_n 9.39239e-19 $X=7.555 $Y=2.24 $X2=0
+ $Y2=0
cc_597 N_RESET_B_c_557_n N_VPWR_c_1803_n 0.00515964f $X=10.81 $Y=2.37 $X2=0
+ $Y2=0
cc_598 N_RESET_B_M1034_g N_A_413_90#_c_1985_n 0.0147713f $X=3.58 $Y=0.65 $X2=0
+ $Y2=0
cc_599 N_RESET_B_M1034_g N_A_413_90#_c_1986_n 0.028357f $X=3.58 $Y=0.65 $X2=0
+ $Y2=0
cc_600 N_RESET_B_c_553_n N_A_413_90#_c_1986_n 0.00430128f $X=3.595 $Y=2.245
+ $X2=0 $Y2=0
cc_601 N_RESET_B_c_559_n N_A_413_90#_c_1986_n 0.00108246f $X=4.225 $Y=2.035
+ $X2=0 $Y2=0
cc_602 N_RESET_B_c_565_n N_A_413_90#_c_1986_n 0.0146661f $X=3.595 $Y=2.032 $X2=0
+ $Y2=0
cc_603 N_RESET_B_c_566_n N_A_413_90#_c_1986_n 0.0228178f $X=3.95 $Y=1.985 $X2=0
+ $Y2=0
cc_604 N_RESET_B_c_553_n N_A_413_90#_c_1994_n 0.00864976f $X=3.595 $Y=2.245
+ $X2=0 $Y2=0
cc_605 N_RESET_B_c_558_n N_A_413_90#_c_1995_n 0.0279449f $X=7.775 $Y=2.035 $X2=0
+ $Y2=0
cc_606 N_RESET_B_c_559_n N_A_413_90#_c_1995_n 0.0071452f $X=4.225 $Y=2.035 $X2=0
+ $Y2=0
cc_607 N_RESET_B_c_565_n N_A_413_90#_c_1995_n 0.00213778f $X=3.595 $Y=2.032
+ $X2=0 $Y2=0
cc_608 N_RESET_B_c_566_n N_A_413_90#_c_1995_n 0.00970518f $X=3.95 $Y=1.985 $X2=0
+ $Y2=0
cc_609 N_RESET_B_c_558_n N_A_413_90#_c_1996_n 0.0199642f $X=7.775 $Y=2.035 $X2=0
+ $Y2=0
cc_610 N_RESET_B_c_558_n N_A_413_90#_c_1990_n 0.0113119f $X=7.775 $Y=2.035 $X2=0
+ $Y2=0
cc_611 N_RESET_B_c_553_n N_A_413_90#_c_1999_n 0.0117793f $X=3.595 $Y=2.245 $X2=0
+ $Y2=0
cc_612 N_RESET_B_c_559_n N_A_413_90#_c_1999_n 0.00119344f $X=4.225 $Y=2.035
+ $X2=0 $Y2=0
cc_613 N_RESET_B_c_565_n N_A_413_90#_c_1999_n 0.00736185f $X=3.595 $Y=2.032
+ $X2=0 $Y2=0
cc_614 N_RESET_B_c_566_n N_A_413_90#_c_1999_n 0.0145688f $X=3.95 $Y=1.985 $X2=0
+ $Y2=0
cc_615 N_RESET_B_c_558_n N_A_413_90#_c_2000_n 0.0131914f $X=7.775 $Y=2.035 $X2=0
+ $Y2=0
cc_616 N_RESET_B_M1034_g N_VGND_c_2175_n 0.00305751f $X=3.58 $Y=0.65 $X2=0 $Y2=0
cc_617 N_RESET_B_M1017_g N_VGND_c_2177_n 0.00166614f $X=7.31 $Y=0.695 $X2=0
+ $Y2=0
cc_618 N_RESET_B_M1007_g N_VGND_c_2178_n 0.0110663f $X=10.545 $Y=0.58 $X2=0
+ $Y2=0
cc_619 N_RESET_B_M1034_g N_VGND_c_2181_n 0.00527445f $X=3.58 $Y=0.65 $X2=0 $Y2=0
cc_620 N_RESET_B_M1017_g N_VGND_c_2186_n 0.00378369f $X=7.31 $Y=0.695 $X2=0
+ $Y2=0
cc_621 N_RESET_B_M1007_g N_VGND_c_2188_n 0.00383152f $X=10.545 $Y=0.58 $X2=0
+ $Y2=0
cc_622 N_RESET_B_M1034_g N_VGND_c_2190_n 0.00523671f $X=3.58 $Y=0.65 $X2=0 $Y2=0
cc_623 N_RESET_B_M1017_g N_VGND_c_2190_n 0.00509887f $X=7.31 $Y=0.695 $X2=0
+ $Y2=0
cc_624 N_RESET_B_M1007_g N_VGND_c_2190_n 0.0075694f $X=10.545 $Y=0.58 $X2=0
+ $Y2=0
cc_625 N_RESET_B_M1034_g N_noxref_25_c_2316_n 0.00190287f $X=3.58 $Y=0.65 $X2=0
+ $Y2=0
cc_626 N_CLK_c_766_n N_A_1023_74#_c_822_n 6.38919e-19 $X=4.645 $Y=1.745 $X2=0
+ $Y2=0
cc_627 N_CLK_c_765_n N_A_850_74#_c_1245_n 0.0170522f $X=4.61 $Y=1.22 $X2=0 $Y2=0
cc_628 N_CLK_c_766_n N_A_850_74#_c_1246_n 0.0755118f $X=4.645 $Y=1.745 $X2=0
+ $Y2=0
cc_629 N_CLK_c_768_n N_A_850_74#_c_1246_n 2.13741e-19 $X=4.48 $Y=1.385 $X2=0
+ $Y2=0
cc_630 N_CLK_c_767_n N_A_850_74#_c_1255_n 0.00175971f $X=4.535 $Y=1.385 $X2=0
+ $Y2=0
cc_631 N_CLK_c_768_n N_A_850_74#_c_1255_n 0.021751f $X=4.48 $Y=1.385 $X2=0 $Y2=0
cc_632 N_CLK_c_765_n N_A_850_74#_c_1256_n 8.26992e-19 $X=4.61 $Y=1.22 $X2=0
+ $Y2=0
cc_633 N_CLK_c_765_n N_A_850_74#_c_1299_n 0.0107807f $X=4.61 $Y=1.22 $X2=0 $Y2=0
cc_634 N_CLK_c_768_n N_A_850_74#_c_1299_n 0.0102243f $X=4.48 $Y=1.385 $X2=0
+ $Y2=0
cc_635 N_CLK_c_766_n N_A_850_74#_c_1274_n 0.0112467f $X=4.645 $Y=1.745 $X2=0
+ $Y2=0
cc_636 N_CLK_c_768_n N_A_850_74#_c_1274_n 0.0028392f $X=4.48 $Y=1.385 $X2=0
+ $Y2=0
cc_637 N_CLK_c_765_n N_A_850_74#_c_1257_n 0.00452733f $X=4.61 $Y=1.22 $X2=0
+ $Y2=0
cc_638 N_CLK_c_768_n N_A_850_74#_c_1257_n 0.00946739f $X=4.48 $Y=1.385 $X2=0
+ $Y2=0
cc_639 N_CLK_c_766_n N_A_850_74#_c_1258_n 0.00390175f $X=4.645 $Y=1.745 $X2=0
+ $Y2=0
cc_640 N_CLK_c_766_n N_A_850_74#_c_1276_n 0.00502987f $X=4.645 $Y=1.745 $X2=0
+ $Y2=0
cc_641 N_CLK_c_767_n N_A_850_74#_c_1276_n 0.00482708f $X=4.535 $Y=1.385 $X2=0
+ $Y2=0
cc_642 N_CLK_c_768_n N_A_850_74#_c_1276_n 0.0135888f $X=4.48 $Y=1.385 $X2=0
+ $Y2=0
cc_643 N_CLK_c_766_n N_A_850_74#_c_1259_n 0.00422605f $X=4.645 $Y=1.745 $X2=0
+ $Y2=0
cc_644 N_CLK_c_768_n N_A_850_74#_c_1259_n 0.0214634f $X=4.48 $Y=1.385 $X2=0
+ $Y2=0
cc_645 N_CLK_c_766_n N_VPWR_c_1806_n 0.0182454f $X=4.645 $Y=1.745 $X2=0 $Y2=0
cc_646 N_CLK_c_766_n N_VPWR_c_1814_n 0.00505726f $X=4.645 $Y=1.745 $X2=0 $Y2=0
cc_647 N_CLK_c_766_n N_VPWR_c_1803_n 0.00489105f $X=4.645 $Y=1.745 $X2=0 $Y2=0
cc_648 N_CLK_c_767_n N_A_413_90#_c_1986_n 3.90147e-19 $X=4.535 $Y=1.385 $X2=0
+ $Y2=0
cc_649 N_CLK_c_768_n N_A_413_90#_c_1986_n 0.0173888f $X=4.48 $Y=1.385 $X2=0
+ $Y2=0
cc_650 N_CLK_c_766_n N_A_413_90#_c_1994_n 0.0107559f $X=4.645 $Y=1.745 $X2=0
+ $Y2=0
cc_651 N_CLK_c_766_n N_A_413_90#_c_1995_n 0.0146251f $X=4.645 $Y=1.745 $X2=0
+ $Y2=0
cc_652 N_CLK_c_766_n N_A_413_90#_c_1999_n 0.00178667f $X=4.645 $Y=1.745 $X2=0
+ $Y2=0
cc_653 N_CLK_c_765_n N_VGND_c_2175_n 0.00241532f $X=4.61 $Y=1.22 $X2=0 $Y2=0
cc_654 N_CLK_c_768_n N_VGND_c_2175_n 0.00156407f $X=4.48 $Y=1.385 $X2=0 $Y2=0
cc_655 N_CLK_c_765_n N_VGND_c_2176_n 0.0082347f $X=4.61 $Y=1.22 $X2=0 $Y2=0
cc_656 N_CLK_c_765_n N_VGND_c_2183_n 0.00383152f $X=4.61 $Y=1.22 $X2=0 $Y2=0
cc_657 N_CLK_c_765_n N_VGND_c_2190_n 0.00388966f $X=4.61 $Y=1.22 $X2=0 $Y2=0
cc_658 N_A_1023_74#_c_825_n N_A_1369_71#_M1041_d 0.00176461f $X=8.78 $Y=0.34
+ $X2=-0.19 $Y2=-0.245
cc_659 N_A_1023_74#_M1004_g N_A_1369_71#_M1016_g 0.0338256f $X=6.53 $Y=0.695
+ $X2=0 $Y2=0
cc_660 N_A_1023_74#_c_819_n N_A_1369_71#_M1016_g 0.0112527f $X=7.015 $Y=0.34
+ $X2=0 $Y2=0
cc_661 N_A_1023_74#_c_824_n N_A_1369_71#_M1016_g 0.00185656f $X=7.1 $Y=0.595
+ $X2=0 $Y2=0
cc_662 N_A_1023_74#_c_833_n N_A_1369_71#_c_1031_n 0.00179782f $X=6.115 $Y=2.15
+ $X2=0 $Y2=0
cc_663 N_A_1023_74#_c_832_n N_A_1369_71#_c_1031_n 0.00146462f $X=6.055 $Y=1.65
+ $X2=0 $Y2=0
cc_664 N_A_1023_74#_c_834_n N_A_1369_71#_c_1032_n 0.00179782f $X=6.115 $Y=2.24
+ $X2=0 $Y2=0
cc_665 N_A_1023_74#_c_813_n N_A_1369_71#_c_1024_n 0.0338256f $X=6.455 $Y=1.65
+ $X2=0 $Y2=0
cc_666 N_A_1023_74#_c_863_p N_A_1369_71#_c_1024_n 4.39545e-19 $X=7.185 $Y=0.68
+ $X2=0 $Y2=0
cc_667 N_A_1023_74#_c_832_n N_A_1369_71#_c_1024_n 4.00257e-19 $X=6.055 $Y=1.65
+ $X2=0 $Y2=0
cc_668 N_A_1023_74#_c_848_n N_A_1369_71#_c_1025_n 0.0615902f $X=7.94 $Y=0.68
+ $X2=0 $Y2=0
cc_669 N_A_1023_74#_c_825_n N_A_1369_71#_c_1025_n 0.0034413f $X=8.78 $Y=0.34
+ $X2=0 $Y2=0
cc_670 N_A_1023_74#_c_863_p N_A_1369_71#_c_1026_n 0.0134072f $X=7.185 $Y=0.68
+ $X2=0 $Y2=0
cc_671 N_A_1023_74#_c_815_n N_A_1369_71#_c_1068_n 0.0041679f $X=8.66 $Y=1.085
+ $X2=0 $Y2=0
cc_672 N_A_1023_74#_c_825_n N_A_1369_71#_c_1068_n 0.0158584f $X=8.78 $Y=0.34
+ $X2=0 $Y2=0
cc_673 N_A_1023_74#_c_817_n N_A_1369_71#_c_1027_n 0.00444121f $X=8.735 $Y=1.16
+ $X2=0 $Y2=0
cc_674 N_A_1023_74#_c_827_n N_A_1369_71#_c_1027_n 0.00425045f $X=9.27 $Y=1.345
+ $X2=0 $Y2=0
cc_675 N_A_1023_74#_c_817_n N_A_1369_71#_c_1028_n 0.010636f $X=8.735 $Y=1.16
+ $X2=0 $Y2=0
cc_676 N_A_1023_74#_c_827_n N_A_1369_71#_c_1028_n 0.00854237f $X=9.27 $Y=1.345
+ $X2=0 $Y2=0
cc_677 N_A_1023_74#_c_829_n N_A_1369_71#_c_1028_n 0.011663f $X=9.27 $Y=1.07
+ $X2=0 $Y2=0
cc_678 N_A_1023_74#_c_831_n N_A_1369_71#_c_1028_n 0.00620138f $X=9.63 $Y=1.46
+ $X2=0 $Y2=0
cc_679 N_A_1023_74#_c_839_n N_A_1369_71#_c_1029_n 0.00513948f $X=9.67 $Y=2.065
+ $X2=0 $Y2=0
cc_680 N_A_1023_74#_c_831_n N_A_1369_71#_c_1029_n 0.0132001f $X=9.63 $Y=1.46
+ $X2=0 $Y2=0
cc_681 N_A_1023_74#_c_815_n N_A_1369_71#_c_1030_n 0.00251445f $X=8.66 $Y=1.085
+ $X2=0 $Y2=0
cc_682 N_A_1023_74#_c_817_n N_A_1369_71#_c_1030_n 8.10451e-19 $X=8.735 $Y=1.16
+ $X2=0 $Y2=0
cc_683 N_A_1023_74#_c_827_n N_A_1369_71#_c_1030_n 9.81795e-19 $X=9.27 $Y=1.345
+ $X2=0 $Y2=0
cc_684 N_A_1023_74#_c_829_n N_A_1369_71#_c_1030_n 0.00881609f $X=9.27 $Y=1.07
+ $X2=0 $Y2=0
cc_685 N_A_1023_74#_c_815_n N_A_1221_97#_M1041_g 0.0262081f $X=8.66 $Y=1.085
+ $X2=0 $Y2=0
cc_686 N_A_1023_74#_c_825_n N_A_1221_97#_M1041_g 0.0116741f $X=8.78 $Y=0.34
+ $X2=0 $Y2=0
cc_687 N_A_1023_74#_c_813_n N_A_1221_97#_c_1131_n 5.54149e-19 $X=6.455 $Y=1.65
+ $X2=0 $Y2=0
cc_688 N_A_1023_74#_M1004_g N_A_1221_97#_c_1131_n 0.0157041f $X=6.53 $Y=0.695
+ $X2=0 $Y2=0
cc_689 N_A_1023_74#_c_819_n N_A_1221_97#_c_1131_n 0.0438127f $X=7.015 $Y=0.34
+ $X2=0 $Y2=0
cc_690 N_A_1023_74#_c_834_n N_A_1221_97#_c_1138_n 0.00408911f $X=6.115 $Y=2.24
+ $X2=0 $Y2=0
cc_691 N_A_1023_74#_c_813_n N_A_1221_97#_c_1138_n 9.38112e-19 $X=6.455 $Y=1.65
+ $X2=0 $Y2=0
cc_692 N_A_1023_74#_c_833_n N_A_1221_97#_c_1132_n 3.98198e-19 $X=6.115 $Y=2.15
+ $X2=0 $Y2=0
cc_693 N_A_1023_74#_M1004_g N_A_1221_97#_c_1132_n 0.00803125f $X=6.53 $Y=0.695
+ $X2=0 $Y2=0
cc_694 N_A_1023_74#_c_817_n N_A_1221_97#_c_1136_n 0.00320051f $X=8.735 $Y=1.16
+ $X2=0 $Y2=0
cc_695 N_A_1023_74#_c_820_n N_A_850_74#_c_1245_n 0.00266901f $X=5.42 $Y=0.34
+ $X2=0 $Y2=0
cc_696 N_A_1023_74#_c_821_n N_A_850_74#_c_1245_n 9.82309e-19 $X=5.535 $Y=1.575
+ $X2=0 $Y2=0
cc_697 N_A_1023_74#_c_828_n N_A_850_74#_c_1245_n 4.31798e-19 $X=5.535 $Y=1.045
+ $X2=0 $Y2=0
cc_698 N_A_1023_74#_c_821_n N_A_850_74#_c_1246_n 0.00138121f $X=5.535 $Y=1.575
+ $X2=0 $Y2=0
cc_699 N_A_1023_74#_c_822_n N_A_850_74#_c_1246_n 0.0097467f $X=5.62 $Y=1.74
+ $X2=0 $Y2=0
cc_700 N_A_1023_74#_c_828_n N_A_850_74#_c_1246_n 0.00772817f $X=5.535 $Y=1.045
+ $X2=0 $Y2=0
cc_701 N_A_1023_74#_c_821_n N_A_850_74#_c_1247_n 0.00548452f $X=5.535 $Y=1.575
+ $X2=0 $Y2=0
cc_702 N_A_1023_74#_c_822_n N_A_850_74#_c_1247_n 9.56646e-19 $X=5.62 $Y=1.74
+ $X2=0 $Y2=0
cc_703 N_A_1023_74#_c_828_n N_A_850_74#_c_1247_n 0.00143808f $X=5.535 $Y=1.045
+ $X2=0 $Y2=0
cc_704 N_A_1023_74#_c_833_n N_A_850_74#_c_1248_n 0.011534f $X=6.115 $Y=2.15
+ $X2=0 $Y2=0
cc_705 N_A_1023_74#_c_834_n N_A_850_74#_c_1248_n 0.0128825f $X=6.115 $Y=2.24
+ $X2=0 $Y2=0
cc_706 N_A_1023_74#_c_821_n N_A_850_74#_c_1248_n 0.0125279f $X=5.535 $Y=1.575
+ $X2=0 $Y2=0
cc_707 N_A_1023_74#_c_822_n N_A_850_74#_c_1248_n 0.0156362f $X=5.62 $Y=1.74
+ $X2=0 $Y2=0
cc_708 N_A_1023_74#_c_823_n N_A_850_74#_c_1248_n 0.00862606f $X=6.055 $Y=1.74
+ $X2=0 $Y2=0
cc_709 N_A_1023_74#_c_832_n N_A_850_74#_c_1248_n 0.0213783f $X=6.055 $Y=1.65
+ $X2=0 $Y2=0
cc_710 N_A_1023_74#_c_823_n N_A_850_74#_c_1249_n 0.00713715f $X=6.055 $Y=1.74
+ $X2=0 $Y2=0
cc_711 N_A_1023_74#_c_832_n N_A_850_74#_c_1249_n 0.0122266f $X=6.055 $Y=1.65
+ $X2=0 $Y2=0
cc_712 N_A_1023_74#_c_834_n N_A_850_74#_c_1262_n 0.010344f $X=6.115 $Y=2.24
+ $X2=0 $Y2=0
cc_713 N_A_1023_74#_M1004_g N_A_850_74#_M1012_g 0.0267822f $X=6.53 $Y=0.695
+ $X2=0 $Y2=0
cc_714 N_A_1023_74#_c_818_n N_A_850_74#_M1012_g 0.00361916f $X=5.255 $Y=0.515
+ $X2=0 $Y2=0
cc_715 N_A_1023_74#_c_819_n N_A_850_74#_M1012_g 0.00996885f $X=7.015 $Y=0.34
+ $X2=0 $Y2=0
cc_716 N_A_1023_74#_c_821_n N_A_850_74#_M1012_g 2.69793e-19 $X=5.535 $Y=1.575
+ $X2=0 $Y2=0
cc_717 N_A_1023_74#_c_828_n N_A_850_74#_M1012_g 9.21061e-19 $X=5.535 $Y=1.045
+ $X2=0 $Y2=0
cc_718 N_A_1023_74#_c_834_n N_A_850_74#_c_1264_n 0.00278823f $X=6.115 $Y=2.24
+ $X2=0 $Y2=0
cc_719 N_A_1023_74#_c_834_n N_A_850_74#_c_1266_n 0.0116365f $X=6.115 $Y=2.24
+ $X2=0 $Y2=0
cc_720 N_A_1023_74#_c_813_n N_A_850_74#_c_1266_n 0.0034104f $X=6.455 $Y=1.65
+ $X2=0 $Y2=0
cc_721 N_A_1023_74#_c_836_n N_A_850_74#_c_1268_n 0.00464206f $X=9.77 $Y=2.37
+ $X2=0 $Y2=0
cc_722 N_A_1023_74#_c_836_n N_A_850_74#_M1023_g 0.00689007f $X=9.77 $Y=2.37
+ $X2=0 $Y2=0
cc_723 N_A_1023_74#_c_839_n N_A_850_74#_M1023_g 0.00157762f $X=9.67 $Y=2.065
+ $X2=0 $Y2=0
cc_724 N_A_1023_74#_c_836_n N_A_850_74#_c_1251_n 0.0191375f $X=9.77 $Y=2.37
+ $X2=0 $Y2=0
cc_725 N_A_1023_74#_c_827_n N_A_850_74#_c_1251_n 3.3013e-19 $X=9.27 $Y=1.345
+ $X2=0 $Y2=0
cc_726 N_A_1023_74#_c_839_n N_A_850_74#_c_1251_n 0.00813875f $X=9.67 $Y=2.065
+ $X2=0 $Y2=0
cc_727 N_A_1023_74#_c_830_n N_A_850_74#_c_1251_n 0.0125871f $X=9.27 $Y=1.07
+ $X2=0 $Y2=0
cc_728 N_A_1023_74#_c_831_n N_A_850_74#_c_1251_n 0.0175647f $X=9.63 $Y=1.46
+ $X2=0 $Y2=0
cc_729 N_A_1023_74#_c_816_n N_A_850_74#_c_1252_n 0.0125871f $X=9.105 $Y=1.16
+ $X2=0 $Y2=0
cc_730 N_A_1023_74#_c_827_n N_A_850_74#_M1013_g 0.00266955f $X=9.27 $Y=1.345
+ $X2=0 $Y2=0
cc_731 N_A_1023_74#_c_830_n N_A_850_74#_M1013_g 0.0176907f $X=9.27 $Y=1.07 $X2=0
+ $Y2=0
cc_732 N_A_1023_74#_c_831_n N_A_850_74#_M1013_g 0.00700032f $X=9.63 $Y=1.46
+ $X2=0 $Y2=0
cc_733 N_A_1023_74#_c_821_n N_A_850_74#_c_1254_n 0.00666423f $X=5.535 $Y=1.575
+ $X2=0 $Y2=0
cc_734 N_A_1023_74#_c_822_n N_A_850_74#_c_1274_n 0.00792363f $X=5.62 $Y=1.74
+ $X2=0 $Y2=0
cc_735 N_A_1023_74#_c_821_n N_A_850_74#_c_1257_n 0.00528326f $X=5.535 $Y=1.575
+ $X2=0 $Y2=0
cc_736 N_A_1023_74#_c_828_n N_A_850_74#_c_1257_n 0.00449595f $X=5.535 $Y=1.045
+ $X2=0 $Y2=0
cc_737 N_A_1023_74#_c_822_n N_A_850_74#_c_1258_n 0.00711149f $X=5.62 $Y=1.74
+ $X2=0 $Y2=0
cc_738 N_A_1023_74#_c_822_n N_A_850_74#_c_1276_n 0.00234498f $X=5.62 $Y=1.74
+ $X2=0 $Y2=0
cc_739 N_A_1023_74#_c_821_n N_A_850_74#_c_1259_n 0.021083f $X=5.535 $Y=1.575
+ $X2=0 $Y2=0
cc_740 N_A_1023_74#_c_822_n N_A_850_74#_c_1259_n 0.0140089f $X=5.62 $Y=1.74
+ $X2=0 $Y2=0
cc_741 N_A_1023_74#_c_828_n N_A_850_74#_c_1259_n 0.00826703f $X=5.535 $Y=1.045
+ $X2=0 $Y2=0
cc_742 N_A_1023_74#_c_831_n N_A_2008_48#_M1005_g 2.03511e-19 $X=9.63 $Y=1.46
+ $X2=0 $Y2=0
cc_743 N_A_1023_74#_c_836_n N_A_2008_48#_c_1438_n 0.0294704f $X=9.77 $Y=2.37
+ $X2=0 $Y2=0
cc_744 N_A_1023_74#_c_839_n N_A_2008_48#_c_1438_n 0.0016211f $X=9.67 $Y=2.065
+ $X2=0 $Y2=0
cc_745 N_A_1023_74#_c_836_n N_A_2008_48#_c_1446_n 0.0336986f $X=9.77 $Y=2.37
+ $X2=0 $Y2=0
cc_746 N_A_1023_74#_c_825_n N_A_1747_74#_M1030_d 0.0019485f $X=8.78 $Y=0.34
+ $X2=-0.19 $Y2=-0.245
cc_747 N_A_1023_74#_c_944_p N_A_1747_74#_M1030_d 0.0100293f $X=8.865 $Y=0.905
+ $X2=-0.19 $Y2=-0.245
cc_748 N_A_1023_74#_c_829_n N_A_1747_74#_M1030_d 0.00256528f $X=9.27 $Y=1.07
+ $X2=-0.19 $Y2=-0.245
cc_749 N_A_1023_74#_c_836_n N_A_1747_74#_c_1609_n 0.00430249f $X=9.77 $Y=2.37
+ $X2=0 $Y2=0
cc_750 N_A_1023_74#_c_839_n N_A_1747_74#_c_1609_n 0.0330459f $X=9.67 $Y=2.065
+ $X2=0 $Y2=0
cc_751 N_A_1023_74#_c_831_n N_A_1747_74#_c_1609_n 0.0150349f $X=9.63 $Y=1.46
+ $X2=0 $Y2=0
cc_752 N_A_1023_74#_c_815_n N_A_1747_74#_c_1627_n 7.45707e-19 $X=8.66 $Y=1.085
+ $X2=0 $Y2=0
cc_753 N_A_1023_74#_c_825_n N_A_1747_74#_c_1627_n 0.00160036f $X=8.78 $Y=0.34
+ $X2=0 $Y2=0
cc_754 N_A_1023_74#_c_944_p N_A_1747_74#_c_1627_n 0.0234496f $X=8.865 $Y=0.905
+ $X2=0 $Y2=0
cc_755 N_A_1023_74#_c_829_n N_A_1747_74#_c_1627_n 0.0221981f $X=9.27 $Y=1.07
+ $X2=0 $Y2=0
cc_756 N_A_1023_74#_c_830_n N_A_1747_74#_c_1627_n 0.00683469f $X=9.27 $Y=1.07
+ $X2=0 $Y2=0
cc_757 N_A_1023_74#_c_831_n N_A_1747_74#_c_1627_n 0.00536065f $X=9.63 $Y=1.46
+ $X2=0 $Y2=0
cc_758 N_A_1023_74#_c_836_n N_A_1747_74#_c_1594_n 0.0159422f $X=9.77 $Y=2.37
+ $X2=0 $Y2=0
cc_759 N_A_1023_74#_c_839_n N_A_1747_74#_c_1594_n 0.0169381f $X=9.67 $Y=2.065
+ $X2=0 $Y2=0
cc_760 N_A_1023_74#_c_944_p N_A_1747_74#_c_1581_n 0.00463964f $X=8.865 $Y=0.905
+ $X2=0 $Y2=0
cc_761 N_A_1023_74#_c_829_n N_A_1747_74#_c_1581_n 0.00785017f $X=9.27 $Y=1.07
+ $X2=0 $Y2=0
cc_762 N_A_1023_74#_c_830_n N_A_1747_74#_c_1581_n 2.98286e-19 $X=9.27 $Y=1.07
+ $X2=0 $Y2=0
cc_763 N_A_1023_74#_c_836_n N_A_1747_74#_c_1582_n 0.00418565f $X=9.77 $Y=2.37
+ $X2=0 $Y2=0
cc_764 N_A_1023_74#_c_839_n N_A_1747_74#_c_1582_n 0.0483469f $X=9.67 $Y=2.065
+ $X2=0 $Y2=0
cc_765 N_A_1023_74#_c_831_n N_A_1747_74#_c_1582_n 0.0109876f $X=9.63 $Y=1.46
+ $X2=0 $Y2=0
cc_766 N_A_1023_74#_c_827_n N_A_1747_74#_c_1583_n 0.015348f $X=9.27 $Y=1.345
+ $X2=0 $Y2=0
cc_767 N_A_1023_74#_c_829_n N_A_1747_74#_c_1583_n 0.00613506f $X=9.27 $Y=1.07
+ $X2=0 $Y2=0
cc_768 N_A_1023_74#_c_830_n N_A_1747_74#_c_1583_n 0.00101813f $X=9.27 $Y=1.07
+ $X2=0 $Y2=0
cc_769 N_A_1023_74#_c_831_n N_A_1747_74#_c_1583_n 0.0202102f $X=9.63 $Y=1.46
+ $X2=0 $Y2=0
cc_770 N_A_1023_74#_c_836_n N_VPWR_c_1821_n 0.0038628f $X=9.77 $Y=2.37 $X2=0
+ $Y2=0
cc_771 N_A_1023_74#_c_834_n N_VPWR_c_1803_n 9.39239e-19 $X=6.115 $Y=2.24 $X2=0
+ $Y2=0
cc_772 N_A_1023_74#_c_836_n N_VPWR_c_1803_n 0.00515964f $X=9.77 $Y=2.37 $X2=0
+ $Y2=0
cc_773 N_A_1023_74#_M1038_d N_A_413_90#_c_1995_n 0.00696219f $X=5.17 $Y=1.82
+ $X2=0 $Y2=0
cc_774 N_A_1023_74#_c_822_n N_A_413_90#_c_1995_n 0.0232326f $X=5.62 $Y=1.74
+ $X2=0 $Y2=0
cc_775 N_A_1023_74#_c_823_n N_A_413_90#_c_1995_n 0.00177673f $X=6.055 $Y=1.74
+ $X2=0 $Y2=0
cc_776 N_A_1023_74#_M1004_g N_A_413_90#_c_1987_n 8.53322e-19 $X=6.53 $Y=0.695
+ $X2=0 $Y2=0
cc_777 N_A_1023_74#_c_818_n N_A_413_90#_c_1987_n 0.00725699f $X=5.255 $Y=0.515
+ $X2=0 $Y2=0
cc_778 N_A_1023_74#_c_828_n N_A_413_90#_c_1987_n 0.0100776f $X=5.535 $Y=1.045
+ $X2=0 $Y2=0
cc_779 N_A_1023_74#_c_833_n N_A_413_90#_c_1996_n 0.00517622f $X=6.115 $Y=2.15
+ $X2=0 $Y2=0
cc_780 N_A_1023_74#_c_834_n N_A_413_90#_c_1996_n 0.0101047f $X=6.115 $Y=2.24
+ $X2=0 $Y2=0
cc_781 N_A_1023_74#_c_813_n N_A_413_90#_c_1996_n 0.00272338f $X=6.455 $Y=1.65
+ $X2=0 $Y2=0
cc_782 N_A_1023_74#_c_823_n N_A_413_90#_c_1996_n 0.0118264f $X=6.055 $Y=1.74
+ $X2=0 $Y2=0
cc_783 N_A_1023_74#_c_832_n N_A_413_90#_c_1996_n 0.001604f $X=6.055 $Y=1.65
+ $X2=0 $Y2=0
cc_784 N_A_1023_74#_M1004_g N_A_413_90#_c_1988_n 0.00511004f $X=6.53 $Y=0.695
+ $X2=0 $Y2=0
cc_785 N_A_1023_74#_c_819_n N_A_413_90#_c_1988_n 0.00398151f $X=7.015 $Y=0.34
+ $X2=0 $Y2=0
cc_786 N_A_1023_74#_c_823_n N_A_413_90#_c_1988_n 0.00837959f $X=6.055 $Y=1.74
+ $X2=0 $Y2=0
cc_787 N_A_1023_74#_c_832_n N_A_413_90#_c_1988_n 0.00714825f $X=6.055 $Y=1.65
+ $X2=0 $Y2=0
cc_788 N_A_1023_74#_c_821_n N_A_413_90#_c_1989_n 0.00988314f $X=5.535 $Y=1.575
+ $X2=0 $Y2=0
cc_789 N_A_1023_74#_c_823_n N_A_413_90#_c_1989_n 0.00845438f $X=6.055 $Y=1.74
+ $X2=0 $Y2=0
cc_790 N_A_1023_74#_c_828_n N_A_413_90#_c_1989_n 0.00285927f $X=5.535 $Y=1.045
+ $X2=0 $Y2=0
cc_791 N_A_1023_74#_c_832_n N_A_413_90#_c_1989_n 2.97054e-19 $X=6.055 $Y=1.65
+ $X2=0 $Y2=0
cc_792 N_A_1023_74#_c_833_n N_A_413_90#_c_1990_n 0.00381322f $X=6.115 $Y=2.15
+ $X2=0 $Y2=0
cc_793 N_A_1023_74#_c_813_n N_A_413_90#_c_1990_n 0.0117688f $X=6.455 $Y=1.65
+ $X2=0 $Y2=0
cc_794 N_A_1023_74#_M1004_g N_A_413_90#_c_1990_n 0.00819144f $X=6.53 $Y=0.695
+ $X2=0 $Y2=0
cc_795 N_A_1023_74#_c_823_n N_A_413_90#_c_1990_n 0.0257264f $X=6.055 $Y=1.74
+ $X2=0 $Y2=0
cc_796 N_A_1023_74#_c_832_n N_A_413_90#_c_1990_n 0.00205131f $X=6.055 $Y=1.65
+ $X2=0 $Y2=0
cc_797 N_A_1023_74#_c_818_n N_A_413_90#_c_1992_n 0.0127884f $X=5.255 $Y=0.515
+ $X2=0 $Y2=0
cc_798 N_A_1023_74#_c_819_n N_A_413_90#_c_1992_n 0.0211967f $X=7.015 $Y=0.34
+ $X2=0 $Y2=0
cc_799 N_A_1023_74#_c_834_n N_A_413_90#_c_2000_n 0.0058235f $X=6.115 $Y=2.24
+ $X2=0 $Y2=0
cc_800 N_A_1023_74#_c_822_n N_A_413_90#_c_2000_n 0.00397178f $X=5.62 $Y=1.74
+ $X2=0 $Y2=0
cc_801 N_A_1023_74#_c_823_n N_A_413_90#_c_2000_n 0.0135052f $X=6.055 $Y=1.74
+ $X2=0 $Y2=0
cc_802 N_A_1023_74#_c_832_n N_A_413_90#_c_2000_n 0.0018949f $X=6.055 $Y=1.65
+ $X2=0 $Y2=0
cc_803 N_A_1023_74#_c_848_n N_VGND_M1017_d 0.0173515f $X=7.94 $Y=0.68 $X2=0
+ $Y2=0
cc_804 N_A_1023_74#_c_850_n N_VGND_M1017_d 0.00302969f $X=8.025 $Y=0.595 $X2=0
+ $Y2=0
cc_805 N_A_1023_74#_c_826_n N_VGND_M1017_d 6.57704e-19 $X=8.11 $Y=0.34 $X2=0
+ $Y2=0
cc_806 N_A_1023_74#_c_820_n N_VGND_c_2176_n 0.0112234f $X=5.42 $Y=0.34 $X2=0
+ $Y2=0
cc_807 N_A_1023_74#_c_819_n N_VGND_c_2177_n 0.0113147f $X=7.015 $Y=0.34 $X2=0
+ $Y2=0
cc_808 N_A_1023_74#_c_848_n N_VGND_c_2177_n 0.0246763f $X=7.94 $Y=0.68 $X2=0
+ $Y2=0
cc_809 N_A_1023_74#_c_826_n N_VGND_c_2177_n 0.0148568f $X=8.11 $Y=0.34 $X2=0
+ $Y2=0
cc_810 N_A_1023_74#_M1004_g N_VGND_c_2186_n 7.35405e-19 $X=6.53 $Y=0.695 $X2=0
+ $Y2=0
cc_811 N_A_1023_74#_c_819_n N_VGND_c_2186_n 0.114615f $X=7.015 $Y=0.34 $X2=0
+ $Y2=0
cc_812 N_A_1023_74#_c_820_n N_VGND_c_2186_n 0.0179706f $X=5.42 $Y=0.34 $X2=0
+ $Y2=0
cc_813 N_A_1023_74#_c_848_n N_VGND_c_2186_n 0.0038254f $X=7.94 $Y=0.68 $X2=0
+ $Y2=0
cc_814 N_A_1023_74#_c_815_n N_VGND_c_2187_n 0.00278271f $X=8.66 $Y=1.085 $X2=0
+ $Y2=0
cc_815 N_A_1023_74#_c_848_n N_VGND_c_2187_n 0.00323133f $X=7.94 $Y=0.68 $X2=0
+ $Y2=0
cc_816 N_A_1023_74#_c_825_n N_VGND_c_2187_n 0.0543743f $X=8.78 $Y=0.34 $X2=0
+ $Y2=0
cc_817 N_A_1023_74#_c_826_n N_VGND_c_2187_n 0.0119262f $X=8.11 $Y=0.34 $X2=0
+ $Y2=0
cc_818 N_A_1023_74#_c_815_n N_VGND_c_2190_n 0.00358525f $X=8.66 $Y=1.085 $X2=0
+ $Y2=0
cc_819 N_A_1023_74#_c_819_n N_VGND_c_2190_n 0.0665208f $X=7.015 $Y=0.34 $X2=0
+ $Y2=0
cc_820 N_A_1023_74#_c_820_n N_VGND_c_2190_n 0.00972865f $X=5.42 $Y=0.34 $X2=0
+ $Y2=0
cc_821 N_A_1023_74#_c_848_n N_VGND_c_2190_n 0.0140279f $X=7.94 $Y=0.68 $X2=0
+ $Y2=0
cc_822 N_A_1023_74#_c_825_n N_VGND_c_2190_n 0.0304188f $X=8.78 $Y=0.34 $X2=0
+ $Y2=0
cc_823 N_A_1023_74#_c_826_n N_VGND_c_2190_n 0.00656035f $X=8.11 $Y=0.34 $X2=0
+ $Y2=0
cc_824 N_A_1023_74#_c_863_p A_1399_97# 0.00130995f $X=7.185 $Y=0.68 $X2=-0.19
+ $Y2=-0.245
cc_825 N_A_1369_71#_c_1025_n N_A_1221_97#_M1041_g 0.01067f $X=8.28 $Y=1.02 $X2=0
+ $Y2=0
cc_826 N_A_1369_71#_c_1068_n N_A_1221_97#_M1041_g 0.00970467f $X=8.445 $Y=0.81
+ $X2=0 $Y2=0
cc_827 N_A_1369_71#_c_1027_n N_A_1221_97#_M1041_g 0.0031265f $X=8.525 $Y=1.245
+ $X2=0 $Y2=0
cc_828 N_A_1369_71#_c_1030_n N_A_1221_97#_M1041_g 0.0021525f $X=8.445 $Y=1.02
+ $X2=0 $Y2=0
cc_829 N_A_1369_71#_c_1029_n N_A_1221_97#_c_1137_n 0.00507431f $X=8.77 $Y=1.88
+ $X2=0 $Y2=0
cc_830 N_A_1369_71#_M1016_g N_A_1221_97#_c_1131_n 0.00671859f $X=6.92 $Y=0.695
+ $X2=0 $Y2=0
cc_831 N_A_1369_71#_M1016_g N_A_1221_97#_c_1132_n 0.00680947f $X=6.92 $Y=0.695
+ $X2=0 $Y2=0
cc_832 N_A_1369_71#_c_1031_n N_A_1221_97#_c_1132_n 0.00782496f $X=6.955 $Y=2.15
+ $X2=0 $Y2=0
cc_833 N_A_1369_71#_c_1032_n N_A_1221_97#_c_1132_n 8.9565e-19 $X=6.955 $Y=2.24
+ $X2=0 $Y2=0
cc_834 N_A_1369_71#_c_1023_n N_A_1221_97#_c_1132_n 0.0489555f $X=7.125 $Y=1.595
+ $X2=0 $Y2=0
cc_835 N_A_1369_71#_c_1026_n N_A_1221_97#_c_1132_n 0.0143478f $X=7.235 $Y=1.02
+ $X2=0 $Y2=0
cc_836 N_A_1369_71#_c_1032_n N_A_1221_97#_c_1148_n 0.0106967f $X=6.955 $Y=2.24
+ $X2=0 $Y2=0
cc_837 N_A_1369_71#_c_1023_n N_A_1221_97#_c_1148_n 0.00241061f $X=7.125 $Y=1.595
+ $X2=0 $Y2=0
cc_838 N_A_1369_71#_c_1024_n N_A_1221_97#_c_1148_n 0.00225416f $X=7.125 $Y=1.595
+ $X2=0 $Y2=0
cc_839 N_A_1369_71#_c_1031_n N_A_1221_97#_c_1133_n 0.00354747f $X=6.955 $Y=2.15
+ $X2=0 $Y2=0
cc_840 N_A_1369_71#_c_1032_n N_A_1221_97#_c_1133_n 0.00138556f $X=6.955 $Y=2.24
+ $X2=0 $Y2=0
cc_841 N_A_1369_71#_c_1023_n N_A_1221_97#_c_1133_n 0.0156336f $X=7.125 $Y=1.595
+ $X2=0 $Y2=0
cc_842 N_A_1369_71#_c_1024_n N_A_1221_97#_c_1133_n 0.00141843f $X=7.125 $Y=1.595
+ $X2=0 $Y2=0
cc_843 N_A_1369_71#_c_1023_n N_A_1221_97#_c_1134_n 0.0227604f $X=7.125 $Y=1.595
+ $X2=0 $Y2=0
cc_844 N_A_1369_71#_c_1024_n N_A_1221_97#_c_1134_n 8.70669e-19 $X=7.125 $Y=1.595
+ $X2=0 $Y2=0
cc_845 N_A_1369_71#_c_1025_n N_A_1221_97#_c_1134_n 0.0135118f $X=8.28 $Y=1.02
+ $X2=0 $Y2=0
cc_846 N_A_1369_71#_c_1025_n N_A_1221_97#_c_1135_n 0.0516286f $X=8.28 $Y=1.02
+ $X2=0 $Y2=0
cc_847 N_A_1369_71#_c_1028_n N_A_1221_97#_c_1135_n 0.0120015f $X=8.81 $Y=1.415
+ $X2=0 $Y2=0
cc_848 N_A_1369_71#_c_1029_n N_A_1221_97#_c_1135_n 0.00540759f $X=8.77 $Y=1.88
+ $X2=0 $Y2=0
cc_849 N_A_1369_71#_c_1032_n N_A_1221_97#_c_1141_n 0.00112114f $X=6.955 $Y=2.24
+ $X2=0 $Y2=0
cc_850 N_A_1369_71#_c_1025_n N_A_1221_97#_c_1136_n 0.00505406f $X=8.28 $Y=1.02
+ $X2=0 $Y2=0
cc_851 N_A_1369_71#_c_1028_n N_A_1221_97#_c_1136_n 0.012066f $X=8.81 $Y=1.415
+ $X2=0 $Y2=0
cc_852 N_A_1369_71#_c_1029_n N_A_1221_97#_c_1136_n 0.00632508f $X=8.77 $Y=1.88
+ $X2=0 $Y2=0
cc_853 N_A_1369_71#_c_1030_n N_A_1221_97#_c_1136_n 0.00275569f $X=8.445 $Y=1.02
+ $X2=0 $Y2=0
cc_854 N_A_1369_71#_c_1032_n N_A_850_74#_c_1264_n 0.00322812f $X=6.955 $Y=2.24
+ $X2=0 $Y2=0
cc_855 N_A_1369_71#_c_1032_n N_A_850_74#_c_1266_n 0.0307484f $X=6.955 $Y=2.24
+ $X2=0 $Y2=0
cc_856 N_A_1369_71#_c_1032_n N_A_850_74#_c_1267_n 0.0100502f $X=6.955 $Y=2.24
+ $X2=0 $Y2=0
cc_857 N_A_1369_71#_c_1029_n N_A_850_74#_c_1267_n 0.00262042f $X=8.77 $Y=1.88
+ $X2=0 $Y2=0
cc_858 N_A_1369_71#_c_1029_n N_A_850_74#_c_1268_n 5.08057e-19 $X=8.77 $Y=1.88
+ $X2=0 $Y2=0
cc_859 N_A_1369_71#_c_1029_n N_A_850_74#_M1023_g 0.0124176f $X=8.77 $Y=1.88
+ $X2=0 $Y2=0
cc_860 N_A_1369_71#_c_1029_n N_A_850_74#_c_1252_n 0.00543498f $X=8.77 $Y=1.88
+ $X2=0 $Y2=0
cc_861 N_A_1369_71#_c_1029_n N_A_1747_74#_c_1609_n 0.0261048f $X=8.77 $Y=1.88
+ $X2=0 $Y2=0
cc_862 N_A_1369_71#_c_1029_n N_A_1747_74#_c_1595_n 0.0128087f $X=8.77 $Y=1.88
+ $X2=0 $Y2=0
cc_863 N_A_1369_71#_c_1032_n N_VPWR_c_1807_n 0.00420497f $X=6.955 $Y=2.24 $X2=0
+ $Y2=0
cc_864 N_A_1369_71#_c_1025_n N_VPWR_c_1808_n 2.9437e-19 $X=8.28 $Y=1.02 $X2=0
+ $Y2=0
cc_865 N_A_1369_71#_c_1028_n N_VPWR_c_1808_n 0.00220892f $X=8.81 $Y=1.415 $X2=0
+ $Y2=0
cc_866 N_A_1369_71#_c_1029_n N_VPWR_c_1808_n 0.0670793f $X=8.77 $Y=1.88 $X2=0
+ $Y2=0
cc_867 N_A_1369_71#_c_1030_n N_VPWR_c_1808_n 0.00582847f $X=8.445 $Y=1.02 $X2=0
+ $Y2=0
cc_868 N_A_1369_71#_c_1029_n N_VPWR_c_1821_n 0.00567879f $X=8.77 $Y=1.88 $X2=0
+ $Y2=0
cc_869 N_A_1369_71#_c_1032_n N_VPWR_c_1803_n 9.39239e-19 $X=6.955 $Y=2.24 $X2=0
+ $Y2=0
cc_870 N_A_1369_71#_c_1029_n N_VPWR_c_1803_n 0.00684413f $X=8.77 $Y=1.88 $X2=0
+ $Y2=0
cc_871 N_A_1369_71#_c_1025_n N_VGND_M1017_d 0.00233925f $X=8.28 $Y=1.02 $X2=0
+ $Y2=0
cc_872 N_A_1369_71#_M1016_g N_VGND_c_2186_n 7.35405e-19 $X=6.92 $Y=0.695 $X2=0
+ $Y2=0
cc_873 N_A_1221_97#_c_1138_n N_A_850_74#_c_1262_n 0.00381872f $X=6.675 $Y=2.585
+ $X2=0 $Y2=0
cc_874 N_A_1221_97#_c_1131_n N_A_850_74#_M1012_g 0.00178378f $X=6.675 $Y=0.76
+ $X2=0 $Y2=0
cc_875 N_A_1221_97#_c_1138_n N_A_850_74#_c_1264_n 9.692e-19 $X=6.675 $Y=2.585
+ $X2=0 $Y2=0
cc_876 N_A_1221_97#_c_1138_n N_A_850_74#_c_1266_n 0.0125516f $X=6.675 $Y=2.585
+ $X2=0 $Y2=0
cc_877 N_A_1221_97#_c_1132_n N_A_850_74#_c_1266_n 0.00206435f $X=6.76 $Y=2.32
+ $X2=0 $Y2=0
cc_878 N_A_1221_97#_c_1137_n N_A_850_74#_c_1267_n 0.0103562f $X=8.545 $Y=1.66
+ $X2=0 $Y2=0
cc_879 N_A_1221_97#_c_1148_n N_A_850_74#_c_1267_n 0.00215266f $X=7.405 $Y=2.405
+ $X2=0 $Y2=0
cc_880 N_A_1221_97#_c_1133_n N_A_850_74#_c_1267_n 0.00744895f $X=7.49 $Y=2.32
+ $X2=0 $Y2=0
cc_881 N_A_1221_97#_c_1141_n N_A_850_74#_c_1267_n 0.00202544f $X=6.76 $Y=2.537
+ $X2=0 $Y2=0
cc_882 N_A_1221_97#_c_1137_n N_A_850_74#_c_1268_n 0.00249951f $X=8.545 $Y=1.66
+ $X2=0 $Y2=0
cc_883 N_A_1221_97#_c_1137_n N_A_850_74#_M1023_g 0.00575058f $X=8.545 $Y=1.66
+ $X2=0 $Y2=0
cc_884 N_A_1221_97#_c_1136_n N_A_850_74#_c_1252_n 0.0067924f $X=8.23 $Y=1.452
+ $X2=0 $Y2=0
cc_885 N_A_1221_97#_c_1148_n N_VPWR_M1018_d 0.00766967f $X=7.405 $Y=2.405 $X2=0
+ $Y2=0
cc_886 N_A_1221_97#_c_1148_n N_VPWR_c_1807_n 0.0241478f $X=7.405 $Y=2.405 $X2=0
+ $Y2=0
cc_887 N_A_1221_97#_c_1133_n N_VPWR_c_1807_n 0.00784846f $X=7.49 $Y=2.32 $X2=0
+ $Y2=0
cc_888 N_A_1221_97#_c_1141_n N_VPWR_c_1807_n 0.00363331f $X=6.76 $Y=2.537 $X2=0
+ $Y2=0
cc_889 N_A_1221_97#_c_1137_n N_VPWR_c_1808_n 0.0151329f $X=8.545 $Y=1.66 $X2=0
+ $Y2=0
cc_890 N_A_1221_97#_c_1133_n N_VPWR_c_1808_n 0.0313215f $X=7.49 $Y=2.32 $X2=0
+ $Y2=0
cc_891 N_A_1221_97#_c_1135_n N_VPWR_c_1808_n 0.00271335f $X=8.105 $Y=1.41 $X2=0
+ $Y2=0
cc_892 N_A_1221_97#_c_1136_n N_VPWR_c_1808_n 0.00677043f $X=8.23 $Y=1.452 $X2=0
+ $Y2=0
cc_893 N_A_1221_97#_c_1138_n N_VPWR_c_1816_n 0.0105518f $X=6.675 $Y=2.585 $X2=0
+ $Y2=0
cc_894 N_A_1221_97#_c_1141_n N_VPWR_c_1816_n 0.00389335f $X=6.76 $Y=2.537 $X2=0
+ $Y2=0
cc_895 N_A_1221_97#_c_1133_n N_VPWR_c_1820_n 0.00731736f $X=7.49 $Y=2.32 $X2=0
+ $Y2=0
cc_896 N_A_1221_97#_c_1137_n N_VPWR_c_1803_n 8.51577e-19 $X=8.545 $Y=1.66 $X2=0
+ $Y2=0
cc_897 N_A_1221_97#_c_1138_n N_VPWR_c_1803_n 0.0131649f $X=6.675 $Y=2.585 $X2=0
+ $Y2=0
cc_898 N_A_1221_97#_c_1148_n N_VPWR_c_1803_n 0.00805206f $X=7.405 $Y=2.405 $X2=0
+ $Y2=0
cc_899 N_A_1221_97#_c_1133_n N_VPWR_c_1803_n 0.0152718f $X=7.49 $Y=2.32 $X2=0
+ $Y2=0
cc_900 N_A_1221_97#_c_1141_n N_VPWR_c_1803_n 0.00470184f $X=6.76 $Y=2.537 $X2=0
+ $Y2=0
cc_901 N_A_1221_97#_c_1131_n N_A_413_90#_c_1987_n 0.00540476f $X=6.675 $Y=0.76
+ $X2=0 $Y2=0
cc_902 N_A_1221_97#_c_1138_n N_A_413_90#_c_1996_n 0.0212263f $X=6.675 $Y=2.585
+ $X2=0 $Y2=0
cc_903 N_A_1221_97#_c_1132_n N_A_413_90#_c_1996_n 0.0137556f $X=6.76 $Y=2.32
+ $X2=0 $Y2=0
cc_904 N_A_1221_97#_c_1131_n N_A_413_90#_c_1988_n 0.0292368f $X=6.675 $Y=0.76
+ $X2=0 $Y2=0
cc_905 N_A_1221_97#_c_1132_n N_A_413_90#_c_1988_n 0.013608f $X=6.76 $Y=2.32
+ $X2=0 $Y2=0
cc_906 N_A_1221_97#_c_1132_n N_A_413_90#_c_1990_n 0.0586249f $X=6.76 $Y=2.32
+ $X2=0 $Y2=0
cc_907 N_A_1221_97#_c_1138_n N_A_413_90#_c_2000_n 0.0247482f $X=6.675 $Y=2.585
+ $X2=0 $Y2=0
cc_908 N_A_1221_97#_M1041_g N_VGND_c_2177_n 0.00117551f $X=8.23 $Y=0.69 $X2=0
+ $Y2=0
cc_909 N_A_1221_97#_M1041_g N_VGND_c_2187_n 0.00278271f $X=8.23 $Y=0.69 $X2=0
+ $Y2=0
cc_910 N_A_1221_97#_M1041_g N_VGND_c_2190_n 0.00358525f $X=8.23 $Y=0.69 $X2=0
+ $Y2=0
cc_911 N_A_1221_97#_c_1131_n A_1321_97# 0.00136908f $X=6.675 $Y=0.76 $X2=-0.19
+ $Y2=-0.245
cc_912 N_A_850_74#_M1013_g N_A_2008_48#_M1005_g 0.0422064f $X=9.755 $Y=0.58
+ $X2=0 $Y2=0
cc_913 N_A_850_74#_c_1251_n N_A_2008_48#_c_1438_n 0.0427595f $X=9.68 $Y=1.585
+ $X2=0 $Y2=0
cc_914 N_A_850_74#_M1023_g N_A_1747_74#_c_1609_n 2.44304e-19 $X=8.995 $Y=2.235
+ $X2=0 $Y2=0
cc_915 N_A_850_74#_c_1251_n N_A_1747_74#_c_1609_n 0.00473791f $X=9.68 $Y=1.585
+ $X2=0 $Y2=0
cc_916 N_A_850_74#_M1013_g N_A_1747_74#_c_1627_n 0.0150881f $X=9.755 $Y=0.58
+ $X2=0 $Y2=0
cc_917 N_A_850_74#_M1023_g N_A_1747_74#_c_1595_n 0.00211239f $X=8.995 $Y=2.235
+ $X2=0 $Y2=0
cc_918 N_A_850_74#_M1013_g N_A_1747_74#_c_1581_n 0.00884302f $X=9.755 $Y=0.58
+ $X2=0 $Y2=0
cc_919 N_A_850_74#_M1013_g N_A_1747_74#_c_1582_n 0.0014557f $X=9.755 $Y=0.58
+ $X2=0 $Y2=0
cc_920 N_A_850_74#_c_1251_n N_A_1747_74#_c_1583_n 4.03784e-19 $X=9.68 $Y=1.585
+ $X2=0 $Y2=0
cc_921 N_A_850_74#_M1013_g N_A_1747_74#_c_1583_n 0.0141061f $X=9.755 $Y=0.58
+ $X2=0 $Y2=0
cc_922 N_A_850_74#_c_1274_n N_VPWR_M1025_d 0.00226298f $X=4.815 $Y=1.885 $X2=0
+ $Y2=0
cc_923 N_A_850_74#_c_1246_n N_VPWR_c_1806_n 0.00919622f $X=5.095 $Y=1.745 $X2=0
+ $Y2=0
cc_924 N_A_850_74#_c_1248_n N_VPWR_c_1806_n 0.00475591f $X=5.605 $Y=3.075 $X2=0
+ $Y2=0
cc_925 N_A_850_74#_c_1264_n N_VPWR_c_1807_n 0.00607321f $X=6.565 $Y=2.9 $X2=0
+ $Y2=0
cc_926 N_A_850_74#_c_1267_n N_VPWR_c_1807_n 0.0253641f $X=8.905 $Y=3.15 $X2=0
+ $Y2=0
cc_927 N_A_850_74#_c_1267_n N_VPWR_c_1808_n 0.0213056f $X=8.905 $Y=3.15 $X2=0
+ $Y2=0
cc_928 N_A_850_74#_c_1268_n N_VPWR_c_1808_n 0.00613773f $X=8.995 $Y=2.9 $X2=0
+ $Y2=0
cc_929 N_A_850_74#_M1023_g N_VPWR_c_1808_n 6.49178e-19 $X=8.995 $Y=2.235 $X2=0
+ $Y2=0
cc_930 N_A_850_74#_c_1246_n N_VPWR_c_1816_n 0.00505726f $X=5.095 $Y=1.745 $X2=0
+ $Y2=0
cc_931 N_A_850_74#_c_1263_n N_VPWR_c_1816_n 0.0467845f $X=5.68 $Y=3.15 $X2=0
+ $Y2=0
cc_932 N_A_850_74#_c_1267_n N_VPWR_c_1820_n 0.0250026f $X=8.905 $Y=3.15 $X2=0
+ $Y2=0
cc_933 N_A_850_74#_c_1267_n N_VPWR_c_1821_n 0.0193014f $X=8.905 $Y=3.15 $X2=0
+ $Y2=0
cc_934 N_A_850_74#_c_1246_n N_VPWR_c_1803_n 0.00489105f $X=5.095 $Y=1.745 $X2=0
+ $Y2=0
cc_935 N_A_850_74#_c_1262_n N_VPWR_c_1803_n 0.0238273f $X=6.475 $Y=3.15 $X2=0
+ $Y2=0
cc_936 N_A_850_74#_c_1263_n N_VPWR_c_1803_n 0.0070819f $X=5.68 $Y=3.15 $X2=0
+ $Y2=0
cc_937 N_A_850_74#_c_1267_n N_VPWR_c_1803_n 0.0676231f $X=8.905 $Y=3.15 $X2=0
+ $Y2=0
cc_938 N_A_850_74#_c_1273_n N_VPWR_c_1803_n 0.00495695f $X=6.565 $Y=3.15 $X2=0
+ $Y2=0
cc_939 N_A_850_74#_c_1255_n N_A_413_90#_c_1985_n 0.00301448f $X=4.355 $Y=0.84
+ $X2=0 $Y2=0
cc_940 N_A_850_74#_M1025_s N_A_413_90#_c_1995_n 0.0083322f $X=4.275 $Y=1.82
+ $X2=0 $Y2=0
cc_941 N_A_850_74#_c_1246_n N_A_413_90#_c_1995_n 0.0126314f $X=5.095 $Y=1.745
+ $X2=0 $Y2=0
cc_942 N_A_850_74#_c_1248_n N_A_413_90#_c_1995_n 0.0130181f $X=5.605 $Y=3.075
+ $X2=0 $Y2=0
cc_943 N_A_850_74#_c_1274_n N_A_413_90#_c_1995_n 0.00842051f $X=4.815 $Y=1.885
+ $X2=0 $Y2=0
cc_944 N_A_850_74#_c_1276_n N_A_413_90#_c_1995_n 0.0136272f $X=4.46 $Y=1.885
+ $X2=0 $Y2=0
cc_945 N_A_850_74#_M1012_g N_A_413_90#_c_1987_n 0.00810667f $X=6.03 $Y=0.695
+ $X2=0 $Y2=0
cc_946 N_A_850_74#_c_1266_n N_A_413_90#_c_1996_n 0.00175546f $X=6.565 $Y=2.81
+ $X2=0 $Y2=0
cc_947 N_A_850_74#_c_1249_n N_A_413_90#_c_1988_n 0.00322497f $X=5.955 $Y=1.26
+ $X2=0 $Y2=0
cc_948 N_A_850_74#_M1012_g N_A_413_90#_c_1988_n 0.00583375f $X=6.03 $Y=0.695
+ $X2=0 $Y2=0
cc_949 N_A_850_74#_c_1249_n N_A_413_90#_c_1989_n 0.00532557f $X=5.955 $Y=1.26
+ $X2=0 $Y2=0
cc_950 N_A_850_74#_M1012_g N_A_413_90#_c_1989_n 0.00172798f $X=6.03 $Y=0.695
+ $X2=0 $Y2=0
cc_951 N_A_850_74#_c_1248_n N_A_413_90#_c_1990_n 0.00316493f $X=5.605 $Y=3.075
+ $X2=0 $Y2=0
cc_952 N_A_850_74#_c_1249_n N_A_413_90#_c_1990_n 0.00148483f $X=5.955 $Y=1.26
+ $X2=0 $Y2=0
cc_953 N_A_850_74#_M1012_g N_A_413_90#_c_1992_n 0.00243646f $X=6.03 $Y=0.695
+ $X2=0 $Y2=0
cc_954 N_A_850_74#_c_1254_n N_A_413_90#_c_1992_n 0.00454513f $X=5.605 $Y=1.26
+ $X2=0 $Y2=0
cc_955 N_A_850_74#_c_1248_n N_A_413_90#_c_2000_n 0.0127799f $X=5.605 $Y=3.075
+ $X2=0 $Y2=0
cc_956 N_A_850_74#_c_1262_n N_A_413_90#_c_2000_n 0.00413072f $X=6.475 $Y=3.15
+ $X2=0 $Y2=0
cc_957 N_A_850_74#_c_1299_n N_VGND_M1035_d 0.00449457f $X=4.815 $Y=0.925 $X2=0
+ $Y2=0
cc_958 N_A_850_74#_c_1257_n N_VGND_M1035_d 0.00112082f $X=4.9 $Y=1.3 $X2=0 $Y2=0
cc_959 N_A_850_74#_c_1256_n N_VGND_c_2175_n 0.0264125f $X=4.395 $Y=0.515 $X2=0
+ $Y2=0
cc_960 N_A_850_74#_c_1245_n N_VGND_c_2176_n 0.00734828f $X=5.04 $Y=1.185 $X2=0
+ $Y2=0
cc_961 N_A_850_74#_c_1256_n N_VGND_c_2176_n 0.0121972f $X=4.395 $Y=0.515 $X2=0
+ $Y2=0
cc_962 N_A_850_74#_c_1299_n N_VGND_c_2176_n 0.0170468f $X=4.815 $Y=0.925 $X2=0
+ $Y2=0
cc_963 N_A_850_74#_M1013_g N_VGND_c_2178_n 0.00177088f $X=9.755 $Y=0.58 $X2=0
+ $Y2=0
cc_964 N_A_850_74#_c_1256_n N_VGND_c_2183_n 0.0110419f $X=4.395 $Y=0.515 $X2=0
+ $Y2=0
cc_965 N_A_850_74#_c_1245_n N_VGND_c_2186_n 0.00383152f $X=5.04 $Y=1.185 $X2=0
+ $Y2=0
cc_966 N_A_850_74#_M1012_g N_VGND_c_2186_n 7.35405e-19 $X=6.03 $Y=0.695 $X2=0
+ $Y2=0
cc_967 N_A_850_74#_M1013_g N_VGND_c_2187_n 0.00358451f $X=9.755 $Y=0.58 $X2=0
+ $Y2=0
cc_968 N_A_850_74#_c_1245_n N_VGND_c_2190_n 0.00762539f $X=5.04 $Y=1.185 $X2=0
+ $Y2=0
cc_969 N_A_850_74#_M1013_g N_VGND_c_2190_n 0.00569641f $X=9.755 $Y=0.58 $X2=0
+ $Y2=0
cc_970 N_A_850_74#_c_1256_n N_VGND_c_2190_n 0.00915013f $X=4.395 $Y=0.515 $X2=0
+ $Y2=0
cc_971 N_A_850_74#_c_1299_n N_VGND_c_2190_n 0.00638302f $X=4.815 $Y=0.925 $X2=0
+ $Y2=0
cc_972 N_A_2008_48#_c_1442_n N_A_1747_74#_c_1573_n 0.0023753f $X=11.76 $Y=1.63
+ $X2=0 $Y2=0
cc_973 N_A_2008_48#_c_1443_n N_A_1747_74#_c_1573_n 0.00741302f $X=11.12 $Y=0.55
+ $X2=0 $Y2=0
cc_974 N_A_2008_48#_c_1440_n N_A_1747_74#_c_1574_n 0.00406259f $X=11.675
+ $Y=0.665 $X2=0 $Y2=0
cc_975 N_A_2008_48#_c_1442_n N_A_1747_74#_c_1574_n 0.00385495f $X=11.76 $Y=1.63
+ $X2=0 $Y2=0
cc_976 N_A_2008_48#_c_1443_n N_A_1747_74#_c_1574_n 0.00768727f $X=11.12 $Y=0.55
+ $X2=0 $Y2=0
cc_977 N_A_2008_48#_c_1450_n N_A_1747_74#_c_1585_n 0.00562099f $X=11.02 $Y=2.655
+ $X2=0 $Y2=0
cc_978 N_A_2008_48#_c_1454_n N_A_1747_74#_c_1585_n 0.00739298f $X=11.13 $Y=2.405
+ $X2=0 $Y2=0
cc_979 N_A_2008_48#_c_1451_n N_A_1747_74#_c_1586_n 0.0105765f $X=11.32 $Y=2.32
+ $X2=0 $Y2=0
cc_980 N_A_2008_48#_c_1452_n N_A_1747_74#_c_1586_n 0.00277596f $X=11.675
+ $Y=1.715 $X2=0 $Y2=0
cc_981 N_A_2008_48#_c_1441_n N_A_1747_74#_c_1586_n 0.00167941f $X=11.405
+ $Y=1.715 $X2=0 $Y2=0
cc_982 N_A_2008_48#_c_1451_n N_A_1747_74#_c_1587_n 6.41559e-19 $X=11.32 $Y=2.32
+ $X2=0 $Y2=0
cc_983 N_A_2008_48#_c_1452_n N_A_1747_74#_c_1587_n 3.71546e-19 $X=11.675
+ $Y=1.715 $X2=0 $Y2=0
cc_984 N_A_2008_48#_c_1442_n N_A_1747_74#_c_1576_n 0.00507794f $X=11.76 $Y=1.63
+ $X2=0 $Y2=0
cc_985 N_A_2008_48#_c_1443_n N_A_1747_74#_c_1576_n 0.00413357f $X=11.12 $Y=0.55
+ $X2=0 $Y2=0
cc_986 N_A_2008_48#_c_1440_n N_A_1747_74#_c_1578_n 0.00447579f $X=11.675
+ $Y=0.665 $X2=0 $Y2=0
cc_987 N_A_2008_48#_c_1452_n N_A_1747_74#_c_1578_n 0.0228154f $X=11.675 $Y=1.715
+ $X2=0 $Y2=0
cc_988 N_A_2008_48#_c_1441_n N_A_1747_74#_c_1578_n 0.00406088f $X=11.405
+ $Y=1.715 $X2=0 $Y2=0
cc_989 N_A_2008_48#_c_1442_n N_A_1747_74#_c_1578_n 0.0258377f $X=11.76 $Y=1.63
+ $X2=0 $Y2=0
cc_990 N_A_2008_48#_c_1451_n N_A_1747_74#_c_1592_n 0.00434917f $X=11.32 $Y=2.32
+ $X2=0 $Y2=0
cc_991 N_A_2008_48#_c_1454_n N_A_1747_74#_c_1592_n 0.00686891f $X=11.13 $Y=2.405
+ $X2=0 $Y2=0
cc_992 N_A_2008_48#_M1005_g N_A_1747_74#_c_1627_n 0.00100268f $X=10.115 $Y=0.58
+ $X2=0 $Y2=0
cc_993 N_A_2008_48#_c_1446_n N_A_1747_74#_c_1594_n 0.00888546f $X=10.16 $Y=2.37
+ $X2=0 $Y2=0
cc_994 N_A_2008_48#_c_1449_n N_A_1747_74#_c_1594_n 0.00364065f $X=10.525
+ $Y=2.405 $X2=0 $Y2=0
cc_995 N_A_2008_48#_M1005_g N_A_1747_74#_c_1581_n 0.00151652f $X=10.115 $Y=0.58
+ $X2=0 $Y2=0
cc_996 N_A_2008_48#_M1005_g N_A_1747_74#_c_1582_n 0.00175137f $X=10.115 $Y=0.58
+ $X2=0 $Y2=0
cc_997 N_A_2008_48#_c_1438_n N_A_1747_74#_c_1582_n 0.0146343f $X=10.16 $Y=1.98
+ $X2=0 $Y2=0
cc_998 N_A_2008_48#_c_1445_n N_A_1747_74#_c_1582_n 0.0045792f $X=10.16 $Y=2.28
+ $X2=0 $Y2=0
cc_999 N_A_2008_48#_c_1446_n N_A_1747_74#_c_1582_n 0.00266565f $X=10.16 $Y=2.37
+ $X2=0 $Y2=0
cc_1000 N_A_2008_48#_c_1439_n N_A_1747_74#_c_1582_n 0.0472402f $X=10.36 $Y=1.815
+ $X2=0 $Y2=0
cc_1001 N_A_2008_48#_c_1449_n N_A_1747_74#_c_1582_n 0.00840223f $X=10.525
+ $Y=2.405 $X2=0 $Y2=0
cc_1002 N_A_2008_48#_M1005_g N_A_1747_74#_c_1583_n 0.00782885f $X=10.115 $Y=0.58
+ $X2=0 $Y2=0
cc_1003 N_A_2008_48#_M1005_g N_A_1747_74#_c_1584_n 0.0151836f $X=10.115 $Y=0.58
+ $X2=0 $Y2=0
cc_1004 N_A_2008_48#_c_1438_n N_A_1747_74#_c_1584_n 0.00516648f $X=10.16 $Y=1.98
+ $X2=0 $Y2=0
cc_1005 N_A_2008_48#_c_1439_n N_A_1747_74#_c_1584_n 0.0174506f $X=10.36 $Y=1.815
+ $X2=0 $Y2=0
cc_1006 N_A_2008_48#_c_1440_n N_A_1747_74#_c_1584_n 0.00792529f $X=11.675
+ $Y=0.665 $X2=0 $Y2=0
cc_1007 N_A_2008_48#_c_1452_n N_A_1747_74#_c_1584_n 0.00127707f $X=11.675
+ $Y=1.715 $X2=0 $Y2=0
cc_1008 N_A_2008_48#_c_1441_n N_A_1747_74#_c_1584_n 0.0125719f $X=11.405
+ $Y=1.715 $X2=0 $Y2=0
cc_1009 N_A_2008_48#_c_1442_n N_A_1747_74#_c_1584_n 0.0245935f $X=11.76 $Y=1.63
+ $X2=0 $Y2=0
cc_1010 N_A_2008_48#_c_1443_n N_A_1747_74#_c_1584_n 0.017591f $X=11.12 $Y=0.55
+ $X2=0 $Y2=0
cc_1011 N_A_2008_48#_c_1448_n N_VPWR_M1003_d 0.00157126f $X=10.855 $Y=2.405
+ $X2=0 $Y2=0
cc_1012 N_A_2008_48#_c_1449_n N_VPWR_M1003_d 0.00330343f $X=10.525 $Y=2.405
+ $X2=0 $Y2=0
cc_1013 N_A_2008_48#_c_1454_n N_VPWR_M1031_d 7.76434e-19 $X=11.13 $Y=2.405 $X2=0
+ $Y2=0
cc_1014 N_A_2008_48#_c_1438_n N_VPWR_c_1809_n 6.38002e-19 $X=10.16 $Y=1.98 $X2=0
+ $Y2=0
cc_1015 N_A_2008_48#_c_1446_n N_VPWR_c_1809_n 0.0080003f $X=10.16 $Y=2.37 $X2=0
+ $Y2=0
cc_1016 N_A_2008_48#_c_1448_n N_VPWR_c_1809_n 0.00951507f $X=10.855 $Y=2.405
+ $X2=0 $Y2=0
cc_1017 N_A_2008_48#_c_1449_n N_VPWR_c_1809_n 0.0187155f $X=10.525 $Y=2.405
+ $X2=0 $Y2=0
cc_1018 N_A_2008_48#_c_1450_n N_VPWR_c_1809_n 0.0152062f $X=11.02 $Y=2.655 $X2=0
+ $Y2=0
cc_1019 N_A_2008_48#_c_1450_n N_VPWR_c_1923_n 0.00796791f $X=11.02 $Y=2.655
+ $X2=0 $Y2=0
cc_1020 N_A_2008_48#_c_1451_n N_VPWR_c_1923_n 0.0240111f $X=11.32 $Y=2.32 $X2=0
+ $Y2=0
cc_1021 N_A_2008_48#_c_1452_n N_VPWR_c_1923_n 0.019153f $X=11.675 $Y=1.715 $X2=0
+ $Y2=0
cc_1022 N_A_2008_48#_c_1454_n N_VPWR_c_1923_n 0.0135229f $X=11.13 $Y=2.405 $X2=0
+ $Y2=0
cc_1023 N_A_2008_48#_c_1450_n N_VPWR_c_1818_n 0.00744123f $X=11.02 $Y=2.655
+ $X2=0 $Y2=0
cc_1024 N_A_2008_48#_c_1454_n N_VPWR_c_1818_n 0.00211481f $X=11.13 $Y=2.405
+ $X2=0 $Y2=0
cc_1025 N_A_2008_48#_c_1446_n N_VPWR_c_1821_n 0.00502154f $X=10.16 $Y=2.37 $X2=0
+ $Y2=0
cc_1026 N_A_2008_48#_c_1450_n N_VPWR_c_1822_n 0.0103547f $X=11.02 $Y=2.655 $X2=0
+ $Y2=0
cc_1027 N_A_2008_48#_c_1446_n N_VPWR_c_1803_n 0.00515964f $X=10.16 $Y=2.37 $X2=0
+ $Y2=0
cc_1028 N_A_2008_48#_c_1448_n N_VPWR_c_1803_n 0.00704664f $X=10.855 $Y=2.405
+ $X2=0 $Y2=0
cc_1029 N_A_2008_48#_c_1449_n N_VPWR_c_1803_n 0.00241369f $X=10.525 $Y=2.405
+ $X2=0 $Y2=0
cc_1030 N_A_2008_48#_c_1450_n N_VPWR_c_1803_n 0.011288f $X=11.02 $Y=2.655 $X2=0
+ $Y2=0
cc_1031 N_A_2008_48#_c_1454_n N_VPWR_c_1803_n 0.00672753f $X=11.13 $Y=2.405
+ $X2=0 $Y2=0
cc_1032 N_A_2008_48#_c_1451_n Q_N 0.00264229f $X=11.32 $Y=2.32 $X2=0 $Y2=0
cc_1033 N_A_2008_48#_c_1452_n Q_N 0.0140768f $X=11.675 $Y=1.715 $X2=0 $Y2=0
cc_1034 N_A_2008_48#_c_1442_n Q_N 0.0510002f $X=11.76 $Y=1.63 $X2=0 $Y2=0
cc_1035 N_A_2008_48#_c_1440_n N_VGND_M1008_s 0.00795702f $X=11.675 $Y=0.665
+ $X2=0 $Y2=0
cc_1036 N_A_2008_48#_c_1442_n N_VGND_M1008_s 0.00751007f $X=11.76 $Y=1.63 $X2=0
+ $Y2=0
cc_1037 N_A_2008_48#_M1005_g N_VGND_c_2178_n 0.0106684f $X=10.115 $Y=0.58 $X2=0
+ $Y2=0
cc_1038 N_A_2008_48#_c_1443_n N_VGND_c_2178_n 0.0133829f $X=11.12 $Y=0.55 $X2=0
+ $Y2=0
cc_1039 N_A_2008_48#_M1005_g N_VGND_c_2187_n 0.00383152f $X=10.115 $Y=0.58 $X2=0
+ $Y2=0
cc_1040 N_A_2008_48#_c_1440_n N_VGND_c_2188_n 0.00463151f $X=11.675 $Y=0.665
+ $X2=0 $Y2=0
cc_1041 N_A_2008_48#_c_1443_n N_VGND_c_2188_n 0.0140232f $X=11.12 $Y=0.55 $X2=0
+ $Y2=0
cc_1042 N_A_2008_48#_M1005_g N_VGND_c_2190_n 0.0075694f $X=10.115 $Y=0.58 $X2=0
+ $Y2=0
cc_1043 N_A_2008_48#_c_1440_n N_VGND_c_2190_n 0.00869887f $X=11.675 $Y=0.665
+ $X2=0 $Y2=0
cc_1044 N_A_2008_48#_c_1443_n N_VGND_c_2190_n 0.0117897f $X=11.12 $Y=0.55 $X2=0
+ $Y2=0
cc_1045 N_A_2008_48#_c_1440_n N_VGND_c_2194_n 0.0253659f $X=11.675 $Y=0.665
+ $X2=0 $Y2=0
cc_1046 N_A_2008_48#_c_1443_n N_VGND_c_2194_n 0.00410713f $X=11.12 $Y=0.55 $X2=0
+ $Y2=0
cc_1047 N_A_1747_74#_M1002_g N_A_2513_424#_M1039_g 0.0206457f $X=12.93 $Y=0.645
+ $X2=0 $Y2=0
cc_1048 N_A_1747_74#_c_1590_n N_A_2513_424#_c_1754_n 0.00504987f $X=12.915
+ $Y=1.955 $X2=0 $Y2=0
cc_1049 N_A_1747_74#_c_1591_n N_A_2513_424#_c_1754_n 0.00577491f $X=12.915
+ $Y=2.045 $X2=0 $Y2=0
cc_1050 N_A_1747_74#_M1002_g N_A_2513_424#_c_1754_n 0.0214527f $X=12.93 $Y=0.645
+ $X2=0 $Y2=0
cc_1051 N_A_1747_74#_c_1580_n N_A_2513_424#_c_1754_n 0.00491452f $X=12.915
+ $Y=1.52 $X2=0 $Y2=0
cc_1052 N_A_1747_74#_c_1576_n N_A_2513_424#_c_1755_n 0.00194375f $X=11.965
+ $Y=1.235 $X2=0 $Y2=0
cc_1053 N_A_1747_74#_M1002_g N_A_2513_424#_c_1755_n 0.0144342f $X=12.93 $Y=0.645
+ $X2=0 $Y2=0
cc_1054 N_A_1747_74#_c_1577_n N_A_2513_424#_c_1759_n 0.00842101f $X=12.825
+ $Y=1.52 $X2=0 $Y2=0
cc_1055 N_A_1747_74#_c_1590_n N_A_2513_424#_c_1759_n 0.00946828f $X=12.915
+ $Y=1.955 $X2=0 $Y2=0
cc_1056 N_A_1747_74#_c_1591_n N_A_2513_424#_c_1759_n 0.0176712f $X=12.915
+ $Y=2.045 $X2=0 $Y2=0
cc_1057 N_A_1747_74#_c_1580_n N_A_2513_424#_c_1759_n 0.00107618f $X=12.915
+ $Y=1.52 $X2=0 $Y2=0
cc_1058 N_A_1747_74#_M1002_g N_A_2513_424#_c_1756_n 0.00833371f $X=12.93
+ $Y=0.645 $X2=0 $Y2=0
cc_1059 N_A_1747_74#_c_1580_n N_A_2513_424#_c_1756_n 0.0134227f $X=12.915
+ $Y=1.52 $X2=0 $Y2=0
cc_1060 N_A_1747_74#_c_1577_n N_A_2513_424#_c_1757_n 0.0160046f $X=12.825
+ $Y=1.52 $X2=0 $Y2=0
cc_1061 N_A_1747_74#_c_1578_n N_A_2513_424#_c_1757_n 2.29508e-19 $X=12.04
+ $Y=1.52 $X2=0 $Y2=0
cc_1062 N_A_1747_74#_M1002_g N_A_2513_424#_c_1757_n 0.00105416f $X=12.93
+ $Y=0.645 $X2=0 $Y2=0
cc_1063 N_A_1747_74#_c_1580_n N_A_2513_424#_c_1757_n 7.76856e-19 $X=12.915
+ $Y=1.52 $X2=0 $Y2=0
cc_1064 N_A_1747_74#_c_1594_n N_VPWR_c_1809_n 0.00666746f $X=9.925 $Y=2.59 $X2=0
+ $Y2=0
cc_1065 N_A_1747_74#_c_1587_n N_VPWR_c_1810_n 0.007084f $X=11.925 $Y=1.765 $X2=0
+ $Y2=0
cc_1066 N_A_1747_74#_c_1585_n N_VPWR_c_1923_n 0.00224083f $X=11.245 $Y=2.37
+ $X2=0 $Y2=0
cc_1067 N_A_1747_74#_c_1586_n N_VPWR_c_1923_n 0.00306886f $X=11.35 $Y=2.22 $X2=0
+ $Y2=0
cc_1068 N_A_1747_74#_c_1578_n N_VPWR_c_1923_n 0.00131549f $X=12.04 $Y=1.52 $X2=0
+ $Y2=0
cc_1069 N_A_1747_74#_c_1590_n N_VPWR_c_1811_n 0.00204598f $X=12.915 $Y=1.955
+ $X2=0 $Y2=0
cc_1070 N_A_1747_74#_c_1591_n N_VPWR_c_1811_n 0.00440242f $X=12.915 $Y=2.045
+ $X2=0 $Y2=0
cc_1071 N_A_1747_74#_c_1585_n N_VPWR_c_1818_n 0.00493443f $X=11.245 $Y=2.37
+ $X2=0 $Y2=0
cc_1072 N_A_1747_74#_c_1592_n N_VPWR_c_1818_n 0.00100251f $X=11.35 $Y=2.295
+ $X2=0 $Y2=0
cc_1073 N_A_1747_74#_c_1594_n N_VPWR_c_1821_n 0.0144557f $X=9.925 $Y=2.59 $X2=0
+ $Y2=0
cc_1074 N_A_1747_74#_c_1595_n N_VPWR_c_1821_n 0.00507318f $X=9.325 $Y=2.59 $X2=0
+ $Y2=0
cc_1075 N_A_1747_74#_c_1585_n N_VPWR_c_1822_n 0.00497687f $X=11.245 $Y=2.37
+ $X2=0 $Y2=0
cc_1076 N_A_1747_74#_c_1587_n N_VPWR_c_1823_n 0.00461464f $X=11.925 $Y=1.765
+ $X2=0 $Y2=0
cc_1077 N_A_1747_74#_c_1591_n N_VPWR_c_1823_n 0.00445602f $X=12.915 $Y=2.045
+ $X2=0 $Y2=0
cc_1078 N_A_1747_74#_c_1585_n N_VPWR_c_1803_n 0.00515964f $X=11.245 $Y=2.37
+ $X2=0 $Y2=0
cc_1079 N_A_1747_74#_c_1587_n N_VPWR_c_1803_n 0.00917882f $X=11.925 $Y=1.765
+ $X2=0 $Y2=0
cc_1080 N_A_1747_74#_c_1591_n N_VPWR_c_1803_n 0.00862843f $X=12.915 $Y=2.045
+ $X2=0 $Y2=0
cc_1081 N_A_1747_74#_c_1594_n N_VPWR_c_1803_n 0.023611f $X=9.925 $Y=2.59 $X2=0
+ $Y2=0
cc_1082 N_A_1747_74#_c_1595_n N_VPWR_c_1803_n 0.00697584f $X=9.325 $Y=2.59 $X2=0
+ $Y2=0
cc_1083 N_A_1747_74#_c_1594_n A_1969_489# 0.0021089f $X=9.925 $Y=2.59 $X2=-0.19
+ $Y2=-0.245
cc_1084 N_A_1747_74#_c_1587_n Q_N 0.00308691f $X=11.925 $Y=1.765 $X2=0 $Y2=0
cc_1085 N_A_1747_74#_c_1576_n Q_N 0.0192064f $X=11.965 $Y=1.235 $X2=0 $Y2=0
cc_1086 N_A_1747_74#_c_1577_n Q_N 0.0275523f $X=12.825 $Y=1.52 $X2=0 $Y2=0
cc_1087 N_A_1747_74#_c_1578_n Q_N 0.0123682f $X=12.04 $Y=1.52 $X2=0 $Y2=0
cc_1088 N_A_1747_74#_c_1590_n Q_N 0.00153041f $X=12.915 $Y=1.955 $X2=0 $Y2=0
cc_1089 N_A_1747_74#_c_1591_n Q_N 0.00229735f $X=12.915 $Y=2.045 $X2=0 $Y2=0
cc_1090 N_A_1747_74#_M1002_g Q_N 0.00438444f $X=12.93 $Y=0.645 $X2=0 $Y2=0
cc_1091 N_A_1747_74#_c_1573_n N_VGND_c_2178_n 0.00170773f $X=10.905 $Y=0.87
+ $X2=0 $Y2=0
cc_1092 N_A_1747_74#_c_1627_n N_VGND_c_2178_n 0.0133993f $X=9.605 $Y=0.57 $X2=0
+ $Y2=0
cc_1093 N_A_1747_74#_c_1581_n N_VGND_c_2178_n 8.97539e-19 $X=9.69 $Y=1.005 $X2=0
+ $Y2=0
cc_1094 N_A_1747_74#_c_1584_n N_VGND_c_2178_n 0.0179642f $X=11.26 $Y=1.27 $X2=0
+ $Y2=0
cc_1095 N_A_1747_74#_c_1576_n N_VGND_c_2179_n 0.00434272f $X=11.965 $Y=1.235
+ $X2=0 $Y2=0
cc_1096 N_A_1747_74#_M1002_g N_VGND_c_2179_n 0.00461464f $X=12.93 $Y=0.645 $X2=0
+ $Y2=0
cc_1097 N_A_1747_74#_M1002_g N_VGND_c_2180_n 0.0103391f $X=12.93 $Y=0.645 $X2=0
+ $Y2=0
cc_1098 N_A_1747_74#_c_1627_n N_VGND_c_2187_n 0.0207002f $X=9.605 $Y=0.57 $X2=0
+ $Y2=0
cc_1099 N_A_1747_74#_c_1573_n N_VGND_c_2188_n 0.00434272f $X=10.905 $Y=0.87
+ $X2=0 $Y2=0
cc_1100 N_A_1747_74#_c_1573_n N_VGND_c_2190_n 0.00825669f $X=10.905 $Y=0.87
+ $X2=0 $Y2=0
cc_1101 N_A_1747_74#_c_1576_n N_VGND_c_2190_n 0.0083017f $X=11.965 $Y=1.235
+ $X2=0 $Y2=0
cc_1102 N_A_1747_74#_M1002_g N_VGND_c_2190_n 0.00914946f $X=12.93 $Y=0.645 $X2=0
+ $Y2=0
cc_1103 N_A_1747_74#_c_1627_n N_VGND_c_2190_n 0.0219224f $X=9.605 $Y=0.57 $X2=0
+ $Y2=0
cc_1104 N_A_1747_74#_c_1573_n N_VGND_c_2194_n 0.00289541f $X=10.905 $Y=0.87
+ $X2=0 $Y2=0
cc_1105 N_A_1747_74#_c_1576_n N_VGND_c_2194_n 0.00583402f $X=11.965 $Y=1.235
+ $X2=0 $Y2=0
cc_1106 N_A_2513_424#_c_1754_n N_VPWR_c_1811_n 0.00624321f $X=13.435 $Y=1.765
+ $X2=0 $Y2=0
cc_1107 N_A_2513_424#_c_1759_n N_VPWR_c_1811_n 0.0507962f $X=12.69 $Y=2.265
+ $X2=0 $Y2=0
cc_1108 N_A_2513_424#_c_1756_n N_VPWR_c_1811_n 0.0222736f $X=13.38 $Y=1.465
+ $X2=0 $Y2=0
cc_1109 N_A_2513_424#_c_1759_n N_VPWR_c_1823_n 0.0125859f $X=12.69 $Y=2.265
+ $X2=0 $Y2=0
cc_1110 N_A_2513_424#_c_1754_n N_VPWR_c_1824_n 0.00461464f $X=13.435 $Y=1.765
+ $X2=0 $Y2=0
cc_1111 N_A_2513_424#_c_1754_n N_VPWR_c_1803_n 0.0091238f $X=13.435 $Y=1.765
+ $X2=0 $Y2=0
cc_1112 N_A_2513_424#_c_1759_n N_VPWR_c_1803_n 0.0103846f $X=12.69 $Y=2.265
+ $X2=0 $Y2=0
cc_1113 N_A_2513_424#_c_1755_n Q_N 0.0571733f $X=12.715 $Y=0.645 $X2=0 $Y2=0
cc_1114 N_A_2513_424#_c_1759_n Q_N 0.0895806f $X=12.69 $Y=2.265 $X2=0 $Y2=0
cc_1115 N_A_2513_424#_c_1757_n Q_N 0.0215198f $X=12.712 $Y=1.465 $X2=0 $Y2=0
cc_1116 N_A_2513_424#_M1039_g Q 0.00811057f $X=13.42 $Y=0.74 $X2=0 $Y2=0
cc_1117 N_A_2513_424#_M1039_g Q 0.00301691f $X=13.42 $Y=0.74 $X2=0 $Y2=0
cc_1118 N_A_2513_424#_c_1754_n Q 0.00230594f $X=13.435 $Y=1.765 $X2=0 $Y2=0
cc_1119 N_A_2513_424#_c_1756_n Q 0.00111755f $X=13.38 $Y=1.465 $X2=0 $Y2=0
cc_1120 N_A_2513_424#_c_1754_n Q 0.00190204f $X=13.435 $Y=1.765 $X2=0 $Y2=0
cc_1121 N_A_2513_424#_M1039_g N_Q_c_2156_n 0.0040915f $X=13.42 $Y=0.74 $X2=0
+ $Y2=0
cc_1122 N_A_2513_424#_c_1754_n N_Q_c_2156_n 0.0129497f $X=13.435 $Y=1.765 $X2=0
+ $Y2=0
cc_1123 N_A_2513_424#_c_1756_n N_Q_c_2156_n 0.0250949f $X=13.38 $Y=1.465 $X2=0
+ $Y2=0
cc_1124 N_A_2513_424#_c_1755_n N_VGND_c_2179_n 0.00778672f $X=12.715 $Y=0.645
+ $X2=0 $Y2=0
cc_1125 N_A_2513_424#_M1039_g N_VGND_c_2180_n 0.00330159f $X=13.42 $Y=0.74 $X2=0
+ $Y2=0
cc_1126 N_A_2513_424#_c_1754_n N_VGND_c_2180_n 0.00172388f $X=13.435 $Y=1.765
+ $X2=0 $Y2=0
cc_1127 N_A_2513_424#_c_1755_n N_VGND_c_2180_n 0.035427f $X=12.715 $Y=0.645
+ $X2=0 $Y2=0
cc_1128 N_A_2513_424#_c_1756_n N_VGND_c_2180_n 0.0145561f $X=13.38 $Y=1.465
+ $X2=0 $Y2=0
cc_1129 N_A_2513_424#_M1039_g N_VGND_c_2189_n 0.00434272f $X=13.42 $Y=0.74 $X2=0
+ $Y2=0
cc_1130 N_A_2513_424#_M1039_g N_VGND_c_2190_n 0.00824587f $X=13.42 $Y=0.74 $X2=0
+ $Y2=0
cc_1131 N_A_2513_424#_c_1755_n N_VGND_c_2190_n 0.00976756f $X=12.715 $Y=0.645
+ $X2=0 $Y2=0
cc_1132 N_VPWR_c_1805_n N_A_413_90#_c_1994_n 0.0213404f $X=3.265 $Y=2.815 $X2=0
+ $Y2=0
cc_1133 N_VPWR_c_1814_n N_A_413_90#_c_1994_n 0.0171392f $X=4.705 $Y=3.33 $X2=0
+ $Y2=0
cc_1134 N_VPWR_c_1803_n N_A_413_90#_c_1994_n 0.013307f $X=13.68 $Y=3.33 $X2=0
+ $Y2=0
cc_1135 N_VPWR_M1025_d N_A_413_90#_c_1995_n 0.00454038f $X=4.72 $Y=1.82 $X2=0
+ $Y2=0
cc_1136 N_VPWR_c_1806_n N_A_413_90#_c_1995_n 0.0162763f $X=4.87 $Y=2.785 $X2=0
+ $Y2=0
cc_1137 N_VPWR_c_1803_n N_A_413_90#_c_1995_n 0.0489602f $X=13.68 $Y=3.33 $X2=0
+ $Y2=0
cc_1138 N_VPWR_c_1804_n N_A_413_90#_c_1998_n 0.0180232f $X=1.39 $Y=2.475 $X2=0
+ $Y2=0
cc_1139 N_VPWR_c_1805_n N_A_413_90#_c_1998_n 0.00657188f $X=3.265 $Y=2.815 $X2=0
+ $Y2=0
cc_1140 N_VPWR_c_1819_n N_A_413_90#_c_1998_n 0.0156984f $X=3.085 $Y=3.33 $X2=0
+ $Y2=0
cc_1141 N_VPWR_c_1803_n N_A_413_90#_c_1998_n 0.0120809f $X=13.68 $Y=3.33 $X2=0
+ $Y2=0
cc_1142 N_VPWR_M1032_d N_A_413_90#_c_2004_n 0.0114582f $X=3.1 $Y=2.32 $X2=0
+ $Y2=0
cc_1143 N_VPWR_c_1805_n N_A_413_90#_c_2004_n 0.0236929f $X=3.265 $Y=2.815 $X2=0
+ $Y2=0
cc_1144 N_VPWR_c_1803_n N_A_413_90#_c_2004_n 0.0235866f $X=13.68 $Y=3.33 $X2=0
+ $Y2=0
cc_1145 N_VPWR_M1032_d N_A_413_90#_c_1999_n 0.00148356f $X=3.1 $Y=2.32 $X2=0
+ $Y2=0
cc_1146 N_VPWR_c_1803_n N_A_413_90#_c_1999_n 0.00583441f $X=13.68 $Y=3.33 $X2=0
+ $Y2=0
cc_1147 N_VPWR_c_1816_n N_A_413_90#_c_2000_n 0.00570315f $X=7.09 $Y=3.33 $X2=0
+ $Y2=0
cc_1148 N_VPWR_c_1803_n N_A_413_90#_c_2000_n 0.00689183f $X=13.68 $Y=3.33 $X2=0
+ $Y2=0
cc_1149 N_VPWR_c_1810_n Q_N 0.00144265f $X=11.592 $Y=3.245 $X2=0 $Y2=0
cc_1150 N_VPWR_c_1823_n Q_N 0.0146357f $X=13.045 $Y=3.33 $X2=0 $Y2=0
cc_1151 N_VPWR_c_1803_n Q_N 0.0121141f $X=13.68 $Y=3.33 $X2=0 $Y2=0
cc_1152 N_VPWR_c_1811_n Q 0.00249543f $X=13.21 $Y=1.985 $X2=0 $Y2=0
cc_1153 N_VPWR_c_1824_n Q 0.0124046f $X=13.68 $Y=3.33 $X2=0 $Y2=0
cc_1154 N_VPWR_c_1803_n Q 0.0102675f $X=13.68 $Y=3.33 $X2=0 $Y2=0
cc_1155 N_A_413_90#_c_2004_n A_512_464# 0.0137346f $X=3.445 $Y=2.44 $X2=-0.19
+ $Y2=-0.245
cc_1156 N_A_413_90#_c_1985_n N_noxref_25_c_2314_n 0.0184085f $X=3.445 $Y=1.005
+ $X2=0 $Y2=0
cc_1157 N_A_413_90#_c_1991_n N_noxref_25_c_2314_n 0.0224658f $X=2.435 $Y=0.76
+ $X2=0 $Y2=0
cc_1158 N_A_413_90#_c_1985_n N_noxref_25_c_2316_n 0.0246695f $X=3.445 $Y=1.005
+ $X2=0 $Y2=0
cc_1159 Q_N N_VGND_c_2179_n 0.0145639f $X=12.155 $Y=0.47 $X2=0 $Y2=0
cc_1160 Q_N N_VGND_c_2190_n 0.0119984f $X=12.155 $Y=0.47 $X2=0 $Y2=0
cc_1161 Q_N N_VGND_c_2194_n 0.00297405f $X=12.155 $Y=0.47 $X2=0 $Y2=0
cc_1162 Q N_VGND_c_2180_n 0.0297276f $X=13.595 $Y=0.47 $X2=0 $Y2=0
cc_1163 Q N_VGND_c_2189_n 0.0161257f $X=13.595 $Y=0.47 $X2=0 $Y2=0
cc_1164 Q N_VGND_c_2190_n 0.013291f $X=13.595 $Y=0.47 $X2=0 $Y2=0
cc_1165 N_VGND_c_2174_n N_noxref_25_c_2313_n 0.0253895f $X=0.71 $Y=0.58 $X2=0
+ $Y2=0
cc_1166 N_VGND_c_2181_n N_noxref_25_c_2314_n 0.11689f $X=3.67 $Y=0 $X2=0 $Y2=0
cc_1167 N_VGND_c_2190_n N_noxref_25_c_2314_n 0.068236f $X=13.68 $Y=0 $X2=0 $Y2=0
cc_1168 N_VGND_c_2174_n N_noxref_25_c_2315_n 0.0121617f $X=0.71 $Y=0.58 $X2=0
+ $Y2=0
cc_1169 N_VGND_c_2181_n N_noxref_25_c_2315_n 0.0176516f $X=3.67 $Y=0 $X2=0 $Y2=0
cc_1170 N_VGND_c_2190_n N_noxref_25_c_2315_n 0.00966868f $X=13.68 $Y=0 $X2=0
+ $Y2=0
cc_1171 N_VGND_c_2175_n N_noxref_25_c_2316_n 0.0153137f $X=3.835 $Y=0.585 $X2=0
+ $Y2=0
cc_1172 N_VGND_c_2181_n N_noxref_25_c_2316_n 0.0229596f $X=3.67 $Y=0 $X2=0 $Y2=0
cc_1173 N_VGND_c_2190_n N_noxref_25_c_2316_n 0.0126481f $X=13.68 $Y=0 $X2=0
+ $Y2=0
