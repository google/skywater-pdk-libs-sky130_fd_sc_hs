* NGSPICE file created from sky130_fd_sc_hs__dlclkp_4.ext - technology: sky130A

.subckt sky130_fd_sc_hs__dlclkp_4 CLK GATE VGND VNB VPB VPWR GCLK
M1000 VGND a_27_74# a_491_124# VNB nlowvt w=420000u l=150000u
+  ad=1.78525e+12p pd=1.468e+07u as=2.3775e+11p ps=2.39e+06u
M1001 VPWR a_1044_368# GCLK VPB pshort w=1.12e+06u l=150000u
+  ad=3.1894e+12p pd=1.939e+07u as=6.888e+11p ps=5.71e+06u
M1002 a_283_392# GATE VPWR VPB pshort w=1e+06u l=150000u
+  ad=2.7e+11p pd=2.54e+06u as=0p ps=0u
M1003 a_524_508# a_334_54# a_84_48# VPB pshort w=420000u l=150000u
+  ad=1.134e+11p pd=1.38e+06u as=4.204e+11p ps=3.27e+06u
M1004 a_334_338# a_334_54# VPWR VPB pshort w=840000u l=150000u
+  ad=2.478e+11p pd=2.27e+06u as=0p ps=0u
M1005 a_1047_74# CLK VGND VNB nlowvt w=740000u l=150000u
+  ad=1.776e+11p pd=1.96e+06u as=0p ps=0u
M1006 GCLK a_1044_368# VGND VNB nlowvt w=740000u l=150000u
+  ad=4.144e+11p pd=4.08e+06u as=0p ps=0u
M1007 VPWR a_27_74# a_1044_368# VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=3.752e+11p ps=2.91e+06u
M1008 VGND a_1044_368# GCLK VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_84_48# a_334_338# a_283_392# VPB pshort w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VPWR a_27_74# a_524_508# VPB pshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VPWR a_84_48# a_27_74# VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=3.304e+11p ps=2.83e+06u
M1012 a_491_124# a_334_338# a_84_48# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=2.587e+11p ps=2.25e+06u
M1013 VGND a_1044_368# GCLK VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_1044_368# CLK VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 GCLK a_1044_368# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VPWR CLK a_334_54# VPB pshort w=840000u l=150000u
+  ad=0p pd=0u as=2.478e+11p ps=2.27e+06u
M1017 a_286_80# GATE VGND VNB nlowvt w=640000u l=150000u
+  ad=1.536e+11p pd=1.76e+06u as=0p ps=0u
M1018 a_84_48# a_334_54# a_286_80# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VGND CLK a_334_54# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.333e+11p ps=2.19e+06u
M1020 GCLK a_1044_368# VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 VGND a_84_48# a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1022 GCLK a_1044_368# VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_1044_368# a_27_74# a_1047_74# VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1024 VPWR a_1044_368# GCLK VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 a_334_338# a_334_54# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.675e+11p pd=2.66e+06u as=0p ps=0u
.ends

