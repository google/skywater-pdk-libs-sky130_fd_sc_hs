* File: sky130_fd_sc_hs__o211ai_4.spice
* Created: Tue Sep  1 20:14:06 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hs__o211ai_4.pex.spice"
.subckt sky130_fd_sc_hs__o211ai_4  VNB VPB A1 A2 B1 C1 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* C1	C1
* B1	B1
* A2	A2
* A1	A1
* VPB	VPB
* VNB	VNB
MM1010 N_A_27_74#_M1010_d N_A1_M1010_g N_VGND_M1010_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.1295 PD=2.05 PS=1.09 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75000.2
+ SB=75005.1 A=0.111 P=1.78 MULT=1
MM1014 N_A_27_74#_M1014_d N_A1_M1014_g N_VGND_M1010_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1295 PD=1.02 PS=1.09 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.7
+ SB=75004.6 A=0.111 P=1.78 MULT=1
MM1019 N_A_27_74#_M1014_d N_A1_M1019_g N_VGND_M1019_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1295 PD=1.02 PS=1.09 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75001.1
+ SB=75004.2 A=0.111 P=1.78 MULT=1
MM1023 N_A_27_74#_M1023_d N_A1_M1023_g N_VGND_M1019_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1295 PD=1.02 PS=1.09 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.6
+ SB=75003.7 A=0.111 P=1.78 MULT=1
MM1006 N_VGND_M1006_d N_A2_M1006_g N_A_27_74#_M1023_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75002.1
+ SB=75003.2 A=0.111 P=1.78 MULT=1
MM1007 N_VGND_M1006_d N_A2_M1007_g N_A_27_74#_M1007_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75002.5
+ SB=75002.8 A=0.111 P=1.78 MULT=1
MM1009 N_VGND_M1009_d N_A2_M1009_g N_A_27_74#_M1007_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.111 AS=0.1036 PD=1.04 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75002.9
+ SB=75002.4 A=0.111 P=1.78 MULT=1
MM1012 N_VGND_M1009_d N_A2_M1012_g N_A_27_74#_M1012_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.111 AS=0.1036 PD=1.04 PS=1.02 NRD=3.24 NRS=0 M=1 R=4.93333 SA=75003.4
+ SB=75001.9 A=0.111 P=1.78 MULT=1
MM1008 N_A_834_74#_M1008_d N_B1_M1008_g N_A_27_74#_M1012_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75003.8 SB=75001.5 A=0.111 P=1.78 MULT=1
MM1011 N_A_834_74#_M1008_d N_B1_M1011_g N_A_27_74#_M1011_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75004.2 SB=75001.1 A=0.111 P=1.78 MULT=1
MM1016 N_A_834_74#_M1016_d N_B1_M1016_g N_A_27_74#_M1011_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75004.7 SB=75000.6 A=0.111 P=1.78 MULT=1
MM1017 N_A_834_74#_M1016_d N_B1_M1017_g N_A_27_74#_M1017_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.2109 PD=1.02 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75005.1 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1002 N_Y_M1002_d N_C1_M1002_g N_A_834_74#_M1002_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.2109 PD=1.02 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75001.5 A=0.111 P=1.78 MULT=1
MM1005 N_Y_M1002_d N_C1_M1005_g N_A_834_74#_M1005_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.6
+ SB=75001.1 A=0.111 P=1.78 MULT=1
MM1013 N_Y_M1013_d N_C1_M1013_g N_A_834_74#_M1005_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.1
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1015 N_Y_M1013_d N_C1_M1015_g N_A_834_74#_M1015_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.2109 PD=1.02 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.5
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1020 N_VPWR_M1020_d N_A1_M1020_g N_A_30_368#_M1020_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.3304 PD=1.42 PS=2.83 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75003.5 A=0.168 P=2.54 MULT=1
MM1021 N_VPWR_M1020_d N_A1_M1021_g N_A_30_368#_M1021_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.7 SB=75003.1 A=0.168 P=2.54 MULT=1
MM1024 N_VPWR_M1024_d N_A1_M1024_g N_A_30_368#_M1021_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.1 SB=75002.6 A=0.168 P=2.54 MULT=1
MM1026 N_VPWR_M1024_d N_A1_M1026_g N_A_30_368#_M1026_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.196 PD=1.42 PS=1.47 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.6 SB=75002.2 A=0.168 P=2.54 MULT=1
MM1000 N_A_30_368#_M1026_s N_A2_M1000_g N_Y_M1000_s VPB PSHORT L=0.15 W=1.12
+ AD=0.196 AS=0.168 PD=1.47 PS=1.42 NRD=10.5395 NRS=1.7533 M=1 R=7.46667
+ SA=75002.1 SB=75001.7 A=0.168 P=2.54 MULT=1
MM1003 N_A_30_368#_M1003_d N_A2_M1003_g N_Y_M1000_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75002.5 SB=75001.2 A=0.168 P=2.54 MULT=1
MM1004 N_A_30_368#_M1003_d N_A2_M1004_g N_Y_M1004_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.196 PD=1.42 PS=1.47 NRD=1.7533 NRS=10.5395 M=1 R=7.46667
+ SA=75003 SB=75000.8 A=0.168 P=2.54 MULT=1
MM1027 N_A_30_368#_M1027_d N_A2_M1027_g N_Y_M1004_s VPB PSHORT L=0.15 W=1.12
+ AD=0.3864 AS=0.196 PD=2.93 PS=1.47 NRD=10.5395 NRS=1.7533 M=1 R=7.46667
+ SA=75003.5 SB=75000.3 A=0.168 P=2.54 MULT=1
MM1001 N_VPWR_M1001_d N_B1_M1001_g N_Y_M1001_s VPB PSHORT L=0.15 W=1.12
+ AD=0.3304 AS=0.2184 PD=2.83 PS=1.51 NRD=1.7533 NRS=10.5395 M=1 R=7.46667
+ SA=75000.2 SB=75002.3 A=0.168 P=2.54 MULT=1
MM1018 N_VPWR_M1018_d N_B1_M1018_g N_Y_M1001_s VPB PSHORT L=0.15 W=1.12
+ AD=0.2016 AS=0.2184 PD=1.48 PS=1.51 NRD=3.5066 NRS=8.7862 M=1 R=7.46667
+ SA=75000.8 SB=75001.7 A=0.168 P=2.54 MULT=1
MM1022 N_Y_M1022_d N_C1_M1022_g N_VPWR_M1018_d VPB PSHORT L=0.15 W=1.12 AD=0.168
+ AS=0.2016 PD=1.42 PS=1.48 NRD=1.7533 NRS=10.5395 M=1 R=7.46667 SA=75001.3
+ SB=75001.2 A=0.168 P=2.54 MULT=1
MM1025 N_Y_M1022_d N_C1_M1025_g N_VPWR_M1025_s VPB PSHORT L=0.15 W=1.12 AD=0.168
+ AS=0.9688 PD=1.42 PS=3.97 NRD=1.7533 NRS=1.7533 M=1 R=7.46667 SA=75001.7
+ SB=75000.8 A=0.168 P=2.54 MULT=1
DX28_noxref VNB VPB NWDIODE A=15.8844 P=20.8
c_76 VNB 0 1.29151e-19 $X=0 $Y=0
*
.include "sky130_fd_sc_hs__o211ai_4.pxi.spice"
*
.ends
*
*
