# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_hs__or4bb_2
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_hs__or4bb_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.800000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.485000 1.470000 3.925000 1.800000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.150000 0.255000 3.715000 0.570000 ;
        RECT 3.485000 0.570000 3.715000 0.670000 ;
    END
  END B
  PIN C_N
    ANTENNAGATEAREA  0.208500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.435000 1.300000 4.695000 1.780000 ;
    END
  END C_N
  PIN D_N
    ANTENNAGATEAREA  0.208500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.350000 0.550000 1.780000 ;
    END
  END D_N
  PIN X
    ANTENNADIFFAREA  0.543200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.060000 0.440000 1.315000 1.180000 ;
        RECT 1.060000 1.180000 1.230000 1.850000 ;
        RECT 1.060000 1.850000 1.390000 2.100000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 4.800000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 4.800000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.800000 0.085000 ;
      RECT 0.000000  3.245000 4.800000 3.415000 ;
      RECT 0.105000  2.100000 0.890000 2.270000 ;
      RECT 0.105000  2.270000 2.265000 2.440000 ;
      RECT 0.105000  2.440000 0.435000 2.980000 ;
      RECT 0.120000  0.670000 0.450000 1.010000 ;
      RECT 0.120000  1.010000 0.890000 1.180000 ;
      RECT 0.605000  2.610000 0.935000 3.245000 ;
      RECT 0.630000  0.085000 0.880000 0.840000 ;
      RECT 0.720000  1.180000 0.890000 2.100000 ;
      RECT 1.400000  1.350000 1.730000 1.680000 ;
      RECT 1.510000  2.610000 1.840000 3.245000 ;
      RECT 1.560000  1.130000 3.735000 1.300000 ;
      RECT 1.560000  1.300000 1.730000 1.350000 ;
      RECT 1.575000  0.085000 2.035000 0.910000 ;
      RECT 1.970000  1.470000 2.265000 2.270000 ;
      RECT 2.050000  2.610000 2.605000 2.780000 ;
      RECT 2.050000  2.780000 2.380000 2.980000 ;
      RECT 2.310000  0.580000 2.640000 1.130000 ;
      RECT 2.435000  1.300000 2.605000 2.610000 ;
      RECT 2.775000  1.470000 3.070000 1.970000 ;
      RECT 2.775000  1.970000 4.690000 2.140000 ;
      RECT 2.810000  0.085000 2.980000 0.740000 ;
      RECT 2.810000  0.740000 3.195000 0.960000 ;
      RECT 3.405000  0.840000 3.735000 1.130000 ;
      RECT 3.820000  2.310000 4.150000 3.245000 ;
      RECT 3.925000  0.085000 4.255000 0.790000 ;
      RECT 4.095000  0.960000 4.685000 1.130000 ;
      RECT 4.095000  1.130000 4.265000 1.950000 ;
      RECT 4.095000  1.950000 4.690000 1.970000 ;
      RECT 4.360000  2.140000 4.690000 2.820000 ;
      RECT 4.435000  0.435000 4.685000 0.960000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
  END
END sky130_fd_sc_hs__or4bb_2
