* File: sky130_fd_sc_hs__sdlclkp_1.pex.spice
* Created: Thu Aug 27 21:10:34 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HS__SDLCLKP_1%SCE 2 5 7 9 10 13 14
r35 13 15 45.1558 $w=3.75e-07 $l=1.65e-07 $layer=POLY_cond $X=0.407 $Y=1.455
+ $X2=0.407 $Y2=1.29
r36 13 14 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.385
+ $Y=1.455 $X2=0.385 $Y2=1.455
r37 10 14 2.58853 $w=6.68e-07 $l=1.45e-07 $layer=LI1_cond $X=0.24 $Y=1.625
+ $X2=0.385 $Y2=1.625
r38 7 9 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=0.505 $Y=2.045
+ $X2=0.505 $Y2=2.54
r39 5 15 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=0.495 $Y=0.835
+ $X2=0.495 $Y2=1.29
r40 2 7 41.7529 $w=3.14e-07 $l=3.17238e-07 $layer=POLY_cond $X=0.407 $Y=1.773
+ $X2=0.505 $Y2=2.045
r41 1 13 3.26277 $w=3.75e-07 $l=2.2e-08 $layer=POLY_cond $X=0.407 $Y=1.477
+ $X2=0.407 $Y2=1.455
r42 1 2 43.8991 $w=3.75e-07 $l=2.96e-07 $layer=POLY_cond $X=0.407 $Y=1.477
+ $X2=0.407 $Y2=1.773
.ends

.subckt PM_SKY130_FD_SC_HS__SDLCLKP_1%GATE 1 3 6 8 12
r40 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.97
+ $Y=1.795 $X2=0.97 $Y2=1.795
r41 8 12 5.98039 $w=4.78e-07 $l=2.4e-07 $layer=LI1_cond $X=1.045 $Y=2.035
+ $X2=1.045 $Y2=1.795
r42 4 11 38.5562 $w=2.99e-07 $l=1.86145e-07 $layer=POLY_cond $X=0.925 $Y=1.63
+ $X2=0.97 $Y2=1.795
r43 4 6 407.649 $w=1.5e-07 $l=7.95e-07 $layer=POLY_cond $X=0.925 $Y=1.63
+ $X2=0.925 $Y2=0.835
r44 1 11 52.2586 $w=2.99e-07 $l=2.85044e-07 $layer=POLY_cond $X=0.895 $Y=2.045
+ $X2=0.97 $Y2=1.795
r45 1 3 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=0.895 $Y=2.045
+ $X2=0.895 $Y2=2.54
.ends

.subckt PM_SKY130_FD_SC_HS__SDLCLKP_1%A_318_74# 1 2 7 9 12 15 16 19 25 27 33
c77 33 0 6.25246e-20 $X=3 $Y=1.602
c78 27 0 8.55408e-20 $X=2.79 $Y=1.55
c79 7 0 1.13986e-19 $X=3 $Y=1.82
r80 33 34 35.2022 $w=3.56e-07 $l=2.6e-07 $layer=POLY_cond $X=3 $Y=1.602 $X2=3.26
+ $Y2=1.602
r81 28 33 28.4326 $w=3.56e-07 $l=2.1e-07 $layer=POLY_cond $X=2.79 $Y=1.602 $X2=3
+ $Y2=1.602
r82 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.79
+ $Y=1.55 $X2=2.79 $Y2=1.55
r83 24 25 10.1887 $w=6.03e-07 $l=1.65e-07 $layer=LI1_cond $X=2.215 $Y=1.847
+ $X2=2.38 $Y2=1.847
r84 19 20 8.06167 $w=2.27e-07 $l=1.5e-07 $layer=LI1_cond $X=1.73 $Y=1 $X2=1.88
+ $Y2=1
r85 16 27 3.35256 $w=2.73e-07 $l=8e-08 $layer=LI1_cond $X=2.762 $Y=1.63
+ $X2=2.762 $Y2=1.55
r86 16 25 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=2.625 $Y=1.63
+ $X2=2.38 $Y2=1.63
r87 15 24 6.62291 $w=6.03e-07 $l=3.35e-07 $layer=LI1_cond $X=1.88 $Y=1.847
+ $X2=2.215 $Y2=1.847
r88 14 20 2.43258 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=1.88 $Y=1.12 $X2=1.88
+ $Y2=1
r89 14 15 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=1.88 $Y=1.12
+ $X2=1.88 $Y2=1.545
r90 10 34 23.0368 $w=1.5e-07 $l=2.17e-07 $layer=POLY_cond $X=3.26 $Y=1.385
+ $X2=3.26 $Y2=1.602
r91 10 12 397.394 $w=1.5e-07 $l=7.75e-07 $layer=POLY_cond $X=3.26 $Y=1.385
+ $X2=3.26 $Y2=0.61
r92 7 33 23.0368 $w=1.5e-07 $l=2.18e-07 $layer=POLY_cond $X=3 $Y=1.82 $X2=3
+ $Y2=1.602
r93 7 9 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=3 $Y=1.82 $X2=3
+ $Y2=2.315
r94 2 24 600 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=2.065
+ $Y=1.84 $X2=2.215 $Y2=1.985
r95 1 19 182 $w=1.7e-07 $l=6.61306e-07 $layer=licon1_NDIFF $count=1 $X=1.59
+ $Y=0.37 $X2=1.73 $Y2=0.965
.ends

.subckt PM_SKY130_FD_SC_HS__SDLCLKP_1%A_288_48# 1 2 7 9 10 11 13 14 15 16 19 20
+ 21 22 23 24 26 27 29 30 33 34 35 37 38 39 41 42 43 47 49 51 54 58
c172 37 0 1.99229e-19 $X=3.495 $Y=0.88
c173 27 0 7.6749e-20 $X=3.535 $Y=2.955
c174 24 0 3.05753e-20 $X=2.755 $Y=0.995
r175 55 58 4.88915 $w=3.28e-07 $l=1.4e-07 $layer=LI1_cond $X=5.075 $Y=2.16
+ $X2=5.215 $Y2=2.16
r176 51 53 18.7692 $w=2.47e-07 $l=3.8e-07 $layer=LI1_cond $X=2.25 $Y=1.195
+ $X2=2.63 $Y2=1.195
r177 51 52 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.25
+ $Y=1.195 $X2=2.25 $Y2=1.195
r178 49 55 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.075 $Y=1.995
+ $X2=5.075 $Y2=2.16
r179 49 54 56.4332 $w=1.68e-07 $l=8.65e-07 $layer=LI1_cond $X=5.075 $Y=1.995
+ $X2=5.075 $Y2=1.13
r180 45 54 7.20219 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=5.065 $Y=0.965
+ $X2=5.065 $Y2=1.13
r181 45 47 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=5.065 $Y=0.965
+ $X2=5.065 $Y2=0.515
r182 44 47 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=5.065 $Y=0.425
+ $X2=5.065 $Y2=0.515
r183 42 44 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.9 $Y=0.34
+ $X2=5.065 $Y2=0.425
r184 42 43 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=4.9 $Y=0.34 $X2=4.26
+ $Y2=0.34
r185 40 43 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.175 $Y=0.425
+ $X2=4.26 $Y2=0.34
r186 40 41 29.6845 $w=1.68e-07 $l=4.55e-07 $layer=LI1_cond $X=4.175 $Y=0.425
+ $X2=4.175 $Y2=0.88
r187 38 41 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.09 $Y=0.965
+ $X2=4.175 $Y2=0.88
r188 38 39 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=4.09 $Y=0.965
+ $X2=3.58 $Y2=0.965
r189 37 39 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.495 $Y=0.88
+ $X2=3.58 $Y2=0.965
r190 36 37 29.6845 $w=1.68e-07 $l=4.55e-07 $layer=LI1_cond $X=3.495 $Y=0.425
+ $X2=3.495 $Y2=0.88
r191 34 36 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.41 $Y=0.34
+ $X2=3.495 $Y2=0.425
r192 34 35 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=3.41 $Y=0.34
+ $X2=2.715 $Y2=0.34
r193 33 53 2.92482 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.63 $Y=1.03
+ $X2=2.63 $Y2=1.195
r194 32 35 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.63 $Y=0.425
+ $X2=2.715 $Y2=0.34
r195 32 33 39.4706 $w=1.68e-07 $l=6.05e-07 $layer=LI1_cond $X=2.63 $Y=0.425
+ $X2=2.63 $Y2=1.03
r196 27 30 77.9482 $w=1.8e-07 $l=1.95e-07 $layer=POLY_cond $X=3.535 $Y=2.955
+ $X2=3.535 $Y2=3.15
r197 27 29 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=3.535 $Y=2.955
+ $X2=3.535 $Y2=2.67
r198 24 26 112.467 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=2.755 $Y=0.995
+ $X2=2.755 $Y2=0.645
r199 23 52 38.6443 $w=2.87e-07 $l=2.11849e-07 $layer=POLY_cond $X=2.415 $Y=1.07
+ $X2=2.25 $Y2=1.177
r200 22 24 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.68 $Y=1.07
+ $X2=2.755 $Y2=0.995
r201 22 23 135.883 $w=1.5e-07 $l=2.65e-07 $layer=POLY_cond $X=2.68 $Y=1.07
+ $X2=2.415 $Y2=1.07
r202 20 30 7.1379 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=3.445 $Y=3.15
+ $X2=3.535 $Y2=3.15
r203 20 21 699.926 $w=1.5e-07 $l=1.365e-06 $layer=POLY_cond $X=3.445 $Y=3.15
+ $X2=2.08 $Y2=3.15
r204 17 19 253.819 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=1.99 $Y=2.755
+ $X2=1.99 $Y2=2.26
r205 16 19 253.819 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=1.99 $Y=1.765
+ $X2=1.99 $Y2=2.26
r206 15 21 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=1.99 $Y=3.075
+ $X2=2.08 $Y2=3.15
r207 14 17 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=1.99 $Y=2.845
+ $X2=1.99 $Y2=2.755
r208 14 15 89.4032 $w=1.8e-07 $l=2.3e-07 $layer=POLY_cond $X=1.99 $Y=2.845
+ $X2=1.99 $Y2=3.075
r209 13 16 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=1.99 $Y=1.675
+ $X2=1.99 $Y2=1.765
r210 12 52 43.6655 $w=2.87e-07 $l=3.39382e-07 $layer=POLY_cond $X=1.99 $Y=1.36
+ $X2=2.25 $Y2=1.177
r211 12 13 122.444 $w=1.8e-07 $l=3.15e-07 $layer=POLY_cond $X=1.99 $Y=1.36
+ $X2=1.99 $Y2=1.675
r212 10 12 26.0485 $w=2.87e-07 $l=1.21861e-07 $layer=POLY_cond $X=1.9 $Y=1.285
+ $X2=1.99 $Y2=1.36
r213 10 11 158.957 $w=1.5e-07 $l=3.1e-07 $layer=POLY_cond $X=1.9 $Y=1.285
+ $X2=1.59 $Y2=1.285
r214 7 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.515 $Y=1.21
+ $X2=1.59 $Y2=1.285
r215 7 9 151.027 $w=1.5e-07 $l=4.7e-07 $layer=POLY_cond $X=1.515 $Y=1.21
+ $X2=1.515 $Y2=0.74
r216 2 58 600 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=5.07
+ $Y=2.015 $X2=5.215 $Y2=2.16
r217 1 47 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=4.925
+ $Y=0.37 $X2=5.065 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__SDLCLKP_1%A_709_54# 1 2 9 12 13 15 16 18 20 21 23 24
+ 31 34 36 37 40 41 43 44 51 52 57
c131 52 0 1.28225e-19 $X=6.205 $Y=1.385
c132 51 0 1.17701e-19 $X=6.205 $Y=1.385
c133 37 0 2.48952e-19 $X=5.83 $Y=2.58
c134 24 0 2.5326e-19 $X=4.49 $Y=1.93
c135 9 0 8.55408e-20 $X=3.62 $Y=0.61
r136 52 61 57.0592 $w=3.21e-07 $l=3.8e-07 $layer=POLY_cond $X=6.205 $Y=1.385
+ $X2=6.585 $Y2=1.385
r137 52 59 13.514 $w=3.21e-07 $l=9e-08 $layer=POLY_cond $X=6.205 $Y=1.385
+ $X2=6.115 $Y2=1.385
r138 51 52 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.205
+ $Y=1.385 $X2=6.205 $Y2=1.385
r139 48 51 10.1275 $w=3.28e-07 $l=2.9e-07 $layer=LI1_cond $X=5.915 $Y=1.385
+ $X2=6.205 $Y2=1.385
r140 44 46 5.41299 $w=3.28e-07 $l=1.55e-07 $layer=LI1_cond $X=4.655 $Y=2.58
+ $X2=4.655 $Y2=2.735
r141 39 48 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.915 $Y=1.55
+ $X2=5.915 $Y2=1.385
r142 39 40 61.6524 $w=1.68e-07 $l=9.45e-07 $layer=LI1_cond $X=5.915 $Y=1.55
+ $X2=5.915 $Y2=2.495
r143 38 44 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.82 $Y=2.58
+ $X2=4.655 $Y2=2.58
r144 37 40 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.83 $Y=2.58
+ $X2=5.915 $Y2=2.495
r145 37 38 65.8931 $w=1.68e-07 $l=1.01e-06 $layer=LI1_cond $X=5.83 $Y=2.58
+ $X2=4.82 $Y2=2.58
r146 36 44 2.96841 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=4.655 $Y=2.495
+ $X2=4.655 $Y2=2.58
r147 35 43 6.99524 $w=2.6e-07 $l=1.9e-07 $layer=LI1_cond $X=4.655 $Y=2.12
+ $X2=4.655 $Y2=1.93
r148 35 36 13.0959 $w=3.28e-07 $l=3.75e-07 $layer=LI1_cond $X=4.655 $Y=2.12
+ $X2=4.655 $Y2=2.495
r149 34 43 6.99524 $w=2.6e-07 $l=2.22261e-07 $layer=LI1_cond $X=4.585 $Y=1.74
+ $X2=4.655 $Y2=1.93
r150 34 41 40.2775 $w=1.88e-07 $l=6.9e-07 $layer=LI1_cond $X=4.585 $Y=1.74
+ $X2=4.585 $Y2=1.05
r151 29 41 6.45386 $w=2.48e-07 $l=1.25e-07 $layer=LI1_cond $X=4.555 $Y=0.925
+ $X2=4.555 $Y2=1.05
r152 29 31 4.84026 $w=2.48e-07 $l=1.05e-07 $layer=LI1_cond $X=4.555 $Y=0.925
+ $X2=4.555 $Y2=0.82
r153 27 57 27.9778 $w=3.3e-07 $l=1.6e-07 $layer=POLY_cond $X=3.765 $Y=1.955
+ $X2=3.925 $Y2=1.955
r154 27 54 25.3549 $w=3.3e-07 $l=1.45e-07 $layer=POLY_cond $X=3.765 $Y=1.955
+ $X2=3.62 $Y2=1.955
r155 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.765
+ $Y=1.955 $X2=3.765 $Y2=1.955
r156 24 43 0.0189998 $w=3.8e-07 $l=1.65e-07 $layer=LI1_cond $X=4.49 $Y=1.93
+ $X2=4.655 $Y2=1.93
r157 24 26 21.9874 $w=3.78e-07 $l=7.25e-07 $layer=LI1_cond $X=4.49 $Y=1.93
+ $X2=3.765 $Y2=1.93
r158 21 23 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=6.585 $Y=1.94
+ $X2=6.585 $Y2=2.435
r159 20 21 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=6.585 $Y=1.85
+ $X2=6.585 $Y2=1.94
r160 19 61 16.2883 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=6.585 $Y=1.55
+ $X2=6.585 $Y2=1.385
r161 19 20 116.613 $w=1.8e-07 $l=3e-07 $layer=POLY_cond $X=6.585 $Y=1.55
+ $X2=6.585 $Y2=1.85
r162 16 59 20.5661 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.115 $Y=1.22
+ $X2=6.115 $Y2=1.385
r163 16 18 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=6.115 $Y=1.22
+ $X2=6.115 $Y2=0.79
r164 13 15 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=3.925 $Y=2.385
+ $X2=3.925 $Y2=2.67
r165 12 13 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=3.925 $Y=2.295
+ $X2=3.925 $Y2=2.385
r166 11 57 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=3.925 $Y=2.12
+ $X2=3.925 $Y2=1.955
r167 11 12 68.0242 $w=1.8e-07 $l=1.75e-07 $layer=POLY_cond $X=3.925 $Y=2.12
+ $X2=3.925 $Y2=2.295
r168 7 54 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.62 $Y=1.79
+ $X2=3.62 $Y2=1.955
r169 7 9 605.064 $w=1.5e-07 $l=1.18e-06 $layer=POLY_cond $X=3.62 $Y=1.79
+ $X2=3.62 $Y2=0.61
r170 2 46 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=4.505
+ $Y=1.76 $X2=4.655 $Y2=2.735
r171 2 43 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=4.505
+ $Y=1.76 $X2=4.655 $Y2=1.905
r172 1 31 182 $w=1.7e-07 $l=5.15267e-07 $layer=licon1_NDIFF $count=1 $X=4.375
+ $Y=0.37 $X2=4.515 $Y2=0.82
.ends

.subckt PM_SKY130_FD_SC_HS__SDLCLKP_1%A_566_74# 1 2 7 9 10 12 14 18 21 27 30 33
c78 27 0 3.05753e-20 $X=3.155 $Y=0.76
c79 10 0 8.61783e-20 $X=4.43 $Y=1.685
c80 7 0 1.99229e-19 $X=4.3 $Y=1.22
r81 30 31 5.76222 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=3.225 $Y=2.59
+ $X2=3.225 $Y2=2.425
r82 25 27 6.46067 $w=3.28e-07 $l=1.85e-07 $layer=LI1_cond $X=2.97 $Y=0.76
+ $X2=3.155 $Y2=0.76
r83 21 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.155
+ $Y=1.385 $X2=4.155 $Y2=1.385
r84 19 33 0.295496 $w=3.3e-07 $l=1.6e-07 $layer=LI1_cond $X=3.39 $Y=1.385
+ $X2=3.23 $Y2=1.385
r85 19 21 26.7157 $w=3.28e-07 $l=7.65e-07 $layer=LI1_cond $X=3.39 $Y=1.385
+ $X2=4.155 $Y2=1.385
r86 18 31 13.5052 $w=3.18e-07 $l=3.75e-07 $layer=LI1_cond $X=3.23 $Y=2.05
+ $X2=3.23 $Y2=2.425
r87 15 33 6.56857 $w=2.45e-07 $l=1.65e-07 $layer=LI1_cond $X=3.23 $Y=1.55
+ $X2=3.23 $Y2=1.385
r88 15 18 18.0069 $w=3.18e-07 $l=5e-07 $layer=LI1_cond $X=3.23 $Y=1.55 $X2=3.23
+ $Y2=2.05
r89 14 33 6.56857 $w=2.45e-07 $l=1.98997e-07 $layer=LI1_cond $X=3.155 $Y=1.22
+ $X2=3.23 $Y2=1.385
r90 13 27 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.155 $Y=0.925
+ $X2=3.155 $Y2=0.76
r91 13 14 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=3.155 $Y=0.925
+ $X2=3.155 $Y2=1.22
r92 10 22 55.3768 $w=4.28e-07 $l=3.77492e-07 $layer=POLY_cond $X=4.43 $Y=1.685
+ $X2=4.255 $Y2=1.385
r93 10 12 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=4.43 $Y=1.685
+ $X2=4.43 $Y2=2.32
r94 7 22 40.1736 $w=4.28e-07 $l=1.86145e-07 $layer=POLY_cond $X=4.3 $Y=1.22
+ $X2=4.255 $Y2=1.385
r95 7 9 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=4.3 $Y=1.22 $X2=4.3
+ $Y2=0.74
r96 2 30 600 $w=1.7e-07 $l=7.66339e-07 $layer=licon1_PDIFF $count=1 $X=3.075
+ $Y=1.895 $X2=3.225 $Y2=2.59
r97 2 18 600 $w=1.7e-07 $l=2.17428e-07 $layer=licon1_PDIFF $count=1 $X=3.075
+ $Y=1.895 $X2=3.225 $Y2=2.05
r98 1 25 182 $w=1.7e-07 $l=4.54643e-07 $layer=licon1_NDIFF $count=1 $X=2.83
+ $Y=0.37 $X2=2.97 $Y2=0.76
.ends

.subckt PM_SKY130_FD_SC_HS__SDLCLKP_1%CLK 3 5 7 10 12 13 14 16 17 23
c61 23 0 1.28225e-19 $X=5.495 $Y=1.52
c62 10 0 1.13508e-19 $X=5.755 $Y=0.79
r63 22 24 23.8705 $w=5.25e-07 $l=2.6e-07 $layer=POLY_cond $X=5.495 $Y=1.647
+ $X2=5.755 $Y2=1.647
r64 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.495
+ $Y=1.52 $X2=5.495 $Y2=1.52
r65 20 22 5.04952 $w=5.25e-07 $l=5.5e-08 $layer=POLY_cond $X=5.44 $Y=1.647
+ $X2=5.495 $Y2=1.647
r66 19 20 14.6895 $w=5.25e-07 $l=1.6e-07 $layer=POLY_cond $X=5.28 $Y=1.647
+ $X2=5.44 $Y2=1.647
r67 17 23 5.06376 $w=3.28e-07 $l=1.45e-07 $layer=LI1_cond $X=5.495 $Y=1.665
+ $X2=5.495 $Y2=1.52
r68 14 16 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=6.135 $Y=1.94
+ $X2=6.135 $Y2=2.435
r69 13 24 34.3153 $w=5.25e-07 $l=2.52733e-07 $layer=POLY_cond $X=5.83 $Y=1.865
+ $X2=5.755 $Y2=1.647
r70 12 14 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=6.06 $Y=1.865
+ $X2=6.135 $Y2=1.94
r71 12 13 117.936 $w=1.5e-07 $l=2.3e-07 $layer=POLY_cond $X=6.06 $Y=1.865
+ $X2=5.83 $Y2=1.865
r72 8 24 32.6451 $w=1.5e-07 $l=2.92e-07 $layer=POLY_cond $X=5.755 $Y=1.355
+ $X2=5.755 $Y2=1.647
r73 8 10 289.713 $w=1.5e-07 $l=5.65e-07 $layer=POLY_cond $X=5.755 $Y=1.355
+ $X2=5.755 $Y2=0.79
r74 5 20 32.6451 $w=1.5e-07 $l=2.93e-07 $layer=POLY_cond $X=5.44 $Y=1.94
+ $X2=5.44 $Y2=1.647
r75 5 7 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=5.44 $Y=1.94 $X2=5.44
+ $Y2=2.435
r76 1 19 32.6451 $w=1.5e-07 $l=2.92e-07 $layer=POLY_cond $X=5.28 $Y=1.355
+ $X2=5.28 $Y2=1.647
r77 1 3 315.351 $w=1.5e-07 $l=6.15e-07 $layer=POLY_cond $X=5.28 $Y=1.355
+ $X2=5.28 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HS__SDLCLKP_1%A_1238_94# 1 2 7 9 12 13 14 15 16 18 21 24
+ 25 28
c65 21 0 2.79353e-20 $X=6.56 $Y=1.3
c66 16 0 8.55731e-20 $X=6.36 $Y=1.89
c67 13 0 1.17701e-19 $X=7.09 $Y=1.36
c68 7 0 1.41593e-19 $X=7.09 $Y=1.765
r69 28 30 16.1243 $w=4.78e-07 $l=4.35e-07 $layer=LI1_cond $X=6.405 $Y=0.615
+ $X2=6.405 $Y2=1.05
r70 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.08
+ $Y=1.465 $X2=7.08 $Y2=1.465
r71 22 24 15.1913 $w=3.28e-07 $l=4.35e-07 $layer=LI1_cond $X=6.645 $Y=1.465
+ $X2=7.08 $Y2=1.465
r72 21 22 9.30874 $w=2.5e-07 $l=2.03101e-07 $layer=LI1_cond $X=6.56 $Y=1.3
+ $X2=6.475 $Y2=1.465
r73 21 30 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=6.56 $Y=1.3 $X2=6.56
+ $Y2=1.05
r74 16 22 16.4581 $w=3.3e-07 $l=4.79062e-07 $layer=LI1_cond $X=6.36 $Y=1.89
+ $X2=6.475 $Y2=1.465
r75 16 18 9.42908 $w=3.28e-07 $l=2.7e-07 $layer=LI1_cond $X=6.36 $Y=1.89
+ $X2=6.36 $Y2=2.16
r76 15 25 14.0139 $w=3.5e-07 $l=8.5e-08 $layer=POLY_cond $X=7.09 $Y=1.55
+ $X2=7.09 $Y2=1.465
r77 13 25 17.3113 $w=3.5e-07 $l=1.05e-07 $layer=POLY_cond $X=7.09 $Y=1.36
+ $X2=7.09 $Y2=1.465
r78 13 14 48.0802 $w=3.5e-07 $l=1.75e-07 $layer=POLY_cond $X=7.09 $Y=1.36
+ $X2=7.09 $Y2=1.185
r79 12 14 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=7.19 $Y=0.74
+ $X2=7.19 $Y2=1.185
r80 7 15 32.5881 $w=3.18e-07 $l=2.15e-07 $layer=POLY_cond $X=7.09 $Y=1.765
+ $X2=7.09 $Y2=1.55
r81 7 9 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=7.09 $Y=1.765
+ $X2=7.09 $Y2=2.4
r82 2 18 300 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=2 $X=6.21
+ $Y=2.015 $X2=6.36 $Y2=2.16
r83 1 28 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=6.19
+ $Y=0.47 $X2=6.33 $Y2=0.615
.ends

.subckt PM_SKY130_FD_SC_HS__SDLCLKP_1%VPWR 1 2 3 4 5 16 18 22 26 30 34 37 38 40
+ 41 42 44 49 68 69 75 78
c88 40 0 1.62774e-19 $X=6.695 $Y=3.33
r89 78 79 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r90 75 76 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r91 72 73 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r92 68 69 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r93 66 69 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=7.44 $Y2=3.33
r94 65 66 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r95 63 66 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=6.48 $Y2=3.33
r96 62 63 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r97 60 63 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=5.52 $Y2=3.33
r98 60 79 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=4.08 $Y2=3.33
r99 59 62 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=4.56 $Y=3.33 $X2=5.52
+ $Y2=3.33
r100 59 60 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r101 57 78 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.315 $Y=3.33
+ $X2=4.15 $Y2=3.33
r102 57 59 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=4.315 $Y=3.33
+ $X2=4.56 $Y2=3.33
r103 55 56 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r104 53 56 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=3.6 $Y2=3.33
r105 53 76 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.68 $Y2=3.33
r106 52 55 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=2.16 $Y=3.33
+ $X2=3.6 $Y2=3.33
r107 52 53 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r108 50 75 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.845 $Y=3.33
+ $X2=1.68 $Y2=3.33
r109 50 52 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=1.845 $Y=3.33
+ $X2=2.16 $Y2=3.33
r110 49 78 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.985 $Y=3.33
+ $X2=4.15 $Y2=3.33
r111 49 55 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=3.985 $Y=3.33
+ $X2=3.6 $Y2=3.33
r112 48 76 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=1.68 $Y2=3.33
r113 48 73 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.24 $Y2=3.33
r114 47 48 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r115 45 72 4.73185 $w=1.7e-07 $l=2.23e-07 $layer=LI1_cond $X=0.445 $Y=3.33
+ $X2=0.222 $Y2=3.33
r116 45 47 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=0.445 $Y=3.33
+ $X2=1.2 $Y2=3.33
r117 44 75 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.515 $Y=3.33
+ $X2=1.68 $Y2=3.33
r118 44 47 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=1.515 $Y=3.33
+ $X2=1.2 $Y2=3.33
r119 42 79 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=3.84 $Y=3.33
+ $X2=4.08 $Y2=3.33
r120 42 56 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=3.84 $Y=3.33
+ $X2=3.6 $Y2=3.33
r121 40 65 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=6.695 $Y=3.33
+ $X2=6.48 $Y2=3.33
r122 40 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.695 $Y=3.33
+ $X2=6.86 $Y2=3.33
r123 39 68 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=7.025 $Y=3.33
+ $X2=7.44 $Y2=3.33
r124 39 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.025 $Y=3.33
+ $X2=6.86 $Y2=3.33
r125 37 62 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=5.585 $Y=3.33
+ $X2=5.52 $Y2=3.33
r126 37 38 9.89127 $w=1.7e-07 $l=2.02e-07 $layer=LI1_cond $X=5.585 $Y=3.33
+ $X2=5.787 $Y2=3.33
r127 36 65 31.9679 $w=1.68e-07 $l=4.9e-07 $layer=LI1_cond $X=5.99 $Y=3.33
+ $X2=6.48 $Y2=3.33
r128 36 38 9.89127 $w=1.7e-07 $l=2.03e-07 $layer=LI1_cond $X=5.99 $Y=3.33
+ $X2=5.787 $Y2=3.33
r129 32 41 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.86 $Y=3.245
+ $X2=6.86 $Y2=3.33
r130 32 34 35.621 $w=3.28e-07 $l=1.02e-06 $layer=LI1_cond $X=6.86 $Y=3.245
+ $X2=6.86 $Y2=2.225
r131 28 38 1.50354 $w=4.05e-07 $l=8.5e-08 $layer=LI1_cond $X=5.787 $Y=3.245
+ $X2=5.787 $Y2=3.33
r132 28 30 6.97157 $w=4.03e-07 $l=2.45e-07 $layer=LI1_cond $X=5.787 $Y=3.245
+ $X2=5.787 $Y2=3
r133 24 78 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.15 $Y=3.245
+ $X2=4.15 $Y2=3.33
r134 24 26 20.0804 $w=3.28e-07 $l=5.75e-07 $layer=LI1_cond $X=4.15 $Y=3.245
+ $X2=4.15 $Y2=2.67
r135 20 75 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.68 $Y=3.245
+ $X2=1.68 $Y2=3.33
r136 20 22 14.6675 $w=3.28e-07 $l=4.2e-07 $layer=LI1_cond $X=1.68 $Y=3.245
+ $X2=1.68 $Y2=2.825
r137 16 72 3.03433 $w=3.3e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.28 $Y=3.245
+ $X2=0.222 $Y2=3.33
r138 16 18 33.1764 $w=3.28e-07 $l=9.5e-07 $layer=LI1_cond $X=0.28 $Y=3.245
+ $X2=0.28 $Y2=2.295
r139 5 34 300 $w=1.7e-07 $l=2.93428e-07 $layer=licon1_PDIFF $count=2 $X=6.66
+ $Y=2.015 $X2=6.86 $Y2=2.225
r140 4 30 600 $w=1.7e-07 $l=1.11183e-06 $layer=licon1_PDIFF $count=1 $X=5.515
+ $Y=2.015 $X2=5.785 $Y2=3
r141 3 26 600 $w=1.7e-07 $l=2.74955e-07 $layer=licon1_PDIFF $count=1 $X=4
+ $Y=2.46 $X2=4.15 $Y2=2.67
r142 2 22 600 $w=1.7e-07 $l=1.05501e-06 $layer=licon1_PDIFF $count=1 $X=1.535
+ $Y=1.84 $X2=1.68 $Y2=2.825
r143 1 18 300 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=2.12 $X2=0.28 $Y2=2.295
.ends

.subckt PM_SKY130_FD_SC_HS__SDLCLKP_1%A_114_112# 1 2 3 4 16 18 20 21 22 26 27 28
+ 31 33 35 39 40
r103 39 40 8.78489 $w=4.28e-07 $l=1.65e-07 $layer=LI1_cond $X=2.29 $Y=0.565
+ $X2=2.125 $Y2=0.565
r104 35 37 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=1.12 $Y=2.405
+ $X2=1.54 $Y2=2.405
r105 29 31 12.4464 $w=2.48e-07 $l=2.7e-07 $layer=LI1_cond $X=2.735 $Y=2.32
+ $X2=2.735 $Y2=2.05
r106 28 37 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=1.625 $Y=2.405
+ $X2=1.54 $Y2=2.405
r107 27 29 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=2.61 $Y=2.405
+ $X2=2.735 $Y2=2.32
r108 27 28 64.262 $w=1.68e-07 $l=9.85e-07 $layer=LI1_cond $X=2.61 $Y=2.405
+ $X2=1.625 $Y2=2.405
r109 26 37 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.54 $Y=2.32
+ $X2=1.54 $Y2=2.405
r110 25 26 56.107 $w=1.68e-07 $l=8.6e-07 $layer=LI1_cond $X=1.54 $Y=1.46
+ $X2=1.54 $Y2=2.32
r111 21 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.455 $Y=1.375
+ $X2=1.54 $Y2=1.46
r112 21 22 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=1.455 $Y=1.375
+ $X2=0.885 $Y2=1.375
r113 20 40 80.8984 $w=1.68e-07 $l=1.24e-06 $layer=LI1_cond $X=0.885 $Y=0.625
+ $X2=2.125 $Y2=0.625
r114 18 22 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.8 $Y=1.29
+ $X2=0.885 $Y2=1.375
r115 18 33 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=0.8 $Y=1.29 $X2=0.8
+ $Y2=1.12
r116 14 33 8.64139 $w=3.38e-07 $l=1.7e-07 $layer=LI1_cond $X=0.715 $Y=0.95
+ $X2=0.715 $Y2=1.12
r117 14 16 4.06745 $w=3.38e-07 $l=1.2e-07 $layer=LI1_cond $X=0.715 $Y=0.95
+ $X2=0.715 $Y2=0.83
r118 13 20 7.85115 $w=1.7e-07 $l=2.08207e-07 $layer=LI1_cond $X=0.715 $Y=0.71
+ $X2=0.885 $Y2=0.625
r119 13 16 4.06745 $w=3.38e-07 $l=1.2e-07 $layer=LI1_cond $X=0.715 $Y=0.71
+ $X2=0.715 $Y2=0.83
r120 4 31 300 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_PDIFF $count=2 $X=2.63
+ $Y=1.895 $X2=2.775 $Y2=2.05
r121 3 35 300 $w=1.7e-07 $l=3.52101e-07 $layer=licon1_PDIFF $count=2 $X=0.97
+ $Y=2.12 $X2=1.12 $Y2=2.405
r122 2 39 182 $w=1.7e-07 $l=2.57488e-07 $layer=licon1_NDIFF $count=1 $X=2.145
+ $Y=0.37 $X2=2.29 $Y2=0.565
r123 1 16 182 $w=1.7e-07 $l=3.32716e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.56 $X2=0.71 $Y2=0.83
.ends

.subckt PM_SKY130_FD_SC_HS__SDLCLKP_1%GCLK 1 2 9 13 14 15 16 23 32
c21 32 0 1.41593e-19 $X=7.41 $Y=1.82
r22 21 23 1.31708 $w=3.48e-07 $l=4e-08 $layer=LI1_cond $X=7.41 $Y=1.995 $X2=7.41
+ $Y2=2.035
r23 15 16 12.183 $w=3.48e-07 $l=3.7e-07 $layer=LI1_cond $X=7.41 $Y=2.405
+ $X2=7.41 $Y2=2.775
r24 14 21 0.75732 $w=3.48e-07 $l=2.3e-08 $layer=LI1_cond $X=7.41 $Y=1.972
+ $X2=7.41 $Y2=1.995
r25 14 32 8.06043 $w=3.48e-07 $l=1.52e-07 $layer=LI1_cond $X=7.41 $Y=1.972
+ $X2=7.41 $Y2=1.82
r26 14 15 11.4586 $w=3.48e-07 $l=3.48e-07 $layer=LI1_cond $X=7.41 $Y=2.057
+ $X2=7.41 $Y2=2.405
r27 14 23 0.724393 $w=3.48e-07 $l=2.2e-08 $layer=LI1_cond $X=7.41 $Y=2.057
+ $X2=7.41 $Y2=2.035
r28 13 32 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=7.5 $Y=1.13 $X2=7.5
+ $Y2=1.82
r29 7 13 8.71323 $w=3.43e-07 $l=1.72e-07 $layer=LI1_cond $X=7.412 $Y=0.958
+ $X2=7.412 $Y2=1.13
r30 7 9 14.798 $w=3.43e-07 $l=4.43e-07 $layer=LI1_cond $X=7.412 $Y=0.958
+ $X2=7.412 $Y2=0.515
r31 2 14 400 $w=1.7e-07 $l=2.98831e-07 $layer=licon1_PDIFF $count=1 $X=7.165
+ $Y=1.84 $X2=7.4 $Y2=1.985
r32 2 16 400 $w=1.7e-07 $l=1.08616e-06 $layer=licon1_PDIFF $count=1 $X=7.165
+ $Y=1.84 $X2=7.4 $Y2=2.815
r33 1 9 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=7.265
+ $Y=0.37 $X2=7.405 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__SDLCLKP_1%VGND 1 2 3 4 5 16 18 22 26 30 33 34 35 37
+ 49 56 63 64 71 77 80
r85 80 81 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=0 $X2=6.96
+ $Y2=0
r86 77 78 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r87 71 74 9.95292 $w=3.28e-07 $l=2.85e-07 $layer=LI1_cond $X=1.22 $Y=0 $X2=1.22
+ $Y2=0.285
r88 71 72 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r89 67 68 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r90 64 81 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=0 $X2=6.96
+ $Y2=0
r91 63 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=0 $X2=7.44
+ $Y2=0
r92 61 80 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.065 $Y=0 $X2=6.94
+ $Y2=0
r93 61 63 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=7.065 $Y=0 $X2=7.44
+ $Y2=0
r94 60 81 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=0 $X2=6.96
+ $Y2=0
r95 60 78 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.48 $Y=0 $X2=5.52
+ $Y2=0
r96 59 60 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.48 $Y=0 $X2=6.48
+ $Y2=0
r97 57 77 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.66 $Y=0 $X2=5.535
+ $Y2=0
r98 57 59 53.4973 $w=1.68e-07 $l=8.2e-07 $layer=LI1_cond $X=5.66 $Y=0 $X2=6.48
+ $Y2=0
r99 56 80 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.815 $Y=0 $X2=6.94
+ $Y2=0
r100 56 59 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=6.815 $Y=0
+ $X2=6.48 $Y2=0
r101 55 78 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=5.52
+ $Y2=0
r102 54 55 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r103 52 55 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=5.04
+ $Y2=0
r104 51 54 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=4.08 $Y=0 $X2=5.04
+ $Y2=0
r105 51 52 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r106 49 77 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.41 $Y=0 $X2=5.535
+ $Y2=0
r107 49 54 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=5.41 $Y=0 $X2=5.04
+ $Y2=0
r108 47 48 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r109 45 48 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=1.68 $Y=0 $X2=3.6
+ $Y2=0
r110 45 72 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r111 44 47 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=1.68 $Y=0 $X2=3.6
+ $Y2=0
r112 44 45 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.68 $Y=0
+ $X2=1.68 $Y2=0
r113 42 71 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.385 $Y=0 $X2=1.22
+ $Y2=0
r114 42 44 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=1.385 $Y=0 $X2=1.68
+ $Y2=0
r115 41 72 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r116 41 68 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r117 40 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r118 38 67 4.00981 $w=1.7e-07 $l=1.83e-07 $layer=LI1_cond $X=0.365 $Y=0
+ $X2=0.182 $Y2=0
r119 38 40 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=0.365 $Y=0
+ $X2=0.72 $Y2=0
r120 37 71 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.055 $Y=0 $X2=1.22
+ $Y2=0
r121 37 40 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=1.055 $Y=0
+ $X2=0.72 $Y2=0
r122 35 52 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=3.84 $Y=0
+ $X2=4.08 $Y2=0
r123 35 48 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=3.84 $Y=0 $X2=3.6
+ $Y2=0
r124 33 47 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=3.75 $Y=0 $X2=3.6
+ $Y2=0
r125 33 34 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.75 $Y=0 $X2=3.835
+ $Y2=0
r126 32 51 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=3.92 $Y=0 $X2=4.08
+ $Y2=0
r127 32 34 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.92 $Y=0 $X2=3.835
+ $Y2=0
r128 28 80 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.94 $Y=0.085
+ $X2=6.94 $Y2=0
r129 28 30 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=6.94 $Y=0.085
+ $X2=6.94 $Y2=0.515
r130 24 77 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.535 $Y=0.085
+ $X2=5.535 $Y2=0
r131 24 26 24.4318 $w=2.48e-07 $l=5.3e-07 $layer=LI1_cond $X=5.535 $Y=0.085
+ $X2=5.535 $Y2=0.615
r132 20 34 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.835 $Y=0.085
+ $X2=3.835 $Y2=0
r133 20 22 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=3.835 $Y=0.085
+ $X2=3.835 $Y2=0.545
r134 16 67 3.13335 $w=2.5e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.24 $Y=0.085
+ $X2=0.182 $Y2=0
r135 16 18 34.3428 $w=2.48e-07 $l=7.45e-07 $layer=LI1_cond $X=0.24 $Y=0.085
+ $X2=0.24 $Y2=0.83
r136 5 30 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=6.755
+ $Y=0.37 $X2=6.9 $Y2=0.515
r137 4 26 91 $w=1.7e-07 $l=3.07124e-07 $layer=licon1_NDIFF $count=2 $X=5.355
+ $Y=0.37 $X2=5.495 $Y2=0.615
r138 3 22 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=3.695
+ $Y=0.4 $X2=3.835 $Y2=0.545
r139 2 74 182 $w=1.7e-07 $l=3.68951e-07 $layer=licon1_NDIFF $count=1 $X=1
+ $Y=0.56 $X2=1.22 $Y2=0.285
r140 1 18 182 $w=1.7e-07 $l=3.34739e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.56 $X2=0.28 $Y2=0.83
.ends

