* File: sky130_fd_sc_hs__o31ai_4.spice
* Created: Thu Aug 27 21:03:10 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hs__o31ai_4.pex.spice"
.subckt sky130_fd_sc_hs__o31ai_4  VNB VPB A1 A2 A3 B1 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* B1	B1
* A3	A3
* A2	A2
* A1	A1
* VPB	VPB
* VNB	VNB
MM1000 N_VGND_M1000_d N_A1_M1000_g N_A_27_82#_M1000_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1295 AS=0.2109 PD=1.09 PS=2.05 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75007.9 A=0.111 P=1.78 MULT=1
MM1004 N_VGND_M1000_d N_A1_M1004_g N_A_27_82#_M1004_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1295 AS=0.1036 PD=1.09 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.7
+ SB=75007.4 A=0.111 P=1.78 MULT=1
MM1022 N_VGND_M1022_d N_A1_M1022_g N_A_27_82#_M1004_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1295 AS=0.1036 PD=1.09 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.1
+ SB=75006.9 A=0.111 P=1.78 MULT=1
MM1029 N_VGND_M1022_d N_A1_M1029_g N_A_27_82#_M1029_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1295 AS=0.1036 PD=1.09 PS=1.02 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75001.6
+ SB=75006.4 A=0.111 P=1.78 MULT=1
MM1001 N_VGND_M1001_d N_A2_M1001_g N_A_27_82#_M1029_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.2183 AS=0.1036 PD=1.33 PS=1.02 NRD=25.128 NRS=0 M=1 R=4.93333 SA=75002.1
+ SB=75006 A=0.111 P=1.78 MULT=1
MM1002 N_VGND_M1001_d N_A2_M1002_g N_A_27_82#_M1002_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.2183 AS=0.1295 PD=1.33 PS=1.09 NRD=25.128 NRS=0 M=1 R=4.93333 SA=75002.8
+ SB=75005.3 A=0.111 P=1.78 MULT=1
MM1005 N_VGND_M1005_d N_A2_M1005_g N_A_27_82#_M1002_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1295 PD=1.02 PS=1.09 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75003.3
+ SB=75004.8 A=0.111 P=1.78 MULT=1
MM1020 N_VGND_M1005_d N_A2_M1020_g N_A_27_82#_M1020_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75003.7
+ SB=75004.3 A=0.111 P=1.78 MULT=1
MM1006 N_A_27_82#_M1020_s N_A3_M1006_g N_VGND_M1006_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.3627 PD=1.02 PS=1.75 NRD=0 NRS=70.56 M=1 R=4.93333 SA=75004.2
+ SB=75003.9 A=0.111 P=1.78 MULT=1
MM1019 N_A_27_82#_M1019_d N_A3_M1019_g N_VGND_M1006_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.3627 PD=1.02 PS=1.75 NRD=0 NRS=70.56 M=1 R=4.93333 SA=75005.1
+ SB=75003 A=0.111 P=1.78 MULT=1
MM1023 N_A_27_82#_M1019_d N_A3_M1023_g N_VGND_M1023_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.201 PD=1.02 PS=1.42 NRD=0 NRS=35.124 M=1 R=4.93333 SA=75005.5
+ SB=75002.5 A=0.111 P=1.78 MULT=1
MM1026 N_A_27_82#_M1026_d N_A3_M1026_g N_VGND_M1023_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.201 PD=1.02 PS=1.42 NRD=0 NRS=35.124 M=1 R=4.93333 SA=75006.1
+ SB=75001.9 A=0.111 P=1.78 MULT=1
MM1018 N_Y_M1018_d N_B1_M1018_g N_A_27_82#_M1026_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75006.6
+ SB=75001.5 A=0.111 P=1.78 MULT=1
MM1021 N_Y_M1018_d N_B1_M1021_g N_A_27_82#_M1021_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75007
+ SB=75001.1 A=0.111 P=1.78 MULT=1
MM1024 N_Y_M1024_d N_B1_M1024_g N_A_27_82#_M1021_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75007.4
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1025 N_Y_M1024_d N_B1_M1025_g N_A_27_82#_M1025_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.2109 PD=1.02 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333 SA=75007.9
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1011 N_A_28_368#_M1011_d N_A1_M1011_g N_VPWR_M1011_s VPB PSHORT L=0.15 W=1.12
+ AD=0.3304 AS=0.168 PD=2.83 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75003.8 A=0.168 P=2.54 MULT=1
MM1012 N_A_28_368#_M1012_d N_A1_M1012_g N_VPWR_M1011_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.7 SB=75003.3 A=0.168 P=2.54 MULT=1
MM1013 N_A_28_368#_M1012_d N_A1_M1013_g N_VPWR_M1013_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.196 PD=1.42 PS=1.47 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.1 SB=75002.9 A=0.168 P=2.54 MULT=1
MM1014 N_A_28_368#_M1014_d N_A1_M1014_g N_VPWR_M1013_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.196 PD=1.42 PS=1.47 NRD=1.7533 NRS=10.5395 M=1 R=7.46667
+ SA=75001.6 SB=75002.4 A=0.168 P=2.54 MULT=1
MM1010 N_A_487_368#_M1010_d N_A2_M1010_g N_A_28_368#_M1014_d VPB PSHORT L=0.15
+ W=1.12 AD=0.196 AS=0.168 PD=1.47 PS=1.42 NRD=10.5395 NRS=1.7533 M=1 R=7.46667
+ SA=75002.1 SB=75001.9 A=0.168 P=2.54 MULT=1
MM1015 N_A_487_368#_M1010_d N_A2_M1015_g N_A_28_368#_M1015_s VPB PSHORT L=0.15
+ W=1.12 AD=0.196 AS=0.3192 PD=1.47 PS=1.69 NRD=1.7533 NRS=10.5395 M=1 R=7.46667
+ SA=75002.6 SB=75001.4 A=0.168 P=2.54 MULT=1
MM1016 N_A_487_368#_M1016_d N_A2_M1016_g N_A_28_368#_M1015_s VPB PSHORT L=0.15
+ W=1.12 AD=0.168 AS=0.3192 PD=1.42 PS=1.69 NRD=1.7533 NRS=40.4441 M=1 R=7.46667
+ SA=75003.3 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1017 N_A_487_368#_M1016_d N_A2_M1017_g N_A_28_368#_M1017_s VPB PSHORT L=0.15
+ W=1.12 AD=0.168 AS=0.3864 PD=1.42 PS=2.93 NRD=1.7533 NRS=10.5395 M=1 R=7.46667
+ SA=75003.7 SB=75000.3 A=0.168 P=2.54 MULT=1
MM1003 N_Y_M1003_d N_A3_M1003_g N_A_487_368#_M1003_s VPB PSHORT L=0.15 W=1.12
+ AD=0.3304 AS=0.168 PD=2.83 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75003.3 A=0.168 P=2.54 MULT=1
MM1007 N_Y_M1007_d N_A3_M1007_g N_A_487_368#_M1003_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.7 SB=75002.8 A=0.168 P=2.54 MULT=1
MM1009 N_Y_M1007_d N_A3_M1009_g N_A_487_368#_M1009_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.1 SB=75002.4 A=0.168 P=2.54 MULT=1
MM1027 N_Y_M1027_d N_A3_M1027_g N_A_487_368#_M1009_s VPB PSHORT L=0.15 W=1.12
+ AD=0.196 AS=0.168 PD=1.47 PS=1.42 NRD=10.5395 NRS=1.7533 M=1 R=7.46667
+ SA=75001.6 SB=75001.9 A=0.168 P=2.54 MULT=1
MM1008 N_VPWR_M1008_d N_B1_M1008_g N_Y_M1027_d VPB PSHORT L=0.15 W=1.12
+ AD=0.5852 AS=0.196 PD=2.165 PS=1.47 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75002.1 SB=75001.4 A=0.168 P=2.54 MULT=1
MM1028 N_VPWR_M1008_d N_B1_M1028_g N_Y_M1028_s VPB PSHORT L=0.15 W=1.12
+ AD=0.5852 AS=0.3304 PD=2.165 PS=2.83 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75003.3 SB=75000.2 A=0.168 P=2.54 MULT=1
DX30_noxref VNB VPB NWDIODE A=16.7772 P=21.76
*
.include "sky130_fd_sc_hs__o31ai_4.pxi.spice"
*
.ends
*
*
