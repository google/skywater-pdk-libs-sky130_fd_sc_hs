* File: sky130_fd_sc_hs__a221o_2.pex.spice
* Created: Thu Aug 27 20:25:42 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HS__A221O_2%A_89_260# 1 2 3 10 12 15 19 21 23 24 30 31
+ 32 34 35 36 37 38 41 47 55
c128 24 0 1.42045e-19 $X=1.025 $Y=1.465
c129 19 0 1.97451e-19 $X=0.985 $Y=0.74
r130 55 56 0.599503 $w=4.02e-07 $l=5e-09 $layer=POLY_cond $X=0.985 $Y=1.532
+ $X2=0.99 $Y2=1.532
r131 52 53 1.79851 $w=4.02e-07 $l=1.5e-08 $layer=POLY_cond $X=0.54 $Y=1.532
+ $X2=0.555 $Y2=1.532
r132 45 47 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=4.055 $Y=0.84
+ $X2=4.055 $Y2=0.515
r133 41 43 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=4.05 $Y=2.105
+ $X2=4.05 $Y2=2.815
r134 39 41 7.50834 $w=3.28e-07 $l=2.15e-07 $layer=LI1_cond $X=4.05 $Y=1.89
+ $X2=4.05 $Y2=2.105
r135 37 39 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.885 $Y=1.805
+ $X2=4.05 $Y2=1.89
r136 37 38 51.2139 $w=1.68e-07 $l=7.85e-07 $layer=LI1_cond $X=3.885 $Y=1.805
+ $X2=3.1 $Y2=1.805
r137 35 45 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.89 $Y=0.925
+ $X2=4.055 $Y2=0.84
r138 35 36 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=3.89 $Y=0.925
+ $X2=3.1 $Y2=0.925
r139 34 38 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.015 $Y=1.72
+ $X2=3.1 $Y2=1.805
r140 33 36 9.48932 $w=6.84e-07 $l=2.43824e-07 $layer=LI1_cond $X=3.015 $Y=1.13
+ $X2=3.1 $Y2=0.925
r141 33 50 5.17251 $w=6.84e-07 $l=5.14976e-07 $layer=LI1_cond $X=3.015 $Y=1.13
+ $X2=2.725 $Y2=0.74
r142 33 34 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=3.015 $Y=1.13
+ $X2=3.015 $Y2=1.72
r143 31 50 20.5478 $w=6.84e-07 $l=8.26952e-07 $layer=LI1_cond $X=2.02 $Y=1.005
+ $X2=2.725 $Y2=0.74
r144 31 32 53.8235 $w=1.68e-07 $l=8.25e-07 $layer=LI1_cond $X=2.02 $Y=1.005
+ $X2=1.195 $Y2=1.005
r145 29 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.11 $Y=1.09
+ $X2=1.195 $Y2=1.005
r146 29 30 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=1.11 $Y=1.09
+ $X2=1.11 $Y2=1.3
r147 27 55 4.19652 $w=4.02e-07 $l=3.5e-08 $layer=POLY_cond $X=0.95 $Y=1.532
+ $X2=0.985 $Y2=1.532
r148 27 53 47.3607 $w=4.02e-07 $l=3.95e-07 $layer=POLY_cond $X=0.95 $Y=1.532
+ $X2=0.555 $Y2=1.532
r149 26 27 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.95
+ $Y=1.465 $X2=0.95 $Y2=1.465
r150 24 30 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.025 $Y=1.465
+ $X2=1.11 $Y2=1.3
r151 24 26 2.61919 $w=3.28e-07 $l=7.5e-08 $layer=LI1_cond $X=1.025 $Y=1.465
+ $X2=0.95 $Y2=1.465
r152 21 56 25.9839 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=0.99 $Y=1.765
+ $X2=0.99 $Y2=1.532
r153 21 23 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.99 $Y=1.765
+ $X2=0.99 $Y2=2.4
r154 17 55 25.9839 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=0.985 $Y=1.3
+ $X2=0.985 $Y2=1.532
r155 17 19 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=0.985 $Y=1.3
+ $X2=0.985 $Y2=0.74
r156 13 53 25.9839 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=0.555 $Y=1.3
+ $X2=0.555 $Y2=1.532
r157 13 15 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=0.555 $Y=1.3
+ $X2=0.555 $Y2=0.74
r158 10 52 25.9839 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=0.54 $Y=1.765
+ $X2=0.54 $Y2=1.532
r159 10 12 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.54 $Y=1.765
+ $X2=0.54 $Y2=2.4
r160 3 43 400 $w=1.7e-07 $l=9.26971e-07 $layer=licon1_PDIFF $count=1 $X=3.9
+ $Y=1.96 $X2=4.05 $Y2=2.815
r161 3 41 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=3.9
+ $Y=1.96 $X2=4.05 $Y2=2.105
r162 2 47 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.915
+ $Y=0.37 $X2=4.055 $Y2=0.515
r163 1 50 45.5 $w=1.7e-07 $l=7.48999e-07 $layer=licon1_NDIFF $count=4 $X=2.045
+ $Y=0.37 $X2=2.725 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__A221O_2%A2 2 3 5 8 10 13 14
c45 14 0 3.97653e-20 $X=1.52 $Y=1.425
c46 13 0 1.38754e-19 $X=1.52 $Y=1.425
c47 2 0 3.12249e-19 $X=1.505 $Y=1.795
r48 13 16 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.52 $Y=1.425
+ $X2=1.52 $Y2=1.59
r49 13 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.52 $Y=1.425
+ $X2=1.52 $Y2=1.26
r50 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.52
+ $Y=1.425 $X2=1.52 $Y2=1.425
r51 10 14 6.91466 $w=3.98e-07 $l=2.4e-07 $layer=LI1_cond $X=1.565 $Y=1.665
+ $X2=1.565 $Y2=1.425
r52 8 15 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=1.61 $Y=0.74 $X2=1.61
+ $Y2=1.26
r53 3 5 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=1.505 $Y=1.885
+ $X2=1.505 $Y2=2.46
r54 2 3 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=1.505 $Y=1.795 $X2=1.505
+ $Y2=1.885
r55 2 16 79.6855 $w=1.8e-07 $l=2.05e-07 $layer=POLY_cond $X=1.505 $Y=1.795
+ $X2=1.505 $Y2=1.59
.ends

.subckt PM_SKY130_FD_SC_HS__A221O_2%A1 1 3 6 8
c33 8 0 3.08958e-19 $X=2.16 $Y=1.665
r34 8 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.08
+ $Y=1.615 $X2=2.08 $Y2=1.615
r35 4 11 38.5325 $w=3.12e-07 $l=2.03101e-07 $layer=POLY_cond $X=1.97 $Y=1.45
+ $X2=2.055 $Y2=1.615
r36 4 6 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=1.97 $Y=1.45 $X2=1.97
+ $Y2=0.74
r37 1 11 54.7537 $w=3.12e-07 $l=3.1607e-07 $layer=POLY_cond $X=1.955 $Y=1.885
+ $X2=2.055 $Y2=1.615
r38 1 3 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=1.955 $Y=1.885
+ $X2=1.955 $Y2=2.46
.ends

.subckt PM_SKY130_FD_SC_HS__A221O_2%B1 1 3 6 8 9 10
c44 10 0 2.05981e-19 $X=2.64 $Y=1.665
r45 10 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.62
+ $Y=1.615 $X2=2.62 $Y2=1.615
r46 8 13 37.5952 $w=3.3e-07 $l=2.15e-07 $layer=POLY_cond $X=2.835 $Y=1.615
+ $X2=2.62 $Y2=1.615
r47 8 9 5.03009 $w=3.3e-07 $l=1.13049e-07 $layer=POLY_cond $X=2.835 $Y=1.615
+ $X2=2.925 $Y2=1.667
r48 4 9 37.0704 $w=1.5e-07 $l=2.24375e-07 $layer=POLY_cond $X=2.94 $Y=1.45
+ $X2=2.925 $Y2=1.667
r49 4 6 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=2.94 $Y=1.45 $X2=2.94
+ $Y2=0.74
r50 1 9 37.0704 $w=1.5e-07 $l=2.18e-07 $layer=POLY_cond $X=2.925 $Y=1.885
+ $X2=2.925 $Y2=1.667
r51 1 3 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=2.925 $Y=1.885
+ $X2=2.925 $Y2=2.46
.ends

.subckt PM_SKY130_FD_SC_HS__A221O_2%B2 3 5 6 8 9 12 14
c40 14 0 2.7314e-20 $X=3.39 $Y=1.22
c41 5 0 6.88407e-20 $X=3.375 $Y=1.795
r42 12 15 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.39 $Y=1.385
+ $X2=3.39 $Y2=1.55
r43 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.39 $Y=1.385
+ $X2=3.39 $Y2=1.22
r44 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.39
+ $Y=1.385 $X2=3.39 $Y2=1.385
r45 9 13 6.54089 $w=3.68e-07 $l=2.1e-07 $layer=LI1_cond $X=3.6 $Y=1.365 $X2=3.39
+ $Y2=1.365
r46 6 8 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=3.375 $Y=1.885
+ $X2=3.375 $Y2=2.46
r47 5 6 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=3.375 $Y=1.795 $X2=3.375
+ $Y2=1.885
r48 5 15 95.2339 $w=1.8e-07 $l=2.45e-07 $layer=POLY_cond $X=3.375 $Y=1.795
+ $X2=3.375 $Y2=1.55
r49 3 14 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=3.3 $Y=0.74 $X2=3.3
+ $Y2=1.22
.ends

.subckt PM_SKY130_FD_SC_HS__A221O_2%C1 3 4 6 9 10 11 16
c30 11 0 2.7314e-20 $X=4.08 $Y=1.295
r31 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.03
+ $Y=1.385 $X2=4.03 $Y2=1.385
r32 13 16 33.2236 $w=3.3e-07 $l=1.9e-07 $layer=POLY_cond $X=3.84 $Y=1.385
+ $X2=4.03 $Y2=1.385
r33 11 17 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=4.03 $Y=1.295 $X2=4.03
+ $Y2=1.385
r34 9 10 41.3838 $w=1.65e-07 $l=9.5e-08 $layer=POLY_cond $X=3.832 $Y=1.79
+ $X2=3.832 $Y2=1.885
r35 7 13 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.84 $Y=1.55
+ $X2=3.84 $Y2=1.385
r36 7 9 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=3.84 $Y=1.55 $X2=3.84
+ $Y2=1.79
r37 4 13 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.84 $Y=1.22
+ $X2=3.84 $Y2=1.385
r38 4 6 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=3.84 $Y=1.22 $X2=3.84
+ $Y2=0.74
r39 3 10 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=3.825 $Y=2.46
+ $X2=3.825 $Y2=1.885
.ends

.subckt PM_SKY130_FD_SC_HS__A221O_2%VPWR 1 2 3 10 12 14 18 24 26 28 38 39 45 48
r59 45 46 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r60 43 46 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=1.2 $Y2=3.33
r61 42 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r62 38 39 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r63 36 39 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=4.08 $Y2=3.33
r64 35 38 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=2.64 $Y=3.33
+ $X2=4.08 $Y2=3.33
r65 35 36 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r66 33 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.345 $Y=3.33
+ $X2=2.18 $Y2=3.33
r67 33 35 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=2.345 $Y=3.33
+ $X2=2.64 $Y2=3.33
r68 32 46 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r69 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r70 29 45 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.38 $Y=3.33
+ $X2=1.255 $Y2=3.33
r71 29 31 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=1.38 $Y=3.33 $X2=1.68
+ $Y2=3.33
r72 28 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.015 $Y=3.33
+ $X2=2.18 $Y2=3.33
r73 28 31 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=2.015 $Y=3.33
+ $X2=1.68 $Y2=3.33
r74 26 36 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r75 26 32 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.68 $Y2=3.33
r76 26 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r77 22 48 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.18 $Y=3.245
+ $X2=2.18 $Y2=3.33
r78 22 24 30.3826 $w=3.28e-07 $l=8.7e-07 $layer=LI1_cond $X=2.18 $Y=3.245
+ $X2=2.18 $Y2=2.375
r79 18 21 32.2684 $w=2.48e-07 $l=7e-07 $layer=LI1_cond $X=1.255 $Y=2.115
+ $X2=1.255 $Y2=2.815
r80 16 45 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.255 $Y=3.245
+ $X2=1.255 $Y2=3.33
r81 16 21 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=1.255 $Y=3.245
+ $X2=1.255 $Y2=2.815
r82 15 42 3.96842 $w=1.7e-07 $l=2e-07 $layer=LI1_cond $X=0.4 $Y=3.33 $X2=0.2
+ $Y2=3.33
r83 14 45 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.13 $Y=3.33
+ $X2=1.255 $Y2=3.33
r84 14 15 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=1.13 $Y=3.33 $X2=0.4
+ $Y2=3.33
r85 10 42 3.17474 $w=2.5e-07 $l=1.16619e-07 $layer=LI1_cond $X=0.275 $Y=3.245
+ $X2=0.2 $Y2=3.33
r86 10 12 43.3319 $w=2.48e-07 $l=9.4e-07 $layer=LI1_cond $X=0.275 $Y=3.245
+ $X2=0.275 $Y2=2.305
r87 3 24 300 $w=1.7e-07 $l=4.84226e-07 $layer=licon1_PDIFF $count=2 $X=2.03
+ $Y=1.96 $X2=2.18 $Y2=2.375
r88 2 21 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=1.065
+ $Y=1.84 $X2=1.215 $Y2=2.815
r89 2 18 400 $w=1.7e-07 $l=3.4187e-07 $layer=licon1_PDIFF $count=1 $X=1.065
+ $Y=1.84 $X2=1.215 $Y2=2.115
r90 1 12 300 $w=1.7e-07 $l=5.23784e-07 $layer=licon1_PDIFF $count=2 $X=0.19
+ $Y=1.84 $X2=0.315 $Y2=2.305
.ends

.subckt PM_SKY130_FD_SC_HS__A221O_2%X 1 2 8 9 10 11 12 15 17 18 19 24 27
c46 9 0 1.57686e-19 $X=0.605 $Y=1.045
r47 24 27 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=0.765 $Y=1.97
+ $X2=0.765 $Y2=1.985
r48 18 19 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=0.765 $Y=2.405
+ $X2=0.765 $Y2=2.775
r49 17 24 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.765 $Y=1.885
+ $X2=0.765 $Y2=1.97
r50 17 18 12.5721 $w=3.28e-07 $l=3.6e-07 $layer=LI1_cond $X=0.765 $Y=2.045
+ $X2=0.765 $Y2=2.405
r51 17 27 2.09535 $w=3.28e-07 $l=6e-08 $layer=LI1_cond $X=0.765 $Y=2.045
+ $X2=0.765 $Y2=1.985
r52 13 15 20.5135 $w=2.48e-07 $l=4.45e-07 $layer=LI1_cond $X=0.73 $Y=0.96
+ $X2=0.73 $Y2=0.515
r53 11 17 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.6 $Y=1.885
+ $X2=0.765 $Y2=1.885
r54 11 12 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.6 $Y=1.885
+ $X2=0.335 $Y2=1.885
r55 9 13 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.605 $Y=1.045
+ $X2=0.73 $Y2=0.96
r56 9 10 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=0.605 $Y=1.045
+ $X2=0.335 $Y2=1.045
r57 8 12 7.04737 $w=1.7e-07 $l=1.54771e-07 $layer=LI1_cond $X=0.217 $Y=1.8
+ $X2=0.335 $Y2=1.885
r58 7 10 7.04737 $w=1.7e-07 $l=1.54771e-07 $layer=LI1_cond $X=0.217 $Y=1.13
+ $X2=0.335 $Y2=1.045
r59 7 8 32.8569 $w=2.33e-07 $l=6.7e-07 $layer=LI1_cond $X=0.217 $Y=1.13
+ $X2=0.217 $Y2=1.8
r60 2 19 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=0.615
+ $Y=1.84 $X2=0.765 $Y2=2.815
r61 2 27 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=0.615
+ $Y=1.84 $X2=0.765 $Y2=1.985
r62 1 15 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=0.63
+ $Y=0.37 $X2=0.77 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__A221O_2%A_316_392# 1 2 7 9 11 13 19 24
r42 19 21 6.42105 $w=1.88e-07 $l=1.1e-07 $layer=LI1_cond $X=2.635 $Y=2.035
+ $X2=2.635 $Y2=2.145
r43 14 21 1.386 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=2.73 $Y=2.145 $X2=2.635
+ $Y2=2.145
r44 13 24 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.985 $Y=2.145
+ $X2=3.15 $Y2=2.145
r45 13 14 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=2.985 $Y=2.145
+ $X2=2.73 $Y2=2.145
r46 12 18 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.815 $Y=2.035
+ $X2=1.69 $Y2=2.035
r47 11 19 1.386 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=2.54 $Y=2.035 $X2=2.635
+ $Y2=2.035
r48 11 12 47.2995 $w=1.68e-07 $l=7.25e-07 $layer=LI1_cond $X=2.54 $Y=2.035
+ $X2=1.815 $Y2=2.035
r49 7 18 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.69 $Y=2.12 $X2=1.69
+ $Y2=2.035
r50 7 9 32.0379 $w=2.48e-07 $l=6.95e-07 $layer=LI1_cond $X=1.69 $Y=2.12 $X2=1.69
+ $Y2=2.815
r51 2 24 300 $w=1.7e-07 $l=2.48948e-07 $layer=licon1_PDIFF $count=2 $X=3 $Y=1.96
+ $X2=3.15 $Y2=2.145
r52 1 18 400 $w=1.7e-07 $l=2.17428e-07 $layer=licon1_PDIFF $count=1 $X=1.58
+ $Y=1.96 $X2=1.73 $Y2=2.115
r53 1 9 400 $w=1.7e-07 $l=9.26971e-07 $layer=licon1_PDIFF $count=1 $X=1.58
+ $Y=1.96 $X2=1.73 $Y2=2.815
.ends

.subckt PM_SKY130_FD_SC_HS__A221O_2%A_515_392# 1 2 9 11 12 15
c30 9 0 1.3714e-19 $X=2.7 $Y=2.565
r31 13 15 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=3.6 $Y=2.905 $X2=3.6
+ $Y2=2.225
r32 11 13 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.515 $Y=2.99
+ $X2=3.6 $Y2=2.905
r33 11 12 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=3.515 $Y=2.99
+ $X2=2.785 $Y2=2.99
r34 7 12 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=2.66 $Y=2.905
+ $X2=2.785 $Y2=2.99
r35 7 9 15.6732 $w=2.48e-07 $l=3.4e-07 $layer=LI1_cond $X=2.66 $Y=2.905 $X2=2.66
+ $Y2=2.565
r36 2 15 300 $w=1.7e-07 $l=3.31625e-07 $layer=licon1_PDIFF $count=2 $X=3.45
+ $Y=1.96 $X2=3.6 $Y2=2.225
r37 1 9 600 $w=1.7e-07 $l=6.64568e-07 $layer=licon1_PDIFF $count=1 $X=2.575
+ $Y=1.96 $X2=2.7 $Y2=2.565
.ends

.subckt PM_SKY130_FD_SC_HS__A221O_2%VGND 1 2 3 10 12 16 20 22 24 29 39 40 46 49
r55 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r56 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r57 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r58 40 50 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=3.6
+ $Y2=0
r59 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r60 37 49 9.31531 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=3.72 $Y=0 $X2=3.535
+ $Y2=0
r61 37 39 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=3.72 $Y=0 $X2=4.08
+ $Y2=0
r62 36 50 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=3.6
+ $Y2=0
r63 35 36 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r64 33 47 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r65 32 35 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.68 $Y=0 $X2=3.12
+ $Y2=0
r66 32 33 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r67 30 46 11.6267 $w=1.7e-07 $l=2.63e-07 $layer=LI1_cond $X=1.56 $Y=0 $X2=1.297
+ $Y2=0
r68 30 32 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=1.56 $Y=0 $X2=1.68
+ $Y2=0
r69 29 49 9.31531 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=3.35 $Y=0 $X2=3.535
+ $Y2=0
r70 29 35 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=3.35 $Y=0 $X2=3.12
+ $Y2=0
r71 28 47 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r72 28 44 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r73 27 28 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r74 25 43 3.94169 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=0.425 $Y=0 $X2=0.212
+ $Y2=0
r75 25 27 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.425 $Y=0 $X2=0.72
+ $Y2=0
r76 24 46 11.6267 $w=1.7e-07 $l=2.62e-07 $layer=LI1_cond $X=1.035 $Y=0 $X2=1.297
+ $Y2=0
r77 24 27 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=1.035 $Y=0 $X2=0.72
+ $Y2=0
r78 22 36 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=3.12
+ $Y2=0
r79 22 33 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.68
+ $Y2=0
r80 18 49 1.24149 $w=3.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.535 $Y=0.085
+ $X2=3.535 $Y2=0
r81 18 20 14.4834 $w=3.68e-07 $l=4.65e-07 $layer=LI1_cond $X=3.535 $Y=0.085
+ $X2=3.535 $Y2=0.55
r82 14 46 2.19831 $w=5.25e-07 $l=8.5e-08 $layer=LI1_cond $X=1.297 $Y=0.085
+ $X2=1.297 $Y2=0
r83 14 16 11.9608 $w=5.23e-07 $l=5.25e-07 $layer=LI1_cond $X=1.297 $Y=0.085
+ $X2=1.297 $Y2=0.61
r84 10 43 3.20147 $w=2.5e-07 $l=1.23386e-07 $layer=LI1_cond $X=0.3 $Y=0.085
+ $X2=0.212 $Y2=0
r85 10 12 24.8928 $w=2.48e-07 $l=5.4e-07 $layer=LI1_cond $X=0.3 $Y=0.085 $X2=0.3
+ $Y2=0.625
r86 3 20 182 $w=1.7e-07 $l=2.47386e-07 $layer=licon1_NDIFF $count=1 $X=3.375
+ $Y=0.37 $X2=3.535 $Y2=0.55
r87 2 16 182 $w=1.7e-07 $l=3.37639e-07 $layer=licon1_NDIFF $count=1 $X=1.06
+ $Y=0.37 $X2=1.295 $Y2=0.61
r88 1 12 182 $w=1.7e-07 $l=3.11288e-07 $layer=licon1_NDIFF $count=1 $X=0.215
+ $Y=0.37 $X2=0.34 $Y2=0.625
.ends

