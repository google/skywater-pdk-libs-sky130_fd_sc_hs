* File: sky130_fd_sc_hs__nand4bb_2.spice
* Created: Tue Sep  1 20:10:31 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hs__nand4bb_2.pex.spice"
.subckt sky130_fd_sc_hs__nand4bb_2  VNB VPB A_N B_N C D VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* D	D
* C	C
* B_N	B_N
* A_N	A_N
* VPB	VPB
* VNB	VNB
MM1018 N_VGND_M1018_d N_A_N_M1018_g N_A_27_368#_M1018_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.1344 AS=0.1824 PD=1.06 PS=1.85 NRD=13.116 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75000.8 A=0.096 P=1.58 MULT=1
MM1001 N_A_231_74#_M1001_d N_B_N_M1001_g N_VGND_M1018_d VNB NLOWVT L=0.15 W=0.64
+ AD=0.1824 AS=0.1344 PD=1.85 PS=1.06 NRD=0 NRS=13.116 M=1 R=4.26667 SA=75000.8
+ SB=75000.2 A=0.096 P=1.58 MULT=1
MM1005 N_A_373_74#_M1005_d N_A_27_368#_M1005_g N_Y_M1005_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.2442 AS=0.11285 PD=2.14 PS=1.045 NRD=7.296 NRS=4.044 M=1 R=4.93333
+ SA=75000.3 SB=75001.7 A=0.111 P=1.78 MULT=1
MM1016 N_A_373_74#_M1016_d N_A_27_368#_M1016_g N_Y_M1005_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1773 AS=0.11285 PD=1.28 PS=1.045 NRD=13.776 NRS=0 M=1 R=4.93333
+ SA=75000.7 SB=75001.3 A=0.111 P=1.78 MULT=1
MM1000 N_A_373_74#_M1016_d N_A_231_74#_M1000_g N_A_678_74#_M1000_s VNB NLOWVT
+ L=0.15 W=0.74 AD=0.1773 AS=0.1036 PD=1.28 PS=1.02 NRD=13.776 NRS=0 M=1
+ R=4.93333 SA=75001.3 SB=75000.7 A=0.111 P=1.78 MULT=1
MM1013 N_A_373_74#_M1013_d N_A_231_74#_M1013_g N_A_678_74#_M1000_s VNB NLOWVT
+ L=0.15 W=0.74 AD=0.2516 AS=0.1036 PD=2.16 PS=1.02 NRD=4.044 NRS=0 M=1
+ R=4.93333 SA=75001.7 SB=75000.3 A=0.111 P=1.78 MULT=1
MM1010 N_A_886_74#_M1010_d N_C_M1010_g N_A_678_74#_M1010_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.2109 AS=0.1295 PD=2.05 PS=1.09 NRD=0 NRS=11.34 M=1 R=4.93333
+ SA=75000.2 SB=75001.6 A=0.111 P=1.78 MULT=1
MM1019 N_A_886_74#_M1019_d N_C_M1019_g N_A_678_74#_M1010_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.1295 PD=1.02 PS=1.09 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.7 SB=75001.1 A=0.111 P=1.78 MULT=1
MM1002 N_A_886_74#_M1019_d N_D_M1002_g N_VGND_M1002_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1295 PD=1.02 PS=1.09 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75001.1
+ SB=75000.7 A=0.111 P=1.78 MULT=1
MM1003 N_A_886_74#_M1003_d N_D_M1003_g N_VGND_M1002_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.1295 PD=2.05 PS=1.09 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.6
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1008 N_VPWR_M1008_d N_A_N_M1008_g N_A_27_368#_M1008_s VPB PSHORT L=0.15 W=1
+ AD=0.24225 AS=0.295 PD=1.52 PS=2.59 NRD=18.715 NRS=1.9503 M=1 R=6.66667
+ SA=75000.2 SB=75000.9 A=0.15 P=2.3 MULT=1
MM1007 N_A_231_74#_M1007_d N_B_N_M1007_g N_VPWR_M1008_d VPB PSHORT L=0.15 W=1
+ AD=0.395 AS=0.24225 PD=2.79 PS=1.52 NRD=11.8003 NRS=18.715 M=1 R=6.66667
+ SA=75000.8 SB=75000.3 A=0.15 P=2.3 MULT=1
MM1012 N_Y_M1012_d N_A_27_368#_M1012_g N_VPWR_M1012_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.3864 PD=1.42 PS=2.93 NRD=1.7533 NRS=10.5395 M=1 R=7.46667
+ SA=75000.3 SB=75004.1 A=0.168 P=2.54 MULT=1
MM1015 N_Y_M1012_d N_A_27_368#_M1015_g N_VPWR_M1015_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.224 PD=1.42 PS=1.52 NRD=1.7533 NRS=10.5395 M=1 R=7.46667
+ SA=75000.7 SB=75003.7 A=0.168 P=2.54 MULT=1
MM1011 N_Y_M1011_d N_A_231_74#_M1011_g N_VPWR_M1015_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.224 PD=1.42 PS=1.52 NRD=1.7533 NRS=10.5395 M=1 R=7.46667
+ SA=75001.3 SB=75003.1 A=0.168 P=2.54 MULT=1
MM1014 N_Y_M1011_d N_A_231_74#_M1014_g N_VPWR_M1014_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.4648 PD=1.42 PS=1.95 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.7 SB=75002.7 A=0.168 P=2.54 MULT=1
MM1004 N_Y_M1004_d N_C_M1004_g N_VPWR_M1014_s VPB PSHORT L=0.15 W=1.12 AD=0.168
+ AS=0.4648 PD=1.42 PS=1.95 NRD=1.7533 NRS=1.7533 M=1 R=7.46667 SA=75002.7
+ SB=75001.7 A=0.168 P=2.54 MULT=1
MM1009 N_Y_M1004_d N_C_M1009_g N_VPWR_M1009_s VPB PSHORT L=0.15 W=1.12 AD=0.168
+ AS=0.224 PD=1.42 PS=1.52 NRD=1.7533 NRS=10.5395 M=1 R=7.46667 SA=75003.1
+ SB=75001.3 A=0.168 P=2.54 MULT=1
MM1006 N_Y_M1006_d N_D_M1006_g N_VPWR_M1009_s VPB PSHORT L=0.15 W=1.12 AD=0.1904
+ AS=0.224 PD=1.46 PS=1.52 NRD=1.7533 NRS=10.5395 M=1 R=7.46667 SA=75003.7
+ SB=75000.7 A=0.168 P=2.54 MULT=1
MM1017 N_Y_M1006_d N_D_M1017_g N_VPWR_M1017_s VPB PSHORT L=0.15 W=1.12 AD=0.1904
+ AS=0.3416 PD=1.46 PS=2.85 NRD=8.7862 NRS=3.5066 M=1 R=7.46667 SA=75004.2
+ SB=75000.2 A=0.168 P=2.54 MULT=1
DX20_noxref VNB VPB NWDIODE A=13.206 P=17.92
*
.include "sky130_fd_sc_hs__nand4bb_2.pxi.spice"
*
.ends
*
*
