* File: sky130_fd_sc_hs__and3b_4.pex.spice
* Created: Thu Aug 27 20:32:55 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HS__AND3B_4%A_N 3 5 7 8
c31 8 0 1.93105e-19 $X=0.72 $Y=1.295
r32 8 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.67
+ $Y=1.345 $X2=0.67 $Y2=1.345
r33 5 11 72.8115 $w=3.63e-07 $l=5.01159e-07 $layer=POLY_cond $X=0.865 $Y=1.765
+ $X2=0.687 $Y2=1.345
r34 5 7 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=0.865 $Y=1.765
+ $X2=0.865 $Y2=2.34
r35 1 11 38.952 $w=3.63e-07 $l=2.61809e-07 $layer=POLY_cond $X=0.495 $Y=1.18
+ $X2=0.687 $Y2=1.345
r36 1 3 251.255 $w=1.5e-07 $l=4.9e-07 $layer=POLY_cond $X=0.495 $Y=1.18
+ $X2=0.495 $Y2=0.69
.ends

.subckt PM_SKY130_FD_SC_HS__AND3B_4%A_27_74# 1 2 7 9 12 14 16 19 23 26 27 28 31
+ 35 37 38 40 46
c86 46 0 1.93105e-19 $X=1.865 $Y=1.542
c87 19 0 4.59863e-20 $X=1.985 $Y=0.81
c88 14 0 1.18537e-19 $X=1.865 $Y=1.765
r89 45 46 41.9719 $w=3.56e-07 $l=3.1e-07 $layer=POLY_cond $X=1.555 $Y=1.542
+ $X2=1.865 $Y2=1.542
r90 44 45 18.9551 $w=3.56e-07 $l=1.4e-07 $layer=POLY_cond $X=1.415 $Y=1.542
+ $X2=1.555 $Y2=1.542
r91 41 44 7.44663 $w=3.56e-07 $l=5.5e-08 $layer=POLY_cond $X=1.36 $Y=1.542
+ $X2=1.415 $Y2=1.542
r92 40 41 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.36
+ $Y=1.485 $X2=1.36 $Y2=1.485
r93 36 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.805 $Y=1.765
+ $X2=0.64 $Y2=1.765
r94 35 40 11.1634 $w=3.06e-07 $l=3.64692e-07 $layer=LI1_cond $X=1.135 $Y=1.765
+ $X2=1.33 $Y2=1.485
r95 35 36 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=1.135 $Y=1.765
+ $X2=0.805 $Y2=1.765
r96 31 33 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=0.64 $Y=1.985
+ $X2=0.64 $Y2=2.695
r97 29 38 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.64 $Y=1.85 $X2=0.64
+ $Y2=1.765
r98 29 31 4.71454 $w=3.28e-07 $l=1.35e-07 $layer=LI1_cond $X=0.64 $Y=1.85
+ $X2=0.64 $Y2=1.985
r99 27 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.475 $Y=1.765
+ $X2=0.64 $Y2=1.765
r100 27 28 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=0.475 $Y=1.765
+ $X2=0.285 $Y2=1.765
r101 26 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.2 $Y=1.68
+ $X2=0.285 $Y2=1.765
r102 26 37 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=0.2 $Y=1.68 $X2=0.2
+ $Y2=1.01
r103 21 37 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=0.28 $Y=0.845
+ $X2=0.28 $Y2=1.01
r104 21 23 12.2229 $w=3.28e-07 $l=3.5e-07 $layer=LI1_cond $X=0.28 $Y=0.845
+ $X2=0.28 $Y2=0.495
r105 17 46 16.2472 $w=3.56e-07 $l=2.75543e-07 $layer=POLY_cond $X=1.985 $Y=1.32
+ $X2=1.865 $Y2=1.542
r106 17 19 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=1.985 $Y=1.32
+ $X2=1.985 $Y2=0.81
r107 14 46 23.0368 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=1.865 $Y=1.765
+ $X2=1.865 $Y2=1.542
r108 14 16 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=1.865 $Y=1.765
+ $X2=1.865 $Y2=2.34
r109 10 45 23.0368 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=1.555 $Y=1.32
+ $X2=1.555 $Y2=1.542
r110 10 12 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=1.555 $Y=1.32
+ $X2=1.555 $Y2=0.81
r111 7 44 23.0368 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=1.415 $Y=1.765
+ $X2=1.415 $Y2=1.542
r112 7 9 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=1.415 $Y=1.765
+ $X2=1.415 $Y2=2.34
r113 2 33 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=0.495
+ $Y=1.84 $X2=0.64 $Y2=2.695
r114 2 31 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.495
+ $Y=1.84 $X2=0.64 $Y2=1.985
r115 1 23 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_HS__AND3B_4%B 3 5 7 8 10 13 15 16 23
c56 16 0 1.18537e-19 $X=2.64 $Y=1.665
c57 13 0 7.05897e-20 $X=2.915 $Y=0.81
c58 8 0 1.52362e-19 $X=2.865 $Y=1.765
c59 5 0 8.80901e-20 $X=2.415 $Y=1.765
c60 3 0 1.67143e-19 $X=2.415 $Y=0.81
r61 23 24 6.5847 $w=3.66e-07 $l=5e-08 $layer=POLY_cond $X=2.865 $Y=1.557
+ $X2=2.915 $Y2=1.557
r62 21 23 49.3852 $w=3.66e-07 $l=3.75e-07 $layer=POLY_cond $X=2.49 $Y=1.557
+ $X2=2.865 $Y2=1.557
r63 21 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.49
+ $Y=1.515 $X2=2.49 $Y2=1.515
r64 19 21 9.87705 $w=3.66e-07 $l=7.5e-08 $layer=POLY_cond $X=2.415 $Y=1.557
+ $X2=2.49 $Y2=1.557
r65 16 22 4.02015 $w=4.28e-07 $l=1.5e-07 $layer=LI1_cond $X=2.64 $Y=1.565
+ $X2=2.49 $Y2=1.565
r66 15 22 8.84433 $w=4.28e-07 $l=3.3e-07 $layer=LI1_cond $X=2.16 $Y=1.565
+ $X2=2.49 $Y2=1.565
r67 11 24 23.7042 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.915 $Y=1.35
+ $X2=2.915 $Y2=1.557
r68 11 13 276.894 $w=1.5e-07 $l=5.4e-07 $layer=POLY_cond $X=2.915 $Y=1.35
+ $X2=2.915 $Y2=0.81
r69 8 23 23.7042 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=2.865 $Y=1.765
+ $X2=2.865 $Y2=1.557
r70 8 10 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=2.865 $Y=1.765
+ $X2=2.865 $Y2=2.34
r71 5 19 23.7042 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=2.415 $Y=1.765
+ $X2=2.415 $Y2=1.557
r72 5 7 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=2.415 $Y=1.765
+ $X2=2.415 $Y2=2.34
r73 1 19 23.7042 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.415 $Y=1.35
+ $X2=2.415 $Y2=1.557
r74 1 3 276.894 $w=1.5e-07 $l=5.4e-07 $layer=POLY_cond $X=2.415 $Y=1.35
+ $X2=2.415 $Y2=0.81
.ends

.subckt PM_SKY130_FD_SC_HS__AND3B_4%C 1 3 4 6 7 9 10 11 12 14 15 19
c58 19 0 1.52362e-19 $X=3.395 $Y=1.515
c59 7 0 8.87337e-20 $X=3.925 $Y=1.765
c60 4 0 1.44963e-19 $X=3.905 $Y=1.205
r61 21 22 1.87914 $w=5.13e-07 $l=2e-08 $layer=POLY_cond $X=3.905 $Y=1.485
+ $X2=3.925 $Y2=1.485
r62 20 21 40.4016 $w=5.13e-07 $l=4.3e-07 $layer=POLY_cond $X=3.475 $Y=1.485
+ $X2=3.905 $Y2=1.485
r63 18 20 7.51657 $w=5.13e-07 $l=8e-08 $layer=POLY_cond $X=3.395 $Y=1.485
+ $X2=3.475 $Y2=1.485
r64 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.395
+ $Y=1.515 $X2=3.395 $Y2=1.515
r65 15 19 7.37028 $w=4.28e-07 $l=2.75e-07 $layer=LI1_cond $X=3.12 $Y=1.565
+ $X2=3.395 $Y2=1.565
r66 12 14 133.353 $w=1.5e-07 $l=4.15e-07 $layer=POLY_cond $X=4.335 $Y=1.205
+ $X2=4.335 $Y2=0.79
r67 11 22 35.2164 $w=5.13e-07 $l=2.45917e-07 $layer=POLY_cond $X=4.015 $Y=1.28
+ $X2=3.925 $Y2=1.485
r68 10 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.26 $Y=1.28
+ $X2=4.335 $Y2=1.205
r69 10 11 125.628 $w=1.5e-07 $l=2.45e-07 $layer=POLY_cond $X=4.26 $Y=1.28
+ $X2=4.015 $Y2=1.28
r70 7 22 32.0577 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=3.925 $Y=1.765
+ $X2=3.925 $Y2=1.485
r71 7 9 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=3.925 $Y=1.765
+ $X2=3.925 $Y2=2.34
r72 4 21 32.0577 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=3.905 $Y=1.205
+ $X2=3.905 $Y2=1.485
r73 4 6 133.353 $w=1.5e-07 $l=4.15e-07 $layer=POLY_cond $X=3.905 $Y=1.205
+ $X2=3.905 $Y2=0.79
r74 1 20 32.0577 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=3.475 $Y=1.765
+ $X2=3.475 $Y2=1.485
r75 1 3 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=3.475 $Y=1.765
+ $X2=3.475 $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_HS__AND3B_4%A_298_368# 1 2 3 4 13 15 16 17 20 22 24 27
+ 29 31 34 36 38 41 45 49 53 57 59 63 66 68 71 74 78 79 82 84 86 87 95
c178 79 0 1.28172e-19 $X=1.67 $Y=1.82
c179 78 0 8.80901e-20 $X=1.64 $Y=1.985
c180 41 0 1.61033e-19 $X=6.225 $Y=0.74
c181 29 0 1.88161e-19 $X=5.51 $Y=1.765
c182 20 0 1.64454e-19 $X=4.845 $Y=0.74
r183 94 95 19.6856 $w=4.04e-07 $l=1.65e-07 $layer=POLY_cond $X=5.795 $Y=1.532
+ $X2=5.96 $Y2=1.532
r184 91 92 19.6856 $w=4.04e-07 $l=1.65e-07 $layer=POLY_cond $X=5.345 $Y=1.532
+ $X2=5.51 $Y2=1.532
r185 90 91 45.9332 $w=4.04e-07 $l=3.85e-07 $layer=POLY_cond $X=4.96 $Y=1.532
+ $X2=5.345 $Y2=1.532
r186 80 81 2.81784 $w=3.88e-07 $l=8.5e-08 $layer=LI1_cond $X=1.67 $Y=2.035
+ $X2=1.67 $Y2=2.12
r187 79 82 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.78 $Y=1.82
+ $X2=1.78 $Y2=1.15
r188 78 80 1.47749 $w=3.88e-07 $l=5e-08 $layer=LI1_cond $X=1.67 $Y=1.985
+ $X2=1.67 $Y2=2.035
r189 78 79 8.60763 $w=3.88e-07 $l=1.65e-07 $layer=LI1_cond $X=1.67 $Y=1.985
+ $X2=1.67 $Y2=1.82
r190 75 94 23.2649 $w=4.04e-07 $l=1.95e-07 $layer=POLY_cond $X=5.6 $Y=1.532
+ $X2=5.795 $Y2=1.532
r191 75 92 10.7376 $w=4.04e-07 $l=9e-08 $layer=POLY_cond $X=5.6 $Y=1.532
+ $X2=5.51 $Y2=1.532
r192 74 75 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=5.6
+ $Y=1.465 $X2=5.6 $Y2=1.465
r193 72 90 4.77228 $w=4.04e-07 $l=4e-08 $layer=POLY_cond $X=4.92 $Y=1.532
+ $X2=4.96 $Y2=1.532
r194 72 88 8.94802 $w=4.04e-07 $l=7.5e-08 $layer=POLY_cond $X=4.92 $Y=1.532
+ $X2=4.845 $Y2=1.532
r195 71 87 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=4.92 $Y=1.465
+ $X2=4.755 $Y2=1.465
r196 71 74 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=4.92 $Y=1.465
+ $X2=5.6 $Y2=1.465
r197 71 72 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=4.92
+ $Y=1.465 $X2=4.92 $Y2=1.465
r198 68 87 55.7807 $w=1.68e-07 $l=8.55e-07 $layer=LI1_cond $X=3.9 $Y=1.545
+ $X2=4.755 $Y2=1.545
r199 66 86 3.49088 $w=2.67e-07 $l=1.33918e-07 $layer=LI1_cond $X=3.815 $Y=1.95
+ $X2=3.717 $Y2=2.035
r200 65 68 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.815 $Y=1.63
+ $X2=3.9 $Y2=1.545
r201 65 66 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=3.815 $Y=1.63
+ $X2=3.815 $Y2=1.95
r202 61 86 3.49088 $w=2.67e-07 $l=8.5e-08 $layer=LI1_cond $X=3.717 $Y=2.12
+ $X2=3.717 $Y2=2.035
r203 61 63 18.7864 $w=3.63e-07 $l=5.95e-07 $layer=LI1_cond $X=3.717 $Y=2.12
+ $X2=3.717 $Y2=2.715
r204 60 84 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.805 $Y=2.035
+ $X2=2.64 $Y2=2.035
r205 59 86 3.01551 $w=1.7e-07 $l=1.82e-07 $layer=LI1_cond $X=3.535 $Y=2.035
+ $X2=3.717 $Y2=2.035
r206 59 60 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=3.535 $Y=2.035
+ $X2=2.805 $Y2=2.035
r207 55 84 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.64 $Y=2.12
+ $X2=2.64 $Y2=2.035
r208 55 57 20.7789 $w=3.28e-07 $l=5.95e-07 $layer=LI1_cond $X=2.64 $Y=2.12
+ $X2=2.64 $Y2=2.715
r209 54 80 5.6248 $w=1.7e-07 $l=1.95e-07 $layer=LI1_cond $X=1.865 $Y=2.035
+ $X2=1.67 $Y2=2.035
r210 53 84 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.475 $Y=2.035
+ $X2=2.64 $Y2=2.035
r211 53 54 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=2.475 $Y=2.035
+ $X2=1.865 $Y2=2.035
r212 47 82 5.59224 $w=1.78e-07 $l=9e-08 $layer=LI1_cond $X=1.775 $Y=1.06
+ $X2=1.775 $Y2=1.15
r213 47 49 11.7071 $w=1.78e-07 $l=1.9e-07 $layer=LI1_cond $X=1.775 $Y=1.06
+ $X2=1.775 $Y2=0.87
r214 45 81 20.0804 $w=3.28e-07 $l=5.75e-07 $layer=LI1_cond $X=1.64 $Y=2.695
+ $X2=1.64 $Y2=2.12
r215 39 95 31.6163 $w=4.04e-07 $l=3.62912e-07 $layer=POLY_cond $X=6.225 $Y=1.3
+ $X2=5.96 $Y2=1.532
r216 39 41 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=6.225 $Y=1.3
+ $X2=6.225 $Y2=0.74
r217 36 95 26.1054 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=5.96 $Y=1.765
+ $X2=5.96 $Y2=1.532
r218 36 38 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=5.96 $Y=1.765
+ $X2=5.96 $Y2=2.4
r219 32 94 26.1054 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=5.795 $Y=1.3
+ $X2=5.795 $Y2=1.532
r220 32 34 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=5.795 $Y=1.3
+ $X2=5.795 $Y2=0.74
r221 29 92 26.1054 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=5.51 $Y=1.765
+ $X2=5.51 $Y2=1.532
r222 29 31 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=5.51 $Y=1.765
+ $X2=5.51 $Y2=2.4
r223 25 91 26.1054 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=5.345 $Y=1.3
+ $X2=5.345 $Y2=1.532
r224 25 27 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=5.345 $Y=1.3
+ $X2=5.345 $Y2=0.74
r225 22 90 26.1054 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=4.96 $Y=1.765
+ $X2=4.96 $Y2=1.532
r226 22 24 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=4.96 $Y=1.765
+ $X2=4.96 $Y2=2.4
r227 18 88 26.1054 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=4.845 $Y=1.3
+ $X2=4.845 $Y2=1.532
r228 18 20 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=4.845 $Y=1.3
+ $X2=4.845 $Y2=0.74
r229 16 88 30.7166 $w=4.04e-07 $l=1.77381e-07 $layer=POLY_cond $X=4.755 $Y=1.67
+ $X2=4.845 $Y2=1.532
r230 16 17 79.4787 $w=1.5e-07 $l=1.55e-07 $layer=POLY_cond $X=4.755 $Y=1.67
+ $X2=4.6 $Y2=1.67
r231 13 17 26.9307 $w=1.5e-07 $l=1.32571e-07 $layer=POLY_cond $X=4.51 $Y=1.765
+ $X2=4.6 $Y2=1.67
r232 13 15 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=4.51 $Y=1.765
+ $X2=4.51 $Y2=2.4
r233 4 86 400 $w=1.7e-07 $l=2.59374e-07 $layer=licon1_PDIFF $count=1 $X=3.55
+ $Y=1.84 $X2=3.7 $Y2=2.035
r234 4 63 400 $w=1.7e-07 $l=9.47035e-07 $layer=licon1_PDIFF $count=1 $X=3.55
+ $Y=1.84 $X2=3.7 $Y2=2.715
r235 3 84 400 $w=1.7e-07 $l=2.59374e-07 $layer=licon1_PDIFF $count=1 $X=2.49
+ $Y=1.84 $X2=2.64 $Y2=2.035
r236 3 57 400 $w=1.7e-07 $l=9.47035e-07 $layer=licon1_PDIFF $count=1 $X=2.49
+ $Y=1.84 $X2=2.64 $Y2=2.715
r237 2 78 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=1.49
+ $Y=1.84 $X2=1.64 $Y2=1.985
r238 2 45 400 $w=1.7e-07 $l=9.26971e-07 $layer=licon1_PDIFF $count=1 $X=1.49
+ $Y=1.84 $X2=1.64 $Y2=2.695
r239 1 49 182 $w=1.7e-07 $l=4.44522e-07 $layer=licon1_NDIFF $count=1 $X=1.63
+ $Y=0.49 $X2=1.77 $Y2=0.87
.ends

.subckt PM_SKY130_FD_SC_HS__AND3B_4%VPWR 1 2 3 4 5 6 21 25 29 31 35 41 45 48 49
+ 51 52 53 55 60 65 78 79 82 85 88 91
c98 6 0 1.43861e-19 $X=6.035 $Y=1.84
r99 91 92 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r100 88 89 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r101 85 86 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r102 82 83 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r103 78 79 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r104 76 79 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=3.33 $X2=6.48
+ $Y2=3.33
r105 75 76 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r106 73 76 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.04 $Y=3.33 $X2=6
+ $Y2=3.33
r107 73 92 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=4.08 $Y2=3.33
r108 72 73 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r109 70 91 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.4 $Y=3.33
+ $X2=4.235 $Y2=3.33
r110 70 72 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=4.4 $Y=3.33 $X2=5.04
+ $Y2=3.33
r111 69 89 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r112 69 86 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=2.16 $Y2=3.33
r113 68 69 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r114 66 85 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.305 $Y=3.33
+ $X2=2.14 $Y2=3.33
r115 66 68 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=2.305 $Y=3.33
+ $X2=2.64 $Y2=3.33
r116 65 88 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.975 $Y=3.33
+ $X2=3.14 $Y2=3.33
r117 65 68 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=2.975 $Y=3.33
+ $X2=2.64 $Y2=3.33
r118 64 86 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r119 64 83 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r120 63 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r121 61 82 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.305 $Y=3.33
+ $X2=1.14 $Y2=3.33
r122 61 63 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=1.305 $Y=3.33
+ $X2=1.68 $Y2=3.33
r123 60 85 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.975 $Y=3.33
+ $X2=2.14 $Y2=3.33
r124 60 63 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=1.975 $Y=3.33
+ $X2=1.68 $Y2=3.33
r125 58 83 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r126 57 58 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r127 55 82 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.975 $Y=3.33
+ $X2=1.14 $Y2=3.33
r128 55 57 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.975 $Y=3.33
+ $X2=0.72 $Y2=3.33
r129 53 92 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=3.36 $Y=3.33
+ $X2=4.08 $Y2=3.33
r130 53 89 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=3.36 $Y=3.33
+ $X2=3.12 $Y2=3.33
r131 51 75 4.56684 $w=1.68e-07 $l=7e-08 $layer=LI1_cond $X=6.07 $Y=3.33 $X2=6
+ $Y2=3.33
r132 51 52 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.07 $Y=3.33
+ $X2=6.235 $Y2=3.33
r133 50 78 5.21925 $w=1.68e-07 $l=8e-08 $layer=LI1_cond $X=6.4 $Y=3.33 $X2=6.48
+ $Y2=3.33
r134 50 52 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.4 $Y=3.33
+ $X2=6.235 $Y2=3.33
r135 48 72 1.95722 $w=1.68e-07 $l=3e-08 $layer=LI1_cond $X=5.07 $Y=3.33 $X2=5.04
+ $Y2=3.33
r136 48 49 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.07 $Y=3.33
+ $X2=5.235 $Y2=3.33
r137 47 75 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=5.4 $Y=3.33 $X2=6
+ $Y2=3.33
r138 47 49 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.4 $Y=3.33
+ $X2=5.235 $Y2=3.33
r139 43 52 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.235 $Y=3.245
+ $X2=6.235 $Y2=3.33
r140 43 45 34.7479 $w=3.28e-07 $l=9.95e-07 $layer=LI1_cond $X=6.235 $Y=3.245
+ $X2=6.235 $Y2=2.25
r141 39 49 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.235 $Y=3.245
+ $X2=5.235 $Y2=3.33
r142 39 41 34.7479 $w=3.28e-07 $l=9.95e-07 $layer=LI1_cond $X=5.235 $Y=3.245
+ $X2=5.235 $Y2=2.25
r143 35 38 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=4.235 $Y=1.985
+ $X2=4.235 $Y2=2.815
r144 33 91 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.235 $Y=3.245
+ $X2=4.235 $Y2=3.33
r145 33 38 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=4.235 $Y=3.245
+ $X2=4.235 $Y2=2.815
r146 32 88 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.305 $Y=3.33
+ $X2=3.14 $Y2=3.33
r147 31 91 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.07 $Y=3.33
+ $X2=4.235 $Y2=3.33
r148 31 32 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=4.07 $Y=3.33
+ $X2=3.305 $Y2=3.33
r149 27 88 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.14 $Y=3.245
+ $X2=3.14 $Y2=3.33
r150 27 29 30.3826 $w=3.28e-07 $l=8.7e-07 $layer=LI1_cond $X=3.14 $Y=3.245
+ $X2=3.14 $Y2=2.375
r151 23 85 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.14 $Y=3.245
+ $X2=2.14 $Y2=3.33
r152 23 25 30.3826 $w=3.28e-07 $l=8.7e-07 $layer=LI1_cond $X=2.14 $Y=3.245
+ $X2=2.14 $Y2=2.375
r153 19 82 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.14 $Y=3.245
+ $X2=1.14 $Y2=3.33
r154 19 21 38.2402 $w=3.28e-07 $l=1.095e-06 $layer=LI1_cond $X=1.14 $Y=3.245
+ $X2=1.14 $Y2=2.15
r155 6 45 300 $w=1.7e-07 $l=5.001e-07 $layer=licon1_PDIFF $count=2 $X=6.035
+ $Y=1.84 $X2=6.235 $Y2=2.25
r156 5 41 300 $w=1.7e-07 $l=5.001e-07 $layer=licon1_PDIFF $count=2 $X=5.035
+ $Y=1.84 $X2=5.235 $Y2=2.25
r157 4 38 600 $w=1.7e-07 $l=1.08616e-06 $layer=licon1_PDIFF $count=1 $X=4
+ $Y=1.84 $X2=4.235 $Y2=2.815
r158 4 35 300 $w=1.7e-07 $l=2.98831e-07 $layer=licon1_PDIFF $count=2 $X=4
+ $Y=1.84 $X2=4.235 $Y2=1.985
r159 3 29 300 $w=1.7e-07 $l=6.27077e-07 $layer=licon1_PDIFF $count=2 $X=2.94
+ $Y=1.84 $X2=3.14 $Y2=2.375
r160 2 25 300 $w=1.7e-07 $l=6.27077e-07 $layer=licon1_PDIFF $count=2 $X=1.94
+ $Y=1.84 $X2=2.14 $Y2=2.375
r161 1 21 300 $w=1.7e-07 $l=3.97618e-07 $layer=licon1_PDIFF $count=2 $X=0.94
+ $Y=1.84 $X2=1.14 $Y2=2.15
.ends

.subckt PM_SKY130_FD_SC_HS__AND3B_4%X 1 2 3 4 15 19 20 23 25 26 29 35 38 39 41
+ 42 43
c85 42 0 1.61033e-19 $X=6.015 $Y=1.045
c86 41 0 1.43861e-19 $X=5.837 $Y=1.885
c87 38 0 1.88161e-19 $X=6.02 $Y=1.8
c88 20 0 8.87337e-20 $X=4.9 $Y=1.885
r89 43 48 11.0234 $w=2.28e-07 $l=2.2e-07 $layer=LI1_cond $X=6.48 $Y=1.665
+ $X2=6.48 $Y2=1.885
r90 40 41 4.30018 $w=1.7e-07 $l=2.68e-07 $layer=LI1_cond $X=6.105 $Y=1.885
+ $X2=5.837 $Y2=1.885
r91 39 48 2.50919 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=6.365 $Y=1.885
+ $X2=6.48 $Y2=1.885
r92 39 40 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=6.365 $Y=1.885
+ $X2=6.105 $Y2=1.885
r93 38 41 1.96316 $w=1.7e-07 $l=2.21459e-07 $layer=LI1_cond $X=6.02 $Y=1.8
+ $X2=5.837 $Y2=1.885
r94 37 42 5.04255 $w=1.75e-07 $l=8.74643e-08 $layer=LI1_cond $X=6.02 $Y=1.13
+ $X2=6.015 $Y2=1.045
r95 37 38 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=6.02 $Y=1.13
+ $X2=6.02 $Y2=1.8
r96 33 42 5.04255 $w=1.75e-07 $l=8.5e-08 $layer=LI1_cond $X=6.015 $Y=0.96
+ $X2=6.015 $Y2=1.045
r97 33 35 27.4192 $w=1.78e-07 $l=4.45e-07 $layer=LI1_cond $X=6.015 $Y=0.96
+ $X2=6.015 $Y2=0.515
r98 29 31 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=5.735 $Y=1.985
+ $X2=5.735 $Y2=2.815
r99 27 41 1.96316 $w=3.3e-07 $l=1.38109e-07 $layer=LI1_cond $X=5.735 $Y=1.97
+ $X2=5.837 $Y2=1.885
r100 27 29 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=5.735 $Y=1.97
+ $X2=5.735 $Y2=1.985
r101 25 42 1.44715 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=5.925 $Y=1.045
+ $X2=6.015 $Y2=1.045
r102 25 26 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=5.925 $Y=1.045
+ $X2=5.215 $Y2=1.045
r103 21 26 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=5.09 $Y=0.96
+ $X2=5.215 $Y2=1.045
r104 21 23 20.5135 $w=2.48e-07 $l=4.45e-07 $layer=LI1_cond $X=5.09 $Y=0.96
+ $X2=5.09 $Y2=0.515
r105 19 41 4.30018 $w=1.7e-07 $l=2.67e-07 $layer=LI1_cond $X=5.57 $Y=1.885
+ $X2=5.837 $Y2=1.885
r106 19 20 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.57 $Y=1.885
+ $X2=4.9 $Y2=1.885
r107 15 17 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=4.735 $Y=1.985
+ $X2=4.735 $Y2=2.815
r108 13 20 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.735 $Y=1.97
+ $X2=4.9 $Y2=1.885
r109 13 15 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=4.735 $Y=1.97
+ $X2=4.735 $Y2=1.985
r110 4 31 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=5.585
+ $Y=1.84 $X2=5.735 $Y2=2.815
r111 4 29 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=5.585
+ $Y=1.84 $X2=5.735 $Y2=1.985
r112 3 17 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=4.585
+ $Y=1.84 $X2=4.735 $Y2=2.815
r113 3 15 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=4.585
+ $Y=1.84 $X2=4.735 $Y2=1.985
r114 2 35 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=5.87
+ $Y=0.37 $X2=6.01 $Y2=0.515
r115 1 23 91 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=2 $X=4.92
+ $Y=0.37 $X2=5.13 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__AND3B_4%VGND 1 2 3 4 5 18 22 26 32 34 36 38 40 45 50
+ 55 60 66 69 72 75 79
c92 79 0 3.3892e-20 $X=6.48 $Y=0
r93 78 79 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=0 $X2=6.48
+ $Y2=0
r94 75 76 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r95 72 73 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r96 69 70 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r97 66 67 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r98 64 79 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=0 $X2=6.48
+ $Y2=0
r99 64 76 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=0 $X2=5.52
+ $Y2=0
r100 63 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=0 $X2=6 $Y2=0
r101 61 75 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.725 $Y=0 $X2=5.56
+ $Y2=0
r102 61 63 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=5.725 $Y=0 $X2=6
+ $Y2=0
r103 60 78 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=6.275 $Y=0
+ $X2=6.497 $Y2=0
r104 60 63 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=6.275 $Y=0 $X2=6
+ $Y2=0
r105 59 76 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=5.52
+ $Y2=0
r106 59 73 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=4.56
+ $Y2=0
r107 58 59 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r108 56 72 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.795 $Y=0 $X2=4.63
+ $Y2=0
r109 56 58 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=4.795 $Y=0 $X2=5.04
+ $Y2=0
r110 55 75 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.395 $Y=0 $X2=5.56
+ $Y2=0
r111 55 58 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=5.395 $Y=0
+ $X2=5.04 $Y2=0
r112 54 73 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=4.56
+ $Y2=0
r113 54 70 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=3.6
+ $Y2=0
r114 53 54 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r115 51 69 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.855 $Y=0 $X2=3.69
+ $Y2=0
r116 51 53 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=3.855 $Y=0
+ $X2=4.08 $Y2=0
r117 50 72 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.465 $Y=0 $X2=4.63
+ $Y2=0
r118 50 53 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=4.465 $Y=0
+ $X2=4.08 $Y2=0
r119 49 67 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r120 48 49 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r121 46 66 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=0.875 $Y=0 $X2=0.745
+ $Y2=0
r122 46 48 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.875 $Y=0 $X2=1.2
+ $Y2=0
r123 45 69 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.525 $Y=0 $X2=3.69
+ $Y2=0
r124 45 48 151.684 $w=1.68e-07 $l=2.325e-06 $layer=LI1_cond $X=3.525 $Y=0
+ $X2=1.2 $Y2=0
r125 43 67 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r126 42 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r127 40 66 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=0.615 $Y=0 $X2=0.745
+ $Y2=0
r128 40 42 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=0.615 $Y=0
+ $X2=0.24 $Y2=0
r129 38 70 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=3.36 $Y=0 $X2=3.6
+ $Y2=0
r130 38 49 0.602067 $w=4.9e-07 $l=2.16e-06 $layer=MET1_cond $X=3.36 $Y=0 $X2=1.2
+ $Y2=0
r131 34 78 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=6.44 $Y=0.085
+ $X2=6.497 $Y2=0
r132 34 36 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=6.44 $Y=0.085
+ $X2=6.44 $Y2=0.515
r133 30 75 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.56 $Y=0.085
+ $X2=5.56 $Y2=0
r134 30 32 18.8582 $w=3.28e-07 $l=5.4e-07 $layer=LI1_cond $X=5.56 $Y=0.085
+ $X2=5.56 $Y2=0.625
r135 26 28 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=4.63 $Y=0.515
+ $X2=4.63 $Y2=0.965
r136 24 72 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.63 $Y=0.085
+ $X2=4.63 $Y2=0
r137 24 26 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=4.63 $Y=0.085
+ $X2=4.63 $Y2=0.515
r138 20 69 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.69 $Y=0.085
+ $X2=3.69 $Y2=0
r139 20 22 20.6043 $w=3.28e-07 $l=5.9e-07 $layer=LI1_cond $X=3.69 $Y=0.085
+ $X2=3.69 $Y2=0.675
r140 16 66 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=0.745 $Y=0.085
+ $X2=0.745 $Y2=0
r141 16 18 18.1731 $w=2.58e-07 $l=4.1e-07 $layer=LI1_cond $X=0.745 $Y=0.085
+ $X2=0.745 $Y2=0.495
r142 5 36 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=6.3
+ $Y=0.37 $X2=6.44 $Y2=0.515
r143 4 32 182 $w=1.7e-07 $l=3.17372e-07 $layer=licon1_NDIFF $count=1 $X=5.42
+ $Y=0.37 $X2=5.56 $Y2=0.625
r144 3 28 182 $w=1.7e-07 $l=5.94916e-07 $layer=licon1_NDIFF $count=1 $X=4.41
+ $Y=0.47 $X2=4.63 $Y2=0.965
r145 3 26 182 $w=1.7e-07 $l=2.41454e-07 $layer=licon1_NDIFF $count=1 $X=4.41
+ $Y=0.47 $X2=4.63 $Y2=0.515
r146 2 22 182 $w=1.7e-07 $l=2.67862e-07 $layer=licon1_NDIFF $count=1 $X=3.545
+ $Y=0.47 $X2=3.69 $Y2=0.675
r147 1 18 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=0.57
+ $Y=0.37 $X2=0.71 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_HS__AND3B_4%A_239_98# 1 2 3 12 14 15 20 22 26
c45 26 0 7.05897e-20 $X=2.2 $Y=0.635
c46 20 0 1.20944e-20 $X=3.13 $Y=0.635
c47 14 0 3.89712e-20 $X=2.035 $Y=0.34
r48 24 26 1.3969 $w=3.28e-07 $l=4e-08 $layer=LI1_cond $X=2.2 $Y=0.595 $X2=2.2
+ $Y2=0.635
r49 22 24 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=2.2 $Y=0.34 $X2=2.2
+ $Y2=0.595
r50 18 24 2.36532 $w=2.5e-07 $l=1.65e-07 $layer=LI1_cond $X=2.365 $Y=0.595
+ $X2=2.2 $Y2=0.595
r51 18 20 35.2648 $w=2.48e-07 $l=7.65e-07 $layer=LI1_cond $X=2.365 $Y=0.595
+ $X2=3.13 $Y2=0.595
r52 14 22 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.035 $Y=0.34
+ $X2=2.2 $Y2=0.34
r53 14 15 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=2.035 $Y=0.34
+ $X2=1.505 $Y2=0.34
r54 10 15 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.34 $Y=0.425
+ $X2=1.505 $Y2=0.34
r55 10 12 7.33373 $w=3.28e-07 $l=2.1e-07 $layer=LI1_cond $X=1.34 $Y=0.425
+ $X2=1.34 $Y2=0.635
r56 3 20 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=2.99
+ $Y=0.49 $X2=3.13 $Y2=0.635
r57 2 26 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.06
+ $Y=0.49 $X2=2.2 $Y2=0.635
r58 1 12 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=1.195
+ $Y=0.49 $X2=1.34 $Y2=0.635
.ends

.subckt PM_SKY130_FD_SC_HS__AND3B_4%A_498_98# 1 2 7 11 14
c30 11 0 3.09417e-19 $X=4.12 $Y=0.615
r31 14 16 4.01609 $w=3.28e-07 $l=1.15e-07 $layer=LI1_cond $X=2.7 $Y=0.98 $X2=2.7
+ $Y2=1.095
r32 9 11 18.2086 $w=2.48e-07 $l=3.95e-07 $layer=LI1_cond $X=4.16 $Y=1.01
+ $X2=4.16 $Y2=0.615
r33 8 16 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.865 $Y=1.095
+ $X2=2.7 $Y2=1.095
r34 7 9 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=4.035 $Y=1.095
+ $X2=4.16 $Y2=1.01
r35 7 8 76.3316 $w=1.68e-07 $l=1.17e-06 $layer=LI1_cond $X=4.035 $Y=1.095
+ $X2=2.865 $Y2=1.095
r36 2 11 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.98
+ $Y=0.47 $X2=4.12 $Y2=0.615
r37 1 14 182 $w=1.7e-07 $l=5.85662e-07 $layer=licon1_NDIFF $count=1 $X=2.49
+ $Y=0.49 $X2=2.7 $Y2=0.98
.ends

