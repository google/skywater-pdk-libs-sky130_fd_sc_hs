* File: sky130_fd_sc_hs__clkbuf_16.spice
* Created: Tue Sep  1 19:57:30 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hs__clkbuf_16.pex.spice"
.subckt sky130_fd_sc_hs__clkbuf_16  VNB VPB A VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A	A
* VPB	VPB
* VNB	VNB
MM1000 N_A_114_74#_M1000_d N_A_M1000_g N_VGND_M1000_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.0588 AS=0.1197 PD=0.7 PS=1.41 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2 SB=75008.8
+ A=0.063 P=1.14 MULT=1
MM1028 N_A_114_74#_M1000_d N_A_M1028_g N_VGND_M1028_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.0588 AS=0.063 PD=0.7 PS=0.72 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6 SB=75008.4
+ A=0.063 P=1.14 MULT=1
MM1034 N_A_114_74#_M1034_d N_A_M1034_g N_VGND_M1028_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.0588 AS=0.063 PD=0.7 PS=0.72 NRD=0 NRS=5.712 M=1 R=2.8 SA=75001.1
+ SB=75007.9 A=0.063 P=1.14 MULT=1
MM1035 N_A_114_74#_M1034_d N_A_M1035_g N_VGND_M1035_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.0588 AS=0.0735 PD=0.7 PS=0.77 NRD=0 NRS=0 M=1 R=2.8 SA=75001.5 SB=75007.5
+ A=0.063 P=1.14 MULT=1
MM1001 N_VGND_M1035_s N_A_114_74#_M1001_g N_X_M1001_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.0735 AS=0.0588 PD=0.77 PS=0.7 NRD=19.992 NRS=0 M=1 R=2.8 SA=75002
+ SB=75007 A=0.063 P=1.14 MULT=1
MM1003 N_VGND_M1003_d N_A_114_74#_M1003_g N_X_M1001_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75002.4 SB=75006.6
+ A=0.063 P=1.14 MULT=1
MM1009 N_VGND_M1003_d N_A_114_74#_M1009_g N_X_M1009_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75002.9 SB=75006.1
+ A=0.063 P=1.14 MULT=1
MM1012 N_VGND_M1012_d N_A_114_74#_M1012_g N_X_M1009_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75003.3 SB=75005.7
+ A=0.063 P=1.14 MULT=1
MM1016 N_VGND_M1012_d N_A_114_74#_M1016_g N_X_M1016_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75003.7 SB=75005.3
+ A=0.063 P=1.14 MULT=1
MM1018 N_VGND_M1018_d N_A_114_74#_M1018_g N_X_M1016_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.0735 AS=0.0588 PD=0.77 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75004.2 SB=75004.9
+ A=0.063 P=1.14 MULT=1
MM1019 N_VGND_M1018_d N_A_114_74#_M1019_g N_X_M1019_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.0735 AS=0.0588 PD=0.77 PS=0.7 NRD=19.992 NRS=0 M=1 R=2.8 SA=75004.7
+ SB=75004.4 A=0.063 P=1.14 MULT=1
MM1020 N_VGND_M1020_d N_A_114_74#_M1020_g N_X_M1019_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.0735 AS=0.0588 PD=0.77 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75005.1 SB=75003.9
+ A=0.063 P=1.14 MULT=1
MM1022 N_VGND_M1020_d N_A_114_74#_M1022_g N_X_M1022_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.0735 AS=0.0588 PD=0.77 PS=0.7 NRD=19.992 NRS=0 M=1 R=2.8 SA=75005.6
+ SB=75003.4 A=0.063 P=1.14 MULT=1
MM1024 N_VGND_M1024_d N_A_114_74#_M1024_g N_X_M1022_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.0735 AS=0.0588 PD=0.77 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75006 SB=75003
+ A=0.063 P=1.14 MULT=1
MM1025 N_VGND_M1024_d N_A_114_74#_M1025_g N_X_M1025_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.0735 AS=0.0588 PD=0.77 PS=0.7 NRD=19.992 NRS=0 M=1 R=2.8 SA=75006.5
+ SB=75002.5 A=0.063 P=1.14 MULT=1
MM1026 N_VGND_M1026_d N_A_114_74#_M1026_g N_X_M1025_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.0735 AS=0.0588 PD=0.77 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75007 SB=75002.1
+ A=0.063 P=1.14 MULT=1
MM1031 N_VGND_M1026_d N_A_114_74#_M1031_g N_X_M1031_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.0735 AS=0.0588 PD=0.77 PS=0.7 NRD=19.992 NRS=0 M=1 R=2.8 SA=75007.5
+ SB=75001.6 A=0.063 P=1.14 MULT=1
MM1032 N_VGND_M1032_d N_A_114_74#_M1032_g N_X_M1031_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.0735 AS=0.0588 PD=0.77 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75007.9 SB=75001.1
+ A=0.063 P=1.14 MULT=1
MM1036 N_VGND_M1032_d N_A_114_74#_M1036_g N_X_M1036_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.0735 AS=0.0588 PD=0.77 PS=0.7 NRD=19.992 NRS=0 M=1 R=2.8 SA=75008.4
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1038 N_VGND_M1038_d N_A_114_74#_M1038_g N_X_M1036_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.1197 AS=0.0588 PD=1.41 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75008.8 SB=75000.2
+ A=0.063 P=1.14 MULT=1
MM1013 N_VPWR_M1013_d N_A_M1013_g N_A_114_74#_M1013_s VPB PSHORT L=0.15 W=1.12
+ AD=0.3304 AS=0.168 PD=2.83 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75008.8 A=0.168 P=2.54 MULT=1
MM1015 N_VPWR_M1015_d N_A_M1015_g N_A_114_74#_M1013_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.7 SB=75008.3 A=0.168 P=2.54 MULT=1
MM1017 N_VPWR_M1015_d N_A_M1017_g N_A_114_74#_M1017_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.1 SB=75007.9 A=0.168 P=2.54 MULT=1
MM1021 N_VPWR_M1021_d N_A_M1021_g N_A_114_74#_M1017_s VPB PSHORT L=0.15 W=1.12
+ AD=0.1736 AS=0.168 PD=1.43 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.6 SB=75007.4 A=0.168 P=2.54 MULT=1
MM1002 N_X_M1002_d N_A_114_74#_M1002_g N_VPWR_M1021_d VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.1736 PD=1.42 PS=1.43 NRD=1.7533 NRS=3.5066 M=1 R=7.46667
+ SA=75002 SB=75007 A=0.168 P=2.54 MULT=1
MM1004 N_X_M1002_d N_A_114_74#_M1004_g N_VPWR_M1004_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75002.5 SB=75006.5 A=0.168 P=2.54 MULT=1
MM1005 N_X_M1005_d N_A_114_74#_M1005_g N_VPWR_M1004_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75002.9 SB=75006.1 A=0.168 P=2.54 MULT=1
MM1006 N_X_M1005_d N_A_114_74#_M1006_g N_VPWR_M1006_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75003.4 SB=75005.6 A=0.168 P=2.54 MULT=1
MM1007 N_X_M1007_d N_A_114_74#_M1007_g N_VPWR_M1006_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75003.8 SB=75005.2 A=0.168 P=2.54 MULT=1
MM1008 N_X_M1007_d N_A_114_74#_M1008_g N_VPWR_M1008_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75004.3 SB=75004.7 A=0.168 P=2.54 MULT=1
MM1010 N_X_M1010_d N_A_114_74#_M1010_g N_VPWR_M1008_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75004.7 SB=75004.3 A=0.168 P=2.54 MULT=1
MM1011 N_X_M1010_d N_A_114_74#_M1011_g N_VPWR_M1011_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75005.2 SB=75003.8 A=0.168 P=2.54 MULT=1
MM1014 N_X_M1014_d N_A_114_74#_M1014_g N_VPWR_M1011_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75005.6 SB=75003.4 A=0.168 P=2.54 MULT=1
MM1023 N_X_M1014_d N_A_114_74#_M1023_g N_VPWR_M1023_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75006.1 SB=75002.9 A=0.168 P=2.54 MULT=1
MM1027 N_X_M1027_d N_A_114_74#_M1027_g N_VPWR_M1023_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75006.5 SB=75002.5 A=0.168 P=2.54 MULT=1
MM1029 N_X_M1027_d N_A_114_74#_M1029_g N_VPWR_M1029_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667 SA=75007
+ SB=75002 A=0.168 P=2.54 MULT=1
MM1030 N_X_M1030_d N_A_114_74#_M1030_g N_VPWR_M1029_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75007.4 SB=75001.6 A=0.168 P=2.54 MULT=1
MM1033 N_X_M1030_d N_A_114_74#_M1033_g N_VPWR_M1033_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.1792 PD=1.42 PS=1.44 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75007.9 SB=75001.1 A=0.168 P=2.54 MULT=1
MM1037 N_X_M1037_d N_A_114_74#_M1037_g N_VPWR_M1033_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.1792 PD=1.42 PS=1.44 NRD=1.7533 NRS=5.2599 M=1 R=7.46667
+ SA=75008.3 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1039 N_X_M1037_d N_A_114_74#_M1039_g N_VPWR_M1039_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.3304 PD=1.42 PS=2.83 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75008.8 SB=75000.2 A=0.168 P=2.54 MULT=1
DX40_noxref VNB VPB NWDIODE A=18.5628 P=23.68
*
.include "sky130_fd_sc_hs__clkbuf_16.pxi.spice"
*
.ends
*
*
