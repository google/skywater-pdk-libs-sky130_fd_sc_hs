* File: sky130_fd_sc_hs__xnor3_4.pxi.spice
* Created: Tue Sep  1 20:25:42 2020
* 
x_PM_SKY130_FD_SC_HS__XNOR3_4%A_75_227# N_A_75_227#_M1002_d N_A_75_227#_M1011_d
+ N_A_75_227#_M1023_d N_A_75_227#_M1009_d N_A_75_227#_c_190_n
+ N_A_75_227#_c_200_n N_A_75_227#_M1026_g N_A_75_227#_M1016_g
+ N_A_75_227#_c_191_n N_A_75_227#_c_192_n N_A_75_227#_c_210_p
+ N_A_75_227#_c_261_p N_A_75_227#_c_211_p N_A_75_227#_c_202_n
+ N_A_75_227#_c_217_p N_A_75_227#_c_203_n N_A_75_227#_c_204_n
+ N_A_75_227#_c_193_n N_A_75_227#_c_194_n N_A_75_227#_c_195_n
+ N_A_75_227#_c_196_n N_A_75_227#_c_197_n N_A_75_227#_c_205_n
+ N_A_75_227#_c_198_n PM_SKY130_FD_SC_HS__XNOR3_4%A_75_227#
x_PM_SKY130_FD_SC_HS__XNOR3_4%A N_A_c_324_n N_A_M1023_g N_A_M1002_g A
+ N_A_c_326_n PM_SKY130_FD_SC_HS__XNOR3_4%A
x_PM_SKY130_FD_SC_HS__XNOR3_4%A_386_23# N_A_386_23#_M1021_s N_A_386_23#_M1022_s
+ N_A_386_23#_M1006_g N_A_386_23#_c_369_n N_A_386_23#_c_370_n
+ N_A_386_23#_c_371_n N_A_386_23#_c_372_n N_A_386_23#_c_381_n
+ N_A_386_23#_M1019_g N_A_386_23#_M1011_g N_A_386_23#_c_374_n
+ N_A_386_23#_M1009_g N_A_386_23#_c_375_n N_A_386_23#_c_376_n
+ N_A_386_23#_c_384_n N_A_386_23#_c_377_n N_A_386_23#_c_378_n
+ N_A_386_23#_c_385_n N_A_386_23#_c_386_n N_A_386_23#_c_379_n
+ PM_SKY130_FD_SC_HS__XNOR3_4%A_386_23#
x_PM_SKY130_FD_SC_HS__XNOR3_4%B N_B_M1025_g N_B_c_503_n N_B_c_504_n N_B_c_497_n
+ N_B_M1007_g N_B_c_507_n N_B_c_508_n N_B_M1004_g N_B_c_509_n N_B_c_510_n
+ N_B_M1020_g N_B_c_512_n N_B_c_513_n N_B_M1021_g N_B_c_514_n N_B_M1022_g
+ N_B_c_500_n N_B_c_516_n B N_B_c_501_n N_B_c_502_n
+ PM_SKY130_FD_SC_HS__XNOR3_4%B
x_PM_SKY130_FD_SC_HS__XNOR3_4%A_1024_300# N_A_1024_300#_M1017_s
+ N_A_1024_300#_M1018_s N_A_1024_300#_M1027_g N_A_1024_300#_c_650_n
+ N_A_1024_300#_M1000_g N_A_1024_300#_c_651_n N_A_1024_300#_c_652_n
+ N_A_1024_300#_c_658_n N_A_1024_300#_c_653_n N_A_1024_300#_c_654_n
+ N_A_1024_300#_c_655_n N_A_1024_300#_c_661_n
+ PM_SKY130_FD_SC_HS__XNOR3_4%A_1024_300#
x_PM_SKY130_FD_SC_HS__XNOR3_4%C N_C_M1012_g N_C_c_732_n N_C_c_739_n N_C_M1024_g
+ N_C_c_733_n N_C_c_734_n N_C_c_735_n N_C_M1017_g N_C_c_736_n N_C_M1018_g C
+ N_C_c_737_n PM_SKY130_FD_SC_HS__XNOR3_4%C
x_PM_SKY130_FD_SC_HS__XNOR3_4%A_1057_74# N_A_1057_74#_M1027_d
+ N_A_1057_74#_M1000_d N_A_1057_74#_c_820_n N_A_1057_74#_M1005_g
+ N_A_1057_74#_c_806_n N_A_1057_74#_M1001_g N_A_1057_74#_c_821_n
+ N_A_1057_74#_M1008_g N_A_1057_74#_c_807_n N_A_1057_74#_M1003_g
+ N_A_1057_74#_c_822_n N_A_1057_74#_M1010_g N_A_1057_74#_c_808_n
+ N_A_1057_74#_M1013_g N_A_1057_74#_c_823_n N_A_1057_74#_M1015_g
+ N_A_1057_74#_c_809_n N_A_1057_74#_M1014_g N_A_1057_74#_c_810_n
+ N_A_1057_74#_c_811_n N_A_1057_74#_c_812_n N_A_1057_74#_c_824_n
+ N_A_1057_74#_c_813_n N_A_1057_74#_c_814_n N_A_1057_74#_c_815_n
+ N_A_1057_74#_c_932_p N_A_1057_74#_c_846_n N_A_1057_74#_c_848_n
+ N_A_1057_74#_c_825_n N_A_1057_74#_c_816_n N_A_1057_74#_c_826_n
+ N_A_1057_74#_c_866_p N_A_1057_74#_c_827_n N_A_1057_74#_c_861_p
+ N_A_1057_74#_c_817_n N_A_1057_74#_c_818_n N_A_1057_74#_c_819_n
+ PM_SKY130_FD_SC_HS__XNOR3_4%A_1057_74#
x_PM_SKY130_FD_SC_HS__XNOR3_4%A_27_373# N_A_27_373#_M1016_s N_A_27_373#_M1006_d
+ N_A_27_373#_M1026_s N_A_27_373#_M1019_d N_A_27_373#_c_965_n
+ N_A_27_373#_c_971_n N_A_27_373#_c_972_n N_A_27_373#_c_966_n
+ N_A_27_373#_c_973_n N_A_27_373#_c_967_n N_A_27_373#_c_968_n
+ N_A_27_373#_c_969_n N_A_27_373#_c_975_n N_A_27_373#_c_996_n
+ N_A_27_373#_c_1003_n N_A_27_373#_c_1006_n N_A_27_373#_c_970_n
+ N_A_27_373#_c_977_n PM_SKY130_FD_SC_HS__XNOR3_4%A_27_373#
x_PM_SKY130_FD_SC_HS__XNOR3_4%VPWR N_VPWR_M1026_d N_VPWR_M1022_d N_VPWR_M1018_d
+ N_VPWR_M1008_s N_VPWR_M1015_s N_VPWR_c_1078_n N_VPWR_c_1079_n N_VPWR_c_1080_n
+ N_VPWR_c_1081_n N_VPWR_c_1082_n N_VPWR_c_1083_n N_VPWR_c_1084_n
+ N_VPWR_c_1085_n N_VPWR_c_1147_n VPWR N_VPWR_c_1086_n N_VPWR_c_1087_n
+ N_VPWR_c_1088_n N_VPWR_c_1089_n N_VPWR_c_1090_n N_VPWR_c_1091_n
+ N_VPWR_c_1092_n N_VPWR_c_1093_n N_VPWR_c_1077_n
+ PM_SKY130_FD_SC_HS__XNOR3_4%VPWR
x_PM_SKY130_FD_SC_HS__XNOR3_4%A_324_373# N_A_324_373#_M1004_d
+ N_A_324_373#_M1012_d N_A_324_373#_M1007_d N_A_324_373#_M1000_s
+ N_A_324_373#_c_1192_n N_A_324_373#_c_1184_n N_A_324_373#_c_1185_n
+ N_A_324_373#_c_1186_n N_A_324_373#_c_1187_n N_A_324_373#_c_1188_n
+ N_A_324_373#_c_1189_n N_A_324_373#_c_1190_n N_A_324_373#_c_1210_n
+ N_A_324_373#_c_1191_n N_A_324_373#_c_1195_n N_A_324_373#_c_1219_n
+ N_A_324_373#_c_1196_n N_A_324_373#_c_1197_n N_A_324_373#_c_1220_n
+ PM_SKY130_FD_SC_HS__XNOR3_4%A_324_373#
x_PM_SKY130_FD_SC_HS__XNOR3_4%A_321_77# N_A_321_77#_M1025_d N_A_321_77#_M1027_s
+ N_A_321_77#_M1020_d N_A_321_77#_M1024_d N_A_321_77#_c_1312_n
+ N_A_321_77#_c_1339_n N_A_321_77#_c_1318_n N_A_321_77#_c_1329_n
+ N_A_321_77#_c_1313_n N_A_321_77#_c_1320_n N_A_321_77#_c_1321_n
+ N_A_321_77#_c_1314_n N_A_321_77#_c_1315_n N_A_321_77#_c_1316_n
+ N_A_321_77#_c_1317_n N_A_321_77#_c_1387_n
+ PM_SKY130_FD_SC_HS__XNOR3_4%A_321_77#
x_PM_SKY130_FD_SC_HS__XNOR3_4%X N_X_M1001_d N_X_M1013_d N_X_M1005_d N_X_M1010_d
+ N_X_c_1446_n N_X_c_1443_n N_X_c_1444_n N_X_c_1459_n N_X_c_1447_n N_X_c_1448_n
+ N_X_c_1469_n N_X_c_1472_n X X X X X X X X PM_SKY130_FD_SC_HS__XNOR3_4%X
x_PM_SKY130_FD_SC_HS__XNOR3_4%VGND N_VGND_M1016_d N_VGND_M1021_d N_VGND_M1017_d
+ N_VGND_M1003_s N_VGND_M1014_s N_VGND_c_1501_n N_VGND_c_1502_n N_VGND_c_1503_n
+ N_VGND_c_1553_n N_VGND_c_1504_n N_VGND_c_1505_n N_VGND_c_1506_n
+ N_VGND_c_1507_n N_VGND_c_1508_n VGND N_VGND_c_1509_n N_VGND_c_1510_n
+ N_VGND_c_1511_n N_VGND_c_1512_n N_VGND_c_1513_n N_VGND_c_1514_n
+ PM_SKY130_FD_SC_HS__XNOR3_4%VGND
cc_1 VNB N_A_75_227#_c_190_n 0.0109153f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.7
cc_2 VNB N_A_75_227#_c_191_n 0.00126892f $X=-0.19 $Y=-0.245 $X2=0.62 $Y2=1.95
cc_3 VNB N_A_75_227#_c_192_n 0.0202598f $X=-0.19 $Y=-0.245 $X2=1.175 $Y2=1.12
cc_4 VNB N_A_75_227#_c_193_n 0.00307726f $X=-0.19 $Y=-0.245 $X2=1.425 $Y2=0.34
cc_5 VNB N_A_75_227#_c_194_n 0.00348554f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=1.12
cc_6 VNB N_A_75_227#_c_195_n 0.0344825f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=1.3
cc_7 VNB N_A_75_227#_c_196_n 0.00538013f $X=-0.19 $Y=-0.245 $X2=3.365 $Y2=0.36
cc_8 VNB N_A_75_227#_c_197_n 0.0120995f $X=-0.19 $Y=-0.245 $X2=3.2 $Y2=0.35
cc_9 VNB N_A_75_227#_c_198_n 0.0210495f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=1.135
cc_10 VNB N_A_c_324_n 0.0235524f $X=-0.19 $Y=-0.245 $X2=1.12 $Y2=0.385
cc_11 VNB N_A_M1002_g 0.0285621f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_c_326_n 0.00424938f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_386_23#_M1006_g 0.0336344f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_386_23#_c_369_n 0.076486f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_386_23#_c_370_n 0.0126012f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_386_23#_c_371_n 0.0246414f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.465
cc_17 VNB N_A_386_23#_c_372_n 0.00984973f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.7
cc_18 VNB N_A_386_23#_M1011_g 0.0355421f $X=-0.19 $Y=-0.245 $X2=0.62 $Y2=1.465
cc_19 VNB N_A_386_23#_c_374_n 0.0259245f $X=-0.19 $Y=-0.245 $X2=0.62 $Y2=1.95
cc_20 VNB N_A_386_23#_c_375_n 0.00697882f $X=-0.19 $Y=-0.245 $X2=1.23 $Y2=2.72
cc_21 VNB N_A_386_23#_c_376_n 0.00682553f $X=-0.19 $Y=-0.245 $X2=3.35 $Y2=2.99
cc_22 VNB N_A_386_23#_c_377_n 0.00457202f $X=-0.19 $Y=-0.245 $X2=1.425 $Y2=0.34
cc_23 VNB N_A_386_23#_c_378_n 2.44385e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_386_23#_c_379_n 9.51668e-19 $X=-0.19 $Y=-0.245 $X2=1.23 $Y2=2.035
cc_25 VNB N_B_M1025_g 0.0423531f $X=-0.19 $Y=-0.245 $X2=1.08 $Y2=1.865
cc_26 VNB N_B_c_497_n 0.00197862f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_B_M1004_g 0.0281997f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.79
cc_28 VNB N_B_M1021_g 0.0230134f $X=-0.19 $Y=-0.245 $X2=1.23 $Y2=2.72
cc_29 VNB N_B_c_500_n 0.00360444f $X=-0.19 $Y=-0.245 $X2=3.2 $Y2=0.34
cc_30 VNB N_B_c_501_n 0.00212715f $X=-0.19 $Y=-0.245 $X2=1.23 $Y2=2.035
cc_31 VNB N_B_c_502_n 0.0518963f $X=-0.19 $Y=-0.245 $X2=1.23 $Y2=2.035
cc_32 VNB N_A_1024_300#_M1027_g 0.0461186f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_1024_300#_c_650_n 0.0174851f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_1024_300#_c_651_n 0.00616832f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.7
cc_35 VNB N_A_1024_300#_c_652_n 0.00342923f $X=-0.19 $Y=-0.245 $X2=0.505
+ $Y2=2.365
cc_36 VNB N_A_1024_300#_c_653_n 8.68163e-19 $X=-0.19 $Y=-0.245 $X2=0.705
+ $Y2=1.12
cc_37 VNB N_A_1024_300#_c_654_n 0.00169209f $X=-0.19 $Y=-0.245 $X2=0.705
+ $Y2=2.035
cc_38 VNB N_A_1024_300#_c_655_n 6.55071e-19 $X=-0.19 $Y=-0.245 $X2=1.23 $Y2=2.72
cc_39 VNB N_C_M1012_g 0.0354923f $X=-0.19 $Y=-0.245 $X2=1.08 $Y2=1.865
cc_40 VNB N_C_c_732_n 0.0101334f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_C_c_733_n 0.04531f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_C_c_734_n 0.0171482f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_C_c_735_n 0.0214513f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_C_c_736_n 0.0308399f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.79
cc_45 VNB N_C_c_737_n 0.00271543f $X=-0.19 $Y=-0.245 $X2=0.705 $Y2=2.035
cc_46 VNB N_A_1057_74#_c_806_n 0.0199489f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_1057_74#_c_807_n 0.0157326f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.365
cc_48 VNB N_A_1057_74#_c_808_n 0.0156085f $X=-0.19 $Y=-0.245 $X2=0.62 $Y2=1.95
cc_49 VNB N_A_1057_74#_c_809_n 0.0188693f $X=-0.19 $Y=-0.245 $X2=1.23 $Y2=2.905
cc_50 VNB N_A_1057_74#_c_810_n 0.00252995f $X=-0.19 $Y=-0.245 $X2=1.3 $Y2=0.53
cc_51 VNB N_A_1057_74#_c_811_n 0.0159551f $X=-0.19 $Y=-0.245 $X2=3.35 $Y2=2.99
cc_52 VNB N_A_1057_74#_c_812_n 0.00425762f $X=-0.19 $Y=-0.245 $X2=1.395 $Y2=2.99
cc_53 VNB N_A_1057_74#_c_813_n 0.010379f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_A_1057_74#_c_814_n 0.00552332f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=1.3
cc_55 VNB N_A_1057_74#_c_815_n 0.00330549f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=1.3
cc_56 VNB N_A_1057_74#_c_816_n 0.00511152f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_A_1057_74#_c_817_n 0.00222251f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_A_1057_74#_c_818_n 0.0537622f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_A_1057_74#_c_819_n 0.0815845f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_A_27_373#_c_965_n 0.00716946f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.79
cc_61 VNB N_A_27_373#_c_966_n 0.0244142f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=0.705
cc_62 VNB N_A_27_373#_c_967_n 0.0368156f $X=-0.19 $Y=-0.245 $X2=0.705 $Y2=1.12
cc_63 VNB N_A_27_373#_c_968_n 0.00352767f $X=-0.19 $Y=-0.245 $X2=1.065 $Y2=2.035
cc_64 VNB N_A_27_373#_c_969_n 0.00265022f $X=-0.19 $Y=-0.245 $X2=1.23 $Y2=2.72
cc_65 VNB N_A_27_373#_c_970_n 0.00139242f $X=-0.19 $Y=-0.245 $X2=1.23 $Y2=2.035
cc_66 VNB N_VPWR_c_1077_n 0.422413f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_A_324_373#_c_1184_n 0.00693911f $X=-0.19 $Y=-0.245 $X2=0.505
+ $Y2=1.79
cc_68 VNB N_A_324_373#_c_1185_n 0.00253978f $X=-0.19 $Y=-0.245 $X2=0.505
+ $Y2=2.365
cc_69 VNB N_A_324_373#_c_1186_n 0.00224367f $X=-0.19 $Y=-0.245 $X2=0.545
+ $Y2=1.135
cc_70 VNB N_A_324_373#_c_1187_n 0.00579396f $X=-0.19 $Y=-0.245 $X2=0.545
+ $Y2=0.705
cc_71 VNB N_A_324_373#_c_1188_n 0.00395107f $X=-0.19 $Y=-0.245 $X2=0.62 $Y2=1.95
cc_72 VNB N_A_324_373#_c_1189_n 0.00883735f $X=-0.19 $Y=-0.245 $X2=1.175
+ $Y2=1.12
cc_73 VNB N_A_324_373#_c_1190_n 0.00776468f $X=-0.19 $Y=-0.245 $X2=1.065
+ $Y2=2.035
cc_74 VNB N_A_324_373#_c_1191_n 0.00689628f $X=-0.19 $Y=-0.245 $X2=1.3 $Y2=0.53
cc_75 VNB N_A_321_77#_c_1312_n 0.0080413f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.79
cc_76 VNB N_A_321_77#_c_1313_n 0.0120329f $X=-0.19 $Y=-0.245 $X2=0.705 $Y2=1.12
cc_77 VNB N_A_321_77#_c_1314_n 6.15911e-19 $X=-0.19 $Y=-0.245 $X2=1.3 $Y2=0.425
cc_78 VNB N_A_321_77#_c_1315_n 0.00292969f $X=-0.19 $Y=-0.245 $X2=1.395 $Y2=2.99
cc_79 VNB N_A_321_77#_c_1316_n 2.71919e-19 $X=-0.19 $Y=-0.245 $X2=3.2 $Y2=0.34
cc_80 VNB N_A_321_77#_c_1317_n 0.0234999f $X=-0.19 $Y=-0.245 $X2=1.425 $Y2=0.34
cc_81 VNB N_X_c_1443_n 0.00292847f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=0.705
cc_82 VNB N_X_c_1444_n 0.0010385f $X=-0.19 $Y=-0.245 $X2=0.62 $Y2=1.95
cc_83 VNB X 0.00279061f $X=-0.19 $Y=-0.245 $X2=1.3 $Y2=1.035
cc_84 VNB N_VGND_c_1501_n 0.00734311f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=0.705
cc_85 VNB N_VGND_c_1502_n 0.0123225f $X=-0.19 $Y=-0.245 $X2=0.705 $Y2=1.12
cc_86 VNB N_VGND_c_1503_n 0.0566559f $X=-0.19 $Y=-0.245 $X2=0.705 $Y2=2.035
cc_87 VNB N_VGND_c_1504_n 0.0198695f $X=-0.19 $Y=-0.245 $X2=1.3 $Y2=1.035
cc_88 VNB N_VGND_c_1505_n 0.043087f $X=-0.19 $Y=-0.245 $X2=1.3 $Y2=0.53
cc_89 VNB N_VGND_c_1506_n 0.0181352f $X=-0.19 $Y=-0.245 $X2=1.395 $Y2=2.99
cc_90 VNB N_VGND_c_1507_n 0.010678f $X=-0.19 $Y=-0.245 $X2=1.425 $Y2=0.34
cc_91 VNB N_VGND_c_1508_n 0.0540788f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_92 VNB N_VGND_c_1509_n 0.0779513f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=1.465
cc_93 VNB N_VGND_c_1510_n 0.0197463f $X=-0.19 $Y=-0.245 $X2=3.515 $Y2=2.795
cc_94 VNB N_VGND_c_1511_n 0.0264817f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=1.465
cc_95 VNB N_VGND_c_1512_n 0.00631318f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_96 VNB N_VGND_c_1513_n 0.00326991f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_97 VNB N_VGND_c_1514_n 0.537672f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_98 VPB N_A_75_227#_c_190_n 0.00219432f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.7
cc_99 VPB N_A_75_227#_c_200_n 0.0238838f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.79
cc_100 VPB N_A_75_227#_c_191_n 0.00163357f $X=-0.19 $Y=1.66 $X2=0.62 $Y2=1.95
cc_101 VPB N_A_75_227#_c_202_n 0.00186702f $X=-0.19 $Y=1.66 $X2=1.23 $Y2=2.72
cc_102 VPB N_A_75_227#_c_203_n 0.0337106f $X=-0.19 $Y=1.66 $X2=3.35 $Y2=2.99
cc_103 VPB N_A_75_227#_c_204_n 0.00324785f $X=-0.19 $Y=1.66 $X2=1.395 $Y2=2.99
cc_104 VPB N_A_75_227#_c_205_n 0.00854849f $X=-0.19 $Y=1.66 $X2=3.515 $Y2=2.795
cc_105 VPB N_A_c_324_n 0.0284084f $X=-0.19 $Y=1.66 $X2=1.12 $Y2=0.385
cc_106 VPB N_A_c_326_n 0.00248131f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_107 VPB N_A_386_23#_c_372_n 0.00208407f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.7
cc_108 VPB N_A_386_23#_c_381_n 0.0198381f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.79
cc_109 VPB N_A_386_23#_c_374_n 0.0287255f $X=-0.19 $Y=1.66 $X2=0.62 $Y2=1.95
cc_110 VPB N_A_386_23#_c_375_n 0.00410146f $X=-0.19 $Y=1.66 $X2=1.23 $Y2=2.72
cc_111 VPB N_A_386_23#_c_384_n 0.00171425f $X=-0.19 $Y=1.66 $X2=3.2 $Y2=0.34
cc_112 VPB N_A_386_23#_c_385_n 7.04287e-19 $X=-0.19 $Y=1.66 $X2=0.54 $Y2=1.3
cc_113 VPB N_A_386_23#_c_386_n 0.00142402f $X=-0.19 $Y=1.66 $X2=0.58 $Y2=1.465
cc_114 VPB N_B_c_503_n 0.00917022f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_115 VPB N_B_c_504_n 0.0148751f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_116 VPB N_B_c_497_n 0.00876872f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_117 VPB N_B_M1007_g 0.0101419f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_118 VPB N_B_c_507_n 0.0652391f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_119 VPB N_B_c_508_n 0.0140946f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_120 VPB N_B_c_509_n 0.00645762f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.365
cc_121 VPB N_B_c_510_n 0.0330065f $X=-0.19 $Y=1.66 $X2=0.545 $Y2=1.135
cc_122 VPB N_B_M1020_g 0.00809147f $X=-0.19 $Y=1.66 $X2=0.62 $Y2=1.95
cc_123 VPB N_B_c_512_n 0.0774316f $X=-0.19 $Y=1.66 $X2=1.175 $Y2=1.12
cc_124 VPB N_B_c_513_n 0.0790893f $X=-0.19 $Y=1.66 $X2=0.705 $Y2=2.035
cc_125 VPB N_B_c_514_n 0.0182219f $X=-0.19 $Y=1.66 $X2=1.3 $Y2=0.425
cc_126 VPB N_B_c_500_n 0.0108706f $X=-0.19 $Y=1.66 $X2=3.2 $Y2=0.34
cc_127 VPB N_B_c_516_n 0.00898834f $X=-0.19 $Y=1.66 $X2=0.58 $Y2=1.12
cc_128 VPB N_B_c_501_n 0.00296974f $X=-0.19 $Y=1.66 $X2=1.23 $Y2=2.035
cc_129 VPB N_B_c_502_n 0.0187088f $X=-0.19 $Y=1.66 $X2=1.23 $Y2=2.035
cc_130 VPB N_A_1024_300#_c_650_n 0.0425638f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_131 VPB N_A_1024_300#_c_651_n 0.0138344f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.7
cc_132 VPB N_A_1024_300#_c_658_n 0.00779343f $X=-0.19 $Y=1.66 $X2=0.545
+ $Y2=0.705
cc_133 VPB N_A_1024_300#_c_653_n 0.00172452f $X=-0.19 $Y=1.66 $X2=0.705 $Y2=1.12
cc_134 VPB N_A_1024_300#_c_655_n 0.00270666f $X=-0.19 $Y=1.66 $X2=1.23 $Y2=2.72
cc_135 VPB N_A_1024_300#_c_661_n 0.0147801f $X=-0.19 $Y=1.66 $X2=1.3 $Y2=0.53
cc_136 VPB N_C_c_732_n 0.0110455f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_137 VPB N_C_c_739_n 0.0266295f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_138 VPB N_C_c_736_n 0.0334285f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.79
cc_139 VPB N_C_c_737_n 0.00326488f $X=-0.19 $Y=1.66 $X2=0.705 $Y2=2.035
cc_140 VPB N_A_1057_74#_c_820_n 0.0170451f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_141 VPB N_A_1057_74#_c_821_n 0.0152778f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.465
cc_142 VPB N_A_1057_74#_c_822_n 0.0152843f $X=-0.19 $Y=1.66 $X2=0.545 $Y2=0.705
cc_143 VPB N_A_1057_74#_c_823_n 0.0174296f $X=-0.19 $Y=1.66 $X2=1.065 $Y2=2.035
cc_144 VPB N_A_1057_74#_c_824_n 0.0377701f $X=-0.19 $Y=1.66 $X2=3.2 $Y2=0.34
cc_145 VPB N_A_1057_74#_c_825_n 0.0180278f $X=-0.19 $Y=1.66 $X2=3.365 $Y2=0.36
cc_146 VPB N_A_1057_74#_c_826_n 0.00377141f $X=-0.19 $Y=1.66 $X2=3.515 $Y2=2.795
cc_147 VPB N_A_1057_74#_c_827_n 0.00954227f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_148 VPB N_A_1057_74#_c_818_n 0.0234566f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_149 VPB N_A_1057_74#_c_819_n 0.0551131f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_150 VPB N_A_27_373#_c_971_n 0.00863818f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.365
cc_151 VPB N_A_27_373#_c_972_n 0.00105534f $X=-0.19 $Y=1.66 $X2=0.545 $Y2=1.135
cc_152 VPB N_A_27_373#_c_973_n 0.00886453f $X=-0.19 $Y=1.66 $X2=1.175 $Y2=1.12
cc_153 VPB N_A_27_373#_c_967_n 0.00903323f $X=-0.19 $Y=1.66 $X2=0.705 $Y2=1.12
cc_154 VPB N_A_27_373#_c_975_n 0.002215f $X=-0.19 $Y=1.66 $X2=1.26 $Y2=0.53
cc_155 VPB N_A_27_373#_c_970_n 0.00139459f $X=-0.19 $Y=1.66 $X2=1.23 $Y2=2.035
cc_156 VPB N_A_27_373#_c_977_n 0.0375515f $X=-0.19 $Y=1.66 $X2=3.2 $Y2=0.35
cc_157 VPB N_VPWR_c_1078_n 0.0111985f $X=-0.19 $Y=1.66 $X2=0.545 $Y2=1.135
cc_158 VPB N_VPWR_c_1079_n 0.0137669f $X=-0.19 $Y=1.66 $X2=0.62 $Y2=1.95
cc_159 VPB N_VPWR_c_1080_n 0.013306f $X=-0.19 $Y=1.66 $X2=1.065 $Y2=2.035
cc_160 VPB N_VPWR_c_1081_n 0.0024682f $X=-0.19 $Y=1.66 $X2=1.23 $Y2=2.905
cc_161 VPB N_VPWR_c_1082_n 0.0194151f $X=-0.19 $Y=1.66 $X2=1.23 $Y2=2.72
cc_162 VPB N_VPWR_c_1083_n 0.00935081f $X=-0.19 $Y=1.66 $X2=1.26 $Y2=0.53
cc_163 VPB N_VPWR_c_1084_n 0.0108116f $X=-0.19 $Y=1.66 $X2=1.425 $Y2=0.34
cc_164 VPB N_VPWR_c_1085_n 0.0585173f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_165 VPB N_VPWR_c_1086_n 0.0183206f $X=-0.19 $Y=1.66 $X2=3.2 $Y2=0.35
cc_166 VPB N_VPWR_c_1087_n 0.0861107f $X=-0.19 $Y=1.66 $X2=3.515 $Y2=2.99
cc_167 VPB N_VPWR_c_1088_n 0.0707383f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_168 VPB N_VPWR_c_1089_n 0.0204088f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_169 VPB N_VPWR_c_1090_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_170 VPB N_VPWR_c_1091_n 0.00614151f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_171 VPB N_VPWR_c_1092_n 0.0119958f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_172 VPB N_VPWR_c_1093_n 0.00324402f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_173 VPB N_VPWR_c_1077_n 0.110645f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_174 VPB N_A_324_373#_c_1192_n 0.00150474f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.7
cc_175 VPB N_A_324_373#_c_1184_n 0.00266963f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.79
cc_176 VPB N_A_324_373#_c_1187_n 0.00645585f $X=-0.19 $Y=1.66 $X2=0.545
+ $Y2=0.705
cc_177 VPB N_A_324_373#_c_1195_n 0.00346709f $X=-0.19 $Y=1.66 $X2=3.35 $Y2=2.99
cc_178 VPB N_A_324_373#_c_1196_n 0.0028297f $X=-0.19 $Y=1.66 $X2=0.54 $Y2=1.3
cc_179 VPB N_A_324_373#_c_1197_n 0.00757294f $X=-0.19 $Y=1.66 $X2=0.54 $Y2=1.3
cc_180 VPB N_A_321_77#_c_1318_n 0.00340067f $X=-0.19 $Y=1.66 $X2=0.62 $Y2=1.465
cc_181 VPB N_A_321_77#_c_1313_n 0.00361327f $X=-0.19 $Y=1.66 $X2=0.705 $Y2=1.12
cc_182 VPB N_A_321_77#_c_1320_n 0.00837164f $X=-0.19 $Y=1.66 $X2=1.065 $Y2=2.035
cc_183 VPB N_A_321_77#_c_1321_n 0.00209491f $X=-0.19 $Y=1.66 $X2=1.23 $Y2=2.72
cc_184 VPB N_X_c_1446_n 0.00257348f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.79
cc_185 VPB N_X_c_1447_n 0.00105539f $X=-0.19 $Y=1.66 $X2=1.23 $Y2=2.905
cc_186 VPB N_X_c_1448_n 0.00161844f $X=-0.19 $Y=1.66 $X2=1.23 $Y2=2.72
cc_187 VPB X 0.00257348f $X=-0.19 $Y=1.66 $X2=0.54 $Y2=1.465
cc_188 N_A_75_227#_c_190_n N_A_c_324_n 0.0115699f $X=0.505 $Y=1.7 $X2=-0.19
+ $Y2=-0.245
cc_189 N_A_75_227#_c_200_n N_A_c_324_n 0.0252355f $X=0.505 $Y=1.79 $X2=-0.19
+ $Y2=-0.245
cc_190 N_A_75_227#_c_191_n N_A_c_324_n 0.0054287f $X=0.62 $Y=1.95 $X2=-0.19
+ $Y2=-0.245
cc_191 N_A_75_227#_c_192_n N_A_c_324_n 0.00131609f $X=1.175 $Y=1.12 $X2=-0.19
+ $Y2=-0.245
cc_192 N_A_75_227#_c_210_p N_A_c_324_n 0.0122144f $X=1.065 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_193 N_A_75_227#_c_211_p N_A_c_324_n 0.00129198f $X=1.23 $Y=2.12 $X2=-0.19
+ $Y2=-0.245
cc_194 N_A_75_227#_c_202_n N_A_c_324_n 0.00947394f $X=1.23 $Y=2.72 $X2=-0.19
+ $Y2=-0.245
cc_195 N_A_75_227#_c_204_n N_A_c_324_n 0.00242403f $X=1.395 $Y=2.99 $X2=-0.19
+ $Y2=-0.245
cc_196 N_A_75_227#_c_194_n N_A_c_324_n 3.13863e-19 $X=0.58 $Y=1.12 $X2=-0.19
+ $Y2=-0.245
cc_197 N_A_75_227#_c_195_n N_A_c_324_n 0.00548466f $X=0.54 $Y=1.3 $X2=-0.19
+ $Y2=-0.245
cc_198 N_A_75_227#_c_192_n N_A_M1002_g 0.0141792f $X=1.175 $Y=1.12 $X2=0 $Y2=0
cc_199 N_A_75_227#_c_217_p N_A_M1002_g 2.2106e-19 $X=1.26 $Y=0.53 $X2=0 $Y2=0
cc_200 N_A_75_227#_c_193_n N_A_M1002_g 0.00116563f $X=1.425 $Y=0.34 $X2=0 $Y2=0
cc_201 N_A_75_227#_c_194_n N_A_M1002_g 0.00121602f $X=0.58 $Y=1.12 $X2=0 $Y2=0
cc_202 N_A_75_227#_c_195_n N_A_M1002_g 0.0119439f $X=0.54 $Y=1.3 $X2=0 $Y2=0
cc_203 N_A_75_227#_c_198_n N_A_M1002_g 0.0203508f $X=0.54 $Y=1.135 $X2=0 $Y2=0
cc_204 N_A_75_227#_c_190_n N_A_c_326_n 3.40563e-19 $X=0.505 $Y=1.7 $X2=0 $Y2=0
cc_205 N_A_75_227#_c_192_n N_A_c_326_n 0.031511f $X=1.175 $Y=1.12 $X2=0 $Y2=0
cc_206 N_A_75_227#_c_210_p N_A_c_326_n 0.00930675f $X=1.065 $Y=2.035 $X2=0 $Y2=0
cc_207 N_A_75_227#_c_211_p N_A_c_326_n 0.0173128f $X=1.23 $Y=2.12 $X2=0 $Y2=0
cc_208 N_A_75_227#_c_194_n N_A_c_326_n 0.0261391f $X=0.58 $Y=1.12 $X2=0 $Y2=0
cc_209 N_A_75_227#_c_195_n N_A_c_326_n 3.13185e-19 $X=0.54 $Y=1.3 $X2=0 $Y2=0
cc_210 N_A_75_227#_c_197_n N_A_386_23#_M1006_g 0.00804191f $X=3.2 $Y=0.35 $X2=0
+ $Y2=0
cc_211 N_A_75_227#_c_197_n N_A_386_23#_c_369_n 0.0211522f $X=3.2 $Y=0.35 $X2=0
+ $Y2=0
cc_212 N_A_75_227#_c_197_n N_A_386_23#_c_370_n 0.00150581f $X=3.2 $Y=0.35 $X2=0
+ $Y2=0
cc_213 N_A_75_227#_c_203_n N_A_386_23#_c_381_n 4.13058e-19 $X=3.35 $Y=2.99 $X2=0
+ $Y2=0
cc_214 N_A_75_227#_c_196_n N_A_386_23#_M1011_g 8.00488e-19 $X=3.365 $Y=0.36
+ $X2=0 $Y2=0
cc_215 N_A_75_227#_c_197_n N_A_386_23#_M1011_g 0.0115799f $X=3.2 $Y=0.35 $X2=0
+ $Y2=0
cc_216 N_A_75_227#_c_203_n N_A_386_23#_c_374_n 0.00155596f $X=3.35 $Y=2.99 $X2=0
+ $Y2=0
cc_217 N_A_75_227#_c_205_n N_A_386_23#_c_374_n 0.00326052f $X=3.515 $Y=2.795
+ $X2=0 $Y2=0
cc_218 N_A_75_227#_M1009_d N_A_386_23#_c_384_n 0.00112948f $X=3.28 $Y=1.865
+ $X2=0 $Y2=0
cc_219 N_A_75_227#_M1009_d N_A_386_23#_c_385_n 0.00367614f $X=3.28 $Y=1.865
+ $X2=0 $Y2=0
cc_220 N_A_75_227#_c_192_n N_B_M1025_g 0.00470939f $X=1.175 $Y=1.12 $X2=0 $Y2=0
cc_221 N_A_75_227#_c_217_p N_B_M1025_g 2.28462e-19 $X=1.26 $Y=0.53 $X2=0 $Y2=0
cc_222 N_A_75_227#_c_197_n N_B_M1025_g 0.013294f $X=3.2 $Y=0.35 $X2=0 $Y2=0
cc_223 N_A_75_227#_c_202_n N_B_c_503_n 0.00351671f $X=1.23 $Y=2.72 $X2=0 $Y2=0
cc_224 N_A_75_227#_c_203_n N_B_c_504_n 0.0171103f $X=3.35 $Y=2.99 $X2=0 $Y2=0
cc_225 N_A_75_227#_c_211_p N_B_M1007_g 0.00128638f $X=1.23 $Y=2.12 $X2=0 $Y2=0
cc_226 N_A_75_227#_c_202_n N_B_M1007_g 0.00645319f $X=1.23 $Y=2.72 $X2=0 $Y2=0
cc_227 N_A_75_227#_c_203_n N_B_c_507_n 0.0165357f $X=3.35 $Y=2.99 $X2=0 $Y2=0
cc_228 N_A_75_227#_c_197_n N_B_M1004_g 0.00112634f $X=3.2 $Y=0.35 $X2=0 $Y2=0
cc_229 N_A_75_227#_c_203_n N_B_c_510_n 0.0165978f $X=3.35 $Y=2.99 $X2=0 $Y2=0
cc_230 N_A_75_227#_c_205_n N_B_c_510_n 0.00238787f $X=3.515 $Y=2.795 $X2=0 $Y2=0
cc_231 N_A_75_227#_c_203_n N_B_c_512_n 0.00871983f $X=3.35 $Y=2.99 $X2=0 $Y2=0
cc_232 N_A_75_227#_c_205_n N_B_c_512_n 0.00899965f $X=3.515 $Y=2.795 $X2=0 $Y2=0
cc_233 N_A_75_227#_c_205_n N_B_c_513_n 0.0137302f $X=3.515 $Y=2.795 $X2=0 $Y2=0
cc_234 N_A_75_227#_c_196_n N_B_M1021_g 0.00356999f $X=3.365 $Y=0.36 $X2=0 $Y2=0
cc_235 N_A_75_227#_c_203_n N_A_27_373#_c_971_n 0.038228f $X=3.35 $Y=2.99 $X2=0
+ $Y2=0
cc_236 N_A_75_227#_c_202_n N_A_27_373#_c_972_n 0.0140536f $X=1.23 $Y=2.72 $X2=0
+ $Y2=0
cc_237 N_A_75_227#_c_203_n N_A_27_373#_c_972_n 0.0152397f $X=3.35 $Y=2.99 $X2=0
+ $Y2=0
cc_238 N_A_75_227#_c_194_n N_A_27_373#_c_966_n 0.00252896f $X=0.58 $Y=1.12 $X2=0
+ $Y2=0
cc_239 N_A_75_227#_c_195_n N_A_27_373#_c_966_n 0.0023718f $X=0.54 $Y=1.3 $X2=0
+ $Y2=0
cc_240 N_A_75_227#_c_198_n N_A_27_373#_c_966_n 0.00804959f $X=0.54 $Y=1.135
+ $X2=0 $Y2=0
cc_241 N_A_75_227#_c_200_n N_A_27_373#_c_973_n 0.00715343f $X=0.505 $Y=1.79
+ $X2=0 $Y2=0
cc_242 N_A_75_227#_c_191_n N_A_27_373#_c_973_n 0.00733813f $X=0.62 $Y=1.95 $X2=0
+ $Y2=0
cc_243 N_A_75_227#_c_261_p N_A_27_373#_c_973_n 0.0115538f $X=0.705 $Y=2.035
+ $X2=0 $Y2=0
cc_244 N_A_75_227#_c_190_n N_A_27_373#_c_967_n 0.00708041f $X=0.505 $Y=1.7 $X2=0
+ $Y2=0
cc_245 N_A_75_227#_c_200_n N_A_27_373#_c_967_n 0.0011211f $X=0.505 $Y=1.79 $X2=0
+ $Y2=0
cc_246 N_A_75_227#_c_191_n N_A_27_373#_c_967_n 0.0205539f $X=0.62 $Y=1.95 $X2=0
+ $Y2=0
cc_247 N_A_75_227#_c_194_n N_A_27_373#_c_967_n 0.0324438f $X=0.58 $Y=1.12 $X2=0
+ $Y2=0
cc_248 N_A_75_227#_c_195_n N_A_27_373#_c_967_n 0.00816612f $X=0.54 $Y=1.3 $X2=0
+ $Y2=0
cc_249 N_A_75_227#_c_198_n N_A_27_373#_c_967_n 0.00650851f $X=0.54 $Y=1.135
+ $X2=0 $Y2=0
cc_250 N_A_75_227#_c_192_n N_A_27_373#_c_968_n 0.00352449f $X=1.175 $Y=1.12
+ $X2=0 $Y2=0
cc_251 N_A_75_227#_c_203_n N_A_27_373#_c_975_n 0.031064f $X=3.35 $Y=2.99 $X2=0
+ $Y2=0
cc_252 N_A_75_227#_c_205_n N_A_27_373#_c_975_n 7.42852e-19 $X=3.515 $Y=2.795
+ $X2=0 $Y2=0
cc_253 N_A_75_227#_M1023_d N_A_27_373#_c_996_n 0.0053736f $X=1.08 $Y=1.865 $X2=0
+ $Y2=0
cc_254 N_A_75_227#_c_200_n N_A_27_373#_c_996_n 0.00674706f $X=0.505 $Y=1.79
+ $X2=0 $Y2=0
cc_255 N_A_75_227#_c_210_p N_A_27_373#_c_996_n 0.0252266f $X=1.065 $Y=2.035
+ $X2=0 $Y2=0
cc_256 N_A_75_227#_c_261_p N_A_27_373#_c_996_n 0.0127006f $X=0.705 $Y=2.035
+ $X2=0 $Y2=0
cc_257 N_A_75_227#_c_211_p N_A_27_373#_c_996_n 0.0302905f $X=1.23 $Y=2.12 $X2=0
+ $Y2=0
cc_258 N_A_75_227#_c_194_n N_A_27_373#_c_996_n 0.00231569f $X=0.58 $Y=1.12 $X2=0
+ $Y2=0
cc_259 N_A_75_227#_c_195_n N_A_27_373#_c_996_n 5.88073e-19 $X=0.54 $Y=1.3 $X2=0
+ $Y2=0
cc_260 N_A_75_227#_c_191_n N_A_27_373#_c_1003_n 8.60777e-19 $X=0.62 $Y=1.95
+ $X2=0 $Y2=0
cc_261 N_A_75_227#_c_261_p N_A_27_373#_c_1003_n 8.91026e-19 $X=0.705 $Y=2.035
+ $X2=0 $Y2=0
cc_262 N_A_75_227#_c_195_n N_A_27_373#_c_1003_n 2.18873e-19 $X=0.54 $Y=1.3 $X2=0
+ $Y2=0
cc_263 N_A_75_227#_c_211_p N_A_27_373#_c_1006_n 8.00194e-19 $X=1.23 $Y=2.12
+ $X2=0 $Y2=0
cc_264 N_A_75_227#_c_202_n N_A_27_373#_c_1006_n 7.80159e-19 $X=1.23 $Y=2.72
+ $X2=0 $Y2=0
cc_265 N_A_75_227#_c_211_p N_A_27_373#_c_970_n 0.0116148f $X=1.23 $Y=2.12 $X2=0
+ $Y2=0
cc_266 N_A_75_227#_c_202_n N_A_27_373#_c_970_n 0.0329334f $X=1.23 $Y=2.72 $X2=0
+ $Y2=0
cc_267 N_A_75_227#_c_191_n N_VPWR_M1026_d 0.00101413f $X=0.62 $Y=1.95 $X2=-0.19
+ $Y2=-0.245
cc_268 N_A_75_227#_c_210_p N_VPWR_M1026_d 0.00814722f $X=1.065 $Y=2.035
+ $X2=-0.19 $Y2=-0.245
cc_269 N_A_75_227#_c_261_p N_VPWR_M1026_d 7.41438e-19 $X=0.705 $Y=2.035
+ $X2=-0.19 $Y2=-0.245
cc_270 N_A_75_227#_c_200_n N_VPWR_c_1078_n 0.013136f $X=0.505 $Y=1.79 $X2=0
+ $Y2=0
cc_271 N_A_75_227#_c_210_p N_VPWR_c_1078_n 0.0122582f $X=1.065 $Y=2.035 $X2=0
+ $Y2=0
cc_272 N_A_75_227#_c_261_p N_VPWR_c_1078_n 0.00657661f $X=0.705 $Y=2.035 $X2=0
+ $Y2=0
cc_273 N_A_75_227#_c_202_n N_VPWR_c_1078_n 0.0246613f $X=1.23 $Y=2.72 $X2=0
+ $Y2=0
cc_274 N_A_75_227#_c_204_n N_VPWR_c_1078_n 0.0146282f $X=1.395 $Y=2.99 $X2=0
+ $Y2=0
cc_275 N_A_75_227#_c_200_n N_VPWR_c_1086_n 0.00458208f $X=0.505 $Y=1.79 $X2=0
+ $Y2=0
cc_276 N_A_75_227#_c_203_n N_VPWR_c_1087_n 0.124833f $X=3.35 $Y=2.99 $X2=0 $Y2=0
cc_277 N_A_75_227#_c_204_n N_VPWR_c_1087_n 0.0236566f $X=1.395 $Y=2.99 $X2=0
+ $Y2=0
cc_278 N_A_75_227#_c_205_n N_VPWR_c_1087_n 0.0213919f $X=3.515 $Y=2.795 $X2=0
+ $Y2=0
cc_279 N_A_75_227#_c_200_n N_VPWR_c_1077_n 0.00467808f $X=0.505 $Y=1.79 $X2=0
+ $Y2=0
cc_280 N_A_75_227#_c_203_n N_VPWR_c_1077_n 0.0656561f $X=3.35 $Y=2.99 $X2=0
+ $Y2=0
cc_281 N_A_75_227#_c_204_n N_VPWR_c_1077_n 0.0128296f $X=1.395 $Y=2.99 $X2=0
+ $Y2=0
cc_282 N_A_75_227#_c_205_n N_VPWR_c_1077_n 0.0110564f $X=3.515 $Y=2.795 $X2=0
+ $Y2=0
cc_283 N_A_75_227#_M1009_d N_A_324_373#_c_1195_n 0.00581751f $X=3.28 $Y=1.865
+ $X2=0 $Y2=0
cc_284 N_A_75_227#_c_197_n N_A_321_77#_M1025_d 0.00205163f $X=3.2 $Y=0.35
+ $X2=-0.19 $Y2=-0.245
cc_285 N_A_75_227#_M1011_d N_A_321_77#_c_1312_n 0.0106006f $X=3.145 $Y=0.605
+ $X2=0 $Y2=0
cc_286 N_A_75_227#_c_196_n N_A_321_77#_c_1312_n 0.0228577f $X=3.365 $Y=0.36
+ $X2=0 $Y2=0
cc_287 N_A_75_227#_c_197_n N_A_321_77#_c_1312_n 0.0252875f $X=3.2 $Y=0.35 $X2=0
+ $Y2=0
cc_288 N_A_75_227#_M1009_d N_A_321_77#_c_1318_n 0.00927554f $X=3.28 $Y=1.865
+ $X2=0 $Y2=0
cc_289 N_A_75_227#_c_203_n N_A_321_77#_c_1318_n 0.00653625f $X=3.35 $Y=2.99
+ $X2=0 $Y2=0
cc_290 N_A_75_227#_c_205_n N_A_321_77#_c_1318_n 0.0241281f $X=3.515 $Y=2.795
+ $X2=0 $Y2=0
cc_291 N_A_75_227#_c_203_n N_A_321_77#_c_1329_n 0.00921841f $X=3.35 $Y=2.99
+ $X2=0 $Y2=0
cc_292 N_A_75_227#_c_197_n N_A_321_77#_c_1314_n 0.0214403f $X=3.2 $Y=0.35 $X2=0
+ $Y2=0
cc_293 N_A_75_227#_c_197_n N_A_321_77#_c_1315_n 0.0532333f $X=3.2 $Y=0.35 $X2=0
+ $Y2=0
cc_294 N_A_75_227#_c_192_n N_VGND_c_1501_n 0.0211827f $X=1.175 $Y=1.12 $X2=0
+ $Y2=0
cc_295 N_A_75_227#_c_193_n N_VGND_c_1501_n 0.0118948f $X=1.425 $Y=0.34 $X2=0
+ $Y2=0
cc_296 N_A_75_227#_c_194_n N_VGND_c_1501_n 0.00299742f $X=0.58 $Y=1.12 $X2=0
+ $Y2=0
cc_297 N_A_75_227#_c_195_n N_VGND_c_1501_n 2.06276e-19 $X=0.54 $Y=1.3 $X2=0
+ $Y2=0
cc_298 N_A_75_227#_c_198_n N_VGND_c_1501_n 0.00578941f $X=0.54 $Y=1.135 $X2=0
+ $Y2=0
cc_299 N_A_75_227#_c_193_n N_VGND_c_1509_n 0.0179217f $X=1.425 $Y=0.34 $X2=0
+ $Y2=0
cc_300 N_A_75_227#_c_197_n N_VGND_c_1509_n 0.131374f $X=3.2 $Y=0.35 $X2=0 $Y2=0
cc_301 N_A_75_227#_c_198_n N_VGND_c_1511_n 0.00540915f $X=0.54 $Y=1.135 $X2=0
+ $Y2=0
cc_302 N_A_75_227#_M1011_d N_VGND_c_1514_n 0.00251887f $X=3.145 $Y=0.605 $X2=0
+ $Y2=0
cc_303 N_A_75_227#_c_193_n N_VGND_c_1514_n 0.00971942f $X=1.425 $Y=0.34 $X2=0
+ $Y2=0
cc_304 N_A_75_227#_c_197_n N_VGND_c_1514_n 0.0734849f $X=3.2 $Y=0.35 $X2=0 $Y2=0
cc_305 N_A_75_227#_c_198_n N_VGND_c_1514_n 0.0054106f $X=0.54 $Y=1.135 $X2=0
+ $Y2=0
cc_306 N_A_c_324_n N_B_M1025_g 0.0194584f $X=1.005 $Y=1.79 $X2=0 $Y2=0
cc_307 N_A_M1002_g N_B_M1025_g 0.0160975f $X=1.045 $Y=0.705 $X2=0 $Y2=0
cc_308 N_A_c_326_n N_B_M1025_g 0.00288099f $X=1.08 $Y=1.54 $X2=0 $Y2=0
cc_309 N_A_c_324_n N_B_c_503_n 0.0047983f $X=1.005 $Y=1.79 $X2=0 $Y2=0
cc_310 N_A_c_324_n N_B_c_497_n 0.00252664f $X=1.005 $Y=1.79 $X2=0 $Y2=0
cc_311 N_A_c_324_n N_B_M1007_g 0.0137835f $X=1.005 $Y=1.79 $X2=0 $Y2=0
cc_312 N_A_M1002_g N_A_27_373#_c_968_n 8.13749e-19 $X=1.045 $Y=0.705 $X2=0 $Y2=0
cc_313 N_A_c_326_n N_A_27_373#_c_968_n 0.00584677f $X=1.08 $Y=1.54 $X2=0 $Y2=0
cc_314 N_A_c_326_n N_A_27_373#_c_996_n 0.00309875f $X=1.08 $Y=1.54 $X2=0 $Y2=0
cc_315 N_A_c_324_n N_A_27_373#_c_970_n 9.79361e-19 $X=1.005 $Y=1.79 $X2=0 $Y2=0
cc_316 N_A_c_326_n N_A_27_373#_c_970_n 0.017717f $X=1.08 $Y=1.54 $X2=0 $Y2=0
cc_317 N_A_c_324_n N_VPWR_c_1078_n 0.00418559f $X=1.005 $Y=1.79 $X2=0 $Y2=0
cc_318 N_A_c_324_n N_VPWR_c_1087_n 0.00467123f $X=1.005 $Y=1.79 $X2=0 $Y2=0
cc_319 N_A_c_324_n N_VPWR_c_1077_n 0.00464368f $X=1.005 $Y=1.79 $X2=0 $Y2=0
cc_320 N_A_M1002_g N_VGND_c_1501_n 0.00984806f $X=1.045 $Y=0.705 $X2=0 $Y2=0
cc_321 N_A_M1002_g N_VGND_c_1509_n 0.00471276f $X=1.045 $Y=0.705 $X2=0 $Y2=0
cc_322 N_A_M1002_g N_VGND_c_1514_n 0.0045449f $X=1.045 $Y=0.705 $X2=0 $Y2=0
cc_323 N_A_386_23#_c_370_n N_B_M1025_g 0.0305639f $X=2.08 $Y=0.19 $X2=0 $Y2=0
cc_324 N_A_386_23#_c_372_n N_B_M1025_g 0.00272004f $X=2.245 $Y=1.7 $X2=0 $Y2=0
cc_325 N_A_386_23#_c_372_n N_B_c_497_n 0.00268134f $X=2.245 $Y=1.7 $X2=0 $Y2=0
cc_326 N_A_386_23#_c_381_n N_B_M1007_g 0.0108552f $X=2.245 $Y=1.79 $X2=0 $Y2=0
cc_327 N_A_386_23#_c_381_n N_B_c_507_n 0.00313886f $X=2.245 $Y=1.79 $X2=0 $Y2=0
cc_328 N_A_386_23#_M1006_g N_B_M1004_g 0.017105f $X=2.005 $Y=0.815 $X2=0 $Y2=0
cc_329 N_A_386_23#_c_369_n N_B_M1004_g 0.00976806f $X=2.995 $Y=0.19 $X2=0 $Y2=0
cc_330 N_A_386_23#_c_371_n N_B_M1004_g 0.014943f $X=2.245 $Y=1.47 $X2=0 $Y2=0
cc_331 N_A_386_23#_M1011_g N_B_M1004_g 0.0325534f $X=3.07 $Y=0.925 $X2=0 $Y2=0
cc_332 N_A_386_23#_c_375_n N_B_M1004_g 3.10708e-19 $X=3.6 $Y=1.54 $X2=0 $Y2=0
cc_333 N_A_386_23#_c_381_n N_B_c_509_n 0.00242326f $X=2.245 $Y=1.79 $X2=0 $Y2=0
cc_334 N_A_386_23#_c_374_n N_B_c_509_n 0.00938363f $X=3.205 $Y=1.79 $X2=0 $Y2=0
cc_335 N_A_386_23#_c_381_n N_B_M1020_g 0.0198117f $X=2.245 $Y=1.79 $X2=0 $Y2=0
cc_336 N_A_386_23#_c_374_n N_B_M1020_g 0.0131325f $X=3.205 $Y=1.79 $X2=0 $Y2=0
cc_337 N_A_386_23#_c_374_n N_B_c_512_n 0.00737859f $X=3.205 $Y=1.79 $X2=0 $Y2=0
cc_338 N_A_386_23#_c_374_n N_B_c_513_n 0.0273147f $X=3.205 $Y=1.79 $X2=0 $Y2=0
cc_339 N_A_386_23#_c_384_n N_B_c_513_n 0.00685915f $X=3.685 $Y=1.95 $X2=0 $Y2=0
cc_340 N_A_386_23#_c_385_n N_B_c_513_n 0.00395133f $X=3.77 $Y=2.075 $X2=0 $Y2=0
cc_341 N_A_386_23#_c_386_n N_B_c_513_n 0.0128367f $X=4.105 $Y=2.115 $X2=0 $Y2=0
cc_342 N_A_386_23#_c_379_n N_B_c_513_n 6.38429e-19 $X=3.685 $Y=1.54 $X2=0 $Y2=0
cc_343 N_A_386_23#_c_376_n N_B_M1021_g 0.00370096f $X=3.685 $Y=1.375 $X2=0 $Y2=0
cc_344 N_A_386_23#_c_378_n N_B_M1021_g 0.00328266f $X=3.925 $Y=1.04 $X2=0 $Y2=0
cc_345 N_A_386_23#_c_384_n N_B_c_514_n 4.82877e-19 $X=3.685 $Y=1.95 $X2=0 $Y2=0
cc_346 N_A_386_23#_c_386_n N_B_c_514_n 0.00232542f $X=4.105 $Y=2.115 $X2=0 $Y2=0
cc_347 N_A_386_23#_c_372_n N_B_c_500_n 0.014943f $X=2.245 $Y=1.7 $X2=0 $Y2=0
cc_348 N_A_386_23#_c_374_n N_B_c_500_n 0.00791823f $X=3.205 $Y=1.79 $X2=0 $Y2=0
cc_349 N_A_386_23#_c_375_n N_B_c_500_n 3.16617e-19 $X=3.6 $Y=1.54 $X2=0 $Y2=0
cc_350 N_A_386_23#_c_376_n N_B_c_501_n 0.00184128f $X=3.685 $Y=1.375 $X2=0 $Y2=0
cc_351 N_A_386_23#_c_384_n N_B_c_501_n 0.00562831f $X=3.685 $Y=1.95 $X2=0 $Y2=0
cc_352 N_A_386_23#_c_378_n N_B_c_501_n 0.00730998f $X=3.925 $Y=1.04 $X2=0 $Y2=0
cc_353 N_A_386_23#_c_386_n N_B_c_501_n 0.0220612f $X=4.105 $Y=2.115 $X2=0 $Y2=0
cc_354 N_A_386_23#_c_379_n N_B_c_501_n 0.0271008f $X=3.685 $Y=1.54 $X2=0 $Y2=0
cc_355 N_A_386_23#_c_374_n N_B_c_502_n 0.00670177f $X=3.205 $Y=1.79 $X2=0 $Y2=0
cc_356 N_A_386_23#_c_376_n N_B_c_502_n 6.03443e-19 $X=3.685 $Y=1.375 $X2=0 $Y2=0
cc_357 N_A_386_23#_c_378_n N_B_c_502_n 0.00585644f $X=3.925 $Y=1.04 $X2=0 $Y2=0
cc_358 N_A_386_23#_c_386_n N_B_c_502_n 0.00339088f $X=4.105 $Y=2.115 $X2=0 $Y2=0
cc_359 N_A_386_23#_c_379_n N_B_c_502_n 0.00767005f $X=3.685 $Y=1.54 $X2=0 $Y2=0
cc_360 N_A_386_23#_M1006_g N_A_27_373#_c_965_n 0.00779425f $X=2.005 $Y=0.815
+ $X2=0 $Y2=0
cc_361 N_A_386_23#_c_371_n N_A_27_373#_c_965_n 0.00339009f $X=2.245 $Y=1.47
+ $X2=0 $Y2=0
cc_362 N_A_386_23#_c_381_n N_A_27_373#_c_971_n 0.00649349f $X=2.245 $Y=1.79
+ $X2=0 $Y2=0
cc_363 N_A_386_23#_c_371_n N_A_27_373#_c_968_n 0.00307815f $X=2.245 $Y=1.47
+ $X2=0 $Y2=0
cc_364 N_A_386_23#_M1006_g N_A_27_373#_c_969_n 0.0046962f $X=2.005 $Y=0.815
+ $X2=0 $Y2=0
cc_365 N_A_386_23#_c_371_n N_A_27_373#_c_969_n 0.00729644f $X=2.245 $Y=1.47
+ $X2=0 $Y2=0
cc_366 N_A_386_23#_c_381_n N_A_27_373#_c_975_n 0.00730153f $X=2.245 $Y=1.79
+ $X2=0 $Y2=0
cc_367 N_A_386_23#_c_374_n N_A_27_373#_c_975_n 8.80245e-19 $X=3.205 $Y=1.79
+ $X2=0 $Y2=0
cc_368 N_A_386_23#_c_372_n N_A_27_373#_c_970_n 0.00120455f $X=2.245 $Y=1.7 $X2=0
+ $Y2=0
cc_369 N_A_386_23#_c_381_n N_A_27_373#_c_970_n 0.0049847f $X=2.245 $Y=1.79 $X2=0
+ $Y2=0
cc_370 N_A_386_23#_c_372_n N_A_324_373#_c_1192_n 8.31271e-19 $X=2.245 $Y=1.7
+ $X2=0 $Y2=0
cc_371 N_A_386_23#_c_381_n N_A_324_373#_c_1192_n 0.00829068f $X=2.245 $Y=1.79
+ $X2=0 $Y2=0
cc_372 N_A_386_23#_c_372_n N_A_324_373#_c_1184_n 0.00574458f $X=2.245 $Y=1.7
+ $X2=0 $Y2=0
cc_373 N_A_386_23#_c_374_n N_A_324_373#_c_1184_n 6.38604e-19 $X=3.205 $Y=1.79
+ $X2=0 $Y2=0
cc_374 N_A_386_23#_c_375_n N_A_324_373#_c_1184_n 0.0115248f $X=3.6 $Y=1.54 $X2=0
+ $Y2=0
cc_375 N_A_386_23#_c_371_n N_A_324_373#_c_1185_n 0.00642326f $X=2.245 $Y=1.47
+ $X2=0 $Y2=0
cc_376 N_A_386_23#_c_372_n N_A_324_373#_c_1185_n 0.00506743f $X=2.245 $Y=1.7
+ $X2=0 $Y2=0
cc_377 N_A_386_23#_c_371_n N_A_324_373#_c_1186_n 0.0012074f $X=2.245 $Y=1.47
+ $X2=0 $Y2=0
cc_378 N_A_386_23#_M1011_g N_A_324_373#_c_1186_n 0.00329076f $X=3.07 $Y=0.925
+ $X2=0 $Y2=0
cc_379 N_A_386_23#_c_374_n N_A_324_373#_c_1186_n 4.48181e-19 $X=3.205 $Y=1.79
+ $X2=0 $Y2=0
cc_380 N_A_386_23#_c_375_n N_A_324_373#_c_1186_n 0.00801193f $X=3.6 $Y=1.54
+ $X2=0 $Y2=0
cc_381 N_A_386_23#_M1011_g N_A_324_373#_c_1210_n 0.00577182f $X=3.07 $Y=0.925
+ $X2=0 $Y2=0
cc_382 N_A_386_23#_c_375_n N_A_324_373#_c_1210_n 0.00180109f $X=3.6 $Y=1.54
+ $X2=0 $Y2=0
cc_383 N_A_386_23#_c_376_n N_A_324_373#_c_1210_n 0.00238919f $X=3.685 $Y=1.375
+ $X2=0 $Y2=0
cc_384 N_A_386_23#_c_377_n N_A_324_373#_c_1210_n 0.00562748f $X=3.77 $Y=1.04
+ $X2=0 $Y2=0
cc_385 N_A_386_23#_c_381_n N_A_324_373#_c_1195_n 0.00157986f $X=2.245 $Y=1.79
+ $X2=0 $Y2=0
cc_386 N_A_386_23#_c_374_n N_A_324_373#_c_1195_n 0.00526178f $X=3.205 $Y=1.79
+ $X2=0 $Y2=0
cc_387 N_A_386_23#_c_375_n N_A_324_373#_c_1195_n 0.0136422f $X=3.6 $Y=1.54 $X2=0
+ $Y2=0
cc_388 N_A_386_23#_c_385_n N_A_324_373#_c_1195_n 0.0167115f $X=3.77 $Y=2.075
+ $X2=0 $Y2=0
cc_389 N_A_386_23#_c_386_n N_A_324_373#_c_1195_n 0.0247711f $X=4.105 $Y=2.115
+ $X2=0 $Y2=0
cc_390 N_A_386_23#_c_381_n N_A_324_373#_c_1219_n 0.00333007f $X=2.245 $Y=1.79
+ $X2=0 $Y2=0
cc_391 N_A_386_23#_c_381_n N_A_324_373#_c_1220_n 0.00406253f $X=2.245 $Y=1.79
+ $X2=0 $Y2=0
cc_392 N_A_386_23#_M1021_s N_A_321_77#_c_1312_n 0.00721616f $X=3.78 $Y=0.445
+ $X2=0 $Y2=0
cc_393 N_A_386_23#_c_369_n N_A_321_77#_c_1312_n 8.21484e-19 $X=2.995 $Y=0.19
+ $X2=0 $Y2=0
cc_394 N_A_386_23#_M1011_g N_A_321_77#_c_1312_n 0.0143626f $X=3.07 $Y=0.925
+ $X2=0 $Y2=0
cc_395 N_A_386_23#_c_374_n N_A_321_77#_c_1312_n 0.00309509f $X=3.205 $Y=1.79
+ $X2=0 $Y2=0
cc_396 N_A_386_23#_c_375_n N_A_321_77#_c_1312_n 0.0162608f $X=3.6 $Y=1.54 $X2=0
+ $Y2=0
cc_397 N_A_386_23#_c_377_n N_A_321_77#_c_1312_n 0.0143583f $X=3.77 $Y=1.04 $X2=0
+ $Y2=0
cc_398 N_A_386_23#_c_378_n N_A_321_77#_c_1312_n 0.0189364f $X=3.925 $Y=1.04
+ $X2=0 $Y2=0
cc_399 N_A_386_23#_c_374_n N_A_321_77#_c_1339_n 0.0111604f $X=3.205 $Y=1.79
+ $X2=0 $Y2=0
cc_400 N_A_386_23#_c_375_n N_A_321_77#_c_1339_n 0.0088044f $X=3.6 $Y=1.54 $X2=0
+ $Y2=0
cc_401 N_A_386_23#_c_384_n N_A_321_77#_c_1339_n 0.00251225f $X=3.685 $Y=1.95
+ $X2=0 $Y2=0
cc_402 N_A_386_23#_c_385_n N_A_321_77#_c_1339_n 0.00707185f $X=3.77 $Y=2.075
+ $X2=0 $Y2=0
cc_403 N_A_386_23#_M1022_s N_A_321_77#_c_1318_n 0.00688029f $X=3.96 $Y=1.84
+ $X2=0 $Y2=0
cc_404 N_A_386_23#_c_374_n N_A_321_77#_c_1318_n 0.0105228f $X=3.205 $Y=1.79
+ $X2=0 $Y2=0
cc_405 N_A_386_23#_c_375_n N_A_321_77#_c_1318_n 0.00439452f $X=3.6 $Y=1.54 $X2=0
+ $Y2=0
cc_406 N_A_386_23#_c_385_n N_A_321_77#_c_1318_n 0.0129068f $X=3.77 $Y=2.075
+ $X2=0 $Y2=0
cc_407 N_A_386_23#_c_386_n N_A_321_77#_c_1318_n 0.0301886f $X=4.105 $Y=2.115
+ $X2=0 $Y2=0
cc_408 N_A_386_23#_c_374_n N_A_321_77#_c_1329_n 5.24026e-19 $X=3.205 $Y=1.79
+ $X2=0 $Y2=0
cc_409 N_A_386_23#_c_376_n N_A_321_77#_c_1313_n 0.00632457f $X=3.685 $Y=1.375
+ $X2=0 $Y2=0
cc_410 N_A_386_23#_c_384_n N_A_321_77#_c_1313_n 0.0026521f $X=3.685 $Y=1.95
+ $X2=0 $Y2=0
cc_411 N_A_386_23#_c_378_n N_A_321_77#_c_1313_n 0.00409526f $X=3.925 $Y=1.04
+ $X2=0 $Y2=0
cc_412 N_A_386_23#_c_386_n N_A_321_77#_c_1313_n 0.0116478f $X=4.105 $Y=2.115
+ $X2=0 $Y2=0
cc_413 N_A_386_23#_M1006_g N_A_321_77#_c_1314_n 0.00590709f $X=2.005 $Y=0.815
+ $X2=0 $Y2=0
cc_414 N_A_386_23#_M1006_g N_A_321_77#_c_1315_n 0.00973001f $X=2.005 $Y=0.815
+ $X2=0 $Y2=0
cc_415 N_A_386_23#_c_369_n N_A_321_77#_c_1315_n 0.00193544f $X=2.995 $Y=0.19
+ $X2=0 $Y2=0
cc_416 N_A_386_23#_c_371_n N_A_321_77#_c_1315_n 6.21063e-19 $X=2.245 $Y=1.47
+ $X2=0 $Y2=0
cc_417 N_A_386_23#_M1011_g N_A_321_77#_c_1316_n 2.29766e-19 $X=3.07 $Y=0.925
+ $X2=0 $Y2=0
cc_418 N_A_386_23#_c_378_n N_A_321_77#_c_1317_n 0.00363019f $X=3.925 $Y=1.04
+ $X2=0 $Y2=0
cc_419 N_A_386_23#_c_370_n N_VGND_c_1509_n 0.0257161f $X=2.08 $Y=0.19 $X2=0
+ $Y2=0
cc_420 N_A_386_23#_c_369_n N_VGND_c_1514_n 0.0275023f $X=2.995 $Y=0.19 $X2=0
+ $Y2=0
cc_421 N_A_386_23#_c_370_n N_VGND_c_1514_n 0.00588169f $X=2.08 $Y=0.19 $X2=0
+ $Y2=0
cc_422 N_B_c_502_n N_A_1024_300#_M1027_g 0.00132172f $X=4.14 $Y=1.557 $X2=0
+ $Y2=0
cc_423 N_B_c_514_n N_A_1024_300#_c_650_n 5.47802e-19 $X=4.33 $Y=1.765 $X2=0
+ $Y2=0
cc_424 N_B_c_502_n N_A_1024_300#_c_650_n 0.00253621f $X=4.14 $Y=1.557 $X2=0
+ $Y2=0
cc_425 N_B_c_509_n N_A_27_373#_c_971_n 3.74241e-19 $X=2.695 $Y=2.67 $X2=0 $Y2=0
cc_426 N_B_c_503_n N_A_27_373#_c_972_n 4.31853e-19 $X=1.545 $Y=2.87 $X2=0 $Y2=0
cc_427 N_B_M1007_g N_A_27_373#_c_972_n 0.00652967f $X=1.545 $Y=2.285 $X2=0 $Y2=0
cc_428 N_B_M1025_g N_A_27_373#_c_968_n 0.0103289f $X=1.53 $Y=0.705 $X2=0 $Y2=0
cc_429 N_B_M1004_g N_A_27_373#_c_969_n 0.00447538f $X=2.62 $Y=0.925 $X2=0 $Y2=0
cc_430 N_B_M1007_g N_A_27_373#_c_975_n 4.51847e-19 $X=1.545 $Y=2.285 $X2=0 $Y2=0
cc_431 N_B_c_509_n N_A_27_373#_c_975_n 0.00412427f $X=2.695 $Y=2.67 $X2=0 $Y2=0
cc_432 N_B_c_510_n N_A_27_373#_c_975_n 0.00466697f $X=2.695 $Y=3.075 $X2=0 $Y2=0
cc_433 N_B_M1020_g N_A_27_373#_c_975_n 0.00839352f $X=2.695 $Y=2.185 $X2=0 $Y2=0
cc_434 N_B_c_500_n N_A_27_373#_c_975_n 0.00136831f $X=2.695 $Y=1.715 $X2=0 $Y2=0
cc_435 N_B_c_497_n N_A_27_373#_c_996_n 4.16621e-19 $X=1.545 $Y=1.79 $X2=0 $Y2=0
cc_436 N_B_M1007_g N_A_27_373#_c_996_n 0.00640406f $X=1.545 $Y=2.285 $X2=0 $Y2=0
cc_437 N_B_M1007_g N_A_27_373#_c_1006_n 0.0036739f $X=1.545 $Y=2.285 $X2=0 $Y2=0
cc_438 N_B_M1025_g N_A_27_373#_c_970_n 0.00413342f $X=1.53 $Y=0.705 $X2=0 $Y2=0
cc_439 N_B_c_497_n N_A_27_373#_c_970_n 0.00517832f $X=1.545 $Y=1.79 $X2=0 $Y2=0
cc_440 N_B_M1007_g N_A_27_373#_c_970_n 0.0197153f $X=1.545 $Y=2.285 $X2=0 $Y2=0
cc_441 N_B_c_504_n N_VPWR_c_1078_n 2.99406e-19 $X=1.545 $Y=3.075 $X2=0 $Y2=0
cc_442 N_B_c_508_n N_VPWR_c_1078_n 0.00248898f $X=1.635 $Y=3.15 $X2=0 $Y2=0
cc_443 N_B_c_512_n N_VPWR_c_1079_n 0.00232909f $X=3.735 $Y=3.15 $X2=0 $Y2=0
cc_444 N_B_c_513_n N_VPWR_c_1079_n 0.00167614f $X=3.81 $Y=3.075 $X2=0 $Y2=0
cc_445 N_B_c_514_n N_VPWR_c_1079_n 0.00992346f $X=4.33 $Y=1.765 $X2=0 $Y2=0
cc_446 N_B_c_508_n N_VPWR_c_1087_n 0.055167f $X=1.635 $Y=3.15 $X2=0 $Y2=0
cc_447 N_B_c_514_n N_VPWR_c_1087_n 0.00413917f $X=4.33 $Y=1.765 $X2=0 $Y2=0
cc_448 N_B_c_507_n N_VPWR_c_1077_n 0.0228018f $X=2.605 $Y=3.15 $X2=0 $Y2=0
cc_449 N_B_c_508_n N_VPWR_c_1077_n 0.00675277f $X=1.635 $Y=3.15 $X2=0 $Y2=0
cc_450 N_B_c_512_n N_VPWR_c_1077_n 0.0296846f $X=3.735 $Y=3.15 $X2=0 $Y2=0
cc_451 N_B_c_514_n N_VPWR_c_1077_n 0.00403814f $X=4.33 $Y=1.765 $X2=0 $Y2=0
cc_452 N_B_c_516_n N_VPWR_c_1077_n 0.00442127f $X=2.695 $Y=3.15 $X2=0 $Y2=0
cc_453 N_B_c_497_n N_A_324_373#_c_1192_n 3.43991e-19 $X=1.545 $Y=1.79 $X2=0
+ $Y2=0
cc_454 N_B_M1007_g N_A_324_373#_c_1192_n 5.15093e-19 $X=1.545 $Y=2.285 $X2=0
+ $Y2=0
cc_455 N_B_M1020_g N_A_324_373#_c_1192_n 8.10277e-19 $X=2.695 $Y=2.185 $X2=0
+ $Y2=0
cc_456 N_B_c_500_n N_A_324_373#_c_1192_n 6.40682e-19 $X=2.695 $Y=1.715 $X2=0
+ $Y2=0
cc_457 N_B_M1004_g N_A_324_373#_c_1184_n 0.00418594f $X=2.62 $Y=0.925 $X2=0
+ $Y2=0
cc_458 N_B_c_500_n N_A_324_373#_c_1184_n 0.00716062f $X=2.695 $Y=1.715 $X2=0
+ $Y2=0
cc_459 N_B_M1025_g N_A_324_373#_c_1185_n 4.38234e-19 $X=1.53 $Y=0.705 $X2=0
+ $Y2=0
cc_460 N_B_M1004_g N_A_324_373#_c_1186_n 0.00852261f $X=2.62 $Y=0.925 $X2=0
+ $Y2=0
cc_461 N_B_M1004_g N_A_324_373#_c_1210_n 0.00693619f $X=2.62 $Y=0.925 $X2=0
+ $Y2=0
cc_462 N_B_c_500_n N_A_324_373#_c_1210_n 0.00106073f $X=2.695 $Y=1.715 $X2=0
+ $Y2=0
cc_463 N_B_c_509_n N_A_324_373#_c_1195_n 3.42112e-19 $X=2.695 $Y=2.67 $X2=0
+ $Y2=0
cc_464 N_B_M1020_g N_A_324_373#_c_1195_n 0.00766022f $X=2.695 $Y=2.185 $X2=0
+ $Y2=0
cc_465 N_B_c_514_n N_A_324_373#_c_1195_n 0.00915107f $X=4.33 $Y=1.765 $X2=0
+ $Y2=0
cc_466 N_B_c_500_n N_A_324_373#_c_1195_n 0.00239994f $X=2.695 $Y=1.715 $X2=0
+ $Y2=0
cc_467 N_B_c_501_n N_A_324_373#_c_1195_n 0.00263994f $X=4.105 $Y=1.515 $X2=0
+ $Y2=0
cc_468 N_B_c_502_n N_A_324_373#_c_1195_n 3.7045e-19 $X=4.14 $Y=1.557 $X2=0 $Y2=0
cc_469 N_B_M1020_g N_A_324_373#_c_1219_n 4.63222e-19 $X=2.695 $Y=2.185 $X2=0
+ $Y2=0
cc_470 N_B_M1007_g N_A_324_373#_c_1220_n 5.55941e-19 $X=1.545 $Y=2.285 $X2=0
+ $Y2=0
cc_471 N_B_M1020_g N_A_324_373#_c_1220_n 6.25756e-19 $X=2.695 $Y=2.185 $X2=0
+ $Y2=0
cc_472 N_B_M1021_g N_A_321_77#_c_1312_n 0.017085f $X=4.14 $Y=0.815 $X2=0 $Y2=0
cc_473 N_B_c_501_n N_A_321_77#_c_1312_n 0.00418899f $X=4.105 $Y=1.515 $X2=0
+ $Y2=0
cc_474 N_B_c_502_n N_A_321_77#_c_1312_n 0.00409034f $X=4.14 $Y=1.557 $X2=0 $Y2=0
cc_475 N_B_M1020_g N_A_321_77#_c_1339_n 0.00749405f $X=2.695 $Y=2.185 $X2=0
+ $Y2=0
cc_476 N_B_c_513_n N_A_321_77#_c_1339_n 0.00111742f $X=3.81 $Y=3.075 $X2=0 $Y2=0
cc_477 N_B_c_512_n N_A_321_77#_c_1318_n 0.00102485f $X=3.735 $Y=3.15 $X2=0 $Y2=0
cc_478 N_B_c_513_n N_A_321_77#_c_1318_n 0.0131221f $X=3.81 $Y=3.075 $X2=0 $Y2=0
cc_479 N_B_c_514_n N_A_321_77#_c_1318_n 0.014514f $X=4.33 $Y=1.765 $X2=0 $Y2=0
cc_480 N_B_M1020_g N_A_321_77#_c_1329_n 0.00137779f $X=2.695 $Y=2.185 $X2=0
+ $Y2=0
cc_481 N_B_M1021_g N_A_321_77#_c_1313_n 0.00689761f $X=4.14 $Y=0.815 $X2=0 $Y2=0
cc_482 N_B_c_514_n N_A_321_77#_c_1313_n 0.0115781f $X=4.33 $Y=1.765 $X2=0 $Y2=0
cc_483 N_B_c_501_n N_A_321_77#_c_1313_n 0.0322749f $X=4.105 $Y=1.515 $X2=0 $Y2=0
cc_484 N_B_c_502_n N_A_321_77#_c_1313_n 0.00633841f $X=4.14 $Y=1.557 $X2=0 $Y2=0
cc_485 N_B_M1004_g N_A_321_77#_c_1314_n 8.232e-19 $X=2.62 $Y=0.925 $X2=0 $Y2=0
cc_486 N_B_M1004_g N_A_321_77#_c_1315_n 0.00343798f $X=2.62 $Y=0.925 $X2=0 $Y2=0
cc_487 N_B_M1004_g N_A_321_77#_c_1316_n 0.00788426f $X=2.62 $Y=0.925 $X2=0 $Y2=0
cc_488 N_B_M1021_g N_A_321_77#_c_1317_n 0.0123212f $X=4.14 $Y=0.815 $X2=0 $Y2=0
cc_489 N_B_M1021_g N_VGND_c_1502_n 0.00546687f $X=4.14 $Y=0.815 $X2=0 $Y2=0
cc_490 N_B_M1025_g N_VGND_c_1509_n 0.00388395f $X=1.53 $Y=0.705 $X2=0 $Y2=0
cc_491 N_B_M1021_g N_VGND_c_1509_n 0.00399972f $X=4.14 $Y=0.815 $X2=0 $Y2=0
cc_492 N_B_M1025_g N_VGND_c_1514_n 0.0054106f $X=1.53 $Y=0.705 $X2=0 $Y2=0
cc_493 N_B_M1021_g N_VGND_c_1514_n 0.0052212f $X=4.14 $Y=0.815 $X2=0 $Y2=0
cc_494 N_A_1024_300#_M1027_g N_C_M1012_g 0.025185f $X=5.21 $Y=0.69 $X2=0 $Y2=0
cc_495 N_A_1024_300#_c_652_n N_C_M1012_g 6.18081e-19 $X=6.5 $Y=1.55 $X2=0 $Y2=0
cc_496 N_A_1024_300#_c_654_n N_C_M1012_g 6.75097e-19 $X=6.555 $Y=1.085 $X2=0
+ $Y2=0
cc_497 N_A_1024_300#_c_650_n N_C_c_732_n 0.00966088f $X=5.34 $Y=1.915 $X2=0
+ $Y2=0
cc_498 N_A_1024_300#_c_651_n N_C_c_732_n 0.0159955f $X=6.39 $Y=1.635 $X2=0 $Y2=0
cc_499 N_A_1024_300#_c_652_n N_C_c_732_n 0.00100646f $X=6.5 $Y=1.55 $X2=0 $Y2=0
cc_500 N_A_1024_300#_c_658_n N_C_c_732_n 0.00537101f $X=6.525 $Y=1.99 $X2=0
+ $Y2=0
cc_501 N_A_1024_300#_c_653_n N_C_c_732_n 3.42292e-19 $X=5.45 $Y=1.665 $X2=0
+ $Y2=0
cc_502 N_A_1024_300#_c_650_n N_C_c_739_n 0.0266962f $X=5.34 $Y=1.915 $X2=0 $Y2=0
cc_503 N_A_1024_300#_c_658_n N_C_c_739_n 0.00153883f $X=6.525 $Y=1.99 $X2=0
+ $Y2=0
cc_504 N_A_1024_300#_c_661_n N_C_c_739_n 0.00104631f $X=6.795 $Y=2.235 $X2=0
+ $Y2=0
cc_505 N_A_1024_300#_c_651_n N_C_c_733_n 0.0113645f $X=6.39 $Y=1.635 $X2=0 $Y2=0
cc_506 N_A_1024_300#_c_652_n N_C_c_733_n 0.0202007f $X=6.5 $Y=1.55 $X2=0 $Y2=0
cc_507 N_A_1024_300#_c_661_n N_C_c_733_n 0.00325694f $X=6.795 $Y=2.235 $X2=0
+ $Y2=0
cc_508 N_A_1024_300#_c_651_n N_C_c_734_n 0.00546398f $X=6.39 $Y=1.635 $X2=0
+ $Y2=0
cc_509 N_A_1024_300#_c_652_n N_C_c_735_n 0.00567584f $X=6.5 $Y=1.55 $X2=0 $Y2=0
cc_510 N_A_1024_300#_c_654_n N_C_c_735_n 0.00308441f $X=6.555 $Y=1.085 $X2=0
+ $Y2=0
cc_511 N_A_1024_300#_c_652_n N_C_c_736_n 6.32325e-19 $X=6.5 $Y=1.55 $X2=0 $Y2=0
cc_512 N_A_1024_300#_c_658_n N_C_c_736_n 0.00592164f $X=6.525 $Y=1.99 $X2=0
+ $Y2=0
cc_513 N_A_1024_300#_c_655_n N_C_c_736_n 0.00198816f $X=6.5 $Y=1.635 $X2=0 $Y2=0
cc_514 N_A_1024_300#_c_661_n N_C_c_736_n 0.0124065f $X=6.795 $Y=2.235 $X2=0
+ $Y2=0
cc_515 N_A_1024_300#_c_652_n N_C_c_737_n 0.0147109f $X=6.5 $Y=1.55 $X2=0 $Y2=0
cc_516 N_A_1024_300#_c_658_n N_C_c_737_n 0.00471921f $X=6.525 $Y=1.99 $X2=0
+ $Y2=0
cc_517 N_A_1024_300#_c_655_n N_C_c_737_n 0.0145003f $X=6.5 $Y=1.635 $X2=0 $Y2=0
cc_518 N_A_1024_300#_c_661_n N_C_c_737_n 0.0110904f $X=6.795 $Y=2.235 $X2=0
+ $Y2=0
cc_519 N_A_1024_300#_M1027_g N_A_1057_74#_c_812_n 0.00371279f $X=5.21 $Y=0.69
+ $X2=0 $Y2=0
cc_520 N_A_1024_300#_c_661_n N_A_1057_74#_c_824_n 0.0197653f $X=6.795 $Y=2.235
+ $X2=0 $Y2=0
cc_521 N_A_1024_300#_M1017_s N_A_1057_74#_c_814_n 0.00131178f $X=6.41 $Y=0.81
+ $X2=0 $Y2=0
cc_522 N_A_1024_300#_c_654_n N_A_1057_74#_c_814_n 0.0125593f $X=6.555 $Y=1.085
+ $X2=0 $Y2=0
cc_523 N_A_1024_300#_M1017_s N_A_1057_74#_c_815_n 9.85725e-19 $X=6.41 $Y=0.81
+ $X2=0 $Y2=0
cc_524 N_A_1024_300#_c_654_n N_A_1057_74#_c_815_n 0.00979215f $X=6.555 $Y=1.085
+ $X2=0 $Y2=0
cc_525 N_A_1024_300#_c_661_n N_A_1057_74#_c_825_n 0.0160153f $X=6.795 $Y=2.235
+ $X2=0 $Y2=0
cc_526 N_A_1024_300#_c_650_n N_A_1057_74#_c_827_n 0.00663705f $X=5.34 $Y=1.915
+ $X2=0 $Y2=0
cc_527 N_A_1024_300#_c_650_n N_VPWR_c_1079_n 0.0057683f $X=5.34 $Y=1.915 $X2=0
+ $Y2=0
cc_528 N_A_1024_300#_c_650_n N_VPWR_c_1088_n 0.00487664f $X=5.34 $Y=1.915 $X2=0
+ $Y2=0
cc_529 N_A_1024_300#_c_650_n N_VPWR_c_1077_n 0.00505379f $X=5.34 $Y=1.915 $X2=0
+ $Y2=0
cc_530 N_A_1024_300#_M1027_g N_A_324_373#_c_1187_n 0.00287206f $X=5.21 $Y=0.69
+ $X2=0 $Y2=0
cc_531 N_A_1024_300#_c_650_n N_A_324_373#_c_1187_n 0.00708613f $X=5.34 $Y=1.915
+ $X2=0 $Y2=0
cc_532 N_A_1024_300#_c_653_n N_A_324_373#_c_1187_n 0.0179619f $X=5.45 $Y=1.665
+ $X2=0 $Y2=0
cc_533 N_A_1024_300#_M1027_g N_A_324_373#_c_1189_n 8.88219e-19 $X=5.21 $Y=0.69
+ $X2=0 $Y2=0
cc_534 N_A_1024_300#_c_651_n N_A_324_373#_c_1189_n 0.0375039f $X=6.39 $Y=1.635
+ $X2=0 $Y2=0
cc_535 N_A_1024_300#_c_652_n N_A_324_373#_c_1189_n 0.0135138f $X=6.5 $Y=1.55
+ $X2=0 $Y2=0
cc_536 N_A_1024_300#_M1027_g N_A_324_373#_c_1190_n 8.1639e-19 $X=5.21 $Y=0.69
+ $X2=0 $Y2=0
cc_537 N_A_1024_300#_c_654_n N_A_324_373#_c_1190_n 0.0120836f $X=6.555 $Y=1.085
+ $X2=0 $Y2=0
cc_538 N_A_1024_300#_M1027_g N_A_324_373#_c_1191_n 0.0163205f $X=5.21 $Y=0.69
+ $X2=0 $Y2=0
cc_539 N_A_1024_300#_c_650_n N_A_324_373#_c_1191_n 0.00484029f $X=5.34 $Y=1.915
+ $X2=0 $Y2=0
cc_540 N_A_1024_300#_c_653_n N_A_324_373#_c_1191_n 0.0375039f $X=5.45 $Y=1.665
+ $X2=0 $Y2=0
cc_541 N_A_1024_300#_c_650_n N_A_324_373#_c_1196_n 0.00273737f $X=5.34 $Y=1.915
+ $X2=0 $Y2=0
cc_542 N_A_1024_300#_c_653_n N_A_324_373#_c_1196_n 0.00182723f $X=5.45 $Y=1.665
+ $X2=0 $Y2=0
cc_543 N_A_1024_300#_c_650_n N_A_324_373#_c_1197_n 0.011034f $X=5.34 $Y=1.915
+ $X2=0 $Y2=0
cc_544 N_A_1024_300#_c_653_n N_A_324_373#_c_1197_n 0.0113204f $X=5.45 $Y=1.665
+ $X2=0 $Y2=0
cc_545 N_A_1024_300#_M1027_g N_A_321_77#_c_1313_n 0.00491664f $X=5.21 $Y=0.69
+ $X2=0 $Y2=0
cc_546 N_A_1024_300#_c_650_n N_A_321_77#_c_1313_n 0.00229792f $X=5.34 $Y=1.915
+ $X2=0 $Y2=0
cc_547 N_A_1024_300#_c_650_n N_A_321_77#_c_1320_n 0.0170812f $X=5.34 $Y=1.915
+ $X2=0 $Y2=0
cc_548 N_A_1024_300#_c_651_n N_A_321_77#_c_1320_n 0.0137123f $X=6.39 $Y=1.635
+ $X2=0 $Y2=0
cc_549 N_A_1024_300#_c_653_n N_A_321_77#_c_1320_n 0.00368243f $X=5.45 $Y=1.665
+ $X2=0 $Y2=0
cc_550 N_A_1024_300#_c_661_n N_A_321_77#_c_1320_n 0.00981823f $X=6.795 $Y=2.235
+ $X2=0 $Y2=0
cc_551 N_A_1024_300#_c_650_n N_A_321_77#_c_1321_n 0.0018396f $X=5.34 $Y=1.915
+ $X2=0 $Y2=0
cc_552 N_A_1024_300#_c_651_n N_A_321_77#_c_1321_n 0.0158088f $X=6.39 $Y=1.635
+ $X2=0 $Y2=0
cc_553 N_A_1024_300#_c_658_n N_A_321_77#_c_1321_n 0.00155139f $X=6.525 $Y=1.99
+ $X2=0 $Y2=0
cc_554 N_A_1024_300#_c_661_n N_A_321_77#_c_1321_n 0.0332586f $X=6.795 $Y=2.235
+ $X2=0 $Y2=0
cc_555 N_A_1024_300#_M1027_g N_A_321_77#_c_1317_n 0.00867986f $X=5.21 $Y=0.69
+ $X2=0 $Y2=0
cc_556 N_A_1024_300#_c_650_n N_A_321_77#_c_1387_n 4.98334e-19 $X=5.34 $Y=1.915
+ $X2=0 $Y2=0
cc_557 N_A_1024_300#_M1027_g N_VGND_c_1502_n 0.00294228f $X=5.21 $Y=0.69 $X2=0
+ $Y2=0
cc_558 N_A_1024_300#_M1027_g N_VGND_c_1503_n 0.00433139f $X=5.21 $Y=0.69 $X2=0
+ $Y2=0
cc_559 N_A_1024_300#_M1027_g N_VGND_c_1514_n 0.00823742f $X=5.21 $Y=0.69 $X2=0
+ $Y2=0
cc_560 N_C_M1012_g N_A_1057_74#_c_811_n 0.014965f $X=5.765 $Y=0.69 $X2=0 $Y2=0
cc_561 N_C_c_739_n N_A_1057_74#_c_824_n 0.007953f $X=5.96 $Y=1.915 $X2=0 $Y2=0
cc_562 N_C_c_736_n N_A_1057_74#_c_824_n 0.00527616f $X=7.02 $Y=1.765 $X2=0 $Y2=0
cc_563 N_C_M1012_g N_A_1057_74#_c_813_n 0.00287215f $X=5.765 $Y=0.69 $X2=0 $Y2=0
cc_564 N_C_c_733_n N_A_1057_74#_c_814_n 3.54962e-19 $X=6.695 $Y=1.425 $X2=0
+ $Y2=0
cc_565 N_C_c_735_n N_A_1057_74#_c_814_n 0.0148447f $X=6.77 $Y=1.35 $X2=0 $Y2=0
cc_566 N_C_c_737_n N_A_1057_74#_c_814_n 0.00258247f $X=6.945 $Y=1.515 $X2=0
+ $Y2=0
cc_567 N_C_c_733_n N_A_1057_74#_c_815_n 0.00209722f $X=6.695 $Y=1.425 $X2=0
+ $Y2=0
cc_568 N_C_c_736_n N_A_1057_74#_c_846_n 3.39557e-19 $X=7.02 $Y=1.765 $X2=0 $Y2=0
cc_569 N_C_c_737_n N_A_1057_74#_c_846_n 0.00367584f $X=6.945 $Y=1.515 $X2=0
+ $Y2=0
cc_570 N_C_c_736_n N_A_1057_74#_c_848_n 0.0012636f $X=7.02 $Y=1.765 $X2=0 $Y2=0
cc_571 N_C_c_737_n N_A_1057_74#_c_848_n 0.0135553f $X=6.945 $Y=1.515 $X2=0 $Y2=0
cc_572 N_C_c_736_n N_A_1057_74#_c_825_n 0.0119226f $X=7.02 $Y=1.765 $X2=0 $Y2=0
cc_573 N_C_c_735_n N_A_1057_74#_c_816_n 0.00395023f $X=6.77 $Y=1.35 $X2=0 $Y2=0
cc_574 N_C_c_736_n N_A_1057_74#_c_826_n 0.00745017f $X=7.02 $Y=1.765 $X2=0 $Y2=0
cc_575 N_C_c_737_n N_A_1057_74#_c_826_n 0.007086f $X=6.945 $Y=1.515 $X2=0 $Y2=0
cc_576 N_C_c_739_n N_A_1057_74#_c_827_n 0.00513011f $X=5.96 $Y=1.915 $X2=0 $Y2=0
cc_577 N_C_c_736_n N_A_1057_74#_c_817_n 0.00122161f $X=7.02 $Y=1.765 $X2=0 $Y2=0
cc_578 N_C_c_737_n N_A_1057_74#_c_817_n 0.0215512f $X=6.945 $Y=1.515 $X2=0 $Y2=0
cc_579 N_C_c_736_n N_A_1057_74#_c_818_n 0.0209673f $X=7.02 $Y=1.765 $X2=0 $Y2=0
cc_580 N_C_c_737_n N_A_1057_74#_c_818_n 4.00288e-19 $X=6.945 $Y=1.515 $X2=0
+ $Y2=0
cc_581 N_C_c_736_n N_VPWR_c_1081_n 8.86484e-19 $X=7.02 $Y=1.765 $X2=0 $Y2=0
cc_582 N_C_c_739_n N_VPWR_c_1088_n 7.08494e-19 $X=5.96 $Y=1.915 $X2=0 $Y2=0
cc_583 N_C_M1012_g N_A_324_373#_c_1189_n 0.0147025f $X=5.765 $Y=0.69 $X2=0 $Y2=0
cc_584 N_C_c_733_n N_A_324_373#_c_1189_n 0.00362102f $X=6.695 $Y=1.425 $X2=0
+ $Y2=0
cc_585 N_C_c_734_n N_A_324_373#_c_1189_n 0.00755929f $X=6.05 $Y=1.425 $X2=0
+ $Y2=0
cc_586 N_C_M1012_g N_A_324_373#_c_1190_n 0.0112653f $X=5.765 $Y=0.69 $X2=0 $Y2=0
cc_587 N_C_c_734_n N_A_324_373#_c_1190_n 0.00111739f $X=6.05 $Y=1.425 $X2=0
+ $Y2=0
cc_588 N_C_c_735_n N_A_324_373#_c_1190_n 0.0035702f $X=6.77 $Y=1.35 $X2=0 $Y2=0
cc_589 N_C_c_739_n N_A_324_373#_c_1197_n 0.00116795f $X=5.96 $Y=1.915 $X2=0
+ $Y2=0
cc_590 N_C_c_739_n N_A_321_77#_c_1320_n 0.0153593f $X=5.96 $Y=1.915 $X2=0 $Y2=0
cc_591 N_C_c_736_n N_A_321_77#_c_1320_n 0.00281324f $X=7.02 $Y=1.765 $X2=0 $Y2=0
cc_592 N_C_c_739_n N_A_321_77#_c_1321_n 0.0102291f $X=5.96 $Y=1.915 $X2=0 $Y2=0
cc_593 N_C_c_736_n N_A_321_77#_c_1321_n 5.12614e-19 $X=7.02 $Y=1.765 $X2=0 $Y2=0
cc_594 N_C_M1012_g N_A_321_77#_c_1317_n 2.05732e-19 $X=5.765 $Y=0.69 $X2=0 $Y2=0
cc_595 N_C_M1012_g N_VGND_c_1503_n 0.00278271f $X=5.765 $Y=0.69 $X2=0 $Y2=0
cc_596 N_C_c_735_n N_VGND_c_1503_n 5.51389e-19 $X=6.77 $Y=1.35 $X2=0 $Y2=0
cc_597 N_C_c_735_n N_VGND_c_1505_n 7.66361e-19 $X=6.77 $Y=1.35 $X2=0 $Y2=0
cc_598 N_C_M1012_g N_VGND_c_1514_n 0.00359569f $X=5.765 $Y=0.69 $X2=0 $Y2=0
cc_599 N_A_1057_74#_c_825_n N_VPWR_M1018_d 0.00836264f $X=7.222 $Y=2.905 $X2=0
+ $Y2=0
cc_600 N_A_1057_74#_c_826_n N_VPWR_M1018_d 0.00390247f $X=7.405 $Y=1.95 $X2=0
+ $Y2=0
cc_601 N_A_1057_74#_c_861_p N_VPWR_M1018_d 0.0188982f $X=7.405 $Y=2.035 $X2=0
+ $Y2=0
cc_602 N_A_1057_74#_c_820_n N_VPWR_c_1080_n 0.0131912f $X=8.22 $Y=1.765 $X2=0
+ $Y2=0
cc_603 N_A_1057_74#_c_824_n N_VPWR_c_1080_n 0.0156625f $X=7.13 $Y=2.99 $X2=0
+ $Y2=0
cc_604 N_A_1057_74#_c_825_n N_VPWR_c_1081_n 0.00750254f $X=7.222 $Y=2.905 $X2=0
+ $Y2=0
cc_605 N_A_1057_74#_c_826_n N_VPWR_c_1081_n 0.00774637f $X=7.405 $Y=1.95 $X2=0
+ $Y2=0
cc_606 N_A_1057_74#_c_866_p N_VPWR_c_1081_n 0.0339891f $X=8.165 $Y=1.505 $X2=0
+ $Y2=0
cc_607 N_A_1057_74#_c_861_p N_VPWR_c_1081_n 0.0125379f $X=7.405 $Y=2.035 $X2=0
+ $Y2=0
cc_608 N_A_1057_74#_c_818_n N_VPWR_c_1081_n 0.00979007f $X=8.13 $Y=1.505 $X2=0
+ $Y2=0
cc_609 N_A_1057_74#_c_820_n N_VPWR_c_1082_n 0.00445602f $X=8.22 $Y=1.765 $X2=0
+ $Y2=0
cc_610 N_A_1057_74#_c_821_n N_VPWR_c_1082_n 0.00411612f $X=8.67 $Y=1.765 $X2=0
+ $Y2=0
cc_611 N_A_1057_74#_c_821_n N_VPWR_c_1083_n 0.00615208f $X=8.67 $Y=1.765 $X2=0
+ $Y2=0
cc_612 N_A_1057_74#_c_822_n N_VPWR_c_1083_n 0.00665541f $X=9.12 $Y=1.765 $X2=0
+ $Y2=0
cc_613 N_A_1057_74#_c_819_n N_VPWR_c_1083_n 0.00439943f $X=9.57 $Y=1.552 $X2=0
+ $Y2=0
cc_614 N_A_1057_74#_c_823_n N_VPWR_c_1085_n 0.00963415f $X=9.57 $Y=1.765 $X2=0
+ $Y2=0
cc_615 N_A_1057_74#_c_825_n N_VPWR_c_1147_n 0.0502413f $X=7.222 $Y=2.905 $X2=0
+ $Y2=0
cc_616 N_A_1057_74#_c_866_p N_VPWR_c_1147_n 0.00580119f $X=8.165 $Y=1.505 $X2=0
+ $Y2=0
cc_617 N_A_1057_74#_c_818_n N_VPWR_c_1147_n 0.00332899f $X=8.13 $Y=1.505 $X2=0
+ $Y2=0
cc_618 N_A_1057_74#_c_824_n N_VPWR_c_1088_n 0.097943f $X=7.13 $Y=2.99 $X2=0
+ $Y2=0
cc_619 N_A_1057_74#_c_827_n N_VPWR_c_1088_n 0.0223614f $X=5.65 $Y=2.895 $X2=0
+ $Y2=0
cc_620 N_A_1057_74#_c_822_n N_VPWR_c_1089_n 0.00445602f $X=9.12 $Y=1.765 $X2=0
+ $Y2=0
cc_621 N_A_1057_74#_c_823_n N_VPWR_c_1089_n 0.00417277f $X=9.57 $Y=1.765 $X2=0
+ $Y2=0
cc_622 N_A_1057_74#_c_820_n N_VPWR_c_1077_n 0.00861719f $X=8.22 $Y=1.765 $X2=0
+ $Y2=0
cc_623 N_A_1057_74#_c_821_n N_VPWR_c_1077_n 0.00747529f $X=8.67 $Y=1.765 $X2=0
+ $Y2=0
cc_624 N_A_1057_74#_c_822_n N_VPWR_c_1077_n 0.00857589f $X=9.12 $Y=1.765 $X2=0
+ $Y2=0
cc_625 N_A_1057_74#_c_823_n N_VPWR_c_1077_n 0.00769383f $X=9.57 $Y=1.765 $X2=0
+ $Y2=0
cc_626 N_A_1057_74#_c_824_n N_VPWR_c_1077_n 0.0566295f $X=7.13 $Y=2.99 $X2=0
+ $Y2=0
cc_627 N_A_1057_74#_c_827_n N_VPWR_c_1077_n 0.0125377f $X=5.65 $Y=2.895 $X2=0
+ $Y2=0
cc_628 N_A_1057_74#_c_811_n N_A_324_373#_M1012_d 0.00294181f $X=6.33 $Y=0.34
+ $X2=0 $Y2=0
cc_629 N_A_1057_74#_c_810_n N_A_324_373#_c_1189_n 0.0200764f $X=5.495 $Y=0.515
+ $X2=0 $Y2=0
cc_630 N_A_1057_74#_c_811_n N_A_324_373#_c_1190_n 0.0204002f $X=6.33 $Y=0.34
+ $X2=0 $Y2=0
cc_631 N_A_1057_74#_c_813_n N_A_324_373#_c_1190_n 0.00511586f $X=6.415 $Y=0.66
+ $X2=0 $Y2=0
cc_632 N_A_1057_74#_c_815_n N_A_324_373#_c_1190_n 0.0150383f $X=6.5 $Y=0.745
+ $X2=0 $Y2=0
cc_633 N_A_1057_74#_c_810_n N_A_324_373#_c_1191_n 0.00496574f $X=5.495 $Y=0.515
+ $X2=0 $Y2=0
cc_634 N_A_1057_74#_M1000_d N_A_321_77#_c_1320_n 0.0124053f $X=5.415 $Y=1.99
+ $X2=0 $Y2=0
cc_635 N_A_1057_74#_c_824_n N_A_321_77#_c_1320_n 0.0232623f $X=7.13 $Y=2.99
+ $X2=0 $Y2=0
cc_636 N_A_1057_74#_c_827_n N_A_321_77#_c_1320_n 0.0248462f $X=5.65 $Y=2.895
+ $X2=0 $Y2=0
cc_637 N_A_1057_74#_c_812_n N_A_321_77#_c_1317_n 0.00373319f $X=5.66 $Y=0.34
+ $X2=0 $Y2=0
cc_638 N_A_1057_74#_c_820_n N_X_c_1446_n 0.0103178f $X=8.22 $Y=1.765 $X2=0 $Y2=0
cc_639 N_A_1057_74#_c_821_n N_X_c_1446_n 0.0120855f $X=8.67 $Y=1.765 $X2=0 $Y2=0
cc_640 N_A_1057_74#_c_806_n N_X_c_1443_n 0.0063516f $X=8.295 $Y=1.34 $X2=0 $Y2=0
cc_641 N_A_1057_74#_c_807_n N_X_c_1443_n 0.00605329f $X=8.725 $Y=1.34 $X2=0
+ $Y2=0
cc_642 N_A_1057_74#_c_808_n N_X_c_1443_n 4.95297e-19 $X=9.155 $Y=1.34 $X2=0
+ $Y2=0
cc_643 N_A_1057_74#_c_806_n N_X_c_1444_n 0.00383504f $X=8.295 $Y=1.34 $X2=0
+ $Y2=0
cc_644 N_A_1057_74#_c_807_n N_X_c_1444_n 0.00350884f $X=8.725 $Y=1.34 $X2=0
+ $Y2=0
cc_645 N_A_1057_74#_c_866_p N_X_c_1444_n 0.00606139f $X=8.165 $Y=1.505 $X2=0
+ $Y2=0
cc_646 N_A_1057_74#_c_819_n N_X_c_1444_n 0.00673421f $X=9.57 $Y=1.552 $X2=0
+ $Y2=0
cc_647 N_A_1057_74#_c_819_n N_X_c_1459_n 0.0417832f $X=9.57 $Y=1.552 $X2=0 $Y2=0
cc_648 N_A_1057_74#_c_820_n N_X_c_1447_n 0.00198186f $X=8.22 $Y=1.765 $X2=0
+ $Y2=0
cc_649 N_A_1057_74#_c_821_n N_X_c_1447_n 0.00206972f $X=8.67 $Y=1.765 $X2=0
+ $Y2=0
cc_650 N_A_1057_74#_c_866_p N_X_c_1447_n 0.00126392f $X=8.165 $Y=1.505 $X2=0
+ $Y2=0
cc_651 N_A_1057_74#_c_819_n N_X_c_1447_n 0.00500154f $X=9.57 $Y=1.552 $X2=0
+ $Y2=0
cc_652 N_A_1057_74#_c_820_n N_X_c_1448_n 0.00153296f $X=8.22 $Y=1.765 $X2=0
+ $Y2=0
cc_653 N_A_1057_74#_c_821_n N_X_c_1448_n 0.00178133f $X=8.67 $Y=1.765 $X2=0
+ $Y2=0
cc_654 N_A_1057_74#_c_822_n N_X_c_1448_n 4.94911e-19 $X=9.12 $Y=1.765 $X2=0
+ $Y2=0
cc_655 N_A_1057_74#_c_866_p N_X_c_1448_n 0.00331766f $X=8.165 $Y=1.505 $X2=0
+ $Y2=0
cc_656 N_A_1057_74#_c_819_n N_X_c_1448_n 0.0103003f $X=9.57 $Y=1.552 $X2=0 $Y2=0
cc_657 N_A_1057_74#_c_806_n N_X_c_1469_n 0.00239522f $X=8.295 $Y=1.34 $X2=0
+ $Y2=0
cc_658 N_A_1057_74#_c_807_n N_X_c_1469_n 0.0017052f $X=8.725 $Y=1.34 $X2=0 $Y2=0
cc_659 N_A_1057_74#_c_819_n N_X_c_1469_n 3.01015e-19 $X=9.57 $Y=1.552 $X2=0
+ $Y2=0
cc_660 N_A_1057_74#_c_866_p N_X_c_1472_n 0.0173534f $X=8.165 $Y=1.505 $X2=0
+ $Y2=0
cc_661 N_A_1057_74#_c_819_n N_X_c_1472_n 0.00868505f $X=9.57 $Y=1.552 $X2=0
+ $Y2=0
cc_662 N_A_1057_74#_c_807_n X 5.03719e-19 $X=8.725 $Y=1.34 $X2=0 $Y2=0
cc_663 N_A_1057_74#_c_808_n X 0.0128066f $X=9.155 $Y=1.34 $X2=0 $Y2=0
cc_664 N_A_1057_74#_c_809_n X 0.015578f $X=9.585 $Y=1.34 $X2=0 $Y2=0
cc_665 N_A_1057_74#_c_819_n X 0.0101134f $X=9.57 $Y=1.552 $X2=0 $Y2=0
cc_666 N_A_1057_74#_c_819_n X 0.0173378f $X=9.57 $Y=1.552 $X2=0 $Y2=0
cc_667 N_A_1057_74#_c_821_n X 5.09553e-19 $X=8.67 $Y=1.765 $X2=0 $Y2=0
cc_668 N_A_1057_74#_c_822_n X 0.0146405f $X=9.12 $Y=1.765 $X2=0 $Y2=0
cc_669 N_A_1057_74#_c_823_n X 0.0183129f $X=9.57 $Y=1.765 $X2=0 $Y2=0
cc_670 N_A_1057_74#_c_819_n X 0.0205548f $X=9.57 $Y=1.552 $X2=0 $Y2=0
cc_671 N_A_1057_74#_c_814_n N_VGND_M1017_d 0.00369417f $X=6.89 $Y=0.745 $X2=0
+ $Y2=0
cc_672 N_A_1057_74#_c_932_p N_VGND_M1017_d 0.00687894f $X=6.975 $Y=1.01 $X2=0
+ $Y2=0
cc_673 N_A_1057_74#_c_846_n N_VGND_M1017_d 0.0211435f $X=7.32 $Y=1.095 $X2=0
+ $Y2=0
cc_674 N_A_1057_74#_c_848_n N_VGND_M1017_d 0.00276146f $X=7.06 $Y=1.095 $X2=0
+ $Y2=0
cc_675 N_A_1057_74#_c_816_n N_VGND_M1017_d 0.00260794f $X=7.405 $Y=1.34 $X2=0
+ $Y2=0
cc_676 N_A_1057_74#_c_811_n N_VGND_c_1503_n 0.0546988f $X=6.33 $Y=0.34 $X2=0
+ $Y2=0
cc_677 N_A_1057_74#_c_812_n N_VGND_c_1503_n 0.0236566f $X=5.66 $Y=0.34 $X2=0
+ $Y2=0
cc_678 N_A_1057_74#_c_814_n N_VGND_c_1503_n 0.00691154f $X=6.89 $Y=0.745 $X2=0
+ $Y2=0
cc_679 N_A_1057_74#_c_846_n N_VGND_c_1553_n 0.00671835f $X=7.32 $Y=1.095 $X2=0
+ $Y2=0
cc_680 N_A_1057_74#_c_866_p N_VGND_c_1553_n 0.0203974f $X=8.165 $Y=1.505 $X2=0
+ $Y2=0
cc_681 N_A_1057_74#_c_818_n N_VGND_c_1553_n 0.00584701f $X=8.13 $Y=1.505 $X2=0
+ $Y2=0
cc_682 N_A_1057_74#_c_806_n N_VGND_c_1504_n 0.00473385f $X=8.295 $Y=1.34 $X2=0
+ $Y2=0
cc_683 N_A_1057_74#_c_807_n N_VGND_c_1504_n 0.00473385f $X=8.725 $Y=1.34 $X2=0
+ $Y2=0
cc_684 N_A_1057_74#_c_806_n N_VGND_c_1505_n 0.00558707f $X=8.295 $Y=1.34 $X2=0
+ $Y2=0
cc_685 N_A_1057_74#_c_811_n N_VGND_c_1505_n 0.00877697f $X=6.33 $Y=0.34 $X2=0
+ $Y2=0
cc_686 N_A_1057_74#_c_813_n N_VGND_c_1505_n 0.00301164f $X=6.415 $Y=0.66 $X2=0
+ $Y2=0
cc_687 N_A_1057_74#_c_814_n N_VGND_c_1505_n 0.028714f $X=6.89 $Y=0.745 $X2=0
+ $Y2=0
cc_688 N_A_1057_74#_c_932_p N_VGND_c_1505_n 7.77107e-19 $X=6.975 $Y=1.01 $X2=0
+ $Y2=0
cc_689 N_A_1057_74#_c_846_n N_VGND_c_1505_n 0.0285331f $X=7.32 $Y=1.095 $X2=0
+ $Y2=0
cc_690 N_A_1057_74#_c_866_p N_VGND_c_1505_n 0.0151658f $X=8.165 $Y=1.505 $X2=0
+ $Y2=0
cc_691 N_A_1057_74#_c_818_n N_VGND_c_1505_n 0.00862364f $X=8.13 $Y=1.505 $X2=0
+ $Y2=0
cc_692 N_A_1057_74#_c_807_n N_VGND_c_1506_n 0.0031573f $X=8.725 $Y=1.34 $X2=0
+ $Y2=0
cc_693 N_A_1057_74#_c_808_n N_VGND_c_1506_n 0.00265542f $X=9.155 $Y=1.34 $X2=0
+ $Y2=0
cc_694 N_A_1057_74#_c_819_n N_VGND_c_1506_n 0.00256759f $X=9.57 $Y=1.552 $X2=0
+ $Y2=0
cc_695 N_A_1057_74#_c_809_n N_VGND_c_1508_n 0.00595876f $X=9.585 $Y=1.34 $X2=0
+ $Y2=0
cc_696 N_A_1057_74#_c_808_n N_VGND_c_1510_n 0.00472938f $X=9.155 $Y=1.34 $X2=0
+ $Y2=0
cc_697 N_A_1057_74#_c_809_n N_VGND_c_1510_n 0.00472938f $X=9.585 $Y=1.34 $X2=0
+ $Y2=0
cc_698 N_A_1057_74#_c_806_n N_VGND_c_1514_n 0.00508379f $X=8.295 $Y=1.34 $X2=0
+ $Y2=0
cc_699 N_A_1057_74#_c_807_n N_VGND_c_1514_n 0.00508379f $X=8.725 $Y=1.34 $X2=0
+ $Y2=0
cc_700 N_A_1057_74#_c_808_n N_VGND_c_1514_n 0.00508379f $X=9.155 $Y=1.34 $X2=0
+ $Y2=0
cc_701 N_A_1057_74#_c_809_n N_VGND_c_1514_n 0.00508379f $X=9.585 $Y=1.34 $X2=0
+ $Y2=0
cc_702 N_A_1057_74#_c_811_n N_VGND_c_1514_n 0.0310803f $X=6.33 $Y=0.34 $X2=0
+ $Y2=0
cc_703 N_A_1057_74#_c_812_n N_VGND_c_1514_n 0.0128296f $X=5.66 $Y=0.34 $X2=0
+ $Y2=0
cc_704 N_A_1057_74#_c_814_n N_VGND_c_1514_n 0.0119702f $X=6.89 $Y=0.745 $X2=0
+ $Y2=0
cc_705 N_A_27_373#_c_996_n N_VPWR_c_1078_n 0.00272936f $X=1.535 $Y=2.035 $X2=0
+ $Y2=0
cc_706 N_A_27_373#_c_977_n N_VPWR_c_1078_n 0.0402722f $X=0.28 $Y=2.01 $X2=0
+ $Y2=0
cc_707 N_A_27_373#_c_977_n N_VPWR_c_1086_n 0.00895579f $X=0.28 $Y=2.01 $X2=0
+ $Y2=0
cc_708 N_A_27_373#_c_977_n N_VPWR_c_1077_n 0.0096603f $X=0.28 $Y=2.01 $X2=0
+ $Y2=0
cc_709 N_A_27_373#_c_971_n N_A_324_373#_M1007_d 0.00394167f $X=2.305 $Y=2.65
+ $X2=0 $Y2=0
cc_710 N_A_27_373#_c_1006_n N_A_324_373#_M1007_d 0.00254092f $X=1.68 $Y=2.035
+ $X2=0 $Y2=0
cc_711 N_A_27_373#_c_970_n N_A_324_373#_M1007_d 0.00744138f $X=1.68 $Y=2.035
+ $X2=0 $Y2=0
cc_712 N_A_27_373#_c_1006_n N_A_324_373#_c_1192_n 3.43164e-19 $X=1.68 $Y=2.035
+ $X2=0 $Y2=0
cc_713 N_A_27_373#_c_970_n N_A_324_373#_c_1192_n 0.0222951f $X=1.68 $Y=2.035
+ $X2=0 $Y2=0
cc_714 N_A_27_373#_c_969_n N_A_324_373#_c_1184_n 0.0103721f $X=2.3 $Y=1.1 $X2=0
+ $Y2=0
cc_715 N_A_27_373#_c_975_n N_A_324_373#_c_1184_n 0.00424218f $X=2.47 $Y=2.38
+ $X2=0 $Y2=0
cc_716 N_A_27_373#_c_965_n N_A_324_373#_c_1185_n 0.0158636f $X=2.135 $Y=1.25
+ $X2=0 $Y2=0
cc_717 N_A_27_373#_c_969_n N_A_324_373#_c_1185_n 0.00867013f $X=2.3 $Y=1.1 $X2=0
+ $Y2=0
cc_718 N_A_27_373#_c_970_n N_A_324_373#_c_1185_n 0.0145177f $X=1.68 $Y=2.035
+ $X2=0 $Y2=0
cc_719 N_A_27_373#_c_969_n N_A_324_373#_c_1186_n 0.0096475f $X=2.3 $Y=1.1 $X2=0
+ $Y2=0
cc_720 N_A_27_373#_c_969_n N_A_324_373#_c_1210_n 0.0194434f $X=2.3 $Y=1.1 $X2=0
+ $Y2=0
cc_721 N_A_27_373#_M1019_d N_A_324_373#_c_1195_n 0.00558234f $X=2.32 $Y=1.865
+ $X2=0 $Y2=0
cc_722 N_A_27_373#_c_975_n N_A_324_373#_c_1195_n 0.012913f $X=2.47 $Y=2.38 $X2=0
+ $Y2=0
cc_723 N_A_27_373#_c_965_n N_A_324_373#_c_1219_n 3.65365e-19 $X=2.135 $Y=1.25
+ $X2=0 $Y2=0
cc_724 N_A_27_373#_c_971_n N_A_324_373#_c_1219_n 0.00486f $X=2.305 $Y=2.65 $X2=0
+ $Y2=0
cc_725 N_A_27_373#_c_969_n N_A_324_373#_c_1219_n 4.49084e-19 $X=2.3 $Y=1.1 $X2=0
+ $Y2=0
cc_726 N_A_27_373#_c_1006_n N_A_324_373#_c_1219_n 0.0210157f $X=1.68 $Y=2.035
+ $X2=0 $Y2=0
cc_727 N_A_27_373#_c_970_n N_A_324_373#_c_1219_n 2.03155e-19 $X=1.68 $Y=2.035
+ $X2=0 $Y2=0
cc_728 N_A_27_373#_c_971_n N_A_324_373#_c_1220_n 0.00936303f $X=2.305 $Y=2.65
+ $X2=0 $Y2=0
cc_729 N_A_27_373#_c_1006_n N_A_324_373#_c_1220_n 0.00151832f $X=1.68 $Y=2.035
+ $X2=0 $Y2=0
cc_730 N_A_27_373#_c_970_n N_A_324_373#_c_1220_n 0.0126015f $X=1.68 $Y=2.035
+ $X2=0 $Y2=0
cc_731 N_A_27_373#_c_975_n N_A_321_77#_c_1339_n 0.00615406f $X=2.47 $Y=2.38
+ $X2=0 $Y2=0
cc_732 N_A_27_373#_c_975_n N_A_321_77#_c_1329_n 0.0146685f $X=2.47 $Y=2.38 $X2=0
+ $Y2=0
cc_733 N_A_27_373#_c_965_n N_A_321_77#_c_1314_n 0.0124306f $X=2.135 $Y=1.25
+ $X2=0 $Y2=0
cc_734 N_A_27_373#_c_968_n N_A_321_77#_c_1314_n 0.0108039f $X=1.665 $Y=1.475
+ $X2=0 $Y2=0
cc_735 N_A_27_373#_M1006_d N_A_321_77#_c_1315_n 0.00731496f $X=2.08 $Y=0.605
+ $X2=0 $Y2=0
cc_736 N_A_27_373#_c_965_n N_A_321_77#_c_1315_n 0.00539878f $X=2.135 $Y=1.25
+ $X2=0 $Y2=0
cc_737 N_A_27_373#_c_969_n N_A_321_77#_c_1315_n 0.0192566f $X=2.3 $Y=1.1 $X2=0
+ $Y2=0
cc_738 N_A_27_373#_c_966_n N_VGND_c_1501_n 0.0201853f $X=0.33 $Y=0.615 $X2=0
+ $Y2=0
cc_739 N_A_27_373#_c_966_n N_VGND_c_1511_n 0.016911f $X=0.33 $Y=0.615 $X2=0
+ $Y2=0
cc_740 N_A_27_373#_c_966_n N_VGND_c_1514_n 0.0148316f $X=0.33 $Y=0.615 $X2=0
+ $Y2=0
cc_741 N_VPWR_M1022_d N_A_324_373#_c_1195_n 0.00553803f $X=4.405 $Y=1.84 $X2=0
+ $Y2=0
cc_742 N_VPWR_c_1079_n N_A_321_77#_c_1318_n 9.02477e-19 $X=4.555 $Y=2.815 $X2=0
+ $Y2=0
cc_743 N_VPWR_c_1077_n N_A_321_77#_c_1318_n 0.0246512f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_744 N_VPWR_M1022_d N_A_321_77#_c_1313_n 0.00866885f $X=4.405 $Y=1.84 $X2=0
+ $Y2=0
cc_745 N_VPWR_M1022_d N_A_321_77#_c_1320_n 0.00305933f $X=4.405 $Y=1.84 $X2=0
+ $Y2=0
cc_746 N_VPWR_c_1079_n N_A_321_77#_c_1320_n 0.0086438f $X=4.555 $Y=2.815 $X2=0
+ $Y2=0
cc_747 N_VPWR_c_1077_n N_A_321_77#_c_1320_n 0.0291527f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_748 N_VPWR_M1022_d N_A_321_77#_c_1387_n 0.00227128f $X=4.405 $Y=1.84 $X2=0
+ $Y2=0
cc_749 N_VPWR_c_1079_n N_A_321_77#_c_1387_n 0.01289f $X=4.555 $Y=2.815 $X2=0
+ $Y2=0
cc_750 N_VPWR_c_1077_n N_A_321_77#_c_1387_n 6.84279e-19 $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_751 N_VPWR_c_1082_n N_X_c_1446_n 0.0158009f $X=8.81 $Y=3.33 $X2=0 $Y2=0
cc_752 N_VPWR_c_1077_n N_X_c_1446_n 0.0129424f $X=9.84 $Y=3.33 $X2=0 $Y2=0
cc_753 N_VPWR_c_1083_n N_X_c_1459_n 0.0123804f $X=8.895 $Y=1.985 $X2=0 $Y2=0
cc_754 N_VPWR_c_1080_n N_X_c_1447_n 0.0441815f $X=7.797 $Y=3.245 $X2=0 $Y2=0
cc_755 N_VPWR_c_1083_n N_X_c_1448_n 0.0861314f $X=8.895 $Y=1.985 $X2=0 $Y2=0
cc_756 N_VPWR_c_1083_n X 0.076043f $X=8.895 $Y=1.985 $X2=0 $Y2=0
cc_757 N_VPWR_c_1085_n X 0.0867368f $X=9.795 $Y=1.985 $X2=0 $Y2=0
cc_758 N_VPWR_c_1089_n X 0.0155928f $X=9.71 $Y=3.33 $X2=0 $Y2=0
cc_759 N_VPWR_c_1077_n X 0.0127818f $X=9.84 $Y=3.33 $X2=0 $Y2=0
cc_760 N_VPWR_c_1085_n N_VGND_c_1508_n 0.00977564f $X=9.795 $Y=1.985 $X2=0 $Y2=0
cc_761 N_A_324_373#_c_1195_n N_A_321_77#_M1020_d 0.00894192f $X=4.895 $Y=2.035
+ $X2=0 $Y2=0
cc_762 N_A_324_373#_M1004_d N_A_321_77#_c_1312_n 0.00368186f $X=2.695 $Y=0.605
+ $X2=0 $Y2=0
cc_763 N_A_324_373#_c_1192_n N_A_321_77#_c_1339_n 0.00170998f $X=2.09 $Y=1.965
+ $X2=0 $Y2=0
cc_764 N_A_324_373#_c_1210_n N_A_321_77#_c_1339_n 0.00214892f $X=2.845 $Y=1.04
+ $X2=0 $Y2=0
cc_765 N_A_324_373#_c_1195_n N_A_321_77#_c_1339_n 0.0281991f $X=4.895 $Y=2.035
+ $X2=0 $Y2=0
cc_766 N_A_324_373#_c_1219_n N_A_321_77#_c_1339_n 0.0020436f $X=2.305 $Y=2.035
+ $X2=0 $Y2=0
cc_767 N_A_324_373#_c_1220_n N_A_321_77#_c_1339_n 0.00169507f $X=2.02 $Y=1.99
+ $X2=0 $Y2=0
cc_768 N_A_324_373#_c_1195_n N_A_321_77#_c_1318_n 0.0222067f $X=4.895 $Y=2.035
+ $X2=0 $Y2=0
cc_769 N_A_324_373#_c_1187_n N_A_321_77#_c_1313_n 0.0425792f $X=4.865 $Y=1.95
+ $X2=0 $Y2=0
cc_770 N_A_324_373#_c_1188_n N_A_321_77#_c_1313_n 0.014358f $X=4.95 $Y=1.295
+ $X2=0 $Y2=0
cc_771 N_A_324_373#_c_1195_n N_A_321_77#_c_1313_n 0.0225247f $X=4.895 $Y=2.035
+ $X2=0 $Y2=0
cc_772 N_A_324_373#_c_1196_n N_A_321_77#_c_1313_n 5.02359e-19 $X=5.04 $Y=2.035
+ $X2=0 $Y2=0
cc_773 N_A_324_373#_c_1197_n N_A_321_77#_c_1313_n 0.0200577f $X=5.04 $Y=2.035
+ $X2=0 $Y2=0
cc_774 N_A_324_373#_M1000_s N_A_321_77#_c_1320_n 0.00784776f $X=4.97 $Y=1.99
+ $X2=0 $Y2=0
cc_775 N_A_324_373#_c_1195_n N_A_321_77#_c_1320_n 0.00753536f $X=4.895 $Y=2.035
+ $X2=0 $Y2=0
cc_776 N_A_324_373#_c_1196_n N_A_321_77#_c_1320_n 0.00183698f $X=5.04 $Y=2.035
+ $X2=0 $Y2=0
cc_777 N_A_324_373#_c_1197_n N_A_321_77#_c_1320_n 0.0313734f $X=5.04 $Y=2.035
+ $X2=0 $Y2=0
cc_778 N_A_324_373#_c_1210_n N_A_321_77#_c_1316_n 0.0254466f $X=2.845 $Y=1.04
+ $X2=0 $Y2=0
cc_779 N_A_324_373#_c_1188_n N_A_321_77#_c_1317_n 0.015131f $X=4.95 $Y=1.295
+ $X2=0 $Y2=0
cc_780 N_A_324_373#_c_1190_n N_A_321_77#_c_1317_n 5.07708e-19 $X=5.995 $Y=0.81
+ $X2=0 $Y2=0
cc_781 N_A_324_373#_c_1191_n N_A_321_77#_c_1317_n 0.0167867f $X=5.405 $Y=1.28
+ $X2=0 $Y2=0
cc_782 N_A_321_77#_c_1312_n N_VGND_M1021_d 0.00524428f $X=4.44 $Y=0.7 $X2=0
+ $Y2=0
cc_783 N_A_321_77#_c_1313_n N_VGND_M1021_d 0.00315635f $X=4.525 $Y=2.37 $X2=0
+ $Y2=0
cc_784 N_A_321_77#_c_1317_n N_VGND_M1021_d 0.00804534f $X=4.525 $Y=0.69 $X2=0
+ $Y2=0
cc_785 N_A_321_77#_c_1312_n N_VGND_c_1502_n 0.0127357f $X=4.44 $Y=0.7 $X2=0
+ $Y2=0
cc_786 N_A_321_77#_c_1317_n N_VGND_c_1502_n 0.0197889f $X=4.525 $Y=0.69 $X2=0
+ $Y2=0
cc_787 N_A_321_77#_c_1317_n N_VGND_c_1503_n 0.019328f $X=4.525 $Y=0.69 $X2=0
+ $Y2=0
cc_788 N_A_321_77#_c_1312_n N_VGND_c_1509_n 0.0126356f $X=4.44 $Y=0.7 $X2=0
+ $Y2=0
cc_789 N_A_321_77#_c_1312_n N_VGND_c_1514_n 0.0238176f $X=4.44 $Y=0.7 $X2=0
+ $Y2=0
cc_790 N_A_321_77#_c_1317_n N_VGND_c_1514_n 0.0198891f $X=4.525 $Y=0.69 $X2=0
+ $Y2=0
cc_791 N_X_c_1443_n N_VGND_c_1504_n 0.00971834f $X=8.51 $Y=0.635 $X2=0 $Y2=0
cc_792 N_X_c_1443_n N_VGND_c_1505_n 0.0141711f $X=8.51 $Y=0.635 $X2=0 $Y2=0
cc_793 N_X_c_1443_n N_VGND_c_1506_n 0.0290583f $X=8.51 $Y=0.635 $X2=0 $Y2=0
cc_794 N_X_c_1459_n N_VGND_c_1506_n 0.0137224f $X=9.18 $Y=1.522 $X2=0 $Y2=0
cc_795 X N_VGND_c_1506_n 0.0314886f $X=9.275 $Y=0.47 $X2=0 $Y2=0
cc_796 X N_VGND_c_1508_n 0.0316368f $X=9.275 $Y=0.47 $X2=0 $Y2=0
cc_797 X N_VGND_c_1510_n 0.0105983f $X=9.275 $Y=0.47 $X2=0 $Y2=0
cc_798 N_X_c_1443_n N_VGND_c_1514_n 0.0111609f $X=8.51 $Y=0.635 $X2=0 $Y2=0
cc_799 X N_VGND_c_1514_n 0.0113894f $X=9.275 $Y=0.47 $X2=0 $Y2=0
