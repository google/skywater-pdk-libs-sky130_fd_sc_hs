* File: sky130_fd_sc_hs__dlrbn_1.pxi.spice
* Created: Tue Sep  1 20:01:39 2020
* 
x_PM_SKY130_FD_SC_HS__DLRBN_1%D N_D_c_155_n N_D_M1009_g N_D_c_160_n N_D_M1019_g
+ D N_D_c_158_n PM_SKY130_FD_SC_HS__DLRBN_1%D
x_PM_SKY130_FD_SC_HS__DLRBN_1%GATE_N N_GATE_N_M1003_g N_GATE_N_c_189_n
+ N_GATE_N_c_193_n N_GATE_N_M1015_g GATE_N N_GATE_N_c_190_n N_GATE_N_c_191_n
+ PM_SKY130_FD_SC_HS__DLRBN_1%GATE_N
x_PM_SKY130_FD_SC_HS__DLRBN_1%A_231_74# N_A_231_74#_M1003_d N_A_231_74#_M1015_d
+ N_A_231_74#_M1013_g N_A_231_74#_c_223_n N_A_231_74#_c_235_n
+ N_A_231_74#_M1005_g N_A_231_74#_M1002_g N_A_231_74#_c_236_n
+ N_A_231_74#_M1021_g N_A_231_74#_c_237_n N_A_231_74#_c_238_n
+ N_A_231_74#_c_224_n N_A_231_74#_c_266_p N_A_231_74#_c_225_n
+ N_A_231_74#_c_240_n N_A_231_74#_c_241_n N_A_231_74#_c_242_n
+ N_A_231_74#_c_226_n N_A_231_74#_c_243_n N_A_231_74#_c_227_n
+ N_A_231_74#_c_228_n N_A_231_74#_c_229_n N_A_231_74#_c_271_p
+ N_A_231_74#_c_230_n N_A_231_74#_c_231_n N_A_231_74#_c_232_n
+ N_A_231_74#_c_233_n N_A_231_74#_c_245_n PM_SKY130_FD_SC_HS__DLRBN_1%A_231_74#
x_PM_SKY130_FD_SC_HS__DLRBN_1%A_27_424# N_A_27_424#_M1009_s N_A_27_424#_M1019_s
+ N_A_27_424#_M1001_g N_A_27_424#_c_384_n N_A_27_424#_M1008_g
+ N_A_27_424#_c_385_n N_A_27_424#_c_386_n N_A_27_424#_c_391_n
+ N_A_27_424#_c_392_n N_A_27_424#_c_405_n N_A_27_424#_c_393_n
+ N_A_27_424#_c_413_n N_A_27_424#_c_439_n N_A_27_424#_c_394_n
+ N_A_27_424#_c_387_n N_A_27_424#_c_395_n N_A_27_424#_c_396_n
+ N_A_27_424#_c_388_n PM_SKY130_FD_SC_HS__DLRBN_1%A_27_424#
x_PM_SKY130_FD_SC_HS__DLRBN_1%A_373_74# N_A_373_74#_M1013_s N_A_373_74#_M1005_s
+ N_A_373_74#_c_498_n N_A_373_74#_M1012_g N_A_373_74#_c_499_n
+ N_A_373_74#_c_500_n N_A_373_74#_c_491_n N_A_373_74#_M1011_g
+ N_A_373_74#_c_492_n N_A_373_74#_c_493_n N_A_373_74#_c_525_n
+ N_A_373_74#_c_494_n N_A_373_74#_c_495_n N_A_373_74#_c_496_n
+ N_A_373_74#_c_503_n N_A_373_74#_c_497_n PM_SKY130_FD_SC_HS__DLRBN_1%A_373_74#
x_PM_SKY130_FD_SC_HS__DLRBN_1%A_889_92# N_A_889_92#_M1014_s N_A_889_92#_M1017_d
+ N_A_889_92#_M1022_g N_A_889_92#_c_601_n N_A_889_92#_M1016_g
+ N_A_889_92#_c_591_n N_A_889_92#_M1018_g N_A_889_92#_c_602_n
+ N_A_889_92#_M1004_g N_A_889_92#_c_592_n N_A_889_92#_M1000_g
+ N_A_889_92#_c_593_n N_A_889_92#_M1010_g N_A_889_92#_c_594_n
+ N_A_889_92#_c_595_n N_A_889_92#_c_596_n N_A_889_92#_c_597_n
+ N_A_889_92#_c_607_n N_A_889_92#_c_651_p N_A_889_92#_c_608_n
+ N_A_889_92#_c_598_n N_A_889_92#_c_609_n N_A_889_92#_c_624_p
+ N_A_889_92#_c_599_n PM_SKY130_FD_SC_HS__DLRBN_1%A_889_92#
x_PM_SKY130_FD_SC_HS__DLRBN_1%A_686_74# N_A_686_74#_M1002_d N_A_686_74#_M1012_d
+ N_A_686_74#_c_718_n N_A_686_74#_M1017_g N_A_686_74#_c_719_n
+ N_A_686_74#_M1014_g N_A_686_74#_c_720_n N_A_686_74#_c_721_n
+ N_A_686_74#_c_727_n N_A_686_74#_c_728_n N_A_686_74#_c_722_n
+ N_A_686_74#_c_729_n N_A_686_74#_c_730_n N_A_686_74#_c_723_n
+ N_A_686_74#_c_724_n PM_SKY130_FD_SC_HS__DLRBN_1%A_686_74#
x_PM_SKY130_FD_SC_HS__DLRBN_1%RESET_B N_RESET_B_c_811_n N_RESET_B_M1006_g
+ N_RESET_B_c_812_n N_RESET_B_M1007_g RESET_B
+ PM_SKY130_FD_SC_HS__DLRBN_1%RESET_B
x_PM_SKY130_FD_SC_HS__DLRBN_1%A_1437_112# N_A_1437_112#_M1010_s
+ N_A_1437_112#_M1000_s N_A_1437_112#_M1020_g N_A_1437_112#_c_843_n
+ N_A_1437_112#_M1023_g N_A_1437_112#_c_844_n N_A_1437_112#_c_847_n
+ N_A_1437_112#_c_845_n N_A_1437_112#_c_855_n
+ PM_SKY130_FD_SC_HS__DLRBN_1%A_1437_112#
x_PM_SKY130_FD_SC_HS__DLRBN_1%VPWR N_VPWR_M1019_d N_VPWR_M1005_d N_VPWR_M1016_d
+ N_VPWR_M1007_d N_VPWR_M1000_d N_VPWR_c_881_n N_VPWR_c_882_n N_VPWR_c_883_n
+ N_VPWR_c_884_n N_VPWR_c_885_n N_VPWR_c_886_n VPWR N_VPWR_c_887_n
+ N_VPWR_c_888_n N_VPWR_c_889_n N_VPWR_c_890_n N_VPWR_c_891_n N_VPWR_c_880_n
+ N_VPWR_c_893_n N_VPWR_c_894_n N_VPWR_c_895_n N_VPWR_c_896_n
+ PM_SKY130_FD_SC_HS__DLRBN_1%VPWR
x_PM_SKY130_FD_SC_HS__DLRBN_1%Q N_Q_M1018_d N_Q_M1004_d N_Q_c_991_n N_Q_c_989_n
+ Q Q Q Q N_Q_c_990_n PM_SKY130_FD_SC_HS__DLRBN_1%Q
x_PM_SKY130_FD_SC_HS__DLRBN_1%Q_N N_Q_N_M1020_d N_Q_N_M1023_d N_Q_N_c_1022_n
+ N_Q_N_c_1023_n Q_N Q_N Q_N Q_N N_Q_N_c_1024_n PM_SKY130_FD_SC_HS__DLRBN_1%Q_N
x_PM_SKY130_FD_SC_HS__DLRBN_1%VGND N_VGND_M1009_d N_VGND_M1013_d N_VGND_M1022_d
+ N_VGND_M1006_d N_VGND_M1010_d N_VGND_c_1040_n N_VGND_c_1041_n N_VGND_c_1042_n
+ N_VGND_c_1043_n N_VGND_c_1044_n N_VGND_c_1045_n N_VGND_c_1046_n
+ N_VGND_c_1047_n VGND N_VGND_c_1048_n N_VGND_c_1049_n N_VGND_c_1050_n
+ N_VGND_c_1051_n N_VGND_c_1052_n N_VGND_c_1053_n N_VGND_c_1054_n
+ N_VGND_c_1055_n PM_SKY130_FD_SC_HS__DLRBN_1%VGND
cc_1 VNB N_D_c_155_n 0.016305f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.755
cc_2 VNB N_D_M1009_g 0.0253435f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=0.835
cc_3 VNB D 0.00308426f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_4 VNB N_D_c_158_n 0.0195483f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=1.425
cc_5 VNB N_GATE_N_M1003_g 0.0254204f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=1.26
cc_6 VNB N_GATE_N_c_189_n 0.0177003f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_7 VNB N_GATE_N_c_190_n 0.0194684f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=1.425
cc_8 VNB N_GATE_N_c_191_n 0.00167584f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=1.425
cc_9 VNB N_A_231_74#_c_223_n 5.11773e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_231_74#_c_224_n 0.0174423f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_231_74#_c_225_n 0.00208626f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_231_74#_c_226_n 0.0188951f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_231_74#_c_227_n 0.0104397f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_231_74#_c_228_n 0.0064596f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_231_74#_c_229_n 0.0370968f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_231_74#_c_230_n 0.00340824f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_231_74#_c_231_n 0.0320407f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_231_74#_c_232_n 0.0230031f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_231_74#_c_233_n 0.0221259f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_27_424#_M1001_g 0.0371673f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.54
cc_21 VNB N_A_27_424#_c_384_n 0.0120422f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_27_424#_c_385_n 0.0184896f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=1.425
cc_23 VNB N_A_27_424#_c_386_n 0.0265823f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.58
cc_24 VNB N_A_27_424#_c_387_n 0.00694384f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_27_424#_c_388_n 0.00166816f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_373_74#_c_491_n 0.00724087f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=1.425
cc_27 VNB N_A_373_74#_c_492_n 0.00635466f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_373_74#_c_493_n 0.00994104f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_373_74#_c_494_n 0.00282738f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_373_74#_c_495_n 0.0327142f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_373_74#_c_496_n 0.00156078f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_373_74#_c_497_n 0.0168064f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_889_92#_M1022_g 0.0372568f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.54
cc_34 VNB N_A_889_92#_c_591_n 0.0227136f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=1.425
cc_35 VNB N_A_889_92#_c_592_n 0.0323972f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_889_92#_c_593_n 0.0200296f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_889_92#_c_594_n 0.00949791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_889_92#_c_595_n 0.0509359f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_889_92#_c_596_n 0.00790367f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_889_92#_c_597_n 0.00260448f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_889_92#_c_598_n 0.0014379f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_889_92#_c_599_n 0.0051572f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_686_74#_c_718_n 0.0157995f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.045
cc_44 VNB N_A_686_74#_c_719_n 0.0190214f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_45 VNB N_A_686_74#_c_720_n 0.0514805f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=1.425
cc_46 VNB N_A_686_74#_c_721_n 0.0106362f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.26
cc_47 VNB N_A_686_74#_c_722_n 0.00299392f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_686_74#_c_723_n 0.00867816f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A_686_74#_c_724_n 0.00125564f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_RESET_B_c_811_n 0.0172017f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.435
cc_51 VNB N_RESET_B_c_812_n 0.0267414f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=0.835
cc_52 VNB RESET_B 0.00303071f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.045
cc_53 VNB N_A_1437_112#_M1020_g 0.028717f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.54
cc_54 VNB N_A_1437_112#_c_843_n 0.0343466f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_A_1437_112#_c_844_n 0.00396499f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=1.58
cc_56 VNB N_A_1437_112#_c_845_n 0.00736448f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_VPWR_c_880_n 0.362705f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_Q_c_989_n 0.00298795f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.425
cc_59 VNB N_Q_c_990_n 0.0172723f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_Q_N_c_1022_n 0.0270633f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.54
cc_61 VNB N_Q_N_c_1023_n 0.0103149f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=1.425
cc_62 VNB N_Q_N_c_1024_n 0.0249555f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_VGND_c_1040_n 0.0168478f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.58
cc_64 VNB N_VGND_c_1041_n 0.0241173f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_VGND_c_1042_n 0.00650089f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_VGND_c_1043_n 0.014346f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_VGND_c_1044_n 0.0488481f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_VGND_c_1045_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_VGND_c_1046_n 0.0312541f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_VGND_c_1047_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_VGND_c_1048_n 0.0202939f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_VGND_c_1049_n 0.0372375f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_VGND_c_1050_n 0.0382617f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_VGND_c_1051_n 0.0177539f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_VGND_c_1052_n 0.501058f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_VGND_c_1053_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_VGND_c_1054_n 0.0198288f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_VGND_c_1055_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VPB N_D_c_155_n 0.0336057f $X=-0.19 $Y=1.66 $X2=0.59 $Y2=1.755
cc_80 VPB N_D_c_160_n 0.0210174f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.045
cc_81 VPB D 0.00211207f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_82 VPB N_GATE_N_c_189_n 0.0346399f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_83 VPB N_GATE_N_c_193_n 0.0215124f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.045
cc_84 VPB N_A_231_74#_c_223_n 0.0131119f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_85 VPB N_A_231_74#_c_235_n 0.0238423f $X=-0.19 $Y=1.66 $X2=0.59 $Y2=1.425
cc_86 VPB N_A_231_74#_c_236_n 0.0165629f $X=-0.19 $Y=1.66 $X2=0.72 $Y2=1.58
cc_87 VPB N_A_231_74#_c_237_n 0.0107577f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_88 VPB N_A_231_74#_c_238_n 0.00257062f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_89 VPB N_A_231_74#_c_225_n 0.00404331f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_90 VPB N_A_231_74#_c_240_n 0.00654345f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_91 VPB N_A_231_74#_c_241_n 0.00215416f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_92 VPB N_A_231_74#_c_242_n 0.00470036f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_93 VPB N_A_231_74#_c_243_n 0.00989579f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_94 VPB N_A_231_74#_c_227_n 0.0107174f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_95 VPB N_A_231_74#_c_245_n 0.0515704f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_96 VPB N_A_27_424#_c_384_n 0.0448413f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_97 VPB N_A_27_424#_c_386_n 0.0193028f $X=-0.19 $Y=1.66 $X2=0.72 $Y2=1.58
cc_98 VPB N_A_27_424#_c_391_n 0.0305297f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_99 VPB N_A_27_424#_c_392_n 0.0108668f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_100 VPB N_A_27_424#_c_393_n 0.00609515f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_101 VPB N_A_27_424#_c_394_n 0.00104736f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_102 VPB N_A_27_424#_c_395_n 0.0114606f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_103 VPB N_A_27_424#_c_396_n 0.00651473f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_104 VPB N_A_373_74#_c_498_n 0.0149057f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.045
cc_105 VPB N_A_373_74#_c_499_n 0.0356235f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_106 VPB N_A_373_74#_c_500_n 0.0101843f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_107 VPB N_A_373_74#_c_491_n 0.00831806f $X=-0.19 $Y=1.66 $X2=0.6 $Y2=1.425
cc_108 VPB N_A_373_74#_c_493_n 0.00388309f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_109 VPB N_A_373_74#_c_503_n 0.0113467f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_110 VPB N_A_889_92#_M1022_g 0.00809253f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.54
cc_111 VPB N_A_889_92#_c_601_n 0.0993444f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_112 VPB N_A_889_92#_c_602_n 0.019376f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_113 VPB N_A_889_92#_c_592_n 0.0421727f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_114 VPB N_A_889_92#_c_594_n 0.00641303f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_115 VPB N_A_889_92#_c_595_n 0.0159011f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_116 VPB N_A_889_92#_c_597_n 0.00263986f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_117 VPB N_A_889_92#_c_607_n 0.00328008f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_118 VPB N_A_889_92#_c_608_n 0.00191836f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_119 VPB N_A_889_92#_c_609_n 0.0144596f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_120 VPB N_A_889_92#_c_599_n 3.8003e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_121 VPB N_A_686_74#_c_718_n 0.0228889f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.045
cc_122 VPB N_A_686_74#_c_720_n 0.0131665f $X=-0.19 $Y=1.66 $X2=0.6 $Y2=1.425
cc_123 VPB N_A_686_74#_c_727_n 0.0138866f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_124 VPB N_A_686_74#_c_728_n 0.00347407f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_125 VPB N_A_686_74#_c_729_n 8.46624e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_126 VPB N_A_686_74#_c_730_n 0.0101313f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_127 VPB N_A_686_74#_c_723_n 0.00776532f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_128 VPB N_RESET_B_c_812_n 0.0273801f $X=-0.19 $Y=1.66 $X2=0.5 $Y2=0.835
cc_129 VPB RESET_B 0.00114307f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.045
cc_130 VPB N_A_1437_112#_c_843_n 0.0292273f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_131 VPB N_A_1437_112#_c_847_n 0.00420072f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_132 VPB N_VPWR_c_881_n 0.00687615f $X=-0.19 $Y=1.66 $X2=0.72 $Y2=1.58
cc_133 VPB N_VPWR_c_882_n 0.0128946f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_134 VPB N_VPWR_c_883_n 0.0173003f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_135 VPB N_VPWR_c_884_n 0.0197353f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_136 VPB N_VPWR_c_885_n 0.0192774f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_137 VPB N_VPWR_c_886_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_138 VPB N_VPWR_c_887_n 0.0178711f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_139 VPB N_VPWR_c_888_n 0.0424939f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_140 VPB N_VPWR_c_889_n 0.0468561f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_141 VPB N_VPWR_c_890_n 0.0374389f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_142 VPB N_VPWR_c_891_n 0.0195898f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_143 VPB N_VPWR_c_880_n 0.129666f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_144 VPB N_VPWR_c_893_n 0.00614127f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_145 VPB N_VPWR_c_894_n 0.00631222f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_146 VPB N_VPWR_c_895_n 0.0342281f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_147 VPB N_VPWR_c_896_n 0.00507132f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_148 VPB N_Q_c_991_n 0.00313558f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_149 VPB N_Q_c_989_n 0.00117511f $X=-0.19 $Y=1.66 $X2=0.59 $Y2=1.425
cc_150 VPB Q 0.0187021f $X=-0.19 $Y=1.66 $X2=0.59 $Y2=1.26
cc_151 VPB Q_N 0.0121283f $X=-0.19 $Y=1.66 $X2=0.6 $Y2=1.425
cc_152 VPB Q_N 0.0407407f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_153 VPB N_Q_N_c_1024_n 0.00762538f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_154 N_D_M1009_g N_GATE_N_M1003_g 0.0178869f $X=0.5 $Y=0.835 $X2=0 $Y2=0
cc_155 N_D_c_155_n N_GATE_N_c_189_n 0.0209699f $X=0.59 $Y=1.755 $X2=0 $Y2=0
cc_156 N_D_c_160_n N_GATE_N_c_193_n 0.00955736f $X=0.505 $Y=2.045 $X2=0 $Y2=0
cc_157 D N_GATE_N_c_190_n 0.0039472f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_158 N_D_c_158_n N_GATE_N_c_190_n 0.0178913f $X=0.6 $Y=1.425 $X2=0 $Y2=0
cc_159 D N_GATE_N_c_191_n 0.0514478f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_160 N_D_c_158_n N_GATE_N_c_191_n 7.01786e-19 $X=0.6 $Y=1.425 $X2=0 $Y2=0
cc_161 N_D_M1009_g N_A_27_424#_c_385_n 0.00592841f $X=0.5 $Y=0.835 $X2=0 $Y2=0
cc_162 N_D_M1009_g N_A_27_424#_c_386_n 0.00413599f $X=0.5 $Y=0.835 $X2=0 $Y2=0
cc_163 D N_A_27_424#_c_386_n 0.0488225f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_164 N_D_c_158_n N_A_27_424#_c_386_n 0.0192244f $X=0.6 $Y=1.425 $X2=0 $Y2=0
cc_165 N_D_c_160_n N_A_27_424#_c_391_n 0.00906535f $X=0.505 $Y=2.045 $X2=0 $Y2=0
cc_166 N_D_c_155_n N_A_27_424#_c_392_n 0.00576977f $X=0.59 $Y=1.755 $X2=0 $Y2=0
cc_167 N_D_c_160_n N_A_27_424#_c_392_n 0.014991f $X=0.505 $Y=2.045 $X2=0 $Y2=0
cc_168 D N_A_27_424#_c_392_n 0.031434f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_169 N_D_c_160_n N_A_27_424#_c_405_n 0.00232873f $X=0.505 $Y=2.045 $X2=0 $Y2=0
cc_170 N_D_M1009_g N_A_27_424#_c_387_n 0.00423024f $X=0.5 $Y=0.835 $X2=0 $Y2=0
cc_171 D N_A_27_424#_c_387_n 0.00115505f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_172 N_D_c_160_n N_VPWR_c_881_n 0.0132659f $X=0.505 $Y=2.045 $X2=0 $Y2=0
cc_173 N_D_c_160_n N_VPWR_c_887_n 0.00413917f $X=0.505 $Y=2.045 $X2=0 $Y2=0
cc_174 N_D_c_160_n N_VPWR_c_880_n 0.00821221f $X=0.505 $Y=2.045 $X2=0 $Y2=0
cc_175 N_D_M1009_g N_VGND_c_1040_n 0.00658895f $X=0.5 $Y=0.835 $X2=0 $Y2=0
cc_176 D N_VGND_c_1040_n 0.0179355f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_177 N_D_c_158_n N_VGND_c_1040_n 0.0035943f $X=0.6 $Y=1.425 $X2=0 $Y2=0
cc_178 N_D_M1009_g N_VGND_c_1048_n 0.0043356f $X=0.5 $Y=0.835 $X2=0 $Y2=0
cc_179 N_D_M1009_g N_VGND_c_1052_n 0.00487769f $X=0.5 $Y=0.835 $X2=0 $Y2=0
cc_180 N_GATE_N_M1003_g N_A_231_74#_c_226_n 0.00912459f $X=1.08 $Y=0.74 $X2=0
+ $Y2=0
cc_181 N_GATE_N_c_190_n N_A_231_74#_c_226_n 0.00224336f $X=1.17 $Y=1.425 $X2=0
+ $Y2=0
cc_182 N_GATE_N_c_191_n N_A_231_74#_c_226_n 0.0149863f $X=1.17 $Y=1.425 $X2=0
+ $Y2=0
cc_183 N_GATE_N_c_193_n N_A_231_74#_c_243_n 0.00271601f $X=1.265 $Y=2.045 $X2=0
+ $Y2=0
cc_184 N_GATE_N_M1003_g N_A_231_74#_c_227_n 0.0044988f $X=1.08 $Y=0.74 $X2=0
+ $Y2=0
cc_185 N_GATE_N_c_193_n N_A_231_74#_c_227_n 0.0014507f $X=1.265 $Y=2.045 $X2=0
+ $Y2=0
cc_186 N_GATE_N_c_190_n N_A_231_74#_c_227_n 0.0200944f $X=1.17 $Y=1.425 $X2=0
+ $Y2=0
cc_187 N_GATE_N_c_191_n N_A_231_74#_c_227_n 0.0480239f $X=1.17 $Y=1.425 $X2=0
+ $Y2=0
cc_188 N_GATE_N_c_189_n N_A_27_424#_c_392_n 0.0052319f $X=1.18 $Y=1.755 $X2=0
+ $Y2=0
cc_189 N_GATE_N_c_193_n N_A_27_424#_c_392_n 0.00610303f $X=1.265 $Y=2.045 $X2=0
+ $Y2=0
cc_190 N_GATE_N_c_191_n N_A_27_424#_c_392_n 0.0195412f $X=1.17 $Y=1.425 $X2=0
+ $Y2=0
cc_191 N_GATE_N_c_193_n N_A_27_424#_c_405_n 0.013736f $X=1.265 $Y=2.045 $X2=0
+ $Y2=0
cc_192 N_GATE_N_c_193_n N_A_27_424#_c_393_n 0.0114517f $X=1.265 $Y=2.045 $X2=0
+ $Y2=0
cc_193 N_GATE_N_c_193_n N_A_27_424#_c_413_n 0.0034415f $X=1.265 $Y=2.045 $X2=0
+ $Y2=0
cc_194 N_GATE_N_c_193_n N_A_27_424#_c_396_n 0.00306552f $X=1.265 $Y=2.045 $X2=0
+ $Y2=0
cc_195 N_GATE_N_M1003_g N_A_373_74#_c_492_n 5.03894e-19 $X=1.08 $Y=0.74 $X2=0
+ $Y2=0
cc_196 N_GATE_N_c_193_n N_VPWR_c_881_n 0.00588137f $X=1.265 $Y=2.045 $X2=0 $Y2=0
cc_197 N_GATE_N_c_193_n N_VPWR_c_888_n 0.00302115f $X=1.265 $Y=2.045 $X2=0 $Y2=0
cc_198 N_GATE_N_c_193_n N_VPWR_c_880_n 0.00377517f $X=1.265 $Y=2.045 $X2=0 $Y2=0
cc_199 N_GATE_N_M1003_g N_VGND_c_1040_n 0.0103395f $X=1.08 $Y=0.74 $X2=0 $Y2=0
cc_200 N_GATE_N_M1003_g N_VGND_c_1049_n 0.00434272f $X=1.08 $Y=0.74 $X2=0 $Y2=0
cc_201 N_GATE_N_M1003_g N_VGND_c_1052_n 0.00830058f $X=1.08 $Y=0.74 $X2=0 $Y2=0
cc_202 N_A_231_74#_c_224_n N_A_27_424#_M1001_g 0.010715f $X=3.28 $Y=1.215 $X2=0
+ $Y2=0
cc_203 N_A_231_74#_c_225_n N_A_27_424#_M1001_g 6.03382e-19 $X=3.365 $Y=1.97
+ $X2=0 $Y2=0
cc_204 N_A_231_74#_c_228_n N_A_27_424#_M1001_g 0.00366726f $X=2.37 $Y=1.215
+ $X2=0 $Y2=0
cc_205 N_A_231_74#_c_229_n N_A_27_424#_M1001_g 0.00724447f $X=2.35 $Y=1.385
+ $X2=0 $Y2=0
cc_206 N_A_231_74#_c_230_n N_A_27_424#_M1001_g 0.00115954f $X=3.445 $Y=1.215
+ $X2=0 $Y2=0
cc_207 N_A_231_74#_c_232_n N_A_27_424#_M1001_g 0.0173949f $X=2.332 $Y=1.22 $X2=0
+ $Y2=0
cc_208 N_A_231_74#_c_233_n N_A_27_424#_M1001_g 0.0659836f $X=3.445 $Y=1.12 $X2=0
+ $Y2=0
cc_209 N_A_231_74#_c_223_n N_A_27_424#_c_384_n 0.0102232f $X=2.36 $Y=1.795 $X2=0
+ $Y2=0
cc_210 N_A_231_74#_c_235_n N_A_27_424#_c_384_n 0.0249404f $X=2.36 $Y=1.885 $X2=0
+ $Y2=0
cc_211 N_A_231_74#_c_237_n N_A_27_424#_c_384_n 5.39985e-19 $X=2.385 $Y=2.305
+ $X2=0 $Y2=0
cc_212 N_A_231_74#_c_238_n N_A_27_424#_c_384_n 0.00106107f $X=2.47 $Y=2.22 $X2=0
+ $Y2=0
cc_213 N_A_231_74#_c_224_n N_A_27_424#_c_384_n 0.001253f $X=3.28 $Y=1.215 $X2=0
+ $Y2=0
cc_214 N_A_231_74#_c_266_p N_A_27_424#_c_384_n 0.0083189f $X=3.205 $Y=2.905
+ $X2=0 $Y2=0
cc_215 N_A_231_74#_c_225_n N_A_27_424#_c_384_n 0.00655083f $X=3.365 $Y=1.97
+ $X2=0 $Y2=0
cc_216 N_A_231_74#_c_241_n N_A_27_424#_c_384_n 0.00170343f $X=3.29 $Y=2.99 $X2=0
+ $Y2=0
cc_217 N_A_231_74#_c_228_n N_A_27_424#_c_384_n 0.00204989f $X=2.37 $Y=1.215
+ $X2=0 $Y2=0
cc_218 N_A_231_74#_c_229_n N_A_27_424#_c_384_n 0.00459342f $X=2.35 $Y=1.385
+ $X2=0 $Y2=0
cc_219 N_A_231_74#_c_271_p N_A_27_424#_c_384_n 0.00131666f $X=3.365 $Y=2.055
+ $X2=0 $Y2=0
cc_220 N_A_231_74#_c_243_n N_A_27_424#_c_392_n 0.0113988f $X=1.54 $Y=2.305 $X2=0
+ $Y2=0
cc_221 N_A_231_74#_c_227_n N_A_27_424#_c_392_n 0.00166419f $X=1.54 $Y=2.1 $X2=0
+ $Y2=0
cc_222 N_A_231_74#_c_243_n N_A_27_424#_c_405_n 0.0232648f $X=1.54 $Y=2.305 $X2=0
+ $Y2=0
cc_223 N_A_231_74#_M1015_d N_A_27_424#_c_393_n 0.00696f $X=1.34 $Y=2.12 $X2=0
+ $Y2=0
cc_224 N_A_231_74#_c_237_n N_A_27_424#_c_393_n 0.00792524f $X=2.385 $Y=2.305
+ $X2=0 $Y2=0
cc_225 N_A_231_74#_c_243_n N_A_27_424#_c_393_n 0.0209187f $X=1.54 $Y=2.305 $X2=0
+ $Y2=0
cc_226 N_A_231_74#_c_235_n N_A_27_424#_c_439_n 0.0132063f $X=2.36 $Y=1.885 $X2=0
+ $Y2=0
cc_227 N_A_231_74#_c_237_n N_A_27_424#_c_439_n 0.0310283f $X=2.385 $Y=2.305
+ $X2=0 $Y2=0
cc_228 N_A_231_74#_c_266_p N_A_27_424#_c_439_n 0.0113396f $X=3.205 $Y=2.905
+ $X2=0 $Y2=0
cc_229 N_A_231_74#_c_235_n N_A_27_424#_c_394_n 0.00487321f $X=2.36 $Y=1.885
+ $X2=0 $Y2=0
cc_230 N_A_231_74#_c_237_n N_A_27_424#_c_394_n 0.0129839f $X=2.385 $Y=2.305
+ $X2=0 $Y2=0
cc_231 N_A_231_74#_c_238_n N_A_27_424#_c_394_n 0.0263033f $X=2.47 $Y=2.22 $X2=0
+ $Y2=0
cc_232 N_A_231_74#_c_266_p N_A_27_424#_c_394_n 0.0250344f $X=3.205 $Y=2.905
+ $X2=0 $Y2=0
cc_233 N_A_231_74#_c_225_n N_A_27_424#_c_394_n 0.00653634f $X=3.365 $Y=1.97
+ $X2=0 $Y2=0
cc_234 N_A_231_74#_c_271_p N_A_27_424#_c_394_n 0.0106133f $X=3.365 $Y=2.055
+ $X2=0 $Y2=0
cc_235 N_A_231_74#_c_235_n N_A_27_424#_c_396_n 0.00588648f $X=2.36 $Y=1.885
+ $X2=0 $Y2=0
cc_236 N_A_231_74#_c_237_n N_A_27_424#_c_396_n 0.0131009f $X=2.385 $Y=2.305
+ $X2=0 $Y2=0
cc_237 N_A_231_74#_c_223_n N_A_27_424#_c_388_n 2.68633e-19 $X=2.36 $Y=1.795
+ $X2=0 $Y2=0
cc_238 N_A_231_74#_c_224_n N_A_27_424#_c_388_n 0.0249535f $X=3.28 $Y=1.215 $X2=0
+ $Y2=0
cc_239 N_A_231_74#_c_225_n N_A_27_424#_c_388_n 0.0211654f $X=3.365 $Y=1.97 $X2=0
+ $Y2=0
cc_240 N_A_231_74#_c_228_n N_A_27_424#_c_388_n 0.0263033f $X=2.37 $Y=1.215 $X2=0
+ $Y2=0
cc_241 N_A_231_74#_c_237_n N_A_373_74#_M1005_s 0.00877025f $X=2.385 $Y=2.305
+ $X2=0 $Y2=0
cc_242 N_A_231_74#_c_236_n N_A_373_74#_c_498_n 0.0128379f $X=3.935 $Y=2.465
+ $X2=0 $Y2=0
cc_243 N_A_231_74#_c_225_n N_A_373_74#_c_498_n 0.00218987f $X=3.365 $Y=1.97
+ $X2=0 $Y2=0
cc_244 N_A_231_74#_c_240_n N_A_373_74#_c_498_n 0.0132479f $X=3.96 $Y=2.99 $X2=0
+ $Y2=0
cc_245 N_A_231_74#_c_242_n N_A_373_74#_c_498_n 4.82699e-19 $X=4.125 $Y=2.215
+ $X2=0 $Y2=0
cc_246 N_A_231_74#_c_271_p N_A_373_74#_c_498_n 0.0101569f $X=3.365 $Y=2.055
+ $X2=0 $Y2=0
cc_247 N_A_231_74#_c_245_n N_A_373_74#_c_498_n 0.00937594f $X=3.935 $Y=2.257
+ $X2=0 $Y2=0
cc_248 N_A_231_74#_c_242_n N_A_373_74#_c_499_n 2.66559e-19 $X=4.125 $Y=2.215
+ $X2=0 $Y2=0
cc_249 N_A_231_74#_c_245_n N_A_373_74#_c_499_n 0.0128426f $X=3.935 $Y=2.257
+ $X2=0 $Y2=0
cc_250 N_A_231_74#_c_225_n N_A_373_74#_c_500_n 0.00711042f $X=3.365 $Y=1.97
+ $X2=0 $Y2=0
cc_251 N_A_231_74#_c_230_n N_A_373_74#_c_500_n 0.00105979f $X=3.445 $Y=1.215
+ $X2=0 $Y2=0
cc_252 N_A_231_74#_c_231_n N_A_373_74#_c_500_n 0.0159928f $X=3.445 $Y=1.285
+ $X2=0 $Y2=0
cc_253 N_A_231_74#_c_225_n N_A_373_74#_c_491_n 0.00470863f $X=3.365 $Y=1.97
+ $X2=0 $Y2=0
cc_254 N_A_231_74#_c_226_n N_A_373_74#_c_492_n 0.0371737f $X=1.295 $Y=0.515
+ $X2=0 $Y2=0
cc_255 N_A_231_74#_c_232_n N_A_373_74#_c_492_n 0.011043f $X=2.332 $Y=1.22 $X2=0
+ $Y2=0
cc_256 N_A_231_74#_c_223_n N_A_373_74#_c_493_n 0.00335444f $X=2.36 $Y=1.795
+ $X2=0 $Y2=0
cc_257 N_A_231_74#_c_238_n N_A_373_74#_c_493_n 0.00679791f $X=2.47 $Y=2.22 $X2=0
+ $Y2=0
cc_258 N_A_231_74#_c_226_n N_A_373_74#_c_493_n 0.0580967f $X=1.295 $Y=0.515
+ $X2=0 $Y2=0
cc_259 N_A_231_74#_c_228_n N_A_373_74#_c_493_n 0.0318045f $X=2.37 $Y=1.215 $X2=0
+ $Y2=0
cc_260 N_A_231_74#_c_232_n N_A_373_74#_c_493_n 0.0137414f $X=2.332 $Y=1.22 $X2=0
+ $Y2=0
cc_261 N_A_231_74#_c_224_n N_A_373_74#_c_525_n 0.0445673f $X=3.28 $Y=1.215 $X2=0
+ $Y2=0
cc_262 N_A_231_74#_c_228_n N_A_373_74#_c_525_n 0.0259664f $X=2.37 $Y=1.215 $X2=0
+ $Y2=0
cc_263 N_A_231_74#_c_229_n N_A_373_74#_c_525_n 0.00107295f $X=2.35 $Y=1.385
+ $X2=0 $Y2=0
cc_264 N_A_231_74#_c_230_n N_A_373_74#_c_525_n 0.0226425f $X=3.445 $Y=1.215
+ $X2=0 $Y2=0
cc_265 N_A_231_74#_c_231_n N_A_373_74#_c_525_n 0.00113748f $X=3.445 $Y=1.285
+ $X2=0 $Y2=0
cc_266 N_A_231_74#_c_232_n N_A_373_74#_c_525_n 0.00990074f $X=2.332 $Y=1.22
+ $X2=0 $Y2=0
cc_267 N_A_231_74#_c_233_n N_A_373_74#_c_525_n 0.012479f $X=3.445 $Y=1.12 $X2=0
+ $Y2=0
cc_268 N_A_231_74#_c_230_n N_A_373_74#_c_494_n 0.0173696f $X=3.445 $Y=1.215
+ $X2=0 $Y2=0
cc_269 N_A_231_74#_c_231_n N_A_373_74#_c_494_n 0.00125982f $X=3.445 $Y=1.285
+ $X2=0 $Y2=0
cc_270 N_A_231_74#_c_233_n N_A_373_74#_c_494_n 0.00324092f $X=3.445 $Y=1.12
+ $X2=0 $Y2=0
cc_271 N_A_231_74#_c_230_n N_A_373_74#_c_495_n 0.00125982f $X=3.445 $Y=1.215
+ $X2=0 $Y2=0
cc_272 N_A_231_74#_c_231_n N_A_373_74#_c_495_n 0.0151253f $X=3.445 $Y=1.285
+ $X2=0 $Y2=0
cc_273 N_A_231_74#_c_245_n N_A_373_74#_c_495_n 0.0024768f $X=3.935 $Y=2.257
+ $X2=0 $Y2=0
cc_274 N_A_231_74#_c_226_n N_A_373_74#_c_496_n 0.0164674f $X=1.295 $Y=0.515
+ $X2=0 $Y2=0
cc_275 N_A_231_74#_c_232_n N_A_373_74#_c_496_n 0.00194281f $X=2.332 $Y=1.22
+ $X2=0 $Y2=0
cc_276 N_A_231_74#_c_223_n N_A_373_74#_c_503_n 0.00380229f $X=2.36 $Y=1.795
+ $X2=0 $Y2=0
cc_277 N_A_231_74#_c_235_n N_A_373_74#_c_503_n 0.00360146f $X=2.36 $Y=1.885
+ $X2=0 $Y2=0
cc_278 N_A_231_74#_c_237_n N_A_373_74#_c_503_n 0.0284063f $X=2.385 $Y=2.305
+ $X2=0 $Y2=0
cc_279 N_A_231_74#_c_238_n N_A_373_74#_c_503_n 0.0249181f $X=2.47 $Y=2.22 $X2=0
+ $Y2=0
cc_280 N_A_231_74#_c_227_n N_A_373_74#_c_503_n 0.0263647f $X=1.54 $Y=2.1 $X2=0
+ $Y2=0
cc_281 N_A_231_74#_c_228_n N_A_373_74#_c_503_n 0.00234718f $X=2.37 $Y=1.215
+ $X2=0 $Y2=0
cc_282 N_A_231_74#_c_229_n N_A_373_74#_c_503_n 0.00180929f $X=2.35 $Y=1.385
+ $X2=0 $Y2=0
cc_283 N_A_231_74#_c_233_n N_A_373_74#_c_497_n 0.0102577f $X=3.445 $Y=1.12 $X2=0
+ $Y2=0
cc_284 N_A_231_74#_c_236_n N_A_889_92#_c_601_n 0.00984643f $X=3.935 $Y=2.465
+ $X2=0 $Y2=0
cc_285 N_A_231_74#_c_240_n N_A_889_92#_c_601_n 0.00177437f $X=3.96 $Y=2.99 $X2=0
+ $Y2=0
cc_286 N_A_231_74#_c_242_n N_A_889_92#_c_601_n 0.00787719f $X=4.125 $Y=2.215
+ $X2=0 $Y2=0
cc_287 N_A_231_74#_c_245_n N_A_889_92#_c_601_n 0.0198046f $X=3.935 $Y=2.257
+ $X2=0 $Y2=0
cc_288 N_A_231_74#_c_242_n N_A_889_92#_c_609_n 0.0144629f $X=4.125 $Y=2.215
+ $X2=0 $Y2=0
cc_289 N_A_231_74#_c_245_n N_A_889_92#_c_609_n 9.29575e-19 $X=3.935 $Y=2.257
+ $X2=0 $Y2=0
cc_290 N_A_231_74#_c_240_n N_A_686_74#_M1012_d 0.00334086f $X=3.96 $Y=2.99 $X2=0
+ $Y2=0
cc_291 N_A_231_74#_c_233_n N_A_686_74#_c_721_n 0.0100959f $X=3.445 $Y=1.12 $X2=0
+ $Y2=0
cc_292 N_A_231_74#_c_242_n N_A_686_74#_c_727_n 0.018783f $X=4.125 $Y=2.215 $X2=0
+ $Y2=0
cc_293 N_A_231_74#_c_245_n N_A_686_74#_c_727_n 0.00213123f $X=3.935 $Y=2.257
+ $X2=0 $Y2=0
cc_294 N_A_231_74#_c_225_n N_A_686_74#_c_728_n 0.0135296f $X=3.365 $Y=1.97 $X2=0
+ $Y2=0
cc_295 N_A_231_74#_c_236_n N_A_686_74#_c_729_n 0.00229161f $X=3.935 $Y=2.465
+ $X2=0 $Y2=0
cc_296 N_A_231_74#_c_240_n N_A_686_74#_c_729_n 0.0201163f $X=3.96 $Y=2.99 $X2=0
+ $Y2=0
cc_297 N_A_231_74#_c_225_n N_A_686_74#_c_730_n 0.0126059f $X=3.365 $Y=1.97 $X2=0
+ $Y2=0
cc_298 N_A_231_74#_c_242_n N_A_686_74#_c_730_n 0.052421f $X=4.125 $Y=2.215 $X2=0
+ $Y2=0
cc_299 N_A_231_74#_c_271_p N_A_686_74#_c_730_n 0.0124673f $X=3.365 $Y=2.055
+ $X2=0 $Y2=0
cc_300 N_A_231_74#_c_245_n N_A_686_74#_c_730_n 0.00391663f $X=3.935 $Y=2.257
+ $X2=0 $Y2=0
cc_301 N_A_231_74#_c_237_n N_VPWR_M1005_d 0.00232895f $X=2.385 $Y=2.305 $X2=0
+ $Y2=0
cc_302 N_A_231_74#_c_238_n N_VPWR_M1005_d 0.00239219f $X=2.47 $Y=2.22 $X2=0
+ $Y2=0
cc_303 N_A_231_74#_c_235_n N_VPWR_c_882_n 8.65703e-19 $X=2.36 $Y=1.885 $X2=0
+ $Y2=0
cc_304 N_A_231_74#_c_266_p N_VPWR_c_882_n 2.36327e-19 $X=3.205 $Y=2.905 $X2=0
+ $Y2=0
cc_305 N_A_231_74#_c_241_n N_VPWR_c_882_n 0.0102734f $X=3.29 $Y=2.99 $X2=0 $Y2=0
cc_306 N_A_231_74#_c_235_n N_VPWR_c_888_n 0.00358037f $X=2.36 $Y=1.885 $X2=0
+ $Y2=0
cc_307 N_A_231_74#_c_236_n N_VPWR_c_889_n 0.00278223f $X=3.935 $Y=2.465 $X2=0
+ $Y2=0
cc_308 N_A_231_74#_c_240_n N_VPWR_c_889_n 0.0658254f $X=3.96 $Y=2.99 $X2=0 $Y2=0
cc_309 N_A_231_74#_c_241_n N_VPWR_c_889_n 0.0121867f $X=3.29 $Y=2.99 $X2=0 $Y2=0
cc_310 N_A_231_74#_c_235_n N_VPWR_c_880_n 0.0049649f $X=2.36 $Y=1.885 $X2=0
+ $Y2=0
cc_311 N_A_231_74#_c_236_n N_VPWR_c_880_n 0.00356419f $X=3.935 $Y=2.465 $X2=0
+ $Y2=0
cc_312 N_A_231_74#_c_240_n N_VPWR_c_880_n 0.0366416f $X=3.96 $Y=2.99 $X2=0 $Y2=0
cc_313 N_A_231_74#_c_241_n N_VPWR_c_880_n 0.00660921f $X=3.29 $Y=2.99 $X2=0
+ $Y2=0
cc_314 N_A_231_74#_c_236_n N_VPWR_c_895_n 4.88458e-19 $X=3.935 $Y=2.465 $X2=0
+ $Y2=0
cc_315 N_A_231_74#_c_240_n N_VPWR_c_895_n 0.00800512f $X=3.96 $Y=2.99 $X2=0
+ $Y2=0
cc_316 N_A_231_74#_c_242_n N_VPWR_c_895_n 0.0166602f $X=4.125 $Y=2.215 $X2=0
+ $Y2=0
cc_317 N_A_231_74#_c_266_p A_611_392# 0.0112873f $X=3.205 $Y=2.905 $X2=-0.19
+ $Y2=-0.245
cc_318 N_A_231_74#_c_241_n A_611_392# 6.51498e-19 $X=3.29 $Y=2.99 $X2=-0.19
+ $Y2=-0.245
cc_319 N_A_231_74#_c_271_p A_611_392# 0.00506284f $X=3.365 $Y=2.055 $X2=-0.19
+ $Y2=-0.245
cc_320 N_A_231_74#_c_240_n A_802_508# 0.00100794f $X=3.96 $Y=2.99 $X2=-0.19
+ $Y2=-0.245
cc_321 N_A_231_74#_c_242_n A_802_508# 0.00636757f $X=4.125 $Y=2.215 $X2=-0.19
+ $Y2=-0.245
cc_322 N_A_231_74#_c_226_n N_VGND_c_1040_n 0.0307709f $X=1.295 $Y=0.515 $X2=0
+ $Y2=0
cc_323 N_A_231_74#_c_233_n N_VGND_c_1044_n 0.00433387f $X=3.445 $Y=1.12 $X2=0
+ $Y2=0
cc_324 N_A_231_74#_c_226_n N_VGND_c_1049_n 0.0241574f $X=1.295 $Y=0.515 $X2=0
+ $Y2=0
cc_325 N_A_231_74#_c_232_n N_VGND_c_1049_n 0.00434272f $X=2.332 $Y=1.22 $X2=0
+ $Y2=0
cc_326 N_A_231_74#_c_226_n N_VGND_c_1052_n 0.019939f $X=1.295 $Y=0.515 $X2=0
+ $Y2=0
cc_327 N_A_231_74#_c_232_n N_VGND_c_1052_n 0.00439653f $X=2.332 $Y=1.22 $X2=0
+ $Y2=0
cc_328 N_A_231_74#_c_233_n N_VGND_c_1052_n 0.00439408f $X=3.445 $Y=1.12 $X2=0
+ $Y2=0
cc_329 N_A_231_74#_c_232_n N_VGND_c_1054_n 0.00578246f $X=2.332 $Y=1.22 $X2=0
+ $Y2=0
cc_330 N_A_231_74#_c_233_n N_VGND_c_1054_n 0.0012862f $X=3.445 $Y=1.12 $X2=0
+ $Y2=0
cc_331 N_A_27_424#_c_439_n N_A_373_74#_M1005_s 0.00713378f $X=2.74 $Y=2.645
+ $X2=0 $Y2=0
cc_332 N_A_27_424#_c_396_n N_A_373_74#_M1005_s 0.00394145f $X=1.93 $Y=2.645
+ $X2=0 $Y2=0
cc_333 N_A_27_424#_c_384_n N_A_373_74#_c_498_n 0.0467931f $X=2.98 $Y=1.885 $X2=0
+ $Y2=0
cc_334 N_A_27_424#_c_394_n N_A_373_74#_c_498_n 3.6024e-19 $X=2.825 $Y=2.56 $X2=0
+ $Y2=0
cc_335 N_A_27_424#_c_384_n N_A_373_74#_c_500_n 0.0101838f $X=2.98 $Y=1.885 $X2=0
+ $Y2=0
cc_336 N_A_27_424#_M1001_g N_A_373_74#_c_525_n 0.0124889f $X=2.965 $Y=0.69 $X2=0
+ $Y2=0
cc_337 N_A_27_424#_M1001_g N_A_686_74#_c_721_n 7.17942e-19 $X=2.965 $Y=0.69
+ $X2=0 $Y2=0
cc_338 N_A_27_424#_c_392_n N_VPWR_M1019_d 0.0108651f $X=1.065 $Y=2.155 $X2=-0.19
+ $Y2=-0.245
cc_339 N_A_27_424#_c_405_n N_VPWR_M1019_d 0.00557572f $X=1.15 $Y=2.73 $X2=-0.19
+ $Y2=-0.245
cc_340 N_A_27_424#_c_413_n N_VPWR_M1019_d 0.00259674f $X=1.235 $Y=2.815
+ $X2=-0.19 $Y2=-0.245
cc_341 N_A_27_424#_c_439_n N_VPWR_M1005_d 0.0124927f $X=2.74 $Y=2.645 $X2=0
+ $Y2=0
cc_342 N_A_27_424#_c_394_n N_VPWR_M1005_d 0.00609494f $X=2.825 $Y=2.56 $X2=0
+ $Y2=0
cc_343 N_A_27_424#_c_391_n N_VPWR_c_881_n 0.038474f $X=0.28 $Y=2.265 $X2=0 $Y2=0
cc_344 N_A_27_424#_c_392_n N_VPWR_c_881_n 0.0219335f $X=1.065 $Y=2.155 $X2=0
+ $Y2=0
cc_345 N_A_27_424#_c_405_n N_VPWR_c_881_n 0.0244185f $X=1.15 $Y=2.73 $X2=0 $Y2=0
cc_346 N_A_27_424#_c_413_n N_VPWR_c_881_n 0.0144778f $X=1.235 $Y=2.815 $X2=0
+ $Y2=0
cc_347 N_A_27_424#_c_384_n N_VPWR_c_882_n 0.00437408f $X=2.98 $Y=1.885 $X2=0
+ $Y2=0
cc_348 N_A_27_424#_c_439_n N_VPWR_c_882_n 0.0254173f $X=2.74 $Y=2.645 $X2=0
+ $Y2=0
cc_349 N_A_27_424#_c_391_n N_VPWR_c_887_n 0.0119584f $X=0.28 $Y=2.265 $X2=0
+ $Y2=0
cc_350 N_A_27_424#_c_393_n N_VPWR_c_888_n 0.0174377f $X=1.845 $Y=2.815 $X2=0
+ $Y2=0
cc_351 N_A_27_424#_c_413_n N_VPWR_c_888_n 0.00461086f $X=1.235 $Y=2.815 $X2=0
+ $Y2=0
cc_352 N_A_27_424#_c_439_n N_VPWR_c_888_n 0.00813902f $X=2.74 $Y=2.645 $X2=0
+ $Y2=0
cc_353 N_A_27_424#_c_396_n N_VPWR_c_888_n 0.00539346f $X=1.93 $Y=2.645 $X2=0
+ $Y2=0
cc_354 N_A_27_424#_c_384_n N_VPWR_c_889_n 0.00456824f $X=2.98 $Y=1.885 $X2=0
+ $Y2=0
cc_355 N_A_27_424#_c_439_n N_VPWR_c_889_n 9.62119e-19 $X=2.74 $Y=2.645 $X2=0
+ $Y2=0
cc_356 N_A_27_424#_c_384_n N_VPWR_c_880_n 0.00896864f $X=2.98 $Y=1.885 $X2=0
+ $Y2=0
cc_357 N_A_27_424#_c_391_n N_VPWR_c_880_n 0.00989813f $X=0.28 $Y=2.265 $X2=0
+ $Y2=0
cc_358 N_A_27_424#_c_393_n N_VPWR_c_880_n 0.0198563f $X=1.845 $Y=2.815 $X2=0
+ $Y2=0
cc_359 N_A_27_424#_c_413_n N_VPWR_c_880_n 0.00574357f $X=1.235 $Y=2.815 $X2=0
+ $Y2=0
cc_360 N_A_27_424#_c_439_n N_VPWR_c_880_n 0.0182435f $X=2.74 $Y=2.645 $X2=0
+ $Y2=0
cc_361 N_A_27_424#_c_396_n N_VPWR_c_880_n 0.00574775f $X=1.93 $Y=2.645 $X2=0
+ $Y2=0
cc_362 N_A_27_424#_c_385_n N_VGND_c_1040_n 0.0206573f $X=0.272 $Y=0.913 $X2=0
+ $Y2=0
cc_363 N_A_27_424#_M1001_g N_VGND_c_1044_n 0.00384553f $X=2.965 $Y=0.69 $X2=0
+ $Y2=0
cc_364 N_A_27_424#_c_385_n N_VGND_c_1048_n 0.00870476f $X=0.272 $Y=0.913 $X2=0
+ $Y2=0
cc_365 N_A_27_424#_M1001_g N_VGND_c_1052_n 0.00371083f $X=2.965 $Y=0.69 $X2=0
+ $Y2=0
cc_366 N_A_27_424#_c_385_n N_VGND_c_1052_n 0.0113983f $X=0.272 $Y=0.913 $X2=0
+ $Y2=0
cc_367 N_A_27_424#_M1001_g N_VGND_c_1054_n 0.0137918f $X=2.965 $Y=0.69 $X2=0
+ $Y2=0
cc_368 N_A_373_74#_c_491_n N_A_889_92#_M1022_g 0.00512524f $X=3.95 $Y=1.69 $X2=0
+ $Y2=0
cc_369 N_A_373_74#_c_494_n N_A_889_92#_M1022_g 5.60778e-19 $X=4.04 $Y=1.285
+ $X2=0 $Y2=0
cc_370 N_A_373_74#_c_497_n N_A_889_92#_M1022_g 0.0516229f $X=4.04 $Y=1.12 $X2=0
+ $Y2=0
cc_371 N_A_373_74#_c_499_n N_A_889_92#_c_601_n 0.00512524f $X=3.875 $Y=1.765
+ $X2=0 $Y2=0
cc_372 N_A_373_74#_c_525_n N_A_686_74#_M1002_d 0.0144935f $X=3.875 $Y=0.865
+ $X2=-0.19 $Y2=-0.245
cc_373 N_A_373_74#_c_494_n N_A_686_74#_M1002_d 9.37577e-19 $X=4.04 $Y=1.285
+ $X2=-0.19 $Y2=-0.245
cc_374 N_A_373_74#_c_525_n N_A_686_74#_c_721_n 0.0510609f $X=3.875 $Y=0.865
+ $X2=0 $Y2=0
cc_375 N_A_373_74#_c_495_n N_A_686_74#_c_721_n 5.49906e-19 $X=4.04 $Y=1.285
+ $X2=0 $Y2=0
cc_376 N_A_373_74#_c_497_n N_A_686_74#_c_721_n 0.0110691f $X=4.04 $Y=1.12 $X2=0
+ $Y2=0
cc_377 N_A_373_74#_c_499_n N_A_686_74#_c_727_n 0.00881468f $X=3.875 $Y=1.765
+ $X2=0 $Y2=0
cc_378 N_A_373_74#_c_491_n N_A_686_74#_c_727_n 0.00526469f $X=3.95 $Y=1.69 $X2=0
+ $Y2=0
cc_379 N_A_373_74#_c_525_n N_A_686_74#_c_727_n 0.00229912f $X=3.875 $Y=0.865
+ $X2=0 $Y2=0
cc_380 N_A_373_74#_c_494_n N_A_686_74#_c_727_n 0.0256239f $X=4.04 $Y=1.285 $X2=0
+ $Y2=0
cc_381 N_A_373_74#_c_495_n N_A_686_74#_c_727_n 7.13049e-19 $X=4.04 $Y=1.285
+ $X2=0 $Y2=0
cc_382 N_A_373_74#_c_499_n N_A_686_74#_c_728_n 0.0056327f $X=3.875 $Y=1.765
+ $X2=0 $Y2=0
cc_383 N_A_373_74#_c_525_n N_A_686_74#_c_728_n 0.00523357f $X=3.875 $Y=0.865
+ $X2=0 $Y2=0
cc_384 N_A_373_74#_c_498_n N_A_686_74#_c_729_n 0.00390285f $X=3.4 $Y=1.885 $X2=0
+ $Y2=0
cc_385 N_A_373_74#_c_499_n N_A_686_74#_c_729_n 0.00262654f $X=3.875 $Y=1.765
+ $X2=0 $Y2=0
cc_386 N_A_373_74#_c_498_n N_A_686_74#_c_730_n 0.0060239f $X=3.4 $Y=1.885 $X2=0
+ $Y2=0
cc_387 N_A_373_74#_c_499_n N_A_686_74#_c_730_n 0.00639693f $X=3.875 $Y=1.765
+ $X2=0 $Y2=0
cc_388 N_A_373_74#_c_500_n N_A_686_74#_c_730_n 9.34794e-19 $X=3.49 $Y=1.765
+ $X2=0 $Y2=0
cc_389 N_A_373_74#_c_491_n N_A_686_74#_c_723_n 0.00359753f $X=3.95 $Y=1.69 $X2=0
+ $Y2=0
cc_390 N_A_373_74#_c_495_n N_A_686_74#_c_723_n 0.00141263f $X=4.04 $Y=1.285
+ $X2=0 $Y2=0
cc_391 N_A_373_74#_c_525_n N_A_686_74#_c_724_n 0.0133619f $X=3.875 $Y=0.865
+ $X2=0 $Y2=0
cc_392 N_A_373_74#_c_494_n N_A_686_74#_c_724_n 0.0383881f $X=4.04 $Y=1.285 $X2=0
+ $Y2=0
cc_393 N_A_373_74#_c_497_n N_A_686_74#_c_724_n 0.00535323f $X=4.04 $Y=1.12 $X2=0
+ $Y2=0
cc_394 N_A_373_74#_c_498_n N_VPWR_c_889_n 0.00278271f $X=3.4 $Y=1.885 $X2=0
+ $Y2=0
cc_395 N_A_373_74#_c_498_n N_VPWR_c_880_n 0.00354422f $X=3.4 $Y=1.885 $X2=0
+ $Y2=0
cc_396 N_A_373_74#_c_525_n N_VGND_M1013_d 0.0119294f $X=3.875 $Y=0.865 $X2=0
+ $Y2=0
cc_397 N_A_373_74#_c_497_n N_VGND_c_1044_n 6.60767e-19 $X=4.04 $Y=1.12 $X2=0
+ $Y2=0
cc_398 N_A_373_74#_c_492_n N_VGND_c_1049_n 0.0145091f $X=2.01 $Y=0.515 $X2=0
+ $Y2=0
cc_399 N_A_373_74#_c_492_n N_VGND_c_1052_n 0.0119768f $X=2.01 $Y=0.515 $X2=0
+ $Y2=0
cc_400 N_A_373_74#_c_525_n N_VGND_c_1052_n 0.0241286f $X=3.875 $Y=0.865 $X2=0
+ $Y2=0
cc_401 N_A_373_74#_c_492_n N_VGND_c_1054_n 0.0102391f $X=2.01 $Y=0.515 $X2=0
+ $Y2=0
cc_402 N_A_373_74#_c_525_n N_VGND_c_1054_n 0.0376298f $X=3.875 $Y=0.865 $X2=0
+ $Y2=0
cc_403 N_A_373_74#_c_525_n A_608_74# 0.00377716f $X=3.875 $Y=0.865 $X2=-0.19
+ $Y2=-0.245
cc_404 N_A_889_92#_c_601_n N_A_686_74#_c_718_n 0.00435947f $X=4.62 $Y=2.465
+ $X2=0 $Y2=0
cc_405 N_A_889_92#_c_597_n N_A_686_74#_c_718_n 0.0110373f $X=5.375 $Y=1.72 $X2=0
+ $Y2=0
cc_406 N_A_889_92#_c_607_n N_A_686_74#_c_718_n 0.0130233f $X=5.78 $Y=2.685 $X2=0
+ $Y2=0
cc_407 N_A_889_92#_c_624_p N_A_686_74#_c_718_n 0.0333962f $X=5.945 $Y=2.005
+ $X2=0 $Y2=0
cc_408 N_A_889_92#_c_596_n N_A_686_74#_c_719_n 0.00480714f $X=5.375 $Y=0.515
+ $X2=0 $Y2=0
cc_409 N_A_889_92#_M1022_g N_A_686_74#_c_720_n 0.0177129f $X=4.52 $Y=0.8 $X2=0
+ $Y2=0
cc_410 N_A_889_92#_c_601_n N_A_686_74#_c_720_n 5.38205e-19 $X=4.62 $Y=2.465
+ $X2=0 $Y2=0
cc_411 N_A_889_92#_c_597_n N_A_686_74#_c_720_n 0.0163508f $X=5.375 $Y=1.72 $X2=0
+ $Y2=0
cc_412 N_A_889_92#_c_598_n N_A_686_74#_c_720_n 0.00349862f $X=5.335 $Y=1.05
+ $X2=0 $Y2=0
cc_413 N_A_889_92#_c_609_n N_A_686_74#_c_720_n 0.010421f $X=5.29 $Y=2.005 $X2=0
+ $Y2=0
cc_414 N_A_889_92#_c_624_p N_A_686_74#_c_720_n 7.95602e-19 $X=5.945 $Y=2.005
+ $X2=0 $Y2=0
cc_415 N_A_889_92#_M1022_g N_A_686_74#_c_721_n 0.00557158f $X=4.52 $Y=0.8 $X2=0
+ $Y2=0
cc_416 N_A_889_92#_M1022_g N_A_686_74#_c_727_n 4.11677e-19 $X=4.52 $Y=0.8 $X2=0
+ $Y2=0
cc_417 N_A_889_92#_M1022_g N_A_686_74#_c_722_n 3.51925e-19 $X=4.52 $Y=0.8 $X2=0
+ $Y2=0
cc_418 N_A_889_92#_c_601_n N_A_686_74#_c_722_n 0.00230517f $X=4.62 $Y=2.465
+ $X2=0 $Y2=0
cc_419 N_A_889_92#_c_597_n N_A_686_74#_c_722_n 0.0238893f $X=5.375 $Y=1.72 $X2=0
+ $Y2=0
cc_420 N_A_889_92#_c_609_n N_A_686_74#_c_722_n 0.0161469f $X=5.29 $Y=2.005 $X2=0
+ $Y2=0
cc_421 N_A_889_92#_c_601_n N_A_686_74#_c_730_n 2.02023e-19 $X=4.62 $Y=2.465
+ $X2=0 $Y2=0
cc_422 N_A_889_92#_M1022_g N_A_686_74#_c_723_n 0.0163869f $X=4.52 $Y=0.8 $X2=0
+ $Y2=0
cc_423 N_A_889_92#_c_601_n N_A_686_74#_c_723_n 0.0133556f $X=4.62 $Y=2.465 $X2=0
+ $Y2=0
cc_424 N_A_889_92#_c_597_n N_A_686_74#_c_723_n 0.00593094f $X=5.375 $Y=1.72
+ $X2=0 $Y2=0
cc_425 N_A_889_92#_c_609_n N_A_686_74#_c_723_n 0.01548f $X=5.29 $Y=2.005 $X2=0
+ $Y2=0
cc_426 N_A_889_92#_c_624_p N_A_686_74#_c_723_n 0.00252314f $X=5.945 $Y=2.005
+ $X2=0 $Y2=0
cc_427 N_A_889_92#_M1022_g N_A_686_74#_c_724_n 0.0177045f $X=4.52 $Y=0.8 $X2=0
+ $Y2=0
cc_428 N_A_889_92#_c_598_n N_A_686_74#_c_724_n 5.24568e-19 $X=5.335 $Y=1.05
+ $X2=0 $Y2=0
cc_429 N_A_889_92#_c_591_n N_RESET_B_c_811_n 0.0162015f $X=6.52 $Y=1.22
+ $X2=-0.19 $Y2=-0.245
cc_430 N_A_889_92#_c_602_n N_RESET_B_c_812_n 0.0234066f $X=6.535 $Y=1.635 $X2=0
+ $Y2=0
cc_431 N_A_889_92#_c_594_n N_RESET_B_c_812_n 0.0200527f $X=6.535 $Y=1.427 $X2=0
+ $Y2=0
cc_432 N_A_889_92#_c_597_n N_RESET_B_c_812_n 0.00128592f $X=5.375 $Y=1.72 $X2=0
+ $Y2=0
cc_433 N_A_889_92#_c_607_n N_RESET_B_c_812_n 0.00595515f $X=5.78 $Y=2.685 $X2=0
+ $Y2=0
cc_434 N_A_889_92#_c_651_p N_RESET_B_c_812_n 0.0138341f $X=6.35 $Y=1.805 $X2=0
+ $Y2=0
cc_435 N_A_889_92#_c_608_n N_RESET_B_c_812_n 0.00326465f $X=6.435 $Y=1.72 $X2=0
+ $Y2=0
cc_436 N_A_889_92#_c_624_p N_RESET_B_c_812_n 0.0063419f $X=5.945 $Y=2.005 $X2=0
+ $Y2=0
cc_437 N_A_889_92#_c_599_n N_RESET_B_c_812_n 0.00213331f $X=6.645 $Y=1.385 $X2=0
+ $Y2=0
cc_438 N_A_889_92#_c_591_n RESET_B 8.62312e-19 $X=6.52 $Y=1.22 $X2=0 $Y2=0
cc_439 N_A_889_92#_c_594_n RESET_B 3.28967e-19 $X=6.535 $Y=1.427 $X2=0 $Y2=0
cc_440 N_A_889_92#_c_597_n RESET_B 0.0130859f $X=5.375 $Y=1.72 $X2=0 $Y2=0
cc_441 N_A_889_92#_c_624_p RESET_B 0.0183033f $X=5.945 $Y=2.005 $X2=0 $Y2=0
cc_442 N_A_889_92#_c_599_n RESET_B 0.0264685f $X=6.645 $Y=1.385 $X2=0 $Y2=0
cc_443 N_A_889_92#_c_593_n N_A_1437_112#_M1020_g 0.0156195f $X=7.61 $Y=1.22
+ $X2=0 $Y2=0
cc_444 N_A_889_92#_c_592_n N_A_1437_112#_c_843_n 0.0402949f $X=7.595 $Y=1.845
+ $X2=0 $Y2=0
cc_445 N_A_889_92#_c_591_n N_A_1437_112#_c_844_n 5.99084e-19 $X=6.52 $Y=1.22
+ $X2=0 $Y2=0
cc_446 N_A_889_92#_c_592_n N_A_1437_112#_c_844_n 0.00823277f $X=7.595 $Y=1.845
+ $X2=0 $Y2=0
cc_447 N_A_889_92#_c_593_n N_A_1437_112#_c_844_n 0.0139026f $X=7.61 $Y=1.22
+ $X2=0 $Y2=0
cc_448 N_A_889_92#_c_592_n N_A_1437_112#_c_847_n 0.0296909f $X=7.595 $Y=1.845
+ $X2=0 $Y2=0
cc_449 N_A_889_92#_c_592_n N_A_1437_112#_c_845_n 0.0185974f $X=7.595 $Y=1.845
+ $X2=0 $Y2=0
cc_450 N_A_889_92#_c_592_n N_A_1437_112#_c_855_n 0.0140961f $X=7.595 $Y=1.845
+ $X2=0 $Y2=0
cc_451 N_A_889_92#_c_597_n N_VPWR_M1016_d 5.28397e-19 $X=5.375 $Y=1.72 $X2=0
+ $Y2=0
cc_452 N_A_889_92#_c_609_n N_VPWR_M1016_d 0.00385976f $X=5.29 $Y=2.005 $X2=0
+ $Y2=0
cc_453 N_A_889_92#_c_624_p N_VPWR_M1016_d 0.00643476f $X=5.945 $Y=2.005 $X2=0
+ $Y2=0
cc_454 N_A_889_92#_c_651_p N_VPWR_M1007_d 0.00906914f $X=6.35 $Y=1.805 $X2=0
+ $Y2=0
cc_455 N_A_889_92#_c_602_n N_VPWR_c_883_n 0.0041816f $X=6.535 $Y=1.635 $X2=0
+ $Y2=0
cc_456 N_A_889_92#_c_607_n N_VPWR_c_883_n 0.021803f $X=5.78 $Y=2.685 $X2=0 $Y2=0
cc_457 N_A_889_92#_c_651_p N_VPWR_c_883_n 0.0217974f $X=6.35 $Y=1.805 $X2=0
+ $Y2=0
cc_458 N_A_889_92#_c_592_n N_VPWR_c_884_n 0.0106689f $X=7.595 $Y=1.845 $X2=0
+ $Y2=0
cc_459 N_A_889_92#_c_607_n N_VPWR_c_885_n 0.00938905f $X=5.78 $Y=2.685 $X2=0
+ $Y2=0
cc_460 N_A_889_92#_c_601_n N_VPWR_c_889_n 0.00415318f $X=4.62 $Y=2.465 $X2=0
+ $Y2=0
cc_461 N_A_889_92#_c_602_n N_VPWR_c_890_n 0.00487664f $X=6.535 $Y=1.635 $X2=0
+ $Y2=0
cc_462 N_A_889_92#_c_592_n N_VPWR_c_890_n 0.00435405f $X=7.595 $Y=1.845 $X2=0
+ $Y2=0
cc_463 N_A_889_92#_c_601_n N_VPWR_c_880_n 0.00857361f $X=4.62 $Y=2.465 $X2=0
+ $Y2=0
cc_464 N_A_889_92#_c_602_n N_VPWR_c_880_n 0.00505379f $X=6.535 $Y=1.635 $X2=0
+ $Y2=0
cc_465 N_A_889_92#_c_592_n N_VPWR_c_880_n 0.00484898f $X=7.595 $Y=1.845 $X2=0
+ $Y2=0
cc_466 N_A_889_92#_c_607_n N_VPWR_c_880_n 0.0110215f $X=5.78 $Y=2.685 $X2=0
+ $Y2=0
cc_467 N_A_889_92#_c_601_n N_VPWR_c_895_n 0.0185391f $X=4.62 $Y=2.465 $X2=0
+ $Y2=0
cc_468 N_A_889_92#_c_607_n N_VPWR_c_895_n 0.0132644f $X=5.78 $Y=2.685 $X2=0
+ $Y2=0
cc_469 N_A_889_92#_c_609_n N_VPWR_c_895_n 0.0510813f $X=5.29 $Y=2.005 $X2=0
+ $Y2=0
cc_470 N_A_889_92#_c_602_n N_Q_c_991_n 0.00886342f $X=6.535 $Y=1.635 $X2=0 $Y2=0
cc_471 N_A_889_92#_c_592_n N_Q_c_991_n 0.00272082f $X=7.595 $Y=1.845 $X2=0 $Y2=0
cc_472 N_A_889_92#_c_595_n N_Q_c_991_n 0.00747257f $X=7.275 $Y=1.4 $X2=0 $Y2=0
cc_473 N_A_889_92#_c_651_p N_Q_c_991_n 0.0142718f $X=6.35 $Y=1.805 $X2=0 $Y2=0
cc_474 N_A_889_92#_c_599_n N_Q_c_991_n 0.00693673f $X=6.645 $Y=1.385 $X2=0 $Y2=0
cc_475 N_A_889_92#_c_591_n N_Q_c_989_n 0.00323908f $X=6.52 $Y=1.22 $X2=0 $Y2=0
cc_476 N_A_889_92#_c_602_n N_Q_c_989_n 3.02598e-19 $X=6.535 $Y=1.635 $X2=0 $Y2=0
cc_477 N_A_889_92#_c_592_n N_Q_c_989_n 0.00204262f $X=7.595 $Y=1.845 $X2=0 $Y2=0
cc_478 N_A_889_92#_c_594_n N_Q_c_989_n 5.03321e-19 $X=6.535 $Y=1.427 $X2=0 $Y2=0
cc_479 N_A_889_92#_c_595_n N_Q_c_989_n 0.0240419f $X=7.275 $Y=1.4 $X2=0 $Y2=0
cc_480 N_A_889_92#_c_608_n N_Q_c_989_n 0.00420451f $X=6.435 $Y=1.72 $X2=0 $Y2=0
cc_481 N_A_889_92#_c_599_n N_Q_c_989_n 0.0240318f $X=6.645 $Y=1.385 $X2=0 $Y2=0
cc_482 N_A_889_92#_c_592_n Q 0.00131091f $X=7.595 $Y=1.845 $X2=0 $Y2=0
cc_483 N_A_889_92#_c_591_n N_Q_c_990_n 0.0109023f $X=6.52 $Y=1.22 $X2=0 $Y2=0
cc_484 N_A_889_92#_c_593_n N_Q_c_990_n 0.00401054f $X=7.61 $Y=1.22 $X2=0 $Y2=0
cc_485 N_A_889_92#_c_595_n N_Q_c_990_n 0.00731765f $X=7.275 $Y=1.4 $X2=0 $Y2=0
cc_486 N_A_889_92#_c_599_n N_Q_c_990_n 0.0145705f $X=6.645 $Y=1.385 $X2=0 $Y2=0
cc_487 N_A_889_92#_M1022_g N_VGND_c_1041_n 0.0115863f $X=4.52 $Y=0.8 $X2=0 $Y2=0
cc_488 N_A_889_92#_c_596_n N_VGND_c_1041_n 0.0439255f $X=5.375 $Y=0.515 $X2=0
+ $Y2=0
cc_489 N_A_889_92#_c_591_n N_VGND_c_1042_n 0.00884467f $X=6.52 $Y=1.22 $X2=0
+ $Y2=0
cc_490 N_A_889_92#_c_596_n N_VGND_c_1042_n 0.00946037f $X=5.375 $Y=0.515 $X2=0
+ $Y2=0
cc_491 N_A_889_92#_c_599_n N_VGND_c_1042_n 6.69379e-19 $X=6.645 $Y=1.385 $X2=0
+ $Y2=0
cc_492 N_A_889_92#_c_593_n N_VGND_c_1043_n 0.00677853f $X=7.61 $Y=1.22 $X2=0
+ $Y2=0
cc_493 N_A_889_92#_M1022_g N_VGND_c_1044_n 0.0018875f $X=4.52 $Y=0.8 $X2=0 $Y2=0
cc_494 N_A_889_92#_c_596_n N_VGND_c_1046_n 0.0110735f $X=5.375 $Y=0.515 $X2=0
+ $Y2=0
cc_495 N_A_889_92#_c_591_n N_VGND_c_1050_n 0.00428607f $X=6.52 $Y=1.22 $X2=0
+ $Y2=0
cc_496 N_A_889_92#_c_593_n N_VGND_c_1050_n 0.0043356f $X=7.61 $Y=1.22 $X2=0
+ $Y2=0
cc_497 N_A_889_92#_M1022_g N_VGND_c_1052_n 0.00159737f $X=4.52 $Y=0.8 $X2=0
+ $Y2=0
cc_498 N_A_889_92#_c_591_n N_VGND_c_1052_n 0.00808641f $X=6.52 $Y=1.22 $X2=0
+ $Y2=0
cc_499 N_A_889_92#_c_593_n N_VGND_c_1052_n 0.00487769f $X=7.61 $Y=1.22 $X2=0
+ $Y2=0
cc_500 N_A_889_92#_c_596_n N_VGND_c_1052_n 0.00916237f $X=5.375 $Y=0.515 $X2=0
+ $Y2=0
cc_501 N_A_686_74#_c_719_n N_RESET_B_c_811_n 0.0495768f $X=5.59 $Y=1.22
+ $X2=-0.19 $Y2=-0.245
cc_502 N_A_686_74#_c_718_n N_RESET_B_c_812_n 0.0330408f $X=5.545 $Y=1.635 $X2=0
+ $Y2=0
cc_503 N_A_686_74#_c_718_n RESET_B 0.00152604f $X=5.545 $Y=1.635 $X2=0 $Y2=0
cc_504 N_A_686_74#_c_719_n RESET_B 3.10559e-19 $X=5.59 $Y=1.22 $X2=0 $Y2=0
cc_505 N_A_686_74#_c_718_n N_VPWR_c_885_n 0.00484296f $X=5.545 $Y=1.635 $X2=0
+ $Y2=0
cc_506 N_A_686_74#_c_718_n N_VPWR_c_880_n 0.00505379f $X=5.545 $Y=1.635 $X2=0
+ $Y2=0
cc_507 N_A_686_74#_c_718_n N_VPWR_c_895_n 0.00408456f $X=5.545 $Y=1.635 $X2=0
+ $Y2=0
cc_508 N_A_686_74#_c_719_n N_VGND_c_1041_n 0.00375089f $X=5.59 $Y=1.22 $X2=0
+ $Y2=0
cc_509 N_A_686_74#_c_720_n N_VGND_c_1041_n 0.00320573f $X=5.455 $Y=1.385 $X2=0
+ $Y2=0
cc_510 N_A_686_74#_c_721_n N_VGND_c_1041_n 0.0197029f $X=4.375 $Y=0.485 $X2=0
+ $Y2=0
cc_511 N_A_686_74#_c_722_n N_VGND_c_1041_n 0.0196947f $X=5.005 $Y=1.385 $X2=0
+ $Y2=0
cc_512 N_A_686_74#_c_724_n N_VGND_c_1041_n 0.0284738f $X=4.55 $Y=1.22 $X2=0
+ $Y2=0
cc_513 N_A_686_74#_c_719_n N_VGND_c_1042_n 0.00250149f $X=5.59 $Y=1.22 $X2=0
+ $Y2=0
cc_514 N_A_686_74#_c_721_n N_VGND_c_1044_n 0.0458338f $X=4.375 $Y=0.485 $X2=0
+ $Y2=0
cc_515 N_A_686_74#_c_719_n N_VGND_c_1046_n 0.00461464f $X=5.59 $Y=1.22 $X2=0
+ $Y2=0
cc_516 N_A_686_74#_c_719_n N_VGND_c_1052_n 0.00914027f $X=5.59 $Y=1.22 $X2=0
+ $Y2=0
cc_517 N_A_686_74#_c_721_n N_VGND_c_1052_n 0.0405628f $X=4.375 $Y=0.485 $X2=0
+ $Y2=0
cc_518 N_A_686_74#_c_721_n N_VGND_c_1054_n 0.00836069f $X=4.375 $Y=0.485 $X2=0
+ $Y2=0
cc_519 N_A_686_74#_c_721_n A_841_118# 0.00447747f $X=4.375 $Y=0.485 $X2=-0.19
+ $Y2=-0.245
cc_520 N_A_686_74#_c_724_n A_841_118# 0.00388189f $X=4.55 $Y=1.22 $X2=-0.19
+ $Y2=-0.245
cc_521 N_RESET_B_c_812_n N_VPWR_c_883_n 0.00637166f $X=6.005 $Y=1.635 $X2=0
+ $Y2=0
cc_522 N_RESET_B_c_812_n N_VPWR_c_885_n 0.00475875f $X=6.005 $Y=1.635 $X2=0
+ $Y2=0
cc_523 N_RESET_B_c_812_n N_VPWR_c_880_n 0.00505379f $X=6.005 $Y=1.635 $X2=0
+ $Y2=0
cc_524 N_RESET_B_c_811_n N_VGND_c_1042_n 0.0164371f $X=5.98 $Y=1.22 $X2=0 $Y2=0
cc_525 N_RESET_B_c_812_n N_VGND_c_1042_n 0.00182516f $X=6.005 $Y=1.635 $X2=0
+ $Y2=0
cc_526 RESET_B N_VGND_c_1042_n 0.0102211f $X=5.915 $Y=1.21 $X2=0 $Y2=0
cc_527 N_RESET_B_c_811_n N_VGND_c_1046_n 0.00383152f $X=5.98 $Y=1.22 $X2=0 $Y2=0
cc_528 N_RESET_B_c_811_n N_VGND_c_1052_n 0.0075725f $X=5.98 $Y=1.22 $X2=0 $Y2=0
cc_529 N_A_1437_112#_c_843_n N_VPWR_c_884_n 0.00802746f $X=8.135 $Y=1.765 $X2=0
+ $Y2=0
cc_530 N_A_1437_112#_c_847_n N_VPWR_c_884_n 0.061164f $X=7.37 $Y=2.065 $X2=0
+ $Y2=0
cc_531 N_A_1437_112#_c_845_n N_VPWR_c_884_n 0.0210261f $X=8.06 $Y=1.465 $X2=0
+ $Y2=0
cc_532 N_A_1437_112#_c_847_n N_VPWR_c_890_n 0.00602538f $X=7.37 $Y=2.065 $X2=0
+ $Y2=0
cc_533 N_A_1437_112#_c_843_n N_VPWR_c_891_n 0.00445602f $X=8.135 $Y=1.765 $X2=0
+ $Y2=0
cc_534 N_A_1437_112#_c_843_n N_VPWR_c_880_n 0.00865549f $X=8.135 $Y=1.765 $X2=0
+ $Y2=0
cc_535 N_A_1437_112#_c_847_n N_VPWR_c_880_n 0.00799129f $X=7.37 $Y=2.065 $X2=0
+ $Y2=0
cc_536 N_A_1437_112#_c_847_n N_Q_c_989_n 0.0937326f $X=7.37 $Y=2.065 $X2=0 $Y2=0
cc_537 N_A_1437_112#_c_855_n N_Q_c_989_n 0.0253248f $X=7.422 $Y=1.465 $X2=0
+ $Y2=0
cc_538 N_A_1437_112#_c_844_n N_Q_c_990_n 0.0620552f $X=7.395 $Y=0.835 $X2=0
+ $Y2=0
cc_539 N_A_1437_112#_M1020_g N_Q_N_c_1022_n 0.0020582f $X=8.125 $Y=0.74 $X2=0
+ $Y2=0
cc_540 N_A_1437_112#_c_843_n Q_N 0.00332348f $X=8.135 $Y=1.765 $X2=0 $Y2=0
cc_541 N_A_1437_112#_c_843_n Q_N 0.0114556f $X=8.135 $Y=1.765 $X2=0 $Y2=0
cc_542 N_A_1437_112#_M1020_g N_Q_N_c_1024_n 0.00413599f $X=8.125 $Y=0.74 $X2=0
+ $Y2=0
cc_543 N_A_1437_112#_c_843_n N_Q_N_c_1024_n 0.0127956f $X=8.135 $Y=1.765 $X2=0
+ $Y2=0
cc_544 N_A_1437_112#_c_845_n N_Q_N_c_1024_n 0.0262113f $X=8.06 $Y=1.465 $X2=0
+ $Y2=0
cc_545 N_A_1437_112#_M1020_g N_VGND_c_1043_n 0.017651f $X=8.125 $Y=0.74 $X2=0
+ $Y2=0
cc_546 N_A_1437_112#_c_843_n N_VGND_c_1043_n 0.00361906f $X=8.135 $Y=1.765 $X2=0
+ $Y2=0
cc_547 N_A_1437_112#_c_844_n N_VGND_c_1043_n 0.0423984f $X=7.395 $Y=0.835 $X2=0
+ $Y2=0
cc_548 N_A_1437_112#_c_845_n N_VGND_c_1043_n 0.0281682f $X=8.06 $Y=1.465 $X2=0
+ $Y2=0
cc_549 N_A_1437_112#_c_844_n N_VGND_c_1050_n 0.00677257f $X=7.395 $Y=0.835 $X2=0
+ $Y2=0
cc_550 N_A_1437_112#_M1020_g N_VGND_c_1051_n 0.00383152f $X=8.125 $Y=0.74 $X2=0
+ $Y2=0
cc_551 N_A_1437_112#_M1020_g N_VGND_c_1052_n 0.00761264f $X=8.125 $Y=0.74 $X2=0
+ $Y2=0
cc_552 N_A_1437_112#_c_844_n N_VGND_c_1052_n 0.00885099f $X=7.395 $Y=0.835 $X2=0
+ $Y2=0
cc_553 N_VPWR_c_883_n Q 0.0257679f $X=6.28 $Y=2.145 $X2=0 $Y2=0
cc_554 N_VPWR_c_884_n Q 0.0023223f $X=7.91 $Y=1.985 $X2=0 $Y2=0
cc_555 N_VPWR_c_890_n Q 0.0123381f $X=7.745 $Y=3.33 $X2=0 $Y2=0
cc_556 N_VPWR_c_880_n Q 0.0143507f $X=8.4 $Y=3.33 $X2=0 $Y2=0
cc_557 N_VPWR_c_884_n Q_N 0.0421732f $X=7.91 $Y=1.985 $X2=0 $Y2=0
cc_558 N_VPWR_c_891_n Q_N 0.0148169f $X=8.4 $Y=3.33 $X2=0 $Y2=0
cc_559 N_VPWR_c_880_n Q_N 0.0122313f $X=8.4 $Y=3.33 $X2=0 $Y2=0
cc_560 N_Q_c_990_n N_VGND_c_1042_n 0.0461224f $X=6.735 $Y=0.515 $X2=0 $Y2=0
cc_561 N_Q_c_990_n N_VGND_c_1043_n 0.00656611f $X=6.735 $Y=0.515 $X2=0 $Y2=0
cc_562 N_Q_c_990_n N_VGND_c_1050_n 0.0244012f $X=6.735 $Y=0.515 $X2=0 $Y2=0
cc_563 N_Q_c_990_n N_VGND_c_1052_n 0.0201135f $X=6.735 $Y=0.515 $X2=0 $Y2=0
cc_564 N_Q_N_c_1022_n N_VGND_c_1043_n 0.0308138f $X=8.34 $Y=0.515 $X2=0 $Y2=0
cc_565 N_Q_N_c_1022_n N_VGND_c_1051_n 0.0126277f $X=8.34 $Y=0.515 $X2=0 $Y2=0
cc_566 N_Q_N_c_1022_n N_VGND_c_1052_n 0.0104521f $X=8.34 $Y=0.515 $X2=0 $Y2=0
