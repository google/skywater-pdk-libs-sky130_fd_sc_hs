* File: sky130_fd_sc_hs__xnor2_1.pxi.spice
* Created: Thu Aug 27 21:12:02 2020
* 
x_PM_SKY130_FD_SC_HS__XNOR2_1%B N_B_c_60_n N_B_M1005_g N_B_c_61_n N_B_M1004_g
+ N_B_c_62_n N_B_M1003_g N_B_M1009_g N_B_c_68_n N_B_c_80_p N_B_c_116_p
+ N_B_c_69_n N_B_c_64_n B N_B_c_65_n PM_SKY130_FD_SC_HS__XNOR2_1%B
x_PM_SKY130_FD_SC_HS__XNOR2_1%A N_A_M1008_g N_A_c_149_n N_A_M1001_g N_A_c_143_n
+ N_A_c_144_n N_A_c_145_n N_A_M1007_g N_A_M1000_g N_A_c_151_n A N_A_c_147_n
+ PM_SKY130_FD_SC_HS__XNOR2_1%A
x_PM_SKY130_FD_SC_HS__XNOR2_1%A_138_385# N_A_138_385#_M1005_d
+ N_A_138_385#_M1001_d N_A_138_385#_c_204_n N_A_138_385#_M1002_g
+ N_A_138_385#_M1006_g N_A_138_385#_c_206_n N_A_138_385#_c_207_n
+ N_A_138_385#_c_208_n N_A_138_385#_c_212_n N_A_138_385#_c_209_n
+ N_A_138_385#_c_210_n PM_SKY130_FD_SC_HS__XNOR2_1%A_138_385#
x_PM_SKY130_FD_SC_HS__XNOR2_1%VPWR N_VPWR_M1001_s N_VPWR_M1004_d N_VPWR_M1002_d
+ N_VPWR_c_287_n N_VPWR_c_288_n N_VPWR_c_289_n N_VPWR_c_290_n N_VPWR_c_291_n
+ N_VPWR_c_292_n N_VPWR_c_293_n VPWR N_VPWR_c_294_n N_VPWR_c_295_n
+ N_VPWR_c_296_n N_VPWR_c_286_n PM_SKY130_FD_SC_HS__XNOR2_1%VPWR
x_PM_SKY130_FD_SC_HS__XNOR2_1%Y N_Y_M1006_d N_Y_M1003_d N_Y_c_343_n N_Y_c_340_n
+ N_Y_c_337_n N_Y_c_338_n N_Y_c_339_n Y N_Y_c_342_n
+ PM_SKY130_FD_SC_HS__XNOR2_1%Y
x_PM_SKY130_FD_SC_HS__XNOR2_1%VGND N_VGND_M1008_s N_VGND_M1000_d N_VGND_c_371_n
+ N_VGND_c_372_n N_VGND_c_373_n VGND N_VGND_c_374_n N_VGND_c_375_n
+ N_VGND_c_376_n N_VGND_c_377_n PM_SKY130_FD_SC_HS__XNOR2_1%VGND
x_PM_SKY130_FD_SC_HS__XNOR2_1%A_293_74# N_A_293_74#_M1000_s N_A_293_74#_M1009_d
+ N_A_293_74#_c_410_n N_A_293_74#_c_409_n N_A_293_74#_c_413_n
+ PM_SKY130_FD_SC_HS__XNOR2_1%A_293_74#
cc_1 VNB N_B_c_60_n 0.0162445f $X=-0.19 $Y=-0.245 $X2=0.845 $Y2=1.31
cc_2 VNB N_B_c_61_n 0.0403496f $X=-0.19 $Y=-0.245 $X2=1.065 $Y2=1.85
cc_3 VNB N_B_c_62_n 0.0222957f $X=-0.19 $Y=-0.245 $X2=2.225 $Y2=1.765
cc_4 VNB N_B_M1009_g 0.0257826f $X=-0.19 $Y=-0.245 $X2=2.39 $Y2=0.74
cc_5 VNB N_B_c_64_n 0.0050024f $X=-0.19 $Y=-0.245 $X2=2.3 $Y2=1.515
cc_6 VNB N_B_c_65_n 0.00348558f $X=-0.19 $Y=-0.245 $X2=1.26 $Y2=1.607
cc_7 VNB N_A_M1008_g 0.0615073f $X=-0.19 $Y=-0.245 $X2=1.065 $Y2=1.85
cc_8 VNB N_A_c_143_n 0.10165f $X=-0.19 $Y=-0.245 $X2=2.225 $Y2=2.4
cc_9 VNB N_A_c_144_n 0.011606f $X=-0.19 $Y=-0.245 $X2=2.225 $Y2=2.4
cc_10 VNB N_A_c_145_n 0.0300955f $X=-0.19 $Y=-0.245 $X2=2.39 $Y2=1.35
cc_11 VNB N_A_M1000_g 0.0193389f $X=-0.19 $Y=-0.245 $X2=2.015 $Y2=2.035
cc_12 VNB N_A_c_147_n 0.00208705f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_138_385#_c_204_n 0.0343974f $X=-0.19 $Y=-0.245 $X2=2.225 $Y2=1.765
cc_14 VNB N_A_138_385#_M1006_g 0.0249763f $X=-0.19 $Y=-0.245 $X2=2.39 $Y2=0.74
cc_15 VNB N_A_138_385#_c_206_n 0.00745634f $X=-0.19 $Y=-0.245 $X2=2.1 $Y2=1.515
cc_16 VNB N_A_138_385#_c_207_n 0.0267453f $X=-0.19 $Y=-0.245 $X2=2.3 $Y2=1.515
cc_17 VNB N_A_138_385#_c_208_n 0.00354512f $X=-0.19 $Y=-0.245 $X2=2.3 $Y2=1.515
cc_18 VNB N_A_138_385#_c_209_n 0.00494238f $X=-0.19 $Y=-0.245 $X2=1.022 $Y2=1.6
cc_19 VNB N_A_138_385#_c_210_n 0.00608349f $X=-0.19 $Y=-0.245 $X2=1.11 $Y2=1.6
cc_20 VNB N_VPWR_c_286_n 0.143779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_Y_c_337_n 0.027697f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_Y_c_338_n 0.0247615f $X=-0.19 $Y=-0.245 $X2=2.015 $Y2=2.035
cc_23 VNB N_Y_c_339_n 0.0105427f $X=-0.19 $Y=-0.245 $X2=2.1 $Y2=1.95
cc_24 VNB N_VGND_c_371_n 0.0106846f $X=-0.19 $Y=-0.245 $X2=2.225 $Y2=1.765
cc_25 VNB N_VGND_c_372_n 0.0498887f $X=-0.19 $Y=-0.245 $X2=2.225 $Y2=2.4
cc_26 VNB N_VGND_c_373_n 0.00813052f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_VGND_c_374_n 0.0423941f $X=-0.19 $Y=-0.245 $X2=1.345 $Y2=2.035
cc_28 VNB N_VGND_c_375_n 0.0320561f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_376_n 0.196578f $X=-0.19 $Y=-0.245 $X2=1.022 $Y2=1.6
cc_30 VNB N_VGND_c_377_n 0.00631651f $X=-0.19 $Y=-0.245 $X2=1.2 $Y2=1.607
cc_31 VNB N_A_293_74#_c_409_n 0.00381723f $X=-0.19 $Y=-0.245 $X2=2.39 $Y2=1.35
cc_32 VPB N_B_c_61_n 0.0350078f $X=-0.19 $Y=1.66 $X2=1.065 $Y2=1.85
cc_33 VPB N_B_c_62_n 0.0272375f $X=-0.19 $Y=1.66 $X2=2.225 $Y2=1.765
cc_34 VPB N_B_c_68_n 0.00300914f $X=-0.19 $Y=1.66 $X2=1.26 $Y2=1.95
cc_35 VPB N_B_c_69_n 0.00145233f $X=-0.19 $Y=1.66 $X2=2.1 $Y2=1.95
cc_36 VPB N_B_c_64_n 6.49643e-19 $X=-0.19 $Y=1.66 $X2=2.3 $Y2=1.515
cc_37 VPB N_B_c_65_n 0.00310283f $X=-0.19 $Y=1.66 $X2=1.26 $Y2=1.607
cc_38 VPB N_A_M1008_g 0.00332562f $X=-0.19 $Y=1.66 $X2=1.065 $Y2=1.85
cc_39 VPB N_A_c_149_n 0.0169138f $X=-0.19 $Y=1.66 $X2=1.065 $Y2=2.345
cc_40 VPB N_A_c_145_n 0.0303831f $X=-0.19 $Y=1.66 $X2=2.39 $Y2=1.35
cc_41 VPB N_A_c_151_n 0.0247479f $X=-0.19 $Y=1.66 $X2=2.1 $Y2=1.95
cc_42 VPB N_A_c_147_n 0.0026218f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_43 VPB N_A_138_385#_c_204_n 0.0260147f $X=-0.19 $Y=1.66 $X2=2.225 $Y2=1.765
cc_44 VPB N_A_138_385#_c_212_n 0.00351449f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_45 VPB N_A_138_385#_c_209_n 0.0020675f $X=-0.19 $Y=1.66 $X2=1.022 $Y2=1.6
cc_46 VPB N_VPWR_c_287_n 0.0185202f $X=-0.19 $Y=1.66 $X2=2.39 $Y2=0.74
cc_47 VPB N_VPWR_c_288_n 0.00626527f $X=-0.19 $Y=1.66 $X2=1.26 $Y2=1.78
cc_48 VPB N_VPWR_c_289_n 0.0141048f $X=-0.19 $Y=1.66 $X2=1.26 $Y2=1.95
cc_49 VPB N_VPWR_c_290_n 0.041775f $X=-0.19 $Y=1.66 $X2=1.345 $Y2=2.035
cc_50 VPB N_VPWR_c_291_n 0.0140747f $X=-0.19 $Y=1.66 $X2=2.1 $Y2=1.515
cc_51 VPB N_VPWR_c_292_n 0.0139245f $X=-0.19 $Y=1.66 $X2=2.3 $Y2=1.515
cc_52 VPB N_VPWR_c_293_n 0.0395112f $X=-0.19 $Y=1.66 $X2=1.115 $Y2=1.58
cc_53 VPB N_VPWR_c_294_n 0.0271489f $X=-0.19 $Y=1.66 $X2=2.3 $Y2=1.515
cc_54 VPB N_VPWR_c_295_n 0.0299529f $X=-0.19 $Y=1.66 $X2=1.26 $Y2=1.607
cc_55 VPB N_VPWR_c_296_n 0.00614127f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_56 VPB N_VPWR_c_286_n 0.0826623f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_57 VPB N_Y_c_340_n 0.0114589f $X=-0.19 $Y=1.66 $X2=2.225 $Y2=2.4
cc_58 VPB N_Y_c_338_n 0.00939981f $X=-0.19 $Y=1.66 $X2=2.015 $Y2=2.035
cc_59 VPB N_Y_c_342_n 0.00459573f $X=-0.19 $Y=1.66 $X2=1.115 $Y2=1.58
cc_60 N_B_c_60_n N_A_M1008_g 0.0574491f $X=0.845 $Y=1.31 $X2=0 $Y2=0
cc_61 N_B_c_61_n N_A_M1008_g 0.00613719f $X=1.065 $Y=1.85 $X2=0 $Y2=0
cc_62 N_B_c_61_n N_A_c_149_n 0.0131595f $X=1.065 $Y=1.85 $X2=0 $Y2=0
cc_63 N_B_c_60_n N_A_c_143_n 0.0103003f $X=0.845 $Y=1.31 $X2=0 $Y2=0
cc_64 N_B_M1009_g N_A_c_143_n 0.0302512f $X=2.39 $Y=0.74 $X2=0 $Y2=0
cc_65 N_B_c_61_n N_A_c_145_n 0.0319744f $X=1.065 $Y=1.85 $X2=0 $Y2=0
cc_66 N_B_c_62_n N_A_c_145_n 0.0802925f $X=2.225 $Y=1.765 $X2=0 $Y2=0
cc_67 N_B_c_68_n N_A_c_145_n 0.00154773f $X=1.26 $Y=1.95 $X2=0 $Y2=0
cc_68 N_B_c_80_p N_A_c_145_n 0.0177621f $X=2.015 $Y=2.035 $X2=0 $Y2=0
cc_69 N_B_c_69_n N_A_c_145_n 0.00244625f $X=2.1 $Y=1.95 $X2=0 $Y2=0
cc_70 N_B_c_64_n N_A_c_145_n 0.0022979f $X=2.3 $Y=1.515 $X2=0 $Y2=0
cc_71 N_B_c_65_n N_A_c_145_n 0.00178335f $X=1.26 $Y=1.607 $X2=0 $Y2=0
cc_72 N_B_c_61_n N_A_c_151_n 0.00732589f $X=1.065 $Y=1.85 $X2=0 $Y2=0
cc_73 N_B_c_61_n N_A_c_147_n 0.00121542f $X=1.065 $Y=1.85 $X2=0 $Y2=0
cc_74 N_B_c_62_n N_A_c_147_n 4.00099e-19 $X=2.225 $Y=1.765 $X2=0 $Y2=0
cc_75 N_B_c_80_p N_A_c_147_n 0.0234061f $X=2.015 $Y=2.035 $X2=0 $Y2=0
cc_76 N_B_c_69_n N_A_c_147_n 0.00747766f $X=2.1 $Y=1.95 $X2=0 $Y2=0
cc_77 N_B_c_64_n N_A_c_147_n 0.0267388f $X=2.3 $Y=1.515 $X2=0 $Y2=0
cc_78 N_B_c_65_n N_A_c_147_n 0.028107f $X=1.26 $Y=1.607 $X2=0 $Y2=0
cc_79 N_B_c_62_n N_A_138_385#_c_204_n 0.0355782f $X=2.225 $Y=1.765 $X2=0 $Y2=0
cc_80 N_B_M1009_g N_A_138_385#_c_204_n 0.0210954f $X=2.39 $Y=0.74 $X2=0 $Y2=0
cc_81 N_B_c_69_n N_A_138_385#_c_204_n 8.64876e-19 $X=2.1 $Y=1.95 $X2=0 $Y2=0
cc_82 N_B_c_64_n N_A_138_385#_c_204_n 5.22561e-19 $X=2.3 $Y=1.515 $X2=0 $Y2=0
cc_83 N_B_M1009_g N_A_138_385#_M1006_g 0.0296051f $X=2.39 $Y=0.74 $X2=0 $Y2=0
cc_84 N_B_c_60_n N_A_138_385#_c_206_n 0.00760958f $X=0.845 $Y=1.31 $X2=0 $Y2=0
cc_85 N_B_c_61_n N_A_138_385#_c_207_n 0.00130476f $X=1.065 $Y=1.85 $X2=0 $Y2=0
cc_86 N_B_c_62_n N_A_138_385#_c_207_n 0.00465926f $X=2.225 $Y=1.765 $X2=0 $Y2=0
cc_87 N_B_M1009_g N_A_138_385#_c_207_n 0.0111001f $X=2.39 $Y=0.74 $X2=0 $Y2=0
cc_88 N_B_c_64_n N_A_138_385#_c_207_n 0.0337543f $X=2.3 $Y=1.515 $X2=0 $Y2=0
cc_89 N_B_c_65_n N_A_138_385#_c_207_n 0.00695518f $X=1.26 $Y=1.607 $X2=0 $Y2=0
cc_90 N_B_c_60_n N_A_138_385#_c_208_n 0.0161471f $X=0.845 $Y=1.31 $X2=0 $Y2=0
cc_91 N_B_c_61_n N_A_138_385#_c_208_n 0.00963497f $X=1.065 $Y=1.85 $X2=0 $Y2=0
cc_92 N_B_c_65_n N_A_138_385#_c_208_n 0.0226832f $X=1.26 $Y=1.607 $X2=0 $Y2=0
cc_93 N_B_c_61_n N_A_138_385#_c_212_n 0.024424f $X=1.065 $Y=1.85 $X2=0 $Y2=0
cc_94 N_B_c_65_n N_A_138_385#_c_212_n 0.00291112f $X=1.26 $Y=1.607 $X2=0 $Y2=0
cc_95 N_B_c_60_n N_A_138_385#_c_209_n 3.17485e-19 $X=0.845 $Y=1.31 $X2=0 $Y2=0
cc_96 N_B_c_61_n N_A_138_385#_c_209_n 0.00854012f $X=1.065 $Y=1.85 $X2=0 $Y2=0
cc_97 N_B_c_68_n N_A_138_385#_c_209_n 0.00497997f $X=1.26 $Y=1.95 $X2=0 $Y2=0
cc_98 N_B_c_65_n N_A_138_385#_c_209_n 0.0262595f $X=1.26 $Y=1.607 $X2=0 $Y2=0
cc_99 N_B_c_62_n N_A_138_385#_c_210_n 9.00083e-19 $X=2.225 $Y=1.765 $X2=0 $Y2=0
cc_100 N_B_M1009_g N_A_138_385#_c_210_n 0.00363004f $X=2.39 $Y=0.74 $X2=0 $Y2=0
cc_101 N_B_c_64_n N_A_138_385#_c_210_n 0.0226425f $X=2.3 $Y=1.515 $X2=0 $Y2=0
cc_102 N_B_c_68_n N_VPWR_M1004_d 3.73937e-19 $X=1.26 $Y=1.95 $X2=0 $Y2=0
cc_103 N_B_c_80_p N_VPWR_M1004_d 0.0151476f $X=2.015 $Y=2.035 $X2=0 $Y2=0
cc_104 N_B_c_116_p N_VPWR_M1004_d 0.00742686f $X=1.345 $Y=2.035 $X2=0 $Y2=0
cc_105 N_B_c_61_n N_VPWR_c_291_n 0.00739883f $X=1.065 $Y=1.85 $X2=0 $Y2=0
cc_106 N_B_c_62_n N_VPWR_c_291_n 0.0011771f $X=2.225 $Y=1.765 $X2=0 $Y2=0
cc_107 N_B_c_80_p N_VPWR_c_291_n 0.0219335f $X=2.015 $Y=2.035 $X2=0 $Y2=0
cc_108 N_B_c_62_n N_VPWR_c_293_n 9.74585e-19 $X=2.225 $Y=1.765 $X2=0 $Y2=0
cc_109 N_B_c_61_n N_VPWR_c_294_n 0.00438163f $X=1.065 $Y=1.85 $X2=0 $Y2=0
cc_110 N_B_c_62_n N_VPWR_c_295_n 0.00291649f $X=2.225 $Y=1.765 $X2=0 $Y2=0
cc_111 N_B_c_61_n N_VPWR_c_286_n 0.00486331f $X=1.065 $Y=1.85 $X2=0 $Y2=0
cc_112 N_B_c_62_n N_VPWR_c_286_n 0.00360376f $X=2.225 $Y=1.765 $X2=0 $Y2=0
cc_113 N_B_c_80_p A_376_368# 0.00764317f $X=2.015 $Y=2.035 $X2=-0.19 $Y2=-0.245
cc_114 N_B_c_69_n A_376_368# 0.00150831f $X=2.1 $Y=1.95 $X2=-0.19 $Y2=-0.245
cc_115 N_B_c_62_n N_Y_c_343_n 0.00295532f $X=2.225 $Y=1.765 $X2=0 $Y2=0
cc_116 N_B_c_64_n N_Y_c_343_n 0.00869105f $X=2.3 $Y=1.515 $X2=0 $Y2=0
cc_117 N_B_c_64_n N_Y_c_338_n 0.00136308f $X=2.3 $Y=1.515 $X2=0 $Y2=0
cc_118 N_B_c_62_n N_Y_c_342_n 0.0297741f $X=2.225 $Y=1.765 $X2=0 $Y2=0
cc_119 N_B_c_80_p N_Y_c_342_n 0.0069951f $X=2.015 $Y=2.035 $X2=0 $Y2=0
cc_120 N_B_c_64_n N_Y_c_342_n 0.00390307f $X=2.3 $Y=1.515 $X2=0 $Y2=0
cc_121 N_B_c_60_n N_VGND_c_372_n 0.00207013f $X=0.845 $Y=1.31 $X2=0 $Y2=0
cc_122 N_B_M1009_g N_VGND_c_373_n 0.00452091f $X=2.39 $Y=0.74 $X2=0 $Y2=0
cc_123 N_B_M1009_g N_VGND_c_375_n 0.00327917f $X=2.39 $Y=0.74 $X2=0 $Y2=0
cc_124 N_B_c_60_n N_VGND_c_376_n 9.39239e-19 $X=0.845 $Y=1.31 $X2=0 $Y2=0
cc_125 N_B_M1009_g N_VGND_c_376_n 0.00415199f $X=2.39 $Y=0.74 $X2=0 $Y2=0
cc_126 N_B_M1009_g N_A_293_74#_c_410_n 0.00969414f $X=2.39 $Y=0.74 $X2=0 $Y2=0
cc_127 N_B_c_60_n N_A_293_74#_c_409_n 0.00216277f $X=0.845 $Y=1.31 $X2=0 $Y2=0
cc_128 N_B_M1009_g N_A_293_74#_c_409_n 5.82005e-19 $X=2.39 $Y=0.74 $X2=0 $Y2=0
cc_129 N_B_M1009_g N_A_293_74#_c_413_n 0.00488999f $X=2.39 $Y=0.74 $X2=0 $Y2=0
cc_130 N_A_M1008_g N_A_138_385#_c_206_n 0.00118315f $X=0.485 $Y=0.915 $X2=0
+ $Y2=0
cc_131 N_A_c_143_n N_A_138_385#_c_206_n 0.00622038f $X=1.74 $Y=0.18 $X2=0 $Y2=0
cc_132 N_A_M1000_g N_A_138_385#_c_206_n 0.0040271f $X=1.815 $Y=0.74 $X2=0 $Y2=0
cc_133 N_A_c_145_n N_A_138_385#_c_207_n 0.00177098f $X=1.805 $Y=1.765 $X2=0
+ $Y2=0
cc_134 N_A_M1000_g N_A_138_385#_c_207_n 0.0145692f $X=1.815 $Y=0.74 $X2=0 $Y2=0
cc_135 N_A_c_147_n N_A_138_385#_c_207_n 0.0248926f $X=1.68 $Y=1.515 $X2=0 $Y2=0
cc_136 N_A_M1008_g N_A_138_385#_c_208_n 8.41489e-19 $X=0.485 $Y=0.915 $X2=0
+ $Y2=0
cc_137 N_A_M1000_g N_A_138_385#_c_208_n 0.00210586f $X=1.815 $Y=0.74 $X2=0 $Y2=0
cc_138 N_A_c_149_n N_A_138_385#_c_212_n 0.0149566f $X=0.615 $Y=1.85 $X2=0 $Y2=0
cc_139 N_A_M1008_g N_A_138_385#_c_209_n 0.0112389f $X=0.485 $Y=0.915 $X2=0 $Y2=0
cc_140 N_A_c_149_n N_A_138_385#_c_209_n 0.00372929f $X=0.615 $Y=1.85 $X2=0 $Y2=0
cc_141 N_A_c_151_n N_A_138_385#_c_209_n 0.0106014f $X=0.615 $Y=1.775 $X2=0 $Y2=0
cc_142 N_A_c_149_n N_VPWR_c_287_n 0.00815516f $X=0.615 $Y=1.85 $X2=0 $Y2=0
cc_143 N_A_c_151_n N_VPWR_c_287_n 5.52212e-19 $X=0.615 $Y=1.775 $X2=0 $Y2=0
cc_144 N_A_c_151_n N_VPWR_c_288_n 0.00249294f $X=0.615 $Y=1.775 $X2=0 $Y2=0
cc_145 N_A_c_149_n N_VPWR_c_290_n 0.0144862f $X=0.615 $Y=1.85 $X2=0 $Y2=0
cc_146 N_A_c_145_n N_VPWR_c_291_n 0.0136884f $X=1.805 $Y=1.765 $X2=0 $Y2=0
cc_147 N_A_c_149_n N_VPWR_c_294_n 0.00438163f $X=0.615 $Y=1.85 $X2=0 $Y2=0
cc_148 N_A_c_145_n N_VPWR_c_295_n 0.00413917f $X=1.805 $Y=1.765 $X2=0 $Y2=0
cc_149 N_A_c_149_n N_VPWR_c_286_n 0.00486331f $X=0.615 $Y=1.85 $X2=0 $Y2=0
cc_150 N_A_c_145_n N_VPWR_c_286_n 0.00817532f $X=1.805 $Y=1.765 $X2=0 $Y2=0
cc_151 N_A_c_145_n N_Y_c_342_n 0.00570246f $X=1.805 $Y=1.765 $X2=0 $Y2=0
cc_152 N_A_M1008_g N_VGND_c_372_n 0.0288731f $X=0.485 $Y=0.915 $X2=0 $Y2=0
cc_153 N_A_c_144_n N_VGND_c_372_n 0.00763335f $X=0.56 $Y=0.18 $X2=0 $Y2=0
cc_154 N_A_c_143_n N_VGND_c_373_n 0.0100525f $X=1.74 $Y=0.18 $X2=0 $Y2=0
cc_155 N_A_c_144_n N_VGND_c_374_n 0.0440575f $X=0.56 $Y=0.18 $X2=0 $Y2=0
cc_156 N_A_c_143_n N_VGND_c_376_n 0.0504593f $X=1.74 $Y=0.18 $X2=0 $Y2=0
cc_157 N_A_c_144_n N_VGND_c_376_n 0.00749832f $X=0.56 $Y=0.18 $X2=0 $Y2=0
cc_158 N_A_M1000_g N_A_293_74#_c_410_n 0.00987582f $X=1.815 $Y=0.74 $X2=0 $Y2=0
cc_159 N_A_c_143_n N_A_293_74#_c_409_n 0.00435764f $X=1.74 $Y=0.18 $X2=0 $Y2=0
cc_160 N_A_M1000_g N_A_293_74#_c_409_n 0.00493339f $X=1.815 $Y=0.74 $X2=0 $Y2=0
cc_161 N_A_M1000_g N_A_293_74#_c_413_n 5.82005e-19 $X=1.815 $Y=0.74 $X2=0 $Y2=0
cc_162 N_A_138_385#_c_212_n N_VPWR_c_287_n 0.00955207f $X=0.84 $Y=2.115 $X2=0
+ $Y2=0
cc_163 N_A_138_385#_c_209_n N_VPWR_c_287_n 0.0159937f $X=0.805 $Y=1.95 $X2=0
+ $Y2=0
cc_164 N_A_138_385#_c_212_n N_VPWR_c_290_n 0.0193641f $X=0.84 $Y=2.115 $X2=0
+ $Y2=0
cc_165 N_A_138_385#_c_212_n N_VPWR_c_291_n 0.019538f $X=0.84 $Y=2.115 $X2=0
+ $Y2=0
cc_166 N_A_138_385#_c_204_n N_VPWR_c_293_n 0.01542f $X=2.795 $Y=1.765 $X2=0
+ $Y2=0
cc_167 N_A_138_385#_c_212_n N_VPWR_c_294_n 0.00804153f $X=0.84 $Y=2.115 $X2=0
+ $Y2=0
cc_168 N_A_138_385#_c_204_n N_VPWR_c_295_n 0.00413917f $X=2.795 $Y=1.765 $X2=0
+ $Y2=0
cc_169 N_A_138_385#_c_204_n N_VPWR_c_286_n 0.00818781f $X=2.795 $Y=1.765 $X2=0
+ $Y2=0
cc_170 N_A_138_385#_c_212_n N_VPWR_c_286_n 0.0105967f $X=0.84 $Y=2.115 $X2=0
+ $Y2=0
cc_171 N_A_138_385#_c_207_n N_Y_c_343_n 0.00498172f $X=2.635 $Y=1.095 $X2=0
+ $Y2=0
cc_172 N_A_138_385#_c_210_n N_Y_c_343_n 0.00285479f $X=2.785 $Y=1.095 $X2=0
+ $Y2=0
cc_173 N_A_138_385#_c_204_n N_Y_c_340_n 0.0196526f $X=2.795 $Y=1.765 $X2=0 $Y2=0
cc_174 N_A_138_385#_c_210_n N_Y_c_340_n 0.0124313f $X=2.785 $Y=1.095 $X2=0 $Y2=0
cc_175 N_A_138_385#_M1006_g N_Y_c_337_n 0.0105687f $X=2.82 $Y=0.74 $X2=0 $Y2=0
cc_176 N_A_138_385#_c_204_n N_Y_c_338_n 0.014688f $X=2.795 $Y=1.765 $X2=0 $Y2=0
cc_177 N_A_138_385#_M1006_g N_Y_c_338_n 0.00330707f $X=2.82 $Y=0.74 $X2=0 $Y2=0
cc_178 N_A_138_385#_c_210_n N_Y_c_338_n 0.0329445f $X=2.785 $Y=1.095 $X2=0 $Y2=0
cc_179 N_A_138_385#_c_204_n N_Y_c_339_n 0.0012888f $X=2.795 $Y=1.765 $X2=0 $Y2=0
cc_180 N_A_138_385#_c_210_n N_Y_c_339_n 0.00984957f $X=2.785 $Y=1.095 $X2=0
+ $Y2=0
cc_181 N_A_138_385#_c_204_n N_Y_c_342_n 0.0043432f $X=2.795 $Y=1.765 $X2=0 $Y2=0
cc_182 N_A_138_385#_c_207_n N_VGND_M1000_d 0.00367023f $X=2.635 $Y=1.095 $X2=0
+ $Y2=0
cc_183 N_A_138_385#_c_206_n N_VGND_c_372_n 0.0145372f $X=1.06 $Y=0.74 $X2=0
+ $Y2=0
cc_184 N_A_138_385#_c_208_n N_VGND_c_372_n 0.00994413f $X=1.225 $Y=1.095 $X2=0
+ $Y2=0
cc_185 N_A_138_385#_c_206_n N_VGND_c_374_n 0.00749462f $X=1.06 $Y=0.74 $X2=0
+ $Y2=0
cc_186 N_A_138_385#_M1006_g N_VGND_c_375_n 0.00437532f $X=2.82 $Y=0.74 $X2=0
+ $Y2=0
cc_187 N_A_138_385#_M1006_g N_VGND_c_376_n 0.00829339f $X=2.82 $Y=0.74 $X2=0
+ $Y2=0
cc_188 N_A_138_385#_c_206_n N_VGND_c_376_n 0.00907254f $X=1.06 $Y=0.74 $X2=0
+ $Y2=0
cc_189 N_A_138_385#_c_208_n A_112_119# 0.00433061f $X=1.225 $Y=1.095 $X2=-0.19
+ $Y2=-0.245
cc_190 N_A_138_385#_c_207_n N_A_293_74#_M1000_s 0.00283795f $X=2.635 $Y=1.095
+ $X2=-0.19 $Y2=-0.245
cc_191 N_A_138_385#_c_207_n N_A_293_74#_M1009_d 0.00119058f $X=2.635 $Y=1.095
+ $X2=0 $Y2=0
cc_192 N_A_138_385#_c_210_n N_A_293_74#_M1009_d 5.84861e-19 $X=2.785 $Y=1.095
+ $X2=0 $Y2=0
cc_193 N_A_138_385#_c_207_n N_A_293_74#_c_410_n 0.039534f $X=2.635 $Y=1.095
+ $X2=0 $Y2=0
cc_194 N_A_138_385#_c_206_n N_A_293_74#_c_409_n 0.0190291f $X=1.06 $Y=0.74 $X2=0
+ $Y2=0
cc_195 N_A_138_385#_c_207_n N_A_293_74#_c_409_n 0.0207364f $X=2.635 $Y=1.095
+ $X2=0 $Y2=0
cc_196 N_A_138_385#_M1006_g N_A_293_74#_c_413_n 0.00452712f $X=2.82 $Y=0.74
+ $X2=0 $Y2=0
cc_197 N_A_138_385#_c_207_n N_A_293_74#_c_413_n 0.0103265f $X=2.635 $Y=1.095
+ $X2=0 $Y2=0
cc_198 N_A_138_385#_c_210_n N_A_293_74#_c_413_n 0.00637681f $X=2.785 $Y=1.095
+ $X2=0 $Y2=0
cc_199 N_VPWR_M1002_d N_Y_c_340_n 0.00829565f $X=2.87 $Y=1.84 $X2=0 $Y2=0
cc_200 N_VPWR_c_293_n N_Y_c_340_n 0.0226146f $X=3.02 $Y=2.3 $X2=0 $Y2=0
cc_201 N_VPWR_c_291_n N_Y_c_342_n 0.0365779f $X=1.58 $Y=2.415 $X2=0 $Y2=0
cc_202 N_VPWR_c_293_n N_Y_c_342_n 0.0267695f $X=3.02 $Y=2.3 $X2=0 $Y2=0
cc_203 N_VPWR_c_295_n N_Y_c_342_n 0.0280192f $X=2.855 $Y=3.33 $X2=0 $Y2=0
cc_204 N_VPWR_c_286_n N_Y_c_342_n 0.0229087f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_205 N_VPWR_c_287_n N_VGND_c_372_n 0.00899431f $X=0.34 $Y=2.07 $X2=0 $Y2=0
cc_206 A_376_368# N_Y_c_342_n 0.00786584f $X=1.88 $Y=1.84 $X2=1.115 $Y2=1.58
cc_207 N_Y_c_337_n N_VGND_c_375_n 0.013297f $X=3.06 $Y=0.515 $X2=0 $Y2=0
cc_208 N_Y_c_337_n N_VGND_c_376_n 0.0110061f $X=3.06 $Y=0.515 $X2=0 $Y2=0
cc_209 N_Y_c_337_n N_A_293_74#_c_413_n 0.0220168f $X=3.06 $Y=0.515 $X2=0 $Y2=0
cc_210 N_VGND_M1000_d N_A_293_74#_c_410_n 0.00697375f $X=1.89 $Y=0.37 $X2=0
+ $Y2=0
cc_211 N_VGND_c_373_n N_A_293_74#_c_410_n 0.0239631f $X=2.1 $Y=0.37 $X2=0 $Y2=0
cc_212 N_VGND_c_374_n N_A_293_74#_c_410_n 0.00227739f $X=1.935 $Y=0 $X2=0 $Y2=0
cc_213 N_VGND_c_375_n N_A_293_74#_c_410_n 0.00232204f $X=3.12 $Y=0 $X2=0 $Y2=0
cc_214 N_VGND_c_376_n N_A_293_74#_c_410_n 0.00980247f $X=3.12 $Y=0 $X2=0 $Y2=0
cc_215 N_VGND_c_374_n N_A_293_74#_c_409_n 0.00745853f $X=1.935 $Y=0 $X2=0 $Y2=0
cc_216 N_VGND_c_376_n N_A_293_74#_c_409_n 0.00921561f $X=3.12 $Y=0 $X2=0 $Y2=0
cc_217 N_VGND_c_375_n N_A_293_74#_c_413_n 0.00677194f $X=3.12 $Y=0 $X2=0 $Y2=0
cc_218 N_VGND_c_376_n N_A_293_74#_c_413_n 0.0103183f $X=3.12 $Y=0 $X2=0 $Y2=0
