* File: sky130_fd_sc_hs__a32o_2.spice
* Created: Tue Sep  1 19:53:30 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hs__a32o_2.pex.spice"
.subckt sky130_fd_sc_hs__a32o_2  VNB VPB A3 A2 A1 B1 B2 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* B2	B2
* B1	B1
* A1	A1
* A2	A2
* A3	A3
* VPB	VPB
* VNB	VNB
MM1003 N_VGND_M1003_d N_A_45_264#_M1003_g N_X_M1003_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.259 AS=0.1073 PD=2.18 PS=1.03 NRD=10.536 NRS=0.804 M=1 R=4.93333
+ SA=75000.3 SB=75003.4 A=0.111 P=1.78 MULT=1
MM1012 N_VGND_M1012_d N_A_45_264#_M1012_g N_X_M1003_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.2035 AS=0.1073 PD=1.29 PS=1.03 NRD=21.888 NRS=0.804 M=1 R=4.93333
+ SA=75000.7 SB=75003 A=0.111 P=1.78 MULT=1
MM1008 A_355_74# N_A3_M1008_g N_VGND_M1012_d VNB NLOWVT L=0.15 W=0.74 AD=0.0888
+ AS=0.2035 PD=0.98 PS=1.29 NRD=10.536 NRS=21.888 M=1 R=4.93333 SA=75001.4
+ SB=75002.3 A=0.111 P=1.78 MULT=1
MM1007 A_433_74# N_A2_M1007_g A_355_74# VNB NLOWVT L=0.15 W=0.74 AD=0.1554
+ AS=0.0888 PD=1.16 PS=0.98 NRD=25.128 NRS=10.536 M=1 R=4.93333 SA=75001.8
+ SB=75001.9 A=0.111 P=1.78 MULT=1
MM1013 N_A_45_264#_M1013_d N_A1_M1013_g A_433_74# VNB NLOWVT L=0.15 W=0.74
+ AD=0.1554 AS=0.1554 PD=1.16 PS=1.16 NRD=10.536 NRS=25.128 M=1 R=4.93333
+ SA=75002.4 SB=75001.4 A=0.111 P=1.78 MULT=1
MM1001 A_661_74# N_B1_M1001_g N_A_45_264#_M1013_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.1554 AS=0.1554 PD=1.16 PS=1.16 NRD=25.128 NRS=12.156 M=1 R=4.93333
+ SA=75002.9 SB=75000.8 A=0.111 P=1.78 MULT=1
MM1009 N_VGND_M1009_d N_B2_M1009_g A_661_74# VNB NLOWVT L=0.15 W=0.74 AD=0.2109
+ AS=0.1554 PD=2.05 PS=1.16 NRD=0 NRS=25.128 M=1 R=4.93333 SA=75003.5 SB=75000.2
+ A=0.111 P=1.78 MULT=1
MM1010 N_VPWR_M1010_d N_A_45_264#_M1010_g N_X_M1010_s VPB PSHORT L=0.15 W=1.12
+ AD=0.3304 AS=0.168 PD=2.83 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75003.2 A=0.168 P=2.54 MULT=1
MM1011 N_VPWR_M1011_d N_A_45_264#_M1011_g N_X_M1010_s VPB PSHORT L=0.15 W=1.12
+ AD=0.319728 AS=0.168 PD=1.76453 PS=1.42 NRD=23.7385 NRS=1.7533 M=1 R=7.46667
+ SA=75000.7 SB=75002.8 A=0.168 P=2.54 MULT=1
MM1000 N_A_346_368#_M1000_d N_A3_M1000_g N_VPWR_M1011_d VPB PSHORT L=0.15 W=1
+ AD=0.15 AS=0.285472 PD=1.3 PS=1.57547 NRD=1.9503 NRS=27.5603 M=1 R=6.66667
+ SA=75001.4 SB=75002.4 A=0.15 P=2.3 MULT=1
MM1002 N_VPWR_M1002_d N_A2_M1002_g N_A_346_368#_M1000_d VPB PSHORT L=0.15 W=1
+ AD=0.28 AS=0.15 PD=1.56 PS=1.3 NRD=27.5603 NRS=1.9503 M=1 R=6.66667 SA=75001.8
+ SB=75001.9 A=0.15 P=2.3 MULT=1
MM1005 N_A_346_368#_M1005_d N_A1_M1005_g N_VPWR_M1002_d VPB PSHORT L=0.15 W=1
+ AD=0.15 AS=0.28 PD=1.3 PS=1.56 NRD=1.9503 NRS=27.5603 M=1 R=6.66667 SA=75002.5
+ SB=75001.2 A=0.15 P=2.3 MULT=1
MM1006 N_A_45_264#_M1006_d N_B1_M1006_g N_A_346_368#_M1005_d VPB PSHORT L=0.15
+ W=1 AD=0.2 AS=0.15 PD=1.4 PS=1.3 NRD=11.8003 NRS=1.9503 M=1 R=6.66667 SA=75003
+ SB=75000.8 A=0.15 P=2.3 MULT=1
MM1004 N_A_346_368#_M1004_d N_B2_M1004_g N_A_45_264#_M1006_d VPB PSHORT L=0.15
+ W=1 AD=0.295 AS=0.2 PD=2.59 PS=1.4 NRD=1.9503 NRS=11.8003 M=1 R=6.66667
+ SA=75003.5 SB=75000.2 A=0.15 P=2.3 MULT=1
DX14_noxref VNB VPB NWDIODE A=8.742 P=13.12
*
.include "sky130_fd_sc_hs__a32o_2.pxi.spice"
*
.ends
*
*
