# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_hs__xor2_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__xor2_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  8.640000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  1.638000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.440000 1.420000 1.110000 1.750000 ;
        RECT 0.515000 0.580000 1.445000 0.600000 ;
        RECT 0.515000 0.600000 3.040000 0.750000 ;
        RECT 0.515000 0.750000 0.685000 1.420000 ;
        RECT 1.275000 0.750000 3.040000 0.770000 ;
        RECT 2.870000 0.770000 3.040000 1.020000 ;
        RECT 2.870000 1.020000 3.935000 1.190000 ;
        RECT 3.765000 1.190000 3.935000 1.350000 ;
        RECT 3.765000 1.350000 5.635000 1.520000 ;
        RECT 3.965000 1.520000 5.635000 1.775000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  1.638000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.030000 1.470000 2.360000 1.850000 ;
        RECT 2.030000 1.850000 3.655000 1.945000 ;
        RECT 2.030000 1.945000 5.975000 2.020000 ;
        RECT 3.485000 2.020000 5.975000 2.115000 ;
        RECT 5.805000 1.550000 8.165000 1.780000 ;
        RECT 5.805000 1.780000 5.975000 1.945000 ;
        RECT 5.885000 1.350000 8.165000 1.550000 ;
    END
  END B
  PIN X
    ANTENNADIFFAREA  1.504500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.985000 2.190000 3.315000 2.285000 ;
        RECT 2.985000 2.285000 6.315000 2.455000 ;
        RECT 2.985000 2.455000 3.315000 2.735000 ;
        RECT 3.210000 0.470000 3.540000 0.680000 ;
        RECT 3.210000 0.680000 4.275000 0.850000 ;
        RECT 3.885000 2.455000 4.215000 2.735000 ;
        RECT 4.105000 0.850000 4.275000 1.010000 ;
        RECT 4.105000 1.010000 8.505000 1.180000 ;
        RECT 6.145000 1.950000 8.505000 2.120000 ;
        RECT 6.145000 2.120000 6.315000 2.285000 ;
        RECT 6.835000 0.595000 7.165000 1.010000 ;
        RECT 7.845000 0.595000 8.015000 1.010000 ;
        RECT 8.335000 1.180000 8.505000 1.950000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 8.640000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 8.640000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 8.640000 0.085000 ;
      RECT 0.000000  3.245000 8.640000 3.415000 ;
      RECT 0.095000  0.085000 0.345000 1.250000 ;
      RECT 0.160000  1.920000 1.360000 2.090000 ;
      RECT 0.160000  2.090000 0.490000 2.980000 ;
      RECT 0.690000  2.260000 0.940000 3.245000 ;
      RECT 0.855000  0.920000 1.105000 0.940000 ;
      RECT 0.855000  0.940000 2.700000 1.190000 ;
      RECT 0.855000  1.190000 1.105000 1.250000 ;
      RECT 1.110000  2.090000 1.360000 2.905000 ;
      RECT 1.110000  2.905000 2.340000 3.075000 ;
      RECT 1.285000  0.085000 1.615000 0.410000 ;
      RECT 1.560000  1.190000 1.810000 2.735000 ;
      RECT 2.010000  2.190000 2.340000 2.905000 ;
      RECT 2.415000  0.085000 2.745000 0.430000 ;
      RECT 2.530000  1.190000 2.700000 1.360000 ;
      RECT 2.530000  1.360000 3.595000 1.680000 ;
      RECT 2.535000  2.190000 2.785000 2.905000 ;
      RECT 2.535000  2.905000 4.665000 3.075000 ;
      RECT 3.515000  2.625000 3.685000 2.905000 ;
      RECT 3.720000  0.085000 4.135000 0.510000 ;
      RECT 4.415000  2.625000 6.655000 2.795000 ;
      RECT 4.415000  2.795000 4.665000 2.905000 ;
      RECT 4.445000  0.350000 4.695000 0.670000 ;
      RECT 4.445000  0.670000 6.655000 0.840000 ;
      RECT 4.855000  2.965000 5.185000 3.245000 ;
      RECT 4.875000  0.085000 5.205000 0.500000 ;
      RECT 5.375000  2.795000 5.705000 2.980000 ;
      RECT 5.385000  0.350000 5.715000 0.670000 ;
      RECT 5.890000  2.965000 6.220000 3.245000 ;
      RECT 5.895000  0.085000 6.225000 0.500000 ;
      RECT 6.405000  0.255000 8.525000 0.425000 ;
      RECT 6.405000  0.425000 6.655000 0.670000 ;
      RECT 6.485000  2.290000 8.535000 2.460000 ;
      RECT 6.485000  2.460000 6.655000 2.625000 ;
      RECT 6.485000  2.795000 6.655000 2.980000 ;
      RECT 6.855000  2.630000 7.105000 3.245000 ;
      RECT 7.305000  2.460000 7.635000 2.980000 ;
      RECT 7.335000  0.425000 7.665000 0.840000 ;
      RECT 7.835000  2.630000 8.005000 3.245000 ;
      RECT 8.195000  0.425000 8.525000 0.840000 ;
      RECT 8.205000  2.460000 8.535000 2.980000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
      RECT 7.835000 -0.085000 8.005000 0.085000 ;
      RECT 7.835000  3.245000 8.005000 3.415000 ;
      RECT 8.315000 -0.085000 8.485000 0.085000 ;
      RECT 8.315000  3.245000 8.485000 3.415000 ;
  END
END sky130_fd_sc_hs__xor2_4
END LIBRARY
