* File: sky130_fd_sc_hs__nand3b_4.pxi.spice
* Created: Tue Sep  1 20:09:43 2020
* 
x_PM_SKY130_FD_SC_HS__NAND3B_4%A_N N_A_N_M1000_g N_A_N_c_105_n N_A_N_M1003_g
+ N_A_N_c_102_n N_A_N_c_107_n N_A_N_M1006_g A_N N_A_N_c_103_n N_A_N_c_104_n
+ PM_SKY130_FD_SC_HS__NAND3B_4%A_N
x_PM_SKY130_FD_SC_HS__NAND3B_4%C N_C_c_152_n N_C_M1004_g N_C_c_153_n N_C_c_154_n
+ N_C_c_155_n N_C_M1009_g N_C_c_156_n N_C_M1011_g N_C_c_162_n N_C_M1010_g
+ N_C_c_163_n N_C_M1012_g N_C_c_157_n N_C_M1013_g N_C_c_158_n C C C N_C_c_160_n
+ N_C_c_161_n PM_SKY130_FD_SC_HS__NAND3B_4%C
x_PM_SKY130_FD_SC_HS__NAND3B_4%A_89_172# N_A_89_172#_M1000_s N_A_89_172#_M1003_d
+ N_A_89_172#_c_248_n N_A_89_172#_M1014_g N_A_89_172#_c_234_n
+ N_A_89_172#_M1002_g N_A_89_172#_c_249_n N_A_89_172#_M1015_g
+ N_A_89_172#_c_235_n N_A_89_172#_M1016_g N_A_89_172#_c_236_n
+ N_A_89_172#_c_237_n N_A_89_172#_c_238_n N_A_89_172#_M1017_g
+ N_A_89_172#_c_239_n N_A_89_172#_c_240_n N_A_89_172#_M1020_g
+ N_A_89_172#_c_241_n N_A_89_172#_c_242_n N_A_89_172#_c_256_n
+ N_A_89_172#_c_243_n N_A_89_172#_c_244_n N_A_89_172#_c_245_n
+ N_A_89_172#_c_246_n N_A_89_172#_c_287_n N_A_89_172#_c_247_n
+ PM_SKY130_FD_SC_HS__NAND3B_4%A_89_172#
x_PM_SKY130_FD_SC_HS__NAND3B_4%B N_B_c_374_n N_B_M1007_g N_B_c_366_n N_B_c_367_n
+ N_B_M1001_g N_B_c_377_n N_B_M1008_g N_B_M1005_g N_B_M1018_g N_B_M1019_g B B B
+ N_B_c_372_n N_B_c_373_n PM_SKY130_FD_SC_HS__NAND3B_4%B
x_PM_SKY130_FD_SC_HS__NAND3B_4%VPWR N_VPWR_M1003_s N_VPWR_M1006_s N_VPWR_M1012_s
+ N_VPWR_M1015_d N_VPWR_M1008_s N_VPWR_c_438_n N_VPWR_c_439_n N_VPWR_c_440_n
+ N_VPWR_c_441_n VPWR N_VPWR_c_442_n N_VPWR_c_443_n N_VPWR_c_444_n
+ N_VPWR_c_445_n N_VPWR_c_446_n N_VPWR_c_447_n N_VPWR_c_448_n N_VPWR_c_437_n
+ PM_SKY130_FD_SC_HS__NAND3B_4%VPWR
x_PM_SKY130_FD_SC_HS__NAND3B_4%Y N_Y_M1002_s N_Y_M1017_s N_Y_M1010_d N_Y_M1014_s
+ N_Y_M1007_d N_Y_c_509_n N_Y_c_510_n N_Y_c_506_n N_Y_c_511_n N_Y_c_514_n
+ N_Y_c_560_n Y Y Y N_Y_c_508_n PM_SKY130_FD_SC_HS__NAND3B_4%Y
x_PM_SKY130_FD_SC_HS__NAND3B_4%VGND N_VGND_M1000_d N_VGND_M1009_s N_VGND_M1013_s
+ N_VGND_c_576_n N_VGND_c_577_n N_VGND_c_578_n N_VGND_c_579_n VGND
+ N_VGND_c_580_n N_VGND_c_581_n N_VGND_c_582_n N_VGND_c_583_n
+ PM_SKY130_FD_SC_HS__NAND3B_4%VGND
x_PM_SKY130_FD_SC_HS__NAND3B_4%A_297_82# N_A_297_82#_M1004_d N_A_297_82#_M1011_d
+ N_A_297_82#_M1001_s N_A_297_82#_M1018_s N_A_297_82#_c_643_n
+ N_A_297_82#_c_644_n N_A_297_82#_c_658_n N_A_297_82#_c_650_n
+ N_A_297_82#_c_716_n N_A_297_82#_c_660_n N_A_297_82#_c_727_n
+ N_A_297_82#_c_669_n N_A_297_82#_c_683_n N_A_297_82#_c_701_n
+ N_A_297_82#_c_651_n N_A_297_82#_c_652_n N_A_297_82#_c_645_n
+ N_A_297_82#_c_646_n N_A_297_82#_c_647_n N_A_297_82#_c_648_n
+ PM_SKY130_FD_SC_HS__NAND3B_4%A_297_82#
x_PM_SKY130_FD_SC_HS__NAND3B_4%A_744_74# N_A_744_74#_M1002_d N_A_744_74#_M1016_d
+ N_A_744_74#_M1020_d N_A_744_74#_M1005_d N_A_744_74#_M1019_d
+ N_A_744_74#_c_769_n N_A_744_74#_c_770_n N_A_744_74#_c_771_n
+ N_A_744_74#_c_772_n PM_SKY130_FD_SC_HS__NAND3B_4%A_744_74#
cc_1 VNB N_A_N_M1000_g 0.0287326f $X=-0.19 $Y=-0.245 $X2=0.805 $Y2=0.78
cc_2 VNB N_A_N_c_102_n 0.0105482f $X=-0.19 $Y=-0.245 $X2=1.27 $Y2=1.69
cc_3 VNB N_A_N_c_103_n 0.00482071f $X=-0.19 $Y=-0.245 $X2=0.93 $Y2=1.515
cc_4 VNB N_A_N_c_104_n 0.0526834f $X=-0.19 $Y=-0.245 $X2=1.095 $Y2=1.557
cc_5 VNB N_C_c_152_n 0.0150735f $X=-0.19 $Y=-0.245 $X2=0.805 $Y2=1.35
cc_6 VNB N_C_c_153_n 0.0210958f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_7 VNB N_C_c_154_n 0.00896832f $X=-0.19 $Y=-0.245 $X2=0.895 $Y2=1.765
cc_8 VNB N_C_c_155_n 0.0158871f $X=-0.19 $Y=-0.245 $X2=0.895 $Y2=2.26
cc_9 VNB N_C_c_156_n 0.0164552f $X=-0.19 $Y=-0.245 $X2=1.095 $Y2=1.69
cc_10 VNB N_C_c_157_n 0.0168136f $X=-0.19 $Y=-0.245 $X2=0.93 $Y2=1.557
cc_11 VNB N_C_c_158_n 0.0132043f $X=-0.19 $Y=-0.245 $X2=0.76 $Y2=1.515
cc_12 VNB C 0.00633246f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_C_c_160_n 0.0375955f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_C_c_161_n 0.042969f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_89_172#_c_234_n 0.0173647f $X=-0.19 $Y=-0.245 $X2=1.345 $Y2=1.765
cc_16 VNB N_A_89_172#_c_235_n 0.0152147f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_89_172#_c_236_n 0.015184f $X=-0.19 $Y=-0.245 $X2=0.93 $Y2=1.515
cc_18 VNB N_A_89_172#_c_237_n 0.104014f $X=-0.19 $Y=-0.245 $X2=0.93 $Y2=1.515
cc_19 VNB N_A_89_172#_c_238_n 0.014791f $X=-0.19 $Y=-0.245 $X2=1.095 $Y2=1.557
cc_20 VNB N_A_89_172#_c_239_n 0.0241507f $X=-0.19 $Y=-0.245 $X2=0.76 $Y2=1.665
cc_21 VNB N_A_89_172#_c_240_n 0.015888f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_89_172#_c_241_n 0.00678911f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_89_172#_c_242_n 0.00339641f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_89_172#_c_243_n 0.00551243f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_89_172#_c_244_n 0.03265f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_89_172#_c_245_n 0.00351706f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_89_172#_c_246_n 0.00467773f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_89_172#_c_247_n 0.00586556f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_B_c_366_n 0.0105482f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_B_c_367_n 0.0100568f $X=-0.19 $Y=-0.245 $X2=0.895 $Y2=1.765
cc_31 VNB N_B_M1001_g 0.0220707f $X=-0.19 $Y=-0.245 $X2=1.27 $Y2=1.69
cc_32 VNB N_B_M1005_g 0.0209473f $X=-0.19 $Y=-0.245 $X2=0.805 $Y2=1.557
cc_33 VNB N_B_M1018_g 0.0209424f $X=-0.19 $Y=-0.245 $X2=0.93 $Y2=1.515
cc_34 VNB N_B_M1019_g 0.0278788f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_B_c_372_n 0.0849184f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_B_c_373_n 0.00991188f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_VPWR_c_437_n 0.322901f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_Y_c_506_n 0.0100981f $X=-0.19 $Y=-0.245 $X2=0.76 $Y2=1.665
cc_39 VNB Y 0.00834423f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_Y_c_508_n 0.00413956f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_576_n 0.0145618f $X=-0.19 $Y=-0.245 $X2=1.345 $Y2=2.26
cc_42 VNB N_VGND_c_577_n 0.0450868f $X=-0.19 $Y=-0.245 $X2=0.805 $Y2=1.557
cc_43 VNB N_VGND_c_578_n 0.0184795f $X=-0.19 $Y=-0.245 $X2=0.76 $Y2=1.515
cc_44 VNB N_VGND_c_579_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_VGND_c_580_n 0.0179406f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_VGND_c_581_n 0.10598f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_VGND_c_582_n 0.422046f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_VGND_c_583_n 0.0209864f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A_297_82#_c_643_n 0.0446775f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_A_297_82#_c_644_n 0.0100851f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_A_297_82#_c_645_n 0.0200968f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_A_297_82#_c_646_n 0.0103159f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_A_297_82#_c_647_n 0.00255379f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_A_297_82#_c_648_n 0.00296506f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_A_744_74#_c_769_n 0.00258449f $X=-0.19 $Y=-0.245 $X2=0.93 $Y2=1.515
cc_56 VNB N_A_744_74#_c_770_n 0.0237054f $X=-0.19 $Y=-0.245 $X2=0.76 $Y2=1.665
cc_57 VNB N_A_744_74#_c_771_n 0.00534237f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_A_744_74#_c_772_n 0.00766753f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VPB N_A_N_c_105_n 0.0171679f $X=-0.19 $Y=1.66 $X2=0.895 $Y2=1.765
cc_60 VPB N_A_N_c_102_n 0.00897523f $X=-0.19 $Y=1.66 $X2=1.27 $Y2=1.69
cc_61 VPB N_A_N_c_107_n 0.0162478f $X=-0.19 $Y=1.66 $X2=1.345 $Y2=1.765
cc_62 VPB N_A_N_c_103_n 0.00525699f $X=-0.19 $Y=1.66 $X2=0.93 $Y2=1.515
cc_63 VPB N_A_N_c_104_n 0.0224408f $X=-0.19 $Y=1.66 $X2=1.095 $Y2=1.557
cc_64 VPB N_C_c_162_n 0.018852f $X=-0.19 $Y=1.66 $X2=1.345 $Y2=2.26
cc_65 VPB N_C_c_163_n 0.0161874f $X=-0.19 $Y=1.66 $X2=0.805 $Y2=1.557
cc_66 VPB N_C_c_158_n 0.00490368f $X=-0.19 $Y=1.66 $X2=0.76 $Y2=1.515
cc_67 VPB C 0.0181503f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_68 VPB N_C_c_160_n 0.0183479f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_69 VPB N_C_c_161_n 0.0211909f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_70 VPB N_A_89_172#_c_248_n 0.0186178f $X=-0.19 $Y=1.66 $X2=0.895 $Y2=2.26
cc_71 VPB N_A_89_172#_c_249_n 0.0198069f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_72 VPB N_A_89_172#_c_237_n 0.0169144f $X=-0.19 $Y=1.66 $X2=0.93 $Y2=1.515
cc_73 VPB N_A_89_172#_c_243_n 0.00295021f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_74 VPB N_B_c_374_n 0.017318f $X=-0.19 $Y=1.66 $X2=0.805 $Y2=1.35
cc_75 VPB N_B_c_366_n 0.00534307f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_76 VPB N_B_c_367_n 0.00602487f $X=-0.19 $Y=1.66 $X2=0.895 $Y2=1.765
cc_77 VPB N_B_c_377_n 0.0185177f $X=-0.19 $Y=1.66 $X2=1.345 $Y2=1.765
cc_78 VPB N_B_c_372_n 0.0468933f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_79 VPB N_VPWR_c_438_n 0.0121909f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_80 VPB N_VPWR_c_439_n 0.0528769f $X=-0.19 $Y=1.66 $X2=0.93 $Y2=1.557
cc_81 VPB N_VPWR_c_440_n 0.0043993f $X=-0.19 $Y=1.66 $X2=0.76 $Y2=1.515
cc_82 VPB N_VPWR_c_441_n 0.0165163f $X=-0.19 $Y=1.66 $X2=0.76 $Y2=1.665
cc_83 VPB N_VPWR_c_442_n 0.017758f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_84 VPB N_VPWR_c_443_n 0.0331904f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_85 VPB N_VPWR_c_444_n 0.0459336f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_86 VPB N_VPWR_c_445_n 0.00913469f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_87 VPB N_VPWR_c_446_n 0.0298504f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_88 VPB N_VPWR_c_447_n 0.0232358f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_89 VPB N_VPWR_c_448_n 0.0935916f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_90 VPB N_VPWR_c_437_n 0.0823877f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_91 VPB N_Y_c_509_n 0.00809783f $X=-0.19 $Y=1.66 $X2=0.93 $Y2=1.515
cc_92 VPB N_Y_c_510_n 8.85038e-19 $X=-0.19 $Y=1.66 $X2=1.095 $Y2=1.557
cc_93 VPB N_Y_c_511_n 0.00603019f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_94 VPB Y 0.00477667f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_95 VPB N_A_297_82#_c_643_n 0.0127478f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_96 VPB N_A_297_82#_c_650_n 0.00866242f $X=-0.19 $Y=1.66 $X2=0.93 $Y2=1.557
cc_97 VPB N_A_297_82#_c_651_n 0.0080099f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_98 VPB N_A_297_82#_c_652_n 0.00120419f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_99 VPB N_A_297_82#_c_645_n 0.0102237f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_100 N_A_N_M1000_g N_C_c_152_n 0.0258441f $X=0.805 $Y=0.78 $X2=-0.19
+ $Y2=-0.245
cc_101 N_A_N_c_102_n N_C_c_154_n 0.00554926f $X=1.27 $Y=1.69 $X2=0 $Y2=0
cc_102 N_A_N_c_104_n N_C_c_154_n 0.00139393f $X=1.095 $Y=1.557 $X2=0 $Y2=0
cc_103 N_A_N_c_102_n N_C_c_158_n 0.00248024f $X=1.27 $Y=1.69 $X2=0 $Y2=0
cc_104 N_A_N_c_104_n N_C_c_158_n 0.00268185f $X=1.095 $Y=1.557 $X2=0 $Y2=0
cc_105 N_A_N_c_102_n C 0.00239145f $X=1.27 $Y=1.69 $X2=0 $Y2=0
cc_106 N_A_N_M1000_g N_A_89_172#_c_242_n 0.00915372f $X=0.805 $Y=0.78 $X2=0
+ $Y2=0
cc_107 N_A_N_c_102_n N_A_89_172#_c_242_n 0.0048418f $X=1.27 $Y=1.69 $X2=0 $Y2=0
cc_108 N_A_N_c_103_n N_A_89_172#_c_242_n 0.0256619f $X=0.93 $Y=1.515 $X2=0 $Y2=0
cc_109 N_A_N_c_104_n N_A_89_172#_c_242_n 0.00149069f $X=1.095 $Y=1.557 $X2=0
+ $Y2=0
cc_110 N_A_N_c_105_n N_A_89_172#_c_256_n 0.00226148f $X=0.895 $Y=1.765 $X2=0
+ $Y2=0
cc_111 N_A_N_c_107_n N_A_89_172#_c_256_n 0.0075089f $X=1.345 $Y=1.765 $X2=0
+ $Y2=0
cc_112 N_A_N_c_103_n N_A_89_172#_c_256_n 0.00895896f $X=0.93 $Y=1.515 $X2=0
+ $Y2=0
cc_113 N_A_N_c_104_n N_A_89_172#_c_256_n 0.00315336f $X=1.095 $Y=1.557 $X2=0
+ $Y2=0
cc_114 N_A_N_M1000_g N_A_89_172#_c_243_n 0.00291514f $X=0.805 $Y=0.78 $X2=0
+ $Y2=0
cc_115 N_A_N_c_105_n N_A_89_172#_c_243_n 0.00112646f $X=0.895 $Y=1.765 $X2=0
+ $Y2=0
cc_116 N_A_N_c_102_n N_A_89_172#_c_243_n 0.00853049f $X=1.27 $Y=1.69 $X2=0 $Y2=0
cc_117 N_A_N_c_107_n N_A_89_172#_c_243_n 0.00544149f $X=1.345 $Y=1.765 $X2=0
+ $Y2=0
cc_118 N_A_N_c_103_n N_A_89_172#_c_243_n 0.0336678f $X=0.93 $Y=1.515 $X2=0 $Y2=0
cc_119 N_A_N_c_104_n N_A_89_172#_c_243_n 0.00302054f $X=1.095 $Y=1.557 $X2=0
+ $Y2=0
cc_120 N_A_N_M1000_g N_A_89_172#_c_246_n 0.0040074f $X=0.805 $Y=0.78 $X2=0 $Y2=0
cc_121 N_A_N_c_103_n N_A_89_172#_c_246_n 0.0261451f $X=0.93 $Y=1.515 $X2=0 $Y2=0
cc_122 N_A_N_c_104_n N_A_89_172#_c_246_n 0.00220658f $X=1.095 $Y=1.557 $X2=0
+ $Y2=0
cc_123 N_A_N_c_105_n N_VPWR_c_439_n 0.0106969f $X=0.895 $Y=1.765 $X2=0 $Y2=0
cc_124 N_A_N_c_105_n N_VPWR_c_443_n 0.00402388f $X=0.895 $Y=1.765 $X2=0 $Y2=0
cc_125 N_A_N_c_107_n N_VPWR_c_443_n 0.00402388f $X=1.345 $Y=1.765 $X2=0 $Y2=0
cc_126 N_A_N_c_107_n N_VPWR_c_444_n 0.00728857f $X=1.345 $Y=1.765 $X2=0 $Y2=0
cc_127 N_A_N_c_105_n N_VPWR_c_437_n 0.00462577f $X=0.895 $Y=1.765 $X2=0 $Y2=0
cc_128 N_A_N_c_107_n N_VPWR_c_437_n 0.00462577f $X=1.345 $Y=1.765 $X2=0 $Y2=0
cc_129 N_A_N_M1000_g N_VGND_c_577_n 0.00798327f $X=0.805 $Y=0.78 $X2=0 $Y2=0
cc_130 N_A_N_M1000_g N_VGND_c_582_n 0.00533081f $X=0.805 $Y=0.78 $X2=0 $Y2=0
cc_131 N_A_N_M1000_g N_A_297_82#_c_643_n 0.00747069f $X=0.805 $Y=0.78 $X2=0
+ $Y2=0
cc_132 N_A_N_c_105_n N_A_297_82#_c_643_n 0.00389051f $X=0.895 $Y=1.765 $X2=0
+ $Y2=0
cc_133 N_A_N_c_103_n N_A_297_82#_c_643_n 0.0342298f $X=0.93 $Y=1.515 $X2=0 $Y2=0
cc_134 N_A_N_c_104_n N_A_297_82#_c_643_n 0.0108353f $X=1.095 $Y=1.557 $X2=0
+ $Y2=0
cc_135 N_A_N_c_103_n N_A_297_82#_c_658_n 0.0289512f $X=0.93 $Y=1.515 $X2=0 $Y2=0
cc_136 N_A_N_c_104_n N_A_297_82#_c_658_n 0.00245611f $X=1.095 $Y=1.557 $X2=0
+ $Y2=0
cc_137 N_A_N_c_105_n N_A_297_82#_c_660_n 0.0145748f $X=0.895 $Y=1.765 $X2=0
+ $Y2=0
cc_138 N_A_N_c_107_n N_A_297_82#_c_660_n 0.0138613f $X=1.345 $Y=1.765 $X2=0
+ $Y2=0
cc_139 N_A_N_c_103_n N_A_297_82#_c_660_n 0.00458213f $X=0.93 $Y=1.515 $X2=0
+ $Y2=0
cc_140 N_A_N_M1000_g N_A_297_82#_c_646_n 0.0144512f $X=0.805 $Y=0.78 $X2=0 $Y2=0
cc_141 N_A_N_M1000_g N_A_297_82#_c_647_n 0.00116196f $X=0.805 $Y=0.78 $X2=0
+ $Y2=0
cc_142 N_C_c_163_n N_A_89_172#_c_248_n 0.0334767f $X=3.075 $Y=1.765 $X2=0 $Y2=0
cc_143 C N_A_89_172#_c_248_n 3.17149e-19 $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_144 N_C_c_157_n N_A_89_172#_c_237_n 0.0161146f $X=3.09 $Y=1.225 $X2=0 $Y2=0
cc_145 C N_A_89_172#_c_237_n 0.0056892f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_146 N_C_c_152_n N_A_89_172#_c_243_n 0.00135568f $X=1.41 $Y=1.225 $X2=0 $Y2=0
cc_147 N_C_c_154_n N_A_89_172#_c_243_n 0.00965829f $X=1.485 $Y=1.3 $X2=0 $Y2=0
cc_148 N_C_c_155_n N_A_89_172#_c_243_n 2.47368e-19 $X=1.84 $Y=1.225 $X2=0 $Y2=0
cc_149 N_C_c_158_n N_A_89_172#_c_243_n 0.00106338f $X=1.84 $Y=1.452 $X2=0 $Y2=0
cc_150 C N_A_89_172#_c_243_n 0.020564f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_151 N_C_c_152_n N_A_89_172#_c_244_n 0.00544416f $X=1.41 $Y=1.225 $X2=0 $Y2=0
cc_152 N_C_c_153_n N_A_89_172#_c_244_n 0.00392416f $X=1.765 $Y=1.3 $X2=0 $Y2=0
cc_153 N_C_c_155_n N_A_89_172#_c_244_n 0.0118156f $X=1.84 $Y=1.225 $X2=0 $Y2=0
cc_154 N_C_c_156_n N_A_89_172#_c_244_n 0.0121942f $X=2.59 $Y=1.225 $X2=0 $Y2=0
cc_155 N_C_c_157_n N_A_89_172#_c_244_n 0.0164035f $X=3.09 $Y=1.225 $X2=0 $Y2=0
cc_156 C N_A_89_172#_c_244_n 0.111296f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_157 N_C_c_160_n N_A_89_172#_c_244_n 0.0116694f $X=2.515 $Y=1.452 $X2=0 $Y2=0
cc_158 N_C_c_161_n N_A_89_172#_c_244_n 0.00472334f $X=3.075 $Y=1.495 $X2=0 $Y2=0
cc_159 N_C_c_152_n N_A_89_172#_c_246_n 4.85079e-19 $X=1.41 $Y=1.225 $X2=0 $Y2=0
cc_160 N_C_c_152_n N_A_89_172#_c_287_n 0.00624968f $X=1.41 $Y=1.225 $X2=0 $Y2=0
cc_161 N_C_c_157_n N_A_89_172#_c_247_n 0.00169516f $X=3.09 $Y=1.225 $X2=0 $Y2=0
cc_162 C N_A_89_172#_c_247_n 0.0127818f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_163 N_C_c_161_n N_A_89_172#_c_247_n 3.15585e-19 $X=3.075 $Y=1.495 $X2=0 $Y2=0
cc_164 N_C_c_162_n N_VPWR_c_440_n 0.00129917f $X=2.625 $Y=1.765 $X2=0 $Y2=0
cc_165 N_C_c_163_n N_VPWR_c_440_n 0.0156039f $X=3.075 $Y=1.765 $X2=0 $Y2=0
cc_166 N_C_c_162_n N_VPWR_c_442_n 0.00413917f $X=2.625 $Y=1.765 $X2=0 $Y2=0
cc_167 N_C_c_163_n N_VPWR_c_442_n 0.00413917f $X=3.075 $Y=1.765 $X2=0 $Y2=0
cc_168 N_C_c_162_n N_VPWR_c_444_n 0.0113214f $X=2.625 $Y=1.765 $X2=0 $Y2=0
cc_169 N_C_c_163_n N_VPWR_c_444_n 0.00129417f $X=3.075 $Y=1.765 $X2=0 $Y2=0
cc_170 N_C_c_162_n N_VPWR_c_437_n 0.00415095f $X=2.625 $Y=1.765 $X2=0 $Y2=0
cc_171 N_C_c_163_n N_VPWR_c_437_n 0.00416762f $X=3.075 $Y=1.765 $X2=0 $Y2=0
cc_172 N_C_c_163_n N_Y_c_510_n 5.61466e-19 $X=3.075 $Y=1.765 $X2=0 $Y2=0
cc_173 N_C_c_162_n N_Y_c_514_n 0.009084f $X=2.625 $Y=1.765 $X2=0 $Y2=0
cc_174 N_C_c_163_n N_Y_c_514_n 0.00990295f $X=3.075 $Y=1.765 $X2=0 $Y2=0
cc_175 C N_Y_c_514_n 0.0366527f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_176 N_C_c_161_n N_Y_c_514_n 0.0013173f $X=3.075 $Y=1.495 $X2=0 $Y2=0
cc_177 N_C_c_156_n N_VGND_c_576_n 6.53784e-19 $X=2.59 $Y=1.225 $X2=0 $Y2=0
cc_178 N_C_c_157_n N_VGND_c_576_n 0.0110145f $X=3.09 $Y=1.225 $X2=0 $Y2=0
cc_179 N_C_c_152_n N_VGND_c_577_n 0.00345905f $X=1.41 $Y=1.225 $X2=0 $Y2=0
cc_180 N_C_c_156_n N_VGND_c_578_n 0.00419934f $X=2.59 $Y=1.225 $X2=0 $Y2=0
cc_181 N_C_c_157_n N_VGND_c_578_n 0.00455951f $X=3.09 $Y=1.225 $X2=0 $Y2=0
cc_182 N_C_c_152_n N_VGND_c_580_n 0.00411482f $X=1.41 $Y=1.225 $X2=0 $Y2=0
cc_183 N_C_c_155_n N_VGND_c_580_n 0.00418922f $X=1.84 $Y=1.225 $X2=0 $Y2=0
cc_184 N_C_c_152_n N_VGND_c_582_n 0.00533081f $X=1.41 $Y=1.225 $X2=0 $Y2=0
cc_185 N_C_c_155_n N_VGND_c_582_n 0.00533081f $X=1.84 $Y=1.225 $X2=0 $Y2=0
cc_186 N_C_c_156_n N_VGND_c_582_n 0.00533081f $X=2.59 $Y=1.225 $X2=0 $Y2=0
cc_187 N_C_c_157_n N_VGND_c_582_n 0.00447788f $X=3.09 $Y=1.225 $X2=0 $Y2=0
cc_188 N_C_c_155_n N_VGND_c_583_n 0.00458735f $X=1.84 $Y=1.225 $X2=0 $Y2=0
cc_189 N_C_c_156_n N_VGND_c_583_n 0.00456635f $X=2.59 $Y=1.225 $X2=0 $Y2=0
cc_190 N_C_c_162_n N_A_297_82#_c_660_n 0.015556f $X=2.625 $Y=1.765 $X2=0 $Y2=0
cc_191 N_C_c_163_n N_A_297_82#_c_660_n 0.0127451f $X=3.075 $Y=1.765 $X2=0 $Y2=0
cc_192 N_C_c_158_n N_A_297_82#_c_660_n 0.00335948f $X=1.84 $Y=1.452 $X2=0 $Y2=0
cc_193 C N_A_297_82#_c_660_n 0.0307225f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_194 N_C_c_155_n N_A_297_82#_c_669_n 0.00974223f $X=1.84 $Y=1.225 $X2=0 $Y2=0
cc_195 N_C_c_156_n N_A_297_82#_c_669_n 0.0102985f $X=2.59 $Y=1.225 $X2=0 $Y2=0
cc_196 N_C_c_152_n N_A_297_82#_c_646_n 0.00922607f $X=1.41 $Y=1.225 $X2=0 $Y2=0
cc_197 N_C_c_152_n N_A_297_82#_c_647_n 0.00749188f $X=1.41 $Y=1.225 $X2=0 $Y2=0
cc_198 N_C_c_155_n N_A_297_82#_c_647_n 0.0106036f $X=1.84 $Y=1.225 $X2=0 $Y2=0
cc_199 N_C_c_156_n N_A_297_82#_c_648_n 0.0108343f $X=2.59 $Y=1.225 $X2=0 $Y2=0
cc_200 N_C_c_157_n N_A_297_82#_c_648_n 0.00240868f $X=3.09 $Y=1.225 $X2=0 $Y2=0
cc_201 N_C_c_157_n N_A_744_74#_c_771_n 7.1746e-19 $X=3.09 $Y=1.225 $X2=0 $Y2=0
cc_202 N_A_89_172#_c_239_n N_B_c_367_n 0.00681889f $X=5.32 $Y=1.26 $X2=0 $Y2=0
cc_203 N_A_89_172#_c_240_n N_B_M1001_g 0.0315164f $X=5.395 $Y=1.185 $X2=0 $Y2=0
cc_204 N_A_89_172#_c_239_n N_B_c_372_n 8.25902e-19 $X=5.32 $Y=1.26 $X2=0 $Y2=0
cc_205 N_A_89_172#_c_240_n N_B_c_373_n 7.20156e-19 $X=5.395 $Y=1.185 $X2=0 $Y2=0
cc_206 N_A_89_172#_c_248_n N_VPWR_c_440_n 0.0274173f $X=3.69 $Y=1.765 $X2=0
+ $Y2=0
cc_207 N_A_89_172#_c_248_n N_VPWR_c_446_n 0.00413917f $X=3.69 $Y=1.765 $X2=0
+ $Y2=0
cc_208 N_A_89_172#_c_249_n N_VPWR_c_446_n 0.00413917f $X=4.52 $Y=1.765 $X2=0
+ $Y2=0
cc_209 N_A_89_172#_c_249_n N_VPWR_c_447_n 0.023816f $X=4.52 $Y=1.765 $X2=0 $Y2=0
cc_210 N_A_89_172#_c_248_n N_VPWR_c_437_n 0.0041937f $X=3.69 $Y=1.765 $X2=0
+ $Y2=0
cc_211 N_A_89_172#_c_249_n N_VPWR_c_437_n 0.00417703f $X=4.52 $Y=1.765 $X2=0
+ $Y2=0
cc_212 N_A_89_172#_c_249_n N_Y_c_509_n 0.0168336f $X=4.52 $Y=1.765 $X2=0 $Y2=0
cc_213 N_A_89_172#_c_236_n N_Y_c_509_n 0.00943567f $X=4.89 $Y=1.26 $X2=0 $Y2=0
cc_214 N_A_89_172#_c_237_n N_Y_c_509_n 9.28586e-19 $X=4.61 $Y=1.26 $X2=0 $Y2=0
cc_215 N_A_89_172#_c_248_n N_Y_c_510_n 0.00389498f $X=3.69 $Y=1.765 $X2=0 $Y2=0
cc_216 N_A_89_172#_c_237_n N_Y_c_510_n 0.0167298f $X=4.61 $Y=1.26 $X2=0 $Y2=0
cc_217 N_A_89_172#_c_245_n N_Y_c_510_n 0.0603472f $X=4.445 $Y=1.465 $X2=0 $Y2=0
cc_218 N_A_89_172#_c_247_n N_Y_c_510_n 0.00138986f $X=3.685 $Y=1.095 $X2=0 $Y2=0
cc_219 N_A_89_172#_c_234_n N_Y_c_506_n 0.011661f $X=4.08 $Y=1.185 $X2=0 $Y2=0
cc_220 N_A_89_172#_c_235_n N_Y_c_506_n 0.0131408f $X=4.535 $Y=1.185 $X2=0 $Y2=0
cc_221 N_A_89_172#_c_236_n N_Y_c_506_n 0.00420528f $X=4.89 $Y=1.26 $X2=0 $Y2=0
cc_222 N_A_89_172#_c_237_n N_Y_c_506_n 0.0034731f $X=4.61 $Y=1.26 $X2=0 $Y2=0
cc_223 N_A_89_172#_c_238_n N_Y_c_506_n 0.0069204f $X=4.965 $Y=1.185 $X2=0 $Y2=0
cc_224 N_A_89_172#_c_245_n N_Y_c_506_n 0.0372722f $X=4.445 $Y=1.465 $X2=0 $Y2=0
cc_225 N_A_89_172#_c_247_n N_Y_c_506_n 0.00525886f $X=3.685 $Y=1.095 $X2=0 $Y2=0
cc_226 N_A_89_172#_c_239_n N_Y_c_511_n 0.00683915f $X=5.32 $Y=1.26 $X2=0 $Y2=0
cc_227 N_A_89_172#_c_248_n N_Y_c_514_n 0.00997679f $X=3.69 $Y=1.765 $X2=0 $Y2=0
cc_228 N_A_89_172#_c_247_n N_Y_c_514_n 0.00651328f $X=3.685 $Y=1.095 $X2=0 $Y2=0
cc_229 N_A_89_172#_c_249_n Y 0.00161596f $X=4.52 $Y=1.765 $X2=0 $Y2=0
cc_230 N_A_89_172#_c_235_n Y 3.1248e-19 $X=4.535 $Y=1.185 $X2=0 $Y2=0
cc_231 N_A_89_172#_c_237_n Y 0.00608482f $X=4.61 $Y=1.26 $X2=0 $Y2=0
cc_232 N_A_89_172#_c_238_n Y 0.00164483f $X=4.965 $Y=1.185 $X2=0 $Y2=0
cc_233 N_A_89_172#_c_239_n Y 0.00822151f $X=5.32 $Y=1.26 $X2=0 $Y2=0
cc_234 N_A_89_172#_c_240_n Y 0.00114729f $X=5.395 $Y=1.185 $X2=0 $Y2=0
cc_235 N_A_89_172#_c_241_n Y 0.0104475f $X=4.965 $Y=1.26 $X2=0 $Y2=0
cc_236 N_A_89_172#_c_245_n Y 0.0167252f $X=4.445 $Y=1.465 $X2=0 $Y2=0
cc_237 N_A_89_172#_c_238_n N_Y_c_508_n 0.00625476f $X=4.965 $Y=1.185 $X2=0 $Y2=0
cc_238 N_A_89_172#_c_239_n N_Y_c_508_n 0.00319434f $X=5.32 $Y=1.26 $X2=0 $Y2=0
cc_239 N_A_89_172#_c_240_n N_Y_c_508_n 0.0088709f $X=5.395 $Y=1.185 $X2=0 $Y2=0
cc_240 N_A_89_172#_c_242_n N_VGND_M1000_d 0.00489649f $X=1.265 $Y=1.095
+ $X2=-0.19 $Y2=-0.245
cc_241 N_A_89_172#_c_244_n N_VGND_M1009_s 0.00702535f $X=3.6 $Y=1.095 $X2=0
+ $Y2=0
cc_242 N_A_89_172#_c_244_n N_VGND_M1013_s 0.00259019f $X=3.6 $Y=1.095 $X2=0
+ $Y2=0
cc_243 N_A_89_172#_c_234_n N_VGND_c_576_n 0.00715259f $X=4.08 $Y=1.185 $X2=0
+ $Y2=0
cc_244 N_A_89_172#_c_244_n N_VGND_c_576_n 0.0220913f $X=3.6 $Y=1.095 $X2=0 $Y2=0
cc_245 N_A_89_172#_c_234_n N_VGND_c_581_n 0.00291649f $X=4.08 $Y=1.185 $X2=0
+ $Y2=0
cc_246 N_A_89_172#_c_235_n N_VGND_c_581_n 0.00291649f $X=4.535 $Y=1.185 $X2=0
+ $Y2=0
cc_247 N_A_89_172#_c_238_n N_VGND_c_581_n 0.00291649f $X=4.965 $Y=1.185 $X2=0
+ $Y2=0
cc_248 N_A_89_172#_c_240_n N_VGND_c_581_n 0.00291649f $X=5.395 $Y=1.185 $X2=0
+ $Y2=0
cc_249 N_A_89_172#_c_234_n N_VGND_c_582_n 0.00364365f $X=4.08 $Y=1.185 $X2=0
+ $Y2=0
cc_250 N_A_89_172#_c_235_n N_VGND_c_582_n 0.00359366f $X=4.535 $Y=1.185 $X2=0
+ $Y2=0
cc_251 N_A_89_172#_c_238_n N_VGND_c_582_n 0.00359121f $X=4.965 $Y=1.185 $X2=0
+ $Y2=0
cc_252 N_A_89_172#_c_240_n N_VGND_c_582_n 0.00359833f $X=5.395 $Y=1.185 $X2=0
+ $Y2=0
cc_253 N_A_89_172#_c_244_n N_A_297_82#_M1004_d 0.00176891f $X=3.6 $Y=1.095
+ $X2=-0.19 $Y2=-0.245
cc_254 N_A_89_172#_c_244_n N_A_297_82#_M1011_d 0.00250873f $X=3.6 $Y=1.095 $X2=0
+ $Y2=0
cc_255 N_A_89_172#_c_246_n N_A_297_82#_c_643_n 0.020614f $X=0.59 $Y=1.005 $X2=0
+ $Y2=0
cc_256 N_A_89_172#_M1003_d N_A_297_82#_c_660_n 0.00562653f $X=0.97 $Y=1.84 $X2=0
+ $Y2=0
cc_257 N_A_89_172#_c_248_n N_A_297_82#_c_660_n 0.0141361f $X=3.69 $Y=1.765 $X2=0
+ $Y2=0
cc_258 N_A_89_172#_c_249_n N_A_297_82#_c_660_n 0.0153446f $X=4.52 $Y=1.765 $X2=0
+ $Y2=0
cc_259 N_A_89_172#_c_256_n N_A_297_82#_c_660_n 0.0259986f $X=1.265 $Y=2.045
+ $X2=0 $Y2=0
cc_260 N_A_89_172#_c_240_n N_A_297_82#_c_683_n 5.14228e-19 $X=5.395 $Y=1.185
+ $X2=0 $Y2=0
cc_261 N_A_89_172#_M1000_s N_A_297_82#_c_646_n 0.00566964f $X=0.445 $Y=0.86
+ $X2=0 $Y2=0
cc_262 N_A_89_172#_c_242_n N_A_297_82#_c_646_n 0.0234296f $X=1.265 $Y=1.095
+ $X2=0 $Y2=0
cc_263 N_A_89_172#_c_244_n N_A_297_82#_c_646_n 0.0011585f $X=3.6 $Y=1.095 $X2=0
+ $Y2=0
cc_264 N_A_89_172#_c_246_n N_A_297_82#_c_646_n 0.0203761f $X=0.59 $Y=1.005 $X2=0
+ $Y2=0
cc_265 N_A_89_172#_c_287_n N_A_297_82#_c_646_n 0.00618821f $X=1.35 $Y=1.095
+ $X2=0 $Y2=0
cc_266 N_A_89_172#_c_244_n N_A_297_82#_c_647_n 0.0688738f $X=3.6 $Y=1.095 $X2=0
+ $Y2=0
cc_267 N_A_89_172#_c_244_n N_A_297_82#_c_648_n 0.0203381f $X=3.6 $Y=1.095 $X2=0
+ $Y2=0
cc_268 N_A_89_172#_c_247_n N_A_744_74#_M1002_d 0.00139751f $X=3.685 $Y=1.095
+ $X2=-0.19 $Y2=-0.245
cc_269 N_A_89_172#_c_234_n N_A_744_74#_c_771_n 0.0024281f $X=4.08 $Y=1.185 $X2=0
+ $Y2=0
cc_270 N_A_89_172#_c_237_n N_A_744_74#_c_771_n 0.00449869f $X=4.61 $Y=1.26 $X2=0
+ $Y2=0
cc_271 N_A_89_172#_c_245_n N_A_744_74#_c_771_n 0.00585628f $X=4.445 $Y=1.465
+ $X2=0 $Y2=0
cc_272 N_A_89_172#_c_247_n N_A_744_74#_c_771_n 0.00332029f $X=3.685 $Y=1.095
+ $X2=0 $Y2=0
cc_273 N_A_89_172#_c_234_n N_A_744_74#_c_772_n 0.0122631f $X=4.08 $Y=1.185 $X2=0
+ $Y2=0
cc_274 N_A_89_172#_c_235_n N_A_744_74#_c_772_n 0.0106216f $X=4.535 $Y=1.185
+ $X2=0 $Y2=0
cc_275 N_A_89_172#_c_238_n N_A_744_74#_c_772_n 0.0102551f $X=4.965 $Y=1.185
+ $X2=0 $Y2=0
cc_276 N_A_89_172#_c_240_n N_A_744_74#_c_772_n 0.0175315f $X=5.395 $Y=1.185
+ $X2=0 $Y2=0
cc_277 N_B_c_374_n N_VPWR_c_441_n 0.00261496f $X=5.46 $Y=1.765 $X2=0 $Y2=0
cc_278 N_B_c_377_n N_VPWR_c_441_n 0.00261496f $X=5.91 $Y=1.765 $X2=0 $Y2=0
cc_279 N_B_c_374_n N_VPWR_c_447_n 0.0113144f $X=5.46 $Y=1.765 $X2=0 $Y2=0
cc_280 N_B_c_377_n N_VPWR_c_447_n 0.00129368f $X=5.91 $Y=1.765 $X2=0 $Y2=0
cc_281 N_B_c_374_n N_VPWR_c_448_n 0.00129839f $X=5.46 $Y=1.765 $X2=0 $Y2=0
cc_282 N_B_c_377_n N_VPWR_c_448_n 0.0174135f $X=5.91 $Y=1.765 $X2=0 $Y2=0
cc_283 N_B_c_374_n N_VPWR_c_437_n 0.00415095f $X=5.46 $Y=1.765 $X2=0 $Y2=0
cc_284 N_B_c_377_n N_VPWR_c_437_n 0.00415095f $X=5.91 $Y=1.765 $X2=0 $Y2=0
cc_285 N_B_c_374_n N_Y_c_511_n 0.0187241f $X=5.46 $Y=1.765 $X2=0 $Y2=0
cc_286 N_B_c_366_n N_Y_c_511_n 0.0111614f $X=5.74 $Y=1.65 $X2=0 $Y2=0
cc_287 N_B_c_367_n N_Y_c_511_n 0.00128859f $X=5.55 $Y=1.65 $X2=0 $Y2=0
cc_288 N_B_c_377_n N_Y_c_511_n 0.00414619f $X=5.91 $Y=1.765 $X2=0 $Y2=0
cc_289 N_B_c_372_n N_Y_c_511_n 4.5915e-19 $X=6.965 $Y=1.485 $X2=0 $Y2=0
cc_290 N_B_c_373_n N_Y_c_511_n 0.00236962f $X=6.965 $Y=1.485 $X2=0 $Y2=0
cc_291 N_B_c_374_n Y 0.00179663f $X=5.46 $Y=1.765 $X2=0 $Y2=0
cc_292 N_B_c_367_n Y 0.00669648f $X=5.55 $Y=1.65 $X2=0 $Y2=0
cc_293 N_B_c_372_n Y 0.00471144f $X=6.965 $Y=1.485 $X2=0 $Y2=0
cc_294 N_B_c_373_n Y 0.0127966f $X=6.965 $Y=1.485 $X2=0 $Y2=0
cc_295 N_B_M1001_g N_Y_c_508_n 0.00141517f $X=5.895 $Y=0.74 $X2=0 $Y2=0
cc_296 N_B_M1001_g N_VGND_c_581_n 0.00291649f $X=5.895 $Y=0.74 $X2=0 $Y2=0
cc_297 N_B_M1005_g N_VGND_c_581_n 0.00291649f $X=6.325 $Y=0.74 $X2=0 $Y2=0
cc_298 N_B_M1018_g N_VGND_c_581_n 0.00291649f $X=6.755 $Y=0.74 $X2=0 $Y2=0
cc_299 N_B_M1019_g N_VGND_c_581_n 0.00291649f $X=7.185 $Y=0.74 $X2=0 $Y2=0
cc_300 N_B_M1001_g N_VGND_c_582_n 0.00359833f $X=5.895 $Y=0.74 $X2=0 $Y2=0
cc_301 N_B_M1005_g N_VGND_c_582_n 0.00359121f $X=6.325 $Y=0.74 $X2=0 $Y2=0
cc_302 N_B_M1018_g N_VGND_c_582_n 0.00359121f $X=6.755 $Y=0.74 $X2=0 $Y2=0
cc_303 N_B_M1019_g N_VGND_c_582_n 0.00362779f $X=7.185 $Y=0.74 $X2=0 $Y2=0
cc_304 N_B_c_374_n N_A_297_82#_c_660_n 0.0139026f $X=5.46 $Y=1.765 $X2=0 $Y2=0
cc_305 N_B_c_377_n N_A_297_82#_c_660_n 0.0151556f $X=5.91 $Y=1.765 $X2=0 $Y2=0
cc_306 N_B_c_372_n N_A_297_82#_c_660_n 0.00100114f $X=6.965 $Y=1.485 $X2=0 $Y2=0
cc_307 N_B_c_373_n N_A_297_82#_c_660_n 0.00437833f $X=6.965 $Y=1.485 $X2=0 $Y2=0
cc_308 N_B_M1001_g N_A_297_82#_c_683_n 0.00384298f $X=5.895 $Y=0.74 $X2=0 $Y2=0
cc_309 N_B_M1005_g N_A_297_82#_c_683_n 0.00843705f $X=6.325 $Y=0.74 $X2=0 $Y2=0
cc_310 N_B_M1018_g N_A_297_82#_c_683_n 0.00843705f $X=6.755 $Y=0.74 $X2=0 $Y2=0
cc_311 N_B_M1019_g N_A_297_82#_c_683_n 0.0129826f $X=7.185 $Y=0.74 $X2=0 $Y2=0
cc_312 N_B_c_372_n N_A_297_82#_c_683_n 0.00149218f $X=6.965 $Y=1.485 $X2=0 $Y2=0
cc_313 N_B_c_373_n N_A_297_82#_c_683_n 0.0772269f $X=6.965 $Y=1.485 $X2=0 $Y2=0
cc_314 N_B_c_377_n N_A_297_82#_c_701_n 0.00974114f $X=5.91 $Y=1.765 $X2=0 $Y2=0
cc_315 N_B_c_372_n N_A_297_82#_c_651_n 0.0303401f $X=6.965 $Y=1.485 $X2=0 $Y2=0
cc_316 N_B_c_373_n N_A_297_82#_c_651_n 0.0652259f $X=6.965 $Y=1.485 $X2=0 $Y2=0
cc_317 N_B_c_377_n N_A_297_82#_c_652_n 0.00397137f $X=5.91 $Y=1.765 $X2=0 $Y2=0
cc_318 N_B_c_372_n N_A_297_82#_c_652_n 0.00473088f $X=6.965 $Y=1.485 $X2=0 $Y2=0
cc_319 N_B_c_373_n N_A_297_82#_c_652_n 0.0146559f $X=6.965 $Y=1.485 $X2=0 $Y2=0
cc_320 N_B_M1018_g N_A_297_82#_c_645_n 7.10626e-19 $X=6.755 $Y=0.74 $X2=0 $Y2=0
cc_321 N_B_M1019_g N_A_297_82#_c_645_n 0.00947193f $X=7.185 $Y=0.74 $X2=0 $Y2=0
cc_322 N_B_c_372_n N_A_297_82#_c_645_n 0.0137996f $X=6.965 $Y=1.485 $X2=0 $Y2=0
cc_323 N_B_c_373_n N_A_297_82#_c_645_n 0.036909f $X=6.965 $Y=1.485 $X2=0 $Y2=0
cc_324 N_B_M1001_g N_A_744_74#_c_769_n 0.00118092f $X=5.895 $Y=0.74 $X2=0 $Y2=0
cc_325 N_B_c_372_n N_A_744_74#_c_769_n 0.00131386f $X=6.965 $Y=1.485 $X2=0 $Y2=0
cc_326 N_B_c_373_n N_A_744_74#_c_769_n 0.00389228f $X=6.965 $Y=1.485 $X2=0 $Y2=0
cc_327 N_B_M1001_g N_A_744_74#_c_770_n 0.0122981f $X=5.895 $Y=0.74 $X2=0 $Y2=0
cc_328 N_B_M1005_g N_A_744_74#_c_770_n 0.0120586f $X=6.325 $Y=0.74 $X2=0 $Y2=0
cc_329 N_B_M1018_g N_A_744_74#_c_770_n 0.0120586f $X=6.755 $Y=0.74 $X2=0 $Y2=0
cc_330 N_B_M1019_g N_A_744_74#_c_770_n 0.0122066f $X=7.185 $Y=0.74 $X2=0 $Y2=0
cc_331 N_VPWR_M1015_d N_Y_c_509_n 0.00542137f $X=4.595 $Y=1.84 $X2=0 $Y2=0
cc_332 N_VPWR_M1015_d N_Y_c_511_n 0.00267983f $X=4.595 $Y=1.84 $X2=0 $Y2=0
cc_333 N_VPWR_M1012_s N_Y_c_514_n 0.0176366f $X=3.15 $Y=1.84 $X2=0 $Y2=0
cc_334 N_VPWR_M1015_d N_Y_c_560_n 0.00637067f $X=4.595 $Y=1.84 $X2=0 $Y2=0
cc_335 N_VPWR_M1003_s N_A_297_82#_c_643_n 0.00244688f $X=0.135 $Y=1.84 $X2=0
+ $Y2=0
cc_336 N_VPWR_M1003_s N_A_297_82#_c_658_n 0.0224863f $X=0.135 $Y=1.84 $X2=0
+ $Y2=0
cc_337 N_VPWR_c_439_n N_A_297_82#_c_658_n 0.0153403f $X=0.28 $Y=2.495 $X2=0
+ $Y2=0
cc_338 N_VPWR_M1003_s N_A_297_82#_c_650_n 0.00244603f $X=0.135 $Y=1.84 $X2=0
+ $Y2=0
cc_339 N_VPWR_c_439_n N_A_297_82#_c_650_n 0.0125546f $X=0.28 $Y=2.495 $X2=0
+ $Y2=0
cc_340 N_VPWR_M1003_s N_A_297_82#_c_716_n 0.00696858f $X=0.135 $Y=1.84 $X2=0
+ $Y2=0
cc_341 N_VPWR_c_439_n N_A_297_82#_c_716_n 0.00149212f $X=0.28 $Y=2.495 $X2=0
+ $Y2=0
cc_342 N_VPWR_M1006_s N_A_297_82#_c_660_n 0.0408923f $X=1.42 $Y=1.84 $X2=0 $Y2=0
cc_343 N_VPWR_M1012_s N_A_297_82#_c_660_n 0.00839998f $X=3.15 $Y=1.84 $X2=0
+ $Y2=0
cc_344 N_VPWR_M1015_d N_A_297_82#_c_660_n 0.0183068f $X=4.595 $Y=1.84 $X2=0
+ $Y2=0
cc_345 N_VPWR_M1008_s N_A_297_82#_c_660_n 0.00482931f $X=5.985 $Y=1.84 $X2=0
+ $Y2=0
cc_346 N_VPWR_c_440_n N_A_297_82#_c_660_n 0.0300427f $X=3.38 $Y=2.815 $X2=0
+ $Y2=0
cc_347 N_VPWR_c_444_n N_A_297_82#_c_660_n 0.0805718f $X=2.565 $Y=3.032 $X2=0
+ $Y2=0
cc_348 N_VPWR_c_447_n N_A_297_82#_c_660_n 0.0557237f $X=5.4 $Y=3.032 $X2=0 $Y2=0
cc_349 N_VPWR_c_448_n N_A_297_82#_c_660_n 0.0327426f $X=7.4 $Y=2.325 $X2=0 $Y2=0
cc_350 N_VPWR_c_437_n N_A_297_82#_c_660_n 0.0974071f $X=7.44 $Y=3.33 $X2=0 $Y2=0
cc_351 N_VPWR_M1003_s N_A_297_82#_c_727_n 0.00556166f $X=0.135 $Y=1.84 $X2=0
+ $Y2=0
cc_352 N_VPWR_c_439_n N_A_297_82#_c_727_n 0.0144778f $X=0.28 $Y=2.495 $X2=0
+ $Y2=0
cc_353 N_VPWR_c_437_n N_A_297_82#_c_727_n 0.00648262f $X=7.44 $Y=3.33 $X2=0
+ $Y2=0
cc_354 N_VPWR_M1008_s N_A_297_82#_c_701_n 0.0131509f $X=5.985 $Y=1.84 $X2=0
+ $Y2=0
cc_355 N_VPWR_c_448_n N_A_297_82#_c_701_n 0.0121673f $X=7.4 $Y=2.325 $X2=0 $Y2=0
cc_356 N_VPWR_M1008_s N_A_297_82#_c_651_n 0.0309213f $X=5.985 $Y=1.84 $X2=0
+ $Y2=0
cc_357 N_VPWR_c_448_n N_A_297_82#_c_651_n 0.0889948f $X=7.4 $Y=2.325 $X2=0 $Y2=0
cc_358 N_VPWR_M1008_s N_A_297_82#_c_652_n 0.00279262f $X=5.985 $Y=1.84 $X2=0
+ $Y2=0
cc_359 N_Y_c_506_n N_VGND_c_576_n 0.00115716f $X=4.925 $Y=0.965 $X2=0 $Y2=0
cc_360 N_Y_M1010_d N_A_297_82#_c_660_n 0.0055969f $X=2.7 $Y=1.84 $X2=0 $Y2=0
cc_361 N_Y_M1014_s N_A_297_82#_c_660_n 0.0200688f $X=3.765 $Y=1.84 $X2=0 $Y2=0
cc_362 N_Y_M1007_d N_A_297_82#_c_660_n 0.00557657f $X=5.535 $Y=1.84 $X2=0 $Y2=0
cc_363 N_Y_c_511_n N_A_297_82#_c_660_n 0.0390088f $X=5.685 $Y=2.02 $X2=0 $Y2=0
cc_364 N_Y_c_514_n N_A_297_82#_c_660_n 0.135302f $X=3.75 $Y=1.98 $X2=0 $Y2=0
cc_365 N_Y_c_560_n N_A_297_82#_c_660_n 0.0187125f $X=5.04 $Y=1.98 $X2=0 $Y2=0
cc_366 N_Y_c_508_n N_A_297_82#_c_683_n 0.00497712f $X=5.04 $Y=1.13 $X2=0 $Y2=0
cc_367 N_Y_c_511_n N_A_297_82#_c_701_n 0.00990771f $X=5.685 $Y=2.02 $X2=0 $Y2=0
cc_368 N_Y_c_511_n N_A_297_82#_c_652_n 0.0125669f $X=5.685 $Y=2.02 $X2=0 $Y2=0
cc_369 N_Y_c_506_n N_A_744_74#_M1016_d 0.00189973f $X=4.925 $Y=0.965 $X2=0 $Y2=0
cc_370 N_Y_M1002_s N_A_744_74#_c_772_n 0.00207408f $X=4.155 $Y=0.37 $X2=0 $Y2=0
cc_371 N_Y_M1017_s N_A_744_74#_c_772_n 0.00168993f $X=5.04 $Y=0.37 $X2=0 $Y2=0
cc_372 N_Y_c_506_n N_A_744_74#_c_772_n 0.0365346f $X=4.925 $Y=0.965 $X2=0 $Y2=0
cc_373 N_Y_c_508_n N_A_744_74#_c_772_n 0.0233947f $X=5.04 $Y=1.13 $X2=0 $Y2=0
cc_374 N_VGND_c_577_n N_A_297_82#_c_644_n 0.00387622f $X=0.935 $Y=0 $X2=0 $Y2=0
cc_375 N_VGND_c_582_n N_A_297_82#_c_644_n 0.00537088f $X=7.44 $Y=0 $X2=0 $Y2=0
cc_376 N_VGND_M1009_s N_A_297_82#_c_669_n 0.0117523f $X=1.915 $Y=0.41 $X2=0
+ $Y2=0
cc_377 N_VGND_c_578_n N_A_297_82#_c_669_n 0.00237563f $X=3.14 $Y=0 $X2=0 $Y2=0
cc_378 N_VGND_c_580_n N_A_297_82#_c_669_n 0.00236949f $X=1.97 $Y=0 $X2=0 $Y2=0
cc_379 N_VGND_c_582_n N_A_297_82#_c_669_n 0.011866f $X=7.44 $Y=0 $X2=0 $Y2=0
cc_380 N_VGND_c_583_n N_A_297_82#_c_669_n 0.0374471f $X=2.16 $Y=0 $X2=0 $Y2=0
cc_381 N_VGND_M1000_d N_A_297_82#_c_646_n 0.00852962f $X=0.88 $Y=0.41 $X2=0
+ $Y2=0
cc_382 N_VGND_c_577_n N_A_297_82#_c_646_n 0.0381142f $X=0.935 $Y=0 $X2=0 $Y2=0
cc_383 N_VGND_c_580_n N_A_297_82#_c_646_n 0.00294479f $X=1.97 $Y=0 $X2=0 $Y2=0
cc_384 N_VGND_c_582_n N_A_297_82#_c_646_n 0.0271405f $X=7.44 $Y=0 $X2=0 $Y2=0
cc_385 N_VGND_c_577_n N_A_297_82#_c_647_n 0.00145202f $X=0.935 $Y=0 $X2=0 $Y2=0
cc_386 N_VGND_c_580_n N_A_297_82#_c_647_n 0.0121348f $X=1.97 $Y=0 $X2=0 $Y2=0
cc_387 N_VGND_c_582_n N_A_297_82#_c_647_n 0.0116628f $X=7.44 $Y=0 $X2=0 $Y2=0
cc_388 N_VGND_c_583_n N_A_297_82#_c_647_n 0.00469436f $X=2.16 $Y=0 $X2=0 $Y2=0
cc_389 N_VGND_c_576_n N_A_297_82#_c_648_n 0.0176756f $X=3.305 $Y=0.615 $X2=0
+ $Y2=0
cc_390 N_VGND_c_578_n N_A_297_82#_c_648_n 0.0121755f $X=3.14 $Y=0 $X2=0 $Y2=0
cc_391 N_VGND_c_582_n N_A_297_82#_c_648_n 0.0116241f $X=7.44 $Y=0 $X2=0 $Y2=0
cc_392 N_VGND_c_583_n N_A_297_82#_c_648_n 0.00474851f $X=2.16 $Y=0 $X2=0 $Y2=0
cc_393 N_VGND_c_576_n N_A_744_74#_c_771_n 0.0197752f $X=3.305 $Y=0.615 $X2=0
+ $Y2=0
cc_394 N_VGND_c_581_n N_A_744_74#_c_771_n 0.158354f $X=7.44 $Y=0 $X2=0 $Y2=0
cc_395 N_VGND_c_582_n N_A_744_74#_c_771_n 0.132997f $X=7.44 $Y=0 $X2=0 $Y2=0
cc_396 N_A_297_82#_c_683_n N_A_744_74#_M1005_d 0.00333133f $X=7.245 $Y=0.925
+ $X2=0 $Y2=0
cc_397 N_A_297_82#_c_683_n N_A_744_74#_M1019_d 0.00874113f $X=7.245 $Y=0.925
+ $X2=0 $Y2=0
cc_398 N_A_297_82#_c_645_n N_A_744_74#_M1019_d 0.0037774f $X=7.33 $Y=1.82 $X2=0
+ $Y2=0
cc_399 N_A_297_82#_M1001_s N_A_744_74#_c_770_n 0.00172259f $X=5.97 $Y=0.37 $X2=0
+ $Y2=0
cc_400 N_A_297_82#_M1018_s N_A_744_74#_c_770_n 0.00172259f $X=6.83 $Y=0.37 $X2=0
+ $Y2=0
cc_401 N_A_297_82#_c_683_n N_A_744_74#_c_770_n 0.0780631f $X=7.245 $Y=0.925
+ $X2=0 $Y2=0
