# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_hs__nand4bb_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__nand4bb_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  10.08000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A_N
    ANTENNAGATEAREA  0.363000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.440000 1.450000 0.835000 1.780000 ;
    END
  END A_N
  PIN B_N
    ANTENNAGATEAREA  0.363000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.465000 1.550000 1.795000 1.880000 ;
    END
  END B_N
  PIN C
    ANTENNAGATEAREA  1.116000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.185000 1.320000 7.610000 1.650000 ;
        RECT 6.845000 1.650000 7.075000 1.780000 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  1.116000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.265000 1.300000 9.955000 1.780000 ;
    END
  END D
  PIN Y
    ANTENNADIFFAREA  3.236100 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.320000 0.595000 2.650000 0.870000 ;
        RECT 2.320000 0.870000 3.505000 1.040000 ;
        RECT 2.525000 2.060000 4.815000 2.230000 ;
        RECT 2.525000 2.230000 2.965000 2.990000 ;
        RECT 3.335000 0.595000 3.505000 0.870000 ;
        RECT 3.335000 1.040000 3.505000 1.090000 ;
        RECT 3.335000 1.090000 5.685000 1.260000 ;
        RECT 3.635000 2.230000 3.865000 2.990000 ;
        RECT 4.485000 1.850000 6.665000 1.950000 ;
        RECT 4.485000 1.950000 9.515000 1.990000 ;
        RECT 4.485000 1.990000 5.685000 2.020000 ;
        RECT 4.485000 2.020000 4.815000 2.060000 ;
        RECT 4.535000 2.230000 4.815000 2.980000 ;
        RECT 5.515000 1.260000 5.685000 1.820000 ;
        RECT 5.515000 1.820000 6.665000 1.850000 ;
        RECT 5.515000 2.020000 5.685000 2.980000 ;
        RECT 6.335000 1.990000 9.515000 2.120000 ;
        RECT 6.335000 2.120000 6.665000 2.980000 ;
        RECT 7.335000 1.820000 7.665000 1.950000 ;
        RECT 7.335000 2.120000 7.665000 2.980000 ;
        RECT 8.285000 2.120000 8.615000 2.980000 ;
        RECT 9.185000 2.120000 9.515000 2.980000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 10.080000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 10.080000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 10.080000 0.085000 ;
      RECT 0.000000  3.245000 10.080000 3.415000 ;
      RECT 0.100000  0.550000  0.445000 0.660000 ;
      RECT 0.100000  0.660000  1.760000 0.830000 ;
      RECT 0.100000  0.830000  0.445000 1.280000 ;
      RECT 0.100000  1.280000  0.270000 1.950000 ;
      RECT 0.100000  1.950000  0.815000 2.120000 ;
      RECT 0.115000  2.290000  0.445000 3.245000 ;
      RECT 0.625000  0.085000  0.955000 0.490000 ;
      RECT 0.645000  2.120000  0.815000 2.980000 ;
      RECT 1.015000  2.390000  1.345000 3.245000 ;
      RECT 1.125000  1.000000  1.420000 1.330000 ;
      RECT 1.125000  1.330000  1.295000 2.050000 ;
      RECT 1.125000  2.050000  2.135000 2.220000 ;
      RECT 1.515000  2.220000  1.795000 2.980000 ;
      RECT 1.590000  0.830000  1.760000 1.210000 ;
      RECT 1.590000  1.210000  3.165000 1.380000 ;
      RECT 1.930000  0.255000  3.935000 0.425000 ;
      RECT 1.930000  0.425000  2.100000 1.040000 ;
      RECT 1.965000  1.720000  4.315000 1.890000 ;
      RECT 1.965000  1.890000  2.135000 2.050000 ;
      RECT 2.005000  2.390000  2.335000 3.245000 ;
      RECT 2.155000  1.380000  3.165000 1.550000 ;
      RECT 2.820000  0.425000  3.150000 0.700000 ;
      RECT 3.135000  2.400000  3.465000 3.245000 ;
      RECT 3.685000  0.425000  3.935000 0.750000 ;
      RECT 3.685000  0.750000  5.895000 0.920000 ;
      RECT 4.035000  2.400000  4.365000 3.245000 ;
      RECT 4.115000  0.255000  7.745000 0.425000 ;
      RECT 4.115000  0.425000  5.385000 0.580000 ;
      RECT 4.145000  1.430000  5.345000 1.680000 ;
      RECT 4.145000  1.680000  4.315000 1.720000 ;
      RECT 4.985000  2.190000  5.315000 3.245000 ;
      RECT 5.565000  0.595000  5.895000 0.750000 ;
      RECT 5.885000  2.160000  6.135000 3.245000 ;
      RECT 6.125000  0.595000  6.375000 0.980000 ;
      RECT 6.125000  0.980000  9.965000 1.130000 ;
      RECT 6.125000  1.130000  8.095000 1.150000 ;
      RECT 6.555000  0.425000  6.885000 0.810000 ;
      RECT 6.835000  2.290000  7.165000 3.245000 ;
      RECT 7.065000  0.595000  7.235000 0.980000 ;
      RECT 7.415000  0.425000  7.745000 0.810000 ;
      RECT 7.865000  2.290000  8.115000 3.245000 ;
      RECT 7.925000  0.350000  8.095000 0.960000 ;
      RECT 7.925000  0.960000  9.965000 0.980000 ;
      RECT 8.275000  0.085000  8.605000 0.790000 ;
      RECT 8.785000  0.350000  8.955000 0.960000 ;
      RECT 8.815000  2.290000  8.985000 3.245000 ;
      RECT 9.135000  0.085000  9.465000 0.790000 ;
      RECT 9.635000  0.350000  9.965000 0.960000 ;
      RECT 9.715000  1.950000  9.965000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
      RECT 7.835000 -0.085000 8.005000 0.085000 ;
      RECT 7.835000  3.245000 8.005000 3.415000 ;
      RECT 8.315000 -0.085000 8.485000 0.085000 ;
      RECT 8.315000  3.245000 8.485000 3.415000 ;
      RECT 8.795000 -0.085000 8.965000 0.085000 ;
      RECT 8.795000  3.245000 8.965000 3.415000 ;
      RECT 9.275000 -0.085000 9.445000 0.085000 ;
      RECT 9.275000  3.245000 9.445000 3.415000 ;
      RECT 9.755000 -0.085000 9.925000 0.085000 ;
      RECT 9.755000  3.245000 9.925000 3.415000 ;
  END
END sky130_fd_sc_hs__nand4bb_4
END LIBRARY
