* File: sky130_fd_sc_hs__sdfxbp_2.spice
* Created: Tue Sep  1 20:23:36 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hs__sdfxbp_2.pex.spice"
.subckt sky130_fd_sc_hs__sdfxbp_2  VNB VPB SCE D SCD CLK VPWR Q Q_N VGND
* 
* VGND	VGND
* Q_N	Q_N
* Q	Q
* VPWR	VPWR
* CLK	CLK
* SCD	SCD
* D	D
* SCE	SCE
* VPB	VPB
* VNB	VNB
MM1036 N_VGND_M1036_d N_SCE_M1036_g N_A_36_74#_M1036_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.0735 AS=0.1197 PD=0.77 PS=1.41 NRD=19.992 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75002.7 A=0.063 P=1.14 MULT=1
MM1016 A_223_74# N_A_36_74#_M1016_g N_VGND_M1036_d VNB NLOWVT L=0.15 W=0.42
+ AD=0.0504 AS=0.0735 PD=0.66 PS=0.77 NRD=18.564 NRS=0 M=1 R=2.8 SA=75000.7
+ SB=75002.2 A=0.063 P=1.14 MULT=1
MM1017 N_A_301_74#_M1017_d N_D_M1017_g A_223_74# VNB NLOWVT L=0.15 W=0.42
+ AD=0.12495 AS=0.0504 PD=1.015 PS=0.66 NRD=44.28 NRS=18.564 M=1 R=2.8
+ SA=75001.1 SB=75001.9 A=0.063 P=1.14 MULT=1
MM1031 A_450_74# N_SCE_M1031_g N_A_301_74#_M1017_d VNB NLOWVT L=0.15 W=0.42
+ AD=0.0504 AS=0.12495 PD=0.66 PS=1.015 NRD=18.564 NRS=45.708 M=1 R=2.8
+ SA=75001.8 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1026 N_VGND_M1026_d N_SCD_M1026_g A_450_74# VNB NLOWVT L=0.15 W=0.42
+ AD=0.0877655 AS=0.0504 PD=0.796552 PS=0.66 NRD=22.848 NRS=18.564 M=1 R=2.8
+ SA=75002.2 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1004 N_A_630_74#_M1004_d N_CLK_M1004_g N_VGND_M1026_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.154634 PD=2.05 PS=1.40345 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.6
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1015 N_A_828_74#_M1015_d N_A_630_74#_M1015_g N_VGND_M1015_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1998 AS=0.2109 PD=2.02 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1020 N_A_1021_97#_M1020_d N_A_630_74#_M1020_g N_A_301_74#_M1020_s VNB NLOWVT
+ L=0.15 W=0.42 AD=0.1281 AS=0.1155 PD=1.03 PS=1.39 NRD=94.284 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75003.7 A=0.063 P=1.14 MULT=1
MM1033 A_1173_97# N_A_828_74#_M1033_g N_A_1021_97#_M1020_d VNB NLOWVT L=0.15
+ W=0.42 AD=0.082125 AS=0.1281 PD=0.885 PS=1.03 NRD=40.152 NRS=0 M=1 R=2.8
+ SA=75001 SB=75002.9 A=0.063 P=1.14 MULT=1
MM1018 N_VGND_M1018_d N_A_1243_48#_M1018_g A_1173_97# VNB NLOWVT L=0.15 W=0.42
+ AD=0.125004 AS=0.082125 PD=1.00454 PS=0.885 NRD=0 NRS=40.152 M=1 R=2.8
+ SA=75001.1 SB=75003.4 A=0.063 P=1.14 MULT=1
MM1021 N_A_1243_48#_M1021_d N_A_1021_97#_M1021_g N_VGND_M1018_d VNB NLOWVT
+ L=0.15 W=0.55 AD=0.077 AS=0.163696 PD=0.83 PS=1.31546 NRD=0 NRS=72 M=1
+ R=3.66667 SA=75001.5 SB=75002.2 A=0.0825 P=1.4 MULT=1
MM1037 N_A_1511_74#_M1037_d N_A_828_74#_M1037_g N_A_1243_48#_M1021_d VNB NLOWVT
+ L=0.15 W=0.55 AD=0.163696 AS=0.077 PD=1.31546 PS=0.83 NRD=72 NRS=0 M=1
+ R=3.66667 SA=75001.9 SB=75001.8 A=0.0825 P=1.4 MULT=1
MM1011 A_1663_74# N_A_630_74#_M1011_g N_A_1511_74#_M1037_d VNB NLOWVT L=0.15
+ W=0.42 AD=0.0504 AS=0.125004 PD=0.66 PS=1.00454 NRD=18.564 NRS=0 M=1 R=2.8
+ SA=75003.1 SB=75001.5 A=0.063 P=1.14 MULT=1
MM1012 N_VGND_M1012_d N_A_1711_48#_M1012_g A_1663_74# VNB NLOWVT L=0.15 W=0.42
+ AD=0.139976 AS=0.0504 PD=1.06448 PS=0.66 NRD=79.5 NRS=18.564 M=1 R=2.8
+ SA=75003.4 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1029 N_A_1711_48#_M1029_d N_A_1511_74#_M1029_g N_VGND_M1012_d VNB NLOWVT
+ L=0.15 W=0.74 AD=0.2109 AS=0.246624 PD=2.05 PS=1.87552 NRD=0 NRS=45.12 M=1
+ R=4.93333 SA=75002.5 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1000 N_VGND_M1000_d N_A_1711_48#_M1000_g N_Q_M1000_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.2627 AS=0.1036 PD=2.19 PS=1.02 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75000.3
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1024 N_VGND_M1024_d N_A_1711_48#_M1024_g N_Q_M1000_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.1036 PD=2.05 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.7
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1023 N_VGND_M1023_d N_A_1711_48#_M1023_g N_A_2322_368#_M1023_s VNB NLOWVT
+ L=0.15 W=0.64 AD=0.12007 AS=0.1824 PD=1.02029 PS=1.85 NRD=12.648 NRS=0 M=1
+ R=4.26667 SA=75000.2 SB=75001.1 A=0.096 P=1.58 MULT=1
MM1001 N_VGND_M1023_d N_A_2322_368#_M1001_g N_Q_N_M1001_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.13883 AS=0.10915 PD=1.17971 PS=1.035 NRD=2.424 NRS=0.804 M=1
+ R=4.93333 SA=75000.7 SB=75000.6 A=0.111 P=1.78 MULT=1
MM1022 N_VGND_M1022_d N_A_2322_368#_M1022_g N_Q_N_M1001_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1962 AS=0.10915 PD=2.05 PS=1.035 NRD=0 NRS=1.62 M=1 R=4.93333
+ SA=75001.1 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1010 N_VPWR_M1010_d N_SCE_M1010_g N_A_36_74#_M1010_s VPB PSHORT L=0.15 W=0.64
+ AD=0.096 AS=0.2432 PD=0.94 PS=2.04 NRD=3.0732 NRS=29.2348 M=1 R=4.26667
+ SA=75000.3 SB=75003 A=0.096 P=1.58 MULT=1
MM1013 A_238_453# N_SCE_M1013_g N_VPWR_M1010_d VPB PSHORT L=0.15 W=0.64
+ AD=0.0864 AS=0.096 PD=0.91 PS=0.94 NRD=24.625 NRS=3.0732 M=1 R=4.26667
+ SA=75000.8 SB=75002.6 A=0.096 P=1.58 MULT=1
MM1003 N_A_301_74#_M1003_d N_D_M1003_g A_238_453# VPB PSHORT L=0.15 W=0.64
+ AD=0.1136 AS=0.0864 PD=0.995 PS=0.91 NRD=19.9955 NRS=24.625 M=1 R=4.26667
+ SA=75001.2 SB=75002.1 A=0.096 P=1.58 MULT=1
MM1030 A_423_453# N_A_36_74#_M1030_g N_A_301_74#_M1003_d VPB PSHORT L=0.15
+ W=0.64 AD=0.1072 AS=0.1136 PD=0.975 PS=0.995 NRD=34.6129 NRS=3.0732 M=1
+ R=4.26667 SA=75001.7 SB=75001.6 A=0.096 P=1.58 MULT=1
MM1019 N_VPWR_M1019_d N_SCD_M1019_g A_423_453# VPB PSHORT L=0.15 W=0.64
+ AD=0.188973 AS=0.1072 PD=1.26545 PS=0.975 NRD=44.6205 NRS=34.6129 M=1
+ R=4.26667 SA=75002.2 SB=75001.1 A=0.096 P=1.58 MULT=1
MM1028 N_A_630_74#_M1028_d N_CLK_M1028_g N_VPWR_M1019_d VPB PSHORT L=0.15 W=1.12
+ AD=0.5656 AS=0.330702 PD=3.25 PS=2.21455 NRD=2.6201 NRS=25.4918 M=1 R=7.46667
+ SA=75001.7 SB=75000.4 A=0.168 P=2.54 MULT=1
MM1035 N_A_828_74#_M1035_d N_A_630_74#_M1035_g N_VPWR_M1035_s VPB PSHORT L=0.15
+ W=1.12 AD=0.3304 AS=0.3304 PD=2.83 PS=2.83 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75000.2 A=0.168 P=2.54 MULT=1
MM1007 N_A_1021_97#_M1007_d N_A_828_74#_M1007_g N_A_301_74#_M1007_s VPB PSHORT
+ L=0.15 W=0.42 AD=0.08085 AS=0.1239 PD=0.805 PS=1.43 NRD=4.6886 NRS=4.6886 M=1
+ R=2.8 SA=75000.2 SB=75004.1 A=0.063 P=1.14 MULT=1
MM1014 A_1217_499# N_A_630_74#_M1014_g N_A_1021_97#_M1007_d VPB PSHORT L=0.15
+ W=0.42 AD=0.0567 AS=0.08085 PD=0.69 PS=0.805 NRD=37.5088 NRS=44.5417 M=1 R=2.8
+ SA=75000.8 SB=75003.6 A=0.063 P=1.14 MULT=1
MM1038 N_VPWR_M1038_d N_A_1243_48#_M1038_g A_1217_499# VPB PSHORT L=0.15 W=0.42
+ AD=0.126375 AS=0.0567 PD=1.02333 PS=0.69 NRD=115.324 NRS=37.5088 M=1 R=2.8
+ SA=75001.2 SB=75003.1 A=0.063 P=1.14 MULT=1
MM1027 N_A_1243_48#_M1027_d N_A_1021_97#_M1027_g N_VPWR_M1038_d VPB PSHORT
+ L=0.15 W=0.84 AD=0.2709 AS=0.25275 PD=1.485 PS=2.04667 NRD=5.8509 NRS=57.6619
+ M=1 R=5.6 SA=75001 SB=75001.9 A=0.126 P=1.98 MULT=1
MM1008 N_A_1511_74#_M1008_d N_A_630_74#_M1008_g N_A_1243_48#_M1027_d VPB PSHORT
+ L=0.15 W=0.84 AD=0.1904 AS=0.2709 PD=1.63333 PS=1.485 NRD=2.3443 NRS=79.7259
+ M=1 R=5.6 SA=75001.8 SB=75001.1 A=0.126 P=1.98 MULT=1
MM1005 A_1691_508# N_A_828_74#_M1005_g N_A_1511_74#_M1008_d VPB PSHORT L=0.15
+ W=0.42 AD=0.0567 AS=0.0952 PD=0.69 PS=0.816667 NRD=37.5088 NRS=44.5417 M=1
+ R=2.8 SA=75003 SB=75001.4 A=0.063 P=1.14 MULT=1
MM1009 N_VPWR_M1009_d N_A_1711_48#_M1009_g A_1691_508# VPB PSHORT L=0.15 W=0.42
+ AD=0.118754 AS=0.0567 PD=0.940563 PS=0.69 NRD=60.9715 NRS=37.5088 M=1 R=2.8
+ SA=75003.4 SB=75000.9 A=0.063 P=1.14 MULT=1
MM1025 N_A_1711_48#_M1025_d N_A_1511_74#_M1025_g N_VPWR_M1009_d VPB PSHORT
+ L=0.15 W=1 AD=0.285 AS=0.282746 PD=2.57 PS=2.23944 NRD=1.9503 NRS=35.4403 M=1
+ R=6.66667 SA=75001.8 SB=75000.2 A=0.15 P=2.3 MULT=1
MM1032 N_Q_M1032_d N_A_1711_48#_M1032_g N_VPWR_M1032_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.3192 PD=1.42 PS=2.81 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1034 N_Q_M1032_d N_A_1711_48#_M1034_g N_VPWR_M1034_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.3192 PD=1.42 PS=2.81 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.7 SB=75000.2 A=0.168 P=2.54 MULT=1
MM1039 N_VPWR_M1039_d N_A_1711_48#_M1039_g N_A_2322_368#_M1039_s VPB PSHORT
+ L=0.15 W=1 AD=0.193019 AS=0.285 PD=1.41038 PS=2.57 NRD=17.0602 NRS=1.9503 M=1
+ R=6.66667 SA=75000.2 SB=75001.2 A=0.15 P=2.3 MULT=1
MM1002 N_Q_N_M1002_d N_A_2322_368#_M1002_g N_VPWR_M1039_d VPB PSHORT L=0.15
+ W=1.12 AD=0.168 AS=0.216181 PD=1.42 PS=1.57962 NRD=1.7533 NRS=1.7533 M=1
+ R=7.46667 SA=75000.7 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1006 N_Q_N_M1002_d N_A_2322_368#_M1006_g N_VPWR_M1006_s VPB PSHORT L=0.15
+ W=1.12 AD=0.168 AS=0.3192 PD=1.42 PS=2.81 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.1 SB=75000.2 A=0.168 P=2.54 MULT=1
DX40_noxref VNB VPB NWDIODE A=25.7052 P=31.36
c_145 VNB 0 1.47924e-19 $X=0 $Y=0
*
.include "sky130_fd_sc_hs__sdfxbp_2.pxi.spice"
*
.ends
*
*
