* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hs__dlygate4sd3_1 A VGND VNB VPB VPWR X
M1000 a_289_74# a_28_74# VGND VNB nlowvt w=420000u l=180000u
+  ad=1.092e+11p pd=1.36e+06u as=5.279e+11p ps=4.43e+06u
M1001 VPWR a_289_74# a_405_138# VPB pshort w=1e+06u l=500000u
+  ad=6.905e+11p pd=5.7e+06u as=2.6e+11p ps=2.52e+06u
M1002 X a_405_138# VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=3.136e+11p pd=2.8e+06u as=0p ps=0u
M1003 a_289_74# a_28_74# VPWR VPB pshort w=1e+06u l=500000u
+  ad=2.6e+11p pd=2.52e+06u as=0p ps=0u
M1004 VGND A a_28_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1005 VGND a_289_74# a_405_138# VNB nlowvt w=420000u l=180000u
+  ad=0p pd=0u as=2.436e+11p ps=2e+06u
M1006 X a_405_138# VGND VNB nlowvt w=740000u l=150000u
+  ad=1.961e+11p pd=2.01e+06u as=0p ps=0u
M1007 VPWR A a_28_74# VPB pshort w=420000u l=150000u
+  ad=0p pd=0u as=1.176e+11p ps=1.4e+06u
.ends
