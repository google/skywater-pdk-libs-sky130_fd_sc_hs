* File: sky130_fd_sc_hs__sdfrtp_2.pex.spice
* Created: Tue Sep  1 20:22:45 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HS__SDFRTP_2%A_27_74# 1 2 7 9 11 12 14 17 20 23 27 30 32
+ 33 35 40
c80 35 0 1.02897e-20 $X=2.54 $Y=1.995
c81 9 0 3.56444e-20 $X=1.485 $Y=0.935
r82 35 38 3.31764 $w=3.28e-07 $l=9.5e-08 $layer=LI1_cond $X=2.54 $Y=1.995
+ $X2=2.54 $Y2=2.09
r83 35 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.54
+ $Y=1.995 $X2=2.54 $Y2=1.995
r84 31 33 2.76166 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.445 $Y=2.09
+ $X2=0.28 $Y2=2.09
r85 30 38 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.375 $Y=2.09
+ $X2=2.54 $Y2=2.09
r86 30 31 125.914 $w=1.68e-07 $l=1.93e-06 $layer=LI1_cond $X=2.375 $Y=2.09
+ $X2=0.445 $Y2=2.09
r87 28 40 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=0.975 $Y=1.1 $X2=0.975
+ $Y2=1.01
r88 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.975
+ $Y=1.1 $X2=0.975 $Y2=1.1
r89 25 32 0.221902 $w=3.3e-07 $l=1.25e-07 $layer=LI1_cond $X=0.365 $Y=1.1
+ $X2=0.24 $Y2=1.1
r90 25 27 21.3027 $w=3.28e-07 $l=6.1e-07 $layer=LI1_cond $X=0.365 $Y=1.1
+ $X2=0.975 $Y2=1.1
r91 21 33 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.28 $Y=2.175
+ $X2=0.28 $Y2=2.09
r92 21 23 10.1275 $w=3.28e-07 $l=2.9e-07 $layer=LI1_cond $X=0.28 $Y=2.175
+ $X2=0.28 $Y2=2.465
r93 20 33 3.70735 $w=2.5e-07 $l=1.18427e-07 $layer=LI1_cond $X=0.2 $Y=2.005
+ $X2=0.28 $Y2=2.09
r94 19 32 7.38875 $w=2.1e-07 $l=1.83916e-07 $layer=LI1_cond $X=0.2 $Y=1.265
+ $X2=0.24 $Y2=1.1
r95 19 20 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=0.2 $Y=1.265 $X2=0.2
+ $Y2=2.005
r96 15 32 7.38875 $w=2.1e-07 $l=1.65e-07 $layer=LI1_cond $X=0.24 $Y=0.935
+ $X2=0.24 $Y2=1.1
r97 15 17 16.3647 $w=2.48e-07 $l=3.55e-07 $layer=LI1_cond $X=0.24 $Y=0.935
+ $X2=0.24 $Y2=0.58
r98 12 36 52.2586 $w=2.99e-07 $l=2.7157e-07 $layer=POLY_cond $X=2.495 $Y=2.245
+ $X2=2.54 $Y2=1.995
r99 12 14 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=2.495 $Y=2.245
+ $X2=2.495 $Y2=2.64
r100 9 11 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.485 $Y=0.935
+ $X2=1.485 $Y2=0.615
r101 8 40 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.14 $Y=1.01
+ $X2=0.975 $Y2=1.01
r102 7 9 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.41 $Y=1.01
+ $X2=1.485 $Y2=0.935
r103 7 8 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=1.41 $Y=1.01 $X2=1.14
+ $Y2=1.01
r104 2 23 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=2.32 $X2=0.28 $Y2=2.465
r105 1 17 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_HS__SDFRTP_2%SCE 2 5 7 9 11 12 14 17 20 21 22 25 30 31
+ 32 45 47 56 58
r84 47 56 1.90404 $w=3.43e-07 $l=5.7e-08 $layer=LI1_cond $X=1.623 $Y=1.662
+ $X2=1.68 $Y2=1.662
r85 41 42 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.45
+ $Y=1.67 $X2=1.45 $Y2=1.67
r86 38 41 118.906 $w=3.3e-07 $l=6.8e-07 $layer=POLY_cond $X=0.77 $Y=1.67
+ $X2=1.45 $Y2=1.67
r87 32 58 6.34154 $w=3.43e-07 $l=1.01e-07 $layer=LI1_cond $X=1.694 $Y=1.662
+ $X2=1.795 $Y2=1.662
r88 32 56 0.467658 $w=3.43e-07 $l=1.4e-08 $layer=LI1_cond $X=1.694 $Y=1.662
+ $X2=1.68 $Y2=1.662
r89 32 47 0.467658 $w=3.43e-07 $l=1.4e-08 $layer=LI1_cond $X=1.609 $Y=1.662
+ $X2=1.623 $Y2=1.662
r90 32 42 5.31126 $w=3.43e-07 $l=1.59e-07 $layer=LI1_cond $X=1.609 $Y=1.662
+ $X2=1.45 $Y2=1.662
r91 31 42 8.35104 $w=3.43e-07 $l=2.5e-07 $layer=LI1_cond $X=1.2 $Y=1.662
+ $X2=1.45 $Y2=1.662
r92 30 31 16.034 $w=3.43e-07 $l=4.8e-07 $layer=LI1_cond $X=0.72 $Y=1.662 $X2=1.2
+ $Y2=1.662
r93 30 38 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=0.77
+ $Y=1.67 $X2=0.77 $Y2=1.67
r94 26 45 20.9834 $w=3.3e-07 $l=1.2e-07 $layer=POLY_cond $X=2.54 $Y=1.425
+ $X2=2.66 $Y2=1.425
r95 25 28 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=2.54 $Y=1.425
+ $X2=2.54 $Y2=1.575
r96 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.54
+ $Y=1.425 $X2=2.54 $Y2=1.425
r97 22 28 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.375 $Y=1.575
+ $X2=2.54 $Y2=1.575
r98 22 58 37.8396 $w=1.68e-07 $l=5.8e-07 $layer=LI1_cond $X=2.375 $Y=1.575
+ $X2=1.795 $Y2=1.575
r99 21 41 14.8632 $w=3.3e-07 $l=8.5e-08 $layer=POLY_cond $X=1.535 $Y=1.67
+ $X2=1.45 $Y2=1.67
r100 19 38 30.6007 $w=3.3e-07 $l=1.75e-07 $layer=POLY_cond $X=0.595 $Y=1.67
+ $X2=0.77 $Y2=1.67
r101 19 20 3.90195 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=0.595 $Y=1.67
+ $X2=0.505 $Y2=1.67
r102 15 45 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.66 $Y=1.26
+ $X2=2.66 $Y2=1.425
r103 15 17 330.734 $w=1.5e-07 $l=6.45e-07 $layer=POLY_cond $X=2.66 $Y=1.26
+ $X2=2.66 $Y2=0.615
r104 12 14 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=1.625 $Y=2.245
+ $X2=1.625 $Y2=2.64
r105 11 12 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=1.625 $Y=2.155
+ $X2=1.625 $Y2=2.245
r106 10 21 30.0773 $w=3.3e-07 $l=2.05122e-07 $layer=POLY_cond $X=1.625 $Y=1.835
+ $X2=1.535 $Y2=1.67
r107 10 11 124.387 $w=1.8e-07 $l=3.2e-07 $layer=POLY_cond $X=1.625 $Y=1.835
+ $X2=1.625 $Y2=2.155
r108 7 9 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=0.505 $Y=2.245
+ $X2=0.505 $Y2=2.64
r109 3 20 34.7346 $w=1.65e-07 $l=1.69926e-07 $layer=POLY_cond $X=0.495 $Y=1.505
+ $X2=0.505 $Y2=1.67
r110 3 5 474.309 $w=1.5e-07 $l=9.25e-07 $layer=POLY_cond $X=0.495 $Y=1.505
+ $X2=0.495 $Y2=0.58
r111 2 7 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=0.505 $Y=2.155
+ $X2=0.505 $Y2=2.245
r112 1 20 34.7346 $w=1.65e-07 $l=1.65e-07 $layer=POLY_cond $X=0.505 $Y=1.835
+ $X2=0.505 $Y2=1.67
r113 1 2 124.387 $w=1.8e-07 $l=3.2e-07 $layer=POLY_cond $X=0.505 $Y=1.835
+ $X2=0.505 $Y2=2.155
.ends

.subckt PM_SKY130_FD_SC_HS__SDFRTP_2%D 1 3 5 6 8 9 15 16
c45 6 0 1.02897e-20 $X=2.045 $Y=2.245
r46 14 16 19.2347 $w=3.3e-07 $l=1.1e-07 $layer=POLY_cond $X=1.935 $Y=1.1
+ $X2=2.045 $Y2=1.1
r47 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.935
+ $Y=1.1 $X2=1.935 $Y2=1.1
r48 11 14 10.4917 $w=3.3e-07 $l=6e-08 $layer=POLY_cond $X=1.875 $Y=1.1 $X2=1.935
+ $Y2=1.1
r49 9 15 6.7033 $w=4.53e-07 $l=2.55e-07 $layer=LI1_cond $X=1.68 $Y=1.037
+ $X2=1.935 $Y2=1.037
r50 6 8 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=2.045 $Y=2.245
+ $X2=2.045 $Y2=2.64
r51 5 6 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=2.045 $Y=2.155 $X2=2.045
+ $Y2=2.245
r52 4 16 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=2.045 $Y=1.265
+ $X2=2.045 $Y2=1.1
r53 4 5 345.952 $w=1.8e-07 $l=8.9e-07 $layer=POLY_cond $X=2.045 $Y=1.265
+ $X2=2.045 $Y2=2.155
r54 1 11 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.875 $Y=0.935
+ $X2=1.875 $Y2=1.1
r55 1 3 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.875 $Y=0.935
+ $X2=1.875 $Y2=0.615
.ends

.subckt PM_SKY130_FD_SC_HS__SDFRTP_2%SCD 1 3 6 10 11 12 16
r49 11 12 13.6198 $w=3.28e-07 $l=3.9e-07 $layer=LI1_cond $X=3.11 $Y=1.645
+ $X2=3.11 $Y2=2.035
r50 11 16 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.11
+ $Y=1.645 $X2=3.11 $Y2=1.645
r51 10 16 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=3.11 $Y=1.985
+ $X2=3.11 $Y2=1.645
r52 9 16 41.8716 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.11 $Y=1.48
+ $X2=3.11 $Y2=1.645
r53 6 9 443.543 $w=1.5e-07 $l=8.65e-07 $layer=POLY_cond $X=3.05 $Y=0.615
+ $X2=3.05 $Y2=1.48
r54 1 10 45.5709 $w=2.75e-07 $l=2.95127e-07 $layer=POLY_cond $X=3.035 $Y=2.245
+ $X2=3.11 $Y2=1.985
r55 1 3 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=3.035 $Y=2.245
+ $X2=3.035 $Y2=2.64
.ends

.subckt PM_SKY130_FD_SC_HS__SDFRTP_2%RESET_B 3 5 7 8 10 11 13 15 18 21 22 24 27
+ 29 30 31 32 39 40 43 46 48 54 65
c197 22 0 1.84389e-19 $X=11.35 $Y=2.465
c198 3 0 7.57672e-20 $X=3.595 $Y=0.615
r199 54 56 11.8137 $w=3.06e-07 $l=7.5e-08 $layer=POLY_cond $X=11.275 $Y=2.07
+ $X2=11.35 $Y2=2.07
r200 54 65 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=11.275
+ $Y=2.07 $X2=11.275 $Y2=2.07
r201 52 54 22.0523 $w=3.06e-07 $l=1.4e-07 $layer=POLY_cond $X=11.135 $Y=2.07
+ $X2=11.275 $Y2=2.07
r202 50 51 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.975
+ $Y=1.96 $X2=7.975 $Y2=1.96
r203 48 50 44.8056 $w=3.55e-07 $l=3.3e-07 $layer=POLY_cond $X=7.645 $Y=2.002
+ $X2=7.975 $Y2=2.002
r204 47 48 2.03662 $w=3.55e-07 $l=1.5e-08 $layer=POLY_cond $X=7.63 $Y=2.002
+ $X2=7.645 $Y2=2.002
r205 45 46 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.95
+ $Y=1.995 $X2=3.95 $Y2=1.995
r206 43 45 46.8423 $w=3.55e-07 $l=3.45e-07 $layer=POLY_cond $X=3.605 $Y=2.037
+ $X2=3.95 $Y2=2.037
r207 42 43 1.35775 $w=3.55e-07 $l=1e-08 $layer=POLY_cond $X=3.595 $Y=2.037
+ $X2=3.605 $Y2=2.037
r208 40 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.28 $Y=2.035
+ $X2=11.28 $Y2=2.035
r209 39 51 13.7969 $w=3.53e-07 $l=4.25e-07 $layer=LI1_cond $X=8.4 $Y=1.972
+ $X2=7.975 $Y2=1.972
r210 38 39 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=2.035
+ $X2=8.4 $Y2=2.035
r211 34 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=2.035
+ $X2=4.08 $Y2=2.035
r212 32 38 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=8.545 $Y=2.035
+ $X2=8.4 $Y2=2.035
r213 31 40 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=11.135 $Y=2.035
+ $X2=11.28 $Y2=2.035
r214 31 32 3.20544 $w=1.4e-07 $l=2.59e-06 $layer=MET1_cond $X=11.135 $Y=2.035
+ $X2=8.545 $Y2=2.035
r215 30 34 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.225 $Y=2.035
+ $X2=4.08 $Y2=2.035
r216 29 38 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=8.255 $Y=2.035
+ $X2=8.4 $Y2=2.035
r217 29 30 4.98761 $w=1.4e-07 $l=4.03e-06 $layer=MET1_cond $X=8.255 $Y=2.035
+ $X2=4.225 $Y2=2.035
r218 25 27 87.1702 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=7.475 $Y=1.26
+ $X2=7.645 $Y2=1.26
r219 22 24 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=11.35 $Y=2.465
+ $X2=11.35 $Y2=2.75
r220 21 22 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=11.35 $Y=2.375
+ $X2=11.35 $Y2=2.465
r221 20 56 15.178 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=11.35 $Y=2.235
+ $X2=11.35 $Y2=2.07
r222 20 21 54.4194 $w=1.8e-07 $l=1.4e-07 $layer=POLY_cond $X=11.35 $Y=2.235
+ $X2=11.35 $Y2=2.375
r223 16 52 19.4347 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=11.135 $Y=1.905
+ $X2=11.135 $Y2=2.07
r224 16 18 679.415 $w=1.5e-07 $l=1.325e-06 $layer=POLY_cond $X=11.135 $Y=1.905
+ $X2=11.135 $Y2=0.58
r225 15 48 22.9692 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=7.645 $Y=1.795
+ $X2=7.645 $Y2=2.002
r226 14 27 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.645 $Y=1.335
+ $X2=7.645 $Y2=1.26
r227 14 15 235.872 $w=1.5e-07 $l=4.6e-07 $layer=POLY_cond $X=7.645 $Y=1.335
+ $X2=7.645 $Y2=1.795
r228 11 47 22.9692 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=7.63 $Y=2.21
+ $X2=7.63 $Y2=2.002
r229 11 13 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=7.63 $Y=2.21
+ $X2=7.63 $Y2=2.495
r230 8 25 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.475 $Y=1.185
+ $X2=7.475 $Y2=1.26
r231 8 10 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=7.475 $Y=1.185
+ $X2=7.475 $Y2=0.9
r232 5 43 22.9692 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=3.605 $Y=2.245
+ $X2=3.605 $Y2=2.037
r233 5 7 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=3.605 $Y=2.245
+ $X2=3.605 $Y2=2.64
r234 1 42 22.9692 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.595 $Y=1.83
+ $X2=3.595 $Y2=2.037
r235 1 3 623.011 $w=1.5e-07 $l=1.215e-06 $layer=POLY_cond $X=3.595 $Y=1.83
+ $X2=3.595 $Y2=0.615
.ends

.subckt PM_SKY130_FD_SC_HS__SDFRTP_2%CLK 1 3 6 9 12 15 22
c55 9 0 5.70693e-20 $X=4.555 $Y=1.425
c56 6 0 7.24462e-20 $X=4.69 $Y=0.74
r57 15 22 3.70473 $w=4.08e-07 $l=1.15e-07 $layer=LI1_cond $X=4.08 $Y=1.385
+ $X2=4.195 $Y2=1.385
r58 12 22 9.95292 $w=3.28e-07 $l=2.85e-07 $layer=LI1_cond $X=4.48 $Y=1.425
+ $X2=4.195 $Y2=1.425
r59 12 13 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.48
+ $Y=1.425 $X2=4.48 $Y2=1.425
r60 9 13 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=4.555 $Y=1.425
+ $X2=4.48 $Y2=1.425
r61 4 9 42.9986 $w=1.99e-07 $l=1.79374e-07 $layer=POLY_cond $X=4.69 $Y=1.26
+ $X2=4.66 $Y2=1.425
r62 4 6 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=4.69 $Y=1.26 $X2=4.69
+ $Y2=0.74
r63 1 9 85.3855 $w=1.99e-07 $l=3.47419e-07 $layer=POLY_cond $X=4.645 $Y=1.765
+ $X2=4.66 $Y2=1.425
r64 1 3 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=4.645 $Y=1.765
+ $X2=4.645 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_HS__SDFRTP_2%A_1034_368# 1 2 8 9 11 12 14 16 18 20 21 22
+ 23 25 30 32 33 34 37 40 43 44 45 47 48 49 52 55 58 61 62 66
c202 61 0 1.4646e-20 $X=5.442 $Y=1.125
c203 52 0 8.16714e-20 $X=9.645 $Y=1.17
c204 49 0 6.41644e-20 $X=9.26 $Y=1.17
c205 48 0 1.18082e-19 $X=9.785 $Y=1.17
c206 34 0 5.78002e-20 $X=5.645 $Y=0.415
c207 23 0 4.68929e-20 $X=10.11 $Y=2.465
c208 21 0 2.95884e-20 $X=9.48 $Y=1.26
r209 62 64 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=7.125 $Y=0.415
+ $X2=7.125 $Y2=0.665
r210 58 60 9.55422 $w=3.32e-07 $l=2.6e-07 $layer=LI1_cond $X=5.4 $Y=1.8 $X2=5.4
+ $Y2=2.06
r211 55 56 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.95
+ $Y=2.165 $X2=9.95 $Y2=2.165
r212 53 55 36.0954 $w=2.63e-07 $l=8.3e-07 $layer=LI1_cond $X=9.917 $Y=1.335
+ $X2=9.917 $Y2=2.165
r213 52 72 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=9.645 $Y=1.17
+ $X2=9.645 $Y2=1.26
r214 51 52 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.645
+ $Y=1.17 $X2=9.645 $Y2=1.17
r215 49 51 13.4452 $w=3.28e-07 $l=3.85e-07 $layer=LI1_cond $X=9.26 $Y=1.17
+ $X2=9.645 $Y2=1.17
r216 48 53 6.92284 $w=3.3e-07 $l=2.21371e-07 $layer=LI1_cond $X=9.785 $Y=1.17
+ $X2=9.917 $Y2=1.335
r217 48 51 4.88915 $w=3.28e-07 $l=1.4e-07 $layer=LI1_cond $X=9.785 $Y=1.17
+ $X2=9.645 $Y2=1.17
r218 47 49 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=9.175 $Y=1.005
+ $X2=9.26 $Y2=1.17
r219 46 47 37.8396 $w=1.68e-07 $l=5.8e-07 $layer=LI1_cond $X=9.175 $Y=0.425
+ $X2=9.175 $Y2=1.005
r220 44 46 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.09 $Y=0.34
+ $X2=9.175 $Y2=0.425
r221 44 45 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=9.09 $Y=0.34
+ $X2=8.42 $Y2=0.34
r222 42 45 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.335 $Y=0.425
+ $X2=8.42 $Y2=0.34
r223 42 43 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=8.335 $Y=0.425
+ $X2=8.335 $Y2=0.58
r224 41 64 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.21 $Y=0.665
+ $X2=7.125 $Y2=0.665
r225 40 43 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.25 $Y=0.665
+ $X2=8.335 $Y2=0.58
r226 40 41 67.8503 $w=1.68e-07 $l=1.04e-06 $layer=LI1_cond $X=8.25 $Y=0.665
+ $X2=7.21 $Y2=0.665
r227 38 69 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.065 $Y=1.8
+ $X2=6.065 $Y2=1.965
r228 38 66 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=6.065 $Y=1.8
+ $X2=6.065 $Y2=1.71
r229 37 38 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.065
+ $Y=1.8 $X2=6.065 $Y2=1.8
r230 35 58 0.753319 $w=3.3e-07 $l=2.45e-07 $layer=LI1_cond $X=5.645 $Y=1.8
+ $X2=5.4 $Y2=1.8
r231 35 37 14.6675 $w=3.28e-07 $l=4.2e-07 $layer=LI1_cond $X=5.645 $Y=1.8
+ $X2=6.065 $Y2=1.8
r232 33 62 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.04 $Y=0.415
+ $X2=7.125 $Y2=0.415
r233 33 34 91.0107 $w=1.68e-07 $l=1.395e-06 $layer=LI1_cond $X=7.04 $Y=0.415
+ $X2=5.645 $Y2=0.415
r234 32 58 8.95967 $w=3.32e-07 $l=2.31571e-07 $layer=LI1_cond $X=5.56 $Y=1.635
+ $X2=5.4 $Y2=1.8
r235 32 61 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=5.56 $Y=1.635
+ $X2=5.56 $Y2=1.125
r236 28 61 9.72165 $w=4.03e-07 $l=2.02e-07 $layer=LI1_cond $X=5.442 $Y=0.923
+ $X2=5.442 $Y2=1.125
r237 28 30 11.6098 $w=4.03e-07 $l=4.08e-07 $layer=LI1_cond $X=5.442 $Y=0.923
+ $X2=5.442 $Y2=0.515
r238 27 34 8.41448 $w=1.7e-07 $l=2.41793e-07 $layer=LI1_cond $X=5.442 $Y=0.5
+ $X2=5.645 $Y2=0.415
r239 27 30 0.426831 $w=4.03e-07 $l=1.5e-08 $layer=LI1_cond $X=5.442 $Y=0.5
+ $X2=5.442 $Y2=0.515
r240 23 56 57.5457 $w=3.46e-07 $l=3.54119e-07 $layer=POLY_cond $X=10.11 $Y=2.465
+ $X2=9.992 $Y2=2.165
r241 23 25 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=10.11 $Y=2.465
+ $X2=10.11 $Y2=2.75
r242 21 72 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.48 $Y=1.26
+ $X2=9.645 $Y2=1.26
r243 21 22 184.596 $w=1.5e-07 $l=3.6e-07 $layer=POLY_cond $X=9.48 $Y=1.26
+ $X2=9.12 $Y2=1.26
r244 18 22 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=9.045 $Y=1.185
+ $X2=9.12 $Y2=1.26
r245 18 20 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=9.045 $Y=1.185
+ $X2=9.045 $Y2=0.74
r246 14 26 93.1232 $w=1.88e-07 $l=3.8151e-07 $layer=POLY_cond $X=6.695 $Y=1.355
+ $X2=6.64 $Y2=1.71
r247 14 16 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=6.695 $Y=1.355
+ $X2=6.695 $Y2=0.9
r248 13 66 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.23 $Y=1.71
+ $X2=6.065 $Y2=1.71
r249 12 26 8.14712 $w=1.5e-07 $l=1.3e-07 $layer=POLY_cond $X=6.51 $Y=1.71
+ $X2=6.64 $Y2=1.71
r250 12 13 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=6.51 $Y=1.71
+ $X2=6.23 $Y2=1.71
r251 9 11 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=6.135 $Y=2.21
+ $X2=6.135 $Y2=2.495
r252 8 9 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=6.135 $Y=2.12 $X2=6.135
+ $Y2=2.21
r253 8 69 60.25 $w=1.8e-07 $l=1.55e-07 $layer=POLY_cond $X=6.135 $Y=2.12
+ $X2=6.135 $Y2=1.965
r254 2 60 600 $w=1.7e-07 $l=2.85307e-07 $layer=licon1_PDIFF $count=1 $X=5.17
+ $Y=1.84 $X2=5.32 $Y2=2.06
r255 1 30 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=5.265
+ $Y=0.37 $X2=5.405 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__SDFRTP_2%A_1383_349# 1 2 7 9 12 16 19 20 25 28 33 34
c90 12 0 3.01223e-20 $X=7.085 $Y=0.9
r91 33 34 8.52431 $w=3.63e-07 $l=1.65e-07 $layer=LI1_cond $X=8.932 $Y=1.88
+ $X2=8.932 $Y2=1.715
r92 31 34 38.1658 $w=1.68e-07 $l=5.85e-07 $layer=LI1_cond $X=8.835 $Y=1.13
+ $X2=8.835 $Y2=1.715
r93 30 31 7.06528 $w=3.28e-07 $l=1.25e-07 $layer=LI1_cond $X=8.755 $Y=1.005
+ $X2=8.755 $Y2=1.13
r94 28 30 5.06376 $w=3.28e-07 $l=1.45e-07 $layer=LI1_cond $X=8.755 $Y=0.86
+ $X2=8.755 $Y2=1.005
r95 23 33 0.536754 $w=3.63e-07 $l=1.7e-08 $layer=LI1_cond $X=8.932 $Y=1.897
+ $X2=8.932 $Y2=1.88
r96 23 25 10.6719 $w=3.63e-07 $l=3.38e-07 $layer=LI1_cond $X=8.932 $Y=1.897
+ $X2=8.932 $Y2=2.235
r97 19 30 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.59 $Y=1.005
+ $X2=8.755 $Y2=1.005
r98 19 20 83.1818 $w=1.68e-07 $l=1.275e-06 $layer=LI1_cond $X=8.59 $Y=1.005
+ $X2=7.315 $Y2=1.005
r99 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.165
+ $Y=1.91 $X2=7.165 $Y2=1.91
r100 14 20 7.32204 $w=1.7e-07 $l=1.75425e-07 $layer=LI1_cond $X=7.177 $Y=1.09
+ $X2=7.315 $Y2=1.005
r101 14 16 34.3638 $w=2.73e-07 $l=8.2e-07 $layer=LI1_cond $X=7.177 $Y=1.09
+ $X2=7.177 $Y2=1.91
r102 10 17 38.7394 $w=3.46e-07 $l=1.82565e-07 $layer=POLY_cond $X=7.085 $Y=1.745
+ $X2=7.122 $Y2=1.91
r103 10 12 433.287 $w=1.5e-07 $l=8.45e-07 $layer=POLY_cond $X=7.085 $Y=1.745
+ $X2=7.085 $Y2=0.9
r104 7 17 57.5457 $w=3.46e-07 $l=3.53695e-07 $layer=POLY_cond $X=7.005 $Y=2.21
+ $X2=7.122 $Y2=1.91
r105 7 9 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=7.005 $Y=2.21
+ $X2=7.005 $Y2=2.495
r106 2 33 600 $w=1.7e-07 $l=2.98831e-07 $layer=licon1_PDIFF $count=1 $X=8.715
+ $Y=1.735 $X2=8.95 $Y2=1.88
r107 2 25 300 $w=1.7e-07 $l=6.06218e-07 $layer=licon1_PDIFF $count=2 $X=8.715
+ $Y=1.735 $X2=8.95 $Y2=2.235
r108 1 28 182 $w=1.7e-07 $l=5.55608e-07 $layer=licon1_NDIFF $count=1 $X=8.615
+ $Y=0.37 $X2=8.755 $Y2=0.86
.ends

.subckt PM_SKY130_FD_SC_HS__SDFRTP_2%A_1242_457# 1 2 3 12 14 16 18 19 24 25 28
+ 29 31 35 37
c120 28 0 1.23597e-19 $X=7.57 $Y=2.32
c121 24 0 6.99242e-20 $X=6.785 $Y=2.32
c122 12 0 6.41644e-20 $X=8.54 $Y=0.74
r123 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.255
+ $Y=1.41 $X2=8.255 $Y2=1.41
r124 29 31 21.9513 $w=3.13e-07 $l=6e-07 $layer=LI1_cond $X=7.655 $Y=1.417
+ $X2=8.255 $Y2=1.417
r125 28 40 11.0732 $w=3.14e-07 $l=3.72552e-07 $layer=LI1_cond $X=7.57 $Y=2.32
+ $X2=7.855 $Y2=2.522
r126 27 29 7.64049 $w=3.15e-07 $l=1.95944e-07 $layer=LI1_cond $X=7.57 $Y=1.575
+ $X2=7.655 $Y2=1.417
r127 27 28 48.6043 $w=1.68e-07 $l=7.45e-07 $layer=LI1_cond $X=7.57 $Y=1.575
+ $X2=7.57 $Y2=2.32
r128 26 37 4.3182 $w=2.1e-07 $l=1.53734e-07 $layer=LI1_cond $X=6.87 $Y=2.405
+ $X2=6.785 $Y2=2.522
r129 25 28 5.85116 $w=3.14e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.485 $Y=2.405
+ $X2=7.57 $Y2=2.32
r130 25 26 40.123 $w=1.68e-07 $l=6.15e-07 $layer=LI1_cond $X=7.485 $Y=2.405
+ $X2=6.87 $Y2=2.405
r131 24 37 2.11342 $w=1.7e-07 $l=2.02e-07 $layer=LI1_cond $X=6.785 $Y=2.32
+ $X2=6.785 $Y2=2.522
r132 23 35 10.9764 $w=3.39e-07 $l=4.03194e-07 $layer=LI1_cond $X=6.785 $Y=1.125
+ $X2=6.48 $Y2=0.897
r133 23 24 77.9626 $w=1.68e-07 $l=1.195e-06 $layer=LI1_cond $X=6.785 $Y=1.125
+ $X2=6.785 $Y2=2.32
r134 19 37 4.3182 $w=2.1e-07 $l=1.17707e-07 $layer=LI1_cond $X=6.7 $Y=2.6
+ $X2=6.785 $Y2=2.522
r135 19 21 15.6732 $w=2.48e-07 $l=3.4e-07 $layer=LI1_cond $X=6.7 $Y=2.6 $X2=6.36
+ $Y2=2.6
r136 18 32 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=8.465 $Y=1.41
+ $X2=8.255 $Y2=1.41
r137 14 18 64.0286 $w=1.97e-07 $l=2.70647e-07 $layer=POLY_cond $X=8.64 $Y=1.66
+ $X2=8.597 $Y2=1.41
r138 14 16 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=8.64 $Y=1.66
+ $X2=8.64 $Y2=2.235
r139 10 18 43.2316 $w=1.97e-07 $l=1.9139e-07 $layer=POLY_cond $X=8.54 $Y=1.245
+ $X2=8.597 $Y2=1.41
r140 10 12 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=8.54 $Y=1.245
+ $X2=8.54 $Y2=0.74
r141 3 40 600 $w=1.7e-07 $l=3.00791e-07 $layer=licon1_PDIFF $count=1 $X=7.705
+ $Y=2.285 $X2=7.855 $Y2=2.52
r142 2 21 600 $w=1.7e-07 $l=3.4187e-07 $layer=licon1_PDIFF $count=1 $X=6.21
+ $Y=2.285 $X2=6.36 $Y2=2.56
r143 1 35 182 $w=1.7e-07 $l=2.95212e-07 $layer=licon1_NDIFF $count=1 $X=6.27
+ $Y=0.69 $X2=6.48 $Y2=0.895
.ends

.subckt PM_SKY130_FD_SC_HS__SDFRTP_2%A_855_368# 1 2 7 9 12 14 17 18 20 21 24 26
+ 27 28 30 31 36 37 38 40 43 45 46 47 51 55 57 58 59 62 64 65 73
c197 62 0 1.84505e-19 $X=4.9 $Y=1.295
c198 18 0 6.99242e-20 $X=6.12 $Y=1.32
r199 74 76 23.3495 $w=2.89e-07 $l=1.4e-07 $layer=POLY_cond $X=5.14 $Y=1.46
+ $X2=5.14 $Y2=1.32
r200 73 74 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.14
+ $Y=1.46 $X2=5.14 $Y2=1.46
r201 70 73 8.3814 $w=3.28e-07 $l=2.4e-07 $layer=LI1_cond $X=4.9 $Y=1.46 $X2=5.14
+ $Y2=1.46
r202 65 68 5.30124 $w=2.48e-07 $l=1.15e-07 $layer=LI1_cond $X=4.46 $Y=1.905
+ $X2=4.46 $Y2=2.02
r203 63 70 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.9 $Y=1.625
+ $X2=4.9 $Y2=1.46
r204 63 64 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=4.9 $Y=1.625
+ $X2=4.9 $Y2=1.82
r205 62 70 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.9 $Y=1.295
+ $X2=4.9 $Y2=1.46
r206 61 62 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=4.9 $Y=1.09
+ $X2=4.9 $Y2=1.295
r207 60 65 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.585 $Y=1.905
+ $X2=4.46 $Y2=1.905
r208 59 64 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.815 $Y=1.905
+ $X2=4.9 $Y2=1.82
r209 59 60 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=4.815 $Y=1.905
+ $X2=4.585 $Y2=1.905
r210 57 61 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.815 $Y=1.005
+ $X2=4.9 $Y2=1.09
r211 57 58 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=4.815 $Y=1.005
+ $X2=4.56 $Y2=1.005
r212 53 58 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.475 $Y=0.92
+ $X2=4.56 $Y2=1.005
r213 53 55 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=4.475 $Y=0.92
+ $X2=4.475 $Y2=0.515
r214 49 51 97.4255 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=10.125 $Y=1.055
+ $X2=10.315 $Y2=1.055
r215 41 51 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=10.315 $Y=0.98
+ $X2=10.315 $Y2=1.055
r216 41 43 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=10.315 $Y=0.98
+ $X2=10.315 $Y2=0.58
r217 39 49 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=10.125 $Y=1.13
+ $X2=10.125 $Y2=1.055
r218 39 40 228.181 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=10.125 $Y=1.13
+ $X2=10.125 $Y2=1.575
r219 37 40 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=10.05 $Y=1.65
+ $X2=10.125 $Y2=1.575
r220 37 38 358.936 $w=1.5e-07 $l=7e-07 $layer=POLY_cond $X=10.05 $Y=1.65
+ $X2=9.35 $Y2=1.65
r221 34 47 97.3837 $w=1.8e-07 $l=2.45e-07 $layer=POLY_cond $X=9.26 $Y=2.905
+ $X2=9.26 $Y2=3.15
r222 34 36 294.84 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=9.26 $Y=2.905
+ $X2=9.26 $Y2=2.33
r223 33 38 26.9307 $w=1.5e-07 $l=1.43091e-07 $layer=POLY_cond $X=9.26 $Y=1.755
+ $X2=9.35 $Y2=1.65
r224 33 36 294.84 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=9.26 $Y=1.755
+ $X2=9.26 $Y2=2.33
r225 32 46 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=6.675 $Y=3.15
+ $X2=6.585 $Y2=3.15
r226 31 47 7.1379 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=9.17 $Y=3.15 $X2=9.26
+ $Y2=3.15
r227 31 32 1279.35 $w=1.5e-07 $l=2.495e-06 $layer=POLY_cond $X=9.17 $Y=3.15
+ $X2=6.675 $Y2=3.15
r228 28 30 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=6.585 $Y=2.78
+ $X2=6.585 $Y2=2.495
r229 27 46 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=6.585 $Y=3.075
+ $X2=6.585 $Y2=3.15
r230 26 28 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=6.585 $Y=2.87
+ $X2=6.585 $Y2=2.78
r231 26 27 79.6855 $w=1.8e-07 $l=2.05e-07 $layer=POLY_cond $X=6.585 $Y=2.87
+ $X2=6.585 $Y2=3.075
r232 22 24 176.904 $w=1.5e-07 $l=3.45e-07 $layer=POLY_cond $X=6.195 $Y=1.245
+ $X2=6.195 $Y2=0.9
r233 20 46 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=6.495 $Y=3.15
+ $X2=6.585 $Y2=3.15
r234 20 21 412.777 $w=1.5e-07 $l=8.05e-07 $layer=POLY_cond $X=6.495 $Y=3.15
+ $X2=5.69 $Y2=3.15
r235 19 45 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.69 $Y=1.32
+ $X2=5.615 $Y2=1.32
r236 18 22 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=6.12 $Y=1.32
+ $X2=6.195 $Y2=1.245
r237 18 19 220.489 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=6.12 $Y=1.32
+ $X2=5.69 $Y2=1.32
r238 17 21 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.615 $Y=3.075
+ $X2=5.69 $Y2=3.15
r239 16 45 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.615 $Y=1.395
+ $X2=5.615 $Y2=1.32
r240 16 17 861.447 $w=1.5e-07 $l=1.68e-06 $layer=POLY_cond $X=5.615 $Y=1.395
+ $X2=5.615 $Y2=3.075
r241 15 76 18.0918 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.305 $Y=1.32
+ $X2=5.14 $Y2=1.32
r242 14 45 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.54 $Y=1.32
+ $X2=5.615 $Y2=1.32
r243 14 15 120.5 $w=1.5e-07 $l=2.35e-07 $layer=POLY_cond $X=5.54 $Y=1.32
+ $X2=5.305 $Y2=1.32
r244 10 76 23.6143 $w=2.89e-07 $l=9.68246e-08 $layer=POLY_cond $X=5.19 $Y=1.245
+ $X2=5.14 $Y2=1.32
r245 10 12 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=5.19 $Y=1.245
+ $X2=5.19 $Y2=0.74
r246 7 74 61.9742 $w=2.89e-07 $l=3.26726e-07 $layer=POLY_cond $X=5.095 $Y=1.765
+ $X2=5.14 $Y2=1.46
r247 7 9 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=5.095 $Y=1.765
+ $X2=5.095 $Y2=2.4
r248 2 68 600 $w=1.7e-07 $l=2.41868e-07 $layer=licon1_PDIFF $count=1 $X=4.275
+ $Y=1.84 $X2=4.42 $Y2=2.02
r249 1 55 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=4.33
+ $Y=0.37 $X2=4.475 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__SDFRTP_2%A_2082_446# 1 2 7 9 12 14 18 19 20 22 23 26
+ 30 32 33 35 37 38
c122 23 0 4.68929e-20 $X=10.85 $Y=2.475
c123 18 0 2.97873e-19 $X=10.685 $Y=2.215
c124 12 0 1.18082e-19 $X=10.705 $Y=0.58
r125 38 41 5.42589 $w=4.1e-07 $l=4e-08 $layer=POLY_cond $X=10.645 $Y=1.535
+ $X2=10.645 $Y2=1.575
r126 38 44 45.9078 $w=4.1e-07 $l=1.65e-07 $layer=POLY_cond $X=10.645 $Y=1.535
+ $X2=10.645 $Y2=1.37
r127 37 40 5.16612 $w=2.88e-07 $l=1.3e-07 $layer=LI1_cond $X=10.705 $Y=1.535
+ $X2=10.705 $Y2=1.665
r128 37 38 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=10.685
+ $Y=1.535 $X2=10.685 $Y2=1.535
r129 34 35 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=12.145 $Y=0.94
+ $X2=12.145 $Y2=1.58
r130 32 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=12.06 $Y=0.855
+ $X2=12.145 $Y2=0.94
r131 32 33 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=12.06 $Y=0.855
+ $X2=11.875 $Y2=0.855
r132 28 33 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=11.71 $Y=0.77
+ $X2=11.875 $Y2=0.855
r133 28 30 6.63528 $w=3.28e-07 $l=1.9e-07 $layer=LI1_cond $X=11.71 $Y=0.77
+ $X2=11.71 $Y2=0.58
r134 24 26 6.63528 $w=3.28e-07 $l=1.9e-07 $layer=LI1_cond $X=11.575 $Y=2.56
+ $X2=11.575 $Y2=2.75
r135 22 24 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=11.41 $Y=2.475
+ $X2=11.575 $Y2=2.56
r136 22 23 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=11.41 $Y=2.475
+ $X2=10.85 $Y2=2.475
r137 21 40 3.86198 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=10.85 $Y=1.665
+ $X2=10.705 $Y2=1.665
r138 20 35 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=12.06 $Y=1.665
+ $X2=12.145 $Y2=1.58
r139 20 21 78.9412 $w=1.68e-07 $l=1.21e-06 $layer=LI1_cond $X=12.06 $Y=1.665
+ $X2=10.85 $Y2=1.665
r140 19 41 86.8143 $w=4.1e-07 $l=6.4e-07 $layer=POLY_cond $X=10.645 $Y=2.215
+ $X2=10.645 $Y2=1.575
r141 18 19 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=10.685
+ $Y=2.215 $X2=10.685 $Y2=2.215
r142 16 23 7.43784 $w=1.7e-07 $l=1.8262e-07 $layer=LI1_cond $X=10.705 $Y=2.39
+ $X2=10.85 $Y2=2.475
r143 16 18 6.9544 $w=2.88e-07 $l=1.75e-07 $layer=LI1_cond $X=10.705 $Y=2.39
+ $X2=10.705 $Y2=2.215
r144 15 40 3.37785 $w=2.88e-07 $l=8.5e-08 $layer=LI1_cond $X=10.705 $Y=1.75
+ $X2=10.705 $Y2=1.665
r145 15 18 18.4788 $w=2.88e-07 $l=4.65e-07 $layer=LI1_cond $X=10.705 $Y=1.75
+ $X2=10.705 $Y2=2.215
r146 14 19 2.03471 $w=4.1e-07 $l=1.5e-08 $layer=POLY_cond $X=10.645 $Y=2.23
+ $X2=10.645 $Y2=2.215
r147 12 44 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=10.705 $Y=0.58
+ $X2=10.705 $Y2=1.37
r148 7 14 32.8319 $w=3.45e-07 $l=2.98831e-07 $layer=POLY_cond $X=10.5 $Y=2.465
+ $X2=10.645 $Y2=2.23
r149 7 9 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=10.5 $Y=2.465 $X2=10.5
+ $Y2=2.75
r150 2 26 600 $w=1.7e-07 $l=2.74955e-07 $layer=licon1_PDIFF $count=1 $X=11.425
+ $Y=2.54 $X2=11.575 $Y2=2.75
r151 1 30 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=11.57
+ $Y=0.37 $X2=11.71 $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_HS__SDFRTP_2%A_1824_74# 1 2 9 11 12 13 15 18 19 21 22 24
+ 25 27 28 29 32 34 38 39 43 45 50 53 54 55
c144 53 0 6.53658e-20 $X=10.305 $Y=1.115
c145 43 0 1.63056e-20 $X=10.305 $Y=1.03
c146 32 0 2.95884e-20 $X=9.485 $Y=2.005
c147 28 0 6.36774e-20 $X=11.8 $Y=1.665
r148 54 55 8.67671 $w=2.98e-07 $l=1.7e-07 $layer=LI1_cond $X=11.02 $Y=1.22
+ $X2=11.19 $Y2=1.22
r149 51 58 15.7174 $w=2.76e-07 $l=9e-08 $layer=POLY_cond $X=11.725 $Y=1.26
+ $X2=11.815 $Y2=1.26
r150 50 55 20.5519 $w=2.98e-07 $l=5.35e-07 $layer=LI1_cond $X=11.725 $Y=1.26
+ $X2=11.19 $Y2=1.26
r151 50 51 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=11.725
+ $Y=1.26 $X2=11.725 $Y2=1.26
r152 47 53 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.39 $Y=1.115
+ $X2=10.305 $Y2=1.115
r153 47 54 41.1016 $w=1.68e-07 $l=6.3e-07 $layer=LI1_cond $X=10.39 $Y=1.115
+ $X2=11.02 $Y2=1.115
r154 44 53 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.305 $Y=1.2
+ $X2=10.305 $Y2=1.115
r155 44 45 86.1176 $w=1.68e-07 $l=1.32e-06 $layer=LI1_cond $X=10.305 $Y=1.2
+ $X2=10.305 $Y2=2.52
r156 43 53 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.305 $Y=1.03
+ $X2=10.305 $Y2=1.115
r157 42 43 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=10.305 $Y=0.81
+ $X2=10.305 $Y2=1.03
r158 39 41 9.95292 $w=3.28e-07 $l=2.85e-07 $layer=LI1_cond $X=9.6 $Y=2.685
+ $X2=9.885 $Y2=2.685
r159 38 45 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=10.22 $Y=2.685
+ $X2=10.305 $Y2=2.52
r160 38 41 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=10.22 $Y=2.685
+ $X2=9.885 $Y2=2.685
r161 34 42 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=10.22 $Y=0.645
+ $X2=10.305 $Y2=0.81
r162 34 36 4.1907 $w=3.28e-07 $l=1.2e-07 $layer=LI1_cond $X=10.22 $Y=0.645
+ $X2=10.1 $Y2=0.645
r163 30 39 6.87623 $w=3.3e-07 $l=2.24332e-07 $layer=LI1_cond $X=9.46 $Y=2.52
+ $X2=9.6 $Y2=2.685
r164 30 32 21.1967 $w=2.78e-07 $l=5.15e-07 $layer=LI1_cond $X=9.46 $Y=2.52
+ $X2=9.46 $Y2=2.005
r165 25 29 34.7346 $w=1.65e-07 $l=1.9e-07 $layer=POLY_cond $X=12.485 $Y=1.095
+ $X2=12.295 $Y2=1.095
r166 25 27 130.14 $w=1.5e-07 $l=4.05e-07 $layer=POLY_cond $X=12.485 $Y=1.095
+ $X2=12.485 $Y2=0.69
r167 22 24 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=12.385 $Y=1.885
+ $X2=12.385 $Y2=2.46
r168 21 22 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=12.385 $Y=1.795
+ $X2=12.385 $Y2=1.885
r169 20 29 34.7346 $w=1.65e-07 $l=3.7229e-07 $layer=POLY_cond $X=12.385 $Y=1.425
+ $X2=12.295 $Y2=1.095
r170 20 21 143.823 $w=1.8e-07 $l=3.7e-07 $layer=POLY_cond $X=12.385 $Y=1.425
+ $X2=12.385 $Y2=1.795
r171 19 58 12.3868 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=11.89 $Y=1.26
+ $X2=11.815 $Y2=1.26
r172 18 29 3.90195 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=12.295 $Y=1.26
+ $X2=12.295 $Y2=1.095
r173 18 19 70.8188 $w=3.3e-07 $l=4.05e-07 $layer=POLY_cond $X=12.295 $Y=1.26
+ $X2=11.89 $Y2=1.26
r174 16 58 17.0164 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=11.815 $Y=1.425
+ $X2=11.815 $Y2=1.26
r175 16 28 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=11.815 $Y=1.425
+ $X2=11.815 $Y2=1.665
r176 13 15 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=11.8 $Y=2.465
+ $X2=11.8 $Y2=2.75
r177 12 13 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=11.8 $Y=2.375
+ $X2=11.8 $Y2=2.465
r178 11 28 37.1337 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=11.8 $Y=1.755
+ $X2=11.8 $Y2=1.665
r179 11 12 241 $w=1.8e-07 $l=6.2e-07 $layer=POLY_cond $X=11.8 $Y=1.755 $X2=11.8
+ $Y2=2.375
r180 7 51 40.1667 $w=2.76e-07 $l=3.01413e-07 $layer=POLY_cond $X=11.495 $Y=1.095
+ $X2=11.725 $Y2=1.26
r181 7 9 264.074 $w=1.5e-07 $l=5.15e-07 $layer=POLY_cond $X=11.495 $Y=1.095
+ $X2=11.495 $Y2=0.58
r182 2 41 300 $w=1.7e-07 $l=1.09603e-06 $layer=licon1_PDIFF $count=2 $X=9.335
+ $Y=1.83 $X2=9.885 $Y2=2.685
r183 2 32 300 $w=1.7e-07 $l=2.38485e-07 $layer=licon1_PDIFF $count=2 $X=9.335
+ $Y=1.83 $X2=9.485 $Y2=2.005
r184 1 36 91 $w=1.7e-07 $l=1.10901e-06 $layer=licon1_NDIFF $count=2 $X=9.12
+ $Y=0.37 $X2=10.1 $Y2=0.645
.ends

.subckt PM_SKY130_FD_SC_HS__SDFRTP_2%A_2492_392# 1 2 7 9 12 14 16 19 23 25 29 35
+ 38 39 43
r62 43 44 7.77419 $w=3.72e-07 $l=6e-08 $layer=POLY_cond $X=13.845 $Y=1.532
+ $X2=13.905 $Y2=1.532
r63 42 43 47.9409 $w=3.72e-07 $l=3.7e-07 $layer=POLY_cond $X=13.475 $Y=1.532
+ $X2=13.845 $Y2=1.532
r64 41 42 10.3656 $w=3.72e-07 $l=8e-08 $layer=POLY_cond $X=13.395 $Y=1.532
+ $X2=13.475 $Y2=1.532
r65 36 41 26.5618 $w=3.72e-07 $l=2.05e-07 $layer=POLY_cond $X=13.19 $Y=1.532
+ $X2=13.395 $Y2=1.532
r66 35 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=13.19
+ $Y=1.465 $X2=13.19 $Y2=1.465
r67 33 39 0.144206 $w=3.3e-07 $l=1.3e-07 $layer=LI1_cond $X=12.865 $Y=1.465
+ $X2=12.735 $Y2=1.465
r68 33 35 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=12.865 $Y=1.465
+ $X2=13.19 $Y2=1.465
r69 31 39 7.25953 $w=2.15e-07 $l=1.86145e-07 $layer=LI1_cond $X=12.69 $Y=1.63
+ $X2=12.735 $Y2=1.465
r70 31 38 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=12.69 $Y=1.63
+ $X2=12.69 $Y2=1.94
r71 27 39 7.25953 $w=2.15e-07 $l=1.65e-07 $layer=LI1_cond $X=12.735 $Y=1.3
+ $X2=12.735 $Y2=1.465
r72 27 29 34.7949 $w=2.58e-07 $l=7.85e-07 $layer=LI1_cond $X=12.735 $Y=1.3
+ $X2=12.735 $Y2=0.515
r73 23 38 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=12.61 $Y=2.105
+ $X2=12.61 $Y2=1.94
r74 23 25 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=12.61 $Y=2.105
+ $X2=12.61 $Y2=2.815
r75 17 44 24.0971 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=13.905 $Y=1.3
+ $X2=13.905 $Y2=1.532
r76 17 19 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=13.905 $Y=1.3
+ $X2=13.905 $Y2=0.74
r77 14 43 24.0971 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=13.845 $Y=1.765
+ $X2=13.845 $Y2=1.532
r78 14 16 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=13.845 $Y=1.765
+ $X2=13.845 $Y2=2.4
r79 10 42 24.0971 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=13.475 $Y=1.3
+ $X2=13.475 $Y2=1.532
r80 10 12 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=13.475 $Y=1.3
+ $X2=13.475 $Y2=0.74
r81 7 41 24.0971 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=13.395 $Y=1.765
+ $X2=13.395 $Y2=1.532
r82 7 9 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=13.395 $Y=1.765
+ $X2=13.395 $Y2=2.4
r83 2 25 400 $w=1.7e-07 $l=9.26971e-07 $layer=licon1_PDIFF $count=1 $X=12.46
+ $Y=1.96 $X2=12.61 $Y2=2.815
r84 2 23 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=12.46
+ $Y=1.96 $X2=12.61 $Y2=2.105
r85 1 29 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=12.56
+ $Y=0.37 $X2=12.7 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__SDFRTP_2%VPWR 1 2 3 4 5 6 7 8 9 30 34 38 42 46 52 56
+ 58 63 64 66 67 69 70 71 73 78 96 100 112 116 122 129 132 135 142 146
c175 4 0 1.23597e-19 $X=7.08 $Y=2.285
c176 2 0 1.19423e-19 $X=3.11 $Y=2.32
r177 145 146 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=14.16 $Y=3.33
+ $X2=14.16 $Y2=3.33
r178 142 143 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.2 $Y=3.33
+ $X2=13.2 $Y2=3.33
r179 138 139 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.8 $Y=3.33
+ $X2=10.8 $Y2=3.33
r180 135 138 9.05853 $w=6.78e-07 $l=5.15e-07 $layer=LI1_cond $X=10.9 $Y=2.815
+ $X2=10.9 $Y2=3.33
r181 132 133 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=3.33
+ $X2=8.4 $Y2=3.33
r182 129 130 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r183 125 126 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r184 122 125 11.1084 $w=9.48e-07 $l=8.65e-07 $layer=LI1_cond $X=1.09 $Y=2.465
+ $X2=1.09 $Y2=3.33
r185 120 146 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=13.68 $Y=3.33
+ $X2=14.16 $Y2=3.33
r186 120 143 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=13.68 $Y=3.33
+ $X2=13.2 $Y2=3.33
r187 119 120 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.68 $Y=3.33
+ $X2=13.68 $Y2=3.33
r188 117 142 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=13.335 $Y=3.33
+ $X2=13.17 $Y2=3.33
r189 117 119 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=13.335 $Y=3.33
+ $X2=13.68 $Y2=3.33
r190 116 145 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=13.955 $Y=3.33
+ $X2=14.177 $Y2=3.33
r191 116 119 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=13.955 $Y=3.33
+ $X2=13.68 $Y2=3.33
r192 115 143 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.72 $Y=3.33
+ $X2=13.2 $Y2=3.33
r193 114 115 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=12.72 $Y=3.33
+ $X2=12.72 $Y2=3.33
r194 112 142 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=13.005 $Y=3.33
+ $X2=13.17 $Y2=3.33
r195 112 114 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=13.005 $Y=3.33
+ $X2=12.72 $Y2=3.33
r196 111 115 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=11.76 $Y=3.33
+ $X2=12.72 $Y2=3.33
r197 111 139 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=11.76 $Y=3.33
+ $X2=10.8 $Y2=3.33
r198 110 111 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=11.76 $Y=3.33
+ $X2=11.76 $Y2=3.33
r199 108 138 9.13095 $w=1.7e-07 $l=3.4e-07 $layer=LI1_cond $X=11.24 $Y=3.33
+ $X2=10.9 $Y2=3.33
r200 108 110 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=11.24 $Y=3.33
+ $X2=11.76 $Y2=3.33
r201 107 139 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.32 $Y=3.33
+ $X2=10.8 $Y2=3.33
r202 106 107 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.32 $Y=3.33
+ $X2=10.32 $Y2=3.33
r203 104 107 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=8.88 $Y=3.33
+ $X2=10.32 $Y2=3.33
r204 104 133 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=3.33
+ $X2=8.4 $Y2=3.33
r205 103 106 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=8.88 $Y=3.33
+ $X2=10.32 $Y2=3.33
r206 103 104 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r207 101 132 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.58 $Y=3.33
+ $X2=8.415 $Y2=3.33
r208 101 103 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=8.58 $Y=3.33
+ $X2=8.88 $Y2=3.33
r209 100 138 9.13095 $w=1.7e-07 $l=3.4e-07 $layer=LI1_cond $X=10.56 $Y=3.33
+ $X2=10.9 $Y2=3.33
r210 100 106 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=10.56 $Y=3.33
+ $X2=10.32 $Y2=3.33
r211 99 133 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=3.33
+ $X2=8.4 $Y2=3.33
r212 98 99 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r213 96 132 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.25 $Y=3.33
+ $X2=8.415 $Y2=3.33
r214 96 98 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=8.25 $Y=3.33
+ $X2=7.92 $Y2=3.33
r215 94 95 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r216 92 95 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=6.96 $Y2=3.33
r217 91 94 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=5.04 $Y=3.33
+ $X2=6.96 $Y2=3.33
r218 91 92 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r219 89 92 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=5.04 $Y2=3.33
r220 88 89 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r221 86 89 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.56 $Y2=3.33
r222 86 130 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=3.12 $Y2=3.33
r223 85 88 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=3.6 $Y=3.33 $X2=4.56
+ $Y2=3.33
r224 85 86 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r225 83 129 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.425 $Y=3.33
+ $X2=3.26 $Y2=3.33
r226 83 85 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=3.425 $Y=3.33
+ $X2=3.6 $Y2=3.33
r227 82 130 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=3.12 $Y2=3.33
r228 82 126 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r229 81 82 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r230 79 125 11.3727 $w=1.7e-07 $l=4.75e-07 $layer=LI1_cond $X=1.565 $Y=3.33
+ $X2=1.09 $Y2=3.33
r231 79 81 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=1.565 $Y=3.33
+ $X2=1.68 $Y2=3.33
r232 78 129 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.095 $Y=3.33
+ $X2=3.26 $Y2=3.33
r233 78 81 92.3155 $w=1.68e-07 $l=1.415e-06 $layer=LI1_cond $X=3.095 $Y=3.33
+ $X2=1.68 $Y2=3.33
r234 76 126 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=1.2 $Y2=3.33
r235 75 76 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r236 73 125 11.3727 $w=1.7e-07 $l=4.75e-07 $layer=LI1_cond $X=0.615 $Y=3.33
+ $X2=1.09 $Y2=3.33
r237 73 75 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=0.615 $Y=3.33
+ $X2=0.24 $Y2=3.33
r238 71 99 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=7.2 $Y=3.33
+ $X2=7.92 $Y2=3.33
r239 71 95 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=7.2 $Y=3.33
+ $X2=6.96 $Y2=3.33
r240 69 110 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=11.945 $Y=3.33
+ $X2=11.76 $Y2=3.33
r241 69 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.945 $Y=3.33
+ $X2=12.11 $Y2=3.33
r242 68 114 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=12.275 $Y=3.33
+ $X2=12.72 $Y2=3.33
r243 68 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12.275 $Y=3.33
+ $X2=12.11 $Y2=3.33
r244 66 94 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=7.15 $Y=3.33
+ $X2=6.96 $Y2=3.33
r245 66 67 8.70163 $w=1.7e-07 $l=1.67e-07 $layer=LI1_cond $X=7.15 $Y=3.33
+ $X2=7.317 $Y2=3.33
r246 65 98 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=7.485 $Y=3.33
+ $X2=7.92 $Y2=3.33
r247 65 67 8.70163 $w=1.7e-07 $l=1.68e-07 $layer=LI1_cond $X=7.485 $Y=3.33
+ $X2=7.317 $Y2=3.33
r248 63 88 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=4.705 $Y=3.33
+ $X2=4.56 $Y2=3.33
r249 63 64 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.705 $Y=3.33
+ $X2=4.87 $Y2=3.33
r250 62 91 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=5.035 $Y=3.33
+ $X2=5.04 $Y2=3.33
r251 62 64 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.035 $Y=3.33
+ $X2=4.87 $Y2=3.33
r252 58 61 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=14.12 $Y=1.985
+ $X2=14.12 $Y2=2.815
r253 56 145 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=14.12 $Y=3.245
+ $X2=14.177 $Y2=3.33
r254 56 61 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=14.12 $Y=3.245
+ $X2=14.12 $Y2=2.815
r255 52 55 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=13.17 $Y=1.985
+ $X2=13.17 $Y2=2.815
r256 50 142 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=13.17 $Y=3.245
+ $X2=13.17 $Y2=3.33
r257 50 55 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=13.17 $Y=3.245
+ $X2=13.17 $Y2=2.815
r258 46 49 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=12.11 $Y=2.105
+ $X2=12.11 $Y2=2.815
r259 44 70 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=12.11 $Y=3.245
+ $X2=12.11 $Y2=3.33
r260 44 49 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=12.11 $Y=3.245
+ $X2=12.11 $Y2=2.815
r261 40 132 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.415 $Y=3.245
+ $X2=8.415 $Y2=3.33
r262 40 42 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=8.415 $Y=3.245
+ $X2=8.415 $Y2=2.535
r263 36 67 0.942324 $w=3.35e-07 $l=8.5e-08 $layer=LI1_cond $X=7.317 $Y=3.245
+ $X2=7.317 $Y2=3.33
r264 36 38 14.4485 $w=3.33e-07 $l=4.2e-07 $layer=LI1_cond $X=7.317 $Y=3.245
+ $X2=7.317 $Y2=2.825
r265 32 64 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.87 $Y=3.245
+ $X2=4.87 $Y2=3.33
r266 32 34 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=4.87 $Y=3.245
+ $X2=4.87 $Y2=2.815
r267 28 129 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.26 $Y=3.245
+ $X2=3.26 $Y2=3.33
r268 28 30 15.8897 $w=3.28e-07 $l=4.55e-07 $layer=LI1_cond $X=3.26 $Y=3.245
+ $X2=3.26 $Y2=2.79
r269 9 61 400 $w=1.7e-07 $l=1.07034e-06 $layer=licon1_PDIFF $count=1 $X=13.92
+ $Y=1.84 $X2=14.12 $Y2=2.815
r270 9 58 400 $w=1.7e-07 $l=2.62678e-07 $layer=licon1_PDIFF $count=1 $X=13.92
+ $Y=1.84 $X2=14.12 $Y2=1.985
r271 8 55 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=13.025
+ $Y=1.84 $X2=13.17 $Y2=2.815
r272 8 52 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=13.025
+ $Y=1.84 $X2=13.17 $Y2=1.985
r273 7 49 600 $w=1.7e-07 $l=3.745e-07 $layer=licon1_PDIFF $count=1 $X=11.875
+ $Y=2.54 $X2=12.11 $Y2=2.815
r274 7 46 300 $w=1.7e-07 $l=5.39861e-07 $layer=licon1_PDIFF $count=2 $X=11.875
+ $Y=2.54 $X2=12.11 $Y2=2.105
r275 6 135 300 $w=1.7e-07 $l=6.22495e-07 $layer=licon1_PDIFF $count=2 $X=10.575
+ $Y=2.54 $X2=11.075 $Y2=2.815
r276 5 42 600 $w=1.7e-07 $l=2.57488e-07 $layer=licon1_PDIFF $count=1 $X=8.27
+ $Y=2.34 $X2=8.415 $Y2=2.535
r277 4 38 600 $w=1.7e-07 $l=6.46916e-07 $layer=licon1_PDIFF $count=1 $X=7.08
+ $Y=2.285 $X2=7.315 $Y2=2.825
r278 3 34 600 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=4.72
+ $Y=1.84 $X2=4.87 $Y2=2.815
r279 2 30 600 $w=1.7e-07 $l=5.39815e-07 $layer=licon1_PDIFF $count=1 $X=3.11
+ $Y=2.32 $X2=3.26 $Y2=2.79
r280 1 122 150 $w=1.7e-07 $l=8.8955e-07 $layer=licon1_PDIFF $count=4 $X=0.58
+ $Y=2.32 $X2=1.4 $Y2=2.465
.ends

.subckt PM_SKY130_FD_SC_HS__SDFRTP_2%A_390_81# 1 2 3 4 5 18 22 25 26 27 29 30 32
+ 33 36 38 40 41 43 45 50
c151 29 0 1.19423e-19 $X=3.53 $Y=2.33
c152 26 0 5.70693e-20 $X=3.445 $Y=1.225
c153 18 0 7.57672e-20 $X=2.875 $Y=0.72
r154 52 54 0.921954 $w=2.48e-07 $l=2e-08 $layer=LI1_cond $X=5.87 $Y=2.475
+ $X2=5.87 $Y2=2.495
r155 50 52 11.7549 $w=2.48e-07 $l=2.55e-07 $layer=LI1_cond $X=5.87 $Y=2.22
+ $X2=5.87 $Y2=2.475
r156 42 43 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=6.445 $Y=1.465
+ $X2=6.445 $Y2=2.135
r157 40 42 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.36 $Y=1.38
+ $X2=6.445 $Y2=1.465
r158 40 41 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=6.36 $Y=1.38
+ $X2=6.145 $Y2=1.38
r159 39 50 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.995 $Y=2.22
+ $X2=5.87 $Y2=2.22
r160 38 43 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.36 $Y=2.22
+ $X2=6.445 $Y2=2.135
r161 38 39 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=6.36 $Y=2.22
+ $X2=5.995 $Y2=2.22
r162 34 41 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=5.98 $Y=1.295
+ $X2=6.145 $Y2=1.38
r163 34 36 13.7944 $w=3.28e-07 $l=3.95e-07 $layer=LI1_cond $X=5.98 $Y=1.295
+ $X2=5.98 $Y2=0.9
r164 33 49 9.90656 $w=2.16e-07 $l=1.79374e-07 $layer=LI1_cond $X=3.995 $Y=2.475
+ $X2=3.83 $Y2=2.445
r165 32 52 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.745 $Y=2.475
+ $X2=5.87 $Y2=2.475
r166 32 33 114.171 $w=1.68e-07 $l=1.75e-06 $layer=LI1_cond $X=5.745 $Y=2.475
+ $X2=3.995 $Y2=2.475
r167 30 49 1.41204 $w=2.16e-07 $l=2.5e-08 $layer=LI1_cond $X=3.805 $Y=2.445
+ $X2=3.83 $Y2=2.445
r168 30 46 15.5324 $w=2.16e-07 $l=2.75e-07 $layer=LI1_cond $X=3.805 $Y=2.445
+ $X2=3.53 $Y2=2.445
r169 29 46 2.14224 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=3.53 $Y=2.33
+ $X2=3.53 $Y2=2.445
r170 28 29 66.5455 $w=1.68e-07 $l=1.02e-06 $layer=LI1_cond $X=3.53 $Y=1.31
+ $X2=3.53 $Y2=2.33
r171 26 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.445 $Y=1.225
+ $X2=3.53 $Y2=1.31
r172 26 27 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=3.445 $Y=1.225
+ $X2=3.045 $Y2=1.225
r173 25 27 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.96 $Y=1.14
+ $X2=3.045 $Y2=1.225
r174 24 25 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=2.96 $Y=0.845
+ $X2=2.96 $Y2=1.14
r175 23 45 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.435 $Y=2.43
+ $X2=2.27 $Y2=2.43
r176 22 46 5.38804 $w=2.16e-07 $l=9.21954e-08 $layer=LI1_cond $X=3.445 $Y=2.43
+ $X2=3.53 $Y2=2.445
r177 22 23 65.8931 $w=1.68e-07 $l=1.01e-06 $layer=LI1_cond $X=3.445 $Y=2.43
+ $X2=2.435 $Y2=2.43
r178 18 24 7.14316 $w=2.5e-07 $l=1.62019e-07 $layer=LI1_cond $X=2.875 $Y=0.72
+ $X2=2.96 $Y2=0.845
r179 18 20 20.0525 $w=2.48e-07 $l=4.35e-07 $layer=LI1_cond $X=2.875 $Y=0.72
+ $X2=2.44 $Y2=0.72
r180 5 54 600 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_PDIFF $count=1 $X=5.765
+ $Y=2.285 $X2=5.91 $Y2=2.495
r181 4 49 300 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=2 $X=3.68
+ $Y=2.32 $X2=3.83 $Y2=2.465
r182 3 45 300 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=2 $X=2.12
+ $Y=2.32 $X2=2.27 $Y2=2.465
r183 2 36 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=5.835
+ $Y=0.69 $X2=5.98 $Y2=0.9
r184 1 20 182 $w=1.7e-07 $l=6.1225e-07 $layer=licon1_NDIFF $count=1 $X=1.95
+ $Y=0.405 $X2=2.44 $Y2=0.68
.ends

.subckt PM_SKY130_FD_SC_HS__SDFRTP_2%Q 1 2 9 13 14 15 29
r21 20 29 1.74613 $w=3.28e-07 $l=5e-08 $layer=LI1_cond $X=13.69 $Y=1.245
+ $X2=13.69 $Y2=1.295
r22 15 31 3.97298 $w=3.28e-07 $l=9.8e-08 $layer=LI1_cond $X=13.69 $Y=1.312
+ $X2=13.69 $Y2=1.41
r23 15 29 0.593683 $w=3.28e-07 $l=1.7e-08 $layer=LI1_cond $X=13.69 $Y=1.312
+ $X2=13.69 $Y2=1.295
r24 15 20 0.628605 $w=3.28e-07 $l=1.8e-08 $layer=LI1_cond $X=13.69 $Y=1.227
+ $X2=13.69 $Y2=1.245
r25 14 15 10.5466 $w=3.28e-07 $l=3.02e-07 $layer=LI1_cond $X=13.69 $Y=0.925
+ $X2=13.69 $Y2=1.227
r26 13 14 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=13.69 $Y=0.515
+ $X2=13.69 $Y2=0.925
r27 9 11 36.7895 $w=2.58e-07 $l=8.3e-07 $layer=LI1_cond $X=13.655 $Y=1.985
+ $X2=13.655 $Y2=2.815
r28 9 31 25.4867 $w=2.58e-07 $l=5.75e-07 $layer=LI1_cond $X=13.655 $Y=1.985
+ $X2=13.655 $Y2=1.41
r29 2 11 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=13.47
+ $Y=1.84 $X2=13.62 $Y2=2.815
r30 2 9 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=13.47
+ $Y=1.84 $X2=13.62 $Y2=1.985
r31 1 13 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=13.55
+ $Y=0.37 $X2=13.69 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__SDFRTP_2%VGND 1 2 3 4 5 6 7 8 27 31 35 39 43 47 49
+ 51 54 55 56 58 70 74 79 84 89 94 100 103 113 116 119 123
c137 123 0 6.57667e-20 $X=14.16 $Y=0
c138 3 0 1.84505e-19 $X=4.765 $Y=0.37
r139 122 123 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=14.16 $Y=0
+ $X2=14.16 $Y2=0
r140 119 120 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.2 $Y=0
+ $X2=13.2 $Y2=0
r141 116 117 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.24 $Y=0
+ $X2=12.24 $Y2=0
r142 113 114 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=10.8 $Y=0
+ $X2=10.8 $Y2=0
r143 103 104 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=5.04 $Y=0
+ $X2=5.04 $Y2=0
r144 100 101 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0
+ $X2=0.72 $Y2=0
r145 98 123 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=13.68 $Y=0
+ $X2=14.16 $Y2=0
r146 98 120 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=13.68 $Y=0
+ $X2=13.2 $Y2=0
r147 97 98 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.68 $Y=0
+ $X2=13.68 $Y2=0
r148 95 119 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=13.345 $Y=0
+ $X2=13.22 $Y2=0
r149 95 97 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=13.345 $Y=0
+ $X2=13.68 $Y2=0
r150 94 122 4.01252 $w=1.7e-07 $l=1.82e-07 $layer=LI1_cond $X=14.035 $Y=0
+ $X2=14.217 $Y2=0
r151 94 97 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=14.035 $Y=0
+ $X2=13.68 $Y2=0
r152 93 120 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.72 $Y=0
+ $X2=13.2 $Y2=0
r153 93 117 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.72 $Y=0
+ $X2=12.24 $Y2=0
r154 92 93 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.72 $Y=0
+ $X2=12.72 $Y2=0
r155 90 116 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12.435 $Y=0
+ $X2=12.27 $Y2=0
r156 90 92 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=12.435 $Y=0
+ $X2=12.72 $Y2=0
r157 89 119 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=13.095 $Y=0
+ $X2=13.22 $Y2=0
r158 89 92 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=13.095 $Y=0
+ $X2=12.72 $Y2=0
r159 88 117 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.76 $Y=0
+ $X2=12.24 $Y2=0
r160 88 114 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=11.76 $Y=0
+ $X2=10.8 $Y2=0
r161 87 88 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=11.76 $Y=0
+ $X2=11.76 $Y2=0
r162 85 113 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.085 $Y=0
+ $X2=10.92 $Y2=0
r163 85 87 44.0374 $w=1.68e-07 $l=6.75e-07 $layer=LI1_cond $X=11.085 $Y=0
+ $X2=11.76 $Y2=0
r164 84 116 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12.105 $Y=0
+ $X2=12.27 $Y2=0
r165 84 87 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=12.105 $Y=0
+ $X2=11.76 $Y2=0
r166 83 114 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=8.4 $Y=0 $X2=10.8
+ $Y2=0
r167 83 108 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=0 $X2=7.92
+ $Y2=0
r168 82 83 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r169 80 82 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=8.08 $Y=0 $X2=8.4
+ $Y2=0
r170 79 113 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.755 $Y=0
+ $X2=10.92 $Y2=0
r171 79 82 153.642 $w=1.68e-07 $l=2.355e-06 $layer=LI1_cond $X=10.755 $Y=0
+ $X2=8.4 $Y2=0
r172 78 108 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=0
+ $X2=7.92 $Y2=0
r173 77 78 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=7.44 $Y=0 $X2=7.44
+ $Y2=0
r174 75 103 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.07 $Y=0
+ $X2=4.905 $Y2=0
r175 75 77 154.62 $w=1.68e-07 $l=2.37e-06 $layer=LI1_cond $X=5.07 $Y=0 $X2=7.44
+ $Y2=0
r176 74 110 8.18369 $w=4.73e-07 $l=3.25e-07 $layer=LI1_cond $X=7.842 $Y=0
+ $X2=7.842 $Y2=0.325
r177 74 80 6.83586 $w=1.7e-07 $l=2.38e-07 $layer=LI1_cond $X=7.842 $Y=0 $X2=8.08
+ $Y2=0
r178 74 108 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=0 $X2=7.92
+ $Y2=0
r179 74 77 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=7.605 $Y=0
+ $X2=7.44 $Y2=0
r180 73 104 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0
+ $X2=5.04 $Y2=0
r181 72 73 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r182 70 103 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.74 $Y=0
+ $X2=4.905 $Y2=0
r183 70 72 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=4.74 $Y=0 $X2=4.56
+ $Y2=0
r184 69 73 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.56
+ $Y2=0
r185 68 69 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r186 66 69 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=1.2 $Y=0 $X2=3.6
+ $Y2=0
r187 66 101 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r188 65 68 156.578 $w=1.68e-07 $l=2.4e-06 $layer=LI1_cond $X=1.2 $Y=0 $X2=3.6
+ $Y2=0
r189 65 66 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r190 63 100 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.875 $Y=0
+ $X2=0.71 $Y2=0
r191 63 65 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.875 $Y=0 $X2=1.2
+ $Y2=0
r192 61 101 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0
+ $X2=0.72 $Y2=0
r193 60 61 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r194 58 100 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.545 $Y=0
+ $X2=0.71 $Y2=0
r195 58 60 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.545 $Y=0
+ $X2=0.24 $Y2=0
r196 56 78 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=7.2 $Y=0 $X2=7.44
+ $Y2=0
r197 56 104 0.602067 $w=4.9e-07 $l=2.16e-06 $layer=MET1_cond $X=7.2 $Y=0
+ $X2=5.04 $Y2=0
r198 54 68 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=3.715 $Y=0 $X2=3.6
+ $Y2=0
r199 54 55 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.715 $Y=0 $X2=3.88
+ $Y2=0
r200 53 72 33.5989 $w=1.68e-07 $l=5.15e-07 $layer=LI1_cond $X=4.045 $Y=0
+ $X2=4.56 $Y2=0
r201 53 55 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.045 $Y=0 $X2=3.88
+ $Y2=0
r202 49 122 3.13065 $w=2.5e-07 $l=1.09864e-07 $layer=LI1_cond $X=14.16 $Y=0.085
+ $X2=14.217 $Y2=0
r203 49 51 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=14.16 $Y=0.085
+ $X2=14.16 $Y2=0.515
r204 45 119 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=13.22 $Y=0.085
+ $X2=13.22 $Y2=0
r205 45 47 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=13.22 $Y=0.085
+ $X2=13.22 $Y2=0.515
r206 41 116 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=12.27 $Y=0.085
+ $X2=12.27 $Y2=0
r207 41 43 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=12.27 $Y=0.085
+ $X2=12.27 $Y2=0.515
r208 37 113 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=10.92 $Y=0.085
+ $X2=10.92 $Y2=0
r209 37 39 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=10.92 $Y=0.085
+ $X2=10.92 $Y2=0.58
r210 33 103 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.905 $Y=0.085
+ $X2=4.905 $Y2=0
r211 33 35 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=4.905 $Y=0.085
+ $X2=4.905 $Y2=0.55
r212 29 55 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.88 $Y=0.085
+ $X2=3.88 $Y2=0
r213 29 31 18.5089 $w=3.28e-07 $l=5.3e-07 $layer=LI1_cond $X=3.88 $Y=0.085
+ $X2=3.88 $Y2=0.615
r214 25 100 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.71 $Y=0.085
+ $X2=0.71 $Y2=0
r215 25 27 16.4136 $w=3.28e-07 $l=4.7e-07 $layer=LI1_cond $X=0.71 $Y=0.085
+ $X2=0.71 $Y2=0.555
r216 8 51 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=13.98
+ $Y=0.37 $X2=14.12 $Y2=0.515
r217 7 47 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=13.115
+ $Y=0.37 $X2=13.26 $Y2=0.515
r218 6 43 182 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=1 $X=12.125
+ $Y=0.37 $X2=12.27 $Y2=0.515
r219 5 39 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=10.78
+ $Y=0.37 $X2=10.92 $Y2=0.58
r220 4 110 182 $w=1.7e-07 $l=4.88953e-07 $layer=licon1_NDIFF $count=1 $X=7.55
+ $Y=0.69 $X2=7.84 $Y2=0.325
r221 3 35 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=4.765
+ $Y=0.37 $X2=4.905 $Y2=0.55
r222 2 31 182 $w=1.7e-07 $l=2.96985e-07 $layer=licon1_NDIFF $count=1 $X=3.67
+ $Y=0.405 $X2=3.88 $Y2=0.615
r223 1 27 182 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.37 $X2=0.71 $Y2=0.555
.ends

.subckt PM_SKY130_FD_SC_HS__SDFRTP_2%noxref_24 1 2 7 11 13
r30 13 16 7.33373 $w=3.28e-07 $l=2.1e-07 $layer=LI1_cond $X=1.27 $Y=0.34
+ $X2=1.27 $Y2=0.55
r31 9 11 6.63528 $w=3.28e-07 $l=1.9e-07 $layer=LI1_cond $X=3.38 $Y=0.425
+ $X2=3.38 $Y2=0.615
r32 8 13 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.435 $Y=0.34
+ $X2=1.27 $Y2=0.34
r33 7 9 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.215 $Y=0.34
+ $X2=3.38 $Y2=0.425
r34 7 8 116.128 $w=1.68e-07 $l=1.78e-06 $layer=LI1_cond $X=3.215 $Y=0.34
+ $X2=1.435 $Y2=0.34
r35 2 11 182 $w=1.7e-07 $l=3.44347e-07 $layer=licon1_NDIFF $count=1 $X=3.125
+ $Y=0.405 $X2=3.38 $Y2=0.615
r36 1 16 182 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=1 $X=1.125
+ $Y=0.405 $X2=1.27 $Y2=0.55
.ends

