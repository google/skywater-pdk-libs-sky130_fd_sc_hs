* File: sky130_fd_sc_hs__o41a_2.pxi.spice
* Created: Tue Sep  1 20:19:16 2020
* 
x_PM_SKY130_FD_SC_HS__O41A_2%A1 N_A1_M1011_g N_A1_c_73_n N_A1_M1007_g A1
+ N_A1_c_74_n PM_SKY130_FD_SC_HS__O41A_2%A1
x_PM_SKY130_FD_SC_HS__O41A_2%A2 N_A2_c_97_n N_A2_M1001_g N_A2_M1013_g
+ N_A2_c_99_n A2 A2 A2 PM_SKY130_FD_SC_HS__O41A_2%A2
x_PM_SKY130_FD_SC_HS__O41A_2%A3 N_A3_M1006_g N_A3_c_133_n N_A3_M1012_g A3 A3 A3
+ A3 PM_SKY130_FD_SC_HS__O41A_2%A3
x_PM_SKY130_FD_SC_HS__O41A_2%A4 N_A4_c_167_n N_A4_M1010_g N_A4_M1004_g A4
+ N_A4_c_169_n PM_SKY130_FD_SC_HS__O41A_2%A4
x_PM_SKY130_FD_SC_HS__O41A_2%B1 N_B1_c_195_n N_B1_M1000_g N_B1_M1009_g B1 B1
+ PM_SKY130_FD_SC_HS__O41A_2%B1
x_PM_SKY130_FD_SC_HS__O41A_2%A_428_368# N_A_428_368#_M1009_d
+ N_A_428_368#_M1010_d N_A_428_368#_M1005_g N_A_428_368#_c_238_n
+ N_A_428_368#_M1002_g N_A_428_368#_M1008_g N_A_428_368#_c_239_n
+ N_A_428_368#_M1003_g N_A_428_368#_c_243_n N_A_428_368#_c_240_n
+ N_A_428_368#_c_250_n N_A_428_368#_c_232_n N_A_428_368#_c_233_n
+ N_A_428_368#_c_234_n N_A_428_368#_c_235_n N_A_428_368#_c_236_n
+ N_A_428_368#_c_237_n PM_SKY130_FD_SC_HS__O41A_2%A_428_368#
x_PM_SKY130_FD_SC_HS__O41A_2%VPWR N_VPWR_M1007_s N_VPWR_M1000_d N_VPWR_M1003_s
+ N_VPWR_c_309_n N_VPWR_c_310_n N_VPWR_c_311_n N_VPWR_c_312_n VPWR
+ N_VPWR_c_313_n N_VPWR_c_314_n N_VPWR_c_315_n N_VPWR_c_308_n
+ PM_SKY130_FD_SC_HS__O41A_2%VPWR
x_PM_SKY130_FD_SC_HS__O41A_2%X N_X_M1005_d N_X_M1002_d N_X_c_360_n N_X_c_361_n
+ N_X_c_362_n X PM_SKY130_FD_SC_HS__O41A_2%X
x_PM_SKY130_FD_SC_HS__O41A_2%A_27_74# N_A_27_74#_M1011_s N_A_27_74#_M1013_d
+ N_A_27_74#_M1004_d N_A_27_74#_c_383_n N_A_27_74#_c_384_n N_A_27_74#_c_385_n
+ N_A_27_74#_c_386_n N_A_27_74#_c_387_n N_A_27_74#_c_388_n N_A_27_74#_c_389_n
+ PM_SKY130_FD_SC_HS__O41A_2%A_27_74#
x_PM_SKY130_FD_SC_HS__O41A_2%VGND N_VGND_M1011_d N_VGND_M1006_d N_VGND_M1005_s
+ N_VGND_M1008_s N_VGND_c_436_n N_VGND_c_437_n N_VGND_c_438_n N_VGND_c_439_n
+ N_VGND_c_440_n N_VGND_c_441_n VGND N_VGND_c_442_n N_VGND_c_443_n
+ N_VGND_c_444_n N_VGND_c_445_n N_VGND_c_446_n N_VGND_c_447_n N_VGND_c_448_n
+ PM_SKY130_FD_SC_HS__O41A_2%VGND
cc_1 VNB N_A1_M1011_g 0.0348798f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_2 VNB N_A1_c_73_n 0.0276543f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.765
cc_3 VNB N_A1_c_74_n 0.0155193f $X=-0.19 $Y=-0.245 $X2=0.43 $Y2=1.515
cc_4 VNB N_A2_c_97_n 0.0269678f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.35
cc_5 VNB N_A2_M1013_g 0.0257807f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_6 VNB N_A2_c_99_n 0.00167106f $X=-0.19 $Y=-0.245 $X2=0.43 $Y2=1.515
cc_7 VNB N_A3_M1006_g 0.0273614f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_8 VNB N_A3_c_133_n 0.022392f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.765
cc_9 VNB A3 0.00465445f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_10 VNB N_A4_c_167_n 0.0269778f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.35
cc_11 VNB N_A4_M1004_g 0.0275785f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_12 VNB N_A4_c_169_n 0.00166777f $X=-0.19 $Y=-0.245 $X2=0.43 $Y2=1.515
cc_13 VNB N_B1_c_195_n 0.0267626f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.35
cc_14 VNB N_B1_M1009_g 0.0281622f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_15 VNB B1 0.00953293f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_428_368#_M1005_g 0.0224767f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_428_368#_M1008_g 0.0265448f $X=-0.19 $Y=-0.245 $X2=0.43 $Y2=1.565
cc_18 VNB N_A_428_368#_c_232_n 0.0104431f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_428_368#_c_233_n 0.01612f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_428_368#_c_234_n 0.00406491f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_428_368#_c_235_n 4.08426e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_428_368#_c_236_n 0.00840116f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_428_368#_c_237_n 0.0985742f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_VPWR_c_308_n 0.203486f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_X_c_360_n 0.00240191f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_X_c_361_n 0.00415351f $X=-0.19 $Y=-0.245 $X2=0.43 $Y2=1.515
cc_27 VNB N_X_c_362_n 4.65031e-19 $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.565
cc_28 VNB N_A_27_74#_c_383_n 0.0277086f $X=-0.19 $Y=-0.245 $X2=0.43 $Y2=1.515
cc_29 VNB N_A_27_74#_c_384_n 0.00948616f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_27_74#_c_385_n 0.00995328f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_27_74#_c_386_n 0.00240191f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_27_74#_c_387_n 0.0188114f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_27_74#_c_388_n 0.00253059f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_27_74#_c_389_n 0.0100545f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_436_n 0.00900728f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_437_n 0.0186948f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_438_n 0.0109596f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_439_n 0.0139769f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_440_n 0.0131032f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_441_n 0.0117082f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_442_n 0.0191515f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_443_n 0.0339528f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_444_n 0.0186948f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_445_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_VGND_c_446_n 0.00980973f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_VGND_c_447_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_VGND_c_448_n 0.285003f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VPB N_A1_c_73_n 0.0305897f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.765
cc_49 VPB N_A1_c_74_n 0.00889413f $X=-0.19 $Y=1.66 $X2=0.43 $Y2=1.515
cc_50 VPB N_A2_c_97_n 0.0271752f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.35
cc_51 VPB N_A2_c_99_n 0.00213487f $X=-0.19 $Y=1.66 $X2=0.43 $Y2=1.515
cc_52 VPB N_A3_c_133_n 0.0292972f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.765
cc_53 VPB A3 0.00181505f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_54 VPB N_A4_c_167_n 0.0299902f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.35
cc_55 VPB N_A4_c_169_n 0.00284535f $X=-0.19 $Y=1.66 $X2=0.43 $Y2=1.515
cc_56 VPB N_B1_c_195_n 0.0303605f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.35
cc_57 VPB B1 0.00773518f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_58 VPB N_A_428_368#_c_238_n 0.0171963f $X=-0.19 $Y=1.66 $X2=0.43 $Y2=1.515
cc_59 VPB N_A_428_368#_c_239_n 0.0186863f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_60 VPB N_A_428_368#_c_240_n 0.00384301f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_61 VPB N_A_428_368#_c_235_n 0.00340738f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_62 VPB N_A_428_368#_c_237_n 0.017335f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_63 VPB N_VPWR_c_309_n 0.0120106f $X=-0.19 $Y=1.66 $X2=0.43 $Y2=1.515
cc_64 VPB N_VPWR_c_310_n 0.0489067f $X=-0.19 $Y=1.66 $X2=0.43 $Y2=1.515
cc_65 VPB N_VPWR_c_311_n 0.0120106f $X=-0.19 $Y=1.66 $X2=0.43 $Y2=1.565
cc_66 VPB N_VPWR_c_312_n 0.0651399f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_67 VPB N_VPWR_c_313_n 0.0641878f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_68 VPB N_VPWR_c_314_n 0.0163631f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_69 VPB N_VPWR_c_315_n 0.0366166f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_70 VPB N_VPWR_c_308_n 0.0866974f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_71 VPB N_X_c_362_n 0.00506469f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=1.565
cc_72 N_A1_c_73_n N_A2_c_97_n 0.0801924f $X=0.505 $Y=1.765 $X2=-0.19 $Y2=-0.245
cc_73 N_A1_c_74_n N_A2_c_97_n 0.00154471f $X=0.43 $Y=1.515 $X2=-0.19 $Y2=-0.245
cc_74 N_A1_M1011_g N_A2_M1013_g 0.0260254f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_75 N_A1_c_73_n N_A2_c_99_n 0.00473801f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_76 N_A1_c_74_n N_A2_c_99_n 0.0252745f $X=0.43 $Y=1.515 $X2=0 $Y2=0
cc_77 N_A1_c_73_n N_VPWR_c_310_n 0.0207642f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_78 N_A1_c_74_n N_VPWR_c_310_n 0.0255179f $X=0.43 $Y=1.515 $X2=0 $Y2=0
cc_79 N_A1_c_73_n N_VPWR_c_313_n 0.00413917f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_80 N_A1_c_73_n N_VPWR_c_308_n 0.00817532f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_81 N_A1_M1011_g N_A_27_74#_c_383_n 0.0103339f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_82 N_A1_M1011_g N_A_27_74#_c_384_n 0.0117984f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_83 N_A1_c_73_n N_A_27_74#_c_384_n 6.16197e-19 $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_84 N_A1_c_74_n N_A_27_74#_c_384_n 0.0110042f $X=0.43 $Y=1.515 $X2=0 $Y2=0
cc_85 N_A1_M1011_g N_A_27_74#_c_385_n 0.00214722f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_86 N_A1_c_73_n N_A_27_74#_c_385_n 0.00361626f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_87 N_A1_c_74_n N_A_27_74#_c_385_n 0.0279713f $X=0.43 $Y=1.515 $X2=0 $Y2=0
cc_88 N_A1_M1011_g N_A_27_74#_c_386_n 6.28869e-19 $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_89 N_A1_M1011_g N_VGND_c_436_n 0.00622602f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_90 N_A1_M1011_g N_VGND_c_442_n 0.00434272f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_91 N_A1_M1011_g N_VGND_c_448_n 0.0082497f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_92 N_A2_M1013_g N_A3_M1006_g 0.019972f $X=1.065 $Y=0.74 $X2=0 $Y2=0
cc_93 N_A2_c_97_n N_A3_c_133_n 0.0522582f $X=0.925 $Y=1.765 $X2=0 $Y2=0
cc_94 N_A2_c_99_n N_A3_c_133_n 0.00251729f $X=1 $Y=1.515 $X2=0 $Y2=0
cc_95 A2 N_A3_c_133_n 0.00959387f $X=1.115 $Y=1.95 $X2=0 $Y2=0
cc_96 N_A2_c_97_n A3 0.00211252f $X=0.925 $Y=1.765 $X2=0 $Y2=0
cc_97 N_A2_c_99_n A3 0.0286223f $X=1 $Y=1.515 $X2=0 $Y2=0
cc_98 A2 A3 0.0562235f $X=1.115 $Y=1.95 $X2=0 $Y2=0
cc_99 N_A2_c_97_n N_VPWR_c_310_n 0.00195604f $X=0.925 $Y=1.765 $X2=0 $Y2=0
cc_100 N_A2_c_97_n N_VPWR_c_313_n 0.00303293f $X=0.925 $Y=1.765 $X2=0 $Y2=0
cc_101 A2 N_VPWR_c_313_n 0.0138369f $X=1.115 $Y=2.32 $X2=0 $Y2=0
cc_102 N_A2_c_97_n N_VPWR_c_308_n 0.00372936f $X=0.925 $Y=1.765 $X2=0 $Y2=0
cc_103 A2 N_VPWR_c_308_n 0.0159188f $X=1.115 $Y=2.32 $X2=0 $Y2=0
cc_104 N_A2_c_99_n A_200_368# 9.9932e-19 $X=1 $Y=1.515 $X2=-0.19 $Y2=-0.245
cc_105 A2 A_200_368# 0.0108532f $X=1.115 $Y=1.95 $X2=-0.19 $Y2=-0.245
cc_106 A2 A_200_368# 0.0161826f $X=1.115 $Y=2.32 $X2=-0.19 $Y2=-0.245
cc_107 N_A2_M1013_g N_A_27_74#_c_383_n 6.28869e-19 $X=1.065 $Y=0.74 $X2=0 $Y2=0
cc_108 N_A2_c_97_n N_A_27_74#_c_384_n 0.00107205f $X=0.925 $Y=1.765 $X2=0 $Y2=0
cc_109 N_A2_M1013_g N_A_27_74#_c_384_n 0.0117933f $X=1.065 $Y=0.74 $X2=0 $Y2=0
cc_110 N_A2_c_99_n N_A_27_74#_c_384_n 0.0217949f $X=1 $Y=1.515 $X2=0 $Y2=0
cc_111 N_A2_M1013_g N_A_27_74#_c_386_n 0.00966073f $X=1.065 $Y=0.74 $X2=0 $Y2=0
cc_112 N_A2_M1013_g N_A_27_74#_c_389_n 0.0015571f $X=1.065 $Y=0.74 $X2=0 $Y2=0
cc_113 N_A2_c_99_n N_A_27_74#_c_389_n 0.00425598f $X=1 $Y=1.515 $X2=0 $Y2=0
cc_114 N_A2_M1013_g N_VGND_c_436_n 0.00484409f $X=1.065 $Y=0.74 $X2=0 $Y2=0
cc_115 N_A2_M1013_g N_VGND_c_437_n 0.00434272f $X=1.065 $Y=0.74 $X2=0 $Y2=0
cc_116 N_A2_M1013_g N_VGND_c_448_n 0.0082141f $X=1.065 $Y=0.74 $X2=0 $Y2=0
cc_117 N_A3_c_133_n N_A4_c_167_n 0.0519601f $X=1.495 $Y=1.765 $X2=-0.19
+ $Y2=-0.245
cc_118 A3 N_A4_c_167_n 0.0146009f $X=1.595 $Y=1.58 $X2=-0.19 $Y2=-0.245
cc_119 N_A3_M1006_g N_A4_M1004_g 0.018224f $X=1.495 $Y=0.74 $X2=0 $Y2=0
cc_120 N_A3_c_133_n N_A4_c_169_n 4.85968e-19 $X=1.495 $Y=1.765 $X2=0 $Y2=0
cc_121 A3 N_A4_c_169_n 0.0327491f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_122 A3 N_A_428_368#_c_243_n 0.00817432f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_123 N_A3_c_133_n N_A_428_368#_c_240_n 0.00102748f $X=1.495 $Y=1.765 $X2=0
+ $Y2=0
cc_124 A3 N_A_428_368#_c_240_n 0.0349229f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_125 N_A3_c_133_n N_VPWR_c_313_n 0.00457246f $X=1.495 $Y=1.765 $X2=0 $Y2=0
cc_126 A3 N_VPWR_c_313_n 0.0063665f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_127 N_A3_c_133_n N_VPWR_c_308_n 0.00893363f $X=1.495 $Y=1.765 $X2=0 $Y2=0
cc_128 A3 N_VPWR_c_308_n 0.00792965f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_129 A3 A_314_368# 0.0166298f $X=1.595 $Y=1.58 $X2=-0.19 $Y2=-0.245
cc_130 N_A3_M1006_g N_A_27_74#_c_386_n 0.0145272f $X=1.495 $Y=0.74 $X2=0 $Y2=0
cc_131 N_A3_M1006_g N_A_27_74#_c_387_n 0.0122944f $X=1.495 $Y=0.74 $X2=0 $Y2=0
cc_132 N_A3_c_133_n N_A_27_74#_c_387_n 0.00371567f $X=1.495 $Y=1.765 $X2=0 $Y2=0
cc_133 A3 N_A_27_74#_c_387_n 0.0260507f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_134 N_A3_M1006_g N_A_27_74#_c_389_n 0.00155819f $X=1.495 $Y=0.74 $X2=0 $Y2=0
cc_135 N_A3_c_133_n N_A_27_74#_c_389_n 3.65737e-19 $X=1.495 $Y=1.765 $X2=0 $Y2=0
cc_136 A3 N_A_27_74#_c_389_n 0.00326062f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_137 N_A3_M1006_g N_VGND_c_437_n 0.00434272f $X=1.495 $Y=0.74 $X2=0 $Y2=0
cc_138 N_A3_M1006_g N_VGND_c_438_n 0.00586574f $X=1.495 $Y=0.74 $X2=0 $Y2=0
cc_139 N_A3_M1006_g N_VGND_c_448_n 0.00822442f $X=1.495 $Y=0.74 $X2=0 $Y2=0
cc_140 N_A4_c_167_n N_B1_c_195_n 0.0363251f $X=2.065 $Y=1.765 $X2=-0.19
+ $Y2=-0.245
cc_141 N_A4_c_169_n N_B1_c_195_n 7.80108e-19 $X=2.14 $Y=1.515 $X2=-0.19
+ $Y2=-0.245
cc_142 N_A4_M1004_g N_B1_M1009_g 0.0193383f $X=2.23 $Y=0.74 $X2=0 $Y2=0
cc_143 N_A4_c_167_n B1 0.00251621f $X=2.065 $Y=1.765 $X2=0 $Y2=0
cc_144 N_A4_c_169_n B1 0.0302881f $X=2.14 $Y=1.515 $X2=0 $Y2=0
cc_145 N_A4_c_167_n N_A_428_368#_c_243_n 0.00328702f $X=2.065 $Y=1.765 $X2=0
+ $Y2=0
cc_146 N_A4_c_169_n N_A_428_368#_c_243_n 0.0131798f $X=2.14 $Y=1.515 $X2=0 $Y2=0
cc_147 N_A4_c_167_n N_A_428_368#_c_240_n 0.012525f $X=2.065 $Y=1.765 $X2=0 $Y2=0
cc_148 N_A4_c_167_n N_VPWR_c_313_n 0.00445602f $X=2.065 $Y=1.765 $X2=0 $Y2=0
cc_149 N_A4_c_167_n N_VPWR_c_315_n 0.00318675f $X=2.065 $Y=1.765 $X2=0 $Y2=0
cc_150 N_A4_c_167_n N_VPWR_c_308_n 0.00864208f $X=2.065 $Y=1.765 $X2=0 $Y2=0
cc_151 N_A4_c_167_n N_A_27_74#_c_387_n 0.00124693f $X=2.065 $Y=1.765 $X2=0 $Y2=0
cc_152 N_A4_M1004_g N_A_27_74#_c_387_n 0.0145711f $X=2.23 $Y=0.74 $X2=0 $Y2=0
cc_153 N_A4_c_169_n N_A_27_74#_c_387_n 0.0247664f $X=2.14 $Y=1.515 $X2=0 $Y2=0
cc_154 N_A4_M1004_g N_A_27_74#_c_388_n 0.013702f $X=2.23 $Y=0.74 $X2=0 $Y2=0
cc_155 N_A4_M1004_g N_VGND_c_438_n 0.00757529f $X=2.23 $Y=0.74 $X2=0 $Y2=0
cc_156 N_A4_M1004_g N_VGND_c_443_n 0.00451267f $X=2.23 $Y=0.74 $X2=0 $Y2=0
cc_157 N_A4_M1004_g N_VGND_c_448_n 0.00877274f $X=2.23 $Y=0.74 $X2=0 $Y2=0
cc_158 N_B1_c_195_n N_A_428_368#_c_240_n 0.0109555f $X=2.635 $Y=1.765 $X2=0
+ $Y2=0
cc_159 N_B1_c_195_n N_A_428_368#_c_250_n 0.0180748f $X=2.635 $Y=1.765 $X2=0
+ $Y2=0
cc_160 B1 N_A_428_368#_c_250_n 0.052208f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_161 N_B1_M1009_g N_A_428_368#_c_232_n 0.00161219f $X=2.675 $Y=0.74 $X2=0
+ $Y2=0
cc_162 B1 N_A_428_368#_c_233_n 0.00887071f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_163 N_B1_c_195_n N_A_428_368#_c_234_n 0.00186365f $X=2.635 $Y=1.765 $X2=0
+ $Y2=0
cc_164 N_B1_M1009_g N_A_428_368#_c_234_n 0.00162779f $X=2.675 $Y=0.74 $X2=0
+ $Y2=0
cc_165 B1 N_A_428_368#_c_234_n 0.0294134f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_166 N_B1_c_195_n N_A_428_368#_c_235_n 0.00425882f $X=2.635 $Y=1.765 $X2=0
+ $Y2=0
cc_167 B1 N_A_428_368#_c_235_n 0.0271533f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_168 N_B1_M1009_g N_A_428_368#_c_236_n 0.00273312f $X=2.675 $Y=0.74 $X2=0
+ $Y2=0
cc_169 B1 N_A_428_368#_c_236_n 0.00969568f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_170 N_B1_c_195_n N_A_428_368#_c_237_n 0.00488449f $X=2.635 $Y=1.765 $X2=0
+ $Y2=0
cc_171 N_B1_M1009_g N_A_428_368#_c_237_n 6.21883e-19 $X=2.675 $Y=0.74 $X2=0
+ $Y2=0
cc_172 B1 N_A_428_368#_c_237_n 0.00239357f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_173 N_B1_c_195_n N_VPWR_c_313_n 0.00444645f $X=2.635 $Y=1.765 $X2=0 $Y2=0
cc_174 N_B1_c_195_n N_VPWR_c_315_n 0.0113047f $X=2.635 $Y=1.765 $X2=0 $Y2=0
cc_175 N_B1_c_195_n N_VPWR_c_308_n 0.00460931f $X=2.635 $Y=1.765 $X2=0 $Y2=0
cc_176 N_B1_c_195_n N_A_27_74#_c_387_n 0.00145533f $X=2.635 $Y=1.765 $X2=0 $Y2=0
cc_177 N_B1_M1009_g N_A_27_74#_c_387_n 0.00302367f $X=2.675 $Y=0.74 $X2=0 $Y2=0
cc_178 B1 N_A_27_74#_c_387_n 0.00856196f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_179 N_B1_M1009_g N_A_27_74#_c_388_n 0.0082268f $X=2.675 $Y=0.74 $X2=0 $Y2=0
cc_180 N_B1_M1009_g N_VGND_c_439_n 0.00327253f $X=2.675 $Y=0.74 $X2=0 $Y2=0
cc_181 N_B1_M1009_g N_VGND_c_443_n 0.00434272f $X=2.675 $Y=0.74 $X2=0 $Y2=0
cc_182 N_B1_M1009_g N_VGND_c_448_n 0.00826504f $X=2.675 $Y=0.74 $X2=0 $Y2=0
cc_183 N_A_428_368#_c_250_n N_VPWR_M1000_d 0.0290021f $X=3.405 $Y=2.035 $X2=0
+ $Y2=0
cc_184 N_A_428_368#_c_235_n N_VPWR_M1000_d 0.00398391f $X=3.57 $Y=1.95 $X2=0
+ $Y2=0
cc_185 N_A_428_368#_c_238_n N_VPWR_c_312_n 6.79505e-19 $X=3.845 $Y=1.765 $X2=0
+ $Y2=0
cc_186 N_A_428_368#_c_239_n N_VPWR_c_312_n 0.0186805f $X=4.295 $Y=1.765 $X2=0
+ $Y2=0
cc_187 N_A_428_368#_c_237_n N_VPWR_c_312_n 7.4439e-19 $X=4.235 $Y=1.532 $X2=0
+ $Y2=0
cc_188 N_A_428_368#_c_240_n N_VPWR_c_313_n 0.0145938f $X=2.29 $Y=2.815 $X2=0
+ $Y2=0
cc_189 N_A_428_368#_c_238_n N_VPWR_c_314_n 0.004307f $X=3.845 $Y=1.765 $X2=0
+ $Y2=0
cc_190 N_A_428_368#_c_239_n N_VPWR_c_314_n 0.00413917f $X=4.295 $Y=1.765 $X2=0
+ $Y2=0
cc_191 N_A_428_368#_c_238_n N_VPWR_c_315_n 0.013111f $X=3.845 $Y=1.765 $X2=0
+ $Y2=0
cc_192 N_A_428_368#_c_239_n N_VPWR_c_315_n 4.9724e-19 $X=4.295 $Y=1.765 $X2=0
+ $Y2=0
cc_193 N_A_428_368#_c_240_n N_VPWR_c_315_n 0.043685f $X=2.29 $Y=2.815 $X2=0
+ $Y2=0
cc_194 N_A_428_368#_c_250_n N_VPWR_c_315_n 0.0806194f $X=3.405 $Y=2.035 $X2=0
+ $Y2=0
cc_195 N_A_428_368#_c_237_n N_VPWR_c_315_n 9.63724e-19 $X=4.235 $Y=1.532 $X2=0
+ $Y2=0
cc_196 N_A_428_368#_c_238_n N_VPWR_c_308_n 0.00847721f $X=3.845 $Y=1.765 $X2=0
+ $Y2=0
cc_197 N_A_428_368#_c_239_n N_VPWR_c_308_n 0.00817726f $X=4.295 $Y=1.765 $X2=0
+ $Y2=0
cc_198 N_A_428_368#_c_240_n N_VPWR_c_308_n 0.0120466f $X=2.29 $Y=2.815 $X2=0
+ $Y2=0
cc_199 N_A_428_368#_M1005_g N_X_c_360_n 0.0124354f $X=3.805 $Y=0.74 $X2=0 $Y2=0
cc_200 N_A_428_368#_M1008_g N_X_c_360_n 0.00772833f $X=4.235 $Y=0.74 $X2=0 $Y2=0
cc_201 N_A_428_368#_M1005_g N_X_c_361_n 0.006795f $X=3.805 $Y=0.74 $X2=0 $Y2=0
cc_202 N_A_428_368#_M1008_g N_X_c_361_n 0.0150748f $X=4.235 $Y=0.74 $X2=0 $Y2=0
cc_203 N_A_428_368#_c_236_n N_X_c_361_n 0.0214332f $X=3.57 $Y=1.465 $X2=0 $Y2=0
cc_204 N_A_428_368#_c_237_n N_X_c_361_n 0.0128724f $X=4.235 $Y=1.532 $X2=0 $Y2=0
cc_205 N_A_428_368#_c_238_n N_X_c_362_n 0.00101636f $X=3.845 $Y=1.765 $X2=0
+ $Y2=0
cc_206 N_A_428_368#_c_239_n N_X_c_362_n 0.00556772f $X=4.295 $Y=1.765 $X2=0
+ $Y2=0
cc_207 N_A_428_368#_c_235_n N_X_c_362_n 0.0241031f $X=3.57 $Y=1.95 $X2=0 $Y2=0
cc_208 N_A_428_368#_c_236_n N_X_c_362_n 0.0032852f $X=3.57 $Y=1.465 $X2=0 $Y2=0
cc_209 N_A_428_368#_c_237_n N_X_c_362_n 0.0259109f $X=4.235 $Y=1.532 $X2=0 $Y2=0
cc_210 N_A_428_368#_c_234_n N_A_27_74#_c_387_n 0.0104256f $X=3.125 $Y=1.095
+ $X2=0 $Y2=0
cc_211 N_A_428_368#_c_232_n N_A_27_74#_c_388_n 0.0255177f $X=2.89 $Y=0.515 $X2=0
+ $Y2=0
cc_212 N_A_428_368#_c_233_n N_VGND_M1005_s 4.82091e-19 $X=3.405 $Y=1.095 $X2=0
+ $Y2=0
cc_213 N_A_428_368#_c_236_n N_VGND_M1005_s 0.00397467f $X=3.57 $Y=1.465 $X2=0
+ $Y2=0
cc_214 N_A_428_368#_M1005_g N_VGND_c_439_n 0.00545191f $X=3.805 $Y=0.74 $X2=0
+ $Y2=0
cc_215 N_A_428_368#_c_232_n N_VGND_c_439_n 0.0316872f $X=2.89 $Y=0.515 $X2=0
+ $Y2=0
cc_216 N_A_428_368#_c_233_n N_VGND_c_439_n 0.00369599f $X=3.405 $Y=1.095 $X2=0
+ $Y2=0
cc_217 N_A_428_368#_c_236_n N_VGND_c_439_n 0.0181094f $X=3.57 $Y=1.465 $X2=0
+ $Y2=0
cc_218 N_A_428_368#_c_237_n N_VGND_c_439_n 0.00141269f $X=4.235 $Y=1.532 $X2=0
+ $Y2=0
cc_219 N_A_428_368#_M1008_g N_VGND_c_441_n 0.00364571f $X=4.235 $Y=0.74 $X2=0
+ $Y2=0
cc_220 N_A_428_368#_c_237_n N_VGND_c_441_n 7.78919e-19 $X=4.235 $Y=1.532 $X2=0
+ $Y2=0
cc_221 N_A_428_368#_c_232_n N_VGND_c_443_n 0.0146357f $X=2.89 $Y=0.515 $X2=0
+ $Y2=0
cc_222 N_A_428_368#_M1005_g N_VGND_c_444_n 0.00434272f $X=3.805 $Y=0.74 $X2=0
+ $Y2=0
cc_223 N_A_428_368#_M1008_g N_VGND_c_444_n 0.00434272f $X=4.235 $Y=0.74 $X2=0
+ $Y2=0
cc_224 N_A_428_368#_M1005_g N_VGND_c_448_n 0.00825059f $X=3.805 $Y=0.74 $X2=0
+ $Y2=0
cc_225 N_A_428_368#_M1008_g N_VGND_c_448_n 0.00823934f $X=4.235 $Y=0.74 $X2=0
+ $Y2=0
cc_226 N_A_428_368#_c_232_n N_VGND_c_448_n 0.0121141f $X=2.89 $Y=0.515 $X2=0
+ $Y2=0
cc_227 N_VPWR_c_312_n N_X_c_362_n 0.0766785f $X=4.52 $Y=1.985 $X2=0 $Y2=0
cc_228 N_VPWR_c_314_n N_X_c_362_n 0.00905805f $X=4.355 $Y=3.33 $X2=0 $Y2=0
cc_229 N_VPWR_c_315_n N_X_c_362_n 0.0296638f $X=3.215 $Y=2.375 $X2=0 $Y2=0
cc_230 N_VPWR_c_308_n N_X_c_362_n 0.00749747f $X=4.56 $Y=3.33 $X2=0 $Y2=0
cc_231 N_X_c_360_n N_VGND_c_439_n 0.018426f $X=4.02 $Y=0.515 $X2=0 $Y2=0
cc_232 N_X_c_360_n N_VGND_c_441_n 0.0238012f $X=4.02 $Y=0.515 $X2=0 $Y2=0
cc_233 N_X_c_360_n N_VGND_c_444_n 0.0144922f $X=4.02 $Y=0.515 $X2=0 $Y2=0
cc_234 N_X_c_360_n N_VGND_c_448_n 0.0118826f $X=4.02 $Y=0.515 $X2=0 $Y2=0
cc_235 N_A_27_74#_c_384_n N_VGND_M1011_d 0.00358162f $X=1.115 $Y=1.095 $X2=-0.19
+ $Y2=-0.245
cc_236 N_A_27_74#_c_387_n N_VGND_M1006_d 0.00654166f $X=2.295 $Y=1.095 $X2=0
+ $Y2=0
cc_237 N_A_27_74#_c_383_n N_VGND_c_436_n 0.0191765f $X=0.28 $Y=0.515 $X2=0 $Y2=0
cc_238 N_A_27_74#_c_384_n N_VGND_c_436_n 0.0248957f $X=1.115 $Y=1.095 $X2=0
+ $Y2=0
cc_239 N_A_27_74#_c_386_n N_VGND_c_436_n 0.0191765f $X=1.28 $Y=0.515 $X2=0 $Y2=0
cc_240 N_A_27_74#_c_386_n N_VGND_c_437_n 0.0144922f $X=1.28 $Y=0.515 $X2=0 $Y2=0
cc_241 N_A_27_74#_c_386_n N_VGND_c_438_n 0.0182921f $X=1.28 $Y=0.515 $X2=0 $Y2=0
cc_242 N_A_27_74#_c_387_n N_VGND_c_438_n 0.0345921f $X=2.295 $Y=1.095 $X2=0
+ $Y2=0
cc_243 N_A_27_74#_c_388_n N_VGND_c_438_n 0.0182921f $X=2.46 $Y=0.515 $X2=0 $Y2=0
cc_244 N_A_27_74#_c_383_n N_VGND_c_442_n 0.0145639f $X=0.28 $Y=0.515 $X2=0 $Y2=0
cc_245 N_A_27_74#_c_388_n N_VGND_c_443_n 0.014537f $X=2.46 $Y=0.515 $X2=0 $Y2=0
cc_246 N_A_27_74#_c_383_n N_VGND_c_448_n 0.0119984f $X=0.28 $Y=0.515 $X2=0 $Y2=0
cc_247 N_A_27_74#_c_386_n N_VGND_c_448_n 0.0118826f $X=1.28 $Y=0.515 $X2=0 $Y2=0
cc_248 N_A_27_74#_c_388_n N_VGND_c_448_n 0.011955f $X=2.46 $Y=0.515 $X2=0 $Y2=0
