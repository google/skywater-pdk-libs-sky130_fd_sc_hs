* File: sky130_fd_sc_hs__dfxbp_2.pxi.spice
* Created: Thu Aug 27 20:39:49 2020
* 
x_PM_SKY130_FD_SC_HS__DFXBP_2%CLK N_CLK_c_221_n N_CLK_M1025_g N_CLK_c_222_n
+ N_CLK_M1017_g CLK N_CLK_c_223_n PM_SKY130_FD_SC_HS__DFXBP_2%CLK
x_PM_SKY130_FD_SC_HS__DFXBP_2%A_27_74# N_A_27_74#_M1025_s N_A_27_74#_M1017_s
+ N_A_27_74#_c_248_n N_A_27_74#_M1016_g N_A_27_74#_c_249_n N_A_27_74#_M1011_g
+ N_A_27_74#_c_250_n N_A_27_74#_M1026_g N_A_27_74#_c_251_n N_A_27_74#_c_280_n
+ N_A_27_74#_M1029_g N_A_27_74#_c_281_n N_A_27_74#_M1000_g N_A_27_74#_c_252_n
+ N_A_27_74#_c_253_n N_A_27_74#_c_254_n N_A_27_74#_M1002_g N_A_27_74#_c_256_n
+ N_A_27_74#_c_257_n N_A_27_74#_c_258_n N_A_27_74#_c_259_n N_A_27_74#_c_285_n
+ N_A_27_74#_c_296_n N_A_27_74#_c_260_n N_A_27_74#_c_286_n N_A_27_74#_c_287_n
+ N_A_27_74#_c_261_n N_A_27_74#_c_262_n N_A_27_74#_c_263_n N_A_27_74#_c_264_n
+ N_A_27_74#_c_265_n N_A_27_74#_c_266_n N_A_27_74#_c_267_n N_A_27_74#_c_268_n
+ N_A_27_74#_c_269_n N_A_27_74#_c_334_p N_A_27_74#_c_270_n N_A_27_74#_c_271_n
+ N_A_27_74#_c_272_n N_A_27_74#_c_273_n N_A_27_74#_c_375_p N_A_27_74#_c_274_n
+ N_A_27_74#_c_290_n N_A_27_74#_c_331_p N_A_27_74#_c_275_n N_A_27_74#_c_276_n
+ N_A_27_74#_c_277_n PM_SKY130_FD_SC_HS__DFXBP_2%A_27_74#
x_PM_SKY130_FD_SC_HS__DFXBP_2%D N_D_c_517_n N_D_M1022_g N_D_c_513_n N_D_M1024_g
+ N_D_c_518_n N_D_c_519_n N_D_c_520_n D D N_D_c_515_n D
+ PM_SKY130_FD_SC_HS__DFXBP_2%D
x_PM_SKY130_FD_SC_HS__DFXBP_2%A_206_368# N_A_206_368#_M1011_d
+ N_A_206_368#_M1016_d N_A_206_368#_c_570_n N_A_206_368#_c_571_n
+ N_A_206_368#_c_581_n N_A_206_368#_c_582_n N_A_206_368#_c_583_n
+ N_A_206_368#_M1028_g N_A_206_368#_M1014_g N_A_206_368#_M1012_g
+ N_A_206_368#_c_584_n N_A_206_368#_M1030_g N_A_206_368#_c_585_n
+ N_A_206_368#_c_574_n N_A_206_368#_c_586_n N_A_206_368#_c_575_n
+ N_A_206_368#_c_588_n N_A_206_368#_c_589_n N_A_206_368#_c_576_n
+ N_A_206_368#_c_577_n N_A_206_368#_c_578_n N_A_206_368#_c_579_n
+ N_A_206_368#_c_592_n N_A_206_368#_c_580_n
+ PM_SKY130_FD_SC_HS__DFXBP_2%A_206_368#
x_PM_SKY130_FD_SC_HS__DFXBP_2%A_753_284# N_A_753_284#_M1007_d
+ N_A_753_284#_M1031_d N_A_753_284#_c_759_n N_A_753_284#_c_760_n
+ N_A_753_284#_c_766_n N_A_753_284#_M1005_g N_A_753_284#_M1004_g
+ N_A_753_284#_c_762_n N_A_753_284#_c_763_n N_A_753_284#_c_764_n
+ PM_SKY130_FD_SC_HS__DFXBP_2%A_753_284#
x_PM_SKY130_FD_SC_HS__DFXBP_2%A_558_445# N_A_558_445#_M1026_d
+ N_A_558_445#_M1028_d N_A_558_445#_M1007_g N_A_558_445#_c_817_n
+ N_A_558_445#_M1031_g N_A_558_445#_c_818_n N_A_558_445#_c_819_n
+ N_A_558_445#_c_820_n N_A_558_445#_c_846_n N_A_558_445#_c_859_n
+ N_A_558_445#_c_824_n N_A_558_445#_c_821_n
+ PM_SKY130_FD_SC_HS__DFXBP_2%A_558_445#
x_PM_SKY130_FD_SC_HS__DFXBP_2%A_1290_102# N_A_1290_102#_M1021_s
+ N_A_1290_102#_M1015_d N_A_1290_102#_c_894_n N_A_1290_102#_M1010_g
+ N_A_1290_102#_c_913_n N_A_1290_102#_c_914_n N_A_1290_102#_c_915_n
+ N_A_1290_102#_M1032_g N_A_1290_102#_M1003_g N_A_1290_102#_c_896_n
+ N_A_1290_102#_c_917_n N_A_1290_102#_M1001_g N_A_1290_102#_c_897_n
+ N_A_1290_102#_M1013_g N_A_1290_102#_c_899_n N_A_1290_102#_M1009_g
+ N_A_1290_102#_c_919_n N_A_1290_102#_M1019_g N_A_1290_102#_M1027_g
+ N_A_1290_102#_c_901_n N_A_1290_102#_c_902_n N_A_1290_102#_c_903_n
+ N_A_1290_102#_c_904_n N_A_1290_102#_c_905_n N_A_1290_102#_c_906_n
+ N_A_1290_102#_c_907_n N_A_1290_102#_c_908_n N_A_1290_102#_c_909_n
+ N_A_1290_102#_c_910_n N_A_1290_102#_c_923_n N_A_1290_102#_c_911_n
+ N_A_1290_102#_c_925_n N_A_1290_102#_c_938_p N_A_1290_102#_c_912_n
+ PM_SKY130_FD_SC_HS__DFXBP_2%A_1290_102#
x_PM_SKY130_FD_SC_HS__DFXBP_2%A_1000_424# N_A_1000_424#_M1012_d
+ N_A_1000_424#_M1000_d N_A_1000_424#_c_1067_n N_A_1000_424#_M1015_g
+ N_A_1000_424#_c_1068_n N_A_1000_424#_M1020_g N_A_1000_424#_M1021_g
+ N_A_1000_424#_c_1069_n N_A_1000_424#_c_1059_n N_A_1000_424#_c_1060_n
+ N_A_1000_424#_c_1061_n N_A_1000_424#_c_1072_n N_A_1000_424#_c_1062_n
+ N_A_1000_424#_c_1063_n N_A_1000_424#_c_1064_n N_A_1000_424#_c_1065_n
+ N_A_1000_424#_c_1066_n PM_SKY130_FD_SC_HS__DFXBP_2%A_1000_424#
x_PM_SKY130_FD_SC_HS__DFXBP_2%A_1835_368# N_A_1835_368#_M1027_s
+ N_A_1835_368#_M1019_s N_A_1835_368#_c_1174_n N_A_1835_368#_M1018_g
+ N_A_1835_368#_M1006_g N_A_1835_368#_c_1175_n N_A_1835_368#_M1023_g
+ N_A_1835_368#_M1008_g N_A_1835_368#_c_1170_n N_A_1835_368#_c_1176_n
+ N_A_1835_368#_c_1171_n N_A_1835_368#_c_1172_n N_A_1835_368#_c_1173_n
+ PM_SKY130_FD_SC_HS__DFXBP_2%A_1835_368#
x_PM_SKY130_FD_SC_HS__DFXBP_2%VPWR N_VPWR_M1017_d N_VPWR_M1022_s N_VPWR_M1005_d
+ N_VPWR_M1032_d N_VPWR_M1020_s N_VPWR_M1009_s N_VPWR_M1019_d N_VPWR_M1023_s
+ N_VPWR_c_1238_n N_VPWR_c_1239_n N_VPWR_c_1240_n N_VPWR_c_1241_n
+ N_VPWR_c_1242_n N_VPWR_c_1243_n N_VPWR_c_1244_n N_VPWR_c_1245_n
+ N_VPWR_c_1246_n N_VPWR_c_1247_n N_VPWR_c_1248_n VPWR N_VPWR_c_1249_n
+ N_VPWR_c_1250_n N_VPWR_c_1251_n N_VPWR_c_1252_n N_VPWR_c_1253_n
+ N_VPWR_c_1254_n N_VPWR_c_1255_n N_VPWR_c_1256_n N_VPWR_c_1257_n
+ N_VPWR_c_1258_n N_VPWR_c_1237_n PM_SKY130_FD_SC_HS__DFXBP_2%VPWR
x_PM_SKY130_FD_SC_HS__DFXBP_2%A_451_503# N_A_451_503#_M1024_d
+ N_A_451_503#_M1022_d N_A_451_503#_c_1355_n N_A_451_503#_c_1356_n
+ N_A_451_503#_c_1359_n N_A_451_503#_c_1357_n
+ PM_SKY130_FD_SC_HS__DFXBP_2%A_451_503#
x_PM_SKY130_FD_SC_HS__DFXBP_2%Q N_Q_M1003_d N_Q_M1001_d N_Q_c_1396_n Q
+ PM_SKY130_FD_SC_HS__DFXBP_2%Q
x_PM_SKY130_FD_SC_HS__DFXBP_2%Q_N N_Q_N_M1006_d N_Q_N_M1018_d N_Q_N_c_1417_n
+ N_Q_N_c_1418_n Q_N Q_N Q_N Q_N N_Q_N_c_1419_n PM_SKY130_FD_SC_HS__DFXBP_2%Q_N
x_PM_SKY130_FD_SC_HS__DFXBP_2%VGND N_VGND_M1025_d N_VGND_M1024_s N_VGND_M1004_d
+ N_VGND_M1010_d N_VGND_M1021_d N_VGND_M1013_s N_VGND_M1027_d N_VGND_M1008_s
+ N_VGND_c_1447_n N_VGND_c_1448_n N_VGND_c_1449_n N_VGND_c_1450_n
+ N_VGND_c_1451_n N_VGND_c_1452_n N_VGND_c_1453_n N_VGND_c_1454_n
+ N_VGND_c_1455_n N_VGND_c_1456_n N_VGND_c_1457_n N_VGND_c_1458_n
+ N_VGND_c_1459_n N_VGND_c_1460_n N_VGND_c_1461_n N_VGND_c_1462_n VGND
+ N_VGND_c_1463_n N_VGND_c_1464_n N_VGND_c_1465_n N_VGND_c_1466_n
+ N_VGND_c_1467_n N_VGND_c_1468_n N_VGND_c_1469_n N_VGND_c_1470_n
+ N_VGND_c_1471_n PM_SKY130_FD_SC_HS__DFXBP_2%VGND
cc_1 VNB N_CLK_c_221_n 0.0248291f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.22
cc_2 VNB N_CLK_c_222_n 0.0454833f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.765
cc_3 VNB N_CLK_c_223_n 0.0186611f $X=-0.19 $Y=-0.245 $X2=0.42 $Y2=1.385
cc_4 VNB N_A_27_74#_c_248_n 0.0455305f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_5 VNB N_A_27_74#_c_249_n 0.0201109f $X=-0.19 $Y=-0.245 $X2=0.42 $Y2=1.385
cc_6 VNB N_A_27_74#_c_250_n 0.014006f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_7 VNB N_A_27_74#_c_251_n 0.028028f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_A_27_74#_c_252_n 0.0110465f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A_27_74#_c_253_n 0.0107485f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_27_74#_c_254_n 0.0250517f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_27_74#_M1002_g 0.00825398f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_27_74#_c_256_n 0.0170488f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_27_74#_c_257_n 0.0187971f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_27_74#_c_258_n 0.0772123f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_27_74#_c_259_n 0.0170752f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_27_74#_c_260_n 0.0120699f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_27_74#_c_261_n 0.00193848f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_27_74#_c_262_n 0.00103927f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_27_74#_c_263_n 0.00517734f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_27_74#_c_264_n 0.00279668f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_27_74#_c_265_n 0.0233946f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_27_74#_c_266_n 0.00145623f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_27_74#_c_267_n 6.70789e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_27_74#_c_268_n 0.0113863f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_27_74#_c_269_n 0.0080865f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_27_74#_c_270_n 0.00804801f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_27_74#_c_271_n 0.00266108f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_27_74#_c_272_n 0.00984407f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_27_74#_c_273_n 0.00361919f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_27_74#_c_274_n 0.00323288f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_27_74#_c_275_n 9.09959e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_27_74#_c_276_n 0.00328754f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_27_74#_c_277_n 0.0334971f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_D_c_513_n 0.0167887f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.765
cc_35 VNB D 0.00853968f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_D_c_515_n 0.0483977f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB D 0.00104288f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_206_368#_c_570_n 0.125066f $X=-0.19 $Y=-0.245 $X2=0.425 $Y2=1.385
cc_39 VNB N_A_206_368#_c_571_n 0.0124378f $X=-0.19 $Y=-0.245 $X2=0.42 $Y2=1.385
cc_40 VNB N_A_206_368#_M1014_g 0.0271426f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_206_368#_M1012_g 0.02346f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_206_368#_c_574_n 0.00615862f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_206_368#_c_575_n 0.00564079f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_206_368#_c_576_n 0.00410678f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_A_206_368#_c_577_n 0.0191451f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_A_206_368#_c_578_n 0.00426517f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_206_368#_c_579_n 0.0377215f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_206_368#_c_580_n 0.0783778f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A_753_284#_c_759_n 0.0424085f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_50 VNB N_A_753_284#_c_760_n 0.0254986f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_A_753_284#_M1004_g 0.0202168f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_A_753_284#_c_762_n 0.0153406f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_A_753_284#_c_763_n 2.0776e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_A_753_284#_c_764_n 0.0101325f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_A_558_445#_M1007_g 0.0503954f $X=-0.19 $Y=-0.245 $X2=0.425 $Y2=1.385
cc_56 VNB N_A_558_445#_c_817_n 0.0320978f $X=-0.19 $Y=-0.245 $X2=0.42 $Y2=1.385
cc_57 VNB N_A_558_445#_c_818_n 0.00109969f $X=-0.19 $Y=-0.245 $X2=0.42 $Y2=1.365
cc_58 VNB N_A_558_445#_c_819_n 0.00668477f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_A_558_445#_c_820_n 0.0033222f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_A_558_445#_c_821_n 0.00185469f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_A_1290_102#_c_894_n 0.0184985f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_62 VNB N_A_1290_102#_M1003_g 0.021048f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_A_1290_102#_c_896_n 0.00974444f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_A_1290_102#_c_897_n 0.0138996f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_A_1290_102#_M1013_g 0.0221515f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_A_1290_102#_c_899_n 0.0102557f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_A_1290_102#_M1027_g 0.026822f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_A_1290_102#_c_901_n 0.0130894f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_A_1290_102#_c_902_n 0.0134612f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_A_1290_102#_c_903_n 0.00607022f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_A_1290_102#_c_904_n 0.0836964f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_A_1290_102#_c_905_n 0.0105969f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_A_1290_102#_c_906_n 0.00740382f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_A_1290_102#_c_907_n 0.0461614f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_A_1290_102#_c_908_n 0.0115974f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_A_1290_102#_c_909_n 0.00737837f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_A_1290_102#_c_910_n 0.00289355f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_A_1290_102#_c_911_n 0.00524712f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VNB N_A_1290_102#_c_912_n 0.00462034f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_A_1000_424#_M1021_g 0.042928f $X=-0.19 $Y=-0.245 $X2=0.42 $Y2=1.365
cc_81 VNB N_A_1000_424#_c_1059_n 0.00264572f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_82 VNB N_A_1000_424#_c_1060_n 0.00411523f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_83 VNB N_A_1000_424#_c_1061_n 0.00766825f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_84 VNB N_A_1000_424#_c_1062_n 2.98211e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_85 VNB N_A_1000_424#_c_1063_n 2.4818e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_86 VNB N_A_1000_424#_c_1064_n 0.00530038f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_87 VNB N_A_1000_424#_c_1065_n 0.00280538f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_88 VNB N_A_1000_424#_c_1066_n 0.00926369f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_89 VNB N_A_1835_368#_M1006_g 0.0228003f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.365
cc_90 VNB N_A_1835_368#_M1008_g 0.0260188f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_91 VNB N_A_1835_368#_c_1170_n 0.00552991f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_92 VNB N_A_1835_368#_c_1171_n 0.00834609f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_93 VNB N_A_1835_368#_c_1172_n 3.4825e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_94 VNB N_A_1835_368#_c_1173_n 0.0739491f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_95 VNB N_VPWR_c_1237_n 0.462217f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_96 VNB N_A_451_503#_c_1355_n 0.00636495f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_97 VNB N_A_451_503#_c_1356_n 0.00230704f $X=-0.19 $Y=-0.245 $X2=0.42
+ $Y2=1.385
cc_98 VNB N_A_451_503#_c_1357_n 0.00615407f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_99 VNB N_Q_c_1396_n 0.00444959f $X=-0.19 $Y=-0.245 $X2=0.425 $Y2=1.385
cc_100 VNB N_Q_N_c_1417_n 0.00240191f $X=-0.19 $Y=-0.245 $X2=0.425 $Y2=1.385
cc_101 VNB N_Q_N_c_1418_n 0.00429087f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_102 VNB N_Q_N_c_1419_n 0.00142046f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_103 VNB N_VGND_c_1447_n 0.00900288f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_104 VNB N_VGND_c_1448_n 0.00444947f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_105 VNB N_VGND_c_1449_n 0.0446419f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_106 VNB N_VGND_c_1450_n 0.00821481f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_107 VNB N_VGND_c_1451_n 0.020982f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_108 VNB N_VGND_c_1452_n 0.0104237f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_109 VNB N_VGND_c_1453_n 0.0240648f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_110 VNB N_VGND_c_1454_n 0.0147061f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_111 VNB N_VGND_c_1455_n 0.010678f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_112 VNB N_VGND_c_1456_n 0.0505285f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_113 VNB N_VGND_c_1457_n 0.0571046f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_114 VNB N_VGND_c_1458_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_115 VNB N_VGND_c_1459_n 0.0190497f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_116 VNB N_VGND_c_1460_n 0.00630956f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_117 VNB N_VGND_c_1461_n 0.0181728f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_118 VNB N_VGND_c_1462_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_119 VNB N_VGND_c_1463_n 0.0187989f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_120 VNB N_VGND_c_1464_n 0.0228203f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_121 VNB N_VGND_c_1465_n 0.0231643f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_122 VNB N_VGND_c_1466_n 0.0192531f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_123 VNB N_VGND_c_1467_n 0.00737741f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_124 VNB N_VGND_c_1468_n 0.0043669f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_125 VNB N_VGND_c_1469_n 0.00640372f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_126 VNB N_VGND_c_1470_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_127 VNB N_VGND_c_1471_n 0.600453f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_128 VPB N_CLK_c_222_n 0.0283447f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.765
cc_129 VPB N_A_27_74#_c_248_n 0.0236139f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.21
cc_130 VPB N_A_27_74#_c_251_n 0.00416232f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_131 VPB N_A_27_74#_c_280_n 0.015388f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_132 VPB N_A_27_74#_c_281_n 0.019741f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_133 VPB N_A_27_74#_c_252_n 0.0368428f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_134 VPB N_A_27_74#_c_253_n 0.00212274f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_135 VPB N_A_27_74#_c_257_n 0.00706385f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_136 VPB N_A_27_74#_c_285_n 0.0441294f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_137 VPB N_A_27_74#_c_286_n 0.00546222f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_138 VPB N_A_27_74#_c_287_n 0.0100637f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_139 VPB N_A_27_74#_c_262_n 5.62538e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_140 VPB N_A_27_74#_c_268_n 0.00556198f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_141 VPB N_A_27_74#_c_290_n 0.0525507f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_142 VPB N_D_c_517_n 0.0208791f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.22
cc_143 VPB N_D_c_518_n 0.00463479f $X=-0.19 $Y=1.66 $X2=0.42 $Y2=1.385
cc_144 VPB N_D_c_519_n 0.0523228f $X=-0.19 $Y=1.66 $X2=0.42 $Y2=1.385
cc_145 VPB N_D_c_520_n 0.00514898f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=1.365
cc_146 VPB N_A_206_368#_c_581_n 0.0591271f $X=-0.19 $Y=1.66 $X2=0.42 $Y2=1.385
cc_147 VPB N_A_206_368#_c_582_n 0.0154119f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_148 VPB N_A_206_368#_c_583_n 0.022034f $X=-0.19 $Y=1.66 $X2=0.42 $Y2=1.365
cc_149 VPB N_A_206_368#_c_584_n 0.0620045f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_150 VPB N_A_206_368#_c_585_n 0.0212579f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_151 VPB N_A_206_368#_c_586_n 0.0258394f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_152 VPB N_A_206_368#_c_575_n 0.00309425f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_153 VPB N_A_206_368#_c_588_n 0.0125057f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_154 VPB N_A_206_368#_c_589_n 0.00241053f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_155 VPB N_A_206_368#_c_576_n 0.0226329f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_156 VPB N_A_206_368#_c_577_n 0.0179103f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_157 VPB N_A_206_368#_c_592_n 0.00147829f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_158 VPB N_A_753_284#_c_760_n 0.00694019f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_159 VPB N_A_753_284#_c_766_n 0.0211462f $X=-0.19 $Y=1.66 $X2=0.425 $Y2=1.385
cc_160 VPB N_A_753_284#_c_764_n 0.00275013f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_161 VPB N_A_558_445#_c_817_n 0.0312556f $X=-0.19 $Y=1.66 $X2=0.42 $Y2=1.385
cc_162 VPB N_A_558_445#_c_818_n 0.00500181f $X=-0.19 $Y=1.66 $X2=0.42 $Y2=1.365
cc_163 VPB N_A_558_445#_c_824_n 0.00262443f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_164 VPB N_A_558_445#_c_821_n 0.00101928f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_165 VPB N_A_1290_102#_c_913_n 0.00656714f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=1.365
cc_166 VPB N_A_1290_102#_c_914_n 0.0235663f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_167 VPB N_A_1290_102#_c_915_n 0.0233244f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_168 VPB N_A_1290_102#_c_896_n 6.7296e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_169 VPB N_A_1290_102#_c_917_n 0.0210074f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_170 VPB N_A_1290_102#_c_899_n 0.0234374f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_171 VPB N_A_1290_102#_c_919_n 0.017871f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_172 VPB N_A_1290_102#_c_902_n 0.00542996f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_173 VPB N_A_1290_102#_c_905_n 0.00858094f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_174 VPB N_A_1290_102#_c_910_n 0.00321692f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_175 VPB N_A_1290_102#_c_923_n 0.00585896f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_176 VPB N_A_1290_102#_c_911_n 0.00723663f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_177 VPB N_A_1290_102#_c_925_n 0.00256516f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_178 VPB N_A_1000_424#_c_1067_n 0.0165346f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.21
cc_179 VPB N_A_1000_424#_c_1068_n 0.0164849f $X=-0.19 $Y=1.66 $X2=0.42 $Y2=1.385
cc_180 VPB N_A_1000_424#_c_1069_n 0.0130476f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_181 VPB N_A_1000_424#_c_1059_n 0.00736567f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_182 VPB N_A_1000_424#_c_1060_n 2.81715e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_183 VPB N_A_1000_424#_c_1072_n 0.0122882f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_184 VPB N_A_1000_424#_c_1063_n 0.00177415f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_185 VPB N_A_1000_424#_c_1064_n 0.00628421f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_186 VPB N_A_1000_424#_c_1065_n 0.0050355f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_187 VPB N_A_1000_424#_c_1066_n 0.0550712f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_188 VPB N_A_1835_368#_c_1174_n 0.0163067f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.21
cc_189 VPB N_A_1835_368#_c_1175_n 0.017361f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_190 VPB N_A_1835_368#_c_1176_n 0.00417913f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_191 VPB N_A_1835_368#_c_1173_n 0.0168942f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_192 VPB N_VPWR_c_1238_n 0.00571271f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_193 VPB N_VPWR_c_1239_n 0.014158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_194 VPB N_VPWR_c_1240_n 0.00592663f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_195 VPB N_VPWR_c_1241_n 0.0136488f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_196 VPB N_VPWR_c_1242_n 0.0157532f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_197 VPB N_VPWR_c_1243_n 0.0106521f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_198 VPB N_VPWR_c_1244_n 0.0645004f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_199 VPB N_VPWR_c_1245_n 0.0594915f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_200 VPB N_VPWR_c_1246_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_201 VPB N_VPWR_c_1247_n 0.0177589f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_202 VPB N_VPWR_c_1248_n 0.00614127f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_203 VPB N_VPWR_c_1249_n 0.0518591f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_204 VPB N_VPWR_c_1250_n 0.0217179f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_205 VPB N_VPWR_c_1251_n 0.0227498f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_206 VPB N_VPWR_c_1252_n 0.0204898f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_207 VPB N_VPWR_c_1253_n 0.0247087f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_208 VPB N_VPWR_c_1254_n 0.0182228f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_209 VPB N_VPWR_c_1255_n 0.0179606f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_210 VPB N_VPWR_c_1256_n 0.0173402f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_211 VPB N_VPWR_c_1257_n 0.00614127f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_212 VPB N_VPWR_c_1258_n 0.0047828f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_213 VPB N_VPWR_c_1237_n 0.154642f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_214 VPB N_A_451_503#_c_1355_n 0.00457508f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_215 VPB N_A_451_503#_c_1359_n 0.00497685f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_216 VPB Q_N 0.00201765f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_217 VPB Q_N 0.00257348f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_218 VPB N_Q_N_c_1419_n 0.00105273f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_219 N_CLK_c_222_n N_A_27_74#_c_248_n 0.0526417f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_220 N_CLK_c_223_n N_A_27_74#_c_248_n 3.658e-19 $X=0.42 $Y=1.385 $X2=0 $Y2=0
cc_221 N_CLK_c_221_n N_A_27_74#_c_249_n 0.0182726f $X=0.495 $Y=1.22 $X2=0 $Y2=0
cc_222 N_CLK_c_221_n N_A_27_74#_c_259_n 0.00687376f $X=0.495 $Y=1.22 $X2=0 $Y2=0
cc_223 N_CLK_c_222_n N_A_27_74#_c_285_n 0.0140455f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_224 N_CLK_c_221_n N_A_27_74#_c_296_n 0.0128696f $X=0.495 $Y=1.22 $X2=0 $Y2=0
cc_225 N_CLK_c_223_n N_A_27_74#_c_296_n 0.00994571f $X=0.42 $Y=1.385 $X2=0 $Y2=0
cc_226 N_CLK_c_221_n N_A_27_74#_c_260_n 9.65763e-19 $X=0.495 $Y=1.22 $X2=0 $Y2=0
cc_227 N_CLK_c_222_n N_A_27_74#_c_260_n 0.00100741f $X=0.505 $Y=1.765 $X2=0
+ $Y2=0
cc_228 N_CLK_c_223_n N_A_27_74#_c_260_n 0.0251668f $X=0.42 $Y=1.385 $X2=0 $Y2=0
cc_229 N_CLK_c_222_n N_A_27_74#_c_286_n 0.012687f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_230 N_CLK_c_223_n N_A_27_74#_c_286_n 0.0100567f $X=0.42 $Y=1.385 $X2=0 $Y2=0
cc_231 N_CLK_c_222_n N_A_27_74#_c_287_n 0.00722743f $X=0.505 $Y=1.765 $X2=0
+ $Y2=0
cc_232 N_CLK_c_223_n N_A_27_74#_c_287_n 0.0276095f $X=0.42 $Y=1.385 $X2=0 $Y2=0
cc_233 N_CLK_c_221_n N_A_27_74#_c_261_n 0.0044736f $X=0.495 $Y=1.22 $X2=0 $Y2=0
cc_234 N_CLK_c_222_n N_A_27_74#_c_261_n 0.00545248f $X=0.505 $Y=1.765 $X2=0
+ $Y2=0
cc_235 N_CLK_c_223_n N_A_27_74#_c_261_n 0.0302146f $X=0.42 $Y=1.385 $X2=0 $Y2=0
cc_236 N_CLK_c_222_n N_VPWR_c_1238_n 0.0069311f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_237 N_CLK_c_222_n N_VPWR_c_1253_n 0.00445602f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_238 N_CLK_c_222_n N_VPWR_c_1237_n 0.00861168f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_239 N_CLK_c_221_n N_VGND_c_1447_n 0.00482202f $X=0.495 $Y=1.22 $X2=0 $Y2=0
cc_240 N_CLK_c_221_n N_VGND_c_1463_n 0.00329783f $X=0.495 $Y=1.22 $X2=0 $Y2=0
cc_241 N_CLK_c_221_n N_VGND_c_1471_n 0.00427564f $X=0.495 $Y=1.22 $X2=0 $Y2=0
cc_242 N_A_27_74#_c_250_n N_D_c_513_n 0.00797244f $X=3 $Y=1.09 $X2=0 $Y2=0
cc_243 N_A_27_74#_c_263_n N_D_c_513_n 0.00696197f $X=2.36 $Y=0.815 $X2=0 $Y2=0
cc_244 N_A_27_74#_c_264_n N_D_c_513_n 0.00767546f $X=2.445 $Y=0.73 $X2=0 $Y2=0
cc_245 N_A_27_74#_c_265_n N_D_c_513_n 0.00171466f $X=3.47 $Y=0.34 $X2=0 $Y2=0
cc_246 N_A_27_74#_c_263_n D 0.0248035f $X=2.36 $Y=0.815 $X2=0 $Y2=0
cc_247 N_A_27_74#_c_251_n N_D_c_515_n 0.00275881f $X=3.12 $Y=1.735 $X2=0 $Y2=0
cc_248 N_A_27_74#_c_256_n N_D_c_515_n 0.00797244f $X=3.12 $Y=1.165 $X2=0 $Y2=0
cc_249 N_A_27_74#_c_263_n N_D_c_515_n 0.0055481f $X=2.36 $Y=0.815 $X2=0 $Y2=0
cc_250 N_A_27_74#_c_263_n N_A_206_368#_M1011_d 0.00986221f $X=2.36 $Y=0.815
+ $X2=-0.19 $Y2=-0.245
cc_251 N_A_27_74#_c_250_n N_A_206_368#_c_570_n 0.00882199f $X=3 $Y=1.09 $X2=0
+ $Y2=0
cc_252 N_A_27_74#_c_263_n N_A_206_368#_c_570_n 0.00387758f $X=2.36 $Y=0.815
+ $X2=0 $Y2=0
cc_253 N_A_27_74#_c_265_n N_A_206_368#_c_570_n 0.015696f $X=3.47 $Y=0.34 $X2=0
+ $Y2=0
cc_254 N_A_27_74#_c_266_n N_A_206_368#_c_570_n 0.0035998f $X=2.53 $Y=0.34 $X2=0
+ $Y2=0
cc_255 N_A_27_74#_c_249_n N_A_206_368#_c_571_n 0.015168f $X=1.14 $Y=1.22 $X2=0
+ $Y2=0
cc_256 N_A_27_74#_c_251_n N_A_206_368#_c_581_n 0.0103492f $X=3.12 $Y=1.735 $X2=0
+ $Y2=0
cc_257 N_A_27_74#_c_290_n N_A_206_368#_c_582_n 0.0103492f $X=3.39 $Y=1.9 $X2=0
+ $Y2=0
cc_258 N_A_27_74#_c_280_n N_A_206_368#_c_583_n 0.0107162f $X=3.435 $Y=2.15 $X2=0
+ $Y2=0
cc_259 N_A_27_74#_c_290_n N_A_206_368#_c_583_n 0.00118235f $X=3.39 $Y=1.9 $X2=0
+ $Y2=0
cc_260 N_A_27_74#_c_250_n N_A_206_368#_M1014_g 0.0114381f $X=3 $Y=1.09 $X2=0
+ $Y2=0
cc_261 N_A_27_74#_c_265_n N_A_206_368#_M1014_g 0.0102075f $X=3.47 $Y=0.34 $X2=0
+ $Y2=0
cc_262 N_A_27_74#_c_267_n N_A_206_368#_M1014_g 0.0094249f $X=3.555 $Y=0.78 $X2=0
+ $Y2=0
cc_263 N_A_27_74#_c_268_n N_A_206_368#_M1014_g 0.00494932f $X=3.555 $Y=1.75
+ $X2=0 $Y2=0
cc_264 N_A_27_74#_c_290_n N_A_206_368#_M1014_g 0.00171256f $X=3.39 $Y=1.9 $X2=0
+ $Y2=0
cc_265 N_A_27_74#_c_331_p N_A_206_368#_M1014_g 0.00450183f $X=3.555 $Y=0.865
+ $X2=0 $Y2=0
cc_266 N_A_27_74#_c_258_n N_A_206_368#_M1012_g 0.00590495f $X=6.09 $Y=0.365
+ $X2=0 $Y2=0
cc_267 N_A_27_74#_c_269_n N_A_206_368#_M1012_g 0.00266787f $X=4.645 $Y=0.865
+ $X2=0 $Y2=0
cc_268 N_A_27_74#_c_334_p N_A_206_368#_M1012_g 0.00317769f $X=4.73 $Y=0.78 $X2=0
+ $Y2=0
cc_269 N_A_27_74#_c_270_n N_A_206_368#_M1012_g 0.0179567f $X=5.445 $Y=0.392
+ $X2=0 $Y2=0
cc_270 N_A_27_74#_c_272_n N_A_206_368#_M1012_g 0.0126463f $X=5.53 $Y=1.17 $X2=0
+ $Y2=0
cc_271 N_A_27_74#_c_254_n N_A_206_368#_c_584_n 0.00448785f $X=6.09 $Y=1.245
+ $X2=0 $Y2=0
cc_272 N_A_27_74#_c_248_n N_A_206_368#_c_585_n 0.00552026f $X=0.955 $Y=1.765
+ $X2=0 $Y2=0
cc_273 N_A_27_74#_c_285_n N_A_206_368#_c_585_n 0.00194382f $X=0.28 $Y=1.985
+ $X2=0 $Y2=0
cc_274 N_A_27_74#_c_249_n N_A_206_368#_c_574_n 0.00419009f $X=1.14 $Y=1.22 $X2=0
+ $Y2=0
cc_275 N_A_27_74#_c_261_n N_A_206_368#_c_574_n 0.0311215f $X=0.927 $Y=1.378
+ $X2=0 $Y2=0
cc_276 N_A_27_74#_c_263_n N_A_206_368#_c_574_n 0.0266632f $X=2.36 $Y=0.815 $X2=0
+ $Y2=0
cc_277 N_A_27_74#_c_280_n N_A_206_368#_c_586_n 0.0107841f $X=3.435 $Y=2.15 $X2=0
+ $Y2=0
cc_278 N_A_27_74#_c_281_n N_A_206_368#_c_586_n 0.0157771f $X=4.925 $Y=2.045
+ $X2=0 $Y2=0
cc_279 N_A_27_74#_c_290_n N_A_206_368#_c_586_n 3.12175e-19 $X=3.39 $Y=1.9 $X2=0
+ $Y2=0
cc_280 N_A_27_74#_c_281_n N_A_206_368#_c_575_n 0.0116285f $X=4.925 $Y=2.045
+ $X2=0 $Y2=0
cc_281 N_A_27_74#_c_252_n N_A_206_368#_c_575_n 0.0118097f $X=5.515 $Y=1.765
+ $X2=0 $Y2=0
cc_282 N_A_27_74#_c_253_n N_A_206_368#_c_575_n 3.49966e-19 $X=5.59 $Y=1.69 $X2=0
+ $Y2=0
cc_283 N_A_27_74#_c_257_n N_A_206_368#_c_575_n 0.00502964f $X=4.925 $Y=1.765
+ $X2=0 $Y2=0
cc_284 N_A_27_74#_c_277_n N_A_206_368#_c_575_n 0.00512619f $X=5.68 $Y=1.245
+ $X2=0 $Y2=0
cc_285 N_A_27_74#_c_248_n N_A_206_368#_c_576_n 0.00982303f $X=0.955 $Y=1.765
+ $X2=0 $Y2=0
cc_286 N_A_27_74#_c_285_n N_A_206_368#_c_576_n 0.00259477f $X=0.28 $Y=1.985
+ $X2=0 $Y2=0
cc_287 N_A_27_74#_c_286_n N_A_206_368#_c_576_n 0.0111365f $X=0.755 $Y=1.805
+ $X2=0 $Y2=0
cc_288 N_A_27_74#_c_262_n N_A_206_368#_c_576_n 0.00791807f $X=0.84 $Y=1.72 $X2=0
+ $Y2=0
cc_289 N_A_27_74#_c_263_n N_A_206_368#_c_576_n 0.00579075f $X=2.36 $Y=0.815
+ $X2=0 $Y2=0
cc_290 N_A_27_74#_c_274_n N_A_206_368#_c_576_n 0.00539842f $X=0.97 $Y=1.385
+ $X2=0 $Y2=0
cc_291 N_A_27_74#_c_248_n N_A_206_368#_c_577_n 0.00865081f $X=0.955 $Y=1.765
+ $X2=0 $Y2=0
cc_292 N_A_27_74#_c_263_n N_A_206_368#_c_577_n 6.88622e-19 $X=2.36 $Y=0.815
+ $X2=0 $Y2=0
cc_293 N_A_27_74#_c_252_n N_A_206_368#_c_578_n 4.4812e-19 $X=5.515 $Y=1.765
+ $X2=0 $Y2=0
cc_294 N_A_27_74#_c_257_n N_A_206_368#_c_578_n 3.39287e-19 $X=4.925 $Y=1.765
+ $X2=0 $Y2=0
cc_295 N_A_27_74#_c_270_n N_A_206_368#_c_578_n 0.00746249f $X=5.445 $Y=0.392
+ $X2=0 $Y2=0
cc_296 N_A_27_74#_c_272_n N_A_206_368#_c_578_n 0.00372092f $X=5.53 $Y=1.17 $X2=0
+ $Y2=0
cc_297 N_A_27_74#_c_276_n N_A_206_368#_c_578_n 0.0222442f $X=5.68 $Y=1.335 $X2=0
+ $Y2=0
cc_298 N_A_27_74#_c_277_n N_A_206_368#_c_578_n 2.85311e-19 $X=5.68 $Y=1.245
+ $X2=0 $Y2=0
cc_299 N_A_27_74#_c_257_n N_A_206_368#_c_579_n 0.0207373f $X=4.925 $Y=1.765
+ $X2=0 $Y2=0
cc_300 N_A_27_74#_c_270_n N_A_206_368#_c_579_n 0.00160029f $X=5.445 $Y=0.392
+ $X2=0 $Y2=0
cc_301 N_A_27_74#_c_272_n N_A_206_368#_c_579_n 0.00118555f $X=5.53 $Y=1.17 $X2=0
+ $Y2=0
cc_302 N_A_27_74#_c_276_n N_A_206_368#_c_579_n 0.00171869f $X=5.68 $Y=1.335
+ $X2=0 $Y2=0
cc_303 N_A_27_74#_c_277_n N_A_206_368#_c_579_n 0.0176236f $X=5.68 $Y=1.245 $X2=0
+ $Y2=0
cc_304 N_A_27_74#_c_281_n N_A_206_368#_c_592_n 0.0034289f $X=4.925 $Y=2.045
+ $X2=0 $Y2=0
cc_305 N_A_27_74#_c_248_n N_A_206_368#_c_580_n 0.015168f $X=0.955 $Y=1.765 $X2=0
+ $Y2=0
cc_306 N_A_27_74#_c_261_n N_A_206_368#_c_580_n 3.53314e-19 $X=0.927 $Y=1.378
+ $X2=0 $Y2=0
cc_307 N_A_27_74#_c_263_n N_A_206_368#_c_580_n 0.0164129f $X=2.36 $Y=0.815 $X2=0
+ $Y2=0
cc_308 N_A_27_74#_c_264_n N_A_206_368#_c_580_n 0.00273349f $X=2.445 $Y=0.73
+ $X2=0 $Y2=0
cc_309 N_A_27_74#_c_375_p N_A_206_368#_c_580_n 5.01237e-19 $X=0.927 $Y=0.87
+ $X2=0 $Y2=0
cc_310 N_A_27_74#_c_269_n N_A_753_284#_M1007_d 0.00781679f $X=4.645 $Y=0.865
+ $X2=-0.19 $Y2=-0.245
cc_311 N_A_27_74#_c_334_p N_A_753_284#_M1007_d 0.00748701f $X=4.73 $Y=0.78
+ $X2=-0.19 $Y2=-0.245
cc_312 N_A_27_74#_c_270_n N_A_753_284#_M1007_d 0.00270947f $X=5.445 $Y=0.392
+ $X2=-0.19 $Y2=-0.245
cc_313 N_A_27_74#_c_271_n N_A_753_284#_M1007_d 0.00253073f $X=4.815 $Y=0.392
+ $X2=-0.19 $Y2=-0.245
cc_314 N_A_27_74#_c_251_n N_A_753_284#_c_759_n 0.00410905f $X=3.12 $Y=1.735
+ $X2=0 $Y2=0
cc_315 N_A_27_74#_c_256_n N_A_753_284#_c_759_n 0.00430052f $X=3.12 $Y=1.165
+ $X2=0 $Y2=0
cc_316 N_A_27_74#_c_268_n N_A_753_284#_c_759_n 0.010166f $X=3.555 $Y=1.75 $X2=0
+ $Y2=0
cc_317 N_A_27_74#_c_269_n N_A_753_284#_c_759_n 0.00579297f $X=4.645 $Y=0.865
+ $X2=0 $Y2=0
cc_318 N_A_27_74#_c_268_n N_A_753_284#_c_760_n 0.00334484f $X=3.555 $Y=1.75
+ $X2=0 $Y2=0
cc_319 N_A_27_74#_c_290_n N_A_753_284#_c_760_n 0.0196919f $X=3.39 $Y=1.9 $X2=0
+ $Y2=0
cc_320 N_A_27_74#_c_280_n N_A_753_284#_c_766_n 0.0306527f $X=3.435 $Y=2.15 $X2=0
+ $Y2=0
cc_321 N_A_27_74#_c_290_n N_A_753_284#_c_766_n 0.00487061f $X=3.39 $Y=1.9 $X2=0
+ $Y2=0
cc_322 N_A_27_74#_c_265_n N_A_753_284#_M1004_g 4.07545e-19 $X=3.47 $Y=0.34 $X2=0
+ $Y2=0
cc_323 N_A_27_74#_c_267_n N_A_753_284#_M1004_g 0.00137293f $X=3.555 $Y=0.78
+ $X2=0 $Y2=0
cc_324 N_A_27_74#_c_268_n N_A_753_284#_M1004_g 0.00316409f $X=3.555 $Y=1.75
+ $X2=0 $Y2=0
cc_325 N_A_27_74#_c_269_n N_A_753_284#_M1004_g 0.0117681f $X=4.645 $Y=0.865
+ $X2=0 $Y2=0
cc_326 N_A_27_74#_c_268_n N_A_753_284#_c_762_n 0.0262118f $X=3.555 $Y=1.75 $X2=0
+ $Y2=0
cc_327 N_A_27_74#_c_269_n N_A_753_284#_c_762_n 0.0628209f $X=4.645 $Y=0.865
+ $X2=0 $Y2=0
cc_328 N_A_27_74#_c_269_n N_A_753_284#_c_763_n 0.0153523f $X=4.645 $Y=0.865
+ $X2=0 $Y2=0
cc_329 N_A_27_74#_c_281_n N_A_753_284#_c_764_n 0.00415934f $X=4.925 $Y=2.045
+ $X2=0 $Y2=0
cc_330 N_A_27_74#_c_257_n N_A_753_284#_c_764_n 0.00322002f $X=4.925 $Y=1.765
+ $X2=0 $Y2=0
cc_331 N_A_27_74#_c_269_n N_A_558_445#_M1007_g 0.0123068f $X=4.645 $Y=0.865
+ $X2=0 $Y2=0
cc_332 N_A_27_74#_c_334_p N_A_558_445#_M1007_g 0.00458856f $X=4.73 $Y=0.78 $X2=0
+ $Y2=0
cc_333 N_A_27_74#_c_271_n N_A_558_445#_M1007_g 0.00279328f $X=4.815 $Y=0.392
+ $X2=0 $Y2=0
cc_334 N_A_27_74#_c_281_n N_A_558_445#_c_817_n 0.0287818f $X=4.925 $Y=2.045
+ $X2=0 $Y2=0
cc_335 N_A_27_74#_c_257_n N_A_558_445#_c_817_n 0.0147796f $X=4.925 $Y=1.765
+ $X2=0 $Y2=0
cc_336 N_A_27_74#_c_251_n N_A_558_445#_c_818_n 0.00442182f $X=3.12 $Y=1.735
+ $X2=0 $Y2=0
cc_337 N_A_27_74#_c_280_n N_A_558_445#_c_818_n 0.00265258f $X=3.435 $Y=2.15
+ $X2=0 $Y2=0
cc_338 N_A_27_74#_c_268_n N_A_558_445#_c_818_n 0.0290653f $X=3.555 $Y=1.75 $X2=0
+ $Y2=0
cc_339 N_A_27_74#_c_290_n N_A_558_445#_c_818_n 0.00899012f $X=3.39 $Y=1.9 $X2=0
+ $Y2=0
cc_340 N_A_27_74#_c_251_n N_A_558_445#_c_819_n 0.0136932f $X=3.12 $Y=1.735 $X2=0
+ $Y2=0
cc_341 N_A_27_74#_c_256_n N_A_558_445#_c_819_n 0.00498074f $X=3.12 $Y=1.165
+ $X2=0 $Y2=0
cc_342 N_A_27_74#_c_268_n N_A_558_445#_c_819_n 0.0192438f $X=3.555 $Y=1.75 $X2=0
+ $Y2=0
cc_343 N_A_27_74#_c_290_n N_A_558_445#_c_819_n 0.0028568f $X=3.39 $Y=1.9 $X2=0
+ $Y2=0
cc_344 N_A_27_74#_c_250_n N_A_558_445#_c_820_n 0.00664794f $X=3 $Y=1.09 $X2=0
+ $Y2=0
cc_345 N_A_27_74#_c_251_n N_A_558_445#_c_820_n 0.00663545f $X=3.12 $Y=1.735
+ $X2=0 $Y2=0
cc_346 N_A_27_74#_c_256_n N_A_558_445#_c_820_n 0.00770505f $X=3.12 $Y=1.165
+ $X2=0 $Y2=0
cc_347 N_A_27_74#_c_265_n N_A_558_445#_c_820_n 0.0168877f $X=3.47 $Y=0.34 $X2=0
+ $Y2=0
cc_348 N_A_27_74#_c_267_n N_A_558_445#_c_820_n 0.0133535f $X=3.555 $Y=0.78 $X2=0
+ $Y2=0
cc_349 N_A_27_74#_c_268_n N_A_558_445#_c_820_n 0.0351378f $X=3.555 $Y=1.75 $X2=0
+ $Y2=0
cc_350 N_A_27_74#_c_331_p N_A_558_445#_c_820_n 0.0137305f $X=3.555 $Y=0.865
+ $X2=0 $Y2=0
cc_351 N_A_27_74#_c_280_n N_A_558_445#_c_846_n 0.0116472f $X=3.435 $Y=2.15 $X2=0
+ $Y2=0
cc_352 N_A_27_74#_c_268_n N_A_558_445#_c_846_n 0.0215727f $X=3.555 $Y=1.75 $X2=0
+ $Y2=0
cc_353 N_A_27_74#_c_290_n N_A_558_445#_c_846_n 0.00905466f $X=3.39 $Y=1.9 $X2=0
+ $Y2=0
cc_354 N_A_27_74#_c_268_n N_A_558_445#_c_821_n 0.0150504f $X=3.555 $Y=1.75 $X2=0
+ $Y2=0
cc_355 N_A_27_74#_c_258_n N_A_1290_102#_c_894_n 0.0256002f $X=6.09 $Y=0.365
+ $X2=0 $Y2=0
cc_356 N_A_27_74#_M1002_g N_A_1290_102#_c_901_n 0.0256002f $X=6.165 $Y=0.85
+ $X2=0 $Y2=0
cc_357 N_A_27_74#_c_277_n N_A_1290_102#_c_901_n 0.00247443f $X=5.68 $Y=1.245
+ $X2=0 $Y2=0
cc_358 N_A_27_74#_c_254_n N_A_1290_102#_c_906_n 4.08739e-19 $X=6.09 $Y=1.245
+ $X2=0 $Y2=0
cc_359 N_A_27_74#_c_270_n N_A_1000_424#_M1012_d 0.00473057f $X=5.445 $Y=0.392
+ $X2=-0.19 $Y2=-0.245
cc_360 N_A_27_74#_c_272_n N_A_1000_424#_M1012_d 0.00942711f $X=5.53 $Y=1.17
+ $X2=-0.19 $Y2=-0.245
cc_361 N_A_27_74#_c_252_n N_A_1000_424#_c_1069_n 0.00982957f $X=5.515 $Y=1.765
+ $X2=0 $Y2=0
cc_362 N_A_27_74#_c_254_n N_A_1000_424#_c_1059_n 0.00207122f $X=6.09 $Y=1.245
+ $X2=0 $Y2=0
cc_363 N_A_27_74#_c_276_n N_A_1000_424#_c_1059_n 0.010353f $X=5.68 $Y=1.335
+ $X2=0 $Y2=0
cc_364 N_A_27_74#_c_277_n N_A_1000_424#_c_1059_n 0.00332694f $X=5.68 $Y=1.245
+ $X2=0 $Y2=0
cc_365 N_A_27_74#_c_252_n N_A_1000_424#_c_1060_n 0.00882714f $X=5.515 $Y=1.765
+ $X2=0 $Y2=0
cc_366 N_A_27_74#_c_253_n N_A_1000_424#_c_1060_n 0.00599434f $X=5.59 $Y=1.69
+ $X2=0 $Y2=0
cc_367 N_A_27_74#_c_276_n N_A_1000_424#_c_1060_n 0.0212885f $X=5.68 $Y=1.335
+ $X2=0 $Y2=0
cc_368 N_A_27_74#_c_277_n N_A_1000_424#_c_1060_n 9.89943e-19 $X=5.68 $Y=1.245
+ $X2=0 $Y2=0
cc_369 N_A_27_74#_c_253_n N_A_1000_424#_c_1061_n 0.00336429f $X=5.59 $Y=1.69
+ $X2=0 $Y2=0
cc_370 N_A_27_74#_c_254_n N_A_1000_424#_c_1061_n 0.0103862f $X=6.09 $Y=1.245
+ $X2=0 $Y2=0
cc_371 N_A_27_74#_M1002_g N_A_1000_424#_c_1061_n 0.00656427f $X=6.165 $Y=0.85
+ $X2=0 $Y2=0
cc_372 N_A_27_74#_c_272_n N_A_1000_424#_c_1061_n 0.00900667f $X=5.53 $Y=1.17
+ $X2=0 $Y2=0
cc_373 N_A_27_74#_c_276_n N_A_1000_424#_c_1061_n 0.0207508f $X=5.68 $Y=1.335
+ $X2=0 $Y2=0
cc_374 N_A_27_74#_c_277_n N_A_1000_424#_c_1061_n 0.00179411f $X=5.68 $Y=1.245
+ $X2=0 $Y2=0
cc_375 N_A_27_74#_M1002_g N_A_1000_424#_c_1062_n 0.00675215f $X=6.165 $Y=0.85
+ $X2=0 $Y2=0
cc_376 N_A_27_74#_c_258_n N_A_1000_424#_c_1062_n 0.00302649f $X=6.09 $Y=0.365
+ $X2=0 $Y2=0
cc_377 N_A_27_74#_c_272_n N_A_1000_424#_c_1062_n 0.01939f $X=5.53 $Y=1.17 $X2=0
+ $Y2=0
cc_378 N_A_27_74#_c_273_n N_A_1000_424#_c_1062_n 0.0264072f $X=6.075 $Y=0.365
+ $X2=0 $Y2=0
cc_379 N_A_27_74#_c_276_n N_A_1000_424#_c_1062_n 0.00372461f $X=5.68 $Y=1.335
+ $X2=0 $Y2=0
cc_380 N_A_27_74#_c_277_n N_A_1000_424#_c_1062_n 0.00286745f $X=5.68 $Y=1.245
+ $X2=0 $Y2=0
cc_381 N_A_27_74#_c_254_n N_A_1000_424#_c_1064_n 0.00169205f $X=6.09 $Y=1.245
+ $X2=0 $Y2=0
cc_382 N_A_27_74#_c_286_n N_VPWR_M1017_d 0.00224397f $X=0.755 $Y=1.805 $X2=-0.19
+ $Y2=-0.245
cc_383 N_A_27_74#_c_248_n N_VPWR_c_1238_n 0.0181688f $X=0.955 $Y=1.765 $X2=0
+ $Y2=0
cc_384 N_A_27_74#_c_285_n N_VPWR_c_1238_n 0.0617165f $X=0.28 $Y=1.985 $X2=0
+ $Y2=0
cc_385 N_A_27_74#_c_286_n N_VPWR_c_1238_n 0.0161054f $X=0.755 $Y=1.805 $X2=0
+ $Y2=0
cc_386 N_A_27_74#_c_281_n N_VPWR_c_1245_n 0.00314961f $X=4.925 $Y=2.045 $X2=0
+ $Y2=0
cc_387 N_A_27_74#_c_280_n N_VPWR_c_1249_n 6.43532e-19 $X=3.435 $Y=2.15 $X2=0
+ $Y2=0
cc_388 N_A_27_74#_c_285_n N_VPWR_c_1253_n 0.0145938f $X=0.28 $Y=1.985 $X2=0
+ $Y2=0
cc_389 N_A_27_74#_c_248_n N_VPWR_c_1254_n 0.00413917f $X=0.955 $Y=1.765 $X2=0
+ $Y2=0
cc_390 N_A_27_74#_c_248_n N_VPWR_c_1255_n 0.00285153f $X=0.955 $Y=1.765 $X2=0
+ $Y2=0
cc_391 N_A_27_74#_c_248_n N_VPWR_c_1237_n 0.00822528f $X=0.955 $Y=1.765 $X2=0
+ $Y2=0
cc_392 N_A_27_74#_c_281_n N_VPWR_c_1237_n 0.00395887f $X=4.925 $Y=2.045 $X2=0
+ $Y2=0
cc_393 N_A_27_74#_c_285_n N_VPWR_c_1237_n 0.0120466f $X=0.28 $Y=1.985 $X2=0
+ $Y2=0
cc_394 N_A_27_74#_c_251_n N_A_451_503#_c_1355_n 0.00281437f $X=3.12 $Y=1.735
+ $X2=0 $Y2=0
cc_395 N_A_27_74#_c_250_n N_A_451_503#_c_1356_n 5.15818e-19 $X=3 $Y=1.09 $X2=0
+ $Y2=0
cc_396 N_A_27_74#_c_265_n N_A_451_503#_c_1356_n 0.0125903f $X=3.47 $Y=0.34 $X2=0
+ $Y2=0
cc_397 N_A_27_74#_c_250_n N_A_451_503#_c_1357_n 0.00136449f $X=3 $Y=1.09 $X2=0
+ $Y2=0
cc_398 N_A_27_74#_c_265_n N_A_451_503#_c_1357_n 0.00426655f $X=3.47 $Y=0.34
+ $X2=0 $Y2=0
cc_399 N_A_27_74#_c_296_n N_VGND_M1025_d 0.00654624f $X=0.755 $Y=0.87 $X2=-0.19
+ $Y2=-0.245
cc_400 N_A_27_74#_c_261_n N_VGND_M1025_d 0.00147064f $X=0.927 $Y=1.378 $X2=-0.19
+ $Y2=-0.245
cc_401 N_A_27_74#_c_375_p N_VGND_M1025_d 0.00474637f $X=0.927 $Y=0.87 $X2=-0.19
+ $Y2=-0.245
cc_402 N_A_27_74#_c_263_n N_VGND_M1024_s 0.017344f $X=2.36 $Y=0.815 $X2=0 $Y2=0
cc_403 N_A_27_74#_c_264_n N_VGND_M1024_s 0.00216437f $X=2.445 $Y=0.73 $X2=0
+ $Y2=0
cc_404 N_A_27_74#_c_269_n N_VGND_M1004_d 0.00284628f $X=4.645 $Y=0.865 $X2=0
+ $Y2=0
cc_405 N_A_27_74#_c_248_n N_VGND_c_1447_n 6.03634e-19 $X=0.955 $Y=1.765 $X2=0
+ $Y2=0
cc_406 N_A_27_74#_c_249_n N_VGND_c_1447_n 0.00520561f $X=1.14 $Y=1.22 $X2=0
+ $Y2=0
cc_407 N_A_27_74#_c_259_n N_VGND_c_1447_n 0.00830381f $X=0.28 $Y=0.515 $X2=0
+ $Y2=0
cc_408 N_A_27_74#_c_296_n N_VGND_c_1447_n 0.0103246f $X=0.755 $Y=0.87 $X2=0
+ $Y2=0
cc_409 N_A_27_74#_c_375_p N_VGND_c_1447_n 0.0218924f $X=0.927 $Y=0.87 $X2=0
+ $Y2=0
cc_410 N_A_27_74#_c_263_n N_VGND_c_1448_n 0.025747f $X=2.36 $Y=0.815 $X2=0 $Y2=0
cc_411 N_A_27_74#_c_264_n N_VGND_c_1448_n 0.0104593f $X=2.445 $Y=0.73 $X2=0
+ $Y2=0
cc_412 N_A_27_74#_c_266_n N_VGND_c_1448_n 0.0148933f $X=2.53 $Y=0.34 $X2=0 $Y2=0
cc_413 N_A_27_74#_c_263_n N_VGND_c_1449_n 0.00241577f $X=2.36 $Y=0.815 $X2=0
+ $Y2=0
cc_414 N_A_27_74#_c_265_n N_VGND_c_1449_n 0.0721609f $X=3.47 $Y=0.34 $X2=0 $Y2=0
cc_415 N_A_27_74#_c_266_n N_VGND_c_1449_n 0.0115448f $X=2.53 $Y=0.34 $X2=0 $Y2=0
cc_416 N_A_27_74#_c_265_n N_VGND_c_1450_n 0.00845988f $X=3.47 $Y=0.34 $X2=0
+ $Y2=0
cc_417 N_A_27_74#_c_267_n N_VGND_c_1450_n 0.00372338f $X=3.555 $Y=0.78 $X2=0
+ $Y2=0
cc_418 N_A_27_74#_c_269_n N_VGND_c_1450_n 0.0220573f $X=4.645 $Y=0.865 $X2=0
+ $Y2=0
cc_419 N_A_27_74#_c_334_p N_VGND_c_1450_n 0.00406641f $X=4.73 $Y=0.78 $X2=0
+ $Y2=0
cc_420 N_A_27_74#_c_271_n N_VGND_c_1450_n 0.0159558f $X=4.815 $Y=0.392 $X2=0
+ $Y2=0
cc_421 N_A_27_74#_c_258_n N_VGND_c_1451_n 0.00286833f $X=6.09 $Y=0.365 $X2=0
+ $Y2=0
cc_422 N_A_27_74#_c_273_n N_VGND_c_1451_n 0.0117193f $X=6.075 $Y=0.365 $X2=0
+ $Y2=0
cc_423 N_A_27_74#_c_258_n N_VGND_c_1457_n 0.0125151f $X=6.09 $Y=0.365 $X2=0
+ $Y2=0
cc_424 N_A_27_74#_c_270_n N_VGND_c_1457_n 0.0414454f $X=5.445 $Y=0.392 $X2=0
+ $Y2=0
cc_425 N_A_27_74#_c_271_n N_VGND_c_1457_n 0.012207f $X=4.815 $Y=0.392 $X2=0
+ $Y2=0
cc_426 N_A_27_74#_c_273_n N_VGND_c_1457_n 0.0396429f $X=6.075 $Y=0.365 $X2=0
+ $Y2=0
cc_427 N_A_27_74#_c_275_n N_VGND_c_1457_n 0.0120286f $X=5.53 $Y=0.392 $X2=0
+ $Y2=0
cc_428 N_A_27_74#_c_259_n N_VGND_c_1463_n 0.0145323f $X=0.28 $Y=0.515 $X2=0
+ $Y2=0
cc_429 N_A_27_74#_c_296_n N_VGND_c_1463_n 0.00211533f $X=0.755 $Y=0.87 $X2=0
+ $Y2=0
cc_430 N_A_27_74#_c_249_n N_VGND_c_1464_n 0.00336054f $X=1.14 $Y=1.22 $X2=0
+ $Y2=0
cc_431 N_A_27_74#_c_263_n N_VGND_c_1464_n 0.0102896f $X=2.36 $Y=0.815 $X2=0
+ $Y2=0
cc_432 N_A_27_74#_c_375_p N_VGND_c_1464_n 9.24443e-19 $X=0.927 $Y=0.87 $X2=0
+ $Y2=0
cc_433 N_A_27_74#_c_249_n N_VGND_c_1471_n 0.00439202f $X=1.14 $Y=1.22 $X2=0
+ $Y2=0
cc_434 N_A_27_74#_c_258_n N_VGND_c_1471_n 0.0174291f $X=6.09 $Y=0.365 $X2=0
+ $Y2=0
cc_435 N_A_27_74#_c_259_n N_VGND_c_1471_n 0.0119861f $X=0.28 $Y=0.515 $X2=0
+ $Y2=0
cc_436 N_A_27_74#_c_296_n N_VGND_c_1471_n 0.00479362f $X=0.755 $Y=0.87 $X2=0
+ $Y2=0
cc_437 N_A_27_74#_c_263_n N_VGND_c_1471_n 0.0237784f $X=2.36 $Y=0.815 $X2=0
+ $Y2=0
cc_438 N_A_27_74#_c_265_n N_VGND_c_1471_n 0.0376224f $X=3.47 $Y=0.34 $X2=0 $Y2=0
cc_439 N_A_27_74#_c_266_n N_VGND_c_1471_n 0.00582224f $X=2.53 $Y=0.34 $X2=0
+ $Y2=0
cc_440 N_A_27_74#_c_269_n N_VGND_c_1471_n 0.0244708f $X=4.645 $Y=0.865 $X2=0
+ $Y2=0
cc_441 N_A_27_74#_c_270_n N_VGND_c_1471_n 0.0238428f $X=5.445 $Y=0.392 $X2=0
+ $Y2=0
cc_442 N_A_27_74#_c_271_n N_VGND_c_1471_n 0.00661303f $X=4.815 $Y=0.392 $X2=0
+ $Y2=0
cc_443 N_A_27_74#_c_273_n N_VGND_c_1471_n 0.0208588f $X=6.075 $Y=0.365 $X2=0
+ $Y2=0
cc_444 N_A_27_74#_c_375_p N_VGND_c_1471_n 0.00350516f $X=0.927 $Y=0.87 $X2=0
+ $Y2=0
cc_445 N_A_27_74#_c_275_n N_VGND_c_1471_n 0.0064033f $X=5.53 $Y=0.392 $X2=0
+ $Y2=0
cc_446 N_A_27_74#_c_269_n A_717_102# 0.002402f $X=4.645 $Y=0.865 $X2=-0.19
+ $Y2=-0.245
cc_447 N_D_c_513_n N_A_206_368#_c_570_n 0.00903828f $X=2.57 $Y=1.125 $X2=0 $Y2=0
cc_448 N_D_c_518_n N_A_206_368#_c_581_n 0.00106267f $X=1.99 $Y=2.19 $X2=0 $Y2=0
cc_449 N_D_c_519_n N_A_206_368#_c_581_n 0.02828f $X=1.99 $Y=2.19 $X2=0 $Y2=0
cc_450 N_D_c_520_n N_A_206_368#_c_581_n 0.00324039f $X=1.99 $Y=2.025 $X2=0 $Y2=0
cc_451 N_D_c_515_n N_A_206_368#_c_581_n 0.0308807f $X=2.21 $Y=1.29 $X2=0 $Y2=0
cc_452 D N_A_206_368#_c_581_n 0.0163967f $X=2.16 $Y=1.665 $X2=0 $Y2=0
cc_453 N_D_c_519_n N_A_206_368#_c_582_n 0.00403951f $X=1.99 $Y=2.19 $X2=0 $Y2=0
cc_454 N_D_c_520_n N_A_206_368#_c_582_n 0.00107077f $X=1.99 $Y=2.025 $X2=0 $Y2=0
cc_455 N_D_c_517_n N_A_206_368#_c_583_n 0.0089361f $X=2.18 $Y=2.44 $X2=0 $Y2=0
cc_456 N_D_c_519_n N_A_206_368#_c_583_n 0.0050378f $X=1.99 $Y=2.19 $X2=0 $Y2=0
cc_457 N_D_c_517_n N_A_206_368#_c_585_n 0.00412021f $X=2.18 $Y=2.44 $X2=0 $Y2=0
cc_458 N_D_c_518_n N_A_206_368#_c_585_n 0.0142713f $X=1.99 $Y=2.19 $X2=0 $Y2=0
cc_459 N_D_c_519_n N_A_206_368#_c_585_n 0.00885036f $X=1.99 $Y=2.19 $X2=0 $Y2=0
cc_460 N_D_c_520_n N_A_206_368#_c_585_n 0.00131293f $X=1.99 $Y=2.025 $X2=0 $Y2=0
cc_461 D N_A_206_368#_c_574_n 0.0171608f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_462 N_D_c_517_n N_A_206_368#_c_586_n 0.0168782f $X=2.18 $Y=2.44 $X2=0 $Y2=0
cc_463 N_D_c_518_n N_A_206_368#_c_586_n 0.0159503f $X=1.99 $Y=2.19 $X2=0 $Y2=0
cc_464 N_D_c_519_n N_A_206_368#_c_586_n 0.00157307f $X=1.99 $Y=2.19 $X2=0 $Y2=0
cc_465 N_D_c_520_n N_A_206_368#_c_576_n 0.00611417f $X=1.99 $Y=2.025 $X2=0 $Y2=0
cc_466 D N_A_206_368#_c_576_n 0.0267182f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_467 D N_A_206_368#_c_577_n 0.0013489f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_468 N_D_c_513_n N_A_206_368#_c_580_n 0.00936782f $X=2.57 $Y=1.125 $X2=0 $Y2=0
cc_469 D N_A_206_368#_c_580_n 0.00337034f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_470 N_D_c_515_n N_A_206_368#_c_580_n 0.0165052f $X=2.21 $Y=1.29 $X2=0 $Y2=0
cc_471 N_D_c_513_n N_A_558_445#_c_820_n 2.71632e-19 $X=2.57 $Y=1.125 $X2=0 $Y2=0
cc_472 N_D_c_517_n N_VPWR_c_1249_n 0.00418282f $X=2.18 $Y=2.44 $X2=0 $Y2=0
cc_473 N_D_c_517_n N_VPWR_c_1255_n 0.00427869f $X=2.18 $Y=2.44 $X2=0 $Y2=0
cc_474 N_D_c_517_n N_VPWR_c_1237_n 0.00537853f $X=2.18 $Y=2.44 $X2=0 $Y2=0
cc_475 N_D_c_519_n N_A_451_503#_c_1355_n 0.00146835f $X=1.99 $Y=2.19 $X2=0 $Y2=0
cc_476 N_D_c_520_n N_A_451_503#_c_1355_n 0.0173578f $X=1.99 $Y=2.025 $X2=0 $Y2=0
cc_477 D N_A_451_503#_c_1355_n 0.0413916f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_478 N_D_c_515_n N_A_451_503#_c_1355_n 0.0047987f $X=2.21 $Y=1.29 $X2=0 $Y2=0
cc_479 N_D_c_513_n N_A_451_503#_c_1356_n 0.0014192f $X=2.57 $Y=1.125 $X2=0 $Y2=0
cc_480 N_D_c_517_n N_A_451_503#_c_1359_n 3.9836e-19 $X=2.18 $Y=2.44 $X2=0 $Y2=0
cc_481 N_D_c_518_n N_A_451_503#_c_1359_n 0.0120068f $X=1.99 $Y=2.19 $X2=0 $Y2=0
cc_482 N_D_c_519_n N_A_451_503#_c_1359_n 0.00402689f $X=1.99 $Y=2.19 $X2=0 $Y2=0
cc_483 D N_A_451_503#_c_1359_n 0.00201546f $X=2.16 $Y=1.665 $X2=0 $Y2=0
cc_484 N_D_c_513_n N_A_451_503#_c_1357_n 0.00573263f $X=2.57 $Y=1.125 $X2=0
+ $Y2=0
cc_485 D N_A_451_503#_c_1357_n 0.00870101f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_486 N_D_c_515_n N_A_451_503#_c_1357_n 0.00400841f $X=2.21 $Y=1.29 $X2=0 $Y2=0
cc_487 N_D_c_513_n N_VGND_c_1448_n 3.10895e-19 $X=2.57 $Y=1.125 $X2=0 $Y2=0
cc_488 N_A_206_368#_c_586_n N_A_753_284#_M1031_d 0.00483417f $X=5.035 $Y=2.71
+ $X2=0 $Y2=0
cc_489 N_A_206_368#_c_586_n N_A_753_284#_c_766_n 0.0105026f $X=5.035 $Y=2.71
+ $X2=0 $Y2=0
cc_490 N_A_206_368#_M1014_g N_A_753_284#_M1004_g 0.0346499f $X=3.51 $Y=0.72
+ $X2=0 $Y2=0
cc_491 N_A_206_368#_c_578_n N_A_753_284#_c_763_n 0.0270425f $X=5.14 $Y=1.285
+ $X2=0 $Y2=0
cc_492 N_A_206_368#_c_579_n N_A_753_284#_c_763_n 0.00328335f $X=5.14 $Y=1.285
+ $X2=0 $Y2=0
cc_493 N_A_206_368#_c_586_n N_A_753_284#_c_764_n 0.0160525f $X=5.035 $Y=2.71
+ $X2=0 $Y2=0
cc_494 N_A_206_368#_c_575_n N_A_753_284#_c_764_n 0.041391f $X=5.12 $Y=2.625
+ $X2=0 $Y2=0
cc_495 N_A_206_368#_c_586_n N_A_558_445#_M1028_d 0.00583843f $X=5.035 $Y=2.71
+ $X2=0 $Y2=0
cc_496 N_A_206_368#_M1012_g N_A_558_445#_M1007_g 0.0270846f $X=5.015 $Y=0.655
+ $X2=0 $Y2=0
cc_497 N_A_206_368#_c_578_n N_A_558_445#_M1007_g 2.57251e-19 $X=5.14 $Y=1.285
+ $X2=0 $Y2=0
cc_498 N_A_206_368#_c_586_n N_A_558_445#_c_817_n 0.0157601f $X=5.035 $Y=2.71
+ $X2=0 $Y2=0
cc_499 N_A_206_368#_c_581_n N_A_558_445#_c_818_n 0.00354143f $X=2.625 $Y=1.74
+ $X2=0 $Y2=0
cc_500 N_A_206_368#_c_583_n N_A_558_445#_c_818_n 0.00129974f $X=2.715 $Y=2.15
+ $X2=0 $Y2=0
cc_501 N_A_206_368#_M1014_g N_A_558_445#_c_820_n 0.00326752f $X=3.51 $Y=0.72
+ $X2=0 $Y2=0
cc_502 N_A_206_368#_c_586_n N_A_558_445#_c_846_n 0.0755489f $X=5.035 $Y=2.71
+ $X2=0 $Y2=0
cc_503 N_A_206_368#_c_583_n N_A_558_445#_c_859_n 0.00182039f $X=2.715 $Y=2.15
+ $X2=0 $Y2=0
cc_504 N_A_206_368#_c_586_n N_A_558_445#_c_859_n 0.0137412f $X=5.035 $Y=2.71
+ $X2=0 $Y2=0
cc_505 N_A_206_368#_c_586_n N_A_558_445#_c_821_n 0.00283163f $X=5.035 $Y=2.71
+ $X2=0 $Y2=0
cc_506 N_A_206_368#_c_584_n N_A_1290_102#_c_914_n 0.0180126f $X=5.965 $Y=2.32
+ $X2=0 $Y2=0
cc_507 N_A_206_368#_c_589_n N_A_1290_102#_c_914_n 0.00180132f $X=6.04 $Y=2.07
+ $X2=0 $Y2=0
cc_508 N_A_206_368#_c_584_n N_A_1290_102#_c_915_n 0.016453f $X=5.965 $Y=2.32
+ $X2=0 $Y2=0
cc_509 N_A_206_368#_c_588_n N_A_1290_102#_c_915_n 0.00143078f $X=5.875 $Y=2.88
+ $X2=0 $Y2=0
cc_510 N_A_206_368#_c_589_n N_A_1290_102#_c_915_n 0.00678087f $X=6.04 $Y=2.07
+ $X2=0 $Y2=0
cc_511 N_A_206_368#_c_575_n N_A_1000_424#_M1000_d 0.00788988f $X=5.12 $Y=2.625
+ $X2=0 $Y2=0
cc_512 N_A_206_368#_c_588_n N_A_1000_424#_M1000_d 0.0163467f $X=5.875 $Y=2.88
+ $X2=0 $Y2=0
cc_513 N_A_206_368#_c_592_n N_A_1000_424#_M1000_d 0.00389937f $X=5.12 $Y=2.71
+ $X2=0 $Y2=0
cc_514 N_A_206_368#_c_584_n N_A_1000_424#_c_1069_n 0.0117519f $X=5.965 $Y=2.32
+ $X2=0 $Y2=0
cc_515 N_A_206_368#_c_575_n N_A_1000_424#_c_1069_n 0.0647087f $X=5.12 $Y=2.625
+ $X2=0 $Y2=0
cc_516 N_A_206_368#_c_588_n N_A_1000_424#_c_1069_n 0.0254969f $X=5.875 $Y=2.88
+ $X2=0 $Y2=0
cc_517 N_A_206_368#_c_589_n N_A_1000_424#_c_1069_n 0.0439164f $X=6.04 $Y=2.07
+ $X2=0 $Y2=0
cc_518 N_A_206_368#_c_584_n N_A_1000_424#_c_1059_n 0.00172034f $X=5.965 $Y=2.32
+ $X2=0 $Y2=0
cc_519 N_A_206_368#_c_589_n N_A_1000_424#_c_1059_n 0.0110698f $X=6.04 $Y=2.07
+ $X2=0 $Y2=0
cc_520 N_A_206_368#_c_575_n N_A_1000_424#_c_1060_n 0.0135294f $X=5.12 $Y=2.625
+ $X2=0 $Y2=0
cc_521 N_A_206_368#_c_584_n N_A_1000_424#_c_1063_n 0.00203097f $X=5.965 $Y=2.32
+ $X2=0 $Y2=0
cc_522 N_A_206_368#_c_589_n N_A_1000_424#_c_1063_n 0.0151551f $X=6.04 $Y=2.07
+ $X2=0 $Y2=0
cc_523 N_A_206_368#_c_584_n N_A_1000_424#_c_1064_n 2.27652e-19 $X=5.965 $Y=2.32
+ $X2=0 $Y2=0
cc_524 N_A_206_368#_c_589_n N_A_1000_424#_c_1064_n 0.00148051f $X=6.04 $Y=2.07
+ $X2=0 $Y2=0
cc_525 N_A_206_368#_c_584_n N_A_1000_424#_c_1065_n 7.279e-19 $X=5.965 $Y=2.32
+ $X2=0 $Y2=0
cc_526 N_A_206_368#_c_586_n N_VPWR_M1022_s 0.0188104f $X=5.035 $Y=2.71 $X2=0
+ $Y2=0
cc_527 N_A_206_368#_c_586_n N_VPWR_M1005_d 0.00808693f $X=5.035 $Y=2.71 $X2=0
+ $Y2=0
cc_528 N_A_206_368#_c_585_n N_VPWR_c_1238_n 0.0624043f $X=1.267 $Y=2.625 $X2=0
+ $Y2=0
cc_529 N_A_206_368#_c_584_n N_VPWR_c_1239_n 4.96348e-19 $X=5.965 $Y=2.32 $X2=0
+ $Y2=0
cc_530 N_A_206_368#_c_588_n N_VPWR_c_1239_n 0.00769846f $X=5.875 $Y=2.88 $X2=0
+ $Y2=0
cc_531 N_A_206_368#_c_589_n N_VPWR_c_1239_n 0.0170546f $X=6.04 $Y=2.07 $X2=0
+ $Y2=0
cc_532 N_A_206_368#_c_584_n N_VPWR_c_1245_n 7.88928e-19 $X=5.965 $Y=2.32 $X2=0
+ $Y2=0
cc_533 N_A_206_368#_c_586_n N_VPWR_c_1245_n 0.0133099f $X=5.035 $Y=2.71 $X2=0
+ $Y2=0
cc_534 N_A_206_368#_c_588_n N_VPWR_c_1245_n 0.0393823f $X=5.875 $Y=2.88 $X2=0
+ $Y2=0
cc_535 N_A_206_368#_c_592_n N_VPWR_c_1245_n 0.00707028f $X=5.12 $Y=2.71 $X2=0
+ $Y2=0
cc_536 N_A_206_368#_c_583_n N_VPWR_c_1249_n 6.43532e-19 $X=2.715 $Y=2.15 $X2=0
+ $Y2=0
cc_537 N_A_206_368#_c_586_n N_VPWR_c_1249_n 0.0433683f $X=5.035 $Y=2.71 $X2=0
+ $Y2=0
cc_538 N_A_206_368#_c_585_n N_VPWR_c_1254_n 0.0135613f $X=1.267 $Y=2.625 $X2=0
+ $Y2=0
cc_539 N_A_206_368#_c_586_n N_VPWR_c_1254_n 0.0030692f $X=5.035 $Y=2.71 $X2=0
+ $Y2=0
cc_540 N_A_206_368#_c_585_n N_VPWR_c_1255_n 9.55366e-19 $X=1.267 $Y=2.625 $X2=0
+ $Y2=0
cc_541 N_A_206_368#_c_586_n N_VPWR_c_1255_n 0.0337559f $X=5.035 $Y=2.71 $X2=0
+ $Y2=0
cc_542 N_A_206_368#_c_586_n N_VPWR_c_1256_n 0.0242244f $X=5.035 $Y=2.71 $X2=0
+ $Y2=0
cc_543 N_A_206_368#_c_585_n N_VPWR_c_1237_n 0.0123337f $X=1.267 $Y=2.625 $X2=0
+ $Y2=0
cc_544 N_A_206_368#_c_586_n N_VPWR_c_1237_n 0.0893229f $X=5.035 $Y=2.71 $X2=0
+ $Y2=0
cc_545 N_A_206_368#_c_588_n N_VPWR_c_1237_n 0.0355191f $X=5.875 $Y=2.88 $X2=0
+ $Y2=0
cc_546 N_A_206_368#_c_592_n N_VPWR_c_1237_n 0.00614846f $X=5.12 $Y=2.71 $X2=0
+ $Y2=0
cc_547 N_A_206_368#_c_586_n N_A_451_503#_M1022_d 0.00666725f $X=5.035 $Y=2.71
+ $X2=0 $Y2=0
cc_548 N_A_206_368#_c_581_n N_A_451_503#_c_1355_n 0.0103793f $X=2.625 $Y=1.74
+ $X2=0 $Y2=0
cc_549 N_A_206_368#_c_582_n N_A_451_503#_c_1355_n 0.00725576f $X=2.715 $Y=2.06
+ $X2=0 $Y2=0
cc_550 N_A_206_368#_c_583_n N_A_451_503#_c_1355_n 0.00365258f $X=2.715 $Y=2.15
+ $X2=0 $Y2=0
cc_551 N_A_206_368#_c_581_n N_A_451_503#_c_1359_n 0.00593995f $X=2.625 $Y=1.74
+ $X2=0 $Y2=0
cc_552 N_A_206_368#_c_583_n N_A_451_503#_c_1359_n 0.00503159f $X=2.715 $Y=2.15
+ $X2=0 $Y2=0
cc_553 N_A_206_368#_c_586_n N_A_451_503#_c_1359_n 0.0244923f $X=5.035 $Y=2.71
+ $X2=0 $Y2=0
cc_554 N_A_206_368#_c_581_n N_A_451_503#_c_1357_n 0.00309542f $X=2.625 $Y=1.74
+ $X2=0 $Y2=0
cc_555 N_A_206_368#_c_586_n A_702_445# 0.00166235f $X=5.035 $Y=2.71 $X2=-0.19
+ $Y2=-0.245
cc_556 N_A_206_368#_c_588_n A_1208_479# 2.57859e-19 $X=5.875 $Y=2.88 $X2=-0.19
+ $Y2=-0.245
cc_557 N_A_206_368#_c_589_n A_1208_479# 0.00503041f $X=6.04 $Y=2.07 $X2=-0.19
+ $Y2=-0.245
cc_558 N_A_206_368#_c_571_n N_VGND_c_1447_n 0.00253706f $X=1.805 $Y=0.18 $X2=0
+ $Y2=0
cc_559 N_A_206_368#_c_570_n N_VGND_c_1448_n 0.0234399f $X=3.435 $Y=0.18 $X2=0
+ $Y2=0
cc_560 N_A_206_368#_c_580_n N_VGND_c_1448_n 0.0118196f $X=1.65 $Y=1.485 $X2=0
+ $Y2=0
cc_561 N_A_206_368#_c_570_n N_VGND_c_1449_n 0.0298589f $X=3.435 $Y=0.18 $X2=0
+ $Y2=0
cc_562 N_A_206_368#_c_570_n N_VGND_c_1450_n 0.00302245f $X=3.435 $Y=0.18 $X2=0
+ $Y2=0
cc_563 N_A_206_368#_M1014_g N_VGND_c_1450_n 8.10696e-19 $X=3.51 $Y=0.72 $X2=0
+ $Y2=0
cc_564 N_A_206_368#_M1012_g N_VGND_c_1450_n 2.55276e-19 $X=5.015 $Y=0.655 $X2=0
+ $Y2=0
cc_565 N_A_206_368#_M1012_g N_VGND_c_1457_n 0.00390708f $X=5.015 $Y=0.655 $X2=0
+ $Y2=0
cc_566 N_A_206_368#_c_571_n N_VGND_c_1464_n 0.00596402f $X=1.805 $Y=0.18 $X2=0
+ $Y2=0
cc_567 N_A_206_368#_c_570_n N_VGND_c_1471_n 0.0372044f $X=3.435 $Y=0.18 $X2=0
+ $Y2=0
cc_568 N_A_206_368#_c_571_n N_VGND_c_1471_n 0.0067234f $X=1.805 $Y=0.18 $X2=0
+ $Y2=0
cc_569 N_A_206_368#_M1012_g N_VGND_c_1471_n 0.00542671f $X=5.015 $Y=0.655 $X2=0
+ $Y2=0
cc_570 N_A_753_284#_c_759_n N_A_558_445#_M1007_g 0.0289342f $X=3.855 $Y=1.51
+ $X2=0 $Y2=0
cc_571 N_A_753_284#_M1004_g N_A_558_445#_M1007_g 0.0170503f $X=3.9 $Y=0.72 $X2=0
+ $Y2=0
cc_572 N_A_753_284#_c_762_n N_A_558_445#_M1007_g 0.0174442f $X=4.645 $Y=1.285
+ $X2=0 $Y2=0
cc_573 N_A_753_284#_c_764_n N_A_558_445#_M1007_g 0.00629652f $X=4.73 $Y=2.18
+ $X2=0 $Y2=0
cc_574 N_A_753_284#_c_760_n N_A_558_445#_c_817_n 0.0241275f $X=3.855 $Y=2.06
+ $X2=0 $Y2=0
cc_575 N_A_753_284#_c_766_n N_A_558_445#_c_817_n 0.0140158f $X=3.855 $Y=2.15
+ $X2=0 $Y2=0
cc_576 N_A_753_284#_c_762_n N_A_558_445#_c_817_n 0.00423325f $X=4.645 $Y=1.285
+ $X2=0 $Y2=0
cc_577 N_A_753_284#_c_764_n N_A_558_445#_c_817_n 0.00896627f $X=4.73 $Y=2.18
+ $X2=0 $Y2=0
cc_578 N_A_753_284#_c_766_n N_A_558_445#_c_846_n 0.01555f $X=3.855 $Y=2.15 $X2=0
+ $Y2=0
cc_579 N_A_753_284#_c_764_n N_A_558_445#_c_846_n 0.0119043f $X=4.73 $Y=2.18
+ $X2=0 $Y2=0
cc_580 N_A_753_284#_c_760_n N_A_558_445#_c_824_n 0.00289887f $X=3.855 $Y=2.06
+ $X2=0 $Y2=0
cc_581 N_A_753_284#_c_766_n N_A_558_445#_c_824_n 0.00282149f $X=3.855 $Y=2.15
+ $X2=0 $Y2=0
cc_582 N_A_753_284#_c_764_n N_A_558_445#_c_824_n 0.0169832f $X=4.73 $Y=2.18
+ $X2=0 $Y2=0
cc_583 N_A_753_284#_c_760_n N_A_558_445#_c_821_n 0.0012793f $X=3.855 $Y=2.06
+ $X2=0 $Y2=0
cc_584 N_A_753_284#_c_762_n N_A_558_445#_c_821_n 0.0244168f $X=4.645 $Y=1.285
+ $X2=0 $Y2=0
cc_585 N_A_753_284#_c_764_n N_A_558_445#_c_821_n 0.0247407f $X=4.73 $Y=2.18
+ $X2=0 $Y2=0
cc_586 N_A_753_284#_c_766_n N_VPWR_c_1249_n 6.43532e-19 $X=3.855 $Y=2.15 $X2=0
+ $Y2=0
cc_587 N_A_753_284#_M1004_g N_VGND_c_1449_n 0.00481372f $X=3.9 $Y=0.72 $X2=0
+ $Y2=0
cc_588 N_A_753_284#_M1004_g N_VGND_c_1450_n 0.00211756f $X=3.9 $Y=0.72 $X2=0
+ $Y2=0
cc_589 N_A_753_284#_M1004_g N_VGND_c_1471_n 0.00502397f $X=3.9 $Y=0.72 $X2=0
+ $Y2=0
cc_590 N_A_558_445#_c_846_n N_VPWR_M1005_d 0.0135279f $X=4.155 $Y=2.37 $X2=0
+ $Y2=0
cc_591 N_A_558_445#_c_824_n N_VPWR_M1005_d 0.00485809f $X=4.24 $Y=2.285 $X2=0
+ $Y2=0
cc_592 N_A_558_445#_c_817_n N_VPWR_c_1245_n 0.00314961f $X=4.475 $Y=2.045 $X2=0
+ $Y2=0
cc_593 N_A_558_445#_c_817_n N_VPWR_c_1256_n 0.0051324f $X=4.475 $Y=2.045 $X2=0
+ $Y2=0
cc_594 N_A_558_445#_c_817_n N_VPWR_c_1237_n 0.00395238f $X=4.475 $Y=2.045 $X2=0
+ $Y2=0
cc_595 N_A_558_445#_c_818_n N_A_451_503#_c_1355_n 0.0449172f $X=2.97 $Y=2.285
+ $X2=0 $Y2=0
cc_596 N_A_558_445#_c_819_n N_A_451_503#_c_1355_n 0.0136278f $X=3.175 $Y=1.41
+ $X2=0 $Y2=0
cc_597 N_A_558_445#_c_820_n N_A_451_503#_c_1355_n 0.00752852f $X=3.215 $Y=0.815
+ $X2=0 $Y2=0
cc_598 N_A_558_445#_c_820_n N_A_451_503#_c_1356_n 0.0182668f $X=3.215 $Y=0.815
+ $X2=0 $Y2=0
cc_599 N_A_558_445#_c_818_n N_A_451_503#_c_1359_n 0.00592774f $X=2.97 $Y=2.285
+ $X2=0 $Y2=0
cc_600 N_A_558_445#_c_859_n N_A_451_503#_c_1359_n 0.0141909f $X=3.055 $Y=2.37
+ $X2=0 $Y2=0
cc_601 N_A_558_445#_c_820_n N_A_451_503#_c_1357_n 0.0124921f $X=3.215 $Y=0.815
+ $X2=0 $Y2=0
cc_602 N_A_558_445#_c_846_n A_702_445# 0.00568771f $X=4.155 $Y=2.37 $X2=-0.19
+ $Y2=-0.245
cc_603 N_A_558_445#_M1007_g N_VGND_c_1450_n 0.00781439f $X=4.425 $Y=0.655 $X2=0
+ $Y2=0
cc_604 N_A_558_445#_M1007_g N_VGND_c_1457_n 0.00493442f $X=4.425 $Y=0.655 $X2=0
+ $Y2=0
cc_605 N_A_558_445#_M1007_g N_VGND_c_1471_n 0.00473933f $X=4.425 $Y=0.655 $X2=0
+ $Y2=0
cc_606 N_A_1290_102#_c_914_n N_A_1000_424#_c_1067_n 0.00935642f $X=6.54 $Y=2.23
+ $X2=0 $Y2=0
cc_607 N_A_1290_102#_c_915_n N_A_1000_424#_c_1067_n 0.00976736f $X=6.54 $Y=2.32
+ $X2=0 $Y2=0
cc_608 N_A_1290_102#_c_925_n N_A_1000_424#_c_1067_n 0.0083953f $X=7.325 $Y=2.295
+ $X2=0 $Y2=0
cc_609 N_A_1290_102#_c_938_p N_A_1000_424#_c_1067_n 0.00573072f $X=7.925 $Y=2.27
+ $X2=0 $Y2=0
cc_610 N_A_1290_102#_c_917_n N_A_1000_424#_c_1068_n 0.022868f $X=8.085 $Y=1.765
+ $X2=0 $Y2=0
cc_611 N_A_1290_102#_c_910_n N_A_1000_424#_c_1068_n 0.00193983f $X=7.84 $Y=2.13
+ $X2=0 $Y2=0
cc_612 N_A_1290_102#_c_925_n N_A_1000_424#_c_1068_n 0.00949091f $X=7.325
+ $Y=2.295 $X2=0 $Y2=0
cc_613 N_A_1290_102#_c_938_p N_A_1000_424#_c_1068_n 0.0168326f $X=7.925 $Y=2.27
+ $X2=0 $Y2=0
cc_614 N_A_1290_102#_M1003_g N_A_1000_424#_M1021_g 0.0135422f $X=8.07 $Y=0.76
+ $X2=0 $Y2=0
cc_615 N_A_1290_102#_c_907_n N_A_1000_424#_M1021_g 0.00657776f $X=6.88 $Y=1.335
+ $X2=0 $Y2=0
cc_616 N_A_1290_102#_c_908_n N_A_1000_424#_M1021_g 0.00282836f $X=7.38 $Y=0.535
+ $X2=0 $Y2=0
cc_617 N_A_1290_102#_c_909_n N_A_1000_424#_M1021_g 0.0160542f $X=7.755 $Y=1.415
+ $X2=0 $Y2=0
cc_618 N_A_1290_102#_c_910_n N_A_1000_424#_M1021_g 0.00660122f $X=7.84 $Y=2.13
+ $X2=0 $Y2=0
cc_619 N_A_1290_102#_c_912_n N_A_1000_424#_M1021_g 0.00544313f $X=7.34 $Y=1.335
+ $X2=0 $Y2=0
cc_620 N_A_1290_102#_c_894_n N_A_1000_424#_c_1061_n 0.00177877f $X=6.525 $Y=1.17
+ $X2=0 $Y2=0
cc_621 N_A_1290_102#_c_901_n N_A_1000_424#_c_1061_n 0.00591361f $X=6.525
+ $Y=1.335 $X2=0 $Y2=0
cc_622 N_A_1290_102#_c_906_n N_A_1000_424#_c_1061_n 0.010473f $X=7.215 $Y=1.335
+ $X2=0 $Y2=0
cc_623 N_A_1290_102#_c_913_n N_A_1000_424#_c_1072_n 0.00251658f $X=6.54 $Y=1.83
+ $X2=0 $Y2=0
cc_624 N_A_1290_102#_c_914_n N_A_1000_424#_c_1072_n 0.00610334f $X=6.54 $Y=2.23
+ $X2=0 $Y2=0
cc_625 N_A_1290_102#_c_902_n N_A_1000_424#_c_1072_n 0.004253f $X=6.54 $Y=1.74
+ $X2=0 $Y2=0
cc_626 N_A_1290_102#_c_906_n N_A_1000_424#_c_1072_n 0.0398263f $X=7.215 $Y=1.335
+ $X2=0 $Y2=0
cc_627 N_A_1290_102#_c_907_n N_A_1000_424#_c_1072_n 0.0103313f $X=6.88 $Y=1.335
+ $X2=0 $Y2=0
cc_628 N_A_1290_102#_c_909_n N_A_1000_424#_c_1072_n 0.00864935f $X=7.755
+ $Y=1.415 $X2=0 $Y2=0
cc_629 N_A_1290_102#_c_910_n N_A_1000_424#_c_1072_n 0.0228576f $X=7.84 $Y=2.13
+ $X2=0 $Y2=0
cc_630 N_A_1290_102#_c_938_p N_A_1000_424#_c_1072_n 0.0274136f $X=7.925 $Y=2.27
+ $X2=0 $Y2=0
cc_631 N_A_1290_102#_c_912_n N_A_1000_424#_c_1072_n 0.0210596f $X=7.34 $Y=1.335
+ $X2=0 $Y2=0
cc_632 N_A_1290_102#_c_894_n N_A_1000_424#_c_1062_n 7.94759e-19 $X=6.525 $Y=1.17
+ $X2=0 $Y2=0
cc_633 N_A_1290_102#_c_913_n N_A_1000_424#_c_1065_n 0.00264146f $X=6.54 $Y=1.83
+ $X2=0 $Y2=0
cc_634 N_A_1290_102#_c_914_n N_A_1000_424#_c_1065_n 0.0070396f $X=6.54 $Y=2.23
+ $X2=0 $Y2=0
cc_635 N_A_1290_102#_c_902_n N_A_1000_424#_c_1065_n 0.0105968f $X=6.54 $Y=1.74
+ $X2=0 $Y2=0
cc_636 N_A_1290_102#_c_913_n N_A_1000_424#_c_1066_n 0.00875666f $X=6.54 $Y=1.83
+ $X2=0 $Y2=0
cc_637 N_A_1290_102#_c_896_n N_A_1000_424#_c_1066_n 0.0135422f $X=8.085 $Y=1.675
+ $X2=0 $Y2=0
cc_638 N_A_1290_102#_c_917_n N_A_1000_424#_c_1066_n 0.00776282f $X=8.085
+ $Y=1.765 $X2=0 $Y2=0
cc_639 N_A_1290_102#_c_902_n N_A_1000_424#_c_1066_n 0.00180154f $X=6.54 $Y=1.74
+ $X2=0 $Y2=0
cc_640 N_A_1290_102#_c_906_n N_A_1000_424#_c_1066_n 9.22454e-19 $X=7.215
+ $Y=1.335 $X2=0 $Y2=0
cc_641 N_A_1290_102#_c_907_n N_A_1000_424#_c_1066_n 0.00131525f $X=6.88 $Y=1.335
+ $X2=0 $Y2=0
cc_642 N_A_1290_102#_c_909_n N_A_1000_424#_c_1066_n 0.00148667f $X=7.755
+ $Y=1.415 $X2=0 $Y2=0
cc_643 N_A_1290_102#_c_910_n N_A_1000_424#_c_1066_n 0.00198529f $X=7.84 $Y=2.13
+ $X2=0 $Y2=0
cc_644 N_A_1290_102#_c_938_p N_A_1000_424#_c_1066_n 0.00570252f $X=7.925 $Y=2.27
+ $X2=0 $Y2=0
cc_645 N_A_1290_102#_c_912_n N_A_1000_424#_c_1066_n 0.00536859f $X=7.34 $Y=1.335
+ $X2=0 $Y2=0
cc_646 N_A_1290_102#_c_919_n N_A_1835_368#_c_1174_n 0.0152051f $X=9.545 $Y=1.765
+ $X2=0 $Y2=0
cc_647 N_A_1290_102#_M1027_g N_A_1835_368#_M1006_g 0.0144461f $X=9.56 $Y=0.79
+ $X2=0 $Y2=0
cc_648 N_A_1290_102#_M1013_g N_A_1835_368#_c_1170_n 0.00442778f $X=8.5 $Y=0.76
+ $X2=0 $Y2=0
cc_649 N_A_1290_102#_M1027_g N_A_1835_368#_c_1170_n 0.0204222f $X=9.56 $Y=0.79
+ $X2=0 $Y2=0
cc_650 N_A_1290_102#_c_899_n N_A_1835_368#_c_1176_n 0.00553801f $X=8.535
+ $Y=1.765 $X2=0 $Y2=0
cc_651 N_A_1290_102#_c_919_n N_A_1835_368#_c_1176_n 0.013769f $X=9.545 $Y=1.765
+ $X2=0 $Y2=0
cc_652 N_A_1290_102#_c_904_n N_A_1835_368#_c_1176_n 0.00608934f $X=9.455
+ $Y=1.485 $X2=0 $Y2=0
cc_653 N_A_1290_102#_c_905_n N_A_1835_368#_c_1176_n 0.00519786f $X=9.545
+ $Y=1.542 $X2=0 $Y2=0
cc_654 N_A_1290_102#_c_923_n N_A_1835_368#_c_1176_n 0.0120391f $X=8.685 $Y=2.325
+ $X2=0 $Y2=0
cc_655 N_A_1290_102#_c_911_n N_A_1835_368#_c_1176_n 0.0406944f $X=8.85 $Y=1.485
+ $X2=0 $Y2=0
cc_656 N_A_1290_102#_M1027_g N_A_1835_368#_c_1171_n 0.0062929f $X=9.56 $Y=0.79
+ $X2=0 $Y2=0
cc_657 N_A_1290_102#_c_905_n N_A_1835_368#_c_1171_n 0.0122689f $X=9.545 $Y=1.542
+ $X2=0 $Y2=0
cc_658 N_A_1290_102#_M1013_g N_A_1835_368#_c_1172_n 4.85699e-19 $X=8.5 $Y=0.76
+ $X2=0 $Y2=0
cc_659 N_A_1290_102#_M1027_g N_A_1835_368#_c_1172_n 4.11505e-19 $X=9.56 $Y=0.79
+ $X2=0 $Y2=0
cc_660 N_A_1290_102#_c_904_n N_A_1835_368#_c_1172_n 0.0154839f $X=9.455 $Y=1.485
+ $X2=0 $Y2=0
cc_661 N_A_1290_102#_c_905_n N_A_1835_368#_c_1172_n 0.00290339f $X=9.545
+ $Y=1.542 $X2=0 $Y2=0
cc_662 N_A_1290_102#_c_911_n N_A_1835_368#_c_1172_n 0.0201139f $X=8.85 $Y=1.485
+ $X2=0 $Y2=0
cc_663 N_A_1290_102#_M1027_g N_A_1835_368#_c_1173_n 0.0215705f $X=9.56 $Y=0.79
+ $X2=0 $Y2=0
cc_664 N_A_1290_102#_c_905_n N_A_1835_368#_c_1173_n 0.00509043f $X=9.545
+ $Y=1.542 $X2=0 $Y2=0
cc_665 N_A_1290_102#_c_910_n N_VPWR_M1020_s 0.00792577f $X=7.84 $Y=2.13 $X2=0
+ $Y2=0
cc_666 N_A_1290_102#_c_923_n N_VPWR_M1020_s 0.00131722f $X=8.685 $Y=2.325 $X2=0
+ $Y2=0
cc_667 N_A_1290_102#_c_938_p N_VPWR_M1020_s 0.00674665f $X=7.925 $Y=2.27 $X2=0
+ $Y2=0
cc_668 N_A_1290_102#_c_923_n N_VPWR_M1009_s 0.00396902f $X=8.685 $Y=2.325 $X2=0
+ $Y2=0
cc_669 N_A_1290_102#_c_911_n N_VPWR_M1009_s 0.00765323f $X=8.85 $Y=1.485 $X2=0
+ $Y2=0
cc_670 N_A_1290_102#_c_915_n N_VPWR_c_1239_n 0.0119957f $X=6.54 $Y=2.32 $X2=0
+ $Y2=0
cc_671 N_A_1290_102#_c_925_n N_VPWR_c_1239_n 0.0351127f $X=7.325 $Y=2.295 $X2=0
+ $Y2=0
cc_672 N_A_1290_102#_c_938_p N_VPWR_c_1239_n 0.0022175f $X=7.925 $Y=2.27 $X2=0
+ $Y2=0
cc_673 N_A_1290_102#_c_917_n N_VPWR_c_1240_n 0.0111353f $X=8.085 $Y=1.765 $X2=0
+ $Y2=0
cc_674 N_A_1290_102#_c_899_n N_VPWR_c_1240_n 0.0015077f $X=8.535 $Y=1.765 $X2=0
+ $Y2=0
cc_675 N_A_1290_102#_c_925_n N_VPWR_c_1240_n 0.0269155f $X=7.325 $Y=2.295 $X2=0
+ $Y2=0
cc_676 N_A_1290_102#_c_938_p N_VPWR_c_1240_n 0.0225477f $X=7.925 $Y=2.27 $X2=0
+ $Y2=0
cc_677 N_A_1290_102#_c_917_n N_VPWR_c_1241_n 0.0015077f $X=8.085 $Y=1.765 $X2=0
+ $Y2=0
cc_678 N_A_1290_102#_c_899_n N_VPWR_c_1241_n 0.0121397f $X=8.535 $Y=1.765 $X2=0
+ $Y2=0
cc_679 N_A_1290_102#_c_919_n N_VPWR_c_1241_n 0.0034303f $X=9.545 $Y=1.765 $X2=0
+ $Y2=0
cc_680 N_A_1290_102#_c_923_n N_VPWR_c_1241_n 0.0240652f $X=8.685 $Y=2.325 $X2=0
+ $Y2=0
cc_681 N_A_1290_102#_c_919_n N_VPWR_c_1242_n 0.0121299f $X=9.545 $Y=1.765 $X2=0
+ $Y2=0
cc_682 N_A_1290_102#_c_915_n N_VPWR_c_1245_n 0.00429349f $X=6.54 $Y=2.32 $X2=0
+ $Y2=0
cc_683 N_A_1290_102#_c_917_n N_VPWR_c_1247_n 0.00413917f $X=8.085 $Y=1.765 $X2=0
+ $Y2=0
cc_684 N_A_1290_102#_c_899_n N_VPWR_c_1247_n 0.00413917f $X=8.535 $Y=1.765 $X2=0
+ $Y2=0
cc_685 N_A_1290_102#_c_925_n N_VPWR_c_1250_n 0.0143676f $X=7.325 $Y=2.295 $X2=0
+ $Y2=0
cc_686 N_A_1290_102#_c_919_n N_VPWR_c_1251_n 0.00481995f $X=9.545 $Y=1.765 $X2=0
+ $Y2=0
cc_687 N_A_1290_102#_c_915_n N_VPWR_c_1237_n 0.00454161f $X=6.54 $Y=2.32 $X2=0
+ $Y2=0
cc_688 N_A_1290_102#_c_917_n N_VPWR_c_1237_n 0.00817726f $X=8.085 $Y=1.765 $X2=0
+ $Y2=0
cc_689 N_A_1290_102#_c_899_n N_VPWR_c_1237_n 0.00817726f $X=8.535 $Y=1.765 $X2=0
+ $Y2=0
cc_690 N_A_1290_102#_c_919_n N_VPWR_c_1237_n 0.00508379f $X=9.545 $Y=1.765 $X2=0
+ $Y2=0
cc_691 N_A_1290_102#_c_925_n N_VPWR_c_1237_n 0.0119073f $X=7.325 $Y=2.295 $X2=0
+ $Y2=0
cc_692 N_A_1290_102#_c_923_n N_Q_M1001_d 0.00907415f $X=8.685 $Y=2.325 $X2=0
+ $Y2=0
cc_693 N_A_1290_102#_M1003_g N_Q_c_1396_n 0.0054598f $X=8.07 $Y=0.76 $X2=0 $Y2=0
cc_694 N_A_1290_102#_c_896_n N_Q_c_1396_n 0.00181021f $X=8.085 $Y=1.675 $X2=0
+ $Y2=0
cc_695 N_A_1290_102#_c_897_n N_Q_c_1396_n 0.0116828f $X=8.425 $Y=1.395 $X2=0
+ $Y2=0
cc_696 N_A_1290_102#_M1013_g N_Q_c_1396_n 0.0185282f $X=8.5 $Y=0.76 $X2=0 $Y2=0
cc_697 N_A_1290_102#_c_899_n N_Q_c_1396_n 0.00518992f $X=8.535 $Y=1.765 $X2=0
+ $Y2=0
cc_698 N_A_1290_102#_c_903_n N_Q_c_1396_n 0.00194151f $X=8.085 $Y=1.395 $X2=0
+ $Y2=0
cc_699 N_A_1290_102#_c_909_n N_Q_c_1396_n 0.0117241f $X=7.755 $Y=1.415 $X2=0
+ $Y2=0
cc_700 N_A_1290_102#_c_910_n N_Q_c_1396_n 0.0351199f $X=7.84 $Y=2.13 $X2=0 $Y2=0
cc_701 N_A_1290_102#_c_911_n N_Q_c_1396_n 0.0132169f $X=8.85 $Y=1.485 $X2=0
+ $Y2=0
cc_702 N_A_1290_102#_c_896_n Q 0.00288356f $X=8.085 $Y=1.675 $X2=0 $Y2=0
cc_703 N_A_1290_102#_c_917_n Q 0.00684029f $X=8.085 $Y=1.765 $X2=0 $Y2=0
cc_704 N_A_1290_102#_c_899_n Q 0.0158485f $X=8.535 $Y=1.765 $X2=0 $Y2=0
cc_705 N_A_1290_102#_c_923_n Q 0.0201391f $X=8.685 $Y=2.325 $X2=0 $Y2=0
cc_706 N_A_1290_102#_c_911_n Q 0.0406991f $X=8.85 $Y=1.485 $X2=0 $Y2=0
cc_707 N_A_1290_102#_c_894_n N_VGND_c_1451_n 0.0120389f $X=6.525 $Y=1.17 $X2=0
+ $Y2=0
cc_708 N_A_1290_102#_c_906_n N_VGND_c_1451_n 0.0222475f $X=7.215 $Y=1.335 $X2=0
+ $Y2=0
cc_709 N_A_1290_102#_c_907_n N_VGND_c_1451_n 0.008037f $X=6.88 $Y=1.335 $X2=0
+ $Y2=0
cc_710 N_A_1290_102#_c_908_n N_VGND_c_1451_n 0.0415998f $X=7.38 $Y=0.535 $X2=0
+ $Y2=0
cc_711 N_A_1290_102#_M1003_g N_VGND_c_1452_n 0.00239046f $X=8.07 $Y=0.76 $X2=0
+ $Y2=0
cc_712 N_A_1290_102#_c_908_n N_VGND_c_1452_n 0.0294122f $X=7.38 $Y=0.535 $X2=0
+ $Y2=0
cc_713 N_A_1290_102#_c_909_n N_VGND_c_1452_n 0.0238954f $X=7.755 $Y=1.415 $X2=0
+ $Y2=0
cc_714 N_A_1290_102#_M1013_g N_VGND_c_1453_n 0.0184827f $X=8.5 $Y=0.76 $X2=0
+ $Y2=0
cc_715 N_A_1290_102#_M1027_g N_VGND_c_1453_n 0.00494501f $X=9.56 $Y=0.79 $X2=0
+ $Y2=0
cc_716 N_A_1290_102#_c_904_n N_VGND_c_1453_n 0.00301484f $X=9.455 $Y=1.485 $X2=0
+ $Y2=0
cc_717 N_A_1290_102#_c_911_n N_VGND_c_1453_n 0.0234476f $X=8.85 $Y=1.485 $X2=0
+ $Y2=0
cc_718 N_A_1290_102#_M1027_g N_VGND_c_1454_n 0.00884549f $X=9.56 $Y=0.79 $X2=0
+ $Y2=0
cc_719 N_A_1290_102#_c_894_n N_VGND_c_1457_n 0.00407505f $X=6.525 $Y=1.17 $X2=0
+ $Y2=0
cc_720 N_A_1290_102#_c_908_n N_VGND_c_1459_n 0.0102427f $X=7.38 $Y=0.535 $X2=0
+ $Y2=0
cc_721 N_A_1290_102#_M1003_g N_VGND_c_1461_n 0.00563421f $X=8.07 $Y=0.76 $X2=0
+ $Y2=0
cc_722 N_A_1290_102#_M1013_g N_VGND_c_1461_n 0.00537471f $X=8.5 $Y=0.76 $X2=0
+ $Y2=0
cc_723 N_A_1290_102#_M1027_g N_VGND_c_1465_n 0.00485498f $X=9.56 $Y=0.79 $X2=0
+ $Y2=0
cc_724 N_A_1290_102#_c_894_n N_VGND_c_1471_n 0.00465306f $X=6.525 $Y=1.17 $X2=0
+ $Y2=0
cc_725 N_A_1290_102#_M1003_g N_VGND_c_1471_n 0.00539454f $X=8.07 $Y=0.76 $X2=0
+ $Y2=0
cc_726 N_A_1290_102#_M1013_g N_VGND_c_1471_n 0.00539454f $X=8.5 $Y=0.76 $X2=0
+ $Y2=0
cc_727 N_A_1290_102#_M1027_g N_VGND_c_1471_n 0.00514438f $X=9.56 $Y=0.79 $X2=0
+ $Y2=0
cc_728 N_A_1290_102#_c_908_n N_VGND_c_1471_n 0.00904831f $X=7.38 $Y=0.535 $X2=0
+ $Y2=0
cc_729 N_A_1000_424#_c_1067_n N_VPWR_c_1239_n 0.0104868f $X=7.1 $Y=2.045 $X2=0
+ $Y2=0
cc_730 N_A_1000_424#_c_1072_n N_VPWR_c_1239_n 0.0149687f $X=7.42 $Y=1.795 $X2=0
+ $Y2=0
cc_731 N_A_1000_424#_c_1068_n N_VPWR_c_1240_n 0.00667613f $X=7.55 $Y=2.045 $X2=0
+ $Y2=0
cc_732 N_A_1000_424#_c_1067_n N_VPWR_c_1250_n 0.00445602f $X=7.1 $Y=2.045 $X2=0
+ $Y2=0
cc_733 N_A_1000_424#_c_1068_n N_VPWR_c_1250_n 0.00445602f $X=7.55 $Y=2.045 $X2=0
+ $Y2=0
cc_734 N_A_1000_424#_c_1067_n N_VPWR_c_1237_n 0.00863063f $X=7.1 $Y=2.045 $X2=0
+ $Y2=0
cc_735 N_A_1000_424#_c_1068_n N_VPWR_c_1237_n 0.00858495f $X=7.55 $Y=2.045 $X2=0
+ $Y2=0
cc_736 N_A_1000_424#_M1021_g N_Q_c_1396_n 3.10397e-19 $X=7.595 $Y=0.76 $X2=0
+ $Y2=0
cc_737 N_A_1000_424#_M1021_g N_VGND_c_1451_n 0.00284645f $X=7.595 $Y=0.76 $X2=0
+ $Y2=0
cc_738 N_A_1000_424#_c_1072_n N_VGND_c_1451_n 0.00182479f $X=7.42 $Y=1.795 $X2=0
+ $Y2=0
cc_739 N_A_1000_424#_M1021_g N_VGND_c_1452_n 0.0142125f $X=7.595 $Y=0.76 $X2=0
+ $Y2=0
cc_740 N_A_1000_424#_M1021_g N_VGND_c_1459_n 0.00468165f $X=7.595 $Y=0.76 $X2=0
+ $Y2=0
cc_741 N_A_1000_424#_M1021_g N_VGND_c_1471_n 0.00453141f $X=7.595 $Y=0.76 $X2=0
+ $Y2=0
cc_742 N_A_1835_368#_c_1176_n N_VPWR_c_1241_n 0.0146469f $X=9.32 $Y=1.985 $X2=0
+ $Y2=0
cc_743 N_A_1835_368#_c_1174_n N_VPWR_c_1242_n 0.00900997f $X=10.08 $Y=1.765
+ $X2=0 $Y2=0
cc_744 N_A_1835_368#_c_1176_n N_VPWR_c_1242_n 0.0670842f $X=9.32 $Y=1.985 $X2=0
+ $Y2=0
cc_745 N_A_1835_368#_c_1171_n N_VPWR_c_1242_n 0.0198836f $X=10.01 $Y=1.465 $X2=0
+ $Y2=0
cc_746 N_A_1835_368#_c_1173_n N_VPWR_c_1242_n 0.0021679f $X=10.53 $Y=1.532 $X2=0
+ $Y2=0
cc_747 N_A_1835_368#_c_1175_n N_VPWR_c_1244_n 0.00947143f $X=10.53 $Y=1.765
+ $X2=0 $Y2=0
cc_748 N_A_1835_368#_c_1176_n N_VPWR_c_1251_n 0.00739961f $X=9.32 $Y=1.985 $X2=0
+ $Y2=0
cc_749 N_A_1835_368#_c_1174_n N_VPWR_c_1252_n 0.00445602f $X=10.08 $Y=1.765
+ $X2=0 $Y2=0
cc_750 N_A_1835_368#_c_1175_n N_VPWR_c_1252_n 0.00405947f $X=10.53 $Y=1.765
+ $X2=0 $Y2=0
cc_751 N_A_1835_368#_c_1174_n N_VPWR_c_1237_n 0.00862391f $X=10.08 $Y=1.765
+ $X2=0 $Y2=0
cc_752 N_A_1835_368#_c_1175_n N_VPWR_c_1237_n 0.00732808f $X=10.53 $Y=1.765
+ $X2=0 $Y2=0
cc_753 N_A_1835_368#_c_1176_n N_VPWR_c_1237_n 0.00845774f $X=9.32 $Y=1.985 $X2=0
+ $Y2=0
cc_754 N_A_1835_368#_M1006_g N_Q_N_c_1417_n 0.00760237f $X=10.115 $Y=0.74 $X2=0
+ $Y2=0
cc_755 N_A_1835_368#_M1008_g N_Q_N_c_1417_n 0.0081896f $X=10.545 $Y=0.74 $X2=0
+ $Y2=0
cc_756 N_A_1835_368#_M1006_g N_Q_N_c_1418_n 0.00299567f $X=10.115 $Y=0.74 $X2=0
+ $Y2=0
cc_757 N_A_1835_368#_M1008_g N_Q_N_c_1418_n 0.00215589f $X=10.545 $Y=0.74 $X2=0
+ $Y2=0
cc_758 N_A_1835_368#_c_1173_n N_Q_N_c_1418_n 0.00244427f $X=10.53 $Y=1.532 $X2=0
+ $Y2=0
cc_759 N_A_1835_368#_c_1174_n Q_N 0.00233133f $X=10.08 $Y=1.765 $X2=0 $Y2=0
cc_760 N_A_1835_368#_c_1175_n Q_N 0.00248981f $X=10.53 $Y=1.765 $X2=0 $Y2=0
cc_761 N_A_1835_368#_c_1171_n Q_N 0.00179727f $X=10.01 $Y=1.465 $X2=0 $Y2=0
cc_762 N_A_1835_368#_c_1173_n Q_N 0.00819215f $X=10.53 $Y=1.532 $X2=0 $Y2=0
cc_763 N_A_1835_368#_c_1174_n Q_N 0.0110815f $X=10.08 $Y=1.765 $X2=0 $Y2=0
cc_764 N_A_1835_368#_c_1175_n Q_N 0.0134273f $X=10.53 $Y=1.765 $X2=0 $Y2=0
cc_765 N_A_1835_368#_M1006_g N_Q_N_c_1419_n 0.0025553f $X=10.115 $Y=0.74 $X2=0
+ $Y2=0
cc_766 N_A_1835_368#_c_1175_n N_Q_N_c_1419_n 0.00304427f $X=10.53 $Y=1.765 $X2=0
+ $Y2=0
cc_767 N_A_1835_368#_M1008_g N_Q_N_c_1419_n 0.00866774f $X=10.545 $Y=0.74 $X2=0
+ $Y2=0
cc_768 N_A_1835_368#_c_1171_n N_Q_N_c_1419_n 0.0249855f $X=10.01 $Y=1.465 $X2=0
+ $Y2=0
cc_769 N_A_1835_368#_c_1173_n N_Q_N_c_1419_n 0.0358413f $X=10.53 $Y=1.532 $X2=0
+ $Y2=0
cc_770 N_A_1835_368#_c_1170_n N_VGND_c_1453_n 0.0391375f $X=9.345 $Y=0.835 $X2=0
+ $Y2=0
cc_771 N_A_1835_368#_M1006_g N_VGND_c_1454_n 0.00500238f $X=10.115 $Y=0.74 $X2=0
+ $Y2=0
cc_772 N_A_1835_368#_c_1170_n N_VGND_c_1454_n 0.0411583f $X=9.345 $Y=0.835 $X2=0
+ $Y2=0
cc_773 N_A_1835_368#_c_1171_n N_VGND_c_1454_n 0.0213646f $X=10.01 $Y=1.465 $X2=0
+ $Y2=0
cc_774 N_A_1835_368#_c_1173_n N_VGND_c_1454_n 0.0032381f $X=10.53 $Y=1.532 $X2=0
+ $Y2=0
cc_775 N_A_1835_368#_M1008_g N_VGND_c_1456_n 0.00646793f $X=10.545 $Y=0.74 $X2=0
+ $Y2=0
cc_776 N_A_1835_368#_c_1170_n N_VGND_c_1465_n 0.0086032f $X=9.345 $Y=0.835 $X2=0
+ $Y2=0
cc_777 N_A_1835_368#_M1006_g N_VGND_c_1466_n 0.00434272f $X=10.115 $Y=0.74 $X2=0
+ $Y2=0
cc_778 N_A_1835_368#_M1008_g N_VGND_c_1466_n 0.00422942f $X=10.545 $Y=0.74 $X2=0
+ $Y2=0
cc_779 N_A_1835_368#_M1006_g N_VGND_c_1471_n 0.00825283f $X=10.115 $Y=0.74 $X2=0
+ $Y2=0
cc_780 N_A_1835_368#_M1008_g N_VGND_c_1471_n 0.00787255f $X=10.545 $Y=0.74 $X2=0
+ $Y2=0
cc_781 N_A_1835_368#_c_1170_n N_VGND_c_1471_n 0.00943069f $X=9.345 $Y=0.835
+ $X2=0 $Y2=0
cc_782 N_VPWR_c_1242_n Q_N 0.0783991f $X=9.855 $Y=1.985 $X2=0 $Y2=0
cc_783 N_VPWR_c_1244_n Q_N 0.0888504f $X=10.76 $Y=1.985 $X2=0 $Y2=0
cc_784 N_VPWR_c_1252_n Q_N 0.0160091f $X=10.675 $Y=3.33 $X2=0 $Y2=0
cc_785 N_VPWR_c_1237_n Q_N 0.0131029f $X=10.8 $Y=3.33 $X2=0 $Y2=0
cc_786 N_Q_c_1396_n N_VGND_c_1452_n 0.0310987f $X=8.285 $Y=0.535 $X2=0 $Y2=0
cc_787 N_Q_c_1396_n N_VGND_c_1453_n 0.0304975f $X=8.285 $Y=0.535 $X2=0 $Y2=0
cc_788 N_Q_c_1396_n N_VGND_c_1461_n 0.0124447f $X=8.285 $Y=0.535 $X2=0 $Y2=0
cc_789 N_Q_c_1396_n N_VGND_c_1471_n 0.0110345f $X=8.285 $Y=0.535 $X2=0 $Y2=0
cc_790 N_Q_N_c_1417_n N_VGND_c_1454_n 0.0295042f $X=10.33 $Y=0.515 $X2=0 $Y2=0
cc_791 N_Q_N_c_1417_n N_VGND_c_1456_n 0.0308798f $X=10.33 $Y=0.515 $X2=0 $Y2=0
cc_792 N_Q_N_c_1417_n N_VGND_c_1466_n 0.0149085f $X=10.33 $Y=0.515 $X2=0 $Y2=0
cc_793 N_Q_N_c_1417_n N_VGND_c_1471_n 0.0122037f $X=10.33 $Y=0.515 $X2=0 $Y2=0
