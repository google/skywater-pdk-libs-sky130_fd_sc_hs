* File: sky130_fd_sc_hs__sdfstp_4.spice
* Created: Thu Aug 27 21:09:43 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hs__sdfstp_4.pex.spice"
.subckt sky130_fd_sc_hs__sdfstp_4  VNB VPB SCE D SCD CLK SET_B VPWR Q VGND
* 
* VGND	VGND
* Q	Q
* VPWR	VPWR
* SET_B	SET_B
* CLK	CLK
* SCD	SCD
* D	D
* SCE	SCE
* VPB	VPB
* VNB	VNB
MM1043 N_VGND_M1043_d N_SCE_M1043_g N_A_27_74#_M1043_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.0819 AS=0.1197 PD=0.81 PS=1.41 NRD=19.992 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75002.1 A=0.063 P=1.14 MULT=1
MM1039 A_222_74# N_A_27_74#_M1039_g N_VGND_M1043_d VNB NLOWVT L=0.15 W=0.42
+ AD=0.0504 AS=0.0819 PD=0.66 PS=0.81 NRD=18.564 NRS=11.424 M=1 R=2.8 SA=75000.7
+ SB=75001.6 A=0.063 P=1.14 MULT=1
MM1040 N_A_288_464#_M1040_d N_D_M1040_g A_222_74# VNB NLOWVT L=0.15 W=0.42
+ AD=0.09135 AS=0.0504 PD=0.855 PS=0.66 NRD=21.42 NRS=18.564 M=1 R=2.8
+ SA=75001.1 SB=75001.2 A=0.063 P=1.14 MULT=1
MM1015 A_417_74# N_SCE_M1015_g N_A_288_464#_M1040_d VNB NLOWVT L=0.15 W=0.42
+ AD=0.0504 AS=0.09135 PD=0.66 PS=0.855 NRD=18.564 NRS=22.848 M=1 R=2.8
+ SA=75001.7 SB=75000.6 A=0.063 P=1.14 MULT=1
MM1016 N_VGND_M1016_d N_SCD_M1016_g A_417_74# VNB NLOWVT L=0.15 W=0.42 AD=0.1197
+ AS=0.0504 PD=1.41 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75002.1 SB=75000.2
+ A=0.063 P=1.14 MULT=1
MM1026 N_VGND_M1026_d N_CLK_M1026_g N_A_616_74#_M1026_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1295 AS=0.2109 PD=1.09 PS=2.05 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75000.7 A=0.111 P=1.78 MULT=1
MM1020 N_A_803_74#_M1020_d N_A_616_74#_M1020_g N_VGND_M1026_d VNB NLOWVT L=0.15
+ W=0.74 AD=0.2109 AS=0.1295 PD=2.05 PS=1.09 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.7 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1003 N_A_1017_81#_M1003_d N_A_616_74#_M1003_g N_A_288_464#_M1003_s VNB NLOWVT
+ L=0.15 W=0.42 AD=0.1113 AS=0.1765 PD=0.95 PS=1.73 NRD=71.424 NRS=24.276 M=1
+ R=2.8 SA=75000.3 SB=75001.4 A=0.063 P=1.14 MULT=1
MM1019 A_1153_81# N_A_803_74#_M1019_g N_A_1017_81#_M1003_d VNB NLOWVT L=0.15
+ W=0.42 AD=0.0504 AS=0.1113 PD=0.66 PS=0.95 NRD=18.564 NRS=0 M=1 R=2.8 SA=75001
+ SB=75000.7 A=0.063 P=1.14 MULT=1
MM1017 N_VGND_M1017_d N_A_1201_55#_M1017_g A_1153_81# VNB NLOWVT L=0.15 W=0.42
+ AD=0.2084 AS=0.0504 PD=1.95 PS=0.66 NRD=24.276 NRS=18.564 M=1 R=2.8 SA=75001.4
+ SB=75000.3 A=0.063 P=1.14 MULT=1
MM1023 A_1445_74# N_A_1017_81#_M1023_g N_A_1201_55#_M1023_s VNB NLOWVT L=0.15
+ W=0.42 AD=0.0504 AS=0.1197 PD=0.66 PS=1.41 NRD=18.564 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75001.8 A=0.063 P=1.14 MULT=1
MM1004 N_VGND_M1004_d N_SET_B_M1004_g A_1445_74# VNB NLOWVT L=0.15 W=0.42
+ AD=0.136302 AS=0.0504 PD=0.998491 PS=0.66 NRD=98.568 NRS=18.564 M=1 R=2.8
+ SA=75000.6 SB=75001.4 A=0.063 P=1.14 MULT=1
MM1013 N_VGND_M1004_d N_A_1017_81#_M1013_g N_A_1677_74#_M1013_s VNB NLOWVT
+ L=0.15 W=0.64 AD=0.207698 AS=0.0896 PD=1.52151 PS=0.92 NRD=0 NRS=0 M=1
+ R=4.26667 SA=75001 SB=75000.6 A=0.096 P=1.58 MULT=1
MM1049 N_VGND_M1049_d N_A_1017_81#_M1049_g N_A_1677_74#_M1013_s VNB NLOWVT
+ L=0.15 W=0.64 AD=0.1824 AS=0.0896 PD=1.85 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75001.4 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1012 N_A_1823_524#_M1012_d N_A_803_74#_M1012_g N_A_1677_74#_M1012_s VNB NLOWVT
+ L=0.15 W=0.64 AD=0.1824 AS=0.0896 PD=1.85 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75002 A=0.096 P=1.58 MULT=1
MM1034 N_A_1823_524#_M1034_d N_A_803_74#_M1034_g N_A_1677_74#_M1012_s VNB NLOWVT
+ L=0.15 W=0.64 AD=0.129147 AS=0.0896 PD=1.20755 PS=0.92 NRD=0 NRS=0 M=1
+ R=4.26667 SA=75000.6 SB=75001.6 A=0.096 P=1.58 MULT=1
MM1028 A_2149_74# N_A_616_74#_M1028_g N_A_1823_524#_M1034_d VNB NLOWVT L=0.15
+ W=0.42 AD=0.0504 AS=0.0847528 PD=0.66 PS=0.792453 NRD=18.564 NRS=23.568 M=1
+ R=2.8 SA=75001.1 SB=75001.8 A=0.063 P=1.14 MULT=1
MM1009 A_2227_74# N_A_2191_180#_M1009_g A_2149_74# VNB NLOWVT L=0.15 W=0.42
+ AD=0.0819 AS=0.0504 PD=0.81 PS=0.66 NRD=39.996 NRS=18.564 M=1 R=2.8 SA=75001.5
+ SB=75001.4 A=0.063 P=1.14 MULT=1
MM1036 N_VGND_M1036_d N_SET_B_M1036_g A_2227_74# VNB NLOWVT L=0.15 W=0.42
+ AD=0.1092 AS=0.0819 PD=0.94 PS=0.81 NRD=24.276 NRS=39.996 M=1 R=2.8 SA=75002.1
+ SB=75000.9 A=0.063 P=1.14 MULT=1
MM1037 N_A_2191_180#_M1037_d N_A_1823_524#_M1037_g N_VGND_M1036_d VNB NLOWVT
+ L=0.15 W=0.42 AD=0.1197 AS=0.1092 PD=1.41 PS=0.94 NRD=0 NRS=44.28 M=1 R=2.8
+ SA=75002.8 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1010 N_VGND_M1010_d N_A_1823_524#_M1010_g N_A_2580_74#_M1010_s VNB NLOWVT
+ L=0.15 W=0.74 AD=0.1295 AS=0.2109 PD=1.09 PS=2.05 NRD=11.34 NRS=0 M=1
+ R=4.93333 SA=75000.2 SB=75002.3 A=0.111 P=1.78 MULT=1
MM1001 N_Q_M1001_d N_A_2580_74#_M1001_g N_VGND_M1010_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.16095 AS=0.1295 PD=1.175 PS=1.09 NRD=13.776 NRS=0 M=1 R=4.93333
+ SA=75000.7 SB=75001.8 A=0.111 P=1.78 MULT=1
MM1014 N_Q_M1001_d N_A_2580_74#_M1014_g N_VGND_M1014_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.16095 AS=0.1295 PD=1.175 PS=1.09 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75001.3
+ SB=75001.2 A=0.111 P=1.78 MULT=1
MM1021 N_Q_M1021_d N_A_2580_74#_M1021_g N_VGND_M1014_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1295 PD=1.02 PS=1.09 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75001.8
+ SB=75000.7 A=0.111 P=1.78 MULT=1
MM1030 N_Q_M1021_d N_A_2580_74#_M1030_g N_VGND_M1030_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.25955 PD=1.02 PS=2.19 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75002.2
+ SB=75000.3 A=0.111 P=1.78 MULT=1
MM1046 N_VPWR_M1046_d N_SCE_M1046_g N_A_27_74#_M1046_s VPB PSHORT L=0.15 W=0.64
+ AD=0.096 AS=0.1824 PD=0.94 PS=1.85 NRD=3.0732 NRS=3.0732 M=1 R=4.26667
+ SA=75000.2 SB=75002.2 A=0.096 P=1.58 MULT=1
MM1047 A_204_464# N_SCE_M1047_g N_VPWR_M1046_d VPB PSHORT L=0.15 W=0.64
+ AD=0.0864 AS=0.096 PD=0.91 PS=0.94 NRD=24.625 NRS=3.0732 M=1 R=4.26667
+ SA=75000.7 SB=75001.8 A=0.096 P=1.58 MULT=1
MM1005 N_A_288_464#_M1005_d N_D_M1005_g A_204_464# VPB PSHORT L=0.15 W=0.64
+ AD=0.1536 AS=0.0864 PD=1.12 PS=0.91 NRD=30.7714 NRS=24.625 M=1 R=4.26667
+ SA=75001.1 SB=75001.4 A=0.096 P=1.58 MULT=1
MM1041 A_414_464# N_A_27_74#_M1041_g N_A_288_464#_M1005_d VPB PSHORT L=0.15
+ W=0.64 AD=0.0864 AS=0.1536 PD=0.91 PS=1.12 NRD=24.625 NRS=30.7714 M=1
+ R=4.26667 SA=75001.7 SB=75000.7 A=0.096 P=1.58 MULT=1
MM1000 N_VPWR_M1000_d N_SCD_M1000_g A_414_464# VPB PSHORT L=0.15 W=0.64
+ AD=0.2954 AS=0.0864 PD=2.4 PS=0.91 NRD=30.7714 NRS=24.625 M=1 R=4.26667
+ SA=75002.1 SB=75000.3 A=0.096 P=1.58 MULT=1
MM1006 N_VPWR_M1006_d N_CLK_M1006_g N_A_616_74#_M1006_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.3304 PD=1.42 PS=2.83 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1011 N_A_803_74#_M1011_d N_A_616_74#_M1011_g N_VPWR_M1006_d VPB PSHORT L=0.15
+ W=1.12 AD=0.3256 AS=0.168 PD=2.93 PS=1.42 NRD=10.5395 NRS=1.7533 M=1 R=7.46667
+ SA=75000.7 SB=75000.2 A=0.168 P=2.54 MULT=1
MM1029 N_A_1017_81#_M1029_d N_A_803_74#_M1029_g N_A_288_464#_M1029_s VPB PSHORT
+ L=0.15 W=0.42 AD=0.097475 AS=0.1239 PD=0.995 PS=1.43 NRD=4.6886 NRS=4.6886 M=1
+ R=2.8 SA=75000.2 SB=75002.1 A=0.063 P=1.14 MULT=1
MM1048 A_1140_495# N_A_616_74#_M1048_g N_A_1017_81#_M1029_d VPB PSHORT L=0.15
+ W=0.42 AD=0.091175 AS=0.097475 PD=0.965 PS=0.995 NRD=76.0223 NRS=46.886 M=1
+ R=2.8 SA=75000.5 SB=75001.8 A=0.063 P=1.14 MULT=1
MM1042 N_VPWR_M1042_d N_A_1201_55#_M1042_g A_1140_495# VPB PSHORT L=0.15 W=0.42
+ AD=0.156925 AS=0.091175 PD=1.24 PS=0.965 NRD=149.444 NRS=76.0223 M=1 R=2.8
+ SA=75000.8 SB=75002.6 A=0.063 P=1.14 MULT=1
MM1038 N_A_1201_55#_M1038_d N_A_1017_81#_M1038_g N_VPWR_M1042_d VPB PSHORT
+ L=0.15 W=0.42 AD=0.0693 AS=0.156925 PD=0.75 PS=1.24 NRD=18.7544 NRS=149.444
+ M=1 R=2.8 SA=75001.5 SB=75001.8 A=0.063 P=1.14 MULT=1
MM1035 N_VPWR_M1035_d N_SET_B_M1035_g N_A_1201_55#_M1038_d VPB PSHORT L=0.15
+ W=0.42 AD=0.1113 AS=0.0693 PD=0.913333 PS=0.75 NRD=112.566 NRS=4.6886 M=1
+ R=2.8 SA=75002 SB=75001.3 A=0.063 P=1.14 MULT=1
MM1002 N_A_1620_373#_M1002_d N_A_1017_81#_M1002_g N_VPWR_M1035_d VPB PSHORT
+ L=0.15 W=0.84 AD=0.126 AS=0.2226 PD=1.14 PS=1.82667 NRD=2.3443 NRS=2.3443 M=1
+ R=5.6 SA=75001.4 SB=75000.7 A=0.126 P=1.98 MULT=1
MM1008 N_A_1620_373#_M1002_d N_A_1017_81#_M1008_g N_VPWR_M1008_s VPB PSHORT
+ L=0.15 W=0.84 AD=0.126 AS=0.23175 PD=1.14 PS=2.27 NRD=2.3443 NRS=2.3443 M=1
+ R=5.6 SA=75001.9 SB=75000.2 A=0.126 P=1.98 MULT=1
MM1022 N_A_1620_373#_M1022_d N_A_616_74#_M1022_g N_A_1823_524#_M1022_s VPB
+ PSHORT L=0.15 W=0.84 AD=0.126 AS=0.2328 PD=1.14 PS=2.27 NRD=2.3443 NRS=2.3443
+ M=1 R=5.6 SA=75000.2 SB=75001.4 A=0.126 P=1.98 MULT=1
MM1024 N_A_1620_373#_M1022_d N_A_616_74#_M1024_g N_A_1823_524#_M1024_s VPB
+ PSHORT L=0.15 W=0.84 AD=0.126 AS=0.1736 PD=1.14 PS=1.59333 NRD=2.3443
+ NRS=14.0658 M=1 R=5.6 SA=75000.7 SB=75001 A=0.126 P=1.98 MULT=1
MM1045 A_2103_508# N_A_803_74#_M1045_g N_A_1823_524#_M1024_s VPB PSHORT L=0.15
+ W=0.42 AD=0.09975 AS=0.0868 PD=0.895 PS=0.796667 NRD=44.5417 NRS=7.0329 M=1
+ R=2.8 SA=75001.2 SB=75001.3 A=0.063 P=1.14 MULT=1
MM1025 N_VPWR_M1025_d N_A_2191_180#_M1025_g A_2103_508# VPB PSHORT L=0.15 W=0.42
+ AD=0.063 AS=0.09975 PD=0.72 PS=0.895 NRD=4.6886 NRS=46.886 M=1 R=2.8
+ SA=75001.8 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1031 N_A_1823_524#_M1031_d N_SET_B_M1031_g N_VPWR_M1025_d VPB PSHORT L=0.15
+ W=0.42 AD=0.1239 AS=0.063 PD=1.43 PS=0.72 NRD=4.6886 NRS=4.6886 M=1 R=2.8
+ SA=75002.2 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1018 N_VPWR_M1018_d N_A_1823_524#_M1018_g N_A_2191_180#_M1018_s VPB PSHORT
+ L=0.15 W=0.42 AD=0.0868 AS=0.1239 PD=0.796667 PS=1.43 NRD=30.4759 NRS=4.6886
+ M=1 R=2.8 SA=75000.2 SB=75003 A=0.063 P=1.14 MULT=1
MM1044 N_A_2580_74#_M1044_d N_A_1823_524#_M1044_g N_VPWR_M1018_d VPB PSHORT
+ L=0.15 W=0.84 AD=0.126 AS=0.1736 PD=1.14 PS=1.59333 NRD=2.3443 NRS=2.3443 M=1
+ R=5.6 SA=75000.5 SB=75002.5 A=0.126 P=1.98 MULT=1
MM1050 N_A_2580_74#_M1044_d N_A_1823_524#_M1050_g N_VPWR_M1050_s VPB PSHORT
+ L=0.15 W=0.84 AD=0.126 AS=0.1596 PD=1.14 PS=1.26429 NRD=2.3443 NRS=2.3443 M=1
+ R=5.6 SA=75000.9 SB=75002.1 A=0.126 P=1.98 MULT=1
MM1007 N_VPWR_M1050_s N_A_2580_74#_M1007_g N_Q_M1007_s VPB PSHORT L=0.15 W=1.12
+ AD=0.2128 AS=0.168 PD=1.68571 PS=1.42 NRD=11.426 NRS=1.7533 M=1 R=7.46667
+ SA=75001.1 SB=75001.6 A=0.168 P=2.54 MULT=1
MM1027 N_VPWR_M1027_d N_A_2580_74#_M1027_g N_Q_M1007_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.6 SB=75001.1 A=0.168 P=2.54 MULT=1
MM1032 N_VPWR_M1027_d N_A_2580_74#_M1032_g N_Q_M1032_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667 SA=75002
+ SB=75000.7 A=0.168 P=2.54 MULT=1
MM1033 N_VPWR_M1033_d N_A_2580_74#_M1033_g N_Q_M1032_s VPB PSHORT L=0.15 W=1.12
+ AD=0.3304 AS=0.168 PD=2.83 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75002.5 SB=75000.2 A=0.168 P=2.54 MULT=1
DX51_noxref VNB VPB NWDIODE A=30.1692 P=36.16
c_165 VNB 0 7.95967e-20 $X=0 $Y=0
*
.include "sky130_fd_sc_hs__sdfstp_4.pxi.spice"
*
.ends
*
*
