* NGSPICE file created from sky130_fd_sc_hs__and4b_1.ext - technology: sky130A

.subckt sky130_fd_sc_hs__and4b_1 A_N B C D VGND VNB VPB VPWR X
M1000 VGND D a_526_139# VNB nlowvt w=640000u l=150000u
+  ad=4.5645e+11p pd=3.97e+06u as=3.418e+11p ps=2.55e+06u
M1001 a_226_424# C VPWR VPB pshort w=840000u l=150000u
+  ad=6.132e+11p pd=4.82e+06u as=1.6114e+12p ps=9.26e+06u
M1002 VPWR D a_226_424# VPB pshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1003 a_448_139# B a_353_124# VNB nlowvt w=640000u l=150000u
+  ad=1.536e+11p pd=1.76e+06u as=2.21125e+11p ps=2.08e+06u
M1004 X a_226_424# VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=3.304e+11p pd=2.83e+06u as=0p ps=0u
M1005 VPWR B a_226_424# VPB pshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_353_124# a_27_74# a_226_424# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=1.824e+11p ps=1.85e+06u
M1007 X a_226_424# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1008 a_226_424# a_27_74# VPWR VPB pshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VPWR A_N a_27_74# VPB pshort w=840000u l=150000u
+  ad=0p pd=0u as=2.478e+11p ps=2.27e+06u
M1010 VGND A_N a_27_74# VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=1.5675e+11p ps=1.67e+06u
M1011 a_526_139# C a_448_139# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

