# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_hs__dfrbp_2
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_hs__dfrbp_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  13.92000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 0.810000 0.515000 1.570000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.543200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 12.975000 1.820000 13.305000 2.980000 ;
        RECT 13.060000 0.330000 13.390000 1.130000 ;
        RECT 13.135000 1.130000 13.305000 1.820000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.543200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 10.895000 1.320000 11.875000 1.410000 ;
        RECT 10.895000 1.410000 11.725000 1.540000 ;
        RECT 10.895000 1.540000 11.065000 2.900000 ;
        RECT 11.195000 0.350000 11.455000 0.770000 ;
        RECT 11.195000 0.770000 11.875000 1.320000 ;
    END
  END Q_N
  PIN RESET_B
    ANTENNAGATEAREA  0.378000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.025000 1.450000 1.315000 1.780000 ;
        RECT 2.385000 1.445000 2.755000 1.775000 ;
        RECT 9.540000 1.450000 9.955000 1.780000 ;
      LAYER mcon ;
        RECT 1.115000 1.580000 1.285000 1.750000 ;
        RECT 2.555000 1.580000 2.725000 1.750000 ;
        RECT 9.755000 1.580000 9.925000 1.750000 ;
      LAYER met1 ;
        RECT 1.055000 1.550000 1.345000 1.595000 ;
        RECT 1.055000 1.595000 9.985000 1.735000 ;
        RECT 1.055000 1.735000 1.345000 1.780000 ;
        RECT 2.495000 1.550000 2.785000 1.595000 ;
        RECT 2.495000 1.735000 2.785000 1.780000 ;
        RECT 9.695000 1.550000 9.985000 1.595000 ;
        RECT 9.695000 1.735000 9.985000 1.780000 ;
    END
  END RESET_B
  PIN CLK
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 6.705000 1.180000 7.045000 1.670000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT  0.000000 -0.085000 13.920000 0.085000 ;
        RECT  1.145000  0.085000  1.475000 0.810000 ;
        RECT  2.205000  0.085000  2.535000 0.780000 ;
        RECT  5.605000  0.085000  5.855000 0.490000 ;
        RECT  9.415000  0.085000  9.745000 0.720000 ;
        RECT 10.845000  0.085000 11.015000 1.100000 ;
        RECT 11.625000  0.085000 11.965000 0.600000 ;
        RECT 12.630000  0.085000 12.880000 1.130000 ;
        RECT 13.560000  0.085000 13.820000 1.130000 ;
      LAYER mcon ;
        RECT  0.155000 -0.085000  0.325000 0.085000 ;
        RECT  0.635000 -0.085000  0.805000 0.085000 ;
        RECT  1.115000 -0.085000  1.285000 0.085000 ;
        RECT  1.595000 -0.085000  1.765000 0.085000 ;
        RECT  2.075000 -0.085000  2.245000 0.085000 ;
        RECT  2.555000 -0.085000  2.725000 0.085000 ;
        RECT  3.035000 -0.085000  3.205000 0.085000 ;
        RECT  3.515000 -0.085000  3.685000 0.085000 ;
        RECT  3.995000 -0.085000  4.165000 0.085000 ;
        RECT  4.475000 -0.085000  4.645000 0.085000 ;
        RECT  4.955000 -0.085000  5.125000 0.085000 ;
        RECT  5.435000 -0.085000  5.605000 0.085000 ;
        RECT  5.915000 -0.085000  6.085000 0.085000 ;
        RECT  6.395000 -0.085000  6.565000 0.085000 ;
        RECT  6.875000 -0.085000  7.045000 0.085000 ;
        RECT  7.355000 -0.085000  7.525000 0.085000 ;
        RECT  7.835000 -0.085000  8.005000 0.085000 ;
        RECT  8.315000 -0.085000  8.485000 0.085000 ;
        RECT  8.795000 -0.085000  8.965000 0.085000 ;
        RECT  9.275000 -0.085000  9.445000 0.085000 ;
        RECT  9.755000 -0.085000  9.925000 0.085000 ;
        RECT 10.235000 -0.085000 10.405000 0.085000 ;
        RECT 10.715000 -0.085000 10.885000 0.085000 ;
        RECT 11.195000 -0.085000 11.365000 0.085000 ;
        RECT 11.675000 -0.085000 11.845000 0.085000 ;
        RECT 12.155000 -0.085000 12.325000 0.085000 ;
        RECT 12.635000 -0.085000 12.805000 0.085000 ;
        RECT 13.115000 -0.085000 13.285000 0.085000 ;
        RECT 13.595000 -0.085000 13.765000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.245000 13.920000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT  0.000000 3.245000 13.920000 3.415000 ;
        RECT  0.115000 1.940000  0.510000 2.965000 ;
        RECT  0.115000 2.965000  1.435000 3.245000 ;
        RECT  2.945000 2.625000  3.195000 3.245000 ;
        RECT  5.990000 2.765000  6.500000 3.245000 ;
        RECT  9.265000 2.290000  9.625000 3.245000 ;
        RECT 10.365000 2.290000 10.695000 3.245000 ;
        RECT 11.265000 1.740000 11.595000 3.245000 ;
        RECT 12.475000 1.820000 12.805000 3.245000 ;
        RECT 13.475000 1.820000 13.805000 3.245000 ;
      LAYER mcon ;
        RECT  0.155000 3.245000  0.325000 3.415000 ;
        RECT  0.635000 3.245000  0.805000 3.415000 ;
        RECT  1.115000 3.245000  1.285000 3.415000 ;
        RECT  1.595000 3.245000  1.765000 3.415000 ;
        RECT  2.075000 3.245000  2.245000 3.415000 ;
        RECT  2.555000 3.245000  2.725000 3.415000 ;
        RECT  3.035000 3.245000  3.205000 3.415000 ;
        RECT  3.515000 3.245000  3.685000 3.415000 ;
        RECT  3.995000 3.245000  4.165000 3.415000 ;
        RECT  4.475000 3.245000  4.645000 3.415000 ;
        RECT  4.955000 3.245000  5.125000 3.415000 ;
        RECT  5.435000 3.245000  5.605000 3.415000 ;
        RECT  5.915000 3.245000  6.085000 3.415000 ;
        RECT  6.395000 3.245000  6.565000 3.415000 ;
        RECT  6.875000 3.245000  7.045000 3.415000 ;
        RECT  7.355000 3.245000  7.525000 3.415000 ;
        RECT  7.835000 3.245000  8.005000 3.415000 ;
        RECT  8.315000 3.245000  8.485000 3.415000 ;
        RECT  8.795000 3.245000  8.965000 3.415000 ;
        RECT  9.275000 3.245000  9.445000 3.415000 ;
        RECT  9.755000 3.245000  9.925000 3.415000 ;
        RECT 10.235000 3.245000 10.405000 3.415000 ;
        RECT 10.715000 3.245000 10.885000 3.415000 ;
        RECT 11.195000 3.245000 11.365000 3.415000 ;
        RECT 11.675000 3.245000 11.845000 3.415000 ;
        RECT 12.155000 3.245000 12.325000 3.415000 ;
        RECT 12.635000 3.245000 12.805000 3.415000 ;
        RECT 13.115000 3.245000 13.285000 3.415000 ;
        RECT 13.595000 3.245000 13.765000 3.415000 ;
      LAYER met1 ;
        RECT 0.000000 3.085000 13.920000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.325000 0.390000  0.855000 0.640000 ;
      RECT  0.680000 1.950000  1.010000 2.625000 ;
      RECT  0.680000 2.625000  1.775000 2.795000 ;
      RECT  0.685000 0.640000  0.855000 1.950000 ;
      RECT  1.485000 1.015000  3.095000 1.185000 ;
      RECT  1.485000 1.185000  1.655000 2.285000 ;
      RECT  1.485000 2.285000  1.970000 2.455000 ;
      RECT  1.605000 2.795000  1.775000 2.905000 ;
      RECT  1.605000 2.905000  2.775000 3.075000 ;
      RECT  1.645000 0.350000  1.975000 1.015000 ;
      RECT  1.825000 1.470000  2.155000 1.945000 ;
      RECT  1.825000 1.945000  4.120000 2.115000 ;
      RECT  2.185000 2.115000  2.435000 2.735000 ;
      RECT  2.605000 2.285000  3.535000 2.455000 ;
      RECT  2.605000 2.455000  2.775000 2.905000 ;
      RECT  2.705000 0.255000  5.235000 0.425000 ;
      RECT  2.705000 0.425000  2.875000 1.015000 ;
      RECT  2.925000 1.185000  3.095000 1.555000 ;
      RECT  2.925000 1.555000  3.255000 1.775000 ;
      RECT  3.045000 0.595000  4.895000 0.765000 ;
      RECT  3.345000 0.935000  4.475000 1.105000 ;
      RECT  3.345000 1.105000  3.715000 1.385000 ;
      RECT  3.365000 2.455000  3.535000 2.905000 ;
      RECT  3.365000 2.905000  4.460000 3.075000 ;
      RECT  3.790000 2.115000  4.120000 2.735000 ;
      RECT  3.885000 1.275000  4.135000 1.610000 ;
      RECT  3.885000 1.610000  4.120000 1.945000 ;
      RECT  4.290000 2.410000  4.475000 2.485000 ;
      RECT  4.290000 2.485000  4.960000 2.815000 ;
      RECT  4.290000 2.815000  4.460000 2.905000 ;
      RECT  4.305000 1.105000  4.475000 2.410000 ;
      RECT  4.645000 0.765000  4.895000 1.600000 ;
      RECT  4.645000 1.910000  5.785000 2.240000 ;
      RECT  5.065000 0.425000  5.235000 0.660000 ;
      RECT  5.065000 0.660000  6.195000 0.830000 ;
      RECT  5.095000 1.000000  5.425000 1.840000 ;
      RECT  5.095000 1.840000  5.785000 1.910000 ;
      RECT  5.425000 2.240000  5.785000 2.425000 ;
      RECT  5.425000 2.425000  7.505000 2.595000 ;
      RECT  5.425000 2.595000  5.785000 2.980000 ;
      RECT  5.595000 1.340000  6.535000 1.670000 ;
      RECT  6.025000 0.255000  8.780000 0.425000 ;
      RECT  6.025000 0.425000  6.195000 0.660000 ;
      RECT  6.095000 1.670000  6.265000 1.840000 ;
      RECT  6.095000 1.840000  7.505000 2.170000 ;
      RECT  6.365000 0.635000  6.960000 0.965000 ;
      RECT  6.365000 0.965000  6.535000 1.340000 ;
      RECT  6.705000 2.170000  7.035000 2.255000 ;
      RECT  7.215000 0.425000  7.385000 1.355000 ;
      RECT  7.215000 1.355000  7.880000 1.525000 ;
      RECT  7.315000 2.595000  7.505000 2.905000 ;
      RECT  7.315000 2.905000  8.220000 3.075000 ;
      RECT  7.555000 0.595000  9.235000 0.765000 ;
      RECT  7.555000 0.765000  7.725000 1.185000 ;
      RECT  7.710000 1.525000  7.880000 2.735000 ;
      RECT  7.905000 0.935000 10.335000 1.105000 ;
      RECT  8.050000 1.275000  8.555000 1.605000 ;
      RECT  8.050000 1.605000  8.220000 2.905000 ;
      RECT  8.390000 1.925000  8.895000 2.095000 ;
      RECT  8.390000 2.095000  8.640000 2.385000 ;
      RECT  8.725000 1.105000 10.335000 1.265000 ;
      RECT  8.725000 1.265000  8.895000 1.925000 ;
      RECT  8.985000 0.350000  9.235000 0.595000 ;
      RECT  9.065000 1.455000  9.330000 1.950000 ;
      RECT  9.065000 1.950000 10.675000 2.120000 ;
      RECT  9.830000 2.120000 10.160000 2.385000 ;
      RECT 10.205000 0.350000 10.675000 0.765000 ;
      RECT 10.505000 0.765000 10.675000 1.950000 ;
      RECT 11.895000 1.740000 12.305000 2.780000 ;
      RECT 12.135000 0.350000 12.430000 1.300000 ;
      RECT 12.135000 1.300000 12.965000 1.630000 ;
      RECT 12.135000 1.630000 12.305000 1.740000 ;
  END
END sky130_fd_sc_hs__dfrbp_2
