* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hs__and4b_4 A_N B C D VGND VNB VPB VPWR X
M1000 a_664_125# C a_751_125# VNB nlowvt w=640000u l=150000u
+  ad=5.37125e+11p pd=5.53e+06u as=3.872e+11p ps=3.77e+06u
M1001 X a_199_294# VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=7.952e+11p pd=5.9e+06u as=2.8072e+12p ps=2.011e+07u
M1002 a_199_294# C VPWR VPB pshort w=1e+06u l=150000u
+  ad=1.76e+12p pd=1.152e+07u as=0p ps=0u
M1003 VPWR C a_199_294# VPB pshort w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_664_125# B a_1136_125# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=4.992e+11p ps=4.12e+06u
M1005 VPWR D a_199_294# VPB pshort w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VGND a_199_294# X VNB nlowvt w=740000u l=150000u
+  ad=1.25925e+12p pd=9.57e+06u as=4.144e+11p ps=4.08e+06u
M1007 VPWR a_199_294# X VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VGND D a_751_125# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VPWR a_199_294# X VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_199_294# D VPWR VPB pshort w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 X a_199_294# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VPWR A_N a_27_368# VPB pshort w=1e+06u l=150000u
+  ad=0p pd=0u as=2.95e+11p ps=2.59e+06u
M1013 VGND A_N a_27_368# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=1.824e+11p ps=1.85e+06u
M1014 a_1136_125# a_27_368# a_199_294# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=1.792e+11p ps=1.84e+06u
M1015 a_199_294# B VPWR VPB pshort w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_751_125# C a_664_125# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_1136_125# B a_664_125# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_751_125# D VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VPWR a_27_368# a_199_294# VPB pshort w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 VGND a_199_294# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_199_294# a_27_368# VPWR VPB pshort w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_199_294# a_27_368# a_1136_125# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 X a_199_294# VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 X a_199_294# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 VPWR B a_199_294# VPB pshort w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
