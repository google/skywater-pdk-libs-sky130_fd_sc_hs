* File: sky130_fd_sc_hs__o221a_1.spice
* Created: Thu Aug 27 20:59:10 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hs__o221a_1.pex.spice"
.subckt sky130_fd_sc_hs__o221a_1  VNB VPB A1 A2 B2 B1 C1 X VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* X	X
* C1	C1
* B1	B1
* B2	B2
* A2	A2
* A1	A1
* VPB	VPB
* VNB	VNB
MM1003 N_VGND_M1003_d N_A_83_264#_M1003_g N_X_M1003_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.166607 AS=0.2109 PD=1.25478 PS=2.05 NRD=11.34 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75001.2 A=0.111 P=1.78 MULT=1
MM1002 N_A_245_94#_M1002_d N_A1_M1002_g N_VGND_M1003_d VNB NLOWVT L=0.15 W=0.64
+ AD=0.112 AS=0.144093 PD=0.99 PS=1.08522 NRD=0 NRS=15.468 M=1 R=4.26667
+ SA=75000.8 SB=75000.7 A=0.096 P=1.58 MULT=1
MM1000 N_VGND_M1000_d N_A2_M1000_g N_A_245_94#_M1002_d VNB NLOWVT L=0.15 W=0.64
+ AD=0.1824 AS=0.112 PD=1.85 PS=0.99 NRD=0 NRS=13.116 M=1 R=4.26667 SA=75001.3
+ SB=75000.2 A=0.096 P=1.58 MULT=1
MM1001 N_A_245_94#_M1001_d N_B2_M1001_g N_A_456_74#_M1001_s VNB NLOWVT L=0.15
+ W=0.64 AD=0.0896 AS=0.2336 PD=0.92 PS=2.01 NRD=0 NRS=7.488 M=1 R=4.26667
+ SA=75000.3 SB=75001.3 A=0.096 P=1.58 MULT=1
MM1007 N_A_456_74#_M1007_d N_B1_M1007_g N_A_245_94#_M1001_d VNB NLOWVT L=0.15
+ W=0.64 AD=0.112 AS=0.0896 PD=0.99 PS=0.92 NRD=13.116 NRS=0 M=1 R=4.26667
+ SA=75000.7 SB=75000.9 A=0.096 P=1.58 MULT=1
MM1005 N_A_83_264#_M1005_d N_C1_M1005_g N_A_456_74#_M1007_d VNB NLOWVT L=0.15
+ W=0.64 AD=0.2944 AS=0.112 PD=2.2 PS=0.99 NRD=13.116 NRS=0 M=1 R=4.26667
+ SA=75001.2 SB=75000.4 A=0.096 P=1.58 MULT=1
MM1009 N_VPWR_M1009_d N_A_83_264#_M1009_g N_X_M1009_s VPB PSHORT L=0.15 W=1.12
+ AD=0.328498 AS=0.3304 PD=1.80679 PS=2.83 NRD=26.3783 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75003.2 A=0.168 P=2.54 MULT=1
MM1004 A_264_392# N_A1_M1004_g N_VPWR_M1009_d VPB PSHORT L=0.15 W=1 AD=0.135
+ AS=0.293302 PD=1.27 PS=1.61321 NRD=15.7403 NRS=31.5003 M=1 R=6.66667 SA=75001
+ SB=75002.8 A=0.15 P=2.3 MULT=1
MM1006 N_A_83_264#_M1006_d N_A2_M1006_g A_264_392# VPB PSHORT L=0.15 W=1 AD=0.21
+ AS=0.135 PD=1.42 PS=1.27 NRD=1.9503 NRS=15.7403 M=1 R=6.66667 SA=75001.4
+ SB=75002.4 A=0.15 P=2.3 MULT=1
MM1010 A_462_392# N_B2_M1010_g N_A_83_264#_M1006_d VPB PSHORT L=0.15 W=1 AD=0.21
+ AS=0.21 PD=1.42 PS=1.42 NRD=30.5153 NRS=25.5903 M=1 R=6.66667 SA=75001.9
+ SB=75001.8 A=0.15 P=2.3 MULT=1
MM1008 N_VPWR_M1008_d N_B1_M1008_g A_462_392# VPB PSHORT L=0.15 W=1 AD=0.43
+ AS=0.21 PD=1.86 PS=1.42 NRD=1.9503 NRS=30.5153 M=1 R=6.66667 SA=75002.5
+ SB=75001.2 A=0.15 P=2.3 MULT=1
MM1011 N_A_83_264#_M1011_d N_C1_M1011_g N_VPWR_M1008_d VPB PSHORT L=0.15 W=1
+ AD=0.295 AS=0.43 PD=2.59 PS=1.86 NRD=1.9503 NRS=11.8003 M=1 R=6.66667
+ SA=75003.5 SB=75000.2 A=0.15 P=2.3 MULT=1
DX12_noxref VNB VPB NWDIODE A=8.742 P=13.12
c_42 VNB 0 1.2498e-19 $X=0 $Y=0
*
.include "sky130_fd_sc_hs__o221a_1.pxi.spice"
*
.ends
*
*
