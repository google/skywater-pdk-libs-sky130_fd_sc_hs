* NGSPICE file created from sky130_fd_sc_hs__and3_2.ext - technology: sky130A

.subckt sky130_fd_sc_hs__and3_2 A B C VGND VNB VPB VPWR X
M1000 X a_41_384# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.368e+11p pd=2.12e+06u as=6.9565e+11p ps=5.12e+06u
M1001 a_41_384# B VPWR VPB pshort w=840000u l=150000u
+  ad=4.998e+11p pd=4.55e+06u as=1.3306e+12p ps=8.87e+06u
M1002 VPWR A a_41_384# VPB pshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1003 VPWR C a_41_384# VPB pshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 X a_41_384# VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=3.36e+11p pd=2.84e+06u as=0p ps=0u
M1005 VPWR a_41_384# X VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VGND C a_247_136# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=1.536e+11p ps=1.76e+06u
M1007 a_247_136# B a_133_136# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=2.688e+11p ps=2.12e+06u
M1008 a_133_136# A a_41_384# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=1.824e+11p ps=1.85e+06u
M1009 VGND a_41_384# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

