* File: sky130_fd_sc_hs__and4bb_4.pxi.spice
* Created: Thu Aug 27 20:34:05 2020
* 
x_PM_SKY130_FD_SC_HS__AND4BB_4%B_N N_B_N_M1020_g N_B_N_c_153_n N_B_N_M1010_g B_N
+ B_N PM_SKY130_FD_SC_HS__AND4BB_4%B_N
x_PM_SKY130_FD_SC_HS__AND4BB_4%A_N N_A_N_M1021_g N_A_N_c_180_n N_A_N_M1005_g A_N
+ PM_SKY130_FD_SC_HS__AND4BB_4%A_N
x_PM_SKY130_FD_SC_HS__AND4BB_4%A_200_74# N_A_200_74#_M1021_d N_A_200_74#_M1005_d
+ N_A_200_74#_c_208_n N_A_200_74#_c_214_n N_A_200_74#_M1004_g
+ N_A_200_74#_c_209_n N_A_200_74#_M1007_g N_A_200_74#_c_215_n
+ N_A_200_74#_M1024_g N_A_200_74#_M1027_g N_A_200_74#_c_216_n
+ N_A_200_74#_c_217_n N_A_200_74#_c_211_n N_A_200_74#_c_218_n
+ N_A_200_74#_c_212_n N_A_200_74#_c_213_n PM_SKY130_FD_SC_HS__AND4BB_4%A_200_74#
x_PM_SKY130_FD_SC_HS__AND4BB_4%A_27_74# N_A_27_74#_M1020_s N_A_27_74#_M1010_s
+ N_A_27_74#_M1000_g N_A_27_74#_c_301_n N_A_27_74#_c_318_n N_A_27_74#_M1012_g
+ N_A_27_74#_M1002_g N_A_27_74#_c_303_n N_A_27_74#_c_320_n N_A_27_74#_M1026_g
+ N_A_27_74#_c_304_n N_A_27_74#_c_305_n N_A_27_74#_c_306_n N_A_27_74#_c_321_n
+ N_A_27_74#_c_322_n N_A_27_74#_c_307_n N_A_27_74#_c_308_n N_A_27_74#_c_323_n
+ N_A_27_74#_c_309_n N_A_27_74#_c_310_n N_A_27_74#_c_311_n N_A_27_74#_c_312_n
+ N_A_27_74#_c_313_n N_A_27_74#_c_314_n N_A_27_74#_c_315_n N_A_27_74#_c_316_n
+ PM_SKY130_FD_SC_HS__AND4BB_4%A_27_74#
x_PM_SKY130_FD_SC_HS__AND4BB_4%C N_C_c_439_n N_C_M1019_g N_C_c_435_n N_C_M1001_g
+ N_C_c_440_n N_C_M1025_g N_C_c_436_n N_C_M1022_g C C N_C_c_438_n
+ PM_SKY130_FD_SC_HS__AND4BB_4%C
x_PM_SKY130_FD_SC_HS__AND4BB_4%D N_D_c_493_n N_D_M1003_g N_D_M1008_g N_D_M1023_g
+ N_D_c_494_n N_D_M1017_g D N_D_c_491_n N_D_c_492_n
+ PM_SKY130_FD_SC_HS__AND4BB_4%D
x_PM_SKY130_FD_SC_HS__AND4BB_4%A_472_388# N_A_472_388#_M1007_d
+ N_A_472_388#_M1004_d N_A_472_388#_M1012_d N_A_472_388#_M1019_d
+ N_A_472_388#_M1003_s N_A_472_388#_M1006_g N_A_472_388#_c_553_n
+ N_A_472_388#_M1011_g N_A_472_388#_M1009_g N_A_472_388#_c_554_n
+ N_A_472_388#_M1013_g N_A_472_388#_M1014_g N_A_472_388#_c_555_n
+ N_A_472_388#_M1015_g N_A_472_388#_c_556_n N_A_472_388#_M1016_g
+ N_A_472_388#_M1018_g N_A_472_388#_c_557_n N_A_472_388#_c_546_n
+ N_A_472_388#_c_547_n N_A_472_388#_c_559_n N_A_472_388#_c_548_n
+ N_A_472_388#_c_586_n N_A_472_388#_c_561_n N_A_472_388#_c_601_n
+ N_A_472_388#_c_609_n N_A_472_388#_c_562_n N_A_472_388#_c_549_n
+ N_A_472_388#_c_668_p N_A_472_388#_c_574_n N_A_472_388#_c_550_n
+ N_A_472_388#_c_551_n N_A_472_388#_c_604_n N_A_472_388#_c_563_n
+ N_A_472_388#_c_552_n PM_SKY130_FD_SC_HS__AND4BB_4%A_472_388#
x_PM_SKY130_FD_SC_HS__AND4BB_4%VPWR N_VPWR_M1010_d N_VPWR_M1004_s N_VPWR_M1024_s
+ N_VPWR_M1026_s N_VPWR_M1025_s N_VPWR_M1017_d N_VPWR_M1013_s N_VPWR_M1016_s
+ N_VPWR_c_719_n N_VPWR_c_720_n N_VPWR_c_721_n N_VPWR_c_722_n N_VPWR_c_723_n
+ N_VPWR_c_724_n N_VPWR_c_725_n N_VPWR_c_726_n N_VPWR_c_727_n N_VPWR_c_728_n
+ VPWR N_VPWR_c_729_n N_VPWR_c_730_n N_VPWR_c_731_n N_VPWR_c_732_n
+ N_VPWR_c_733_n N_VPWR_c_734_n N_VPWR_c_735_n N_VPWR_c_736_n N_VPWR_c_737_n
+ N_VPWR_c_738_n N_VPWR_c_739_n N_VPWR_c_740_n N_VPWR_c_741_n N_VPWR_c_718_n
+ PM_SKY130_FD_SC_HS__AND4BB_4%VPWR
x_PM_SKY130_FD_SC_HS__AND4BB_4%X N_X_M1006_s N_X_M1014_s N_X_M1011_d N_X_M1015_d
+ N_X_c_838_n N_X_c_845_n N_X_c_846_n N_X_c_839_n N_X_c_847_n N_X_c_840_n
+ N_X_c_841_n N_X_c_842_n X X X X N_X_c_844_n N_X_c_849_n
+ PM_SKY130_FD_SC_HS__AND4BB_4%X
x_PM_SKY130_FD_SC_HS__AND4BB_4%VGND N_VGND_M1020_d N_VGND_M1008_d N_VGND_M1023_d
+ N_VGND_M1009_d N_VGND_M1018_d N_VGND_c_902_n N_VGND_c_903_n N_VGND_c_904_n
+ N_VGND_c_905_n N_VGND_c_906_n N_VGND_c_907_n VGND N_VGND_c_908_n
+ N_VGND_c_909_n N_VGND_c_910_n N_VGND_c_911_n N_VGND_c_912_n N_VGND_c_913_n
+ N_VGND_c_914_n N_VGND_c_915_n N_VGND_c_916_n N_VGND_c_917_n
+ PM_SKY130_FD_SC_HS__AND4BB_4%VGND
x_PM_SKY130_FD_SC_HS__AND4BB_4%A_412_140# N_A_412_140#_M1007_s
+ N_A_412_140#_M1027_s N_A_412_140#_M1002_s N_A_412_140#_c_999_n
+ N_A_412_140#_c_1005_n N_A_412_140#_c_1009_n N_A_412_140#_c_1000_n
+ N_A_412_140#_c_1001_n N_A_412_140#_c_1002_n
+ PM_SKY130_FD_SC_HS__AND4BB_4%A_412_140#
x_PM_SKY130_FD_SC_HS__AND4BB_4%A_685_140# N_A_685_140#_M1000_d
+ N_A_685_140#_M1001_d N_A_685_140#_c_1045_n N_A_685_140#_c_1043_n
+ N_A_685_140#_c_1044_n PM_SKY130_FD_SC_HS__AND4BB_4%A_685_140#
x_PM_SKY130_FD_SC_HS__AND4BB_4%A_882_137# N_A_882_137#_M1001_s
+ N_A_882_137#_M1022_s N_A_882_137#_M1008_s N_A_882_137#_c_1078_n
+ N_A_882_137#_c_1072_n N_A_882_137#_c_1073_n N_A_882_137#_c_1074_n
+ N_A_882_137#_c_1075_n N_A_882_137#_c_1076_n
+ PM_SKY130_FD_SC_HS__AND4BB_4%A_882_137#
cc_1 VNB N_B_N_M1020_g 0.0436373f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.69
cc_2 VNB N_B_N_c_153_n 0.0204677f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.885
cc_3 VNB B_N 0.013883f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_4 VNB N_A_N_M1021_g 0.0402643f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.69
cc_5 VNB N_A_N_c_180_n 0.030448f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.885
cc_6 VNB A_N 0.00304223f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_7 VNB N_A_200_74#_c_208_n 0.0937102f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.46
cc_8 VNB N_A_200_74#_c_209_n 0.0162121f $X=-0.19 $Y=-0.245 $X2=0.41 $Y2=1.615
cc_9 VNB N_A_200_74#_M1027_g 0.0207625f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_200_74#_c_211_n 0.0148435f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_200_74#_c_212_n 0.0498318f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_200_74#_c_213_n 0.0701538f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_27_74#_M1000_g 0.00909884f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_27_74#_c_301_n 0.00938867f $X=-0.19 $Y=-0.245 $X2=0.41 $Y2=1.615
cc_15 VNB N_A_27_74#_M1002_g 0.0133109f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.615
cc_16 VNB N_A_27_74#_c_303_n 0.0099697f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_27_74#_c_304_n 0.00952495f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_27_74#_c_305_n 0.0143436f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_27_74#_c_306_n 0.0316008f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_27_74#_c_307_n 0.0193765f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_27_74#_c_308_n 0.00966715f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_27_74#_c_309_n 0.0127305f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_27_74#_c_310_n 0.00971798f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_27_74#_c_311_n 0.00538949f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_27_74#_c_312_n 0.00200673f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_27_74#_c_313_n 0.0201993f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_27_74#_c_314_n 0.0513599f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_27_74#_c_315_n 0.0134686f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_27_74#_c_316_n 0.0104154f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_C_c_435_n 0.0233589f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_C_c_436_n 0.0226967f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB C 0.00956749f $X=-0.19 $Y=-0.245 $X2=0.405 $Y2=1.615
cc_33 VNB N_C_c_438_n 0.0767249f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_D_M1008_g 0.0268913f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.46
cc_35 VNB N_D_M1023_g 0.0235388f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_D_c_491_n 0.0460295f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_D_c_492_n 0.00206152f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_472_388#_M1006_g 0.0234624f $X=-0.19 $Y=-0.245 $X2=0.405 $Y2=1.615
cc_39 VNB N_A_472_388#_M1009_g 0.0230515f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_472_388#_M1014_g 0.0236662f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_472_388#_M1018_g 0.0249674f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_472_388#_c_546_n 5.136e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_472_388#_c_547_n 0.00304539f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_472_388#_c_548_n 0.00464291f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_A_472_388#_c_549_n 0.00432957f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_A_472_388#_c_550_n 6.67308e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_472_388#_c_551_n 0.00259817f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_472_388#_c_552_n 0.103037f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_VPWR_c_718_n 0.382608f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_X_c_838_n 0.00240191f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.615
cc_51 VNB N_X_c_839_n 0.00230427f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_X_c_840_n 0.00203361f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_X_c_841_n 0.00139918f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_X_c_842_n 0.00300669f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB X 0.0253531f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_X_c_844_n 0.0158674f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_VGND_c_902_n 0.00396467f $X=-0.19 $Y=-0.245 $X2=0.405 $Y2=1.615
cc_58 VNB N_VGND_c_903_n 0.0238866f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_VGND_c_904_n 0.015906f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_VGND_c_905_n 0.00827016f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_VGND_c_906_n 0.0120978f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_VGND_c_907_n 0.0186272f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_VGND_c_908_n 0.0173909f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_VGND_c_909_n 0.1283f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_VGND_c_910_n 0.0177559f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_VGND_c_911_n 0.0186948f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_VGND_c_912_n 0.0188203f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_VGND_c_913_n 0.00604233f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_VGND_c_914_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_VGND_c_915_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_VGND_c_916_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_VGND_c_917_n 0.501346f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_A_412_140#_c_999_n 0.0022256f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_A_412_140#_c_1000_n 0.00269654f $X=-0.19 $Y=-0.245 $X2=0.405
+ $Y2=1.615
cc_75 VNB N_A_412_140#_c_1001_n 0.00229683f $X=-0.19 $Y=-0.245 $X2=0.72
+ $Y2=1.615
cc_76 VNB N_A_412_140#_c_1002_n 0.00574873f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_A_685_140#_c_1043_n 0.00377366f $X=-0.19 $Y=-0.245 $X2=0.405
+ $Y2=1.615
cc_78 VNB N_A_685_140#_c_1044_n 0.00951282f $X=-0.19 $Y=-0.245 $X2=0.24
+ $Y2=1.615
cc_79 VNB N_A_882_137#_c_1072_n 0.00720517f $X=-0.19 $Y=-0.245 $X2=0.405
+ $Y2=1.615
cc_80 VNB N_A_882_137#_c_1073_n 0.0195894f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_81 VNB N_A_882_137#_c_1074_n 0.00241395f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_82 VNB N_A_882_137#_c_1075_n 0.00490447f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_83 VNB N_A_882_137#_c_1076_n 0.00192273f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_84 VPB N_B_N_c_153_n 0.0451326f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.885
cc_85 VPB B_N 0.00939185f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_86 VPB N_A_N_c_180_n 0.0487003f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.885
cc_87 VPB A_N 0.00175299f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_88 VPB N_A_200_74#_c_214_n 0.0178531f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_89 VPB N_A_200_74#_c_215_n 0.0154174f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=1.615
cc_90 VPB N_A_200_74#_c_216_n 0.0274802f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_91 VPB N_A_200_74#_c_217_n 0.00172799f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_92 VPB N_A_200_74#_c_218_n 0.014605f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_93 VPB N_A_200_74#_c_213_n 0.0396065f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_94 VPB N_A_27_74#_c_301_n 6.75661e-19 $X=-0.19 $Y=1.66 $X2=0.41 $Y2=1.615
cc_95 VPB N_A_27_74#_c_318_n 0.0217f $X=-0.19 $Y=1.66 $X2=0.405 $Y2=1.615
cc_96 VPB N_A_27_74#_c_303_n 6.52919e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_97 VPB N_A_27_74#_c_320_n 0.0215602f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_98 VPB N_A_27_74#_c_321_n 0.00944206f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_99 VPB N_A_27_74#_c_322_n 0.035396f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_100 VPB N_A_27_74#_c_323_n 0.0128354f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_101 VPB N_A_27_74#_c_309_n 0.00660483f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_102 VPB N_C_c_439_n 0.0151591f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.45
cc_103 VPB N_C_c_440_n 0.0166678f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.46
cc_104 VPB C 0.00595846f $X=-0.19 $Y=1.66 $X2=0.405 $Y2=1.615
cc_105 VPB N_C_c_438_n 0.04197f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_106 VPB N_D_c_493_n 0.0194893f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.45
cc_107 VPB N_D_c_494_n 0.0159081f $X=-0.19 $Y=1.66 $X2=0.41 $Y2=1.615
cc_108 VPB N_D_c_491_n 0.0327994f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_109 VPB N_D_c_492_n 0.00482061f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_110 VPB N_A_472_388#_c_553_n 0.0167625f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_111 VPB N_A_472_388#_c_554_n 0.0148977f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_112 VPB N_A_472_388#_c_555_n 0.0148878f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_113 VPB N_A_472_388#_c_556_n 0.017194f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_114 VPB N_A_472_388#_c_557_n 0.00590147f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_115 VPB N_A_472_388#_c_547_n 0.00265889f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_116 VPB N_A_472_388#_c_559_n 0.00464832f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_117 VPB N_A_472_388#_c_548_n 0.00445015f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_118 VPB N_A_472_388#_c_561_n 0.0026622f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_119 VPB N_A_472_388#_c_562_n 0.00139165f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_120 VPB N_A_472_388#_c_563_n 9.411e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_121 VPB N_A_472_388#_c_552_n 0.0258073f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_122 VPB N_VPWR_c_719_n 0.00970163f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_123 VPB N_VPWR_c_720_n 0.0106927f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_124 VPB N_VPWR_c_721_n 0.0097085f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_125 VPB N_VPWR_c_722_n 0.012167f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_126 VPB N_VPWR_c_723_n 0.00810709f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_127 VPB N_VPWR_c_724_n 0.00261791f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_128 VPB N_VPWR_c_725_n 0.0120106f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_129 VPB N_VPWR_c_726_n 0.0341743f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_130 VPB N_VPWR_c_727_n 0.0274458f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_131 VPB N_VPWR_c_728_n 0.00638169f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_132 VPB N_VPWR_c_729_n 0.0191515f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_133 VPB N_VPWR_c_730_n 0.0209682f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_134 VPB N_VPWR_c_731_n 0.0187421f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_135 VPB N_VPWR_c_732_n 0.0204795f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_136 VPB N_VPWR_c_733_n 0.0164465f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_137 VPB N_VPWR_c_734_n 0.0177589f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_138 VPB N_VPWR_c_735_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_139 VPB N_VPWR_c_736_n 0.00628551f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_140 VPB N_VPWR_c_737_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_141 VPB N_VPWR_c_738_n 0.0187933f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_142 VPB N_VPWR_c_739_n 0.0397224f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_143 VPB N_VPWR_c_740_n 0.00614127f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_144 VPB N_VPWR_c_741_n 0.00601644f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_145 VPB N_VPWR_c_718_n 0.136431f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_146 VPB N_X_c_845_n 0.00118063f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_147 VPB N_X_c_846_n 0.00180921f $X=-0.19 $Y=1.66 $X2=0.72 $Y2=1.615
cc_148 VPB N_X_c_847_n 0.00511057f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_149 VPB X 0.00790433f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_150 VPB N_X_c_849_n 0.0137315f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_151 N_B_N_M1020_g N_A_N_M1021_g 0.0205581f $X=0.495 $Y=0.69 $X2=0 $Y2=0
cc_152 N_B_N_c_153_n N_A_N_c_180_n 0.0535272f $X=0.505 $Y=1.885 $X2=0 $Y2=0
cc_153 B_N N_A_N_c_180_n 0.00334101f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_154 N_B_N_c_153_n A_N 2.20145e-19 $X=0.505 $Y=1.885 $X2=0 $Y2=0
cc_155 B_N A_N 0.0277562f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_156 N_B_N_M1020_g N_A_27_74#_c_306_n 0.00446473f $X=0.495 $Y=0.69 $X2=0 $Y2=0
cc_157 N_B_N_c_153_n N_A_27_74#_c_321_n 0.00515127f $X=0.505 $Y=1.885 $X2=0
+ $Y2=0
cc_158 B_N N_A_27_74#_c_321_n 0.0273936f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_159 N_B_N_c_153_n N_A_27_74#_c_322_n 0.0104164f $X=0.505 $Y=1.885 $X2=0 $Y2=0
cc_160 N_B_N_M1020_g N_A_27_74#_c_307_n 0.0156808f $X=0.495 $Y=0.69 $X2=0 $Y2=0
cc_161 N_B_N_c_153_n N_A_27_74#_c_307_n 0.00123751f $X=0.505 $Y=1.885 $X2=0
+ $Y2=0
cc_162 B_N N_A_27_74#_c_307_n 0.0358185f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_163 N_B_N_c_153_n N_A_27_74#_c_308_n 0.00291196f $X=0.505 $Y=1.885 $X2=0
+ $Y2=0
cc_164 B_N N_A_27_74#_c_308_n 0.0207147f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_165 N_B_N_c_153_n N_A_27_74#_c_323_n 0.0124102f $X=0.505 $Y=1.885 $X2=0 $Y2=0
cc_166 B_N N_A_27_74#_c_323_n 0.0298654f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_167 N_B_N_c_153_n N_VPWR_c_719_n 0.00737447f $X=0.505 $Y=1.885 $X2=0 $Y2=0
cc_168 N_B_N_c_153_n N_VPWR_c_729_n 0.00445602f $X=0.505 $Y=1.885 $X2=0 $Y2=0
cc_169 N_B_N_c_153_n N_VPWR_c_718_n 0.00861319f $X=0.505 $Y=1.885 $X2=0 $Y2=0
cc_170 N_B_N_M1020_g N_VGND_c_902_n 0.0134383f $X=0.495 $Y=0.69 $X2=0 $Y2=0
cc_171 N_B_N_M1020_g N_VGND_c_908_n 0.00383152f $X=0.495 $Y=0.69 $X2=0 $Y2=0
cc_172 N_B_N_M1020_g N_VGND_c_917_n 0.00761198f $X=0.495 $Y=0.69 $X2=0 $Y2=0
cc_173 N_A_N_M1021_g N_A_200_74#_c_211_n 0.00908685f $X=0.925 $Y=0.69 $X2=0
+ $Y2=0
cc_174 N_A_N_c_180_n N_A_200_74#_c_218_n 0.00733793f $X=1.055 $Y=1.885 $X2=0
+ $Y2=0
cc_175 N_A_N_M1021_g N_A_200_74#_c_212_n 0.00993237f $X=0.925 $Y=0.69 $X2=0
+ $Y2=0
cc_176 N_A_N_c_180_n N_A_200_74#_c_213_n 0.00470986f $X=1.055 $Y=1.885 $X2=0
+ $Y2=0
cc_177 N_A_N_c_180_n N_A_27_74#_c_322_n 9.09193e-19 $X=1.055 $Y=1.885 $X2=0
+ $Y2=0
cc_178 N_A_N_M1021_g N_A_27_74#_c_307_n 0.0182295f $X=0.925 $Y=0.69 $X2=0 $Y2=0
cc_179 N_A_N_c_180_n N_A_27_74#_c_307_n 0.00248776f $X=1.055 $Y=1.885 $X2=0
+ $Y2=0
cc_180 A_N N_A_27_74#_c_307_n 0.0247729f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_181 N_A_N_c_180_n N_A_27_74#_c_323_n 0.0232501f $X=1.055 $Y=1.885 $X2=0 $Y2=0
cc_182 A_N N_A_27_74#_c_323_n 0.0243089f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_183 N_A_N_M1021_g N_A_27_74#_c_309_n 0.00408509f $X=0.925 $Y=0.69 $X2=0 $Y2=0
cc_184 N_A_N_c_180_n N_A_27_74#_c_309_n 0.00820947f $X=1.055 $Y=1.885 $X2=0
+ $Y2=0
cc_185 A_N N_A_27_74#_c_309_n 0.0248017f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_186 N_A_N_c_180_n N_VPWR_c_719_n 0.00737447f $X=1.055 $Y=1.885 $X2=0 $Y2=0
cc_187 N_A_N_c_180_n N_VPWR_c_727_n 0.00445602f $X=1.055 $Y=1.885 $X2=0 $Y2=0
cc_188 N_A_N_c_180_n N_VPWR_c_718_n 0.00862626f $X=1.055 $Y=1.885 $X2=0 $Y2=0
cc_189 N_A_N_M1021_g N_VGND_c_902_n 0.00978617f $X=0.925 $Y=0.69 $X2=0 $Y2=0
cc_190 N_A_N_M1021_g N_VGND_c_909_n 0.00383152f $X=0.925 $Y=0.69 $X2=0 $Y2=0
cc_191 N_A_N_M1021_g N_VGND_c_917_n 0.00758333f $X=0.925 $Y=0.69 $X2=0 $Y2=0
cc_192 N_A_200_74#_M1027_g N_A_27_74#_M1000_g 0.014235f $X=2.92 $Y=1.02 $X2=0
+ $Y2=0
cc_193 N_A_200_74#_c_213_n N_A_27_74#_c_301_n 0.0131467f $X=2.905 $Y=1.642 $X2=0
+ $Y2=0
cc_194 N_A_200_74#_c_215_n N_A_27_74#_c_318_n 0.00695262f $X=2.905 $Y=1.865
+ $X2=0 $Y2=0
cc_195 N_A_200_74#_c_213_n N_A_27_74#_c_304_n 0.014235f $X=2.905 $Y=1.642 $X2=0
+ $Y2=0
cc_196 N_A_200_74#_c_211_n N_A_27_74#_c_307_n 0.0398614f $X=1.525 $Y=0.42 $X2=0
+ $Y2=0
cc_197 N_A_200_74#_c_212_n N_A_27_74#_c_307_n 5.61223e-19 $X=1.525 $Y=0.255
+ $X2=0 $Y2=0
cc_198 N_A_200_74#_M1005_d N_A_27_74#_c_323_n 0.00354207f $X=1.13 $Y=1.96 $X2=0
+ $Y2=0
cc_199 N_A_200_74#_c_214_n N_A_27_74#_c_323_n 7.60268e-19 $X=2.285 $Y=1.865
+ $X2=0 $Y2=0
cc_200 N_A_200_74#_c_216_n N_A_27_74#_c_323_n 0.0187077f $X=1.93 $Y=2.375 $X2=0
+ $Y2=0
cc_201 N_A_200_74#_c_217_n N_A_27_74#_c_323_n 0.0110431f $X=2.095 $Y=1.615 $X2=0
+ $Y2=0
cc_202 N_A_200_74#_c_218_n N_A_27_74#_c_323_n 0.0221794f $X=1.28 $Y=2.455 $X2=0
+ $Y2=0
cc_203 N_A_200_74#_c_214_n N_A_27_74#_c_309_n 3.21515e-19 $X=2.285 $Y=1.865
+ $X2=0 $Y2=0
cc_204 N_A_200_74#_c_217_n N_A_27_74#_c_309_n 0.028437f $X=2.095 $Y=1.615 $X2=0
+ $Y2=0
cc_205 N_A_200_74#_c_213_n N_A_27_74#_c_309_n 0.00491283f $X=2.905 $Y=1.642
+ $X2=0 $Y2=0
cc_206 N_A_200_74#_c_209_n N_A_27_74#_c_310_n 3.77207e-19 $X=2.49 $Y=1.42 $X2=0
+ $Y2=0
cc_207 N_A_200_74#_c_211_n N_A_27_74#_c_310_n 0.00123224f $X=1.525 $Y=0.42 $X2=0
+ $Y2=0
cc_208 N_A_200_74#_c_209_n N_A_27_74#_c_311_n 0.00462012f $X=2.49 $Y=1.42 $X2=0
+ $Y2=0
cc_209 N_A_200_74#_c_211_n N_A_27_74#_c_311_n 0.00878228f $X=1.525 $Y=0.42 $X2=0
+ $Y2=0
cc_210 N_A_200_74#_c_208_n N_A_27_74#_c_312_n 0.0070675f $X=2.845 $Y=0.255 $X2=0
+ $Y2=0
cc_211 N_A_200_74#_c_211_n N_A_27_74#_c_312_n 0.0289714f $X=1.525 $Y=0.42 $X2=0
+ $Y2=0
cc_212 N_A_200_74#_c_212_n N_A_27_74#_c_312_n 0.00201826f $X=1.525 $Y=0.255
+ $X2=0 $Y2=0
cc_213 N_A_200_74#_c_208_n N_A_27_74#_c_313_n 0.0267676f $X=2.845 $Y=0.255 $X2=0
+ $Y2=0
cc_214 N_A_200_74#_c_209_n N_A_27_74#_c_313_n 0.00435912f $X=2.49 $Y=1.42 $X2=0
+ $Y2=0
cc_215 N_A_200_74#_M1027_g N_A_27_74#_c_313_n 0.0124453f $X=2.92 $Y=1.02 $X2=0
+ $Y2=0
cc_216 N_A_200_74#_c_208_n N_A_27_74#_c_314_n 0.014235f $X=2.845 $Y=0.255 $X2=0
+ $Y2=0
cc_217 N_A_200_74#_c_211_n N_A_27_74#_c_315_n 0.00515294f $X=1.525 $Y=0.42 $X2=0
+ $Y2=0
cc_218 N_A_200_74#_c_212_n N_A_27_74#_c_315_n 8.53526e-19 $X=1.525 $Y=0.255
+ $X2=0 $Y2=0
cc_219 N_A_200_74#_c_208_n N_A_27_74#_c_316_n 0.00186169f $X=2.845 $Y=0.255
+ $X2=0 $Y2=0
cc_220 N_A_200_74#_c_209_n N_A_27_74#_c_316_n 7.68543e-19 $X=2.49 $Y=1.42 $X2=0
+ $Y2=0
cc_221 N_A_200_74#_c_217_n N_A_27_74#_c_316_n 0.00336014f $X=2.095 $Y=1.615
+ $X2=0 $Y2=0
cc_222 N_A_200_74#_c_211_n N_A_27_74#_c_316_n 0.0145405f $X=1.525 $Y=0.42 $X2=0
+ $Y2=0
cc_223 N_A_200_74#_c_213_n N_A_27_74#_c_316_n 0.0018084f $X=2.905 $Y=1.642 $X2=0
+ $Y2=0
cc_224 N_A_200_74#_c_214_n N_A_472_388#_c_557_n 0.0138478f $X=2.285 $Y=1.865
+ $X2=0 $Y2=0
cc_225 N_A_200_74#_c_215_n N_A_472_388#_c_557_n 0.0123168f $X=2.905 $Y=1.865
+ $X2=0 $Y2=0
cc_226 N_A_200_74#_c_216_n N_A_472_388#_c_557_n 0.0140085f $X=1.93 $Y=2.375
+ $X2=0 $Y2=0
cc_227 N_A_200_74#_c_217_n N_A_472_388#_c_557_n 0.0408423f $X=2.095 $Y=1.615
+ $X2=0 $Y2=0
cc_228 N_A_200_74#_c_213_n N_A_472_388#_c_557_n 0.0123033f $X=2.905 $Y=1.642
+ $X2=0 $Y2=0
cc_229 N_A_200_74#_c_209_n N_A_472_388#_c_546_n 0.00328475f $X=2.49 $Y=1.42
+ $X2=0 $Y2=0
cc_230 N_A_200_74#_c_217_n N_A_472_388#_c_546_n 0.00705931f $X=2.095 $Y=1.615
+ $X2=0 $Y2=0
cc_231 N_A_200_74#_c_213_n N_A_472_388#_c_546_n 0.0125008f $X=2.905 $Y=1.642
+ $X2=0 $Y2=0
cc_232 N_A_200_74#_c_213_n N_A_472_388#_c_547_n 0.0198065f $X=2.905 $Y=1.642
+ $X2=0 $Y2=0
cc_233 N_A_200_74#_c_217_n N_A_472_388#_c_574_n 0.0135702f $X=2.095 $Y=1.615
+ $X2=0 $Y2=0
cc_234 N_A_200_74#_c_213_n N_A_472_388#_c_574_n 0.0111343f $X=2.905 $Y=1.642
+ $X2=0 $Y2=0
cc_235 N_A_200_74#_c_209_n N_A_472_388#_c_550_n 0.00617901f $X=2.49 $Y=1.42
+ $X2=0 $Y2=0
cc_236 N_A_200_74#_M1027_g N_A_472_388#_c_550_n 0.0034006f $X=2.92 $Y=1.02 $X2=0
+ $Y2=0
cc_237 N_A_200_74#_c_216_n N_VPWR_M1004_s 0.00565233f $X=1.93 $Y=2.375 $X2=0
+ $Y2=0
cc_238 N_A_200_74#_c_217_n N_VPWR_M1004_s 0.0110629f $X=2.095 $Y=1.615 $X2=0
+ $Y2=0
cc_239 N_A_200_74#_c_218_n N_VPWR_c_719_n 0.0202646f $X=1.28 $Y=2.455 $X2=0
+ $Y2=0
cc_240 N_A_200_74#_c_214_n N_VPWR_c_720_n 0.00884708f $X=2.285 $Y=1.865 $X2=0
+ $Y2=0
cc_241 N_A_200_74#_c_215_n N_VPWR_c_720_n 5.48865e-19 $X=2.905 $Y=1.865 $X2=0
+ $Y2=0
cc_242 N_A_200_74#_c_216_n N_VPWR_c_720_n 0.0243403f $X=1.93 $Y=2.375 $X2=0
+ $Y2=0
cc_243 N_A_200_74#_c_218_n N_VPWR_c_720_n 0.0144807f $X=1.28 $Y=2.455 $X2=0
+ $Y2=0
cc_244 N_A_200_74#_c_214_n N_VPWR_c_721_n 6.92486e-19 $X=2.285 $Y=1.865 $X2=0
+ $Y2=0
cc_245 N_A_200_74#_c_215_n N_VPWR_c_721_n 0.0150347f $X=2.905 $Y=1.865 $X2=0
+ $Y2=0
cc_246 N_A_200_74#_c_213_n N_VPWR_c_721_n 4.60757e-19 $X=2.905 $Y=1.642 $X2=0
+ $Y2=0
cc_247 N_A_200_74#_c_218_n N_VPWR_c_727_n 0.0146094f $X=1.28 $Y=2.455 $X2=0
+ $Y2=0
cc_248 N_A_200_74#_c_214_n N_VPWR_c_730_n 0.00505726f $X=2.285 $Y=1.865 $X2=0
+ $Y2=0
cc_249 N_A_200_74#_c_215_n N_VPWR_c_730_n 0.00505726f $X=2.905 $Y=1.865 $X2=0
+ $Y2=0
cc_250 N_A_200_74#_c_214_n N_VPWR_c_718_n 0.00489105f $X=2.285 $Y=1.865 $X2=0
+ $Y2=0
cc_251 N_A_200_74#_c_215_n N_VPWR_c_718_n 0.00489105f $X=2.905 $Y=1.865 $X2=0
+ $Y2=0
cc_252 N_A_200_74#_c_218_n N_VPWR_c_718_n 0.0120527f $X=1.28 $Y=2.455 $X2=0
+ $Y2=0
cc_253 N_A_200_74#_c_211_n N_VGND_c_902_n 0.0310975f $X=1.525 $Y=0.42 $X2=0
+ $Y2=0
cc_254 N_A_200_74#_c_212_n N_VGND_c_902_n 0.00139083f $X=1.525 $Y=0.255 $X2=0
+ $Y2=0
cc_255 N_A_200_74#_c_211_n N_VGND_c_909_n 0.044552f $X=1.525 $Y=0.42 $X2=0 $Y2=0
cc_256 N_A_200_74#_c_212_n N_VGND_c_909_n 0.0311384f $X=1.525 $Y=0.255 $X2=0
+ $Y2=0
cc_257 N_A_200_74#_c_208_n N_VGND_c_917_n 0.0339501f $X=2.845 $Y=0.255 $X2=0
+ $Y2=0
cc_258 N_A_200_74#_c_211_n N_VGND_c_917_n 0.0234606f $X=1.525 $Y=0.42 $X2=0
+ $Y2=0
cc_259 N_A_200_74#_c_212_n N_VGND_c_917_n 0.00902231f $X=1.525 $Y=0.255 $X2=0
+ $Y2=0
cc_260 N_A_200_74#_c_217_n N_A_412_140#_c_999_n 0.0173419f $X=2.095 $Y=1.615
+ $X2=0 $Y2=0
cc_261 N_A_200_74#_c_213_n N_A_412_140#_c_999_n 0.00993336f $X=2.905 $Y=1.642
+ $X2=0 $Y2=0
cc_262 N_A_200_74#_c_208_n N_A_412_140#_c_1005_n 7.84051e-19 $X=2.845 $Y=0.255
+ $X2=0 $Y2=0
cc_263 N_A_200_74#_c_209_n N_A_412_140#_c_1005_n 0.0135536f $X=2.49 $Y=1.42
+ $X2=0 $Y2=0
cc_264 N_A_200_74#_M1027_g N_A_412_140#_c_1005_n 0.0112505f $X=2.92 $Y=1.02
+ $X2=0 $Y2=0
cc_265 N_A_200_74#_c_213_n N_A_412_140#_c_1005_n 3.49041e-19 $X=2.905 $Y=1.642
+ $X2=0 $Y2=0
cc_266 N_A_200_74#_c_208_n N_A_412_140#_c_1009_n 7.05474e-19 $X=2.845 $Y=0.255
+ $X2=0 $Y2=0
cc_267 N_A_200_74#_M1027_g N_A_412_140#_c_1001_n 0.00134031f $X=2.92 $Y=1.02
+ $X2=0 $Y2=0
cc_268 N_A_27_74#_c_320_n N_C_c_439_n 0.0250405f $X=3.855 $Y=1.865 $X2=-0.19
+ $Y2=-0.245
cc_269 N_A_27_74#_c_305_n N_C_c_438_n 0.0150711f $X=3.825 $Y=1.565 $X2=0 $Y2=0
cc_270 N_A_27_74#_c_304_n N_A_472_388#_c_546_n 5.80494e-19 $X=3.37 $Y=1.565
+ $X2=0 $Y2=0
cc_271 N_A_27_74#_c_301_n N_A_472_388#_c_547_n 0.0147184f $X=3.375 $Y=1.775
+ $X2=0 $Y2=0
cc_272 N_A_27_74#_c_304_n N_A_472_388#_c_547_n 3.10926e-19 $X=3.37 $Y=1.565
+ $X2=0 $Y2=0
cc_273 N_A_27_74#_c_301_n N_A_472_388#_c_559_n 0.00292666f $X=3.375 $Y=1.775
+ $X2=0 $Y2=0
cc_274 N_A_27_74#_c_318_n N_A_472_388#_c_559_n 0.00225222f $X=3.375 $Y=1.865
+ $X2=0 $Y2=0
cc_275 N_A_27_74#_c_303_n N_A_472_388#_c_559_n 2.35363e-19 $X=3.855 $Y=1.775
+ $X2=0 $Y2=0
cc_276 N_A_27_74#_c_320_n N_A_472_388#_c_559_n 0.0156499f $X=3.855 $Y=1.865
+ $X2=0 $Y2=0
cc_277 N_A_27_74#_c_303_n N_A_472_388#_c_548_n 0.0132561f $X=3.855 $Y=1.775
+ $X2=0 $Y2=0
cc_278 N_A_27_74#_c_303_n N_A_472_388#_c_586_n 3.06637e-19 $X=3.855 $Y=1.775
+ $X2=0 $Y2=0
cc_279 N_A_27_74#_c_320_n N_A_472_388#_c_586_n 2.1541e-19 $X=3.855 $Y=1.865
+ $X2=0 $Y2=0
cc_280 N_A_27_74#_c_301_n N_A_472_388#_c_551_n 0.00215191f $X=3.375 $Y=1.775
+ $X2=0 $Y2=0
cc_281 N_A_27_74#_c_303_n N_A_472_388#_c_551_n 0.00306703f $X=3.855 $Y=1.775
+ $X2=0 $Y2=0
cc_282 N_A_27_74#_c_305_n N_A_472_388#_c_551_n 0.00193587f $X=3.825 $Y=1.565
+ $X2=0 $Y2=0
cc_283 N_A_27_74#_c_323_n N_VPWR_M1010_d 0.00339226f $X=1.505 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_284 N_A_27_74#_c_322_n N_VPWR_c_719_n 0.0266809f $X=0.28 $Y=2.815 $X2=0 $Y2=0
cc_285 N_A_27_74#_c_323_n N_VPWR_c_719_n 0.0232685f $X=1.505 $Y=2.035 $X2=0
+ $Y2=0
cc_286 N_A_27_74#_c_318_n N_VPWR_c_721_n 0.00231206f $X=3.375 $Y=1.865 $X2=0
+ $Y2=0
cc_287 N_A_27_74#_c_320_n N_VPWR_c_722_n 0.00800839f $X=3.855 $Y=1.865 $X2=0
+ $Y2=0
cc_288 N_A_27_74#_c_322_n N_VPWR_c_729_n 0.0145938f $X=0.28 $Y=2.815 $X2=0 $Y2=0
cc_289 N_A_27_74#_c_318_n N_VPWR_c_731_n 0.00563421f $X=3.375 $Y=1.865 $X2=0
+ $Y2=0
cc_290 N_A_27_74#_c_320_n N_VPWR_c_731_n 0.00548284f $X=3.855 $Y=1.865 $X2=0
+ $Y2=0
cc_291 N_A_27_74#_c_318_n N_VPWR_c_718_n 0.00539454f $X=3.375 $Y=1.865 $X2=0
+ $Y2=0
cc_292 N_A_27_74#_c_320_n N_VPWR_c_718_n 0.00539454f $X=3.855 $Y=1.865 $X2=0
+ $Y2=0
cc_293 N_A_27_74#_c_322_n N_VPWR_c_718_n 0.0120466f $X=0.28 $Y=2.815 $X2=0 $Y2=0
cc_294 N_A_27_74#_c_306_n N_VGND_c_902_n 0.0218743f $X=0.28 $Y=0.515 $X2=0 $Y2=0
cc_295 N_A_27_74#_c_307_n N_VGND_c_902_n 0.0216087f $X=1.505 $Y=1.195 $X2=0
+ $Y2=0
cc_296 N_A_27_74#_c_306_n N_VGND_c_908_n 0.011066f $X=0.28 $Y=0.515 $X2=0 $Y2=0
cc_297 N_A_27_74#_c_312_n N_VGND_c_909_n 0.0113382f $X=2.03 $Y=0.42 $X2=0 $Y2=0
cc_298 N_A_27_74#_c_313_n N_VGND_c_909_n 0.102136f $X=3.44 $Y=0.42 $X2=0 $Y2=0
cc_299 N_A_27_74#_c_314_n N_VGND_c_909_n 0.0140245f $X=3.44 $Y=0.42 $X2=0 $Y2=0
cc_300 N_A_27_74#_c_316_n N_VGND_c_909_n 0.00231009f $X=1.945 $Y=0.84 $X2=0
+ $Y2=0
cc_301 N_A_27_74#_c_306_n N_VGND_c_917_n 0.00915947f $X=0.28 $Y=0.515 $X2=0
+ $Y2=0
cc_302 N_A_27_74#_c_312_n N_VGND_c_917_n 0.00578038f $X=2.03 $Y=0.42 $X2=0 $Y2=0
cc_303 N_A_27_74#_c_313_n N_VGND_c_917_n 0.0554621f $X=3.44 $Y=0.42 $X2=0 $Y2=0
cc_304 N_A_27_74#_c_314_n N_VGND_c_917_n 0.0195747f $X=3.44 $Y=0.42 $X2=0 $Y2=0
cc_305 N_A_27_74#_c_316_n N_VGND_c_917_n 0.00356149f $X=1.945 $Y=0.84 $X2=0
+ $Y2=0
cc_306 N_A_27_74#_c_310_n N_A_412_140#_c_999_n 0.00892866f $X=1.785 $Y=1.11
+ $X2=0 $Y2=0
cc_307 N_A_27_74#_c_313_n N_A_412_140#_c_999_n 0.00576807f $X=3.44 $Y=0.42 $X2=0
+ $Y2=0
cc_308 N_A_27_74#_c_315_n N_A_412_140#_c_999_n 0.0149304f $X=1.785 $Y=1.195
+ $X2=0 $Y2=0
cc_309 N_A_27_74#_c_313_n N_A_412_140#_c_1005_n 0.0562084f $X=3.44 $Y=0.42 $X2=0
+ $Y2=0
cc_310 N_A_27_74#_c_313_n N_A_412_140#_c_1009_n 0.0130786f $X=3.44 $Y=0.42 $X2=0
+ $Y2=0
cc_311 N_A_27_74#_c_316_n N_A_412_140#_c_1009_n 0.014633f $X=1.945 $Y=0.84 $X2=0
+ $Y2=0
cc_312 N_A_27_74#_M1000_g N_A_412_140#_c_1000_n 0.00951876f $X=3.35 $Y=1.02
+ $X2=0 $Y2=0
cc_313 N_A_27_74#_M1002_g N_A_412_140#_c_1000_n 0.00665652f $X=3.78 $Y=1.02
+ $X2=0 $Y2=0
cc_314 N_A_27_74#_c_304_n N_A_412_140#_c_1000_n 0.00355459f $X=3.37 $Y=1.565
+ $X2=0 $Y2=0
cc_315 N_A_27_74#_c_305_n N_A_412_140#_c_1000_n 0.00164533f $X=3.825 $Y=1.565
+ $X2=0 $Y2=0
cc_316 N_A_27_74#_c_313_n N_A_412_140#_c_1000_n 0.00373775f $X=3.44 $Y=0.42
+ $X2=0 $Y2=0
cc_317 N_A_27_74#_M1000_g N_A_412_140#_c_1002_n 5.2012e-19 $X=3.35 $Y=1.02 $X2=0
+ $Y2=0
cc_318 N_A_27_74#_M1002_g N_A_412_140#_c_1002_n 0.00555614f $X=3.78 $Y=1.02
+ $X2=0 $Y2=0
cc_319 N_A_27_74#_c_305_n N_A_412_140#_c_1002_n 0.00376118f $X=3.825 $Y=1.565
+ $X2=0 $Y2=0
cc_320 N_A_27_74#_M1000_g N_A_685_140#_c_1045_n 0.00403483f $X=3.35 $Y=1.02
+ $X2=0 $Y2=0
cc_321 N_A_27_74#_c_313_n N_A_685_140#_c_1045_n 0.0131248f $X=3.44 $Y=0.42 $X2=0
+ $Y2=0
cc_322 N_A_27_74#_c_314_n N_A_685_140#_c_1045_n 0.00230414f $X=3.44 $Y=0.42
+ $X2=0 $Y2=0
cc_323 N_A_27_74#_M1002_g N_A_685_140#_c_1044_n 0.0125952f $X=3.78 $Y=1.02 $X2=0
+ $Y2=0
cc_324 N_A_27_74#_c_305_n N_A_685_140#_c_1044_n 2.4493e-19 $X=3.825 $Y=1.565
+ $X2=0 $Y2=0
cc_325 N_A_27_74#_M1002_g N_A_882_137#_c_1075_n 4.96257e-19 $X=3.78 $Y=1.02
+ $X2=0 $Y2=0
cc_326 C N_D_c_491_n 0.0050985f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_327 N_C_c_438_n N_D_c_491_n 0.00607386f $X=5.27 $Y=1.657 $X2=0 $Y2=0
cc_328 C N_D_c_492_n 0.021868f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_329 N_C_c_439_n N_A_472_388#_c_559_n 4.21309e-19 $X=4.405 $Y=1.865 $X2=0
+ $Y2=0
cc_330 N_C_c_438_n N_A_472_388#_c_559_n 3.21583e-19 $X=5.27 $Y=1.657 $X2=0 $Y2=0
cc_331 C N_A_472_388#_c_548_n 0.0143906f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_332 N_C_c_438_n N_A_472_388#_c_548_n 0.0253852f $X=5.27 $Y=1.657 $X2=0 $Y2=0
cc_333 N_C_c_439_n N_A_472_388#_c_586_n 0.00241623f $X=4.405 $Y=1.865 $X2=0
+ $Y2=0
cc_334 N_C_c_440_n N_A_472_388#_c_586_n 0.0044102f $X=4.855 $Y=1.865 $X2=0 $Y2=0
cc_335 C N_A_472_388#_c_586_n 0.00107985f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_336 N_C_c_438_n N_A_472_388#_c_586_n 0.0158057f $X=5.27 $Y=1.657 $X2=0 $Y2=0
cc_337 N_C_c_439_n N_A_472_388#_c_561_n 0.0084427f $X=4.405 $Y=1.865 $X2=0 $Y2=0
cc_338 N_C_c_440_n N_A_472_388#_c_561_n 0.0142651f $X=4.855 $Y=1.865 $X2=0 $Y2=0
cc_339 N_C_c_440_n N_A_472_388#_c_601_n 0.0159635f $X=4.855 $Y=1.865 $X2=0 $Y2=0
cc_340 C N_A_472_388#_c_601_n 0.08529f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_341 N_C_c_438_n N_A_472_388#_c_601_n 0.01656f $X=5.27 $Y=1.657 $X2=0 $Y2=0
cc_342 N_C_c_439_n N_A_472_388#_c_604_n 0.00163992f $X=4.405 $Y=1.865 $X2=0
+ $Y2=0
cc_343 N_C_c_440_n N_A_472_388#_c_604_n 2.24111e-19 $X=4.855 $Y=1.865 $X2=0
+ $Y2=0
cc_344 N_C_c_439_n N_VPWR_c_722_n 0.00800711f $X=4.405 $Y=1.865 $X2=0 $Y2=0
cc_345 N_C_c_439_n N_VPWR_c_738_n 0.00548284f $X=4.405 $Y=1.865 $X2=0 $Y2=0
cc_346 N_C_c_440_n N_VPWR_c_738_n 0.00548284f $X=4.855 $Y=1.865 $X2=0 $Y2=0
cc_347 N_C_c_440_n N_VPWR_c_739_n 0.0167538f $X=4.855 $Y=1.865 $X2=0 $Y2=0
cc_348 N_C_c_439_n N_VPWR_c_718_n 0.00539454f $X=4.405 $Y=1.865 $X2=0 $Y2=0
cc_349 N_C_c_440_n N_VPWR_c_718_n 0.00539454f $X=4.855 $Y=1.865 $X2=0 $Y2=0
cc_350 N_C_c_436_n N_VGND_c_903_n 0.00297788f $X=5.27 $Y=1.45 $X2=0 $Y2=0
cc_351 N_C_c_435_n N_VGND_c_909_n 0.0030414f $X=4.84 $Y=1.45 $X2=0 $Y2=0
cc_352 N_C_c_436_n N_VGND_c_909_n 0.00370946f $X=5.27 $Y=1.45 $X2=0 $Y2=0
cc_353 N_C_c_435_n N_VGND_c_917_n 0.00453162f $X=4.84 $Y=1.45 $X2=0 $Y2=0
cc_354 N_C_c_436_n N_VGND_c_917_n 0.00453162f $X=5.27 $Y=1.45 $X2=0 $Y2=0
cc_355 N_C_c_435_n N_A_412_140#_c_1002_n 0.00266806f $X=4.84 $Y=1.45 $X2=0 $Y2=0
cc_356 N_C_c_435_n N_A_685_140#_c_1043_n 0.00584349f $X=4.84 $Y=1.45 $X2=0 $Y2=0
cc_357 N_C_c_436_n N_A_685_140#_c_1043_n 0.00397428f $X=5.27 $Y=1.45 $X2=0 $Y2=0
cc_358 N_C_c_435_n N_A_685_140#_c_1044_n 0.0103912f $X=4.84 $Y=1.45 $X2=0 $Y2=0
cc_359 N_C_c_438_n N_A_685_140#_c_1044_n 0.00187539f $X=5.27 $Y=1.657 $X2=0
+ $Y2=0
cc_360 N_C_c_435_n N_A_882_137#_c_1078_n 0.0141065f $X=4.84 $Y=1.45 $X2=0 $Y2=0
cc_361 N_C_c_436_n N_A_882_137#_c_1078_n 0.011974f $X=5.27 $Y=1.45 $X2=0 $Y2=0
cc_362 C N_A_882_137#_c_1078_n 0.0274003f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_363 N_C_c_438_n N_A_882_137#_c_1078_n 0.00224206f $X=5.27 $Y=1.657 $X2=0
+ $Y2=0
cc_364 N_C_c_436_n N_A_882_137#_c_1072_n 4.61883e-19 $X=5.27 $Y=1.45 $X2=0 $Y2=0
cc_365 C N_A_882_137#_c_1073_n 0.0267022f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_366 N_C_c_435_n N_A_882_137#_c_1075_n 0.00165863f $X=4.84 $Y=1.45 $X2=0 $Y2=0
cc_367 N_C_c_438_n N_A_882_137#_c_1075_n 0.00883774f $X=5.27 $Y=1.657 $X2=0
+ $Y2=0
cc_368 C N_A_882_137#_c_1076_n 0.0204877f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_369 N_C_c_438_n N_A_882_137#_c_1076_n 0.00544331f $X=5.27 $Y=1.657 $X2=0
+ $Y2=0
cc_370 N_D_M1023_g N_A_472_388#_M1006_g 0.0208933f $X=6.69 $Y=0.79 $X2=0 $Y2=0
cc_371 N_D_c_494_n N_A_472_388#_c_553_n 0.0219014f $X=6.73 $Y=1.765 $X2=0 $Y2=0
cc_372 N_D_c_493_n N_A_472_388#_c_601_n 0.0215942f $X=6.225 $Y=1.865 $X2=0 $Y2=0
cc_373 N_D_c_494_n N_A_472_388#_c_609_n 0.0127538f $X=6.73 $Y=1.765 $X2=0 $Y2=0
cc_374 N_D_c_491_n N_A_472_388#_c_609_n 2.24055e-19 $X=6.71 $Y=1.515 $X2=0 $Y2=0
cc_375 N_D_c_492_n N_A_472_388#_c_609_n 0.0136865f $X=6.71 $Y=1.515 $X2=0 $Y2=0
cc_376 N_D_c_494_n N_A_472_388#_c_562_n 0.00335443f $X=6.73 $Y=1.765 $X2=0 $Y2=0
cc_377 N_D_c_491_n N_A_472_388#_c_562_n 3.49588e-19 $X=6.71 $Y=1.515 $X2=0 $Y2=0
cc_378 N_D_c_492_n N_A_472_388#_c_562_n 0.00966496f $X=6.71 $Y=1.515 $X2=0 $Y2=0
cc_379 N_D_M1023_g N_A_472_388#_c_549_n 7.24231e-19 $X=6.69 $Y=0.79 $X2=0 $Y2=0
cc_380 N_D_c_491_n N_A_472_388#_c_549_n 0.0012231f $X=6.71 $Y=1.515 $X2=0 $Y2=0
cc_381 N_D_c_492_n N_A_472_388#_c_549_n 0.0240042f $X=6.71 $Y=1.515 $X2=0 $Y2=0
cc_382 N_D_c_494_n N_A_472_388#_c_563_n 0.0125816f $X=6.73 $Y=1.765 $X2=0 $Y2=0
cc_383 N_D_c_491_n N_A_472_388#_c_563_n 0.00240335f $X=6.71 $Y=1.515 $X2=0 $Y2=0
cc_384 N_D_c_492_n N_A_472_388#_c_563_n 0.0238486f $X=6.71 $Y=1.515 $X2=0 $Y2=0
cc_385 N_D_c_491_n N_A_472_388#_c_552_n 0.0182475f $X=6.71 $Y=1.515 $X2=0 $Y2=0
cc_386 N_D_c_492_n N_A_472_388#_c_552_n 6.29709e-19 $X=6.71 $Y=1.515 $X2=0 $Y2=0
cc_387 N_D_c_493_n N_VPWR_c_723_n 0.00265483f $X=6.225 $Y=1.865 $X2=0 $Y2=0
cc_388 N_D_c_494_n N_VPWR_c_723_n 0.00829628f $X=6.73 $Y=1.765 $X2=0 $Y2=0
cc_389 N_D_c_493_n N_VPWR_c_732_n 0.00505726f $X=6.225 $Y=1.865 $X2=0 $Y2=0
cc_390 N_D_c_494_n N_VPWR_c_732_n 0.00486301f $X=6.73 $Y=1.765 $X2=0 $Y2=0
cc_391 N_D_c_493_n N_VPWR_c_739_n 0.016669f $X=6.225 $Y=1.865 $X2=0 $Y2=0
cc_392 N_D_c_494_n N_VPWR_c_739_n 7.35957e-19 $X=6.73 $Y=1.765 $X2=0 $Y2=0
cc_393 N_D_c_493_n N_VPWR_c_718_n 0.00485508f $X=6.225 $Y=1.865 $X2=0 $Y2=0
cc_394 N_D_c_494_n N_VPWR_c_718_n 0.00508379f $X=6.73 $Y=1.765 $X2=0 $Y2=0
cc_395 N_D_M1023_g N_X_c_838_n 2.04021e-19 $X=6.69 $Y=0.79 $X2=0 $Y2=0
cc_396 N_D_M1008_g N_VGND_c_903_n 0.00354008f $X=6.26 $Y=0.79 $X2=0 $Y2=0
cc_397 N_D_M1008_g N_VGND_c_904_n 5.55326e-19 $X=6.26 $Y=0.79 $X2=0 $Y2=0
cc_398 N_D_M1023_g N_VGND_c_904_n 0.0117856f $X=6.69 $Y=0.79 $X2=0 $Y2=0
cc_399 N_D_c_491_n N_VGND_c_904_n 0.00266105f $X=6.71 $Y=1.515 $X2=0 $Y2=0
cc_400 N_D_c_492_n N_VGND_c_904_n 0.00937578f $X=6.71 $Y=1.515 $X2=0 $Y2=0
cc_401 N_D_M1008_g N_VGND_c_910_n 0.00485498f $X=6.26 $Y=0.79 $X2=0 $Y2=0
cc_402 N_D_M1023_g N_VGND_c_910_n 0.00421418f $X=6.69 $Y=0.79 $X2=0 $Y2=0
cc_403 N_D_M1008_g N_VGND_c_917_n 0.00514438f $X=6.26 $Y=0.79 $X2=0 $Y2=0
cc_404 N_D_M1023_g N_VGND_c_917_n 0.00432128f $X=6.69 $Y=0.79 $X2=0 $Y2=0
cc_405 N_D_M1008_g N_A_882_137#_c_1072_n 0.00294371f $X=6.26 $Y=0.79 $X2=0 $Y2=0
cc_406 N_D_M1008_g N_A_882_137#_c_1073_n 0.0190642f $X=6.26 $Y=0.79 $X2=0 $Y2=0
cc_407 N_D_M1023_g N_A_882_137#_c_1073_n 0.00144374f $X=6.69 $Y=0.79 $X2=0 $Y2=0
cc_408 N_D_c_491_n N_A_882_137#_c_1073_n 0.0043782f $X=6.71 $Y=1.515 $X2=0 $Y2=0
cc_409 N_D_c_492_n N_A_882_137#_c_1073_n 0.0167507f $X=6.71 $Y=1.515 $X2=0 $Y2=0
cc_410 N_D_M1008_g N_A_882_137#_c_1074_n 0.00846733f $X=6.26 $Y=0.79 $X2=0 $Y2=0
cc_411 N_D_M1008_g N_A_882_137#_c_1076_n 0.00280711f $X=6.26 $Y=0.79 $X2=0 $Y2=0
cc_412 N_A_472_388#_c_601_n N_VPWR_M1025_s 0.0297742f $X=6.335 $Y=2.035 $X2=0
+ $Y2=0
cc_413 N_A_472_388#_c_609_n N_VPWR_M1017_d 0.0108309f $X=7.065 $Y=2.035 $X2=0
+ $Y2=0
cc_414 N_A_472_388#_c_562_n N_VPWR_M1017_d 0.00135409f $X=7.15 $Y=1.95 $X2=0
+ $Y2=0
cc_415 N_A_472_388#_c_557_n N_VPWR_c_720_n 0.0222353f $X=2.595 $Y=2.085 $X2=0
+ $Y2=0
cc_416 N_A_472_388#_c_557_n N_VPWR_c_721_n 0.0689299f $X=2.595 $Y=2.085 $X2=0
+ $Y2=0
cc_417 N_A_472_388#_c_547_n N_VPWR_c_721_n 0.0274961f $X=3.465 $Y=1.68 $X2=0
+ $Y2=0
cc_418 N_A_472_388#_c_559_n N_VPWR_c_721_n 0.00191379f $X=3.63 $Y=2.085 $X2=0
+ $Y2=0
cc_419 N_A_472_388#_c_559_n N_VPWR_c_722_n 0.0394173f $X=3.63 $Y=2.085 $X2=0
+ $Y2=0
cc_420 N_A_472_388#_c_548_n N_VPWR_c_722_n 0.027703f $X=4.465 $Y=1.68 $X2=0
+ $Y2=0
cc_421 N_A_472_388#_c_586_n N_VPWR_c_722_n 6.91732e-19 $X=4.63 $Y=1.95 $X2=0
+ $Y2=0
cc_422 N_A_472_388#_c_561_n N_VPWR_c_722_n 0.0322718f $X=4.63 $Y=2.795 $X2=0
+ $Y2=0
cc_423 N_A_472_388#_c_553_n N_VPWR_c_723_n 0.0119495f $X=7.265 $Y=1.765 $X2=0
+ $Y2=0
cc_424 N_A_472_388#_c_554_n N_VPWR_c_723_n 5.35985e-19 $X=7.715 $Y=1.765 $X2=0
+ $Y2=0
cc_425 N_A_472_388#_c_609_n N_VPWR_c_723_n 0.022569f $X=7.065 $Y=2.035 $X2=0
+ $Y2=0
cc_426 N_A_472_388#_c_563_n N_VPWR_c_723_n 0.0376406f $X=6.5 $Y=2.065 $X2=0
+ $Y2=0
cc_427 N_A_472_388#_c_553_n N_VPWR_c_724_n 5.26866e-19 $X=7.265 $Y=1.765 $X2=0
+ $Y2=0
cc_428 N_A_472_388#_c_554_n N_VPWR_c_724_n 0.0112323f $X=7.715 $Y=1.765 $X2=0
+ $Y2=0
cc_429 N_A_472_388#_c_555_n N_VPWR_c_724_n 0.0160972f $X=8.165 $Y=1.765 $X2=0
+ $Y2=0
cc_430 N_A_472_388#_c_556_n N_VPWR_c_724_n 0.00227565f $X=8.615 $Y=1.765 $X2=0
+ $Y2=0
cc_431 N_A_472_388#_c_555_n N_VPWR_c_726_n 0.00227565f $X=8.165 $Y=1.765 $X2=0
+ $Y2=0
cc_432 N_A_472_388#_c_556_n N_VPWR_c_726_n 0.0169867f $X=8.615 $Y=1.765 $X2=0
+ $Y2=0
cc_433 N_A_472_388#_c_557_n N_VPWR_c_730_n 0.0135468f $X=2.595 $Y=2.085 $X2=0
+ $Y2=0
cc_434 N_A_472_388#_c_559_n N_VPWR_c_731_n 0.0135062f $X=3.63 $Y=2.085 $X2=0
+ $Y2=0
cc_435 N_A_472_388#_c_563_n N_VPWR_c_732_n 0.0092875f $X=6.5 $Y=2.065 $X2=0
+ $Y2=0
cc_436 N_A_472_388#_c_553_n N_VPWR_c_733_n 0.00413917f $X=7.265 $Y=1.765 $X2=0
+ $Y2=0
cc_437 N_A_472_388#_c_554_n N_VPWR_c_733_n 0.00413917f $X=7.715 $Y=1.765 $X2=0
+ $Y2=0
cc_438 N_A_472_388#_c_555_n N_VPWR_c_734_n 0.00413917f $X=8.165 $Y=1.765 $X2=0
+ $Y2=0
cc_439 N_A_472_388#_c_556_n N_VPWR_c_734_n 0.00413917f $X=8.615 $Y=1.765 $X2=0
+ $Y2=0
cc_440 N_A_472_388#_c_561_n N_VPWR_c_738_n 0.0134657f $X=4.63 $Y=2.795 $X2=0
+ $Y2=0
cc_441 N_A_472_388#_c_561_n N_VPWR_c_739_n 0.0261074f $X=4.63 $Y=2.795 $X2=0
+ $Y2=0
cc_442 N_A_472_388#_c_601_n N_VPWR_c_739_n 0.0906832f $X=6.335 $Y=2.035 $X2=0
+ $Y2=0
cc_443 N_A_472_388#_c_553_n N_VPWR_c_718_n 0.00817726f $X=7.265 $Y=1.765 $X2=0
+ $Y2=0
cc_444 N_A_472_388#_c_554_n N_VPWR_c_718_n 0.00817726f $X=7.715 $Y=1.765 $X2=0
+ $Y2=0
cc_445 N_A_472_388#_c_555_n N_VPWR_c_718_n 0.00817726f $X=8.165 $Y=1.765 $X2=0
+ $Y2=0
cc_446 N_A_472_388#_c_556_n N_VPWR_c_718_n 0.00817726f $X=8.615 $Y=1.765 $X2=0
+ $Y2=0
cc_447 N_A_472_388#_c_557_n N_VPWR_c_718_n 0.0119671f $X=2.595 $Y=2.085 $X2=0
+ $Y2=0
cc_448 N_A_472_388#_c_559_n N_VPWR_c_718_n 0.0119552f $X=3.63 $Y=2.085 $X2=0
+ $Y2=0
cc_449 N_A_472_388#_c_561_n N_VPWR_c_718_n 0.0119432f $X=4.63 $Y=2.795 $X2=0
+ $Y2=0
cc_450 N_A_472_388#_c_563_n N_VPWR_c_718_n 0.0111958f $X=6.5 $Y=2.065 $X2=0
+ $Y2=0
cc_451 N_A_472_388#_M1006_g N_X_c_838_n 0.00761489f $X=7.19 $Y=0.74 $X2=0 $Y2=0
cc_452 N_A_472_388#_M1009_g N_X_c_838_n 0.00931022f $X=7.62 $Y=0.74 $X2=0 $Y2=0
cc_453 N_A_472_388#_M1014_g N_X_c_838_n 5.61679e-19 $X=8.15 $Y=0.74 $X2=0 $Y2=0
cc_454 N_A_472_388#_c_553_n N_X_c_845_n 0.00203182f $X=7.265 $Y=1.765 $X2=0
+ $Y2=0
cc_455 N_A_472_388#_c_609_n N_X_c_845_n 0.0148585f $X=7.065 $Y=2.035 $X2=0 $Y2=0
cc_456 N_A_472_388#_c_562_n N_X_c_845_n 0.0102617f $X=7.15 $Y=1.95 $X2=0 $Y2=0
cc_457 N_A_472_388#_c_668_p N_X_c_845_n 0.0143367f $X=8.4 $Y=1.485 $X2=0 $Y2=0
cc_458 N_A_472_388#_c_552_n N_X_c_845_n 0.00443356f $X=8.615 $Y=1.542 $X2=0
+ $Y2=0
cc_459 N_A_472_388#_c_553_n N_X_c_846_n 0.00518554f $X=7.265 $Y=1.765 $X2=0
+ $Y2=0
cc_460 N_A_472_388#_c_554_n N_X_c_846_n 0.00567416f $X=7.715 $Y=1.765 $X2=0
+ $Y2=0
cc_461 N_A_472_388#_M1006_g N_X_c_839_n 0.00277457f $X=7.19 $Y=0.74 $X2=0 $Y2=0
cc_462 N_A_472_388#_M1009_g N_X_c_839_n 0.00121617f $X=7.62 $Y=0.74 $X2=0 $Y2=0
cc_463 N_A_472_388#_c_668_p N_X_c_839_n 0.0276081f $X=8.4 $Y=1.485 $X2=0 $Y2=0
cc_464 N_A_472_388#_c_552_n N_X_c_839_n 0.00232957f $X=8.615 $Y=1.542 $X2=0
+ $Y2=0
cc_465 N_A_472_388#_c_554_n N_X_c_847_n 0.0176877f $X=7.715 $Y=1.765 $X2=0 $Y2=0
cc_466 N_A_472_388#_c_555_n N_X_c_847_n 0.0176407f $X=8.165 $Y=1.765 $X2=0 $Y2=0
cc_467 N_A_472_388#_c_556_n N_X_c_847_n 0.0220078f $X=8.615 $Y=1.765 $X2=0 $Y2=0
cc_468 N_A_472_388#_c_668_p N_X_c_847_n 0.0769748f $X=8.4 $Y=1.485 $X2=0 $Y2=0
cc_469 N_A_472_388#_c_552_n N_X_c_847_n 0.0169459f $X=8.615 $Y=1.542 $X2=0 $Y2=0
cc_470 N_A_472_388#_M1018_g N_X_c_840_n 0.0206679f $X=8.62 $Y=0.74 $X2=0 $Y2=0
cc_471 N_A_472_388#_c_552_n N_X_c_841_n 0.00319865f $X=8.615 $Y=1.542 $X2=0
+ $Y2=0
cc_472 N_A_472_388#_M1009_g N_X_c_842_n 0.0116357f $X=7.62 $Y=0.74 $X2=0 $Y2=0
cc_473 N_A_472_388#_M1014_g N_X_c_842_n 0.014058f $X=8.15 $Y=0.74 $X2=0 $Y2=0
cc_474 N_A_472_388#_c_668_p N_X_c_842_n 0.0751459f $X=8.4 $Y=1.485 $X2=0 $Y2=0
cc_475 N_A_472_388#_c_552_n N_X_c_842_n 0.00452522f $X=8.615 $Y=1.542 $X2=0
+ $Y2=0
cc_476 N_A_472_388#_c_556_n X 0.00212519f $X=8.615 $Y=1.765 $X2=0 $Y2=0
cc_477 N_A_472_388#_M1018_g X 0.0213283f $X=8.62 $Y=0.74 $X2=0 $Y2=0
cc_478 N_A_472_388#_c_668_p X 0.0236873f $X=8.4 $Y=1.485 $X2=0 $Y2=0
cc_479 N_A_472_388#_M1006_g N_VGND_c_904_n 0.00730861f $X=7.19 $Y=0.74 $X2=0
+ $Y2=0
cc_480 N_A_472_388#_M1009_g N_VGND_c_905_n 0.00438574f $X=7.62 $Y=0.74 $X2=0
+ $Y2=0
cc_481 N_A_472_388#_M1014_g N_VGND_c_905_n 0.00260786f $X=8.15 $Y=0.74 $X2=0
+ $Y2=0
cc_482 N_A_472_388#_M1014_g N_VGND_c_907_n 0.00110236f $X=8.15 $Y=0.74 $X2=0
+ $Y2=0
cc_483 N_A_472_388#_M1018_g N_VGND_c_907_n 0.0101865f $X=8.62 $Y=0.74 $X2=0
+ $Y2=0
cc_484 N_A_472_388#_M1006_g N_VGND_c_911_n 0.00434272f $X=7.19 $Y=0.74 $X2=0
+ $Y2=0
cc_485 N_A_472_388#_M1009_g N_VGND_c_911_n 0.00434272f $X=7.62 $Y=0.74 $X2=0
+ $Y2=0
cc_486 N_A_472_388#_M1014_g N_VGND_c_912_n 0.00461464f $X=8.15 $Y=0.74 $X2=0
+ $Y2=0
cc_487 N_A_472_388#_M1018_g N_VGND_c_912_n 0.00383152f $X=8.62 $Y=0.74 $X2=0
+ $Y2=0
cc_488 N_A_472_388#_M1006_g N_VGND_c_917_n 0.00825059f $X=7.19 $Y=0.74 $X2=0
+ $Y2=0
cc_489 N_A_472_388#_M1009_g N_VGND_c_917_n 0.00820974f $X=7.62 $Y=0.74 $X2=0
+ $Y2=0
cc_490 N_A_472_388#_M1014_g N_VGND_c_917_n 0.00908514f $X=8.15 $Y=0.74 $X2=0
+ $Y2=0
cc_491 N_A_472_388#_M1018_g N_VGND_c_917_n 0.00369657f $X=8.62 $Y=0.74 $X2=0
+ $Y2=0
cc_492 N_A_472_388#_M1007_d N_A_412_140#_c_1005_n 0.00319077f $X=2.565 $Y=0.7
+ $X2=0 $Y2=0
cc_493 N_A_472_388#_c_547_n N_A_412_140#_c_1005_n 0.00349748f $X=3.465 $Y=1.68
+ $X2=0 $Y2=0
cc_494 N_A_472_388#_c_574_n N_A_412_140#_c_1005_n 0.00265382f $X=2.595 $Y=1.68
+ $X2=0 $Y2=0
cc_495 N_A_472_388#_c_550_n N_A_412_140#_c_1005_n 0.0167843f $X=2.705 $Y=1.185
+ $X2=0 $Y2=0
cc_496 N_A_472_388#_c_547_n N_A_412_140#_c_1000_n 0.0169856f $X=3.465 $Y=1.68
+ $X2=0 $Y2=0
cc_497 N_A_472_388#_c_548_n N_A_412_140#_c_1000_n 0.00233842f $X=4.465 $Y=1.68
+ $X2=0 $Y2=0
cc_498 N_A_472_388#_c_551_n N_A_412_140#_c_1000_n 0.027396f $X=3.63 $Y=1.68
+ $X2=0 $Y2=0
cc_499 N_A_472_388#_c_546_n N_A_412_140#_c_1001_n 0.00379815f $X=2.65 $Y=1.595
+ $X2=0 $Y2=0
cc_500 N_A_472_388#_c_547_n N_A_412_140#_c_1001_n 0.0143406f $X=3.465 $Y=1.68
+ $X2=0 $Y2=0
cc_501 N_A_472_388#_c_550_n N_A_412_140#_c_1001_n 0.00463069f $X=2.705 $Y=1.185
+ $X2=0 $Y2=0
cc_502 N_A_472_388#_c_548_n N_A_412_140#_c_1002_n 0.0252298f $X=4.465 $Y=1.68
+ $X2=0 $Y2=0
cc_503 N_A_472_388#_c_548_n N_A_685_140#_c_1044_n 0.00641663f $X=4.465 $Y=1.68
+ $X2=0 $Y2=0
cc_504 N_A_472_388#_c_548_n N_A_882_137#_c_1078_n 0.00254662f $X=4.465 $Y=1.68
+ $X2=0 $Y2=0
cc_505 N_A_472_388#_c_601_n N_A_882_137#_c_1078_n 0.00273534f $X=6.335 $Y=2.035
+ $X2=0 $Y2=0
cc_506 N_A_472_388#_c_548_n N_A_882_137#_c_1075_n 0.0198005f $X=4.465 $Y=1.68
+ $X2=0 $Y2=0
cc_507 N_VPWR_c_723_n N_X_c_846_n 0.0449718f $X=7.04 $Y=2.455 $X2=0 $Y2=0
cc_508 N_VPWR_c_724_n N_X_c_846_n 0.0430177f $X=7.94 $Y=2.405 $X2=0 $Y2=0
cc_509 N_VPWR_c_733_n N_X_c_846_n 0.00749631f $X=7.775 $Y=3.33 $X2=0 $Y2=0
cc_510 N_VPWR_c_718_n N_X_c_846_n 0.0062048f $X=8.88 $Y=3.33 $X2=0 $Y2=0
cc_511 N_VPWR_M1013_s N_X_c_847_n 0.00201799f $X=7.79 $Y=1.84 $X2=0 $Y2=0
cc_512 N_VPWR_c_724_n N_X_c_847_n 0.0179913f $X=7.94 $Y=2.405 $X2=0 $Y2=0
cc_513 N_VPWR_c_726_n N_X_c_847_n 0.00256809f $X=8.84 $Y=2.405 $X2=0 $Y2=0
cc_514 N_VPWR_M1016_s N_X_c_849_n 0.00440781f $X=8.69 $Y=1.84 $X2=0 $Y2=0
cc_515 N_VPWR_c_726_n N_X_c_849_n 0.0207257f $X=8.84 $Y=2.405 $X2=0 $Y2=0
cc_516 N_X_c_842_n N_VGND_M1009_d 0.00297044f $X=8.24 $Y=0.96 $X2=0 $Y2=0
cc_517 N_X_c_844_n N_VGND_M1018_d 0.00445656f $X=8.88 $Y=1.15 $X2=0 $Y2=0
cc_518 N_X_c_838_n N_VGND_c_904_n 0.0243921f $X=7.405 $Y=0.515 $X2=0 $Y2=0
cc_519 N_X_c_839_n N_VGND_c_904_n 0.00711243f $X=7.57 $Y=1.065 $X2=0 $Y2=0
cc_520 N_X_c_838_n N_VGND_c_905_n 0.0180508f $X=7.405 $Y=0.515 $X2=0 $Y2=0
cc_521 N_X_c_842_n N_VGND_c_905_n 0.0216414f $X=8.24 $Y=0.96 $X2=0 $Y2=0
cc_522 N_X_c_840_n N_VGND_c_907_n 0.00288208f $X=8.765 $Y=0.96 $X2=0 $Y2=0
cc_523 N_X_c_844_n N_VGND_c_907_n 0.0201316f $X=8.88 $Y=1.15 $X2=0 $Y2=0
cc_524 N_X_c_838_n N_VGND_c_911_n 0.0144922f $X=7.405 $Y=0.515 $X2=0 $Y2=0
cc_525 N_X_c_838_n N_VGND_c_917_n 0.0118826f $X=7.405 $Y=0.515 $X2=0 $Y2=0
cc_526 N_X_c_840_n N_VGND_c_917_n 3.49881e-19 $X=8.765 $Y=0.96 $X2=0 $Y2=0
cc_527 N_X_c_841_n N_VGND_c_917_n 0.0160493f $X=8.43 $Y=0.96 $X2=0 $Y2=0
cc_528 N_X_c_844_n N_VGND_c_917_n 9.31328e-19 $X=8.88 $Y=1.15 $X2=0 $Y2=0
cc_529 N_X_c_839_n N_A_882_137#_c_1073_n 6.08693e-19 $X=7.57 $Y=1.065 $X2=0
+ $Y2=0
cc_530 N_VGND_c_909_n N_A_685_140#_c_1045_n 6.22085e-19 $X=5.88 $Y=0 $X2=0 $Y2=0
cc_531 N_VGND_c_917_n N_A_685_140#_c_1045_n 0.00153572f $X=8.88 $Y=0 $X2=0 $Y2=0
cc_532 N_VGND_c_909_n N_A_685_140#_c_1043_n 0.00575291f $X=5.88 $Y=0 $X2=0 $Y2=0
cc_533 N_VGND_c_917_n N_A_685_140#_c_1043_n 0.00933739f $X=8.88 $Y=0 $X2=0 $Y2=0
cc_534 N_VGND_c_909_n N_A_685_140#_c_1044_n 0.0156902f $X=5.88 $Y=0 $X2=0 $Y2=0
cc_535 N_VGND_c_917_n N_A_685_140#_c_1044_n 0.0319574f $X=8.88 $Y=0 $X2=0 $Y2=0
cc_536 N_VGND_c_903_n N_A_882_137#_c_1072_n 0.0113125f $X=6.045 $Y=0.645 $X2=0
+ $Y2=0
cc_537 N_VGND_c_909_n N_A_882_137#_c_1072_n 0.00468849f $X=5.88 $Y=0 $X2=0 $Y2=0
cc_538 N_VGND_c_917_n N_A_882_137#_c_1072_n 0.00732591f $X=8.88 $Y=0 $X2=0 $Y2=0
cc_539 N_VGND_M1008_d N_A_882_137#_c_1073_n 0.00299905f $X=5.9 $Y=0.47 $X2=0
+ $Y2=0
cc_540 N_VGND_c_903_n N_A_882_137#_c_1073_n 0.0201545f $X=6.045 $Y=0.645 $X2=0
+ $Y2=0
cc_541 N_VGND_c_904_n N_A_882_137#_c_1073_n 0.00517071f $X=6.905 $Y=0.615 $X2=0
+ $Y2=0
cc_542 N_VGND_c_903_n N_A_882_137#_c_1074_n 0.0141239f $X=6.045 $Y=0.645 $X2=0
+ $Y2=0
cc_543 N_VGND_c_904_n N_A_882_137#_c_1074_n 0.0207991f $X=6.905 $Y=0.615 $X2=0
+ $Y2=0
cc_544 N_VGND_c_910_n N_A_882_137#_c_1074_n 0.0078096f $X=6.74 $Y=0 $X2=0 $Y2=0
cc_545 N_VGND_c_917_n N_A_882_137#_c_1074_n 0.0085649f $X=8.88 $Y=0 $X2=0 $Y2=0
cc_546 N_A_412_140#_c_1000_n N_A_685_140#_M1000_d 0.00168967f $X=3.83 $Y=1.34
+ $X2=-0.19 $Y2=-0.245
cc_547 N_A_412_140#_c_1000_n N_A_685_140#_c_1045_n 0.0144331f $X=3.83 $Y=1.34
+ $X2=0 $Y2=0
cc_548 N_A_412_140#_M1002_s N_A_685_140#_c_1044_n 0.00785889f $X=3.855 $Y=0.7
+ $X2=0 $Y2=0
cc_549 N_A_412_140#_c_1000_n N_A_685_140#_c_1044_n 0.00496071f $X=3.83 $Y=1.34
+ $X2=0 $Y2=0
cc_550 N_A_412_140#_c_1002_n N_A_685_140#_c_1044_n 0.0207078f $X=3.995 $Y=1.185
+ $X2=0 $Y2=0
cc_551 N_A_412_140#_c_1002_n N_A_882_137#_c_1075_n 0.0174387f $X=3.995 $Y=1.185
+ $X2=0 $Y2=0
cc_552 N_A_685_140#_c_1044_n N_A_882_137#_M1001_s 0.0103513f $X=4.89 $Y=0.802
+ $X2=-0.19 $Y2=-0.245
cc_553 N_A_685_140#_M1001_d N_A_882_137#_c_1078_n 0.00330913f $X=4.915 $Y=0.685
+ $X2=0 $Y2=0
cc_554 N_A_685_140#_c_1043_n N_A_882_137#_c_1078_n 0.0159532f $X=5.055 $Y=0.84
+ $X2=0 $Y2=0
cc_555 N_A_685_140#_c_1044_n N_A_882_137#_c_1078_n 0.0078857f $X=4.89 $Y=0.802
+ $X2=0 $Y2=0
cc_556 N_A_685_140#_c_1043_n N_A_882_137#_c_1072_n 0.0112424f $X=5.055 $Y=0.84
+ $X2=0 $Y2=0
cc_557 N_A_685_140#_c_1044_n N_A_882_137#_c_1075_n 0.0238397f $X=4.89 $Y=0.802
+ $X2=0 $Y2=0
