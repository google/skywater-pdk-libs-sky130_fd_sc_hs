* File: sky130_fd_sc_hs__a21bo_4.pxi.spice
* Created: Tue Sep  1 19:49:10 2020
* 
x_PM_SKY130_FD_SC_HS__A21BO_4%B1_N N_B1_N_c_117_n N_B1_N_c_123_n N_B1_N_M1018_g
+ N_B1_N_M1005_g N_B1_N_c_119_n B1_N N_B1_N_c_121_n
+ PM_SKY130_FD_SC_HS__A21BO_4%B1_N
x_PM_SKY130_FD_SC_HS__A21BO_4%A_187_338# N_A_187_338#_M1015_s
+ N_A_187_338#_M1006_s N_A_187_338#_M1014_d N_A_187_338#_c_164_n
+ N_A_187_338#_M1004_g N_A_187_338#_c_152_n N_A_187_338#_M1001_g
+ N_A_187_338#_c_165_n N_A_187_338#_M1007_g N_A_187_338#_c_153_n
+ N_A_187_338#_M1003_g N_A_187_338#_c_166_n N_A_187_338#_M1011_g
+ N_A_187_338#_c_154_n N_A_187_338#_M1008_g N_A_187_338#_c_167_n
+ N_A_187_338#_M1013_g N_A_187_338#_c_155_n N_A_187_338#_M1010_g
+ N_A_187_338#_c_198_p N_A_187_338#_c_156_n N_A_187_338#_c_157_n
+ N_A_187_338#_c_158_n N_A_187_338#_c_159_n N_A_187_338#_c_160_n
+ N_A_187_338#_c_161_n N_A_187_338#_c_162_n N_A_187_338#_c_163_n
+ PM_SKY130_FD_SC_HS__A21BO_4%A_187_338#
x_PM_SKY130_FD_SC_HS__A21BO_4%A_29_392# N_A_29_392#_M1005_s N_A_29_392#_M1018_s
+ N_A_29_392#_M1015_g N_A_29_392#_c_314_n N_A_29_392#_M1014_g
+ N_A_29_392#_c_308_n N_A_29_392#_M1021_g N_A_29_392#_c_310_n
+ N_A_29_392#_c_317_n N_A_29_392#_M1016_g N_A_29_392#_c_311_n
+ N_A_29_392#_c_319_n N_A_29_392#_c_328_n N_A_29_392#_c_379_p
+ N_A_29_392#_c_320_n N_A_29_392#_c_362_n N_A_29_392#_c_312_n
+ N_A_29_392#_c_313_n N_A_29_392#_c_322_n PM_SKY130_FD_SC_HS__A21BO_4%A_29_392#
x_PM_SKY130_FD_SC_HS__A21BO_4%A1 N_A1_c_424_n N_A1_M1000_g N_A1_M1006_g
+ N_A1_c_425_n N_A1_M1019_g N_A1_M1012_g A1 A1 N_A1_c_423_n
+ PM_SKY130_FD_SC_HS__A21BO_4%A1
x_PM_SKY130_FD_SC_HS__A21BO_4%A2 N_A2_c_467_n N_A2_c_468_n N_A2_c_477_n
+ N_A2_M1002_g N_A2_M1009_g N_A2_c_470_n N_A2_c_471_n N_A2_c_472_n N_A2_c_479_n
+ N_A2_M1017_g N_A2_M1020_g A2 N_A2_c_474_n N_A2_c_475_n
+ PM_SKY130_FD_SC_HS__A21BO_4%A2
x_PM_SKY130_FD_SC_HS__A21BO_4%VPWR N_VPWR_M1018_d N_VPWR_M1007_s N_VPWR_M1013_s
+ N_VPWR_M1002_s N_VPWR_M1019_d N_VPWR_c_541_n N_VPWR_c_542_n N_VPWR_c_543_n
+ N_VPWR_c_544_n N_VPWR_c_545_n N_VPWR_c_546_n N_VPWR_c_547_n N_VPWR_c_548_n
+ N_VPWR_c_549_n VPWR N_VPWR_c_550_n N_VPWR_c_551_n N_VPWR_c_552_n
+ N_VPWR_c_553_n N_VPWR_c_540_n N_VPWR_c_555_n N_VPWR_c_556_n N_VPWR_c_557_n
+ PM_SKY130_FD_SC_HS__A21BO_4%VPWR
x_PM_SKY130_FD_SC_HS__A21BO_4%X N_X_M1001_d N_X_M1008_d N_X_M1004_d N_X_M1011_d
+ N_X_c_628_n N_X_c_629_n N_X_c_642_n N_X_c_647_n N_X_c_630_n N_X_c_653_n
+ N_X_c_631_n N_X_c_657_n X PM_SKY130_FD_SC_HS__A21BO_4%X
x_PM_SKY130_FD_SC_HS__A21BO_4%A_596_392# N_A_596_392#_M1014_s
+ N_A_596_392#_M1016_s N_A_596_392#_M1000_s N_A_596_392#_M1017_d
+ N_A_596_392#_c_683_n N_A_596_392#_c_684_n N_A_596_392#_c_685_n
+ N_A_596_392#_c_686_n N_A_596_392#_c_700_n N_A_596_392#_c_687_n
+ N_A_596_392#_c_688_n N_A_596_392#_c_689_n N_A_596_392#_c_690_n
+ N_A_596_392#_c_691_n N_A_596_392#_c_692_n
+ PM_SKY130_FD_SC_HS__A21BO_4%A_596_392#
x_PM_SKY130_FD_SC_HS__A21BO_4%VGND N_VGND_M1005_d N_VGND_M1003_s N_VGND_M1010_s
+ N_VGND_M1021_d N_VGND_M1020_d N_VGND_c_754_n N_VGND_c_755_n N_VGND_c_756_n
+ N_VGND_c_757_n N_VGND_c_758_n N_VGND_c_759_n N_VGND_c_760_n N_VGND_c_761_n
+ N_VGND_c_762_n N_VGND_c_763_n N_VGND_c_764_n N_VGND_c_765_n VGND
+ N_VGND_c_766_n N_VGND_c_767_n N_VGND_c_768_n N_VGND_c_769_n
+ PM_SKY130_FD_SC_HS__A21BO_4%VGND
x_PM_SKY130_FD_SC_HS__A21BO_4%A_864_123# N_A_864_123#_M1009_s
+ N_A_864_123#_M1012_d N_A_864_123#_c_841_n N_A_864_123#_c_842_n
+ N_A_864_123#_c_843_n N_A_864_123#_c_844_n
+ PM_SKY130_FD_SC_HS__A21BO_4%A_864_123#
cc_1 VNB N_B1_N_c_117_n 0.0124344f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.795
cc_2 VNB N_B1_N_M1005_g 0.00796521f $X=-0.19 $Y=-0.245 $X2=0.665 $Y2=0.935
cc_3 VNB N_B1_N_c_119_n 0.0214147f $X=-0.19 $Y=-0.245 $X2=0.665 $Y2=1.405
cc_4 VNB B1_N 0.0230286f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.47
cc_5 VNB N_B1_N_c_121_n 0.0578415f $X=-0.19 $Y=-0.245 $X2=0.665 $Y2=0.34
cc_6 VNB N_A_187_338#_c_152_n 0.0173822f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_7 VNB N_A_187_338#_c_153_n 0.015779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_A_187_338#_c_154_n 0.0162345f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A_187_338#_c_155_n 0.0173813f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_187_338#_c_156_n 0.0824931f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_187_338#_c_157_n 0.00321807f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_187_338#_c_158_n 0.00349665f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_187_338#_c_159_n 0.00300874f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_187_338#_c_160_n 0.0131087f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_187_338#_c_161_n 0.00490329f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_187_338#_c_162_n 0.00145889f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_187_338#_c_163_n 0.0030898f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_29_392#_M1015_g 0.0218255f $X=-0.19 $Y=-0.245 $X2=0.665 $Y2=0.935
cc_19 VNB N_A_29_392#_c_308_n 0.0402881f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.47
cc_20 VNB N_A_29_392#_M1021_g 0.0230599f $X=-0.19 $Y=-0.245 $X2=0.46 $Y2=0.34
cc_21 VNB N_A_29_392#_c_310_n 0.00299868f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_29_392#_c_311_n 0.0190292f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_29_392#_c_312_n 8.33235e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_29_392#_c_313_n 0.0246733f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A1_M1006_g 0.0198169f $X=-0.19 $Y=-0.245 $X2=0.665 $Y2=0.505
cc_26 VNB N_A1_M1012_g 0.0183217f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB A1 0.00366019f $X=-0.19 $Y=-0.245 $X2=0.46 $Y2=0.34
cc_28 VNB N_A1_c_423_n 0.0258387f $X=-0.19 $Y=-0.245 $X2=0.46 $Y2=0.462
cc_29 VNB N_A2_c_467_n 0.00698561f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.48
cc_30 VNB N_A2_c_468_n 0.0138626f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.795
cc_31 VNB N_A2_M1009_g 0.0110175f $X=-0.19 $Y=-0.245 $X2=0.665 $Y2=0.935
cc_32 VNB N_A2_c_470_n 0.0959582f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.405
cc_33 VNB N_A2_c_471_n 0.00840425f $X=-0.19 $Y=-0.245 $X2=0.665 $Y2=1.405
cc_34 VNB N_A2_c_472_n 0.0203569f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A2_M1020_g 0.0257185f $X=-0.19 $Y=-0.245 $X2=0.665 $Y2=0.34
cc_36 VNB N_A2_c_474_n 0.0512238f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A2_c_475_n 7.54705e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_VPWR_c_540_n 0.263193f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_X_c_628_n 0.00252572f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_X_c_629_n 0.00107068f $X=-0.19 $Y=-0.245 $X2=0.46 $Y2=0.34
cc_41 VNB N_X_c_630_n 0.00252589f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_X_c_631_n 0.00690082f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_754_n 0.0185583f $X=-0.19 $Y=-0.245 $X2=0.46 $Y2=0.34
cc_44 VNB N_VGND_c_755_n 0.0122133f $X=-0.19 $Y=-0.245 $X2=0.46 $Y2=0.462
cc_45 VNB N_VGND_c_756_n 0.0178473f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_VGND_c_757_n 0.015487f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_VGND_c_758_n 0.022222f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_VGND_c_759_n 0.0189061f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_VGND_c_760_n 0.0154628f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_VGND_c_761_n 0.0536926f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_VGND_c_762_n 0.0225119f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_VGND_c_763_n 0.00480499f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_VGND_c_764_n 0.0200603f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_VGND_c_765_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_VGND_c_766_n 0.0481317f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_VGND_c_767_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_VGND_c_768_n 0.00326658f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_VGND_c_769_n 0.367636f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_A_864_123#_c_841_n 0.00391695f $X=-0.19 $Y=-0.245 $X2=0.665
+ $Y2=0.935
cc_60 VNB N_A_864_123#_c_842_n 0.00824493f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_A_864_123#_c_843_n 9.0125e-19 $X=-0.19 $Y=-0.245 $X2=0.665 $Y2=1.405
cc_62 VNB N_A_864_123#_c_844_n 0.00549412f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VPB N_B1_N_c_117_n 0.00926301f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.795
cc_64 VPB N_B1_N_c_123_n 0.0275745f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.885
cc_65 VPB N_A_187_338#_c_164_n 0.0148939f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.405
cc_66 VPB N_A_187_338#_c_165_n 0.0147839f $X=-0.19 $Y=1.66 $X2=0.46 $Y2=0.34
cc_67 VPB N_A_187_338#_c_166_n 0.0151052f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=0.462
cc_68 VPB N_A_187_338#_c_167_n 0.0177347f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_69 VPB N_A_187_338#_c_156_n 0.051951f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_70 VPB N_A_187_338#_c_159_n 0.00203648f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_71 VPB N_A_187_338#_c_163_n 0.00170132f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_72 VPB N_A_29_392#_c_314_n 0.017331f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_73 VPB N_A_29_392#_c_308_n 0.0270234f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=0.47
cc_74 VPB N_A_29_392#_c_310_n 0.00679201f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_75 VPB N_A_29_392#_c_317_n 0.0203788f $X=-0.19 $Y=1.66 $X2=0.665 $Y2=0.34
cc_76 VPB N_A_29_392#_c_311_n 0.0244627f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_77 VPB N_A_29_392#_c_319_n 0.0236291f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_78 VPB N_A_29_392#_c_320_n 0.0119625f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_79 VPB N_A_29_392#_c_312_n 9.8204e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_80 VPB N_A_29_392#_c_322_n 0.00717518f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_81 VPB N_A1_c_424_n 0.0157872f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.48
cc_82 VPB N_A1_c_425_n 0.0157872f $X=-0.19 $Y=1.66 $X2=0.665 $Y2=0.935
cc_83 VPB A1 0.00266425f $X=-0.19 $Y=1.66 $X2=0.46 $Y2=0.34
cc_84 VPB N_A1_c_423_n 0.0318087f $X=-0.19 $Y=1.66 $X2=0.46 $Y2=0.462
cc_85 VPB N_A2_c_468_n 0.00755845f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.795
cc_86 VPB N_A2_c_477_n 0.021209f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.885
cc_87 VPB N_A2_c_472_n 0.0114819f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_88 VPB N_A2_c_479_n 0.0284588f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=0.47
cc_89 VPB N_VPWR_c_541_n 0.00591026f $X=-0.19 $Y=1.66 $X2=0.46 $Y2=0.34
cc_90 VPB N_VPWR_c_542_n 0.00261791f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=0.462
cc_91 VPB N_VPWR_c_543_n 0.00953806f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_92 VPB N_VPWR_c_544_n 0.00571271f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_93 VPB N_VPWR_c_545_n 0.00571271f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_94 VPB N_VPWR_c_546_n 0.0376026f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_95 VPB N_VPWR_c_547_n 0.00460249f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_96 VPB N_VPWR_c_548_n 0.0206041f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_97 VPB N_VPWR_c_549_n 0.00460249f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_98 VPB N_VPWR_c_550_n 0.0193106f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_99 VPB N_VPWR_c_551_n 0.0177589f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_100 VPB N_VPWR_c_552_n 0.0177589f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_101 VPB N_VPWR_c_553_n 0.0229598f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_102 VPB N_VPWR_c_540_n 0.109144f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_103 VPB N_VPWR_c_555_n 0.00614127f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_104 VPB N_VPWR_c_556_n 0.00601644f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_105 VPB N_VPWR_c_557_n 0.00614127f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_106 VPB N_X_c_631_n 0.00290489f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_107 VPB N_A_596_392#_c_683_n 0.00812364f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_108 VPB N_A_596_392#_c_684_n 0.00478015f $X=-0.19 $Y=1.66 $X2=0.46 $Y2=0.34
cc_109 VPB N_A_596_392#_c_685_n 0.00424137f $X=-0.19 $Y=1.66 $X2=0.46 $Y2=0.34
cc_110 VPB N_A_596_392#_c_686_n 0.00318119f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_111 VPB N_A_596_392#_c_687_n 0.00462722f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_112 VPB N_A_596_392#_c_688_n 0.00257348f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_113 VPB N_A_596_392#_c_689_n 0.00649597f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_114 VPB N_A_596_392#_c_690_n 0.0121739f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_115 VPB N_A_596_392#_c_691_n 0.0345863f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_116 VPB N_A_596_392#_c_692_n 0.00183558f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_117 N_B1_N_c_123_n N_A_187_338#_c_164_n 0.0333479f $X=0.495 $Y=1.885 $X2=0
+ $Y2=0
cc_118 N_B1_N_c_121_n N_A_187_338#_c_152_n 0.0189708f $X=0.665 $Y=0.34 $X2=0
+ $Y2=0
cc_119 N_B1_N_c_117_n N_A_187_338#_c_156_n 0.00900137f $X=0.495 $Y=1.795 $X2=0
+ $Y2=0
cc_120 N_B1_N_c_119_n N_A_187_338#_c_156_n 0.00934283f $X=0.665 $Y=1.405 $X2=0
+ $Y2=0
cc_121 B1_N N_A_29_392#_M1005_s 0.00103744f $X=0.155 $Y=0.47 $X2=-0.19
+ $Y2=-0.245
cc_122 N_B1_N_c_117_n N_A_29_392#_c_311_n 0.0101392f $X=0.495 $Y=1.795 $X2=0
+ $Y2=0
cc_123 N_B1_N_c_123_n N_A_29_392#_c_311_n 0.00992502f $X=0.495 $Y=1.885 $X2=0
+ $Y2=0
cc_124 N_B1_N_c_119_n N_A_29_392#_c_311_n 0.00715308f $X=0.665 $Y=1.405 $X2=0
+ $Y2=0
cc_125 N_B1_N_c_123_n N_A_29_392#_c_319_n 0.00736778f $X=0.495 $Y=1.885 $X2=0
+ $Y2=0
cc_126 N_B1_N_c_123_n N_A_29_392#_c_328_n 0.0161899f $X=0.495 $Y=1.885 $X2=0
+ $Y2=0
cc_127 N_B1_N_M1005_g N_A_29_392#_c_313_n 0.00631428f $X=0.665 $Y=0.935 $X2=0
+ $Y2=0
cc_128 N_B1_N_c_119_n N_A_29_392#_c_313_n 0.00826526f $X=0.665 $Y=1.405 $X2=0
+ $Y2=0
cc_129 B1_N N_A_29_392#_c_313_n 0.0288538f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_130 N_B1_N_c_121_n N_A_29_392#_c_313_n 0.00169755f $X=0.665 $Y=0.34 $X2=0
+ $Y2=0
cc_131 N_B1_N_c_123_n N_A_29_392#_c_322_n 2.24111e-19 $X=0.495 $Y=1.885 $X2=0
+ $Y2=0
cc_132 N_B1_N_c_123_n N_VPWR_c_541_n 0.00513915f $X=0.495 $Y=1.885 $X2=0 $Y2=0
cc_133 N_B1_N_c_123_n N_VPWR_c_550_n 0.00445602f $X=0.495 $Y=1.885 $X2=0 $Y2=0
cc_134 N_B1_N_c_123_n N_VPWR_c_540_n 0.0086135f $X=0.495 $Y=1.885 $X2=0 $Y2=0
cc_135 N_B1_N_M1005_g N_X_c_629_n 9.78852e-19 $X=0.665 $Y=0.935 $X2=0 $Y2=0
cc_136 N_B1_N_c_117_n N_X_c_631_n 0.00373183f $X=0.495 $Y=1.795 $X2=0 $Y2=0
cc_137 N_B1_N_c_123_n N_X_c_631_n 0.00147493f $X=0.495 $Y=1.885 $X2=0 $Y2=0
cc_138 N_B1_N_c_119_n N_X_c_631_n 0.00721533f $X=0.665 $Y=1.405 $X2=0 $Y2=0
cc_139 B1_N N_VGND_c_754_n 0.0255983f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_140 N_B1_N_c_121_n N_VGND_c_754_n 0.0135756f $X=0.665 $Y=0.34 $X2=0 $Y2=0
cc_141 B1_N N_VGND_c_762_n 0.0328545f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_142 N_B1_N_c_121_n N_VGND_c_762_n 0.010364f $X=0.665 $Y=0.34 $X2=0 $Y2=0
cc_143 B1_N N_VGND_c_769_n 0.0175703f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_144 N_B1_N_c_121_n N_VGND_c_769_n 0.0170572f $X=0.665 $Y=0.34 $X2=0 $Y2=0
cc_145 N_A_187_338#_c_155_n N_A_29_392#_M1015_g 0.0160601f $X=2.545 $Y=1.35
+ $X2=0 $Y2=0
cc_146 N_A_187_338#_c_157_n N_A_29_392#_M1015_g 0.0106037f $X=3.085 $Y=1.195
+ $X2=0 $Y2=0
cc_147 N_A_187_338#_c_158_n N_A_29_392#_M1015_g 0.008147f $X=3.25 $Y=0.76 $X2=0
+ $Y2=0
cc_148 N_A_187_338#_c_159_n N_A_29_392#_M1015_g 9.01637e-19 $X=3.555 $Y=2.115
+ $X2=0 $Y2=0
cc_149 N_A_187_338#_c_161_n N_A_29_392#_M1015_g 0.00113175f $X=3.72 $Y=1.195
+ $X2=0 $Y2=0
cc_150 N_A_187_338#_c_163_n N_A_29_392#_M1015_g 0.00539532f $X=2.67 $Y=1.195
+ $X2=0 $Y2=0
cc_151 N_A_187_338#_c_159_n N_A_29_392#_c_314_n 0.00652065f $X=3.555 $Y=2.115
+ $X2=0 $Y2=0
cc_152 N_A_187_338#_c_167_n N_A_29_392#_c_308_n 3.7888e-19 $X=2.36 $Y=1.765
+ $X2=0 $Y2=0
cc_153 N_A_187_338#_c_156_n N_A_29_392#_c_308_n 0.0183453f $X=2.435 $Y=1.515
+ $X2=0 $Y2=0
cc_154 N_A_187_338#_c_159_n N_A_29_392#_c_308_n 0.0156825f $X=3.555 $Y=2.115
+ $X2=0 $Y2=0
cc_155 N_A_187_338#_c_161_n N_A_29_392#_c_308_n 0.00816026f $X=3.72 $Y=1.195
+ $X2=0 $Y2=0
cc_156 N_A_187_338#_c_158_n N_A_29_392#_M1021_g 0.0118095f $X=3.25 $Y=0.76 $X2=0
+ $Y2=0
cc_157 N_A_187_338#_c_159_n N_A_29_392#_M1021_g 0.00612122f $X=3.555 $Y=2.115
+ $X2=0 $Y2=0
cc_158 N_A_187_338#_c_161_n N_A_29_392#_M1021_g 0.0152251f $X=3.72 $Y=1.195
+ $X2=0 $Y2=0
cc_159 N_A_187_338#_c_159_n N_A_29_392#_c_310_n 0.00528271f $X=3.555 $Y=2.115
+ $X2=0 $Y2=0
cc_160 N_A_187_338#_c_159_n N_A_29_392#_c_317_n 0.0133621f $X=3.555 $Y=2.115
+ $X2=0 $Y2=0
cc_161 N_A_187_338#_c_164_n N_A_29_392#_c_311_n 7.86349e-19 $X=1.01 $Y=1.765
+ $X2=0 $Y2=0
cc_162 N_A_187_338#_c_156_n N_A_29_392#_c_311_n 0.00109545f $X=2.435 $Y=1.515
+ $X2=0 $Y2=0
cc_163 N_A_187_338#_c_164_n N_A_29_392#_c_319_n 8.09587e-19 $X=1.01 $Y=1.765
+ $X2=0 $Y2=0
cc_164 N_A_187_338#_c_164_n N_A_29_392#_c_328_n 0.0149727f $X=1.01 $Y=1.765
+ $X2=0 $Y2=0
cc_165 N_A_187_338#_c_165_n N_A_29_392#_c_328_n 0.014686f $X=1.46 $Y=1.765 $X2=0
+ $Y2=0
cc_166 N_A_187_338#_c_166_n N_A_29_392#_c_328_n 0.0146364f $X=1.91 $Y=1.765
+ $X2=0 $Y2=0
cc_167 N_A_187_338#_c_167_n N_A_29_392#_c_328_n 0.0174699f $X=2.36 $Y=1.765
+ $X2=0 $Y2=0
cc_168 N_A_187_338#_c_198_p N_A_29_392#_c_328_n 0.00392008f $X=2.585 $Y=1.515
+ $X2=0 $Y2=0
cc_169 N_A_187_338#_c_156_n N_A_29_392#_c_328_n 7.25681e-19 $X=2.435 $Y=1.515
+ $X2=0 $Y2=0
cc_170 N_A_187_338#_c_157_n N_A_29_392#_c_320_n 0.00665025f $X=3.085 $Y=1.195
+ $X2=0 $Y2=0
cc_171 N_A_187_338#_c_159_n N_A_29_392#_c_320_n 0.0132509f $X=3.555 $Y=2.115
+ $X2=0 $Y2=0
cc_172 N_A_187_338#_c_163_n N_A_29_392#_c_320_n 0.00935958f $X=2.67 $Y=1.195
+ $X2=0 $Y2=0
cc_173 N_A_187_338#_c_198_p N_A_29_392#_c_362_n 0.00842244f $X=2.585 $Y=1.515
+ $X2=0 $Y2=0
cc_174 N_A_187_338#_c_156_n N_A_29_392#_c_362_n 0.00336158f $X=2.435 $Y=1.515
+ $X2=0 $Y2=0
cc_175 N_A_187_338#_c_163_n N_A_29_392#_c_362_n 0.00469696f $X=2.67 $Y=1.195
+ $X2=0 $Y2=0
cc_176 N_A_187_338#_c_167_n N_A_29_392#_c_312_n 0.00185317f $X=2.36 $Y=1.765
+ $X2=0 $Y2=0
cc_177 N_A_187_338#_c_156_n N_A_29_392#_c_312_n 6.99374e-19 $X=2.435 $Y=1.515
+ $X2=0 $Y2=0
cc_178 N_A_187_338#_c_157_n N_A_29_392#_c_312_n 0.0252564f $X=3.085 $Y=1.195
+ $X2=0 $Y2=0
cc_179 N_A_187_338#_c_159_n N_A_29_392#_c_312_n 0.0290314f $X=3.555 $Y=2.115
+ $X2=0 $Y2=0
cc_180 N_A_187_338#_c_163_n N_A_29_392#_c_312_n 0.0150195f $X=2.67 $Y=1.195
+ $X2=0 $Y2=0
cc_181 N_A_187_338#_c_160_n N_A1_M1006_g 0.0121855f $X=4.785 $Y=1.195 $X2=0
+ $Y2=0
cc_182 N_A_187_338#_c_162_n N_A1_M1006_g 0.00709401f $X=4.95 $Y=0.76 $X2=0 $Y2=0
cc_183 N_A_187_338#_c_160_n N_A1_M1012_g 3.19858e-19 $X=4.785 $Y=1.195 $X2=0
+ $Y2=0
cc_184 N_A_187_338#_c_160_n A1 0.0466358f $X=4.785 $Y=1.195 $X2=0 $Y2=0
cc_185 N_A_187_338#_c_160_n N_A1_c_423_n 0.00413199f $X=4.785 $Y=1.195 $X2=0
+ $Y2=0
cc_186 N_A_187_338#_c_159_n N_A2_c_467_n 0.00225412f $X=3.555 $Y=2.115 $X2=-0.19
+ $Y2=-0.245
cc_187 N_A_187_338#_c_160_n N_A2_c_467_n 0.00106972f $X=4.785 $Y=1.195 $X2=-0.19
+ $Y2=-0.245
cc_188 N_A_187_338#_c_159_n N_A2_c_468_n 0.00207123f $X=3.555 $Y=2.115 $X2=0
+ $Y2=0
cc_189 N_A_187_338#_c_159_n N_A2_c_477_n 3.18071e-19 $X=3.555 $Y=2.115 $X2=0
+ $Y2=0
cc_190 N_A_187_338#_c_159_n N_A2_M1009_g 9.04115e-19 $X=3.555 $Y=2.115 $X2=0
+ $Y2=0
cc_191 N_A_187_338#_c_160_n N_A2_M1009_g 0.0169245f $X=4.785 $Y=1.195 $X2=0
+ $Y2=0
cc_192 N_A_187_338#_c_162_n N_A2_M1009_g 8.96234e-19 $X=4.95 $Y=0.76 $X2=0 $Y2=0
cc_193 N_A_187_338#_c_162_n N_A2_c_470_n 0.00126713f $X=4.95 $Y=0.76 $X2=0 $Y2=0
cc_194 N_A_187_338#_c_160_n N_A2_c_474_n 8.68147e-19 $X=4.785 $Y=1.195 $X2=0
+ $Y2=0
cc_195 N_A_187_338#_c_160_n N_A2_c_475_n 0.0100199f $X=4.785 $Y=1.195 $X2=0
+ $Y2=0
cc_196 N_A_187_338#_c_164_n N_VPWR_c_541_n 0.010481f $X=1.01 $Y=1.765 $X2=0
+ $Y2=0
cc_197 N_A_187_338#_c_165_n N_VPWR_c_541_n 0.0014191f $X=1.46 $Y=1.765 $X2=0
+ $Y2=0
cc_198 N_A_187_338#_c_164_n N_VPWR_c_542_n 0.0014191f $X=1.01 $Y=1.765 $X2=0
+ $Y2=0
cc_199 N_A_187_338#_c_165_n N_VPWR_c_542_n 0.0105066f $X=1.46 $Y=1.765 $X2=0
+ $Y2=0
cc_200 N_A_187_338#_c_166_n N_VPWR_c_542_n 0.0105066f $X=1.91 $Y=1.765 $X2=0
+ $Y2=0
cc_201 N_A_187_338#_c_167_n N_VPWR_c_542_n 0.0014191f $X=2.36 $Y=1.765 $X2=0
+ $Y2=0
cc_202 N_A_187_338#_c_166_n N_VPWR_c_543_n 0.0014191f $X=1.91 $Y=1.765 $X2=0
+ $Y2=0
cc_203 N_A_187_338#_c_167_n N_VPWR_c_543_n 0.0114975f $X=2.36 $Y=1.765 $X2=0
+ $Y2=0
cc_204 N_A_187_338#_c_164_n N_VPWR_c_551_n 0.00413917f $X=1.01 $Y=1.765 $X2=0
+ $Y2=0
cc_205 N_A_187_338#_c_165_n N_VPWR_c_551_n 0.00413917f $X=1.46 $Y=1.765 $X2=0
+ $Y2=0
cc_206 N_A_187_338#_c_166_n N_VPWR_c_552_n 0.00413917f $X=1.91 $Y=1.765 $X2=0
+ $Y2=0
cc_207 N_A_187_338#_c_167_n N_VPWR_c_552_n 0.00413917f $X=2.36 $Y=1.765 $X2=0
+ $Y2=0
cc_208 N_A_187_338#_c_164_n N_VPWR_c_540_n 0.00817726f $X=1.01 $Y=1.765 $X2=0
+ $Y2=0
cc_209 N_A_187_338#_c_165_n N_VPWR_c_540_n 0.00817726f $X=1.46 $Y=1.765 $X2=0
+ $Y2=0
cc_210 N_A_187_338#_c_166_n N_VPWR_c_540_n 0.00817726f $X=1.91 $Y=1.765 $X2=0
+ $Y2=0
cc_211 N_A_187_338#_c_167_n N_VPWR_c_540_n 0.00817726f $X=2.36 $Y=1.765 $X2=0
+ $Y2=0
cc_212 N_A_187_338#_c_152_n N_X_c_628_n 0.00905582f $X=1.255 $Y=1.35 $X2=0 $Y2=0
cc_213 N_A_187_338#_c_152_n N_X_c_629_n 0.00393613f $X=1.255 $Y=1.35 $X2=0 $Y2=0
cc_214 N_A_187_338#_c_153_n N_X_c_629_n 0.00331437f $X=1.685 $Y=1.35 $X2=0 $Y2=0
cc_215 N_A_187_338#_c_198_p N_X_c_629_n 0.0120778f $X=2.585 $Y=1.515 $X2=0 $Y2=0
cc_216 N_A_187_338#_c_156_n N_X_c_629_n 0.00746874f $X=2.435 $Y=1.515 $X2=0
+ $Y2=0
cc_217 N_A_187_338#_c_165_n N_X_c_642_n 0.0103777f $X=1.46 $Y=1.765 $X2=0 $Y2=0
cc_218 N_A_187_338#_c_166_n N_X_c_642_n 0.010767f $X=1.91 $Y=1.765 $X2=0 $Y2=0
cc_219 N_A_187_338#_c_167_n N_X_c_642_n 0.0028671f $X=2.36 $Y=1.765 $X2=0 $Y2=0
cc_220 N_A_187_338#_c_198_p N_X_c_642_n 0.0468148f $X=2.585 $Y=1.515 $X2=0 $Y2=0
cc_221 N_A_187_338#_c_156_n N_X_c_642_n 0.0139419f $X=2.435 $Y=1.515 $X2=0 $Y2=0
cc_222 N_A_187_338#_c_153_n N_X_c_647_n 0.0120233f $X=1.685 $Y=1.35 $X2=0 $Y2=0
cc_223 N_A_187_338#_c_154_n N_X_c_647_n 0.01168f $X=2.115 $Y=1.35 $X2=0 $Y2=0
cc_224 N_A_187_338#_c_198_p N_X_c_647_n 0.0547785f $X=2.585 $Y=1.515 $X2=0 $Y2=0
cc_225 N_A_187_338#_c_156_n N_X_c_647_n 0.00534379f $X=2.435 $Y=1.515 $X2=0
+ $Y2=0
cc_226 N_A_187_338#_c_153_n N_X_c_630_n 6.0186e-19 $X=1.685 $Y=1.35 $X2=0 $Y2=0
cc_227 N_A_187_338#_c_154_n N_X_c_630_n 0.00736569f $X=2.115 $Y=1.35 $X2=0 $Y2=0
cc_228 N_A_187_338#_c_152_n N_X_c_653_n 0.00253172f $X=1.255 $Y=1.35 $X2=0 $Y2=0
cc_229 N_A_187_338#_c_156_n N_X_c_653_n 0.00340569f $X=2.435 $Y=1.515 $X2=0
+ $Y2=0
cc_230 N_A_187_338#_c_164_n N_X_c_631_n 0.0119494f $X=1.01 $Y=1.765 $X2=0 $Y2=0
cc_231 N_A_187_338#_c_156_n N_X_c_631_n 0.0247194f $X=2.435 $Y=1.515 $X2=0 $Y2=0
cc_232 N_A_187_338#_c_165_n N_X_c_657_n 0.00397284f $X=1.46 $Y=1.765 $X2=0 $Y2=0
cc_233 N_A_187_338#_c_166_n N_X_c_657_n 4.10023e-19 $X=1.91 $Y=1.765 $X2=0 $Y2=0
cc_234 N_A_187_338#_c_198_p N_X_c_657_n 0.014306f $X=2.585 $Y=1.515 $X2=0 $Y2=0
cc_235 N_A_187_338#_c_156_n N_X_c_657_n 0.0113643f $X=2.435 $Y=1.515 $X2=0 $Y2=0
cc_236 N_A_187_338#_c_167_n N_A_596_392#_c_683_n 0.00507436f $X=2.36 $Y=1.765
+ $X2=0 $Y2=0
cc_237 N_A_187_338#_c_159_n N_A_596_392#_c_683_n 0.0365429f $X=3.555 $Y=2.115
+ $X2=0 $Y2=0
cc_238 N_A_187_338#_M1014_d N_A_596_392#_c_684_n 0.00222494f $X=3.405 $Y=1.96
+ $X2=0 $Y2=0
cc_239 N_A_187_338#_c_159_n N_A_596_392#_c_684_n 0.0144323f $X=3.555 $Y=2.115
+ $X2=0 $Y2=0
cc_240 N_A_187_338#_c_167_n N_A_596_392#_c_685_n 5.75404e-19 $X=2.36 $Y=1.765
+ $X2=0 $Y2=0
cc_241 N_A_187_338#_c_159_n N_A_596_392#_c_686_n 0.0128198f $X=3.555 $Y=2.115
+ $X2=0 $Y2=0
cc_242 N_A_187_338#_c_160_n N_A_596_392#_c_686_n 0.00555366f $X=4.785 $Y=1.195
+ $X2=0 $Y2=0
cc_243 N_A_187_338#_c_159_n N_A_596_392#_c_700_n 0.039183f $X=3.555 $Y=2.115
+ $X2=0 $Y2=0
cc_244 N_A_187_338#_c_160_n N_A_596_392#_c_687_n 0.00911997f $X=4.785 $Y=1.195
+ $X2=0 $Y2=0
cc_245 N_A_187_338#_c_157_n N_VGND_M1010_s 0.00354182f $X=3.085 $Y=1.195 $X2=0
+ $Y2=0
cc_246 N_A_187_338#_c_163_n N_VGND_M1010_s 0.00119952f $X=2.67 $Y=1.195 $X2=0
+ $Y2=0
cc_247 N_A_187_338#_c_160_n N_VGND_M1021_d 0.0117991f $X=4.785 $Y=1.195 $X2=0
+ $Y2=0
cc_248 N_A_187_338#_c_161_n N_VGND_M1021_d 0.00130751f $X=3.72 $Y=1.195 $X2=0
+ $Y2=0
cc_249 N_A_187_338#_c_152_n N_VGND_c_754_n 0.00937327f $X=1.255 $Y=1.35 $X2=0
+ $Y2=0
cc_250 N_A_187_338#_c_156_n N_VGND_c_754_n 0.00306734f $X=2.435 $Y=1.515 $X2=0
+ $Y2=0
cc_251 N_A_187_338#_c_152_n N_VGND_c_755_n 6.55754e-19 $X=1.255 $Y=1.35 $X2=0
+ $Y2=0
cc_252 N_A_187_338#_c_153_n N_VGND_c_755_n 0.00771743f $X=1.685 $Y=1.35 $X2=0
+ $Y2=0
cc_253 N_A_187_338#_c_154_n N_VGND_c_755_n 0.00159705f $X=2.115 $Y=1.35 $X2=0
+ $Y2=0
cc_254 N_A_187_338#_c_154_n N_VGND_c_756_n 0.00467453f $X=2.115 $Y=1.35 $X2=0
+ $Y2=0
cc_255 N_A_187_338#_c_155_n N_VGND_c_756_n 0.00405273f $X=2.545 $Y=1.35 $X2=0
+ $Y2=0
cc_256 N_A_187_338#_c_154_n N_VGND_c_757_n 4.82422e-19 $X=2.115 $Y=1.35 $X2=0
+ $Y2=0
cc_257 N_A_187_338#_c_155_n N_VGND_c_757_n 0.0108453f $X=2.545 $Y=1.35 $X2=0
+ $Y2=0
cc_258 N_A_187_338#_c_157_n N_VGND_c_757_n 0.00724091f $X=3.085 $Y=1.195 $X2=0
+ $Y2=0
cc_259 N_A_187_338#_c_158_n N_VGND_c_757_n 0.0201182f $X=3.25 $Y=0.76 $X2=0
+ $Y2=0
cc_260 N_A_187_338#_c_163_n N_VGND_c_757_n 0.00881517f $X=2.67 $Y=1.195 $X2=0
+ $Y2=0
cc_261 N_A_187_338#_c_158_n N_VGND_c_758_n 0.00697494f $X=3.25 $Y=0.76 $X2=0
+ $Y2=0
cc_262 N_A_187_338#_c_158_n N_VGND_c_759_n 0.0130518f $X=3.25 $Y=0.76 $X2=0
+ $Y2=0
cc_263 N_A_187_338#_c_161_n N_VGND_c_759_n 0.0135504f $X=3.72 $Y=1.195 $X2=0
+ $Y2=0
cc_264 N_A_187_338#_c_152_n N_VGND_c_764_n 0.00421137f $X=1.255 $Y=1.35 $X2=0
+ $Y2=0
cc_265 N_A_187_338#_c_153_n N_VGND_c_764_n 0.00405273f $X=1.685 $Y=1.35 $X2=0
+ $Y2=0
cc_266 N_A_187_338#_c_152_n N_VGND_c_769_n 0.00505379f $X=1.255 $Y=1.35 $X2=0
+ $Y2=0
cc_267 N_A_187_338#_c_153_n N_VGND_c_769_n 0.00424518f $X=1.685 $Y=1.35 $X2=0
+ $Y2=0
cc_268 N_A_187_338#_c_154_n N_VGND_c_769_n 0.00505379f $X=2.115 $Y=1.35 $X2=0
+ $Y2=0
cc_269 N_A_187_338#_c_155_n N_VGND_c_769_n 0.00424518f $X=2.545 $Y=1.35 $X2=0
+ $Y2=0
cc_270 N_A_187_338#_c_158_n N_VGND_c_769_n 0.0100676f $X=3.25 $Y=0.76 $X2=0
+ $Y2=0
cc_271 N_A_187_338#_c_160_n N_A_864_123#_M1009_s 0.00402642f $X=4.785 $Y=1.195
+ $X2=-0.19 $Y2=-0.245
cc_272 N_A_187_338#_c_160_n N_A_864_123#_c_841_n 0.013595f $X=4.785 $Y=1.195
+ $X2=0 $Y2=0
cc_273 N_A_187_338#_c_162_n N_A_864_123#_c_841_n 0.0125368f $X=4.95 $Y=0.76
+ $X2=0 $Y2=0
cc_274 N_A_187_338#_c_162_n N_A_864_123#_c_842_n 0.0195074f $X=4.95 $Y=0.76
+ $X2=0 $Y2=0
cc_275 N_A_187_338#_c_160_n N_A_864_123#_c_844_n 0.00679079f $X=4.785 $Y=1.195
+ $X2=0 $Y2=0
cc_276 N_A_187_338#_c_162_n N_A_864_123#_c_844_n 0.0191862f $X=4.95 $Y=0.76
+ $X2=0 $Y2=0
cc_277 N_A_29_392#_M1021_g N_A2_c_467_n 0.00162326f $X=3.465 $Y=0.935 $X2=-0.19
+ $Y2=-0.245
cc_278 N_A_29_392#_c_308_n N_A2_c_468_n 0.0104141f $X=3.465 $Y=1.45 $X2=0 $Y2=0
cc_279 N_A_29_392#_c_310_n N_A2_c_477_n 0.0104141f $X=3.78 $Y=1.795 $X2=0 $Y2=0
cc_280 N_A_29_392#_c_317_n N_A2_c_477_n 0.00782861f $X=3.78 $Y=1.885 $X2=0 $Y2=0
cc_281 N_A_29_392#_M1021_g N_A2_M1009_g 0.00962689f $X=3.465 $Y=0.935 $X2=0
+ $Y2=0
cc_282 N_A_29_392#_M1021_g N_A2_c_474_n 4.60391e-19 $X=3.465 $Y=0.935 $X2=0
+ $Y2=0
cc_283 N_A_29_392#_c_328_n N_VPWR_M1018_d 0.00538936f $X=2.47 $Y=2.355 $X2=-0.19
+ $Y2=-0.245
cc_284 N_A_29_392#_c_328_n N_VPWR_M1007_s 0.00378491f $X=2.47 $Y=2.355 $X2=0
+ $Y2=0
cc_285 N_A_29_392#_c_328_n N_VPWR_M1013_s 0.00408194f $X=2.47 $Y=2.355 $X2=0
+ $Y2=0
cc_286 N_A_29_392#_c_379_p N_VPWR_M1013_s 0.00466061f $X=2.555 $Y=2.27 $X2=0
+ $Y2=0
cc_287 N_A_29_392#_c_320_n N_VPWR_M1013_s 0.00270092f $X=2.96 $Y=1.935 $X2=0
+ $Y2=0
cc_288 N_A_29_392#_c_362_n N_VPWR_M1013_s 0.00263202f $X=2.64 $Y=1.935 $X2=0
+ $Y2=0
cc_289 N_A_29_392#_c_319_n N_VPWR_c_541_n 0.0137183f $X=0.27 $Y=2.815 $X2=0
+ $Y2=0
cc_290 N_A_29_392#_c_328_n N_VPWR_c_541_n 0.0214453f $X=2.47 $Y=2.355 $X2=0
+ $Y2=0
cc_291 N_A_29_392#_c_328_n N_VPWR_c_542_n 0.0171814f $X=2.47 $Y=2.355 $X2=0
+ $Y2=0
cc_292 N_A_29_392#_c_314_n N_VPWR_c_543_n 0.00133712f $X=3.33 $Y=1.885 $X2=0
+ $Y2=0
cc_293 N_A_29_392#_c_328_n N_VPWR_c_543_n 0.0142293f $X=2.47 $Y=2.355 $X2=0
+ $Y2=0
cc_294 N_A_29_392#_c_320_n N_VPWR_c_543_n 0.00361115f $X=2.96 $Y=1.935 $X2=0
+ $Y2=0
cc_295 N_A_29_392#_c_314_n N_VPWR_c_546_n 0.00278257f $X=3.33 $Y=1.885 $X2=0
+ $Y2=0
cc_296 N_A_29_392#_c_317_n N_VPWR_c_546_n 0.00278271f $X=3.78 $Y=1.885 $X2=0
+ $Y2=0
cc_297 N_A_29_392#_c_319_n N_VPWR_c_550_n 0.0145938f $X=0.27 $Y=2.815 $X2=0
+ $Y2=0
cc_298 N_A_29_392#_c_314_n N_VPWR_c_540_n 0.00358623f $X=3.33 $Y=1.885 $X2=0
+ $Y2=0
cc_299 N_A_29_392#_c_317_n N_VPWR_c_540_n 0.00353907f $X=3.78 $Y=1.885 $X2=0
+ $Y2=0
cc_300 N_A_29_392#_c_319_n N_VPWR_c_540_n 0.0120466f $X=0.27 $Y=2.815 $X2=0
+ $Y2=0
cc_301 N_A_29_392#_c_328_n N_X_M1004_d 0.00890288f $X=2.47 $Y=2.355 $X2=0 $Y2=0
cc_302 N_A_29_392#_c_328_n N_X_M1011_d 0.00890462f $X=2.47 $Y=2.355 $X2=0 $Y2=0
cc_303 N_A_29_392#_c_328_n N_X_c_642_n 0.047273f $X=2.47 $Y=2.355 $X2=0 $Y2=0
cc_304 N_A_29_392#_c_311_n N_X_c_631_n 0.0429777f $X=0.27 $Y=2.105 $X2=0 $Y2=0
cc_305 N_A_29_392#_c_328_n N_X_c_631_n 0.0398874f $X=2.47 $Y=2.355 $X2=0 $Y2=0
cc_306 N_A_29_392#_c_313_n N_X_c_631_n 6.64223e-19 $X=0.45 $Y=1.055 $X2=0 $Y2=0
cc_307 N_A_29_392#_c_328_n N_X_c_657_n 0.00896998f $X=2.47 $Y=2.355 $X2=0 $Y2=0
cc_308 N_A_29_392#_c_320_n N_A_596_392#_M1014_s 0.00266517f $X=2.96 $Y=1.935
+ $X2=-0.19 $Y2=-0.245
cc_309 N_A_29_392#_c_314_n N_A_596_392#_c_683_n 0.0103116f $X=3.33 $Y=1.885
+ $X2=0 $Y2=0
cc_310 N_A_29_392#_c_308_n N_A_596_392#_c_683_n 0.00119613f $X=3.465 $Y=1.45
+ $X2=0 $Y2=0
cc_311 N_A_29_392#_c_317_n N_A_596_392#_c_683_n 6.4534e-19 $X=3.78 $Y=1.885
+ $X2=0 $Y2=0
cc_312 N_A_29_392#_c_328_n N_A_596_392#_c_683_n 0.0097999f $X=2.47 $Y=2.355
+ $X2=0 $Y2=0
cc_313 N_A_29_392#_c_379_p N_A_596_392#_c_683_n 0.00413595f $X=2.555 $Y=2.27
+ $X2=0 $Y2=0
cc_314 N_A_29_392#_c_320_n N_A_596_392#_c_683_n 0.023946f $X=2.96 $Y=1.935 $X2=0
+ $Y2=0
cc_315 N_A_29_392#_c_314_n N_A_596_392#_c_684_n 0.0107904f $X=3.33 $Y=1.885
+ $X2=0 $Y2=0
cc_316 N_A_29_392#_c_317_n N_A_596_392#_c_684_n 0.012504f $X=3.78 $Y=1.885 $X2=0
+ $Y2=0
cc_317 N_A_29_392#_c_314_n N_A_596_392#_c_685_n 0.00262934f $X=3.33 $Y=1.885
+ $X2=0 $Y2=0
cc_318 N_A_29_392#_c_317_n N_A_596_392#_c_686_n 8.64891e-19 $X=3.78 $Y=1.885
+ $X2=0 $Y2=0
cc_319 N_A_29_392#_c_313_n N_VGND_c_754_n 0.0173641f $X=0.45 $Y=1.055 $X2=0
+ $Y2=0
cc_320 N_A_29_392#_M1015_g N_VGND_c_757_n 0.00548634f $X=3.035 $Y=0.935 $X2=0
+ $Y2=0
cc_321 N_A_29_392#_M1015_g N_VGND_c_758_n 0.00404905f $X=3.035 $Y=0.935 $X2=0
+ $Y2=0
cc_322 N_A_29_392#_M1021_g N_VGND_c_758_n 0.00404905f $X=3.465 $Y=0.935 $X2=0
+ $Y2=0
cc_323 N_A_29_392#_M1021_g N_VGND_c_759_n 0.00323233f $X=3.465 $Y=0.935 $X2=0
+ $Y2=0
cc_324 N_A_29_392#_M1015_g N_VGND_c_769_n 0.00472204f $X=3.035 $Y=0.935 $X2=0
+ $Y2=0
cc_325 N_A_29_392#_M1021_g N_VGND_c_769_n 0.00472204f $X=3.465 $Y=0.935 $X2=0
+ $Y2=0
cc_326 N_A_29_392#_c_313_n N_VGND_c_769_n 0.00195038f $X=0.45 $Y=1.055 $X2=0
+ $Y2=0
cc_327 A1 N_A2_c_468_n 0.00954291f $X=4.955 $Y=1.58 $X2=0 $Y2=0
cc_328 N_A1_c_423_n N_A2_c_468_n 0.0199126f $X=5.13 $Y=1.667 $X2=0 $Y2=0
cc_329 N_A1_c_424_n N_A2_c_477_n 0.0201493f $X=4.68 $Y=1.885 $X2=0 $Y2=0
cc_330 N_A1_M1006_g N_A2_c_470_n 0.00977419f $X=4.735 $Y=0.935 $X2=0 $Y2=0
cc_331 N_A1_M1012_g N_A2_c_470_n 0.00977211f $X=5.165 $Y=0.935 $X2=0 $Y2=0
cc_332 N_A1_M1012_g N_A2_c_471_n 0.00774781f $X=5.165 $Y=0.935 $X2=0 $Y2=0
cc_333 A1 N_A2_c_472_n 0.00197413f $X=4.955 $Y=1.58 $X2=0 $Y2=0
cc_334 N_A1_c_423_n N_A2_c_472_n 0.0229759f $X=5.13 $Y=1.667 $X2=0 $Y2=0
cc_335 N_A1_c_425_n N_A2_c_479_n 0.0201493f $X=5.13 $Y=1.885 $X2=0 $Y2=0
cc_336 N_A1_M1012_g N_A2_M1020_g 0.00949913f $X=5.165 $Y=0.935 $X2=0 $Y2=0
cc_337 N_A1_M1006_g N_A2_c_474_n 0.0269452f $X=4.735 $Y=0.935 $X2=0 $Y2=0
cc_338 N_A1_c_424_n N_VPWR_c_544_n 0.00526215f $X=4.68 $Y=1.885 $X2=0 $Y2=0
cc_339 N_A1_c_425_n N_VPWR_c_545_n 0.00526215f $X=5.13 $Y=1.885 $X2=0 $Y2=0
cc_340 N_A1_c_424_n N_VPWR_c_548_n 0.00445602f $X=4.68 $Y=1.885 $X2=0 $Y2=0
cc_341 N_A1_c_425_n N_VPWR_c_548_n 0.00445602f $X=5.13 $Y=1.885 $X2=0 $Y2=0
cc_342 N_A1_c_424_n N_VPWR_c_540_n 0.00857673f $X=4.68 $Y=1.885 $X2=0 $Y2=0
cc_343 N_A1_c_425_n N_VPWR_c_540_n 0.00857673f $X=5.13 $Y=1.885 $X2=0 $Y2=0
cc_344 N_A1_c_424_n N_A_596_392#_c_687_n 0.0119563f $X=4.68 $Y=1.885 $X2=0 $Y2=0
cc_345 A1 N_A_596_392#_c_687_n 0.0222304f $X=4.955 $Y=1.58 $X2=0 $Y2=0
cc_346 N_A1_c_423_n N_A_596_392#_c_687_n 4.03117e-19 $X=5.13 $Y=1.667 $X2=0
+ $Y2=0
cc_347 N_A1_c_424_n N_A_596_392#_c_688_n 0.0105452f $X=4.68 $Y=1.885 $X2=0 $Y2=0
cc_348 N_A1_c_425_n N_A_596_392#_c_688_n 0.0105452f $X=5.13 $Y=1.885 $X2=0 $Y2=0
cc_349 N_A1_c_425_n N_A_596_392#_c_689_n 0.012109f $X=5.13 $Y=1.885 $X2=0 $Y2=0
cc_350 A1 N_A_596_392#_c_689_n 0.00924974f $X=4.955 $Y=1.58 $X2=0 $Y2=0
cc_351 N_A1_c_423_n N_A_596_392#_c_689_n 0.00115835f $X=5.13 $Y=1.667 $X2=0
+ $Y2=0
cc_352 N_A1_c_424_n N_A_596_392#_c_692_n 5.56417e-19 $X=4.68 $Y=1.885 $X2=0
+ $Y2=0
cc_353 N_A1_c_425_n N_A_596_392#_c_692_n 5.56417e-19 $X=5.13 $Y=1.885 $X2=0
+ $Y2=0
cc_354 A1 N_A_596_392#_c_692_n 0.0276944f $X=4.955 $Y=1.58 $X2=0 $Y2=0
cc_355 N_A1_c_423_n N_A_596_392#_c_692_n 0.0078875f $X=5.13 $Y=1.667 $X2=0 $Y2=0
cc_356 N_A1_M1006_g N_A_864_123#_c_841_n 0.00160839f $X=4.735 $Y=0.935 $X2=0
+ $Y2=0
cc_357 N_A1_M1006_g N_A_864_123#_c_842_n 0.00321922f $X=4.735 $Y=0.935 $X2=0
+ $Y2=0
cc_358 N_A1_M1012_g N_A_864_123#_c_842_n 0.00299942f $X=5.165 $Y=0.935 $X2=0
+ $Y2=0
cc_359 N_A1_M1006_g N_A_864_123#_c_844_n 5.55256e-19 $X=4.735 $Y=0.935 $X2=0
+ $Y2=0
cc_360 N_A1_M1012_g N_A_864_123#_c_844_n 0.0115123f $X=5.165 $Y=0.935 $X2=0
+ $Y2=0
cc_361 N_A2_c_477_n N_VPWR_c_544_n 0.00996098f $X=4.23 $Y=1.885 $X2=0 $Y2=0
cc_362 N_A2_c_479_n N_VPWR_c_545_n 0.0135832f $X=5.58 $Y=1.885 $X2=0 $Y2=0
cc_363 N_A2_c_477_n N_VPWR_c_546_n 0.00413917f $X=4.23 $Y=1.885 $X2=0 $Y2=0
cc_364 N_A2_c_479_n N_VPWR_c_553_n 0.00413917f $X=5.58 $Y=1.885 $X2=0 $Y2=0
cc_365 N_A2_c_477_n N_VPWR_c_540_n 0.0081781f $X=4.23 $Y=1.885 $X2=0 $Y2=0
cc_366 N_A2_c_479_n N_VPWR_c_540_n 0.00821632f $X=5.58 $Y=1.885 $X2=0 $Y2=0
cc_367 N_A2_c_477_n N_A_596_392#_c_684_n 0.00125031f $X=4.23 $Y=1.885 $X2=0
+ $Y2=0
cc_368 N_A2_c_477_n N_A_596_392#_c_686_n 2.39049e-19 $X=4.23 $Y=1.885 $X2=0
+ $Y2=0
cc_369 N_A2_c_477_n N_A_596_392#_c_687_n 0.0160233f $X=4.23 $Y=1.885 $X2=0 $Y2=0
cc_370 N_A2_c_477_n N_A_596_392#_c_688_n 6.69308e-19 $X=4.23 $Y=1.885 $X2=0
+ $Y2=0
cc_371 N_A2_c_479_n N_A_596_392#_c_688_n 6.69308e-19 $X=5.58 $Y=1.885 $X2=0
+ $Y2=0
cc_372 N_A2_c_479_n N_A_596_392#_c_689_n 0.0179777f $X=5.58 $Y=1.885 $X2=0 $Y2=0
cc_373 N_A2_c_479_n N_A_596_392#_c_690_n 4.02768e-19 $X=5.58 $Y=1.885 $X2=0
+ $Y2=0
cc_374 N_A2_c_479_n N_A_596_392#_c_691_n 0.0043207f $X=5.58 $Y=1.885 $X2=0 $Y2=0
cc_375 N_A2_c_475_n N_VGND_M1021_d 0.00358673f $X=4.1 $Y=0.34 $X2=0 $Y2=0
cc_376 N_A2_M1009_g N_VGND_c_759_n 0.00283851f $X=4.245 $Y=0.935 $X2=0 $Y2=0
cc_377 N_A2_c_474_n N_VGND_c_759_n 0.0095538f $X=4.127 $Y=0.2 $X2=0 $Y2=0
cc_378 N_A2_c_475_n N_VGND_c_759_n 0.0317133f $X=4.1 $Y=0.34 $X2=0 $Y2=0
cc_379 N_A2_c_470_n N_VGND_c_761_n 0.0136213f $X=5.52 $Y=0.2 $X2=0 $Y2=0
cc_380 N_A2_c_474_n N_VGND_c_766_n 0.0401489f $X=4.127 $Y=0.2 $X2=0 $Y2=0
cc_381 N_A2_c_475_n N_VGND_c_766_n 0.0215843f $X=4.1 $Y=0.34 $X2=0 $Y2=0
cc_382 N_A2_c_470_n N_VGND_c_769_n 0.0424251f $X=5.52 $Y=0.2 $X2=0 $Y2=0
cc_383 N_A2_c_474_n N_VGND_c_769_n 0.0133751f $X=4.127 $Y=0.2 $X2=0 $Y2=0
cc_384 N_A2_c_475_n N_VGND_c_769_n 0.0110944f $X=4.1 $Y=0.34 $X2=0 $Y2=0
cc_385 N_A2_c_474_n N_A_864_123#_c_841_n 0.00608522f $X=4.127 $Y=0.2 $X2=0 $Y2=0
cc_386 N_A2_c_475_n N_A_864_123#_c_841_n 0.0182646f $X=4.1 $Y=0.34 $X2=0 $Y2=0
cc_387 N_A2_c_470_n N_A_864_123#_c_842_n 0.0216348f $X=5.52 $Y=0.2 $X2=0 $Y2=0
cc_388 N_A2_M1020_g N_A_864_123#_c_842_n 0.00523557f $X=5.595 $Y=0.935 $X2=0
+ $Y2=0
cc_389 N_A2_c_470_n N_A_864_123#_c_843_n 0.00594104f $X=5.52 $Y=0.2 $X2=0 $Y2=0
cc_390 N_A2_c_474_n N_A_864_123#_c_843_n 0.00385041f $X=4.127 $Y=0.2 $X2=0 $Y2=0
cc_391 N_A2_c_475_n N_A_864_123#_c_843_n 0.0142455f $X=4.1 $Y=0.34 $X2=0 $Y2=0
cc_392 N_A2_c_471_n N_A_864_123#_c_844_n 0.00117013f $X=5.58 $Y=1.42 $X2=0 $Y2=0
cc_393 N_A2_M1020_g N_A_864_123#_c_844_n 0.0129429f $X=5.595 $Y=0.935 $X2=0
+ $Y2=0
cc_394 N_VPWR_M1007_s N_X_c_642_n 0.00358101f $X=1.535 $Y=1.84 $X2=0 $Y2=0
cc_395 N_VPWR_M1018_d N_X_c_631_n 0.00434025f $X=0.57 $Y=1.96 $X2=0 $Y2=0
cc_396 N_VPWR_c_543_n N_A_596_392#_c_683_n 0.0226773f $X=2.585 $Y=2.775 $X2=0
+ $Y2=0
cc_397 N_VPWR_c_544_n N_A_596_392#_c_684_n 0.0123543f $X=4.455 $Y=2.455 $X2=0
+ $Y2=0
cc_398 N_VPWR_c_546_n N_A_596_392#_c_684_n 0.0531736f $X=4.29 $Y=3.33 $X2=0
+ $Y2=0
cc_399 N_VPWR_c_540_n N_A_596_392#_c_684_n 0.0297434f $X=6 $Y=3.33 $X2=0 $Y2=0
cc_400 N_VPWR_c_543_n N_A_596_392#_c_685_n 0.0139f $X=2.585 $Y=2.775 $X2=0 $Y2=0
cc_401 N_VPWR_c_546_n N_A_596_392#_c_685_n 0.0236039f $X=4.29 $Y=3.33 $X2=0
+ $Y2=0
cc_402 N_VPWR_c_540_n N_A_596_392#_c_685_n 0.012761f $X=6 $Y=3.33 $X2=0 $Y2=0
cc_403 N_VPWR_c_544_n N_A_596_392#_c_700_n 0.039183f $X=4.455 $Y=2.455 $X2=0
+ $Y2=0
cc_404 N_VPWR_M1002_s N_A_596_392#_c_687_n 0.00222494f $X=4.305 $Y=1.96 $X2=0
+ $Y2=0
cc_405 N_VPWR_c_544_n N_A_596_392#_c_687_n 0.0154248f $X=4.455 $Y=2.455 $X2=0
+ $Y2=0
cc_406 N_VPWR_c_544_n N_A_596_392#_c_688_n 0.0462948f $X=4.455 $Y=2.455 $X2=0
+ $Y2=0
cc_407 N_VPWR_c_545_n N_A_596_392#_c_688_n 0.0462948f $X=5.355 $Y=2.455 $X2=0
+ $Y2=0
cc_408 N_VPWR_c_548_n N_A_596_392#_c_688_n 0.014552f $X=5.27 $Y=3.33 $X2=0 $Y2=0
cc_409 N_VPWR_c_540_n N_A_596_392#_c_688_n 0.0119791f $X=6 $Y=3.33 $X2=0 $Y2=0
cc_410 N_VPWR_M1019_d N_A_596_392#_c_689_n 0.00222494f $X=5.205 $Y=1.96 $X2=0
+ $Y2=0
cc_411 N_VPWR_c_545_n N_A_596_392#_c_689_n 0.0154248f $X=5.355 $Y=2.455 $X2=0
+ $Y2=0
cc_412 N_VPWR_c_545_n N_A_596_392#_c_691_n 0.0453479f $X=5.355 $Y=2.455 $X2=0
+ $Y2=0
cc_413 N_VPWR_c_553_n N_A_596_392#_c_691_n 0.011066f $X=6 $Y=3.33 $X2=0 $Y2=0
cc_414 N_VPWR_c_540_n N_A_596_392#_c_691_n 0.00915947f $X=6 $Y=3.33 $X2=0 $Y2=0
cc_415 N_X_c_647_n N_VGND_M1003_s 0.00330483f $X=2.165 $Y=1.095 $X2=0 $Y2=0
cc_416 N_X_c_628_n N_VGND_c_754_n 0.0346633f $X=1.47 $Y=0.645 $X2=0 $Y2=0
cc_417 N_X_c_629_n N_VGND_c_754_n 0.00595397f $X=1.335 $Y=1.51 $X2=0 $Y2=0
cc_418 N_X_c_653_n N_VGND_c_754_n 0.0118739f $X=1.402 $Y=1.095 $X2=0 $Y2=0
cc_419 N_X_c_631_n N_VGND_c_754_n 0.0177997f $X=1.25 $Y=1.805 $X2=0 $Y2=0
cc_420 N_X_c_628_n N_VGND_c_755_n 0.0131157f $X=1.47 $Y=0.645 $X2=0 $Y2=0
cc_421 N_X_c_647_n N_VGND_c_755_n 0.0152916f $X=2.165 $Y=1.095 $X2=0 $Y2=0
cc_422 N_X_c_630_n N_VGND_c_755_n 0.0130934f $X=2.33 $Y=0.645 $X2=0 $Y2=0
cc_423 N_X_c_630_n N_VGND_c_756_n 0.00718756f $X=2.33 $Y=0.645 $X2=0 $Y2=0
cc_424 N_X_c_630_n N_VGND_c_757_n 0.0165282f $X=2.33 $Y=0.645 $X2=0 $Y2=0
cc_425 N_X_c_628_n N_VGND_c_764_n 0.00864478f $X=1.47 $Y=0.645 $X2=0 $Y2=0
cc_426 N_X_c_628_n N_VGND_c_769_n 0.0102032f $X=1.47 $Y=0.645 $X2=0 $Y2=0
cc_427 N_X_c_630_n N_VGND_c_769_n 0.0083989f $X=2.33 $Y=0.645 $X2=0 $Y2=0
cc_428 N_A_596_392#_c_690_n N_VGND_c_761_n 0.00876636f $X=5.845 $Y=2.12 $X2=0
+ $Y2=0
cc_429 N_A_596_392#_c_689_n N_A_864_123#_c_844_n 0.0101583f $X=5.72 $Y=2.035
+ $X2=0 $Y2=0
cc_430 N_VGND_c_759_n N_A_864_123#_c_841_n 0.00693182f $X=3.68 $Y=0.775 $X2=0
+ $Y2=0
cc_431 N_VGND_c_761_n N_A_864_123#_c_842_n 0.0133372f $X=5.81 $Y=0.76 $X2=0
+ $Y2=0
cc_432 N_VGND_c_766_n N_A_864_123#_c_842_n 0.0599312f $X=5.725 $Y=0 $X2=0 $Y2=0
cc_433 N_VGND_c_769_n N_A_864_123#_c_842_n 0.0314373f $X=6 $Y=0 $X2=0 $Y2=0
cc_434 N_VGND_c_766_n N_A_864_123#_c_843_n 0.0115954f $X=5.725 $Y=0 $X2=0 $Y2=0
cc_435 N_VGND_c_769_n N_A_864_123#_c_843_n 0.00583261f $X=6 $Y=0 $X2=0 $Y2=0
cc_436 N_VGND_c_761_n N_A_864_123#_c_844_n 0.0383986f $X=5.81 $Y=0.76 $X2=0
+ $Y2=0
