* File: sky130_fd_sc_hs__and4bb_4.pex.spice
* Created: Tue Sep  1 19:56:31 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HS__AND4BB_4%B_N 3 5 7 8 9
r27 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.405
+ $Y=1.615 $X2=0.405 $Y2=1.615
r28 9 14 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=0.72 $Y=1.615
+ $X2=0.405 $Y2=1.615
r29 8 14 5.76222 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=0.24 $Y=1.615
+ $X2=0.405 $Y2=1.615
r30 5 13 56.0674 $w=2.9e-07 $l=3.13927e-07 $layer=POLY_cond $X=0.505 $Y=1.885
+ $X2=0.41 $Y2=1.615
r31 5 7 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=0.505 $Y=1.885
+ $X2=0.505 $Y2=2.46
r32 1 13 38.6157 $w=2.9e-07 $l=2.03101e-07 $layer=POLY_cond $X=0.495 $Y=1.45
+ $X2=0.41 $Y2=1.615
r33 1 3 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=0.495 $Y=1.45
+ $X2=0.495 $Y2=0.69
.ends

.subckt PM_SKY130_FD_SC_HS__AND4BB_4%A_N 3 5 7 8
r29 8 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.17
+ $Y=1.615 $X2=1.17 $Y2=1.615
r30 5 11 52.1213 $w=4.11e-07 $l=2.87906e-07 $layer=POLY_cond $X=1.055 $Y=1.885
+ $X2=1.092 $Y2=1.615
r31 5 7 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=1.055 $Y=1.885
+ $X2=1.055 $Y2=2.46
r32 1 11 39.8074 $w=4.11e-07 $l=2.35465e-07 $layer=POLY_cond $X=0.925 $Y=1.45
+ $X2=1.092 $Y2=1.615
r33 1 3 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=0.925 $Y=1.45
+ $X2=0.925 $Y2=0.69
.ends

.subckt PM_SKY130_FD_SC_HS__AND4BB_4%A_200_74# 1 2 7 9 11 12 14 15 17 21 24 28
+ 32 37 38 45
c92 32 0 6.58453e-20 $X=1.525 $Y=0.42
c93 21 0 9.745e-20 $X=2.92 $Y=1.02
r94 45 46 1.8634 $w=3.88e-07 $l=1.5e-08 $layer=POLY_cond $X=2.905 $Y=1.642
+ $X2=2.92 $Y2=1.642
r95 44 45 51.5541 $w=3.88e-07 $l=4.15e-07 $layer=POLY_cond $X=2.49 $Y=1.642
+ $X2=2.905 $Y2=1.642
r96 43 44 25.4665 $w=3.88e-07 $l=2.05e-07 $layer=POLY_cond $X=2.285 $Y=1.642
+ $X2=2.49 $Y2=1.642
r97 33 38 28.8521 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.525 $Y=0.42
+ $X2=1.525 $Y2=0.255
r98 32 35 9.44306 $w=5.62e-07 $l=4.35e-07 $layer=LI1_cond $X=1.367 $Y=0.42
+ $X2=1.367 $Y2=0.855
r99 32 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.525
+ $Y=0.42 $X2=1.525 $Y2=0.42
r100 29 43 23.6031 $w=3.88e-07 $l=1.9e-07 $layer=POLY_cond $X=2.095 $Y=1.642
+ $X2=2.285 $Y2=1.642
r101 28 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.095
+ $Y=1.615 $X2=2.095 $Y2=1.615
r102 26 28 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=2.095 $Y=2.29
+ $X2=2.095 $Y2=1.615
r103 25 37 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.445 $Y=2.375
+ $X2=1.28 $Y2=2.375
r104 24 26 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.93 $Y=2.375
+ $X2=2.095 $Y2=2.29
r105 24 25 31.6417 $w=1.68e-07 $l=4.85e-07 $layer=LI1_cond $X=1.93 $Y=2.375
+ $X2=1.445 $Y2=2.375
r106 19 46 25.1189 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=2.92 $Y=1.42
+ $X2=2.92 $Y2=1.642
r107 19 21 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=2.92 $Y=1.42 $X2=2.92
+ $Y2=1.02
r108 18 21 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=2.92 $Y=0.33
+ $X2=2.92 $Y2=1.02
r109 15 45 25.1189 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=2.905 $Y=1.865
+ $X2=2.905 $Y2=1.642
r110 15 17 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=2.905 $Y=1.865
+ $X2=2.905 $Y2=2.44
r111 12 44 25.1189 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=2.49 $Y=1.42
+ $X2=2.49 $Y2=1.642
r112 12 14 128.533 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=2.49 $Y=1.42 $X2=2.49
+ $Y2=1.02
r113 9 43 25.1189 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=2.285 $Y=1.865
+ $X2=2.285 $Y2=1.642
r114 9 11 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=2.285 $Y=1.865
+ $X2=2.285 $Y2=2.44
r115 8 38 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.69 $Y=0.255
+ $X2=1.525 $Y2=0.255
r116 7 18 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.845 $Y=0.255
+ $X2=2.92 $Y2=0.33
r117 7 8 592.245 $w=1.5e-07 $l=1.155e-06 $layer=POLY_cond $X=2.845 $Y=0.255
+ $X2=1.69 $Y2=0.255
r118 2 37 300 $w=1.7e-07 $l=5.65044e-07 $layer=licon1_PDIFF $count=2 $X=1.13
+ $Y=1.96 $X2=1.28 $Y2=2.455
r119 1 35 182 $w=1.7e-07 $l=5.80582e-07 $layer=licon1_NDIFF $count=1 $X=1
+ $Y=0.37 $X2=1.21 $Y2=0.855
.ends

.subckt PM_SKY130_FD_SC_HS__AND4BB_4%A_27_74# 1 2 10 12 13 15 19 21 22 24 26 28
+ 31 33 35 37 38 39 42 44 46 47 49 50 55 59
c135 44 0 2.63371e-20 $X=1.785 $Y=1.11
c136 26 0 3.95433e-21 $X=3.37 $Y=1.565
c137 12 0 1.75904e-19 $X=3.375 $Y=1.775
c138 10 0 2.67594e-19 $X=3.35 $Y=1.02
r139 57 59 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=1.785 $Y=0.84
+ $X2=1.945 $Y2=0.84
r140 54 55 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=1.59 $Y=1.195
+ $X2=1.785 $Y2=1.195
r141 50 61 17.2143 $w=2.52e-07 $l=9e-08 $layer=POLY_cond $X=3.44 $Y=0.42
+ $X2=3.35 $Y2=0.42
r142 49 50 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.44
+ $Y=0.42 $X2=3.44 $Y2=0.42
r143 47 49 49.2407 $w=3.28e-07 $l=1.41e-06 $layer=LI1_cond $X=2.03 $Y=0.42
+ $X2=3.44 $Y2=0.42
r144 46 59 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.945 $Y=0.755
+ $X2=1.945 $Y2=0.84
r145 45 47 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.945 $Y=0.585
+ $X2=2.03 $Y2=0.42
r146 45 46 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=1.945 $Y=0.585
+ $X2=1.945 $Y2=0.755
r147 44 55 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.785 $Y=1.11
+ $X2=1.785 $Y2=1.195
r148 43 57 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.785 $Y=0.925
+ $X2=1.785 $Y2=0.84
r149 43 44 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=1.785 $Y=0.925
+ $X2=1.785 $Y2=1.11
r150 41 54 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.59 $Y=1.28
+ $X2=1.59 $Y2=1.195
r151 41 42 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.59 $Y=1.28
+ $X2=1.59 $Y2=1.95
r152 40 53 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.445 $Y=2.035
+ $X2=0.28 $Y2=2.035
r153 39 42 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.505 $Y=2.035
+ $X2=1.59 $Y2=1.95
r154 39 40 69.1551 $w=1.68e-07 $l=1.06e-06 $layer=LI1_cond $X=1.505 $Y=2.035
+ $X2=0.445 $Y2=2.035
r155 37 54 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=1.505 $Y=1.195
+ $X2=1.59 $Y2=1.195
r156 37 38 74.3743 $w=1.68e-07 $l=1.14e-06 $layer=LI1_cond $X=1.505 $Y=1.195
+ $X2=0.365 $Y2=1.195
r157 33 53 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.28 $Y=2.12 $X2=0.28
+ $Y2=2.035
r158 33 35 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=0.28 $Y=2.12
+ $X2=0.28 $Y2=2.815
r159 29 38 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.24 $Y=1.11
+ $X2=0.365 $Y2=1.195
r160 29 31 27.4281 $w=2.48e-07 $l=5.95e-07 $layer=LI1_cond $X=0.24 $Y=1.11
+ $X2=0.24 $Y2=0.515
r161 27 28 60.4563 $w=1.8e-07 $l=1.5e-07 $layer=POLY_cond $X=3.825 $Y=1.415
+ $X2=3.825 $Y2=1.565
r162 25 26 60.4563 $w=1.8e-07 $l=1.5e-07 $layer=POLY_cond $X=3.37 $Y=1.415
+ $X2=3.37 $Y2=1.565
r163 22 24 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=3.855 $Y=1.865
+ $X2=3.855 $Y2=2.44
r164 21 22 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=3.855 $Y=1.775
+ $X2=3.855 $Y2=1.865
r165 21 28 81.629 $w=1.8e-07 $l=2.1e-07 $layer=POLY_cond $X=3.855 $Y=1.775
+ $X2=3.855 $Y2=1.565
r166 19 27 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=3.78 $Y=1.02
+ $X2=3.78 $Y2=1.415
r167 16 50 65.0317 $w=2.52e-07 $l=4.14367e-07 $layer=POLY_cond $X=3.78 $Y=0.585
+ $X2=3.44 $Y2=0.42
r168 16 19 223.053 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.78 $Y=0.585
+ $X2=3.78 $Y2=1.02
r169 13 15 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=3.375 $Y=1.865
+ $X2=3.375 $Y2=2.44
r170 12 13 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=3.375 $Y=1.775
+ $X2=3.375 $Y2=1.865
r171 12 26 81.629 $w=1.8e-07 $l=2.1e-07 $layer=POLY_cond $X=3.375 $Y=1.775
+ $X2=3.375 $Y2=1.565
r172 10 25 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=3.35 $Y=1.02
+ $X2=3.35 $Y2=1.415
r173 7 61 14.904 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.35 $Y=0.585
+ $X2=3.35 $Y2=0.42
r174 7 10 223.053 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.35 $Y=0.585
+ $X2=3.35 $Y2=1.02
r175 2 53 400 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.96 $X2=0.28 $Y2=2.115
r176 2 35 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.96 $X2=0.28 $Y2=2.815
r177 1 31 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__AND4BB_4%C 1 3 4 6 7 9 10 12 13 14 20
r54 20 22 27.3088 $w=3.53e-07 $l=2e-07 $layer=POLY_cond $X=5.27 $Y=1.657
+ $X2=5.47 $Y2=1.657
r55 19 20 56.6657 $w=3.53e-07 $l=4.15e-07 $layer=POLY_cond $X=4.855 $Y=1.657
+ $X2=5.27 $Y2=1.657
r56 18 19 2.04816 $w=3.53e-07 $l=1.5e-08 $layer=POLY_cond $X=4.84 $Y=1.657
+ $X2=4.855 $Y2=1.657
r57 17 18 59.3966 $w=3.53e-07 $l=4.35e-07 $layer=POLY_cond $X=4.405 $Y=1.657
+ $X2=4.84 $Y2=1.657
r58 13 14 18.5089 $w=3.28e-07 $l=5.3e-07 $layer=LI1_cond $X=5.47 $Y=1.615 $X2=6
+ $Y2=1.615
r59 13 22 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.47
+ $Y=1.615 $X2=5.47 $Y2=1.615
r60 10 20 22.8335 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=5.27 $Y=1.45
+ $X2=5.27 $Y2=1.657
r61 10 12 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=5.27 $Y=1.45
+ $X2=5.27 $Y2=1.005
r62 7 19 22.8335 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=4.855 $Y=1.865
+ $X2=4.855 $Y2=1.657
r63 7 9 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=4.855 $Y=1.865
+ $X2=4.855 $Y2=2.44
r64 4 18 22.8335 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.84 $Y=1.45
+ $X2=4.84 $Y2=1.657
r65 4 6 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=4.84 $Y=1.45 $X2=4.84
+ $Y2=1.005
r66 1 17 22.8335 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=4.405 $Y=1.865
+ $X2=4.405 $Y2=1.657
r67 1 3 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=4.405 $Y=1.865
+ $X2=4.405 $Y2=2.44
.ends

.subckt PM_SKY130_FD_SC_HS__AND4BB_4%D 1 3 6 10 12 14 15 21 22
c53 22 0 4.3247e-20 $X=6.71 $Y=1.515
c54 10 0 2.51603e-19 $X=6.69 $Y=0.79
r55 21 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.71
+ $Y=1.515 $X2=6.71 $Y2=1.515
r56 19 21 2.44051 $w=3.95e-07 $l=2e-08 $layer=POLY_cond $X=6.69 $Y=1.607
+ $X2=6.71 $Y2=1.607
r57 18 19 52.4709 $w=3.95e-07 $l=4.3e-07 $layer=POLY_cond $X=6.26 $Y=1.607
+ $X2=6.69 $Y2=1.607
r58 17 18 4.27089 $w=3.95e-07 $l=3.5e-08 $layer=POLY_cond $X=6.225 $Y=1.607
+ $X2=6.26 $Y2=1.607
r59 15 22 6.16423 $w=4.28e-07 $l=2.3e-07 $layer=LI1_cond $X=6.48 $Y=1.565
+ $X2=6.71 $Y2=1.565
r60 12 21 2.44051 $w=3.95e-07 $l=2e-08 $layer=POLY_cond $X=6.73 $Y=1.607
+ $X2=6.71 $Y2=1.607
r61 12 14 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=6.73 $Y=1.765
+ $X2=6.73 $Y2=2.34
r62 8 19 25.5547 $w=1.5e-07 $l=2.57e-07 $layer=POLY_cond $X=6.69 $Y=1.35
+ $X2=6.69 $Y2=1.607
r63 8 10 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=6.69 $Y=1.35 $X2=6.69
+ $Y2=0.79
r64 4 18 25.5547 $w=1.5e-07 $l=2.57e-07 $layer=POLY_cond $X=6.26 $Y=1.35
+ $X2=6.26 $Y2=1.607
r65 4 6 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=6.26 $Y=1.35 $X2=6.26
+ $Y2=0.79
r66 1 17 25.5547 $w=1.5e-07 $l=2.58e-07 $layer=POLY_cond $X=6.225 $Y=1.865
+ $X2=6.225 $Y2=1.607
r67 1 3 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=6.225 $Y=1.865
+ $X2=6.225 $Y2=2.44
.ends

.subckt PM_SKY130_FD_SC_HS__AND4BB_4%A_472_388# 1 2 3 4 5 18 20 22 25 27 29 32
+ 34 36 37 39 42 46 51 52 56 60 63 66 68 72 75 76 81 84 86 89 91 93 102
c176 86 0 1.54641e-19 $X=2.705 $Y=1.185
c177 75 0 5.63592e-20 $X=7.15 $Y=1.95
c178 51 0 2.58135e-19 $X=2.65 $Y=1.595
c179 46 0 5.70593e-20 $X=2.595 $Y=2.085
c180 20 0 4.3247e-20 $X=7.265 $Y=1.765
r181 102 103 0.644385 $w=3.74e-07 $l=5e-09 $layer=POLY_cond $X=8.615 $Y=1.542
+ $X2=8.62 $Y2=1.542
r182 99 100 1.93316 $w=3.74e-07 $l=1.5e-08 $layer=POLY_cond $X=8.15 $Y=1.542
+ $X2=8.165 $Y2=1.542
r183 98 99 56.0615 $w=3.74e-07 $l=4.35e-07 $layer=POLY_cond $X=7.715 $Y=1.542
+ $X2=8.15 $Y2=1.542
r184 97 98 12.2433 $w=3.74e-07 $l=9.5e-08 $layer=POLY_cond $X=7.62 $Y=1.542
+ $X2=7.715 $Y2=1.542
r185 94 95 9.66578 $w=3.74e-07 $l=7.5e-08 $layer=POLY_cond $X=7.19 $Y=1.542
+ $X2=7.265 $Y2=1.542
r186 86 88 7.39493 $w=3.28e-07 $l=1.75e-07 $layer=LI1_cond $X=2.705 $Y=1.185
+ $X2=2.705 $Y2=1.36
r187 82 102 27.7086 $w=3.74e-07 $l=2.15e-07 $layer=POLY_cond $X=8.4 $Y=1.542
+ $X2=8.615 $Y2=1.542
r188 82 100 30.2861 $w=3.74e-07 $l=2.35e-07 $layer=POLY_cond $X=8.4 $Y=1.542
+ $X2=8.165 $Y2=1.542
r189 81 82 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=8.4
+ $Y=1.485 $X2=8.4 $Y2=1.485
r190 79 97 30.9305 $w=3.74e-07 $l=2.4e-07 $layer=POLY_cond $X=7.38 $Y=1.542
+ $X2=7.62 $Y2=1.542
r191 79 95 14.8209 $w=3.74e-07 $l=1.15e-07 $layer=POLY_cond $X=7.38 $Y=1.542
+ $X2=7.265 $Y2=1.542
r192 78 81 35.621 $w=3.28e-07 $l=1.02e-06 $layer=LI1_cond $X=7.38 $Y=1.485
+ $X2=8.4 $Y2=1.485
r193 78 79 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=7.38
+ $Y=1.485 $X2=7.38 $Y2=1.485
r194 76 78 5.06376 $w=3.28e-07 $l=1.45e-07 $layer=LI1_cond $X=7.235 $Y=1.485
+ $X2=7.38 $Y2=1.485
r195 74 76 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=7.15 $Y=1.65
+ $X2=7.235 $Y2=1.485
r196 74 75 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=7.15 $Y=1.65 $X2=7.15
+ $Y2=1.95
r197 73 93 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.665 $Y=2.035
+ $X2=6.5 $Y2=2.035
r198 72 75 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.065 $Y=2.035
+ $X2=7.15 $Y2=1.95
r199 72 73 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=7.065 $Y=2.035
+ $X2=6.665 $Y2=2.035
r200 69 91 3.80956 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.795 $Y=2.035
+ $X2=4.63 $Y2=2.035
r201 68 93 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.335 $Y=2.035
+ $X2=6.5 $Y2=2.035
r202 68 69 100.471 $w=1.68e-07 $l=1.54e-06 $layer=LI1_cond $X=6.335 $Y=2.035
+ $X2=4.795 $Y2=2.035
r203 64 91 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.63 $Y=2.12
+ $X2=4.63 $Y2=2.035
r204 64 66 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=4.63 $Y=2.12
+ $X2=4.63 $Y2=2.795
r205 63 91 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.63 $Y=1.95
+ $X2=4.63 $Y2=2.035
r206 62 63 6.46067 $w=3.28e-07 $l=1.85e-07 $layer=LI1_cond $X=4.63 $Y=1.765
+ $X2=4.63 $Y2=1.95
r207 61 89 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.795 $Y=1.68
+ $X2=3.63 $Y2=1.68
r208 60 62 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.465 $Y=1.68
+ $X2=4.63 $Y2=1.765
r209 60 61 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.465 $Y=1.68
+ $X2=3.795 $Y2=1.68
r210 56 58 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=3.63 $Y=2.085
+ $X2=3.63 $Y2=2.795
r211 54 89 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.63 $Y=1.765
+ $X2=3.63 $Y2=1.68
r212 54 56 11.1752 $w=3.28e-07 $l=3.2e-07 $layer=LI1_cond $X=3.63 $Y=1.765
+ $X2=3.63 $Y2=2.085
r213 53 84 3.11956 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.76 $Y=1.68
+ $X2=2.595 $Y2=1.68
r214 52 89 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.465 $Y=1.68
+ $X2=3.63 $Y2=1.68
r215 52 53 45.9947 $w=1.68e-07 $l=7.05e-07 $layer=LI1_cond $X=3.465 $Y=1.68
+ $X2=2.76 $Y2=1.68
r216 51 84 3.40559 $w=2.75e-07 $l=1.09087e-07 $layer=LI1_cond $X=2.65 $Y=1.595
+ $X2=2.595 $Y2=1.68
r217 51 88 12.3102 $w=2.18e-07 $l=2.35e-07 $layer=LI1_cond $X=2.65 $Y=1.595
+ $X2=2.65 $Y2=1.36
r218 46 48 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=2.595 $Y=2.085
+ $X2=2.595 $Y2=2.795
r219 44 84 3.40559 $w=2.75e-07 $l=8.5e-08 $layer=LI1_cond $X=2.595 $Y=1.765
+ $X2=2.595 $Y2=1.68
r220 44 46 11.1752 $w=3.28e-07 $l=3.2e-07 $layer=LI1_cond $X=2.595 $Y=1.765
+ $X2=2.595 $Y2=2.085
r221 40 103 24.2268 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=8.62 $Y=1.32
+ $X2=8.62 $Y2=1.542
r222 40 42 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=8.62 $Y=1.32
+ $X2=8.62 $Y2=0.74
r223 37 102 24.2268 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=8.615 $Y=1.765
+ $X2=8.615 $Y2=1.542
r224 37 39 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=8.615 $Y=1.765
+ $X2=8.615 $Y2=2.4
r225 34 100 24.2268 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=8.165 $Y=1.765
+ $X2=8.165 $Y2=1.542
r226 34 36 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=8.165 $Y=1.765
+ $X2=8.165 $Y2=2.4
r227 30 99 24.2268 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=8.15 $Y=1.32
+ $X2=8.15 $Y2=1.542
r228 30 32 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=8.15 $Y=1.32
+ $X2=8.15 $Y2=0.74
r229 27 98 24.2268 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=7.715 $Y=1.765
+ $X2=7.715 $Y2=1.542
r230 27 29 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=7.715 $Y=1.765
+ $X2=7.715 $Y2=2.4
r231 23 97 24.2268 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=7.62 $Y=1.32
+ $X2=7.62 $Y2=1.542
r232 23 25 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=7.62 $Y=1.32
+ $X2=7.62 $Y2=0.74
r233 20 95 24.2268 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=7.265 $Y=1.765
+ $X2=7.265 $Y2=1.542
r234 20 22 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=7.265 $Y=1.765
+ $X2=7.265 $Y2=2.4
r235 16 94 24.2268 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=7.19 $Y=1.32
+ $X2=7.19 $Y2=1.542
r236 16 18 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=7.19 $Y=1.32
+ $X2=7.19 $Y2=0.74
r237 5 93 300 $w=1.7e-07 $l=2.54951e-07 $layer=licon1_PDIFF $count=2 $X=6.3
+ $Y=1.94 $X2=6.5 $Y2=2.065
r238 4 91 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=4.48
+ $Y=1.94 $X2=4.63 $Y2=2.085
r239 4 66 400 $w=1.7e-07 $l=9.26971e-07 $layer=licon1_PDIFF $count=1 $X=4.48
+ $Y=1.94 $X2=4.63 $Y2=2.795
r240 3 58 400 $w=1.7e-07 $l=9.40705e-07 $layer=licon1_PDIFF $count=1 $X=3.45
+ $Y=1.94 $X2=3.63 $Y2=2.795
r241 3 56 400 $w=1.7e-07 $l=2.41868e-07 $layer=licon1_PDIFF $count=1 $X=3.45
+ $Y=1.94 $X2=3.63 $Y2=2.085
r242 2 48 400 $w=1.7e-07 $l=9.65376e-07 $layer=licon1_PDIFF $count=1 $X=2.36
+ $Y=1.94 $X2=2.595 $Y2=2.795
r243 2 46 400 $w=1.7e-07 $l=2.98831e-07 $layer=licon1_PDIFF $count=1 $X=2.36
+ $Y=1.94 $X2=2.595 $Y2=2.085
r244 1 86 182 $w=1.7e-07 $l=5.50568e-07 $layer=licon1_NDIFF $count=1 $X=2.565
+ $Y=0.7 $X2=2.705 $Y2=1.185
.ends

.subckt PM_SKY130_FD_SC_HS__AND4BB_4%VPWR 1 2 3 4 5 6 7 8 27 31 35 41 49 55 57
+ 59 62 63 64 66 75 79 84 89 94 100 103 106 111 118 120 123 127
c120 8 0 1.8444e-19 $X=8.69 $Y=1.84
r121 126 127 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r122 123 124 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r123 120 121 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r124 115 118 13.5255 $w=1.123e-06 $l=1.65e-07 $layer=LI1_cond $X=6 $Y=2.852
+ $X2=6.165 $Y2=2.852
r125 115 117 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r126 113 115 9.43467 $w=1.123e-06 $l=8.7e-07 $layer=LI1_cond $X=5.13 $Y=2.852
+ $X2=6 $Y2=2.852
r127 110 117 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=6 $Y2=3.33
r128 109 113 0.976 $w=1.123e-06 $l=9e-08 $layer=LI1_cond $X=5.04 $Y=2.852
+ $X2=5.13 $Y2=2.852
r129 109 111 12.5495 $w=1.123e-06 $l=7.5e-08 $layer=LI1_cond $X=5.04 $Y=2.852
+ $X2=4.965 $Y2=2.852
r130 109 110 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r131 106 107 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r132 103 104 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r133 100 101 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r134 98 127 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=3.33
+ $X2=8.88 $Y2=3.33
r135 98 124 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=3.33
+ $X2=7.92 $Y2=3.33
r136 97 98 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=3.33 $X2=8.4
+ $Y2=3.33
r137 95 123 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.105 $Y=3.33
+ $X2=7.94 $Y2=3.33
r138 95 97 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=8.105 $Y=3.33
+ $X2=8.4 $Y2=3.33
r139 94 126 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=8.675 $Y=3.33
+ $X2=8.897 $Y2=3.33
r140 94 97 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=8.675 $Y=3.33
+ $X2=8.4 $Y2=3.33
r141 93 124 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=7.92 $Y2=3.33
r142 93 121 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=6.96 $Y2=3.33
r143 92 93 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r144 90 120 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.205 $Y=3.33
+ $X2=7.04 $Y2=3.33
r145 90 92 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=7.205 $Y=3.33
+ $X2=7.44 $Y2=3.33
r146 89 123 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.775 $Y=3.33
+ $X2=7.94 $Y2=3.33
r147 89 92 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=7.775 $Y=3.33
+ $X2=7.44 $Y2=3.33
r148 88 121 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=6.96 $Y2=3.33
r149 88 117 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=6 $Y2=3.33
r150 87 118 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=6.48 $Y=3.33
+ $X2=6.165 $Y2=3.33
r151 87 88 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r152 84 120 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.875 $Y=3.33
+ $X2=7.04 $Y2=3.33
r153 84 87 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=6.875 $Y=3.33
+ $X2=6.48 $Y2=3.33
r154 83 107 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.08 $Y2=3.33
r155 83 104 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=3.12 $Y2=3.33
r156 82 83 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r157 80 103 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.295 $Y=3.33
+ $X2=3.13 $Y2=3.33
r158 80 82 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=3.295 $Y=3.33
+ $X2=3.6 $Y2=3.33
r159 79 106 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.965 $Y=3.33
+ $X2=4.13 $Y2=3.33
r160 79 82 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=3.965 $Y=3.33
+ $X2=3.6 $Y2=3.33
r161 78 104 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r162 77 78 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r163 75 103 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.965 $Y=3.33
+ $X2=3.13 $Y2=3.33
r164 75 77 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=2.965 $Y=3.33
+ $X2=2.64 $Y2=3.33
r165 74 78 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.64 $Y2=3.33
r166 74 101 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=0.72 $Y2=3.33
r167 73 74 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r168 71 100 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.945 $Y=3.33
+ $X2=0.78 $Y2=3.33
r169 71 73 47.9519 $w=1.68e-07 $l=7.35e-07 $layer=LI1_cond $X=0.945 $Y=3.33
+ $X2=1.68 $Y2=3.33
r170 69 101 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r171 68 69 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r172 66 100 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.615 $Y=3.33
+ $X2=0.78 $Y2=3.33
r173 66 68 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=0.615 $Y=3.33
+ $X2=0.24 $Y2=3.33
r174 64 110 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=5.04 $Y2=3.33
r175 64 107 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=4.08 $Y2=3.33
r176 62 73 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=1.89 $Y=3.33
+ $X2=1.68 $Y2=3.33
r177 62 63 8.70163 $w=1.7e-07 $l=1.67e-07 $layer=LI1_cond $X=1.89 $Y=3.33
+ $X2=2.057 $Y2=3.33
r178 61 77 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=2.225 $Y=3.33
+ $X2=2.64 $Y2=3.33
r179 61 63 8.70163 $w=1.7e-07 $l=1.68e-07 $layer=LI1_cond $X=2.225 $Y=3.33
+ $X2=2.057 $Y2=3.33
r180 57 126 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=8.84 $Y=3.245
+ $X2=8.897 $Y2=3.33
r181 57 59 29.3349 $w=3.28e-07 $l=8.4e-07 $layer=LI1_cond $X=8.84 $Y=3.245
+ $X2=8.84 $Y2=2.405
r182 53 123 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.94 $Y=3.245
+ $X2=7.94 $Y2=3.33
r183 53 55 29.3349 $w=3.28e-07 $l=8.4e-07 $layer=LI1_cond $X=7.94 $Y=3.245
+ $X2=7.94 $Y2=2.405
r184 49 52 12.5721 $w=3.28e-07 $l=3.6e-07 $layer=LI1_cond $X=7.04 $Y=2.455
+ $X2=7.04 $Y2=2.815
r185 47 120 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.04 $Y=3.245
+ $X2=7.04 $Y2=3.33
r186 47 52 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=7.04 $Y=3.245
+ $X2=7.04 $Y2=2.815
r187 46 106 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.295 $Y=3.33
+ $X2=4.13 $Y2=3.33
r188 46 111 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.295 $Y=3.33
+ $X2=4.965 $Y2=3.33
r189 41 44 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=4.13 $Y=2.1
+ $X2=4.13 $Y2=2.795
r190 39 106 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.13 $Y=3.245
+ $X2=4.13 $Y2=3.33
r191 39 44 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=4.13 $Y=3.245
+ $X2=4.13 $Y2=2.795
r192 35 38 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=3.13 $Y=2.1
+ $X2=3.13 $Y2=2.795
r193 33 103 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.13 $Y=3.245
+ $X2=3.13 $Y2=3.33
r194 33 38 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=3.13 $Y=3.245
+ $X2=3.13 $Y2=2.795
r195 29 63 0.942324 $w=3.35e-07 $l=8.5e-08 $layer=LI1_cond $X=2.057 $Y=3.245
+ $X2=2.057 $Y2=3.33
r196 29 31 17.0286 $w=3.33e-07 $l=4.95e-07 $layer=LI1_cond $X=2.057 $Y=3.245
+ $X2=2.057 $Y2=2.75
r197 25 100 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.78 $Y=3.245
+ $X2=0.78 $Y2=3.33
r198 25 27 27.5888 $w=3.28e-07 $l=7.9e-07 $layer=LI1_cond $X=0.78 $Y=3.245
+ $X2=0.78 $Y2=2.455
r199 8 59 300 $w=1.7e-07 $l=6.3559e-07 $layer=licon1_PDIFF $count=2 $X=8.69
+ $Y=1.84 $X2=8.84 $Y2=2.405
r200 7 55 300 $w=1.7e-07 $l=6.3559e-07 $layer=licon1_PDIFF $count=2 $X=7.79
+ $Y=1.84 $X2=7.94 $Y2=2.405
r201 6 52 600 $w=1.7e-07 $l=1.08616e-06 $layer=licon1_PDIFF $count=1 $X=6.805
+ $Y=1.84 $X2=7.04 $Y2=2.815
r202 6 49 600 $w=1.7e-07 $l=7.23015e-07 $layer=licon1_PDIFF $count=1 $X=6.805
+ $Y=1.84 $X2=7.04 $Y2=2.455
r203 5 115 200 $w=1.7e-07 $l=1.269e-06 $layer=licon1_PDIFF $count=3 $X=4.93
+ $Y=1.94 $X2=6 $Y2=2.375
r204 5 113 200 $w=1.7e-07 $l=5.25571e-07 $layer=licon1_PDIFF $count=3 $X=4.93
+ $Y=1.94 $X2=5.13 $Y2=2.375
r205 4 44 400 $w=1.7e-07 $l=9.4975e-07 $layer=licon1_PDIFF $count=1 $X=3.93
+ $Y=1.94 $X2=4.13 $Y2=2.795
r206 4 41 400 $w=1.7e-07 $l=2.68328e-07 $layer=licon1_PDIFF $count=1 $X=3.93
+ $Y=1.94 $X2=4.13 $Y2=2.1
r207 3 38 400 $w=1.7e-07 $l=9.26971e-07 $layer=licon1_PDIFF $count=1 $X=2.98
+ $Y=1.94 $X2=3.13 $Y2=2.795
r208 3 35 400 $w=1.7e-07 $l=2.22711e-07 $layer=licon1_PDIFF $count=1 $X=2.98
+ $Y=1.94 $X2=3.13 $Y2=2.1
r209 2 31 600 $w=1.7e-07 $l=8.88679e-07 $layer=licon1_PDIFF $count=1 $X=1.89
+ $Y=1.94 $X2=2.055 $Y2=2.75
r210 1 27 300 $w=1.7e-07 $l=5.86536e-07 $layer=licon1_PDIFF $count=2 $X=0.58
+ $Y=1.96 $X2=0.78 $Y2=2.455
.ends

.subckt PM_SKY130_FD_SC_HS__AND4BB_4%X 1 2 3 4 15 17 19 22 23 27 28 33 34 35 36
+ 37 42 43
c64 27 0 1.28179e-19 $X=8.765 $Y=0.96
c65 23 0 1.8444e-19 $X=8.765 $Y=1.985
c66 22 0 1.0664e-19 $X=7.57 $Y=1.065
r67 37 43 4.18573 $w=2.3e-07 $l=1.65e-07 $layer=LI1_cond $X=8.88 $Y=1.985
+ $X2=8.88 $Y2=1.82
r68 36 43 7.76646 $w=2.28e-07 $l=1.55e-07 $layer=LI1_cond $X=8.88 $Y=1.665
+ $X2=8.88 $Y2=1.82
r69 35 36 18.5393 $w=2.28e-07 $l=3.7e-07 $layer=LI1_cond $X=8.88 $Y=1.295
+ $X2=8.88 $Y2=1.665
r70 35 42 7.2654 $w=2.28e-07 $l=1.45e-07 $layer=LI1_cond $X=8.88 $Y=1.295
+ $X2=8.88 $Y2=1.15
r71 34 42 4.58911 $w=2.3e-07 $l=1.9e-07 $layer=LI1_cond $X=8.88 $Y=0.96 $X2=8.88
+ $Y2=1.15
r72 32 33 8.5712 $w=3.78e-07 $l=1.65e-07 $layer=LI1_cond $X=8.405 $Y=0.96
+ $X2=8.24 $Y2=0.96
r73 28 32 0.758186 $w=3.78e-07 $l=2.5e-08 $layer=LI1_cond $X=8.43 $Y=0.96
+ $X2=8.405 $Y2=0.96
r74 27 34 2.77762 $w=3.8e-07 $l=1.15e-07 $layer=LI1_cond $X=8.765 $Y=0.96
+ $X2=8.88 $Y2=0.96
r75 27 28 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=8.765 $Y=0.96
+ $X2=8.43 $Y2=0.96
r76 24 30 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.575 $Y=1.985
+ $X2=7.49 $Y2=1.985
r77 24 26 28.4618 $w=3.28e-07 $l=8.15e-07 $layer=LI1_cond $X=7.575 $Y=1.985
+ $X2=8.39 $Y2=1.985
r78 23 37 2.91733 $w=3.3e-07 $l=1.15e-07 $layer=LI1_cond $X=8.765 $Y=1.985
+ $X2=8.88 $Y2=1.985
r79 23 26 13.0959 $w=3.28e-07 $l=3.75e-07 $layer=LI1_cond $X=8.765 $Y=1.985
+ $X2=8.39 $Y2=1.985
r80 22 33 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=7.57 $Y=1.065
+ $X2=8.24 $Y2=1.065
r81 17 30 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.49 $Y=2.15
+ $X2=7.49 $Y2=1.985
r82 17 19 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=7.49 $Y=2.15
+ $X2=7.49 $Y2=2.4
r83 13 22 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=7.405 $Y=0.98
+ $X2=7.57 $Y2=1.065
r84 13 15 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=7.405 $Y=0.98
+ $X2=7.405 $Y2=0.515
r85 4 26 600 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=8.24
+ $Y=1.84 $X2=8.39 $Y2=1.985
r86 3 30 600 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=7.34
+ $Y=1.84 $X2=7.49 $Y2=1.985
r87 3 19 300 $w=1.7e-07 $l=6.30555e-07 $layer=licon1_PDIFF $count=2 $X=7.34
+ $Y=1.84 $X2=7.49 $Y2=2.4
r88 2 32 182 $w=1.7e-07 $l=6.63928e-07 $layer=licon1_NDIFF $count=1 $X=8.225
+ $Y=0.37 $X2=8.405 $Y2=0.95
r89 1 15 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=7.265
+ $Y=0.37 $X2=7.405 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__AND4BB_4%VGND 1 2 3 4 5 18 22 26 30 32 34 36 38 43
+ 51 56 61 67 70 73 76 80
c97 5 0 1.28179e-19 $X=8.695 $Y=0.37
r98 79 80 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=0 $X2=8.88
+ $Y2=0
r99 76 77 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=0 $X2=7.92
+ $Y2=0
r100 73 74 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=0 $X2=6.96
+ $Y2=0
r101 70 71 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=0 $X2=6 $Y2=0
r102 67 68 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r103 65 80 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=0 $X2=8.88
+ $Y2=0
r104 65 77 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=0 $X2=7.92
+ $Y2=0
r105 64 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r106 62 76 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.07 $Y=0 $X2=7.905
+ $Y2=0
r107 62 64 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=8.07 $Y=0 $X2=8.4
+ $Y2=0
r108 61 79 4.77426 $w=1.7e-07 $l=2.25e-07 $layer=LI1_cond $X=8.67 $Y=0 $X2=8.895
+ $Y2=0
r109 61 64 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=8.67 $Y=0 $X2=8.4
+ $Y2=0
r110 60 77 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=0 $X2=7.92
+ $Y2=0
r111 60 74 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=0 $X2=6.96
+ $Y2=0
r112 59 60 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=0 $X2=7.44
+ $Y2=0
r113 57 73 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.07 $Y=0 $X2=6.905
+ $Y2=0
r114 57 59 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=7.07 $Y=0 $X2=7.44
+ $Y2=0
r115 56 76 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.74 $Y=0 $X2=7.905
+ $Y2=0
r116 56 59 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=7.74 $Y=0 $X2=7.44
+ $Y2=0
r117 55 74 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=0 $X2=6.96
+ $Y2=0
r118 55 71 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=0 $X2=6
+ $Y2=0
r119 54 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=0 $X2=6.48
+ $Y2=0
r120 52 70 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.13 $Y=0 $X2=6.005
+ $Y2=0
r121 52 54 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=6.13 $Y=0 $X2=6.48
+ $Y2=0
r122 51 73 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.74 $Y=0 $X2=6.905
+ $Y2=0
r123 51 54 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=6.74 $Y=0 $X2=6.48
+ $Y2=0
r124 50 71 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=6
+ $Y2=0
r125 49 50 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r126 47 68 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r127 46 49 281.84 $w=1.68e-07 $l=4.32e-06 $layer=LI1_cond $X=1.2 $Y=0 $X2=5.52
+ $Y2=0
r128 46 47 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r129 44 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.875 $Y=0 $X2=0.71
+ $Y2=0
r130 44 46 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.875 $Y=0 $X2=1.2
+ $Y2=0
r131 43 70 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.88 $Y=0 $X2=6.005
+ $Y2=0
r132 43 49 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=5.88 $Y=0 $X2=5.52
+ $Y2=0
r133 41 68 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r134 40 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r135 38 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.545 $Y=0 $X2=0.71
+ $Y2=0
r136 38 40 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.545 $Y=0
+ $X2=0.24 $Y2=0
r137 36 50 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=5.52
+ $Y2=0
r138 36 47 0.936549 $w=4.9e-07 $l=3.36e-06 $layer=MET1_cond $X=4.56 $Y=0 $X2=1.2
+ $Y2=0
r139 32 79 3.03431 $w=3.35e-07 $l=1.1025e-07 $layer=LI1_cond $X=8.837 $Y=0.085
+ $X2=8.895 $Y2=0
r140 32 34 14.7926 $w=3.33e-07 $l=4.3e-07 $layer=LI1_cond $X=8.837 $Y=0.085
+ $X2=8.837 $Y2=0.515
r141 28 76 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.905 $Y=0.085
+ $X2=7.905 $Y2=0
r142 28 30 19.5566 $w=3.28e-07 $l=5.6e-07 $layer=LI1_cond $X=7.905 $Y=0.085
+ $X2=7.905 $Y2=0.645
r143 24 73 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.905 $Y=0.085
+ $X2=6.905 $Y2=0
r144 24 26 18.5089 $w=3.28e-07 $l=5.3e-07 $layer=LI1_cond $X=6.905 $Y=0.085
+ $X2=6.905 $Y2=0.615
r145 20 70 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.005 $Y=0.085
+ $X2=6.005 $Y2=0
r146 20 22 25.8147 $w=2.48e-07 $l=5.6e-07 $layer=LI1_cond $X=6.005 $Y=0.085
+ $X2=6.005 $Y2=0.645
r147 16 67 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.71 $Y=0.085
+ $X2=0.71 $Y2=0
r148 16 18 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=0.71 $Y=0.085
+ $X2=0.71 $Y2=0.495
r149 5 34 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=8.695
+ $Y=0.37 $X2=8.835 $Y2=0.515
r150 4 30 182 $w=1.7e-07 $l=3.65205e-07 $layer=licon1_NDIFF $count=1 $X=7.695
+ $Y=0.37 $X2=7.905 $Y2=0.645
r151 3 26 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=6.765
+ $Y=0.47 $X2=6.905 $Y2=0.615
r152 2 22 182 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_NDIFF $count=1 $X=5.9
+ $Y=0.47 $X2=6.045 $Y2=0.645
r153 1 18 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=0.57
+ $Y=0.37 $X2=0.71 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_HS__AND4BB_4%A_412_140# 1 2 3 11 12 13 18 19 26
c44 26 0 3.95433e-21 $X=3.995 $Y=1.185
c45 13 0 6.58453e-20 $X=2.37 $Y=0.84
r46 26 28 5.41299 $w=3.28e-07 $l=1.55e-07 $layer=LI1_cond $X=3.995 $Y=1.185
+ $X2=3.995 $Y2=1.34
r47 18 28 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.83 $Y=1.34
+ $X2=3.995 $Y2=1.34
r48 18 19 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=3.83 $Y=1.34
+ $X2=3.22 $Y2=1.34
r49 15 19 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.135 $Y=1.255
+ $X2=3.22 $Y2=1.34
r50 15 17 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=3.135 $Y=1.255
+ $X2=3.135 $Y2=1.055
r51 14 17 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=3.135 $Y=0.925
+ $X2=3.135 $Y2=1.055
r52 12 14 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.05 $Y=0.84
+ $X2=3.135 $Y2=0.925
r53 12 13 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=3.05 $Y=0.84
+ $X2=2.37 $Y2=0.84
r54 11 21 4.79607 $w=1.83e-07 $l=8e-08 $layer=LI1_cond $X=2.285 $Y=1.187
+ $X2=2.205 $Y2=1.187
r55 10 13 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.285 $Y=0.925
+ $X2=2.37 $Y2=0.84
r56 10 11 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=2.285 $Y=0.925
+ $X2=2.285 $Y2=1.095
r57 3 26 182 $w=1.7e-07 $l=5.50568e-07 $layer=licon1_NDIFF $count=1 $X=3.855
+ $Y=0.7 $X2=3.995 $Y2=1.185
r58 2 17 182 $w=1.7e-07 $l=4.19196e-07 $layer=licon1_NDIFF $count=1 $X=2.995
+ $Y=0.7 $X2=3.135 $Y2=1.055
r59 1 21 182 $w=1.7e-07 $l=5.52766e-07 $layer=licon1_NDIFF $count=1 $X=2.06
+ $Y=0.7 $X2=2.205 $Y2=1.185
.ends

.subckt PM_SKY130_FD_SC_HS__AND4BB_4%A_685_140# 1 2 11 14 15
c29 11 0 9.745e-20 $X=3.565 $Y=0.92
r30 14 15 8.58424 $w=2.73e-07 $l=1.65e-07 $layer=LI1_cond $X=5.055 $Y=0.802
+ $X2=4.89 $Y2=0.802
r31 8 11 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.65 $Y=0.84
+ $X2=3.525 $Y2=0.84
r32 8 15 80.8984 $w=1.68e-07 $l=1.24e-06 $layer=LI1_cond $X=3.65 $Y=0.84
+ $X2=4.89 $Y2=0.84
r33 2 14 182 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_NDIFF $count=1 $X=4.915
+ $Y=0.685 $X2=5.055 $Y2=0.84
r34 1 11 182 $w=1.7e-07 $l=2.81425e-07 $layer=licon1_NDIFF $count=1 $X=3.425
+ $Y=0.7 $X2=3.565 $Y2=0.92
.ends

.subckt PM_SKY130_FD_SC_HS__AND4BB_4%A_882_137# 1 2 3 10 14 16 20 25 27
c44 20 0 1.44963e-19 $X=6.475 $Y=0.615
r45 23 25 8.79328 $w=2.48e-07 $l=1.65e-07 $layer=LI1_cond $X=4.555 $Y=1.22
+ $X2=4.72 $Y2=1.22
r46 18 20 18.2086 $w=2.48e-07 $l=3.95e-07 $layer=LI1_cond $X=6.435 $Y=1.01
+ $X2=6.435 $Y2=0.615
r47 17 27 7.02821 $w=1.7e-07 $l=1.47902e-07 $layer=LI1_cond $X=5.65 $Y=1.095
+ $X2=5.525 $Y2=1.145
r48 16 18 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=6.31 $Y=1.095
+ $X2=6.435 $Y2=1.01
r49 16 17 43.0588 $w=1.68e-07 $l=6.6e-07 $layer=LI1_cond $X=6.31 $Y=1.095
+ $X2=5.65 $Y2=1.095
r50 12 27 0.00168595 $w=2.5e-07 $l=1.35e-07 $layer=LI1_cond $X=5.525 $Y=1.01
+ $X2=5.525 $Y2=1.145
r51 12 14 8.29759 $w=2.48e-07 $l=1.8e-07 $layer=LI1_cond $X=5.525 $Y=1.01
+ $X2=5.525 $Y2=0.83
r52 10 27 7.02821 $w=1.7e-07 $l=1.47902e-07 $layer=LI1_cond $X=5.4 $Y=1.195
+ $X2=5.525 $Y2=1.145
r53 10 25 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=5.4 $Y=1.195
+ $X2=4.72 $Y2=1.195
r54 3 20 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=6.335
+ $Y=0.47 $X2=6.475 $Y2=0.615
r55 2 27 182 $w=1.7e-07 $l=5.7576e-07 $layer=licon1_NDIFF $count=1 $X=5.345
+ $Y=0.685 $X2=5.485 $Y2=1.195
r56 2 14 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=5.345
+ $Y=0.685 $X2=5.485 $Y2=0.83
r57 1 23 182 $w=1.7e-07 $l=5.6285e-07 $layer=licon1_NDIFF $count=1 $X=4.41
+ $Y=0.685 $X2=4.555 $Y2=1.18
.ends

