# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_hs__xnor2_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.360000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.501000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.515000 1.350000 1.845000 1.780000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.501000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.945000 1.435000 1.345000 1.780000 ;
        RECT 1.175000 1.780000 1.345000 1.950000 ;
        RECT 1.175000 1.950000 2.185000 2.120000 ;
        RECT 2.015000 1.350000 2.465000 1.680000 ;
        RECT 2.015000 1.680000 2.185000 1.950000 ;
    END
  END B
  PIN Y
    ANTENNADIFFAREA  0.699800 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.045000 2.290000 2.685000 2.980000 ;
        RECT 2.355000 1.850000 3.275000 2.020000 ;
        RECT 2.355000 2.020000 2.685000 2.290000 ;
        RECT 2.975000 0.350000 3.275000 1.130000 ;
        RECT 3.105000 1.130000 3.275000 1.850000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 3.360000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 3.360000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.360000 0.085000 ;
      RECT 0.000000  3.245000 3.360000 3.415000 ;
      RECT 0.105000  0.085000 0.435000 1.255000 ;
      RECT 0.175000  1.905000 0.425000 2.290000 ;
      RECT 0.175000  2.290000 0.505000 3.245000 ;
      RECT 0.605000  1.085000 2.805000 1.180000 ;
      RECT 0.605000  1.180000 1.225000 1.255000 ;
      RECT 0.605000  1.255000 0.775000 1.950000 ;
      RECT 0.605000  1.950000 1.005000 2.120000 ;
      RECT 0.675000  2.120000 1.005000 2.785000 ;
      RECT 0.895000  0.575000 1.225000 1.010000 ;
      RECT 0.895000  1.010000 2.805000 1.085000 ;
      RECT 1.415000  2.290000 1.745000 3.245000 ;
      RECT 1.435000  0.510000 1.765000 0.670000 ;
      RECT 1.435000  0.670000 2.770000 0.840000 ;
      RECT 1.935000  0.085000 2.265000 0.500000 ;
      RECT 2.440000  0.510000 2.770000 0.670000 ;
      RECT 2.635000  1.180000 2.805000 1.300000 ;
      RECT 2.635000  1.300000 2.935000 1.630000 ;
      RECT 2.855000  2.190000 3.185000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
  END
END sky130_fd_sc_hs__xnor2_1
