* File: sky130_fd_sc_hs__o211a_4.spice
* Created: Tue Sep  1 20:13:47 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hs__o211a_4.pex.spice"
.subckt sky130_fd_sc_hs__o211a_4  VNB VPB C1 B1 A2 A1 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A1	A1
* A2	A2
* B1	B1
* C1	C1
* VPB	VPB
* VNB	VNB
MM1000 N_VGND_M1000_d N_A_91_48#_M1000_g N_X_M1000_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.1036 PD=2.05 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75001.6 A=0.111 P=1.78 MULT=1
MM1013 N_VGND_M1013_d N_A_91_48#_M1013_g N_X_M1000_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1295 AS=0.1036 PD=1.09 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.6
+ SB=75001.1 A=0.111 P=1.78 MULT=1
MM1016 N_VGND_M1013_d N_A_91_48#_M1016_g N_X_M1016_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1295 AS=0.1036 PD=1.09 PS=1.02 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75001.1
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1017 N_VGND_M1017_d N_A_91_48#_M1017_g N_X_M1016_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.1036 PD=2.05 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.6
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1014 N_A_510_125#_M1014_d N_B1_M1014_g N_A_597_125#_M1014_s VNB NLOWVT L=0.15
+ W=0.64 AD=0.1817 AS=0.0896 PD=1.85 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75003.5 A=0.096 P=1.58 MULT=1
MM1015 N_A_597_125#_M1014_s N_C1_M1015_g N_A_91_48#_M1015_s VNB NLOWVT L=0.15
+ W=0.64 AD=0.0896 AS=0.0896 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.6 SB=75003.1 A=0.096 P=1.58 MULT=1
MM1021 N_A_597_125#_M1021_d N_C1_M1021_g N_A_91_48#_M1015_s VNB NLOWVT L=0.15
+ W=0.64 AD=0.112 AS=0.0896 PD=0.99 PS=0.92 NRD=13.116 NRS=0 M=1 R=4.26667
+ SA=75001.1 SB=75002.7 A=0.096 P=1.58 MULT=1
MM1020 N_A_510_125#_M1020_d N_B1_M1020_g N_A_597_125#_M1021_d VNB NLOWVT L=0.15
+ W=0.64 AD=0.1152 AS=0.112 PD=1 PS=0.99 NRD=0 NRS=0 M=1 R=4.26667 SA=75001.6
+ SB=75002.2 A=0.096 P=1.58 MULT=1
MM1011 N_VGND_M1011_d N_A1_M1011_g N_A_510_125#_M1020_d VNB NLOWVT L=0.15 W=0.64
+ AD=0.0992 AS=0.1152 PD=0.95 PS=1 NRD=0.936 NRS=14.988 M=1 R=4.26667 SA=75002.1
+ SB=75001.7 A=0.096 P=1.58 MULT=1
MM1003 N_A_510_125#_M1003_d N_A2_M1003_g N_VGND_M1011_d VNB NLOWVT L=0.15 W=0.64
+ AD=0.1072 AS=0.0992 PD=0.975 PS=0.95 NRD=10.308 NRS=4.68 M=1 R=4.26667
+ SA=75002.5 SB=75001.2 A=0.096 P=1.58 MULT=1
MM1022 N_A_510_125#_M1003_d N_A2_M1022_g N_VGND_M1022_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.1072 AS=0.112 PD=0.975 PS=0.99 NRD=0 NRS=0 M=1 R=4.26667 SA=75003
+ SB=75000.7 A=0.096 P=1.58 MULT=1
MM1023 N_VGND_M1022_s N_A1_M1023_g N_A_510_125#_M1023_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.112 AS=0.1824 PD=0.99 PS=1.85 NRD=13.116 NRS=0 M=1 R=4.26667 SA=75003.5
+ SB=75000.2 A=0.096 P=1.58 MULT=1
MM1007 N_X_M1007_d N_A_91_48#_M1007_g N_VPWR_M1007_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.3864 PD=1.42 PS=2.93 NRD=1.7533 NRS=10.5395 M=1 R=7.46667
+ SA=75000.3 SB=75004.8 A=0.168 P=2.54 MULT=1
MM1009 N_X_M1007_d N_A_91_48#_M1009_g N_VPWR_M1009_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.224 PD=1.42 PS=1.52 NRD=1.7533 NRS=10.5395 M=1 R=7.46667
+ SA=75000.7 SB=75004.4 A=0.168 P=2.54 MULT=1
MM1010 N_X_M1010_d N_A_91_48#_M1010_g N_VPWR_M1009_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.224 PD=1.42 PS=1.52 NRD=1.7533 NRS=10.5395 M=1 R=7.46667
+ SA=75001.3 SB=75003.8 A=0.168 P=2.54 MULT=1
MM1012 N_X_M1010_d N_A_91_48#_M1012_g N_VPWR_M1012_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.318743 PD=1.42 PS=1.92 NRD=1.7533 NRS=10.5395 M=1 R=7.46667
+ SA=75001.7 SB=75003.4 A=0.168 P=2.54 MULT=1
MM1002 N_A_91_48#_M1002_d N_B1_M1002_g N_VPWR_M1012_s VPB PSHORT L=0.15 W=0.84
+ AD=0.126 AS=0.239057 PD=1.14 PS=1.44 NRD=2.3443 NRS=52.1656 M=1 R=5.6
+ SA=75002.4 SB=75003.7 A=0.126 P=1.98 MULT=1
MM1005 N_VPWR_M1005_d N_C1_M1005_g N_A_91_48#_M1002_d VPB PSHORT L=0.15 W=0.84
+ AD=0.1743 AS=0.126 PD=1.255 PS=1.14 NRD=14.0658 NRS=2.3443 M=1 R=5.6
+ SA=75002.9 SB=75003.3 A=0.126 P=1.98 MULT=1
MM1018 N_VPWR_M1005_d N_C1_M1018_g N_A_91_48#_M1018_s VPB PSHORT L=0.15 W=0.84
+ AD=0.1743 AS=0.126 PD=1.255 PS=1.14 NRD=17.5724 NRS=2.3443 M=1 R=5.6
+ SA=75003.4 SB=75002.7 A=0.126 P=1.98 MULT=1
MM1019 N_A_91_48#_M1018_s N_B1_M1019_g N_VPWR_M1019_s VPB PSHORT L=0.15 W=0.84
+ AD=0.126 AS=0.192013 PD=1.14 PS=1.31022 NRD=2.3443 NRS=22.852 M=1 R=5.6
+ SA=75003.9 SB=75002.3 A=0.126 P=1.98 MULT=1
MM1001 N_A_968_391#_M1001_d N_A1_M1001_g N_VPWR_M1019_s VPB PSHORT L=0.15 W=1
+ AD=0.15 AS=0.228587 PD=1.3 PS=1.55978 NRD=1.9503 NRS=11.8003 M=1 R=6.66667
+ SA=75003.8 SB=75001.7 A=0.15 P=2.3 MULT=1
MM1004 N_A_968_391#_M1001_d N_A2_M1004_g N_A_91_48#_M1004_s VPB PSHORT L=0.15
+ W=1 AD=0.15 AS=0.175 PD=1.3 PS=1.35 NRD=1.9503 NRS=11.8003 M=1 R=6.66667
+ SA=75004.3 SB=75001.2 A=0.15 P=2.3 MULT=1
MM1006 N_A_968_391#_M1006_d N_A2_M1006_g N_A_91_48#_M1004_s VPB PSHORT L=0.15
+ W=1 AD=0.15 AS=0.175 PD=1.3 PS=1.35 NRD=1.9503 NRS=1.9503 M=1 R=6.66667
+ SA=75004.8 SB=75000.7 A=0.15 P=2.3 MULT=1
MM1008 N_A_968_391#_M1006_d N_A1_M1008_g N_VPWR_M1008_s VPB PSHORT L=0.15 W=1
+ AD=0.15 AS=0.345 PD=1.3 PS=2.69 NRD=1.9503 NRS=11.8003 M=1 R=6.66667
+ SA=75005.2 SB=75000.3 A=0.15 P=2.3 MULT=1
DX24_noxref VNB VPB NWDIODE A=13.206 P=17.92
*
.include "sky130_fd_sc_hs__o211a_4.pxi.spice"
*
.ends
*
*
