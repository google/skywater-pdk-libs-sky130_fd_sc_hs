* File: sky130_fd_sc_hs__xor2_2.spice
* Created: Tue Sep  1 20:25:54 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hs__xor2_2.pex.spice"
.subckt sky130_fd_sc_hs__xor2_2  VNB VPB A B VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* B	B
* A	A
* VPB	VPB
* VNB	VNB
MM1004 N_A_183_74#_M1004_d N_A_M1004_g N_VGND_M1004_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.0896 AS=0.5031 PD=0.92 PS=2.9 NRD=0 NRS=137.076 M=1 R=4.26667 SA=75000.6
+ SB=75003.7 A=0.096 P=1.58 MULT=1
MM1000 N_VGND_M1000_d N_B_M1000_g N_A_183_74#_M1004_d VNB NLOWVT L=0.15 W=0.64
+ AD=0.16 AS=0.0896 PD=1.15014 PS=0.92 NRD=13.116 NRS=0 M=1 R=4.26667 SA=75001
+ SB=75003.2 A=0.096 P=1.58 MULT=1
MM1002 N_A_399_74#_M1002_d N_A_M1002_g N_VGND_M1000_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.185 PD=1.02 PS=1.32986 NRD=0 NRS=24.324 M=1 R=4.93333
+ SA=75001.4 SB=75002.6 A=0.111 P=1.78 MULT=1
MM1009 N_A_399_74#_M1002_d N_A_M1009_g N_VGND_M1009_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.3156 PD=1.02 PS=1.7 NRD=0 NRS=60.24 M=1 R=4.93333 SA=75001.9
+ SB=75002.2 A=0.111 P=1.78 MULT=1
MM1014 N_X_M1014_d N_A_183_74#_M1014_g N_VGND_M1009_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.3156 PD=1.02 PS=1.7 NRD=0 NRS=60.24 M=1 R=4.93333 SA=75002.8
+ SB=75001.2 A=0.111 P=1.78 MULT=1
MM1001 N_X_M1014_d N_B_M1001_g N_A_399_74#_M1001_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1794 PD=1.02 PS=1.285 NRD=0 NRS=13.776 M=1 R=4.93333 SA=75003.2
+ SB=75000.8 A=0.111 P=1.78 MULT=1
MM1005 N_X_M1005_d N_B_M1005_g N_A_399_74#_M1001_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.1794 PD=2.05 PS=1.285 NRD=0 NRS=14.592 M=1 R=4.93333 SA=75003.8
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1003 A_116_392# N_A_M1003_g N_VPWR_M1003_s VPB PSHORT L=0.15 W=1 AD=0.135
+ AS=0.295 PD=1.27 PS=2.59 NRD=15.7403 NRS=1.9503 M=1 R=6.66667 SA=75000.2
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1013 N_A_183_74#_M1013_d N_B_M1013_g A_116_392# VPB PSHORT L=0.15 W=1 AD=0.295
+ AS=0.135 PD=2.59 PS=1.27 NRD=1.9503 NRS=15.7403 M=1 R=6.66667 SA=75000.6
+ SB=75000.2 A=0.15 P=2.3 MULT=1
MM1006 N_A_313_368#_M1006_d N_A_M1006_g N_VPWR_M1006_s VPB PSHORT L=0.15 W=1.12
+ AD=0.3304 AS=0.196 PD=2.83 PS=1.47 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75002.6 A=0.168 P=2.54 MULT=1
MM1007 N_A_313_368#_M1007_d N_A_M1007_g N_VPWR_M1006_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.196 PD=1.42 PS=1.47 NRD=1.7533 NRS=10.5395 M=1 R=7.46667
+ SA=75000.7 SB=75002.1 A=0.168 P=2.54 MULT=1
MM1008 N_X_M1008_d N_A_183_74#_M1008_g N_A_313_368#_M1007_d VPB PSHORT L=0.15
+ W=1.12 AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.2 SB=75001.6 A=0.168 P=2.54 MULT=1
MM1010 N_X_M1008_d N_A_183_74#_M1010_g N_A_313_368#_M1010_s VPB PSHORT L=0.15
+ W=1.12 AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.6 SB=75001.2 A=0.168 P=2.54 MULT=1
MM1011 N_A_313_368#_M1010_s N_B_M1011_g N_VPWR_M1011_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.196 PD=1.42 PS=1.47 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75002.1 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1012 N_A_313_368#_M1012_d N_B_M1012_g N_VPWR_M1011_s VPB PSHORT L=0.15 W=1.12
+ AD=0.3416 AS=0.196 PD=2.85 PS=1.47 NRD=2.6201 NRS=10.5395 M=1 R=7.46667
+ SA=75002.6 SB=75000.2 A=0.168 P=2.54 MULT=1
DX15_noxref VNB VPB NWDIODE A=9.6348 P=14.08
*
.include "sky130_fd_sc_hs__xor2_2.pxi.spice"
*
.ends
*
*
