* File: sky130_fd_sc_hs__a21o_4.pxi.spice
* Created: Thu Aug 27 20:25:02 2020
* 
x_PM_SKY130_FD_SC_HS__A21O_4%A_91_48# N_A_91_48#_M1011_d N_A_91_48#_M1009_s
+ N_A_91_48#_M1000_s N_A_91_48#_M1006_g N_A_91_48#_c_120_n N_A_91_48#_M1002_g
+ N_A_91_48#_M1010_g N_A_91_48#_c_121_n N_A_91_48#_M1004_g N_A_91_48#_M1012_g
+ N_A_91_48#_c_122_n N_A_91_48#_M1018_g N_A_91_48#_M1013_g N_A_91_48#_c_123_n
+ N_A_91_48#_M1019_g N_A_91_48#_c_172_p N_A_91_48#_c_112_n N_A_91_48#_c_113_n
+ N_A_91_48#_c_114_n N_A_91_48#_c_115_n N_A_91_48#_c_116_n N_A_91_48#_c_117_n
+ N_A_91_48#_c_118_n N_A_91_48#_c_119_n PM_SKY130_FD_SC_HS__A21O_4%A_91_48#
x_PM_SKY130_FD_SC_HS__A21O_4%B1 N_B1_M1011_g N_B1_M1017_g N_B1_c_244_n
+ N_B1_M1000_g N_B1_c_245_n N_B1_M1016_g B1 N_B1_c_243_n
+ PM_SKY130_FD_SC_HS__A21O_4%B1
x_PM_SKY130_FD_SC_HS__A21O_4%A1 N_A1_c_296_n N_A1_M1003_g N_A1_M1009_g
+ N_A1_c_297_n N_A1_M1005_g N_A1_M1015_g A1 A1 N_A1_c_295_n
+ PM_SKY130_FD_SC_HS__A21O_4%A1
x_PM_SKY130_FD_SC_HS__A21O_4%A2 N_A2_c_351_n N_A2_c_358_n N_A2_M1007_g
+ N_A2_M1001_g N_A2_c_353_n N_A2_c_360_n N_A2_M1008_g N_A2_M1014_g A2
+ N_A2_c_355_n N_A2_c_356_n PM_SKY130_FD_SC_HS__A21O_4%A2
x_PM_SKY130_FD_SC_HS__A21O_4%VPWR N_VPWR_M1002_s N_VPWR_M1004_s N_VPWR_M1019_s
+ N_VPWR_M1003_d N_VPWR_M1007_d N_VPWR_c_400_n N_VPWR_c_401_n N_VPWR_c_402_n
+ N_VPWR_c_403_n N_VPWR_c_404_n N_VPWR_c_405_n N_VPWR_c_406_n N_VPWR_c_407_n
+ N_VPWR_c_408_n N_VPWR_c_409_n VPWR N_VPWR_c_410_n N_VPWR_c_411_n
+ N_VPWR_c_412_n N_VPWR_c_399_n N_VPWR_c_414_n N_VPWR_c_415_n
+ PM_SKY130_FD_SC_HS__A21O_4%VPWR
x_PM_SKY130_FD_SC_HS__A21O_4%X N_X_M1006_d N_X_M1012_d N_X_M1002_d N_X_M1018_d
+ N_X_c_484_n N_X_c_485_n N_X_c_491_n N_X_c_492_n N_X_c_486_n N_X_c_493_n
+ N_X_c_487_n N_X_c_494_n N_X_c_488_n N_X_c_495_n N_X_c_489_n N_X_c_496_n X X
+ PM_SKY130_FD_SC_HS__A21O_4%X
x_PM_SKY130_FD_SC_HS__A21O_4%A_503_392# N_A_503_392#_M1000_d
+ N_A_503_392#_M1016_d N_A_503_392#_M1005_s N_A_503_392#_M1008_s
+ N_A_503_392#_c_559_n N_A_503_392#_c_560_n N_A_503_392#_c_561_n
+ N_A_503_392#_c_562_n N_A_503_392#_c_574_n N_A_503_392#_c_563_n
+ N_A_503_392#_c_564_n N_A_503_392#_c_565_n N_A_503_392#_c_566_n
+ N_A_503_392#_c_567_n N_A_503_392#_c_568_n
+ PM_SKY130_FD_SC_HS__A21O_4%A_503_392#
x_PM_SKY130_FD_SC_HS__A21O_4%VGND N_VGND_M1006_s N_VGND_M1010_s N_VGND_M1013_s
+ N_VGND_M1017_s N_VGND_M1001_s N_VGND_c_619_n N_VGND_c_620_n N_VGND_c_621_n
+ N_VGND_c_622_n N_VGND_c_623_n N_VGND_c_624_n N_VGND_c_625_n N_VGND_c_626_n
+ N_VGND_c_627_n N_VGND_c_628_n N_VGND_c_629_n N_VGND_c_630_n N_VGND_c_631_n
+ N_VGND_c_632_n VGND N_VGND_c_633_n N_VGND_c_634_n
+ PM_SKY130_FD_SC_HS__A21O_4%VGND
x_PM_SKY130_FD_SC_HS__A21O_4%A_700_74# N_A_700_74#_M1009_d N_A_700_74#_M1015_d
+ N_A_700_74#_M1014_d N_A_700_74#_c_706_n N_A_700_74#_c_707_n
+ N_A_700_74#_c_708_n N_A_700_74#_c_709_n N_A_700_74#_c_710_n
+ N_A_700_74#_c_711_n PM_SKY130_FD_SC_HS__A21O_4%A_700_74#
cc_1 VNB N_A_91_48#_M1006_g 0.0232962f $X=-0.19 $Y=-0.245 $X2=0.53 $Y2=0.74
cc_2 VNB N_A_91_48#_M1010_g 0.0203425f $X=-0.19 $Y=-0.245 $X2=0.96 $Y2=0.74
cc_3 VNB N_A_91_48#_M1012_g 0.0209206f $X=-0.19 $Y=-0.245 $X2=1.39 $Y2=0.74
cc_4 VNB N_A_91_48#_M1013_g 0.0218034f $X=-0.19 $Y=-0.245 $X2=1.82 $Y2=0.74
cc_5 VNB N_A_91_48#_c_112_n 0.102873f $X=-0.19 $Y=-0.245 $X2=1.82 $Y2=1.465
cc_6 VNB N_A_91_48#_c_113_n 0.00241395f $X=-0.19 $Y=-0.245 $X2=2.525 $Y2=0.615
cc_7 VNB N_A_91_48#_c_114_n 0.00154126f $X=-0.19 $Y=-0.245 $X2=2.925 $Y2=1.18
cc_8 VNB N_A_91_48#_c_115_n 0.0114549f $X=-0.19 $Y=-0.245 $X2=2.61 $Y2=1.18
cc_9 VNB N_A_91_48#_c_116_n 0.00371113f $X=-0.19 $Y=-0.245 $X2=3.09 $Y2=2.125
cc_10 VNB N_A_91_48#_c_117_n 0.0214012f $X=-0.19 $Y=-0.245 $X2=3.96 $Y2=1.195
cc_11 VNB N_A_91_48#_c_118_n 9.35553e-19 $X=-0.19 $Y=-0.245 $X2=4.055 $Y2=0.76
cc_12 VNB N_A_91_48#_c_119_n 0.00779066f $X=-0.19 $Y=-0.245 $X2=3.09 $Y2=1.187
cc_13 VNB N_B1_M1011_g 0.026748f $X=-0.19 $Y=-0.245 $X2=2.94 $Y2=1.96
cc_14 VNB N_B1_M1017_g 0.0303227f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB B1 9.26387e-19 $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=2.4
cc_16 VNB N_B1_c_243_n 0.0554872f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=2.4
cc_17 VNB N_A1_M1009_g 0.0405164f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A1_M1015_g 0.0321769f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB A1 0.00321331f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=2.4
cc_20 VNB N_A1_c_295_n 0.0271216f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=2.4
cc_21 VNB N_A2_c_351_n 0.00308223f $X=-0.19 $Y=-0.245 $X2=3.915 $Y2=0.37
cc_22 VNB N_A2_M1001_g 0.0233845f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A2_c_353_n 0.00578684f $X=-0.19 $Y=-0.245 $X2=0.53 $Y2=0.74
cc_24 VNB N_A2_M1014_g 0.0324492f $X=-0.19 $Y=-0.245 $X2=0.96 $Y2=1.3
cc_25 VNB N_A2_c_355_n 0.00608101f $X=-0.19 $Y=-0.245 $X2=1.39 $Y2=0.74
cc_26 VNB N_A2_c_356_n 0.0503315f $X=-0.19 $Y=-0.245 $X2=1.445 $Y2=1.765
cc_27 VNB N_VPWR_c_399_n 0.243291f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=1.532
cc_28 VNB N_X_c_484_n 0.00218177f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_X_c_485_n 0.00852127f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=1.765
cc_30 VNB N_X_c_486_n 0.00178908f $X=-0.19 $Y=-0.245 $X2=0.96 $Y2=0.74
cc_31 VNB N_X_c_487_n 0.00467065f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_X_c_488_n 0.00206666f $X=-0.19 $Y=-0.245 $X2=1.82 $Y2=0.74
cc_33 VNB N_X_c_489_n 0.00127131f $X=-0.19 $Y=-0.245 $X2=1.82 $Y2=1.465
cc_34 VNB X 0.0268863f $X=-0.19 $Y=-0.245 $X2=1.82 $Y2=1.465
cc_35 VNB N_VGND_c_619_n 0.0131437f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=2.4
cc_36 VNB N_VGND_c_620_n 0.0253865f $X=-0.19 $Y=-0.245 $X2=0.96 $Y2=0.74
cc_37 VNB N_VGND_c_621_n 0.0040939f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=2.4
cc_38 VNB N_VGND_c_622_n 0.00500784f $X=-0.19 $Y=-0.245 $X2=1.39 $Y2=0.74
cc_39 VNB N_VGND_c_623_n 0.0150374f $X=-0.19 $Y=-0.245 $X2=1.445 $Y2=2.4
cc_40 VNB N_VGND_c_624_n 0.00396467f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_625_n 0.0151736f $X=-0.19 $Y=-0.245 $X2=1.895 $Y2=2.4
cc_42 VNB N_VGND_c_626_n 0.00461913f $X=-0.19 $Y=-0.245 $X2=1.87 $Y2=1.465
cc_43 VNB N_VGND_c_627_n 0.0172524f $X=-0.19 $Y=-0.245 $X2=0.8 $Y2=1.465
cc_44 VNB N_VGND_c_628_n 0.00461913f $X=-0.19 $Y=-0.245 $X2=0.8 $Y2=1.465
cc_45 VNB N_VGND_c_629_n 0.0196652f $X=-0.19 $Y=-0.245 $X2=1.82 $Y2=1.465
cc_46 VNB N_VGND_c_630_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=1.82 $Y2=1.465
cc_47 VNB N_VGND_c_631_n 0.0409245f $X=-0.19 $Y=-0.245 $X2=2.485 $Y2=1.095
cc_48 VNB N_VGND_c_632_n 0.00604233f $X=-0.19 $Y=-0.245 $X2=2.485 $Y2=0.615
cc_49 VNB N_VGND_c_633_n 0.0216869f $X=-0.19 $Y=-0.245 $X2=0.96 $Y2=1.532
cc_50 VNB N_VGND_c_634_n 0.347716f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=1.532
cc_51 VNB N_A_700_74#_c_706_n 0.00629727f $X=-0.19 $Y=-0.245 $X2=0.53 $Y2=0.74
cc_52 VNB N_A_700_74#_c_707_n 0.00449328f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=1.765
cc_53 VNB N_A_700_74#_c_708_n 0.00473324f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=2.4
cc_54 VNB N_A_700_74#_c_709_n 0.0244999f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_A_700_74#_c_710_n 0.0036276f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=1.765
cc_56 VNB N_A_700_74#_c_711_n 0.0237116f $X=-0.19 $Y=-0.245 $X2=1.39 $Y2=1.3
cc_57 VPB N_A_91_48#_c_120_n 0.0172602f $X=-0.19 $Y=1.66 $X2=0.545 $Y2=1.765
cc_58 VPB N_A_91_48#_c_121_n 0.014716f $X=-0.19 $Y=1.66 $X2=0.995 $Y2=1.765
cc_59 VPB N_A_91_48#_c_122_n 0.015247f $X=-0.19 $Y=1.66 $X2=1.445 $Y2=1.765
cc_60 VPB N_A_91_48#_c_123_n 0.0178158f $X=-0.19 $Y=1.66 $X2=1.895 $Y2=1.765
cc_61 VPB N_A_91_48#_c_112_n 0.0263702f $X=-0.19 $Y=1.66 $X2=1.82 $Y2=1.465
cc_62 VPB N_B1_c_244_n 0.018172f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_63 VPB N_B1_c_245_n 0.0145904f $X=-0.19 $Y=1.66 $X2=0.53 $Y2=0.74
cc_64 VPB B1 0.00558514f $X=-0.19 $Y=1.66 $X2=0.545 $Y2=2.4
cc_65 VPB N_B1_c_243_n 0.0621522f $X=-0.19 $Y=1.66 $X2=0.995 $Y2=2.4
cc_66 VPB N_A1_c_296_n 0.0152645f $X=-0.19 $Y=1.66 $X2=2.385 $Y2=0.47
cc_67 VPB N_A1_c_297_n 0.0157745f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_68 VPB A1 0.00258732f $X=-0.19 $Y=1.66 $X2=0.545 $Y2=2.4
cc_69 VPB N_A1_c_295_n 0.0317718f $X=-0.19 $Y=1.66 $X2=0.995 $Y2=2.4
cc_70 VPB N_A2_c_351_n 0.00614586f $X=-0.19 $Y=1.66 $X2=3.915 $Y2=0.37
cc_71 VPB N_A2_c_358_n 0.0209822f $X=-0.19 $Y=1.66 $X2=2.94 $Y2=1.96
cc_72 VPB N_A2_c_353_n 0.0112418f $X=-0.19 $Y=1.66 $X2=0.53 $Y2=0.74
cc_73 VPB N_A2_c_360_n 0.0281896f $X=-0.19 $Y=1.66 $X2=0.53 $Y2=0.74
cc_74 VPB N_A2_c_355_n 0.00467294f $X=-0.19 $Y=1.66 $X2=1.39 $Y2=0.74
cc_75 VPB N_VPWR_c_400_n 0.0132865f $X=-0.19 $Y=1.66 $X2=0.545 $Y2=2.4
cc_76 VPB N_VPWR_c_401_n 0.0415304f $X=-0.19 $Y=1.66 $X2=0.96 $Y2=0.74
cc_77 VPB N_VPWR_c_402_n 0.00504372f $X=-0.19 $Y=1.66 $X2=0.995 $Y2=2.4
cc_78 VPB N_VPWR_c_403_n 0.0182622f $X=-0.19 $Y=1.66 $X2=1.39 $Y2=0.74
cc_79 VPB N_VPWR_c_404_n 0.00501395f $X=-0.19 $Y=1.66 $X2=1.82 $Y2=0.74
cc_80 VPB N_VPWR_c_405_n 0.00339119f $X=-0.19 $Y=1.66 $X2=1.895 $Y2=2.4
cc_81 VPB N_VPWR_c_406_n 0.0376948f $X=-0.19 $Y=1.66 $X2=0.8 $Y2=1.465
cc_82 VPB N_VPWR_c_407_n 0.00460249f $X=-0.19 $Y=1.66 $X2=0.8 $Y2=1.465
cc_83 VPB N_VPWR_c_408_n 0.0185253f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_84 VPB N_VPWR_c_409_n 0.00601644f $X=-0.19 $Y=1.66 $X2=1.82 $Y2=1.465
cc_85 VPB N_VPWR_c_410_n 0.0164465f $X=-0.19 $Y=1.66 $X2=2.485 $Y2=1.095
cc_86 VPB N_VPWR_c_411_n 0.0206041f $X=-0.19 $Y=1.66 $X2=2.61 $Y2=1.18
cc_87 VPB N_VPWR_c_412_n 0.0224824f $X=-0.19 $Y=1.66 $X2=0.96 $Y2=1.532
cc_88 VPB N_VPWR_c_399_n 0.095301f $X=-0.19 $Y=1.66 $X2=0.995 $Y2=1.532
cc_89 VPB N_VPWR_c_414_n 0.00460249f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_90 VPB N_VPWR_c_415_n 0.0047828f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_91 VPB N_X_c_491_n 0.00205681f $X=-0.19 $Y=1.66 $X2=0.545 $Y2=2.4
cc_92 VPB N_X_c_492_n 0.00909169f $X=-0.19 $Y=1.66 $X2=0.545 $Y2=2.4
cc_93 VPB N_X_c_493_n 0.00180921f $X=-0.19 $Y=1.66 $X2=0.995 $Y2=2.4
cc_94 VPB N_X_c_494_n 0.00401098f $X=-0.19 $Y=1.66 $X2=1.445 $Y2=2.4
cc_95 VPB N_X_c_495_n 0.00257348f $X=-0.19 $Y=1.66 $X2=1.895 $Y2=2.4
cc_96 VPB N_X_c_496_n 0.00104376f $X=-0.19 $Y=1.66 $X2=1.82 $Y2=1.465
cc_97 VPB X 0.00713242f $X=-0.19 $Y=1.66 $X2=1.82 $Y2=1.465
cc_98 VPB N_A_503_392#_c_559_n 0.0101892f $X=-0.19 $Y=1.66 $X2=0.545 $Y2=2.4
cc_99 VPB N_A_503_392#_c_560_n 0.00523584f $X=-0.19 $Y=1.66 $X2=0.96 $Y2=0.74
cc_100 VPB N_A_503_392#_c_561_n 0.00376819f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_101 VPB N_A_503_392#_c_562_n 0.00191281f $X=-0.19 $Y=1.66 $X2=0.995 $Y2=1.765
cc_102 VPB N_A_503_392#_c_563_n 0.00233322f $X=-0.19 $Y=1.66 $X2=1.39 $Y2=0.74
cc_103 VPB N_A_503_392#_c_564_n 0.00216998f $X=-0.19 $Y=1.66 $X2=1.445 $Y2=2.4
cc_104 VPB N_A_503_392#_c_565_n 0.00723758f $X=-0.19 $Y=1.66 $X2=1.82 $Y2=1.3
cc_105 VPB N_A_503_392#_c_566_n 0.0178982f $X=-0.19 $Y=1.66 $X2=1.82 $Y2=0.74
cc_106 VPB N_A_503_392#_c_567_n 0.0345863f $X=-0.19 $Y=1.66 $X2=1.895 $Y2=1.765
cc_107 VPB N_A_503_392#_c_568_n 0.00554471f $X=-0.19 $Y=1.66 $X2=0.8 $Y2=1.465
cc_108 N_A_91_48#_M1013_g N_B1_M1011_g 0.0237775f $X=1.82 $Y=0.74 $X2=0 $Y2=0
cc_109 N_A_91_48#_c_112_n N_B1_M1011_g 0.0246033f $X=1.82 $Y=1.465 $X2=0 $Y2=0
cc_110 N_A_91_48#_c_113_n N_B1_M1011_g 0.00945691f $X=2.525 $Y=0.615 $X2=0 $Y2=0
cc_111 N_A_91_48#_c_115_n N_B1_M1011_g 0.0260214f $X=2.61 $Y=1.18 $X2=0 $Y2=0
cc_112 N_A_91_48#_c_114_n N_B1_M1017_g 0.0178404f $X=2.925 $Y=1.18 $X2=0 $Y2=0
cc_113 N_A_91_48#_c_116_n N_B1_M1017_g 0.00609733f $X=3.09 $Y=2.125 $X2=0 $Y2=0
cc_114 N_A_91_48#_c_119_n N_B1_M1017_g 6.5814e-19 $X=3.09 $Y=1.187 $X2=0 $Y2=0
cc_115 N_A_91_48#_c_116_n N_B1_c_244_n 0.0129727f $X=3.09 $Y=2.125 $X2=0 $Y2=0
cc_116 N_A_91_48#_c_116_n N_B1_c_245_n 0.0109026f $X=3.09 $Y=2.125 $X2=0 $Y2=0
cc_117 N_A_91_48#_c_123_n B1 3.99641e-19 $X=1.895 $Y=1.765 $X2=0 $Y2=0
cc_118 N_A_91_48#_c_112_n B1 7.3424e-19 $X=1.82 $Y=1.465 $X2=0 $Y2=0
cc_119 N_A_91_48#_c_114_n B1 0.010543f $X=2.925 $Y=1.18 $X2=0 $Y2=0
cc_120 N_A_91_48#_c_115_n B1 0.029196f $X=2.61 $Y=1.18 $X2=0 $Y2=0
cc_121 N_A_91_48#_c_116_n B1 0.0259517f $X=3.09 $Y=2.125 $X2=0 $Y2=0
cc_122 N_A_91_48#_c_114_n N_B1_c_243_n 0.00454834f $X=2.925 $Y=1.18 $X2=0 $Y2=0
cc_123 N_A_91_48#_c_115_n N_B1_c_243_n 7.91474e-19 $X=2.61 $Y=1.18 $X2=0 $Y2=0
cc_124 N_A_91_48#_c_116_n N_B1_c_243_n 0.0422113f $X=3.09 $Y=2.125 $X2=0 $Y2=0
cc_125 N_A_91_48#_c_117_n N_B1_c_243_n 0.00627271f $X=3.96 $Y=1.195 $X2=0 $Y2=0
cc_126 N_A_91_48#_c_116_n N_A1_c_296_n 3.61165e-19 $X=3.09 $Y=2.125 $X2=-0.19
+ $Y2=-0.245
cc_127 N_A_91_48#_c_116_n N_A1_M1009_g 0.00407816f $X=3.09 $Y=2.125 $X2=0 $Y2=0
cc_128 N_A_91_48#_c_117_n N_A1_M1009_g 0.0163803f $X=3.96 $Y=1.195 $X2=0 $Y2=0
cc_129 N_A_91_48#_c_118_n N_A1_M1009_g 0.00281396f $X=4.055 $Y=0.76 $X2=0 $Y2=0
cc_130 N_A_91_48#_c_119_n N_A1_M1009_g 4.3183e-19 $X=3.09 $Y=1.187 $X2=0 $Y2=0
cc_131 N_A_91_48#_c_117_n N_A1_M1015_g 0.00597757f $X=3.96 $Y=1.195 $X2=0 $Y2=0
cc_132 N_A_91_48#_c_118_n N_A1_M1015_g 0.00720134f $X=4.055 $Y=0.76 $X2=0 $Y2=0
cc_133 N_A_91_48#_c_116_n A1 0.0221389f $X=3.09 $Y=2.125 $X2=0 $Y2=0
cc_134 N_A_91_48#_c_117_n A1 0.0557184f $X=3.96 $Y=1.195 $X2=0 $Y2=0
cc_135 N_A_91_48#_c_116_n N_A1_c_295_n 7.56267e-19 $X=3.09 $Y=2.125 $X2=0 $Y2=0
cc_136 N_A_91_48#_c_117_n N_A1_c_295_n 0.0046592f $X=3.96 $Y=1.195 $X2=0 $Y2=0
cc_137 N_A_91_48#_c_117_n N_A2_M1001_g 7.22688e-19 $X=3.96 $Y=1.195 $X2=0 $Y2=0
cc_138 N_A_91_48#_c_117_n N_A2_c_355_n 0.00139372f $X=3.96 $Y=1.195 $X2=0 $Y2=0
cc_139 N_A_91_48#_c_120_n N_VPWR_c_401_n 0.0176265f $X=0.545 $Y=1.765 $X2=0
+ $Y2=0
cc_140 N_A_91_48#_c_121_n N_VPWR_c_401_n 5.81581e-19 $X=0.995 $Y=1.765 $X2=0
+ $Y2=0
cc_141 N_A_91_48#_c_120_n N_VPWR_c_402_n 5.83721e-19 $X=0.545 $Y=1.765 $X2=0
+ $Y2=0
cc_142 N_A_91_48#_c_121_n N_VPWR_c_402_n 0.0133451f $X=0.995 $Y=1.765 $X2=0
+ $Y2=0
cc_143 N_A_91_48#_c_122_n N_VPWR_c_402_n 0.00630489f $X=1.445 $Y=1.765 $X2=0
+ $Y2=0
cc_144 N_A_91_48#_c_123_n N_VPWR_c_403_n 0.00831688f $X=1.895 $Y=1.765 $X2=0
+ $Y2=0
cc_145 N_A_91_48#_c_115_n N_VPWR_c_403_n 0.00967443f $X=2.61 $Y=1.18 $X2=0 $Y2=0
cc_146 N_A_91_48#_c_120_n N_VPWR_c_410_n 0.00413917f $X=0.545 $Y=1.765 $X2=0
+ $Y2=0
cc_147 N_A_91_48#_c_121_n N_VPWR_c_410_n 0.00413917f $X=0.995 $Y=1.765 $X2=0
+ $Y2=0
cc_148 N_A_91_48#_c_122_n N_VPWR_c_411_n 0.00445602f $X=1.445 $Y=1.765 $X2=0
+ $Y2=0
cc_149 N_A_91_48#_c_123_n N_VPWR_c_411_n 0.00445602f $X=1.895 $Y=1.765 $X2=0
+ $Y2=0
cc_150 N_A_91_48#_c_120_n N_VPWR_c_399_n 0.00817726f $X=0.545 $Y=1.765 $X2=0
+ $Y2=0
cc_151 N_A_91_48#_c_121_n N_VPWR_c_399_n 0.00817726f $X=0.995 $Y=1.765 $X2=0
+ $Y2=0
cc_152 N_A_91_48#_c_122_n N_VPWR_c_399_n 0.00857589f $X=1.445 $Y=1.765 $X2=0
+ $Y2=0
cc_153 N_A_91_48#_c_123_n N_VPWR_c_399_n 0.00862391f $X=1.895 $Y=1.765 $X2=0
+ $Y2=0
cc_154 N_A_91_48#_M1006_g N_X_c_484_n 0.0161282f $X=0.53 $Y=0.74 $X2=0 $Y2=0
cc_155 N_A_91_48#_c_172_p N_X_c_484_n 0.00184167f $X=1.87 $Y=1.465 $X2=0 $Y2=0
cc_156 N_A_91_48#_c_120_n N_X_c_491_n 0.0167603f $X=0.545 $Y=1.765 $X2=0 $Y2=0
cc_157 N_A_91_48#_c_172_p N_X_c_491_n 0.0037202f $X=1.87 $Y=1.465 $X2=0 $Y2=0
cc_158 N_A_91_48#_c_112_n N_X_c_491_n 0.00243093f $X=1.82 $Y=1.465 $X2=0 $Y2=0
cc_159 N_A_91_48#_M1006_g N_X_c_486_n 3.92313e-19 $X=0.53 $Y=0.74 $X2=0 $Y2=0
cc_160 N_A_91_48#_M1010_g N_X_c_486_n 3.92313e-19 $X=0.96 $Y=0.74 $X2=0 $Y2=0
cc_161 N_A_91_48#_c_120_n N_X_c_493_n 0.00624195f $X=0.545 $Y=1.765 $X2=0 $Y2=0
cc_162 N_A_91_48#_c_121_n N_X_c_493_n 0.00438646f $X=0.995 $Y=1.765 $X2=0 $Y2=0
cc_163 N_A_91_48#_M1010_g N_X_c_487_n 0.0124434f $X=0.96 $Y=0.74 $X2=0 $Y2=0
cc_164 N_A_91_48#_M1012_g N_X_c_487_n 0.0120709f $X=1.39 $Y=0.74 $X2=0 $Y2=0
cc_165 N_A_91_48#_c_172_p N_X_c_487_n 0.0657213f $X=1.87 $Y=1.465 $X2=0 $Y2=0
cc_166 N_A_91_48#_c_112_n N_X_c_487_n 0.00457162f $X=1.82 $Y=1.465 $X2=0 $Y2=0
cc_167 N_A_91_48#_c_115_n N_X_c_487_n 0.00226813f $X=2.61 $Y=1.18 $X2=0 $Y2=0
cc_168 N_A_91_48#_c_121_n N_X_c_494_n 0.0131837f $X=0.995 $Y=1.765 $X2=0 $Y2=0
cc_169 N_A_91_48#_c_122_n N_X_c_494_n 0.0129464f $X=1.445 $Y=1.765 $X2=0 $Y2=0
cc_170 N_A_91_48#_c_123_n N_X_c_494_n 0.00787118f $X=1.895 $Y=1.765 $X2=0 $Y2=0
cc_171 N_A_91_48#_c_172_p N_X_c_494_n 0.0754071f $X=1.87 $Y=1.465 $X2=0 $Y2=0
cc_172 N_A_91_48#_c_112_n N_X_c_494_n 0.0173523f $X=1.82 $Y=1.465 $X2=0 $Y2=0
cc_173 N_A_91_48#_M1010_g N_X_c_488_n 6.20738e-19 $X=0.96 $Y=0.74 $X2=0 $Y2=0
cc_174 N_A_91_48#_M1012_g N_X_c_488_n 0.00866629f $X=1.39 $Y=0.74 $X2=0 $Y2=0
cc_175 N_A_91_48#_M1013_g N_X_c_488_n 3.97481e-19 $X=1.82 $Y=0.74 $X2=0 $Y2=0
cc_176 N_A_91_48#_c_121_n N_X_c_495_n 7.68526e-19 $X=0.995 $Y=1.765 $X2=0 $Y2=0
cc_177 N_A_91_48#_c_122_n N_X_c_495_n 0.012705f $X=1.445 $Y=1.765 $X2=0 $Y2=0
cc_178 N_A_91_48#_c_123_n N_X_c_495_n 0.0118573f $X=1.895 $Y=1.765 $X2=0 $Y2=0
cc_179 N_A_91_48#_c_172_p N_X_c_489_n 0.0143381f $X=1.87 $Y=1.465 $X2=0 $Y2=0
cc_180 N_A_91_48#_c_112_n N_X_c_489_n 0.00232957f $X=1.82 $Y=1.465 $X2=0 $Y2=0
cc_181 N_A_91_48#_c_172_p N_X_c_496_n 0.0143367f $X=1.87 $Y=1.465 $X2=0 $Y2=0
cc_182 N_A_91_48#_c_112_n N_X_c_496_n 0.00423635f $X=1.82 $Y=1.465 $X2=0 $Y2=0
cc_183 N_A_91_48#_M1006_g X 0.0217805f $X=0.53 $Y=0.74 $X2=0 $Y2=0
cc_184 N_A_91_48#_c_120_n X 0.00128081f $X=0.545 $Y=1.765 $X2=0 $Y2=0
cc_185 N_A_91_48#_c_172_p X 0.0184026f $X=1.87 $Y=1.465 $X2=0 $Y2=0
cc_186 N_A_91_48#_c_116_n N_A_503_392#_c_559_n 0.0526499f $X=3.09 $Y=2.125 $X2=0
+ $Y2=0
cc_187 N_A_91_48#_M1000_s N_A_503_392#_c_560_n 0.00197722f $X=2.94 $Y=1.96 $X2=0
+ $Y2=0
cc_188 N_A_91_48#_c_116_n N_A_503_392#_c_560_n 0.0160777f $X=3.09 $Y=2.125 $X2=0
+ $Y2=0
cc_189 N_A_91_48#_c_116_n N_A_503_392#_c_562_n 0.0123997f $X=3.09 $Y=2.125 $X2=0
+ $Y2=0
cc_190 N_A_91_48#_c_117_n N_A_503_392#_c_562_n 9.69132e-19 $X=3.96 $Y=1.195
+ $X2=0 $Y2=0
cc_191 N_A_91_48#_c_116_n N_A_503_392#_c_574_n 0.040027f $X=3.09 $Y=2.125 $X2=0
+ $Y2=0
cc_192 N_A_91_48#_c_117_n N_A_503_392#_c_563_n 6.03499e-19 $X=3.96 $Y=1.195
+ $X2=0 $Y2=0
cc_193 N_A_91_48#_c_115_n N_VGND_M1013_s 0.00442076f $X=2.61 $Y=1.18 $X2=0 $Y2=0
cc_194 N_A_91_48#_c_114_n N_VGND_M1017_s 5.5277e-19 $X=2.925 $Y=1.18 $X2=0 $Y2=0
cc_195 N_A_91_48#_c_119_n N_VGND_M1017_s 0.00178584f $X=3.09 $Y=1.187 $X2=0
+ $Y2=0
cc_196 N_A_91_48#_M1006_g N_VGND_c_620_n 0.0111233f $X=0.53 $Y=0.74 $X2=0 $Y2=0
cc_197 N_A_91_48#_M1010_g N_VGND_c_620_n 4.56715e-19 $X=0.96 $Y=0.74 $X2=0 $Y2=0
cc_198 N_A_91_48#_M1006_g N_VGND_c_621_n 4.57991e-19 $X=0.53 $Y=0.74 $X2=0 $Y2=0
cc_199 N_A_91_48#_M1010_g N_VGND_c_621_n 0.00900784f $X=0.96 $Y=0.74 $X2=0 $Y2=0
cc_200 N_A_91_48#_M1012_g N_VGND_c_621_n 0.00183835f $X=1.39 $Y=0.74 $X2=0 $Y2=0
cc_201 N_A_91_48#_M1012_g N_VGND_c_622_n 5.46162e-19 $X=1.39 $Y=0.74 $X2=0 $Y2=0
cc_202 N_A_91_48#_M1013_g N_VGND_c_622_n 0.0127508f $X=1.82 $Y=0.74 $X2=0 $Y2=0
cc_203 N_A_91_48#_c_112_n N_VGND_c_622_n 3.23166e-19 $X=1.82 $Y=1.465 $X2=0
+ $Y2=0
cc_204 N_A_91_48#_c_113_n N_VGND_c_622_n 0.0271353f $X=2.525 $Y=0.615 $X2=0
+ $Y2=0
cc_205 N_A_91_48#_c_115_n N_VGND_c_622_n 0.0167891f $X=2.61 $Y=1.18 $X2=0 $Y2=0
cc_206 N_A_91_48#_c_113_n N_VGND_c_623_n 0.0177526f $X=2.525 $Y=0.615 $X2=0
+ $Y2=0
cc_207 N_A_91_48#_c_114_n N_VGND_c_623_n 0.00606161f $X=2.925 $Y=1.18 $X2=0
+ $Y2=0
cc_208 N_A_91_48#_c_119_n N_VGND_c_623_n 0.0176293f $X=3.09 $Y=1.187 $X2=0 $Y2=0
cc_209 N_A_91_48#_M1006_g N_VGND_c_625_n 0.00383152f $X=0.53 $Y=0.74 $X2=0 $Y2=0
cc_210 N_A_91_48#_M1010_g N_VGND_c_625_n 0.00383152f $X=0.96 $Y=0.74 $X2=0 $Y2=0
cc_211 N_A_91_48#_M1012_g N_VGND_c_627_n 0.00434272f $X=1.39 $Y=0.74 $X2=0 $Y2=0
cc_212 N_A_91_48#_M1013_g N_VGND_c_627_n 0.00383152f $X=1.82 $Y=0.74 $X2=0 $Y2=0
cc_213 N_A_91_48#_c_113_n N_VGND_c_629_n 0.0078096f $X=2.525 $Y=0.615 $X2=0
+ $Y2=0
cc_214 N_A_91_48#_M1006_g N_VGND_c_634_n 0.0075754f $X=0.53 $Y=0.74 $X2=0 $Y2=0
cc_215 N_A_91_48#_M1010_g N_VGND_c_634_n 0.0075754f $X=0.96 $Y=0.74 $X2=0 $Y2=0
cc_216 N_A_91_48#_M1012_g N_VGND_c_634_n 0.00820284f $X=1.39 $Y=0.74 $X2=0 $Y2=0
cc_217 N_A_91_48#_M1013_g N_VGND_c_634_n 0.0075754f $X=1.82 $Y=0.74 $X2=0 $Y2=0
cc_218 N_A_91_48#_c_113_n N_VGND_c_634_n 0.0085649f $X=2.525 $Y=0.615 $X2=0
+ $Y2=0
cc_219 N_A_91_48#_c_117_n N_A_700_74#_c_706_n 0.0244478f $X=3.96 $Y=1.195 $X2=0
+ $Y2=0
cc_220 N_A_91_48#_M1009_s N_A_700_74#_c_707_n 0.00176461f $X=3.915 $Y=0.37 $X2=0
+ $Y2=0
cc_221 N_A_91_48#_c_118_n N_A_700_74#_c_707_n 0.0143157f $X=4.055 $Y=0.76 $X2=0
+ $Y2=0
cc_222 N_A_91_48#_c_118_n N_A_700_74#_c_710_n 0.0094371f $X=4.055 $Y=0.76 $X2=0
+ $Y2=0
cc_223 N_B1_c_245_n N_A1_c_296_n 0.00793765f $X=3.315 $Y=1.885 $X2=-0.19
+ $Y2=-0.245
cc_224 N_B1_c_243_n N_A1_M1009_g 5.97977e-19 $X=2.865 $Y=1.66 $X2=0 $Y2=0
cc_225 N_B1_c_243_n A1 0.00337577f $X=2.865 $Y=1.66 $X2=0 $Y2=0
cc_226 N_B1_c_243_n N_A1_c_295_n 0.0207279f $X=2.865 $Y=1.66 $X2=0 $Y2=0
cc_227 N_B1_c_244_n N_VPWR_c_403_n 8.45076e-19 $X=2.865 $Y=1.885 $X2=0 $Y2=0
cc_228 N_B1_c_243_n N_VPWR_c_403_n 0.00233281f $X=2.865 $Y=1.66 $X2=0 $Y2=0
cc_229 N_B1_c_244_n N_VPWR_c_406_n 0.00278271f $X=2.865 $Y=1.885 $X2=0 $Y2=0
cc_230 N_B1_c_245_n N_VPWR_c_406_n 0.00278271f $X=3.315 $Y=1.885 $X2=0 $Y2=0
cc_231 N_B1_c_244_n N_VPWR_c_399_n 0.00358624f $X=2.865 $Y=1.885 $X2=0 $Y2=0
cc_232 N_B1_c_245_n N_VPWR_c_399_n 0.00353907f $X=3.315 $Y=1.885 $X2=0 $Y2=0
cc_233 N_B1_c_244_n N_A_503_392#_c_559_n 0.00648664f $X=2.865 $Y=1.885 $X2=0
+ $Y2=0
cc_234 B1 N_A_503_392#_c_559_n 0.0221057f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_235 N_B1_c_243_n N_A_503_392#_c_559_n 0.00186824f $X=2.865 $Y=1.66 $X2=0
+ $Y2=0
cc_236 N_B1_c_244_n N_A_503_392#_c_560_n 0.0136485f $X=2.865 $Y=1.885 $X2=0
+ $Y2=0
cc_237 N_B1_c_245_n N_A_503_392#_c_560_n 0.012504f $X=3.315 $Y=1.885 $X2=0 $Y2=0
cc_238 N_B1_c_245_n N_A_503_392#_c_562_n 7.89448e-19 $X=3.315 $Y=1.885 $X2=0
+ $Y2=0
cc_239 N_B1_M1011_g N_VGND_c_622_n 0.005271f $X=2.31 $Y=0.79 $X2=0 $Y2=0
cc_240 N_B1_M1011_g N_VGND_c_623_n 4.92858e-19 $X=2.31 $Y=0.79 $X2=0 $Y2=0
cc_241 N_B1_M1017_g N_VGND_c_623_n 0.0124783f $X=2.74 $Y=0.79 $X2=0 $Y2=0
cc_242 N_B1_c_243_n N_VGND_c_623_n 8.49409e-19 $X=2.865 $Y=1.66 $X2=0 $Y2=0
cc_243 N_B1_M1011_g N_VGND_c_629_n 0.00485498f $X=2.31 $Y=0.79 $X2=0 $Y2=0
cc_244 N_B1_M1017_g N_VGND_c_629_n 0.00421418f $X=2.74 $Y=0.79 $X2=0 $Y2=0
cc_245 N_B1_M1011_g N_VGND_c_634_n 0.00514438f $X=2.31 $Y=0.79 $X2=0 $Y2=0
cc_246 N_B1_M1017_g N_VGND_c_634_n 0.00432128f $X=2.74 $Y=0.79 $X2=0 $Y2=0
cc_247 N_B1_M1017_g N_A_700_74#_c_706_n 0.00129185f $X=2.74 $Y=0.79 $X2=0 $Y2=0
cc_248 N_B1_M1017_g N_A_700_74#_c_708_n 3.66717e-19 $X=2.74 $Y=0.79 $X2=0 $Y2=0
cc_249 N_A1_c_295_n N_A2_c_351_n 0.0234129f $X=4.215 $Y=1.667 $X2=0 $Y2=0
cc_250 N_A1_c_297_n N_A2_c_358_n 0.00843956f $X=4.215 $Y=1.885 $X2=0 $Y2=0
cc_251 N_A1_M1015_g N_A2_M1001_g 0.0162328f $X=4.27 $Y=0.69 $X2=0 $Y2=0
cc_252 N_A1_M1015_g N_A2_c_355_n 0.00606004f $X=4.27 $Y=0.69 $X2=0 $Y2=0
cc_253 A1 N_A2_c_355_n 0.0211953f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_254 N_A1_c_295_n N_A2_c_355_n 0.00162069f $X=4.215 $Y=1.667 $X2=0 $Y2=0
cc_255 N_A1_M1015_g N_A2_c_356_n 0.00931764f $X=4.27 $Y=0.69 $X2=0 $Y2=0
cc_256 A1 N_A2_c_356_n 2.81306e-19 $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_257 N_A1_c_296_n N_VPWR_c_404_n 0.00996098f $X=3.765 $Y=1.885 $X2=0 $Y2=0
cc_258 N_A1_c_297_n N_VPWR_c_404_n 0.00395359f $X=4.215 $Y=1.885 $X2=0 $Y2=0
cc_259 N_A1_c_297_n N_VPWR_c_405_n 5.55114e-19 $X=4.215 $Y=1.885 $X2=0 $Y2=0
cc_260 N_A1_c_296_n N_VPWR_c_406_n 0.00413917f $X=3.765 $Y=1.885 $X2=0 $Y2=0
cc_261 N_A1_c_297_n N_VPWR_c_408_n 0.00445602f $X=4.215 $Y=1.885 $X2=0 $Y2=0
cc_262 N_A1_c_296_n N_VPWR_c_399_n 0.0081781f $X=3.765 $Y=1.885 $X2=0 $Y2=0
cc_263 N_A1_c_297_n N_VPWR_c_399_n 0.00857673f $X=4.215 $Y=1.885 $X2=0 $Y2=0
cc_264 N_A1_c_296_n N_A_503_392#_c_560_n 0.00125031f $X=3.765 $Y=1.885 $X2=0
+ $Y2=0
cc_265 A1 N_A_503_392#_c_562_n 0.0123846f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_266 N_A1_c_296_n N_A_503_392#_c_563_n 0.0127777f $X=3.765 $Y=1.885 $X2=0
+ $Y2=0
cc_267 N_A1_c_297_n N_A_503_392#_c_563_n 0.0139848f $X=4.215 $Y=1.885 $X2=0
+ $Y2=0
cc_268 A1 N_A_503_392#_c_563_n 0.0422401f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_269 N_A1_c_295_n N_A_503_392#_c_563_n 0.00802096f $X=4.215 $Y=1.667 $X2=0
+ $Y2=0
cc_270 N_A1_c_296_n N_A_503_392#_c_564_n 6.71799e-19 $X=3.765 $Y=1.885 $X2=0
+ $Y2=0
cc_271 N_A1_c_297_n N_A_503_392#_c_564_n 0.0104892f $X=4.215 $Y=1.885 $X2=0
+ $Y2=0
cc_272 N_A1_c_297_n N_A_503_392#_c_568_n 0.00111497f $X=4.215 $Y=1.885 $X2=0
+ $Y2=0
cc_273 N_A1_c_295_n N_A_503_392#_c_568_n 0.00241193f $X=4.215 $Y=1.667 $X2=0
+ $Y2=0
cc_274 N_A1_M1009_g N_VGND_c_623_n 0.00188825f $X=3.84 $Y=0.69 $X2=0 $Y2=0
cc_275 N_A1_M1009_g N_VGND_c_631_n 0.00278247f $X=3.84 $Y=0.69 $X2=0 $Y2=0
cc_276 N_A1_M1015_g N_VGND_c_631_n 0.00278271f $X=4.27 $Y=0.69 $X2=0 $Y2=0
cc_277 N_A1_M1009_g N_VGND_c_634_n 0.00358425f $X=3.84 $Y=0.69 $X2=0 $Y2=0
cc_278 N_A1_M1015_g N_VGND_c_634_n 0.00353526f $X=4.27 $Y=0.69 $X2=0 $Y2=0
cc_279 N_A1_M1009_g N_A_700_74#_c_706_n 0.00697945f $X=3.84 $Y=0.69 $X2=0 $Y2=0
cc_280 N_A1_M1015_g N_A_700_74#_c_706_n 4.5114e-19 $X=4.27 $Y=0.69 $X2=0 $Y2=0
cc_281 N_A1_M1009_g N_A_700_74#_c_707_n 0.0100245f $X=3.84 $Y=0.69 $X2=0 $Y2=0
cc_282 N_A1_M1015_g N_A_700_74#_c_707_n 0.0120041f $X=4.27 $Y=0.69 $X2=0 $Y2=0
cc_283 N_A1_M1009_g N_A_700_74#_c_708_n 0.00281658f $X=3.84 $Y=0.69 $X2=0 $Y2=0
cc_284 N_A1_M1015_g N_A_700_74#_c_710_n 6.58764e-19 $X=4.27 $Y=0.69 $X2=0 $Y2=0
cc_285 N_A2_c_358_n N_VPWR_c_405_n 0.0111578f $X=4.665 $Y=1.885 $X2=0 $Y2=0
cc_286 N_A2_c_360_n N_VPWR_c_405_n 0.0141019f $X=5.115 $Y=1.885 $X2=0 $Y2=0
cc_287 N_A2_c_358_n N_VPWR_c_408_n 0.00413917f $X=4.665 $Y=1.885 $X2=0 $Y2=0
cc_288 N_A2_c_360_n N_VPWR_c_412_n 0.00413917f $X=5.115 $Y=1.885 $X2=0 $Y2=0
cc_289 N_A2_c_358_n N_VPWR_c_399_n 0.0081781f $X=4.665 $Y=1.885 $X2=0 $Y2=0
cc_290 N_A2_c_360_n N_VPWR_c_399_n 0.00821601f $X=5.115 $Y=1.885 $X2=0 $Y2=0
cc_291 N_A2_c_358_n N_A_503_392#_c_564_n 0.00605728f $X=4.665 $Y=1.885 $X2=0
+ $Y2=0
cc_292 N_A2_c_358_n N_A_503_392#_c_565_n 0.0136736f $X=4.665 $Y=1.885 $X2=0
+ $Y2=0
cc_293 N_A2_c_360_n N_A_503_392#_c_565_n 0.01884f $X=5.115 $Y=1.885 $X2=0 $Y2=0
cc_294 N_A2_c_355_n N_A_503_392#_c_565_n 0.0299228f $X=4.74 $Y=1.425 $X2=0 $Y2=0
cc_295 N_A2_c_356_n N_A_503_392#_c_565_n 0.00121557f $X=5.13 $Y=1.425 $X2=0
+ $Y2=0
cc_296 N_A2_c_360_n N_A_503_392#_c_566_n 4.02768e-19 $X=5.115 $Y=1.885 $X2=0
+ $Y2=0
cc_297 N_A2_c_360_n N_A_503_392#_c_567_n 0.00634858f $X=5.115 $Y=1.885 $X2=0
+ $Y2=0
cc_298 N_A2_c_355_n N_A_503_392#_c_568_n 0.0072558f $X=4.74 $Y=1.425 $X2=0 $Y2=0
cc_299 N_A2_M1001_g N_VGND_c_624_n 0.00801653f $X=4.7 $Y=0.69 $X2=0 $Y2=0
cc_300 N_A2_M1014_g N_VGND_c_624_n 0.0116536f $X=5.13 $Y=0.69 $X2=0 $Y2=0
cc_301 N_A2_M1001_g N_VGND_c_631_n 0.00383152f $X=4.7 $Y=0.69 $X2=0 $Y2=0
cc_302 N_A2_M1014_g N_VGND_c_633_n 0.00383152f $X=5.13 $Y=0.69 $X2=0 $Y2=0
cc_303 N_A2_M1001_g N_VGND_c_634_n 0.00757637f $X=4.7 $Y=0.69 $X2=0 $Y2=0
cc_304 N_A2_M1014_g N_VGND_c_634_n 0.00761578f $X=5.13 $Y=0.69 $X2=0 $Y2=0
cc_305 N_A2_M1001_g N_A_700_74#_c_707_n 9.48753e-19 $X=4.7 $Y=0.69 $X2=0 $Y2=0
cc_306 N_A2_M1001_g N_A_700_74#_c_709_n 0.0129822f $X=4.7 $Y=0.69 $X2=0 $Y2=0
cc_307 N_A2_M1014_g N_A_700_74#_c_709_n 0.0183911f $X=5.13 $Y=0.69 $X2=0 $Y2=0
cc_308 N_A2_c_355_n N_A_700_74#_c_709_n 0.0255536f $X=4.74 $Y=1.425 $X2=0 $Y2=0
cc_309 N_A2_c_356_n N_A_700_74#_c_709_n 0.00303269f $X=5.13 $Y=1.425 $X2=0 $Y2=0
cc_310 N_A2_c_355_n N_A_700_74#_c_710_n 0.0113888f $X=4.74 $Y=1.425 $X2=0 $Y2=0
cc_311 N_A2_M1014_g N_A_700_74#_c_711_n 4.43891e-19 $X=5.13 $Y=0.69 $X2=0 $Y2=0
cc_312 N_VPWR_M1002_s N_X_c_491_n 6.05921e-19 $X=0.195 $Y=1.84 $X2=0 $Y2=0
cc_313 N_VPWR_c_401_n N_X_c_491_n 0.00570665f $X=0.32 $Y=2.225 $X2=0 $Y2=0
cc_314 N_VPWR_M1002_s N_X_c_492_n 0.00245417f $X=0.195 $Y=1.84 $X2=0 $Y2=0
cc_315 N_VPWR_c_401_n N_X_c_492_n 0.0180801f $X=0.32 $Y=2.225 $X2=0 $Y2=0
cc_316 N_VPWR_c_401_n N_X_c_493_n 0.0547423f $X=0.32 $Y=2.225 $X2=0 $Y2=0
cc_317 N_VPWR_c_402_n N_X_c_493_n 0.0535896f $X=1.22 $Y=2.305 $X2=0 $Y2=0
cc_318 N_VPWR_c_410_n N_X_c_493_n 0.00749631f $X=1.055 $Y=3.33 $X2=0 $Y2=0
cc_319 N_VPWR_c_399_n N_X_c_493_n 0.0062048f $X=5.52 $Y=3.33 $X2=0 $Y2=0
cc_320 N_VPWR_M1004_s N_X_c_494_n 0.00222494f $X=1.07 $Y=1.84 $X2=0 $Y2=0
cc_321 N_VPWR_c_402_n N_X_c_494_n 0.0154248f $X=1.22 $Y=2.305 $X2=0 $Y2=0
cc_322 N_VPWR_c_403_n N_X_c_494_n 0.00142382f $X=2.12 $Y=2.115 $X2=0 $Y2=0
cc_323 N_VPWR_c_402_n N_X_c_495_n 0.0563525f $X=1.22 $Y=2.305 $X2=0 $Y2=0
cc_324 N_VPWR_c_403_n N_X_c_495_n 0.0677182f $X=2.12 $Y=2.115 $X2=0 $Y2=0
cc_325 N_VPWR_c_411_n N_X_c_495_n 0.014552f $X=2.035 $Y=3.33 $X2=0 $Y2=0
cc_326 N_VPWR_c_399_n N_X_c_495_n 0.0119791f $X=5.52 $Y=3.33 $X2=0 $Y2=0
cc_327 N_VPWR_c_403_n N_A_503_392#_c_559_n 0.0704733f $X=2.12 $Y=2.115 $X2=0
+ $Y2=0
cc_328 N_VPWR_c_404_n N_A_503_392#_c_560_n 0.0123543f $X=3.99 $Y=2.455 $X2=0
+ $Y2=0
cc_329 N_VPWR_c_406_n N_A_503_392#_c_560_n 0.0582543f $X=3.825 $Y=3.33 $X2=0
+ $Y2=0
cc_330 N_VPWR_c_399_n N_A_503_392#_c_560_n 0.0326789f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_331 N_VPWR_c_403_n N_A_503_392#_c_561_n 0.0136296f $X=2.12 $Y=2.115 $X2=0
+ $Y2=0
cc_332 N_VPWR_c_406_n N_A_503_392#_c_561_n 0.0179217f $X=3.825 $Y=3.33 $X2=0
+ $Y2=0
cc_333 N_VPWR_c_399_n N_A_503_392#_c_561_n 0.00971942f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_334 N_VPWR_c_404_n N_A_503_392#_c_574_n 0.039183f $X=3.99 $Y=2.455 $X2=0
+ $Y2=0
cc_335 N_VPWR_M1003_d N_A_503_392#_c_563_n 0.00222494f $X=3.84 $Y=1.96 $X2=0
+ $Y2=0
cc_336 N_VPWR_c_404_n N_A_503_392#_c_563_n 0.0154248f $X=3.99 $Y=2.455 $X2=0
+ $Y2=0
cc_337 N_VPWR_c_404_n N_A_503_392#_c_564_n 0.0453479f $X=3.99 $Y=2.455 $X2=0
+ $Y2=0
cc_338 N_VPWR_c_405_n N_A_503_392#_c_564_n 0.0462948f $X=4.89 $Y=2.455 $X2=0
+ $Y2=0
cc_339 N_VPWR_c_408_n N_A_503_392#_c_564_n 0.0110241f $X=4.725 $Y=3.33 $X2=0
+ $Y2=0
cc_340 N_VPWR_c_399_n N_A_503_392#_c_564_n 0.00909194f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_341 N_VPWR_M1007_d N_A_503_392#_c_565_n 0.00197722f $X=4.74 $Y=1.96 $X2=0
+ $Y2=0
cc_342 N_VPWR_c_405_n N_A_503_392#_c_565_n 0.0171814f $X=4.89 $Y=2.455 $X2=0
+ $Y2=0
cc_343 N_VPWR_c_405_n N_A_503_392#_c_567_n 0.0462948f $X=4.89 $Y=2.455 $X2=0
+ $Y2=0
cc_344 N_VPWR_c_412_n N_A_503_392#_c_567_n 0.011066f $X=5.52 $Y=3.33 $X2=0 $Y2=0
cc_345 N_VPWR_c_399_n N_A_503_392#_c_567_n 0.00915947f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_346 N_X_c_484_n N_VGND_M1006_s 4.46468e-19 $X=0.66 $Y=1.045 $X2=-0.19
+ $Y2=-0.245
cc_347 N_X_c_485_n N_VGND_M1006_s 0.00291902f $X=0.355 $Y=1.045 $X2=-0.19
+ $Y2=-0.245
cc_348 N_X_c_487_n N_VGND_M1010_s 0.00176461f $X=1.44 $Y=1.045 $X2=0 $Y2=0
cc_349 N_X_c_484_n N_VGND_c_620_n 0.00524802f $X=0.66 $Y=1.045 $X2=0 $Y2=0
cc_350 N_X_c_485_n N_VGND_c_620_n 0.0184602f $X=0.355 $Y=1.045 $X2=0 $Y2=0
cc_351 N_X_c_486_n N_VGND_c_620_n 0.0164567f $X=0.745 $Y=0.515 $X2=0 $Y2=0
cc_352 N_X_c_486_n N_VGND_c_621_n 0.0157999f $X=0.745 $Y=0.515 $X2=0 $Y2=0
cc_353 N_X_c_487_n N_VGND_c_621_n 0.0152916f $X=1.44 $Y=1.045 $X2=0 $Y2=0
cc_354 N_X_c_488_n N_VGND_c_621_n 0.0158413f $X=1.605 $Y=0.515 $X2=0 $Y2=0
cc_355 N_X_c_488_n N_VGND_c_622_n 0.0204783f $X=1.605 $Y=0.515 $X2=0 $Y2=0
cc_356 N_X_c_486_n N_VGND_c_625_n 0.00749631f $X=0.745 $Y=0.515 $X2=0 $Y2=0
cc_357 N_X_c_488_n N_VGND_c_627_n 0.0109942f $X=1.605 $Y=0.515 $X2=0 $Y2=0
cc_358 N_X_c_486_n N_VGND_c_634_n 0.0062048f $X=0.745 $Y=0.515 $X2=0 $Y2=0
cc_359 N_X_c_488_n N_VGND_c_634_n 0.00904371f $X=1.605 $Y=0.515 $X2=0 $Y2=0
cc_360 N_VGND_c_623_n N_A_700_74#_c_706_n 0.0257494f $X=2.955 $Y=0.76 $X2=0
+ $Y2=0
cc_361 N_VGND_c_624_n N_A_700_74#_c_707_n 0.0112234f $X=4.915 $Y=0.585 $X2=0
+ $Y2=0
cc_362 N_VGND_c_631_n N_A_700_74#_c_707_n 0.050626f $X=4.75 $Y=0 $X2=0 $Y2=0
cc_363 N_VGND_c_634_n N_A_700_74#_c_707_n 0.028285f $X=5.52 $Y=0 $X2=0 $Y2=0
cc_364 N_VGND_c_623_n N_A_700_74#_c_708_n 0.00929004f $X=2.955 $Y=0.76 $X2=0
+ $Y2=0
cc_365 N_VGND_c_631_n N_A_700_74#_c_708_n 0.0235818f $X=4.75 $Y=0 $X2=0 $Y2=0
cc_366 N_VGND_c_634_n N_A_700_74#_c_708_n 0.0127177f $X=5.52 $Y=0 $X2=0 $Y2=0
cc_367 N_VGND_M1001_s N_A_700_74#_c_709_n 0.00176461f $X=4.775 $Y=0.37 $X2=0
+ $Y2=0
cc_368 N_VGND_c_624_n N_A_700_74#_c_709_n 0.0170777f $X=4.915 $Y=0.585 $X2=0
+ $Y2=0
cc_369 N_VGND_c_624_n N_A_700_74#_c_711_n 0.0150645f $X=4.915 $Y=0.585 $X2=0
+ $Y2=0
cc_370 N_VGND_c_633_n N_A_700_74#_c_711_n 0.011066f $X=5.52 $Y=0 $X2=0 $Y2=0
cc_371 N_VGND_c_634_n N_A_700_74#_c_711_n 0.00915947f $X=5.52 $Y=0 $X2=0 $Y2=0
