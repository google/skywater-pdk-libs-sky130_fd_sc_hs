* File: sky130_fd_sc_hs__o22ai_2.pxi.spice
* Created: Tue Sep  1 20:16:28 2020
* 
x_PM_SKY130_FD_SC_HS__O22AI_2%B1 N_B1_M1009_g N_B1_c_83_n N_B1_M1002_g
+ N_B1_c_84_n N_B1_M1006_g N_B1_M1012_g B1 B1 B1 N_B1_c_82_n
+ PM_SKY130_FD_SC_HS__O22AI_2%B1
x_PM_SKY130_FD_SC_HS__O22AI_2%B2 N_B2_c_129_n N_B2_M1005_g N_B2_M1003_g
+ N_B2_c_130_n N_B2_M1008_g N_B2_M1007_g B2 N_B2_c_127_n N_B2_c_128_n
+ PM_SKY130_FD_SC_HS__O22AI_2%B2
x_PM_SKY130_FD_SC_HS__O22AI_2%A2 N_A2_M1010_g N_A2_c_187_n N_A2_M1011_g
+ N_A2_c_188_n N_A2_M1013_g N_A2_M1014_g A2 N_A2_c_185_n N_A2_c_186_n
+ PM_SKY130_FD_SC_HS__O22AI_2%A2
x_PM_SKY130_FD_SC_HS__O22AI_2%A1 N_A1_M1001_g N_A1_c_247_n N_A1_M1000_g
+ N_A1_c_248_n N_A1_M1015_g N_A1_M1004_g A1 A1 N_A1_c_246_n
+ PM_SKY130_FD_SC_HS__O22AI_2%A1
x_PM_SKY130_FD_SC_HS__O22AI_2%A_28_368# N_A_28_368#_M1002_d N_A_28_368#_M1006_d
+ N_A_28_368#_M1008_s N_A_28_368#_c_290_n N_A_28_368#_c_291_n
+ N_A_28_368#_c_297_n N_A_28_368#_c_301_n N_A_28_368#_c_303_n
+ N_A_28_368#_c_292_n N_A_28_368#_c_293_n N_A_28_368#_c_294_n
+ PM_SKY130_FD_SC_HS__O22AI_2%A_28_368#
x_PM_SKY130_FD_SC_HS__O22AI_2%VPWR N_VPWR_M1002_s N_VPWR_M1000_s N_VPWR_c_337_n
+ N_VPWR_c_338_n N_VPWR_c_339_n N_VPWR_c_340_n VPWR N_VPWR_c_341_n
+ N_VPWR_c_342_n N_VPWR_c_336_n N_VPWR_c_344_n PM_SKY130_FD_SC_HS__O22AI_2%VPWR
x_PM_SKY130_FD_SC_HS__O22AI_2%Y N_Y_M1009_s N_Y_M1003_s N_Y_M1005_d N_Y_M1011_d
+ N_Y_c_449_p N_Y_c_386_n N_Y_c_387_n N_Y_c_401_n N_Y_c_402_n N_Y_c_390_n
+ N_Y_c_420_n N_Y_c_404_n N_Y_c_388_n N_Y_c_391_n Y
+ PM_SKY130_FD_SC_HS__O22AI_2%Y
x_PM_SKY130_FD_SC_HS__O22AI_2%A_510_368# N_A_510_368#_M1011_s
+ N_A_510_368#_M1013_s N_A_510_368#_M1015_d N_A_510_368#_c_458_n
+ N_A_510_368#_c_459_n N_A_510_368#_c_460_n N_A_510_368#_c_470_n
+ N_A_510_368#_c_489_n N_A_510_368#_c_471_n N_A_510_368#_c_461_n
+ N_A_510_368#_c_462_n PM_SKY130_FD_SC_HS__O22AI_2%A_510_368#
x_PM_SKY130_FD_SC_HS__O22AI_2%A_27_74# N_A_27_74#_M1009_d N_A_27_74#_M1012_d
+ N_A_27_74#_M1007_d N_A_27_74#_M1014_d N_A_27_74#_M1004_d N_A_27_74#_c_503_n
+ N_A_27_74#_c_504_n N_A_27_74#_c_505_n N_A_27_74#_c_520_n N_A_27_74#_c_506_n
+ N_A_27_74#_c_507_n N_A_27_74#_c_508_n N_A_27_74#_c_509_n N_A_27_74#_c_510_n
+ N_A_27_74#_c_511_n N_A_27_74#_c_512_n N_A_27_74#_c_513_n
+ PM_SKY130_FD_SC_HS__O22AI_2%A_27_74#
x_PM_SKY130_FD_SC_HS__O22AI_2%VGND N_VGND_M1010_s N_VGND_M1001_s N_VGND_c_581_n
+ N_VGND_c_582_n VGND N_VGND_c_583_n N_VGND_c_584_n N_VGND_c_585_n
+ N_VGND_c_586_n N_VGND_c_587_n N_VGND_c_588_n PM_SKY130_FD_SC_HS__O22AI_2%VGND
cc_1 VNB N_B1_M1009_g 0.033015f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_2 VNB N_B1_M1012_g 0.0244807f $X=-0.19 $Y=-0.245 $X2=1.025 $Y2=0.74
cc_3 VNB B1 0.0210388f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.58
cc_4 VNB N_B1_c_82_n 0.0400048f $X=-0.19 $Y=-0.245 $X2=1.01 $Y2=1.557
cc_5 VNB N_B2_M1003_g 0.0240538f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=2.4
cc_6 VNB N_B2_M1007_g 0.0279479f $X=-0.19 $Y=-0.245 $X2=1.025 $Y2=0.74
cc_7 VNB N_B2_c_127_n 0.00143484f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.557
cc_8 VNB N_B2_c_128_n 0.0439325f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=1.557
cc_9 VNB N_A2_M1010_g 0.0239562f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_10 VNB N_A2_M1014_g 0.0219989f $X=-0.19 $Y=-0.245 $X2=1.025 $Y2=0.74
cc_11 VNB A2 0.00755947f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.58
cc_12 VNB N_A2_c_185_n 0.00345565f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=1.557
cc_13 VNB N_A2_c_186_n 0.0626259f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=1.515
cc_14 VNB N_A1_M1001_g 0.0244981f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_15 VNB N_A1_M1004_g 0.0328675f $X=-0.19 $Y=-0.245 $X2=1.025 $Y2=0.74
cc_16 VNB A1 0.0134698f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_17 VNB N_A1_c_246_n 0.0517161f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=1.557
cc_18 VNB N_VPWR_c_336_n 0.203486f $X=-0.19 $Y=-0.245 $X2=1.2 $Y2=1.565
cc_19 VNB N_Y_c_386_n 0.00474786f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.58
cc_20 VNB N_Y_c_387_n 0.00340221f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_Y_c_388_n 0.00615473f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB Y 0.00712626f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_27_74#_c_503_n 0.0302158f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_27_74#_c_504_n 0.00288965f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_27_74#_c_505_n 0.00971634f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.557
cc_26 VNB N_A_27_74#_c_506_n 0.00280532f $X=-0.19 $Y=-0.245 $X2=1.01 $Y2=1.557
cc_27 VNB N_A_27_74#_c_507_n 0.00329829f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.565
cc_28 VNB N_A_27_74#_c_508_n 0.00207407f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_27_74#_c_509_n 0.0132237f $X=-0.19 $Y=-0.245 $X2=1.2 $Y2=1.565
cc_30 VNB N_A_27_74#_c_510_n 0.0266107f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_27_74#_c_511_n 0.00220733f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_27_74#_c_512_n 0.012391f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_27_74#_c_513_n 0.00327131f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_581_n 0.00572435f $X=-0.19 $Y=-0.245 $X2=1.01 $Y2=2.4
cc_35 VNB N_VGND_c_582_n 0.00566037f $X=-0.19 $Y=-0.245 $X2=1.025 $Y2=0.74
cc_36 VNB N_VGND_c_583_n 0.0703081f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.58
cc_37 VNB N_VGND_c_584_n 0.0183651f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=1.515
cc_38 VNB N_VGND_c_585_n 0.0173909f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_586_n 0.276858f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=1.565
cc_40 VNB N_VGND_c_587_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_588_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VPB N_B1_c_83_n 0.0205227f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=1.765
cc_43 VPB N_B1_c_84_n 0.0156228f $X=-0.19 $Y=1.66 $X2=1.01 $Y2=1.765
cc_44 VPB B1 0.0144621f $X=-0.19 $Y=1.66 $X2=1.115 $Y2=1.58
cc_45 VPB N_B1_c_82_n 0.0224364f $X=-0.19 $Y=1.66 $X2=1.01 $Y2=1.557
cc_46 VPB N_B2_c_129_n 0.0148479f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.35
cc_47 VPB N_B2_c_130_n 0.0170112f $X=-0.19 $Y=1.66 $X2=1.01 $Y2=1.765
cc_48 VPB N_B2_c_127_n 0.00425857f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.557
cc_49 VPB N_B2_c_128_n 0.0206707f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=1.557
cc_50 VPB N_A2_c_187_n 0.0173891f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=1.765
cc_51 VPB N_A2_c_188_n 0.0147113f $X=-0.19 $Y=1.66 $X2=1.01 $Y2=1.765
cc_52 VPB A2 0.00500584f $X=-0.19 $Y=1.66 $X2=1.115 $Y2=1.58
cc_53 VPB N_A2_c_186_n 0.0145966f $X=-0.19 $Y=1.66 $X2=0.925 $Y2=1.515
cc_54 VPB N_A1_c_247_n 0.0153896f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=1.765
cc_55 VPB N_A1_c_248_n 0.0208611f $X=-0.19 $Y=1.66 $X2=1.01 $Y2=1.765
cc_56 VPB A1 0.011105f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_57 VPB N_A1_c_246_n 0.0278557f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=1.557
cc_58 VPB N_A_28_368#_c_290_n 0.00739392f $X=-0.19 $Y=1.66 $X2=1.01 $Y2=2.4
cc_59 VPB N_A_28_368#_c_291_n 0.0339313f $X=-0.19 $Y=1.66 $X2=1.025 $Y2=0.74
cc_60 VPB N_A_28_368#_c_292_n 0.00644841f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_61 VPB N_A_28_368#_c_293_n 0.0021839f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.557
cc_62 VPB N_A_28_368#_c_294_n 0.00568479f $X=-0.19 $Y=1.66 $X2=0.925 $Y2=1.515
cc_63 VPB N_VPWR_c_337_n 0.00610411f $X=-0.19 $Y=1.66 $X2=1.01 $Y2=2.4
cc_64 VPB N_VPWR_c_338_n 0.00571271f $X=-0.19 $Y=1.66 $X2=1.025 $Y2=0.74
cc_65 VPB N_VPWR_c_339_n 0.0715292f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_66 VPB N_VPWR_c_340_n 0.00460249f $X=-0.19 $Y=1.66 $X2=1.115 $Y2=1.58
cc_67 VPB N_VPWR_c_341_n 0.0181665f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_68 VPB N_VPWR_c_342_n 0.0209017f $X=-0.19 $Y=1.66 $X2=0.925 $Y2=1.565
cc_69 VPB N_VPWR_c_336_n 0.0831118f $X=-0.19 $Y=1.66 $X2=1.2 $Y2=1.565
cc_70 VPB N_VPWR_c_344_n 0.00613757f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_71 VPB N_Y_c_390_n 0.0228497f $X=-0.19 $Y=1.66 $X2=1.025 $Y2=1.557
cc_72 VPB N_Y_c_391_n 6.30886e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_73 VPB Y 0.00379399f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_74 VPB N_A_510_368#_c_458_n 0.00791255f $X=-0.19 $Y=1.66 $X2=1.025 $Y2=0.74
cc_75 VPB N_A_510_368#_c_459_n 0.00478015f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_76 VPB N_A_510_368#_c_460_n 0.00431238f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_77 VPB N_A_510_368#_c_461_n 0.00723723f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=1.557
cc_78 VPB N_A_510_368#_c_462_n 0.035396f $X=-0.19 $Y=1.66 $X2=0.925 $Y2=1.515
cc_79 N_B1_c_84_n N_B2_c_129_n 0.0126076f $X=1.01 $Y=1.765 $X2=-0.19 $Y2=-0.245
cc_80 N_B1_M1012_g N_B2_M1003_g 0.0279646f $X=1.025 $Y=0.74 $X2=0 $Y2=0
cc_81 B1 N_B2_c_127_n 0.0360516f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_82 N_B1_c_82_n N_B2_c_127_n 3.09177e-19 $X=1.01 $Y=1.557 $X2=0 $Y2=0
cc_83 B1 N_B2_c_128_n 0.00384452f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_84 N_B1_c_82_n N_B2_c_128_n 0.0191318f $X=1.01 $Y=1.557 $X2=0 $Y2=0
cc_85 B1 N_A_28_368#_c_290_n 0.021684f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_86 N_B1_c_83_n N_A_28_368#_c_291_n 0.00634858f $X=0.51 $Y=1.765 $X2=0 $Y2=0
cc_87 N_B1_c_83_n N_A_28_368#_c_297_n 0.0129585f $X=0.51 $Y=1.765 $X2=0 $Y2=0
cc_88 N_B1_c_84_n N_A_28_368#_c_297_n 0.0122806f $X=1.01 $Y=1.765 $X2=0 $Y2=0
cc_89 B1 N_A_28_368#_c_297_n 0.0475354f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_90 N_B1_c_82_n N_A_28_368#_c_297_n 0.00158477f $X=1.01 $Y=1.557 $X2=0 $Y2=0
cc_91 N_B1_c_84_n N_A_28_368#_c_301_n 4.27055e-19 $X=1.01 $Y=1.765 $X2=0 $Y2=0
cc_92 B1 N_A_28_368#_c_301_n 0.0189518f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_93 N_B1_c_83_n N_A_28_368#_c_303_n 7.18055e-19 $X=0.51 $Y=1.765 $X2=0 $Y2=0
cc_94 N_B1_c_84_n N_A_28_368#_c_303_n 0.00898942f $X=1.01 $Y=1.765 $X2=0 $Y2=0
cc_95 N_B1_c_84_n N_A_28_368#_c_293_n 0.00312124f $X=1.01 $Y=1.765 $X2=0 $Y2=0
cc_96 N_B1_c_83_n N_VPWR_c_337_n 0.0140375f $X=0.51 $Y=1.765 $X2=0 $Y2=0
cc_97 N_B1_c_84_n N_VPWR_c_337_n 0.00496464f $X=1.01 $Y=1.765 $X2=0 $Y2=0
cc_98 N_B1_c_84_n N_VPWR_c_339_n 0.0044313f $X=1.01 $Y=1.765 $X2=0 $Y2=0
cc_99 N_B1_c_83_n N_VPWR_c_341_n 0.00413917f $X=0.51 $Y=1.765 $X2=0 $Y2=0
cc_100 N_B1_c_83_n N_VPWR_c_336_n 0.00821237f $X=0.51 $Y=1.765 $X2=0 $Y2=0
cc_101 N_B1_c_84_n N_VPWR_c_336_n 0.00853234f $X=1.01 $Y=1.765 $X2=0 $Y2=0
cc_102 N_B1_M1012_g N_Y_c_386_n 0.012846f $X=1.025 $Y=0.74 $X2=0 $Y2=0
cc_103 B1 N_Y_c_386_n 0.0287022f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_104 N_B1_M1009_g N_Y_c_387_n 0.00241337f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_105 B1 N_Y_c_387_n 0.0280045f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_106 N_B1_c_82_n N_Y_c_387_n 0.00463094f $X=1.01 $Y=1.557 $X2=0 $Y2=0
cc_107 N_B1_M1009_g N_A_27_74#_c_503_n 0.0108851f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_108 N_B1_M1012_g N_A_27_74#_c_503_n 6.35781e-19 $X=1.025 $Y=0.74 $X2=0 $Y2=0
cc_109 B1 N_A_27_74#_c_503_n 0.023775f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_110 N_B1_M1009_g N_A_27_74#_c_504_n 0.0106115f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_111 N_B1_M1012_g N_A_27_74#_c_504_n 0.0118932f $X=1.025 $Y=0.74 $X2=0 $Y2=0
cc_112 N_B1_M1009_g N_A_27_74#_c_505_n 0.00282152f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_113 N_B1_M1009_g N_VGND_c_583_n 0.00278247f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_114 N_B1_M1012_g N_VGND_c_583_n 0.00278271f $X=1.025 $Y=0.74 $X2=0 $Y2=0
cc_115 N_B1_M1009_g N_VGND_c_586_n 0.00357999f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_116 N_B1_M1012_g N_VGND_c_586_n 0.00354801f $X=1.025 $Y=0.74 $X2=0 $Y2=0
cc_117 N_B2_M1007_g N_A2_c_186_n 0.00279892f $X=1.995 $Y=0.74 $X2=0 $Y2=0
cc_118 N_B2_c_128_n N_A2_c_186_n 0.00143843f $X=1.91 $Y=1.557 $X2=0 $Y2=0
cc_119 N_B2_c_129_n N_A_28_368#_c_301_n 0.00228787f $X=1.46 $Y=1.765 $X2=0 $Y2=0
cc_120 N_B2_c_129_n N_A_28_368#_c_303_n 0.00876394f $X=1.46 $Y=1.765 $X2=0 $Y2=0
cc_121 N_B2_c_130_n N_A_28_368#_c_303_n 5.9624e-19 $X=1.91 $Y=1.765 $X2=0 $Y2=0
cc_122 N_B2_c_129_n N_A_28_368#_c_292_n 0.0108414f $X=1.46 $Y=1.765 $X2=0 $Y2=0
cc_123 N_B2_c_130_n N_A_28_368#_c_292_n 0.0134708f $X=1.91 $Y=1.765 $X2=0 $Y2=0
cc_124 N_B2_c_129_n N_A_28_368#_c_293_n 0.00171731f $X=1.46 $Y=1.765 $X2=0 $Y2=0
cc_125 N_B2_c_129_n N_A_28_368#_c_294_n 5.52094e-19 $X=1.46 $Y=1.765 $X2=0 $Y2=0
cc_126 N_B2_c_130_n N_A_28_368#_c_294_n 0.00837677f $X=1.91 $Y=1.765 $X2=0 $Y2=0
cc_127 N_B2_c_129_n N_VPWR_c_339_n 0.00278257f $X=1.46 $Y=1.765 $X2=0 $Y2=0
cc_128 N_B2_c_130_n N_VPWR_c_339_n 0.00278257f $X=1.91 $Y=1.765 $X2=0 $Y2=0
cc_129 N_B2_c_129_n N_VPWR_c_336_n 0.00353905f $X=1.46 $Y=1.765 $X2=0 $Y2=0
cc_130 N_B2_c_130_n N_VPWR_c_336_n 0.00358623f $X=1.91 $Y=1.765 $X2=0 $Y2=0
cc_131 N_B2_M1003_g N_Y_c_386_n 0.014657f $X=1.495 $Y=0.74 $X2=0 $Y2=0
cc_132 N_B2_c_127_n N_Y_c_386_n 0.0249311f $X=1.65 $Y=1.515 $X2=0 $Y2=0
cc_133 N_B2_c_128_n N_Y_c_386_n 0.0020325f $X=1.91 $Y=1.557 $X2=0 $Y2=0
cc_134 N_B2_M1007_g N_Y_c_401_n 0.0068998f $X=1.995 $Y=0.74 $X2=0 $Y2=0
cc_135 N_B2_c_130_n N_Y_c_402_n 0.017676f $X=1.91 $Y=1.765 $X2=0 $Y2=0
cc_136 N_B2_c_128_n N_Y_c_402_n 8.48385e-19 $X=1.91 $Y=1.557 $X2=0 $Y2=0
cc_137 N_B2_c_127_n N_Y_c_404_n 0.0184426f $X=1.65 $Y=1.515 $X2=0 $Y2=0
cc_138 N_B2_c_128_n N_Y_c_404_n 0.00129847f $X=1.91 $Y=1.557 $X2=0 $Y2=0
cc_139 N_B2_M1007_g N_Y_c_388_n 0.0167839f $X=1.995 $Y=0.74 $X2=0 $Y2=0
cc_140 N_B2_c_128_n N_Y_c_388_n 0.00169754f $X=1.91 $Y=1.557 $X2=0 $Y2=0
cc_141 N_B2_c_129_n N_Y_c_391_n 2.7303e-19 $X=1.46 $Y=1.765 $X2=0 $Y2=0
cc_142 N_B2_c_130_n N_Y_c_391_n 0.00144336f $X=1.91 $Y=1.765 $X2=0 $Y2=0
cc_143 N_B2_M1003_g Y 8.02322e-19 $X=1.495 $Y=0.74 $X2=0 $Y2=0
cc_144 N_B2_c_130_n Y 0.00713359f $X=1.91 $Y=1.765 $X2=0 $Y2=0
cc_145 N_B2_M1007_g Y 0.00612352f $X=1.995 $Y=0.74 $X2=0 $Y2=0
cc_146 N_B2_c_127_n Y 0.0261971f $X=1.65 $Y=1.515 $X2=0 $Y2=0
cc_147 N_B2_c_128_n Y 0.0111373f $X=1.91 $Y=1.557 $X2=0 $Y2=0
cc_148 N_B2_c_130_n N_A_510_368#_c_458_n 0.00366099f $X=1.91 $Y=1.765 $X2=0
+ $Y2=0
cc_149 N_B2_c_130_n N_A_510_368#_c_460_n 5.92854e-19 $X=1.91 $Y=1.765 $X2=0
+ $Y2=0
cc_150 N_B2_M1003_g N_A_27_74#_c_520_n 0.00682727f $X=1.495 $Y=0.74 $X2=0 $Y2=0
cc_151 N_B2_M1007_g N_A_27_74#_c_520_n 4.62551e-19 $X=1.995 $Y=0.74 $X2=0 $Y2=0
cc_152 N_B2_M1003_g N_A_27_74#_c_506_n 0.00831967f $X=1.495 $Y=0.74 $X2=0 $Y2=0
cc_153 N_B2_M1007_g N_A_27_74#_c_506_n 0.0132502f $X=1.995 $Y=0.74 $X2=0 $Y2=0
cc_154 N_B2_M1003_g N_A_27_74#_c_511_n 0.00272972f $X=1.495 $Y=0.74 $X2=0 $Y2=0
cc_155 N_B2_M1007_g N_A_27_74#_c_512_n 0.0033343f $X=1.995 $Y=0.74 $X2=0 $Y2=0
cc_156 N_B2_M1003_g N_VGND_c_583_n 0.00278247f $X=1.495 $Y=0.74 $X2=0 $Y2=0
cc_157 N_B2_M1007_g N_VGND_c_583_n 0.00278271f $X=1.995 $Y=0.74 $X2=0 $Y2=0
cc_158 N_B2_M1003_g N_VGND_c_586_n 0.00354543f $X=1.495 $Y=0.74 $X2=0 $Y2=0
cc_159 N_B2_M1007_g N_VGND_c_586_n 0.00359085f $X=1.995 $Y=0.74 $X2=0 $Y2=0
cc_160 N_A2_M1014_g N_A1_M1001_g 0.0167769f $X=3.375 $Y=0.74 $X2=0 $Y2=0
cc_161 A2 N_A1_M1001_g 3.98292e-19 $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_162 N_A2_c_186_n N_A1_M1001_g 0.0215027f $X=3.37 $Y=1.532 $X2=0 $Y2=0
cc_163 N_A2_c_188_n N_A1_c_247_n 0.0113554f $X=3.37 $Y=1.765 $X2=0 $Y2=0
cc_164 A2 A1 0.0315595f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_165 N_A2_c_186_n A1 2.9359e-19 $X=3.37 $Y=1.532 $X2=0 $Y2=0
cc_166 A2 N_A1_c_246_n 0.00386828f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_167 N_A2_c_187_n N_A_28_368#_c_292_n 5.92854e-19 $X=2.92 $Y=1.765 $X2=0 $Y2=0
cc_168 N_A2_c_187_n N_A_28_368#_c_294_n 0.0013063f $X=2.92 $Y=1.765 $X2=0 $Y2=0
cc_169 N_A2_c_187_n N_VPWR_c_339_n 0.00278257f $X=2.92 $Y=1.765 $X2=0 $Y2=0
cc_170 N_A2_c_188_n N_VPWR_c_339_n 0.00278271f $X=3.37 $Y=1.765 $X2=0 $Y2=0
cc_171 N_A2_c_187_n N_VPWR_c_336_n 0.00358623f $X=2.92 $Y=1.765 $X2=0 $Y2=0
cc_172 N_A2_c_188_n N_VPWR_c_336_n 0.00353907f $X=3.37 $Y=1.765 $X2=0 $Y2=0
cc_173 N_A2_c_187_n N_Y_c_390_n 0.014933f $X=2.92 $Y=1.765 $X2=0 $Y2=0
cc_174 N_A2_c_188_n N_Y_c_390_n 0.00381291f $X=3.37 $Y=1.765 $X2=0 $Y2=0
cc_175 A2 N_Y_c_390_n 0.0117965f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_176 N_A2_c_185_n N_Y_c_390_n 0.0383263f $X=3.17 $Y=1.465 $X2=0 $Y2=0
cc_177 N_A2_c_186_n N_Y_c_390_n 0.00988904f $X=3.37 $Y=1.532 $X2=0 $Y2=0
cc_178 N_A2_c_187_n N_Y_c_420_n 0.0064963f $X=2.92 $Y=1.765 $X2=0 $Y2=0
cc_179 N_A2_c_188_n N_Y_c_420_n 0.00983812f $X=3.37 $Y=1.765 $X2=0 $Y2=0
cc_180 N_A2_M1010_g N_Y_c_388_n 0.00158819f $X=2.905 $Y=0.74 $X2=0 $Y2=0
cc_181 N_A2_c_187_n N_Y_c_391_n 0.00376984f $X=2.92 $Y=1.765 $X2=0 $Y2=0
cc_182 N_A2_M1010_g Y 0.00283903f $X=2.905 $Y=0.74 $X2=0 $Y2=0
cc_183 N_A2_c_187_n Y 8.18966e-19 $X=2.92 $Y=1.765 $X2=0 $Y2=0
cc_184 N_A2_c_185_n Y 0.0143507f $X=3.17 $Y=1.465 $X2=0 $Y2=0
cc_185 N_A2_c_186_n Y 0.00464968f $X=3.37 $Y=1.532 $X2=0 $Y2=0
cc_186 N_A2_c_187_n N_A_510_368#_c_458_n 0.0118413f $X=2.92 $Y=1.765 $X2=0 $Y2=0
cc_187 N_A2_c_188_n N_A_510_368#_c_458_n 7.1863e-19 $X=3.37 $Y=1.765 $X2=0 $Y2=0
cc_188 N_A2_c_187_n N_A_510_368#_c_459_n 0.0107904f $X=2.92 $Y=1.765 $X2=0 $Y2=0
cc_189 N_A2_c_188_n N_A_510_368#_c_459_n 0.012504f $X=3.37 $Y=1.765 $X2=0 $Y2=0
cc_190 N_A2_c_187_n N_A_510_368#_c_460_n 0.00262934f $X=2.92 $Y=1.765 $X2=0
+ $Y2=0
cc_191 A2 N_A_510_368#_c_470_n 0.0149894f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_192 A2 N_A_510_368#_c_471_n 0.00175724f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_193 N_A2_M1010_g N_A_27_74#_c_507_n 0.01289f $X=2.905 $Y=0.74 $X2=0 $Y2=0
cc_194 N_A2_M1014_g N_A_27_74#_c_507_n 0.0138493f $X=3.375 $Y=0.74 $X2=0 $Y2=0
cc_195 A2 N_A_27_74#_c_507_n 0.0212066f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_196 N_A2_c_185_n N_A_27_74#_c_507_n 0.0283f $X=3.17 $Y=1.465 $X2=0 $Y2=0
cc_197 N_A2_c_186_n N_A_27_74#_c_507_n 0.00378167f $X=3.37 $Y=1.532 $X2=0 $Y2=0
cc_198 N_A2_M1014_g N_A_27_74#_c_508_n 4.09578e-19 $X=3.375 $Y=0.74 $X2=0 $Y2=0
cc_199 N_A2_M1010_g N_A_27_74#_c_512_n 0.00384249f $X=2.905 $Y=0.74 $X2=0 $Y2=0
cc_200 N_A2_c_185_n N_A_27_74#_c_512_n 0.01012f $X=3.17 $Y=1.465 $X2=0 $Y2=0
cc_201 N_A2_c_186_n N_A_27_74#_c_512_n 0.00279548f $X=3.37 $Y=1.532 $X2=0 $Y2=0
cc_202 N_A2_M1014_g N_A_27_74#_c_513_n 0.00158218f $X=3.375 $Y=0.74 $X2=0 $Y2=0
cc_203 A2 N_A_27_74#_c_513_n 0.0162604f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_204 N_A2_M1010_g N_VGND_c_581_n 0.0092302f $X=2.905 $Y=0.74 $X2=0 $Y2=0
cc_205 N_A2_M1014_g N_VGND_c_581_n 0.00222839f $X=3.375 $Y=0.74 $X2=0 $Y2=0
cc_206 N_A2_M1010_g N_VGND_c_583_n 0.00383152f $X=2.905 $Y=0.74 $X2=0 $Y2=0
cc_207 N_A2_M1014_g N_VGND_c_584_n 0.00461464f $X=3.375 $Y=0.74 $X2=0 $Y2=0
cc_208 N_A2_M1010_g N_VGND_c_586_n 0.00762539f $X=2.905 $Y=0.74 $X2=0 $Y2=0
cc_209 N_A2_M1014_g N_VGND_c_586_n 0.00907921f $X=3.375 $Y=0.74 $X2=0 $Y2=0
cc_210 N_A1_c_247_n N_VPWR_c_338_n 0.00996098f $X=3.82 $Y=1.765 $X2=0 $Y2=0
cc_211 N_A1_c_248_n N_VPWR_c_338_n 0.00526215f $X=4.27 $Y=1.765 $X2=0 $Y2=0
cc_212 N_A1_c_247_n N_VPWR_c_339_n 0.00413917f $X=3.82 $Y=1.765 $X2=0 $Y2=0
cc_213 N_A1_c_248_n N_VPWR_c_342_n 0.00445602f $X=4.27 $Y=1.765 $X2=0 $Y2=0
cc_214 N_A1_c_247_n N_VPWR_c_336_n 0.0081781f $X=3.82 $Y=1.765 $X2=0 $Y2=0
cc_215 N_A1_c_248_n N_VPWR_c_336_n 0.00861164f $X=4.27 $Y=1.765 $X2=0 $Y2=0
cc_216 N_A1_c_247_n N_Y_c_390_n 6.40562e-19 $X=3.82 $Y=1.765 $X2=0 $Y2=0
cc_217 N_A1_c_247_n N_A_510_368#_c_459_n 0.00125031f $X=3.82 $Y=1.765 $X2=0
+ $Y2=0
cc_218 N_A1_c_247_n N_A_510_368#_c_471_n 0.0172359f $X=3.82 $Y=1.765 $X2=0 $Y2=0
cc_219 N_A1_c_248_n N_A_510_368#_c_471_n 0.0119563f $X=4.27 $Y=1.765 $X2=0 $Y2=0
cc_220 A1 N_A_510_368#_c_471_n 0.0289213f $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_221 N_A1_c_246_n N_A_510_368#_c_471_n 0.00131353f $X=4.305 $Y=1.557 $X2=0
+ $Y2=0
cc_222 N_A1_c_248_n N_A_510_368#_c_461_n 4.27055e-19 $X=4.27 $Y=1.765 $X2=0
+ $Y2=0
cc_223 A1 N_A_510_368#_c_461_n 0.0265009f $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_224 N_A1_c_246_n N_A_510_368#_c_461_n 0.00124936f $X=4.305 $Y=1.557 $X2=0
+ $Y2=0
cc_225 N_A1_c_247_n N_A_510_368#_c_462_n 6.69308e-19 $X=3.82 $Y=1.765 $X2=0
+ $Y2=0
cc_226 N_A1_c_248_n N_A_510_368#_c_462_n 0.0106911f $X=4.27 $Y=1.765 $X2=0 $Y2=0
cc_227 N_A1_M1001_g N_A_27_74#_c_508_n 0.00819795f $X=3.805 $Y=0.74 $X2=0 $Y2=0
cc_228 N_A1_M1004_g N_A_27_74#_c_508_n 6.73095e-19 $X=4.305 $Y=0.74 $X2=0 $Y2=0
cc_229 N_A1_M1001_g N_A_27_74#_c_509_n 0.0153304f $X=3.805 $Y=0.74 $X2=0 $Y2=0
cc_230 N_A1_M1004_g N_A_27_74#_c_509_n 0.0140467f $X=4.305 $Y=0.74 $X2=0 $Y2=0
cc_231 A1 N_A_27_74#_c_509_n 0.0606947f $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_232 N_A1_c_246_n N_A_27_74#_c_509_n 0.0084203f $X=4.305 $Y=1.557 $X2=0 $Y2=0
cc_233 N_A1_M1004_g N_A_27_74#_c_510_n 0.00159319f $X=4.305 $Y=0.74 $X2=0 $Y2=0
cc_234 N_A1_M1001_g N_A_27_74#_c_513_n 0.00337157f $X=3.805 $Y=0.74 $X2=0 $Y2=0
cc_235 N_A1_M1004_g N_A_27_74#_c_513_n 2.34371e-19 $X=4.305 $Y=0.74 $X2=0 $Y2=0
cc_236 N_A1_M1001_g N_VGND_c_582_n 0.00429078f $X=3.805 $Y=0.74 $X2=0 $Y2=0
cc_237 N_A1_M1004_g N_VGND_c_582_n 0.0137334f $X=4.305 $Y=0.74 $X2=0 $Y2=0
cc_238 N_A1_M1001_g N_VGND_c_584_n 0.00434272f $X=3.805 $Y=0.74 $X2=0 $Y2=0
cc_239 N_A1_M1004_g N_VGND_c_585_n 0.00383152f $X=4.305 $Y=0.74 $X2=0 $Y2=0
cc_240 N_A1_M1001_g N_VGND_c_586_n 0.00820816f $X=3.805 $Y=0.74 $X2=0 $Y2=0
cc_241 N_A1_M1004_g N_VGND_c_586_n 0.00761198f $X=4.305 $Y=0.74 $X2=0 $Y2=0
cc_242 N_A_28_368#_c_297_n N_VPWR_M1002_s 0.00455969f $X=1.07 $Y=2.035 $X2=-0.19
+ $Y2=1.66
cc_243 N_A_28_368#_c_291_n N_VPWR_c_337_n 0.0462948f $X=0.285 $Y=2.815 $X2=0
+ $Y2=0
cc_244 N_A_28_368#_c_297_n N_VPWR_c_337_n 0.0202249f $X=1.07 $Y=2.035 $X2=0
+ $Y2=0
cc_245 N_A_28_368#_c_293_n N_VPWR_c_337_n 0.0119239f $X=1.4 $Y=2.99 $X2=0 $Y2=0
cc_246 N_A_28_368#_c_292_n N_VPWR_c_339_n 0.0594839f $X=1.97 $Y=2.99 $X2=0 $Y2=0
cc_247 N_A_28_368#_c_293_n N_VPWR_c_339_n 0.0235512f $X=1.4 $Y=2.99 $X2=0 $Y2=0
cc_248 N_A_28_368#_c_291_n N_VPWR_c_341_n 0.011066f $X=0.285 $Y=2.815 $X2=0
+ $Y2=0
cc_249 N_A_28_368#_c_291_n N_VPWR_c_336_n 0.00915947f $X=0.285 $Y=2.815 $X2=0
+ $Y2=0
cc_250 N_A_28_368#_c_292_n N_VPWR_c_336_n 0.0329562f $X=1.97 $Y=2.99 $X2=0 $Y2=0
cc_251 N_A_28_368#_c_293_n N_VPWR_c_336_n 0.0126924f $X=1.4 $Y=2.99 $X2=0 $Y2=0
cc_252 N_A_28_368#_c_292_n N_Y_M1005_d 0.00197722f $X=1.97 $Y=2.99 $X2=0 $Y2=0
cc_253 N_A_28_368#_M1008_s N_Y_c_402_n 4.9676e-19 $X=1.985 $Y=1.84 $X2=0 $Y2=0
cc_254 N_A_28_368#_c_294_n N_Y_c_402_n 0.00126841f $X=2.135 $Y=2.375 $X2=0 $Y2=0
cc_255 N_A_28_368#_M1008_s N_Y_c_390_n 4.31813e-19 $X=1.985 $Y=1.84 $X2=0 $Y2=0
cc_256 N_A_28_368#_c_294_n N_Y_c_390_n 0.00128853f $X=2.135 $Y=2.375 $X2=0 $Y2=0
cc_257 N_A_28_368#_c_292_n N_Y_c_404_n 0.014157f $X=1.97 $Y=2.99 $X2=0 $Y2=0
cc_258 N_A_28_368#_M1008_s N_Y_c_391_n 0.00877927f $X=1.985 $Y=1.84 $X2=0 $Y2=0
cc_259 N_A_28_368#_c_294_n N_Y_c_391_n 0.0205569f $X=2.135 $Y=2.375 $X2=0 $Y2=0
cc_260 N_A_28_368#_c_294_n N_A_510_368#_c_458_n 0.0413951f $X=2.135 $Y=2.375
+ $X2=0 $Y2=0
cc_261 N_A_28_368#_c_292_n N_A_510_368#_c_460_n 0.0128665f $X=1.97 $Y=2.99 $X2=0
+ $Y2=0
cc_262 N_VPWR_c_338_n N_A_510_368#_c_459_n 0.0123543f $X=4.045 $Y=2.455 $X2=0
+ $Y2=0
cc_263 N_VPWR_c_339_n N_A_510_368#_c_459_n 0.0531736f $X=3.88 $Y=3.33 $X2=0
+ $Y2=0
cc_264 N_VPWR_c_336_n N_A_510_368#_c_459_n 0.0297434f $X=4.56 $Y=3.33 $X2=0
+ $Y2=0
cc_265 N_VPWR_c_339_n N_A_510_368#_c_460_n 0.0236039f $X=3.88 $Y=3.33 $X2=0
+ $Y2=0
cc_266 N_VPWR_c_336_n N_A_510_368#_c_460_n 0.012761f $X=4.56 $Y=3.33 $X2=0 $Y2=0
cc_267 N_VPWR_c_338_n N_A_510_368#_c_489_n 0.039183f $X=4.045 $Y=2.455 $X2=0
+ $Y2=0
cc_268 N_VPWR_M1000_s N_A_510_368#_c_471_n 0.00384138f $X=3.895 $Y=1.84 $X2=0
+ $Y2=0
cc_269 N_VPWR_c_338_n N_A_510_368#_c_471_n 0.0154248f $X=4.045 $Y=2.455 $X2=0
+ $Y2=0
cc_270 N_VPWR_c_338_n N_A_510_368#_c_462_n 0.0462948f $X=4.045 $Y=2.455 $X2=0
+ $Y2=0
cc_271 N_VPWR_c_342_n N_A_510_368#_c_462_n 0.0145938f $X=4.56 $Y=3.33 $X2=0
+ $Y2=0
cc_272 N_VPWR_c_336_n N_A_510_368#_c_462_n 0.0120466f $X=4.56 $Y=3.33 $X2=0
+ $Y2=0
cc_273 N_Y_c_390_n N_A_510_368#_M1011_s 0.00335111f $X=3.06 $Y=1.885 $X2=-0.19
+ $Y2=-0.245
cc_274 N_Y_c_390_n N_A_510_368#_c_458_n 0.0219924f $X=3.06 $Y=1.885 $X2=0 $Y2=0
cc_275 N_Y_c_420_n N_A_510_368#_c_458_n 0.0398954f $X=3.145 $Y=1.985 $X2=0 $Y2=0
cc_276 N_Y_M1011_d N_A_510_368#_c_459_n 0.00222494f $X=2.995 $Y=1.84 $X2=0 $Y2=0
cc_277 N_Y_c_420_n N_A_510_368#_c_459_n 0.0144323f $X=3.145 $Y=1.985 $X2=0 $Y2=0
cc_278 N_Y_c_390_n N_A_510_368#_c_470_n 0.00154024f $X=3.06 $Y=1.885 $X2=0 $Y2=0
cc_279 N_Y_c_420_n N_A_510_368#_c_470_n 0.0106867f $X=3.145 $Y=1.985 $X2=0 $Y2=0
cc_280 N_Y_c_420_n N_A_510_368#_c_489_n 0.039183f $X=3.145 $Y=1.985 $X2=0 $Y2=0
cc_281 N_Y_c_386_n N_A_27_74#_M1012_d 0.00218982f $X=1.615 $Y=1.095 $X2=0 $Y2=0
cc_282 N_Y_c_388_n N_A_27_74#_M1007_d 0.00272289f $X=2.16 $Y=1.18 $X2=0 $Y2=0
cc_283 N_Y_c_387_n N_A_27_74#_c_503_n 0.00540984f $X=0.945 $Y=1.095 $X2=0 $Y2=0
cc_284 N_Y_M1009_s N_A_27_74#_c_504_n 0.00288741f $X=0.57 $Y=0.37 $X2=0 $Y2=0
cc_285 N_Y_c_449_p N_A_27_74#_c_504_n 0.0200134f $X=0.78 $Y=0.76 $X2=0 $Y2=0
cc_286 N_Y_c_386_n N_A_27_74#_c_504_n 0.0036669f $X=1.615 $Y=1.095 $X2=0 $Y2=0
cc_287 N_Y_c_386_n N_A_27_74#_c_520_n 0.0183199f $X=1.615 $Y=1.095 $X2=0 $Y2=0
cc_288 N_Y_M1003_s N_A_27_74#_c_506_n 0.00250873f $X=1.57 $Y=0.37 $X2=0 $Y2=0
cc_289 N_Y_c_386_n N_A_27_74#_c_506_n 0.00612372f $X=1.615 $Y=1.095 $X2=0 $Y2=0
cc_290 N_Y_c_401_n N_A_27_74#_c_506_n 0.018913f $X=1.78 $Y=0.76 $X2=0 $Y2=0
cc_291 N_Y_c_401_n N_A_27_74#_c_512_n 0.00573111f $X=1.78 $Y=0.76 $X2=0 $Y2=0
cc_292 N_Y_c_390_n N_A_27_74#_c_512_n 0.00678392f $X=3.06 $Y=1.885 $X2=0 $Y2=0
cc_293 N_Y_c_388_n N_A_27_74#_c_512_n 0.0222436f $X=2.16 $Y=1.18 $X2=0 $Y2=0
cc_294 N_A_27_74#_c_507_n N_VGND_M1010_s 0.00218982f $X=3.505 $Y=1.045 $X2=-0.19
+ $Y2=-0.245
cc_295 N_A_27_74#_c_509_n N_VGND_M1001_s 0.00250873f $X=4.435 $Y=1.095 $X2=0
+ $Y2=0
cc_296 N_A_27_74#_c_507_n N_VGND_c_581_n 0.0185459f $X=3.505 $Y=1.045 $X2=0
+ $Y2=0
cc_297 N_A_27_74#_c_508_n N_VGND_c_581_n 0.00129215f $X=3.59 $Y=0.515 $X2=0
+ $Y2=0
cc_298 N_A_27_74#_c_512_n N_VGND_c_581_n 0.0254844f $X=2.69 $Y=0.965 $X2=0 $Y2=0
cc_299 N_A_27_74#_c_508_n N_VGND_c_582_n 0.0184106f $X=3.59 $Y=0.515 $X2=0 $Y2=0
cc_300 N_A_27_74#_c_509_n N_VGND_c_582_n 0.0209867f $X=4.435 $Y=1.095 $X2=0
+ $Y2=0
cc_301 N_A_27_74#_c_510_n N_VGND_c_582_n 0.0182902f $X=4.52 $Y=0.515 $X2=0 $Y2=0
cc_302 N_A_27_74#_c_504_n N_VGND_c_583_n 0.0423044f $X=1.115 $Y=0.34 $X2=0 $Y2=0
cc_303 N_A_27_74#_c_505_n N_VGND_c_583_n 0.0235688f $X=0.445 $Y=0.34 $X2=0 $Y2=0
cc_304 N_A_27_74#_c_506_n N_VGND_c_583_n 0.0423044f $X=2.115 $Y=0.34 $X2=0 $Y2=0
cc_305 N_A_27_74#_c_511_n N_VGND_c_583_n 0.0233048f $X=1.28 $Y=0.34 $X2=0 $Y2=0
cc_306 N_A_27_74#_c_512_n N_VGND_c_583_n 0.0477547f $X=2.69 $Y=0.965 $X2=0 $Y2=0
cc_307 N_A_27_74#_c_508_n N_VGND_c_584_n 0.0109942f $X=3.59 $Y=0.515 $X2=0 $Y2=0
cc_308 N_A_27_74#_c_510_n N_VGND_c_585_n 0.011066f $X=4.52 $Y=0.515 $X2=0 $Y2=0
cc_309 N_A_27_74#_c_504_n N_VGND_c_586_n 0.0239316f $X=1.115 $Y=0.34 $X2=0 $Y2=0
cc_310 N_A_27_74#_c_505_n N_VGND_c_586_n 0.0127152f $X=0.445 $Y=0.34 $X2=0 $Y2=0
cc_311 N_A_27_74#_c_506_n N_VGND_c_586_n 0.0239316f $X=2.115 $Y=0.34 $X2=0 $Y2=0
cc_312 N_A_27_74#_c_508_n N_VGND_c_586_n 0.00904371f $X=3.59 $Y=0.515 $X2=0
+ $Y2=0
cc_313 N_A_27_74#_c_510_n N_VGND_c_586_n 0.00915947f $X=4.52 $Y=0.515 $X2=0
+ $Y2=0
cc_314 N_A_27_74#_c_511_n N_VGND_c_586_n 0.0126653f $X=1.28 $Y=0.34 $X2=0 $Y2=0
cc_315 N_A_27_74#_c_512_n N_VGND_c_586_n 0.0259963f $X=2.69 $Y=0.965 $X2=0 $Y2=0
