* File: sky130_fd_sc_hs__clkdlyinv5sd1_1.pxi.spice
* Created: Thu Aug 27 20:36:24 2020
* 
x_PM_SKY130_FD_SC_HS__CLKDLYINV5SD1_1%A N_A_M1008_g N_A_c_81_n N_A_c_85_n
+ N_A_M1001_g A A N_A_c_83_n PM_SKY130_FD_SC_HS__CLKDLYINV5SD1_1%A
x_PM_SKY130_FD_SC_HS__CLKDLYINV5SD1_1%A_28_74# N_A_28_74#_M1008_s
+ N_A_28_74#_M1001_s N_A_28_74#_M1009_g N_A_28_74#_M1007_g N_A_28_74#_c_118_n
+ N_A_28_74#_c_119_n N_A_28_74#_c_120_n N_A_28_74#_c_125_n N_A_28_74#_c_126_n
+ N_A_28_74#_c_137_n N_A_28_74#_c_121_n N_A_28_74#_c_122_n N_A_28_74#_c_123_n
+ PM_SKY130_FD_SC_HS__CLKDLYINV5SD1_1%A_28_74#
x_PM_SKY130_FD_SC_HS__CLKDLYINV5SD1_1%A_288_74# N_A_288_74#_M1009_d
+ N_A_288_74#_M1007_d N_A_288_74#_M1003_g N_A_288_74#_M1000_g
+ N_A_288_74#_c_179_n N_A_288_74#_c_180_n N_A_288_74#_c_181_n
+ N_A_288_74#_c_182_n N_A_288_74#_c_183_n N_A_288_74#_c_187_n
+ N_A_288_74#_c_184_n PM_SKY130_FD_SC_HS__CLKDLYINV5SD1_1%A_288_74#
x_PM_SKY130_FD_SC_HS__CLKDLYINV5SD1_1%A_549_74# N_A_549_74#_M1003_d
+ N_A_549_74#_M1000_d N_A_549_74#_M1005_g N_A_549_74#_M1006_g
+ N_A_549_74#_c_223_n N_A_549_74#_c_224_n N_A_549_74#_c_225_n
+ N_A_549_74#_c_226_n N_A_549_74#_c_227_n N_A_549_74#_c_228_n
+ PM_SKY130_FD_SC_HS__CLKDLYINV5SD1_1%A_549_74#
x_PM_SKY130_FD_SC_HS__CLKDLYINV5SD1_1%A_682_74# N_A_682_74#_M1006_s
+ N_A_682_74#_M1005_s N_A_682_74#_M1004_g N_A_682_74#_c_271_n
+ N_A_682_74#_M1002_g N_A_682_74#_c_272_n N_A_682_74#_c_279_n
+ N_A_682_74#_c_273_n N_A_682_74#_c_274_n N_A_682_74#_c_275_n
+ N_A_682_74#_c_276_n N_A_682_74#_c_277_n
+ PM_SKY130_FD_SC_HS__CLKDLYINV5SD1_1%A_682_74#
x_PM_SKY130_FD_SC_HS__CLKDLYINV5SD1_1%VPWR N_VPWR_M1001_d N_VPWR_M1000_s
+ N_VPWR_M1005_d N_VPWR_c_327_n N_VPWR_c_328_n N_VPWR_c_329_n VPWR
+ N_VPWR_c_330_n N_VPWR_c_331_n N_VPWR_c_332_n N_VPWR_c_333_n N_VPWR_c_326_n
+ N_VPWR_c_335_n N_VPWR_c_336_n N_VPWR_c_337_n VPWR
+ PM_SKY130_FD_SC_HS__CLKDLYINV5SD1_1%VPWR
x_PM_SKY130_FD_SC_HS__CLKDLYINV5SD1_1%Y N_Y_M1004_d N_Y_M1002_d Y Y Y Y Y Y Y Y
+ PM_SKY130_FD_SC_HS__CLKDLYINV5SD1_1%Y
x_PM_SKY130_FD_SC_HS__CLKDLYINV5SD1_1%VGND N_VGND_M1008_d N_VGND_M1003_s
+ N_VGND_M1006_d N_VGND_c_393_n N_VGND_c_394_n N_VGND_c_395_n VGND
+ N_VGND_c_396_n N_VGND_c_397_n N_VGND_c_398_n N_VGND_c_399_n N_VGND_c_400_n
+ N_VGND_c_401_n N_VGND_c_402_n N_VGND_c_403_n VGND
+ PM_SKY130_FD_SC_HS__CLKDLYINV5SD1_1%VGND
cc_1 VNB N_A_M1008_g 0.0470676f $X=-0.19 $Y=-0.245 $X2=0.48 $Y2=0.58
cc_2 VNB N_A_c_81_n 0.00995999f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.675
cc_3 VNB A 0.0267916f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_4 VNB N_A_c_83_n 0.0365431f $X=-0.19 $Y=-0.245 $X2=0.57 $Y2=1.355
cc_5 VNB N_A_28_74#_M1009_g 0.0365884f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.4
cc_6 VNB N_A_28_74#_M1007_g 0.0120025f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_7 VNB N_A_28_74#_c_118_n 0.0375823f $X=-0.19 $Y=-0.245 $X2=0.57 $Y2=1.355
cc_8 VNB N_A_28_74#_c_119_n 0.0137526f $X=-0.19 $Y=-0.245 $X2=0.57 $Y2=1.355
cc_9 VNB N_A_28_74#_c_120_n 0.0226356f $X=-0.19 $Y=-0.245 $X2=0.415 $Y2=1.295
cc_10 VNB N_A_28_74#_c_121_n 0.0214092f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_28_74#_c_122_n 0.0121635f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_28_74#_c_123_n 0.00301793f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_288_74#_M1003_g 0.0459218f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.4
cc_14 VNB N_A_288_74#_M1000_g 0.015929f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_288_74#_c_179_n 0.0563825f $X=-0.19 $Y=-0.245 $X2=0.57 $Y2=1.355
cc_16 VNB N_A_288_74#_c_180_n 0.0131921f $X=-0.19 $Y=-0.245 $X2=0.57 $Y2=1.355
cc_17 VNB N_A_288_74#_c_181_n 0.0268697f $X=-0.19 $Y=-0.245 $X2=0.415 $Y2=1.295
cc_18 VNB N_A_288_74#_c_182_n 0.00978917f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_288_74#_c_183_n 0.0255344f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_288_74#_c_184_n 0.00614775f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_549_74#_M1005_g 0.0136178f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.4
cc_22 VNB N_A_549_74#_M1006_g 0.0409871f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_549_74#_c_223_n 0.0419063f $X=-0.19 $Y=-0.245 $X2=0.57 $Y2=1.355
cc_24 VNB N_A_549_74#_c_224_n 0.0134245f $X=-0.19 $Y=-0.245 $X2=0.57 $Y2=1.355
cc_25 VNB N_A_549_74#_c_225_n 0.0155677f $X=-0.19 $Y=-0.245 $X2=0.415 $Y2=1.295
cc_26 VNB N_A_549_74#_c_226_n 0.0111173f $X=-0.19 $Y=-0.245 $X2=0.415 $Y2=1.665
cc_27 VNB N_A_549_74#_c_227_n 0.0372738f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_549_74#_c_228_n 0.00227058f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_682_74#_M1004_g 0.0444659f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.4
cc_30 VNB N_A_682_74#_c_271_n 0.0391593f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_31 VNB N_A_682_74#_c_272_n 0.00817528f $X=-0.19 $Y=-0.245 $X2=0.57 $Y2=1.355
cc_32 VNB N_A_682_74#_c_273_n 0.00706738f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_682_74#_c_274_n 0.00422437f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_682_74#_c_275_n 0.0273095f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_682_74#_c_276_n 0.0067964f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_682_74#_c_277_n 0.00272046f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_VPWR_c_326_n 0.223389f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB Y 0.0204118f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.765
cc_39 VNB Y 0.0466962f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.4
cc_40 VNB N_VGND_c_393_n 0.00990754f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_394_n 0.0149646f $X=-0.19 $Y=-0.245 $X2=0.57 $Y2=1.355
cc_42 VNB N_VGND_c_395_n 0.00662038f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_396_n 0.0180717f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_397_n 0.0296852f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_VGND_c_398_n 0.0621707f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_VGND_c_399_n 0.0189455f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_VGND_c_400_n 0.347307f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_VGND_c_401_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_VGND_c_402_n 0.00673217f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_VGND_c_403_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VPB N_A_c_81_n 0.00100316f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.675
cc_52 VPB N_A_c_85_n 0.0286879f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.765
cc_53 VPB A 0.0108255f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.21
cc_54 VPB N_A_28_74#_M1007_g 0.0334201f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_55 VPB N_A_28_74#_c_125_n 0.0079884f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_56 VPB N_A_28_74#_c_126_n 0.0205617f $X=-0.19 $Y=1.66 $X2=0.415 $Y2=1.665
cc_57 VPB N_A_28_74#_c_123_n 0.00436726f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_58 VPB N_A_288_74#_M1000_g 0.040832f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_59 VPB N_A_288_74#_c_182_n 0.02236f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_60 VPB N_A_288_74#_c_187_n 0.00306613f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_61 VPB N_A_549_74#_M1005_g 0.0358586f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=2.4
cc_62 VPB N_A_549_74#_c_226_n 0.0106835f $X=-0.19 $Y=1.66 $X2=0.415 $Y2=1.665
cc_63 VPB N_A_682_74#_c_271_n 0.0254953f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_64 VPB N_A_682_74#_c_279_n 0.00990629f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_65 VPB N_A_682_74#_c_273_n 0.0212578f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_66 VPB N_A_682_74#_c_274_n 0.00141791f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_67 VPB N_VPWR_c_327_n 0.0103216f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_68 VPB N_VPWR_c_328_n 0.026197f $X=-0.19 $Y=1.66 $X2=0.57 $Y2=1.355
cc_69 VPB N_VPWR_c_329_n 0.00777218f $X=-0.19 $Y=1.66 $X2=0.415 $Y2=1.355
cc_70 VPB N_VPWR_c_330_n 0.018958f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_71 VPB N_VPWR_c_331_n 0.0298867f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_72 VPB N_VPWR_c_332_n 0.0624644f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_73 VPB N_VPWR_c_333_n 0.0184442f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_74 VPB N_VPWR_c_326_n 0.136759f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_75 VPB N_VPWR_c_335_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_76 VPB N_VPWR_c_336_n 0.00670627f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_77 VPB N_VPWR_c_337_n 0.00614127f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_78 VPB Y 0.0121098f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=2.4
cc_79 VPB Y 0.0526708f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.21
cc_80 A N_A_28_74#_M1001_s 0.00256075f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_81 N_A_c_81_n N_A_28_74#_M1007_g 0.00227483f $X=0.495 $Y=1.675 $X2=0 $Y2=0
cc_82 A N_A_28_74#_M1007_g 0.00110625f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_83 N_A_c_83_n N_A_28_74#_M1007_g 8.99867e-19 $X=0.57 $Y=1.355 $X2=0 $Y2=0
cc_84 N_A_M1008_g N_A_28_74#_c_118_n 0.0021171f $X=0.48 $Y=0.58 $X2=0 $Y2=0
cc_85 A N_A_28_74#_c_118_n 0.00102763f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_86 N_A_c_83_n N_A_28_74#_c_118_n 0.0170907f $X=0.57 $Y=1.355 $X2=0 $Y2=0
cc_87 N_A_M1008_g N_A_28_74#_c_120_n 0.0127782f $X=0.48 $Y=0.58 $X2=0 $Y2=0
cc_88 A N_A_28_74#_c_125_n 0.0237727f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_89 N_A_c_85_n N_A_28_74#_c_137_n 0.0152432f $X=0.495 $Y=1.765 $X2=0 $Y2=0
cc_90 A N_A_28_74#_c_137_n 0.0197054f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_91 N_A_c_83_n N_A_28_74#_c_137_n 6.00585e-19 $X=0.57 $Y=1.355 $X2=0 $Y2=0
cc_92 N_A_M1008_g N_A_28_74#_c_121_n 0.0127534f $X=0.48 $Y=0.58 $X2=0 $Y2=0
cc_93 A N_A_28_74#_c_121_n 0.0251751f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_94 N_A_c_83_n N_A_28_74#_c_121_n 0.00146806f $X=0.57 $Y=1.355 $X2=0 $Y2=0
cc_95 N_A_M1008_g N_A_28_74#_c_122_n 0.00415005f $X=0.48 $Y=0.58 $X2=0 $Y2=0
cc_96 A N_A_28_74#_c_122_n 0.0289843f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_97 N_A_M1008_g N_A_28_74#_c_123_n 0.00344321f $X=0.48 $Y=0.58 $X2=0 $Y2=0
cc_98 N_A_c_81_n N_A_28_74#_c_123_n 8.33404e-19 $X=0.495 $Y=1.675 $X2=0 $Y2=0
cc_99 N_A_c_85_n N_A_28_74#_c_123_n 0.0053811f $X=0.495 $Y=1.765 $X2=0 $Y2=0
cc_100 A N_A_28_74#_c_123_n 0.0427389f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_101 N_A_c_83_n N_A_28_74#_c_123_n 0.00146966f $X=0.57 $Y=1.355 $X2=0 $Y2=0
cc_102 A N_VPWR_M1001_d 0.00136529f $X=0.155 $Y=1.21 $X2=-0.19 $Y2=-0.245
cc_103 N_A_c_85_n N_VPWR_c_327_n 0.00571996f $X=0.495 $Y=1.765 $X2=0 $Y2=0
cc_104 N_A_c_85_n N_VPWR_c_330_n 0.00461464f $X=0.495 $Y=1.765 $X2=0 $Y2=0
cc_105 N_A_c_85_n N_VPWR_c_326_n 0.00915869f $X=0.495 $Y=1.765 $X2=0 $Y2=0
cc_106 N_A_M1008_g N_VGND_c_393_n 0.00427883f $X=0.48 $Y=0.58 $X2=0 $Y2=0
cc_107 N_A_M1008_g N_VGND_c_396_n 0.00456766f $X=0.48 $Y=0.58 $X2=0 $Y2=0
cc_108 N_A_M1008_g N_VGND_c_400_n 0.00458574f $X=0.48 $Y=0.58 $X2=0 $Y2=0
cc_109 N_A_28_74#_M1009_g N_A_288_74#_c_181_n 0.0106652f $X=1.365 $Y=0.58 $X2=0
+ $Y2=0
cc_110 N_A_28_74#_c_119_n N_A_288_74#_c_181_n 2.87835e-19 $X=1.367 $Y=1.295
+ $X2=0 $Y2=0
cc_111 N_A_28_74#_c_121_n N_A_288_74#_c_181_n 0.0164122f $X=0.975 $Y=0.92 $X2=0
+ $Y2=0
cc_112 N_A_28_74#_c_123_n N_A_288_74#_c_181_n 0.00916028f $X=1.14 $Y=1.295 $X2=0
+ $Y2=0
cc_113 N_A_28_74#_M1007_g N_A_288_74#_c_182_n 0.0112394f $X=1.37 $Y=2.46 $X2=0
+ $Y2=0
cc_114 N_A_28_74#_c_123_n N_A_288_74#_c_182_n 0.0406706f $X=1.14 $Y=1.295 $X2=0
+ $Y2=0
cc_115 N_A_28_74#_M1007_g N_A_288_74#_c_187_n 0.0065242f $X=1.37 $Y=2.46 $X2=0
+ $Y2=0
cc_116 N_A_28_74#_c_119_n N_A_288_74#_c_184_n 0.0098227f $X=1.367 $Y=1.295 $X2=0
+ $Y2=0
cc_117 N_A_28_74#_c_123_n N_A_288_74#_c_184_n 0.0277877f $X=1.14 $Y=1.295 $X2=0
+ $Y2=0
cc_118 N_A_28_74#_c_137_n N_VPWR_M1001_d 0.0305614f $X=0.975 $Y=2.117 $X2=-0.19
+ $Y2=-0.245
cc_119 N_A_28_74#_c_123_n N_VPWR_M1001_d 0.00158821f $X=1.14 $Y=1.295 $X2=-0.19
+ $Y2=-0.245
cc_120 N_A_28_74#_M1007_g N_VPWR_c_327_n 0.0149559f $X=1.37 $Y=2.46 $X2=0 $Y2=0
cc_121 N_A_28_74#_c_137_n N_VPWR_c_327_n 0.0220956f $X=0.975 $Y=2.117 $X2=0
+ $Y2=0
cc_122 N_A_28_74#_M1007_g N_VPWR_c_328_n 0.00438706f $X=1.37 $Y=2.46 $X2=0 $Y2=0
cc_123 N_A_28_74#_c_126_n N_VPWR_c_330_n 0.00593336f $X=0.265 $Y=2.56 $X2=0
+ $Y2=0
cc_124 N_A_28_74#_M1007_g N_VPWR_c_331_n 0.00430639f $X=1.37 $Y=2.46 $X2=0 $Y2=0
cc_125 N_A_28_74#_M1007_g N_VPWR_c_326_n 0.00815045f $X=1.37 $Y=2.46 $X2=0 $Y2=0
cc_126 N_A_28_74#_c_126_n N_VPWR_c_326_n 0.00940928f $X=0.265 $Y=2.56 $X2=0
+ $Y2=0
cc_127 N_A_28_74#_M1009_g N_VGND_c_393_n 0.00830587f $X=1.365 $Y=0.58 $X2=0
+ $Y2=0
cc_128 N_A_28_74#_c_120_n N_VGND_c_393_n 0.0151665f $X=0.265 $Y=0.58 $X2=0 $Y2=0
cc_129 N_A_28_74#_c_121_n N_VGND_c_393_n 0.0255952f $X=0.975 $Y=0.92 $X2=0 $Y2=0
cc_130 N_A_28_74#_M1009_g N_VGND_c_394_n 0.00244567f $X=1.365 $Y=0.58 $X2=0
+ $Y2=0
cc_131 N_A_28_74#_c_120_n N_VGND_c_396_n 0.0170785f $X=0.265 $Y=0.58 $X2=0 $Y2=0
cc_132 N_A_28_74#_M1009_g N_VGND_c_397_n 0.00461464f $X=1.365 $Y=0.58 $X2=0
+ $Y2=0
cc_133 N_A_28_74#_M1009_g N_VGND_c_400_n 0.00874319f $X=1.365 $Y=0.58 $X2=0
+ $Y2=0
cc_134 N_A_28_74#_c_120_n N_VGND_c_400_n 0.0118627f $X=0.265 $Y=0.58 $X2=0 $Y2=0
cc_135 N_A_28_74#_c_121_n N_VGND_c_400_n 0.0215989f $X=0.975 $Y=0.92 $X2=0 $Y2=0
cc_136 N_A_288_74#_M1003_g N_A_549_74#_c_225_n 0.0162175f $X=2.67 $Y=0.58 $X2=0
+ $Y2=0
cc_137 N_A_288_74#_c_183_n N_A_549_74#_c_225_n 0.00419423f $X=2.425 $Y=1.305
+ $X2=0 $Y2=0
cc_138 N_A_288_74#_c_180_n N_A_549_74#_c_226_n 0.0216563f $X=2.67 $Y=1.305 $X2=0
+ $Y2=0
cc_139 N_A_288_74#_c_183_n N_A_549_74#_c_226_n 0.00419423f $X=2.425 $Y=1.305
+ $X2=0 $Y2=0
cc_140 N_A_288_74#_c_180_n N_A_549_74#_c_228_n 0.00534783f $X=2.67 $Y=1.305
+ $X2=0 $Y2=0
cc_141 N_A_288_74#_c_183_n N_A_549_74#_c_228_n 0.0101411f $X=2.425 $Y=1.305
+ $X2=0 $Y2=0
cc_142 N_A_288_74#_c_187_n N_VPWR_c_327_n 0.00826281f $X=1.58 $Y=2.815 $X2=0
+ $Y2=0
cc_143 N_A_288_74#_M1000_g N_VPWR_c_328_n 0.0237278f $X=2.67 $Y=2.46 $X2=0 $Y2=0
cc_144 N_A_288_74#_c_179_n N_VPWR_c_328_n 3.64176e-19 $X=2.595 $Y=1.305 $X2=0
+ $Y2=0
cc_145 N_A_288_74#_c_182_n N_VPWR_c_328_n 0.0793707f $X=1.58 $Y=2.105 $X2=0
+ $Y2=0
cc_146 N_A_288_74#_c_183_n N_VPWR_c_328_n 0.0151215f $X=2.425 $Y=1.305 $X2=0
+ $Y2=0
cc_147 N_A_288_74#_c_187_n N_VPWR_c_331_n 0.00976575f $X=1.58 $Y=2.815 $X2=0
+ $Y2=0
cc_148 N_A_288_74#_M1000_g N_VPWR_c_332_n 0.00461464f $X=2.67 $Y=2.46 $X2=0
+ $Y2=0
cc_149 N_A_288_74#_M1000_g N_VPWR_c_326_n 0.00919316f $X=2.67 $Y=2.46 $X2=0
+ $Y2=0
cc_150 N_A_288_74#_c_187_n N_VPWR_c_326_n 0.0112865f $X=1.58 $Y=2.815 $X2=0
+ $Y2=0
cc_151 N_A_288_74#_c_181_n N_VGND_c_393_n 0.00689376f $X=1.58 $Y=0.58 $X2=0
+ $Y2=0
cc_152 N_A_288_74#_M1003_g N_VGND_c_394_n 0.0119093f $X=2.67 $Y=0.58 $X2=0 $Y2=0
cc_153 N_A_288_74#_c_179_n N_VGND_c_394_n 3.84795e-19 $X=2.595 $Y=1.305 $X2=0
+ $Y2=0
cc_154 N_A_288_74#_c_181_n N_VGND_c_394_n 0.0326862f $X=1.58 $Y=0.58 $X2=0 $Y2=0
cc_155 N_A_288_74#_c_183_n N_VGND_c_394_n 0.0165176f $X=2.425 $Y=1.305 $X2=0
+ $Y2=0
cc_156 N_A_288_74#_c_181_n N_VGND_c_397_n 0.0132196f $X=1.58 $Y=0.58 $X2=0 $Y2=0
cc_157 N_A_288_74#_M1003_g N_VGND_c_398_n 0.00461464f $X=2.67 $Y=0.58 $X2=0
+ $Y2=0
cc_158 N_A_288_74#_M1003_g N_VGND_c_400_n 0.00919316f $X=2.67 $Y=0.58 $X2=0
+ $Y2=0
cc_159 N_A_288_74#_c_181_n N_VGND_c_400_n 0.00920999f $X=1.58 $Y=0.58 $X2=0
+ $Y2=0
cc_160 N_A_549_74#_M1006_g N_A_682_74#_M1004_g 0.0191451f $X=4.1 $Y=0.58 $X2=0
+ $Y2=0
cc_161 N_A_549_74#_M1005_g N_A_682_74#_c_271_n 0.0182884f $X=4.095 $Y=2.46 $X2=0
+ $Y2=0
cc_162 N_A_549_74#_c_224_n N_A_682_74#_c_271_n 0.0128901f $X=4.02 $Y=1.14 $X2=0
+ $Y2=0
cc_163 N_A_549_74#_c_227_n N_A_682_74#_c_271_n 2.99954e-19 $X=3.84 $Y=1.305
+ $X2=0 $Y2=0
cc_164 N_A_549_74#_M1006_g N_A_682_74#_c_272_n 0.0120746f $X=4.1 $Y=0.58 $X2=0
+ $Y2=0
cc_165 N_A_549_74#_c_225_n N_A_682_74#_c_272_n 0.0198272f $X=2.885 $Y=0.58 $X2=0
+ $Y2=0
cc_166 N_A_549_74#_M1005_g N_A_682_74#_c_279_n 0.0256928f $X=4.095 $Y=2.46 $X2=0
+ $Y2=0
cc_167 N_A_549_74#_c_226_n N_A_682_74#_c_279_n 0.046582f $X=2.885 $Y=2.105 $X2=0
+ $Y2=0
cc_168 N_A_549_74#_M1005_g N_A_682_74#_c_273_n 0.0191499f $X=4.095 $Y=2.46 $X2=0
+ $Y2=0
cc_169 N_A_549_74#_c_223_n N_A_682_74#_c_273_n 0.00866615f $X=4.02 $Y=1.305
+ $X2=0 $Y2=0
cc_170 N_A_549_74#_c_227_n N_A_682_74#_c_273_n 0.02505f $X=3.84 $Y=1.305 $X2=0
+ $Y2=0
cc_171 N_A_549_74#_c_226_n N_A_682_74#_c_274_n 0.0073655f $X=2.885 $Y=2.105
+ $X2=0 $Y2=0
cc_172 N_A_549_74#_c_227_n N_A_682_74#_c_274_n 0.0202705f $X=3.84 $Y=1.305 $X2=0
+ $Y2=0
cc_173 N_A_549_74#_M1006_g N_A_682_74#_c_275_n 0.0191653f $X=4.1 $Y=0.58 $X2=0
+ $Y2=0
cc_174 N_A_549_74#_c_223_n N_A_682_74#_c_275_n 0.00808945f $X=4.02 $Y=1.305
+ $X2=0 $Y2=0
cc_175 N_A_549_74#_c_227_n N_A_682_74#_c_275_n 0.021775f $X=3.84 $Y=1.305 $X2=0
+ $Y2=0
cc_176 N_A_549_74#_c_223_n N_A_682_74#_c_276_n 7.67879e-19 $X=4.02 $Y=1.305
+ $X2=0 $Y2=0
cc_177 N_A_549_74#_c_225_n N_A_682_74#_c_276_n 0.0079307f $X=2.885 $Y=0.58 $X2=0
+ $Y2=0
cc_178 N_A_549_74#_c_227_n N_A_682_74#_c_276_n 0.0276549f $X=3.84 $Y=1.305 $X2=0
+ $Y2=0
cc_179 N_A_549_74#_M1006_g N_A_682_74#_c_277_n 0.00399027f $X=4.1 $Y=0.58 $X2=0
+ $Y2=0
cc_180 N_A_549_74#_c_224_n N_A_682_74#_c_277_n 0.0014721f $X=4.02 $Y=1.14 $X2=0
+ $Y2=0
cc_181 N_A_549_74#_c_227_n N_A_682_74#_c_277_n 0.00545692f $X=3.84 $Y=1.305
+ $X2=0 $Y2=0
cc_182 N_A_549_74#_c_226_n N_VPWR_c_328_n 0.0186311f $X=2.885 $Y=2.105 $X2=0
+ $Y2=0
cc_183 N_A_549_74#_M1005_g N_VPWR_c_329_n 0.0177733f $X=4.095 $Y=2.46 $X2=0
+ $Y2=0
cc_184 N_A_549_74#_M1005_g N_VPWR_c_332_n 0.00461464f $X=4.095 $Y=2.46 $X2=0
+ $Y2=0
cc_185 N_A_549_74#_c_226_n N_VPWR_c_332_n 0.00749631f $X=2.885 $Y=2.105 $X2=0
+ $Y2=0
cc_186 N_A_549_74#_M1005_g N_VPWR_c_326_n 0.00915948f $X=4.095 $Y=2.46 $X2=0
+ $Y2=0
cc_187 N_A_549_74#_c_226_n N_VPWR_c_326_n 0.0062048f $X=2.885 $Y=2.105 $X2=0
+ $Y2=0
cc_188 N_A_549_74#_M1006_g N_VGND_c_395_n 0.00771808f $X=4.1 $Y=0.58 $X2=0 $Y2=0
cc_189 N_A_549_74#_M1006_g N_VGND_c_398_n 0.00461464f $X=4.1 $Y=0.58 $X2=0 $Y2=0
cc_190 N_A_549_74#_c_225_n N_VGND_c_398_n 0.00573605f $X=2.885 $Y=0.58 $X2=0
+ $Y2=0
cc_191 N_A_549_74#_M1006_g N_VGND_c_400_n 0.00915849f $X=4.1 $Y=0.58 $X2=0 $Y2=0
cc_192 N_A_549_74#_c_225_n N_VGND_c_400_n 0.00594877f $X=2.885 $Y=0.58 $X2=0
+ $Y2=0
cc_193 N_A_682_74#_c_271_n N_VPWR_c_329_n 0.0163879f $X=4.72 $Y=1.765 $X2=0
+ $Y2=0
cc_194 N_A_682_74#_c_279_n N_VPWR_c_329_n 0.0299754f $X=3.535 $Y=2.105 $X2=0
+ $Y2=0
cc_195 N_A_682_74#_c_273_n N_VPWR_c_329_n 0.0255637f $X=4.53 $Y=1.645 $X2=0
+ $Y2=0
cc_196 N_A_682_74#_c_279_n N_VPWR_c_332_n 0.0106198f $X=3.535 $Y=2.105 $X2=0
+ $Y2=0
cc_197 N_A_682_74#_c_271_n N_VPWR_c_333_n 0.00413917f $X=4.72 $Y=1.765 $X2=0
+ $Y2=0
cc_198 N_A_682_74#_c_271_n N_VPWR_c_326_n 0.00821389f $X=4.72 $Y=1.765 $X2=0
+ $Y2=0
cc_199 N_A_682_74#_c_279_n N_VPWR_c_326_n 0.00879013f $X=3.535 $Y=2.105 $X2=0
+ $Y2=0
cc_200 N_A_682_74#_M1004_g Y 8.21909e-19 $X=4.71 $Y=0.58 $X2=0 $Y2=0
cc_201 N_A_682_74#_M1004_g Y 0.0124475f $X=4.71 $Y=0.58 $X2=0 $Y2=0
cc_202 N_A_682_74#_c_271_n Y 0.0163621f $X=4.72 $Y=1.765 $X2=0 $Y2=0
cc_203 N_A_682_74#_c_273_n Y 0.0140324f $X=4.53 $Y=1.645 $X2=0 $Y2=0
cc_204 N_A_682_74#_c_275_n Y 0.0133247f $X=4.53 $Y=0.965 $X2=0 $Y2=0
cc_205 N_A_682_74#_c_277_n Y 0.0384675f $X=4.67 $Y=1.46 $X2=0 $Y2=0
cc_206 N_A_682_74#_c_271_n Y 0.00229934f $X=4.72 $Y=1.765 $X2=0 $Y2=0
cc_207 N_A_682_74#_M1004_g N_VGND_c_395_n 0.0112059f $X=4.71 $Y=0.58 $X2=0 $Y2=0
cc_208 N_A_682_74#_c_271_n N_VGND_c_395_n 3.24916e-19 $X=4.72 $Y=1.765 $X2=0
+ $Y2=0
cc_209 N_A_682_74#_c_272_n N_VGND_c_395_n 0.0080629f $X=3.535 $Y=0.565 $X2=0
+ $Y2=0
cc_210 N_A_682_74#_c_275_n N_VGND_c_395_n 0.0218411f $X=4.53 $Y=0.965 $X2=0
+ $Y2=0
cc_211 N_A_682_74#_c_272_n N_VGND_c_398_n 0.0118185f $X=3.535 $Y=0.565 $X2=0
+ $Y2=0
cc_212 N_A_682_74#_M1004_g N_VGND_c_399_n 0.00383152f $X=4.71 $Y=0.58 $X2=0
+ $Y2=0
cc_213 N_A_682_74#_M1004_g N_VGND_c_400_n 0.00761428f $X=4.71 $Y=0.58 $X2=0
+ $Y2=0
cc_214 N_A_682_74#_c_272_n N_VGND_c_400_n 0.0117223f $X=3.535 $Y=0.565 $X2=0
+ $Y2=0
cc_215 N_VPWR_c_329_n Y 0.0476994f $X=4.495 $Y=1.985 $X2=0 $Y2=0
cc_216 N_VPWR_c_333_n Y 0.0234396f $X=5.04 $Y=3.33 $X2=0 $Y2=0
cc_217 N_VPWR_c_326_n Y 0.0138183f $X=5.04 $Y=3.33 $X2=0 $Y2=0
cc_218 Y N_VGND_c_395_n 0.0124097f $X=4.95 $Y=0.47 $X2=0 $Y2=0
cc_219 Y N_VGND_c_399_n 0.0155069f $X=4.95 $Y=0.47 $X2=0 $Y2=0
cc_220 Y N_VGND_c_400_n 0.013122f $X=4.95 $Y=0.47 $X2=0 $Y2=0
