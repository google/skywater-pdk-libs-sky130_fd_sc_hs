* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hs__a31oi_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
M1000 Y A1 a_475_74# VNB nlowvt w=740000u l=150000u
+  ad=9.2695e+11p pd=8.48e+06u as=1.1544e+12p ps=9.04e+06u
M1001 a_475_74# A2 a_30_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=1.03482e+12p ps=1.022e+07u
M1002 a_475_74# A1 Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1003 Y B1 a_27_368# VPB pshort w=1.12e+06u l=150000u
+  ad=6.944e+11p pd=5.72e+06u as=3.696e+12p ps=2.676e+07u
M1004 a_30_74# A2 a_475_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_30_74# A3 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=1.2839e+12p ps=7.91e+06u
M1006 a_27_368# A3 VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=2.296e+12p ps=1.754e+07u
M1007 VGND A3 a_30_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_30_74# A2 a_475_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 Y B1 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VPWR A3 a_27_368# VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VPWR A3 a_27_368# VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_475_74# A1 Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_27_368# A3 VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_27_368# A2 VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_27_368# A1 VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_27_368# A1 VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 Y A1 a_475_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 VPWR A2 a_27_368# VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VPWR A1 a_27_368# VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 VPWR A2 a_27_368# VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_27_368# A2 VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_27_368# B1 Y VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_475_74# A2 a_30_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 VPWR A1 a_27_368# VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 Y B1 a_27_368# VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 a_27_368# B1 Y VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 VGND B1 Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1028 VGND A3 a_30_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1029 a_30_74# A3 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
