* File: sky130_fd_sc_hs__o21ba_4.spice
* Created: Thu Aug 27 20:58:38 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hs__o21ba_4.pex.spice"
.subckt sky130_fd_sc_hs__o21ba_4  VNB VPB B1_N A2 A1 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A1	A1
* A2	A2
* B1_N	B1_N
* VPB	VPB
* VNB	VNB
MM1021 N_VGND_M1021_d N_B1_N_M1021_g N_A_27_368#_M1021_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.13505 AS=0.2109 PD=1.105 PS=2.05 NRD=11.34 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75002 A=0.111 P=1.78 MULT=1
MM1002 N_VGND_M1021_d N_A_193_48#_M1002_g N_X_M1002_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.13505 AS=0.1073 PD=1.105 PS=1.03 NRD=2.424 NRS=0 M=1 R=4.93333 SA=75000.7
+ SB=75001.5 A=0.111 P=1.78 MULT=1
MM1005 N_VGND_M1005_d N_A_193_48#_M1005_g N_X_M1002_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1073 PD=1.02 PS=1.03 NRD=0 NRS=1.62 M=1 R=4.93333 SA=75001.2
+ SB=75001.1 A=0.111 P=1.78 MULT=1
MM1013 N_VGND_M1005_d N_A_193_48#_M1013_g N_X_M1013_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.6
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1020 N_VGND_M1020_d N_A_193_48#_M1020_g N_X_M1013_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.1036 PD=2.05 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75002
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1007 N_A_193_48#_M1007_d N_A_27_368#_M1007_g N_A_618_94#_M1007_s VNB NLOWVT
+ L=0.15 W=0.64 AD=0.0896 AS=0.1824 PD=0.92 PS=1.85 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75002 A=0.096 P=1.58 MULT=1
MM1019 N_A_193_48#_M1007_d N_A_27_368#_M1019_g N_A_618_94#_M1019_s VNB NLOWVT
+ L=0.15 W=0.64 AD=0.0896 AS=0.123625 PD=0.92 PS=1.145 NRD=0 NRS=13.116 M=1
+ R=4.26667 SA=75000.6 SB=75001.6 A=0.096 P=1.58 MULT=1
MM1006 N_A_618_94#_M1019_s N_A1_M1006_g N_VGND_M1006_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.123625 AS=0.112 PD=1.145 PS=0.99 NRD=0 NRS=13.116 M=1 R=4.26667
+ SA=75000.9 SB=75001.6 A=0.096 P=1.58 MULT=1
MM1003 N_VGND_M1006_s N_A2_M1003_g N_A_618_94#_M1003_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.112 AS=0.0896 PD=0.99 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667 SA=75001.4
+ SB=75001.1 A=0.096 P=1.58 MULT=1
MM1009 N_VGND_M1009_d N_A2_M1009_g N_A_618_94#_M1003_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.0896 AS=0.0896 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667 SA=75001.8
+ SB=75000.6 A=0.096 P=1.58 MULT=1
MM1010 N_A_618_94#_M1010_d N_A1_M1010_g N_VGND_M1009_d VNB NLOWVT L=0.15 W=0.64
+ AD=0.1856 AS=0.0896 PD=1.86 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667 SA=75002.3
+ SB=75000.2 A=0.096 P=1.58 MULT=1
MM1016 N_VPWR_M1016_d N_B1_N_M1016_g N_A_27_368#_M1016_s VPB PSHORT L=0.15
+ W=1.12 AD=0.224 AS=0.3304 PD=1.52 PS=2.83 NRD=14.9326 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75004.6 A=0.168 P=2.54 MULT=1
MM1011 N_X_M1011_d N_A_193_48#_M1011_g N_VPWR_M1016_d VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.224 PD=1.42 PS=1.52 NRD=1.7533 NRS=6.1464 M=1 R=7.46667
+ SA=75000.8 SB=75004.1 A=0.168 P=2.54 MULT=1
MM1012 N_X_M1011_d N_A_193_48#_M1012_g N_VPWR_M1012_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.2 SB=75003.6 A=0.168 P=2.54 MULT=1
MM1014 N_X_M1014_d N_A_193_48#_M1014_g N_VPWR_M1012_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.7 SB=75003.2 A=0.168 P=2.54 MULT=1
MM1017 N_X_M1014_d N_A_193_48#_M1017_g N_VPWR_M1017_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.424 PD=1.42 PS=2.18857 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75002.1 SB=75002.7 A=0.168 P=2.54 MULT=1
MM1000 N_A_193_48#_M1000_d N_A_27_368#_M1000_g N_VPWR_M1017_s VPB PSHORT L=0.15
+ W=0.84 AD=0.126 AS=0.318 PD=1.14 PS=1.64143 NRD=2.3443 NRS=22.261 M=1 R=5.6
+ SA=75003.1 SB=75002.6 A=0.126 P=1.98 MULT=1
MM1001 N_A_193_48#_M1000_d N_A_27_368#_M1001_g N_VPWR_M1001_s VPB PSHORT L=0.15
+ W=0.84 AD=0.126 AS=0.18617 PD=1.14 PS=1.31022 NRD=2.3443 NRS=22.261 M=1 R=5.6
+ SA=75003.5 SB=75002.2 A=0.126 P=1.98 MULT=1
MM1004 N_A_892_392#_M1004_d N_A1_M1004_g N_VPWR_M1001_s VPB PSHORT L=0.15 W=1
+ AD=0.15 AS=0.22163 PD=1.3 PS=1.55978 NRD=1.9503 NRS=11.8003 M=1 R=6.66667
+ SA=75003.5 SB=75001.6 A=0.15 P=2.3 MULT=1
MM1008 N_A_193_48#_M1008_d N_A2_M1008_g N_A_892_392#_M1004_d VPB PSHORT L=0.15
+ W=1 AD=0.15 AS=0.15 PD=1.3 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=6.66667
+ SA=75003.9 SB=75001.1 A=0.15 P=2.3 MULT=1
MM1015 N_A_193_48#_M1008_d N_A2_M1015_g N_A_892_392#_M1015_s VPB PSHORT L=0.15
+ W=1 AD=0.15 AS=0.15 PD=1.3 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=6.66667
+ SA=75004.4 SB=75000.7 A=0.15 P=2.3 MULT=1
MM1018 N_A_892_392#_M1015_s N_A1_M1018_g N_VPWR_M1018_s VPB PSHORT L=0.15 W=1
+ AD=0.15 AS=0.295 PD=1.3 PS=2.59 NRD=1.9503 NRS=1.9503 M=1 R=6.66667 SA=75004.8
+ SB=75000.2 A=0.15 P=2.3 MULT=1
DX22_noxref VNB VPB NWDIODE A=12.3132 P=16.96
c_114 VPB 0 4.78765e-20 $X=0 $Y=3.085
*
.include "sky130_fd_sc_hs__o21ba_4.pxi.spice"
*
.ends
*
*
