* File: sky130_fd_sc_hs__or4_4.pxi.spice
* Created: Thu Aug 27 21:06:53 2020
* 
x_PM_SKY130_FD_SC_HS__OR4_4%A_83_264# N_A_83_264#_M1003_d N_A_83_264#_M1015_d
+ N_A_83_264#_M1014_d N_A_83_264#_c_120_n N_A_83_264#_M1010_g
+ N_A_83_264#_M1002_g N_A_83_264#_c_121_n N_A_83_264#_M1011_g
+ N_A_83_264#_M1004_g N_A_83_264#_c_122_n N_A_83_264#_M1012_g
+ N_A_83_264#_M1006_g N_A_83_264#_c_123_n N_A_83_264#_M1016_g
+ N_A_83_264#_M1007_g N_A_83_264#_c_112_n N_A_83_264#_c_113_n
+ N_A_83_264#_c_130_p N_A_83_264#_c_256_p N_A_83_264#_c_114_n
+ N_A_83_264#_c_137_p N_A_83_264#_c_115_n N_A_83_264#_c_116_n
+ N_A_83_264#_c_124_n N_A_83_264#_c_117_n N_A_83_264#_c_118_n
+ N_A_83_264#_c_136_p N_A_83_264#_c_119_n N_A_83_264#_c_127_n
+ PM_SKY130_FD_SC_HS__OR4_4%A_83_264#
x_PM_SKY130_FD_SC_HS__OR4_4%B N_B_c_267_n N_B_c_268_n N_B_c_276_n N_B_M1009_g
+ N_B_c_269_n N_B_M1003_g N_B_c_270_n N_B_c_278_n N_B_M1019_g N_B_c_271_n
+ N_B_c_272_n N_B_c_273_n N_B_c_274_n B B PM_SKY130_FD_SC_HS__OR4_4%B
x_PM_SKY130_FD_SC_HS__OR4_4%A N_A_M1013_g N_A_c_357_n N_A_M1000_g N_A_c_358_n
+ N_A_M1001_g A N_A_c_356_n PM_SKY130_FD_SC_HS__OR4_4%A
x_PM_SKY130_FD_SC_HS__OR4_4%C N_C_M1015_g N_C_c_403_n N_C_M1008_g N_C_c_404_n
+ N_C_M1018_g C C C N_C_c_405_n N_C_c_406_n PM_SKY130_FD_SC_HS__OR4_4%C
x_PM_SKY130_FD_SC_HS__OR4_4%D N_D_c_466_n N_D_M1005_g N_D_c_467_n N_D_c_476_n
+ N_D_M1014_g N_D_c_468_n N_D_c_478_n N_D_M1017_g N_D_c_469_n N_D_c_470_n
+ N_D_c_471_n N_D_c_472_n D N_D_c_473_n N_D_c_474_n PM_SKY130_FD_SC_HS__OR4_4%D
x_PM_SKY130_FD_SC_HS__OR4_4%VPWR N_VPWR_M1010_d N_VPWR_M1011_d N_VPWR_M1016_d
+ N_VPWR_M1000_d N_VPWR_c_527_n N_VPWR_c_528_n N_VPWR_c_529_n N_VPWR_c_530_n
+ N_VPWR_c_531_n VPWR N_VPWR_c_532_n N_VPWR_c_533_n N_VPWR_c_534_n
+ N_VPWR_c_535_n N_VPWR_c_526_n N_VPWR_c_537_n N_VPWR_c_538_n N_VPWR_c_539_n
+ PM_SKY130_FD_SC_HS__OR4_4%VPWR
x_PM_SKY130_FD_SC_HS__OR4_4%X N_X_M1002_s N_X_M1006_s N_X_M1010_s N_X_M1012_s
+ N_X_c_612_n N_X_c_613_n N_X_c_617_n N_X_c_614_n N_X_c_618_n N_X_c_615_n X X X
+ X N_X_c_621_n PM_SKY130_FD_SC_HS__OR4_4%X
x_PM_SKY130_FD_SC_HS__OR4_4%A_499_392# N_A_499_392#_M1009_d N_A_499_392#_M1019_d
+ N_A_499_392#_M1018_s N_A_499_392#_c_681_n N_A_499_392#_c_682_n
+ N_A_499_392#_c_699_n N_A_499_392#_c_683_n N_A_499_392#_c_690_n
+ N_A_499_392#_c_684_n N_A_499_392#_c_691_n N_A_499_392#_c_721_n
+ N_A_499_392#_c_685_n PM_SKY130_FD_SC_HS__OR4_4%A_499_392#
x_PM_SKY130_FD_SC_HS__OR4_4%A_588_392# N_A_588_392#_M1009_s N_A_588_392#_M1001_s
+ N_A_588_392#_c_752_n N_A_588_392#_c_750_n N_A_588_392#_c_756_n
+ N_A_588_392#_c_754_n N_A_588_392#_c_751_n PM_SKY130_FD_SC_HS__OR4_4%A_588_392#
x_PM_SKY130_FD_SC_HS__OR4_4%A_962_392# N_A_962_392#_M1008_d N_A_962_392#_M1017_s
+ N_A_962_392#_c_778_n PM_SKY130_FD_SC_HS__OR4_4%A_962_392#
x_PM_SKY130_FD_SC_HS__OR4_4%VGND N_VGND_M1002_d N_VGND_M1004_d N_VGND_M1007_d
+ N_VGND_M1013_d N_VGND_M1005_d N_VGND_c_792_n N_VGND_c_793_n N_VGND_c_794_n
+ N_VGND_c_795_n VGND N_VGND_c_796_n N_VGND_c_797_n N_VGND_c_798_n
+ N_VGND_c_799_n N_VGND_c_800_n N_VGND_c_801_n N_VGND_c_802_n N_VGND_c_803_n
+ N_VGND_c_804_n N_VGND_c_805_n PM_SKY130_FD_SC_HS__OR4_4%VGND
cc_1 VNB N_A_83_264#_M1002_g 0.0272031f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=0.74
cc_2 VNB N_A_83_264#_M1004_g 0.0219865f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=0.74
cc_3 VNB N_A_83_264#_M1006_g 0.0256793f $X=-0.19 $Y=-0.245 $X2=1.495 $Y2=0.74
cc_4 VNB N_A_83_264#_M1007_g 0.0265883f $X=-0.19 $Y=-0.245 $X2=2.25 $Y2=0.74
cc_5 VNB N_A_83_264#_c_112_n 6.71782e-19 $X=-0.19 $Y=-0.245 $X2=2.155 $Y2=1.485
cc_6 VNB N_A_83_264#_c_113_n 0.008967f $X=-0.19 $Y=-0.245 $X2=2.24 $Y2=1.32
cc_7 VNB N_A_83_264#_c_114_n 0.00239713f $X=-0.19 $Y=-0.245 $X2=3.085 $Y2=0.515
cc_8 VNB N_A_83_264#_c_115_n 0.00280366f $X=-0.19 $Y=-0.245 $X2=4.935 $Y2=0.515
cc_9 VNB N_A_83_264#_c_116_n 0.0283703f $X=-0.19 $Y=-0.245 $X2=6.465 $Y2=1.11
cc_10 VNB N_A_83_264#_c_117_n 0.0231448f $X=-0.19 $Y=-0.245 $X2=6.55 $Y2=1.95
cc_11 VNB N_A_83_264#_c_118_n 0.12905f $X=-0.19 $Y=-0.245 $X2=2.16 $Y2=1.485
cc_12 VNB N_A_83_264#_c_119_n 0.00258271f $X=-0.19 $Y=-0.245 $X2=4.935 $Y2=0.875
cc_13 VNB N_B_c_267_n 0.0361519f $X=-0.19 $Y=-0.245 $X2=2.945 $Y2=0.37
cc_14 VNB N_B_c_268_n 0.00142475f $X=-0.19 $Y=-0.245 $X2=4.795 $Y2=0.37
cc_15 VNB N_B_c_269_n 0.0182315f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_B_c_270_n 0.00629716f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.765
cc_17 VNB N_B_c_271_n 0.0154954f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=0.74
cc_18 VNB N_B_c_272_n 0.0151427f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=0.74
cc_19 VNB N_B_c_273_n 0.0060756f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_B_c_274_n 0.0397097f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=1.32
cc_21 VNB N_A_M1013_g 0.0336515f $X=-0.19 $Y=-0.245 $X2=5.31 $Y2=1.96
cc_22 VNB A 0.00304223f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_23 VNB N_A_c_356_n 0.0327983f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_C_M1015_g 0.0306063f $X=-0.19 $Y=-0.245 $X2=5.31 $Y2=1.96
cc_25 VNB N_C_c_403_n 0.017674f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_C_c_404_n 0.0286116f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_C_c_405_n 0.00148209f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=0.74
cc_28 VNB N_C_c_406_n 0.00637831f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_D_c_466_n 0.0169511f $X=-0.19 $Y=-0.245 $X2=2.945 $Y2=0.37
cc_30 VNB N_D_c_467_n 0.00733563f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_D_c_468_n 0.00733563f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.765
cc_32 VNB N_D_c_469_n 0.0176918f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=0.74
cc_33 VNB N_D_c_470_n 0.054246f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_D_c_471_n 0.00909013f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=1.765
cc_35 VNB N_D_c_472_n 0.0403232f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=0.74
cc_36 VNB N_D_c_473_n 0.0691165f $X=-0.19 $Y=-0.245 $X2=1.495 $Y2=0.74
cc_37 VNB N_D_c_474_n 0.00238263f $X=-0.19 $Y=-0.245 $X2=1.495 $Y2=0.74
cc_38 VNB N_VPWR_c_526_n 0.283096f $X=-0.19 $Y=-0.245 $X2=3.25 $Y2=0.875
cc_39 VNB N_X_c_612_n 0.00240191f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=0.74
cc_40 VNB N_X_c_613_n 0.0209897f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=1.765
cc_41 VNB N_X_c_614_n 0.00674496f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=0.74
cc_42 VNB N_X_c_615_n 0.0033365f $X=-0.19 $Y=-0.245 $X2=1.495 $Y2=0.74
cc_43 VNB N_VGND_c_792_n 0.0122168f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_793_n 0.0449905f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=2.4
cc_45 VNB N_VGND_c_794_n 0.00571618f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=0.74
cc_46 VNB N_VGND_c_795_n 0.00950637f $X=-0.19 $Y=-0.245 $X2=1.405 $Y2=2.4
cc_47 VNB N_VGND_c_796_n 0.0186948f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_VGND_c_797_n 0.0269696f $X=-0.19 $Y=-0.245 $X2=2.25 $Y2=0.74
cc_49 VNB N_VGND_c_798_n 0.018096f $X=-0.19 $Y=-0.245 $X2=3.25 $Y2=0.875
cc_50 VNB N_VGND_c_799_n 0.362172f $X=-0.19 $Y=-0.245 $X2=4.935 $Y2=0.79
cc_51 VNB N_VGND_c_800_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=6.465 $Y2=2.035
cc_52 VNB N_VGND_c_801_n 0.00689995f $X=-0.19 $Y=-0.245 $X2=6.55 $Y2=1.95
cc_53 VNB N_VGND_c_802_n 0.0193312f $X=-0.19 $Y=-0.245 $X2=3.085 $Y2=0.875
cc_54 VNB N_VGND_c_803_n 0.0378507f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=1.542
cc_55 VNB N_VGND_c_804_n 0.0176133f $X=-0.19 $Y=-0.245 $X2=1.405 $Y2=1.542
cc_56 VNB N_VGND_c_805_n 0.0344666f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VPB N_A_83_264#_c_120_n 0.0173785f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.765
cc_58 VPB N_A_83_264#_c_121_n 0.0146723f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=1.765
cc_59 VPB N_A_83_264#_c_122_n 0.0149018f $X=-0.19 $Y=1.66 $X2=1.405 $Y2=1.765
cc_60 VPB N_A_83_264#_c_123_n 0.0186231f $X=-0.19 $Y=1.66 $X2=1.855 $Y2=1.765
cc_61 VPB N_A_83_264#_c_124_n 0.018368f $X=-0.19 $Y=1.66 $X2=6.465 $Y2=2.035
cc_62 VPB N_A_83_264#_c_117_n 0.0141625f $X=-0.19 $Y=1.66 $X2=6.55 $Y2=1.95
cc_63 VPB N_A_83_264#_c_118_n 0.0290242f $X=-0.19 $Y=1.66 $X2=2.16 $Y2=1.485
cc_64 VPB N_A_83_264#_c_127_n 0.00247553f $X=-0.19 $Y=1.66 $X2=5.625 $Y2=2.07
cc_65 VPB N_B_c_268_n 0.0115109f $X=-0.19 $Y=1.66 $X2=4.795 $Y2=0.37
cc_66 VPB N_B_c_276_n 0.0252174f $X=-0.19 $Y=1.66 $X2=5.31 $Y2=1.96
cc_67 VPB N_B_c_270_n 0.00778116f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.765
cc_68 VPB N_B_c_278_n 0.0228675f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.4
cc_69 VPB N_A_c_357_n 0.0154387f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_70 VPB N_A_c_358_n 0.0155883f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_71 VPB A 0.002495f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.4
cc_72 VPB N_A_c_356_n 0.0335137f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_73 VPB N_C_c_403_n 0.0354219f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_74 VPB N_C_c_404_n 0.0386564f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_75 VPB N_C_c_405_n 0.0043287f $X=-0.19 $Y=1.66 $X2=0.995 $Y2=0.74
cc_76 VPB N_C_c_406_n 0.0070921f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_77 VPB N_D_c_467_n 0.00590321f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_78 VPB N_D_c_476_n 0.0221638f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_79 VPB N_D_c_468_n 0.00582344f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.765
cc_80 VPB N_D_c_478_n 0.0214349f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.4
cc_81 VPB N_VPWR_c_527_n 0.0120106f $X=-0.19 $Y=1.66 $X2=0.565 $Y2=1.32
cc_82 VPB N_VPWR_c_528_n 0.0341837f $X=-0.19 $Y=1.66 $X2=0.565 $Y2=0.74
cc_83 VPB N_VPWR_c_529_n 0.00261791f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=2.4
cc_84 VPB N_VPWR_c_530_n 0.0122845f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_85 VPB N_VPWR_c_531_n 0.00396467f $X=-0.19 $Y=1.66 $X2=1.495 $Y2=1.32
cc_86 VPB N_VPWR_c_532_n 0.0159778f $X=-0.19 $Y=1.66 $X2=1.855 $Y2=1.765
cc_87 VPB N_VPWR_c_533_n 0.0159778f $X=-0.19 $Y=1.66 $X2=2.25 $Y2=0.74
cc_88 VPB N_VPWR_c_534_n 0.0313938f $X=-0.19 $Y=1.66 $X2=1.48 $Y2=1.485
cc_89 VPB N_VPWR_c_535_n 0.0810424f $X=-0.19 $Y=1.66 $X2=4.77 $Y2=0.875
cc_90 VPB N_VPWR_c_526_n 0.0881624f $X=-0.19 $Y=1.66 $X2=3.25 $Y2=0.875
cc_91 VPB N_VPWR_c_537_n 0.00601644f $X=-0.19 $Y=1.66 $X2=5.1 $Y2=1.11
cc_92 VPB N_VPWR_c_538_n 0.00614127f $X=-0.19 $Y=1.66 $X2=6.55 $Y2=1.195
cc_93 VPB N_VPWR_c_539_n 0.00601668f $X=-0.19 $Y=1.66 $X2=2.16 $Y2=1.485
cc_94 VPB N_X_c_613_n 0.0208972f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=1.765
cc_95 VPB N_X_c_617_n 0.00233217f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=2.4
cc_96 VPB N_X_c_618_n 0.00233217f $X=-0.19 $Y=1.66 $X2=1.405 $Y2=2.4
cc_97 VPB X 0.00141215f $X=-0.19 $Y=1.66 $X2=2.25 $Y2=1.32
cc_98 VPB X 0.00770046f $X=-0.19 $Y=1.66 $X2=2.25 $Y2=0.74
cc_99 VPB N_X_c_621_n 0.00400014f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_100 VPB N_A_499_392#_c_681_n 0.00752808f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.765
cc_101 VPB N_A_499_392#_c_682_n 0.0104513f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.4
cc_102 VPB N_A_499_392#_c_683_n 0.0095708f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_103 VPB N_A_499_392#_c_684_n 0.00289722f $X=-0.19 $Y=1.66 $X2=0.995 $Y2=1.32
cc_104 VPB N_A_499_392#_c_685_n 0.03008f $X=-0.19 $Y=1.66 $X2=1.855 $Y2=2.4
cc_105 VPB N_A_588_392#_c_750_n 0.00242717f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_106 VPB N_A_588_392#_c_751_n 0.00244088f $X=-0.19 $Y=1.66 $X2=0.565 $Y2=0.74
cc_107 VPB N_A_962_392#_c_778_n 0.00792862f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.4
cc_108 N_A_83_264#_M1007_g N_B_c_267_n 0.0139171f $X=2.25 $Y=0.74 $X2=-0.19
+ $Y2=-0.245
cc_109 N_A_83_264#_c_113_n N_B_c_267_n 9.47471e-19 $X=2.24 $Y=1.32 $X2=-0.19
+ $Y2=-0.245
cc_110 N_A_83_264#_c_130_p N_B_c_267_n 8.97023e-19 $X=2.92 $Y=0.875 $X2=-0.19
+ $Y2=-0.245
cc_111 N_A_83_264#_c_118_n N_B_c_267_n 0.00225496f $X=2.16 $Y=1.485 $X2=-0.19
+ $Y2=-0.245
cc_112 N_A_83_264#_M1007_g N_B_c_269_n 0.0204288f $X=2.25 $Y=0.74 $X2=0 $Y2=0
cc_113 N_A_83_264#_c_113_n N_B_c_269_n 0.00101364f $X=2.24 $Y=1.32 $X2=0 $Y2=0
cc_114 N_A_83_264#_c_130_p N_B_c_269_n 0.0092233f $X=2.92 $Y=0.875 $X2=0 $Y2=0
cc_115 N_A_83_264#_c_114_n N_B_c_269_n 0.00689388f $X=3.085 $Y=0.515 $X2=0 $Y2=0
cc_116 N_A_83_264#_c_136_p N_B_c_269_n 7.15033e-19 $X=3.085 $Y=0.875 $X2=0 $Y2=0
cc_117 N_A_83_264#_c_137_p N_B_c_271_n 0.0574059f $X=4.77 $Y=0.875 $X2=0 $Y2=0
cc_118 N_A_83_264#_c_136_p N_B_c_271_n 0.00109891f $X=3.085 $Y=0.875 $X2=0 $Y2=0
cc_119 N_A_83_264#_M1007_g N_B_c_272_n 0.00140149f $X=2.25 $Y=0.74 $X2=0 $Y2=0
cc_120 N_A_83_264#_c_113_n N_B_c_272_n 0.0283182f $X=2.24 $Y=1.32 $X2=0 $Y2=0
cc_121 N_A_83_264#_c_130_p N_B_c_272_n 0.02837f $X=2.92 $Y=0.875 $X2=0 $Y2=0
cc_122 N_A_83_264#_c_118_n N_B_c_272_n 5.52866e-19 $X=2.16 $Y=1.485 $X2=0 $Y2=0
cc_123 N_A_83_264#_c_136_p N_B_c_272_n 0.0223159f $X=3.085 $Y=0.875 $X2=0 $Y2=0
cc_124 N_A_83_264#_c_137_p N_B_c_273_n 0.0261968f $X=4.77 $Y=0.875 $X2=0 $Y2=0
cc_125 N_A_83_264#_c_119_n N_B_c_273_n 0.00285444f $X=4.935 $Y=0.875 $X2=0 $Y2=0
cc_126 N_A_83_264#_c_137_p N_B_c_274_n 0.00181437f $X=4.77 $Y=0.875 $X2=0 $Y2=0
cc_127 N_A_83_264#_c_114_n N_A_M1013_g 0.010756f $X=3.085 $Y=0.515 $X2=0 $Y2=0
cc_128 N_A_83_264#_c_137_p N_A_M1013_g 0.0104279f $X=4.77 $Y=0.875 $X2=0 $Y2=0
cc_129 N_A_83_264#_c_136_p N_A_M1013_g 7.15645e-19 $X=3.085 $Y=0.875 $X2=0 $Y2=0
cc_130 N_A_83_264#_c_137_p N_C_M1015_g 0.0120241f $X=4.77 $Y=0.875 $X2=0 $Y2=0
cc_131 N_A_83_264#_c_115_n N_C_M1015_g 0.0114883f $X=4.935 $Y=0.515 $X2=0 $Y2=0
cc_132 N_A_83_264#_c_119_n N_C_M1015_g 0.0106918f $X=4.935 $Y=0.875 $X2=0 $Y2=0
cc_133 N_A_83_264#_c_119_n N_C_c_403_n 9.10599e-19 $X=4.935 $Y=0.875 $X2=0 $Y2=0
cc_134 N_A_83_264#_c_127_n N_C_c_403_n 7.2065e-19 $X=5.625 $Y=2.07 $X2=0 $Y2=0
cc_135 N_A_83_264#_c_116_n N_C_c_404_n 0.0033708f $X=6.465 $Y=1.11 $X2=0 $Y2=0
cc_136 N_A_83_264#_c_124_n N_C_c_404_n 0.0174437f $X=6.465 $Y=2.035 $X2=0 $Y2=0
cc_137 N_A_83_264#_c_117_n N_C_c_404_n 0.0150067f $X=6.55 $Y=1.95 $X2=0 $Y2=0
cc_138 N_A_83_264#_c_127_n N_C_c_404_n 3.28132e-19 $X=5.625 $Y=2.07 $X2=0 $Y2=0
cc_139 N_A_83_264#_c_116_n N_C_c_405_n 0.0715147f $X=6.465 $Y=1.11 $X2=0 $Y2=0
cc_140 N_A_83_264#_c_117_n N_C_c_405_n 0.0315994f $X=6.55 $Y=1.95 $X2=0 $Y2=0
cc_141 N_A_83_264#_c_127_n N_C_c_405_n 0.0736416f $X=5.625 $Y=2.07 $X2=0 $Y2=0
cc_142 N_A_83_264#_c_137_p N_C_c_406_n 0.00546445f $X=4.77 $Y=0.875 $X2=0 $Y2=0
cc_143 N_A_83_264#_c_116_n N_C_c_406_n 0.01791f $X=6.465 $Y=1.11 $X2=0 $Y2=0
cc_144 N_A_83_264#_c_119_n N_C_c_406_n 0.0293972f $X=4.935 $Y=0.875 $X2=0 $Y2=0
cc_145 N_A_83_264#_c_127_n N_C_c_406_n 0.00355534f $X=5.625 $Y=2.07 $X2=0 $Y2=0
cc_146 N_A_83_264#_c_115_n N_D_c_466_n 0.00358648f $X=4.935 $Y=0.515 $X2=-0.19
+ $Y2=-0.245
cc_147 N_A_83_264#_c_116_n N_D_c_466_n 0.0113592f $X=6.465 $Y=1.11 $X2=-0.19
+ $Y2=-0.245
cc_148 N_A_83_264#_c_119_n N_D_c_466_n 4.42511e-19 $X=4.935 $Y=0.875 $X2=-0.19
+ $Y2=-0.245
cc_149 N_A_83_264#_c_127_n N_D_c_476_n 0.00538238f $X=5.625 $Y=2.07 $X2=0 $Y2=0
cc_150 N_A_83_264#_c_124_n N_D_c_478_n 0.00868026f $X=6.465 $Y=2.035 $X2=0 $Y2=0
cc_151 N_A_83_264#_c_127_n N_D_c_478_n 0.00241381f $X=5.625 $Y=2.07 $X2=0 $Y2=0
cc_152 N_A_83_264#_c_116_n N_D_c_469_n 0.0105003f $X=6.465 $Y=1.11 $X2=0 $Y2=0
cc_153 N_A_83_264#_c_116_n N_D_c_470_n 0.0192499f $X=6.465 $Y=1.11 $X2=0 $Y2=0
cc_154 N_A_83_264#_c_116_n N_D_c_472_n 0.0120613f $X=6.465 $Y=1.11 $X2=0 $Y2=0
cc_155 N_A_83_264#_c_117_n N_D_c_472_n 0.00405285f $X=6.55 $Y=1.95 $X2=0 $Y2=0
cc_156 N_A_83_264#_c_127_n N_D_c_472_n 3.42297e-19 $X=5.625 $Y=2.07 $X2=0 $Y2=0
cc_157 N_A_83_264#_c_116_n N_D_c_474_n 0.0272875f $X=6.465 $Y=1.11 $X2=0 $Y2=0
cc_158 N_A_83_264#_c_120_n N_VPWR_c_528_n 0.0116616f $X=0.505 $Y=1.765 $X2=0
+ $Y2=0
cc_159 N_A_83_264#_c_121_n N_VPWR_c_528_n 4.98648e-19 $X=0.955 $Y=1.765 $X2=0
+ $Y2=0
cc_160 N_A_83_264#_c_120_n N_VPWR_c_529_n 4.98648e-19 $X=0.505 $Y=1.765 $X2=0
+ $Y2=0
cc_161 N_A_83_264#_c_121_n N_VPWR_c_529_n 0.0105176f $X=0.955 $Y=1.765 $X2=0
+ $Y2=0
cc_162 N_A_83_264#_c_122_n N_VPWR_c_529_n 0.0105176f $X=1.405 $Y=1.765 $X2=0
+ $Y2=0
cc_163 N_A_83_264#_c_123_n N_VPWR_c_529_n 4.98648e-19 $X=1.855 $Y=1.765 $X2=0
+ $Y2=0
cc_164 N_A_83_264#_c_122_n N_VPWR_c_530_n 4.98648e-19 $X=1.405 $Y=1.765 $X2=0
+ $Y2=0
cc_165 N_A_83_264#_c_123_n N_VPWR_c_530_n 0.0116621f $X=1.855 $Y=1.765 $X2=0
+ $Y2=0
cc_166 N_A_83_264#_c_120_n N_VPWR_c_532_n 0.00413917f $X=0.505 $Y=1.765 $X2=0
+ $Y2=0
cc_167 N_A_83_264#_c_121_n N_VPWR_c_532_n 0.00413917f $X=0.955 $Y=1.765 $X2=0
+ $Y2=0
cc_168 N_A_83_264#_c_122_n N_VPWR_c_533_n 0.00413917f $X=1.405 $Y=1.765 $X2=0
+ $Y2=0
cc_169 N_A_83_264#_c_123_n N_VPWR_c_533_n 0.00413917f $X=1.855 $Y=1.765 $X2=0
+ $Y2=0
cc_170 N_A_83_264#_c_120_n N_VPWR_c_526_n 0.00817726f $X=0.505 $Y=1.765 $X2=0
+ $Y2=0
cc_171 N_A_83_264#_c_121_n N_VPWR_c_526_n 0.00817726f $X=0.955 $Y=1.765 $X2=0
+ $Y2=0
cc_172 N_A_83_264#_c_122_n N_VPWR_c_526_n 0.00817726f $X=1.405 $Y=1.765 $X2=0
+ $Y2=0
cc_173 N_A_83_264#_c_123_n N_VPWR_c_526_n 0.00817726f $X=1.855 $Y=1.765 $X2=0
+ $Y2=0
cc_174 N_A_83_264#_M1002_g N_X_c_612_n 0.00788812f $X=0.565 $Y=0.74 $X2=0 $Y2=0
cc_175 N_A_83_264#_M1004_g N_X_c_612_n 0.00926373f $X=0.995 $Y=0.74 $X2=0 $Y2=0
cc_176 N_A_83_264#_M1006_g N_X_c_612_n 6.73969e-19 $X=1.495 $Y=0.74 $X2=0 $Y2=0
cc_177 N_A_83_264#_c_120_n N_X_c_613_n 0.0212877f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_178 N_A_83_264#_M1002_g N_X_c_613_n 0.0189011f $X=0.565 $Y=0.74 $X2=0 $Y2=0
cc_179 N_A_83_264#_c_121_n N_X_c_613_n 0.0066527f $X=0.955 $Y=1.765 $X2=0 $Y2=0
cc_180 N_A_83_264#_M1004_g N_X_c_613_n 0.00535402f $X=0.995 $Y=0.74 $X2=0 $Y2=0
cc_181 N_A_83_264#_M1006_g N_X_c_613_n 5.67152e-19 $X=1.495 $Y=0.74 $X2=0 $Y2=0
cc_182 N_A_83_264#_c_112_n N_X_c_613_n 0.0147894f $X=2.155 $Y=1.485 $X2=0 $Y2=0
cc_183 N_A_83_264#_c_118_n N_X_c_613_n 0.0464636f $X=2.16 $Y=1.485 $X2=0 $Y2=0
cc_184 N_A_83_264#_c_120_n N_X_c_617_n 3.85296e-19 $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_185 N_A_83_264#_c_121_n N_X_c_617_n 3.85296e-19 $X=0.955 $Y=1.765 $X2=0 $Y2=0
cc_186 N_A_83_264#_M1004_g N_X_c_614_n 0.0133465f $X=0.995 $Y=0.74 $X2=0 $Y2=0
cc_187 N_A_83_264#_M1006_g N_X_c_614_n 0.0155759f $X=1.495 $Y=0.74 $X2=0 $Y2=0
cc_188 N_A_83_264#_M1007_g N_X_c_614_n 8.15014e-19 $X=2.25 $Y=0.74 $X2=0 $Y2=0
cc_189 N_A_83_264#_c_112_n N_X_c_614_n 0.0497808f $X=2.155 $Y=1.485 $X2=0 $Y2=0
cc_190 N_A_83_264#_c_113_n N_X_c_614_n 0.00786297f $X=2.24 $Y=1.32 $X2=0 $Y2=0
cc_191 N_A_83_264#_c_118_n N_X_c_614_n 0.0121439f $X=2.16 $Y=1.485 $X2=0 $Y2=0
cc_192 N_A_83_264#_c_122_n N_X_c_618_n 3.85296e-19 $X=1.405 $Y=1.765 $X2=0 $Y2=0
cc_193 N_A_83_264#_c_123_n N_X_c_618_n 3.85296e-19 $X=1.855 $Y=1.765 $X2=0 $Y2=0
cc_194 N_A_83_264#_M1006_g N_X_c_615_n 0.00516826f $X=1.495 $Y=0.74 $X2=0 $Y2=0
cc_195 N_A_83_264#_M1007_g N_X_c_615_n 0.00796805f $X=2.25 $Y=0.74 $X2=0 $Y2=0
cc_196 N_A_83_264#_c_112_n X 0.0193967f $X=2.155 $Y=1.485 $X2=0 $Y2=0
cc_197 N_A_83_264#_c_118_n X 0.00592991f $X=2.16 $Y=1.485 $X2=0 $Y2=0
cc_198 N_A_83_264#_c_123_n X 0.0204061f $X=1.855 $Y=1.765 $X2=0 $Y2=0
cc_199 N_A_83_264#_c_112_n X 0.0317535f $X=2.155 $Y=1.485 $X2=0 $Y2=0
cc_200 N_A_83_264#_c_113_n X 0.0100698f $X=2.24 $Y=1.32 $X2=0 $Y2=0
cc_201 N_A_83_264#_c_118_n X 0.00722452f $X=2.16 $Y=1.485 $X2=0 $Y2=0
cc_202 N_A_83_264#_c_121_n N_X_c_621_n 0.0126739f $X=0.955 $Y=1.765 $X2=0 $Y2=0
cc_203 N_A_83_264#_c_122_n N_X_c_621_n 0.0177404f $X=1.405 $Y=1.765 $X2=0 $Y2=0
cc_204 N_A_83_264#_c_112_n N_X_c_621_n 0.0151717f $X=2.155 $Y=1.485 $X2=0 $Y2=0
cc_205 N_A_83_264#_c_118_n N_X_c_621_n 0.00430664f $X=2.16 $Y=1.485 $X2=0 $Y2=0
cc_206 N_A_83_264#_c_124_n N_A_499_392#_M1018_s 0.00453841f $X=6.465 $Y=2.035
+ $X2=0 $Y2=0
cc_207 N_A_83_264#_c_123_n N_A_499_392#_c_681_n 0.00184119f $X=1.855 $Y=1.765
+ $X2=0 $Y2=0
cc_208 N_A_83_264#_c_123_n N_A_499_392#_c_682_n 0.00309581f $X=1.855 $Y=1.765
+ $X2=0 $Y2=0
cc_209 N_A_83_264#_c_127_n N_A_499_392#_c_683_n 0.0053729f $X=5.625 $Y=2.07
+ $X2=0 $Y2=0
cc_210 N_A_83_264#_c_127_n N_A_499_392#_c_690_n 0.00124609f $X=5.625 $Y=2.07
+ $X2=0 $Y2=0
cc_211 N_A_83_264#_M1014_d N_A_499_392#_c_691_n 0.00393062f $X=5.31 $Y=1.96
+ $X2=0 $Y2=0
cc_212 N_A_83_264#_c_124_n N_A_499_392#_c_691_n 0.0251151f $X=6.465 $Y=2.035
+ $X2=0 $Y2=0
cc_213 N_A_83_264#_c_127_n N_A_499_392#_c_691_n 0.0158852f $X=5.625 $Y=2.07
+ $X2=0 $Y2=0
cc_214 N_A_83_264#_c_124_n N_A_499_392#_c_685_n 0.026091f $X=6.465 $Y=2.035
+ $X2=0 $Y2=0
cc_215 N_A_83_264#_c_124_n N_A_962_392#_M1017_s 0.00230902f $X=6.465 $Y=2.035
+ $X2=0 $Y2=0
cc_216 N_A_83_264#_M1014_d N_A_962_392#_c_778_n 0.00201274f $X=5.31 $Y=1.96
+ $X2=0 $Y2=0
cc_217 N_A_83_264#_c_130_p N_VGND_M1007_d 0.0122153f $X=2.92 $Y=0.875 $X2=0
+ $Y2=0
cc_218 N_A_83_264#_c_137_p N_VGND_M1013_d 0.0370525f $X=4.77 $Y=0.875 $X2=0
+ $Y2=0
cc_219 N_A_83_264#_c_116_n N_VGND_M1005_d 0.00286681f $X=6.465 $Y=1.11 $X2=0
+ $Y2=0
cc_220 N_A_83_264#_M1002_g N_VGND_c_793_n 0.0184904f $X=0.565 $Y=0.74 $X2=0
+ $Y2=0
cc_221 N_A_83_264#_c_118_n N_VGND_c_793_n 2.15299e-19 $X=2.16 $Y=1.485 $X2=0
+ $Y2=0
cc_222 N_A_83_264#_M1004_g N_VGND_c_794_n 0.00417204f $X=0.995 $Y=0.74 $X2=0
+ $Y2=0
cc_223 N_A_83_264#_M1006_g N_VGND_c_794_n 0.0125758f $X=1.495 $Y=0.74 $X2=0
+ $Y2=0
cc_224 N_A_83_264#_M1007_g N_VGND_c_795_n 0.00516167f $X=2.25 $Y=0.74 $X2=0
+ $Y2=0
cc_225 N_A_83_264#_c_130_p N_VGND_c_795_n 0.0282828f $X=2.92 $Y=0.875 $X2=0
+ $Y2=0
cc_226 N_A_83_264#_c_114_n N_VGND_c_795_n 0.0104464f $X=3.085 $Y=0.515 $X2=0
+ $Y2=0
cc_227 N_A_83_264#_M1002_g N_VGND_c_796_n 0.00434272f $X=0.565 $Y=0.74 $X2=0
+ $Y2=0
cc_228 N_A_83_264#_M1004_g N_VGND_c_796_n 0.00434272f $X=0.995 $Y=0.74 $X2=0
+ $Y2=0
cc_229 N_A_83_264#_M1006_g N_VGND_c_797_n 0.00383152f $X=1.495 $Y=0.74 $X2=0
+ $Y2=0
cc_230 N_A_83_264#_M1007_g N_VGND_c_797_n 0.00461464f $X=2.25 $Y=0.74 $X2=0
+ $Y2=0
cc_231 N_A_83_264#_M1002_g N_VGND_c_799_n 0.00823934f $X=0.565 $Y=0.74 $X2=0
+ $Y2=0
cc_232 N_A_83_264#_M1004_g N_VGND_c_799_n 0.00820718f $X=0.995 $Y=0.74 $X2=0
+ $Y2=0
cc_233 N_A_83_264#_M1006_g N_VGND_c_799_n 0.00759969f $X=1.495 $Y=0.74 $X2=0
+ $Y2=0
cc_234 N_A_83_264#_M1007_g N_VGND_c_799_n 0.0045489f $X=2.25 $Y=0.74 $X2=0 $Y2=0
cc_235 N_A_83_264#_c_130_p N_VGND_c_799_n 0.00886098f $X=2.92 $Y=0.875 $X2=0
+ $Y2=0
cc_236 N_A_83_264#_c_256_p N_VGND_c_799_n 0.00583874f $X=2.325 $Y=0.875 $X2=0
+ $Y2=0
cc_237 N_A_83_264#_c_114_n N_VGND_c_799_n 0.0118382f $X=3.085 $Y=0.515 $X2=0
+ $Y2=0
cc_238 N_A_83_264#_c_137_p N_VGND_c_799_n 0.0151942f $X=4.77 $Y=0.875 $X2=0
+ $Y2=0
cc_239 N_A_83_264#_c_115_n N_VGND_c_799_n 0.0119984f $X=4.935 $Y=0.515 $X2=0
+ $Y2=0
cc_240 N_A_83_264#_c_114_n N_VGND_c_802_n 0.014379f $X=3.085 $Y=0.515 $X2=0
+ $Y2=0
cc_241 N_A_83_264#_c_114_n N_VGND_c_803_n 0.010535f $X=3.085 $Y=0.515 $X2=0
+ $Y2=0
cc_242 N_A_83_264#_c_137_p N_VGND_c_803_n 0.091374f $X=4.77 $Y=0.875 $X2=0 $Y2=0
cc_243 N_A_83_264#_c_115_n N_VGND_c_803_n 0.010535f $X=4.935 $Y=0.515 $X2=0
+ $Y2=0
cc_244 N_A_83_264#_c_115_n N_VGND_c_804_n 0.0145639f $X=4.935 $Y=0.515 $X2=0
+ $Y2=0
cc_245 N_A_83_264#_c_115_n N_VGND_c_805_n 0.0146527f $X=4.935 $Y=0.515 $X2=0
+ $Y2=0
cc_246 N_A_83_264#_c_116_n N_VGND_c_805_n 0.0390715f $X=6.465 $Y=1.11 $X2=0
+ $Y2=0
cc_247 N_B_c_269_n N_A_M1013_g 0.013775f $X=2.87 $Y=1.22 $X2=0 $Y2=0
cc_248 N_B_c_271_n N_A_M1013_g 0.0117361f $X=4.065 $Y=1.215 $X2=0 $Y2=0
cc_249 N_B_c_272_n N_A_M1013_g 0.0120208f $X=3.235 $Y=1.215 $X2=0 $Y2=0
cc_250 N_B_c_273_n N_A_M1013_g 9.8879e-19 $X=4.23 $Y=1.215 $X2=0 $Y2=0
cc_251 N_B_c_274_n N_A_M1013_g 0.0040104f $X=4.23 $Y=1.385 $X2=0 $Y2=0
cc_252 N_B_c_276_n N_A_c_357_n 0.0216649f $X=2.865 $Y=1.885 $X2=0 $Y2=0
cc_253 N_B_c_278_n N_A_c_358_n 0.0185807f $X=4.235 $Y=1.885 $X2=0 $Y2=0
cc_254 N_B_c_267_n A 0.00117317f $X=2.865 $Y=1.64 $X2=0 $Y2=0
cc_255 N_B_c_270_n A 0.00124404f $X=4.235 $Y=1.795 $X2=0 $Y2=0
cc_256 N_B_c_271_n A 0.0247729f $X=4.065 $Y=1.215 $X2=0 $Y2=0
cc_257 N_B_c_272_n A 0.00633894f $X=3.235 $Y=1.215 $X2=0 $Y2=0
cc_258 N_B_c_273_n A 0.00352889f $X=4.23 $Y=1.215 $X2=0 $Y2=0
cc_259 N_B_c_274_n A 2.32886e-19 $X=4.23 $Y=1.385 $X2=0 $Y2=0
cc_260 N_B_c_267_n N_A_c_356_n 0.032028f $X=2.865 $Y=1.64 $X2=0 $Y2=0
cc_261 N_B_c_270_n N_A_c_356_n 0.0168757f $X=4.235 $Y=1.795 $X2=0 $Y2=0
cc_262 N_B_c_271_n N_A_c_356_n 0.00697339f $X=4.065 $Y=1.215 $X2=0 $Y2=0
cc_263 N_B_c_272_n N_A_c_356_n 0.00237378f $X=3.235 $Y=1.215 $X2=0 $Y2=0
cc_264 N_B_c_273_n N_A_c_356_n 3.40206e-19 $X=4.23 $Y=1.215 $X2=0 $Y2=0
cc_265 N_B_c_274_n N_A_c_356_n 0.00523467f $X=4.23 $Y=1.385 $X2=0 $Y2=0
cc_266 N_B_c_273_n N_C_M1015_g 0.00316947f $X=4.23 $Y=1.215 $X2=0 $Y2=0
cc_267 N_B_c_274_n N_C_M1015_g 0.0114999f $X=4.23 $Y=1.385 $X2=0 $Y2=0
cc_268 N_B_c_270_n N_C_c_403_n 0.0145288f $X=4.235 $Y=1.795 $X2=0 $Y2=0
cc_269 N_B_c_278_n N_C_c_403_n 0.0212433f $X=4.235 $Y=1.885 $X2=0 $Y2=0
cc_270 N_B_c_274_n N_C_c_403_n 0.00691933f $X=4.23 $Y=1.385 $X2=0 $Y2=0
cc_271 N_B_c_270_n N_C_c_406_n 0.00138903f $X=4.235 $Y=1.795 $X2=0 $Y2=0
cc_272 N_B_c_273_n N_C_c_406_n 0.012807f $X=4.23 $Y=1.215 $X2=0 $Y2=0
cc_273 N_B_c_274_n N_C_c_406_n 8.90064e-19 $X=4.23 $Y=1.385 $X2=0 $Y2=0
cc_274 N_B_c_276_n N_VPWR_c_530_n 0.00383295f $X=2.865 $Y=1.885 $X2=0 $Y2=0
cc_275 N_B_c_276_n N_VPWR_c_531_n 6.09546e-19 $X=2.865 $Y=1.885 $X2=0 $Y2=0
cc_276 N_B_c_278_n N_VPWR_c_531_n 6.07905e-19 $X=4.235 $Y=1.885 $X2=0 $Y2=0
cc_277 N_B_c_276_n N_VPWR_c_534_n 0.00445602f $X=2.865 $Y=1.885 $X2=0 $Y2=0
cc_278 N_B_c_278_n N_VPWR_c_535_n 0.00445602f $X=4.235 $Y=1.885 $X2=0 $Y2=0
cc_279 N_B_c_276_n N_VPWR_c_526_n 0.00863237f $X=2.865 $Y=1.885 $X2=0 $Y2=0
cc_280 N_B_c_278_n N_VPWR_c_526_n 0.00859126f $X=4.235 $Y=1.885 $X2=0 $Y2=0
cc_281 N_B_c_276_n X 0.00389401f $X=2.865 $Y=1.885 $X2=0 $Y2=0
cc_282 N_B_c_267_n N_A_499_392#_c_681_n 0.00111452f $X=2.865 $Y=1.64 $X2=0 $Y2=0
cc_283 N_B_c_276_n N_A_499_392#_c_681_n 0.00352009f $X=2.865 $Y=1.885 $X2=0
+ $Y2=0
cc_284 N_B_c_272_n N_A_499_392#_c_681_n 0.0121282f $X=3.235 $Y=1.215 $X2=0 $Y2=0
cc_285 N_B_c_276_n N_A_499_392#_c_682_n 4.53441e-19 $X=2.865 $Y=1.885 $X2=0
+ $Y2=0
cc_286 N_B_c_276_n N_A_499_392#_c_699_n 0.0127033f $X=2.865 $Y=1.885 $X2=0 $Y2=0
cc_287 N_B_c_278_n N_A_499_392#_c_699_n 0.0164423f $X=4.235 $Y=1.885 $X2=0 $Y2=0
cc_288 N_B_c_271_n N_A_499_392#_c_699_n 0.0116178f $X=4.065 $Y=1.215 $X2=0 $Y2=0
cc_289 N_B_c_272_n N_A_499_392#_c_699_n 0.014934f $X=3.235 $Y=1.215 $X2=0 $Y2=0
cc_290 N_B_c_273_n N_A_499_392#_c_699_n 0.00839278f $X=4.23 $Y=1.215 $X2=0 $Y2=0
cc_291 N_B_c_274_n N_A_499_392#_c_699_n 3.23468e-19 $X=4.23 $Y=1.385 $X2=0 $Y2=0
cc_292 N_B_c_278_n N_A_499_392#_c_683_n 6.05832e-19 $X=4.235 $Y=1.885 $X2=0
+ $Y2=0
cc_293 N_B_c_273_n N_A_499_392#_c_683_n 0.0022688f $X=4.23 $Y=1.215 $X2=0 $Y2=0
cc_294 N_B_c_274_n N_A_499_392#_c_683_n 3.46941e-19 $X=4.23 $Y=1.385 $X2=0 $Y2=0
cc_295 N_B_c_278_n N_A_499_392#_c_684_n 0.00245875f $X=4.235 $Y=1.885 $X2=0
+ $Y2=0
cc_296 N_B_c_276_n N_A_588_392#_c_752_n 0.0022166f $X=2.865 $Y=1.885 $X2=0 $Y2=0
cc_297 N_B_c_276_n N_A_588_392#_c_750_n 0.00450948f $X=2.865 $Y=1.885 $X2=0
+ $Y2=0
cc_298 N_B_c_278_n N_A_588_392#_c_754_n 0.00257852f $X=4.235 $Y=1.885 $X2=0
+ $Y2=0
cc_299 N_B_c_278_n N_A_588_392#_c_751_n 0.00465254f $X=4.235 $Y=1.885 $X2=0
+ $Y2=0
cc_300 N_B_c_269_n N_VGND_c_795_n 0.00508528f $X=2.87 $Y=1.22 $X2=0 $Y2=0
cc_301 N_B_c_269_n N_VGND_c_799_n 0.00436349f $X=2.87 $Y=1.22 $X2=0 $Y2=0
cc_302 N_B_c_269_n N_VGND_c_802_n 0.00434272f $X=2.87 $Y=1.22 $X2=0 $Y2=0
cc_303 N_A_c_357_n N_VPWR_c_531_n 0.00645777f $X=3.315 $Y=1.885 $X2=0 $Y2=0
cc_304 N_A_c_358_n N_VPWR_c_531_n 0.00661395f $X=3.765 $Y=1.885 $X2=0 $Y2=0
cc_305 N_A_c_357_n N_VPWR_c_534_n 0.00413917f $X=3.315 $Y=1.885 $X2=0 $Y2=0
cc_306 N_A_c_358_n N_VPWR_c_535_n 0.00413917f $X=3.765 $Y=1.885 $X2=0 $Y2=0
cc_307 N_A_c_357_n N_VPWR_c_526_n 0.00398725f $X=3.315 $Y=1.885 $X2=0 $Y2=0
cc_308 N_A_c_358_n N_VPWR_c_526_n 0.00398877f $X=3.765 $Y=1.885 $X2=0 $Y2=0
cc_309 N_A_c_357_n N_A_499_392#_c_681_n 3.80443e-19 $X=3.315 $Y=1.885 $X2=0
+ $Y2=0
cc_310 N_A_c_357_n N_A_499_392#_c_699_n 0.0132145f $X=3.315 $Y=1.885 $X2=0 $Y2=0
cc_311 N_A_c_358_n N_A_499_392#_c_699_n 0.0123532f $X=3.765 $Y=1.885 $X2=0 $Y2=0
cc_312 A N_A_499_392#_c_699_n 0.0206598f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_313 N_A_c_356_n N_A_499_392#_c_699_n 0.00171521f $X=3.57 $Y=1.635 $X2=0 $Y2=0
cc_314 N_A_c_357_n N_A_588_392#_c_756_n 0.0107824f $X=3.315 $Y=1.885 $X2=0 $Y2=0
cc_315 N_A_c_358_n N_A_588_392#_c_756_n 0.00993773f $X=3.765 $Y=1.885 $X2=0
+ $Y2=0
cc_316 N_A_c_357_n N_A_588_392#_c_754_n 2.37588e-19 $X=3.315 $Y=1.885 $X2=0
+ $Y2=0
cc_317 N_A_c_358_n N_A_588_392#_c_754_n 0.00167276f $X=3.765 $Y=1.885 $X2=0
+ $Y2=0
cc_318 N_A_c_358_n N_A_588_392#_c_751_n 3.01994e-19 $X=3.765 $Y=1.885 $X2=0
+ $Y2=0
cc_319 N_A_M1013_g N_VGND_c_799_n 0.00439727f $X=3.3 $Y=0.74 $X2=0 $Y2=0
cc_320 N_A_M1013_g N_VGND_c_802_n 0.00434272f $X=3.3 $Y=0.74 $X2=0 $Y2=0
cc_321 N_A_M1013_g N_VGND_c_803_n 0.0103115f $X=3.3 $Y=0.74 $X2=0 $Y2=0
cc_322 N_C_M1015_g N_D_c_466_n 0.0280437f $X=4.72 $Y=0.74 $X2=-0.19 $Y2=-0.245
cc_323 N_C_c_403_n N_D_c_467_n 0.00517616f $X=4.735 $Y=1.885 $X2=0 $Y2=0
cc_324 N_C_c_406_n N_D_c_467_n 0.0154041f $X=5.34 $Y=1.572 $X2=0 $Y2=0
cc_325 N_C_c_403_n N_D_c_476_n 0.0351335f $X=4.735 $Y=1.885 $X2=0 $Y2=0
cc_326 N_C_c_404_n N_D_c_468_n 0.005349f $X=6.135 $Y=1.885 $X2=0 $Y2=0
cc_327 N_C_c_405_n N_D_c_468_n 0.0133602f $X=6.15 $Y=1.53 $X2=0 $Y2=0
cc_328 N_C_c_404_n N_D_c_478_n 0.0371696f $X=6.135 $Y=1.885 $X2=0 $Y2=0
cc_329 N_C_c_404_n N_D_c_470_n 0.00670431f $X=6.135 $Y=1.885 $X2=0 $Y2=0
cc_330 N_C_c_403_n N_D_c_472_n 0.0213325f $X=4.735 $Y=1.885 $X2=0 $Y2=0
cc_331 N_C_c_404_n N_D_c_472_n 0.0268774f $X=6.135 $Y=1.885 $X2=0 $Y2=0
cc_332 N_C_c_405_n N_D_c_472_n 0.0139321f $X=6.15 $Y=1.53 $X2=0 $Y2=0
cc_333 N_C_c_406_n N_D_c_472_n 0.00645108f $X=5.34 $Y=1.572 $X2=0 $Y2=0
cc_334 N_C_c_403_n N_VPWR_c_535_n 0.00445602f $X=4.735 $Y=1.885 $X2=0 $Y2=0
cc_335 N_C_c_404_n N_VPWR_c_535_n 0.00444483f $X=6.135 $Y=1.885 $X2=0 $Y2=0
cc_336 N_C_c_403_n N_VPWR_c_526_n 0.00445519f $X=4.735 $Y=1.885 $X2=0 $Y2=0
cc_337 N_C_c_404_n N_VPWR_c_526_n 0.00449262f $X=6.135 $Y=1.885 $X2=0 $Y2=0
cc_338 N_C_c_403_n N_A_499_392#_c_683_n 0.00495609f $X=4.735 $Y=1.885 $X2=0
+ $Y2=0
cc_339 N_C_c_406_n N_A_499_392#_c_683_n 0.00594841f $X=5.34 $Y=1.572 $X2=0 $Y2=0
cc_340 N_C_c_403_n N_A_499_392#_c_690_n 0.00404604f $X=4.735 $Y=1.885 $X2=0
+ $Y2=0
cc_341 N_C_c_403_n N_A_499_392#_c_684_n 0.00617104f $X=4.735 $Y=1.885 $X2=0
+ $Y2=0
cc_342 N_C_c_403_n N_A_499_392#_c_691_n 0.0114825f $X=4.735 $Y=1.885 $X2=0 $Y2=0
cc_343 N_C_c_404_n N_A_499_392#_c_691_n 0.0136513f $X=6.135 $Y=1.885 $X2=0 $Y2=0
cc_344 N_C_c_406_n N_A_499_392#_c_691_n 0.0163652f $X=5.34 $Y=1.572 $X2=0 $Y2=0
cc_345 N_C_c_403_n N_A_499_392#_c_721_n 2.24111e-19 $X=4.735 $Y=1.885 $X2=0
+ $Y2=0
cc_346 N_C_c_404_n N_A_499_392#_c_685_n 0.00889577f $X=6.135 $Y=1.885 $X2=0
+ $Y2=0
cc_347 N_C_c_403_n N_A_962_392#_c_778_n 0.00155487f $X=4.735 $Y=1.885 $X2=0
+ $Y2=0
cc_348 N_C_c_404_n N_A_962_392#_c_778_n 0.00335044f $X=6.135 $Y=1.885 $X2=0
+ $Y2=0
cc_349 N_C_M1015_g N_VGND_c_799_n 0.00440341f $X=4.72 $Y=0.74 $X2=0 $Y2=0
cc_350 N_C_M1015_g N_VGND_c_803_n 0.00868136f $X=4.72 $Y=0.74 $X2=0 $Y2=0
cc_351 N_C_M1015_g N_VGND_c_804_n 0.00434272f $X=4.72 $Y=0.74 $X2=0 $Y2=0
cc_352 N_C_M1015_g N_VGND_c_805_n 4.32194e-19 $X=4.72 $Y=0.74 $X2=0 $Y2=0
cc_353 N_D_c_476_n N_VPWR_c_535_n 0.00291649f $X=5.235 $Y=1.885 $X2=0 $Y2=0
cc_354 N_D_c_478_n N_VPWR_c_535_n 0.00291649f $X=5.685 $Y=1.885 $X2=0 $Y2=0
cc_355 N_D_c_476_n N_VPWR_c_526_n 0.0036003f $X=5.235 $Y=1.885 $X2=0 $Y2=0
cc_356 N_D_c_478_n N_VPWR_c_526_n 0.00359599f $X=5.685 $Y=1.885 $X2=0 $Y2=0
cc_357 N_D_c_476_n N_A_499_392#_c_683_n 6.22908e-19 $X=5.235 $Y=1.885 $X2=0
+ $Y2=0
cc_358 N_D_c_476_n N_A_499_392#_c_690_n 9.39713e-19 $X=5.235 $Y=1.885 $X2=0
+ $Y2=0
cc_359 N_D_c_476_n N_A_499_392#_c_684_n 6.4283e-19 $X=5.235 $Y=1.885 $X2=0 $Y2=0
cc_360 N_D_c_476_n N_A_499_392#_c_691_n 0.0127059f $X=5.235 $Y=1.885 $X2=0 $Y2=0
cc_361 N_D_c_478_n N_A_499_392#_c_691_n 0.0110457f $X=5.685 $Y=1.885 $X2=0 $Y2=0
cc_362 N_D_c_476_n N_A_962_392#_c_778_n 0.0112102f $X=5.235 $Y=1.885 $X2=0 $Y2=0
cc_363 N_D_c_478_n N_A_962_392#_c_778_n 0.0112134f $X=5.685 $Y=1.885 $X2=0 $Y2=0
cc_364 N_D_c_470_n N_VGND_c_798_n 0.0025954f $X=6.285 $Y=0.85 $X2=0 $Y2=0
cc_365 N_D_c_473_n N_VGND_c_798_n 0.00213166f $X=6.45 $Y=0.42 $X2=0 $Y2=0
cc_366 N_D_c_474_n N_VGND_c_798_n 0.0221582f $X=6.45 $Y=0.42 $X2=0 $Y2=0
cc_367 N_D_c_466_n N_VGND_c_799_n 0.00753637f $X=5.22 $Y=1.185 $X2=0 $Y2=0
cc_368 N_D_c_470_n N_VGND_c_799_n 0.00358943f $X=6.285 $Y=0.85 $X2=0 $Y2=0
cc_369 N_D_c_474_n N_VGND_c_799_n 0.0125166f $X=6.45 $Y=0.42 $X2=0 $Y2=0
cc_370 N_D_c_466_n N_VGND_c_804_n 0.00230732f $X=5.22 $Y=1.185 $X2=0 $Y2=0
cc_371 N_D_c_466_n N_VGND_c_805_n 0.00971517f $X=5.22 $Y=1.185 $X2=0 $Y2=0
cc_372 N_D_c_471_n N_VGND_c_805_n 0.013425f $X=5.775 $Y=0.85 $X2=0 $Y2=0
cc_373 N_D_c_472_n N_VGND_c_805_n 8.10942e-19 $X=5.7 $Y=1.335 $X2=0 $Y2=0
cc_374 N_D_c_473_n N_VGND_c_805_n 0.00987736f $X=6.45 $Y=0.42 $X2=0 $Y2=0
cc_375 N_D_c_474_n N_VGND_c_805_n 0.0357573f $X=6.45 $Y=0.42 $X2=0 $Y2=0
cc_376 N_VPWR_M1010_d N_X_c_613_n 0.00451983f $X=0.135 $Y=1.84 $X2=0 $Y2=0
cc_377 N_VPWR_c_528_n N_X_c_613_n 0.0235383f $X=0.28 $Y=2.405 $X2=0 $Y2=0
cc_378 N_VPWR_c_528_n N_X_c_617_n 0.0255132f $X=0.28 $Y=2.405 $X2=0 $Y2=0
cc_379 N_VPWR_c_529_n N_X_c_617_n 0.0255132f $X=1.18 $Y=2.405 $X2=0 $Y2=0
cc_380 N_VPWR_c_532_n N_X_c_617_n 0.0101736f $X=1.015 $Y=3.33 $X2=0 $Y2=0
cc_381 N_VPWR_c_526_n N_X_c_617_n 0.0084208f $X=6.48 $Y=3.33 $X2=0 $Y2=0
cc_382 N_VPWR_c_529_n N_X_c_618_n 0.0255132f $X=1.18 $Y=2.405 $X2=0 $Y2=0
cc_383 N_VPWR_c_530_n N_X_c_618_n 0.0255132f $X=2.08 $Y=2.405 $X2=0 $Y2=0
cc_384 N_VPWR_c_533_n N_X_c_618_n 0.0101736f $X=1.915 $Y=3.33 $X2=0 $Y2=0
cc_385 N_VPWR_c_526_n N_X_c_618_n 0.0084208f $X=6.48 $Y=3.33 $X2=0 $Y2=0
cc_386 N_VPWR_M1016_d X 0.00454904f $X=1.93 $Y=1.84 $X2=0 $Y2=0
cc_387 N_VPWR_c_530_n X 0.0230252f $X=2.08 $Y=2.405 $X2=0 $Y2=0
cc_388 N_VPWR_M1011_d N_X_c_621_n 0.00201799f $X=1.03 $Y=1.84 $X2=0 $Y2=0
cc_389 N_VPWR_c_529_n N_X_c_621_n 0.0179913f $X=1.18 $Y=2.405 $X2=0 $Y2=0
cc_390 N_VPWR_c_530_n N_A_499_392#_c_682_n 0.0439499f $X=2.08 $Y=2.405 $X2=0
+ $Y2=0
cc_391 N_VPWR_c_534_n N_A_499_392#_c_682_n 0.0124046f $X=3.375 $Y=3.33 $X2=0
+ $Y2=0
cc_392 N_VPWR_c_526_n N_A_499_392#_c_682_n 0.0102675f $X=6.48 $Y=3.33 $X2=0
+ $Y2=0
cc_393 N_VPWR_M1000_d N_A_499_392#_c_699_n 0.0037709f $X=3.39 $Y=1.96 $X2=0
+ $Y2=0
cc_394 N_VPWR_c_535_n N_A_499_392#_c_684_n 0.0145938f $X=6.48 $Y=3.33 $X2=0
+ $Y2=0
cc_395 N_VPWR_c_526_n N_A_499_392#_c_684_n 0.0120466f $X=6.48 $Y=3.33 $X2=0
+ $Y2=0
cc_396 N_VPWR_c_526_n N_A_499_392#_c_691_n 0.0119345f $X=6.48 $Y=3.33 $X2=0
+ $Y2=0
cc_397 N_VPWR_c_535_n N_A_499_392#_c_685_n 0.0146513f $X=6.48 $Y=3.33 $X2=0
+ $Y2=0
cc_398 N_VPWR_c_526_n N_A_499_392#_c_685_n 0.0121202f $X=6.48 $Y=3.33 $X2=0
+ $Y2=0
cc_399 N_VPWR_c_531_n N_A_588_392#_c_750_n 0.0101517f $X=3.54 $Y=2.815 $X2=0
+ $Y2=0
cc_400 N_VPWR_c_534_n N_A_588_392#_c_750_n 0.0122801f $X=3.375 $Y=3.33 $X2=0
+ $Y2=0
cc_401 N_VPWR_c_526_n N_A_588_392#_c_750_n 0.0101678f $X=6.48 $Y=3.33 $X2=0
+ $Y2=0
cc_402 N_VPWR_M1000_d N_A_588_392#_c_756_n 0.0039506f $X=3.39 $Y=1.96 $X2=0
+ $Y2=0
cc_403 N_VPWR_c_531_n N_A_588_392#_c_756_n 0.0168789f $X=3.54 $Y=2.815 $X2=0
+ $Y2=0
cc_404 N_VPWR_c_526_n N_A_588_392#_c_756_n 0.0101191f $X=6.48 $Y=3.33 $X2=0
+ $Y2=0
cc_405 N_VPWR_c_526_n N_A_588_392#_c_754_n 0.00252518f $X=6.48 $Y=3.33 $X2=0
+ $Y2=0
cc_406 N_VPWR_c_531_n N_A_588_392#_c_751_n 0.00929383f $X=3.54 $Y=2.815 $X2=0
+ $Y2=0
cc_407 N_VPWR_c_535_n N_A_588_392#_c_751_n 0.0123494f $X=6.48 $Y=3.33 $X2=0
+ $Y2=0
cc_408 N_VPWR_c_526_n N_A_588_392#_c_751_n 0.0101947f $X=6.48 $Y=3.33 $X2=0
+ $Y2=0
cc_409 N_VPWR_c_535_n N_A_962_392#_c_778_n 0.0504896f $X=6.48 $Y=3.33 $X2=0
+ $Y2=0
cc_410 N_VPWR_c_526_n N_A_962_392#_c_778_n 0.0426127f $X=6.48 $Y=3.33 $X2=0
+ $Y2=0
cc_411 X N_A_499_392#_c_681_n 0.0172799f $X=2.075 $Y=1.95 $X2=0 $Y2=0
cc_412 N_X_c_614_n N_VGND_M1004_d 0.00250873f $X=1.615 $Y=1.065 $X2=0 $Y2=0
cc_413 N_X_c_612_n N_VGND_c_793_n 0.0243921f $X=0.78 $Y=0.515 $X2=0 $Y2=0
cc_414 N_X_c_613_n N_VGND_c_793_n 0.0370015f $X=0.73 $Y=2.15 $X2=0 $Y2=0
cc_415 N_X_c_612_n N_VGND_c_794_n 0.0180508f $X=0.78 $Y=0.515 $X2=0 $Y2=0
cc_416 N_X_c_614_n N_VGND_c_794_n 0.0210288f $X=1.615 $Y=1.065 $X2=0 $Y2=0
cc_417 N_X_c_615_n N_VGND_c_794_n 0.0180508f $X=1.78 $Y=0.515 $X2=0 $Y2=0
cc_418 N_X_c_615_n N_VGND_c_795_n 0.00585761f $X=1.78 $Y=0.515 $X2=0 $Y2=0
cc_419 N_X_c_612_n N_VGND_c_796_n 0.0144922f $X=0.78 $Y=0.515 $X2=0 $Y2=0
cc_420 N_X_c_615_n N_VGND_c_797_n 0.0146357f $X=1.78 $Y=0.515 $X2=0 $Y2=0
cc_421 N_X_c_612_n N_VGND_c_799_n 0.0118826f $X=0.78 $Y=0.515 $X2=0 $Y2=0
cc_422 N_X_c_615_n N_VGND_c_799_n 0.0121141f $X=1.78 $Y=0.515 $X2=0 $Y2=0
cc_423 N_A_499_392#_c_699_n N_A_588_392#_M1009_s 0.00527111f $X=4.345 $Y=2.055
+ $X2=-0.19 $Y2=1.66
cc_424 N_A_499_392#_c_699_n N_A_588_392#_M1001_s 0.00623879f $X=4.345 $Y=2.055
+ $X2=0 $Y2=0
cc_425 N_A_499_392#_c_699_n N_A_588_392#_c_752_n 0.0132885f $X=4.345 $Y=2.055
+ $X2=0 $Y2=0
cc_426 N_A_499_392#_c_682_n N_A_588_392#_c_750_n 0.0161022f $X=2.64 $Y=2.445
+ $X2=0 $Y2=0
cc_427 N_A_499_392#_c_699_n N_A_588_392#_c_756_n 0.0271649f $X=4.345 $Y=2.055
+ $X2=0 $Y2=0
cc_428 N_A_499_392#_c_699_n N_A_588_392#_c_754_n 0.018856f $X=4.345 $Y=2.055
+ $X2=0 $Y2=0
cc_429 N_A_499_392#_c_684_n N_A_588_392#_c_751_n 0.0161216f $X=4.51 $Y=2.815
+ $X2=0 $Y2=0
cc_430 N_A_499_392#_c_691_n N_A_962_392#_M1008_d 0.00690649f $X=6.245 $Y=2.445
+ $X2=-0.19 $Y2=1.66
cc_431 N_A_499_392#_c_691_n N_A_962_392#_M1017_s 0.00423551f $X=6.245 $Y=2.445
+ $X2=0 $Y2=0
cc_432 N_A_499_392#_c_684_n N_A_962_392#_c_778_n 0.0113199f $X=4.51 $Y=2.815
+ $X2=0 $Y2=0
cc_433 N_A_499_392#_c_691_n N_A_962_392#_c_778_n 0.0660711f $X=6.245 $Y=2.445
+ $X2=0 $Y2=0
cc_434 N_A_499_392#_c_685_n N_A_962_392#_c_778_n 0.0124625f $X=6.41 $Y=2.455
+ $X2=0 $Y2=0
