* File: sky130_fd_sc_hs__a32o_4.spice
* Created: Tue Sep  1 19:53:36 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hs__a32o_4.pex.spice"
.subckt sky130_fd_sc_hs__a32o_4  VNB VPB B2 B1 A2 A1 A3 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A3	A3
* A1	A1
* A2	A2
* B1	B1
* B2	B2
* VPB	VPB
* VNB	VNB
MM1005 N_X_M1005_d N_A_83_283#_M1005_g N_VGND_M1005_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.10915 AS=0.2109 PD=1.035 PS=2.05 NRD=0.804 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75003.5 A=0.111 P=1.78 MULT=1
MM1006 N_X_M1005_d N_A_83_283#_M1006_g N_VGND_M1006_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.10915 AS=0.1591 PD=1.035 PS=1.17 NRD=1.62 NRS=6.48 M=1 R=4.93333
+ SA=75000.7 SB=75003 A=0.111 P=1.78 MULT=1
MM1009 N_X_M1009_d N_A_83_283#_M1009_g N_VGND_M1006_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1591 PD=1.02 PS=1.17 NRD=0 NRS=17.832 M=1 R=4.93333 SA=75001.2
+ SB=75002.4 A=0.111 P=1.78 MULT=1
MM1017 N_X_M1009_d N_A_83_283#_M1017_g N_VGND_M1017_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.274229 PD=1.02 PS=1.6087 NRD=0 NRS=11.34 M=1 R=4.93333
+ SA=75001.7 SB=75002 A=0.111 P=1.78 MULT=1
MM1000 N_A_587_110#_M1000_d N_B2_M1000_g N_VGND_M1017_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.0896 AS=0.237171 PD=0.92 PS=1.3913 NRD=0 NRS=76.872 M=1 R=4.26667
+ SA=75002.6 SB=75001.4 A=0.096 P=1.58 MULT=1
MM1001 N_A_83_283#_M1001_d N_B1_M1001_g N_A_587_110#_M1000_d VNB NLOWVT L=0.15
+ W=0.64 AD=0.127887 AS=0.0896 PD=1.145 PS=0.92 NRD=15.936 NRS=0 M=1 R=4.26667
+ SA=75003 SB=75001 A=0.096 P=1.58 MULT=1
MM1012 N_A_83_283#_M1001_d N_B1_M1012_g N_A_587_110#_M1012_s VNB NLOWVT L=0.15
+ W=0.64 AD=0.127887 AS=0.0896 PD=1.145 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75002.8 SB=75000.7 A=0.096 P=1.58 MULT=1
MM1015 N_A_587_110#_M1012_s N_B2_M1015_g N_VGND_M1015_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.0896 AS=0.192025 PD=0.92 PS=1.99 NRD=0 NRS=13.116 M=1 R=4.26667
+ SA=75003.2 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1007 N_A_992_122#_M1007_d N_A2_M1007_g N_A_1079_122#_M1007_s VNB NLOWVT L=0.15
+ W=0.64 AD=0.1824 AS=0.0896 PD=1.85 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75002.6 A=0.096 P=1.58 MULT=1
MM1026 N_A_83_283#_M1026_d N_A1_M1026_g N_A_1079_122#_M1007_s VNB NLOWVT L=0.15
+ W=0.64 AD=0.0896 AS=0.0896 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.6 SB=75002.1 A=0.096 P=1.58 MULT=1
MM1027 N_A_83_283#_M1026_d N_A1_M1027_g N_A_1079_122#_M1027_s VNB NLOWVT L=0.15
+ W=0.64 AD=0.0896 AS=0.1152 PD=0.92 PS=1 NRD=0 NRS=0 M=1 R=4.26667 SA=75001.1
+ SB=75001.7 A=0.096 P=1.58 MULT=1
MM1024 N_A_992_122#_M1024_d N_A2_M1024_g N_A_1079_122#_M1027_s VNB NLOWVT L=0.15
+ W=0.64 AD=0.096 AS=0.1152 PD=0.94 PS=1 NRD=0 NRS=14.988 M=1 R=4.26667
+ SA=75001.6 SB=75001.2 A=0.096 P=1.58 MULT=1
MM1003 N_A_992_122#_M1024_d N_A3_M1003_g N_VGND_M1003_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.096 AS=0.12 PD=0.94 PS=1.015 NRD=3.744 NRS=1.872 M=1 R=4.26667 SA=75002
+ SB=75000.7 A=0.096 P=1.58 MULT=1
MM1008 N_A_992_122#_M1008_d N_A3_M1008_g N_VGND_M1003_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.1824 AS=0.12 PD=1.85 PS=1.015 NRD=0 NRS=15.936 M=1 R=4.26667 SA=75002.6
+ SB=75000.2 A=0.096 P=1.58 MULT=1
MM1010 N_VPWR_M1010_d N_A_83_283#_M1010_g N_X_M1010_s VPB PSHORT L=0.15 W=1.12
+ AD=0.3304 AS=0.168 PD=2.83 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75001.6 A=0.168 P=2.54 MULT=1
MM1011 N_VPWR_M1011_d N_A_83_283#_M1011_g N_X_M1010_s VPB PSHORT L=0.15 W=1.12
+ AD=0.196 AS=0.168 PD=1.47 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.7 SB=75001.2 A=0.168 P=2.54 MULT=1
MM1013 N_VPWR_M1011_d N_A_83_283#_M1013_g N_X_M1013_s VPB PSHORT L=0.15 W=1.12
+ AD=0.196 AS=0.168 PD=1.47 PS=1.42 NRD=10.5395 NRS=1.7533 M=1 R=7.46667
+ SA=75001.2 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1014 N_VPWR_M1014_d N_A_83_283#_M1014_g N_X_M1013_s VPB PSHORT L=0.15 W=1.12
+ AD=0.3304 AS=0.168 PD=2.83 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.6 SB=75000.2 A=0.168 P=2.54 MULT=1
MM1021 N_A_509_392#_M1021_d N_B2_M1021_g N_A_83_283#_M1021_s VPB PSHORT L=0.15
+ W=1 AD=0.295 AS=0.175 PD=2.59 PS=1.35 NRD=1.9503 NRS=11.8003 M=1 R=6.66667
+ SA=75000.2 SB=75005 A=0.15 P=2.3 MULT=1
MM1020 N_A_83_283#_M1021_s N_B1_M1020_g N_A_509_392#_M1020_s VPB PSHORT L=0.15
+ W=1 AD=0.175 AS=0.175 PD=1.35 PS=1.35 NRD=1.9503 NRS=11.8003 M=1 R=6.66667
+ SA=75000.7 SB=75004.5 A=0.15 P=2.3 MULT=1
MM1023 N_A_83_283#_M1023_d N_B1_M1023_g N_A_509_392#_M1020_s VPB PSHORT L=0.15
+ W=1 AD=0.175 AS=0.175 PD=1.35 PS=1.35 NRD=11.8003 NRS=1.9503 M=1 R=6.66667
+ SA=75001.2 SB=75004 A=0.15 P=2.3 MULT=1
MM1025 N_A_509_392#_M1025_d N_B2_M1025_g N_A_83_283#_M1023_d VPB PSHORT L=0.15
+ W=1 AD=0.2725 AS=0.175 PD=1.545 PS=1.35 NRD=25.5903 NRS=1.9503 M=1 R=6.66667
+ SA=75001.7 SB=75003.5 A=0.15 P=2.3 MULT=1
MM1016 N_A_509_392#_M1025_d N_A2_M1016_g N_VPWR_M1016_s VPB PSHORT L=0.15 W=1
+ AD=0.2725 AS=0.2325 PD=1.545 PS=1.465 NRD=26.5753 NRS=12.7853 M=1 R=6.66667
+ SA=75002.4 SB=75002.8 A=0.15 P=2.3 MULT=1
MM1002 N_A_509_392#_M1002_d N_A1_M1002_g N_VPWR_M1016_s VPB PSHORT L=0.15 W=1
+ AD=0.16 AS=0.2325 PD=1.32 PS=1.465 NRD=1.9503 NRS=23.6203 M=1 R=6.66667
+ SA=75003 SB=75002.1 A=0.15 P=2.3 MULT=1
MM1004 N_A_509_392#_M1002_d N_A1_M1004_g N_VPWR_M1004_s VPB PSHORT L=0.15 W=1
+ AD=0.16 AS=0.18 PD=1.32 PS=1.36 NRD=5.8903 NRS=10.8153 M=1 R=6.66667
+ SA=75003.5 SB=75001.7 A=0.15 P=2.3 MULT=1
MM1018 N_A_509_392#_M1018_d N_A2_M1018_g N_VPWR_M1004_s VPB PSHORT L=0.15 W=1
+ AD=0.15 AS=0.18 PD=1.3 PS=1.36 NRD=1.9503 NRS=4.9053 M=1 R=6.66667 SA=75004
+ SB=75001.2 A=0.15 P=2.3 MULT=1
MM1019 N_A_509_392#_M1018_d N_A3_M1019_g N_VPWR_M1019_s VPB PSHORT L=0.15 W=1
+ AD=0.15 AS=0.175 PD=1.3 PS=1.35 NRD=1.9503 NRS=1.9503 M=1 R=6.66667 SA=75004.5
+ SB=75000.7 A=0.15 P=2.3 MULT=1
MM1022 N_A_509_392#_M1022_d N_A3_M1022_g N_VPWR_M1019_s VPB PSHORT L=0.15 W=1
+ AD=0.295 AS=0.175 PD=2.59 PS=1.35 NRD=1.9503 NRS=11.8003 M=1 R=6.66667
+ SA=75005 SB=75000.2 A=0.15 P=2.3 MULT=1
DX28_noxref VNB VPB NWDIODE A=15.669 P=21.04
*
.include "sky130_fd_sc_hs__a32o_4.pxi.spice"
*
.ends
*
*
