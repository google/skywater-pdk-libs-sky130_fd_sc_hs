* File: sky130_fd_sc_hs__xor3_4.pxi.spice
* Created: Thu Aug 27 21:13:34 2020
* 
x_PM_SKY130_FD_SC_HS__XOR3_4%A_74_294# N_A_74_294#_M1025_d N_A_74_294#_M1027_d
+ N_A_74_294#_M1006_d N_A_74_294#_M1002_d N_A_74_294#_M1012_g
+ N_A_74_294#_c_205_n N_A_74_294#_M1008_g N_A_74_294#_c_206_n
+ N_A_74_294#_c_212_n N_A_74_294#_c_213_n N_A_74_294#_c_214_n
+ N_A_74_294#_c_215_n N_A_74_294#_c_216_n N_A_74_294#_c_207_n
+ N_A_74_294#_c_218_n N_A_74_294#_c_219_n N_A_74_294#_c_220_n
+ N_A_74_294#_c_208_n N_A_74_294#_c_209_n PM_SKY130_FD_SC_HS__XOR3_4%A_74_294#
x_PM_SKY130_FD_SC_HS__XOR3_4%A N_A_c_318_n N_A_M1006_g N_A_c_319_n N_A_M1025_g A
+ PM_SKY130_FD_SC_HS__XOR3_4%A
x_PM_SKY130_FD_SC_HS__XOR3_4%A_397_320# N_A_397_320#_M1026_s
+ N_A_397_320#_M1003_s N_A_397_320#_c_369_n N_A_397_320#_M1011_g
+ N_A_397_320#_c_354_n N_A_397_320#_M1022_g N_A_397_320#_c_371_n
+ N_A_397_320#_M1002_g N_A_397_320#_c_356_n N_A_397_320#_M1027_g
+ N_A_397_320#_c_358_n N_A_397_320#_c_359_n N_A_397_320#_c_360_n
+ N_A_397_320#_c_361_n N_A_397_320#_c_362_n N_A_397_320#_c_363_n
+ N_A_397_320#_c_364_n N_A_397_320#_c_391_n N_A_397_320#_c_365_n
+ N_A_397_320#_c_366_n N_A_397_320#_c_367_n N_A_397_320#_c_368_n
+ PM_SKY130_FD_SC_HS__XOR3_4%A_397_320#
x_PM_SKY130_FD_SC_HS__XOR3_4%B N_B_c_483_n N_B_M1023_g N_B_c_484_n N_B_M1019_g
+ N_B_c_471_n N_B_c_472_n N_B_c_485_n N_B_c_486_n N_B_c_487_n N_B_M1004_g
+ N_B_c_488_n N_B_M1014_g N_B_c_474_n N_B_c_475_n N_B_c_476_n N_B_c_477_n
+ N_B_c_478_n N_B_M1003_g N_B_c_479_n N_B_M1026_g N_B_c_491_n N_B_c_492_n
+ N_B_c_480_n N_B_c_481_n B PM_SKY130_FD_SC_HS__XOR3_4%B
x_PM_SKY130_FD_SC_HS__XOR3_4%A_1155_284# N_A_1155_284#_M1001_s
+ N_A_1155_284#_M1010_s N_A_1155_284#_c_606_n N_A_1155_284#_M1009_g
+ N_A_1155_284#_M1016_g N_A_1155_284#_c_612_n N_A_1155_284#_c_613_n
+ N_A_1155_284#_c_614_n N_A_1155_284#_c_615_n N_A_1155_284#_c_608_n
+ N_A_1155_284#_c_617_n N_A_1155_284#_c_609_n N_A_1155_284#_c_610_n
+ PM_SKY130_FD_SC_HS__XOR3_4%A_1155_284#
x_PM_SKY130_FD_SC_HS__XOR3_4%C N_C_c_692_n N_C_M1020_g N_C_M1021_g N_C_c_694_n
+ N_C_c_695_n N_C_c_696_n N_C_c_702_n N_C_c_703_n N_C_M1010_g N_C_c_697_n
+ N_C_M1001_g N_C_c_698_n N_C_c_699_n C PM_SKY130_FD_SC_HS__XOR3_4%C
x_PM_SKY130_FD_SC_HS__XOR3_4%A_1218_388# N_A_1218_388#_M1016_d
+ N_A_1218_388#_M1009_d N_A_1218_388#_c_778_n N_A_1218_388#_M1000_g
+ N_A_1218_388#_M1007_g N_A_1218_388#_c_779_n N_A_1218_388#_M1005_g
+ N_A_1218_388#_M1017_g N_A_1218_388#_c_780_n N_A_1218_388#_M1013_g
+ N_A_1218_388#_M1018_g N_A_1218_388#_c_781_n N_A_1218_388#_M1015_g
+ N_A_1218_388#_M1024_g N_A_1218_388#_c_774_n N_A_1218_388#_c_792_n
+ N_A_1218_388#_c_864_p N_A_1218_388#_c_783_n N_A_1218_388#_c_784_n
+ N_A_1218_388#_c_785_n N_A_1218_388#_c_817_p N_A_1218_388#_c_775_n
+ N_A_1218_388#_c_776_n N_A_1218_388#_c_777_n
+ PM_SKY130_FD_SC_HS__XOR3_4%A_1218_388#
x_PM_SKY130_FD_SC_HS__XOR3_4%A_27_118# N_A_27_118#_M1012_s N_A_27_118#_M1022_d
+ N_A_27_118#_M1008_s N_A_27_118#_M1011_d N_A_27_118#_c_909_n
+ N_A_27_118#_c_910_n N_A_27_118#_c_918_n N_A_27_118#_c_919_n
+ N_A_27_118#_c_911_n N_A_27_118#_c_912_n N_A_27_118#_c_913_n
+ N_A_27_118#_c_914_n N_A_27_118#_c_915_n N_A_27_118#_c_916_n
+ N_A_27_118#_c_917_n PM_SKY130_FD_SC_HS__XOR3_4%A_27_118#
x_PM_SKY130_FD_SC_HS__XOR3_4%VPWR N_VPWR_M1008_d N_VPWR_M1003_d N_VPWR_M1010_d
+ N_VPWR_M1005_s N_VPWR_M1015_s N_VPWR_c_994_n N_VPWR_c_995_n N_VPWR_c_996_n
+ N_VPWR_c_997_n N_VPWR_c_998_n N_VPWR_c_999_n N_VPWR_c_1000_n N_VPWR_c_1001_n
+ N_VPWR_c_1046_n VPWR N_VPWR_c_1002_n N_VPWR_c_1003_n N_VPWR_c_1004_n
+ N_VPWR_c_1005_n N_VPWR_c_1006_n N_VPWR_c_1007_n N_VPWR_c_1008_n
+ N_VPWR_c_1009_n N_VPWR_c_993_n PM_SKY130_FD_SC_HS__XOR3_4%VPWR
x_PM_SKY130_FD_SC_HS__XOR3_4%A_323_392# N_A_323_392#_M1014_d
+ N_A_323_392#_M1016_s N_A_323_392#_M1023_d N_A_323_392#_M1020_d
+ N_A_323_392#_c_1117_n N_A_323_392#_c_1119_n N_A_323_392#_c_1112_n
+ N_A_323_392#_c_1104_n N_A_323_392#_c_1105_n N_A_323_392#_c_1106_n
+ N_A_323_392#_c_1151_n N_A_323_392#_c_1107_n N_A_323_392#_c_1155_n
+ N_A_323_392#_c_1108_n N_A_323_392#_c_1109_n N_A_323_392#_c_1110_n
+ N_A_323_392#_c_1111_n N_A_323_392#_c_1115_n N_A_323_392#_c_1116_n
+ PM_SKY130_FD_SC_HS__XOR3_4%A_323_392#
x_PM_SKY130_FD_SC_HS__XOR3_4%A_416_118# N_A_416_118#_M1019_d
+ N_A_416_118#_M1021_d N_A_416_118#_M1004_d N_A_416_118#_M1009_s
+ N_A_416_118#_c_1235_n N_A_416_118#_c_1236_n N_A_416_118#_c_1237_n
+ N_A_416_118#_c_1238_n N_A_416_118#_c_1239_n N_A_416_118#_c_1240_n
+ N_A_416_118#_c_1291_n N_A_416_118#_c_1241_n N_A_416_118#_c_1242_n
+ N_A_416_118#_c_1243_n N_A_416_118#_c_1246_n N_A_416_118#_c_1247_n
+ N_A_416_118#_c_1248_n N_A_416_118#_c_1249_n N_A_416_118#_c_1250_n
+ N_A_416_118#_c_1244_n PM_SKY130_FD_SC_HS__XOR3_4%A_416_118#
x_PM_SKY130_FD_SC_HS__XOR3_4%X N_X_M1007_s N_X_M1018_s N_X_M1000_d N_X_M1013_d
+ N_X_c_1360_n N_X_c_1356_n N_X_c_1357_n N_X_c_1373_n N_X_c_1358_n N_X_c_1361_n
+ N_X_c_1359_n N_X_c_1390_n N_X_c_1393_n X X X X N_X_c_1399_n X
+ PM_SKY130_FD_SC_HS__XOR3_4%X
x_PM_SKY130_FD_SC_HS__XOR3_4%VGND N_VGND_M1012_d N_VGND_M1026_d N_VGND_M1001_d
+ N_VGND_M1017_d N_VGND_M1024_d N_VGND_c_1419_n N_VGND_c_1420_n N_VGND_c_1421_n
+ N_VGND_c_1422_n N_VGND_c_1423_n N_VGND_c_1424_n N_VGND_c_1425_n
+ N_VGND_c_1426_n VGND N_VGND_c_1427_n N_VGND_c_1428_n N_VGND_c_1429_n
+ N_VGND_c_1430_n N_VGND_c_1431_n N_VGND_c_1432_n N_VGND_c_1433_n
+ PM_SKY130_FD_SC_HS__XOR3_4%VGND
cc_1 VNB N_A_74_294#_M1012_g 0.0318606f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.91
cc_2 VNB N_A_74_294#_c_205_n 0.0192113f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.885
cc_3 VNB N_A_74_294#_c_206_n 0.00510846f $X=-0.19 $Y=-0.245 $X2=0.535 $Y2=1.635
cc_4 VNB N_A_74_294#_c_207_n 0.00892299f $X=-0.19 $Y=-0.245 $X2=1.54 $Y2=1.085
cc_5 VNB N_A_74_294#_c_208_n 0.00297214f $X=-0.19 $Y=-0.245 $X2=3.99 $Y2=1.905
cc_6 VNB N_A_74_294#_c_209_n 8.73313e-19 $X=-0.19 $Y=-0.245 $X2=4.24 $Y2=1.1
cc_7 VNB N_A_c_318_n 0.0312171f $X=-0.19 $Y=-0.245 $X2=1.24 $Y2=0.59
cc_8 VNB N_A_c_319_n 0.020485f $X=-0.19 $Y=-0.245 $X2=3.28 $Y2=1.895
cc_9 VNB A 0.00502784f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_397_320#_c_354_n 0.00886979f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_397_320#_M1022_g 0.0361557f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.91
cc_12 VNB N_A_397_320#_c_356_n 0.00997588f $X=-0.19 $Y=-0.245 $X2=0.562
+ $Y2=1.635
cc_13 VNB N_A_397_320#_M1027_g 0.0194039f $X=-0.19 $Y=-0.245 $X2=1.065 $Y2=1.925
cc_14 VNB N_A_397_320#_c_358_n 0.00687282f $X=-0.19 $Y=-0.245 $X2=1.23 $Y2=2.01
cc_15 VNB N_A_397_320#_c_359_n 9.55161e-19 $X=-0.19 $Y=-0.245 $X2=1.23 $Y2=2.105
cc_16 VNB N_A_397_320#_c_360_n 0.0168028f $X=-0.19 $Y=-0.245 $X2=1.23 $Y2=2.815
cc_17 VNB N_A_397_320#_c_361_n 0.00840643f $X=-0.19 $Y=-0.245 $X2=1.23 $Y2=2.815
cc_18 VNB N_A_397_320#_c_362_n 0.00123369f $X=-0.19 $Y=-0.245 $X2=1.395 $Y2=2.99
cc_19 VNB N_A_397_320#_c_363_n 0.00538737f $X=-0.19 $Y=-0.245 $X2=1.54 $Y2=1.84
cc_20 VNB N_A_397_320#_c_364_n 3.26207e-19 $X=-0.19 $Y=-0.245 $X2=1.54 $Y2=1.085
cc_21 VNB N_A_397_320#_c_365_n 0.00571645f $X=-0.19 $Y=-0.245 $X2=1.23 $Y2=1.925
cc_22 VNB N_A_397_320#_c_366_n 0.00142557f $X=-0.19 $Y=-0.245 $X2=4.08 $Y2=1.1
cc_23 VNB N_A_397_320#_c_367_n 0.0249124f $X=-0.19 $Y=-0.245 $X2=4.08 $Y2=1.1
cc_24 VNB N_A_397_320#_c_368_n 8.51178e-19 $X=-0.19 $Y=-0.245 $X2=4.24 $Y2=1.1
cc_25 VNB N_B_M1019_g 0.0421415f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_B_c_471_n 0.0647382f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_B_c_472_n 0.012806f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_B_M1014_g 0.0355273f $X=-0.19 $Y=-0.245 $X2=0.562 $Y2=1.635
cc_29 VNB N_B_c_474_n 0.0890197f $X=-0.19 $Y=-0.245 $X2=0.535 $Y2=1.635
cc_30 VNB N_B_c_475_n 0.00530041f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=1.925
cc_31 VNB N_B_c_476_n 0.0679642f $X=-0.19 $Y=-0.245 $X2=1.23 $Y2=2.905
cc_32 VNB N_B_c_477_n 0.0200225f $X=-0.19 $Y=-0.245 $X2=1.23 $Y2=2.105
cc_33 VNB N_B_c_478_n 0.0557702f $X=-0.19 $Y=-0.245 $X2=1.23 $Y2=2.815
cc_34 VNB N_B_c_479_n 0.0201399f $X=-0.19 $Y=-0.245 $X2=1.395 $Y2=2.99
cc_35 VNB N_B_c_480_n 0.00749069f $X=-0.19 $Y=-0.245 $X2=3.74 $Y2=2.905
cc_36 VNB N_B_c_481_n 0.00608976f $X=-0.19 $Y=-0.245 $X2=4.24 $Y2=1.265
cc_37 VNB B 0.00646241f $X=-0.19 $Y=-0.245 $X2=4.24 $Y2=1.905
cc_38 VNB N_A_1155_284#_c_606_n 0.0279689f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_1155_284#_M1016_g 0.0230894f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_1155_284#_c_608_n 0.00167734f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=1.925
cc_41 VNB N_A_1155_284#_c_609_n 0.0188721f $X=-0.19 $Y=-0.245 $X2=1.23 $Y2=2.105
cc_42 VNB N_A_1155_284#_c_610_n 0.00392074f $X=-0.19 $Y=-0.245 $X2=1.54 $Y2=1.84
cc_43 VNB N_C_c_692_n 0.0123259f $X=-0.19 $Y=-0.245 $X2=1.24 $Y2=0.59
cc_44 VNB N_C_M1021_g 0.024649f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_C_c_694_n 0.0238657f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_C_c_695_n 0.0657705f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_C_c_696_n 0.00977486f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_C_c_697_n 0.0210961f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.885
cc_49 VNB N_C_c_698_n 0.0141574f $X=-0.19 $Y=-0.245 $X2=0.535 $Y2=1.635
cc_50 VNB N_C_c_699_n 0.0081686f $X=-0.19 $Y=-0.245 $X2=0.535 $Y2=1.635
cc_51 VNB C 0.00125263f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_A_1218_388#_M1007_g 0.0239049f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_A_1218_388#_M1017_g 0.0182194f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.46
cc_54 VNB N_A_1218_388#_M1018_g 0.0182166f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=1.925
cc_55 VNB N_A_1218_388#_M1024_g 0.0240808f $X=-0.19 $Y=-0.245 $X2=3.655 $Y2=2.99
cc_56 VNB N_A_1218_388#_c_774_n 0.00547693f $X=-0.19 $Y=-0.245 $X2=3.74
+ $Y2=2.755
cc_57 VNB N_A_1218_388#_c_775_n 0.00173929f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_A_1218_388#_c_776_n 0.0696069f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_A_1218_388#_c_777_n 0.135981f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_A_27_118#_c_909_n 0.0117778f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.47
cc_61 VNB N_A_27_118#_c_910_n 0.0125547f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.91
cc_62 VNB N_A_27_118#_c_911_n 0.0100203f $X=-0.19 $Y=-0.245 $X2=0.562 $Y2=1.635
cc_63 VNB N_A_27_118#_c_912_n 0.00247756f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_A_27_118#_c_913_n 9.46905e-19 $X=-0.19 $Y=-0.245 $X2=1.23 $Y2=2.01
cc_65 VNB N_A_27_118#_c_914_n 0.0189945f $X=-0.19 $Y=-0.245 $X2=1.23 $Y2=2.105
cc_66 VNB N_A_27_118#_c_915_n 0.00353847f $X=-0.19 $Y=-0.245 $X2=1.23 $Y2=2.815
cc_67 VNB N_A_27_118#_c_916_n 0.0124576f $X=-0.19 $Y=-0.245 $X2=1.54 $Y2=1.84
cc_68 VNB N_A_27_118#_c_917_n 0.0195252f $X=-0.19 $Y=-0.245 $X2=1.54 $Y2=1.085
cc_69 VNB N_VPWR_c_993_n 0.442315f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_A_323_392#_c_1104_n 0.0108249f $X=-0.19 $Y=-0.245 $X2=0.535
+ $Y2=1.635
cc_71 VNB N_A_323_392#_c_1105_n 0.0225385f $X=-0.19 $Y=-0.245 $X2=0.535
+ $Y2=1.635
cc_72 VNB N_A_323_392#_c_1106_n 0.00289943f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_A_323_392#_c_1107_n 0.00782494f $X=-0.19 $Y=-0.245 $X2=1.23 $Y2=2.01
cc_74 VNB N_A_323_392#_c_1108_n 0.00943365f $X=-0.19 $Y=-0.245 $X2=1.23
+ $Y2=2.815
cc_75 VNB N_A_323_392#_c_1109_n 0.0416477f $X=-0.19 $Y=-0.245 $X2=3.655 $Y2=2.99
cc_76 VNB N_A_323_392#_c_1110_n 0.00510988f $X=-0.19 $Y=-0.245 $X2=1.395
+ $Y2=2.99
cc_77 VNB N_A_323_392#_c_1111_n 0.0159377f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_A_416_118#_c_1235_n 0.00381805f $X=-0.19 $Y=-0.245 $X2=0.495
+ $Y2=0.91
cc_79 VNB N_A_416_118#_c_1236_n 0.0116789f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.46
cc_80 VNB N_A_416_118#_c_1237_n 0.00446241f $X=-0.19 $Y=-0.245 $X2=0.562
+ $Y2=1.84
cc_81 VNB N_A_416_118#_c_1238_n 0.00421867f $X=-0.19 $Y=-0.245 $X2=0.535
+ $Y2=1.635
cc_82 VNB N_A_416_118#_c_1239_n 0.0117566f $X=-0.19 $Y=-0.245 $X2=1.23 $Y2=2.01
cc_83 VNB N_A_416_118#_c_1240_n 0.00432371f $X=-0.19 $Y=-0.245 $X2=1.23
+ $Y2=2.905
cc_84 VNB N_A_416_118#_c_1241_n 0.00331446f $X=-0.19 $Y=-0.245 $X2=1.23
+ $Y2=2.815
cc_85 VNB N_A_416_118#_c_1242_n 0.00111916f $X=-0.19 $Y=-0.245 $X2=1.23
+ $Y2=2.815
cc_86 VNB N_A_416_118#_c_1243_n 0.00389878f $X=-0.19 $Y=-0.245 $X2=1.54
+ $Y2=1.085
cc_87 VNB N_A_416_118#_c_1244_n 0.00833339f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_88 VNB N_X_c_1356_n 0.00240191f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.46
cc_89 VNB N_X_c_1357_n 0.00136893f $X=-0.19 $Y=-0.245 $X2=0.535 $Y2=1.635
cc_90 VNB N_X_c_1358_n 0.00336962f $X=-0.19 $Y=-0.245 $X2=1.23 $Y2=2.105
cc_91 VNB N_X_c_1359_n 6.54478e-19 $X=-0.19 $Y=-0.245 $X2=3.655 $Y2=2.99
cc_92 VNB N_VGND_c_1419_n 0.0106771f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.46
cc_93 VNB N_VGND_c_1420_n 0.0133176f $X=-0.19 $Y=-0.245 $X2=0.535 $Y2=1.635
cc_94 VNB N_VGND_c_1421_n 0.019013f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_95 VNB N_VGND_c_1422_n 0.00877682f $X=-0.19 $Y=-0.245 $X2=1.23 $Y2=2.905
cc_96 VNB N_VGND_c_1423_n 0.0118677f $X=-0.19 $Y=-0.245 $X2=1.23 $Y2=2.105
cc_97 VNB N_VGND_c_1424_n 0.0508226f $X=-0.19 $Y=-0.245 $X2=1.23 $Y2=2.815
cc_98 VNB N_VGND_c_1425_n 0.106119f $X=-0.19 $Y=-0.245 $X2=1.54 $Y2=1.84
cc_99 VNB N_VGND_c_1426_n 0.00478335f $X=-0.19 $Y=-0.245 $X2=1.54 $Y2=1.085
cc_100 VNB N_VGND_c_1427_n 0.0193471f $X=-0.19 $Y=-0.245 $X2=3.74 $Y2=2.755
cc_101 VNB N_VGND_c_1428_n 0.0701054f $X=-0.19 $Y=-0.245 $X2=4.08 $Y2=1.1
cc_102 VNB N_VGND_c_1429_n 0.0172524f $X=-0.19 $Y=-0.245 $X2=0.535 $Y2=1.635
cc_103 VNB N_VGND_c_1430_n 0.0267154f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_104 VNB N_VGND_c_1431_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_105 VNB N_VGND_c_1432_n 0.00326991f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_106 VNB N_VGND_c_1433_n 0.547849f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_107 VPB N_A_74_294#_c_205_n 0.0408211f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.885
cc_108 VPB N_A_74_294#_c_206_n 4.104e-19 $X=-0.19 $Y=1.66 $X2=0.535 $Y2=1.635
cc_109 VPB N_A_74_294#_c_212_n 0.00721425f $X=-0.19 $Y=1.66 $X2=1.065 $Y2=1.925
cc_110 VPB N_A_74_294#_c_213_n 6.94896e-19 $X=-0.19 $Y=1.66 $X2=0.7 $Y2=1.925
cc_111 VPB N_A_74_294#_c_214_n 0.00102784f $X=-0.19 $Y=1.66 $X2=1.23 $Y2=2.105
cc_112 VPB N_A_74_294#_c_215_n 0.0427434f $X=-0.19 $Y=1.66 $X2=3.655 $Y2=2.99
cc_113 VPB N_A_74_294#_c_216_n 0.00233563f $X=-0.19 $Y=1.66 $X2=1.395 $Y2=2.99
cc_114 VPB N_A_74_294#_c_207_n 0.00381963f $X=-0.19 $Y=1.66 $X2=1.54 $Y2=1.085
cc_115 VPB N_A_74_294#_c_218_n 0.0052774f $X=-0.19 $Y=1.66 $X2=3.74 $Y2=2.905
cc_116 VPB N_A_74_294#_c_219_n 0.00848935f $X=-0.19 $Y=1.66 $X2=1.54 $Y2=1.925
cc_117 VPB N_A_74_294#_c_220_n 0.0117238f $X=-0.19 $Y=1.66 $X2=3.74 $Y2=2.07
cc_118 VPB N_A_74_294#_c_208_n 0.0031888f $X=-0.19 $Y=1.66 $X2=3.99 $Y2=1.905
cc_119 VPB N_A_c_318_n 0.0343237f $X=-0.19 $Y=1.66 $X2=1.24 $Y2=0.59
cc_120 VPB A 0.00185801f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_121 VPB N_A_397_320#_c_369_n 0.0140072f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_122 VPB N_A_397_320#_c_354_n 0.0108743f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_123 VPB N_A_397_320#_c_371_n 0.0156432f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.46
cc_124 VPB N_A_397_320#_c_356_n 0.0136064f $X=-0.19 $Y=1.66 $X2=0.562 $Y2=1.635
cc_125 VPB N_A_397_320#_c_358_n 0.0150712f $X=-0.19 $Y=1.66 $X2=1.23 $Y2=2.01
cc_126 VPB N_A_397_320#_c_359_n 0.00801079f $X=-0.19 $Y=1.66 $X2=1.23 $Y2=2.105
cc_127 VPB N_A_397_320#_c_360_n 0.0169171f $X=-0.19 $Y=1.66 $X2=1.23 $Y2=2.815
cc_128 VPB N_A_397_320#_c_361_n 0.00751716f $X=-0.19 $Y=1.66 $X2=1.23 $Y2=2.815
cc_129 VPB N_A_397_320#_c_365_n 0.00527178f $X=-0.19 $Y=1.66 $X2=1.23 $Y2=1.925
cc_130 VPB N_A_397_320#_c_366_n 4.70948e-19 $X=-0.19 $Y=1.66 $X2=4.08 $Y2=1.1
cc_131 VPB N_A_397_320#_c_367_n 0.0142779f $X=-0.19 $Y=1.66 $X2=4.08 $Y2=1.1
cc_132 VPB N_B_c_483_n 0.0169801f $X=-0.19 $Y=1.66 $X2=1.24 $Y2=0.59
cc_133 VPB N_B_c_484_n 0.0634257f $X=-0.19 $Y=1.66 $X2=3.28 $Y2=1.895
cc_134 VPB N_B_c_485_n 0.00953984f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_135 VPB N_B_c_486_n 0.0139787f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.47
cc_136 VPB N_B_c_487_n 0.0142822f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.91
cc_137 VPB N_B_c_488_n 0.115795f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.885
cc_138 VPB N_B_c_475_n 0.0893865f $X=-0.19 $Y=1.66 $X2=0.7 $Y2=1.925
cc_139 VPB N_B_c_478_n 0.026285f $X=-0.19 $Y=1.66 $X2=1.23 $Y2=2.815
cc_140 VPB N_B_c_491_n 0.0285986f $X=-0.19 $Y=1.66 $X2=1.54 $Y2=1.085
cc_141 VPB N_B_c_492_n 0.00898645f $X=-0.19 $Y=1.66 $X2=3.74 $Y2=2.755
cc_142 VPB N_A_1155_284#_c_606_n 0.0459662f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_143 VPB N_A_1155_284#_c_612_n 0.00319492f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.91
cc_144 VPB N_A_1155_284#_c_613_n 0.038282f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_145 VPB N_A_1155_284#_c_614_n 0.00795758f $X=-0.19 $Y=1.66 $X2=0.505
+ $Y2=1.885
cc_146 VPB N_A_1155_284#_c_615_n 0.00552058f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.46
cc_147 VPB N_A_1155_284#_c_608_n 8.26712e-19 $X=-0.19 $Y=1.66 $X2=0.7 $Y2=1.925
cc_148 VPB N_A_1155_284#_c_617_n 0.00589786f $X=-0.19 $Y=1.66 $X2=1.23 $Y2=2.105
cc_149 VPB N_A_1155_284#_c_609_n 0.0039909f $X=-0.19 $Y=1.66 $X2=1.23 $Y2=2.105
cc_150 VPB N_C_c_692_n 0.0313551f $X=-0.19 $Y=1.66 $X2=1.24 $Y2=0.59
cc_151 VPB N_C_c_702_n 0.0383247f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_152 VPB N_C_c_703_n 0.0183557f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.91
cc_153 VPB N_C_c_698_n 0.0143712f $X=-0.19 $Y=1.66 $X2=0.535 $Y2=1.635
cc_154 VPB N_C_c_699_n 0.015802f $X=-0.19 $Y=1.66 $X2=0.535 $Y2=1.635
cc_155 VPB C 0.00204899f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_156 VPB N_A_1218_388#_c_778_n 0.0162423f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_157 VPB N_A_1218_388#_c_779_n 0.0158491f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.91
cc_158 VPB N_A_1218_388#_c_780_n 0.0158704f $X=-0.19 $Y=1.66 $X2=0.562 $Y2=1.635
cc_159 VPB N_A_1218_388#_c_781_n 0.0174349f $X=-0.19 $Y=1.66 $X2=1.23 $Y2=2.905
cc_160 VPB N_A_1218_388#_c_774_n 0.00215497f $X=-0.19 $Y=1.66 $X2=3.74 $Y2=2.755
cc_161 VPB N_A_1218_388#_c_783_n 0.00193385f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_162 VPB N_A_1218_388#_c_784_n 0.00502419f $X=-0.19 $Y=1.66 $X2=4.24 $Y2=1.1
cc_163 VPB N_A_1218_388#_c_785_n 0.00313822f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_164 VPB N_A_1218_388#_c_775_n 0.00459217f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_165 VPB N_A_1218_388#_c_777_n 0.0301352f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_166 VPB N_A_27_118#_c_918_n 0.00536733f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.885
cc_167 VPB N_A_27_118#_c_919_n 0.0279419f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.46
cc_168 VPB N_A_27_118#_c_913_n 0.0027274f $X=-0.19 $Y=1.66 $X2=1.23 $Y2=2.01
cc_169 VPB N_A_27_118#_c_917_n 0.0220788f $X=-0.19 $Y=1.66 $X2=1.54 $Y2=1.085
cc_170 VPB N_VPWR_c_994_n 0.00609828f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.46
cc_171 VPB N_VPWR_c_995_n 0.0274034f $X=-0.19 $Y=1.66 $X2=0.535 $Y2=1.635
cc_172 VPB N_VPWR_c_996_n 0.00158678f $X=-0.19 $Y=1.66 $X2=1.23 $Y2=2.905
cc_173 VPB N_VPWR_c_997_n 0.0131442f $X=-0.19 $Y=1.66 $X2=1.23 $Y2=2.815
cc_174 VPB N_VPWR_c_998_n 0.0218132f $X=-0.19 $Y=1.66 $X2=1.23 $Y2=2.815
cc_175 VPB N_VPWR_c_999_n 0.0096968f $X=-0.19 $Y=1.66 $X2=1.54 $Y2=1.085
cc_176 VPB N_VPWR_c_1000_n 0.0106521f $X=-0.19 $Y=1.66 $X2=3.74 $Y2=2.905
cc_177 VPB N_VPWR_c_1001_n 0.0645756f $X=-0.19 $Y=1.66 $X2=4.24 $Y2=1.905
cc_178 VPB N_VPWR_c_1002_n 0.017793f $X=-0.19 $Y=1.66 $X2=4.08 $Y2=1.1
cc_179 VPB N_VPWR_c_1003_n 0.0972054f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_180 VPB N_VPWR_c_1004_n 0.0684862f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_181 VPB N_VPWR_c_1005_n 0.0206041f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_182 VPB N_VPWR_c_1006_n 0.00613757f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_183 VPB N_VPWR_c_1007_n 0.00614127f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_184 VPB N_VPWR_c_1008_n 0.0106494f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_185 VPB N_VPWR_c_1009_n 0.00324402f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_186 VPB N_VPWR_c_993_n 0.12149f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_187 VPB N_A_323_392#_c_1112_n 0.0058341f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.885
cc_188 VPB N_A_323_392#_c_1104_n 0.00326003f $X=-0.19 $Y=1.66 $X2=0.535
+ $Y2=1.635
cc_189 VPB N_A_323_392#_c_1111_n 0.00151578f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_190 VPB N_A_323_392#_c_1115_n 0.00620953f $X=-0.19 $Y=1.66 $X2=4.24 $Y2=1.905
cc_191 VPB N_A_323_392#_c_1116_n 0.0102751f $X=-0.19 $Y=1.66 $X2=1.54 $Y2=1.925
cc_192 VPB N_A_416_118#_c_1238_n 0.00232832f $X=-0.19 $Y=1.66 $X2=0.535
+ $Y2=1.635
cc_193 VPB N_A_416_118#_c_1246_n 0.0151284f $X=-0.19 $Y=1.66 $X2=1.54 $Y2=1.085
cc_194 VPB N_A_416_118#_c_1247_n 0.00176541f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_195 VPB N_A_416_118#_c_1248_n 0.0062625f $X=-0.19 $Y=1.66 $X2=1.54 $Y2=1.925
cc_196 VPB N_A_416_118#_c_1249_n 0.0157427f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_197 VPB N_A_416_118#_c_1250_n 0.00477874f $X=-0.19 $Y=1.66 $X2=4.08 $Y2=1.1
cc_198 VPB N_A_416_118#_c_1244_n 0.0063041f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_199 VPB N_X_c_1360_n 0.00257348f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.91
cc_200 VPB N_X_c_1361_n 0.00262126f $X=-0.19 $Y=1.66 $X2=1.23 $Y2=2.815
cc_201 VPB N_X_c_1359_n 0.00139158f $X=-0.19 $Y=1.66 $X2=3.655 $Y2=2.99
cc_202 VPB X 0.00257348f $X=-0.19 $Y=1.66 $X2=1.54 $Y2=1.085
cc_203 N_A_74_294#_M1012_g N_A_c_318_n 0.004504f $X=0.495 $Y=0.91 $X2=-0.19
+ $Y2=-0.245
cc_204 N_A_74_294#_c_205_n N_A_c_318_n 0.0479296f $X=0.505 $Y=1.885 $X2=-0.19
+ $Y2=-0.245
cc_205 N_A_74_294#_c_206_n N_A_c_318_n 0.00243884f $X=0.535 $Y=1.635 $X2=-0.19
+ $Y2=-0.245
cc_206 N_A_74_294#_c_212_n N_A_c_318_n 0.012668f $X=1.065 $Y=1.925 $X2=-0.19
+ $Y2=-0.245
cc_207 N_A_74_294#_c_214_n N_A_c_318_n 0.0100974f $X=1.23 $Y=2.105 $X2=-0.19
+ $Y2=-0.245
cc_208 N_A_74_294#_c_216_n N_A_c_318_n 0.00336542f $X=1.395 $Y=2.99 $X2=-0.19
+ $Y2=-0.245
cc_209 N_A_74_294#_c_207_n N_A_c_318_n 0.00474324f $X=1.54 $Y=1.085 $X2=-0.19
+ $Y2=-0.245
cc_210 N_A_74_294#_c_219_n N_A_c_318_n 0.00373208f $X=1.54 $Y=1.925 $X2=-0.19
+ $Y2=-0.245
cc_211 N_A_74_294#_M1012_g N_A_c_319_n 0.019568f $X=0.495 $Y=0.91 $X2=0 $Y2=0
cc_212 N_A_74_294#_c_207_n N_A_c_319_n 0.0085975f $X=1.54 $Y=1.085 $X2=0 $Y2=0
cc_213 N_A_74_294#_M1012_g A 0.00262858f $X=0.495 $Y=0.91 $X2=0 $Y2=0
cc_214 N_A_74_294#_c_205_n A 6.96173e-19 $X=0.505 $Y=1.885 $X2=0 $Y2=0
cc_215 N_A_74_294#_c_206_n A 0.0126253f $X=0.535 $Y=1.635 $X2=0 $Y2=0
cc_216 N_A_74_294#_c_212_n A 0.0285285f $X=1.065 $Y=1.925 $X2=0 $Y2=0
cc_217 N_A_74_294#_c_207_n A 0.0370113f $X=1.54 $Y=1.085 $X2=0 $Y2=0
cc_218 N_A_74_294#_c_215_n N_A_397_320#_c_369_n 4.92401e-19 $X=3.655 $Y=2.99
+ $X2=0 $Y2=0
cc_219 N_A_74_294#_c_219_n N_A_397_320#_c_369_n 7.83506e-19 $X=1.54 $Y=1.925
+ $X2=0 $Y2=0
cc_220 N_A_74_294#_c_215_n N_A_397_320#_c_371_n 0.00115048f $X=3.655 $Y=2.99
+ $X2=0 $Y2=0
cc_221 N_A_74_294#_c_220_n N_A_397_320#_c_371_n 0.0057628f $X=3.74 $Y=2.07 $X2=0
+ $Y2=0
cc_222 N_A_74_294#_c_208_n N_A_397_320#_M1027_g 4.89753e-19 $X=3.99 $Y=1.905
+ $X2=0 $Y2=0
cc_223 N_A_74_294#_c_209_n N_A_397_320#_M1027_g 0.00119421f $X=4.24 $Y=1.1 $X2=0
+ $Y2=0
cc_224 N_A_74_294#_c_207_n N_A_397_320#_c_358_n 0.00512439f $X=1.54 $Y=1.085
+ $X2=0 $Y2=0
cc_225 N_A_74_294#_c_219_n N_A_397_320#_c_358_n 3.88319e-19 $X=1.54 $Y=1.925
+ $X2=0 $Y2=0
cc_226 N_A_74_294#_c_208_n N_A_397_320#_c_362_n 0.00794469f $X=3.99 $Y=1.905
+ $X2=0 $Y2=0
cc_227 N_A_74_294#_M1027_d N_A_397_320#_c_363_n 0.0066978f $X=3.77 $Y=0.625
+ $X2=0 $Y2=0
cc_228 N_A_74_294#_c_209_n N_A_397_320#_c_363_n 0.0252587f $X=4.24 $Y=1.1 $X2=0
+ $Y2=0
cc_229 N_A_74_294#_c_209_n N_A_397_320#_c_391_n 0.0209855f $X=4.24 $Y=1.1 $X2=0
+ $Y2=0
cc_230 N_A_74_294#_c_208_n N_A_397_320#_c_365_n 0.0929586f $X=3.99 $Y=1.905
+ $X2=0 $Y2=0
cc_231 N_A_74_294#_c_220_n N_A_397_320#_c_366_n 0.0250817f $X=3.74 $Y=2.07 $X2=0
+ $Y2=0
cc_232 N_A_74_294#_c_208_n N_A_397_320#_c_366_n 0.0225071f $X=3.99 $Y=1.905
+ $X2=0 $Y2=0
cc_233 N_A_74_294#_c_220_n N_A_397_320#_c_367_n 0.00830593f $X=3.74 $Y=2.07
+ $X2=0 $Y2=0
cc_234 N_A_74_294#_c_208_n N_A_397_320#_c_367_n 0.00135436f $X=3.99 $Y=1.905
+ $X2=0 $Y2=0
cc_235 N_A_74_294#_c_214_n N_B_c_483_n 0.0136841f $X=1.23 $Y=2.105 $X2=-0.19
+ $Y2=-0.245
cc_236 N_A_74_294#_c_207_n N_B_c_483_n 0.00448607f $X=1.54 $Y=1.085 $X2=-0.19
+ $Y2=-0.245
cc_237 N_A_74_294#_c_219_n N_B_c_483_n 0.0124313f $X=1.54 $Y=1.925 $X2=-0.19
+ $Y2=-0.245
cc_238 N_A_74_294#_c_215_n N_B_c_484_n 0.015877f $X=3.655 $Y=2.99 $X2=0 $Y2=0
cc_239 N_A_74_294#_c_207_n N_B_M1019_g 0.00131726f $X=1.54 $Y=1.085 $X2=0 $Y2=0
cc_240 N_A_74_294#_c_215_n N_B_c_486_n 0.0148201f $X=3.655 $Y=2.99 $X2=0 $Y2=0
cc_241 N_A_74_294#_c_215_n N_B_c_488_n 0.0205994f $X=3.655 $Y=2.99 $X2=0 $Y2=0
cc_242 N_A_74_294#_c_220_n N_B_c_488_n 0.00680497f $X=3.74 $Y=2.07 $X2=0 $Y2=0
cc_243 N_A_74_294#_c_215_n N_B_c_475_n 0.00532519f $X=3.655 $Y=2.99 $X2=0 $Y2=0
cc_244 N_A_74_294#_c_218_n N_B_c_475_n 0.00389649f $X=3.74 $Y=2.905 $X2=0 $Y2=0
cc_245 N_A_74_294#_c_220_n N_B_c_475_n 0.0331852f $X=3.74 $Y=2.07 $X2=0 $Y2=0
cc_246 N_A_74_294#_c_208_n N_B_c_475_n 0.00874935f $X=3.99 $Y=1.905 $X2=0 $Y2=0
cc_247 N_A_74_294#_c_208_n N_B_c_476_n 0.00323245f $X=3.99 $Y=1.905 $X2=0 $Y2=0
cc_248 N_A_74_294#_c_209_n N_B_c_476_n 0.00936145f $X=4.24 $Y=1.1 $X2=0 $Y2=0
cc_249 N_A_74_294#_c_214_n N_B_c_491_n 8.31485e-19 $X=1.23 $Y=2.105 $X2=0 $Y2=0
cc_250 N_A_74_294#_c_215_n N_B_c_491_n 0.0177219f $X=3.655 $Y=2.99 $X2=0 $Y2=0
cc_251 N_A_74_294#_c_208_n N_B_c_481_n 0.00487217f $X=3.99 $Y=1.905 $X2=0 $Y2=0
cc_252 N_A_74_294#_c_209_n N_B_c_481_n 2.18267e-19 $X=4.24 $Y=1.1 $X2=0 $Y2=0
cc_253 N_A_74_294#_M1012_g N_A_27_118#_c_909_n 0.00136219f $X=0.495 $Y=0.91
+ $X2=0 $Y2=0
cc_254 N_A_74_294#_M1012_g N_A_27_118#_c_910_n 0.00701795f $X=0.495 $Y=0.91
+ $X2=0 $Y2=0
cc_255 N_A_74_294#_c_205_n N_A_27_118#_c_918_n 0.00472178f $X=0.505 $Y=1.885
+ $X2=0 $Y2=0
cc_256 N_A_74_294#_M1025_d N_A_27_118#_c_911_n 0.0172433f $X=1.24 $Y=0.59 $X2=0
+ $Y2=0
cc_257 N_A_74_294#_M1012_g N_A_27_118#_c_911_n 0.0123984f $X=0.495 $Y=0.91 $X2=0
+ $Y2=0
cc_258 N_A_74_294#_c_207_n N_A_27_118#_c_911_n 0.0136682f $X=1.54 $Y=1.085 $X2=0
+ $Y2=0
cc_259 N_A_74_294#_M1025_d N_A_27_118#_c_912_n 0.00571414f $X=1.24 $Y=0.59 $X2=0
+ $Y2=0
cc_260 N_A_74_294#_c_207_n N_A_27_118#_c_912_n 0.0368226f $X=1.54 $Y=1.085 $X2=0
+ $Y2=0
cc_261 N_A_74_294#_c_207_n N_A_27_118#_c_913_n 0.00809439f $X=1.54 $Y=1.085
+ $X2=0 $Y2=0
cc_262 N_A_74_294#_c_219_n N_A_27_118#_c_913_n 0.00501248f $X=1.54 $Y=1.925
+ $X2=0 $Y2=0
cc_263 N_A_74_294#_c_207_n N_A_27_118#_c_914_n 0.0141893f $X=1.54 $Y=1.085 $X2=0
+ $Y2=0
cc_264 N_A_74_294#_M1012_g N_A_27_118#_c_916_n 0.0045716f $X=0.495 $Y=0.91 $X2=0
+ $Y2=0
cc_265 N_A_74_294#_c_205_n N_A_27_118#_c_916_n 0.00209596f $X=0.505 $Y=1.885
+ $X2=0 $Y2=0
cc_266 N_A_74_294#_c_206_n N_A_27_118#_c_916_n 0.00121581f $X=0.535 $Y=1.635
+ $X2=0 $Y2=0
cc_267 N_A_74_294#_M1012_g N_A_27_118#_c_917_n 0.00407149f $X=0.495 $Y=0.91
+ $X2=0 $Y2=0
cc_268 N_A_74_294#_c_205_n N_A_27_118#_c_917_n 0.0145593f $X=0.505 $Y=1.885
+ $X2=0 $Y2=0
cc_269 N_A_74_294#_c_206_n N_A_27_118#_c_917_n 0.0273872f $X=0.535 $Y=1.635
+ $X2=0 $Y2=0
cc_270 N_A_74_294#_c_213_n N_A_27_118#_c_917_n 0.0117066f $X=0.7 $Y=1.925 $X2=0
+ $Y2=0
cc_271 N_A_74_294#_c_212_n N_VPWR_M1008_d 0.00182839f $X=1.065 $Y=1.925
+ $X2=-0.19 $Y2=-0.245
cc_272 N_A_74_294#_c_213_n N_VPWR_M1008_d 6.813e-19 $X=0.7 $Y=1.925 $X2=-0.19
+ $Y2=-0.245
cc_273 N_A_74_294#_c_205_n N_VPWR_c_994_n 0.0166225f $X=0.505 $Y=1.885 $X2=0
+ $Y2=0
cc_274 N_A_74_294#_c_212_n N_VPWR_c_994_n 0.0140386f $X=1.065 $Y=1.925 $X2=0
+ $Y2=0
cc_275 N_A_74_294#_c_213_n N_VPWR_c_994_n 0.0067086f $X=0.7 $Y=1.925 $X2=0 $Y2=0
cc_276 N_A_74_294#_c_216_n N_VPWR_c_994_n 0.0119239f $X=1.395 $Y=2.99 $X2=0
+ $Y2=0
cc_277 N_A_74_294#_c_205_n N_VPWR_c_1002_n 0.00413917f $X=0.505 $Y=1.885 $X2=0
+ $Y2=0
cc_278 N_A_74_294#_c_215_n N_VPWR_c_1003_n 0.156034f $X=3.655 $Y=2.99 $X2=0
+ $Y2=0
cc_279 N_A_74_294#_c_216_n N_VPWR_c_1003_n 0.0236039f $X=1.395 $Y=2.99 $X2=0
+ $Y2=0
cc_280 N_A_74_294#_c_220_n N_VPWR_c_1003_n 0.0113172f $X=3.74 $Y=2.07 $X2=0
+ $Y2=0
cc_281 N_A_74_294#_c_205_n N_VPWR_c_993_n 0.00821221f $X=0.505 $Y=1.885 $X2=0
+ $Y2=0
cc_282 N_A_74_294#_c_215_n N_VPWR_c_993_n 0.0817155f $X=3.655 $Y=2.99 $X2=0
+ $Y2=0
cc_283 N_A_74_294#_c_216_n N_VPWR_c_993_n 0.012761f $X=1.395 $Y=2.99 $X2=0 $Y2=0
cc_284 N_A_74_294#_c_220_n N_VPWR_c_993_n 0.0137388f $X=3.74 $Y=2.07 $X2=0 $Y2=0
cc_285 N_A_74_294#_c_214_n N_A_323_392#_c_1117_n 0.0121155f $X=1.23 $Y=2.105
+ $X2=0 $Y2=0
cc_286 N_A_74_294#_c_215_n N_A_323_392#_c_1117_n 0.0228238f $X=3.655 $Y=2.99
+ $X2=0 $Y2=0
cc_287 N_A_74_294#_c_214_n N_A_323_392#_c_1119_n 0.0258437f $X=1.23 $Y=2.105
+ $X2=0 $Y2=0
cc_288 N_A_74_294#_c_219_n N_A_323_392#_c_1119_n 0.00100766f $X=1.54 $Y=1.925
+ $X2=0 $Y2=0
cc_289 N_A_74_294#_M1002_d N_A_323_392#_c_1112_n 0.00343339f $X=3.28 $Y=1.895
+ $X2=0 $Y2=0
cc_290 N_A_74_294#_c_215_n N_A_323_392#_c_1112_n 0.10542f $X=3.655 $Y=2.99 $X2=0
+ $Y2=0
cc_291 N_A_74_294#_c_220_n N_A_323_392#_c_1112_n 0.0152397f $X=3.74 $Y=2.07
+ $X2=0 $Y2=0
cc_292 N_A_74_294#_M1002_d N_A_323_392#_c_1104_n 0.010352f $X=3.28 $Y=1.895
+ $X2=0 $Y2=0
cc_293 N_A_74_294#_c_220_n N_A_323_392#_c_1104_n 0.0517893f $X=3.74 $Y=2.07
+ $X2=0 $Y2=0
cc_294 N_A_74_294#_c_208_n N_A_323_392#_c_1104_n 0.00487615f $X=3.99 $Y=1.905
+ $X2=0 $Y2=0
cc_295 N_A_74_294#_M1002_d N_A_416_118#_c_1246_n 0.0102262f $X=3.28 $Y=1.895
+ $X2=0 $Y2=0
cc_296 N_A_74_294#_c_220_n N_A_416_118#_c_1246_n 0.0693533f $X=3.74 $Y=2.07
+ $X2=0 $Y2=0
cc_297 N_A_74_294#_M1012_g N_VGND_c_1427_n 0.00331146f $X=0.495 $Y=0.91 $X2=0
+ $Y2=0
cc_298 N_A_74_294#_M1012_g N_VGND_c_1433_n 0.00479212f $X=0.495 $Y=0.91 $X2=0
+ $Y2=0
cc_299 N_A_c_318_n N_B_c_483_n 0.014046f $X=1.005 $Y=1.885 $X2=-0.19 $Y2=-0.245
cc_300 N_A_c_319_n N_B_M1019_g 0.0104543f $X=1.165 $Y=1.34 $X2=0 $Y2=0
cc_301 N_A_c_318_n N_B_c_491_n 0.00535642f $X=1.005 $Y=1.885 $X2=0 $Y2=0
cc_302 N_A_c_319_n N_A_27_118#_c_910_n 0.00185091f $X=1.165 $Y=1.34 $X2=0 $Y2=0
cc_303 N_A_c_318_n N_A_27_118#_c_911_n 6.365e-19 $X=1.005 $Y=1.885 $X2=0 $Y2=0
cc_304 N_A_c_319_n N_A_27_118#_c_911_n 0.0145958f $X=1.165 $Y=1.34 $X2=0 $Y2=0
cc_305 A N_A_27_118#_c_911_n 0.0101016f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_306 N_A_c_319_n N_A_27_118#_c_912_n 0.00287039f $X=1.165 $Y=1.34 $X2=0 $Y2=0
cc_307 A N_A_27_118#_c_916_n 0.00256975f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_308 A N_A_27_118#_c_917_n 0.00472684f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_309 N_A_c_318_n N_VPWR_c_994_n 0.00554997f $X=1.005 $Y=1.885 $X2=0 $Y2=0
cc_310 N_A_c_318_n N_VPWR_c_1003_n 0.0044313f $X=1.005 $Y=1.885 $X2=0 $Y2=0
cc_311 N_A_c_318_n N_VPWR_c_993_n 0.00853879f $X=1.005 $Y=1.885 $X2=0 $Y2=0
cc_312 A N_VGND_M1012_d 0.00281085f $X=1.115 $Y=1.21 $X2=-0.19 $Y2=-0.245
cc_313 N_A_c_319_n N_VGND_c_1425_n 0.0033127f $X=1.165 $Y=1.34 $X2=0 $Y2=0
cc_314 N_A_c_319_n N_VGND_c_1433_n 0.00479212f $X=1.165 $Y=1.34 $X2=0 $Y2=0
cc_315 N_A_397_320#_c_369_n N_B_c_483_n 0.0133552f $X=2.075 $Y=1.885 $X2=-0.19
+ $Y2=-0.245
cc_316 N_A_397_320#_c_358_n N_B_c_483_n 0.0016228f $X=2.075 $Y=1.675 $X2=-0.19
+ $Y2=-0.245
cc_317 N_A_397_320#_c_369_n N_B_c_484_n 0.004527f $X=2.075 $Y=1.885 $X2=0 $Y2=0
cc_318 N_A_397_320#_M1022_g N_B_M1019_g 0.0108207f $X=2.505 $Y=1.02 $X2=0 $Y2=0
cc_319 N_A_397_320#_c_358_n N_B_M1019_g 0.00516515f $X=2.075 $Y=1.675 $X2=0
+ $Y2=0
cc_320 N_A_397_320#_M1022_g N_B_c_471_n 0.00325348f $X=2.505 $Y=1.02 $X2=0 $Y2=0
cc_321 N_A_397_320#_c_371_n N_B_c_485_n 0.00240207f $X=3.205 $Y=1.82 $X2=0 $Y2=0
cc_322 N_A_397_320#_c_369_n N_B_c_487_n 0.0143735f $X=2.075 $Y=1.885 $X2=0 $Y2=0
cc_323 N_A_397_320#_c_371_n N_B_c_487_n 0.0202957f $X=3.205 $Y=1.82 $X2=0 $Y2=0
cc_324 N_A_397_320#_c_360_n N_B_c_487_n 0.00938742f $X=3.115 $Y=1.71 $X2=0 $Y2=0
cc_325 N_A_397_320#_c_371_n N_B_c_488_n 0.00882199f $X=3.205 $Y=1.82 $X2=0 $Y2=0
cc_326 N_A_397_320#_M1022_g N_B_M1014_g 0.0110201f $X=2.505 $Y=1.02 $X2=0 $Y2=0
cc_327 N_A_397_320#_M1027_g N_B_M1014_g 0.0156701f $X=3.695 $Y=0.945 $X2=0 $Y2=0
cc_328 N_A_397_320#_c_360_n N_B_M1014_g 0.00886845f $X=3.115 $Y=1.71 $X2=0 $Y2=0
cc_329 N_A_397_320#_M1027_g N_B_c_474_n 0.00737859f $X=3.695 $Y=0.945 $X2=0
+ $Y2=0
cc_330 N_A_397_320#_c_365_n N_B_c_475_n 0.0137878f $X=4.62 $Y=1.985 $X2=0 $Y2=0
cc_331 N_A_397_320#_M1027_g N_B_c_476_n 0.0172653f $X=3.695 $Y=0.945 $X2=0 $Y2=0
cc_332 N_A_397_320#_c_362_n N_B_c_476_n 4.02697e-19 $X=3.74 $Y=1.435 $X2=0 $Y2=0
cc_333 N_A_397_320#_c_363_n N_B_c_476_n 0.0149863f $X=4.535 $Y=0.68 $X2=0 $Y2=0
cc_334 N_A_397_320#_c_391_n N_B_c_476_n 0.00774765f $X=4.655 $Y=0.86 $X2=0 $Y2=0
cc_335 N_A_397_320#_c_363_n N_B_c_477_n 0.00220975f $X=4.535 $Y=0.68 $X2=0 $Y2=0
cc_336 N_A_397_320#_c_365_n N_B_c_477_n 0.0140311f $X=4.62 $Y=1.985 $X2=0 $Y2=0
cc_337 N_A_397_320#_c_368_n N_B_c_477_n 0.00142955f $X=4.637 $Y=1.13 $X2=0 $Y2=0
cc_338 N_A_397_320#_c_365_n N_B_c_478_n 0.0125433f $X=4.62 $Y=1.985 $X2=0 $Y2=0
cc_339 N_A_397_320#_c_365_n N_B_c_479_n 0.00147807f $X=4.62 $Y=1.985 $X2=0 $Y2=0
cc_340 N_A_397_320#_c_368_n N_B_c_479_n 7.77673e-19 $X=4.637 $Y=1.13 $X2=0 $Y2=0
cc_341 N_A_397_320#_c_366_n N_B_c_481_n 3.19844e-19 $X=3.82 $Y=1.57 $X2=0 $Y2=0
cc_342 N_A_397_320#_c_367_n N_B_c_481_n 0.0167206f $X=3.82 $Y=1.57 $X2=0 $Y2=0
cc_343 N_A_397_320#_c_365_n B 0.0235521f $X=4.62 $Y=1.985 $X2=0 $Y2=0
cc_344 N_A_397_320#_M1022_g N_A_27_118#_c_912_n 0.00144183f $X=2.505 $Y=1.02
+ $X2=0 $Y2=0
cc_345 N_A_397_320#_c_369_n N_A_27_118#_c_913_n 0.00975662f $X=2.075 $Y=1.885
+ $X2=0 $Y2=0
cc_346 N_A_397_320#_c_354_n N_A_27_118#_c_913_n 0.0153899f $X=2.43 $Y=1.675
+ $X2=0 $Y2=0
cc_347 N_A_397_320#_M1022_g N_A_27_118#_c_913_n 2.63712e-19 $X=2.505 $Y=1.02
+ $X2=0 $Y2=0
cc_348 N_A_397_320#_c_358_n N_A_27_118#_c_913_n 0.00893486f $X=2.075 $Y=1.675
+ $X2=0 $Y2=0
cc_349 N_A_397_320#_c_354_n N_A_27_118#_c_914_n 0.00185617f $X=2.43 $Y=1.675
+ $X2=0 $Y2=0
cc_350 N_A_397_320#_M1022_g N_A_27_118#_c_914_n 0.018906f $X=2.505 $Y=1.02 $X2=0
+ $Y2=0
cc_351 N_A_397_320#_c_358_n N_A_27_118#_c_914_n 0.00992456f $X=2.075 $Y=1.675
+ $X2=0 $Y2=0
cc_352 N_A_397_320#_c_360_n N_A_27_118#_c_914_n 0.00337236f $X=3.115 $Y=1.71
+ $X2=0 $Y2=0
cc_353 N_A_397_320#_M1022_g N_A_27_118#_c_915_n 0.011728f $X=2.505 $Y=1.02 $X2=0
+ $Y2=0
cc_354 N_A_397_320#_c_365_n N_VPWR_c_995_n 0.0743839f $X=4.62 $Y=1.985 $X2=0
+ $Y2=0
cc_355 N_A_397_320#_c_365_n N_VPWR_c_1003_n 0.00749631f $X=4.62 $Y=1.985 $X2=0
+ $Y2=0
cc_356 N_A_397_320#_c_365_n N_VPWR_c_993_n 0.0062048f $X=4.62 $Y=1.985 $X2=0
+ $Y2=0
cc_357 N_A_397_320#_c_369_n N_A_323_392#_c_1119_n 0.00667392f $X=2.075 $Y=1.885
+ $X2=0 $Y2=0
cc_358 N_A_397_320#_c_369_n N_A_323_392#_c_1112_n 0.0143127f $X=2.075 $Y=1.885
+ $X2=0 $Y2=0
cc_359 N_A_397_320#_c_371_n N_A_323_392#_c_1112_n 0.0122153f $X=3.205 $Y=1.82
+ $X2=0 $Y2=0
cc_360 N_A_397_320#_c_371_n N_A_323_392#_c_1104_n 0.0146226f $X=3.205 $Y=1.82
+ $X2=0 $Y2=0
cc_361 N_A_397_320#_c_356_n N_A_323_392#_c_1104_n 0.0147637f $X=3.62 $Y=1.675
+ $X2=0 $Y2=0
cc_362 N_A_397_320#_M1027_g N_A_323_392#_c_1104_n 0.0137034f $X=3.695 $Y=0.945
+ $X2=0 $Y2=0
cc_363 N_A_397_320#_c_361_n N_A_323_392#_c_1104_n 0.00166247f $X=3.295 $Y=1.71
+ $X2=0 $Y2=0
cc_364 N_A_397_320#_c_362_n N_A_323_392#_c_1104_n 0.0471932f $X=3.74 $Y=1.435
+ $X2=0 $Y2=0
cc_365 N_A_397_320#_c_364_n N_A_323_392#_c_1104_n 0.0133618f $X=3.825 $Y=0.68
+ $X2=0 $Y2=0
cc_366 N_A_397_320#_c_366_n N_A_323_392#_c_1104_n 0.0220053f $X=3.82 $Y=1.57
+ $X2=0 $Y2=0
cc_367 N_A_397_320#_M1026_s N_A_323_392#_c_1105_n 0.00237105f $X=4.515 $Y=0.37
+ $X2=0 $Y2=0
cc_368 N_A_397_320#_M1027_g N_A_323_392#_c_1105_n 0.00174767f $X=3.695 $Y=0.945
+ $X2=0 $Y2=0
cc_369 N_A_397_320#_c_363_n N_A_323_392#_c_1105_n 0.0645371f $X=4.535 $Y=0.68
+ $X2=0 $Y2=0
cc_370 N_A_397_320#_c_364_n N_A_323_392#_c_1105_n 0.0129683f $X=3.825 $Y=0.68
+ $X2=0 $Y2=0
cc_371 N_A_397_320#_M1022_g N_A_416_118#_c_1235_n 0.00407278f $X=2.505 $Y=1.02
+ $X2=0 $Y2=0
cc_372 N_A_397_320#_M1022_g N_A_416_118#_c_1236_n 0.00380542f $X=2.505 $Y=1.02
+ $X2=0 $Y2=0
cc_373 N_A_397_320#_M1022_g N_A_416_118#_c_1238_n 0.0014728f $X=2.505 $Y=1.02
+ $X2=0 $Y2=0
cc_374 N_A_397_320#_c_371_n N_A_416_118#_c_1238_n 0.00152837f $X=3.205 $Y=1.82
+ $X2=0 $Y2=0
cc_375 N_A_397_320#_c_360_n N_A_416_118#_c_1238_n 0.0104838f $X=3.115 $Y=1.71
+ $X2=0 $Y2=0
cc_376 N_A_397_320#_c_361_n N_A_416_118#_c_1238_n 0.00501713f $X=3.295 $Y=1.71
+ $X2=0 $Y2=0
cc_377 N_A_397_320#_M1003_s N_A_416_118#_c_1246_n 0.0083057f $X=4.475 $Y=1.84
+ $X2=0 $Y2=0
cc_378 N_A_397_320#_c_371_n N_A_416_118#_c_1246_n 0.00828579f $X=3.205 $Y=1.82
+ $X2=0 $Y2=0
cc_379 N_A_397_320#_c_356_n N_A_416_118#_c_1246_n 0.00475242f $X=3.62 $Y=1.675
+ $X2=0 $Y2=0
cc_380 N_A_397_320#_c_361_n N_A_416_118#_c_1246_n 3.42966e-19 $X=3.295 $Y=1.71
+ $X2=0 $Y2=0
cc_381 N_A_397_320#_c_365_n N_A_416_118#_c_1246_n 0.0204259f $X=4.62 $Y=1.985
+ $X2=0 $Y2=0
cc_382 N_A_397_320#_c_366_n N_A_416_118#_c_1246_n 0.00212633f $X=3.82 $Y=1.57
+ $X2=0 $Y2=0
cc_383 N_A_397_320#_c_359_n N_A_416_118#_c_1247_n 0.00177559f $X=2.505 $Y=1.675
+ $X2=0 $Y2=0
cc_384 N_A_397_320#_c_369_n N_A_416_118#_c_1250_n 5.26654e-19 $X=2.075 $Y=1.885
+ $X2=0 $Y2=0
cc_385 N_A_397_320#_c_371_n N_A_416_118#_c_1250_n 0.00766496f $X=3.205 $Y=1.82
+ $X2=0 $Y2=0
cc_386 N_A_397_320#_c_359_n N_A_416_118#_c_1250_n 0.0108639f $X=2.505 $Y=1.675
+ $X2=0 $Y2=0
cc_387 N_A_397_320#_c_360_n N_A_416_118#_c_1250_n 8.16991e-19 $X=3.115 $Y=1.71
+ $X2=0 $Y2=0
cc_388 N_B_c_478_n N_A_1155_284#_c_606_n 0.00220621f $X=4.845 $Y=1.765 $X2=0
+ $Y2=0
cc_389 N_B_M1019_g N_A_27_118#_c_911_n 0.00615086f $X=2.005 $Y=0.91 $X2=0 $Y2=0
cc_390 N_B_M1019_g N_A_27_118#_c_912_n 0.0164031f $X=2.005 $Y=0.91 $X2=0 $Y2=0
cc_391 N_B_c_483_n N_A_27_118#_c_913_n 7.04891e-19 $X=1.54 $Y=2.875 $X2=0 $Y2=0
cc_392 N_B_c_487_n N_A_27_118#_c_913_n 0.00149913f $X=2.67 $Y=2.805 $X2=0 $Y2=0
cc_393 N_B_M1019_g N_A_27_118#_c_914_n 0.00361406f $X=2.005 $Y=0.91 $X2=0 $Y2=0
cc_394 N_B_c_487_n N_A_27_118#_c_914_n 2.36236e-19 $X=2.67 $Y=2.805 $X2=0 $Y2=0
cc_395 N_B_M1019_g N_A_27_118#_c_915_n 4.4652e-19 $X=2.005 $Y=0.91 $X2=0 $Y2=0
cc_396 N_B_M1014_g N_A_27_118#_c_915_n 0.00190771f $X=3.105 $Y=0.91 $X2=0 $Y2=0
cc_397 N_B_c_491_n N_VPWR_c_994_n 0.00217365f $X=1.54 $Y=3.15 $X2=0 $Y2=0
cc_398 N_B_c_488_n N_VPWR_c_995_n 0.00232909f $X=4.25 $Y=3.15 $X2=0 $Y2=0
cc_399 N_B_c_475_n N_VPWR_c_995_n 8.68538e-19 $X=4.325 $Y=3.075 $X2=0 $Y2=0
cc_400 N_B_c_478_n N_VPWR_c_995_n 0.0210003f $X=4.845 $Y=1.765 $X2=0 $Y2=0
cc_401 B N_VPWR_c_995_n 0.0175404f $X=4.955 $Y=1.21 $X2=0 $Y2=0
cc_402 N_B_c_478_n N_VPWR_c_1003_n 0.00413917f $X=4.845 $Y=1.765 $X2=0 $Y2=0
cc_403 N_B_c_491_n N_VPWR_c_1003_n 0.0655287f $X=1.54 $Y=3.15 $X2=0 $Y2=0
cc_404 N_B_c_484_n N_VPWR_c_993_n 0.0223434f $X=2.58 $Y=3.15 $X2=0 $Y2=0
cc_405 N_B_c_488_n N_VPWR_c_993_n 0.0451072f $X=4.25 $Y=3.15 $X2=0 $Y2=0
cc_406 N_B_c_478_n N_VPWR_c_993_n 0.0081836f $X=4.845 $Y=1.765 $X2=0 $Y2=0
cc_407 N_B_c_491_n N_VPWR_c_993_n 0.00670671f $X=1.54 $Y=3.15 $X2=0 $Y2=0
cc_408 N_B_c_492_n N_VPWR_c_993_n 0.00441537f $X=2.67 $Y=3.15 $X2=0 $Y2=0
cc_409 N_B_c_483_n N_A_323_392#_c_1117_n 0.00196216f $X=1.54 $Y=2.875 $X2=0
+ $Y2=0
cc_410 N_B_c_483_n N_A_323_392#_c_1119_n 0.00418619f $X=1.54 $Y=2.875 $X2=0
+ $Y2=0
cc_411 N_B_c_485_n N_A_323_392#_c_1112_n 7.95665e-19 $X=2.67 $Y=2.895 $X2=0
+ $Y2=0
cc_412 N_B_c_487_n N_A_323_392#_c_1112_n 0.0115759f $X=2.67 $Y=2.805 $X2=0 $Y2=0
cc_413 N_B_M1014_g N_A_323_392#_c_1104_n 0.0083722f $X=3.105 $Y=0.91 $X2=0 $Y2=0
cc_414 N_B_c_474_n N_A_323_392#_c_1105_n 0.0143527f $X=4.29 $Y=0.18 $X2=0 $Y2=0
cc_415 N_B_c_476_n N_A_323_392#_c_1105_n 0.0121287f $X=4.365 $Y=1.4 $X2=0 $Y2=0
cc_416 N_B_c_479_n N_A_323_392#_c_1105_n 0.0134686f $X=4.87 $Y=1.22 $X2=0 $Y2=0
cc_417 N_B_M1014_g N_A_323_392#_c_1106_n 0.00724099f $X=3.105 $Y=0.91 $X2=0
+ $Y2=0
cc_418 N_B_c_474_n N_A_323_392#_c_1106_n 0.00420304f $X=4.29 $Y=0.18 $X2=0 $Y2=0
cc_419 N_B_c_476_n N_A_323_392#_c_1151_n 9.49236e-19 $X=4.365 $Y=1.4 $X2=0 $Y2=0
cc_420 N_B_c_479_n N_A_323_392#_c_1151_n 0.0112116f $X=4.87 $Y=1.22 $X2=0 $Y2=0
cc_421 N_B_c_478_n N_A_323_392#_c_1107_n 9.5528e-19 $X=4.845 $Y=1.765 $X2=0
+ $Y2=0
cc_422 B N_A_323_392#_c_1107_n 0.0100791f $X=4.955 $Y=1.21 $X2=0 $Y2=0
cc_423 N_B_c_478_n N_A_323_392#_c_1155_n 7.4925e-19 $X=4.845 $Y=1.765 $X2=0
+ $Y2=0
cc_424 N_B_c_479_n N_A_323_392#_c_1155_n 0.00655142f $X=4.87 $Y=1.22 $X2=0 $Y2=0
cc_425 B N_A_323_392#_c_1155_n 0.00963599f $X=4.955 $Y=1.21 $X2=0 $Y2=0
cc_426 N_B_M1014_g N_A_416_118#_c_1235_n 3.48096e-19 $X=3.105 $Y=0.91 $X2=0
+ $Y2=0
cc_427 N_B_c_471_n N_A_416_118#_c_1236_n 0.00964413f $X=3.03 $Y=0.18 $X2=0 $Y2=0
cc_428 N_B_M1014_g N_A_416_118#_c_1236_n 0.00881029f $X=3.105 $Y=0.91 $X2=0
+ $Y2=0
cc_429 N_B_M1019_g N_A_416_118#_c_1237_n 0.00628461f $X=2.005 $Y=0.91 $X2=0
+ $Y2=0
cc_430 N_B_c_471_n N_A_416_118#_c_1237_n 0.00478134f $X=3.03 $Y=0.18 $X2=0 $Y2=0
cc_431 N_B_M1014_g N_A_416_118#_c_1238_n 0.0196551f $X=3.105 $Y=0.91 $X2=0 $Y2=0
cc_432 N_B_c_478_n N_A_416_118#_c_1240_n 0.00173686f $X=4.845 $Y=1.765 $X2=0
+ $Y2=0
cc_433 N_B_c_479_n N_A_416_118#_c_1240_n 0.00193183f $X=4.87 $Y=1.22 $X2=0 $Y2=0
cc_434 B N_A_416_118#_c_1240_n 0.00853672f $X=4.955 $Y=1.21 $X2=0 $Y2=0
cc_435 N_B_c_475_n N_A_416_118#_c_1246_n 0.00733464f $X=4.325 $Y=3.075 $X2=0
+ $Y2=0
cc_436 N_B_c_477_n N_A_416_118#_c_1246_n 8.43864e-19 $X=4.755 $Y=1.475 $X2=0
+ $Y2=0
cc_437 N_B_c_478_n N_A_416_118#_c_1246_n 0.0115063f $X=4.845 $Y=1.765 $X2=0
+ $Y2=0
cc_438 B N_A_416_118#_c_1246_n 0.00191389f $X=4.955 $Y=1.21 $X2=0 $Y2=0
cc_439 N_B_c_478_n N_A_416_118#_c_1249_n 0.00127768f $X=4.845 $Y=1.765 $X2=0
+ $Y2=0
cc_440 N_B_c_487_n N_A_416_118#_c_1250_n 0.0186036f $X=2.67 $Y=2.805 $X2=0 $Y2=0
cc_441 N_B_c_478_n N_A_416_118#_c_1244_n 0.0112754f $X=4.845 $Y=1.765 $X2=0
+ $Y2=0
cc_442 B N_A_416_118#_c_1244_n 0.0175916f $X=4.955 $Y=1.21 $X2=0 $Y2=0
cc_443 N_B_c_479_n N_VGND_c_1419_n 0.00229971f $X=4.87 $Y=1.22 $X2=0 $Y2=0
cc_444 N_B_c_472_n N_VGND_c_1425_n 0.0612704f $X=2.08 $Y=0.18 $X2=0 $Y2=0
cc_445 N_B_c_479_n N_VGND_c_1425_n 0.00278237f $X=4.87 $Y=1.22 $X2=0 $Y2=0
cc_446 N_B_c_471_n N_VGND_c_1433_n 0.0253825f $X=3.03 $Y=0.18 $X2=0 $Y2=0
cc_447 N_B_c_472_n N_VGND_c_1433_n 0.0104168f $X=2.08 $Y=0.18 $X2=0 $Y2=0
cc_448 N_B_c_474_n N_VGND_c_1433_n 0.0367763f $X=4.29 $Y=0.18 $X2=0 $Y2=0
cc_449 N_B_c_479_n N_VGND_c_1433_n 0.00359127f $X=4.87 $Y=1.22 $X2=0 $Y2=0
cc_450 N_B_c_480_n N_VGND_c_1433_n 0.00515892f $X=3.105 $Y=0.18 $X2=0 $Y2=0
cc_451 N_A_1155_284#_c_606_n N_C_c_692_n 0.0210593f $X=6.015 $Y=1.865 $X2=-0.19
+ $Y2=-0.245
cc_452 N_A_1155_284#_c_612_n N_C_c_692_n 0.00260005f $X=6.05 $Y=2.905 $X2=-0.19
+ $Y2=-0.245
cc_453 N_A_1155_284#_c_613_n N_C_c_692_n 0.00875865f $X=7.33 $Y=2.99 $X2=-0.19
+ $Y2=-0.245
cc_454 N_A_1155_284#_c_608_n N_C_c_692_n 2.87763e-19 $X=6.05 $Y=1.605 $X2=-0.19
+ $Y2=-0.245
cc_455 N_A_1155_284#_c_617_n N_C_c_692_n 0.00434687f $X=7.495 $Y=2.455 $X2=-0.19
+ $Y2=-0.245
cc_456 N_A_1155_284#_M1016_g N_C_M1021_g 0.0142541f $X=6.09 $Y=0.935 $X2=0 $Y2=0
cc_457 N_A_1155_284#_c_609_n N_C_c_694_n 0.00289177f $X=7.54 $Y=2.29 $X2=0 $Y2=0
cc_458 N_A_1155_284#_c_609_n N_C_c_695_n 0.0149489f $X=7.54 $Y=2.29 $X2=0 $Y2=0
cc_459 N_A_1155_284#_c_610_n N_C_c_695_n 0.0124419f $X=7.985 $Y=0.58 $X2=0 $Y2=0
cc_460 N_A_1155_284#_c_617_n N_C_c_702_n 0.00510622f $X=7.495 $Y=2.455 $X2=0
+ $Y2=0
cc_461 N_A_1155_284#_c_609_n N_C_c_702_n 0.0110404f $X=7.54 $Y=2.29 $X2=0 $Y2=0
cc_462 N_A_1155_284#_c_615_n N_C_c_703_n 0.00249724f $X=7.415 $Y=2.905 $X2=0
+ $Y2=0
cc_463 N_A_1155_284#_c_617_n N_C_c_703_n 0.00987831f $X=7.495 $Y=2.455 $X2=0
+ $Y2=0
cc_464 N_A_1155_284#_c_609_n N_C_c_703_n 0.00899104f $X=7.54 $Y=2.29 $X2=0 $Y2=0
cc_465 N_A_1155_284#_c_609_n N_C_c_697_n 0.00174057f $X=7.54 $Y=2.29 $X2=0 $Y2=0
cc_466 N_A_1155_284#_c_610_n N_C_c_697_n 0.00422628f $X=7.985 $Y=0.58 $X2=0
+ $Y2=0
cc_467 N_A_1155_284#_c_617_n N_C_c_699_n 4.40372e-19 $X=7.495 $Y=2.455 $X2=0
+ $Y2=0
cc_468 N_A_1155_284#_c_606_n N_A_1218_388#_c_774_n 6.14056e-19 $X=6.015 $Y=1.865
+ $X2=0 $Y2=0
cc_469 N_A_1155_284#_M1016_g N_A_1218_388#_c_774_n 0.00664534f $X=6.09 $Y=0.935
+ $X2=0 $Y2=0
cc_470 N_A_1155_284#_c_612_n N_A_1218_388#_c_774_n 0.00797895f $X=6.05 $Y=2.905
+ $X2=0 $Y2=0
cc_471 N_A_1155_284#_c_608_n N_A_1218_388#_c_774_n 0.0131686f $X=6.05 $Y=1.605
+ $X2=0 $Y2=0
cc_472 N_A_1155_284#_c_609_n N_A_1218_388#_c_792_n 0.0262102f $X=7.54 $Y=2.29
+ $X2=0 $Y2=0
cc_473 N_A_1155_284#_c_610_n N_A_1218_388#_c_792_n 0.00649998f $X=7.985 $Y=0.58
+ $X2=0 $Y2=0
cc_474 N_A_1155_284#_M1010_s N_A_1218_388#_c_783_n 0.00136259f $X=7.35 $Y=2.05
+ $X2=0 $Y2=0
cc_475 N_A_1155_284#_c_617_n N_A_1218_388#_c_783_n 0.00927126f $X=7.495 $Y=2.455
+ $X2=0 $Y2=0
cc_476 N_A_1155_284#_c_609_n N_A_1218_388#_c_783_n 0.0234145f $X=7.54 $Y=2.29
+ $X2=0 $Y2=0
cc_477 N_A_1155_284#_c_612_n N_A_1218_388#_c_784_n 0.0015623f $X=6.05 $Y=2.905
+ $X2=0 $Y2=0
cc_478 N_A_1155_284#_c_606_n N_A_1218_388#_c_785_n 0.00306657f $X=6.015 $Y=1.865
+ $X2=0 $Y2=0
cc_479 N_A_1155_284#_c_612_n N_A_1218_388#_c_785_n 0.0333367f $X=6.05 $Y=2.905
+ $X2=0 $Y2=0
cc_480 N_A_1155_284#_c_613_n N_A_1218_388#_c_785_n 0.0233748f $X=7.33 $Y=2.99
+ $X2=0 $Y2=0
cc_481 N_A_1155_284#_c_609_n N_A_1218_388#_c_775_n 0.00818462f $X=7.54 $Y=2.29
+ $X2=0 $Y2=0
cc_482 N_A_1155_284#_c_609_n N_A_1218_388#_c_776_n 0.00380168f $X=7.54 $Y=2.29
+ $X2=0 $Y2=0
cc_483 N_A_1155_284#_c_609_n N_VPWR_c_996_n 0.0297224f $X=7.54 $Y=2.29 $X2=0
+ $Y2=0
cc_484 N_A_1155_284#_c_613_n N_VPWR_c_997_n 0.00791077f $X=7.33 $Y=2.99 $X2=0
+ $Y2=0
cc_485 N_A_1155_284#_c_615_n N_VPWR_c_997_n 0.00787434f $X=7.415 $Y=2.905 $X2=0
+ $Y2=0
cc_486 N_A_1155_284#_c_617_n N_VPWR_c_1046_n 0.0297224f $X=7.495 $Y=2.455 $X2=0
+ $Y2=0
cc_487 N_A_1155_284#_c_606_n N_VPWR_c_1004_n 0.00128574f $X=6.015 $Y=1.865 $X2=0
+ $Y2=0
cc_488 N_A_1155_284#_c_613_n N_VPWR_c_1004_n 0.0891083f $X=7.33 $Y=2.99 $X2=0
+ $Y2=0
cc_489 N_A_1155_284#_c_614_n N_VPWR_c_1004_n 0.0121867f $X=6.135 $Y=2.99 $X2=0
+ $Y2=0
cc_490 N_A_1155_284#_c_617_n N_VPWR_c_1004_n 0.00490018f $X=7.495 $Y=2.455 $X2=0
+ $Y2=0
cc_491 N_A_1155_284#_c_606_n N_VPWR_c_993_n 8.17763e-19 $X=6.015 $Y=1.865 $X2=0
+ $Y2=0
cc_492 N_A_1155_284#_c_613_n N_VPWR_c_993_n 0.0515306f $X=7.33 $Y=2.99 $X2=0
+ $Y2=0
cc_493 N_A_1155_284#_c_614_n N_VPWR_c_993_n 0.00660921f $X=6.135 $Y=2.99 $X2=0
+ $Y2=0
cc_494 N_A_1155_284#_c_617_n N_VPWR_c_993_n 0.00746272f $X=7.495 $Y=2.455 $X2=0
+ $Y2=0
cc_495 N_A_1155_284#_M1016_g N_A_323_392#_c_1108_n 0.00491067f $X=6.09 $Y=0.935
+ $X2=0 $Y2=0
cc_496 N_A_1155_284#_M1016_g N_A_323_392#_c_1109_n 0.00643069f $X=6.09 $Y=0.935
+ $X2=0 $Y2=0
cc_497 N_A_1155_284#_c_610_n N_A_323_392#_c_1109_n 8.32239e-19 $X=7.985 $Y=0.58
+ $X2=0 $Y2=0
cc_498 N_A_1155_284#_c_609_n N_A_323_392#_c_1111_n 0.0886621f $X=7.54 $Y=2.29
+ $X2=0 $Y2=0
cc_499 N_A_1155_284#_c_610_n N_A_323_392#_c_1111_n 0.0265154f $X=7.985 $Y=0.58
+ $X2=0 $Y2=0
cc_500 N_A_1155_284#_c_613_n N_A_323_392#_c_1115_n 0.0190899f $X=7.33 $Y=2.99
+ $X2=0 $Y2=0
cc_501 N_A_1155_284#_c_617_n N_A_323_392#_c_1115_n 0.0285267f $X=7.495 $Y=2.455
+ $X2=0 $Y2=0
cc_502 N_A_1155_284#_c_609_n N_A_323_392#_c_1115_n 0.00602056f $X=7.54 $Y=2.29
+ $X2=0 $Y2=0
cc_503 N_A_1155_284#_M1010_s N_A_323_392#_c_1116_n 0.00102207f $X=7.35 $Y=2.05
+ $X2=0 $Y2=0
cc_504 N_A_1155_284#_c_617_n N_A_323_392#_c_1116_n 0.00583412f $X=7.495 $Y=2.455
+ $X2=0 $Y2=0
cc_505 N_A_1155_284#_c_609_n N_A_323_392#_c_1116_n 0.0121134f $X=7.54 $Y=2.29
+ $X2=0 $Y2=0
cc_506 N_A_1155_284#_c_606_n N_A_416_118#_c_1239_n 0.00597119f $X=6.015 $Y=1.865
+ $X2=0 $Y2=0
cc_507 N_A_1155_284#_M1016_g N_A_416_118#_c_1239_n 0.0161112f $X=6.09 $Y=0.935
+ $X2=0 $Y2=0
cc_508 N_A_1155_284#_c_608_n N_A_416_118#_c_1239_n 0.0263503f $X=6.05 $Y=1.605
+ $X2=0 $Y2=0
cc_509 N_A_1155_284#_M1016_g N_A_416_118#_c_1291_n 0.0131515f $X=6.09 $Y=0.935
+ $X2=0 $Y2=0
cc_510 N_A_1155_284#_M1016_g N_A_416_118#_c_1242_n 0.00531168f $X=6.09 $Y=0.935
+ $X2=0 $Y2=0
cc_511 N_A_1155_284#_M1016_g N_A_416_118#_c_1243_n 2.06791e-19 $X=6.09 $Y=0.935
+ $X2=0 $Y2=0
cc_512 N_A_1155_284#_c_612_n N_A_416_118#_c_1248_n 0.00113479f $X=6.05 $Y=2.905
+ $X2=0 $Y2=0
cc_513 N_A_1155_284#_c_606_n N_A_416_118#_c_1249_n 0.0181742f $X=6.015 $Y=1.865
+ $X2=0 $Y2=0
cc_514 N_A_1155_284#_c_612_n N_A_416_118#_c_1249_n 0.0643787f $X=6.05 $Y=2.905
+ $X2=0 $Y2=0
cc_515 N_A_1155_284#_c_608_n N_A_416_118#_c_1249_n 0.0015883f $X=6.05 $Y=1.605
+ $X2=0 $Y2=0
cc_516 N_A_1155_284#_c_606_n N_A_416_118#_c_1244_n 0.005784f $X=6.015 $Y=1.865
+ $X2=0 $Y2=0
cc_517 N_A_1155_284#_M1016_g N_A_416_118#_c_1244_n 0.0034264f $X=6.09 $Y=0.935
+ $X2=0 $Y2=0
cc_518 N_A_1155_284#_c_612_n N_A_416_118#_c_1244_n 0.00691963f $X=6.05 $Y=2.905
+ $X2=0 $Y2=0
cc_519 N_A_1155_284#_c_608_n N_A_416_118#_c_1244_n 0.0218967f $X=6.05 $Y=1.605
+ $X2=0 $Y2=0
cc_520 N_A_1155_284#_c_609_n N_VGND_c_1420_n 0.00998489f $X=7.54 $Y=2.29 $X2=0
+ $Y2=0
cc_521 N_A_1155_284#_c_610_n N_VGND_c_1428_n 0.0177026f $X=7.985 $Y=0.58 $X2=0
+ $Y2=0
cc_522 N_A_1155_284#_c_610_n N_VGND_c_1433_n 0.0195345f $X=7.985 $Y=0.58 $X2=0
+ $Y2=0
cc_523 N_C_c_697_n N_A_1218_388#_M1007_g 0.0119424f $X=8.2 $Y=0.865 $X2=0 $Y2=0
cc_524 N_C_c_692_n N_A_1218_388#_c_774_n 0.0144668f $X=6.695 $Y=1.865 $X2=0
+ $Y2=0
cc_525 N_C_M1021_g N_A_1218_388#_c_774_n 0.00287028f $X=6.77 $Y=0.935 $X2=0
+ $Y2=0
cc_526 N_C_c_699_n N_A_1218_388#_c_774_n 6.7552e-19 $X=7.28 $Y=1.712 $X2=0 $Y2=0
cc_527 C N_A_1218_388#_c_774_n 0.023122f $X=6.875 $Y=1.58 $X2=0 $Y2=0
cc_528 N_C_c_695_n N_A_1218_388#_c_792_n 0.00183965f $X=8.125 $Y=0.94 $X2=0
+ $Y2=0
cc_529 N_C_c_692_n N_A_1218_388#_c_783_n 0.0116169f $X=6.695 $Y=1.865 $X2=0
+ $Y2=0
cc_530 N_C_c_702_n N_A_1218_388#_c_783_n 0.0103857f $X=7.645 $Y=1.9 $X2=0 $Y2=0
cc_531 N_C_c_703_n N_A_1218_388#_c_783_n 0.00396916f $X=7.72 $Y=1.975 $X2=0
+ $Y2=0
cc_532 C N_A_1218_388#_c_783_n 0.0027894f $X=6.875 $Y=1.58 $X2=0 $Y2=0
cc_533 N_C_c_692_n N_A_1218_388#_c_785_n 0.0105767f $X=6.695 $Y=1.865 $X2=0
+ $Y2=0
cc_534 N_C_c_694_n N_A_1218_388#_c_776_n 0.00633084f $X=7.28 $Y=1.45 $X2=0 $Y2=0
cc_535 N_C_c_695_n N_A_1218_388#_c_776_n 0.0238665f $X=8.125 $Y=0.94 $X2=0 $Y2=0
cc_536 N_C_c_702_n N_VPWR_c_996_n 0.00394244f $X=7.645 $Y=1.9 $X2=0 $Y2=0
cc_537 N_C_c_703_n N_VPWR_c_996_n 0.0170515f $X=7.72 $Y=1.975 $X2=0 $Y2=0
cc_538 N_C_c_692_n N_VPWR_c_1004_n 6.29586e-19 $X=6.695 $Y=1.865 $X2=0 $Y2=0
cc_539 N_C_c_703_n N_VPWR_c_1004_n 0.00342894f $X=7.72 $Y=1.975 $X2=0 $Y2=0
cc_540 N_C_c_703_n N_VPWR_c_993_n 0.00465306f $X=7.72 $Y=1.975 $X2=0 $Y2=0
cc_541 N_C_M1021_g N_A_323_392#_c_1109_n 0.00449889f $X=6.77 $Y=0.935 $X2=0
+ $Y2=0
cc_542 N_C_c_696_n N_A_323_392#_c_1109_n 0.00107968f $X=7.355 $Y=0.94 $X2=0
+ $Y2=0
cc_543 N_C_c_692_n N_A_323_392#_c_1111_n 5.94319e-19 $X=6.695 $Y=1.865 $X2=0
+ $Y2=0
cc_544 N_C_M1021_g N_A_323_392#_c_1111_n 0.00417992f $X=6.77 $Y=0.935 $X2=0
+ $Y2=0
cc_545 N_C_c_694_n N_A_323_392#_c_1111_n 0.0125253f $X=7.28 $Y=1.45 $X2=0 $Y2=0
cc_546 N_C_c_695_n N_A_323_392#_c_1111_n 0.00531516f $X=8.125 $Y=0.94 $X2=0
+ $Y2=0
cc_547 N_C_c_696_n N_A_323_392#_c_1111_n 0.00509903f $X=7.355 $Y=0.94 $X2=0
+ $Y2=0
cc_548 N_C_c_702_n N_A_323_392#_c_1111_n 0.00377414f $X=7.645 $Y=1.9 $X2=0 $Y2=0
cc_549 N_C_c_699_n N_A_323_392#_c_1111_n 0.0161522f $X=7.28 $Y=1.712 $X2=0 $Y2=0
cc_550 C N_A_323_392#_c_1111_n 0.023122f $X=6.875 $Y=1.58 $X2=0 $Y2=0
cc_551 N_C_c_692_n N_A_323_392#_c_1115_n 0.00330358f $X=6.695 $Y=1.865 $X2=0
+ $Y2=0
cc_552 N_C_c_703_n N_A_323_392#_c_1115_n 0.00164413f $X=7.72 $Y=1.975 $X2=0
+ $Y2=0
cc_553 N_C_c_692_n N_A_323_392#_c_1116_n 0.00163539f $X=6.695 $Y=1.865 $X2=0
+ $Y2=0
cc_554 N_C_c_702_n N_A_323_392#_c_1116_n 0.00149593f $X=7.645 $Y=1.9 $X2=0 $Y2=0
cc_555 N_C_c_703_n N_A_323_392#_c_1116_n 8.39033e-19 $X=7.72 $Y=1.975 $X2=0
+ $Y2=0
cc_556 N_C_c_698_n N_A_323_392#_c_1116_n 0.00543944f $X=7.205 $Y=1.615 $X2=0
+ $Y2=0
cc_557 N_C_c_699_n N_A_323_392#_c_1116_n 0.00522443f $X=7.28 $Y=1.712 $X2=0
+ $Y2=0
cc_558 C N_A_323_392#_c_1116_n 0.0157311f $X=6.875 $Y=1.58 $X2=0 $Y2=0
cc_559 N_C_M1021_g N_A_416_118#_c_1291_n 0.00148249f $X=6.77 $Y=0.935 $X2=0
+ $Y2=0
cc_560 N_C_M1021_g N_A_416_118#_c_1241_n 0.0114827f $X=6.77 $Y=0.935 $X2=0 $Y2=0
cc_561 N_C_M1021_g N_A_416_118#_c_1243_n 0.00821222f $X=6.77 $Y=0.935 $X2=0
+ $Y2=0
cc_562 N_C_c_696_n N_A_416_118#_c_1243_n 0.0033372f $X=7.355 $Y=0.94 $X2=0 $Y2=0
cc_563 N_C_c_698_n N_A_416_118#_c_1243_n 0.00105117f $X=7.205 $Y=1.615 $X2=0
+ $Y2=0
cc_564 C N_A_416_118#_c_1243_n 0.0204158f $X=6.875 $Y=1.58 $X2=0 $Y2=0
cc_565 N_C_c_697_n N_VGND_c_1420_n 0.0100812f $X=8.2 $Y=0.865 $X2=0 $Y2=0
cc_566 N_C_c_697_n N_VGND_c_1428_n 0.00434593f $X=8.2 $Y=0.865 $X2=0 $Y2=0
cc_567 N_C_c_696_n N_VGND_c_1433_n 0.00344512f $X=7.355 $Y=0.94 $X2=0 $Y2=0
cc_568 N_C_c_697_n N_VGND_c_1433_n 0.0082439f $X=8.2 $Y=0.865 $X2=0 $Y2=0
cc_569 N_A_1218_388#_c_783_n N_VPWR_M1010_d 0.00918901f $X=8.255 $Y=2.035 $X2=0
+ $Y2=0
cc_570 N_A_1218_388#_c_817_p N_VPWR_M1010_d 0.00645288f $X=8.4 $Y=2.035 $X2=0
+ $Y2=0
cc_571 N_A_1218_388#_c_775_n N_VPWR_M1010_d 0.00643242f $X=8.4 $Y=2.035 $X2=0
+ $Y2=0
cc_572 N_A_1218_388#_c_778_n N_VPWR_c_996_n 0.00299716f $X=8.625 $Y=1.765 $X2=0
+ $Y2=0
cc_573 N_A_1218_388#_c_792_n N_VPWR_c_996_n 0.010165f $X=8.285 $Y=1.42 $X2=0
+ $Y2=0
cc_574 N_A_1218_388#_c_783_n N_VPWR_c_996_n 0.0168569f $X=8.255 $Y=2.035 $X2=0
+ $Y2=0
cc_575 N_A_1218_388#_c_817_p N_VPWR_c_996_n 0.00266295f $X=8.4 $Y=2.035 $X2=0
+ $Y2=0
cc_576 N_A_1218_388#_c_775_n N_VPWR_c_996_n 0.0228911f $X=8.4 $Y=2.035 $X2=0
+ $Y2=0
cc_577 N_A_1218_388#_c_776_n N_VPWR_c_996_n 0.0037797f $X=8.535 $Y=1.42 $X2=0
+ $Y2=0
cc_578 N_A_1218_388#_c_778_n N_VPWR_c_997_n 0.0053874f $X=8.625 $Y=1.765 $X2=0
+ $Y2=0
cc_579 N_A_1218_388#_c_778_n N_VPWR_c_998_n 0.00445602f $X=8.625 $Y=1.765 $X2=0
+ $Y2=0
cc_580 N_A_1218_388#_c_779_n N_VPWR_c_998_n 0.00320971f $X=9.075 $Y=1.765 $X2=0
+ $Y2=0
cc_581 N_A_1218_388#_c_779_n N_VPWR_c_999_n 0.0104311f $X=9.075 $Y=1.765 $X2=0
+ $Y2=0
cc_582 N_A_1218_388#_c_780_n N_VPWR_c_999_n 0.00685194f $X=9.605 $Y=1.765 $X2=0
+ $Y2=0
cc_583 N_A_1218_388#_c_777_n N_VPWR_c_999_n 0.00432997f $X=10.055 $Y=1.51 $X2=0
+ $Y2=0
cc_584 N_A_1218_388#_c_781_n N_VPWR_c_1001_n 0.0100916f $X=10.055 $Y=1.765 $X2=0
+ $Y2=0
cc_585 N_A_1218_388#_c_783_n N_VPWR_c_1046_n 0.00696054f $X=8.255 $Y=2.035 $X2=0
+ $Y2=0
cc_586 N_A_1218_388#_c_817_p N_VPWR_c_1046_n 0.00350284f $X=8.4 $Y=2.035 $X2=0
+ $Y2=0
cc_587 N_A_1218_388#_c_775_n N_VPWR_c_1046_n 0.0141983f $X=8.4 $Y=2.035 $X2=0
+ $Y2=0
cc_588 N_A_1218_388#_c_780_n N_VPWR_c_1005_n 0.00445602f $X=9.605 $Y=1.765 $X2=0
+ $Y2=0
cc_589 N_A_1218_388#_c_781_n N_VPWR_c_1005_n 0.00445602f $X=10.055 $Y=1.765
+ $X2=0 $Y2=0
cc_590 N_A_1218_388#_c_778_n N_VPWR_c_993_n 0.00862055f $X=8.625 $Y=1.765 $X2=0
+ $Y2=0
cc_591 N_A_1218_388#_c_779_n N_VPWR_c_993_n 0.00455513f $X=9.075 $Y=1.765 $X2=0
+ $Y2=0
cc_592 N_A_1218_388#_c_780_n N_VPWR_c_993_n 0.00858307f $X=9.605 $Y=1.765 $X2=0
+ $Y2=0
cc_593 N_A_1218_388#_c_781_n N_VPWR_c_993_n 0.00861084f $X=10.055 $Y=1.765 $X2=0
+ $Y2=0
cc_594 N_A_1218_388#_c_783_n N_A_323_392#_M1020_d 0.00326211f $X=8.255 $Y=2.035
+ $X2=0 $Y2=0
cc_595 N_A_1218_388#_c_774_n N_A_323_392#_c_1111_n 0.0086988f $X=6.555 $Y=1.105
+ $X2=0 $Y2=0
cc_596 N_A_1218_388#_c_783_n N_A_323_392#_c_1111_n 0.00365456f $X=8.255 $Y=2.035
+ $X2=0 $Y2=0
cc_597 N_A_1218_388#_c_783_n N_A_323_392#_c_1115_n 0.00539563f $X=8.255 $Y=2.035
+ $X2=0 $Y2=0
cc_598 N_A_1218_388#_c_784_n N_A_323_392#_c_1115_n 2.21397e-19 $X=6.625 $Y=2.035
+ $X2=0 $Y2=0
cc_599 N_A_1218_388#_c_785_n N_A_323_392#_c_1115_n 0.0418677f $X=6.48 $Y=2.035
+ $X2=0 $Y2=0
cc_600 N_A_1218_388#_c_783_n N_A_323_392#_c_1116_n 0.0340455f $X=8.255 $Y=2.035
+ $X2=0 $Y2=0
cc_601 N_A_1218_388#_c_784_n N_A_323_392#_c_1116_n 2.23197e-19 $X=6.625 $Y=2.035
+ $X2=0 $Y2=0
cc_602 N_A_1218_388#_c_785_n N_A_323_392#_c_1116_n 0.0100311f $X=6.48 $Y=2.035
+ $X2=0 $Y2=0
cc_603 N_A_1218_388#_M1016_d N_A_416_118#_c_1239_n 0.00128304f $X=6.165 $Y=0.615
+ $X2=0 $Y2=0
cc_604 N_A_1218_388#_c_774_n N_A_416_118#_c_1239_n 0.0139392f $X=6.555 $Y=1.105
+ $X2=0 $Y2=0
cc_605 N_A_1218_388#_M1016_d N_A_416_118#_c_1291_n 0.00399932f $X=6.165 $Y=0.615
+ $X2=0 $Y2=0
cc_606 N_A_1218_388#_c_774_n N_A_416_118#_c_1291_n 0.0134008f $X=6.555 $Y=1.105
+ $X2=0 $Y2=0
cc_607 N_A_1218_388#_M1016_d N_A_416_118#_c_1241_n 0.00964f $X=6.165 $Y=0.615
+ $X2=0 $Y2=0
cc_608 N_A_1218_388#_c_774_n N_A_416_118#_c_1241_n 0.0135869f $X=6.555 $Y=1.105
+ $X2=0 $Y2=0
cc_609 N_A_1218_388#_c_774_n N_A_416_118#_c_1243_n 0.012365f $X=6.555 $Y=1.105
+ $X2=0 $Y2=0
cc_610 N_A_1218_388#_c_778_n N_X_c_1360_n 0.0123254f $X=8.625 $Y=1.765 $X2=0
+ $Y2=0
cc_611 N_A_1218_388#_c_779_n N_X_c_1360_n 0.0178977f $X=9.075 $Y=1.765 $X2=0
+ $Y2=0
cc_612 N_A_1218_388#_M1007_g N_X_c_1356_n 0.0065213f $X=8.78 $Y=0.74 $X2=0 $Y2=0
cc_613 N_A_1218_388#_M1017_g N_X_c_1356_n 0.00652624f $X=9.21 $Y=0.74 $X2=0
+ $Y2=0
cc_614 N_A_1218_388#_M1018_g N_X_c_1356_n 5.98536e-19 $X=9.64 $Y=0.74 $X2=0
+ $Y2=0
cc_615 N_A_1218_388#_M1007_g N_X_c_1357_n 0.00385423f $X=8.78 $Y=0.74 $X2=0
+ $Y2=0
cc_616 N_A_1218_388#_M1017_g N_X_c_1357_n 0.0037907f $X=9.21 $Y=0.74 $X2=0 $Y2=0
cc_617 N_A_1218_388#_c_864_p N_X_c_1357_n 0.00336044f $X=8.695 $Y=1.42 $X2=0
+ $Y2=0
cc_618 N_A_1218_388#_c_777_n N_X_c_1357_n 0.00474311f $X=10.055 $Y=1.51 $X2=0
+ $Y2=0
cc_619 N_A_1218_388#_c_777_n N_X_c_1373_n 0.0399195f $X=10.055 $Y=1.51 $X2=0
+ $Y2=0
cc_620 N_A_1218_388#_M1017_g N_X_c_1358_n 6.00118e-19 $X=9.21 $Y=0.74 $X2=0
+ $Y2=0
cc_621 N_A_1218_388#_M1018_g N_X_c_1358_n 0.0124921f $X=9.64 $Y=0.74 $X2=0 $Y2=0
cc_622 N_A_1218_388#_M1024_g N_X_c_1358_n 0.00374969f $X=10.07 $Y=0.74 $X2=0
+ $Y2=0
cc_623 N_A_1218_388#_c_777_n N_X_c_1358_n 0.00637697f $X=10.055 $Y=1.51 $X2=0
+ $Y2=0
cc_624 N_A_1218_388#_c_778_n N_X_c_1361_n 0.00263077f $X=8.625 $Y=1.765 $X2=0
+ $Y2=0
cc_625 N_A_1218_388#_c_779_n N_X_c_1361_n 0.00394322f $X=9.075 $Y=1.765 $X2=0
+ $Y2=0
cc_626 N_A_1218_388#_c_864_p N_X_c_1361_n 0.00648931f $X=8.695 $Y=1.42 $X2=0
+ $Y2=0
cc_627 N_A_1218_388#_c_817_p N_X_c_1361_n 0.00749736f $X=8.4 $Y=2.035 $X2=0
+ $Y2=0
cc_628 N_A_1218_388#_c_775_n N_X_c_1361_n 0.0159487f $X=8.4 $Y=2.035 $X2=0 $Y2=0
cc_629 N_A_1218_388#_c_777_n N_X_c_1361_n 0.0099448f $X=10.055 $Y=1.51 $X2=0
+ $Y2=0
cc_630 N_A_1218_388#_c_778_n N_X_c_1359_n 3.97716e-19 $X=8.625 $Y=1.765 $X2=0
+ $Y2=0
cc_631 N_A_1218_388#_c_779_n N_X_c_1359_n 0.00156626f $X=9.075 $Y=1.765 $X2=0
+ $Y2=0
cc_632 N_A_1218_388#_c_780_n N_X_c_1359_n 5.2193e-19 $X=9.605 $Y=1.765 $X2=0
+ $Y2=0
cc_633 N_A_1218_388#_c_864_p N_X_c_1359_n 0.00864993f $X=8.695 $Y=1.42 $X2=0
+ $Y2=0
cc_634 N_A_1218_388#_c_775_n N_X_c_1359_n 0.00931569f $X=8.4 $Y=2.035 $X2=0
+ $Y2=0
cc_635 N_A_1218_388#_c_777_n N_X_c_1359_n 0.0146992f $X=10.055 $Y=1.51 $X2=0
+ $Y2=0
cc_636 N_A_1218_388#_M1007_g N_X_c_1390_n 0.00284927f $X=8.78 $Y=0.74 $X2=0
+ $Y2=0
cc_637 N_A_1218_388#_M1017_g N_X_c_1390_n 0.0017052f $X=9.21 $Y=0.74 $X2=0 $Y2=0
cc_638 N_A_1218_388#_c_777_n N_X_c_1390_n 4.44413e-19 $X=10.055 $Y=1.51 $X2=0
+ $Y2=0
cc_639 N_A_1218_388#_c_864_p N_X_c_1393_n 0.0143906f $X=8.695 $Y=1.42 $X2=0
+ $Y2=0
cc_640 N_A_1218_388#_c_777_n N_X_c_1393_n 0.00745846f $X=10.055 $Y=1.51 $X2=0
+ $Y2=0
cc_641 N_A_1218_388#_c_779_n X 4.48652e-19 $X=9.075 $Y=1.765 $X2=0 $Y2=0
cc_642 N_A_1218_388#_c_780_n X 0.0148233f $X=9.605 $Y=1.765 $X2=0 $Y2=0
cc_643 N_A_1218_388#_c_781_n X 0.0167069f $X=10.055 $Y=1.765 $X2=0 $Y2=0
cc_644 N_A_1218_388#_c_777_n X 0.00514228f $X=10.055 $Y=1.51 $X2=0 $Y2=0
cc_645 N_A_1218_388#_c_777_n N_X_c_1399_n 0.0455429f $X=10.055 $Y=1.51 $X2=0
+ $Y2=0
cc_646 N_A_1218_388#_M1007_g N_VGND_c_1420_n 0.005585f $X=8.78 $Y=0.74 $X2=0
+ $Y2=0
cc_647 N_A_1218_388#_c_864_p N_VGND_c_1420_n 0.0265884f $X=8.695 $Y=1.42 $X2=0
+ $Y2=0
cc_648 N_A_1218_388#_c_776_n N_VGND_c_1420_n 0.00804883f $X=8.535 $Y=1.42 $X2=0
+ $Y2=0
cc_649 N_A_1218_388#_M1007_g N_VGND_c_1421_n 0.00434272f $X=8.78 $Y=0.74 $X2=0
+ $Y2=0
cc_650 N_A_1218_388#_M1017_g N_VGND_c_1421_n 0.00434272f $X=9.21 $Y=0.74 $X2=0
+ $Y2=0
cc_651 N_A_1218_388#_M1017_g N_VGND_c_1422_n 0.00313962f $X=9.21 $Y=0.74 $X2=0
+ $Y2=0
cc_652 N_A_1218_388#_M1018_g N_VGND_c_1422_n 0.001891f $X=9.64 $Y=0.74 $X2=0
+ $Y2=0
cc_653 N_A_1218_388#_c_777_n N_VGND_c_1422_n 0.00245982f $X=10.055 $Y=1.51 $X2=0
+ $Y2=0
cc_654 N_A_1218_388#_M1018_g N_VGND_c_1424_n 6.14817e-19 $X=9.64 $Y=0.74 $X2=0
+ $Y2=0
cc_655 N_A_1218_388#_M1024_g N_VGND_c_1424_n 0.0160198f $X=10.07 $Y=0.74 $X2=0
+ $Y2=0
cc_656 N_A_1218_388#_M1018_g N_VGND_c_1429_n 0.00434272f $X=9.64 $Y=0.74 $X2=0
+ $Y2=0
cc_657 N_A_1218_388#_M1024_g N_VGND_c_1429_n 0.00383152f $X=10.07 $Y=0.74 $X2=0
+ $Y2=0
cc_658 N_A_1218_388#_M1007_g N_VGND_c_1433_n 0.00821384f $X=8.78 $Y=0.74 $X2=0
+ $Y2=0
cc_659 N_A_1218_388#_M1017_g N_VGND_c_1433_n 0.00820284f $X=9.21 $Y=0.74 $X2=0
+ $Y2=0
cc_660 N_A_1218_388#_M1018_g N_VGND_c_1433_n 0.00820284f $X=9.64 $Y=0.74 $X2=0
+ $Y2=0
cc_661 N_A_1218_388#_M1024_g N_VGND_c_1433_n 0.0075754f $X=10.07 $Y=0.74 $X2=0
+ $Y2=0
cc_662 N_A_27_118#_c_918_n N_VPWR_c_994_n 0.0541024f $X=0.225 $Y=2.32 $X2=0
+ $Y2=0
cc_663 N_A_27_118#_c_919_n N_VPWR_c_1002_n 0.0124046f $X=0.28 $Y=2.345 $X2=0
+ $Y2=0
cc_664 N_A_27_118#_c_919_n N_VPWR_c_993_n 0.0102675f $X=0.28 $Y=2.345 $X2=0
+ $Y2=0
cc_665 N_A_27_118#_c_913_n N_A_323_392#_c_1119_n 0.014161f $X=2.3 $Y=2.21 $X2=0
+ $Y2=0
cc_666 N_A_27_118#_c_914_n N_A_323_392#_c_1119_n 0.00442522f $X=2.68 $Y=1.42
+ $X2=0 $Y2=0
cc_667 N_A_27_118#_M1011_d N_A_323_392#_c_1112_n 0.0076127f $X=2.15 $Y=1.96
+ $X2=0 $Y2=0
cc_668 N_A_27_118#_c_913_n N_A_323_392#_c_1112_n 0.0154248f $X=2.3 $Y=2.21 $X2=0
+ $Y2=0
cc_669 N_A_27_118#_c_912_n N_A_416_118#_c_1235_n 0.0176692f $X=1.88 $Y=1.42
+ $X2=0 $Y2=0
cc_670 N_A_27_118#_c_914_n N_A_416_118#_c_1235_n 0.0209451f $X=2.68 $Y=1.42
+ $X2=0 $Y2=0
cc_671 N_A_27_118#_c_915_n N_A_416_118#_c_1235_n 0.0180573f $X=2.72 $Y=1.02
+ $X2=0 $Y2=0
cc_672 N_A_27_118#_M1022_d N_A_416_118#_c_1236_n 0.00681577f $X=2.58 $Y=0.81
+ $X2=0 $Y2=0
cc_673 N_A_27_118#_c_915_n N_A_416_118#_c_1236_n 0.0199631f $X=2.72 $Y=1.02
+ $X2=0 $Y2=0
cc_674 N_A_27_118#_c_911_n N_A_416_118#_c_1237_n 0.00211437f $X=1.795 $Y=0.665
+ $X2=0 $Y2=0
cc_675 N_A_27_118#_c_913_n N_A_416_118#_c_1238_n 0.00815753f $X=2.3 $Y=2.21
+ $X2=0 $Y2=0
cc_676 N_A_27_118#_c_914_n N_A_416_118#_c_1238_n 0.014189f $X=2.68 $Y=1.42 $X2=0
+ $Y2=0
cc_677 N_A_27_118#_c_915_n N_A_416_118#_c_1238_n 0.0316281f $X=2.72 $Y=1.02
+ $X2=0 $Y2=0
cc_678 N_A_27_118#_M1011_d N_A_416_118#_c_1247_n 0.00114654f $X=2.15 $Y=1.96
+ $X2=0 $Y2=0
cc_679 N_A_27_118#_c_913_n N_A_416_118#_c_1247_n 0.00778267f $X=2.3 $Y=2.21
+ $X2=0 $Y2=0
cc_680 N_A_27_118#_c_914_n N_A_416_118#_c_1247_n 0.00370897f $X=2.68 $Y=1.42
+ $X2=0 $Y2=0
cc_681 N_A_27_118#_c_913_n N_A_416_118#_c_1250_n 0.0276551f $X=2.3 $Y=2.21 $X2=0
+ $Y2=0
cc_682 N_A_27_118#_c_914_n N_A_416_118#_c_1250_n 0.01239f $X=2.68 $Y=1.42 $X2=0
+ $Y2=0
cc_683 N_A_27_118#_c_911_n N_VGND_M1012_d 0.0178489f $X=1.795 $Y=0.665 $X2=-0.19
+ $Y2=-0.245
cc_684 N_A_27_118#_c_911_n N_VGND_c_1425_n 0.0191349f $X=1.795 $Y=0.665 $X2=0
+ $Y2=0
cc_685 N_A_27_118#_c_909_n N_VGND_c_1427_n 0.00833654f $X=0.265 $Y=0.75 $X2=0
+ $Y2=0
cc_686 N_A_27_118#_c_911_n N_VGND_c_1427_n 0.00345394f $X=1.795 $Y=0.665 $X2=0
+ $Y2=0
cc_687 N_A_27_118#_c_911_n N_VGND_c_1430_n 0.0306422f $X=1.795 $Y=0.665 $X2=0
+ $Y2=0
cc_688 N_A_27_118#_c_909_n N_VGND_c_1433_n 0.0114278f $X=0.265 $Y=0.75 $X2=0
+ $Y2=0
cc_689 N_A_27_118#_c_911_n N_VGND_c_1433_n 0.0350406f $X=1.795 $Y=0.665 $X2=0
+ $Y2=0
cc_690 N_VPWR_c_995_n N_A_416_118#_c_1246_n 0.0306649f $X=5.07 $Y=1.985 $X2=0
+ $Y2=0
cc_691 N_VPWR_c_995_n N_A_416_118#_c_1248_n 0.00270171f $X=5.07 $Y=1.985 $X2=0
+ $Y2=0
cc_692 N_VPWR_c_995_n N_A_416_118#_c_1249_n 0.0711484f $X=5.07 $Y=1.985 $X2=0
+ $Y2=0
cc_693 N_VPWR_c_1004_n N_A_416_118#_c_1249_n 0.00994744f $X=7.945 $Y=3.33 $X2=0
+ $Y2=0
cc_694 N_VPWR_c_993_n N_A_416_118#_c_1249_n 0.012708f $X=10.32 $Y=3.33 $X2=0
+ $Y2=0
cc_695 N_VPWR_c_995_n N_A_416_118#_c_1244_n 0.00704007f $X=5.07 $Y=1.985 $X2=0
+ $Y2=0
cc_696 N_VPWR_c_996_n N_X_c_1360_n 0.00524247f $X=8.03 $Y=1.985 $X2=0 $Y2=0
cc_697 N_VPWR_c_997_n N_X_c_1360_n 0.0246224f $X=8.222 $Y=3.245 $X2=0 $Y2=0
cc_698 N_VPWR_c_998_n N_X_c_1360_n 0.0191315f $X=9.295 $Y=3.33 $X2=0 $Y2=0
cc_699 N_VPWR_c_993_n N_X_c_1360_n 0.0155112f $X=10.32 $Y=3.33 $X2=0 $Y2=0
cc_700 N_VPWR_c_999_n N_X_c_1373_n 0.00793475f $X=9.38 $Y=1.985 $X2=0 $Y2=0
cc_701 N_VPWR_c_999_n N_X_c_1361_n 0.0876229f $X=9.38 $Y=1.985 $X2=0 $Y2=0
cc_702 N_VPWR_c_999_n X 0.0756134f $X=9.38 $Y=1.985 $X2=0 $Y2=0
cc_703 N_VPWR_c_1001_n X 0.0778383f $X=10.28 $Y=1.985 $X2=0 $Y2=0
cc_704 N_VPWR_c_1005_n X 0.014552f $X=10.195 $Y=3.33 $X2=0 $Y2=0
cc_705 N_VPWR_c_993_n X 0.0119791f $X=10.32 $Y=3.33 $X2=0 $Y2=0
cc_706 N_A_323_392#_c_1112_n N_A_416_118#_M1004_d 0.00480583f $X=3.315 $Y=2.65
+ $X2=0 $Y2=0
cc_707 N_A_323_392#_c_1104_n N_A_416_118#_c_1236_n 0.0135457f $X=3.4 $Y=0.735
+ $X2=0 $Y2=0
cc_708 N_A_323_392#_c_1104_n N_A_416_118#_c_1238_n 0.0891871f $X=3.4 $Y=0.735
+ $X2=0 $Y2=0
cc_709 N_A_323_392#_M1016_s N_A_416_118#_c_1239_n 0.00302199f $X=5.74 $Y=0.615
+ $X2=0 $Y2=0
cc_710 N_A_323_392#_c_1107_n N_A_416_118#_c_1239_n 0.0281376f $X=5.71 $Y=0.865
+ $X2=0 $Y2=0
cc_711 N_A_323_392#_c_1107_n N_A_416_118#_c_1240_n 0.0143117f $X=5.71 $Y=0.865
+ $X2=0 $Y2=0
cc_712 N_A_323_392#_c_1109_n N_A_416_118#_c_1241_n 0.0363659f $X=7.24 $Y=0.34
+ $X2=0 $Y2=0
cc_713 N_A_323_392#_c_1108_n N_A_416_118#_c_1242_n 0.00792225f $X=5.875 $Y=0.77
+ $X2=0 $Y2=0
cc_714 N_A_323_392#_c_1109_n N_A_416_118#_c_1242_n 0.0133131f $X=7.24 $Y=0.34
+ $X2=0 $Y2=0
cc_715 N_A_323_392#_c_1109_n N_A_416_118#_c_1243_n 0.0196514f $X=7.24 $Y=0.34
+ $X2=0 $Y2=0
cc_716 N_A_323_392#_c_1111_n N_A_416_118#_c_1243_n 0.0513303f $X=7.325 $Y=1.95
+ $X2=0 $Y2=0
cc_717 N_A_323_392#_c_1112_n N_A_416_118#_c_1246_n 0.0063627f $X=3.315 $Y=2.65
+ $X2=0 $Y2=0
cc_718 N_A_323_392#_c_1104_n N_A_416_118#_c_1246_n 0.0187807f $X=3.4 $Y=0.735
+ $X2=0 $Y2=0
cc_719 N_A_323_392#_c_1112_n N_A_416_118#_c_1247_n 0.00319828f $X=3.315 $Y=2.65
+ $X2=0 $Y2=0
cc_720 N_A_323_392#_c_1104_n N_A_416_118#_c_1247_n 3.25096e-19 $X=3.4 $Y=0.735
+ $X2=0 $Y2=0
cc_721 N_A_323_392#_c_1112_n N_A_416_118#_c_1250_n 0.032291f $X=3.315 $Y=2.65
+ $X2=0 $Y2=0
cc_722 N_A_323_392#_c_1104_n N_A_416_118#_c_1250_n 0.0233665f $X=3.4 $Y=0.735
+ $X2=0 $Y2=0
cc_723 N_A_323_392#_c_1105_n N_VGND_M1026_d 0.00138668f $X=4.91 $Y=0.34 $X2=0
+ $Y2=0
cc_724 N_A_323_392#_c_1151_n N_VGND_M1026_d 0.00522053f $X=4.995 $Y=0.78 $X2=0
+ $Y2=0
cc_725 N_A_323_392#_c_1107_n N_VGND_M1026_d 0.0181293f $X=5.71 $Y=0.865 $X2=0
+ $Y2=0
cc_726 N_A_323_392#_c_1155_n N_VGND_M1026_d 7.95616e-19 $X=5.08 $Y=0.865 $X2=0
+ $Y2=0
cc_727 N_A_323_392#_c_1105_n N_VGND_c_1419_n 0.014344f $X=4.91 $Y=0.34 $X2=0
+ $Y2=0
cc_728 N_A_323_392#_c_1151_n N_VGND_c_1419_n 0.0138003f $X=4.995 $Y=0.78 $X2=0
+ $Y2=0
cc_729 N_A_323_392#_c_1107_n N_VGND_c_1419_n 0.0197465f $X=5.71 $Y=0.865 $X2=0
+ $Y2=0
cc_730 N_A_323_392#_c_1108_n N_VGND_c_1419_n 0.0127034f $X=5.875 $Y=0.77 $X2=0
+ $Y2=0
cc_731 N_A_323_392#_c_1110_n N_VGND_c_1419_n 0.0127057f $X=5.96 $Y=0.34 $X2=0
+ $Y2=0
cc_732 N_A_323_392#_c_1105_n N_VGND_c_1425_n 0.103037f $X=4.91 $Y=0.34 $X2=0
+ $Y2=0
cc_733 N_A_323_392#_c_1106_n N_VGND_c_1425_n 0.0115893f $X=3.485 $Y=0.34 $X2=0
+ $Y2=0
cc_734 N_A_323_392#_c_1109_n N_VGND_c_1428_n 0.0945839f $X=7.24 $Y=0.34 $X2=0
+ $Y2=0
cc_735 N_A_323_392#_c_1110_n N_VGND_c_1428_n 0.0179514f $X=5.96 $Y=0.34 $X2=0
+ $Y2=0
cc_736 N_A_323_392#_c_1105_n N_VGND_c_1433_n 0.055579f $X=4.91 $Y=0.34 $X2=0
+ $Y2=0
cc_737 N_A_323_392#_c_1106_n N_VGND_c_1433_n 0.00583135f $X=3.485 $Y=0.34 $X2=0
+ $Y2=0
cc_738 N_A_323_392#_c_1107_n N_VGND_c_1433_n 0.0147576f $X=5.71 $Y=0.865 $X2=0
+ $Y2=0
cc_739 N_A_323_392#_c_1109_n N_VGND_c_1433_n 0.0547264f $X=7.24 $Y=0.34 $X2=0
+ $Y2=0
cc_740 N_A_323_392#_c_1110_n N_VGND_c_1433_n 0.00972504f $X=5.96 $Y=0.34 $X2=0
+ $Y2=0
cc_741 N_A_416_118#_c_1236_n N_VGND_c_1425_n 0.0220173f $X=2.975 $Y=0.535 $X2=0
+ $Y2=0
cc_742 N_A_416_118#_c_1237_n N_VGND_c_1425_n 0.00792677f $X=2.385 $Y=0.535 $X2=0
+ $Y2=0
cc_743 N_A_416_118#_c_1236_n N_VGND_c_1433_n 0.0221125f $X=2.975 $Y=0.535 $X2=0
+ $Y2=0
cc_744 N_A_416_118#_c_1237_n N_VGND_c_1433_n 0.00765673f $X=2.385 $Y=0.535 $X2=0
+ $Y2=0
cc_745 N_X_c_1356_n N_VGND_c_1420_n 0.0283319f $X=8.995 $Y=0.515 $X2=0 $Y2=0
cc_746 N_X_c_1356_n N_VGND_c_1421_n 0.0144922f $X=8.995 $Y=0.515 $X2=0 $Y2=0
cc_747 N_X_c_1356_n N_VGND_c_1422_n 0.0291466f $X=8.995 $Y=0.515 $X2=0 $Y2=0
cc_748 N_X_c_1373_n N_VGND_c_1422_n 0.0135557f $X=9.665 $Y=1.385 $X2=0 $Y2=0
cc_749 N_X_c_1358_n N_VGND_c_1422_n 0.0281649f $X=9.855 $Y=0.515 $X2=0 $Y2=0
cc_750 N_X_c_1358_n N_VGND_c_1424_n 0.0294122f $X=9.855 $Y=0.515 $X2=0 $Y2=0
cc_751 N_X_c_1358_n N_VGND_c_1429_n 0.0109942f $X=9.855 $Y=0.515 $X2=0 $Y2=0
cc_752 N_X_c_1356_n N_VGND_c_1433_n 0.0118826f $X=8.995 $Y=0.515 $X2=0 $Y2=0
cc_753 N_X_c_1358_n N_VGND_c_1433_n 0.00904371f $X=9.855 $Y=0.515 $X2=0 $Y2=0
