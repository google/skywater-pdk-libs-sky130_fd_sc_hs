# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_hs__clkbuf_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__clkbuf_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  1.920000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.231000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.085000 1.010000 1.495000 2.150000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  0.453600 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.545000 0.350000 0.885000 0.790000 ;
        RECT 0.555000 1.820000 0.885000 2.150000 ;
        RECT 0.715000 0.790000 0.885000 1.820000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 1.920000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 1.920000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 1.920000 0.085000 ;
      RECT 0.000000  3.245000 1.920000 3.415000 ;
      RECT 0.105000  2.660000 0.435000 3.245000 ;
      RECT 0.115000  0.085000 0.365000 0.790000 ;
      RECT 0.215000  0.960000 0.545000 1.630000 ;
      RECT 0.215000  1.630000 0.385000 2.320000 ;
      RECT 0.215000  2.320000 1.835000 2.490000 ;
      RECT 1.005000  2.660000 1.335000 3.245000 ;
      RECT 1.055000  0.085000 1.305000 0.810000 ;
      RECT 1.475000  0.350000 1.835000 0.810000 ;
      RECT 1.535000  2.490000 1.835000 2.980000 ;
      RECT 1.665000  0.810000 1.835000 2.320000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
  END
END sky130_fd_sc_hs__clkbuf_2
END LIBRARY
