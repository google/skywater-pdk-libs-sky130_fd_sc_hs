* File: sky130_fd_sc_hs__dlxtn_4.spice
* Created: Thu Aug 27 20:42:51 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hs__dlxtn_4.pex.spice"
.subckt sky130_fd_sc_hs__dlxtn_4  VNB VPB D GATE_N VPWR Q VGND
* 
* VGND	VGND
* Q	Q
* VPWR	VPWR
* GATE_N	GATE_N
* D	D
* VPB	VPB
* VNB	VNB
MM1011 N_VGND_M1011_d N_D_M1011_g N_A_27_115#_M1011_s VNB NLOWVT L=0.15 W=0.55
+ AD=0.171896 AS=0.15675 PD=1.33876 PS=1.67 NRD=56.184 NRS=0 M=1 R=3.66667
+ SA=75000.2 SB=75000.8 A=0.0825 P=1.4 MULT=1
MM1017 N_A_230_424#_M1017_d N_GATE_N_M1017_g N_VGND_M1011_d VNB NLOWVT L=0.15
+ W=0.74 AD=0.2109 AS=0.231279 PD=2.05 PS=1.80124 NRD=0 NRS=41.76 M=1 R=4.93333
+ SA=75000.6 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1007 N_VGND_M1007_d N_A_230_424#_M1007_g N_A_369_392#_M1007_s VNB NLOWVT
+ L=0.15 W=0.74 AD=0.25707 AS=0.2109 PD=1.55507 PS=2.05 NRD=66.48 NRS=0 M=1
+ R=4.93333 SA=75000.2 SB=75003.6 A=0.111 P=1.78 MULT=1
MM1002 A_658_79# N_A_27_115#_M1002_g N_VGND_M1007_d VNB NLOWVT L=0.15 W=0.64
+ AD=0.0768 AS=0.22233 PD=0.88 PS=1.34493 NRD=12.18 NRS=3.744 M=1 R=4.26667
+ SA=75001.1 SB=75003.3 A=0.096 P=1.58 MULT=1
MM1001 N_A_675_392#_M1001_d N_A_230_424#_M1001_g A_658_79# VNB NLOWVT L=0.15
+ W=0.64 AD=0.19677 AS=0.0768 PD=1.5517 PS=0.88 NRD=0 NRS=12.18 M=1 R=4.26667
+ SA=75001.5 SB=75002.9 A=0.096 P=1.58 MULT=1
MM1010 A_895_123# N_A_369_392#_M1010_g N_A_675_392#_M1001_d VNB NLOWVT L=0.15
+ W=0.42 AD=0.0441 AS=0.12913 PD=0.63 PS=1.0183 NRD=14.28 NRS=0 M=1 R=2.8
+ SA=75002.3 SB=75003.5 A=0.063 P=1.14 MULT=1
MM1005 N_VGND_M1005_d N_A_840_395#_M1005_g A_895_123# VNB NLOWVT L=0.15 W=0.42
+ AD=0.0817019 AS=0.0441 PD=0.792453 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8
+ SA=75002.6 SB=75003.1 A=0.063 P=1.14 MULT=1
MM1009 N_VGND_M1005_d N_A_675_392#_M1009_g N_A_840_395#_M1009_s VNB NLOWVT
+ L=0.15 W=0.64 AD=0.124498 AS=0.0896 PD=1.20755 PS=0.92 NRD=14.988 NRS=0 M=1
+ R=4.26667 SA=75002.1 SB=75002.6 A=0.096 P=1.58 MULT=1
MM1024 N_VGND_M1024_d N_A_675_392#_M1024_g N_A_840_395#_M1009_s VNB NLOWVT
+ L=0.15 W=0.64 AD=0.11993 AS=0.0896 PD=1.02493 PS=0.92 NRD=0 NRS=0 M=1
+ R=4.26667 SA=75002.5 SB=75002.2 A=0.096 P=1.58 MULT=1
MM1013 N_Q_M1013_d N_A_840_395#_M1013_g N_VGND_M1024_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.1369 AS=0.13867 PD=1.11 PS=1.18507 NRD=1.62 NRS=13.776 M=1 R=4.93333
+ SA=75002.7 SB=75001.7 A=0.111 P=1.78 MULT=1
MM1016 N_Q_M1013_d N_A_840_395#_M1016_g N_VGND_M1016_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1369 AS=0.1036 PD=1.11 PS=1.02 NRD=12.972 NRS=0 M=1 R=4.93333 SA=75003.2
+ SB=75001.1 A=0.111 P=1.78 MULT=1
MM1023 N_Q_M1023_d N_A_840_395#_M1023_g N_VGND_M1016_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.12025 AS=0.1036 PD=1.065 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75003.6
+ SB=75000.7 A=0.111 P=1.78 MULT=1
MM1025 N_Q_M1023_d N_A_840_395#_M1025_g N_VGND_M1025_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.12025 AS=0.2294 PD=1.065 PS=2.1 NRD=7.296 NRS=4.044 M=1 R=4.93333
+ SA=75004.1 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1004 N_VPWR_M1004_d N_D_M1004_g N_A_27_115#_M1004_s VPB PSHORT L=0.15 W=0.84
+ AD=0.168 AS=0.2478 PD=1.24 PS=2.27 NRD=14.0658 NRS=2.3443 M=1 R=5.6 SA=75000.2
+ SB=75000.8 A=0.126 P=1.98 MULT=1
MM1019 N_A_230_424#_M1019_d N_GATE_N_M1019_g N_VPWR_M1004_d VPB PSHORT L=0.15
+ W=0.84 AD=0.2478 AS=0.168 PD=2.27 PS=1.24 NRD=2.3443 NRS=14.0658 M=1 R=5.6
+ SA=75000.8 SB=75000.2 A=0.126 P=1.98 MULT=1
MM1006 N_VPWR_M1006_d N_A_230_424#_M1006_g N_A_369_392#_M1006_s VPB PSHORT
+ L=0.15 W=0.84 AD=0.228535 AS=0.2478 PD=1.38326 PS=2.27 NRD=38.6908 NRS=2.3443
+ M=1 R=5.6 SA=75000.2 SB=75002.7 A=0.126 P=1.98 MULT=1
MM1014 A_591_392# N_A_27_115#_M1014_g N_VPWR_M1006_d VPB PSHORT L=0.15 W=1
+ AD=0.135 AS=0.272065 PD=1.27 PS=1.64674 NRD=15.7403 NRS=14.7553 M=1 R=6.66667
+ SA=75000.8 SB=75002.5 A=0.15 P=2.3 MULT=1
MM1018 N_A_675_392#_M1018_d N_A_369_392#_M1018_g A_591_392# VPB PSHORT L=0.15
+ W=1 AD=0.244718 AS=0.135 PD=2 PS=1.27 NRD=1.9503 NRS=15.7403 M=1 R=6.66667
+ SA=75001.2 SB=75002 A=0.15 P=2.3 MULT=1
MM1008 A_789_508# N_A_230_424#_M1008_g N_A_675_392#_M1018_d VPB PSHORT L=0.15
+ W=0.42 AD=0.0567 AS=0.102782 PD=0.69 PS=0.84 NRD=37.5088 NRS=63.3158 M=1 R=2.8
+ SA=75001.7 SB=75004 A=0.063 P=1.14 MULT=1
MM1020 N_VPWR_M1020_d N_A_840_395#_M1020_g A_789_508# VPB PSHORT L=0.15 W=0.42
+ AD=0.1463 AS=0.0567 PD=1.08 PS=0.69 NRD=7.0329 NRS=37.5088 M=1 R=2.8
+ SA=75002.1 SB=75003.6 A=0.063 P=1.14 MULT=1
MM1012 N_A_840_395#_M1012_d N_A_675_392#_M1012_g N_VPWR_M1020_d VPB PSHORT
+ L=0.15 W=0.84 AD=0.1491 AS=0.2926 PD=1.195 PS=2.16 NRD=10.5395 NRS=5.8509 M=1
+ R=5.6 SA=75001.6 SB=75002.7 A=0.126 P=1.98 MULT=1
MM1015 N_A_840_395#_M1012_d N_A_675_392#_M1015_g N_VPWR_M1015_s VPB PSHORT
+ L=0.15 W=0.84 AD=0.1491 AS=0.1596 PD=1.195 PS=1.26429 NRD=7.0329 NRS=9.3772
+ M=1 R=5.6 SA=75002.1 SB=75002.1 A=0.126 P=1.98 MULT=1
MM1000 N_VPWR_M1015_s N_A_840_395#_M1000_g N_Q_M1000_s VPB PSHORT L=0.15 W=1.12
+ AD=0.2128 AS=0.21 PD=1.68571 PS=1.495 NRD=6.1464 NRS=6.1464 M=1 R=7.46667
+ SA=75002 SB=75001.6 A=0.168 P=2.54 MULT=1
MM1003 N_VPWR_M1003_d N_A_840_395#_M1003_g N_Q_M1000_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.21 PD=1.42 PS=1.495 NRD=1.7533 NRS=10.5395 M=1 R=7.46667
+ SA=75002.5 SB=75001.1 A=0.168 P=2.54 MULT=1
MM1021 N_VPWR_M1003_d N_A_840_395#_M1021_g N_Q_M1021_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667 SA=75003
+ SB=75000.7 A=0.168 P=2.54 MULT=1
MM1022 N_VPWR_M1022_d N_A_840_395#_M1022_g N_Q_M1021_s VPB PSHORT L=0.15 W=1.12
+ AD=0.3304 AS=0.168 PD=2.83 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75003.4 SB=75000.2 A=0.168 P=2.54 MULT=1
DX26_noxref VNB VPB NWDIODE A=15.8844 P=20.8
c_86 VNB 0 9.68457e-20 $X=0 $Y=0
c_951 A_591_392# 0 1.00461e-19 $X=2.955 $Y=1.96
c_1140 A_658_79# 0 1.82656e-20 $X=3.29 $Y=0.395
*
.include "sky130_fd_sc_hs__dlxtn_4.pxi.spice"
*
.ends
*
*
