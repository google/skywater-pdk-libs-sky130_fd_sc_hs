* File: sky130_fd_sc_hs__o221ai_2.pex.spice
* Created: Tue Sep  1 20:15:51 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HS__O221AI_2%C1 3 5 7 10 12 14 15 19 22
r43 22 23 9.16848 $w=3.68e-07 $l=7e-08 $layer=POLY_cond $X=0.925 $Y=1.532
+ $X2=0.995 $Y2=1.532
r44 21 22 49.7717 $w=3.68e-07 $l=3.8e-07 $layer=POLY_cond $X=0.545 $Y=1.532
+ $X2=0.925 $Y2=1.532
r45 20 21 6.54891 $w=3.68e-07 $l=5e-08 $layer=POLY_cond $X=0.495 $Y=1.532
+ $X2=0.545 $Y2=1.532
r46 18 20 29.4701 $w=3.68e-07 $l=2.25e-07 $layer=POLY_cond $X=0.27 $Y=1.532
+ $X2=0.495 $Y2=1.532
r47 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.27
+ $Y=1.465 $X2=0.27 $Y2=1.465
r48 15 19 6.9845 $w=3.28e-07 $l=2e-07 $layer=LI1_cond $X=0.27 $Y=1.665 $X2=0.27
+ $Y2=1.465
r49 12 23 23.8357 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=0.995 $Y=1.765
+ $X2=0.995 $Y2=1.532
r50 12 14 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.995 $Y=1.765
+ $X2=0.995 $Y2=2.4
r51 8 22 23.8357 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=0.925 $Y=1.3
+ $X2=0.925 $Y2=1.532
r52 8 10 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=0.925 $Y=1.3
+ $X2=0.925 $Y2=0.74
r53 5 21 23.8357 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=0.545 $Y=1.765
+ $X2=0.545 $Y2=1.532
r54 5 7 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.545 $Y=1.765
+ $X2=0.545 $Y2=2.4
r55 1 20 23.8357 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=0.495 $Y=1.3
+ $X2=0.495 $Y2=1.532
r56 1 3 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=0.495 $Y=1.3 $X2=0.495
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HS__O221AI_2%B1 1 3 4 6 7 9 12 14 18 21 22 23 39
c83 12 0 1.19923e-19 $X=3.33 $Y=0.795
c84 7 0 8.34958e-20 $X=3.255 $Y=1.765
c85 1 0 2.73477e-19 $X=1.805 $Y=1.765
r86 28 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.795
+ $Y=1.515 $X2=1.795 $Y2=1.515
r87 23 39 10.4716 $w=7.68e-07 $l=1.15e-07 $layer=LI1_cond $X=2.16 $Y=1.735
+ $X2=2.275 $Y2=1.735
r88 23 29 5.66972 $w=7.68e-07 $l=3.65e-07 $layer=LI1_cond $X=2.16 $Y=1.735
+ $X2=1.795 $Y2=1.735
r89 22 29 1.78635 $w=7.68e-07 $l=1.15e-07 $layer=LI1_cond $X=1.68 $Y=1.735
+ $X2=1.795 $Y2=1.735
r90 21 22 7.45607 $w=7.68e-07 $l=4.8e-07 $layer=LI1_cond $X=1.2 $Y=1.735
+ $X2=1.68 $Y2=1.735
r91 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.24
+ $Y=1.515 $X2=3.24 $Y2=1.515
r92 16 18 15.1913 $w=3.28e-07 $l=4.35e-07 $layer=LI1_cond $X=3.24 $Y=1.95
+ $X2=3.24 $Y2=1.515
r93 14 16 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.075 $Y=2.035
+ $X2=3.24 $Y2=1.95
r94 14 39 52.1925 $w=1.68e-07 $l=8e-07 $layer=LI1_cond $X=3.075 $Y=2.035
+ $X2=2.275 $Y2=2.035
r95 10 19 38.5562 $w=2.99e-07 $l=2.05122e-07 $layer=POLY_cond $X=3.33 $Y=1.35
+ $X2=3.24 $Y2=1.515
r96 10 12 284.585 $w=1.5e-07 $l=5.55e-07 $layer=POLY_cond $X=3.33 $Y=1.35
+ $X2=3.33 $Y2=0.795
r97 7 19 52.2586 $w=2.99e-07 $l=2.57391e-07 $layer=POLY_cond $X=3.255 $Y=1.765
+ $X2=3.24 $Y2=1.515
r98 7 9 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.255 $Y=1.765
+ $X2=3.255 $Y2=2.4
r99 4 28 47.8017 $w=3.12e-07 $l=2.72489e-07 $layer=POLY_cond $X=1.915 $Y=1.29
+ $X2=1.81 $Y2=1.515
r100 4 6 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=1.915 $Y=1.29
+ $X2=1.915 $Y2=0.795
r101 1 28 51.6639 $w=3.12e-07 $l=2.52488e-07 $layer=POLY_cond $X=1.805 $Y=1.765
+ $X2=1.81 $Y2=1.515
r102 1 3 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.805 $Y=1.765
+ $X2=1.805 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_HS__O221AI_2%B2 1 3 6 8 10 13 15 21 22
c51 21 0 1.93102e-19 $X=2.685 $Y=1.515
r52 22 23 2.70028 $w=3.57e-07 $l=2e-08 $layer=POLY_cond $X=2.755 $Y=1.557
+ $X2=2.775 $Y2=1.557
r53 20 22 9.45098 $w=3.57e-07 $l=7e-08 $layer=POLY_cond $X=2.685 $Y=1.557
+ $X2=2.755 $Y2=1.557
r54 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.685
+ $Y=1.515 $X2=2.685 $Y2=1.515
r55 18 20 45.9048 $w=3.57e-07 $l=3.4e-07 $layer=POLY_cond $X=2.345 $Y=1.557
+ $X2=2.685 $Y2=1.557
r56 17 18 7.42577 $w=3.57e-07 $l=5.5e-08 $layer=POLY_cond $X=2.29 $Y=1.557
+ $X2=2.345 $Y2=1.557
r57 15 21 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=2.685 $Y=1.665
+ $X2=2.685 $Y2=1.515
r58 11 23 23.1043 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.775 $Y=1.35
+ $X2=2.775 $Y2=1.557
r59 11 13 284.585 $w=1.5e-07 $l=5.55e-07 $layer=POLY_cond $X=2.775 $Y=1.35
+ $X2=2.775 $Y2=0.795
r60 8 22 23.1043 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=2.755 $Y=1.765
+ $X2=2.755 $Y2=1.557
r61 8 10 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.755 $Y=1.765
+ $X2=2.755 $Y2=2.4
r62 4 18 23.1043 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.345 $Y=1.35
+ $X2=2.345 $Y2=1.557
r63 4 6 284.585 $w=1.5e-07 $l=5.55e-07 $layer=POLY_cond $X=2.345 $Y=1.35
+ $X2=2.345 $Y2=0.795
r64 1 17 23.1043 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=2.29 $Y=1.765
+ $X2=2.29 $Y2=1.557
r65 1 3 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.29 $Y=1.765
+ $X2=2.29 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_HS__O221AI_2%A1 3 5 7 8 10 13 17 20 21 22 29
c80 5 0 8.35221e-20 $X=3.805 $Y=1.765
c81 3 0 2.04231e-19 $X=3.76 $Y=0.795
r82 28 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.28
+ $Y=1.515 $X2=5.28 $Y2=1.515
r83 22 35 6.23308 $w=7.08e-07 $l=3.7e-07 $layer=LI1_cond $X=5.28 $Y=1.665
+ $X2=5.28 $Y2=2.035
r84 22 29 2.52693 $w=7.08e-07 $l=1.5e-07 $layer=LI1_cond $X=5.28 $Y=1.665
+ $X2=5.28 $Y2=1.515
r85 20 35 9.41505 $w=1.7e-07 $l=3.55e-07 $layer=LI1_cond $X=4.925 $Y=2.035
+ $X2=5.28 $Y2=2.035
r86 20 21 61.9786 $w=1.68e-07 $l=9.5e-07 $layer=LI1_cond $X=4.925 $Y=2.035
+ $X2=3.975 $Y2=2.035
r87 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.81
+ $Y=1.515 $X2=3.81 $Y2=1.515
r88 15 21 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.81 $Y=1.95
+ $X2=3.975 $Y2=2.035
r89 15 17 15.1913 $w=3.28e-07 $l=4.35e-07 $layer=LI1_cond $X=3.81 $Y=1.95
+ $X2=3.81 $Y2=1.515
r90 11 28 38.5562 $w=2.99e-07 $l=1.74714e-07 $layer=POLY_cond $X=5.26 $Y=1.35
+ $X2=5.28 $Y2=1.515
r91 11 13 284.585 $w=1.5e-07 $l=5.55e-07 $layer=POLY_cond $X=5.26 $Y=1.35
+ $X2=5.26 $Y2=0.795
r92 8 28 52.2586 $w=2.99e-07 $l=2.85044e-07 $layer=POLY_cond $X=5.205 $Y=1.765
+ $X2=5.28 $Y2=1.515
r93 8 10 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=5.205 $Y=1.765
+ $X2=5.205 $Y2=2.4
r94 5 18 52.2586 $w=2.99e-07 $l=2.52488e-07 $layer=POLY_cond $X=3.805 $Y=1.765
+ $X2=3.81 $Y2=1.515
r95 5 7 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.805 $Y=1.765
+ $X2=3.805 $Y2=2.4
r96 1 18 38.5562 $w=2.99e-07 $l=1.88348e-07 $layer=POLY_cond $X=3.76 $Y=1.35
+ $X2=3.81 $Y2=1.515
r97 1 3 284.585 $w=1.5e-07 $l=5.55e-07 $layer=POLY_cond $X=3.76 $Y=1.35 $X2=3.76
+ $Y2=0.795
.ends

.subckt PM_SKY130_FD_SC_HS__O221AI_2%A2 3 5 7 8 10 13 15 21 22
r54 22 23 1.9127 $w=3.78e-07 $l=1.5e-08 $layer=POLY_cond $X=4.755 $Y=1.557
+ $X2=4.77 $Y2=1.557
r55 20 22 31.2407 $w=3.78e-07 $l=2.45e-07 $layer=POLY_cond $X=4.51 $Y=1.557
+ $X2=4.755 $Y2=1.557
r56 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.51
+ $Y=1.515 $X2=4.51 $Y2=1.515
r57 18 20 26.1402 $w=3.78e-07 $l=2.05e-07 $layer=POLY_cond $X=4.305 $Y=1.557
+ $X2=4.51 $Y2=1.557
r58 17 18 1.9127 $w=3.78e-07 $l=1.5e-08 $layer=POLY_cond $X=4.29 $Y=1.557
+ $X2=4.305 $Y2=1.557
r59 15 21 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=4.51 $Y=1.665
+ $X2=4.51 $Y2=1.515
r60 11 23 24.4846 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.77 $Y=1.35
+ $X2=4.77 $Y2=1.557
r61 11 13 284.585 $w=1.5e-07 $l=5.55e-07 $layer=POLY_cond $X=4.77 $Y=1.35
+ $X2=4.77 $Y2=0.795
r62 8 22 24.4846 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=4.755 $Y=1.765
+ $X2=4.755 $Y2=1.557
r63 8 10 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=4.755 $Y=1.765
+ $X2=4.755 $Y2=2.4
r64 5 18 24.4846 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=4.305 $Y=1.765
+ $X2=4.305 $Y2=1.557
r65 5 7 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=4.305 $Y=1.765
+ $X2=4.305 $Y2=2.4
r66 1 17 24.4846 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.29 $Y=1.35
+ $X2=4.29 $Y2=1.557
r67 1 3 284.585 $w=1.5e-07 $l=5.55e-07 $layer=POLY_cond $X=4.29 $Y=1.35 $X2=4.29
+ $Y2=0.795
.ends

.subckt PM_SKY130_FD_SC_HS__O221AI_2%VPWR 1 2 3 4 13 15 21 23 25 27 29 34 39 51
+ 60 64
r71 63 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r72 60 61 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r73 55 57 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=1.68 $Y2=3.33
r74 54 57 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r75 54 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r76 51 54 9.99847 $w=6.38e-07 $l=5.35e-07 $layer=LI1_cond $X=1.375 $Y=2.795
+ $X2=1.375 $Y2=3.33
r77 48 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r78 46 64 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=5.52 $Y2=3.33
r79 45 46 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r80 43 46 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=5.04 $Y2=3.33
r81 43 61 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=3.6 $Y2=3.33
r82 42 45 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=4.08 $Y=3.33 $X2=5.04
+ $Y2=3.33
r83 42 43 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r84 40 60 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.695 $Y=3.33
+ $X2=3.53 $Y2=3.33
r85 40 42 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=3.695 $Y=3.33
+ $X2=4.08 $Y2=3.33
r86 39 63 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=5.315 $Y=3.33
+ $X2=5.537 $Y2=3.33
r87 39 45 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=5.315 $Y=3.33
+ $X2=5.04 $Y2=3.33
r88 38 61 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=3.6 $Y2=3.33
r89 37 38 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r90 35 54 8.73481 $w=1.7e-07 $l=3.2e-07 $layer=LI1_cond $X=1.695 $Y=3.33
+ $X2=1.375 $Y2=3.33
r91 35 37 92.9679 $w=1.68e-07 $l=1.425e-06 $layer=LI1_cond $X=1.695 $Y=3.33
+ $X2=3.12 $Y2=3.33
r92 34 60 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.365 $Y=3.33
+ $X2=3.53 $Y2=3.33
r93 34 37 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=3.365 $Y=3.33
+ $X2=3.12 $Y2=3.33
r94 33 55 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r95 33 49 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r96 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r97 30 48 3.96192 $w=1.7e-07 $l=2.03e-07 $layer=LI1_cond $X=0.405 $Y=3.33
+ $X2=0.202 $Y2=3.33
r98 30 32 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=0.405 $Y=3.33
+ $X2=0.72 $Y2=3.33
r99 29 54 8.73481 $w=1.7e-07 $l=3.2e-07 $layer=LI1_cond $X=1.055 $Y=3.33
+ $X2=1.375 $Y2=3.33
r100 29 32 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=1.055 $Y=3.33
+ $X2=0.72 $Y2=3.33
r101 27 38 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.88 $Y=3.33
+ $X2=3.12 $Y2=3.33
r102 27 57 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=2.88 $Y=3.33
+ $X2=1.68 $Y2=3.33
r103 23 63 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=5.48 $Y=3.245
+ $X2=5.537 $Y2=3.33
r104 23 25 27.5888 $w=3.28e-07 $l=7.9e-07 $layer=LI1_cond $X=5.48 $Y=3.245
+ $X2=5.48 $Y2=2.455
r105 19 60 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.53 $Y=3.245
+ $X2=3.53 $Y2=3.33
r106 19 21 15.3659 $w=3.28e-07 $l=4.4e-07 $layer=LI1_cond $X=3.53 $Y=3.245
+ $X2=3.53 $Y2=2.805
r107 15 18 32.2684 $w=2.48e-07 $l=7e-07 $layer=LI1_cond $X=0.28 $Y=2.115
+ $X2=0.28 $Y2=2.815
r108 13 48 3.18124 $w=2.5e-07 $l=1.17707e-07 $layer=LI1_cond $X=0.28 $Y=3.245
+ $X2=0.202 $Y2=3.33
r109 13 18 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=0.28 $Y=3.245
+ $X2=0.28 $Y2=2.815
r110 4 25 300 $w=1.7e-07 $l=7.07972e-07 $layer=licon1_PDIFF $count=2 $X=5.28
+ $Y=1.84 $X2=5.48 $Y2=2.455
r111 3 21 600 $w=1.7e-07 $l=1.06029e-06 $layer=licon1_PDIFF $count=1 $X=3.33
+ $Y=1.84 $X2=3.53 $Y2=2.805
r112 2 51 300 $w=1.7e-07 $l=1.18282e-06 $layer=licon1_PDIFF $count=2 $X=1.07
+ $Y=1.84 $X2=1.58 $Y2=2.795
r113 1 18 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=0.175
+ $Y=1.84 $X2=0.32 $Y2=2.815
r114 1 15 400 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_PDIFF $count=1 $X=0.175
+ $Y=1.84 $X2=0.32 $Y2=2.115
.ends

.subckt PM_SKY130_FD_SC_HS__O221AI_2%Y 1 2 3 4 15 17 22 23 24 25 26 27 28 29
r61 28 37 3.58051 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=0.74 $Y=2.375
+ $X2=0.74 $Y2=2.29
r62 28 49 3.58051 $w=2.6e-07 $l=8.9861e-08 $layer=LI1_cond $X=0.74 $Y=2.375
+ $X2=0.73 $Y2=2.46
r63 28 29 13.8293 $w=2.48e-07 $l=3e-07 $layer=LI1_cond $X=0.73 $Y=2.475 $X2=0.73
+ $Y2=2.775
r64 28 49 0.691466 $w=2.48e-07 $l=1.5e-08 $layer=LI1_cond $X=0.73 $Y=2.475
+ $X2=0.73 $Y2=2.46
r65 27 37 13.0183 $w=2.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.74 $Y=1.985
+ $X2=0.74 $Y2=2.29
r66 26 27 13.6586 $w=2.68e-07 $l=3.2e-07 $layer=LI1_cond $X=0.74 $Y=1.665
+ $X2=0.74 $Y2=1.985
r67 25 26 15.7927 $w=2.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.74 $Y=1.295
+ $X2=0.74 $Y2=1.665
r68 24 25 18.5671 $w=2.68e-07 $l=4.35e-07 $layer=LI1_cond $X=0.74 $Y=0.86
+ $X2=0.74 $Y2=1.295
r69 21 23 8.86124 $w=4.43e-07 $l=1.65e-07 $layer=LI1_cond $X=2.53 $Y=2.512
+ $X2=2.695 $Y2=2.512
r70 21 22 8.86124 $w=4.43e-07 $l=1.65e-07 $layer=LI1_cond $X=2.53 $Y=2.512
+ $X2=2.365 $Y2=2.512
r71 17 19 2.44 $w=2.5e-07 $l=5e-08 $layer=LI1_cond $X=4.49 $Y=2.46 $X2=4.49
+ $Y2=2.51
r72 15 17 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=4.365 $Y=2.375
+ $X2=4.49 $Y2=2.46
r73 15 23 108.952 $w=1.68e-07 $l=1.67e-06 $layer=LI1_cond $X=4.365 $Y=2.375
+ $X2=2.695 $Y2=2.375
r74 14 28 2.90867 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=0.875 $Y=2.375
+ $X2=0.74 $Y2=2.375
r75 14 22 97.2086 $w=1.68e-07 $l=1.49e-06 $layer=LI1_cond $X=0.875 $Y=2.375
+ $X2=2.365 $Y2=2.375
r76 4 19 600 $w=1.7e-07 $l=7.41215e-07 $layer=licon1_PDIFF $count=1 $X=4.38
+ $Y=1.84 $X2=4.53 $Y2=2.51
r77 3 21 600 $w=1.7e-07 $l=7.47964e-07 $layer=licon1_PDIFF $count=1 $X=2.365
+ $Y=1.84 $X2=2.53 $Y2=2.51
r78 2 28 300 $w=1.7e-07 $l=6.30555e-07 $layer=licon1_PDIFF $count=2 $X=0.62
+ $Y=1.84 $X2=0.77 $Y2=2.4
r79 2 27 600 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=0.62
+ $Y=1.84 $X2=0.77 $Y2=1.985
r80 1 24 182 $w=1.7e-07 $l=5.55608e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.37 $X2=0.71 $Y2=0.86
.ends

.subckt PM_SKY130_FD_SC_HS__O221AI_2%A_376_368# 1 2 7 10 15
c28 7 0 1.63872e-19 $X=2.865 $Y=2.99
r29 15 17 6.46067 $w=3.28e-07 $l=1.85e-07 $layer=LI1_cond $X=3.03 $Y=2.805
+ $X2=3.03 $Y2=2.99
r30 10 12 6.46067 $w=3.28e-07 $l=1.85e-07 $layer=LI1_cond $X=2.03 $Y=2.805
+ $X2=2.03 $Y2=2.99
r31 8 12 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.195 $Y=2.99
+ $X2=2.03 $Y2=2.99
r32 7 17 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.865 $Y=2.99
+ $X2=3.03 $Y2=2.99
r33 7 8 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.865 $Y=2.99
+ $X2=2.195 $Y2=2.99
r34 2 15 600 $w=1.7e-07 $l=1.06029e-06 $layer=licon1_PDIFF $count=1 $X=2.83
+ $Y=1.84 $X2=3.03 $Y2=2.805
r35 1 10 600 $w=1.7e-07 $l=1.03729e-06 $layer=licon1_PDIFF $count=1 $X=1.88
+ $Y=1.84 $X2=2.03 $Y2=2.805
.ends

.subckt PM_SKY130_FD_SC_HS__O221AI_2%A_776_368# 1 2 7 11 14
c30 7 0 8.35221e-20 $X=4.815 $Y=2.99
r31 14 16 6.46067 $w=3.28e-07 $l=1.85e-07 $layer=LI1_cond $X=4.03 $Y=2.805
+ $X2=4.03 $Y2=2.99
r32 9 11 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=4.98 $Y=2.905
+ $X2=4.98 $Y2=2.455
r33 8 16 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.195 $Y=2.99
+ $X2=4.03 $Y2=2.99
r34 7 9 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.815 $Y=2.99
+ $X2=4.98 $Y2=2.905
r35 7 8 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=4.815 $Y=2.99
+ $X2=4.195 $Y2=2.99
r36 2 11 300 $w=1.7e-07 $l=6.85912e-07 $layer=licon1_PDIFF $count=2 $X=4.83
+ $Y=1.84 $X2=4.98 $Y2=2.455
r37 1 14 600 $w=1.7e-07 $l=1.03729e-06 $layer=licon1_PDIFF $count=1 $X=3.88
+ $Y=1.84 $X2=4.03 $Y2=2.805
.ends

.subckt PM_SKY130_FD_SC_HS__O221AI_2%A_27_74# 1 2 3 4 15 17 18 22 23 24 27 29 33
+ 35
c51 33 0 1.48041e-19 $X=3.085 $Y=0.68
c52 29 0 5.61893e-20 $X=2.895 $Y=1.095
r53 31 33 9.87808 $w=3.83e-07 $l=3.3e-07 $layer=LI1_cond $X=3.087 $Y=1.01
+ $X2=3.087 $Y2=0.68
r54 30 35 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.215 $Y=1.095
+ $X2=2.13 $Y2=1.095
r55 29 31 8.24022 $w=1.7e-07 $l=2.30617e-07 $layer=LI1_cond $X=2.895 $Y=1.095
+ $X2=3.087 $Y2=1.01
r56 29 30 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=2.895 $Y=1.095
+ $X2=2.215 $Y2=1.095
r57 25 35 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.13 $Y=1.01 $X2=2.13
+ $Y2=1.095
r58 25 27 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=2.13 $Y=1.01
+ $X2=2.13 $Y2=0.885
r59 23 35 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.045 $Y=1.095
+ $X2=2.13 $Y2=1.095
r60 23 24 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=2.045 $Y=1.095
+ $X2=1.305 $Y2=1.095
r61 20 24 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.18 $Y=1.01
+ $X2=1.305 $Y2=1.095
r62 20 22 22.8184 $w=2.48e-07 $l=4.95e-07 $layer=LI1_cond $X=1.18 $Y=1.01
+ $X2=1.18 $Y2=0.515
r63 19 22 4.14879 $w=2.48e-07 $l=9e-08 $layer=LI1_cond $X=1.18 $Y=0.425 $X2=1.18
+ $Y2=0.515
r64 17 19 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.055 $Y=0.34
+ $X2=1.18 $Y2=0.425
r65 17 18 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.055 $Y=0.34
+ $X2=0.365 $Y2=0.34
r66 13 18 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.24 $Y=0.425
+ $X2=0.365 $Y2=0.34
r67 13 15 4.14879 $w=2.48e-07 $l=9e-08 $layer=LI1_cond $X=0.24 $Y=0.425 $X2=0.24
+ $Y2=0.515
r68 4 33 91 $w=1.7e-07 $l=3.53483e-07 $layer=licon1_NDIFF $count=2 $X=2.85
+ $Y=0.425 $X2=3.085 $Y2=0.68
r69 3 27 182 $w=1.7e-07 $l=5.25357e-07 $layer=licon1_NDIFF $count=1 $X=1.99
+ $Y=0.425 $X2=2.13 $Y2=0.885
r70 2 22 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1 $Y=0.37
+ $X2=1.14 $Y2=0.515
r71 1 15 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__O221AI_2%A_311_85# 1 2 3 4 5 18 20 21 24 26 31 32 33
+ 36 38 42 44 45
c79 33 0 1.19923e-19 $X=3.71 $Y=1.095
r80 40 42 19.8853 $w=2.53e-07 $l=4.4e-07 $layer=LI1_cond $X=5.517 $Y=1.01
+ $X2=5.517 $Y2=0.57
r81 39 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.71 $Y=1.095
+ $X2=4.545 $Y2=1.095
r82 38 40 7.17723 $w=1.7e-07 $l=1.64085e-07 $layer=LI1_cond $X=5.39 $Y=1.095
+ $X2=5.517 $Y2=1.01
r83 38 39 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=5.39 $Y=1.095
+ $X2=4.71 $Y2=1.095
r84 34 45 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.545 $Y=1.01
+ $X2=4.545 $Y2=1.095
r85 34 36 15.3659 $w=3.28e-07 $l=4.4e-07 $layer=LI1_cond $X=4.545 $Y=1.01
+ $X2=4.545 $Y2=0.57
r86 32 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.38 $Y=1.095
+ $X2=4.545 $Y2=1.095
r87 32 33 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.38 $Y=1.095
+ $X2=3.71 $Y2=1.095
r88 29 33 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=3.585 $Y=1.01
+ $X2=3.71 $Y2=1.095
r89 29 31 20.283 $w=2.48e-07 $l=4.4e-07 $layer=LI1_cond $X=3.585 $Y=1.01
+ $X2=3.585 $Y2=0.57
r90 28 31 6.68417 $w=2.48e-07 $l=1.45e-07 $layer=LI1_cond $X=3.585 $Y=0.425
+ $X2=3.585 $Y2=0.57
r91 27 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.725 $Y=0.34
+ $X2=2.56 $Y2=0.34
r92 26 28 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=3.46 $Y=0.34
+ $X2=3.585 $Y2=0.425
r93 26 27 47.9519 $w=1.68e-07 $l=7.35e-07 $layer=LI1_cond $X=3.46 $Y=0.34
+ $X2=2.725 $Y2=0.34
r94 22 44 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.56 $Y=0.425
+ $X2=2.56 $Y2=0.34
r95 22 24 8.03218 $w=3.28e-07 $l=2.3e-07 $layer=LI1_cond $X=2.56 $Y=0.425
+ $X2=2.56 $Y2=0.655
r96 20 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.395 $Y=0.34
+ $X2=2.56 $Y2=0.34
r97 20 21 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=2.395 $Y=0.34
+ $X2=1.865 $Y2=0.34
r98 16 21 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.7 $Y=0.425
+ $X2=1.865 $Y2=0.34
r99 16 18 8.03218 $w=3.28e-07 $l=2.3e-07 $layer=LI1_cond $X=1.7 $Y=0.425 $X2=1.7
+ $Y2=0.655
r100 5 42 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=5.335
+ $Y=0.425 $X2=5.475 $Y2=0.57
r101 4 36 91 $w=1.7e-07 $l=2.41868e-07 $layer=licon1_NDIFF $count=2 $X=4.365
+ $Y=0.425 $X2=4.545 $Y2=0.57
r102 3 31 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.405
+ $Y=0.425 $X2=3.545 $Y2=0.57
r103 2 24 182 $w=1.7e-07 $l=2.91719e-07 $layer=licon1_NDIFF $count=1 $X=2.42
+ $Y=0.425 $X2=2.56 $Y2=0.655
r104 1 18 182 $w=1.7e-07 $l=2.93684e-07 $layer=licon1_NDIFF $count=1 $X=1.555
+ $Y=0.425 $X2=1.7 $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_HS__O221AI_2%VGND 1 2 9 13 15 17 25 32 33 36 39
r52 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r53 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r54 33 40 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=5.04
+ $Y2=0
r55 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r56 30 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.21 $Y=0 $X2=5.045
+ $Y2=0
r57 30 32 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=5.21 $Y=0 $X2=5.52
+ $Y2=0
r58 29 40 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=5.04
+ $Y2=0
r59 29 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=4.08
+ $Y2=0
r60 28 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r61 26 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.21 $Y=0 $X2=4.045
+ $Y2=0
r62 26 28 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=4.21 $Y=0 $X2=4.56
+ $Y2=0
r63 25 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.88 $Y=0 $X2=5.045
+ $Y2=0
r64 25 28 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=4.88 $Y=0 $X2=4.56
+ $Y2=0
r65 24 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.08
+ $Y2=0
r66 23 24 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r67 19 23 219.209 $w=1.68e-07 $l=3.36e-06 $layer=LI1_cond $X=0.24 $Y=0 $X2=3.6
+ $Y2=0
r68 19 20 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r69 17 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.88 $Y=0 $X2=4.045
+ $Y2=0
r70 17 23 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=3.88 $Y=0 $X2=3.6
+ $Y2=0
r71 15 24 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=2.88 $Y=0 $X2=3.6
+ $Y2=0
r72 15 20 0.73586 $w=4.9e-07 $l=2.64e-06 $layer=MET1_cond $X=2.88 $Y=0 $X2=0.24
+ $Y2=0
r73 11 39 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.045 $Y=0.085
+ $X2=5.045 $Y2=0
r74 11 13 19.9058 $w=3.28e-07 $l=5.7e-07 $layer=LI1_cond $X=5.045 $Y=0.085
+ $X2=5.045 $Y2=0.655
r75 7 36 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.045 $Y=0.085
+ $X2=4.045 $Y2=0
r76 7 9 19.9058 $w=3.28e-07 $l=5.7e-07 $layer=LI1_cond $X=4.045 $Y=0.085
+ $X2=4.045 $Y2=0.655
r77 2 13 182 $w=1.7e-07 $l=3.14484e-07 $layer=licon1_NDIFF $count=1 $X=4.845
+ $Y=0.425 $X2=5.045 $Y2=0.655
r78 1 9 182 $w=1.7e-07 $l=3.18119e-07 $layer=licon1_NDIFF $count=1 $X=3.835
+ $Y=0.425 $X2=4.045 $Y2=0.655
.ends

