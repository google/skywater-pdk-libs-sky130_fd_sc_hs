* NGSPICE file created from sky130_fd_sc_hs__dlrtp_2.ext - technology: sky130A

.subckt sky130_fd_sc_hs__dlrtp_2 D GATE RESET_B VGND VNB VPB VPWR Q
M1000 a_646_74# a_235_74# a_565_392# VPB pshort w=1e+06u l=150000u
+  ad=3.328e+11p pd=2.77e+06u as=2.7e+11p ps=2.54e+06u
M1001 VGND a_235_74# a_347_98# VNB nlowvt w=740000u l=150000u
+  ad=1.38725e+12p pd=1.126e+07u as=2.701e+11p ps=2.21e+06u
M1002 a_568_74# a_27_392# VGND VNB nlowvt w=640000u l=150000u
+  ad=1.536e+11p pd=1.76e+06u as=0p ps=0u
M1003 a_646_74# a_347_98# a_568_74# VNB nlowvt w=640000u l=150000u
+  ad=3.21575e+11p pd=2.36e+06u as=0p ps=0u
M1004 VGND RESET_B a_1060_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=1.776e+11p ps=1.96e+06u
M1005 Q a_832_55# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.146e+11p pd=2.06e+06u as=0p ps=0u
M1006 VPWR D a_27_392# VPB pshort w=840000u l=150000u
+  ad=2.24475e+12p pd=1.588e+07u as=2.478e+11p ps=2.27e+06u
M1007 a_235_74# GATE VPWR VPB pshort w=840000u l=150000u
+  ad=2.478e+11p pd=2.27e+06u as=0p ps=0u
M1008 a_756_508# a_347_98# a_646_74# VPB pshort w=420000u l=150000u
+  ad=2.247e+11p pd=1.91e+06u as=0p ps=0u
M1009 VGND D a_27_392# VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=1.5675e+11p ps=1.67e+06u
M1010 Q a_832_55# VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=3.528e+11p pd=2.87e+06u as=0p ps=0u
M1011 a_832_55# a_646_74# VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=3.36e+11p pd=2.84e+06u as=0p ps=0u
M1012 VPWR RESET_B a_832_55# VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VPWR a_832_55# a_756_508# VPB pshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 VPWR a_235_74# a_347_98# VPB pshort w=840000u l=150000u
+  ad=0p pd=0u as=2.478e+11p ps=2.27e+06u
M1015 VPWR a_832_55# Q VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_1060_74# a_646_74# a_832_55# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1017 a_565_392# a_27_392# VPWR VPB pshort w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 VGND a_832_55# Q VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_784_81# a_235_74# a_646_74# VNB nlowvt w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=0p ps=0u
M1020 VGND a_832_55# a_784_81# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_235_74# GATE VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
.ends

