* File: sky130_fd_sc_hs__a32oi_1.pex.spice
* Created: Thu Aug 27 20:30:18 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HS__A32OI_1%B2 1 3 4 6 7
r21 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.28
+ $Y=1.385 $X2=0.28 $Y2=1.385
r22 7 11 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=0.28 $Y=1.295 $X2=0.28
+ $Y2=1.385
r23 4 10 38.924 $w=3.61e-07 $l=2.33345e-07 $layer=POLY_cond $X=0.52 $Y=1.22
+ $X2=0.355 $Y2=1.385
r24 4 6 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=0.52 $Y=1.22 $X2=0.52
+ $Y2=0.74
r25 1 10 67.6304 $w=3.61e-07 $l=4.48776e-07 $layer=POLY_cond $X=0.505 $Y=1.765
+ $X2=0.355 $Y2=1.385
r26 1 3 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.505 $Y=1.765
+ $X2=0.505 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_HS__A32OI_1%B1 1 3 4 6 7
c28 7 0 1.62524e-19 $X=1.2 $Y=1.295
c29 1 0 1.47908e-19 $X=0.91 $Y=1.22
r30 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.12
+ $Y=1.385 $X2=1.12 $Y2=1.385
r31 7 11 2.88111 $w=3.58e-07 $l=9e-08 $layer=LI1_cond $X=1.135 $Y=1.295
+ $X2=1.135 $Y2=1.385
r32 4 10 68.9212 $w=3.43e-07 $l=4.06571e-07 $layer=POLY_cond $X=1.005 $Y=1.765
+ $X2=1.06 $Y2=1.385
r33 4 6 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.005 $Y=1.765
+ $X2=1.005 $Y2=2.4
r34 1 10 38.7084 $w=3.43e-07 $l=2.2798e-07 $layer=POLY_cond $X=0.91 $Y=1.22
+ $X2=1.06 $Y2=1.385
r35 1 3 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=0.91 $Y=1.22 $X2=0.91
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HS__A32OI_1%A1 1 3 4 6 7
c29 7 0 1.47908e-19 $X=1.68 $Y=1.295
c30 4 0 1.62524e-19 $X=1.88 $Y=1.22
r31 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.69
+ $Y=1.385 $X2=1.69 $Y2=1.385
r32 7 11 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=1.69 $Y=1.295 $X2=1.69
+ $Y2=1.385
r33 4 10 38.6069 $w=3.31e-07 $l=2.24332e-07 $layer=POLY_cond $X=1.88 $Y=1.22
+ $X2=1.74 $Y2=1.385
r34 4 6 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.88 $Y=1.22 $X2=1.88
+ $Y2=0.74
r35 1 10 69.9151 $w=3.31e-07 $l=4.38064e-07 $layer=POLY_cond $X=1.615 $Y=1.765
+ $X2=1.74 $Y2=1.385
r36 1 3 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.615 $Y=1.765
+ $X2=1.615 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_HS__A32OI_1%A2 1 3 4 6 7 8 9
c35 1 0 3.79709e-20 $X=2.27 $Y=1.22
r36 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.36
+ $Y=1.385 $X2=2.36 $Y2=1.385
r37 9 15 2.24265 $w=4.78e-07 $l=9e-08 $layer=LI1_cond $X=2.285 $Y=1.295
+ $X2=2.285 $Y2=1.385
r38 8 9 9.21977 $w=4.78e-07 $l=3.7e-07 $layer=LI1_cond $X=2.285 $Y=0.925
+ $X2=2.285 $Y2=1.295
r39 7 8 9.21977 $w=4.78e-07 $l=3.7e-07 $layer=LI1_cond $X=2.285 $Y=0.555
+ $X2=2.285 $Y2=0.925
r40 4 14 77.2841 $w=2.7e-07 $l=4.01871e-07 $layer=POLY_cond $X=2.405 $Y=1.765
+ $X2=2.36 $Y2=1.385
r41 4 6 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.405 $Y=1.765
+ $X2=2.405 $Y2=2.4
r42 1 14 38.9026 $w=2.7e-07 $l=2.05122e-07 $layer=POLY_cond $X=2.27 $Y=1.22
+ $X2=2.36 $Y2=1.385
r43 1 3 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=2.27 $Y=1.22 $X2=2.27
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HS__A32OI_1%A3 1 3 4 6 7
c24 7 0 3.79709e-20 $X=3.12 $Y=1.295
r25 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.93
+ $Y=1.385 $X2=2.93 $Y2=1.385
r26 7 11 5.91795 $w=3.68e-07 $l=1.9e-07 $layer=LI1_cond $X=3.12 $Y=1.365
+ $X2=2.93 $Y2=1.365
r27 4 10 77.2841 $w=2.7e-07 $l=4.15812e-07 $layer=POLY_cond $X=2.855 $Y=1.765
+ $X2=2.93 $Y2=1.385
r28 4 6 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.855 $Y=1.765
+ $X2=2.855 $Y2=2.4
r29 1 10 38.9026 $w=2.7e-07 $l=2.05122e-07 $layer=POLY_cond $X=2.84 $Y=1.22
+ $X2=2.93 $Y2=1.385
r30 1 3 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=2.84 $Y=1.22 $X2=2.84
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HS__A32OI_1%A_27_368# 1 2 3 12 16 17 18 21 22 26 30 35
r49 33 34 6.99363 $w=3.14e-07 $l=1.8e-07 $layer=LI1_cond $X=1.28 $Y=2.225
+ $X2=1.28 $Y2=2.405
r50 28 35 3.10218 $w=3.05e-07 $l=9.66954e-08 $layer=LI1_cond $X=2.655 $Y=2.49
+ $X2=2.63 $Y2=2.405
r51 28 30 13.3766 $w=2.78e-07 $l=3.25e-07 $layer=LI1_cond $X=2.655 $Y=2.49
+ $X2=2.655 $Y2=2.815
r52 24 35 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.63 $Y=2.32
+ $X2=2.63 $Y2=2.405
r53 24 26 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=2.63 $Y=2.32
+ $X2=2.63 $Y2=1.985
r54 23 34 4.32966 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.445 $Y=2.405
+ $X2=1.28 $Y2=2.405
r55 22 35 3.51065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.465 $Y=2.405
+ $X2=2.63 $Y2=2.405
r56 22 23 66.5455 $w=1.68e-07 $l=1.02e-06 $layer=LI1_cond $X=2.465 $Y=2.405
+ $X2=1.445 $Y2=2.405
r57 19 21 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=1.28 $Y=2.905 $X2=1.28
+ $Y2=2.815
r58 18 34 3.18267 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.28 $Y=2.49 $X2=1.28
+ $Y2=2.405
r59 18 21 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=1.28 $Y=2.49
+ $X2=1.28 $Y2=2.815
r60 16 19 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.115 $Y=2.99
+ $X2=1.28 $Y2=2.905
r61 16 17 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.115 $Y=2.99
+ $X2=0.445 $Y2=2.99
r62 12 15 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=0.28 $Y=1.985
+ $X2=0.28 $Y2=2.815
r63 10 17 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.28 $Y=2.905
+ $X2=0.445 $Y2=2.99
r64 10 15 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=0.28 $Y=2.905 $X2=0.28
+ $Y2=2.815
r65 3 30 600 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=2.48
+ $Y=1.84 $X2=2.63 $Y2=2.815
r66 3 26 300 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=2 $X=2.48
+ $Y=1.84 $X2=2.63 $Y2=1.985
r67 2 33 600 $w=1.7e-07 $l=4.74579e-07 $layer=licon1_PDIFF $count=1 $X=1.08
+ $Y=1.84 $X2=1.28 $Y2=2.225
r68 2 21 600 $w=1.7e-07 $l=1.07034e-06 $layer=licon1_PDIFF $count=1 $X=1.08
+ $Y=1.84 $X2=1.28 $Y2=2.815
r69 1 15 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.815
r70 1 12 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HS__A32OI_1%Y 1 2 8 11 13 15 19 20 23
c48 13 0 1.06273e-19 $X=0.785 $Y=0.68
c49 8 0 1.6439e-20 $X=0.7 $Y=1.72
r50 20 23 19.6393 $w=4.28e-07 $l=5.7e-07 $layer=LI1_cond $X=2.16 $Y=1.935
+ $X2=1.59 $Y2=1.935
r51 18 19 2.76166 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.945 $Y=1.805
+ $X2=0.78 $Y2=1.805
r52 18 23 42.0802 $w=1.68e-07 $l=6.45e-07 $layer=LI1_cond $X=0.945 $Y=1.805
+ $X2=1.59 $Y2=1.805
r53 13 15 15.9477 $w=6.58e-07 $l=8.8e-07 $layer=LI1_cond $X=0.785 $Y=0.68
+ $X2=1.665 $Y2=0.68
r54 9 19 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.78 $Y=1.89 $X2=0.78
+ $Y2=1.805
r55 9 11 3.31764 $w=3.28e-07 $l=9.5e-08 $layer=LI1_cond $X=0.78 $Y=1.89 $X2=0.78
+ $Y2=1.985
r56 8 19 3.70735 $w=2.5e-07 $l=1.18427e-07 $layer=LI1_cond $X=0.7 $Y=1.72
+ $X2=0.78 $Y2=1.805
r57 7 13 10.5067 $w=6.6e-07 $l=3.70068e-07 $layer=LI1_cond $X=0.7 $Y=1.01
+ $X2=0.785 $Y2=0.68
r58 7 8 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=0.7 $Y=1.01 $X2=0.7
+ $Y2=1.72
r59 2 11 300 $w=1.7e-07 $l=2.62678e-07 $layer=licon1_PDIFF $count=2 $X=0.58
+ $Y=1.84 $X2=0.78 $Y2=1.985
r60 1 15 45.5 $w=1.7e-07 $l=7.39865e-07 $layer=licon1_NDIFF $count=4 $X=0.985
+ $Y=0.37 $X2=1.665 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_HS__A32OI_1%VPWR 1 2 7 9 13 15 20 26 36
r40 35 36 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r41 29 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r42 26 29 9.90781 $w=6.68e-07 $l=5.55e-07 $layer=LI1_cond $X=2.01 $Y=2.775
+ $X2=2.01 $Y2=3.33
r43 24 36 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r44 24 32 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=2.16 $Y2=3.33
r45 23 24 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r46 21 29 9.03384 $w=1.7e-07 $l=3.35e-07 $layer=LI1_cond $X=2.345 $Y=3.33
+ $X2=2.01 $Y2=3.33
r47 21 23 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=2.345 $Y=3.33
+ $X2=2.64 $Y2=3.33
r48 20 35 4.01252 $w=1.7e-07 $l=1.82e-07 $layer=LI1_cond $X=2.995 $Y=3.33
+ $X2=3.177 $Y2=3.33
r49 20 23 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=2.995 $Y=3.33
+ $X2=2.64 $Y2=3.33
r50 17 18 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r51 15 29 9.03384 $w=1.7e-07 $l=3.35e-07 $layer=LI1_cond $X=1.675 $Y=3.33
+ $X2=2.01 $Y2=3.33
r52 15 17 93.6203 $w=1.68e-07 $l=1.435e-06 $layer=LI1_cond $X=1.675 $Y=3.33
+ $X2=0.24 $Y2=3.33
r53 13 32 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r54 13 18 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=0.24 $Y2=3.33
r55 13 29 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r56 9 12 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=3.12 $Y=1.985
+ $X2=3.12 $Y2=2.815
r57 7 35 3.13065 $w=2.5e-07 $l=1.09864e-07 $layer=LI1_cond $X=3.12 $Y=3.245
+ $X2=3.177 $Y2=3.33
r58 7 12 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=3.12 $Y=3.245 $X2=3.12
+ $Y2=2.815
r59 2 12 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=2.93
+ $Y=1.84 $X2=3.08 $Y2=2.815
r60 2 9 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=2.93
+ $Y=1.84 $X2=3.08 $Y2=1.985
r61 1 26 300 $w=1.7e-07 $l=1.15429e-06 $layer=licon1_PDIFF $count=2 $X=1.69
+ $Y=1.84 $X2=2.18 $Y2=2.775
.ends

.subckt PM_SKY130_FD_SC_HS__A32OI_1%VGND 1 2 7 9 11 13 15 17 30
r31 29 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r32 26 27 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r33 24 30 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r34 23 24 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r35 21 27 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r36 20 23 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=0.72 $Y=0 $X2=2.64
+ $Y2=0
r37 20 21 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r38 18 26 4.73185 $w=1.7e-07 $l=2.23e-07 $layer=LI1_cond $X=0.445 $Y=0 $X2=0.222
+ $Y2=0
r39 18 20 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=0.445 $Y=0 $X2=0.72
+ $Y2=0
r40 17 29 4.67962 $w=1.7e-07 $l=2.35e-07 $layer=LI1_cond $X=2.89 $Y=0 $X2=3.125
+ $Y2=0
r41 17 23 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=2.89 $Y=0 $X2=2.64
+ $Y2=0
r42 15 24 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.64
+ $Y2=0
r43 15 21 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=0.72
+ $Y2=0
r44 11 29 3.08656 $w=3.3e-07 $l=1.14782e-07 $layer=LI1_cond $X=3.055 $Y=0.085
+ $X2=3.125 $Y2=0
r45 11 13 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=3.055 $Y=0.085
+ $X2=3.055 $Y2=0.515
r46 7 26 3.03433 $w=3.3e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.28 $Y=0.085
+ $X2=0.222 $Y2=0
r47 7 9 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=0.28 $Y=0.085 $X2=0.28
+ $Y2=0.515
r48 2 13 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.915
+ $Y=0.37 $X2=3.055 $Y2=0.515
r49 1 9 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.515
.ends

