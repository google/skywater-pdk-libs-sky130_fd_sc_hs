* File: sky130_fd_sc_hs__sdfrbp_2.spice
* Created: Tue Sep  1 20:22:25 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hs__sdfrbp_2.pex.spice"
.subckt sky130_fd_sc_hs__sdfrbp_2  VNB VPB SCE D SCD RESET_B CLK VPWR Q_N Q VGND
* 
* VGND	VGND
* Q	Q
* Q_N	Q_N
* VPWR	VPWR
* CLK	CLK
* RESET_B	RESET_B
* SCD	SCD
* D	D
* SCE	SCE
* VPB	VPB
* VNB	VNB
MM1033 N_VGND_M1033_d N_SCE_M1033_g N_A_27_79#_M1033_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.1155 AS=0.1197 PD=1.39 PS=1.41 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1014 noxref_26 N_A_27_79#_M1014_g N_noxref_25_M1014_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.0504 AS=0.1197 PD=0.66 PS=1.41 NRD=18.564 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75002.3 A=0.063 P=1.14 MULT=1
MM1029 N_A_388_79#_M1029_d N_D_M1029_g noxref_26 VNB NLOWVT L=0.15 W=0.42
+ AD=0.13545 AS=0.0504 PD=1.065 PS=0.66 NRD=101.424 NRS=18.564 M=1 R=2.8
+ SA=75000.6 SB=75001.9 A=0.063 P=1.14 MULT=1
MM1034 noxref_27 N_SCE_M1034_g N_A_388_79#_M1029_d VNB NLOWVT L=0.15 W=0.42
+ AD=0.0504 AS=0.13545 PD=0.66 PS=1.065 NRD=18.564 NRS=2.856 M=1 R=2.8
+ SA=75001.4 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1015 N_noxref_25_M1015_d N_SCD_M1015_g noxref_27 VNB NLOWVT L=0.15 W=0.42
+ AD=0.0819 AS=0.0504 PD=0.81 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75001.8
+ SB=75000.7 A=0.063 P=1.14 MULT=1
MM1043 N_VGND_M1043_d N_RESET_B_M1043_g N_noxref_25_M1015_d VNB NLOWVT L=0.15
+ W=0.42 AD=0.1197 AS=0.0819 PD=1.41 PS=0.81 NRD=0 NRS=31.428 M=1 R=2.8
+ SA=75002.3 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1004 N_VGND_M1004_d N_CLK_M1004_g N_A_852_74#_M1004_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.2109 PD=1.02 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1006 N_A_1025_74#_M1006_d N_A_852_74#_M1006_g N_VGND_M1004_d VNB NLOWVT L=0.15
+ W=0.74 AD=0.2109 AS=0.1036 PD=2.05 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.6 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1019 N_A_1223_118#_M1019_d N_A_852_74#_M1019_g N_A_388_79#_M1019_s VNB NLOWVT
+ L=0.15 W=0.42 AD=0.0735 AS=0.1197 PD=0.77 PS=1.41 NRD=19.992 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75004.1 A=0.063 P=1.14 MULT=1
MM1020 A_1323_118# N_A_1025_74#_M1020_g N_A_1223_118#_M1019_d VNB NLOWVT L=0.15
+ W=0.42 AD=0.0504 AS=0.0735 PD=0.66 PS=0.77 NRD=18.564 NRS=0 M=1 R=2.8
+ SA=75000.7 SB=75003.6 A=0.063 P=1.14 MULT=1
MM1001 A_1401_118# N_A_1370_289#_M1001_g A_1323_118# VNB NLOWVT L=0.15 W=0.42
+ AD=0.0504 AS=0.0504 PD=0.66 PS=0.66 NRD=18.564 NRS=18.564 M=1 R=2.8 SA=75001.1
+ SB=75003.2 A=0.063 P=1.14 MULT=1
MM1012 N_VGND_M1012_d N_RESET_B_M1012_g A_1401_118# VNB NLOWVT L=0.15 W=0.42
+ AD=0.277973 AS=0.0504 PD=1.43038 PS=0.66 NRD=173.376 NRS=18.564 M=1 R=2.8
+ SA=75001.5 SB=75002.8 A=0.063 P=1.14 MULT=1
MM1003 N_A_1370_289#_M1003_d N_A_1223_118#_M1003_g N_VGND_M1012_d VNB NLOWVT
+ L=0.15 W=0.64 AD=0.0896 AS=0.423577 PD=0.92 PS=2.17962 NRD=0 NRS=113.772 M=1
+ R=4.26667 SA=75002 SB=75002.1 A=0.096 P=1.58 MULT=1
MM1024 N_A_1790_74#_M1024_d N_A_1025_74#_M1024_g N_A_1370_289#_M1003_d VNB
+ NLOWVT L=0.15 W=0.64 AD=0.261434 AS=0.0896 PD=1.85962 PS=0.92 NRD=105.936
+ NRS=0 M=1 R=4.26667 SA=75002.4 SB=75001.6 A=0.096 P=1.58 MULT=1
MM1002 A_2000_74# N_A_852_74#_M1002_g N_A_1790_74#_M1024_d VNB NLOWVT L=0.15
+ W=0.42 AD=0.0441 AS=0.171566 PD=0.63 PS=1.22038 NRD=14.28 NRS=15.708 M=1 R=2.8
+ SA=75003.2 SB=75001.3 A=0.063 P=1.14 MULT=1
MM1045 N_VGND_M1045_d N_A_2006_373#_M1045_g A_2000_74# VNB NLOWVT L=0.15 W=0.42
+ AD=0.0588 AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75003.5
+ SB=75001 A=0.063 P=1.14 MULT=1
MM1027 A_2158_74# N_RESET_B_M1027_g N_VGND_M1045_d VNB NLOWVT L=0.15 W=0.42
+ AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75003.9
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1018 N_A_2006_373#_M1018_d N_A_1790_74#_M1018_g A_2158_74# VNB NLOWVT L=0.15
+ W=0.42 AD=0.1113 AS=0.0441 PD=1.37 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8
+ SA=75004.3 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1028 N_Q_N_M1028_d N_A_1790_74#_M1028_g N_VGND_M1028_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.27675 PD=1.02 PS=2.42 NRD=0 NRS=10.536 M=1 R=4.93333
+ SA=75000.2 SB=75001 A=0.111 P=1.78 MULT=1
MM1039 N_Q_N_M1028_d N_A_1790_74#_M1039_g N_VGND_M1039_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.124942 PD=1.02 PS=1.14217 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.7 SB=75000.6 A=0.111 P=1.78 MULT=1
MM1010 N_A_2604_392#_M1010_d N_A_1790_74#_M1010_g N_VGND_M1039_s VNB NLOWVT
+ L=0.15 W=0.64 AD=0.1696 AS=0.108058 PD=1.81 PS=0.987826 NRD=0 NRS=8.436 M=1
+ R=4.26667 SA=75001.2 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1025 N_Q_M1025_d N_A_2604_392#_M1025_g N_VGND_M1025_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.2183 PD=1.02 PS=2.07 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1040 N_Q_M1025_d N_A_2604_392#_M1040_g N_VGND_M1040_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1998 PD=1.02 PS=2.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.6
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1023 N_VPWR_M1023_d N_SCE_M1023_g N_A_27_79#_M1023_s VPB PSHORT L=0.15 W=0.64
+ AD=0.2576 AS=0.1888 PD=1.445 PS=1.87 NRD=18.4589 NRS=3.0732 M=1 R=4.26667
+ SA=75000.2 SB=75003.3 A=0.096 P=1.58 MULT=1
MM1007 A_307_464# N_SCE_M1007_g N_VPWR_M1023_d VPB PSHORT L=0.15 W=0.64
+ AD=0.0864 AS=0.2576 PD=0.91 PS=1.445 NRD=24.625 NRS=3.0732 M=1 R=4.26667
+ SA=75001.2 SB=75002.4 A=0.096 P=1.58 MULT=1
MM1035 N_A_388_79#_M1035_d N_D_M1035_g A_307_464# VPB PSHORT L=0.15 W=0.64
+ AD=0.1872 AS=0.0864 PD=1.225 PS=0.91 NRD=46.1571 NRS=24.625 M=1 R=4.26667
+ SA=75001.6 SB=75001.9 A=0.096 P=1.58 MULT=1
MM1026 A_538_464# N_A_27_79#_M1026_g N_A_388_79#_M1035_d VPB PSHORT L=0.15
+ W=0.64 AD=0.0864 AS=0.1872 PD=0.91 PS=1.225 NRD=24.625 NRS=47.6937 M=1
+ R=4.26667 SA=75002.3 SB=75001.2 A=0.096 P=1.58 MULT=1
MM1005 N_VPWR_M1005_d N_SCD_M1005_g A_538_464# VPB PSHORT L=0.15 W=0.64
+ AD=0.1344 AS=0.0864 PD=1.06 PS=0.91 NRD=9.2196 NRS=24.625 M=1 R=4.26667
+ SA=75002.8 SB=75000.8 A=0.096 P=1.58 MULT=1
MM1044 N_A_388_79#_M1044_d N_RESET_B_M1044_g N_VPWR_M1005_d VPB PSHORT L=0.15
+ W=0.64 AD=0.1888 AS=0.1344 PD=1.87 PS=1.06 NRD=3.0732 NRS=33.8446 M=1
+ R=4.26667 SA=75003.3 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1022 N_VPWR_M1022_d N_CLK_M1022_g N_A_852_74#_M1022_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.3304 PD=1.42 PS=2.83 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75000.6 A=0.168 P=2.54 MULT=1
MM1032 N_A_1025_74#_M1032_d N_A_852_74#_M1032_g N_VPWR_M1022_d VPB PSHORT L=0.15
+ W=1.12 AD=0.308 AS=0.168 PD=2.79 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.7 SB=75000.2 A=0.168 P=2.54 MULT=1
MM1000 N_A_1223_118#_M1000_d N_A_1025_74#_M1000_g N_A_388_79#_M1000_s VPB PSHORT
+ L=0.15 W=0.42 AD=0.063 AS=0.1176 PD=0.72 PS=1.4 NRD=4.6886 NRS=4.6886 M=1
+ R=2.8 SA=75000.2 SB=75001.6 A=0.063 P=1.14 MULT=1
MM1008 A_1325_457# N_A_852_74#_M1008_g N_A_1223_118#_M1000_d VPB PSHORT L=0.15
+ W=0.42 AD=0.0504 AS=0.063 PD=0.66 PS=0.72 NRD=30.4759 NRS=4.6886 M=1 R=2.8
+ SA=75000.7 SB=75001.2 A=0.063 P=1.14 MULT=1
MM1037 N_VPWR_M1037_d N_A_1370_289#_M1037_g A_1325_457# VPB PSHORT L=0.15 W=0.42
+ AD=0.127687 AS=0.0504 PD=1.14 PS=0.66 NRD=116.782 NRS=30.4759 M=1 R=2.8
+ SA=75001 SB=75000.8 A=0.063 P=1.14 MULT=1
MM1013 N_A_1223_118#_M1013_d N_RESET_B_M1013_g N_VPWR_M1037_d VPB PSHORT L=0.15
+ W=0.42 AD=0.1176 AS=0.127687 PD=1.4 PS=1.14 NRD=4.6886 NRS=116.782 M=1 R=2.8
+ SA=75001.6 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1011 N_A_1370_289#_M1011_d N_A_1223_118#_M1011_g N_VPWR_M1011_s VPB PSHORT
+ L=0.15 W=1 AD=0.15 AS=0.275 PD=1.3 PS=2.55 NRD=1.9503 NRS=1.9503 M=1 R=6.66667
+ SA=75000.2 SB=75002.2 A=0.15 P=2.3 MULT=1
MM1016 N_A_1790_74#_M1016_d N_A_852_74#_M1016_g N_A_1370_289#_M1011_d VPB PSHORT
+ L=0.15 W=1 AD=0.283732 AS=0.15 PD=2.30986 PS=1.3 NRD=40.3653 NRS=1.9503 M=1
+ R=6.66667 SA=75000.6 SB=75001.7 A=0.15 P=2.3 MULT=1
MM1009 A_1955_471# N_A_1025_74#_M1009_g N_A_1790_74#_M1016_d VPB PSHORT L=0.15
+ W=0.42 AD=0.0567 AS=0.119168 PD=0.69 PS=0.970141 NRD=37.5088 NRS=53.9386 M=1
+ R=2.8 SA=75001.3 SB=75003.4 A=0.063 P=1.14 MULT=1
MM1038 N_VPWR_M1038_d N_A_2006_373#_M1038_g A_1955_471# VPB PSHORT L=0.15 W=0.42
+ AD=0.208462 AS=0.0567 PD=1.35 PS=0.69 NRD=107.877 NRS=37.5088 M=1 R=2.8
+ SA=75001.7 SB=75003 A=0.063 P=1.14 MULT=1
MM1036 N_A_2006_373#_M1036_d N_RESET_B_M1036_g N_VPWR_M1038_d VPB PSHORT L=0.15
+ W=0.42 AD=0.063 AS=0.208462 PD=0.72 PS=1.35 NRD=0 NRS=207.008 M=1 R=2.8
+ SA=75002.6 SB=75002.1 A=0.063 P=1.14 MULT=1
MM1041 N_VPWR_M1041_d N_A_1790_74#_M1041_g N_A_2006_373#_M1036_d VPB PSHORT
+ L=0.15 W=0.42 AD=0.0966 AS=0.063 PD=0.820909 PS=0.72 NRD=119.599 NRS=0 M=1
+ R=2.8 SA=75003 SB=75001.7 A=0.063 P=1.14 MULT=1
MM1017 N_Q_N_M1017_d N_A_1790_74#_M1017_g N_VPWR_M1041_d VPB PSHORT L=0.15
+ W=1.12 AD=0.168 AS=0.2576 PD=1.42 PS=2.18909 NRD=1.7533 NRS=1.7533 M=1
+ R=7.46667 SA=75001.5 SB=75001.1 A=0.168 P=2.54 MULT=1
MM1021 N_Q_N_M1017_d N_A_1790_74#_M1021_g N_VPWR_M1021_s VPB PSHORT L=0.15
+ W=1.12 AD=0.168 AS=0.204347 PD=1.42 PS=1.55849 NRD=1.7533 NRS=1.7533 M=1
+ R=7.46667 SA=75001.9 SB=75000.6 A=0.168 P=2.54 MULT=1
MM1042 N_A_2604_392#_M1042_d N_A_1790_74#_M1042_g N_VPWR_M1021_s VPB PSHORT
+ L=0.15 W=1 AD=0.275 AS=0.182453 PD=2.55 PS=1.39151 NRD=1.9503 NRS=12.7853 M=1
+ R=6.66667 SA=75002.6 SB=75000.2 A=0.15 P=2.3 MULT=1
MM1030 N_Q_M1030_d N_A_2604_392#_M1030_g N_VPWR_M1030_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.3304 PD=1.42 PS=2.83 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1031 N_Q_M1030_d N_A_2604_392#_M1031_g N_VPWR_M1031_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.3192 PD=1.42 PS=2.81 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.7 SB=75000.2 A=0.168 P=2.54 MULT=1
DX46_noxref VNB VPB NWDIODE A=28.7406 P=34.45
c_152 VNB 0 7.64129e-20 $X=0 $Y=0
c_2039 A_1955_471# 0 1.03069e-19 $X=9.775 $Y=2.355
*
.include "sky130_fd_sc_hs__sdfrbp_2.pxi.spice"
*
.ends
*
*
