* File: sky130_fd_sc_hs__sdfrbp_2.pxi.spice
* Created: Thu Aug 27 21:08:27 2020
* 
x_PM_SKY130_FD_SC_HS__SDFRBP_2%A_27_79# N_A_27_79#_M1033_s N_A_27_79#_M1023_s
+ N_A_27_79#_M1014_g N_A_27_79#_c_289_n N_A_27_79#_M1026_g N_A_27_79#_c_284_n
+ N_A_27_79#_c_285_n N_A_27_79#_c_286_n N_A_27_79#_c_291_n N_A_27_79#_c_287_n
+ N_A_27_79#_c_303_p N_A_27_79#_c_292_n N_A_27_79#_c_288_n N_A_27_79#_c_293_n
+ PM_SKY130_FD_SC_HS__SDFRBP_2%A_27_79#
x_PM_SKY130_FD_SC_HS__SDFRBP_2%SCE N_SCE_c_366_n N_SCE_c_367_n N_SCE_M1033_g
+ N_SCE_c_375_n N_SCE_M1023_g N_SCE_c_376_n N_SCE_M1007_g N_SCE_M1034_g
+ N_SCE_c_369_n N_SCE_c_370_n N_SCE_c_371_n N_SCE_c_372_n N_SCE_c_373_n SCE SCE
+ SCE N_SCE_c_378_n N_SCE_c_379_n PM_SKY130_FD_SC_HS__SDFRBP_2%SCE
x_PM_SKY130_FD_SC_HS__SDFRBP_2%D N_D_M1029_g N_D_c_452_n N_D_c_457_n N_D_M1035_g
+ D N_D_c_453_n N_D_c_454_n N_D_c_455_n PM_SKY130_FD_SC_HS__SDFRBP_2%D
x_PM_SKY130_FD_SC_HS__SDFRBP_2%SCD N_SCD_c_503_n N_SCD_M1005_g N_SCD_M1015_g
+ N_SCD_c_500_n SCD SCD N_SCD_c_502_n PM_SKY130_FD_SC_HS__SDFRBP_2%SCD
x_PM_SKY130_FD_SC_HS__SDFRBP_2%RESET_B N_RESET_B_M1043_g N_RESET_B_c_551_n
+ N_RESET_B_M1044_g N_RESET_B_c_544_n N_RESET_B_M1012_g N_RESET_B_c_545_n
+ N_RESET_B_c_546_n N_RESET_B_c_552_n N_RESET_B_M1013_g N_RESET_B_c_547_n
+ N_RESET_B_M1027_g N_RESET_B_c_554_n N_RESET_B_c_555_n N_RESET_B_M1036_g
+ N_RESET_B_c_549_n N_RESET_B_c_557_n N_RESET_B_c_558_n N_RESET_B_c_559_n
+ N_RESET_B_c_560_n RESET_B N_RESET_B_c_562_n N_RESET_B_c_563_n
+ N_RESET_B_c_564_n N_RESET_B_c_565_n N_RESET_B_c_566_n
+ PM_SKY130_FD_SC_HS__SDFRBP_2%RESET_B
x_PM_SKY130_FD_SC_HS__SDFRBP_2%CLK N_CLK_c_733_n N_CLK_M1004_g N_CLK_c_734_n
+ N_CLK_M1022_g N_CLK_c_735_n CLK PM_SKY130_FD_SC_HS__SDFRBP_2%CLK
x_PM_SKY130_FD_SC_HS__SDFRBP_2%A_1025_74# N_A_1025_74#_M1006_d
+ N_A_1025_74#_M1032_d N_A_1025_74#_c_806_n N_A_1025_74#_c_807_n
+ N_A_1025_74#_M1000_g N_A_1025_74#_c_785_n N_A_1025_74#_M1020_g
+ N_A_1025_74#_c_787_n N_A_1025_74#_M1024_g N_A_1025_74#_c_788_n
+ N_A_1025_74#_c_789_n N_A_1025_74#_c_808_n N_A_1025_74#_M1009_g
+ N_A_1025_74#_c_790_n N_A_1025_74#_c_791_n N_A_1025_74#_c_792_n
+ N_A_1025_74#_c_793_n N_A_1025_74#_c_794_n N_A_1025_74#_c_795_n
+ N_A_1025_74#_c_796_n N_A_1025_74#_c_964_p N_A_1025_74#_c_797_n
+ N_A_1025_74#_c_798_n N_A_1025_74#_c_799_n N_A_1025_74#_c_800_n
+ N_A_1025_74#_c_801_n N_A_1025_74#_c_802_n N_A_1025_74#_c_803_n
+ N_A_1025_74#_c_811_n N_A_1025_74#_c_804_n N_A_1025_74#_c_805_n
+ PM_SKY130_FD_SC_HS__SDFRBP_2%A_1025_74#
x_PM_SKY130_FD_SC_HS__SDFRBP_2%A_1370_289# N_A_1370_289#_M1003_d
+ N_A_1370_289#_M1011_d N_A_1370_289#_c_995_n N_A_1370_289#_M1001_g
+ N_A_1370_289#_c_996_n N_A_1370_289#_M1037_g N_A_1370_289#_c_990_n
+ N_A_1370_289#_c_991_n N_A_1370_289#_c_1027_n N_A_1370_289#_c_1029_n
+ N_A_1370_289#_c_999_n N_A_1370_289#_c_992_n N_A_1370_289#_c_993_n
+ N_A_1370_289#_c_994_n PM_SKY130_FD_SC_HS__SDFRBP_2%A_1370_289#
x_PM_SKY130_FD_SC_HS__SDFRBP_2%A_1223_118# N_A_1223_118#_M1019_d
+ N_A_1223_118#_M1000_d N_A_1223_118#_M1013_d N_A_1223_118#_M1003_g
+ N_A_1223_118#_c_1087_n N_A_1223_118#_M1011_g N_A_1223_118#_c_1119_n
+ N_A_1223_118#_c_1088_n N_A_1223_118#_c_1101_n N_A_1223_118#_c_1094_n
+ N_A_1223_118#_c_1089_n N_A_1223_118#_c_1090_n N_A_1223_118#_c_1091_n
+ PM_SKY130_FD_SC_HS__SDFRBP_2%A_1223_118#
x_PM_SKY130_FD_SC_HS__SDFRBP_2%A_852_74# N_A_852_74#_M1004_s N_A_852_74#_M1022_s
+ N_A_852_74#_M1006_g N_A_852_74#_c_1191_n N_A_852_74#_M1032_g
+ N_A_852_74#_c_1192_n N_A_852_74#_c_1193_n N_A_852_74#_c_1194_n
+ N_A_852_74#_c_1208_n N_A_852_74#_c_1209_n N_A_852_74#_c_1195_n
+ N_A_852_74#_M1019_g N_A_852_74#_c_1210_n N_A_852_74#_c_1211_n
+ N_A_852_74#_c_1212_n N_A_852_74#_M1008_g N_A_852_74#_c_1213_n
+ N_A_852_74#_c_1214_n N_A_852_74#_c_1215_n N_A_852_74#_M1016_g
+ N_A_852_74#_c_1196_n N_A_852_74#_c_1197_n N_A_852_74#_M1002_g
+ N_A_852_74#_c_1199_n N_A_852_74#_c_1219_n N_A_852_74#_c_1200_n
+ N_A_852_74#_c_1201_n N_A_852_74#_c_1232_n N_A_852_74#_c_1220_n
+ N_A_852_74#_c_1202_n N_A_852_74#_c_1203_n N_A_852_74#_c_1222_n
+ N_A_852_74#_c_1204_n N_A_852_74#_c_1205_n
+ PM_SKY130_FD_SC_HS__SDFRBP_2%A_852_74#
x_PM_SKY130_FD_SC_HS__SDFRBP_2%A_2006_373# N_A_2006_373#_M1018_d
+ N_A_2006_373#_M1036_d N_A_2006_373#_c_1391_n N_A_2006_373#_M1038_g
+ N_A_2006_373#_M1045_g N_A_2006_373#_c_1393_n N_A_2006_373#_c_1385_n
+ N_A_2006_373#_c_1386_n N_A_2006_373#_c_1395_n N_A_2006_373#_c_1396_n
+ N_A_2006_373#_c_1387_n N_A_2006_373#_c_1388_n N_A_2006_373#_c_1389_n
+ N_A_2006_373#_c_1390_n N_A_2006_373#_c_1397_n N_A_2006_373#_c_1398_n
+ PM_SKY130_FD_SC_HS__SDFRBP_2%A_2006_373#
x_PM_SKY130_FD_SC_HS__SDFRBP_2%A_1790_74# N_A_1790_74#_M1024_d
+ N_A_1790_74#_M1016_d N_A_1790_74#_M1018_g N_A_1790_74#_c_1495_n
+ N_A_1790_74#_c_1505_n N_A_1790_74#_c_1506_n N_A_1790_74#_M1041_g
+ N_A_1790_74#_c_1496_n N_A_1790_74#_c_1507_n N_A_1790_74#_M1017_g
+ N_A_1790_74#_M1028_g N_A_1790_74#_c_1508_n N_A_1790_74#_M1021_g
+ N_A_1790_74#_M1039_g N_A_1790_74#_c_1499_n N_A_1790_74#_c_1500_n
+ N_A_1790_74#_c_1511_n N_A_1790_74#_M1042_g N_A_1790_74#_M1010_g
+ N_A_1790_74#_c_1522_n N_A_1790_74#_c_1531_n N_A_1790_74#_c_1502_n
+ N_A_1790_74#_c_1503_n N_A_1790_74#_c_1504_n N_A_1790_74#_c_1541_n
+ PM_SKY130_FD_SC_HS__SDFRBP_2%A_1790_74#
x_PM_SKY130_FD_SC_HS__SDFRBP_2%A_2604_392# N_A_2604_392#_M1010_d
+ N_A_2604_392#_M1042_d N_A_2604_392#_c_1652_n N_A_2604_392#_M1030_g
+ N_A_2604_392#_M1025_g N_A_2604_392#_c_1653_n N_A_2604_392#_M1031_g
+ N_A_2604_392#_M1040_g N_A_2604_392#_c_1647_n N_A_2604_392#_c_1648_n
+ N_A_2604_392#_c_1649_n N_A_2604_392#_c_1650_n N_A_2604_392#_c_1669_p
+ N_A_2604_392#_c_1651_n PM_SKY130_FD_SC_HS__SDFRBP_2%A_2604_392#
x_PM_SKY130_FD_SC_HS__SDFRBP_2%VPWR N_VPWR_M1023_d N_VPWR_M1005_d N_VPWR_M1022_d
+ N_VPWR_M1037_d N_VPWR_M1011_s N_VPWR_M1038_d N_VPWR_M1041_d N_VPWR_M1021_s
+ N_VPWR_M1030_s N_VPWR_M1031_s N_VPWR_c_1697_n N_VPWR_c_1698_n N_VPWR_c_1699_n
+ N_VPWR_c_1700_n N_VPWR_c_1701_n N_VPWR_c_1702_n N_VPWR_c_1703_n
+ N_VPWR_c_1704_n N_VPWR_c_1705_n N_VPWR_c_1706_n N_VPWR_c_1707_n
+ N_VPWR_c_1708_n N_VPWR_c_1709_n N_VPWR_c_1710_n VPWR N_VPWR_c_1711_n
+ N_VPWR_c_1712_n N_VPWR_c_1713_n N_VPWR_c_1714_n N_VPWR_c_1715_n
+ N_VPWR_c_1716_n N_VPWR_c_1717_n N_VPWR_c_1718_n N_VPWR_c_1719_n
+ N_VPWR_c_1720_n N_VPWR_c_1721_n N_VPWR_c_1722_n N_VPWR_c_1723_n
+ N_VPWR_c_1724_n N_VPWR_c_1696_n PM_SKY130_FD_SC_HS__SDFRBP_2%VPWR
x_PM_SKY130_FD_SC_HS__SDFRBP_2%A_388_79# N_A_388_79#_M1029_d N_A_388_79#_M1019_s
+ N_A_388_79#_M1035_d N_A_388_79#_M1044_d N_A_388_79#_M1000_s
+ N_A_388_79#_c_1898_n N_A_388_79#_c_1879_n N_A_388_79#_c_1880_n
+ N_A_388_79#_c_1881_n N_A_388_79#_c_1900_n N_A_388_79#_c_1921_n
+ N_A_388_79#_c_1888_n N_A_388_79#_c_1882_n N_A_388_79#_c_1890_n
+ N_A_388_79#_c_1891_n N_A_388_79#_c_1892_n N_A_388_79#_c_1883_n
+ N_A_388_79#_c_1893_n N_A_388_79#_c_1894_n N_A_388_79#_c_1884_n
+ N_A_388_79#_c_1885_n N_A_388_79#_c_1886_n N_A_388_79#_c_1887_n
+ N_A_388_79#_c_1896_n PM_SKY130_FD_SC_HS__SDFRBP_2%A_388_79#
x_PM_SKY130_FD_SC_HS__SDFRBP_2%Q_N N_Q_N_M1028_d N_Q_N_M1017_d Q_N Q_N Q_N
+ N_Q_N_c_2041_n Q_N PM_SKY130_FD_SC_HS__SDFRBP_2%Q_N
x_PM_SKY130_FD_SC_HS__SDFRBP_2%Q N_Q_M1025_d N_Q_M1030_d Q N_Q_c_2068_n
+ PM_SKY130_FD_SC_HS__SDFRBP_2%Q
x_PM_SKY130_FD_SC_HS__SDFRBP_2%VGND N_VGND_M1033_d N_VGND_M1043_d N_VGND_M1004_d
+ N_VGND_M1012_d N_VGND_M1045_d N_VGND_M1028_s N_VGND_M1039_s N_VGND_M1025_s
+ N_VGND_M1040_s N_VGND_c_2084_n N_VGND_c_2085_n N_VGND_c_2086_n N_VGND_c_2087_n
+ N_VGND_c_2088_n N_VGND_c_2089_n N_VGND_c_2090_n N_VGND_c_2091_n
+ N_VGND_c_2092_n N_VGND_c_2093_n N_VGND_c_2094_n N_VGND_c_2095_n
+ N_VGND_c_2096_n N_VGND_c_2097_n N_VGND_c_2098_n N_VGND_c_2099_n VGND
+ N_VGND_c_2100_n N_VGND_c_2101_n N_VGND_c_2102_n N_VGND_c_2103_n
+ N_VGND_c_2104_n N_VGND_c_2105_n N_VGND_c_2106_n N_VGND_c_2107_n
+ N_VGND_c_2108_n N_VGND_c_2109_n N_VGND_c_2110_n
+ PM_SKY130_FD_SC_HS__SDFRBP_2%VGND
x_PM_SKY130_FD_SC_HS__SDFRBP_2%noxref_25 N_noxref_25_M1014_s N_noxref_25_M1015_d
+ N_noxref_25_c_2241_n N_noxref_25_c_2242_n N_noxref_25_c_2243_n
+ N_noxref_25_c_2244_n PM_SKY130_FD_SC_HS__SDFRBP_2%noxref_25
cc_1 VNB N_A_27_79#_M1014_g 0.0455097f $X=-0.19 $Y=-0.245 $X2=1.475 $Y2=0.605
cc_2 VNB N_A_27_79#_c_284_n 0.0789787f $X=-0.19 $Y=-0.245 $X2=1.4 $Y2=1.415
cc_3 VNB N_A_27_79#_c_285_n 0.0355558f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=0.605
cc_4 VNB N_A_27_79#_c_286_n 0.00354448f $X=-0.19 $Y=-0.245 $X2=0.2 $Y2=2.32
cc_5 VNB N_A_27_79#_c_287_n 0.00484068f $X=-0.19 $Y=-0.245 $X2=1.23 $Y2=1.415
cc_6 VNB N_A_27_79#_c_288_n 0.0159647f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.415
cc_7 VNB N_SCE_c_366_n 0.0443833f $X=-0.19 $Y=-0.245 $X2=0.135 $Y2=2.32
cc_8 VNB N_SCE_c_367_n 0.0211781f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_SCE_M1034_g 0.0363026f $X=-0.19 $Y=-0.245 $X2=1.4 $Y2=1.415
cc_10 VNB N_SCE_c_369_n 0.0216296f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_SCE_c_370_n 0.00133979f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=2.65
cc_12 VNB N_SCE_c_371_n 0.00450757f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_SCE_c_372_n 0.0230028f $X=-0.19 $Y=-0.245 $X2=1.23 $Y2=1.415
cc_14 VNB N_SCE_c_373_n 0.0330707f $X=-0.19 $Y=-0.245 $X2=1.23 $Y2=1.415
cc_15 VNB N_D_c_452_n 0.0238331f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_D_c_453_n 0.0310845f $X=-0.19 $Y=-0.245 $X2=2.615 $Y2=2.64
cc_17 VNB N_D_c_454_n 0.00902418f $X=-0.19 $Y=-0.245 $X2=2.615 $Y2=2.64
cc_18 VNB N_D_c_455_n 0.0162587f $X=-0.19 $Y=-0.245 $X2=1.4 $Y2=1.415
cc_19 VNB N_SCD_M1015_g 0.043102f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_SCD_c_500_n 0.0051095f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB SCD 0.00197778f $X=-0.19 $Y=-0.245 $X2=2.615 $Y2=2.245
cc_22 VNB N_SCD_c_502_n 0.0165348f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=0.605
cc_23 VNB N_RESET_B_M1043_g 0.0661566f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_RESET_B_c_544_n 0.0188088f $X=-0.19 $Y=-0.245 $X2=1.475 $Y2=0.605
cc_25 VNB N_RESET_B_c_545_n 0.0282366f $X=-0.19 $Y=-0.245 $X2=2.615 $Y2=2.245
cc_26 VNB N_RESET_B_c_546_n 0.0118779f $X=-0.19 $Y=-0.245 $X2=2.615 $Y2=2.64
cc_27 VNB N_RESET_B_c_547_n 0.0227742f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=0.605
cc_28 VNB N_RESET_B_M1027_g 0.0456332f $X=-0.19 $Y=-0.245 $X2=0.2 $Y2=2.32
cc_29 VNB N_RESET_B_c_549_n 0.0112292f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_CLK_c_733_n 0.0203282f $X=-0.19 $Y=-0.245 $X2=0.135 $Y2=0.395
cc_31 VNB N_CLK_c_734_n 0.0232936f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_CLK_c_735_n 0.0614545f $X=-0.19 $Y=-0.245 $X2=1.475 $Y2=0.605
cc_33 VNB CLK 0.0142868f $X=-0.19 $Y=-0.245 $X2=1.475 $Y2=0.605
cc_34 VNB N_A_1025_74#_c_785_n 0.0266196f $X=-0.19 $Y=-0.245 $X2=2.615 $Y2=2.64
cc_35 VNB N_A_1025_74#_M1020_g 0.038919f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=0.605
cc_36 VNB N_A_1025_74#_c_787_n 0.016501f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_1025_74#_c_788_n 0.0226212f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=2.49
cc_38 VNB N_A_1025_74#_c_789_n 0.00721388f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=2.65
cc_39 VNB N_A_1025_74#_c_790_n 0.00587392f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_1025_74#_c_791_n 0.0261185f $X=-0.19 $Y=-0.245 $X2=2.275 $Y2=2.405
cc_41 VNB N_A_1025_74#_c_792_n 0.00279409f $X=-0.19 $Y=-0.245 $X2=0.445
+ $Y2=2.405
cc_42 VNB N_A_1025_74#_c_793_n 0.00205192f $X=-0.19 $Y=-0.245 $X2=2.44 $Y2=1.995
cc_43 VNB N_A_1025_74#_c_794_n 9.68255e-19 $X=-0.19 $Y=-0.245 $X2=2.44 $Y2=1.995
cc_44 VNB N_A_1025_74#_c_795_n 0.00204982f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_A_1025_74#_c_796_n 0.00173368f $X=-0.19 $Y=-0.245 $X2=1.23 $Y2=1.415
cc_46 VNB N_A_1025_74#_c_797_n 0.00706005f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_1025_74#_c_798_n 0.00245748f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_1025_74#_c_799_n 0.00157163f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A_1025_74#_c_800_n 0.00699014f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_A_1025_74#_c_801_n 0.00573141f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_A_1025_74#_c_802_n 0.00460249f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_A_1025_74#_c_803_n 0.033082f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_A_1025_74#_c_804_n 0.0048475f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_A_1025_74#_c_805_n 0.0142363f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_A_1370_289#_M1001_g 0.0322358f $X=-0.19 $Y=-0.245 $X2=2.615
+ $Y2=2.245
cc_56 VNB N_A_1370_289#_c_990_n 0.00365613f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_A_1370_289#_c_991_n 0.0259328f $X=-0.19 $Y=-0.245 $X2=0.2 $Y2=1.58
cc_58 VNB N_A_1370_289#_c_992_n 0.00572372f $X=-0.19 $Y=-0.245 $X2=2.44
+ $Y2=1.995
cc_59 VNB N_A_1370_289#_c_993_n 0.00431592f $X=-0.19 $Y=-0.245 $X2=2.44
+ $Y2=1.995
cc_60 VNB N_A_1370_289#_c_994_n 0.00664491f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_A_1223_118#_M1003_g 0.026757f $X=-0.19 $Y=-0.245 $X2=2.615 $Y2=2.64
cc_62 VNB N_A_1223_118#_c_1087_n 0.0288104f $X=-0.19 $Y=-0.245 $X2=1.4 $Y2=1.415
cc_63 VNB N_A_1223_118#_c_1088_n 0.010971f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=2.65
cc_64 VNB N_A_1223_118#_c_1089_n 0.00155425f $X=-0.19 $Y=-0.245 $X2=1.23
+ $Y2=1.415
cc_65 VNB N_A_1223_118#_c_1090_n 0.00407991f $X=-0.19 $Y=-0.245 $X2=1.23
+ $Y2=1.415
cc_66 VNB N_A_1223_118#_c_1091_n 0.00984617f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_A_852_74#_M1006_g 0.0262718f $X=-0.19 $Y=-0.245 $X2=1.475 $Y2=0.605
cc_68 VNB N_A_852_74#_c_1191_n 0.0193778f $X=-0.19 $Y=-0.245 $X2=2.615 $Y2=2.245
cc_69 VNB N_A_852_74#_c_1192_n 0.00997766f $X=-0.19 $Y=-0.245 $X2=1.4 $Y2=1.415
cc_70 VNB N_A_852_74#_c_1193_n 0.00688658f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=0.605
cc_71 VNB N_A_852_74#_c_1194_n 0.0251276f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_A_852_74#_c_1195_n 0.0193173f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=2.65
cc_73 VNB N_A_852_74#_c_1196_n 0.029955f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=2.405
cc_74 VNB N_A_852_74#_c_1197_n 0.00539027f $X=-0.19 $Y=-0.245 $X2=1.23 $Y2=1.415
cc_75 VNB N_A_852_74#_M1002_g 0.0453681f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_A_852_74#_c_1199_n 0.0215149f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_A_852_74#_c_1200_n 0.00740257f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_A_852_74#_c_1201_n 0.00277221f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VNB N_A_852_74#_c_1202_n 4.53969e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_A_852_74#_c_1203_n 0.00281383f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_81 VNB N_A_852_74#_c_1204_n 0.00183723f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_82 VNB N_A_852_74#_c_1205_n 0.00622133f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_83 VNB N_A_2006_373#_M1045_g 0.0481405f $X=-0.19 $Y=-0.245 $X2=2.615 $Y2=2.64
cc_84 VNB N_A_2006_373#_c_1385_n 0.00410394f $X=-0.19 $Y=-0.245 $X2=0.2 $Y2=1.58
cc_85 VNB N_A_2006_373#_c_1386_n 0.00173724f $X=-0.19 $Y=-0.245 $X2=0.2 $Y2=2.32
cc_86 VNB N_A_2006_373#_c_1387_n 0.0070639f $X=-0.19 $Y=-0.245 $X2=0.365
+ $Y2=1.415
cc_87 VNB N_A_2006_373#_c_1388_n 0.00667447f $X=-0.19 $Y=-0.245 $X2=1.23
+ $Y2=1.415
cc_88 VNB N_A_2006_373#_c_1389_n 0.00230863f $X=-0.19 $Y=-0.245 $X2=1.23
+ $Y2=1.415
cc_89 VNB N_A_2006_373#_c_1390_n 0.00172407f $X=-0.19 $Y=-0.245 $X2=2.275
+ $Y2=2.405
cc_90 VNB N_A_1790_74#_M1018_g 0.0262898f $X=-0.19 $Y=-0.245 $X2=1.475 $Y2=0.605
cc_91 VNB N_A_1790_74#_c_1495_n 0.0559917f $X=-0.19 $Y=-0.245 $X2=2.615
+ $Y2=2.245
cc_92 VNB N_A_1790_74#_c_1496_n 0.0318785f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=0.605
cc_93 VNB N_A_1790_74#_M1028_g 0.0197591f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=2.65
cc_94 VNB N_A_1790_74#_M1039_g 0.0192815f $X=-0.19 $Y=-0.245 $X2=2.275 $Y2=2.405
cc_95 VNB N_A_1790_74#_c_1499_n 0.0729414f $X=-0.19 $Y=-0.245 $X2=2.44 $Y2=2.32
cc_96 VNB N_A_1790_74#_c_1500_n 0.00428291f $X=-0.19 $Y=-0.245 $X2=2.44
+ $Y2=1.995
cc_97 VNB N_A_1790_74#_M1010_g 0.027051f $X=-0.19 $Y=-0.245 $X2=1.23 $Y2=1.415
cc_98 VNB N_A_1790_74#_c_1502_n 0.00230536f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_99 VNB N_A_1790_74#_c_1503_n 0.00223918f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_100 VNB N_A_1790_74#_c_1504_n 0.021329f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_101 VNB N_A_2604_392#_M1025_g 0.023917f $X=-0.19 $Y=-0.245 $X2=2.615 $Y2=2.64
cc_102 VNB N_A_2604_392#_M1040_g 0.0268211f $X=-0.19 $Y=-0.245 $X2=0.2 $Y2=1.58
cc_103 VNB N_A_2604_392#_c_1647_n 0.0652038f $X=-0.19 $Y=-0.245 $X2=0.28
+ $Y2=2.49
cc_104 VNB N_A_2604_392#_c_1648_n 0.0587782f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_105 VNB N_A_2604_392#_c_1649_n 0.0102396f $X=-0.19 $Y=-0.245 $X2=1.23
+ $Y2=1.415
cc_106 VNB N_A_2604_392#_c_1650_n 7.2775e-19 $X=-0.19 $Y=-0.245 $X2=2.44
+ $Y2=2.32
cc_107 VNB N_A_2604_392#_c_1651_n 0.00109231f $X=-0.19 $Y=-0.245 $X2=2.49
+ $Y2=1.995
cc_108 VNB N_VPWR_c_1696_n 0.621437f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_109 VNB N_A_388_79#_c_1879_n 0.00214649f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=2.65
cc_110 VNB N_A_388_79#_c_1880_n 0.0244723f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_111 VNB N_A_388_79#_c_1881_n 0.00417762f $X=-0.19 $Y=-0.245 $X2=0.365
+ $Y2=1.415
cc_112 VNB N_A_388_79#_c_1882_n 0.0041886f $X=-0.19 $Y=-0.245 $X2=0.445
+ $Y2=2.405
cc_113 VNB N_A_388_79#_c_1883_n 7.83649e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_114 VNB N_A_388_79#_c_1884_n 0.00627051f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_115 VNB N_A_388_79#_c_1885_n 0.00155859f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_116 VNB N_A_388_79#_c_1886_n 0.00308378f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_117 VNB N_A_388_79#_c_1887_n 0.00186702f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_118 VNB Q_N 0.00143966f $X=-0.19 $Y=-0.245 $X2=1.475 $Y2=0.605
cc_119 VNB N_Q_N_c_2041_n 0.00240191f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=0.605
cc_120 VNB N_Q_c_2068_n 0.0065793f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_121 VNB N_VGND_c_2084_n 0.0153683f $X=-0.19 $Y=-0.245 $X2=2.275 $Y2=2.405
cc_122 VNB N_VGND_c_2085_n 0.0225707f $X=-0.19 $Y=-0.245 $X2=2.44 $Y2=1.995
cc_123 VNB N_VGND_c_2086_n 0.00983072f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=2.405
cc_124 VNB N_VGND_c_2087_n 0.00692506f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_125 VNB N_VGND_c_2088_n 0.00869988f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_126 VNB N_VGND_c_2089_n 0.0114612f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_127 VNB N_VGND_c_2090_n 0.0225701f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_128 VNB N_VGND_c_2091_n 0.00935384f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_129 VNB N_VGND_c_2092_n 0.0108727f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_130 VNB N_VGND_c_2093_n 0.0526431f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_131 VNB N_VGND_c_2094_n 0.0659895f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_132 VNB N_VGND_c_2095_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_133 VNB N_VGND_c_2096_n 0.0221562f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_134 VNB N_VGND_c_2097_n 0.00326991f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_135 VNB N_VGND_c_2098_n 0.0583825f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_136 VNB N_VGND_c_2099_n 0.00604233f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_137 VNB N_VGND_c_2100_n 0.0176416f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_138 VNB N_VGND_c_2101_n 0.0276584f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_139 VNB N_VGND_c_2102_n 0.0209223f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_140 VNB N_VGND_c_2103_n 0.0186734f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_141 VNB N_VGND_c_2104_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_142 VNB N_VGND_c_2105_n 0.0615922f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_143 VNB N_VGND_c_2106_n 0.0213232f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_144 VNB N_VGND_c_2107_n 0.00478044f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_145 VNB N_VGND_c_2108_n 0.00500104f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_146 VNB N_VGND_c_2109_n 0.00326991f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_147 VNB N_VGND_c_2110_n 0.813571f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_148 VNB N_noxref_25_c_2241_n 0.00622698f $X=-0.19 $Y=-0.245 $X2=1.475
+ $Y2=0.605
cc_149 VNB N_noxref_25_c_2242_n 0.0179038f $X=-0.19 $Y=-0.245 $X2=2.615
+ $Y2=2.245
cc_150 VNB N_noxref_25_c_2243_n 0.00386383f $X=-0.19 $Y=-0.245 $X2=2.615
+ $Y2=2.64
cc_151 VNB N_noxref_25_c_2244_n 0.00277566f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.25
cc_152 VPB N_A_27_79#_c_289_n 0.0656313f $X=-0.19 $Y=1.66 $X2=2.615 $Y2=2.245
cc_153 VPB N_A_27_79#_c_286_n 0.031275f $X=-0.19 $Y=1.66 $X2=0.2 $Y2=2.32
cc_154 VPB N_A_27_79#_c_291_n 0.0213374f $X=-0.19 $Y=1.66 $X2=0.28 $Y2=2.65
cc_155 VPB N_A_27_79#_c_292_n 0.00449549f $X=-0.19 $Y=1.66 $X2=2.44 $Y2=1.995
cc_156 VPB N_A_27_79#_c_293_n 0.00957909f $X=-0.19 $Y=1.66 $X2=0.28 $Y2=2.405
cc_157 VPB N_SCE_c_366_n 0.013397f $X=-0.19 $Y=1.66 $X2=0.135 $Y2=2.32
cc_158 VPB N_SCE_c_375_n 0.052364f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_159 VPB N_SCE_c_376_n 0.0413346f $X=-0.19 $Y=1.66 $X2=1.475 $Y2=0.605
cc_160 VPB N_SCE_c_370_n 0.00700226f $X=-0.19 $Y=1.66 $X2=0.28 $Y2=2.65
cc_161 VPB N_SCE_c_378_n 0.0605067f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_162 VPB N_SCE_c_379_n 0.00222208f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_163 VPB N_D_c_452_n 0.0324711f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_164 VPB N_D_c_457_n 0.0243702f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_165 VPB N_SCD_c_503_n 0.0168486f $X=-0.19 $Y=1.66 $X2=0.135 $Y2=0.395
cc_166 VPB N_SCD_c_500_n 0.0502021f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_167 VPB SCD 0.00164561f $X=-0.19 $Y=1.66 $X2=2.615 $Y2=2.245
cc_168 VPB N_RESET_B_M1043_g 0.0118663f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_169 VPB N_RESET_B_c_551_n 0.0217569f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_170 VPB N_RESET_B_c_552_n 0.0164974f $X=-0.19 $Y=1.66 $X2=2.615 $Y2=2.64
cc_171 VPB N_RESET_B_c_547_n 0.009182f $X=-0.19 $Y=1.66 $X2=0.28 $Y2=0.605
cc_172 VPB N_RESET_B_c_554_n 0.0120728f $X=-0.19 $Y=1.66 $X2=0.28 $Y2=2.65
cc_173 VPB N_RESET_B_c_555_n 0.0547375f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_174 VPB N_RESET_B_c_549_n 0.00587573f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_175 VPB N_RESET_B_c_557_n 0.0217181f $X=-0.19 $Y=1.66 $X2=0.445 $Y2=2.405
cc_176 VPB N_RESET_B_c_558_n 0.00332059f $X=-0.19 $Y=1.66 $X2=2.44 $Y2=2.32
cc_177 VPB N_RESET_B_c_559_n 0.00850003f $X=-0.19 $Y=1.66 $X2=2.44 $Y2=1.995
cc_178 VPB N_RESET_B_c_560_n 0.00382672f $X=-0.19 $Y=1.66 $X2=2.44 $Y2=1.995
cc_179 VPB RESET_B 0.00298374f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_180 VPB N_RESET_B_c_562_n 0.0678306f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_181 VPB N_RESET_B_c_563_n 0.00203407f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_182 VPB N_RESET_B_c_564_n 0.0565102f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_183 VPB N_RESET_B_c_565_n 0.00232432f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_184 VPB N_RESET_B_c_566_n 0.0062794f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_185 VPB N_CLK_c_734_n 0.0296847f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_186 VPB N_A_1025_74#_c_806_n 0.0182724f $X=-0.19 $Y=1.66 $X2=1.475 $Y2=0.605
cc_187 VPB N_A_1025_74#_c_807_n 0.0206464f $X=-0.19 $Y=1.66 $X2=1.475 $Y2=0.605
cc_188 VPB N_A_1025_74#_c_808_n 0.0554159f $X=-0.19 $Y=1.66 $X2=0.28 $Y2=2.65
cc_189 VPB N_A_1025_74#_c_794_n 0.00487395f $X=-0.19 $Y=1.66 $X2=2.44 $Y2=1.995
cc_190 VPB N_A_1025_74#_c_795_n 0.00205711f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_191 VPB N_A_1025_74#_c_811_n 0.00662341f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_192 VPB N_A_1025_74#_c_804_n 0.0041865f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_193 VPB N_A_1025_74#_c_805_n 0.0162545f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_194 VPB N_A_1370_289#_c_995_n 0.0248418f $X=-0.19 $Y=1.66 $X2=1.475 $Y2=0.605
cc_195 VPB N_A_1370_289#_c_996_n 0.0209394f $X=-0.19 $Y=1.66 $X2=2.615 $Y2=2.64
cc_196 VPB N_A_1370_289#_c_990_n 0.002138f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_197 VPB N_A_1370_289#_c_991_n 0.0182201f $X=-0.19 $Y=1.66 $X2=0.2 $Y2=1.58
cc_198 VPB N_A_1370_289#_c_999_n 0.0024203f $X=-0.19 $Y=1.66 $X2=0.365 $Y2=1.415
cc_199 VPB N_A_1370_289#_c_994_n 0.00166674f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_200 VPB N_A_1223_118#_c_1087_n 0.0272296f $X=-0.19 $Y=1.66 $X2=1.4 $Y2=1.415
cc_201 VPB N_A_1223_118#_c_1088_n 0.0117144f $X=-0.19 $Y=1.66 $X2=0.28 $Y2=2.65
cc_202 VPB N_A_1223_118#_c_1094_n 0.00341835f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_203 VPB N_A_1223_118#_c_1089_n 0.0153656f $X=-0.19 $Y=1.66 $X2=1.23 $Y2=1.415
cc_204 VPB N_A_1223_118#_c_1091_n 0.00370269f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_205 VPB N_A_852_74#_c_1191_n 0.0264389f $X=-0.19 $Y=1.66 $X2=2.615 $Y2=2.245
cc_206 VPB N_A_852_74#_c_1193_n 0.0768424f $X=-0.19 $Y=1.66 $X2=0.28 $Y2=0.605
cc_207 VPB N_A_852_74#_c_1208_n 0.0543622f $X=-0.19 $Y=1.66 $X2=0.2 $Y2=2.32
cc_208 VPB N_A_852_74#_c_1209_n 0.0123654f $X=-0.19 $Y=1.66 $X2=0.28 $Y2=2.49
cc_209 VPB N_A_852_74#_c_1210_n 0.0070758f $X=-0.19 $Y=1.66 $X2=0.365 $Y2=1.415
cc_210 VPB N_A_852_74#_c_1211_n 0.0191676f $X=-0.19 $Y=1.66 $X2=1.23 $Y2=1.415
cc_211 VPB N_A_852_74#_c_1212_n 0.0146102f $X=-0.19 $Y=1.66 $X2=1.23 $Y2=1.415
cc_212 VPB N_A_852_74#_c_1213_n 0.180093f $X=-0.19 $Y=1.66 $X2=2.275 $Y2=2.405
cc_213 VPB N_A_852_74#_c_1214_n 0.00747951f $X=-0.19 $Y=1.66 $X2=2.44 $Y2=2.32
cc_214 VPB N_A_852_74#_c_1215_n 0.0161081f $X=-0.19 $Y=1.66 $X2=2.44 $Y2=1.995
cc_215 VPB N_A_852_74#_M1016_g 0.00865924f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=1.415
cc_216 VPB N_A_852_74#_c_1196_n 0.0303876f $X=-0.19 $Y=1.66 $X2=0.28 $Y2=2.405
cc_217 VPB N_A_852_74#_c_1197_n 0.00515977f $X=-0.19 $Y=1.66 $X2=1.23 $Y2=1.415
cc_218 VPB N_A_852_74#_c_1219_n 0.0089867f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_219 VPB N_A_852_74#_c_1220_n 9.6535e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_220 VPB N_A_852_74#_c_1202_n 0.00324613f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_221 VPB N_A_852_74#_c_1222_n 0.00197544f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_222 VPB N_A_2006_373#_c_1391_n 0.0154015f $X=-0.19 $Y=1.66 $X2=1.475 $Y2=1.25
cc_223 VPB N_A_2006_373#_M1045_g 0.0146783f $X=-0.19 $Y=1.66 $X2=2.615 $Y2=2.64
cc_224 VPB N_A_2006_373#_c_1393_n 0.0043277f $X=-0.19 $Y=1.66 $X2=0.28 $Y2=0.605
cc_225 VPB N_A_2006_373#_c_1385_n 0.010942f $X=-0.19 $Y=1.66 $X2=0.2 $Y2=1.58
cc_226 VPB N_A_2006_373#_c_1395_n 0.00277764f $X=-0.19 $Y=1.66 $X2=0.28 $Y2=2.49
cc_227 VPB N_A_2006_373#_c_1396_n 2.07695e-19 $X=-0.19 $Y=1.66 $X2=0.28 $Y2=2.65
cc_228 VPB N_A_2006_373#_c_1397_n 0.00608544f $X=-0.19 $Y=1.66 $X2=0.445
+ $Y2=2.405
cc_229 VPB N_A_2006_373#_c_1398_n 0.0572791f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=1.415
cc_230 VPB N_A_1790_74#_c_1505_n 0.0332504f $X=-0.19 $Y=1.66 $X2=2.615 $Y2=2.64
cc_231 VPB N_A_1790_74#_c_1506_n 0.0220882f $X=-0.19 $Y=1.66 $X2=2.615 $Y2=2.64
cc_232 VPB N_A_1790_74#_c_1507_n 0.0159809f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_233 VPB N_A_1790_74#_c_1508_n 0.0160546f $X=-0.19 $Y=1.66 $X2=0.365 $Y2=1.415
cc_234 VPB N_A_1790_74#_c_1499_n 0.0202262f $X=-0.19 $Y=1.66 $X2=2.44 $Y2=2.32
cc_235 VPB N_A_1790_74#_c_1500_n 0.00804325f $X=-0.19 $Y=1.66 $X2=2.44 $Y2=1.995
cc_236 VPB N_A_1790_74#_c_1511_n 0.0246892f $X=-0.19 $Y=1.66 $X2=2.44 $Y2=1.995
cc_237 VPB N_A_1790_74#_c_1503_n 0.00737395f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_238 VPB N_A_2604_392#_c_1652_n 0.0177068f $X=-0.19 $Y=1.66 $X2=1.475 $Y2=1.25
cc_239 VPB N_A_2604_392#_c_1653_n 0.0174134f $X=-0.19 $Y=1.66 $X2=1.4 $Y2=1.415
cc_240 VPB N_A_2604_392#_c_1648_n 0.0176653f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_241 VPB N_A_2604_392#_c_1650_n 0.0195039f $X=-0.19 $Y=1.66 $X2=2.44 $Y2=2.32
cc_242 VPB N_VPWR_c_1697_n 0.00985307f $X=-0.19 $Y=1.66 $X2=2.44 $Y2=1.995
cc_243 VPB N_VPWR_c_1698_n 0.00396467f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=1.415
cc_244 VPB N_VPWR_c_1699_n 0.0080144f $X=-0.19 $Y=1.66 $X2=2.49 $Y2=1.995
cc_245 VPB N_VPWR_c_1700_n 0.0135327f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_246 VPB N_VPWR_c_1701_n 0.0511217f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_247 VPB N_VPWR_c_1702_n 0.0221602f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_248 VPB N_VPWR_c_1703_n 0.0103382f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_249 VPB N_VPWR_c_1704_n 0.0184711f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_250 VPB N_VPWR_c_1705_n 0.0109102f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_251 VPB N_VPWR_c_1706_n 0.0663373f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_252 VPB N_VPWR_c_1707_n 0.0369212f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_253 VPB N_VPWR_c_1708_n 0.00601644f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_254 VPB N_VPWR_c_1709_n 0.059824f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_255 VPB N_VPWR_c_1710_n 0.00330333f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_256 VPB N_VPWR_c_1711_n 0.0474691f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_257 VPB N_VPWR_c_1712_n 0.0237904f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_258 VPB N_VPWR_c_1713_n 0.0217361f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_259 VPB N_VPWR_c_1714_n 0.0193312f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_260 VPB N_VPWR_c_1715_n 0.0206736f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_261 VPB N_VPWR_c_1716_n 0.0174144f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_262 VPB N_VPWR_c_1717_n 0.0191515f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_263 VPB N_VPWR_c_1718_n 0.0263586f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_264 VPB N_VPWR_c_1719_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_265 VPB N_VPWR_c_1720_n 0.00330333f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_266 VPB N_VPWR_c_1721_n 0.0389406f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_267 VPB N_VPWR_c_1722_n 0.0047828f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_268 VPB N_VPWR_c_1723_n 0.00555219f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_269 VPB N_VPWR_c_1724_n 0.00614127f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_270 VPB N_VPWR_c_1696_n 0.131569f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_271 VPB N_A_388_79#_c_1888_n 0.0051238f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_272 VPB N_A_388_79#_c_1882_n 0.00481007f $X=-0.19 $Y=1.66 $X2=0.445 $Y2=2.405
cc_273 VPB N_A_388_79#_c_1890_n 0.0100423f $X=-0.19 $Y=1.66 $X2=2.44 $Y2=2.32
cc_274 VPB N_A_388_79#_c_1891_n 0.0177901f $X=-0.19 $Y=1.66 $X2=2.44 $Y2=1.995
cc_275 VPB N_A_388_79#_c_1892_n 0.00238636f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_276 VPB N_A_388_79#_c_1893_n 0.0058574f $X=-0.19 $Y=1.66 $X2=2.49 $Y2=1.995
cc_277 VPB N_A_388_79#_c_1894_n 0.00141271f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_278 VPB N_A_388_79#_c_1886_n 0.00540609f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_279 VPB N_A_388_79#_c_1896_n 0.00215028f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_280 VPB Q_N 0.00344098f $X=-0.19 $Y=1.66 $X2=1.475 $Y2=0.605
cc_281 VPB N_Q_c_2068_n 0.00405531f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_282 N_A_27_79#_c_284_n N_SCE_c_366_n 0.0181735f $X=1.4 $Y=1.415 $X2=0 $Y2=0
cc_283 N_A_27_79#_c_285_n N_SCE_c_366_n 0.0127444f $X=0.28 $Y=0.605 $X2=0 $Y2=0
cc_284 N_A_27_79#_c_286_n N_SCE_c_366_n 0.0140797f $X=0.2 $Y=2.32 $X2=0 $Y2=0
cc_285 N_A_27_79#_c_287_n N_SCE_c_366_n 0.0179605f $X=1.23 $Y=1.415 $X2=0 $Y2=0
cc_286 N_A_27_79#_c_288_n N_SCE_c_366_n 0.00851213f $X=0.24 $Y=1.415 $X2=0 $Y2=0
cc_287 N_A_27_79#_c_285_n N_SCE_c_367_n 0.00367837f $X=0.28 $Y=0.605 $X2=0 $Y2=0
cc_288 N_A_27_79#_c_286_n N_SCE_c_375_n 0.0112444f $X=0.2 $Y=2.32 $X2=0 $Y2=0
cc_289 N_A_27_79#_c_291_n N_SCE_c_375_n 0.0155777f $X=0.28 $Y=2.65 $X2=0 $Y2=0
cc_290 N_A_27_79#_c_287_n N_SCE_c_375_n 0.00644399f $X=1.23 $Y=1.415 $X2=0 $Y2=0
cc_291 N_A_27_79#_c_303_p N_SCE_c_375_n 0.0138322f $X=2.275 $Y=2.405 $X2=0 $Y2=0
cc_292 N_A_27_79#_c_293_n N_SCE_c_375_n 0.00605135f $X=0.28 $Y=2.405 $X2=0 $Y2=0
cc_293 N_A_27_79#_c_303_p N_SCE_c_376_n 0.0137373f $X=2.275 $Y=2.405 $X2=0 $Y2=0
cc_294 N_A_27_79#_c_285_n N_SCE_c_369_n 0.0100023f $X=0.28 $Y=0.605 $X2=0 $Y2=0
cc_295 N_A_27_79#_c_287_n N_SCE_c_369_n 0.00327315f $X=1.23 $Y=1.415 $X2=0 $Y2=0
cc_296 N_A_27_79#_c_289_n N_SCE_c_370_n 0.00102331f $X=2.615 $Y=2.245 $X2=0
+ $Y2=0
cc_297 N_A_27_79#_c_303_p N_SCE_c_370_n 0.0123483f $X=2.275 $Y=2.405 $X2=0 $Y2=0
cc_298 N_A_27_79#_c_292_n N_SCE_c_370_n 0.0109466f $X=2.44 $Y=1.995 $X2=0 $Y2=0
cc_299 N_A_27_79#_c_284_n N_SCE_c_371_n 0.00219996f $X=1.4 $Y=1.415 $X2=0 $Y2=0
cc_300 N_A_27_79#_c_287_n N_SCE_c_371_n 0.0155382f $X=1.23 $Y=1.415 $X2=0 $Y2=0
cc_301 N_A_27_79#_c_289_n N_SCE_c_372_n 0.00192643f $X=2.615 $Y=2.245 $X2=0
+ $Y2=0
cc_302 N_A_27_79#_c_292_n N_SCE_c_372_n 0.0221869f $X=2.44 $Y=1.995 $X2=0 $Y2=0
cc_303 N_A_27_79#_c_289_n N_SCE_c_373_n 0.0202521f $X=2.615 $Y=2.245 $X2=0 $Y2=0
cc_304 N_A_27_79#_c_292_n N_SCE_c_373_n 7.02495e-19 $X=2.44 $Y=1.995 $X2=0 $Y2=0
cc_305 N_A_27_79#_c_284_n N_SCE_c_378_n 0.0448734f $X=1.4 $Y=1.415 $X2=0 $Y2=0
cc_306 N_A_27_79#_c_287_n N_SCE_c_378_n 0.00247218f $X=1.23 $Y=1.415 $X2=0 $Y2=0
cc_307 N_A_27_79#_c_303_p N_SCE_c_378_n 0.0171512f $X=2.275 $Y=2.405 $X2=0 $Y2=0
cc_308 N_A_27_79#_c_284_n N_SCE_c_379_n 0.00363355f $X=1.4 $Y=1.415 $X2=0 $Y2=0
cc_309 N_A_27_79#_c_286_n N_SCE_c_379_n 0.0192999f $X=0.2 $Y=2.32 $X2=0 $Y2=0
cc_310 N_A_27_79#_c_287_n N_SCE_c_379_n 0.0494351f $X=1.23 $Y=1.415 $X2=0 $Y2=0
cc_311 N_A_27_79#_c_303_p N_SCE_c_379_n 0.0736349f $X=2.275 $Y=2.405 $X2=0 $Y2=0
cc_312 N_A_27_79#_c_289_n N_D_c_452_n 0.0130861f $X=2.615 $Y=2.245 $X2=0 $Y2=0
cc_313 N_A_27_79#_c_284_n N_D_c_452_n 0.0185925f $X=1.4 $Y=1.415 $X2=0 $Y2=0
cc_314 N_A_27_79#_c_287_n N_D_c_452_n 6.63701e-19 $X=1.23 $Y=1.415 $X2=0 $Y2=0
cc_315 N_A_27_79#_c_292_n N_D_c_452_n 0.00129661f $X=2.44 $Y=1.995 $X2=0 $Y2=0
cc_316 N_A_27_79#_c_289_n N_D_c_457_n 0.0173318f $X=2.615 $Y=2.245 $X2=0 $Y2=0
cc_317 N_A_27_79#_c_303_p N_D_c_457_n 0.0174363f $X=2.275 $Y=2.405 $X2=0 $Y2=0
cc_318 N_A_27_79#_c_292_n N_D_c_457_n 0.00352705f $X=2.44 $Y=1.995 $X2=0 $Y2=0
cc_319 N_A_27_79#_M1014_g N_D_c_453_n 0.0200462f $X=1.475 $Y=0.605 $X2=0 $Y2=0
cc_320 N_A_27_79#_M1014_g N_D_c_454_n 0.0109288f $X=1.475 $Y=0.605 $X2=0 $Y2=0
cc_321 N_A_27_79#_M1014_g N_D_c_455_n 0.03521f $X=1.475 $Y=0.605 $X2=0 $Y2=0
cc_322 N_A_27_79#_c_289_n N_SCD_c_503_n 0.0359696f $X=2.615 $Y=2.245 $X2=-0.19
+ $Y2=-0.245
cc_323 N_A_27_79#_c_292_n N_SCD_c_503_n 3.88432e-19 $X=2.44 $Y=1.995 $X2=-0.19
+ $Y2=-0.245
cc_324 N_A_27_79#_c_289_n N_SCD_c_500_n 0.0223785f $X=2.615 $Y=2.245 $X2=0 $Y2=0
cc_325 N_A_27_79#_c_292_n N_SCD_c_500_n 0.00149955f $X=2.44 $Y=1.995 $X2=0 $Y2=0
cc_326 N_A_27_79#_c_289_n SCD 0.00131261f $X=2.615 $Y=2.245 $X2=0 $Y2=0
cc_327 N_A_27_79#_c_292_n SCD 0.0137554f $X=2.44 $Y=1.995 $X2=0 $Y2=0
cc_328 N_A_27_79#_c_303_p N_VPWR_M1023_d 0.0181551f $X=2.275 $Y=2.405 $X2=-0.19
+ $Y2=-0.245
cc_329 N_A_27_79#_c_289_n N_VPWR_c_1711_n 0.00300876f $X=2.615 $Y=2.245 $X2=0
+ $Y2=0
cc_330 N_A_27_79#_c_291_n N_VPWR_c_1717_n 0.0145785f $X=0.28 $Y=2.65 $X2=0 $Y2=0
cc_331 N_A_27_79#_c_291_n N_VPWR_c_1718_n 0.0102732f $X=0.28 $Y=2.65 $X2=0 $Y2=0
cc_332 N_A_27_79#_c_303_p N_VPWR_c_1718_n 0.0418977f $X=2.275 $Y=2.405 $X2=0
+ $Y2=0
cc_333 N_A_27_79#_c_289_n N_VPWR_c_1696_n 0.00370805f $X=2.615 $Y=2.245 $X2=0
+ $Y2=0
cc_334 N_A_27_79#_c_291_n N_VPWR_c_1696_n 0.0120406f $X=0.28 $Y=2.65 $X2=0 $Y2=0
cc_335 N_A_27_79#_c_303_p N_VPWR_c_1696_n 0.0250254f $X=2.275 $Y=2.405 $X2=0
+ $Y2=0
cc_336 N_A_27_79#_c_303_p A_307_464# 0.00479553f $X=2.275 $Y=2.405 $X2=-0.19
+ $Y2=-0.245
cc_337 N_A_27_79#_c_303_p N_A_388_79#_M1035_d 0.0167952f $X=2.275 $Y=2.405 $X2=0
+ $Y2=0
cc_338 N_A_27_79#_c_289_n N_A_388_79#_c_1898_n 0.0181967f $X=2.615 $Y=2.245
+ $X2=0 $Y2=0
cc_339 N_A_27_79#_c_303_p N_A_388_79#_c_1898_n 0.0419607f $X=2.275 $Y=2.405
+ $X2=0 $Y2=0
cc_340 N_A_27_79#_c_289_n N_A_388_79#_c_1900_n 0.00384668f $X=2.615 $Y=2.245
+ $X2=0 $Y2=0
cc_341 N_A_27_79#_c_289_n N_A_388_79#_c_1888_n 0.0012654f $X=2.615 $Y=2.245
+ $X2=0 $Y2=0
cc_342 N_A_27_79#_c_303_p N_A_388_79#_c_1888_n 0.0148585f $X=2.275 $Y=2.405
+ $X2=0 $Y2=0
cc_343 N_A_27_79#_M1014_g N_VGND_c_2084_n 5.90987e-19 $X=1.475 $Y=0.605 $X2=0
+ $Y2=0
cc_344 N_A_27_79#_c_284_n N_VGND_c_2084_n 0.00297438f $X=1.4 $Y=1.415 $X2=0
+ $Y2=0
cc_345 N_A_27_79#_c_285_n N_VGND_c_2084_n 0.0179429f $X=0.28 $Y=0.605 $X2=0
+ $Y2=0
cc_346 N_A_27_79#_c_287_n N_VGND_c_2084_n 0.0148785f $X=1.23 $Y=1.415 $X2=0
+ $Y2=0
cc_347 N_A_27_79#_M1014_g N_VGND_c_2094_n 9.44495e-19 $X=1.475 $Y=0.605 $X2=0
+ $Y2=0
cc_348 N_A_27_79#_c_285_n N_VGND_c_2100_n 0.0100552f $X=0.28 $Y=0.605 $X2=0
+ $Y2=0
cc_349 N_A_27_79#_c_285_n N_VGND_c_2110_n 0.00902019f $X=0.28 $Y=0.605 $X2=0
+ $Y2=0
cc_350 N_A_27_79#_M1014_g N_noxref_25_c_2241_n 7.43016e-19 $X=1.475 $Y=0.605
+ $X2=0 $Y2=0
cc_351 N_A_27_79#_c_284_n N_noxref_25_c_2241_n 0.0048989f $X=1.4 $Y=1.415 $X2=0
+ $Y2=0
cc_352 N_A_27_79#_c_287_n N_noxref_25_c_2241_n 0.0106151f $X=1.23 $Y=1.415 $X2=0
+ $Y2=0
cc_353 N_A_27_79#_M1014_g N_noxref_25_c_2242_n 0.0154771f $X=1.475 $Y=0.605
+ $X2=0 $Y2=0
cc_354 N_SCE_c_376_n N_D_c_452_n 0.0238606f $X=1.46 $Y=2.245 $X2=0 $Y2=0
cc_355 N_SCE_M1034_g N_D_c_452_n 8.48778e-19 $X=2.66 $Y=0.605 $X2=0 $Y2=0
cc_356 N_SCE_c_370_n N_D_c_452_n 0.0202953f $X=1.71 $Y=1.82 $X2=0 $Y2=0
cc_357 N_SCE_c_371_n N_D_c_452_n 0.00239218f $X=1.795 $Y=1.49 $X2=0 $Y2=0
cc_358 N_SCE_c_372_n N_D_c_452_n 0.0188764f $X=2.57 $Y=1.455 $X2=0 $Y2=0
cc_359 N_SCE_c_373_n N_D_c_452_n 0.00894005f $X=2.57 $Y=1.455 $X2=0 $Y2=0
cc_360 N_SCE_c_376_n N_D_c_457_n 0.0403591f $X=1.46 $Y=2.245 $X2=0 $Y2=0
cc_361 N_SCE_M1034_g N_D_c_453_n 0.00730331f $X=2.66 $Y=0.605 $X2=0 $Y2=0
cc_362 N_SCE_c_371_n N_D_c_453_n 7.56204e-19 $X=1.795 $Y=1.49 $X2=0 $Y2=0
cc_363 N_SCE_c_372_n N_D_c_453_n 0.002936f $X=2.57 $Y=1.455 $X2=0 $Y2=0
cc_364 N_SCE_M1034_g N_D_c_454_n 5.42624e-19 $X=2.66 $Y=0.605 $X2=0 $Y2=0
cc_365 N_SCE_c_371_n N_D_c_454_n 0.0150217f $X=1.795 $Y=1.49 $X2=0 $Y2=0
cc_366 N_SCE_c_372_n N_D_c_454_n 0.0224216f $X=2.57 $Y=1.455 $X2=0 $Y2=0
cc_367 N_SCE_c_379_n N_D_c_454_n 0.0020111f $X=1.625 $Y=1.985 $X2=0 $Y2=0
cc_368 N_SCE_M1034_g N_D_c_455_n 0.00705002f $X=2.66 $Y=0.605 $X2=0 $Y2=0
cc_369 N_SCE_M1034_g N_SCD_M1015_g 0.0628756f $X=2.66 $Y=0.605 $X2=0 $Y2=0
cc_370 N_SCE_c_372_n N_SCD_M1015_g 5.04484e-19 $X=2.57 $Y=1.455 $X2=0 $Y2=0
cc_371 N_SCE_c_372_n SCD 0.0120234f $X=2.57 $Y=1.455 $X2=0 $Y2=0
cc_372 N_SCE_c_373_n SCD 2.2546e-19 $X=2.57 $Y=1.455 $X2=0 $Y2=0
cc_373 N_SCE_c_372_n N_SCD_c_502_n 6.19299e-19 $X=2.57 $Y=1.455 $X2=0 $Y2=0
cc_374 N_SCE_c_373_n N_SCD_c_502_n 0.0113035f $X=2.57 $Y=1.455 $X2=0 $Y2=0
cc_375 N_SCE_c_376_n N_VPWR_c_1711_n 0.00413917f $X=1.46 $Y=2.245 $X2=0 $Y2=0
cc_376 N_SCE_c_375_n N_VPWR_c_1717_n 0.00445602f $X=0.505 $Y=2.245 $X2=0 $Y2=0
cc_377 N_SCE_c_375_n N_VPWR_c_1718_n 0.0101493f $X=0.505 $Y=2.245 $X2=0 $Y2=0
cc_378 N_SCE_c_376_n N_VPWR_c_1718_n 0.0101104f $X=1.46 $Y=2.245 $X2=0 $Y2=0
cc_379 N_SCE_c_375_n N_VPWR_c_1696_n 0.00460319f $X=0.505 $Y=2.245 $X2=0 $Y2=0
cc_380 N_SCE_c_376_n N_VPWR_c_1696_n 0.00412661f $X=1.46 $Y=2.245 $X2=0 $Y2=0
cc_381 N_SCE_c_376_n N_A_388_79#_c_1898_n 8.44751e-19 $X=1.46 $Y=2.245 $X2=0
+ $Y2=0
cc_382 N_SCE_M1034_g N_A_388_79#_c_1879_n 0.0103246f $X=2.66 $Y=0.605 $X2=0
+ $Y2=0
cc_383 N_SCE_M1034_g N_A_388_79#_c_1880_n 0.0087327f $X=2.66 $Y=0.605 $X2=0
+ $Y2=0
cc_384 N_SCE_c_372_n N_A_388_79#_c_1880_n 0.00815275f $X=2.57 $Y=1.455 $X2=0
+ $Y2=0
cc_385 N_SCE_M1034_g N_A_388_79#_c_1881_n 0.00327429f $X=2.66 $Y=0.605 $X2=0
+ $Y2=0
cc_386 N_SCE_c_372_n N_A_388_79#_c_1881_n 0.0273677f $X=2.57 $Y=1.455 $X2=0
+ $Y2=0
cc_387 N_SCE_c_373_n N_A_388_79#_c_1881_n 0.00449985f $X=2.57 $Y=1.455 $X2=0
+ $Y2=0
cc_388 N_SCE_c_367_n N_VGND_c_2084_n 0.0143331f $X=0.495 $Y=0.89 $X2=0 $Y2=0
cc_389 N_SCE_M1034_g N_VGND_c_2094_n 9.44495e-19 $X=2.66 $Y=0.605 $X2=0 $Y2=0
cc_390 N_SCE_c_367_n N_VGND_c_2100_n 0.00465077f $X=0.495 $Y=0.89 $X2=0 $Y2=0
cc_391 N_SCE_c_367_n N_VGND_c_2110_n 0.00451796f $X=0.495 $Y=0.89 $X2=0 $Y2=0
cc_392 N_SCE_c_367_n N_noxref_25_c_2241_n 7.27954e-19 $X=0.495 $Y=0.89 $X2=0
+ $Y2=0
cc_393 N_SCE_M1034_g N_noxref_25_c_2242_n 0.0128121f $X=2.66 $Y=0.605 $X2=0
+ $Y2=0
cc_394 N_SCE_c_367_n N_noxref_25_c_2243_n 6.46792e-19 $X=0.495 $Y=0.89 $X2=0
+ $Y2=0
cc_395 N_SCE_M1034_g N_noxref_25_c_2244_n 0.00151906f $X=2.66 $Y=0.605 $X2=0
+ $Y2=0
cc_396 N_D_c_457_n N_VPWR_c_1711_n 0.00445405f $X=1.88 $Y=2.245 $X2=0 $Y2=0
cc_397 N_D_c_457_n N_VPWR_c_1718_n 0.00139022f $X=1.88 $Y=2.245 $X2=0 $Y2=0
cc_398 N_D_c_457_n N_VPWR_c_1696_n 0.00457269f $X=1.88 $Y=2.245 $X2=0 $Y2=0
cc_399 N_D_c_454_n N_A_388_79#_M1029_d 0.00145733f $X=1.925 $Y=1.09 $X2=-0.19
+ $Y2=-0.245
cc_400 N_D_c_457_n N_A_388_79#_c_1898_n 0.00949498f $X=1.88 $Y=2.245 $X2=0 $Y2=0
cc_401 N_D_c_453_n N_A_388_79#_c_1879_n 3.29098e-19 $X=1.925 $Y=1.09 $X2=0 $Y2=0
cc_402 N_D_c_454_n N_A_388_79#_c_1879_n 0.0164816f $X=1.925 $Y=1.09 $X2=0 $Y2=0
cc_403 N_D_c_455_n N_A_388_79#_c_1879_n 0.00523412f $X=1.925 $Y=0.925 $X2=0
+ $Y2=0
cc_404 N_D_c_453_n N_A_388_79#_c_1881_n 7.8315e-19 $X=1.925 $Y=1.09 $X2=0 $Y2=0
cc_405 N_D_c_454_n N_A_388_79#_c_1881_n 0.0148785f $X=1.925 $Y=1.09 $X2=0 $Y2=0
cc_406 N_D_c_455_n N_VGND_c_2094_n 9.44495e-19 $X=1.925 $Y=0.925 $X2=0 $Y2=0
cc_407 N_D_c_454_n N_noxref_25_c_2241_n 0.00134475f $X=1.925 $Y=1.09 $X2=0 $Y2=0
cc_408 N_D_c_453_n N_noxref_25_c_2242_n 5.75063e-19 $X=1.925 $Y=1.09 $X2=0 $Y2=0
cc_409 N_D_c_454_n N_noxref_25_c_2242_n 0.0127007f $X=1.925 $Y=1.09 $X2=0 $Y2=0
cc_410 N_D_c_455_n N_noxref_25_c_2242_n 0.0123465f $X=1.925 $Y=0.925 $X2=0 $Y2=0
cc_411 N_D_c_454_n noxref_26 0.00197445f $X=1.925 $Y=1.09 $X2=-0.19 $Y2=-0.245
cc_412 N_SCD_M1015_g N_RESET_B_M1043_g 0.0270106f $X=3.05 $Y=0.605 $X2=0 $Y2=0
cc_413 SCD N_RESET_B_M1043_g 7.42142e-19 $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_414 N_SCD_c_502_n N_RESET_B_M1043_g 0.0175943f $X=3.11 $Y=1.605 $X2=0 $Y2=0
cc_415 N_SCD_c_503_n N_RESET_B_c_551_n 0.0148831f $X=3.035 $Y=2.245 $X2=0 $Y2=0
cc_416 N_SCD_c_500_n N_RESET_B_c_562_n 0.0213043f $X=3.11 $Y=1.945 $X2=0 $Y2=0
cc_417 N_SCD_c_503_n N_VPWR_c_1697_n 0.00395262f $X=3.035 $Y=2.245 $X2=0 $Y2=0
cc_418 N_SCD_c_503_n N_VPWR_c_1711_n 0.00461464f $X=3.035 $Y=2.245 $X2=0 $Y2=0
cc_419 N_SCD_c_503_n N_VPWR_c_1696_n 0.00463738f $X=3.035 $Y=2.245 $X2=0 $Y2=0
cc_420 N_SCD_M1015_g N_A_388_79#_c_1879_n 0.00151803f $X=3.05 $Y=0.605 $X2=0
+ $Y2=0
cc_421 N_SCD_M1015_g N_A_388_79#_c_1880_n 0.0128888f $X=3.05 $Y=0.605 $X2=0
+ $Y2=0
cc_422 SCD N_A_388_79#_c_1880_n 0.0182456f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_423 N_SCD_c_502_n N_A_388_79#_c_1880_n 0.00113125f $X=3.11 $Y=1.605 $X2=0
+ $Y2=0
cc_424 N_SCD_c_503_n N_A_388_79#_c_1921_n 0.011884f $X=3.035 $Y=2.245 $X2=0
+ $Y2=0
cc_425 N_SCD_c_500_n N_A_388_79#_c_1921_n 8.43385e-19 $X=3.11 $Y=1.945 $X2=0
+ $Y2=0
cc_426 SCD N_A_388_79#_c_1921_n 0.023597f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_427 N_SCD_c_503_n N_A_388_79#_c_1882_n 0.00133602f $X=3.035 $Y=2.245 $X2=0
+ $Y2=0
cc_428 N_SCD_M1015_g N_A_388_79#_c_1882_n 0.00479317f $X=3.05 $Y=0.605 $X2=0
+ $Y2=0
cc_429 N_SCD_c_500_n N_A_388_79#_c_1882_n 0.00183512f $X=3.11 $Y=1.945 $X2=0
+ $Y2=0
cc_430 SCD N_A_388_79#_c_1882_n 0.0534507f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_431 N_SCD_c_502_n N_A_388_79#_c_1882_n 0.003794f $X=3.11 $Y=1.605 $X2=0 $Y2=0
cc_432 N_SCD_c_503_n N_A_388_79#_c_1890_n 3.42916e-19 $X=3.035 $Y=2.245 $X2=0
+ $Y2=0
cc_433 N_SCD_M1015_g N_VGND_c_2085_n 2.31759e-19 $X=3.05 $Y=0.605 $X2=0 $Y2=0
cc_434 N_SCD_M1015_g N_VGND_c_2094_n 9.63557e-19 $X=3.05 $Y=0.605 $X2=0 $Y2=0
cc_435 N_SCD_M1015_g N_noxref_25_c_2242_n 0.0111117f $X=3.05 $Y=0.605 $X2=0
+ $Y2=0
cc_436 N_SCD_M1015_g N_noxref_25_c_2244_n 0.00776653f $X=3.05 $Y=0.605 $X2=0
+ $Y2=0
cc_437 N_RESET_B_c_557_n N_CLK_c_734_n 0.00211211f $X=7.775 $Y=2.035 $X2=0 $Y2=0
cc_438 N_RESET_B_c_562_n N_CLK_c_734_n 0.00402257f $X=3.605 $Y=2.032 $X2=0 $Y2=0
cc_439 N_RESET_B_c_563_n N_CLK_c_734_n 4.17832e-19 $X=3.95 $Y=1.985 $X2=0 $Y2=0
cc_440 N_RESET_B_M1043_g N_CLK_c_735_n 0.0173986f $X=3.59 $Y=0.605 $X2=0 $Y2=0
cc_441 N_RESET_B_c_557_n N_CLK_c_735_n 0.00213186f $X=7.775 $Y=2.035 $X2=0 $Y2=0
cc_442 N_RESET_B_c_562_n N_CLK_c_735_n 0.00970285f $X=3.605 $Y=2.032 $X2=0 $Y2=0
cc_443 N_RESET_B_c_563_n N_CLK_c_735_n 6.11048e-19 $X=3.95 $Y=1.985 $X2=0 $Y2=0
cc_444 N_RESET_B_M1043_g CLK 0.00186105f $X=3.59 $Y=0.605 $X2=0 $Y2=0
cc_445 N_RESET_B_c_557_n CLK 2.97792e-19 $X=7.775 $Y=2.035 $X2=0 $Y2=0
cc_446 N_RESET_B_c_558_n CLK 0.00364034f $X=4.225 $Y=2.035 $X2=0 $Y2=0
cc_447 N_RESET_B_c_562_n CLK 8.03812e-19 $X=3.605 $Y=2.032 $X2=0 $Y2=0
cc_448 N_RESET_B_c_563_n CLK 0.0122967f $X=3.95 $Y=1.985 $X2=0 $Y2=0
cc_449 N_RESET_B_c_557_n N_A_1025_74#_c_806_n 0.00324919f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_450 N_RESET_B_c_557_n N_A_1025_74#_c_785_n 0.00395271f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_451 N_RESET_B_c_559_n N_A_1025_74#_c_808_n 0.00170256f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_452 N_RESET_B_c_557_n N_A_1025_74#_c_794_n 0.0318868f $X=7.775 $Y=2.035 $X2=0
+ $Y2=0
cc_453 N_RESET_B_c_557_n N_A_1025_74#_c_795_n 0.0136592f $X=7.775 $Y=2.035 $X2=0
+ $Y2=0
cc_454 N_RESET_B_c_544_n N_A_1025_74#_c_796_n 0.0115453f $X=7.32 $Y=1.085 $X2=0
+ $Y2=0
cc_455 N_RESET_B_c_545_n N_A_1025_74#_c_796_n 0.00187511f $X=7.66 $Y=1.16 $X2=0
+ $Y2=0
cc_456 N_RESET_B_c_544_n N_A_1025_74#_c_801_n 0.00299808f $X=7.32 $Y=1.085 $X2=0
+ $Y2=0
cc_457 N_RESET_B_c_559_n N_A_1025_74#_c_811_n 0.0277328f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_458 N_RESET_B_c_557_n N_A_1025_74#_c_805_n 0.00369615f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_459 N_RESET_B_c_559_n N_A_1370_289#_M1011_d 0.00455663f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_460 N_RESET_B_c_547_n N_A_1370_289#_c_995_n 0.00171141f $X=7.735 $Y=1.795
+ $X2=0 $Y2=0
cc_461 N_RESET_B_c_557_n N_A_1370_289#_c_995_n 0.0118939f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_462 N_RESET_B_c_564_n N_A_1370_289#_c_995_n 0.00541842f $X=7.735 $Y=2.002
+ $X2=0 $Y2=0
cc_463 N_RESET_B_c_544_n N_A_1370_289#_M1001_g 0.0413638f $X=7.32 $Y=1.085 $X2=0
+ $Y2=0
cc_464 N_RESET_B_c_547_n N_A_1370_289#_M1001_g 0.00134145f $X=7.735 $Y=1.795
+ $X2=0 $Y2=0
cc_465 N_RESET_B_c_552_n N_A_1370_289#_c_996_n 0.0148016f $X=7.525 $Y=2.21 $X2=0
+ $Y2=0
cc_466 N_RESET_B_c_546_n N_A_1370_289#_c_990_n 0.00378904f $X=7.395 $Y=1.16
+ $X2=0 $Y2=0
cc_467 N_RESET_B_c_547_n N_A_1370_289#_c_990_n 4.21074e-19 $X=7.735 $Y=1.795
+ $X2=0 $Y2=0
cc_468 N_RESET_B_c_557_n N_A_1370_289#_c_990_n 0.006336f $X=7.775 $Y=2.035 $X2=0
+ $Y2=0
cc_469 N_RESET_B_c_546_n N_A_1370_289#_c_991_n 0.00184819f $X=7.395 $Y=1.16
+ $X2=0 $Y2=0
cc_470 N_RESET_B_c_547_n N_A_1370_289#_c_991_n 0.00820554f $X=7.735 $Y=1.795
+ $X2=0 $Y2=0
cc_471 N_RESET_B_c_557_n N_A_1370_289#_c_991_n 0.00145503f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_472 N_RESET_B_c_559_n N_A_1370_289#_c_999_n 0.0380147f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_473 N_RESET_B_c_544_n N_A_1370_289#_c_992_n 0.00994147f $X=7.32 $Y=1.085
+ $X2=0 $Y2=0
cc_474 N_RESET_B_c_545_n N_A_1370_289#_c_992_n 0.011861f $X=7.66 $Y=1.16 $X2=0
+ $Y2=0
cc_475 N_RESET_B_c_546_n N_A_1370_289#_c_992_n 0.00476761f $X=7.395 $Y=1.16
+ $X2=0 $Y2=0
cc_476 N_RESET_B_c_545_n N_A_1223_118#_M1003_g 0.00470516f $X=7.66 $Y=1.16 $X2=0
+ $Y2=0
cc_477 N_RESET_B_c_547_n N_A_1223_118#_c_1087_n 0.0123408f $X=7.735 $Y=1.795
+ $X2=0 $Y2=0
cc_478 N_RESET_B_c_559_n N_A_1223_118#_c_1087_n 0.00747349f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_479 N_RESET_B_c_557_n N_A_1223_118#_c_1088_n 0.0243758f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_480 N_RESET_B_c_557_n N_A_1223_118#_c_1101_n 0.0192265f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_481 N_RESET_B_c_557_n N_A_1223_118#_c_1094_n 0.00963546f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_482 N_RESET_B_c_552_n N_A_1223_118#_c_1089_n 0.0169766f $X=7.525 $Y=2.21
+ $X2=0 $Y2=0
cc_483 N_RESET_B_c_547_n N_A_1223_118#_c_1089_n 0.00612906f $X=7.735 $Y=1.795
+ $X2=0 $Y2=0
cc_484 N_RESET_B_c_557_n N_A_1223_118#_c_1089_n 0.0319772f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_485 N_RESET_B_c_560_n N_A_1223_118#_c_1089_n 0.00394987f $X=8.065 $Y=2.035
+ $X2=0 $Y2=0
cc_486 N_RESET_B_c_564_n N_A_1223_118#_c_1089_n 0.0177116f $X=7.735 $Y=2.002
+ $X2=0 $Y2=0
cc_487 N_RESET_B_c_565_n N_A_1223_118#_c_1089_n 0.0379481f $X=7.825 $Y=1.96
+ $X2=0 $Y2=0
cc_488 N_RESET_B_c_546_n N_A_1223_118#_c_1090_n 0.00417742f $X=7.395 $Y=1.16
+ $X2=0 $Y2=0
cc_489 N_RESET_B_c_545_n N_A_1223_118#_c_1091_n 0.00253033f $X=7.66 $Y=1.16
+ $X2=0 $Y2=0
cc_490 N_RESET_B_c_547_n N_A_1223_118#_c_1091_n 0.0179025f $X=7.735 $Y=1.795
+ $X2=0 $Y2=0
cc_491 N_RESET_B_c_557_n N_A_1223_118#_c_1091_n 0.00645679f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_492 N_RESET_B_c_559_n N_A_1223_118#_c_1091_n 0.0108792f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_493 N_RESET_B_c_560_n N_A_1223_118#_c_1091_n 0.00336108f $X=8.065 $Y=2.035
+ $X2=0 $Y2=0
cc_494 N_RESET_B_c_564_n N_A_1223_118#_c_1091_n 0.00671537f $X=7.735 $Y=2.002
+ $X2=0 $Y2=0
cc_495 N_RESET_B_c_565_n N_A_1223_118#_c_1091_n 0.0174718f $X=7.825 $Y=1.96
+ $X2=0 $Y2=0
cc_496 N_RESET_B_c_557_n N_A_852_74#_M1022_s 0.00155813f $X=7.775 $Y=2.035 $X2=0
+ $Y2=0
cc_497 N_RESET_B_c_557_n N_A_852_74#_c_1191_n 0.00462237f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_498 N_RESET_B_c_557_n N_A_852_74#_c_1193_n 0.0014923f $X=7.775 $Y=2.035 $X2=0
+ $Y2=0
cc_499 N_RESET_B_c_557_n N_A_852_74#_c_1212_n 0.00255127f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_500 N_RESET_B_c_552_n N_A_852_74#_c_1213_n 0.00850098f $X=7.525 $Y=2.21 $X2=0
+ $Y2=0
cc_501 N_RESET_B_c_559_n N_A_852_74#_M1016_g 0.00873993f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_502 N_RESET_B_c_559_n N_A_852_74#_c_1196_n 0.00840564f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_503 N_RESET_B_c_559_n N_A_852_74#_c_1197_n 3.03408e-19 $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_504 N_RESET_B_M1043_g N_A_852_74#_c_1200_n 0.00531801f $X=3.59 $Y=0.605 $X2=0
+ $Y2=0
cc_505 N_RESET_B_c_557_n N_A_852_74#_c_1232_n 9.69099e-19 $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_506 N_RESET_B_c_557_n N_A_852_74#_c_1220_n 0.0111029f $X=7.775 $Y=2.035 $X2=0
+ $Y2=0
cc_507 N_RESET_B_c_557_n N_A_852_74#_c_1222_n 0.0150959f $X=7.775 $Y=2.035 $X2=0
+ $Y2=0
cc_508 N_RESET_B_c_558_n N_A_852_74#_c_1222_n 0.00279861f $X=4.225 $Y=2.035
+ $X2=0 $Y2=0
cc_509 N_RESET_B_c_562_n N_A_852_74#_c_1222_n 0.00169098f $X=3.605 $Y=2.032
+ $X2=0 $Y2=0
cc_510 N_RESET_B_c_563_n N_A_852_74#_c_1222_n 0.0240323f $X=3.95 $Y=1.985 $X2=0
+ $Y2=0
cc_511 N_RESET_B_c_557_n N_A_852_74#_c_1204_n 0.00121003f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_512 N_RESET_B_c_557_n N_A_852_74#_c_1205_n 0.00750094f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_513 N_RESET_B_M1027_g N_A_2006_373#_M1045_g 0.0455699f $X=10.715 $Y=0.58
+ $X2=0 $Y2=0
cc_514 N_RESET_B_c_554_n N_A_2006_373#_M1045_g 0.00569933f $X=10.855 $Y=1.82
+ $X2=0 $Y2=0
cc_515 N_RESET_B_c_554_n N_A_2006_373#_c_1393_n 0.00379957f $X=10.855 $Y=1.82
+ $X2=0 $Y2=0
cc_516 N_RESET_B_c_555_n N_A_2006_373#_c_1393_n 0.00369134f $X=11.005 $Y=2.28
+ $X2=0 $Y2=0
cc_517 N_RESET_B_c_559_n N_A_2006_373#_c_1393_n 0.0257703f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_518 RESET_B N_A_2006_373#_c_1393_n 0.00275621f $X=10.715 $Y=1.95 $X2=0 $Y2=0
cc_519 N_RESET_B_c_566_n N_A_2006_373#_c_1393_n 0.0241058f $X=10.8 $Y=2.035
+ $X2=0 $Y2=0
cc_520 N_RESET_B_c_554_n N_A_2006_373#_c_1385_n 0.00306368f $X=10.855 $Y=1.82
+ $X2=0 $Y2=0
cc_521 N_RESET_B_c_555_n N_A_2006_373#_c_1385_n 0.0031248f $X=11.005 $Y=2.28
+ $X2=0 $Y2=0
cc_522 N_RESET_B_c_549_n N_A_2006_373#_c_1385_n 0.012737f $X=10.855 $Y=1.55
+ $X2=0 $Y2=0
cc_523 N_RESET_B_c_559_n N_A_2006_373#_c_1385_n 0.00282721f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_524 RESET_B N_A_2006_373#_c_1385_n 0.00310808f $X=10.715 $Y=1.95 $X2=0 $Y2=0
cc_525 N_RESET_B_c_566_n N_A_2006_373#_c_1385_n 0.0505438f $X=10.8 $Y=2.035
+ $X2=0 $Y2=0
cc_526 N_RESET_B_c_555_n N_A_2006_373#_c_1395_n 0.0144067f $X=11.005 $Y=2.28
+ $X2=0 $Y2=0
cc_527 N_RESET_B_c_549_n N_A_2006_373#_c_1395_n 4.02079e-19 $X=10.855 $Y=1.55
+ $X2=0 $Y2=0
cc_528 N_RESET_B_c_559_n N_A_2006_373#_c_1395_n 0.00318931f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_529 RESET_B N_A_2006_373#_c_1395_n 0.0077273f $X=10.715 $Y=1.95 $X2=0 $Y2=0
cc_530 N_RESET_B_c_566_n N_A_2006_373#_c_1395_n 0.0232665f $X=10.8 $Y=2.035
+ $X2=0 $Y2=0
cc_531 N_RESET_B_M1027_g N_A_2006_373#_c_1387_n 9.65407e-19 $X=10.715 $Y=0.58
+ $X2=0 $Y2=0
cc_532 N_RESET_B_M1027_g N_A_2006_373#_c_1389_n 6.07222e-19 $X=10.715 $Y=0.58
+ $X2=0 $Y2=0
cc_533 N_RESET_B_c_555_n N_A_2006_373#_c_1397_n 0.0117118f $X=11.005 $Y=2.28
+ $X2=0 $Y2=0
cc_534 N_RESET_B_c_566_n N_A_2006_373#_c_1397_n 0.0277898f $X=10.8 $Y=2.035
+ $X2=0 $Y2=0
cc_535 N_RESET_B_c_555_n N_A_2006_373#_c_1398_n 0.0215739f $X=11.005 $Y=2.28
+ $X2=0 $Y2=0
cc_536 N_RESET_B_c_559_n N_A_2006_373#_c_1398_n 0.0142613f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_537 RESET_B N_A_2006_373#_c_1398_n 0.00149024f $X=10.715 $Y=1.95 $X2=0 $Y2=0
cc_538 N_RESET_B_c_566_n N_A_2006_373#_c_1398_n 0.00155699f $X=10.8 $Y=2.035
+ $X2=0 $Y2=0
cc_539 N_RESET_B_c_559_n N_A_1790_74#_M1016_d 0.00975786f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_540 N_RESET_B_M1027_g N_A_1790_74#_M1018_g 0.0556926f $X=10.715 $Y=0.58 $X2=0
+ $Y2=0
cc_541 N_RESET_B_M1027_g N_A_1790_74#_c_1495_n 0.0094439f $X=10.715 $Y=0.58
+ $X2=0 $Y2=0
cc_542 N_RESET_B_c_555_n N_A_1790_74#_c_1495_n 0.00125789f $X=11.005 $Y=2.28
+ $X2=0 $Y2=0
cc_543 N_RESET_B_c_549_n N_A_1790_74#_c_1495_n 0.00511143f $X=10.855 $Y=1.55
+ $X2=0 $Y2=0
cc_544 N_RESET_B_c_554_n N_A_1790_74#_c_1505_n 0.00511143f $X=10.855 $Y=1.82
+ $X2=0 $Y2=0
cc_545 N_RESET_B_c_555_n N_A_1790_74#_c_1505_n 0.0232392f $X=11.005 $Y=2.28
+ $X2=0 $Y2=0
cc_546 N_RESET_B_c_566_n N_A_1790_74#_c_1505_n 0.0083262f $X=10.8 $Y=2.035 $X2=0
+ $Y2=0
cc_547 N_RESET_B_c_555_n N_A_1790_74#_c_1506_n 0.00947913f $X=11.005 $Y=2.28
+ $X2=0 $Y2=0
cc_548 N_RESET_B_c_559_n N_A_1790_74#_c_1522_n 0.0195683f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_549 N_RESET_B_c_559_n N_A_1790_74#_c_1503_n 0.0213448f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_550 N_RESET_B_M1027_g N_A_1790_74#_c_1504_n 0.0184362f $X=10.715 $Y=0.58
+ $X2=0 $Y2=0
cc_551 N_RESET_B_c_549_n N_A_1790_74#_c_1504_n 0.00370089f $X=10.855 $Y=1.55
+ $X2=0 $Y2=0
cc_552 N_RESET_B_c_557_n N_VPWR_M1022_d 0.00289772f $X=7.775 $Y=2.035 $X2=0
+ $Y2=0
cc_553 N_RESET_B_c_559_n N_VPWR_M1011_s 0.00198285f $X=10.655 $Y=2.035 $X2=0
+ $Y2=0
cc_554 N_RESET_B_c_551_n N_VPWR_c_1697_n 0.00579128f $X=3.605 $Y=2.245 $X2=0
+ $Y2=0
cc_555 N_RESET_B_c_552_n N_VPWR_c_1699_n 0.00314968f $X=7.525 $Y=2.21 $X2=0
+ $Y2=0
cc_556 N_RESET_B_c_552_n N_VPWR_c_1700_n 0.00490213f $X=7.525 $Y=2.21 $X2=0
+ $Y2=0
cc_557 N_RESET_B_c_547_n N_VPWR_c_1700_n 4.78591e-19 $X=7.735 $Y=1.795 $X2=0
+ $Y2=0
cc_558 N_RESET_B_c_559_n N_VPWR_c_1700_n 0.0236795f $X=10.655 $Y=2.035 $X2=0
+ $Y2=0
cc_559 N_RESET_B_c_560_n N_VPWR_c_1700_n 0.0027362f $X=8.065 $Y=2.035 $X2=0
+ $Y2=0
cc_560 N_RESET_B_c_564_n N_VPWR_c_1700_n 0.0020516f $X=7.735 $Y=2.002 $X2=0
+ $Y2=0
cc_561 N_RESET_B_c_565_n N_VPWR_c_1700_n 0.0258087f $X=7.825 $Y=1.96 $X2=0 $Y2=0
cc_562 N_RESET_B_c_566_n N_VPWR_c_1702_n 0.0233946f $X=10.8 $Y=2.035 $X2=0 $Y2=0
cc_563 N_RESET_B_c_551_n N_VPWR_c_1707_n 0.00388952f $X=3.605 $Y=2.245 $X2=0
+ $Y2=0
cc_564 N_RESET_B_c_555_n N_VPWR_c_1713_n 0.00443738f $X=11.005 $Y=2.28 $X2=0
+ $Y2=0
cc_565 N_RESET_B_c_555_n N_VPWR_c_1721_n 0.00802674f $X=11.005 $Y=2.28 $X2=0
+ $Y2=0
cc_566 N_RESET_B_c_559_n N_VPWR_c_1721_n 0.00135379f $X=10.655 $Y=2.035 $X2=0
+ $Y2=0
cc_567 N_RESET_B_c_551_n N_VPWR_c_1696_n 0.0042369f $X=3.605 $Y=2.245 $X2=0
+ $Y2=0
cc_568 N_RESET_B_c_552_n N_VPWR_c_1696_n 9.49986e-19 $X=7.525 $Y=2.21 $X2=0
+ $Y2=0
cc_569 N_RESET_B_c_555_n N_VPWR_c_1696_n 0.00489211f $X=11.005 $Y=2.28 $X2=0
+ $Y2=0
cc_570 N_RESET_B_M1043_g N_A_388_79#_c_1880_n 0.0166505f $X=3.59 $Y=0.605 $X2=0
+ $Y2=0
cc_571 N_RESET_B_M1043_g N_A_388_79#_c_1882_n 0.0227291f $X=3.59 $Y=0.605 $X2=0
+ $Y2=0
cc_572 N_RESET_B_c_551_n N_A_388_79#_c_1882_n 0.00392187f $X=3.605 $Y=2.245
+ $X2=0 $Y2=0
cc_573 N_RESET_B_c_558_n N_A_388_79#_c_1882_n 0.00108246f $X=4.225 $Y=2.035
+ $X2=0 $Y2=0
cc_574 N_RESET_B_c_562_n N_A_388_79#_c_1882_n 0.0144658f $X=3.605 $Y=2.032 $X2=0
+ $Y2=0
cc_575 N_RESET_B_c_563_n N_A_388_79#_c_1882_n 0.0228178f $X=3.95 $Y=1.985 $X2=0
+ $Y2=0
cc_576 N_RESET_B_c_551_n N_A_388_79#_c_1890_n 0.010753f $X=3.605 $Y=2.245 $X2=0
+ $Y2=0
cc_577 N_RESET_B_c_557_n N_A_388_79#_c_1891_n 0.0300096f $X=7.775 $Y=2.035 $X2=0
+ $Y2=0
cc_578 N_RESET_B_c_558_n N_A_388_79#_c_1891_n 0.00691285f $X=4.225 $Y=2.035
+ $X2=0 $Y2=0
cc_579 N_RESET_B_c_562_n N_A_388_79#_c_1891_n 0.00197315f $X=3.605 $Y=2.032
+ $X2=0 $Y2=0
cc_580 N_RESET_B_c_563_n N_A_388_79#_c_1891_n 0.00917413f $X=3.95 $Y=1.985 $X2=0
+ $Y2=0
cc_581 N_RESET_B_c_551_n N_A_388_79#_c_1892_n 0.0144438f $X=3.605 $Y=2.245 $X2=0
+ $Y2=0
cc_582 N_RESET_B_c_558_n N_A_388_79#_c_1892_n 0.001474f $X=4.225 $Y=2.035 $X2=0
+ $Y2=0
cc_583 N_RESET_B_c_562_n N_A_388_79#_c_1892_n 0.00751654f $X=3.605 $Y=2.032
+ $X2=0 $Y2=0
cc_584 N_RESET_B_c_563_n N_A_388_79#_c_1892_n 0.0165337f $X=3.95 $Y=1.985 $X2=0
+ $Y2=0
cc_585 N_RESET_B_c_557_n N_A_388_79#_c_1893_n 0.0218218f $X=7.775 $Y=2.035 $X2=0
+ $Y2=0
cc_586 N_RESET_B_c_557_n N_A_388_79#_c_1894_n 0.0125501f $X=7.775 $Y=2.035 $X2=0
+ $Y2=0
cc_587 N_RESET_B_c_557_n N_A_388_79#_c_1886_n 0.00638354f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_588 N_RESET_B_M1043_g N_VGND_c_2085_n 0.0117931f $X=3.59 $Y=0.605 $X2=0 $Y2=0
cc_589 N_RESET_B_M1027_g N_VGND_c_2087_n 0.0122664f $X=10.715 $Y=0.58 $X2=0
+ $Y2=0
cc_590 N_RESET_B_M1043_g N_VGND_c_2094_n 0.00465077f $X=3.59 $Y=0.605 $X2=0
+ $Y2=0
cc_591 N_RESET_B_M1027_g N_VGND_c_2101_n 0.00383152f $X=10.715 $Y=0.58 $X2=0
+ $Y2=0
cc_592 N_RESET_B_c_544_n N_VGND_c_2105_n 0.0033127f $X=7.32 $Y=1.085 $X2=0 $Y2=0
cc_593 N_RESET_B_M1043_g N_VGND_c_2110_n 0.00451796f $X=3.59 $Y=0.605 $X2=0
+ $Y2=0
cc_594 N_RESET_B_c_544_n N_VGND_c_2110_n 0.00479212f $X=7.32 $Y=1.085 $X2=0
+ $Y2=0
cc_595 N_RESET_B_M1027_g N_VGND_c_2110_n 0.0075694f $X=10.715 $Y=0.58 $X2=0
+ $Y2=0
cc_596 N_RESET_B_M1043_g N_noxref_25_c_2242_n 0.00154841f $X=3.59 $Y=0.605 $X2=0
+ $Y2=0
cc_597 N_RESET_B_M1043_g N_noxref_25_c_2244_n 0.00366715f $X=3.59 $Y=0.605 $X2=0
+ $Y2=0
cc_598 N_CLK_c_734_n N_A_1025_74#_c_794_n 6.63932e-19 $X=4.645 $Y=1.765 $X2=0
+ $Y2=0
cc_599 N_CLK_c_733_n N_A_852_74#_M1006_g 0.0113419f $X=4.62 $Y=1.22 $X2=0 $Y2=0
cc_600 N_CLK_c_734_n N_A_852_74#_M1006_g 0.024458f $X=4.645 $Y=1.765 $X2=0 $Y2=0
cc_601 N_CLK_c_734_n N_A_852_74#_c_1191_n 0.0446523f $X=4.645 $Y=1.765 $X2=0
+ $Y2=0
cc_602 N_CLK_c_733_n N_A_852_74#_c_1200_n 0.00627309f $X=4.62 $Y=1.22 $X2=0
+ $Y2=0
cc_603 N_CLK_c_733_n N_A_852_74#_c_1201_n 0.00467636f $X=4.62 $Y=1.22 $X2=0
+ $Y2=0
cc_604 N_CLK_c_734_n N_A_852_74#_c_1201_n 0.00193272f $X=4.645 $Y=1.765 $X2=0
+ $Y2=0
cc_605 N_CLK_c_735_n N_A_852_74#_c_1201_n 0.00630475f $X=4.545 $Y=1.385 $X2=0
+ $Y2=0
cc_606 CLK N_A_852_74#_c_1201_n 0.0109927f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_607 N_CLK_c_734_n N_A_852_74#_c_1232_n 8.07216e-19 $X=4.645 $Y=1.765 $X2=0
+ $Y2=0
cc_608 N_CLK_c_735_n N_A_852_74#_c_1232_n 0.00607893f $X=4.545 $Y=1.385 $X2=0
+ $Y2=0
cc_609 CLK N_A_852_74#_c_1232_n 0.0135702f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_610 N_CLK_c_734_n N_A_852_74#_c_1220_n 0.0091772f $X=4.645 $Y=1.765 $X2=0
+ $Y2=0
cc_611 N_CLK_c_734_n N_A_852_74#_c_1202_n 0.00367016f $X=4.645 $Y=1.765 $X2=0
+ $Y2=0
cc_612 N_CLK_c_733_n N_A_852_74#_c_1203_n 0.00175584f $X=4.62 $Y=1.22 $X2=0
+ $Y2=0
cc_613 N_CLK_c_735_n N_A_852_74#_c_1203_n 0.00690635f $X=4.545 $Y=1.385 $X2=0
+ $Y2=0
cc_614 N_CLK_c_734_n N_A_852_74#_c_1222_n 0.00460814f $X=4.645 $Y=1.765 $X2=0
+ $Y2=0
cc_615 N_CLK_c_735_n N_A_852_74#_c_1222_n 0.00585219f $X=4.545 $Y=1.385 $X2=0
+ $Y2=0
cc_616 N_CLK_c_734_n N_A_852_74#_c_1204_n 0.01381f $X=4.645 $Y=1.765 $X2=0 $Y2=0
cc_617 N_CLK_c_734_n N_A_852_74#_c_1205_n 0.00379234f $X=4.645 $Y=1.765 $X2=0
+ $Y2=0
cc_618 CLK N_A_852_74#_c_1205_n 0.0016136f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_619 N_CLK_c_734_n N_VPWR_c_1698_n 0.0189827f $X=4.645 $Y=1.765 $X2=0 $Y2=0
cc_620 N_CLK_c_734_n N_VPWR_c_1707_n 0.00413917f $X=4.645 $Y=1.765 $X2=0 $Y2=0
cc_621 N_CLK_c_734_n N_VPWR_c_1696_n 0.00412518f $X=4.645 $Y=1.765 $X2=0 $Y2=0
cc_622 N_CLK_c_735_n N_A_388_79#_c_1882_n 0.00130698f $X=4.545 $Y=1.385 $X2=0
+ $Y2=0
cc_623 CLK N_A_388_79#_c_1882_n 0.0174093f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_624 N_CLK_c_734_n N_A_388_79#_c_1890_n 0.0113821f $X=4.645 $Y=1.765 $X2=0
+ $Y2=0
cc_625 N_CLK_c_734_n N_A_388_79#_c_1891_n 0.0145615f $X=4.645 $Y=1.765 $X2=0
+ $Y2=0
cc_626 N_CLK_c_734_n N_A_388_79#_c_1892_n 8.09031e-19 $X=4.645 $Y=1.765 $X2=0
+ $Y2=0
cc_627 N_CLK_c_733_n N_VGND_c_2085_n 0.00361986f $X=4.62 $Y=1.22 $X2=0 $Y2=0
cc_628 N_CLK_c_735_n N_VGND_c_2085_n 4.22243e-19 $X=4.545 $Y=1.385 $X2=0 $Y2=0
cc_629 CLK N_VGND_c_2085_n 0.00344374f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_630 N_CLK_c_733_n N_VGND_c_2086_n 0.0031368f $X=4.62 $Y=1.22 $X2=0 $Y2=0
cc_631 N_CLK_c_733_n N_VGND_c_2096_n 0.00428607f $X=4.62 $Y=1.22 $X2=0 $Y2=0
cc_632 N_CLK_c_733_n N_VGND_c_2110_n 0.00807037f $X=4.62 $Y=1.22 $X2=0 $Y2=0
cc_633 N_A_1025_74#_c_797_n N_A_1370_289#_M1003_d 0.00176891f $X=9.1 $Y=0.34
+ $X2=-0.19 $Y2=-0.245
cc_634 N_A_1025_74#_c_806_n N_A_1370_289#_c_995_n 0.00189178f $X=6.1 $Y=2.12
+ $X2=0 $Y2=0
cc_635 N_A_1025_74#_M1020_g N_A_1370_289#_M1001_g 0.0462918f $X=6.54 $Y=0.8
+ $X2=0 $Y2=0
cc_636 N_A_1025_74#_c_791_n N_A_1370_289#_M1001_g 0.00943625f $X=7 $Y=0.395
+ $X2=0 $Y2=0
cc_637 N_A_1025_74#_c_801_n N_A_1370_289#_M1001_g 0.00547119f $X=7.085 $Y=0.395
+ $X2=0 $Y2=0
cc_638 N_A_1025_74#_c_807_n N_A_1370_289#_c_996_n 0.00189178f $X=6.1 $Y=2.21
+ $X2=0 $Y2=0
cc_639 N_A_1025_74#_M1020_g N_A_1370_289#_c_991_n 0.0107798f $X=6.54 $Y=0.8
+ $X2=0 $Y2=0
cc_640 N_A_1025_74#_c_801_n N_A_1370_289#_c_991_n 3.86554e-19 $X=7.085 $Y=0.395
+ $X2=0 $Y2=0
cc_641 N_A_1025_74#_c_805_n N_A_1370_289#_c_991_n 0.00192454f $X=6.045 $Y=1.575
+ $X2=0 $Y2=0
cc_642 N_A_1025_74#_c_796_n N_A_1370_289#_c_1027_n 0.00146445f $X=8.155 $Y=0.665
+ $X2=0 $Y2=0
cc_643 N_A_1025_74#_c_801_n N_A_1370_289#_c_1027_n 0.00967347f $X=7.085 $Y=0.395
+ $X2=0 $Y2=0
cc_644 N_A_1025_74#_c_808_n N_A_1370_289#_c_1029_n 3.85264e-19 $X=9.7 $Y=2.28
+ $X2=0 $Y2=0
cc_645 N_A_1025_74#_c_811_n N_A_1370_289#_c_1029_n 0.0194918f $X=9.615 $Y=2.03
+ $X2=0 $Y2=0
cc_646 N_A_1025_74#_c_808_n N_A_1370_289#_c_999_n 0.00120571f $X=9.7 $Y=2.28
+ $X2=0 $Y2=0
cc_647 N_A_1025_74#_c_796_n N_A_1370_289#_c_992_n 0.0737203f $X=8.155 $Y=0.665
+ $X2=0 $Y2=0
cc_648 N_A_1025_74#_c_797_n N_A_1370_289#_c_992_n 0.00353238f $X=9.1 $Y=0.34
+ $X2=0 $Y2=0
cc_649 N_A_1025_74#_c_787_n N_A_1370_289#_c_993_n 0.0114651f $X=8.875 $Y=1.085
+ $X2=0 $Y2=0
cc_650 N_A_1025_74#_c_789_n N_A_1370_289#_c_993_n 4.45722e-19 $X=8.95 $Y=1.16
+ $X2=0 $Y2=0
cc_651 N_A_1025_74#_c_797_n N_A_1370_289#_c_993_n 0.0229775f $X=9.1 $Y=0.34
+ $X2=0 $Y2=0
cc_652 N_A_1025_74#_c_799_n N_A_1370_289#_c_993_n 0.0234316f $X=9.185 $Y=0.905
+ $X2=0 $Y2=0
cc_653 N_A_1025_74#_c_802_n N_A_1370_289#_c_993_n 0.0157507f $X=9.475 $Y=1.07
+ $X2=0 $Y2=0
cc_654 N_A_1025_74#_c_789_n N_A_1370_289#_c_994_n 0.006971f $X=8.95 $Y=1.16
+ $X2=0 $Y2=0
cc_655 N_A_1025_74#_c_802_n N_A_1370_289#_c_994_n 0.0107601f $X=9.475 $Y=1.07
+ $X2=0 $Y2=0
cc_656 N_A_1025_74#_c_804_n N_A_1370_289#_c_994_n 0.0194918f $X=9.532 $Y=1.865
+ $X2=0 $Y2=0
cc_657 N_A_1025_74#_c_787_n N_A_1223_118#_M1003_g 0.0264029f $X=8.875 $Y=1.085
+ $X2=0 $Y2=0
cc_658 N_A_1025_74#_c_797_n N_A_1223_118#_M1003_g 0.0116384f $X=9.1 $Y=0.34
+ $X2=0 $Y2=0
cc_659 N_A_1025_74#_c_785_n N_A_1223_118#_c_1119_n 6.10614e-19 $X=6.465 $Y=1.575
+ $X2=0 $Y2=0
cc_660 N_A_1025_74#_M1020_g N_A_1223_118#_c_1119_n 0.0148322f $X=6.54 $Y=0.8
+ $X2=0 $Y2=0
cc_661 N_A_1025_74#_c_791_n N_A_1223_118#_c_1119_n 0.0431682f $X=7 $Y=0.395
+ $X2=0 $Y2=0
cc_662 N_A_1025_74#_c_806_n N_A_1223_118#_c_1088_n 4.7499e-19 $X=6.1 $Y=2.12
+ $X2=0 $Y2=0
cc_663 N_A_1025_74#_M1020_g N_A_1223_118#_c_1088_n 0.00532373f $X=6.54 $Y=0.8
+ $X2=0 $Y2=0
cc_664 N_A_1025_74#_c_807_n N_A_1223_118#_c_1094_n 0.00437093f $X=6.1 $Y=2.21
+ $X2=0 $Y2=0
cc_665 N_A_1025_74#_c_785_n N_A_1223_118#_c_1094_n 0.0010957f $X=6.465 $Y=1.575
+ $X2=0 $Y2=0
cc_666 N_A_1025_74#_c_790_n N_A_852_74#_M1006_g 0.00654973f $X=5.265 $Y=0.515
+ $X2=0 $Y2=0
cc_667 N_A_1025_74#_c_792_n N_A_852_74#_M1006_g 0.00338004f $X=5.43 $Y=0.395
+ $X2=0 $Y2=0
cc_668 N_A_1025_74#_c_793_n N_A_852_74#_M1006_g 0.0029449f $X=5.56 $Y=1.5 $X2=0
+ $Y2=0
cc_669 N_A_1025_74#_c_800_n N_A_852_74#_M1006_g 0.00307434f $X=5.56 $Y=1.075
+ $X2=0 $Y2=0
cc_670 N_A_1025_74#_c_794_n N_A_852_74#_c_1191_n 0.00991617f $X=5.645 $Y=1.665
+ $X2=0 $Y2=0
cc_671 N_A_1025_74#_c_800_n N_A_852_74#_c_1191_n 0.00428164f $X=5.56 $Y=1.075
+ $X2=0 $Y2=0
cc_672 N_A_1025_74#_c_793_n N_A_852_74#_c_1192_n 0.00252518f $X=5.56 $Y=1.5
+ $X2=0 $Y2=0
cc_673 N_A_1025_74#_c_794_n N_A_852_74#_c_1192_n 0.00383968f $X=5.645 $Y=1.665
+ $X2=0 $Y2=0
cc_674 N_A_1025_74#_c_806_n N_A_852_74#_c_1193_n 0.0129259f $X=6.1 $Y=2.12 $X2=0
+ $Y2=0
cc_675 N_A_1025_74#_c_807_n N_A_852_74#_c_1193_n 0.0132885f $X=6.1 $Y=2.21 $X2=0
+ $Y2=0
cc_676 N_A_1025_74#_c_793_n N_A_852_74#_c_1193_n 5.77257e-19 $X=5.56 $Y=1.5
+ $X2=0 $Y2=0
cc_677 N_A_1025_74#_c_794_n N_A_852_74#_c_1193_n 0.0186066f $X=5.645 $Y=1.665
+ $X2=0 $Y2=0
cc_678 N_A_1025_74#_c_795_n N_A_852_74#_c_1193_n 0.00529731f $X=6.045 $Y=1.665
+ $X2=0 $Y2=0
cc_679 N_A_1025_74#_c_805_n N_A_852_74#_c_1193_n 0.0213786f $X=6.045 $Y=1.575
+ $X2=0 $Y2=0
cc_680 N_A_1025_74#_c_795_n N_A_852_74#_c_1194_n 0.00583367f $X=6.045 $Y=1.665
+ $X2=0 $Y2=0
cc_681 N_A_1025_74#_c_805_n N_A_852_74#_c_1194_n 0.0127944f $X=6.045 $Y=1.575
+ $X2=0 $Y2=0
cc_682 N_A_1025_74#_c_807_n N_A_852_74#_c_1208_n 0.00899632f $X=6.1 $Y=2.21
+ $X2=0 $Y2=0
cc_683 N_A_1025_74#_M1020_g N_A_852_74#_c_1195_n 0.0200223f $X=6.54 $Y=0.8 $X2=0
+ $Y2=0
cc_684 N_A_1025_74#_c_790_n N_A_852_74#_c_1195_n 0.00422225f $X=5.265 $Y=0.515
+ $X2=0 $Y2=0
cc_685 N_A_1025_74#_c_791_n N_A_852_74#_c_1195_n 0.00744742f $X=7 $Y=0.395 $X2=0
+ $Y2=0
cc_686 N_A_1025_74#_c_800_n N_A_852_74#_c_1195_n 6.53033e-19 $X=5.56 $Y=1.075
+ $X2=0 $Y2=0
cc_687 N_A_1025_74#_c_807_n N_A_852_74#_c_1210_n 0.00278823f $X=6.1 $Y=2.21
+ $X2=0 $Y2=0
cc_688 N_A_1025_74#_c_807_n N_A_852_74#_c_1212_n 0.0105241f $X=6.1 $Y=2.21 $X2=0
+ $Y2=0
cc_689 N_A_1025_74#_c_785_n N_A_852_74#_c_1212_n 0.00365124f $X=6.465 $Y=1.575
+ $X2=0 $Y2=0
cc_690 N_A_1025_74#_c_808_n N_A_852_74#_c_1214_n 0.00247489f $X=9.7 $Y=2.28
+ $X2=0 $Y2=0
cc_691 N_A_1025_74#_c_808_n N_A_852_74#_M1016_g 0.0185475f $X=9.7 $Y=2.28 $X2=0
+ $Y2=0
cc_692 N_A_1025_74#_c_804_n N_A_852_74#_M1016_g 0.00632245f $X=9.532 $Y=1.865
+ $X2=0 $Y2=0
cc_693 N_A_1025_74#_c_788_n N_A_852_74#_c_1196_n 0.0218467f $X=9.31 $Y=1.16
+ $X2=0 $Y2=0
cc_694 N_A_1025_74#_c_808_n N_A_852_74#_c_1196_n 0.0184752f $X=9.7 $Y=2.28 $X2=0
+ $Y2=0
cc_695 N_A_1025_74#_c_802_n N_A_852_74#_c_1196_n 0.00157771f $X=9.475 $Y=1.07
+ $X2=0 $Y2=0
cc_696 N_A_1025_74#_c_811_n N_A_852_74#_c_1196_n 7.40372e-19 $X=9.615 $Y=2.03
+ $X2=0 $Y2=0
cc_697 N_A_1025_74#_c_804_n N_A_852_74#_c_1196_n 0.0190498f $X=9.532 $Y=1.865
+ $X2=0 $Y2=0
cc_698 N_A_1025_74#_c_789_n N_A_852_74#_c_1197_n 0.0218467f $X=8.95 $Y=1.16
+ $X2=0 $Y2=0
cc_699 N_A_1025_74#_c_804_n N_A_852_74#_c_1197_n 7.05953e-19 $X=9.532 $Y=1.865
+ $X2=0 $Y2=0
cc_700 N_A_1025_74#_c_797_n N_A_852_74#_M1002_g 0.00370958f $X=9.1 $Y=0.34 $X2=0
+ $Y2=0
cc_701 N_A_1025_74#_c_799_n N_A_852_74#_M1002_g 0.00214927f $X=9.185 $Y=0.905
+ $X2=0 $Y2=0
cc_702 N_A_1025_74#_c_802_n N_A_852_74#_M1002_g 0.00105258f $X=9.475 $Y=1.07
+ $X2=0 $Y2=0
cc_703 N_A_1025_74#_c_803_n N_A_852_74#_M1002_g 0.0196932f $X=9.475 $Y=1.07
+ $X2=0 $Y2=0
cc_704 N_A_1025_74#_c_804_n N_A_852_74#_M1002_g 0.00477388f $X=9.532 $Y=1.865
+ $X2=0 $Y2=0
cc_705 N_A_1025_74#_c_791_n N_A_852_74#_c_1199_n 0.00122664f $X=7 $Y=0.395 $X2=0
+ $Y2=0
cc_706 N_A_1025_74#_c_793_n N_A_852_74#_c_1199_n 0.0125452f $X=5.56 $Y=1.5 $X2=0
+ $Y2=0
cc_707 N_A_1025_74#_c_800_n N_A_852_74#_c_1199_n 0.00520589f $X=5.56 $Y=1.075
+ $X2=0 $Y2=0
cc_708 N_A_1025_74#_c_800_n N_A_852_74#_c_1201_n 8.59093e-19 $X=5.56 $Y=1.075
+ $X2=0 $Y2=0
cc_709 N_A_1025_74#_c_794_n N_A_852_74#_c_1220_n 0.00754252f $X=5.645 $Y=1.665
+ $X2=0 $Y2=0
cc_710 N_A_1025_74#_c_794_n N_A_852_74#_c_1202_n 0.00641585f $X=5.645 $Y=1.665
+ $X2=0 $Y2=0
cc_711 N_A_1025_74#_c_794_n N_A_852_74#_c_1222_n 0.00293499f $X=5.645 $Y=1.665
+ $X2=0 $Y2=0
cc_712 N_A_1025_74#_c_793_n N_A_852_74#_c_1205_n 0.0129106f $X=5.56 $Y=1.5 $X2=0
+ $Y2=0
cc_713 N_A_1025_74#_c_794_n N_A_852_74#_c_1205_n 0.024952f $X=5.645 $Y=1.665
+ $X2=0 $Y2=0
cc_714 N_A_1025_74#_c_800_n N_A_852_74#_c_1205_n 0.015315f $X=5.56 $Y=1.075
+ $X2=0 $Y2=0
cc_715 N_A_1025_74#_c_808_n N_A_2006_373#_c_1391_n 0.0292474f $X=9.7 $Y=2.28
+ $X2=0 $Y2=0
cc_716 N_A_1025_74#_c_808_n N_A_2006_373#_c_1398_n 0.0224077f $X=9.7 $Y=2.28
+ $X2=0 $Y2=0
cc_717 N_A_1025_74#_c_811_n N_A_2006_373#_c_1398_n 3.95315e-19 $X=9.615 $Y=2.03
+ $X2=0 $Y2=0
cc_718 N_A_1025_74#_c_797_n N_A_1790_74#_M1024_d 0.00293623f $X=9.1 $Y=0.34
+ $X2=-0.19 $Y2=-0.245
cc_719 N_A_1025_74#_c_799_n N_A_1790_74#_M1024_d 0.0113447f $X=9.185 $Y=0.905
+ $X2=-0.19 $Y2=-0.245
cc_720 N_A_1025_74#_c_802_n N_A_1790_74#_M1024_d 0.00118465f $X=9.475 $Y=1.07
+ $X2=-0.19 $Y2=-0.245
cc_721 N_A_1025_74#_c_808_n N_A_1790_74#_c_1522_n 0.0204256f $X=9.7 $Y=2.28
+ $X2=0 $Y2=0
cc_722 N_A_1025_74#_c_811_n N_A_1790_74#_c_1522_n 0.0316971f $X=9.615 $Y=2.03
+ $X2=0 $Y2=0
cc_723 N_A_1025_74#_c_787_n N_A_1790_74#_c_1531_n 5.95394e-19 $X=8.875 $Y=1.085
+ $X2=0 $Y2=0
cc_724 N_A_1025_74#_c_797_n N_A_1790_74#_c_1531_n 0.00170833f $X=9.1 $Y=0.34
+ $X2=0 $Y2=0
cc_725 N_A_1025_74#_c_799_n N_A_1790_74#_c_1531_n 0.0250265f $X=9.185 $Y=0.905
+ $X2=0 $Y2=0
cc_726 N_A_1025_74#_c_802_n N_A_1790_74#_c_1531_n 0.0155252f $X=9.475 $Y=1.07
+ $X2=0 $Y2=0
cc_727 N_A_1025_74#_c_803_n N_A_1790_74#_c_1531_n 0.00455646f $X=9.475 $Y=1.07
+ $X2=0 $Y2=0
cc_728 N_A_1025_74#_c_799_n N_A_1790_74#_c_1502_n 0.00427034f $X=9.185 $Y=0.905
+ $X2=0 $Y2=0
cc_729 N_A_1025_74#_c_802_n N_A_1790_74#_c_1502_n 0.00683662f $X=9.475 $Y=1.07
+ $X2=0 $Y2=0
cc_730 N_A_1025_74#_c_808_n N_A_1790_74#_c_1503_n 0.00539734f $X=9.7 $Y=2.28
+ $X2=0 $Y2=0
cc_731 N_A_1025_74#_c_811_n N_A_1790_74#_c_1503_n 0.0241297f $X=9.615 $Y=2.03
+ $X2=0 $Y2=0
cc_732 N_A_1025_74#_c_804_n N_A_1790_74#_c_1503_n 0.0288004f $X=9.532 $Y=1.865
+ $X2=0 $Y2=0
cc_733 N_A_1025_74#_c_802_n N_A_1790_74#_c_1541_n 0.0103633f $X=9.475 $Y=1.07
+ $X2=0 $Y2=0
cc_734 N_A_1025_74#_c_803_n N_A_1790_74#_c_1541_n 2.09861e-19 $X=9.475 $Y=1.07
+ $X2=0 $Y2=0
cc_735 N_A_1025_74#_c_804_n N_A_1790_74#_c_1541_n 0.00427046f $X=9.532 $Y=1.865
+ $X2=0 $Y2=0
cc_736 N_A_1025_74#_c_808_n N_VPWR_c_1701_n 0.00349642f $X=9.7 $Y=2.28 $X2=0
+ $Y2=0
cc_737 N_A_1025_74#_c_807_n N_VPWR_c_1696_n 9.49986e-19 $X=6.1 $Y=2.21 $X2=0
+ $Y2=0
cc_738 N_A_1025_74#_c_808_n N_VPWR_c_1696_n 0.00489211f $X=9.7 $Y=2.28 $X2=0
+ $Y2=0
cc_739 N_A_1025_74#_M1032_d N_A_388_79#_c_1891_n 0.00646182f $X=5.17 $Y=1.84
+ $X2=0 $Y2=0
cc_740 N_A_1025_74#_c_794_n N_A_388_79#_c_1891_n 0.0279831f $X=5.645 $Y=1.665
+ $X2=0 $Y2=0
cc_741 N_A_1025_74#_c_795_n N_A_388_79#_c_1891_n 0.00271336f $X=6.045 $Y=1.665
+ $X2=0 $Y2=0
cc_742 N_A_1025_74#_M1020_g N_A_388_79#_c_1883_n 4.31453e-19 $X=6.54 $Y=0.8
+ $X2=0 $Y2=0
cc_743 N_A_1025_74#_c_790_n N_A_388_79#_c_1883_n 0.00733866f $X=5.265 $Y=0.515
+ $X2=0 $Y2=0
cc_744 N_A_1025_74#_c_800_n N_A_388_79#_c_1883_n 0.010339f $X=5.56 $Y=1.075
+ $X2=0 $Y2=0
cc_745 N_A_1025_74#_c_806_n N_A_388_79#_c_1893_n 0.00707608f $X=6.1 $Y=2.12
+ $X2=0 $Y2=0
cc_746 N_A_1025_74#_c_807_n N_A_388_79#_c_1893_n 0.00869011f $X=6.1 $Y=2.21
+ $X2=0 $Y2=0
cc_747 N_A_1025_74#_c_785_n N_A_388_79#_c_1893_n 0.00260393f $X=6.465 $Y=1.575
+ $X2=0 $Y2=0
cc_748 N_A_1025_74#_c_795_n N_A_388_79#_c_1893_n 0.0103323f $X=6.045 $Y=1.665
+ $X2=0 $Y2=0
cc_749 N_A_1025_74#_c_805_n N_A_388_79#_c_1893_n 0.00122453f $X=6.045 $Y=1.575
+ $X2=0 $Y2=0
cc_750 N_A_1025_74#_c_794_n N_A_388_79#_c_1894_n 0.0121841f $X=5.645 $Y=1.665
+ $X2=0 $Y2=0
cc_751 N_A_1025_74#_c_795_n N_A_388_79#_c_1894_n 0.0116438f $X=6.045 $Y=1.665
+ $X2=0 $Y2=0
cc_752 N_A_1025_74#_c_805_n N_A_388_79#_c_1894_n 0.00234227f $X=6.045 $Y=1.575
+ $X2=0 $Y2=0
cc_753 N_A_1025_74#_M1020_g N_A_388_79#_c_1884_n 0.00474699f $X=6.54 $Y=0.8
+ $X2=0 $Y2=0
cc_754 N_A_1025_74#_c_791_n N_A_388_79#_c_1884_n 0.00414539f $X=7 $Y=0.395 $X2=0
+ $Y2=0
cc_755 N_A_1025_74#_c_795_n N_A_388_79#_c_1884_n 0.0102296f $X=6.045 $Y=1.665
+ $X2=0 $Y2=0
cc_756 N_A_1025_74#_c_805_n N_A_388_79#_c_1884_n 0.00755283f $X=6.045 $Y=1.575
+ $X2=0 $Y2=0
cc_757 N_A_1025_74#_c_793_n N_A_388_79#_c_1885_n 0.009798f $X=5.56 $Y=1.5 $X2=0
+ $Y2=0
cc_758 N_A_1025_74#_c_795_n N_A_388_79#_c_1885_n 0.0121259f $X=6.045 $Y=1.665
+ $X2=0 $Y2=0
cc_759 N_A_1025_74#_c_800_n N_A_388_79#_c_1885_n 0.00316754f $X=5.56 $Y=1.075
+ $X2=0 $Y2=0
cc_760 N_A_1025_74#_c_805_n N_A_388_79#_c_1885_n 6.96658e-19 $X=6.045 $Y=1.575
+ $X2=0 $Y2=0
cc_761 N_A_1025_74#_c_806_n N_A_388_79#_c_1886_n 0.00249482f $X=6.1 $Y=2.12
+ $X2=0 $Y2=0
cc_762 N_A_1025_74#_c_785_n N_A_388_79#_c_1886_n 0.0122801f $X=6.465 $Y=1.575
+ $X2=0 $Y2=0
cc_763 N_A_1025_74#_M1020_g N_A_388_79#_c_1886_n 0.00569046f $X=6.54 $Y=0.8
+ $X2=0 $Y2=0
cc_764 N_A_1025_74#_c_793_n N_A_388_79#_c_1886_n 0.00522407f $X=5.56 $Y=1.5
+ $X2=0 $Y2=0
cc_765 N_A_1025_74#_c_794_n N_A_388_79#_c_1886_n 0.00398889f $X=5.645 $Y=1.665
+ $X2=0 $Y2=0
cc_766 N_A_1025_74#_c_795_n N_A_388_79#_c_1886_n 0.0256385f $X=6.045 $Y=1.665
+ $X2=0 $Y2=0
cc_767 N_A_1025_74#_c_805_n N_A_388_79#_c_1886_n 0.00206889f $X=6.045 $Y=1.575
+ $X2=0 $Y2=0
cc_768 N_A_1025_74#_c_790_n N_A_388_79#_c_1887_n 0.0113657f $X=5.265 $Y=0.515
+ $X2=0 $Y2=0
cc_769 N_A_1025_74#_c_791_n N_A_388_79#_c_1887_n 0.0212058f $X=7 $Y=0.395 $X2=0
+ $Y2=0
cc_770 N_A_1025_74#_c_807_n N_A_388_79#_c_1896_n 0.0020657f $X=6.1 $Y=2.21 $X2=0
+ $Y2=0
cc_771 N_A_1025_74#_c_796_n N_VGND_M1012_d 0.0231403f $X=8.155 $Y=0.665 $X2=0
+ $Y2=0
cc_772 N_A_1025_74#_c_964_p N_VGND_M1012_d 0.00612573f $X=8.24 $Y=0.58 $X2=0
+ $Y2=0
cc_773 N_A_1025_74#_c_798_n N_VGND_M1012_d 0.0012599f $X=8.325 $Y=0.34 $X2=0
+ $Y2=0
cc_774 N_A_1025_74#_c_792_n N_VGND_c_2086_n 0.00897876f $X=5.43 $Y=0.395 $X2=0
+ $Y2=0
cc_775 N_A_1025_74#_c_800_n N_VGND_c_2086_n 0.0060955f $X=5.56 $Y=1.075 $X2=0
+ $Y2=0
cc_776 N_A_1025_74#_c_787_n N_VGND_c_2098_n 0.00278271f $X=8.875 $Y=1.085 $X2=0
+ $Y2=0
cc_777 N_A_1025_74#_c_796_n N_VGND_c_2098_n 0.003347f $X=8.155 $Y=0.665 $X2=0
+ $Y2=0
cc_778 N_A_1025_74#_c_797_n N_VGND_c_2098_n 0.0611382f $X=9.1 $Y=0.34 $X2=0
+ $Y2=0
cc_779 N_A_1025_74#_c_798_n N_VGND_c_2098_n 0.0118998f $X=8.325 $Y=0.34 $X2=0
+ $Y2=0
cc_780 N_A_1025_74#_M1020_g N_VGND_c_2105_n 6.21153e-19 $X=6.54 $Y=0.8 $X2=0
+ $Y2=0
cc_781 N_A_1025_74#_c_791_n N_VGND_c_2105_n 0.0752121f $X=7 $Y=0.395 $X2=0 $Y2=0
cc_782 N_A_1025_74#_c_792_n N_VGND_c_2105_n 0.0174472f $X=5.43 $Y=0.395 $X2=0
+ $Y2=0
cc_783 N_A_1025_74#_c_796_n N_VGND_c_2105_n 0.00545957f $X=8.155 $Y=0.665 $X2=0
+ $Y2=0
cc_784 N_A_1025_74#_c_801_n N_VGND_c_2105_n 0.00864403f $X=7.085 $Y=0.395 $X2=0
+ $Y2=0
cc_785 N_A_1025_74#_c_796_n N_VGND_c_2106_n 0.0398776f $X=8.155 $Y=0.665 $X2=0
+ $Y2=0
cc_786 N_A_1025_74#_c_798_n N_VGND_c_2106_n 0.014039f $X=8.325 $Y=0.34 $X2=0
+ $Y2=0
cc_787 N_A_1025_74#_c_801_n N_VGND_c_2106_n 0.00578724f $X=7.085 $Y=0.395 $X2=0
+ $Y2=0
cc_788 N_A_1025_74#_c_787_n N_VGND_c_2110_n 0.00358525f $X=8.875 $Y=1.085 $X2=0
+ $Y2=0
cc_789 N_A_1025_74#_c_791_n N_VGND_c_2110_n 0.0570267f $X=7 $Y=0.395 $X2=0 $Y2=0
cc_790 N_A_1025_74#_c_792_n N_VGND_c_2110_n 0.0123548f $X=5.43 $Y=0.395 $X2=0
+ $Y2=0
cc_791 N_A_1025_74#_c_796_n N_VGND_c_2110_n 0.0159235f $X=8.155 $Y=0.665 $X2=0
+ $Y2=0
cc_792 N_A_1025_74#_c_797_n N_VGND_c_2110_n 0.0343665f $X=9.1 $Y=0.34 $X2=0
+ $Y2=0
cc_793 N_A_1025_74#_c_798_n N_VGND_c_2110_n 0.00655543f $X=8.325 $Y=0.34 $X2=0
+ $Y2=0
cc_794 N_A_1025_74#_c_801_n N_VGND_c_2110_n 0.00626699f $X=7.085 $Y=0.395 $X2=0
+ $Y2=0
cc_795 N_A_1025_74#_c_796_n A_1401_118# 5.60007e-19 $X=8.155 $Y=0.665 $X2=-0.19
+ $Y2=-0.245
cc_796 N_A_1025_74#_c_801_n A_1401_118# 0.00146729f $X=7.085 $Y=0.395 $X2=-0.19
+ $Y2=-0.245
cc_797 N_A_1370_289#_c_992_n N_A_1223_118#_M1003_g 0.0106637f $X=8.495 $Y=0.842
+ $X2=0 $Y2=0
cc_798 N_A_1370_289#_c_993_n N_A_1223_118#_M1003_g 0.0115167f $X=8.845 $Y=0.842
+ $X2=0 $Y2=0
cc_799 N_A_1370_289#_c_994_n N_A_1223_118#_M1003_g 0.00305733f $X=8.785 $Y=1.745
+ $X2=0 $Y2=0
cc_800 N_A_1370_289#_c_1029_n N_A_1223_118#_c_1087_n 0.00358587f $X=8.785
+ $Y=1.89 $X2=0 $Y2=0
cc_801 N_A_1370_289#_c_992_n N_A_1223_118#_c_1087_n 0.00251001f $X=8.495
+ $Y=0.842 $X2=0 $Y2=0
cc_802 N_A_1370_289#_c_993_n N_A_1223_118#_c_1087_n 0.00187812f $X=8.845
+ $Y=0.842 $X2=0 $Y2=0
cc_803 N_A_1370_289#_c_994_n N_A_1223_118#_c_1087_n 0.00588778f $X=8.785
+ $Y=1.745 $X2=0 $Y2=0
cc_804 N_A_1370_289#_M1001_g N_A_1223_118#_c_1088_n 0.00321544f $X=6.93 $Y=0.8
+ $X2=0 $Y2=0
cc_805 N_A_1370_289#_c_996_n N_A_1223_118#_c_1088_n 0.00107886f $X=6.94 $Y=2.21
+ $X2=0 $Y2=0
cc_806 N_A_1370_289#_c_990_n N_A_1223_118#_c_1088_n 0.0496832f $X=7.105 $Y=1.61
+ $X2=0 $Y2=0
cc_807 N_A_1370_289#_c_991_n N_A_1223_118#_c_1088_n 0.0103879f $X=7.105 $Y=1.61
+ $X2=0 $Y2=0
cc_808 N_A_1370_289#_c_1027_n N_A_1223_118#_c_1088_n 0.00888203f $X=7.21
+ $Y=1.005 $X2=0 $Y2=0
cc_809 N_A_1370_289#_c_996_n N_A_1223_118#_c_1101_n 0.010858f $X=6.94 $Y=2.21
+ $X2=0 $Y2=0
cc_810 N_A_1370_289#_c_990_n N_A_1223_118#_c_1101_n 0.00225012f $X=7.105 $Y=1.61
+ $X2=0 $Y2=0
cc_811 N_A_1370_289#_c_991_n N_A_1223_118#_c_1101_n 0.00231625f $X=7.105 $Y=1.61
+ $X2=0 $Y2=0
cc_812 N_A_1370_289#_c_996_n N_A_1223_118#_c_1094_n 6.94181e-19 $X=6.94 $Y=2.21
+ $X2=0 $Y2=0
cc_813 N_A_1370_289#_c_995_n N_A_1223_118#_c_1089_n 0.00413444f $X=6.94 $Y=2.12
+ $X2=0 $Y2=0
cc_814 N_A_1370_289#_c_996_n N_A_1223_118#_c_1089_n 0.00183889f $X=6.94 $Y=2.21
+ $X2=0 $Y2=0
cc_815 N_A_1370_289#_c_990_n N_A_1223_118#_c_1089_n 0.01449f $X=7.105 $Y=1.61
+ $X2=0 $Y2=0
cc_816 N_A_1370_289#_c_991_n N_A_1223_118#_c_1089_n 0.00176149f $X=7.105 $Y=1.61
+ $X2=0 $Y2=0
cc_817 N_A_1370_289#_M1001_g N_A_1223_118#_c_1090_n 6.9585e-19 $X=6.93 $Y=0.8
+ $X2=0 $Y2=0
cc_818 N_A_1370_289#_c_990_n N_A_1223_118#_c_1090_n 0.0264869f $X=7.105 $Y=1.61
+ $X2=0 $Y2=0
cc_819 N_A_1370_289#_c_991_n N_A_1223_118#_c_1090_n 0.00127349f $X=7.105 $Y=1.61
+ $X2=0 $Y2=0
cc_820 N_A_1370_289#_c_992_n N_A_1223_118#_c_1090_n 0.0136798f $X=8.495 $Y=0.842
+ $X2=0 $Y2=0
cc_821 N_A_1370_289#_c_992_n N_A_1223_118#_c_1091_n 0.0791478f $X=8.495 $Y=0.842
+ $X2=0 $Y2=0
cc_822 N_A_1370_289#_c_994_n N_A_1223_118#_c_1091_n 0.0250137f $X=8.785 $Y=1.745
+ $X2=0 $Y2=0
cc_823 N_A_1370_289#_c_996_n N_A_852_74#_c_1210_n 0.00322542f $X=6.94 $Y=2.21
+ $X2=0 $Y2=0
cc_824 N_A_1370_289#_c_996_n N_A_852_74#_c_1212_n 0.0312132f $X=6.94 $Y=2.21
+ $X2=0 $Y2=0
cc_825 N_A_1370_289#_c_996_n N_A_852_74#_c_1213_n 0.00860132f $X=6.94 $Y=2.21
+ $X2=0 $Y2=0
cc_826 N_A_1370_289#_c_999_n N_A_852_74#_c_1213_n 0.00262042f $X=8.725 $Y=1.91
+ $X2=0 $Y2=0
cc_827 N_A_1370_289#_c_999_n N_A_852_74#_c_1214_n 5.08057e-19 $X=8.725 $Y=1.91
+ $X2=0 $Y2=0
cc_828 N_A_1370_289#_c_1029_n N_A_852_74#_M1016_g 0.00259852f $X=8.785 $Y=1.89
+ $X2=0 $Y2=0
cc_829 N_A_1370_289#_c_999_n N_A_852_74#_M1016_g 0.0157448f $X=8.725 $Y=1.91
+ $X2=0 $Y2=0
cc_830 N_A_1370_289#_c_994_n N_A_852_74#_M1016_g 0.00201426f $X=8.785 $Y=1.745
+ $X2=0 $Y2=0
cc_831 N_A_1370_289#_c_994_n N_A_852_74#_c_1197_n 0.00702349f $X=8.785 $Y=1.745
+ $X2=0 $Y2=0
cc_832 N_A_1370_289#_c_999_n N_A_1790_74#_c_1522_n 0.0268437f $X=8.725 $Y=1.91
+ $X2=0 $Y2=0
cc_833 N_A_1370_289#_c_996_n N_VPWR_c_1699_n 0.00343735f $X=6.94 $Y=2.21 $X2=0
+ $Y2=0
cc_834 N_A_1370_289#_c_1029_n N_VPWR_c_1700_n 0.0654619f $X=8.785 $Y=1.89 $X2=0
+ $Y2=0
cc_835 N_A_1370_289#_c_999_n N_VPWR_c_1701_n 0.00650548f $X=8.725 $Y=1.91 $X2=0
+ $Y2=0
cc_836 N_A_1370_289#_c_996_n N_VPWR_c_1696_n 9.49986e-19 $X=6.94 $Y=2.21 $X2=0
+ $Y2=0
cc_837 N_A_1370_289#_c_999_n N_VPWR_c_1696_n 0.00790777f $X=8.725 $Y=1.91 $X2=0
+ $Y2=0
cc_838 N_A_1370_289#_c_992_n N_VGND_M1012_d 0.010156f $X=8.495 $Y=0.842 $X2=0
+ $Y2=0
cc_839 N_A_1370_289#_M1001_g N_VGND_c_2105_n 6.00448e-19 $X=6.93 $Y=0.8 $X2=0
+ $Y2=0
cc_840 N_A_1370_289#_c_1027_n A_1401_118# 0.00138377f $X=7.21 $Y=1.005 $X2=-0.19
+ $Y2=-0.245
cc_841 N_A_1223_118#_c_1094_n N_A_852_74#_c_1208_n 0.00376247f $X=6.83 $Y=2.425
+ $X2=0 $Y2=0
cc_842 N_A_1223_118#_c_1094_n N_A_852_74#_c_1210_n 0.00100122f $X=6.83 $Y=2.425
+ $X2=0 $Y2=0
cc_843 N_A_1223_118#_c_1088_n N_A_852_74#_c_1212_n 0.00178964f $X=6.745 $Y=2.34
+ $X2=0 $Y2=0
cc_844 N_A_1223_118#_c_1094_n N_A_852_74#_c_1212_n 0.0126538f $X=6.83 $Y=2.425
+ $X2=0 $Y2=0
cc_845 N_A_1223_118#_c_1087_n N_A_852_74#_c_1213_n 0.0103562f $X=8.5 $Y=1.66
+ $X2=0 $Y2=0
cc_846 N_A_1223_118#_c_1101_n N_A_852_74#_c_1213_n 0.00267628f $X=7.38 $Y=2.425
+ $X2=0 $Y2=0
cc_847 N_A_1223_118#_c_1094_n N_A_852_74#_c_1213_n 0.00237118f $X=6.83 $Y=2.425
+ $X2=0 $Y2=0
cc_848 N_A_1223_118#_c_1089_n N_A_852_74#_c_1213_n 0.00749106f $X=7.465 $Y=2.32
+ $X2=0 $Y2=0
cc_849 N_A_1223_118#_c_1087_n N_A_852_74#_c_1214_n 0.00249951f $X=8.5 $Y=1.66
+ $X2=0 $Y2=0
cc_850 N_A_1223_118#_c_1087_n N_A_852_74#_M1016_g 0.00579836f $X=8.5 $Y=1.66
+ $X2=0 $Y2=0
cc_851 N_A_1223_118#_c_1087_n N_A_852_74#_c_1197_n 0.00845345f $X=8.5 $Y=1.66
+ $X2=0 $Y2=0
cc_852 N_A_1223_118#_c_1101_n N_VPWR_M1037_d 0.00731992f $X=7.38 $Y=2.425 $X2=0
+ $Y2=0
cc_853 N_A_1223_118#_c_1089_n N_VPWR_M1037_d 8.72177e-19 $X=7.465 $Y=2.32 $X2=0
+ $Y2=0
cc_854 N_A_1223_118#_c_1101_n N_VPWR_c_1699_n 0.0190336f $X=7.38 $Y=2.425 $X2=0
+ $Y2=0
cc_855 N_A_1223_118#_c_1094_n N_VPWR_c_1699_n 8.68953e-19 $X=6.83 $Y=2.425 $X2=0
+ $Y2=0
cc_856 N_A_1223_118#_c_1089_n N_VPWR_c_1699_n 0.00274183f $X=7.465 $Y=2.32 $X2=0
+ $Y2=0
cc_857 N_A_1223_118#_c_1087_n N_VPWR_c_1700_n 0.0179689f $X=8.5 $Y=1.66 $X2=0
+ $Y2=0
cc_858 N_A_1223_118#_c_1089_n N_VPWR_c_1700_n 0.0295999f $X=7.465 $Y=2.32 $X2=0
+ $Y2=0
cc_859 N_A_1223_118#_c_1091_n N_VPWR_c_1700_n 0.0170777f $X=8.425 $Y=1.41 $X2=0
+ $Y2=0
cc_860 N_A_1223_118#_c_1094_n N_VPWR_c_1709_n 0.00997198f $X=6.83 $Y=2.425 $X2=0
+ $Y2=0
cc_861 N_A_1223_118#_c_1089_n N_VPWR_c_1712_n 0.00745648f $X=7.465 $Y=2.32 $X2=0
+ $Y2=0
cc_862 N_A_1223_118#_c_1087_n N_VPWR_c_1696_n 8.51577e-19 $X=8.5 $Y=1.66 $X2=0
+ $Y2=0
cc_863 N_A_1223_118#_c_1101_n N_VPWR_c_1696_n 0.00974984f $X=7.38 $Y=2.425 $X2=0
+ $Y2=0
cc_864 N_A_1223_118#_c_1094_n N_VPWR_c_1696_n 0.019058f $X=6.83 $Y=2.425 $X2=0
+ $Y2=0
cc_865 N_A_1223_118#_c_1089_n N_VPWR_c_1696_n 0.0153115f $X=7.465 $Y=2.32 $X2=0
+ $Y2=0
cc_866 N_A_1223_118#_c_1094_n N_A_388_79#_c_1891_n 0.0161947f $X=6.83 $Y=2.425
+ $X2=0 $Y2=0
cc_867 N_A_1223_118#_c_1088_n N_A_388_79#_c_1883_n 0.00334791f $X=6.745 $Y=2.34
+ $X2=0 $Y2=0
cc_868 N_A_1223_118#_c_1088_n N_A_388_79#_c_1893_n 0.0130344f $X=6.745 $Y=2.34
+ $X2=0 $Y2=0
cc_869 N_A_1223_118#_c_1094_n N_A_388_79#_c_1893_n 0.0211069f $X=6.83 $Y=2.425
+ $X2=0 $Y2=0
cc_870 N_A_1223_118#_c_1119_n N_A_388_79#_c_1884_n 0.0240423f $X=6.66 $Y=0.8
+ $X2=0 $Y2=0
cc_871 N_A_1223_118#_c_1088_n N_A_388_79#_c_1884_n 0.0135678f $X=6.745 $Y=2.34
+ $X2=0 $Y2=0
cc_872 N_A_1223_118#_c_1088_n N_A_388_79#_c_1886_n 0.0518294f $X=6.745 $Y=2.34
+ $X2=0 $Y2=0
cc_873 N_A_1223_118#_c_1088_n N_A_388_79#_c_1896_n 0.00318798f $X=6.745 $Y=2.34
+ $X2=0 $Y2=0
cc_874 N_A_1223_118#_c_1094_n A_1325_457# 0.00189705f $X=6.83 $Y=2.425 $X2=-0.19
+ $Y2=-0.245
cc_875 N_A_1223_118#_M1003_g N_VGND_c_2098_n 0.00278271f $X=8.445 $Y=0.69 $X2=0
+ $Y2=0
cc_876 N_A_1223_118#_M1003_g N_VGND_c_2106_n 0.00116012f $X=8.445 $Y=0.69 $X2=0
+ $Y2=0
cc_877 N_A_1223_118#_M1003_g N_VGND_c_2110_n 0.00358525f $X=8.445 $Y=0.69 $X2=0
+ $Y2=0
cc_878 N_A_1223_118#_c_1119_n A_1323_118# 0.00139529f $X=6.66 $Y=0.8 $X2=-0.19
+ $Y2=-0.245
cc_879 N_A_852_74#_M1002_g N_A_2006_373#_M1045_g 0.0830829f $X=9.925 $Y=0.58
+ $X2=0 $Y2=0
cc_880 N_A_852_74#_M1016_g N_A_1790_74#_c_1522_n 0.00371138f $X=8.95 $Y=2.235
+ $X2=0 $Y2=0
cc_881 N_A_852_74#_M1002_g N_A_1790_74#_c_1531_n 0.0113037f $X=9.925 $Y=0.58
+ $X2=0 $Y2=0
cc_882 N_A_852_74#_M1002_g N_A_1790_74#_c_1502_n 0.00782202f $X=9.925 $Y=0.58
+ $X2=0 $Y2=0
cc_883 N_A_852_74#_c_1196_n N_A_1790_74#_c_1503_n 0.00624492f $X=9.85 $Y=1.55
+ $X2=0 $Y2=0
cc_884 N_A_852_74#_M1002_g N_A_1790_74#_c_1503_n 0.0034675f $X=9.925 $Y=0.58
+ $X2=0 $Y2=0
cc_885 N_A_852_74#_M1002_g N_A_1790_74#_c_1541_n 0.00668941f $X=9.925 $Y=0.58
+ $X2=0 $Y2=0
cc_886 N_A_852_74#_c_1220_n N_VPWR_M1022_d 0.00219658f $X=4.815 $Y=1.905 $X2=0
+ $Y2=0
cc_887 N_A_852_74#_c_1191_n N_VPWR_c_1698_n 0.00954491f $X=5.095 $Y=1.765 $X2=0
+ $Y2=0
cc_888 N_A_852_74#_c_1193_n N_VPWR_c_1698_n 0.00191176f $X=5.595 $Y=3.075 $X2=0
+ $Y2=0
cc_889 N_A_852_74#_c_1209_n N_VPWR_c_1698_n 0.00241263f $X=5.67 $Y=3.15 $X2=0
+ $Y2=0
cc_890 N_A_852_74#_c_1210_n N_VPWR_c_1699_n 0.00673937f $X=6.55 $Y=2.87 $X2=0
+ $Y2=0
cc_891 N_A_852_74#_c_1213_n N_VPWR_c_1699_n 0.0209699f $X=8.86 $Y=3.15 $X2=0
+ $Y2=0
cc_892 N_A_852_74#_c_1213_n N_VPWR_c_1700_n 0.0213056f $X=8.86 $Y=3.15 $X2=0
+ $Y2=0
cc_893 N_A_852_74#_c_1214_n N_VPWR_c_1700_n 0.00613773f $X=8.95 $Y=2.9 $X2=0
+ $Y2=0
cc_894 N_A_852_74#_M1016_g N_VPWR_c_1700_n 6.31058e-19 $X=8.95 $Y=2.235 $X2=0
+ $Y2=0
cc_895 N_A_852_74#_c_1213_n N_VPWR_c_1701_n 0.0188492f $X=8.86 $Y=3.15 $X2=0
+ $Y2=0
cc_896 N_A_852_74#_c_1191_n N_VPWR_c_1709_n 0.00413917f $X=5.095 $Y=1.765 $X2=0
+ $Y2=0
cc_897 N_A_852_74#_c_1209_n N_VPWR_c_1709_n 0.0483314f $X=5.67 $Y=3.15 $X2=0
+ $Y2=0
cc_898 N_A_852_74#_c_1213_n N_VPWR_c_1712_n 0.0266609f $X=8.86 $Y=3.15 $X2=0
+ $Y2=0
cc_899 N_A_852_74#_c_1191_n N_VPWR_c_1696_n 0.00408177f $X=5.095 $Y=1.765 $X2=0
+ $Y2=0
cc_900 N_A_852_74#_c_1208_n N_VPWR_c_1696_n 0.0232233f $X=6.46 $Y=3.15 $X2=0
+ $Y2=0
cc_901 N_A_852_74#_c_1209_n N_VPWR_c_1696_n 0.00703562f $X=5.67 $Y=3.15 $X2=0
+ $Y2=0
cc_902 N_A_852_74#_c_1213_n N_VPWR_c_1696_n 0.0678746f $X=8.86 $Y=3.15 $X2=0
+ $Y2=0
cc_903 N_A_852_74#_c_1219_n N_VPWR_c_1696_n 0.00503734f $X=6.55 $Y=3.15 $X2=0
+ $Y2=0
cc_904 N_A_852_74#_M1022_s N_A_388_79#_c_1891_n 0.0083322f $X=4.275 $Y=1.84
+ $X2=0 $Y2=0
cc_905 N_A_852_74#_c_1191_n N_A_388_79#_c_1891_n 0.0125138f $X=5.095 $Y=1.765
+ $X2=0 $Y2=0
cc_906 N_A_852_74#_c_1193_n N_A_388_79#_c_1891_n 0.0179108f $X=5.595 $Y=3.075
+ $X2=0 $Y2=0
cc_907 N_A_852_74#_c_1208_n N_A_388_79#_c_1891_n 0.00440485f $X=6.46 $Y=3.15
+ $X2=0 $Y2=0
cc_908 N_A_852_74#_c_1220_n N_A_388_79#_c_1891_n 0.00905317f $X=4.815 $Y=1.905
+ $X2=0 $Y2=0
cc_909 N_A_852_74#_c_1222_n N_A_388_79#_c_1891_n 0.0135649f $X=4.46 $Y=1.905
+ $X2=0 $Y2=0
cc_910 N_A_852_74#_c_1194_n N_A_388_79#_c_1883_n 0.00325896f $X=5.965 $Y=1.185
+ $X2=0 $Y2=0
cc_911 N_A_852_74#_c_1195_n N_A_388_79#_c_1883_n 0.00765017f $X=6.04 $Y=1.11
+ $X2=0 $Y2=0
cc_912 N_A_852_74#_c_1212_n N_A_388_79#_c_1893_n 7.86932e-19 $X=6.55 $Y=2.78
+ $X2=0 $Y2=0
cc_913 N_A_852_74#_c_1193_n N_A_388_79#_c_1894_n 0.00127172f $X=5.595 $Y=3.075
+ $X2=0 $Y2=0
cc_914 N_A_852_74#_c_1194_n N_A_388_79#_c_1884_n 0.00746021f $X=5.965 $Y=1.185
+ $X2=0 $Y2=0
cc_915 N_A_852_74#_c_1194_n N_A_388_79#_c_1885_n 0.0054134f $X=5.965 $Y=1.185
+ $X2=0 $Y2=0
cc_916 N_A_852_74#_c_1199_n N_A_388_79#_c_1886_n 0.00257569f $X=5.58 $Y=1.185
+ $X2=0 $Y2=0
cc_917 N_A_852_74#_M1006_g N_A_388_79#_c_1887_n 4.22867e-19 $X=5.05 $Y=0.74
+ $X2=0 $Y2=0
cc_918 N_A_852_74#_c_1194_n N_A_388_79#_c_1887_n 5.07577e-19 $X=5.965 $Y=1.185
+ $X2=0 $Y2=0
cc_919 N_A_852_74#_c_1195_n N_A_388_79#_c_1887_n 0.00211681f $X=6.04 $Y=1.11
+ $X2=0 $Y2=0
cc_920 N_A_852_74#_c_1199_n N_A_388_79#_c_1887_n 0.00489735f $X=5.58 $Y=1.185
+ $X2=0 $Y2=0
cc_921 N_A_852_74#_c_1193_n N_A_388_79#_c_1896_n 0.0034998f $X=5.595 $Y=3.075
+ $X2=0 $Y2=0
cc_922 N_A_852_74#_c_1200_n N_VGND_c_2085_n 0.0293125f $X=4.405 $Y=0.515 $X2=0
+ $Y2=0
cc_923 N_A_852_74#_M1006_g N_VGND_c_2086_n 0.00246929f $X=5.05 $Y=0.74 $X2=0
+ $Y2=0
cc_924 N_A_852_74#_c_1200_n N_VGND_c_2086_n 0.0295554f $X=4.405 $Y=0.515 $X2=0
+ $Y2=0
cc_925 N_A_852_74#_c_1204_n N_VGND_c_2086_n 0.0129884f $X=4.815 $Y=1.495 $X2=0
+ $Y2=0
cc_926 N_A_852_74#_M1002_g N_VGND_c_2087_n 0.00120934f $X=9.925 $Y=0.58 $X2=0
+ $Y2=0
cc_927 N_A_852_74#_c_1200_n N_VGND_c_2096_n 0.0147561f $X=4.405 $Y=0.515 $X2=0
+ $Y2=0
cc_928 N_A_852_74#_M1002_g N_VGND_c_2098_n 0.00298877f $X=9.925 $Y=0.58 $X2=0
+ $Y2=0
cc_929 N_A_852_74#_M1006_g N_VGND_c_2105_n 0.0043222f $X=5.05 $Y=0.74 $X2=0
+ $Y2=0
cc_930 N_A_852_74#_c_1195_n N_VGND_c_2105_n 6.21153e-19 $X=6.04 $Y=1.11 $X2=0
+ $Y2=0
cc_931 N_A_852_74#_M1006_g N_VGND_c_2110_n 0.00821137f $X=5.05 $Y=0.74 $X2=0
+ $Y2=0
cc_932 N_A_852_74#_M1002_g N_VGND_c_2110_n 0.00370514f $X=9.925 $Y=0.58 $X2=0
+ $Y2=0
cc_933 N_A_852_74#_c_1200_n N_VGND_c_2110_n 0.0121528f $X=4.405 $Y=0.515 $X2=0
+ $Y2=0
cc_934 N_A_2006_373#_c_1387_n N_A_1790_74#_M1018_g 0.00658176f $X=11.29 $Y=0.58
+ $X2=0 $Y2=0
cc_935 N_A_2006_373#_c_1389_n N_A_1790_74#_M1018_g 0.00562994f $X=11.455 $Y=0.79
+ $X2=0 $Y2=0
cc_936 N_A_2006_373#_c_1390_n N_A_1790_74#_M1018_g 0.00311727f $X=11.775 $Y=1.48
+ $X2=0 $Y2=0
cc_937 N_A_2006_373#_c_1385_n N_A_1790_74#_c_1495_n 0.0111503f $X=11.69 $Y=1.565
+ $X2=0 $Y2=0
cc_938 N_A_2006_373#_c_1388_n N_A_1790_74#_c_1495_n 0.00258531f $X=11.69 $Y=0.79
+ $X2=0 $Y2=0
cc_939 N_A_2006_373#_c_1389_n N_A_1790_74#_c_1495_n 0.0075729f $X=11.455 $Y=0.79
+ $X2=0 $Y2=0
cc_940 N_A_2006_373#_c_1390_n N_A_1790_74#_c_1495_n 0.00284108f $X=11.775
+ $Y=1.48 $X2=0 $Y2=0
cc_941 N_A_2006_373#_c_1385_n N_A_1790_74#_c_1505_n 0.00952908f $X=11.69
+ $Y=1.565 $X2=0 $Y2=0
cc_942 N_A_2006_373#_c_1397_n N_A_1790_74#_c_1506_n 0.00686533f $X=11.23
+ $Y=2.405 $X2=0 $Y2=0
cc_943 N_A_2006_373#_c_1385_n N_A_1790_74#_c_1496_n 0.0131208f $X=11.69 $Y=1.565
+ $X2=0 $Y2=0
cc_944 N_A_2006_373#_c_1388_n N_A_1790_74#_c_1496_n 0.00113849f $X=11.69 $Y=0.79
+ $X2=0 $Y2=0
cc_945 N_A_2006_373#_c_1390_n N_A_1790_74#_c_1496_n 0.0180935f $X=11.775 $Y=1.48
+ $X2=0 $Y2=0
cc_946 N_A_2006_373#_c_1387_n N_A_1790_74#_M1028_g 0.00446735f $X=11.29 $Y=0.58
+ $X2=0 $Y2=0
cc_947 N_A_2006_373#_c_1388_n N_A_1790_74#_M1028_g 0.00377396f $X=11.69 $Y=0.79
+ $X2=0 $Y2=0
cc_948 N_A_2006_373#_c_1390_n N_A_1790_74#_M1028_g 0.00455681f $X=11.775 $Y=1.48
+ $X2=0 $Y2=0
cc_949 N_A_2006_373#_c_1385_n N_A_1790_74#_c_1499_n 5.76097e-19 $X=11.69
+ $Y=1.565 $X2=0 $Y2=0
cc_950 N_A_2006_373#_c_1391_n N_A_1790_74#_c_1522_n 0.0150017f $X=10.12 $Y=2.28
+ $X2=0 $Y2=0
cc_951 N_A_2006_373#_c_1396_n N_A_1790_74#_c_1522_n 0.0109254f $X=10.545
+ $Y=2.405 $X2=0 $Y2=0
cc_952 N_A_2006_373#_M1045_g N_A_1790_74#_c_1531_n 0.00245703f $X=10.285 $Y=0.58
+ $X2=0 $Y2=0
cc_953 N_A_2006_373#_M1045_g N_A_1790_74#_c_1502_n 0.00544577f $X=10.285 $Y=0.58
+ $X2=0 $Y2=0
cc_954 N_A_2006_373#_c_1391_n N_A_1790_74#_c_1503_n 0.00156196f $X=10.12 $Y=2.28
+ $X2=0 $Y2=0
cc_955 N_A_2006_373#_M1045_g N_A_1790_74#_c_1503_n 0.0092441f $X=10.285 $Y=0.58
+ $X2=0 $Y2=0
cc_956 N_A_2006_373#_c_1393_n N_A_1790_74#_c_1503_n 0.0474407f $X=10.405 $Y=2.03
+ $X2=0 $Y2=0
cc_957 N_A_2006_373#_c_1386_n N_A_1790_74#_c_1503_n 0.0135848f $X=10.545
+ $Y=1.565 $X2=0 $Y2=0
cc_958 N_A_2006_373#_c_1396_n N_A_1790_74#_c_1503_n 0.00357879f $X=10.545
+ $Y=2.405 $X2=0 $Y2=0
cc_959 N_A_2006_373#_c_1398_n N_A_1790_74#_c_1503_n 0.0108982f $X=10.285
+ $Y=2.072 $X2=0 $Y2=0
cc_960 N_A_2006_373#_M1045_g N_A_1790_74#_c_1504_n 0.0192761f $X=10.285 $Y=0.58
+ $X2=0 $Y2=0
cc_961 N_A_2006_373#_c_1385_n N_A_1790_74#_c_1504_n 0.0718198f $X=11.69 $Y=1.565
+ $X2=0 $Y2=0
cc_962 N_A_2006_373#_c_1386_n N_A_1790_74#_c_1504_n 0.0235777f $X=10.545
+ $Y=1.565 $X2=0 $Y2=0
cc_963 N_A_2006_373#_c_1388_n N_A_1790_74#_c_1504_n 0.00476671f $X=11.69 $Y=0.79
+ $X2=0 $Y2=0
cc_964 N_A_2006_373#_c_1389_n N_A_1790_74#_c_1504_n 0.026725f $X=11.455 $Y=0.79
+ $X2=0 $Y2=0
cc_965 N_A_2006_373#_c_1390_n N_A_1790_74#_c_1504_n 0.0207312f $X=11.775 $Y=1.48
+ $X2=0 $Y2=0
cc_966 N_A_2006_373#_c_1398_n N_A_1790_74#_c_1504_n 0.00394383f $X=10.285
+ $Y=2.072 $X2=0 $Y2=0
cc_967 N_A_2006_373#_c_1395_n N_VPWR_M1038_d 0.00487963f $X=11.065 $Y=2.405
+ $X2=0 $Y2=0
cc_968 N_A_2006_373#_c_1396_n N_VPWR_M1038_d 0.00589954f $X=10.545 $Y=2.405
+ $X2=0 $Y2=0
cc_969 N_A_2006_373#_c_1391_n N_VPWR_c_1701_n 0.00419312f $X=10.12 $Y=2.28 $X2=0
+ $Y2=0
cc_970 N_A_2006_373#_c_1385_n N_VPWR_c_1702_n 0.0223739f $X=11.69 $Y=1.565 $X2=0
+ $Y2=0
cc_971 N_A_2006_373#_c_1397_n N_VPWR_c_1702_n 0.031333f $X=11.23 $Y=2.405 $X2=0
+ $Y2=0
cc_972 N_A_2006_373#_c_1397_n N_VPWR_c_1713_n 0.00802713f $X=11.23 $Y=2.405
+ $X2=0 $Y2=0
cc_973 N_A_2006_373#_c_1391_n N_VPWR_c_1721_n 0.0101552f $X=10.12 $Y=2.28 $X2=0
+ $Y2=0
cc_974 N_A_2006_373#_c_1395_n N_VPWR_c_1721_n 0.0240529f $X=11.065 $Y=2.405
+ $X2=0 $Y2=0
cc_975 N_A_2006_373#_c_1396_n N_VPWR_c_1721_n 0.0238431f $X=10.545 $Y=2.405
+ $X2=0 $Y2=0
cc_976 N_A_2006_373#_c_1397_n N_VPWR_c_1721_n 0.0095412f $X=11.23 $Y=2.405 $X2=0
+ $Y2=0
cc_977 N_A_2006_373#_c_1398_n N_VPWR_c_1721_n 0.00121809f $X=10.285 $Y=2.072
+ $X2=0 $Y2=0
cc_978 N_A_2006_373#_c_1391_n N_VPWR_c_1696_n 0.00489211f $X=10.12 $Y=2.28 $X2=0
+ $Y2=0
cc_979 N_A_2006_373#_c_1395_n N_VPWR_c_1696_n 0.00766785f $X=11.065 $Y=2.405
+ $X2=0 $Y2=0
cc_980 N_A_2006_373#_c_1396_n N_VPWR_c_1696_n 0.00101543f $X=10.545 $Y=2.405
+ $X2=0 $Y2=0
cc_981 N_A_2006_373#_c_1397_n N_VPWR_c_1696_n 0.010512f $X=11.23 $Y=2.405 $X2=0
+ $Y2=0
cc_982 N_A_2006_373#_c_1385_n Q_N 0.0138399f $X=11.69 $Y=1.565 $X2=0 $Y2=0
cc_983 N_A_2006_373#_c_1388_n N_Q_N_c_2041_n 0.00970057f $X=11.69 $Y=0.79 $X2=0
+ $Y2=0
cc_984 N_A_2006_373#_c_1390_n N_Q_N_c_2041_n 0.00199024f $X=11.775 $Y=1.48 $X2=0
+ $Y2=0
cc_985 N_A_2006_373#_c_1390_n Q_N 0.0415299f $X=11.775 $Y=1.48 $X2=0 $Y2=0
cc_986 N_A_2006_373#_c_1388_n N_VGND_M1028_s 0.00517852f $X=11.69 $Y=0.79 $X2=0
+ $Y2=0
cc_987 N_A_2006_373#_c_1390_n N_VGND_M1028_s 0.00675628f $X=11.775 $Y=1.48 $X2=0
+ $Y2=0
cc_988 N_A_2006_373#_M1045_g N_VGND_c_2087_n 0.0105628f $X=10.285 $Y=0.58 $X2=0
+ $Y2=0
cc_989 N_A_2006_373#_c_1387_n N_VGND_c_2087_n 0.0118606f $X=11.29 $Y=0.58 $X2=0
+ $Y2=0
cc_990 N_A_2006_373#_c_1389_n N_VGND_c_2087_n 0.00372607f $X=11.455 $Y=0.79
+ $X2=0 $Y2=0
cc_991 N_A_2006_373#_c_1387_n N_VGND_c_2088_n 0.0139523f $X=11.29 $Y=0.58 $X2=0
+ $Y2=0
cc_992 N_A_2006_373#_c_1388_n N_VGND_c_2088_n 0.0181192f $X=11.69 $Y=0.79 $X2=0
+ $Y2=0
cc_993 N_A_2006_373#_M1045_g N_VGND_c_2098_n 0.00383152f $X=10.285 $Y=0.58 $X2=0
+ $Y2=0
cc_994 N_A_2006_373#_c_1387_n N_VGND_c_2101_n 0.0142949f $X=11.29 $Y=0.58 $X2=0
+ $Y2=0
cc_995 N_A_2006_373#_c_1388_n N_VGND_c_2101_n 0.00298753f $X=11.69 $Y=0.79 $X2=0
+ $Y2=0
cc_996 N_A_2006_373#_M1045_g N_VGND_c_2110_n 0.0075694f $X=10.285 $Y=0.58 $X2=0
+ $Y2=0
cc_997 N_A_2006_373#_c_1387_n N_VGND_c_2110_n 0.011894f $X=11.29 $Y=0.58 $X2=0
+ $Y2=0
cc_998 N_A_2006_373#_c_1388_n N_VGND_c_2110_n 0.00611276f $X=11.69 $Y=0.79 $X2=0
+ $Y2=0
cc_999 N_A_1790_74#_c_1499_n N_A_2604_392#_c_1647_n 0.0166552f $X=12.945
+ $Y=1.585 $X2=0 $Y2=0
cc_1000 N_A_1790_74#_c_1500_n N_A_2604_392#_c_1647_n 0.00200517f $X=12.945
+ $Y=1.795 $X2=0 $Y2=0
cc_1001 N_A_1790_74#_M1010_g N_A_2604_392#_c_1649_n 0.0121223f $X=12.99 $Y=0.69
+ $X2=0 $Y2=0
cc_1002 N_A_1790_74#_c_1500_n N_A_2604_392#_c_1650_n 0.0108738f $X=12.945
+ $Y=1.795 $X2=0 $Y2=0
cc_1003 N_A_1790_74#_c_1511_n N_A_2604_392#_c_1650_n 0.00283082f $X=12.945
+ $Y=1.885 $X2=0 $Y2=0
cc_1004 N_A_1790_74#_c_1499_n N_A_2604_392#_c_1651_n 0.0099279f $X=12.945
+ $Y=1.585 $X2=0 $Y2=0
cc_1005 N_A_1790_74#_c_1500_n N_A_2604_392#_c_1651_n 0.00145958f $X=12.945
+ $Y=1.795 $X2=0 $Y2=0
cc_1006 N_A_1790_74#_c_1522_n N_VPWR_c_1701_n 0.0165613f $X=9.925 $Y=2.53 $X2=0
+ $Y2=0
cc_1007 N_A_1790_74#_c_1505_n N_VPWR_c_1702_n 0.00657334f $X=11.455 $Y=2.19
+ $X2=0 $Y2=0
cc_1008 N_A_1790_74#_c_1506_n N_VPWR_c_1702_n 0.00817866f $X=11.455 $Y=2.28
+ $X2=0 $Y2=0
cc_1009 N_A_1790_74#_c_1496_n N_VPWR_c_1702_n 0.00168841f $X=11.9 $Y=1.422 $X2=0
+ $Y2=0
cc_1010 N_A_1790_74#_c_1507_n N_VPWR_c_1702_n 0.00877379f $X=11.99 $Y=1.765
+ $X2=0 $Y2=0
cc_1011 N_A_1790_74#_c_1508_n N_VPWR_c_1703_n 0.00328506f $X=12.44 $Y=1.765
+ $X2=0 $Y2=0
cc_1012 N_A_1790_74#_c_1499_n N_VPWR_c_1703_n 0.0105801f $X=12.945 $Y=1.585
+ $X2=0 $Y2=0
cc_1013 N_A_1790_74#_c_1511_n N_VPWR_c_1703_n 0.00894992f $X=12.945 $Y=1.885
+ $X2=0 $Y2=0
cc_1014 N_A_1790_74#_c_1511_n N_VPWR_c_1704_n 0.00461748f $X=12.945 $Y=1.885
+ $X2=0 $Y2=0
cc_1015 N_A_1790_74#_c_1506_n N_VPWR_c_1713_n 0.00443738f $X=11.455 $Y=2.28
+ $X2=0 $Y2=0
cc_1016 N_A_1790_74#_c_1507_n N_VPWR_c_1714_n 0.00422942f $X=11.99 $Y=1.765
+ $X2=0 $Y2=0
cc_1017 N_A_1790_74#_c_1508_n N_VPWR_c_1714_n 0.00461464f $X=12.44 $Y=1.765
+ $X2=0 $Y2=0
cc_1018 N_A_1790_74#_c_1511_n N_VPWR_c_1715_n 0.00461464f $X=12.945 $Y=1.885
+ $X2=0 $Y2=0
cc_1019 N_A_1790_74#_c_1522_n N_VPWR_c_1721_n 0.00301353f $X=9.925 $Y=2.53 $X2=0
+ $Y2=0
cc_1020 N_A_1790_74#_c_1506_n N_VPWR_c_1696_n 0.00489211f $X=11.455 $Y=2.28
+ $X2=0 $Y2=0
cc_1021 N_A_1790_74#_c_1507_n N_VPWR_c_1696_n 0.00789017f $X=11.99 $Y=1.765
+ $X2=0 $Y2=0
cc_1022 N_A_1790_74#_c_1508_n N_VPWR_c_1696_n 0.0090856f $X=12.44 $Y=1.765 $X2=0
+ $Y2=0
cc_1023 N_A_1790_74#_c_1511_n N_VPWR_c_1696_n 0.00913697f $X=12.945 $Y=1.885
+ $X2=0 $Y2=0
cc_1024 N_A_1790_74#_c_1522_n N_VPWR_c_1696_n 0.0291224f $X=9.925 $Y=2.53 $X2=0
+ $Y2=0
cc_1025 N_A_1790_74#_c_1522_n A_1955_471# 0.00419128f $X=9.925 $Y=2.53 $X2=-0.19
+ $Y2=-0.245
cc_1026 N_A_1790_74#_c_1505_n Q_N 9.68335e-19 $X=11.455 $Y=2.19 $X2=0 $Y2=0
cc_1027 N_A_1790_74#_c_1507_n Q_N 0.0159647f $X=11.99 $Y=1.765 $X2=0 $Y2=0
cc_1028 N_A_1790_74#_M1028_g Q_N 0.00434424f $X=12.085 $Y=0.74 $X2=0 $Y2=0
cc_1029 N_A_1790_74#_c_1508_n Q_N 0.00257754f $X=12.44 $Y=1.765 $X2=0 $Y2=0
cc_1030 N_A_1790_74#_M1039_g Q_N 0.00444052f $X=12.515 $Y=0.74 $X2=0 $Y2=0
cc_1031 N_A_1790_74#_c_1499_n Q_N 0.0512546f $X=12.945 $Y=1.585 $X2=0 $Y2=0
cc_1032 N_A_1790_74#_c_1500_n Q_N 8.09244e-19 $X=12.945 $Y=1.795 $X2=0 $Y2=0
cc_1033 N_A_1790_74#_M1028_g N_Q_N_c_2041_n 0.0129348f $X=12.085 $Y=0.74 $X2=0
+ $Y2=0
cc_1034 N_A_1790_74#_M1039_g N_Q_N_c_2041_n 0.0062067f $X=12.515 $Y=0.74 $X2=0
+ $Y2=0
cc_1035 N_A_1790_74#_M1010_g N_Q_N_c_2041_n 2.82358e-19 $X=12.99 $Y=0.69 $X2=0
+ $Y2=0
cc_1036 N_A_1790_74#_M1028_g Q_N 0.00845569f $X=12.085 $Y=0.74 $X2=0 $Y2=0
cc_1037 N_A_1790_74#_M1039_g Q_N 0.00357919f $X=12.515 $Y=0.74 $X2=0 $Y2=0
cc_1038 N_A_1790_74#_M1018_g N_VGND_c_2087_n 0.00182072f $X=11.075 $Y=0.58 $X2=0
+ $Y2=0
cc_1039 N_A_1790_74#_c_1531_n N_VGND_c_2087_n 0.0208351f $X=9.925 $Y=0.57 $X2=0
+ $Y2=0
cc_1040 N_A_1790_74#_c_1502_n N_VGND_c_2087_n 0.00424796f $X=10.01 $Y=1.045
+ $X2=0 $Y2=0
cc_1041 N_A_1790_74#_c_1504_n N_VGND_c_2087_n 0.0223381f $X=11.355 $Y=1.175
+ $X2=0 $Y2=0
cc_1042 N_A_1790_74#_M1018_g N_VGND_c_2088_n 0.00310691f $X=11.075 $Y=0.58 $X2=0
+ $Y2=0
cc_1043 N_A_1790_74#_M1028_g N_VGND_c_2088_n 0.00814486f $X=12.085 $Y=0.74 $X2=0
+ $Y2=0
cc_1044 N_A_1790_74#_M1039_g N_VGND_c_2089_n 0.0030832f $X=12.515 $Y=0.74 $X2=0
+ $Y2=0
cc_1045 N_A_1790_74#_c_1499_n N_VGND_c_2089_n 0.00620549f $X=12.945 $Y=1.585
+ $X2=0 $Y2=0
cc_1046 N_A_1790_74#_M1010_g N_VGND_c_2089_n 0.00352391f $X=12.99 $Y=0.69 $X2=0
+ $Y2=0
cc_1047 N_A_1790_74#_M1010_g N_VGND_c_2090_n 0.00461464f $X=12.99 $Y=0.69 $X2=0
+ $Y2=0
cc_1048 N_A_1790_74#_M1010_g N_VGND_c_2091_n 0.00385314f $X=12.99 $Y=0.69 $X2=0
+ $Y2=0
cc_1049 N_A_1790_74#_c_1531_n N_VGND_c_2098_n 0.0202724f $X=9.925 $Y=0.57 $X2=0
+ $Y2=0
cc_1050 N_A_1790_74#_M1018_g N_VGND_c_2101_n 0.00434272f $X=11.075 $Y=0.58 $X2=0
+ $Y2=0
cc_1051 N_A_1790_74#_M1028_g N_VGND_c_2102_n 0.00434272f $X=12.085 $Y=0.74 $X2=0
+ $Y2=0
cc_1052 N_A_1790_74#_M1039_g N_VGND_c_2102_n 0.00434272f $X=12.515 $Y=0.74 $X2=0
+ $Y2=0
cc_1053 N_A_1790_74#_M1018_g N_VGND_c_2110_n 0.00825669f $X=11.075 $Y=0.58 $X2=0
+ $Y2=0
cc_1054 N_A_1790_74#_M1028_g N_VGND_c_2110_n 0.00826269f $X=12.085 $Y=0.74 $X2=0
+ $Y2=0
cc_1055 N_A_1790_74#_M1039_g N_VGND_c_2110_n 0.00820493f $X=12.515 $Y=0.74 $X2=0
+ $Y2=0
cc_1056 N_A_1790_74#_M1010_g N_VGND_c_2110_n 0.00912981f $X=12.99 $Y=0.69 $X2=0
+ $Y2=0
cc_1057 N_A_1790_74#_c_1531_n N_VGND_c_2110_n 0.0221648f $X=9.925 $Y=0.57 $X2=0
+ $Y2=0
cc_1058 N_A_1790_74#_c_1531_n A_2000_74# 0.00371855f $X=9.925 $Y=0.57 $X2=-0.19
+ $Y2=-0.245
cc_1059 N_A_1790_74#_c_1502_n A_2000_74# 5.09211e-19 $X=10.01 $Y=1.045 $X2=-0.19
+ $Y2=-0.245
cc_1060 N_A_2604_392#_c_1650_n N_VPWR_c_1703_n 0.00374141f $X=13.17 $Y=2.105
+ $X2=0 $Y2=0
cc_1061 N_A_2604_392#_c_1652_n N_VPWR_c_1704_n 0.0177685f $X=13.935 $Y=1.765
+ $X2=0 $Y2=0
cc_1062 N_A_2604_392#_c_1653_n N_VPWR_c_1704_n 6.92538e-19 $X=14.385 $Y=1.765
+ $X2=0 $Y2=0
cc_1063 N_A_2604_392#_c_1647_n N_VPWR_c_1704_n 0.00687596f $X=13.845 $Y=1.465
+ $X2=0 $Y2=0
cc_1064 N_A_2604_392#_c_1648_n N_VPWR_c_1704_n 4.36456e-19 $X=14.385 $Y=1.532
+ $X2=0 $Y2=0
cc_1065 N_A_2604_392#_c_1650_n N_VPWR_c_1704_n 0.0792204f $X=13.17 $Y=2.105
+ $X2=0 $Y2=0
cc_1066 N_A_2604_392#_c_1669_p N_VPWR_c_1704_n 0.0253438f $X=13.8 $Y=1.465 $X2=0
+ $Y2=0
cc_1067 N_A_2604_392#_c_1653_n N_VPWR_c_1706_n 0.00508676f $X=14.385 $Y=1.765
+ $X2=0 $Y2=0
cc_1068 N_A_2604_392#_c_1650_n N_VPWR_c_1715_n 0.0115122f $X=13.17 $Y=2.105
+ $X2=0 $Y2=0
cc_1069 N_A_2604_392#_c_1652_n N_VPWR_c_1716_n 0.00413917f $X=13.935 $Y=1.765
+ $X2=0 $Y2=0
cc_1070 N_A_2604_392#_c_1653_n N_VPWR_c_1716_n 0.00445602f $X=14.385 $Y=1.765
+ $X2=0 $Y2=0
cc_1071 N_A_2604_392#_c_1652_n N_VPWR_c_1696_n 0.00817726f $X=13.935 $Y=1.765
+ $X2=0 $Y2=0
cc_1072 N_A_2604_392#_c_1653_n N_VPWR_c_1696_n 0.00860378f $X=14.385 $Y=1.765
+ $X2=0 $Y2=0
cc_1073 N_A_2604_392#_c_1650_n N_VPWR_c_1696_n 0.0095288f $X=13.17 $Y=2.105
+ $X2=0 $Y2=0
cc_1074 N_A_2604_392#_c_1649_n Q_N 0.00105746f $X=13.205 $Y=0.515 $X2=0 $Y2=0
cc_1075 N_A_2604_392#_c_1652_n N_Q_c_2068_n 0.00199967f $X=13.935 $Y=1.765 $X2=0
+ $Y2=0
cc_1076 N_A_2604_392#_M1025_g N_Q_c_2068_n 0.00531072f $X=13.97 $Y=0.74 $X2=0
+ $Y2=0
cc_1077 N_A_2604_392#_c_1653_n N_Q_c_2068_n 0.0153858f $X=14.385 $Y=1.765 $X2=0
+ $Y2=0
cc_1078 N_A_2604_392#_M1040_g N_Q_c_2068_n 0.00534388f $X=14.4 $Y=0.74 $X2=0
+ $Y2=0
cc_1079 N_A_2604_392#_c_1648_n N_Q_c_2068_n 0.045774f $X=14.385 $Y=1.532 $X2=0
+ $Y2=0
cc_1080 N_A_2604_392#_c_1669_p N_Q_c_2068_n 0.0258081f $X=13.8 $Y=1.465 $X2=0
+ $Y2=0
cc_1081 N_A_2604_392#_c_1649_n N_VGND_c_2089_n 0.0303376f $X=13.205 $Y=0.515
+ $X2=0 $Y2=0
cc_1082 N_A_2604_392#_c_1649_n N_VGND_c_2090_n 0.0115122f $X=13.205 $Y=0.515
+ $X2=0 $Y2=0
cc_1083 N_A_2604_392#_M1025_g N_VGND_c_2091_n 0.00508752f $X=13.97 $Y=0.74 $X2=0
+ $Y2=0
cc_1084 N_A_2604_392#_c_1647_n N_VGND_c_2091_n 0.00391367f $X=13.845 $Y=1.465
+ $X2=0 $Y2=0
cc_1085 N_A_2604_392#_c_1649_n N_VGND_c_2091_n 0.0350664f $X=13.205 $Y=0.515
+ $X2=0 $Y2=0
cc_1086 N_A_2604_392#_c_1669_p N_VGND_c_2091_n 0.014168f $X=13.8 $Y=1.465 $X2=0
+ $Y2=0
cc_1087 N_A_2604_392#_M1040_g N_VGND_c_2093_n 0.00543765f $X=14.4 $Y=0.74 $X2=0
+ $Y2=0
cc_1088 N_A_2604_392#_M1025_g N_VGND_c_2103_n 0.00461464f $X=13.97 $Y=0.74 $X2=0
+ $Y2=0
cc_1089 N_A_2604_392#_M1040_g N_VGND_c_2103_n 0.00461464f $X=14.4 $Y=0.74 $X2=0
+ $Y2=0
cc_1090 N_A_2604_392#_M1025_g N_VGND_c_2110_n 0.00913331f $X=13.97 $Y=0.74 $X2=0
+ $Y2=0
cc_1091 N_A_2604_392#_M1040_g N_VGND_c_2110_n 0.00911154f $X=14.4 $Y=0.74 $X2=0
+ $Y2=0
cc_1092 N_A_2604_392#_c_1649_n N_VGND_c_2110_n 0.0095288f $X=13.205 $Y=0.515
+ $X2=0 $Y2=0
cc_1093 N_VPWR_c_1711_n N_A_388_79#_c_1898_n 0.0287061f $X=3.115 $Y=3.33 $X2=0
+ $Y2=0
cc_1094 N_VPWR_c_1718_n N_A_388_79#_c_1898_n 0.00580289f $X=1.4 $Y=3.072 $X2=0
+ $Y2=0
cc_1095 N_VPWR_c_1696_n N_A_388_79#_c_1898_n 0.0336043f $X=14.64 $Y=3.33 $X2=0
+ $Y2=0
cc_1096 N_VPWR_M1005_d N_A_388_79#_c_1921_n 0.0107616f $X=3.11 $Y=2.32 $X2=0
+ $Y2=0
cc_1097 N_VPWR_c_1697_n N_A_388_79#_c_1921_n 0.0220425f $X=3.28 $Y=2.78 $X2=0
+ $Y2=0
cc_1098 N_VPWR_c_1696_n N_A_388_79#_c_1921_n 0.00587028f $X=14.64 $Y=3.33 $X2=0
+ $Y2=0
cc_1099 N_VPWR_c_1697_n N_A_388_79#_c_1890_n 0.0251321f $X=3.28 $Y=2.78 $X2=0
+ $Y2=0
cc_1100 N_VPWR_c_1707_n N_A_388_79#_c_1890_n 0.0166395f $X=4.705 $Y=3.33 $X2=0
+ $Y2=0
cc_1101 N_VPWR_c_1696_n N_A_388_79#_c_1890_n 0.0136379f $X=14.64 $Y=3.33 $X2=0
+ $Y2=0
cc_1102 N_VPWR_M1022_d N_A_388_79#_c_1891_n 0.00447753f $X=4.72 $Y=1.84 $X2=0
+ $Y2=0
cc_1103 N_VPWR_c_1698_n N_A_388_79#_c_1891_n 0.0172192f $X=4.87 $Y=2.795 $X2=0
+ $Y2=0
cc_1104 N_VPWR_c_1709_n N_A_388_79#_c_1891_n 0.00579387f $X=7.07 $Y=3.33 $X2=0
+ $Y2=0
cc_1105 N_VPWR_c_1696_n N_A_388_79#_c_1891_n 0.0543728f $X=14.64 $Y=3.33 $X2=0
+ $Y2=0
cc_1106 N_VPWR_M1005_d N_A_388_79#_c_1892_n 6.64982e-19 $X=3.11 $Y=2.32 $X2=0
+ $Y2=0
cc_1107 N_VPWR_c_1696_n N_A_388_79#_c_1892_n 0.00603182f $X=14.64 $Y=3.33 $X2=0
+ $Y2=0
cc_1108 N_VPWR_c_1702_n Q_N 0.0844051f $X=11.765 $Y=1.985 $X2=0 $Y2=0
cc_1109 N_VPWR_c_1703_n Q_N 0.00150368f $X=12.665 $Y=2.085 $X2=0 $Y2=0
cc_1110 N_VPWR_c_1714_n Q_N 0.014534f $X=12.54 $Y=3.33 $X2=0 $Y2=0
cc_1111 N_VPWR_c_1696_n Q_N 0.0119501f $X=14.64 $Y=3.33 $X2=0 $Y2=0
cc_1112 N_VPWR_c_1704_n N_Q_c_2068_n 0.0430489f $X=13.71 $Y=1.985 $X2=0 $Y2=0
cc_1113 N_VPWR_c_1706_n N_Q_c_2068_n 0.0437503f $X=14.61 $Y=1.985 $X2=0 $Y2=0
cc_1114 N_VPWR_c_1716_n N_Q_c_2068_n 0.0119166f $X=14.495 $Y=3.33 $X2=0 $Y2=0
cc_1115 N_VPWR_c_1696_n N_Q_c_2068_n 0.00983061f $X=14.64 $Y=3.33 $X2=0 $Y2=0
cc_1116 N_A_388_79#_c_1898_n A_538_464# 0.00358318f $X=2.775 $Y=2.785 $X2=-0.19
+ $Y2=-0.245
cc_1117 N_A_388_79#_c_1900_n A_538_464# 0.00186299f $X=2.86 $Y=2.66 $X2=-0.19
+ $Y2=-0.245
cc_1118 N_A_388_79#_c_1888_n A_538_464# 0.00712083f $X=2.945 $Y=2.405 $X2=-0.19
+ $Y2=-0.245
cc_1119 N_A_388_79#_M1029_d N_noxref_25_c_2242_n 0.011077f $X=1.94 $Y=0.395
+ $X2=0 $Y2=0
cc_1120 N_A_388_79#_c_1879_n N_noxref_25_c_2242_n 0.0217278f $X=2.435 $Y=0.68
+ $X2=0 $Y2=0
cc_1121 N_A_388_79#_c_1880_n N_noxref_25_c_2242_n 0.0118204f $X=3.445 $Y=1.09
+ $X2=0 $Y2=0
cc_1122 N_A_388_79#_c_1879_n N_noxref_25_c_2244_n 0.00763776f $X=2.435 $Y=0.68
+ $X2=0 $Y2=0
cc_1123 N_A_388_79#_c_1880_n N_noxref_25_c_2244_n 0.0271448f $X=3.445 $Y=1.09
+ $X2=0 $Y2=0
cc_1124 N_Q_N_c_2041_n N_VGND_c_2088_n 0.010788f $X=12.3 $Y=0.515 $X2=0 $Y2=0
cc_1125 N_Q_N_c_2041_n N_VGND_c_2089_n 0.0272093f $X=12.3 $Y=0.515 $X2=0 $Y2=0
cc_1126 N_Q_N_c_2041_n N_VGND_c_2102_n 0.0144922f $X=12.3 $Y=0.515 $X2=0 $Y2=0
cc_1127 N_Q_N_c_2041_n N_VGND_c_2110_n 0.0118826f $X=12.3 $Y=0.515 $X2=0 $Y2=0
cc_1128 N_Q_c_2068_n N_VGND_c_2091_n 0.00251281f $X=14.185 $Y=0.515 $X2=0 $Y2=0
cc_1129 N_Q_c_2068_n N_VGND_c_2093_n 0.0305242f $X=14.185 $Y=0.515 $X2=0 $Y2=0
cc_1130 N_Q_c_2068_n N_VGND_c_2103_n 0.0119584f $X=14.185 $Y=0.515 $X2=0 $Y2=0
cc_1131 N_Q_c_2068_n N_VGND_c_2110_n 0.00989813f $X=14.185 $Y=0.515 $X2=0 $Y2=0
cc_1132 N_VGND_c_2084_n N_noxref_25_c_2241_n 0.0278855f $X=0.71 $Y=0.605 $X2=0
+ $Y2=0
cc_1133 N_VGND_c_2085_n N_noxref_25_c_2242_n 0.0122221f $X=3.805 $Y=0.605 $X2=0
+ $Y2=0
cc_1134 N_VGND_c_2094_n N_noxref_25_c_2242_n 0.136372f $X=3.64 $Y=0 $X2=0 $Y2=0
cc_1135 N_VGND_c_2110_n N_noxref_25_c_2242_n 0.078753f $X=14.64 $Y=0 $X2=0 $Y2=0
cc_1136 N_VGND_c_2084_n N_noxref_25_c_2243_n 0.0125436f $X=0.71 $Y=0.605 $X2=0
+ $Y2=0
cc_1137 N_VGND_c_2094_n N_noxref_25_c_2243_n 0.0177095f $X=3.64 $Y=0 $X2=0 $Y2=0
cc_1138 N_VGND_c_2110_n N_noxref_25_c_2243_n 0.00967952f $X=14.64 $Y=0 $X2=0
+ $Y2=0
cc_1139 N_VGND_c_2085_n N_noxref_25_c_2244_n 0.0270495f $X=3.805 $Y=0.605 $X2=0
+ $Y2=0
cc_1140 N_noxref_25_c_2242_n noxref_26 0.00198134f $X=3.1 $Y=0.34 $X2=-0.19
+ $Y2=-0.245
cc_1141 N_noxref_25_c_2242_n noxref_27 0.00246354f $X=3.1 $Y=0.34 $X2=-0.19
+ $Y2=-0.245
