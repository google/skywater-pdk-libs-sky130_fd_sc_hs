* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hs__sedfxtp_1 CLK D DE SCD SCE VGND VNB VPB VPWR Q
M1000 a_27_74# a_547_301# a_554_463# VPB pshort w=640000u l=150000u
+  ad=3.744e+11p pd=3.73e+06u as=1.536e+11p ps=1.76e+06u
M1001 a_2385_74# a_1295_74# a_2274_392# VPB pshort w=1e+06u l=150000u
+  ad=3.328e+11p pd=2.77e+06u as=7.85e+11p ps=3.57e+06u
M1002 a_669_111# a_639_85# a_1053_455# VPB pshort w=640000u l=150000u
+  ad=4.696e+11p pd=5.06e+06u as=1.536e+11p ps=1.76e+06u
M1003 VPWR a_1910_71# a_1890_508# VPB pshort w=420000u l=150000u
+  ad=2.66035e+12p pd=2.257e+07u as=1.176e+11p ps=1.4e+06u
M1004 VGND DE a_143_74# VNB nlowvt w=420000u l=150000u
+  ad=1.9208e+12p pd=1.749e+07u as=1.008e+11p ps=1.32e+06u
M1005 a_547_301# a_2385_74# VPWR VPB pshort w=640000u l=150000u
+  ad=1.76e+11p pd=1.83e+06u as=0p ps=0u
M1006 VGND a_2385_74# Q VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1007 a_1492_74# a_1295_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.072e+11p pd=2.04e+06u as=0p ps=0u
M1008 a_669_111# SCE a_27_74# VPB pshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_2274_392# a_1910_71# VPWR VPB pshort w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VGND DE a_159_404# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.197e+11p ps=1.41e+06u
M1011 VPWR a_2385_74# Q VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=3.08e+11p ps=2.79e+06u
M1012 a_505_111# a_159_404# VGND VNB nlowvt w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=0p ps=0u
M1013 a_554_463# DE VPWR VPB pshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_1890_508# a_1295_74# a_1688_97# VPB pshort w=420000u l=150000u
+  ad=0p pd=0u as=1.47e+11p ps=1.54e+06u
M1015 a_1688_97# a_1492_74# a_669_111# VPB pshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_1053_455# SCD VPWR VPB pshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_143_74# D a_27_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=2.982e+11p ps=3.1e+06u
M1018 a_1295_74# CLK VGND VNB nlowvt w=740000u l=150000u
+  ad=2.072e+11p pd=2.04e+06u as=0p ps=0u
M1019 a_547_301# a_2385_74# VGND VNB nlowvt w=420000u l=150000u
+  ad=1.197e+11p pd=1.41e+06u as=0p ps=0u
M1020 a_1295_74# CLK VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=3.08e+11p pd=2.79e+06u as=0p ps=0u
M1021 VPWR a_547_301# a_2568_508# VPB pshort w=420000u l=150000u
+  ad=0p pd=0u as=1.134e+11p ps=1.38e+06u
M1022 a_2313_74# a_1910_71# VGND VNB nlowvt w=640000u l=150000u
+  ad=1.344e+11p pd=1.7e+06u as=0p ps=0u
M1023 VPWR a_159_404# a_114_464# VPB pshort w=640000u l=150000u
+  ad=0p pd=0u as=1.536e+11p ps=1.76e+06u
M1024 a_2385_74# a_1492_74# a_2313_74# VNB nlowvt w=640000u l=150000u
+  ad=2.139e+11p pd=2e+06u as=0p ps=0u
M1025 a_669_111# a_639_85# a_27_74# VNB nlowvt w=420000u l=150000u
+  ad=3.843e+11p pd=4.35e+06u as=0p ps=0u
M1026 a_1688_97# a_1295_74# a_669_111# VNB nlowvt w=420000u l=150000u
+  ad=2.226e+11p pd=1.9e+06u as=0p ps=0u
M1027 VPWR SCE a_639_85# VPB pshort w=640000u l=150000u
+  ad=0p pd=0u as=1.792e+11p ps=1.84e+06u
M1028 a_669_111# SCE a_1026_125# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=8.82e+10p ps=1.26e+06u
M1029 VGND a_1910_71# a_1824_97# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.806e+11p ps=1.7e+06u
M1030 a_1492_74# a_1295_74# VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=3.08e+11p pd=2.79e+06u as=0p ps=0u
M1031 a_1026_125# SCD VGND VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1032 a_1824_97# a_1492_74# a_1688_97# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1033 a_1910_71# a_1688_97# VGND VNB nlowvt w=640000u l=150000u
+  ad=1.824e+11p pd=1.85e+06u as=0p ps=0u
M1034 a_2487_74# a_1295_74# a_2385_74# VNB nlowvt w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=0p ps=0u
M1035 VGND a_547_301# a_2487_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1036 VPWR DE a_159_404# VPB pshort w=640000u l=150000u
+  ad=0p pd=0u as=1.888e+11p ps=1.87e+06u
M1037 a_114_464# D a_27_74# VPB pshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1038 a_27_74# a_547_301# a_505_111# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1039 a_1910_71# a_1688_97# VPWR VPB pshort w=840000u l=150000u
+  ad=2.31e+11p pd=2.23e+06u as=0p ps=0u
M1040 a_2568_508# a_1492_74# a_2385_74# VPB pshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1041 VGND SCE a_639_85# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.176e+11p ps=1.4e+06u
.ends
