* File: sky130_fd_sc_hs__a311o_4.pxi.spice
* Created: Thu Aug 27 20:28:39 2020
* 
x_PM_SKY130_FD_SC_HS__A311O_4%C1 N_C1_c_142_n N_C1_M1006_g N_C1_M1014_g
+ N_C1_c_143_n N_C1_M1007_g N_C1_M1025_g C1 N_C1_c_141_n
+ PM_SKY130_FD_SC_HS__A311O_4%C1
x_PM_SKY130_FD_SC_HS__A311O_4%B1 N_B1_c_202_n N_B1_M1012_g N_B1_M1001_g
+ N_B1_c_203_n N_B1_M1018_g N_B1_M1023_g B1 N_B1_c_201_n
+ PM_SKY130_FD_SC_HS__A311O_4%B1
x_PM_SKY130_FD_SC_HS__A311O_4%A_154_392# N_A_154_392#_M1014_s
+ N_A_154_392#_M1001_s N_A_154_392#_M1004_d N_A_154_392#_M1006_d
+ N_A_154_392#_M1002_g N_A_154_392#_M1008_g N_A_154_392#_c_276_n
+ N_A_154_392#_M1000_g N_A_154_392#_M1015_g N_A_154_392#_c_277_n
+ N_A_154_392#_M1003_g N_A_154_392#_M1020_g N_A_154_392#_c_278_n
+ N_A_154_392#_M1026_g N_A_154_392#_c_264_n N_A_154_392#_c_265_n
+ N_A_154_392#_c_281_n N_A_154_392#_M1027_g N_A_154_392#_c_266_n
+ N_A_154_392#_c_267_n N_A_154_392#_c_268_n N_A_154_392#_c_269_n
+ N_A_154_392#_c_270_n N_A_154_392#_c_271_n N_A_154_392#_c_283_n
+ N_A_154_392#_c_284_n N_A_154_392#_c_361_p N_A_154_392#_c_272_n
+ N_A_154_392#_c_295_n N_A_154_392#_c_273_n N_A_154_392#_c_274_n
+ N_A_154_392#_c_324_p N_A_154_392#_c_275_n
+ PM_SKY130_FD_SC_HS__A311O_4%A_154_392#
x_PM_SKY130_FD_SC_HS__A311O_4%A3 N_A3_c_473_n N_A3_M1009_g N_A3_c_474_n
+ N_A3_c_475_n N_A3_c_476_n N_A3_M1011_g N_A3_c_478_n N_A3_M1013_g N_A3_c_479_n
+ N_A3_M1021_g A3 N_A3_c_477_n N_A3_c_481_n PM_SKY130_FD_SC_HS__A311O_4%A3
x_PM_SKY130_FD_SC_HS__A311O_4%A1 N_A1_c_542_n N_A1_M1022_g N_A1_M1004_g
+ N_A1_c_543_n N_A1_M1024_g N_A1_M1005_g A1 A1 A1 N_A1_c_541_n
+ PM_SKY130_FD_SC_HS__A311O_4%A1
x_PM_SKY130_FD_SC_HS__A311O_4%A2 N_A2_c_599_n N_A2_M1016_g N_A2_M1010_g
+ N_A2_M1019_g N_A2_c_600_n N_A2_M1017_g A2 N_A2_c_598_n
+ PM_SKY130_FD_SC_HS__A311O_4%A2
x_PM_SKY130_FD_SC_HS__A311O_4%A_69_392# N_A_69_392#_M1006_s N_A_69_392#_M1007_s
+ N_A_69_392#_M1018_s N_A_69_392#_c_636_n N_A_69_392#_c_637_n
+ N_A_69_392#_c_638_n N_A_69_392#_c_639_n PM_SKY130_FD_SC_HS__A311O_4%A_69_392#
x_PM_SKY130_FD_SC_HS__A311O_4%A_334_392# N_A_334_392#_M1012_d
+ N_A_334_392#_M1013_d N_A_334_392#_M1022_d N_A_334_392#_M1016_d
+ N_A_334_392#_c_674_n N_A_334_392#_c_692_n N_A_334_392#_c_675_n
+ N_A_334_392#_c_676_n N_A_334_392#_c_677_n N_A_334_392#_c_678_n
+ N_A_334_392#_c_679_n N_A_334_392#_c_682_n N_A_334_392#_c_680_n
+ N_A_334_392#_c_742_p PM_SKY130_FD_SC_HS__A311O_4%A_334_392#
x_PM_SKY130_FD_SC_HS__A311O_4%VPWR N_VPWR_M1000_s N_VPWR_M1003_s N_VPWR_M1027_s
+ N_VPWR_M1021_s N_VPWR_M1024_s N_VPWR_M1017_s N_VPWR_c_758_n N_VPWR_c_759_n
+ N_VPWR_c_760_n N_VPWR_c_761_n N_VPWR_c_762_n N_VPWR_c_763_n N_VPWR_c_764_n
+ N_VPWR_c_765_n N_VPWR_c_766_n VPWR N_VPWR_c_767_n N_VPWR_c_768_n
+ N_VPWR_c_769_n N_VPWR_c_770_n N_VPWR_c_771_n N_VPWR_c_772_n N_VPWR_c_773_n
+ N_VPWR_c_774_n N_VPWR_c_775_n N_VPWR_c_757_n PM_SKY130_FD_SC_HS__A311O_4%VPWR
x_PM_SKY130_FD_SC_HS__A311O_4%X N_X_M1002_s N_X_M1015_s N_X_M1000_d N_X_M1026_d
+ N_X_c_867_n N_X_c_875_n N_X_c_876_n N_X_c_888_n N_X_c_889_n N_X_c_877_n
+ N_X_c_878_n N_X_c_927_n N_X_c_868_n N_X_c_869_n N_X_c_879_n N_X_c_870_n
+ N_X_c_871_n N_X_c_906_n X N_X_c_872_n N_X_c_873_n
+ PM_SKY130_FD_SC_HS__A311O_4%X
x_PM_SKY130_FD_SC_HS__A311O_4%VGND N_VGND_M1014_d N_VGND_M1025_d N_VGND_M1023_d
+ N_VGND_M1008_d N_VGND_M1020_d N_VGND_M1011_s N_VGND_c_999_n N_VGND_c_1000_n
+ N_VGND_c_1001_n N_VGND_c_1002_n N_VGND_c_1003_n N_VGND_c_1004_n
+ N_VGND_c_1005_n N_VGND_c_1006_n N_VGND_c_1007_n N_VGND_c_1008_n
+ N_VGND_c_1009_n N_VGND_c_1010_n N_VGND_c_1011_n VGND N_VGND_c_1012_n
+ N_VGND_c_1013_n N_VGND_c_1014_n N_VGND_c_1015_n N_VGND_c_1016_n
+ N_VGND_c_1017_n PM_SKY130_FD_SC_HS__A311O_4%VGND
x_PM_SKY130_FD_SC_HS__A311O_4%A_888_105# N_A_888_105#_M1009_d
+ N_A_888_105#_M1010_s N_A_888_105#_c_1106_n N_A_888_105#_c_1115_n
+ N_A_888_105#_c_1107_n PM_SKY130_FD_SC_HS__A311O_4%A_888_105#
x_PM_SKY130_FD_SC_HS__A311O_4%A_1081_39# N_A_1081_39#_M1004_s
+ N_A_1081_39#_M1005_s N_A_1081_39#_M1019_d N_A_1081_39#_c_1136_n
+ N_A_1081_39#_c_1137_n N_A_1081_39#_c_1138_n N_A_1081_39#_c_1139_n
+ PM_SKY130_FD_SC_HS__A311O_4%A_1081_39#
cc_1 VNB N_C1_M1014_g 0.0351446f $X=-0.19 $Y=-0.245 $X2=0.775 $Y2=0.73
cc_2 VNB N_C1_M1025_g 0.0281669f $X=-0.19 $Y=-0.245 $X2=1.205 $Y2=0.73
cc_3 VNB C1 0.00185546f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_4 VNB N_C1_c_141_n 0.0414306f $X=-0.19 $Y=-0.245 $X2=1.145 $Y2=1.662
cc_5 VNB N_B1_M1001_g 0.0302599f $X=-0.19 $Y=-0.245 $X2=0.775 $Y2=0.73
cc_6 VNB N_B1_M1023_g 0.0303089f $X=-0.19 $Y=-0.245 $X2=1.205 $Y2=0.73
cc_7 VNB B1 7.52309e-19 $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_8 VNB N_B1_c_201_n 0.0234917f $X=-0.19 $Y=-0.245 $X2=1.145 $Y2=1.662
cc_9 VNB N_A_154_392#_M1002_g 0.0199403f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_10 VNB N_A_154_392#_M1008_g 0.0195521f $X=-0.19 $Y=-0.245 $X2=0.66 $Y2=1.635
cc_11 VNB N_A_154_392#_M1015_g 0.0188157f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_154_392#_M1020_g 0.0201088f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_154_392#_c_264_n 0.0136045f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_154_392#_c_265_n 0.0781868f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_154_392#_c_266_n 0.00349591f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_154_392#_c_267_n 0.00131296f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_154_392#_c_268_n 0.00811861f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_154_392#_c_269_n 0.00336243f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_154_392#_c_270_n 0.00800934f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_154_392#_c_271_n 0.00741641f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_154_392#_c_272_n 0.00604817f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_154_392#_c_273_n 0.00443304f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_154_392#_c_274_n 0.00348695f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_154_392#_c_275_n 0.00364225f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A3_c_473_n 0.0150962f $X=-0.19 $Y=-0.245 $X2=0.695 $Y2=1.885
cc_26 VNB N_A3_c_474_n 0.0137616f $X=-0.19 $Y=-0.245 $X2=0.775 $Y2=1.44
cc_27 VNB N_A3_c_475_n 0.00808421f $X=-0.19 $Y=-0.245 $X2=0.775 $Y2=0.73
cc_28 VNB N_A3_c_476_n 0.0187447f $X=-0.19 $Y=-0.245 $X2=0.775 $Y2=0.73
cc_29 VNB N_A3_c_477_n 0.0576105f $X=-0.19 $Y=-0.245 $X2=0.695 $Y2=1.662
cc_30 VNB N_A1_M1004_g 0.0264016f $X=-0.19 $Y=-0.245 $X2=0.775 $Y2=0.73
cc_31 VNB N_A1_M1005_g 0.0229491f $X=-0.19 $Y=-0.245 $X2=1.205 $Y2=0.73
cc_32 VNB A1 0.0023816f $X=-0.19 $Y=-0.245 $X2=0.66 $Y2=1.662
cc_33 VNB N_A1_c_541_n 0.0271077f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A2_M1010_g 0.0228767f $X=-0.19 $Y=-0.245 $X2=0.775 $Y2=0.73
cc_35 VNB N_A2_M1019_g 0.0283746f $X=-0.19 $Y=-0.245 $X2=1.145 $Y2=2.46
cc_36 VNB A2 0.00431308f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_37 VNB N_A2_c_598_n 0.0477483f $X=-0.19 $Y=-0.245 $X2=0.695 $Y2=1.662
cc_38 VNB N_VPWR_c_757_n 0.322901f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_X_c_867_n 0.0311159f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_X_c_868_n 0.00123375f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_X_c_869_n 0.00225295f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_X_c_870_n 0.00237374f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_X_c_871_n 0.0254155f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_X_c_872_n 0.0025697f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_X_c_873_n 0.0105207f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_VGND_c_999_n 0.0209749f $X=-0.19 $Y=-0.245 $X2=0.775 $Y2=1.662
cc_47 VNB N_VGND_c_1000_n 0.00367233f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_VGND_c_1001_n 0.0155164f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_VGND_c_1002_n 0.00680981f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_VGND_c_1003_n 0.0205594f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_VGND_c_1004_n 0.0101167f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_VGND_c_1005_n 0.0106292f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_VGND_c_1006_n 0.00119403f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_VGND_c_1007_n 0.0101383f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_VGND_c_1008_n 0.014713f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_VGND_c_1009_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_VGND_c_1010_n 0.0155164f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_VGND_c_1011_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_VGND_c_1012_n 0.0176086f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_VGND_c_1013_n 0.0884208f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_VGND_c_1014_n 0.452843f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_VGND_c_1015_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_VGND_c_1016_n 0.00413547f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_VGND_c_1017_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_A_888_105#_c_1106_n 0.0030352f $X=-0.19 $Y=-0.245 $X2=1.205 $Y2=0.73
cc_66 VNB N_A_888_105#_c_1107_n 0.00828173f $X=-0.19 $Y=-0.245 $X2=0.635
+ $Y2=1.58
cc_67 VNB N_A_1081_39#_c_1136_n 0.0519611f $X=-0.19 $Y=-0.245 $X2=1.145 $Y2=2.46
cc_68 VNB N_A_1081_39#_c_1137_n 0.00591587f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_A_1081_39#_c_1138_n 0.0126892f $X=-0.19 $Y=-0.245 $X2=0.66 $Y2=1.635
cc_70 VNB N_A_1081_39#_c_1139_n 0.024407f $X=-0.19 $Y=-0.245 $X2=0.775 $Y2=1.662
cc_71 VPB N_C1_c_142_n 0.0194199f $X=-0.19 $Y=1.66 $X2=0.695 $Y2=1.885
cc_72 VPB N_C1_c_143_n 0.0149839f $X=-0.19 $Y=1.66 $X2=1.145 $Y2=1.885
cc_73 VPB C1 0.00136459f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_74 VPB N_C1_c_141_n 0.0397788f $X=-0.19 $Y=1.66 $X2=1.145 $Y2=1.662
cc_75 VPB N_B1_c_202_n 0.0149109f $X=-0.19 $Y=1.66 $X2=0.695 $Y2=1.885
cc_76 VPB N_B1_c_203_n 0.0172189f $X=-0.19 $Y=1.66 $X2=1.145 $Y2=1.885
cc_77 VPB B1 0.00166024f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_78 VPB N_B1_c_201_n 0.0359908f $X=-0.19 $Y=1.66 $X2=1.145 $Y2=1.662
cc_79 VPB N_A_154_392#_c_276_n 0.018629f $X=-0.19 $Y=1.66 $X2=0.775 $Y2=1.662
cc_80 VPB N_A_154_392#_c_277_n 0.0149083f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_81 VPB N_A_154_392#_c_278_n 0.0149054f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_82 VPB N_A_154_392#_c_264_n 0.0135719f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_83 VPB N_A_154_392#_c_265_n 0.0465105f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_84 VPB N_A_154_392#_c_281_n 0.0155384f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_85 VPB N_A_154_392#_c_267_n 0.00158972f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_86 VPB N_A_154_392#_c_283_n 0.00306022f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_87 VPB N_A_154_392#_c_284_n 0.00722363f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_88 VPB N_A_154_392#_c_272_n 0.00238634f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_89 VPB N_A3_c_478_n 0.0161867f $X=-0.19 $Y=1.66 $X2=1.145 $Y2=2.46
cc_90 VPB N_A3_c_479_n 0.0157503f $X=-0.19 $Y=1.66 $X2=1.205 $Y2=0.73
cc_91 VPB N_A3_c_477_n 0.0337624f $X=-0.19 $Y=1.66 $X2=0.695 $Y2=1.662
cc_92 VPB N_A3_c_481_n 0.0025127f $X=-0.19 $Y=1.66 $X2=0.775 $Y2=1.662
cc_93 VPB N_A1_c_542_n 0.0147747f $X=-0.19 $Y=1.66 $X2=0.695 $Y2=1.885
cc_94 VPB N_A1_c_543_n 0.0153032f $X=-0.19 $Y=1.66 $X2=1.145 $Y2=1.885
cc_95 VPB A1 0.0019514f $X=-0.19 $Y=1.66 $X2=0.66 $Y2=1.662
cc_96 VPB N_A1_c_541_n 0.0339884f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_97 VPB N_A2_c_599_n 0.015326f $X=-0.19 $Y=1.66 $X2=0.695 $Y2=1.885
cc_98 VPB N_A2_c_600_n 0.0188935f $X=-0.19 $Y=1.66 $X2=1.205 $Y2=0.73
cc_99 VPB A2 0.0037002f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_100 VPB N_A2_c_598_n 0.0542196f $X=-0.19 $Y=1.66 $X2=0.695 $Y2=1.662
cc_101 VPB N_A_69_392#_c_636_n 0.00213603f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_102 VPB N_A_69_392#_c_637_n 0.0173694f $X=-0.19 $Y=1.66 $X2=0.66 $Y2=1.635
cc_103 VPB N_A_69_392#_c_638_n 0.00216539f $X=-0.19 $Y=1.66 $X2=0.66 $Y2=1.635
cc_104 VPB N_A_69_392#_c_639_n 0.00675527f $X=-0.19 $Y=1.66 $X2=0.775 $Y2=1.662
cc_105 VPB N_A_334_392#_c_674_n 0.00781107f $X=-0.19 $Y=1.66 $X2=1.205 $Y2=0.73
cc_106 VPB N_A_334_392#_c_675_n 0.00110023f $X=-0.19 $Y=1.66 $X2=0.66 $Y2=1.635
cc_107 VPB N_A_334_392#_c_676_n 0.00180921f $X=-0.19 $Y=1.66 $X2=1.205 $Y2=1.662
cc_108 VPB N_A_334_392#_c_677_n 0.0034066f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_109 VPB N_A_334_392#_c_678_n 0.00110611f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_110 VPB N_A_334_392#_c_679_n 0.00180921f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_111 VPB N_A_334_392#_c_680_n 0.00257417f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_112 VPB N_VPWR_c_758_n 0.00881729f $X=-0.19 $Y=1.66 $X2=0.775 $Y2=1.662
cc_113 VPB N_VPWR_c_759_n 0.0177589f $X=-0.19 $Y=1.66 $X2=1.205 $Y2=1.662
cc_114 VPB N_VPWR_c_760_n 0.00261791f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_115 VPB N_VPWR_c_761_n 0.00591026f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_116 VPB N_VPWR_c_762_n 0.0201268f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_117 VPB N_VPWR_c_763_n 0.00504372f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_118 VPB N_VPWR_c_764_n 0.00261791f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_119 VPB N_VPWR_c_765_n 0.0124891f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_120 VPB N_VPWR_c_766_n 0.0504568f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_121 VPB N_VPWR_c_767_n 0.0667191f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_122 VPB N_VPWR_c_768_n 0.0177589f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_123 VPB N_VPWR_c_769_n 0.0164465f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_124 VPB N_VPWR_c_770_n 0.0164465f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_125 VPB N_VPWR_c_771_n 0.00614127f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_126 VPB N_VPWR_c_772_n 0.00601644f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_127 VPB N_VPWR_c_773_n 0.00614127f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_128 VPB N_VPWR_c_774_n 0.00460249f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_129 VPB N_VPWR_c_775_n 0.00656574f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_130 VPB N_VPWR_c_757_n 0.0895347f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_131 VPB N_X_c_867_n 0.0350668f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_132 VPB N_X_c_875_n 0.00248381f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_133 VPB N_X_c_876_n 0.0113009f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_134 VPB N_X_c_877_n 0.00612414f $X=-0.19 $Y=1.66 $X2=0.775 $Y2=1.662
cc_135 VPB N_X_c_878_n 0.00677331f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_136 VPB N_X_c_879_n 0.00328209f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_137 N_C1_c_143_n N_B1_c_202_n 0.0316207f $X=1.145 $Y=1.885 $X2=-0.19
+ $Y2=-0.245
cc_138 N_C1_M1025_g N_B1_M1001_g 0.0247525f $X=1.205 $Y=0.73 $X2=0 $Y2=0
cc_139 N_C1_c_141_n B1 0.00142809f $X=1.145 $Y=1.662 $X2=0 $Y2=0
cc_140 N_C1_c_141_n N_B1_c_201_n 0.0225347f $X=1.145 $Y=1.662 $X2=0 $Y2=0
cc_141 N_C1_M1014_g N_A_154_392#_c_266_n 0.00158318f $X=0.775 $Y=0.73 $X2=0
+ $Y2=0
cc_142 N_C1_M1025_g N_A_154_392#_c_266_n 0.00145882f $X=1.205 $Y=0.73 $X2=0
+ $Y2=0
cc_143 N_C1_c_142_n N_A_154_392#_c_267_n 0.00244283f $X=0.695 $Y=1.885 $X2=0
+ $Y2=0
cc_144 N_C1_M1014_g N_A_154_392#_c_267_n 0.00296395f $X=0.775 $Y=0.73 $X2=0
+ $Y2=0
cc_145 N_C1_c_143_n N_A_154_392#_c_267_n 0.00335997f $X=1.145 $Y=1.885 $X2=0
+ $Y2=0
cc_146 N_C1_M1025_g N_A_154_392#_c_267_n 0.00344202f $X=1.205 $Y=0.73 $X2=0
+ $Y2=0
cc_147 C1 N_A_154_392#_c_267_n 0.023546f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_148 N_C1_c_141_n N_A_154_392#_c_267_n 0.0221656f $X=1.145 $Y=1.662 $X2=0
+ $Y2=0
cc_149 N_C1_M1025_g N_A_154_392#_c_268_n 0.010261f $X=1.205 $Y=0.73 $X2=0 $Y2=0
cc_150 N_C1_c_142_n N_A_154_392#_c_295_n 0.00331218f $X=0.695 $Y=1.885 $X2=0
+ $Y2=0
cc_151 N_C1_c_143_n N_A_154_392#_c_295_n 0.00405177f $X=1.145 $Y=1.885 $X2=0
+ $Y2=0
cc_152 C1 N_A_154_392#_c_295_n 0.00252338f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_153 N_C1_c_141_n N_A_154_392#_c_295_n 0.00766578f $X=1.145 $Y=1.662 $X2=0
+ $Y2=0
cc_154 N_C1_M1014_g N_A_154_392#_c_273_n 0.00266773f $X=0.775 $Y=0.73 $X2=0
+ $Y2=0
cc_155 N_C1_M1025_g N_A_154_392#_c_273_n 0.00272436f $X=1.205 $Y=0.73 $X2=0
+ $Y2=0
cc_156 N_C1_c_141_n N_A_154_392#_c_273_n 0.00254808f $X=1.145 $Y=1.662 $X2=0
+ $Y2=0
cc_157 N_C1_c_142_n N_A_69_392#_c_637_n 0.0113574f $X=0.695 $Y=1.885 $X2=0 $Y2=0
cc_158 N_C1_c_143_n N_A_69_392#_c_637_n 0.0102143f $X=1.145 $Y=1.885 $X2=0 $Y2=0
cc_159 N_C1_c_142_n N_A_69_392#_c_638_n 4.4235e-19 $X=0.695 $Y=1.885 $X2=0 $Y2=0
cc_160 N_C1_c_143_n N_A_69_392#_c_638_n 0.00386766f $X=1.145 $Y=1.885 $X2=0
+ $Y2=0
cc_161 N_C1_c_142_n N_VPWR_c_767_n 0.00291649f $X=0.695 $Y=1.885 $X2=0 $Y2=0
cc_162 N_C1_c_143_n N_VPWR_c_767_n 0.00290311f $X=1.145 $Y=1.885 $X2=0 $Y2=0
cc_163 N_C1_c_142_n N_VPWR_c_757_n 0.0036349f $X=0.695 $Y=1.885 $X2=0 $Y2=0
cc_164 N_C1_c_143_n N_VPWR_c_757_n 0.0035903f $X=1.145 $Y=1.885 $X2=0 $Y2=0
cc_165 N_C1_c_142_n N_X_c_867_n 0.0119542f $X=0.695 $Y=1.885 $X2=0 $Y2=0
cc_166 N_C1_M1014_g N_X_c_867_n 0.00828409f $X=0.775 $Y=0.73 $X2=0 $Y2=0
cc_167 C1 N_X_c_867_n 0.0219102f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_168 N_C1_c_141_n N_X_c_867_n 0.00600948f $X=1.145 $Y=1.662 $X2=0 $Y2=0
cc_169 N_C1_c_142_n N_X_c_875_n 0.0140796f $X=0.695 $Y=1.885 $X2=0 $Y2=0
cc_170 N_C1_c_143_n N_X_c_875_n 0.0120487f $X=1.145 $Y=1.885 $X2=0 $Y2=0
cc_171 C1 N_X_c_875_n 0.00639388f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_172 N_C1_c_141_n N_X_c_875_n 0.00172654f $X=1.145 $Y=1.662 $X2=0 $Y2=0
cc_173 N_C1_c_143_n N_X_c_888_n 0.00411697f $X=1.145 $Y=1.885 $X2=0 $Y2=0
cc_174 N_C1_c_143_n N_X_c_889_n 0.00127332f $X=1.145 $Y=1.885 $X2=0 $Y2=0
cc_175 N_C1_M1014_g N_X_c_870_n 0.0106431f $X=0.775 $Y=0.73 $X2=0 $Y2=0
cc_176 N_C1_M1025_g N_X_c_870_n 0.00641472f $X=1.205 $Y=0.73 $X2=0 $Y2=0
cc_177 C1 N_X_c_870_n 0.0103097f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_178 N_C1_c_141_n N_X_c_870_n 0.00451519f $X=1.145 $Y=1.662 $X2=0 $Y2=0
cc_179 N_C1_M1014_g N_X_c_871_n 0.001969f $X=0.775 $Y=0.73 $X2=0 $Y2=0
cc_180 N_C1_M1014_g N_X_c_873_n 0.00338785f $X=0.775 $Y=0.73 $X2=0 $Y2=0
cc_181 N_C1_M1014_g N_VGND_c_999_n 0.00806526f $X=0.775 $Y=0.73 $X2=0 $Y2=0
cc_182 N_C1_M1025_g N_VGND_c_999_n 3.98426e-19 $X=1.205 $Y=0.73 $X2=0 $Y2=0
cc_183 N_C1_M1014_g N_VGND_c_1000_n 5.23778e-19 $X=0.775 $Y=0.73 $X2=0 $Y2=0
cc_184 N_C1_M1025_g N_VGND_c_1000_n 0.00953485f $X=1.205 $Y=0.73 $X2=0 $Y2=0
cc_185 N_C1_M1014_g N_VGND_c_1010_n 0.00455951f $X=0.775 $Y=0.73 $X2=0 $Y2=0
cc_186 N_C1_M1025_g N_VGND_c_1010_n 0.00455951f $X=1.205 $Y=0.73 $X2=0 $Y2=0
cc_187 N_C1_M1014_g N_VGND_c_1014_n 0.00447788f $X=0.775 $Y=0.73 $X2=0 $Y2=0
cc_188 N_C1_M1025_g N_VGND_c_1014_n 0.00447788f $X=1.205 $Y=0.73 $X2=0 $Y2=0
cc_189 N_B1_M1023_g N_A_154_392#_M1002_g 0.0163992f $X=2.065 $Y=0.73 $X2=0 $Y2=0
cc_190 B1 N_A_154_392#_c_265_n 5.44412e-19 $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_191 N_B1_c_201_n N_A_154_392#_c_265_n 0.0224918f $X=2.045 $Y=1.677 $X2=0
+ $Y2=0
cc_192 N_B1_c_202_n N_A_154_392#_c_267_n 5.14028e-19 $X=1.595 $Y=1.885 $X2=0
+ $Y2=0
cc_193 N_B1_M1001_g N_A_154_392#_c_267_n 8.44792e-19 $X=1.635 $Y=0.73 $X2=0
+ $Y2=0
cc_194 B1 N_A_154_392#_c_267_n 0.0126148f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_195 N_B1_c_201_n N_A_154_392#_c_267_n 0.00172234f $X=2.045 $Y=1.677 $X2=0
+ $Y2=0
cc_196 N_B1_M1001_g N_A_154_392#_c_268_n 0.0105611f $X=1.635 $Y=0.73 $X2=0 $Y2=0
cc_197 B1 N_A_154_392#_c_268_n 0.0153097f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_198 N_B1_c_201_n N_A_154_392#_c_268_n 0.00109394f $X=2.045 $Y=1.677 $X2=0
+ $Y2=0
cc_199 N_B1_M1001_g N_A_154_392#_c_269_n 0.00145882f $X=1.635 $Y=0.73 $X2=0
+ $Y2=0
cc_200 N_B1_M1023_g N_A_154_392#_c_269_n 0.00137192f $X=2.065 $Y=0.73 $X2=0
+ $Y2=0
cc_201 N_B1_M1001_g N_A_154_392#_c_270_n 9.18327e-19 $X=1.635 $Y=0.73 $X2=0
+ $Y2=0
cc_202 N_B1_M1023_g N_A_154_392#_c_270_n 0.0164591f $X=2.065 $Y=0.73 $X2=0 $Y2=0
cc_203 B1 N_A_154_392#_c_270_n 0.0220632f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_204 N_B1_c_201_n N_A_154_392#_c_270_n 0.00982479f $X=2.045 $Y=1.677 $X2=0
+ $Y2=0
cc_205 N_B1_c_202_n N_A_69_392#_c_636_n 0.0108414f $X=1.595 $Y=1.885 $X2=0 $Y2=0
cc_206 N_B1_c_203_n N_A_69_392#_c_636_n 0.00848139f $X=2.045 $Y=1.885 $X2=0
+ $Y2=0
cc_207 N_B1_c_202_n N_A_69_392#_c_638_n 0.00542024f $X=1.595 $Y=1.885 $X2=0
+ $Y2=0
cc_208 N_B1_c_203_n N_A_69_392#_c_638_n 5.10463e-19 $X=2.045 $Y=1.885 $X2=0
+ $Y2=0
cc_209 N_B1_c_202_n N_A_69_392#_c_639_n 6.04816e-19 $X=1.595 $Y=1.885 $X2=0
+ $Y2=0
cc_210 N_B1_c_203_n N_A_69_392#_c_639_n 0.00703734f $X=2.045 $Y=1.885 $X2=0
+ $Y2=0
cc_211 N_B1_c_203_n N_A_334_392#_c_674_n 0.011674f $X=2.045 $Y=1.885 $X2=0 $Y2=0
cc_212 N_B1_c_202_n N_A_334_392#_c_682_n 0.00436919f $X=1.595 $Y=1.885 $X2=0
+ $Y2=0
cc_213 N_B1_c_203_n N_A_334_392#_c_682_n 0.00392125f $X=2.045 $Y=1.885 $X2=0
+ $Y2=0
cc_214 N_B1_c_203_n N_VPWR_c_758_n 0.00123892f $X=2.045 $Y=1.885 $X2=0 $Y2=0
cc_215 N_B1_c_202_n N_VPWR_c_767_n 0.00278271f $X=1.595 $Y=1.885 $X2=0 $Y2=0
cc_216 N_B1_c_203_n N_VPWR_c_767_n 0.00279479f $X=2.045 $Y=1.885 $X2=0 $Y2=0
cc_217 N_B1_c_202_n N_VPWR_c_757_n 0.00353907f $X=1.595 $Y=1.885 $X2=0 $Y2=0
cc_218 N_B1_c_203_n N_VPWR_c_757_n 0.00357714f $X=2.045 $Y=1.885 $X2=0 $Y2=0
cc_219 N_B1_c_203_n N_X_c_877_n 0.00300008f $X=2.045 $Y=1.885 $X2=0 $Y2=0
cc_220 N_B1_c_201_n N_X_c_877_n 0.00212015f $X=2.045 $Y=1.677 $X2=0 $Y2=0
cc_221 N_B1_M1023_g N_X_c_868_n 5.77553e-19 $X=2.065 $Y=0.73 $X2=0 $Y2=0
cc_222 N_B1_c_202_n N_X_c_879_n 0.014561f $X=1.595 $Y=1.885 $X2=0 $Y2=0
cc_223 N_B1_c_203_n N_X_c_879_n 0.0143156f $X=2.045 $Y=1.885 $X2=0 $Y2=0
cc_224 B1 N_X_c_879_n 0.0219372f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_225 N_B1_c_201_n N_X_c_879_n 0.00356511f $X=2.045 $Y=1.677 $X2=0 $Y2=0
cc_226 N_B1_M1001_g N_X_c_870_n 0.00641498f $X=1.635 $Y=0.73 $X2=0 $Y2=0
cc_227 N_B1_M1023_g N_X_c_870_n 0.00645808f $X=2.065 $Y=0.73 $X2=0 $Y2=0
cc_228 B1 N_X_c_870_n 4.24688e-19 $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_229 N_B1_M1023_g N_X_c_906_n 2.2693e-19 $X=2.065 $Y=0.73 $X2=0 $Y2=0
cc_230 N_B1_M1023_g N_X_c_872_n 3.3543e-19 $X=2.065 $Y=0.73 $X2=0 $Y2=0
cc_231 N_B1_M1001_g N_VGND_c_1000_n 0.00953485f $X=1.635 $Y=0.73 $X2=0 $Y2=0
cc_232 N_B1_M1023_g N_VGND_c_1000_n 5.23778e-19 $X=2.065 $Y=0.73 $X2=0 $Y2=0
cc_233 N_B1_M1001_g N_VGND_c_1001_n 0.00455951f $X=1.635 $Y=0.73 $X2=0 $Y2=0
cc_234 N_B1_M1023_g N_VGND_c_1001_n 0.00455951f $X=2.065 $Y=0.73 $X2=0 $Y2=0
cc_235 N_B1_M1001_g N_VGND_c_1002_n 5.34522e-19 $X=1.635 $Y=0.73 $X2=0 $Y2=0
cc_236 N_B1_M1023_g N_VGND_c_1002_n 0.0113902f $X=2.065 $Y=0.73 $X2=0 $Y2=0
cc_237 N_B1_M1001_g N_VGND_c_1014_n 0.00447788f $X=1.635 $Y=0.73 $X2=0 $Y2=0
cc_238 N_B1_M1023_g N_VGND_c_1014_n 0.00447788f $X=2.065 $Y=0.73 $X2=0 $Y2=0
cc_239 N_A_154_392#_M1020_g N_A3_c_473_n 0.0189143f $X=3.875 $Y=0.795 $X2=-0.19
+ $Y2=-0.245
cc_240 N_A_154_392#_c_271_n N_A3_c_474_n 0.00466849f $X=4.475 $Y=1.565 $X2=0
+ $Y2=0
cc_241 N_A_154_392#_c_284_n N_A3_c_474_n 0.00204554f $X=5.545 $Y=2.035 $X2=0
+ $Y2=0
cc_242 N_A_154_392#_c_264_n N_A3_c_475_n 0.0108244f $X=4.275 $Y=1.675 $X2=0
+ $Y2=0
cc_243 N_A_154_392#_c_265_n N_A3_c_475_n 0.00390388f $X=4.005 $Y=1.675 $X2=0
+ $Y2=0
cc_244 N_A_154_392#_c_271_n N_A3_c_475_n 0.00201387f $X=4.475 $Y=1.565 $X2=0
+ $Y2=0
cc_245 N_A_154_392#_c_324_p N_A3_c_475_n 4.05596e-19 $X=3.905 $Y=1.485 $X2=0
+ $Y2=0
cc_246 N_A_154_392#_c_275_n N_A3_c_476_n 0.00259763f $X=6.02 $Y=1.1 $X2=0 $Y2=0
cc_247 N_A_154_392#_c_281_n N_A3_c_478_n 0.0312898f $X=4.365 $Y=1.765 $X2=0
+ $Y2=0
cc_248 N_A_154_392#_c_283_n N_A3_c_478_n 0.00139691f $X=4.56 $Y=1.95 $X2=0 $Y2=0
cc_249 N_A_154_392#_c_284_n N_A3_c_478_n 0.0144443f $X=5.545 $Y=2.035 $X2=0
+ $Y2=0
cc_250 N_A_154_392#_c_284_n N_A3_c_479_n 0.0137942f $X=5.545 $Y=2.035 $X2=0
+ $Y2=0
cc_251 N_A_154_392#_c_272_n N_A3_c_479_n 0.00138745f $X=5.63 $Y=1.95 $X2=0 $Y2=0
cc_252 N_A_154_392#_c_264_n N_A3_c_477_n 0.00559634f $X=4.275 $Y=1.675 $X2=0
+ $Y2=0
cc_253 N_A_154_392#_c_265_n N_A3_c_477_n 0.00320654f $X=4.005 $Y=1.675 $X2=0
+ $Y2=0
cc_254 N_A_154_392#_c_281_n N_A3_c_477_n 0.00308894f $X=4.365 $Y=1.765 $X2=0
+ $Y2=0
cc_255 N_A_154_392#_c_271_n N_A3_c_477_n 0.00304129f $X=4.475 $Y=1.565 $X2=0
+ $Y2=0
cc_256 N_A_154_392#_c_283_n N_A3_c_477_n 0.00351887f $X=4.56 $Y=1.95 $X2=0 $Y2=0
cc_257 N_A_154_392#_c_284_n N_A3_c_477_n 0.0062513f $X=5.545 $Y=2.035 $X2=0
+ $Y2=0
cc_258 N_A_154_392#_c_272_n N_A3_c_477_n 0.0089252f $X=5.63 $Y=1.95 $X2=0 $Y2=0
cc_259 N_A_154_392#_c_271_n N_A3_c_481_n 0.009987f $X=4.475 $Y=1.565 $X2=0 $Y2=0
cc_260 N_A_154_392#_c_283_n N_A3_c_481_n 0.00672864f $X=4.56 $Y=1.95 $X2=0 $Y2=0
cc_261 N_A_154_392#_c_284_n N_A3_c_481_n 0.028856f $X=5.545 $Y=2.035 $X2=0 $Y2=0
cc_262 N_A_154_392#_c_272_n N_A3_c_481_n 0.0204032f $X=5.63 $Y=1.95 $X2=0 $Y2=0
cc_263 N_A_154_392#_c_284_n N_A1_c_542_n 0.00391862f $X=5.545 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_264 N_A_154_392#_c_272_n N_A1_c_542_n 0.00153688f $X=5.63 $Y=1.95 $X2=-0.19
+ $Y2=-0.245
cc_265 N_A_154_392#_c_272_n N_A1_M1004_g 0.00704871f $X=5.63 $Y=1.95 $X2=0 $Y2=0
cc_266 N_A_154_392#_c_275_n N_A1_M1004_g 0.0200901f $X=6.02 $Y=1.1 $X2=0 $Y2=0
cc_267 N_A_154_392#_c_272_n N_A1_c_543_n 3.01255e-19 $X=5.63 $Y=1.95 $X2=0 $Y2=0
cc_268 N_A_154_392#_c_275_n N_A1_M1005_g 7.51231e-19 $X=6.02 $Y=1.1 $X2=0 $Y2=0
cc_269 N_A_154_392#_c_272_n A1 0.0249855f $X=5.63 $Y=1.95 $X2=0 $Y2=0
cc_270 N_A_154_392#_c_275_n A1 0.0163424f $X=6.02 $Y=1.1 $X2=0 $Y2=0
cc_271 N_A_154_392#_c_272_n N_A1_c_541_n 0.0113411f $X=5.63 $Y=1.95 $X2=0 $Y2=0
cc_272 N_A_154_392#_c_275_n N_A1_c_541_n 0.00306703f $X=6.02 $Y=1.1 $X2=0 $Y2=0
cc_273 N_A_154_392#_M1006_d N_A_69_392#_c_637_n 0.00201274f $X=0.77 $Y=1.96
+ $X2=0 $Y2=0
cc_274 N_A_154_392#_c_276_n N_A_69_392#_c_639_n 8.99459e-19 $X=3.015 $Y=1.765
+ $X2=0 $Y2=0
cc_275 N_A_154_392#_c_284_n N_A_334_392#_M1013_d 0.00197722f $X=5.545 $Y=2.035
+ $X2=0 $Y2=0
cc_276 N_A_154_392#_c_276_n N_A_334_392#_c_674_n 0.0139319f $X=3.015 $Y=1.765
+ $X2=0 $Y2=0
cc_277 N_A_154_392#_c_277_n N_A_334_392#_c_674_n 0.0120114f $X=3.465 $Y=1.765
+ $X2=0 $Y2=0
cc_278 N_A_154_392#_c_278_n N_A_334_392#_c_674_n 0.0120114f $X=3.915 $Y=1.765
+ $X2=0 $Y2=0
cc_279 N_A_154_392#_c_281_n N_A_334_392#_c_674_n 0.0143473f $X=4.365 $Y=1.765
+ $X2=0 $Y2=0
cc_280 N_A_154_392#_c_271_n N_A_334_392#_c_674_n 0.00334363f $X=4.475 $Y=1.565
+ $X2=0 $Y2=0
cc_281 N_A_154_392#_c_284_n N_A_334_392#_c_674_n 0.0146046f $X=5.545 $Y=2.035
+ $X2=0 $Y2=0
cc_282 N_A_154_392#_c_361_p N_A_334_392#_c_674_n 0.0105753f $X=4.645 $Y=2.035
+ $X2=0 $Y2=0
cc_283 N_A_154_392#_c_284_n N_A_334_392#_c_692_n 0.0242083f $X=5.545 $Y=2.035
+ $X2=0 $Y2=0
cc_284 N_A_154_392#_c_284_n N_A_334_392#_c_675_n 0.012862f $X=5.545 $Y=2.035
+ $X2=0 $Y2=0
cc_285 N_A_154_392#_c_281_n N_A_334_392#_c_680_n 6.92625e-19 $X=4.365 $Y=1.765
+ $X2=0 $Y2=0
cc_286 N_A_154_392#_c_284_n N_A_334_392#_c_680_n 0.0173542f $X=5.545 $Y=2.035
+ $X2=0 $Y2=0
cc_287 N_A_154_392#_c_283_n N_VPWR_M1027_s 0.00202354f $X=4.56 $Y=1.95 $X2=0
+ $Y2=0
cc_288 N_A_154_392#_c_284_n N_VPWR_M1027_s 0.00228433f $X=5.545 $Y=2.035 $X2=0
+ $Y2=0
cc_289 N_A_154_392#_c_361_p N_VPWR_M1027_s 0.0029504f $X=4.645 $Y=2.035 $X2=0
+ $Y2=0
cc_290 N_A_154_392#_c_284_n N_VPWR_M1021_s 0.00201643f $X=5.545 $Y=2.035 $X2=0
+ $Y2=0
cc_291 N_A_154_392#_c_276_n N_VPWR_c_758_n 0.0106215f $X=3.015 $Y=1.765 $X2=0
+ $Y2=0
cc_292 N_A_154_392#_c_277_n N_VPWR_c_758_n 0.00127141f $X=3.465 $Y=1.765 $X2=0
+ $Y2=0
cc_293 N_A_154_392#_c_276_n N_VPWR_c_759_n 0.00413917f $X=3.015 $Y=1.765 $X2=0
+ $Y2=0
cc_294 N_A_154_392#_c_277_n N_VPWR_c_759_n 0.00413917f $X=3.465 $Y=1.765 $X2=0
+ $Y2=0
cc_295 N_A_154_392#_c_276_n N_VPWR_c_760_n 0.00127141f $X=3.015 $Y=1.765 $X2=0
+ $Y2=0
cc_296 N_A_154_392#_c_277_n N_VPWR_c_760_n 0.00963065f $X=3.465 $Y=1.765 $X2=0
+ $Y2=0
cc_297 N_A_154_392#_c_278_n N_VPWR_c_760_n 0.00963065f $X=3.915 $Y=1.765 $X2=0
+ $Y2=0
cc_298 N_A_154_392#_c_281_n N_VPWR_c_760_n 0.00127141f $X=4.365 $Y=1.765 $X2=0
+ $Y2=0
cc_299 N_A_154_392#_c_278_n N_VPWR_c_761_n 0.00127141f $X=3.915 $Y=1.765 $X2=0
+ $Y2=0
cc_300 N_A_154_392#_c_281_n N_VPWR_c_761_n 0.00960501f $X=4.365 $Y=1.765 $X2=0
+ $Y2=0
cc_301 N_A_154_392#_c_278_n N_VPWR_c_768_n 0.00413917f $X=3.915 $Y=1.765 $X2=0
+ $Y2=0
cc_302 N_A_154_392#_c_281_n N_VPWR_c_768_n 0.00413917f $X=4.365 $Y=1.765 $X2=0
+ $Y2=0
cc_303 N_A_154_392#_c_276_n N_VPWR_c_757_n 0.00414505f $X=3.015 $Y=1.765 $X2=0
+ $Y2=0
cc_304 N_A_154_392#_c_277_n N_VPWR_c_757_n 0.00414505f $X=3.465 $Y=1.765 $X2=0
+ $Y2=0
cc_305 N_A_154_392#_c_278_n N_VPWR_c_757_n 0.00414505f $X=3.915 $Y=1.765 $X2=0
+ $Y2=0
cc_306 N_A_154_392#_c_281_n N_VPWR_c_757_n 0.00414505f $X=4.365 $Y=1.765 $X2=0
+ $Y2=0
cc_307 N_A_154_392#_c_266_n N_X_c_867_n 0.00256949f $X=0.99 $Y=0.555 $X2=0 $Y2=0
cc_308 N_A_154_392#_c_295_n N_X_c_867_n 0.00608974f $X=1.08 $Y=2.105 $X2=0 $Y2=0
cc_309 N_A_154_392#_c_273_n N_X_c_867_n 0.00582022f $X=1.035 $Y=1.215 $X2=0
+ $Y2=0
cc_310 N_A_154_392#_M1006_d N_X_c_875_n 0.00374176f $X=0.77 $Y=1.96 $X2=0 $Y2=0
cc_311 N_A_154_392#_c_295_n N_X_c_875_n 0.020864f $X=1.08 $Y=2.105 $X2=0 $Y2=0
cc_312 N_A_154_392#_c_295_n N_X_c_888_n 0.0036619f $X=1.08 $Y=2.105 $X2=0 $Y2=0
cc_313 N_A_154_392#_c_267_n N_X_c_889_n 0.00394652f $X=1.08 $Y=2.02 $X2=0 $Y2=0
cc_314 N_A_154_392#_c_268_n N_X_c_889_n 0.00443876f $X=1.755 $Y=1.215 $X2=0
+ $Y2=0
cc_315 N_A_154_392#_c_295_n N_X_c_889_n 0.0100278f $X=1.08 $Y=2.105 $X2=0 $Y2=0
cc_316 N_A_154_392#_c_265_n N_X_c_877_n 0.0117314f $X=4.005 $Y=1.675 $X2=0 $Y2=0
cc_317 N_A_154_392#_c_274_n N_X_c_877_n 0.0686585f $X=3.74 $Y=1.485 $X2=0 $Y2=0
cc_318 N_A_154_392#_c_276_n N_X_c_878_n 0.0165629f $X=3.015 $Y=1.765 $X2=0 $Y2=0
cc_319 N_A_154_392#_c_277_n N_X_c_878_n 0.0131963f $X=3.465 $Y=1.765 $X2=0 $Y2=0
cc_320 N_A_154_392#_c_278_n N_X_c_878_n 0.0131963f $X=3.915 $Y=1.765 $X2=0 $Y2=0
cc_321 N_A_154_392#_c_264_n N_X_c_878_n 0.00623847f $X=4.275 $Y=1.675 $X2=0
+ $Y2=0
cc_322 N_A_154_392#_c_265_n N_X_c_878_n 0.0182271f $X=4.005 $Y=1.675 $X2=0 $Y2=0
cc_323 N_A_154_392#_c_281_n N_X_c_878_n 0.00406588f $X=4.365 $Y=1.765 $X2=0
+ $Y2=0
cc_324 N_A_154_392#_c_283_n N_X_c_878_n 0.00611407f $X=4.56 $Y=1.95 $X2=0 $Y2=0
cc_325 N_A_154_392#_c_324_p N_X_c_878_n 0.0686585f $X=3.905 $Y=1.485 $X2=0 $Y2=0
cc_326 N_A_154_392#_M1008_g N_X_c_927_n 0.0113003f $X=2.97 $Y=0.78 $X2=0 $Y2=0
cc_327 N_A_154_392#_M1015_g N_X_c_927_n 0.0121433f $X=3.445 $Y=0.795 $X2=0 $Y2=0
cc_328 N_A_154_392#_c_265_n N_X_c_927_n 0.00588912f $X=4.005 $Y=1.675 $X2=0
+ $Y2=0
cc_329 N_A_154_392#_c_274_n N_X_c_927_n 0.0554913f $X=3.74 $Y=1.485 $X2=0 $Y2=0
cc_330 N_A_154_392#_M1002_g N_X_c_868_n 0.00454864f $X=2.54 $Y=0.78 $X2=0 $Y2=0
cc_331 N_A_154_392#_M1008_g N_X_c_868_n 7.32094e-19 $X=2.97 $Y=0.78 $X2=0 $Y2=0
cc_332 N_A_154_392#_c_265_n N_X_c_868_n 0.0024556f $X=4.005 $Y=1.675 $X2=0 $Y2=0
cc_333 N_A_154_392#_c_269_n N_X_c_868_n 0.00293534f $X=1.85 $Y=0.555 $X2=0 $Y2=0
cc_334 N_A_154_392#_c_270_n N_X_c_868_n 0.00148317f $X=2.325 $Y=1.485 $X2=0
+ $Y2=0
cc_335 N_A_154_392#_c_274_n N_X_c_868_n 0.0249499f $X=3.74 $Y=1.485 $X2=0 $Y2=0
cc_336 N_A_154_392#_M1008_g N_X_c_869_n 6.24169e-19 $X=2.97 $Y=0.78 $X2=0 $Y2=0
cc_337 N_A_154_392#_M1015_g N_X_c_869_n 0.00799917f $X=3.445 $Y=0.795 $X2=0
+ $Y2=0
cc_338 N_A_154_392#_M1020_g N_X_c_869_n 2.50179e-19 $X=3.875 $Y=0.795 $X2=0
+ $Y2=0
cc_339 N_A_154_392#_c_265_n N_X_c_879_n 0.00158201f $X=4.005 $Y=1.675 $X2=0
+ $Y2=0
cc_340 N_A_154_392#_c_268_n N_X_c_879_n 6.12642e-19 $X=1.755 $Y=1.215 $X2=0
+ $Y2=0
cc_341 N_A_154_392#_c_270_n N_X_c_879_n 0.0164441f $X=2.325 $Y=1.485 $X2=0 $Y2=0
cc_342 N_A_154_392#_c_274_n N_X_c_879_n 0.00982063f $X=3.74 $Y=1.485 $X2=0 $Y2=0
cc_343 N_A_154_392#_M1014_s N_X_c_870_n 0.00599498f $X=0.85 $Y=0.41 $X2=0 $Y2=0
cc_344 N_A_154_392#_M1001_s N_X_c_870_n 0.00438342f $X=1.71 $Y=0.41 $X2=0 $Y2=0
cc_345 N_A_154_392#_M1002_g N_X_c_870_n 0.0014982f $X=2.54 $Y=0.78 $X2=0 $Y2=0
cc_346 N_A_154_392#_c_266_n N_X_c_870_n 0.0232559f $X=0.99 $Y=0.555 $X2=0 $Y2=0
cc_347 N_A_154_392#_c_268_n N_X_c_870_n 0.0189106f $X=1.755 $Y=1.215 $X2=0 $Y2=0
cc_348 N_A_154_392#_c_269_n N_X_c_870_n 0.0197063f $X=1.85 $Y=0.555 $X2=0 $Y2=0
cc_349 N_A_154_392#_c_270_n N_X_c_870_n 0.0134082f $X=2.325 $Y=1.485 $X2=0 $Y2=0
cc_350 N_A_154_392#_c_273_n N_X_c_870_n 0.00402907f $X=1.035 $Y=1.215 $X2=0
+ $Y2=0
cc_351 N_A_154_392#_c_274_n N_X_c_870_n 0.00616549f $X=3.74 $Y=1.485 $X2=0 $Y2=0
cc_352 N_A_154_392#_c_266_n N_X_c_871_n 0.00207279f $X=0.99 $Y=0.555 $X2=0 $Y2=0
cc_353 N_A_154_392#_M1002_g N_X_c_906_n 0.00295692f $X=2.54 $Y=0.78 $X2=0 $Y2=0
cc_354 N_A_154_392#_c_269_n N_X_c_906_n 8.47036e-19 $X=1.85 $Y=0.555 $X2=0 $Y2=0
cc_355 N_A_154_392#_c_274_n N_X_c_906_n 0.00293137f $X=3.74 $Y=1.485 $X2=0 $Y2=0
cc_356 N_A_154_392#_M1002_g N_X_c_872_n 0.00926342f $X=2.54 $Y=0.78 $X2=0 $Y2=0
cc_357 N_A_154_392#_M1008_g N_X_c_872_n 0.00845441f $X=2.97 $Y=0.78 $X2=0 $Y2=0
cc_358 N_A_154_392#_M1015_g N_X_c_872_n 6.25583e-19 $X=3.445 $Y=0.795 $X2=0
+ $Y2=0
cc_359 N_A_154_392#_c_266_n N_X_c_873_n 0.00295826f $X=0.99 $Y=0.555 $X2=0 $Y2=0
cc_360 N_A_154_392#_c_270_n N_VGND_M1023_d 0.00127279f $X=2.325 $Y=1.485 $X2=0
+ $Y2=0
cc_361 N_A_154_392#_c_266_n N_VGND_c_999_n 0.00965289f $X=0.99 $Y=0.555 $X2=0
+ $Y2=0
cc_362 N_A_154_392#_c_266_n N_VGND_c_1000_n 0.0234498f $X=0.99 $Y=0.555 $X2=0
+ $Y2=0
cc_363 N_A_154_392#_c_268_n N_VGND_c_1000_n 0.0194236f $X=1.755 $Y=1.215 $X2=0
+ $Y2=0
cc_364 N_A_154_392#_c_269_n N_VGND_c_1000_n 0.0234498f $X=1.85 $Y=0.555 $X2=0
+ $Y2=0
cc_365 N_A_154_392#_c_269_n N_VGND_c_1001_n 0.00684063f $X=1.85 $Y=0.555 $X2=0
+ $Y2=0
cc_366 N_A_154_392#_M1002_g N_VGND_c_1002_n 0.00516427f $X=2.54 $Y=0.78 $X2=0
+ $Y2=0
cc_367 N_A_154_392#_c_269_n N_VGND_c_1002_n 0.0216242f $X=1.85 $Y=0.555 $X2=0
+ $Y2=0
cc_368 N_A_154_392#_c_270_n N_VGND_c_1002_n 0.0137705f $X=2.325 $Y=1.485 $X2=0
+ $Y2=0
cc_369 N_A_154_392#_c_274_n N_VGND_c_1002_n 0.00120712f $X=3.74 $Y=1.485 $X2=0
+ $Y2=0
cc_370 N_A_154_392#_M1002_g N_VGND_c_1003_n 0.00467156f $X=2.54 $Y=0.78 $X2=0
+ $Y2=0
cc_371 N_A_154_392#_M1008_g N_VGND_c_1003_n 0.00523933f $X=2.97 $Y=0.78 $X2=0
+ $Y2=0
cc_372 N_A_154_392#_M1008_g N_VGND_c_1004_n 0.00322768f $X=2.97 $Y=0.78 $X2=0
+ $Y2=0
cc_373 N_A_154_392#_M1015_g N_VGND_c_1004_n 0.00168511f $X=3.445 $Y=0.795 $X2=0
+ $Y2=0
cc_374 N_A_154_392#_M1015_g N_VGND_c_1005_n 5.1451e-19 $X=3.445 $Y=0.795 $X2=0
+ $Y2=0
cc_375 N_A_154_392#_M1020_g N_VGND_c_1005_n 0.0104924f $X=3.875 $Y=0.795 $X2=0
+ $Y2=0
cc_376 N_A_154_392#_M1020_g N_VGND_c_1006_n 0.00356909f $X=3.875 $Y=0.795 $X2=0
+ $Y2=0
cc_377 N_A_154_392#_c_264_n N_VGND_c_1006_n 0.0016924f $X=4.275 $Y=1.675 $X2=0
+ $Y2=0
cc_378 N_A_154_392#_c_271_n N_VGND_c_1006_n 0.0235203f $X=4.475 $Y=1.565 $X2=0
+ $Y2=0
cc_379 N_A_154_392#_c_271_n N_VGND_c_1007_n 0.0125065f $X=4.475 $Y=1.565 $X2=0
+ $Y2=0
cc_380 N_A_154_392#_c_275_n N_VGND_c_1007_n 0.0128578f $X=6.02 $Y=1.1 $X2=0
+ $Y2=0
cc_381 N_A_154_392#_c_266_n N_VGND_c_1010_n 0.00684063f $X=0.99 $Y=0.555 $X2=0
+ $Y2=0
cc_382 N_A_154_392#_M1015_g N_VGND_c_1012_n 0.00514022f $X=3.445 $Y=0.795 $X2=0
+ $Y2=0
cc_383 N_A_154_392#_M1020_g N_VGND_c_1012_n 0.00447026f $X=3.875 $Y=0.795 $X2=0
+ $Y2=0
cc_384 N_A_154_392#_M1002_g N_VGND_c_1014_n 0.00533081f $X=2.54 $Y=0.78 $X2=0
+ $Y2=0
cc_385 N_A_154_392#_M1008_g N_VGND_c_1014_n 0.00533081f $X=2.97 $Y=0.78 $X2=0
+ $Y2=0
cc_386 N_A_154_392#_M1015_g N_VGND_c_1014_n 0.00528353f $X=3.445 $Y=0.795 $X2=0
+ $Y2=0
cc_387 N_A_154_392#_M1020_g N_VGND_c_1014_n 0.00443817f $X=3.875 $Y=0.795 $X2=0
+ $Y2=0
cc_388 N_A_154_392#_c_266_n N_VGND_c_1014_n 0.00641317f $X=0.99 $Y=0.555 $X2=0
+ $Y2=0
cc_389 N_A_154_392#_c_269_n N_VGND_c_1014_n 0.00641317f $X=1.85 $Y=0.555 $X2=0
+ $Y2=0
cc_390 N_A_154_392#_M1004_d N_A_888_105#_c_1107_n 0.00338281f $X=5.88 $Y=0.585
+ $X2=0 $Y2=0
cc_391 N_A_154_392#_c_275_n N_A_888_105#_c_1107_n 0.0331424f $X=6.02 $Y=1.1
+ $X2=0 $Y2=0
cc_392 N_A_154_392#_c_275_n N_A_1081_39#_M1004_s 0.00591467f $X=6.02 $Y=1.1
+ $X2=-0.19 $Y2=-0.245
cc_393 N_A_154_392#_c_275_n N_A_1081_39#_c_1137_n 0.0112106f $X=6.02 $Y=1.1
+ $X2=0 $Y2=0
cc_394 N_A3_c_479_n N_A1_c_542_n 0.034253f $X=5.33 $Y=1.885 $X2=-0.19 $Y2=-0.245
cc_395 N_A3_c_477_n N_A1_M1004_g 0.00101692f $X=5.13 $Y=1.585 $X2=0 $Y2=0
cc_396 N_A3_c_477_n N_A1_c_541_n 0.0199991f $X=5.13 $Y=1.585 $X2=0 $Y2=0
cc_397 N_A3_c_481_n N_A1_c_541_n 2.79232e-19 $X=5.13 $Y=1.585 $X2=0 $Y2=0
cc_398 N_A3_c_478_n N_A_334_392#_c_674_n 0.00962345f $X=4.88 $Y=1.885 $X2=0
+ $Y2=0
cc_399 N_A3_c_479_n N_A_334_392#_c_692_n 0.0117449f $X=5.33 $Y=1.885 $X2=0 $Y2=0
cc_400 N_A3_c_478_n N_A_334_392#_c_680_n 0.00775168f $X=4.88 $Y=1.885 $X2=0
+ $Y2=0
cc_401 N_A3_c_479_n N_A_334_392#_c_680_n 0.0075092f $X=5.33 $Y=1.885 $X2=0 $Y2=0
cc_402 N_A3_c_478_n N_VPWR_c_761_n 0.00487179f $X=4.88 $Y=1.885 $X2=0 $Y2=0
cc_403 N_A3_c_478_n N_VPWR_c_762_n 0.00445602f $X=4.88 $Y=1.885 $X2=0 $Y2=0
cc_404 N_A3_c_479_n N_VPWR_c_762_n 0.00445602f $X=5.33 $Y=1.885 $X2=0 $Y2=0
cc_405 N_A3_c_479_n N_VPWR_c_763_n 0.00409001f $X=5.33 $Y=1.885 $X2=0 $Y2=0
cc_406 N_A3_c_478_n N_VPWR_c_757_n 0.00453018f $X=4.88 $Y=1.885 $X2=0 $Y2=0
cc_407 N_A3_c_479_n N_VPWR_c_757_n 0.00857673f $X=5.33 $Y=1.885 $X2=0 $Y2=0
cc_408 N_A3_c_478_n N_X_c_878_n 2.64434e-19 $X=4.88 $Y=1.885 $X2=0 $Y2=0
cc_409 N_A3_c_473_n N_VGND_c_1005_n 0.00897916f $X=4.365 $Y=1.24 $X2=0 $Y2=0
cc_410 N_A3_c_473_n N_VGND_c_1006_n 0.0136936f $X=4.365 $Y=1.24 $X2=0 $Y2=0
cc_411 N_A3_c_473_n N_VGND_c_1007_n 0.0036589f $X=4.365 $Y=1.24 $X2=0 $Y2=0
cc_412 N_A3_c_474_n N_VGND_c_1007_n 0.00241111f $X=4.72 $Y=1.315 $X2=0 $Y2=0
cc_413 N_A3_c_476_n N_VGND_c_1007_n 0.0155579f $X=4.795 $Y=1.24 $X2=0 $Y2=0
cc_414 N_A3_c_477_n N_VGND_c_1007_n 0.00777051f $X=5.13 $Y=1.585 $X2=0 $Y2=0
cc_415 N_A3_c_481_n N_VGND_c_1007_n 0.0152955f $X=5.13 $Y=1.585 $X2=0 $Y2=0
cc_416 N_A3_c_473_n N_VGND_c_1013_n 0.00452201f $X=4.365 $Y=1.24 $X2=0 $Y2=0
cc_417 N_A3_c_476_n N_VGND_c_1013_n 0.0035868f $X=4.795 $Y=1.24 $X2=0 $Y2=0
cc_418 N_A3_c_473_n N_VGND_c_1014_n 0.0049796f $X=4.365 $Y=1.24 $X2=0 $Y2=0
cc_419 N_A3_c_476_n N_VGND_c_1014_n 0.0049796f $X=4.795 $Y=1.24 $X2=0 $Y2=0
cc_420 N_A3_c_473_n N_A_888_105#_c_1106_n 0.00395841f $X=4.365 $Y=1.24 $X2=0
+ $Y2=0
cc_421 N_A3_c_476_n N_A_888_105#_c_1106_n 0.00514108f $X=4.795 $Y=1.24 $X2=0
+ $Y2=0
cc_422 N_A3_c_476_n N_A_888_105#_c_1107_n 0.00989589f $X=4.795 $Y=1.24 $X2=0
+ $Y2=0
cc_423 N_A3_c_477_n N_A_888_105#_c_1107_n 0.00530763f $X=5.13 $Y=1.585 $X2=0
+ $Y2=0
cc_424 N_A3_c_481_n N_A_888_105#_c_1107_n 0.0032428f $X=5.13 $Y=1.585 $X2=0
+ $Y2=0
cc_425 N_A3_c_476_n N_A_1081_39#_c_1136_n 8.47669e-19 $X=4.795 $Y=1.24 $X2=0
+ $Y2=0
cc_426 N_A1_c_543_n N_A2_c_599_n 0.0185951f $X=6.23 $Y=1.885 $X2=-0.19
+ $Y2=-0.245
cc_427 N_A1_M1005_g N_A2_M1010_g 0.0320723f $X=6.235 $Y=0.905 $X2=0 $Y2=0
cc_428 A1 A2 0.0261825f $X=6.875 $Y=1.58 $X2=0 $Y2=0
cc_429 A1 N_A2_c_598_n 0.0332813f $X=6.875 $Y=1.58 $X2=0 $Y2=0
cc_430 N_A1_c_541_n N_A2_c_598_n 0.0252795f $X=6.235 $Y=1.667 $X2=0 $Y2=0
cc_431 N_A1_c_542_n N_A_334_392#_c_692_n 0.0166525f $X=5.78 $Y=1.885 $X2=0 $Y2=0
cc_432 A1 N_A_334_392#_c_692_n 6.48131e-19 $X=6.875 $Y=1.58 $X2=0 $Y2=0
cc_433 N_A1_c_541_n N_A_334_392#_c_692_n 8.68446e-19 $X=6.235 $Y=1.667 $X2=0
+ $Y2=0
cc_434 N_A1_c_542_n N_A_334_392#_c_675_n 8.02991e-19 $X=5.78 $Y=1.885 $X2=0
+ $Y2=0
cc_435 A1 N_A_334_392#_c_675_n 0.0143367f $X=6.875 $Y=1.58 $X2=0 $Y2=0
cc_436 N_A1_c_541_n N_A_334_392#_c_675_n 0.00423635f $X=6.235 $Y=1.667 $X2=0
+ $Y2=0
cc_437 N_A1_c_542_n N_A_334_392#_c_676_n 0.00262152f $X=5.78 $Y=1.885 $X2=0
+ $Y2=0
cc_438 N_A1_c_543_n N_A_334_392#_c_676_n 0.00172473f $X=6.23 $Y=1.885 $X2=0
+ $Y2=0
cc_439 N_A1_c_543_n N_A_334_392#_c_677_n 0.0128889f $X=6.23 $Y=1.885 $X2=0 $Y2=0
cc_440 A1 N_A_334_392#_c_677_n 0.056787f $X=6.875 $Y=1.58 $X2=0 $Y2=0
cc_441 N_A1_c_541_n N_A_334_392#_c_677_n 0.00419876f $X=6.235 $Y=1.667 $X2=0
+ $Y2=0
cc_442 A1 N_A_334_392#_c_678_n 0.0143367f $X=6.875 $Y=1.58 $X2=0 $Y2=0
cc_443 N_A1_c_542_n N_A_334_392#_c_680_n 4.96557e-19 $X=5.78 $Y=1.885 $X2=0
+ $Y2=0
cc_444 N_A1_c_542_n N_VPWR_c_763_n 0.00712359f $X=5.78 $Y=1.885 $X2=0 $Y2=0
cc_445 N_A1_c_543_n N_VPWR_c_763_n 4.33728e-19 $X=6.23 $Y=1.885 $X2=0 $Y2=0
cc_446 N_A1_c_542_n N_VPWR_c_764_n 4.8416e-19 $X=5.78 $Y=1.885 $X2=0 $Y2=0
cc_447 N_A1_c_543_n N_VPWR_c_764_n 0.0110903f $X=6.23 $Y=1.885 $X2=0 $Y2=0
cc_448 N_A1_c_542_n N_VPWR_c_769_n 0.00413917f $X=5.78 $Y=1.885 $X2=0 $Y2=0
cc_449 N_A1_c_543_n N_VPWR_c_769_n 0.00413917f $X=6.23 $Y=1.885 $X2=0 $Y2=0
cc_450 N_A1_c_542_n N_VPWR_c_757_n 0.00817726f $X=5.78 $Y=1.885 $X2=0 $Y2=0
cc_451 N_A1_c_543_n N_VPWR_c_757_n 0.00817726f $X=6.23 $Y=1.885 $X2=0 $Y2=0
cc_452 N_A1_M1004_g N_VGND_c_1007_n 0.0012915f $X=5.805 $Y=0.905 $X2=0 $Y2=0
cc_453 N_A1_M1005_g N_A_888_105#_c_1115_n 2.33042e-19 $X=6.235 $Y=0.905 $X2=0
+ $Y2=0
cc_454 N_A1_M1004_g N_A_888_105#_c_1107_n 0.0117891f $X=5.805 $Y=0.905 $X2=0
+ $Y2=0
cc_455 N_A1_M1005_g N_A_888_105#_c_1107_n 0.0138986f $X=6.235 $Y=0.905 $X2=0
+ $Y2=0
cc_456 N_A1_M1004_g N_A_1081_39#_c_1136_n 0.00466389f $X=5.805 $Y=0.905 $X2=0
+ $Y2=0
cc_457 N_A1_M1005_g N_A_1081_39#_c_1136_n 0.00466389f $X=6.235 $Y=0.905 $X2=0
+ $Y2=0
cc_458 N_A1_M1005_g N_A_1081_39#_c_1137_n 0.00368712f $X=6.235 $Y=0.905 $X2=0
+ $Y2=0
cc_459 A1 N_A_1081_39#_c_1137_n 0.0536343f $X=6.875 $Y=1.58 $X2=0 $Y2=0
cc_460 N_A1_c_541_n N_A_1081_39#_c_1137_n 0.0022287f $X=6.235 $Y=1.667 $X2=0
+ $Y2=0
cc_461 N_A2_c_599_n N_A_334_392#_c_677_n 0.0128889f $X=6.71 $Y=1.885 $X2=0 $Y2=0
cc_462 N_A2_c_598_n N_A_334_392#_c_677_n 0.00213288f $X=7.16 $Y=1.667 $X2=0
+ $Y2=0
cc_463 N_A2_c_600_n N_A_334_392#_c_678_n 7.89448e-19 $X=7.16 $Y=1.885 $X2=0
+ $Y2=0
cc_464 N_A2_c_598_n N_A_334_392#_c_678_n 0.00423635f $X=7.16 $Y=1.667 $X2=0
+ $Y2=0
cc_465 N_A2_c_599_n N_A_334_392#_c_679_n 0.00554978f $X=6.71 $Y=1.885 $X2=0
+ $Y2=0
cc_466 N_A2_c_600_n N_A_334_392#_c_679_n 0.00279722f $X=7.16 $Y=1.885 $X2=0
+ $Y2=0
cc_467 N_A2_c_599_n N_VPWR_c_764_n 0.0111121f $X=6.71 $Y=1.885 $X2=0 $Y2=0
cc_468 N_A2_c_600_n N_VPWR_c_764_n 5.3542e-19 $X=7.16 $Y=1.885 $X2=0 $Y2=0
cc_469 N_A2_c_599_n N_VPWR_c_766_n 6.42815e-19 $X=6.71 $Y=1.885 $X2=0 $Y2=0
cc_470 N_A2_c_600_n N_VPWR_c_766_n 0.0161529f $X=7.16 $Y=1.885 $X2=0 $Y2=0
cc_471 A2 N_VPWR_c_766_n 0.0256776f $X=7.355 $Y=1.58 $X2=0 $Y2=0
cc_472 N_A2_c_598_n N_VPWR_c_766_n 0.00304264f $X=7.16 $Y=1.667 $X2=0 $Y2=0
cc_473 N_A2_c_599_n N_VPWR_c_770_n 0.00413917f $X=6.71 $Y=1.885 $X2=0 $Y2=0
cc_474 N_A2_c_600_n N_VPWR_c_770_n 0.00413917f $X=7.16 $Y=1.885 $X2=0 $Y2=0
cc_475 N_A2_c_599_n N_VPWR_c_757_n 0.00817726f $X=6.71 $Y=1.885 $X2=0 $Y2=0
cc_476 N_A2_c_600_n N_VPWR_c_757_n 0.00817726f $X=7.16 $Y=1.885 $X2=0 $Y2=0
cc_477 N_A2_M1010_g N_A_888_105#_c_1115_n 0.00186627f $X=6.725 $Y=0.905 $X2=0
+ $Y2=0
cc_478 N_A2_M1019_g N_A_888_105#_c_1115_n 0.00292963f $X=7.155 $Y=0.905 $X2=0
+ $Y2=0
cc_479 N_A2_M1010_g N_A_888_105#_c_1107_n 0.00727757f $X=6.725 $Y=0.905 $X2=0
+ $Y2=0
cc_480 N_A2_M1010_g N_A_1081_39#_c_1136_n 0.00466389f $X=6.725 $Y=0.905 $X2=0
+ $Y2=0
cc_481 N_A2_M1019_g N_A_1081_39#_c_1136_n 0.0053097f $X=7.155 $Y=0.905 $X2=0
+ $Y2=0
cc_482 N_A2_M1010_g N_A_1081_39#_c_1137_n 0.014894f $X=6.725 $Y=0.905 $X2=0
+ $Y2=0
cc_483 N_A2_M1019_g N_A_1081_39#_c_1137_n 0.017366f $X=7.155 $Y=0.905 $X2=0
+ $Y2=0
cc_484 A2 N_A_1081_39#_c_1137_n 0.00260801f $X=7.355 $Y=1.58 $X2=0 $Y2=0
cc_485 N_A2_c_598_n N_A_1081_39#_c_1137_n 0.00327642f $X=7.16 $Y=1.667 $X2=0
+ $Y2=0
cc_486 A2 N_A_1081_39#_c_1138_n 0.0183965f $X=7.355 $Y=1.58 $X2=0 $Y2=0
cc_487 N_A2_c_598_n N_A_1081_39#_c_1138_n 0.00193272f $X=7.16 $Y=1.667 $X2=0
+ $Y2=0
cc_488 N_A2_M1019_g N_A_1081_39#_c_1139_n 0.00526146f $X=7.155 $Y=0.905 $X2=0
+ $Y2=0
cc_489 N_A_69_392#_c_636_n N_A_334_392#_M1012_d 0.00226014f $X=2.105 $Y=2.99
+ $X2=-0.19 $Y2=1.66
cc_490 N_A_69_392#_M1018_s N_A_334_392#_c_674_n 0.00554861f $X=2.12 $Y=1.96
+ $X2=0 $Y2=0
cc_491 N_A_69_392#_c_636_n N_A_334_392#_c_674_n 0.00405309f $X=2.105 $Y=2.99
+ $X2=0 $Y2=0
cc_492 N_A_69_392#_c_639_n N_A_334_392#_c_674_n 0.0207097f $X=2.27 $Y=2.78 $X2=0
+ $Y2=0
cc_493 N_A_69_392#_c_636_n N_A_334_392#_c_682_n 0.0123386f $X=2.105 $Y=2.99
+ $X2=0 $Y2=0
cc_494 N_A_69_392#_c_638_n N_A_334_392#_c_682_n 0.00235516f $X=1.535 $Y=2.887
+ $X2=0 $Y2=0
cc_495 N_A_69_392#_c_639_n N_A_334_392#_c_682_n 0.00488526f $X=2.27 $Y=2.78
+ $X2=0 $Y2=0
cc_496 N_A_69_392#_c_639_n N_VPWR_c_758_n 0.0319561f $X=2.27 $Y=2.78 $X2=0 $Y2=0
cc_497 N_A_69_392#_c_637_n N_VPWR_c_767_n 0.0367837f $X=1.205 $Y=2.887 $X2=0
+ $Y2=0
cc_498 N_A_69_392#_c_638_n N_VPWR_c_767_n 0.0582926f $X=1.535 $Y=2.887 $X2=0
+ $Y2=0
cc_499 N_A_69_392#_c_639_n N_VPWR_c_767_n 0.0226174f $X=2.27 $Y=2.78 $X2=0 $Y2=0
cc_500 N_A_69_392#_c_637_n N_VPWR_c_757_n 0.0309141f $X=1.205 $Y=2.887 $X2=0
+ $Y2=0
cc_501 N_A_69_392#_c_638_n N_VPWR_c_757_n 0.0326924f $X=1.535 $Y=2.887 $X2=0
+ $Y2=0
cc_502 N_A_69_392#_c_639_n N_VPWR_c_757_n 0.0125293f $X=2.27 $Y=2.78 $X2=0 $Y2=0
cc_503 N_A_69_392#_M1006_s N_X_c_875_n 0.0100063f $X=0.345 $Y=1.96 $X2=0 $Y2=0
cc_504 N_A_69_392#_M1007_s N_X_c_875_n 0.00472114f $X=1.22 $Y=1.96 $X2=0 $Y2=0
cc_505 N_A_69_392#_c_637_n N_X_c_875_n 0.057468f $X=1.205 $Y=2.887 $X2=0 $Y2=0
cc_506 N_A_69_392#_c_638_n N_X_c_875_n 0.0105186f $X=1.535 $Y=2.887 $X2=0 $Y2=0
cc_507 N_A_69_392#_M1007_s N_X_c_888_n 0.00244362f $X=1.22 $Y=1.96 $X2=0 $Y2=0
cc_508 N_A_69_392#_M1007_s N_X_c_889_n 0.0042641f $X=1.22 $Y=1.96 $X2=0 $Y2=0
cc_509 N_A_69_392#_M1018_s N_X_c_879_n 0.00637528f $X=2.12 $Y=1.96 $X2=0 $Y2=0
cc_510 N_A_69_392#_c_638_n N_X_c_879_n 3.91771e-19 $X=1.535 $Y=2.887 $X2=0 $Y2=0
cc_511 N_A_334_392#_c_674_n N_VPWR_M1000_s 0.00527683f $X=4.94 $Y=2.405
+ $X2=-0.19 $Y2=1.66
cc_512 N_A_334_392#_c_674_n N_VPWR_M1003_s 0.00374853f $X=4.94 $Y=2.405 $X2=0
+ $Y2=0
cc_513 N_A_334_392#_c_674_n N_VPWR_M1027_s 0.00553053f $X=4.94 $Y=2.405 $X2=0
+ $Y2=0
cc_514 N_A_334_392#_c_692_n N_VPWR_M1021_s 0.00420431f $X=5.92 $Y=2.375 $X2=0
+ $Y2=0
cc_515 N_A_334_392#_c_677_n N_VPWR_M1024_s 0.00229612f $X=6.85 $Y=2.035 $X2=0
+ $Y2=0
cc_516 N_A_334_392#_c_674_n N_VPWR_c_758_n 0.0215705f $X=4.94 $Y=2.405 $X2=0
+ $Y2=0
cc_517 N_A_334_392#_c_674_n N_VPWR_c_760_n 0.0168032f $X=4.94 $Y=2.405 $X2=0
+ $Y2=0
cc_518 N_A_334_392#_c_674_n N_VPWR_c_761_n 0.0209746f $X=4.94 $Y=2.405 $X2=0
+ $Y2=0
cc_519 N_A_334_392#_c_680_n N_VPWR_c_761_n 0.0119651f $X=5.105 $Y=2.455 $X2=0
+ $Y2=0
cc_520 N_A_334_392#_c_680_n N_VPWR_c_762_n 0.0145674f $X=5.105 $Y=2.455 $X2=0
+ $Y2=0
cc_521 N_A_334_392#_c_692_n N_VPWR_c_763_n 0.0154248f $X=5.92 $Y=2.375 $X2=0
+ $Y2=0
cc_522 N_A_334_392#_c_676_n N_VPWR_c_763_n 0.0223449f $X=6.005 $Y=2.465 $X2=0
+ $Y2=0
cc_523 N_A_334_392#_c_680_n N_VPWR_c_763_n 0.0234974f $X=5.105 $Y=2.455 $X2=0
+ $Y2=0
cc_524 N_A_334_392#_c_676_n N_VPWR_c_764_n 0.034096f $X=6.005 $Y=2.465 $X2=0
+ $Y2=0
cc_525 N_A_334_392#_c_677_n N_VPWR_c_764_n 0.0196221f $X=6.85 $Y=2.035 $X2=0
+ $Y2=0
cc_526 N_A_334_392#_c_679_n N_VPWR_c_764_n 0.0452765f $X=6.935 $Y=2.815 $X2=0
+ $Y2=0
cc_527 N_A_334_392#_c_742_p N_VPWR_c_764_n 0.0124571f $X=6.005 $Y=2.375 $X2=0
+ $Y2=0
cc_528 N_A_334_392#_c_678_n N_VPWR_c_766_n 0.0123997f $X=6.935 $Y=2.12 $X2=0
+ $Y2=0
cc_529 N_A_334_392#_c_679_n N_VPWR_c_766_n 0.0560128f $X=6.935 $Y=2.815 $X2=0
+ $Y2=0
cc_530 N_A_334_392#_c_676_n N_VPWR_c_769_n 0.00749631f $X=6.005 $Y=2.465 $X2=0
+ $Y2=0
cc_531 N_A_334_392#_c_679_n N_VPWR_c_770_n 0.00749631f $X=6.935 $Y=2.815 $X2=0
+ $Y2=0
cc_532 N_A_334_392#_c_674_n N_VPWR_c_757_n 0.0518786f $X=4.94 $Y=2.405 $X2=0
+ $Y2=0
cc_533 N_A_334_392#_c_676_n N_VPWR_c_757_n 0.0062048f $X=6.005 $Y=2.465 $X2=0
+ $Y2=0
cc_534 N_A_334_392#_c_679_n N_VPWR_c_757_n 0.0062048f $X=6.935 $Y=2.815 $X2=0
+ $Y2=0
cc_535 N_A_334_392#_c_680_n N_VPWR_c_757_n 0.0119851f $X=5.105 $Y=2.455 $X2=0
+ $Y2=0
cc_536 N_A_334_392#_c_674_n N_X_M1000_d 0.00553763f $X=4.94 $Y=2.405 $X2=0 $Y2=0
cc_537 N_A_334_392#_c_674_n N_X_M1026_d 0.00553763f $X=4.94 $Y=2.405 $X2=0 $Y2=0
cc_538 N_A_334_392#_c_674_n N_X_c_877_n 0.10342f $X=4.94 $Y=2.405 $X2=0 $Y2=0
cc_539 N_A_334_392#_M1012_d N_X_c_879_n 0.00408401f $X=1.67 $Y=1.96 $X2=0 $Y2=0
cc_540 N_A_334_392#_c_674_n N_X_c_879_n 0.0348102f $X=4.94 $Y=2.405 $X2=0 $Y2=0
cc_541 N_A_334_392#_c_682_n N_X_c_879_n 0.0131605f $X=1.82 $Y=2.405 $X2=0 $Y2=0
cc_542 N_VPWR_c_757_n N_X_c_875_n 0.00179127f $X=7.44 $Y=3.33 $X2=0 $Y2=0
cc_543 N_VPWR_c_757_n N_X_c_876_n 0.00690149f $X=7.44 $Y=3.33 $X2=0 $Y2=0
cc_544 N_VPWR_M1000_s N_X_c_877_n 6.9948e-19 $X=2.665 $Y=1.84 $X2=0 $Y2=0
cc_545 N_VPWR_M1000_s N_X_c_878_n 0.00326831f $X=2.665 $Y=1.84 $X2=0 $Y2=0
cc_546 N_VPWR_M1003_s N_X_c_878_n 0.00202293f $X=3.54 $Y=1.84 $X2=0 $Y2=0
cc_547 N_X_c_870_n N_VGND_M1014_d 0.00713477f $X=2.495 $Y=0.925 $X2=-0.19
+ $Y2=-0.245
cc_548 N_X_c_870_n N_VGND_M1025_d 0.00212101f $X=2.495 $Y=0.925 $X2=0 $Y2=0
cc_549 N_X_c_870_n N_VGND_M1023_d 0.00654612f $X=2.495 $Y=0.925 $X2=0 $Y2=0
cc_550 N_X_c_927_n N_VGND_M1008_d 0.0041598f $X=3.495 $Y=1.065 $X2=0 $Y2=0
cc_551 N_X_c_870_n N_VGND_c_999_n 0.0162807f $X=2.495 $Y=0.925 $X2=0 $Y2=0
cc_552 N_X_c_870_n N_VGND_c_1000_n 0.0241426f $X=2.495 $Y=0.925 $X2=0 $Y2=0
cc_553 N_X_c_870_n N_VGND_c_1002_n 0.0189501f $X=2.495 $Y=0.925 $X2=0 $Y2=0
cc_554 N_X_c_906_n N_VGND_c_1002_n 0.00118216f $X=2.64 $Y=0.925 $X2=0 $Y2=0
cc_555 N_X_c_872_n N_VGND_c_1002_n 0.042245f $X=2.755 $Y=0.555 $X2=0 $Y2=0
cc_556 N_X_c_872_n N_VGND_c_1003_n 0.014429f $X=2.755 $Y=0.555 $X2=0 $Y2=0
cc_557 N_X_c_927_n N_VGND_c_1004_n 0.0171667f $X=3.495 $Y=1.065 $X2=0 $Y2=0
cc_558 N_X_c_869_n N_VGND_c_1004_n 0.0146226f $X=3.66 $Y=0.57 $X2=0 $Y2=0
cc_559 N_X_c_872_n N_VGND_c_1004_n 0.0161242f $X=2.755 $Y=0.555 $X2=0 $Y2=0
cc_560 N_X_c_869_n N_VGND_c_1005_n 0.0188983f $X=3.66 $Y=0.57 $X2=0 $Y2=0
cc_561 N_X_c_869_n N_VGND_c_1012_n 0.00899058f $X=3.66 $Y=0.57 $X2=0 $Y2=0
cc_562 N_X_c_869_n N_VGND_c_1014_n 0.00882735f $X=3.66 $Y=0.57 $X2=0 $Y2=0
cc_563 N_X_c_872_n N_VGND_c_1014_n 0.0137073f $X=2.755 $Y=0.555 $X2=0 $Y2=0
cc_564 N_X_c_873_n N_VGND_c_1014_n 0.00489676f $X=0.24 $Y=0.925 $X2=0 $Y2=0
cc_565 N_VGND_c_1007_n N_A_888_105#_M1009_d 0.00179007f $X=5.01 $Y=1.02
+ $X2=-0.19 $Y2=-0.245
cc_566 N_VGND_c_1005_n N_A_888_105#_c_1106_n 0.0156621f $X=4.09 $Y=0.57 $X2=0
+ $Y2=0
cc_567 N_VGND_c_1006_n N_A_888_105#_c_1106_n 7.25226e-19 $X=4.425 $Y=1.06 $X2=0
+ $Y2=0
cc_568 N_VGND_c_1007_n N_A_888_105#_c_1106_n 0.0429099f $X=5.01 $Y=1.02 $X2=0
+ $Y2=0
cc_569 N_VGND_c_1013_n N_A_888_105#_c_1106_n 0.00828248f $X=7.44 $Y=0 $X2=0
+ $Y2=0
cc_570 N_VGND_c_1014_n N_A_888_105#_c_1106_n 0.0105304f $X=7.44 $Y=0 $X2=0 $Y2=0
cc_571 N_VGND_M1011_s N_A_888_105#_c_1107_n 0.00629528f $X=4.87 $Y=0.525 $X2=0
+ $Y2=0
cc_572 N_VGND_c_1013_n N_A_888_105#_c_1107_n 0.0114112f $X=7.44 $Y=0 $X2=0 $Y2=0
cc_573 N_VGND_c_1014_n N_A_888_105#_c_1107_n 0.0216401f $X=7.44 $Y=0 $X2=0 $Y2=0
cc_574 N_VGND_c_1014_n N_A_1081_39#_M1004_s 0.00243084f $X=7.44 $Y=0 $X2=-0.19
+ $Y2=-0.245
cc_575 N_VGND_c_1013_n N_A_1081_39#_c_1136_n 0.141318f $X=7.44 $Y=0 $X2=0 $Y2=0
cc_576 N_VGND_c_1014_n N_A_1081_39#_c_1136_n 0.0819032f $X=7.44 $Y=0 $X2=0 $Y2=0
cc_577 N_A_888_105#_c_1107_n N_A_1081_39#_M1004_s 0.0104558f $X=6.775 $Y=0.705
+ $X2=-0.19 $Y2=-0.245
cc_578 N_A_888_105#_c_1107_n N_A_1081_39#_M1005_s 0.00495268f $X=6.775 $Y=0.705
+ $X2=0 $Y2=0
cc_579 N_A_888_105#_c_1107_n N_A_1081_39#_c_1136_n 0.107329f $X=6.775 $Y=0.705
+ $X2=0 $Y2=0
cc_580 N_A_888_105#_M1010_s N_A_1081_39#_c_1137_n 0.00179223f $X=6.8 $Y=0.585
+ $X2=0 $Y2=0
cc_581 N_A_888_105#_c_1115_n N_A_1081_39#_c_1137_n 0.016192f $X=6.94 $Y=0.73
+ $X2=0 $Y2=0
cc_582 N_A_888_105#_c_1107_n N_A_1081_39#_c_1137_n 0.0225078f $X=6.775 $Y=0.705
+ $X2=0 $Y2=0
