* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hs__and4b_1 A_N B C D VGND VNB VPB VPWR X
X0 a_526_139# D VGND VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X1 a_353_124# B a_448_139# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X2 VPWR C a_226_424# VPB sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X3 VGND a_226_424# X VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X4 a_448_139# C a_526_139# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X5 a_226_424# D VPWR VPB sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X6 VPWR a_226_424# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X7 a_226_424# a_27_74# a_353_124# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X8 VPWR a_27_74# a_226_424# VPB sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X9 a_27_74# A_N VPWR VPB sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X10 a_226_424# B VPWR VPB sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X11 a_27_74# A_N VGND VNB sky130_fd_pr__nfet_01v8_lvt w=550000u l=150000u
.ends
