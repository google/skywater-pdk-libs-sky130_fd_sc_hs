* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hs__dfxbp_1 CLK D VGND VNB VPB VPWR Q Q_N
X0 VGND D a_420_503# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X1 VPWR a_543_447# a_701_463# VPB sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X2 VGND a_1644_94# Q_N VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X3 VPWR D a_420_503# VPB sky130_fd_pr__pfet_01v8 w=420000u l=150000u
X4 a_1158_482# a_1191_120# VPWR VPB sky130_fd_pr__pfet_01v8 w=420000u l=150000u
X5 a_543_447# a_205_368# a_713_102# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X6 a_713_102# a_701_463# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X7 a_27_74# CLK VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X8 a_1644_94# a_1191_120# VPWR VPB sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X9 VPWR a_1644_94# Q_N VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X10 a_543_447# a_27_74# a_650_508# VPB sky130_fd_pr__pfet_01v8 w=420000u l=150000u
X11 a_1191_120# a_1005_120# VPWR VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=150000u
X12 VPWR a_1191_120# Q VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X13 VGND a_27_74# a_205_368# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X14 a_701_463# a_27_74# a_1005_120# VPB sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X15 a_420_503# a_27_74# a_543_447# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X16 a_1005_120# a_27_74# a_1143_146# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X17 a_650_508# a_701_463# VPWR VPB sky130_fd_pr__pfet_01v8 w=420000u l=150000u
X18 a_1143_146# a_1191_120# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X19 VGND a_1191_120# Q VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X20 a_420_503# a_205_368# a_543_447# VPB sky130_fd_pr__pfet_01v8 w=420000u l=150000u
X21 a_1191_120# a_1005_120# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X22 VPWR a_27_74# a_205_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X23 a_1005_120# a_205_368# a_1158_482# VPB sky130_fd_pr__pfet_01v8 w=420000u l=150000u
X24 a_701_463# a_205_368# a_1005_120# VNB sky130_fd_pr__nfet_01v8_lvt w=550000u l=150000u
X25 a_1644_94# a_1191_120# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X26 VGND a_543_447# a_701_463# VNB sky130_fd_pr__nfet_01v8_lvt w=550000u l=150000u
X27 a_27_74# CLK VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
.ends
