* File: sky130_fd_sc_hs__nand4b_1.pxi.spice
* Created: Thu Aug 27 20:52:06 2020
* 
x_PM_SKY130_FD_SC_HS__NAND4B_1%A_N N_A_N_c_52_n N_A_N_M1007_g N_A_N_c_53_n
+ N_A_N_M1006_g A_N PM_SKY130_FD_SC_HS__NAND4B_1%A_N
x_PM_SKY130_FD_SC_HS__NAND4B_1%D N_D_c_77_n N_D_M1002_g N_D_c_78_n N_D_M1008_g D
+ PM_SKY130_FD_SC_HS__NAND4B_1%D
x_PM_SKY130_FD_SC_HS__NAND4B_1%C N_C_c_106_n N_C_M1009_g N_C_c_107_n N_C_M1004_g
+ C PM_SKY130_FD_SC_HS__NAND4B_1%C
x_PM_SKY130_FD_SC_HS__NAND4B_1%B N_B_c_135_n N_B_M1000_g N_B_c_136_n N_B_M1001_g
+ B PM_SKY130_FD_SC_HS__NAND4B_1%B
x_PM_SKY130_FD_SC_HS__NAND4B_1%A_27_112# N_A_27_112#_M1006_s N_A_27_112#_M1007_s
+ N_A_27_112#_c_165_n N_A_27_112#_M1003_g N_A_27_112#_c_166_n
+ N_A_27_112#_M1005_g N_A_27_112#_c_167_n N_A_27_112#_c_174_n
+ N_A_27_112#_c_168_n N_A_27_112#_c_172_n N_A_27_112#_c_169_n
+ N_A_27_112#_c_180_n N_A_27_112#_c_182_n N_A_27_112#_c_170_n
+ PM_SKY130_FD_SC_HS__NAND4B_1%A_27_112#
x_PM_SKY130_FD_SC_HS__NAND4B_1%VPWR N_VPWR_M1007_d N_VPWR_M1004_d N_VPWR_M1005_d
+ N_VPWR_c_233_n N_VPWR_c_234_n N_VPWR_c_235_n N_VPWR_c_236_n N_VPWR_c_237_n
+ N_VPWR_c_238_n N_VPWR_c_239_n N_VPWR_c_240_n VPWR N_VPWR_c_241_n
+ N_VPWR_c_232_n PM_SKY130_FD_SC_HS__NAND4B_1%VPWR
x_PM_SKY130_FD_SC_HS__NAND4B_1%Y N_Y_M1003_d N_Y_M1002_d N_Y_M1001_d N_Y_c_281_n
+ N_Y_c_282_n N_Y_c_283_n N_Y_c_284_n N_Y_c_278_n N_Y_c_279_n N_Y_c_286_n
+ N_Y_c_287_n N_Y_c_280_n Y PM_SKY130_FD_SC_HS__NAND4B_1%Y
x_PM_SKY130_FD_SC_HS__NAND4B_1%VGND N_VGND_M1006_d N_VGND_c_333_n N_VGND_c_334_n
+ N_VGND_c_335_n VGND N_VGND_c_336_n N_VGND_c_337_n
+ PM_SKY130_FD_SC_HS__NAND4B_1%VGND
cc_1 VNB N_A_N_c_52_n 0.0420363f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.765
cc_2 VNB N_A_N_c_53_n 0.0224562f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=1.22
cc_3 VNB A_N 0.00846479f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_4 VNB N_D_c_77_n 0.0386516f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.765
cc_5 VNB N_D_c_78_n 0.0189071f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=1.22
cc_6 VNB D 0.00411297f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_7 VNB N_C_c_106_n 0.0178699f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.765
cc_8 VNB N_C_c_107_n 0.0385576f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=1.22
cc_9 VNB C 0.00365302f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_10 VNB N_B_c_135_n 0.0191804f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.765
cc_11 VNB N_B_c_136_n 0.0364511f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=1.22
cc_12 VNB B 0.00602028f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_13 VNB N_A_27_112#_c_165_n 0.0220447f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_14 VNB N_A_27_112#_c_166_n 0.0433553f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.385
cc_15 VNB N_A_27_112#_c_167_n 0.0140131f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_27_112#_c_168_n 0.0011463f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_27_112#_c_169_n 0.0298066f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_27_112#_c_170_n 0.0055235f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_VPWR_c_232_n 0.143779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_Y_c_278_n 0.0241427f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_Y_c_279_n 0.028403f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_Y_c_280_n 0.00739565f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_VGND_c_333_n 0.013703f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=0.835
cc_24 VNB N_VGND_c_334_n 0.0271358f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.385
cc_25 VNB N_VGND_c_335_n 0.00616254f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.385
cc_26 VNB N_VGND_c_336_n 0.0683234f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_VGND_c_337_n 0.219095f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VPB N_A_N_c_52_n 0.0286883f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.765
cc_29 VPB N_D_c_77_n 0.024381f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.765
cc_30 VPB N_C_c_107_n 0.0233973f $X=-0.19 $Y=1.66 $X2=0.7 $Y2=1.22
cc_31 VPB N_B_c_136_n 0.0228776f $X=-0.19 $Y=1.66 $X2=0.7 $Y2=1.22
cc_32 VPB N_A_27_112#_c_166_n 0.0240522f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=1.385
cc_33 VPB N_A_27_112#_c_172_n 0.0536112f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_34 VPB N_A_27_112#_c_169_n 0.00809293f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_35 VPB N_VPWR_c_233_n 0.0283042f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=1.365
cc_36 VPB N_VPWR_c_234_n 0.00900819f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_37 VPB N_VPWR_c_235_n 0.0156997f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_38 VPB N_VPWR_c_236_n 0.047631f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_39 VPB N_VPWR_c_237_n 0.0249968f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_40 VPB N_VPWR_c_238_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_41 VPB N_VPWR_c_239_n 0.0186948f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_42 VPB N_VPWR_c_240_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_43 VPB N_VPWR_c_241_n 0.019175f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_44 VPB N_VPWR_c_232_n 0.0710834f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_45 VPB N_Y_c_281_n 0.00963304f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=1.385
cc_46 VPB N_Y_c_282_n 0.00257348f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=1.365
cc_47 VPB N_Y_c_283_n 0.00257348f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_48 VPB N_Y_c_284_n 0.0178895f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_49 VPB N_Y_c_279_n 0.00301454f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_50 VPB N_Y_c_286_n 0.00837886f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_51 VPB N_Y_c_287_n 0.00769224f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_52 N_A_N_c_52_n N_D_c_77_n 0.0483056f $X=0.64 $Y=1.765 $X2=-0.19 $Y2=-0.245
cc_53 A_N N_D_c_77_n 0.00187636f $X=0.635 $Y=1.21 $X2=-0.19 $Y2=-0.245
cc_54 N_A_N_c_53_n N_D_c_78_n 0.019495f $X=0.7 $Y=1.22 $X2=0 $Y2=0
cc_55 N_A_N_c_52_n D 3.7859e-19 $X=0.64 $Y=1.765 $X2=0 $Y2=0
cc_56 A_N D 0.0296943f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_57 N_A_N_c_53_n N_A_27_112#_c_174_n 0.0089549f $X=0.7 $Y=1.22 $X2=0 $Y2=0
cc_58 N_A_N_c_52_n N_A_27_112#_c_172_n 0.0169002f $X=0.64 $Y=1.765 $X2=0 $Y2=0
cc_59 A_N N_A_27_112#_c_172_n 0.00800159f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_60 N_A_N_c_52_n N_A_27_112#_c_169_n 0.0106614f $X=0.64 $Y=1.765 $X2=0 $Y2=0
cc_61 N_A_N_c_53_n N_A_27_112#_c_169_n 0.00457953f $X=0.7 $Y=1.22 $X2=0 $Y2=0
cc_62 A_N N_A_27_112#_c_169_n 0.0282012f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_63 N_A_N_c_52_n N_A_27_112#_c_180_n 0.00105413f $X=0.64 $Y=1.765 $X2=0 $Y2=0
cc_64 A_N N_A_27_112#_c_180_n 0.0250429f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_65 N_A_N_c_53_n N_A_27_112#_c_182_n 0.00455786f $X=0.7 $Y=1.22 $X2=0 $Y2=0
cc_66 N_A_N_c_52_n N_VPWR_c_233_n 0.0116362f $X=0.64 $Y=1.765 $X2=0 $Y2=0
cc_67 A_N N_VPWR_c_233_n 0.00187223f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_68 N_A_N_c_52_n N_VPWR_c_237_n 0.00393873f $X=0.64 $Y=1.765 $X2=0 $Y2=0
cc_69 N_A_N_c_52_n N_VPWR_c_232_n 0.00462577f $X=0.64 $Y=1.765 $X2=0 $Y2=0
cc_70 N_A_N_c_53_n N_VGND_c_333_n 0.00662399f $X=0.7 $Y=1.22 $X2=0 $Y2=0
cc_71 N_A_N_c_53_n N_VGND_c_334_n 0.00434489f $X=0.7 $Y=1.22 $X2=0 $Y2=0
cc_72 N_A_N_c_53_n N_VGND_c_337_n 0.00487769f $X=0.7 $Y=1.22 $X2=0 $Y2=0
cc_73 N_D_c_78_n N_C_c_106_n 0.0541207f $X=1.24 $Y=1.22 $X2=-0.19 $Y2=-0.245
cc_74 N_D_c_77_n N_C_c_107_n 0.0416401f $X=1.225 $Y=1.765 $X2=0 $Y2=0
cc_75 D N_C_c_107_n 0.00114936f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_76 N_D_c_77_n C 0.00114936f $X=1.225 $Y=1.765 $X2=0 $Y2=0
cc_77 N_D_c_78_n C 2.19577e-19 $X=1.24 $Y=1.22 $X2=0 $Y2=0
cc_78 D C 0.0235844f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_79 N_D_c_77_n N_A_27_112#_c_174_n 0.00101144f $X=1.225 $Y=1.765 $X2=0 $Y2=0
cc_80 N_D_c_78_n N_A_27_112#_c_174_n 0.0119277f $X=1.24 $Y=1.22 $X2=0 $Y2=0
cc_81 D N_A_27_112#_c_174_n 0.0228656f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_82 N_D_c_78_n N_A_27_112#_c_182_n 5.7889e-19 $X=1.24 $Y=1.22 $X2=0 $Y2=0
cc_83 N_D_c_77_n N_VPWR_c_233_n 0.0140342f $X=1.225 $Y=1.765 $X2=0 $Y2=0
cc_84 D N_VPWR_c_233_n 0.00773068f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_85 N_D_c_77_n N_VPWR_c_239_n 0.00445602f $X=1.225 $Y=1.765 $X2=0 $Y2=0
cc_86 N_D_c_77_n N_VPWR_c_232_n 0.00861803f $X=1.225 $Y=1.765 $X2=0 $Y2=0
cc_87 N_D_c_77_n N_Y_c_281_n 0.00482258f $X=1.225 $Y=1.765 $X2=0 $Y2=0
cc_88 D N_Y_c_281_n 0.00168052f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_89 N_D_c_77_n N_Y_c_282_n 0.0090468f $X=1.225 $Y=1.765 $X2=0 $Y2=0
cc_90 N_D_c_78_n N_VGND_c_333_n 0.0107451f $X=1.24 $Y=1.22 $X2=0 $Y2=0
cc_91 N_D_c_78_n N_VGND_c_336_n 0.00398535f $X=1.24 $Y=1.22 $X2=0 $Y2=0
cc_92 N_D_c_78_n N_VGND_c_337_n 0.00398847f $X=1.24 $Y=1.22 $X2=0 $Y2=0
cc_93 N_C_c_106_n N_B_c_135_n 0.037909f $X=1.63 $Y=1.22 $X2=-0.19 $Y2=-0.245
cc_94 N_C_c_107_n N_B_c_136_n 0.0573559f $X=1.675 $Y=1.765 $X2=0 $Y2=0
cc_95 C N_B_c_136_n 3.99347e-19 $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_96 N_C_c_107_n B 0.00188716f $X=1.675 $Y=1.765 $X2=0 $Y2=0
cc_97 C B 0.0272327f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_98 N_C_c_106_n N_A_27_112#_c_174_n 0.0119829f $X=1.63 $Y=1.22 $X2=0 $Y2=0
cc_99 N_C_c_107_n N_A_27_112#_c_174_n 8.19833e-19 $X=1.675 $Y=1.765 $X2=0 $Y2=0
cc_100 C N_A_27_112#_c_174_n 0.0218012f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_101 N_C_c_107_n N_VPWR_c_234_n 0.00599602f $X=1.675 $Y=1.765 $X2=0 $Y2=0
cc_102 N_C_c_107_n N_VPWR_c_239_n 0.00445602f $X=1.675 $Y=1.765 $X2=0 $Y2=0
cc_103 N_C_c_107_n N_VPWR_c_232_n 0.00858056f $X=1.675 $Y=1.765 $X2=0 $Y2=0
cc_104 N_C_c_107_n N_Y_c_281_n 0.0252765f $X=1.675 $Y=1.765 $X2=0 $Y2=0
cc_105 C N_Y_c_281_n 0.0223616f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_106 N_C_c_107_n N_Y_c_282_n 0.0106769f $X=1.675 $Y=1.765 $X2=0 $Y2=0
cc_107 N_C_c_107_n N_Y_c_283_n 6.74978e-19 $X=1.675 $Y=1.765 $X2=0 $Y2=0
cc_108 C N_Y_c_286_n 0.00192199f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_109 N_C_c_106_n N_VGND_c_333_n 0.00212642f $X=1.63 $Y=1.22 $X2=0 $Y2=0
cc_110 N_C_c_106_n N_VGND_c_336_n 0.00461464f $X=1.63 $Y=1.22 $X2=0 $Y2=0
cc_111 N_C_c_106_n N_VGND_c_337_n 0.00465092f $X=1.63 $Y=1.22 $X2=0 $Y2=0
cc_112 N_B_c_135_n N_A_27_112#_c_165_n 0.0312011f $X=2.14 $Y=1.22 $X2=0 $Y2=0
cc_113 N_B_c_136_n N_A_27_112#_c_166_n 0.0421628f $X=2.245 $Y=1.765 $X2=0 $Y2=0
cc_114 B N_A_27_112#_c_166_n 3.77186e-19 $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_115 N_B_c_135_n N_A_27_112#_c_174_n 0.0127995f $X=2.14 $Y=1.22 $X2=0 $Y2=0
cc_116 N_B_c_136_n N_A_27_112#_c_174_n 0.00100398f $X=2.245 $Y=1.765 $X2=0 $Y2=0
cc_117 B N_A_27_112#_c_174_n 0.0237469f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_118 N_B_c_135_n N_A_27_112#_c_168_n 0.00162255f $X=2.14 $Y=1.22 $X2=0 $Y2=0
cc_119 B N_A_27_112#_c_168_n 0.00318562f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_120 N_B_c_136_n N_A_27_112#_c_170_n 0.00187066f $X=2.245 $Y=1.765 $X2=0 $Y2=0
cc_121 B N_A_27_112#_c_170_n 0.0264357f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_122 N_B_c_136_n N_VPWR_c_234_n 0.0071356f $X=2.245 $Y=1.765 $X2=0 $Y2=0
cc_123 N_B_c_136_n N_VPWR_c_241_n 0.00422942f $X=2.245 $Y=1.765 $X2=0 $Y2=0
cc_124 N_B_c_136_n N_VPWR_c_232_n 0.0078513f $X=2.245 $Y=1.765 $X2=0 $Y2=0
cc_125 N_B_c_136_n N_Y_c_282_n 6.50327e-19 $X=2.245 $Y=1.765 $X2=0 $Y2=0
cc_126 N_B_c_136_n N_Y_c_283_n 0.0120063f $X=2.245 $Y=1.765 $X2=0 $Y2=0
cc_127 N_B_c_136_n N_Y_c_286_n 0.0197998f $X=2.245 $Y=1.765 $X2=0 $Y2=0
cc_128 B N_Y_c_286_n 0.0190624f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_129 N_B_c_136_n N_Y_c_287_n 0.00442429f $X=2.245 $Y=1.765 $X2=0 $Y2=0
cc_130 B N_Y_c_287_n 0.00908459f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_131 N_B_c_135_n N_VGND_c_336_n 0.00461464f $X=2.14 $Y=1.22 $X2=0 $Y2=0
cc_132 N_B_c_135_n N_VGND_c_337_n 0.00466411f $X=2.14 $Y=1.22 $X2=0 $Y2=0
cc_133 N_A_27_112#_c_172_n N_VPWR_c_233_n 0.0608022f $X=0.415 $Y=1.985 $X2=0
+ $Y2=0
cc_134 N_A_27_112#_c_166_n N_VPWR_c_236_n 0.0227729f $X=2.695 $Y=1.765 $X2=0
+ $Y2=0
cc_135 N_A_27_112#_c_172_n N_VPWR_c_237_n 0.00964662f $X=0.415 $Y=1.985 $X2=0
+ $Y2=0
cc_136 N_A_27_112#_c_166_n N_VPWR_c_241_n 0.00445602f $X=2.695 $Y=1.765 $X2=0
+ $Y2=0
cc_137 N_A_27_112#_c_166_n N_VPWR_c_232_n 0.00860917f $X=2.695 $Y=1.765 $X2=0
+ $Y2=0
cc_138 N_A_27_112#_c_172_n N_VPWR_c_232_n 0.0143899f $X=0.415 $Y=1.985 $X2=0
+ $Y2=0
cc_139 N_A_27_112#_c_166_n N_Y_c_283_n 0.00925663f $X=2.695 $Y=1.765 $X2=0 $Y2=0
cc_140 N_A_27_112#_c_166_n N_Y_c_284_n 0.0175131f $X=2.695 $Y=1.765 $X2=0 $Y2=0
cc_141 N_A_27_112#_c_170_n N_Y_c_284_n 0.0219515f $X=2.77 $Y=1.385 $X2=0 $Y2=0
cc_142 N_A_27_112#_c_165_n N_Y_c_278_n 0.0230379f $X=2.68 $Y=1.22 $X2=0 $Y2=0
cc_143 N_A_27_112#_c_174_n N_Y_c_278_n 0.0140856f $X=2.565 $Y=0.925 $X2=0 $Y2=0
cc_144 N_A_27_112#_c_165_n N_Y_c_279_n 0.00289106f $X=2.68 $Y=1.22 $X2=0 $Y2=0
cc_145 N_A_27_112#_c_166_n N_Y_c_279_n 0.0073612f $X=2.695 $Y=1.765 $X2=0 $Y2=0
cc_146 N_A_27_112#_c_168_n N_Y_c_279_n 0.00669252f $X=2.65 $Y=1.22 $X2=0 $Y2=0
cc_147 N_A_27_112#_c_170_n N_Y_c_279_n 0.0249903f $X=2.77 $Y=1.385 $X2=0 $Y2=0
cc_148 N_A_27_112#_c_166_n N_Y_c_287_n 0.0112884f $X=2.695 $Y=1.765 $X2=0 $Y2=0
cc_149 N_A_27_112#_c_170_n N_Y_c_287_n 0.0059332f $X=2.77 $Y=1.385 $X2=0 $Y2=0
cc_150 N_A_27_112#_c_166_n N_Y_c_280_n 6.75008e-19 $X=2.695 $Y=1.765 $X2=0 $Y2=0
cc_151 N_A_27_112#_c_168_n N_Y_c_280_n 0.00295346f $X=2.65 $Y=1.22 $X2=0 $Y2=0
cc_152 N_A_27_112#_c_170_n N_Y_c_280_n 0.00240045f $X=2.77 $Y=1.385 $X2=0 $Y2=0
cc_153 N_A_27_112#_c_174_n N_VGND_M1006_d 0.0103133f $X=2.565 $Y=0.925 $X2=-0.19
+ $Y2=-0.245
cc_154 N_A_27_112#_c_174_n N_VGND_c_333_n 0.0214267f $X=2.565 $Y=0.925 $X2=0
+ $Y2=0
cc_155 N_A_27_112#_c_167_n N_VGND_c_334_n 0.00300961f $X=0.275 $Y=0.845 $X2=0
+ $Y2=0
cc_156 N_A_27_112#_c_180_n N_VGND_c_334_n 0.00572092f $X=0.485 $Y=0.845 $X2=0
+ $Y2=0
cc_157 N_A_27_112#_c_165_n N_VGND_c_336_n 0.00461464f $X=2.68 $Y=1.22 $X2=0
+ $Y2=0
cc_158 N_A_27_112#_c_165_n N_VGND_c_337_n 0.00528843f $X=2.68 $Y=1.22 $X2=0
+ $Y2=0
cc_159 N_A_27_112#_c_167_n N_VGND_c_337_n 0.00499017f $X=0.275 $Y=0.845 $X2=0
+ $Y2=0
cc_160 N_A_27_112#_c_174_n N_VGND_c_337_n 0.0577132f $X=2.565 $Y=0.925 $X2=0
+ $Y2=0
cc_161 N_A_27_112#_c_180_n N_VGND_c_337_n 0.0105838f $X=0.485 $Y=0.845 $X2=0
+ $Y2=0
cc_162 N_A_27_112#_c_174_n A_263_74# 0.00734082f $X=2.565 $Y=0.925 $X2=-0.19
+ $Y2=-0.245
cc_163 N_A_27_112#_c_174_n A_341_74# 0.0116011f $X=2.565 $Y=0.925 $X2=-0.19
+ $Y2=-0.245
cc_164 N_A_27_112#_c_174_n A_443_74# 0.0127373f $X=2.565 $Y=0.925 $X2=-0.19
+ $Y2=-0.245
cc_165 N_VPWR_M1004_d N_Y_c_281_n 2.5099e-19 $X=1.75 $Y=1.84 $X2=0 $Y2=0
cc_166 N_VPWR_c_233_n N_Y_c_281_n 0.0146948f $X=0.95 $Y=1.985 $X2=0 $Y2=0
cc_167 N_VPWR_c_234_n N_Y_c_281_n 0.00200558f $X=1.95 $Y=2.405 $X2=0 $Y2=0
cc_168 N_VPWR_c_233_n N_Y_c_282_n 0.0318965f $X=0.95 $Y=1.985 $X2=0 $Y2=0
cc_169 N_VPWR_c_234_n N_Y_c_282_n 0.0255553f $X=1.95 $Y=2.405 $X2=0 $Y2=0
cc_170 N_VPWR_c_239_n N_Y_c_282_n 0.014552f $X=1.785 $Y=3.33 $X2=0 $Y2=0
cc_171 N_VPWR_c_232_n N_Y_c_282_n 0.0119791f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_172 N_VPWR_c_234_n N_Y_c_283_n 0.0257793f $X=1.95 $Y=2.405 $X2=0 $Y2=0
cc_173 N_VPWR_c_236_n N_Y_c_283_n 0.032178f $X=2.97 $Y=2.145 $X2=0 $Y2=0
cc_174 N_VPWR_c_241_n N_Y_c_283_n 0.0153846f $X=2.805 $Y=3.33 $X2=0 $Y2=0
cc_175 N_VPWR_c_232_n N_Y_c_283_n 0.0126213f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_176 N_VPWR_M1005_d N_Y_c_284_n 0.00345989f $X=2.77 $Y=1.84 $X2=0 $Y2=0
cc_177 N_VPWR_c_236_n N_Y_c_284_n 0.0252631f $X=2.97 $Y=2.145 $X2=0 $Y2=0
cc_178 N_VPWR_M1004_d N_Y_c_286_n 0.00393632f $X=1.75 $Y=1.84 $X2=0 $Y2=0
cc_179 N_VPWR_c_234_n N_Y_c_286_n 0.0245184f $X=1.95 $Y=2.405 $X2=0 $Y2=0
cc_180 N_Y_c_278_n N_VGND_c_336_n 0.0164394f $X=2.99 $Y=0.515 $X2=0 $Y2=0
cc_181 N_Y_c_278_n N_VGND_c_337_n 0.0135988f $X=2.99 $Y=0.515 $X2=0 $Y2=0
