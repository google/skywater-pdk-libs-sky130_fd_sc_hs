* File: sky130_fd_sc_hs__o21bai_4.pxi.spice
* Created: Thu Aug 27 20:59:01 2020
* 
x_PM_SKY130_FD_SC_HS__O21BAI_4%A1 N_A1_M1006_g N_A1_c_135_n N_A1_M1008_g
+ N_A1_c_136_n N_A1_M1009_g N_A1_M1016_g N_A1_M1019_g N_A1_c_137_n N_A1_M1010_g
+ N_A1_c_129_n N_A1_c_130_n N_A1_M1022_g N_A1_c_132_n N_A1_c_140_n N_A1_M1012_g
+ N_A1_c_133_n A1 A1 A1 A1 PM_SKY130_FD_SC_HS__O21BAI_4%A1
x_PM_SKY130_FD_SC_HS__O21BAI_4%A2 N_A2_M1003_g N_A2_c_212_n N_A2_c_221_n
+ N_A2_M1014_g N_A2_c_213_n N_A2_M1005_g N_A2_c_222_n N_A2_M1017_g N_A2_M1013_g
+ N_A2_c_223_n N_A2_M1020_g N_A2_c_224_n N_A2_M1021_g N_A2_M1023_g N_A2_c_217_n
+ A2 A2 A2 N_A2_c_219_n PM_SKY130_FD_SC_HS__O21BAI_4%A2
x_PM_SKY130_FD_SC_HS__O21BAI_4%A_828_48# N_A_828_48#_M1007_s N_A_828_48#_M1015_d
+ N_A_828_48#_M1001_g N_A_828_48#_M1002_g N_A_828_48#_c_322_n
+ N_A_828_48#_M1000_g N_A_828_48#_M1004_g N_A_828_48#_c_323_n
+ N_A_828_48#_M1024_g N_A_828_48#_M1011_g N_A_828_48#_c_317_n
+ N_A_828_48#_c_318_n N_A_828_48#_c_326_n N_A_828_48#_c_319_n
+ N_A_828_48#_c_327_n N_A_828_48#_c_328_n N_A_828_48#_c_329_n
+ N_A_828_48#_c_320_n N_A_828_48#_c_321_n PM_SKY130_FD_SC_HS__O21BAI_4%A_828_48#
x_PM_SKY130_FD_SC_HS__O21BAI_4%B1_N N_B1_N_c_433_n N_B1_N_M1015_g N_B1_N_c_430_n
+ N_B1_N_c_435_n N_B1_N_c_436_n N_B1_N_M1018_g N_B1_N_M1007_g B1_N B1_N
+ PM_SKY130_FD_SC_HS__O21BAI_4%B1_N
x_PM_SKY130_FD_SC_HS__O21BAI_4%A_28_368# N_A_28_368#_M1008_d N_A_28_368#_M1009_d
+ N_A_28_368#_M1012_d N_A_28_368#_M1017_s N_A_28_368#_M1021_s
+ N_A_28_368#_c_470_n N_A_28_368#_c_471_n N_A_28_368#_c_481_n
+ N_A_28_368#_c_472_n N_A_28_368#_c_488_n N_A_28_368#_c_473_n
+ N_A_28_368#_c_493_n N_A_28_368#_c_474_n N_A_28_368#_c_475_n
+ N_A_28_368#_c_502_n N_A_28_368#_c_476_n N_A_28_368#_c_477_n
+ N_A_28_368#_c_495_n N_A_28_368#_c_478_n PM_SKY130_FD_SC_HS__O21BAI_4%A_28_368#
x_PM_SKY130_FD_SC_HS__O21BAI_4%VPWR N_VPWR_M1008_s N_VPWR_M1010_s N_VPWR_M1000_d
+ N_VPWR_M1015_s N_VPWR_M1018_s N_VPWR_c_552_n N_VPWR_c_553_n N_VPWR_c_554_n
+ N_VPWR_c_555_n N_VPWR_c_556_n N_VPWR_c_557_n N_VPWR_c_558_n N_VPWR_c_559_n
+ VPWR N_VPWR_c_560_n N_VPWR_c_561_n N_VPWR_c_562_n N_VPWR_c_563_n
+ N_VPWR_c_564_n N_VPWR_c_565_n N_VPWR_c_566_n N_VPWR_c_551_n
+ PM_SKY130_FD_SC_HS__O21BAI_4%VPWR
x_PM_SKY130_FD_SC_HS__O21BAI_4%Y N_Y_M1001_d N_Y_M1004_d N_Y_M1014_d N_Y_M1020_d
+ N_Y_M1000_s N_Y_M1024_s N_Y_c_652_n N_Y_c_655_n N_Y_c_657_n N_Y_c_661_n
+ N_Y_c_662_n N_Y_c_645_n N_Y_c_664_n N_Y_c_646_n N_Y_c_642_n N_Y_c_643_n
+ N_Y_c_691_n N_Y_c_695_n N_Y_c_647_n N_Y_c_648_n N_Y_c_667_n N_Y_c_649_n
+ N_Y_c_650_n Y Y PM_SKY130_FD_SC_HS__O21BAI_4%Y
x_PM_SKY130_FD_SC_HS__O21BAI_4%A_27_74# N_A_27_74#_M1006_s N_A_27_74#_M1016_s
+ N_A_27_74#_M1022_s N_A_27_74#_M1005_d N_A_27_74#_M1023_d N_A_27_74#_M1002_s
+ N_A_27_74#_M1011_s N_A_27_74#_c_750_n N_A_27_74#_c_751_n N_A_27_74#_c_752_n
+ N_A_27_74#_c_753_n N_A_27_74#_c_754_n N_A_27_74#_c_755_n N_A_27_74#_c_756_n
+ N_A_27_74#_c_757_n N_A_27_74#_c_791_n N_A_27_74#_c_793_n N_A_27_74#_c_797_n
+ N_A_27_74#_c_758_n N_A_27_74#_c_759_n N_A_27_74#_c_804_n N_A_27_74#_c_760_n
+ N_A_27_74#_c_761_n N_A_27_74#_c_762_n N_A_27_74#_c_763_n N_A_27_74#_c_800_n
+ N_A_27_74#_c_764_n PM_SKY130_FD_SC_HS__O21BAI_4%A_27_74#
x_PM_SKY130_FD_SC_HS__O21BAI_4%VGND N_VGND_M1006_d N_VGND_M1019_d N_VGND_M1003_s
+ N_VGND_M1013_s N_VGND_M1007_d N_VGND_c_864_n N_VGND_c_865_n N_VGND_c_866_n
+ N_VGND_c_867_n N_VGND_c_868_n N_VGND_c_869_n N_VGND_c_870_n N_VGND_c_871_n
+ N_VGND_c_872_n N_VGND_c_873_n VGND N_VGND_c_874_n N_VGND_c_875_n
+ N_VGND_c_876_n N_VGND_c_877_n N_VGND_c_878_n N_VGND_c_879_n
+ PM_SKY130_FD_SC_HS__O21BAI_4%VGND
cc_1 VNB N_A1_M1006_g 0.0325972f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_2 VNB N_A1_M1016_g 0.0238718f $X=-0.19 $Y=-0.245 $X2=0.975 $Y2=0.74
cc_3 VNB N_A1_M1019_g 0.0224921f $X=-0.19 $Y=-0.245 $X2=1.405 $Y2=0.74
cc_4 VNB N_A1_c_129_n 0.00899086f $X=-0.19 $Y=-0.245 $X2=1.76 $Y2=1.425
cc_5 VNB N_A1_c_130_n 0.0524488f $X=-0.19 $Y=-0.245 $X2=1.5 $Y2=1.425
cc_6 VNB N_A1_M1022_g 0.0229971f $X=-0.19 $Y=-0.245 $X2=1.835 $Y2=0.74
cc_7 VNB N_A1_c_132_n 0.00808118f $X=-0.19 $Y=-0.245 $X2=1.86 $Y2=1.675
cc_8 VNB N_A1_c_133_n 0.00678907f $X=-0.19 $Y=-0.245 $X2=1.855 $Y2=1.425
cc_9 VNB A1 0.0166485f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=1.58
cc_10 VNB N_A2_M1003_g 0.0229971f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_11 VNB N_A2_c_212_n 0.00836872f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=2.4
cc_12 VNB N_A2_c_213_n 0.0118957f $X=-0.19 $Y=-0.245 $X2=0.96 $Y2=2.4
cc_13 VNB N_A2_M1005_g 0.0224931f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A2_M1013_g 0.0255099f $X=-0.19 $Y=-0.245 $X2=1.41 $Y2=2.4
cc_15 VNB N_A2_M1023_g 0.0266863f $X=-0.19 $Y=-0.245 $X2=1.86 $Y2=2.4
cc_16 VNB N_A2_c_217_n 0.00773337f $X=-0.19 $Y=-0.245 $X2=1.855 $Y2=1.425
cc_17 VNB A2 0.00177056f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.58
cc_18 VNB N_A2_c_219_n 0.0579573f $X=-0.19 $Y=-0.245 $X2=1.265 $Y2=1.515
cc_19 VNB N_A_828_48#_M1001_g 0.0224958f $X=-0.19 $Y=-0.245 $X2=0.96 $Y2=2.4
cc_20 VNB N_A_828_48#_M1002_g 0.0231786f $X=-0.19 $Y=-0.245 $X2=0.975 $Y2=0.74
cc_21 VNB N_A_828_48#_M1004_g 0.0241972f $X=-0.19 $Y=-0.245 $X2=1.41 $Y2=2.4
cc_22 VNB N_A_828_48#_M1011_g 0.0265982f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_828_48#_c_317_n 0.00283669f $X=-0.19 $Y=-0.245 $X2=1.86 $Y2=1.675
cc_24 VNB N_A_828_48#_c_318_n 0.0744266f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.58
cc_25 VNB N_A_828_48#_c_319_n 0.0180412f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_828_48#_c_320_n 0.00959788f $X=-0.19 $Y=-0.245 $X2=1.265 $Y2=1.557
cc_27 VNB N_A_828_48#_c_321_n 0.0087609f $X=-0.19 $Y=-0.245 $X2=1.265 $Y2=1.515
cc_28 VNB N_B1_N_c_430_n 0.037938f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_B1_N_M1007_g 0.0308777f $X=-0.19 $Y=-0.245 $X2=0.975 $Y2=1.35
cc_30 VNB B1_N 0.0120967f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_VPWR_c_551_n 0.302998f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_Y_c_642_n 0.0053753f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_Y_c_643_n 0.00555178f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.557
cc_34 VNB Y 0.00431708f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_27_74#_c_750_n 0.0266107f $X=-0.19 $Y=-0.245 $X2=1.835 $Y2=1.35
cc_36 VNB N_A_27_74#_c_751_n 0.0035469f $X=-0.19 $Y=-0.245 $X2=1.835 $Y2=0.74
cc_37 VNB N_A_27_74#_c_752_n 0.00998227f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_27_74#_c_753_n 0.00179819f $X=-0.19 $Y=-0.245 $X2=1.86 $Y2=1.765
cc_39 VNB N_A_27_74#_c_754_n 0.0036153f $X=-0.19 $Y=-0.245 $X2=1.86 $Y2=2.4
cc_40 VNB N_A_27_74#_c_755_n 0.00178908f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.58
cc_41 VNB N_A_27_74#_c_756_n 0.00838884f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_27_74#_c_757_n 0.00206666f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.557
cc_43 VNB N_A_27_74#_c_758_n 0.0026202f $X=-0.19 $Y=-0.245 $X2=1.405 $Y2=1.557
cc_44 VNB N_A_27_74#_c_759_n 0.00221459f $X=-0.19 $Y=-0.245 $X2=1.41 $Y2=1.557
cc_45 VNB N_A_27_74#_c_760_n 0.00882952f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.565
cc_46 VNB N_A_27_74#_c_761_n 0.00504363f $X=-0.19 $Y=-0.245 $X2=1.265 $Y2=1.565
cc_47 VNB N_A_27_74#_c_762_n 0.00127131f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_27_74#_c_763_n 0.0037103f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A_27_74#_c_764_n 0.00220733f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_VGND_c_864_n 0.00560659f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_VGND_c_865_n 0.00257504f $X=-0.19 $Y=-0.245 $X2=1.76 $Y2=1.425
cc_52 VNB N_VGND_c_866_n 0.0026136f $X=-0.19 $Y=-0.245 $X2=1.835 $Y2=0.74
cc_53 VNB N_VGND_c_867_n 0.0067113f $X=-0.19 $Y=-0.245 $X2=1.86 $Y2=1.765
cc_54 VNB N_VGND_c_868_n 0.0122168f $X=-0.19 $Y=-0.245 $X2=1.86 $Y2=2.4
cc_55 VNB N_VGND_c_869_n 0.0519799f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_56 VNB N_VGND_c_870_n 0.0151736f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=1.58
cc_57 VNB N_VGND_c_871_n 0.00604233f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_VGND_c_872_n 0.0164978f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_VGND_c_873_n 0.00631651f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_VGND_c_874_n 0.0173909f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.557
cc_61 VNB N_VGND_c_875_n 0.0169227f $X=-0.19 $Y=-0.245 $X2=1.265 $Y2=1.557
cc_62 VNB N_VGND_c_876_n 0.0760195f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_VGND_c_877_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_VGND_c_878_n 0.00604233f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_VGND_c_879_n 0.399316f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VPB N_A1_c_135_n 0.0201401f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=1.765
cc_67 VPB N_A1_c_136_n 0.0155096f $X=-0.19 $Y=1.66 $X2=0.96 $Y2=1.765
cc_68 VPB N_A1_c_137_n 0.0149991f $X=-0.19 $Y=1.66 $X2=1.41 $Y2=1.765
cc_69 VPB N_A1_c_130_n 0.0338836f $X=-0.19 $Y=1.66 $X2=1.5 $Y2=1.425
cc_70 VPB N_A1_c_132_n 7.1155e-19 $X=-0.19 $Y=1.66 $X2=1.86 $Y2=1.675
cc_71 VPB N_A1_c_140_n 0.0207175f $X=-0.19 $Y=1.66 $X2=1.86 $Y2=1.765
cc_72 VPB A1 0.016639f $X=-0.19 $Y=1.66 $X2=1.595 $Y2=1.58
cc_73 VPB N_A2_c_212_n 7.36868e-19 $X=-0.19 $Y=1.66 $X2=0.51 $Y2=2.4
cc_74 VPB N_A2_c_221_n 0.0210455f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=2.4
cc_75 VPB N_A2_c_222_n 0.014659f $X=-0.19 $Y=1.66 $X2=1.405 $Y2=0.74
cc_76 VPB N_A2_c_223_n 0.0150423f $X=-0.19 $Y=1.66 $X2=1.5 $Y2=1.425
cc_77 VPB N_A2_c_224_n 0.0174657f $X=-0.19 $Y=1.66 $X2=1.835 $Y2=0.74
cc_78 VPB A2 0.0088718f $X=-0.19 $Y=1.66 $X2=1.115 $Y2=1.58
cc_79 VPB N_A2_c_219_n 0.0365322f $X=-0.19 $Y=1.66 $X2=1.265 $Y2=1.515
cc_80 VPB N_A_828_48#_c_322_n 0.0181691f $X=-0.19 $Y=1.66 $X2=1.405 $Y2=1.35
cc_81 VPB N_A_828_48#_c_323_n 0.0179703f $X=-0.19 $Y=1.66 $X2=1.76 $Y2=1.425
cc_82 VPB N_A_828_48#_c_317_n 0.00283634f $X=-0.19 $Y=1.66 $X2=1.86 $Y2=1.675
cc_83 VPB N_A_828_48#_c_318_n 0.0509309f $X=-0.19 $Y=1.66 $X2=1.115 $Y2=1.58
cc_84 VPB N_A_828_48#_c_326_n 0.00626665f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_85 VPB N_A_828_48#_c_327_n 0.0103868f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_86 VPB N_A_828_48#_c_328_n 0.0049253f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.557
cc_87 VPB N_A_828_48#_c_329_n 0.00216998f $X=-0.19 $Y=1.66 $X2=0.585 $Y2=1.515
cc_88 VPB N_A_828_48#_c_321_n 2.491e-19 $X=-0.19 $Y=1.66 $X2=1.265 $Y2=1.515
cc_89 VPB N_B1_N_c_433_n 0.0165532f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.35
cc_90 VPB N_B1_N_c_430_n 0.0339388f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_91 VPB N_B1_N_c_435_n 0.0144837f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=1.765
cc_92 VPB N_B1_N_c_436_n 0.0274192f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=2.4
cc_93 VPB B1_N 0.00880174f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_94 VPB N_A_28_368#_c_470_n 0.00739392f $X=-0.19 $Y=1.66 $X2=1.405 $Y2=0.74
cc_95 VPB N_A_28_368#_c_471_n 0.0339313f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_96 VPB N_A_28_368#_c_472_n 0.00216998f $X=-0.19 $Y=1.66 $X2=1.835 $Y2=1.35
cc_97 VPB N_A_28_368#_c_473_n 0.00328381f $X=-0.19 $Y=1.66 $X2=1.86 $Y2=1.5
cc_98 VPB N_A_28_368#_c_474_n 0.00259172f $X=-0.19 $Y=1.66 $X2=1.86 $Y2=2.4
cc_99 VPB N_A_28_368#_c_475_n 0.00218844f $X=-0.19 $Y=1.66 $X2=1.855 $Y2=1.425
cc_100 VPB N_A_28_368#_c_476_n 0.00808706f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_101 VPB N_A_28_368#_c_477_n 0.00561874f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.557
cc_102 VPB N_A_28_368#_c_478_n 0.0021839f $X=-0.19 $Y=1.66 $X2=1.265 $Y2=1.515
cc_103 VPB N_VPWR_c_552_n 0.00501395f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_104 VPB N_VPWR_c_553_n 0.00339119f $X=-0.19 $Y=1.66 $X2=1.76 $Y2=1.425
cc_105 VPB N_VPWR_c_554_n 0.0080007f $X=-0.19 $Y=1.66 $X2=1.835 $Y2=0.74
cc_106 VPB N_VPWR_c_555_n 0.0148531f $X=-0.19 $Y=1.66 $X2=1.86 $Y2=1.765
cc_107 VPB N_VPWR_c_556_n 0.0120106f $X=-0.19 $Y=1.66 $X2=1.86 $Y2=2.4
cc_108 VPB N_VPWR_c_557_n 0.0462325f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_109 VPB N_VPWR_c_558_n 0.0753895f $X=-0.19 $Y=1.66 $X2=1.595 $Y2=1.58
cc_110 VPB N_VPWR_c_559_n 0.00324402f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_111 VPB N_VPWR_c_560_n 0.0181665f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_112 VPB N_VPWR_c_561_n 0.0185253f $X=-0.19 $Y=1.66 $X2=0.585 $Y2=1.515
cc_113 VPB N_VPWR_c_562_n 0.0220105f $X=-0.19 $Y=1.66 $X2=0.72 $Y2=1.565
cc_114 VPB N_VPWR_c_563_n 0.0185253f $X=-0.19 $Y=1.66 $X2=1.265 $Y2=1.565
cc_115 VPB N_VPWR_c_564_n 0.00460249f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_116 VPB N_VPWR_c_565_n 0.00601644f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_117 VPB N_VPWR_c_566_n 0.0047828f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_118 VPB N_VPWR_c_551_n 0.108437f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_119 VPB N_Y_c_645_n 0.0092968f $X=-0.19 $Y=1.66 $X2=1.86 $Y2=2.4
cc_120 VPB N_Y_c_646_n 0.0117037f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_121 VPB N_Y_c_647_n 0.00149646f $X=-0.19 $Y=1.66 $X2=1.265 $Y2=1.557
cc_122 VPB N_Y_c_648_n 0.0122846f $X=-0.19 $Y=1.66 $X2=1.265 $Y2=1.515
cc_123 VPB N_Y_c_649_n 0.00246023f $X=-0.19 $Y=1.66 $X2=1.265 $Y2=1.565
cc_124 VPB N_Y_c_650_n 8.72966e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_125 VPB Y 0.00441084f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_126 N_A1_M1022_g N_A2_M1003_g 0.0190355f $X=1.835 $Y=0.74 $X2=0 $Y2=0
cc_127 N_A1_c_132_n N_A2_c_212_n 0.00595825f $X=1.86 $Y=1.675 $X2=0 $Y2=0
cc_128 A1 N_A2_c_212_n 0.00122929f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_129 N_A1_c_140_n N_A2_c_221_n 0.0154873f $X=1.86 $Y=1.765 $X2=0 $Y2=0
cc_130 N_A1_c_133_n N_A2_c_217_n 0.00964075f $X=1.855 $Y=1.425 $X2=0 $Y2=0
cc_131 A1 N_A2_c_217_n 8.12898e-19 $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_132 N_A1_c_133_n A2 5.93133e-19 $X=1.855 $Y=1.425 $X2=0 $Y2=0
cc_133 A1 N_A_28_368#_c_470_n 0.021684f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_134 N_A1_c_135_n N_A_28_368#_c_471_n 0.00460488f $X=0.51 $Y=1.765 $X2=0 $Y2=0
cc_135 N_A1_c_135_n N_A_28_368#_c_481_n 0.0126853f $X=0.51 $Y=1.765 $X2=0 $Y2=0
cc_136 N_A1_c_136_n N_A_28_368#_c_481_n 0.0120074f $X=0.96 $Y=1.765 $X2=0 $Y2=0
cc_137 N_A1_c_130_n N_A_28_368#_c_481_n 0.00131212f $X=1.5 $Y=1.425 $X2=0 $Y2=0
cc_138 A1 N_A_28_368#_c_481_n 0.0435529f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_139 N_A1_c_135_n N_A_28_368#_c_472_n 6.71799e-19 $X=0.51 $Y=1.765 $X2=0 $Y2=0
cc_140 N_A1_c_136_n N_A_28_368#_c_472_n 0.0106363f $X=0.96 $Y=1.765 $X2=0 $Y2=0
cc_141 N_A1_c_137_n N_A_28_368#_c_472_n 0.00612298f $X=1.41 $Y=1.765 $X2=0 $Y2=0
cc_142 N_A1_c_137_n N_A_28_368#_c_488_n 0.0126342f $X=1.41 $Y=1.765 $X2=0 $Y2=0
cc_143 N_A1_c_129_n N_A_28_368#_c_488_n 3.44942e-19 $X=1.76 $Y=1.425 $X2=0 $Y2=0
cc_144 N_A1_c_140_n N_A_28_368#_c_488_n 0.0168336f $X=1.86 $Y=1.765 $X2=0 $Y2=0
cc_145 A1 N_A_28_368#_c_488_n 0.0344665f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_146 N_A1_c_140_n N_A_28_368#_c_473_n 0.00262483f $X=1.86 $Y=1.765 $X2=0 $Y2=0
cc_147 N_A1_c_140_n N_A_28_368#_c_493_n 0.00544145f $X=1.86 $Y=1.765 $X2=0 $Y2=0
cc_148 N_A1_c_140_n N_A_28_368#_c_475_n 0.00125031f $X=1.86 $Y=1.765 $X2=0 $Y2=0
cc_149 N_A1_c_136_n N_A_28_368#_c_495_n 4.27055e-19 $X=0.96 $Y=1.765 $X2=0 $Y2=0
cc_150 N_A1_c_130_n N_A_28_368#_c_495_n 0.00124229f $X=1.5 $Y=1.425 $X2=0 $Y2=0
cc_151 A1 N_A_28_368#_c_495_n 0.0193936f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_152 N_A1_c_135_n N_VPWR_c_552_n 0.0135832f $X=0.51 $Y=1.765 $X2=0 $Y2=0
cc_153 N_A1_c_136_n N_VPWR_c_552_n 0.00395359f $X=0.96 $Y=1.765 $X2=0 $Y2=0
cc_154 N_A1_c_136_n N_VPWR_c_553_n 5.55114e-19 $X=0.96 $Y=1.765 $X2=0 $Y2=0
cc_155 N_A1_c_137_n N_VPWR_c_553_n 0.0111578f $X=1.41 $Y=1.765 $X2=0 $Y2=0
cc_156 N_A1_c_140_n N_VPWR_c_553_n 0.0102886f $X=1.86 $Y=1.765 $X2=0 $Y2=0
cc_157 N_A1_c_140_n N_VPWR_c_558_n 0.00413917f $X=1.86 $Y=1.765 $X2=0 $Y2=0
cc_158 N_A1_c_135_n N_VPWR_c_560_n 0.00413917f $X=0.51 $Y=1.765 $X2=0 $Y2=0
cc_159 N_A1_c_136_n N_VPWR_c_561_n 0.00445602f $X=0.96 $Y=1.765 $X2=0 $Y2=0
cc_160 N_A1_c_137_n N_VPWR_c_561_n 0.00413917f $X=1.41 $Y=1.765 $X2=0 $Y2=0
cc_161 N_A1_c_135_n N_VPWR_c_551_n 0.00821237f $X=0.51 $Y=1.765 $X2=0 $Y2=0
cc_162 N_A1_c_136_n N_VPWR_c_551_n 0.00857589f $X=0.96 $Y=1.765 $X2=0 $Y2=0
cc_163 N_A1_c_137_n N_VPWR_c_551_n 0.00817726f $X=1.41 $Y=1.765 $X2=0 $Y2=0
cc_164 N_A1_c_140_n N_VPWR_c_551_n 0.0081781f $X=1.86 $Y=1.765 $X2=0 $Y2=0
cc_165 N_A1_M1006_g N_A_27_74#_c_750_n 0.00159319f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_166 N_A1_M1006_g N_A_27_74#_c_751_n 0.0139418f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_167 N_A1_M1016_g N_A_27_74#_c_751_n 0.0141141f $X=0.975 $Y=0.74 $X2=0 $Y2=0
cc_168 N_A1_c_130_n N_A_27_74#_c_751_n 0.00336308f $X=1.5 $Y=1.425 $X2=0 $Y2=0
cc_169 A1 N_A_27_74#_c_751_n 0.055804f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_170 A1 N_A_27_74#_c_752_n 0.0216404f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_171 N_A1_M1016_g N_A_27_74#_c_753_n 4.06088e-19 $X=0.975 $Y=0.74 $X2=0 $Y2=0
cc_172 N_A1_M1019_g N_A_27_74#_c_753_n 3.92313e-19 $X=1.405 $Y=0.74 $X2=0 $Y2=0
cc_173 N_A1_M1019_g N_A_27_74#_c_754_n 0.0130918f $X=1.405 $Y=0.74 $X2=0 $Y2=0
cc_174 N_A1_c_129_n N_A_27_74#_c_754_n 0.00205448f $X=1.76 $Y=1.425 $X2=0 $Y2=0
cc_175 N_A1_M1022_g N_A_27_74#_c_754_n 0.0165853f $X=1.835 $Y=0.74 $X2=0 $Y2=0
cc_176 N_A1_c_133_n N_A_27_74#_c_754_n 0.00161743f $X=1.855 $Y=1.425 $X2=0 $Y2=0
cc_177 A1 N_A_27_74#_c_754_n 0.0390831f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_178 N_A1_M1022_g N_A_27_74#_c_755_n 3.92313e-19 $X=1.835 $Y=0.74 $X2=0 $Y2=0
cc_179 N_A1_c_130_n N_A_27_74#_c_762_n 0.00232957f $X=1.5 $Y=1.425 $X2=0 $Y2=0
cc_180 A1 N_A_27_74#_c_762_n 0.0146029f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_181 N_A1_M1006_g N_VGND_c_864_n 0.0136336f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_182 N_A1_M1016_g N_VGND_c_864_n 0.00238967f $X=0.975 $Y=0.74 $X2=0 $Y2=0
cc_183 N_A1_M1016_g N_VGND_c_865_n 4.78723e-19 $X=0.975 $Y=0.74 $X2=0 $Y2=0
cc_184 N_A1_M1019_g N_VGND_c_865_n 0.010763f $X=1.405 $Y=0.74 $X2=0 $Y2=0
cc_185 N_A1_M1022_g N_VGND_c_865_n 0.0106755f $X=1.835 $Y=0.74 $X2=0 $Y2=0
cc_186 N_A1_M1022_g N_VGND_c_866_n 4.71636e-19 $X=1.835 $Y=0.74 $X2=0 $Y2=0
cc_187 N_A1_M1022_g N_VGND_c_870_n 0.00383152f $X=1.835 $Y=0.74 $X2=0 $Y2=0
cc_188 N_A1_M1006_g N_VGND_c_874_n 0.00383152f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_189 N_A1_M1016_g N_VGND_c_875_n 0.00461464f $X=0.975 $Y=0.74 $X2=0 $Y2=0
cc_190 N_A1_M1019_g N_VGND_c_875_n 0.00383152f $X=1.405 $Y=0.74 $X2=0 $Y2=0
cc_191 N_A1_M1006_g N_VGND_c_879_n 0.00761198f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_192 N_A1_M1016_g N_VGND_c_879_n 0.0090814f $X=0.975 $Y=0.74 $X2=0 $Y2=0
cc_193 N_A1_M1019_g N_VGND_c_879_n 0.0075754f $X=1.405 $Y=0.74 $X2=0 $Y2=0
cc_194 N_A1_M1022_g N_VGND_c_879_n 0.00757637f $X=1.835 $Y=0.74 $X2=0 $Y2=0
cc_195 N_A2_M1023_g N_A_828_48#_M1001_g 0.0166348f $X=3.715 $Y=0.74 $X2=0 $Y2=0
cc_196 A2 N_A_828_48#_c_318_n 2.88328e-19 $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_197 N_A2_c_219_n N_A_828_48#_c_318_n 0.0229362f $X=3.71 $Y=1.557 $X2=0 $Y2=0
cc_198 N_A2_c_221_n N_A_28_368#_c_473_n 0.00336699f $X=2.31 $Y=1.765 $X2=0 $Y2=0
cc_199 N_A2_c_221_n N_A_28_368#_c_493_n 0.00358597f $X=2.31 $Y=1.765 $X2=0 $Y2=0
cc_200 N_A2_c_221_n N_A_28_368#_c_474_n 0.012504f $X=2.31 $Y=1.765 $X2=0 $Y2=0
cc_201 N_A2_c_222_n N_A_28_368#_c_474_n 0.0107904f $X=2.76 $Y=1.765 $X2=0 $Y2=0
cc_202 N_A2_c_221_n N_A_28_368#_c_502_n 6.2388e-19 $X=2.31 $Y=1.765 $X2=0 $Y2=0
cc_203 N_A2_c_222_n N_A_28_368#_c_502_n 0.00786706f $X=2.76 $Y=1.765 $X2=0 $Y2=0
cc_204 N_A2_c_223_n N_A_28_368#_c_502_n 0.00769091f $X=3.21 $Y=1.765 $X2=0 $Y2=0
cc_205 N_A2_c_224_n N_A_28_368#_c_502_n 5.94863e-19 $X=3.71 $Y=1.765 $X2=0 $Y2=0
cc_206 N_A2_c_223_n N_A_28_368#_c_476_n 0.0111147f $X=3.21 $Y=1.765 $X2=0 $Y2=0
cc_207 N_A2_c_224_n N_A_28_368#_c_476_n 0.0152643f $X=3.71 $Y=1.765 $X2=0 $Y2=0
cc_208 N_A2_c_222_n N_A_28_368#_c_478_n 0.00175197f $X=2.76 $Y=1.765 $X2=0 $Y2=0
cc_209 N_A2_c_223_n N_A_28_368#_c_478_n 0.00175197f $X=3.21 $Y=1.765 $X2=0 $Y2=0
cc_210 N_A2_c_221_n N_VPWR_c_558_n 0.00278271f $X=2.31 $Y=1.765 $X2=0 $Y2=0
cc_211 N_A2_c_222_n N_VPWR_c_558_n 0.00278257f $X=2.76 $Y=1.765 $X2=0 $Y2=0
cc_212 N_A2_c_223_n N_VPWR_c_558_n 0.00278257f $X=3.21 $Y=1.765 $X2=0 $Y2=0
cc_213 N_A2_c_224_n N_VPWR_c_558_n 0.00278271f $X=3.71 $Y=1.765 $X2=0 $Y2=0
cc_214 N_A2_c_221_n N_VPWR_c_551_n 0.00353907f $X=2.31 $Y=1.765 $X2=0 $Y2=0
cc_215 N_A2_c_222_n N_VPWR_c_551_n 0.00353822f $X=2.76 $Y=1.765 $X2=0 $Y2=0
cc_216 N_A2_c_223_n N_VPWR_c_551_n 0.00354283f $X=3.21 $Y=1.765 $X2=0 $Y2=0
cc_217 N_A2_c_224_n N_VPWR_c_551_n 0.00359085f $X=3.71 $Y=1.765 $X2=0 $Y2=0
cc_218 N_A2_c_221_n N_Y_c_652_n 0.00243806f $X=2.31 $Y=1.765 $X2=0 $Y2=0
cc_219 N_A2_c_213_n N_Y_c_652_n 0.00361586f $X=2.62 $Y=1.425 $X2=0 $Y2=0
cc_220 A2 N_Y_c_652_n 0.00839776f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_221 N_A2_c_221_n N_Y_c_655_n 0.00783806f $X=2.31 $Y=1.765 $X2=0 $Y2=0
cc_222 N_A2_c_222_n N_Y_c_655_n 0.00576017f $X=2.76 $Y=1.765 $X2=0 $Y2=0
cc_223 N_A2_c_222_n N_Y_c_657_n 0.0126853f $X=2.76 $Y=1.765 $X2=0 $Y2=0
cc_224 N_A2_c_223_n N_Y_c_657_n 0.0151589f $X=3.21 $Y=1.765 $X2=0 $Y2=0
cc_225 A2 N_Y_c_657_n 0.0461979f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_226 N_A2_c_219_n N_Y_c_657_n 0.00150005f $X=3.71 $Y=1.557 $X2=0 $Y2=0
cc_227 N_A2_c_224_n N_Y_c_661_n 0.0135833f $X=3.71 $Y=1.765 $X2=0 $Y2=0
cc_228 N_A2_c_224_n N_Y_c_662_n 0.0160658f $X=3.71 $Y=1.765 $X2=0 $Y2=0
cc_229 A2 N_Y_c_662_n 0.00470872f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_230 N_A2_M1023_g N_Y_c_664_n 8.84124e-19 $X=3.715 $Y=0.74 $X2=0 $Y2=0
cc_231 N_A2_c_224_n N_Y_c_646_n 0.00528409f $X=3.71 $Y=1.765 $X2=0 $Y2=0
cc_232 N_A2_M1023_g N_Y_c_643_n 0.00472032f $X=3.715 $Y=0.74 $X2=0 $Y2=0
cc_233 N_A2_c_224_n N_Y_c_667_n 4.27055e-19 $X=3.71 $Y=1.765 $X2=0 $Y2=0
cc_234 A2 N_Y_c_667_n 0.025478f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_235 N_A2_c_219_n N_Y_c_667_n 0.00168378f $X=3.71 $Y=1.557 $X2=0 $Y2=0
cc_236 N_A2_c_224_n Y 0.00624786f $X=3.71 $Y=1.765 $X2=0 $Y2=0
cc_237 N_A2_M1023_g Y 0.00519773f $X=3.715 $Y=0.74 $X2=0 $Y2=0
cc_238 A2 Y 0.0261148f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_239 N_A2_c_219_n Y 0.00342721f $X=3.71 $Y=1.557 $X2=0 $Y2=0
cc_240 N_A2_M1003_g N_A_27_74#_c_755_n 3.92313e-19 $X=2.265 $Y=0.74 $X2=0 $Y2=0
cc_241 N_A2_M1003_g N_A_27_74#_c_756_n 0.0175066f $X=2.265 $Y=0.74 $X2=0 $Y2=0
cc_242 N_A2_c_213_n N_A_27_74#_c_756_n 0.00334794f $X=2.62 $Y=1.425 $X2=0 $Y2=0
cc_243 N_A2_M1005_g N_A_27_74#_c_756_n 0.0130918f $X=2.695 $Y=0.74 $X2=0 $Y2=0
cc_244 N_A2_M1013_g N_A_27_74#_c_756_n 0.00499651f $X=3.125 $Y=0.74 $X2=0 $Y2=0
cc_245 N_A2_M1023_g N_A_27_74#_c_756_n 7.62044e-19 $X=3.715 $Y=0.74 $X2=0 $Y2=0
cc_246 A2 N_A_27_74#_c_756_n 0.0437388f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_247 N_A2_c_219_n N_A_27_74#_c_756_n 0.00232957f $X=3.71 $Y=1.557 $X2=0 $Y2=0
cc_248 N_A2_M1013_g N_A_27_74#_c_757_n 0.00538884f $X=3.125 $Y=0.74 $X2=0 $Y2=0
cc_249 N_A2_M1023_g N_A_27_74#_c_757_n 7.98198e-19 $X=3.715 $Y=0.74 $X2=0 $Y2=0
cc_250 N_A2_M1013_g N_A_27_74#_c_791_n 0.00337163f $X=3.125 $Y=0.74 $X2=0 $Y2=0
cc_251 N_A2_M1023_g N_A_27_74#_c_791_n 7.65889e-19 $X=3.715 $Y=0.74 $X2=0 $Y2=0
cc_252 N_A2_M1013_g N_A_27_74#_c_793_n 0.0106833f $X=3.125 $Y=0.74 $X2=0 $Y2=0
cc_253 N_A2_M1023_g N_A_27_74#_c_793_n 0.0138896f $X=3.715 $Y=0.74 $X2=0 $Y2=0
cc_254 A2 N_A_27_74#_c_793_n 0.018191f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_255 N_A2_c_219_n N_A_27_74#_c_793_n 0.00451439f $X=3.71 $Y=1.557 $X2=0 $Y2=0
cc_256 N_A2_M1013_g N_A_27_74#_c_797_n 7.80342e-19 $X=3.125 $Y=0.74 $X2=0 $Y2=0
cc_257 N_A2_M1023_g N_A_27_74#_c_797_n 0.0042743f $X=3.715 $Y=0.74 $X2=0 $Y2=0
cc_258 N_A2_M1023_g N_A_27_74#_c_759_n 0.00396171f $X=3.715 $Y=0.74 $X2=0 $Y2=0
cc_259 N_A2_M1013_g N_A_27_74#_c_800_n 9.34275e-19 $X=3.125 $Y=0.74 $X2=0 $Y2=0
cc_260 N_A2_M1003_g N_VGND_c_865_n 4.71636e-19 $X=2.265 $Y=0.74 $X2=0 $Y2=0
cc_261 N_A2_M1003_g N_VGND_c_866_n 0.0106755f $X=2.265 $Y=0.74 $X2=0 $Y2=0
cc_262 N_A2_M1005_g N_VGND_c_866_n 0.0108006f $X=2.695 $Y=0.74 $X2=0 $Y2=0
cc_263 N_A2_M1013_g N_VGND_c_866_n 5.18931e-19 $X=3.125 $Y=0.74 $X2=0 $Y2=0
cc_264 N_A2_M1013_g N_VGND_c_867_n 0.00271269f $X=3.125 $Y=0.74 $X2=0 $Y2=0
cc_265 N_A2_M1023_g N_VGND_c_867_n 0.00231005f $X=3.715 $Y=0.74 $X2=0 $Y2=0
cc_266 N_A2_M1003_g N_VGND_c_870_n 0.00383152f $X=2.265 $Y=0.74 $X2=0 $Y2=0
cc_267 N_A2_M1005_g N_VGND_c_872_n 0.00383152f $X=2.695 $Y=0.74 $X2=0 $Y2=0
cc_268 N_A2_M1013_g N_VGND_c_872_n 0.00324657f $X=3.125 $Y=0.74 $X2=0 $Y2=0
cc_269 N_A2_M1023_g N_VGND_c_876_n 0.00321293f $X=3.715 $Y=0.74 $X2=0 $Y2=0
cc_270 N_A2_M1003_g N_VGND_c_879_n 0.00757637f $X=2.265 $Y=0.74 $X2=0 $Y2=0
cc_271 N_A2_M1005_g N_VGND_c_879_n 0.0075754f $X=2.695 $Y=0.74 $X2=0 $Y2=0
cc_272 N_A2_M1013_g N_VGND_c_879_n 0.0041114f $X=3.125 $Y=0.74 $X2=0 $Y2=0
cc_273 N_A2_M1023_g N_VGND_c_879_n 0.00411864f $X=3.715 $Y=0.74 $X2=0 $Y2=0
cc_274 N_A_828_48#_c_327_n N_B1_N_c_433_n 0.00920906f $X=6.305 $Y=2.035
+ $X2=-0.19 $Y2=-0.245
cc_275 N_A_828_48#_c_329_n N_B1_N_c_433_n 0.01627f $X=6.47 $Y=2.265 $X2=-0.19
+ $Y2=-0.245
cc_276 N_A_828_48#_c_318_n N_B1_N_c_430_n 0.00501947f $X=5.555 $Y=1.515 $X2=0
+ $Y2=0
cc_277 N_A_828_48#_c_326_n N_B1_N_c_430_n 0.00579843f $X=5.88 $Y=1.95 $X2=0
+ $Y2=0
cc_278 N_A_828_48#_c_319_n N_B1_N_c_430_n 0.0116688f $X=6.325 $Y=1.195 $X2=0
+ $Y2=0
cc_279 N_A_828_48#_c_327_n N_B1_N_c_430_n 0.011591f $X=6.305 $Y=2.035 $X2=0
+ $Y2=0
cc_280 N_A_828_48#_c_321_n N_B1_N_c_430_n 0.00511237f $X=5.88 $Y=1.195 $X2=0
+ $Y2=0
cc_281 N_A_828_48#_c_327_n N_B1_N_c_435_n 0.00302426f $X=6.305 $Y=2.035 $X2=0
+ $Y2=0
cc_282 N_A_828_48#_c_327_n N_B1_N_c_436_n 0.00190445f $X=6.305 $Y=2.035 $X2=0
+ $Y2=0
cc_283 N_A_828_48#_c_329_n N_B1_N_c_436_n 0.0037498f $X=6.47 $Y=2.265 $X2=0
+ $Y2=0
cc_284 N_A_828_48#_c_319_n N_B1_N_M1007_g 4.58098e-19 $X=6.325 $Y=1.195 $X2=0
+ $Y2=0
cc_285 N_A_828_48#_c_320_n N_B1_N_M1007_g 0.00159319f $X=6.49 $Y=0.665 $X2=0
+ $Y2=0
cc_286 N_A_828_48#_c_321_n N_B1_N_M1007_g 0.00350542f $X=5.88 $Y=1.195 $X2=0
+ $Y2=0
cc_287 N_A_828_48#_c_319_n B1_N 0.01771f $X=6.325 $Y=1.195 $X2=0 $Y2=0
cc_288 N_A_828_48#_c_327_n B1_N 0.0160253f $X=6.305 $Y=2.035 $X2=0 $Y2=0
cc_289 N_A_828_48#_c_321_n B1_N 0.0137688f $X=5.88 $Y=1.195 $X2=0 $Y2=0
cc_290 N_A_828_48#_c_322_n N_A_28_368#_c_476_n 0.00283598f $X=4.77 $Y=1.765
+ $X2=0 $Y2=0
cc_291 N_A_828_48#_c_322_n N_A_28_368#_c_477_n 0.00106959f $X=4.77 $Y=1.765
+ $X2=0 $Y2=0
cc_292 N_A_828_48#_c_328_n N_VPWR_M1015_s 9.95962e-19 $X=5.965 $Y=2.035 $X2=0
+ $Y2=0
cc_293 N_A_828_48#_c_322_n N_VPWR_c_554_n 0.00552619f $X=4.77 $Y=1.765 $X2=0
+ $Y2=0
cc_294 N_A_828_48#_c_323_n N_VPWR_c_554_n 0.0055495f $X=5.235 $Y=1.765 $X2=0
+ $Y2=0
cc_295 N_A_828_48#_c_323_n N_VPWR_c_555_n 0.00378606f $X=5.235 $Y=1.765 $X2=0
+ $Y2=0
cc_296 N_A_828_48#_c_327_n N_VPWR_c_555_n 0.0114561f $X=6.305 $Y=2.035 $X2=0
+ $Y2=0
cc_297 N_A_828_48#_c_328_n N_VPWR_c_555_n 0.00989481f $X=5.965 $Y=2.035 $X2=0
+ $Y2=0
cc_298 N_A_828_48#_c_329_n N_VPWR_c_555_n 0.0453479f $X=6.47 $Y=2.265 $X2=0
+ $Y2=0
cc_299 N_A_828_48#_c_327_n N_VPWR_c_557_n 0.00149263f $X=6.305 $Y=2.035 $X2=0
+ $Y2=0
cc_300 N_A_828_48#_c_329_n N_VPWR_c_557_n 0.0576594f $X=6.47 $Y=2.265 $X2=0
+ $Y2=0
cc_301 N_A_828_48#_c_322_n N_VPWR_c_558_n 0.00445602f $X=4.77 $Y=1.765 $X2=0
+ $Y2=0
cc_302 N_A_828_48#_c_323_n N_VPWR_c_562_n 0.00445602f $X=5.235 $Y=1.765 $X2=0
+ $Y2=0
cc_303 N_A_828_48#_c_329_n N_VPWR_c_563_n 0.0110241f $X=6.47 $Y=2.265 $X2=0
+ $Y2=0
cc_304 N_A_828_48#_c_322_n N_VPWR_c_551_n 0.00862534f $X=4.77 $Y=1.765 $X2=0
+ $Y2=0
cc_305 N_A_828_48#_c_323_n N_VPWR_c_551_n 0.0086287f $X=5.235 $Y=1.765 $X2=0
+ $Y2=0
cc_306 N_A_828_48#_c_329_n N_VPWR_c_551_n 0.00909194f $X=6.47 $Y=2.265 $X2=0
+ $Y2=0
cc_307 N_A_828_48#_c_317_n N_Y_c_645_n 5.04769e-19 $X=5.795 $Y=1.515 $X2=0 $Y2=0
cc_308 N_A_828_48#_c_318_n N_Y_c_645_n 0.00675205f $X=5.555 $Y=1.515 $X2=0 $Y2=0
cc_309 N_A_828_48#_M1001_g N_Y_c_664_n 0.00661629f $X=4.215 $Y=0.74 $X2=0 $Y2=0
cc_310 N_A_828_48#_M1002_g N_Y_c_664_n 0.00673482f $X=4.645 $Y=0.74 $X2=0 $Y2=0
cc_311 N_A_828_48#_M1004_g N_Y_c_664_n 5.96216e-19 $X=5.145 $Y=0.74 $X2=0 $Y2=0
cc_312 N_A_828_48#_c_322_n N_Y_c_646_n 0.0102048f $X=4.77 $Y=1.765 $X2=0 $Y2=0
cc_313 N_A_828_48#_c_323_n N_Y_c_646_n 3.7226e-19 $X=5.235 $Y=1.765 $X2=0 $Y2=0
cc_314 N_A_828_48#_M1002_g N_Y_c_642_n 0.0093986f $X=4.645 $Y=0.74 $X2=0 $Y2=0
cc_315 N_A_828_48#_M1004_g N_Y_c_642_n 0.0129058f $X=5.145 $Y=0.74 $X2=0 $Y2=0
cc_316 N_A_828_48#_M1011_g N_Y_c_642_n 0.00764453f $X=5.645 $Y=0.74 $X2=0 $Y2=0
cc_317 N_A_828_48#_c_317_n N_Y_c_642_n 0.0273799f $X=5.795 $Y=1.515 $X2=0 $Y2=0
cc_318 N_A_828_48#_c_318_n N_Y_c_642_n 0.00791827f $X=5.555 $Y=1.515 $X2=0 $Y2=0
cc_319 N_A_828_48#_c_321_n N_Y_c_642_n 0.00494448f $X=5.88 $Y=1.195 $X2=0 $Y2=0
cc_320 N_A_828_48#_M1001_g N_Y_c_643_n 0.0135802f $X=4.215 $Y=0.74 $X2=0 $Y2=0
cc_321 N_A_828_48#_M1002_g N_Y_c_643_n 0.00272319f $X=4.645 $Y=0.74 $X2=0 $Y2=0
cc_322 N_A_828_48#_c_317_n N_Y_c_643_n 0.0660757f $X=5.795 $Y=1.515 $X2=0 $Y2=0
cc_323 N_A_828_48#_c_318_n N_Y_c_643_n 0.00224206f $X=5.555 $Y=1.515 $X2=0 $Y2=0
cc_324 N_A_828_48#_c_322_n N_Y_c_691_n 0.0120932f $X=4.77 $Y=1.765 $X2=0 $Y2=0
cc_325 N_A_828_48#_c_323_n N_Y_c_691_n 0.0120932f $X=5.235 $Y=1.765 $X2=0 $Y2=0
cc_326 N_A_828_48#_c_317_n N_Y_c_691_n 0.0383325f $X=5.795 $Y=1.515 $X2=0 $Y2=0
cc_327 N_A_828_48#_c_318_n N_Y_c_691_n 0.00685566f $X=5.555 $Y=1.515 $X2=0 $Y2=0
cc_328 N_A_828_48#_M1011_g N_Y_c_695_n 0.00785289f $X=5.645 $Y=0.74 $X2=0 $Y2=0
cc_329 N_A_828_48#_c_323_n N_Y_c_647_n 4.27055e-19 $X=5.235 $Y=1.765 $X2=0 $Y2=0
cc_330 N_A_828_48#_c_317_n N_Y_c_647_n 0.024645f $X=5.795 $Y=1.515 $X2=0 $Y2=0
cc_331 N_A_828_48#_c_318_n N_Y_c_647_n 0.00743262f $X=5.555 $Y=1.515 $X2=0 $Y2=0
cc_332 N_A_828_48#_c_326_n N_Y_c_647_n 0.00840812f $X=5.88 $Y=1.95 $X2=0 $Y2=0
cc_333 N_A_828_48#_c_328_n N_Y_c_647_n 0.00655874f $X=5.965 $Y=2.035 $X2=0 $Y2=0
cc_334 N_A_828_48#_c_322_n N_Y_c_648_n 6.86372e-19 $X=4.77 $Y=1.765 $X2=0 $Y2=0
cc_335 N_A_828_48#_c_323_n N_Y_c_648_n 0.0122629f $X=5.235 $Y=1.765 $X2=0 $Y2=0
cc_336 N_A_828_48#_c_328_n N_Y_c_648_n 0.00880422f $X=5.965 $Y=2.035 $X2=0 $Y2=0
cc_337 N_A_828_48#_c_322_n N_Y_c_650_n 0.00221578f $X=4.77 $Y=1.765 $X2=0 $Y2=0
cc_338 N_A_828_48#_c_323_n N_Y_c_650_n 2.97171e-19 $X=5.235 $Y=1.765 $X2=0 $Y2=0
cc_339 N_A_828_48#_c_317_n N_Y_c_650_n 0.024645f $X=5.795 $Y=1.515 $X2=0 $Y2=0
cc_340 N_A_828_48#_c_318_n N_Y_c_650_n 0.00764955f $X=5.555 $Y=1.515 $X2=0 $Y2=0
cc_341 N_A_828_48#_M1001_g Y 0.00515227f $X=4.215 $Y=0.74 $X2=0 $Y2=0
cc_342 N_A_828_48#_M1002_g Y 8.76782e-19 $X=4.645 $Y=0.74 $X2=0 $Y2=0
cc_343 N_A_828_48#_c_322_n Y 0.00200263f $X=4.77 $Y=1.765 $X2=0 $Y2=0
cc_344 N_A_828_48#_c_317_n Y 0.0249266f $X=5.795 $Y=1.515 $X2=0 $Y2=0
cc_345 N_A_828_48#_c_318_n Y 0.0127709f $X=5.555 $Y=1.515 $X2=0 $Y2=0
cc_346 N_A_828_48#_c_321_n N_A_27_74#_M1011_s 0.00185913f $X=5.88 $Y=1.195 $X2=0
+ $Y2=0
cc_347 N_A_828_48#_M1001_g N_A_27_74#_c_758_n 0.011188f $X=4.215 $Y=0.74 $X2=0
+ $Y2=0
cc_348 N_A_828_48#_M1002_g N_A_27_74#_c_758_n 0.0112486f $X=4.645 $Y=0.74 $X2=0
+ $Y2=0
cc_349 N_A_828_48#_M1004_g N_A_27_74#_c_804_n 0.0065152f $X=5.145 $Y=0.74 $X2=0
+ $Y2=0
cc_350 N_A_828_48#_M1011_g N_A_27_74#_c_804_n 6.23275e-19 $X=5.645 $Y=0.74 $X2=0
+ $Y2=0
cc_351 N_A_828_48#_M1004_g N_A_27_74#_c_760_n 0.00831967f $X=5.145 $Y=0.74 $X2=0
+ $Y2=0
cc_352 N_A_828_48#_M1011_g N_A_27_74#_c_760_n 0.0149802f $X=5.645 $Y=0.74 $X2=0
+ $Y2=0
cc_353 N_A_828_48#_c_317_n N_A_27_74#_c_761_n 0.00108027f $X=5.795 $Y=1.515
+ $X2=0 $Y2=0
cc_354 N_A_828_48#_c_319_n N_A_27_74#_c_761_n 0.010707f $X=6.325 $Y=1.195 $X2=0
+ $Y2=0
cc_355 N_A_828_48#_c_320_n N_A_27_74#_c_761_n 0.0290538f $X=6.49 $Y=0.665 $X2=0
+ $Y2=0
cc_356 N_A_828_48#_c_321_n N_A_27_74#_c_761_n 0.0151554f $X=5.88 $Y=1.195 $X2=0
+ $Y2=0
cc_357 N_A_828_48#_M1004_g N_A_27_74#_c_764_n 0.00294698f $X=5.145 $Y=0.74 $X2=0
+ $Y2=0
cc_358 N_A_828_48#_c_319_n N_VGND_c_869_n 0.00695774f $X=6.325 $Y=1.195 $X2=0
+ $Y2=0
cc_359 N_A_828_48#_c_320_n N_VGND_c_869_n 0.0225912f $X=6.49 $Y=0.665 $X2=0
+ $Y2=0
cc_360 N_A_828_48#_M1001_g N_VGND_c_876_n 0.00278271f $X=4.215 $Y=0.74 $X2=0
+ $Y2=0
cc_361 N_A_828_48#_M1002_g N_VGND_c_876_n 0.00278271f $X=4.645 $Y=0.74 $X2=0
+ $Y2=0
cc_362 N_A_828_48#_M1004_g N_VGND_c_876_n 0.00278247f $X=5.145 $Y=0.74 $X2=0
+ $Y2=0
cc_363 N_A_828_48#_M1011_g N_VGND_c_876_n 0.00278271f $X=5.645 $Y=0.74 $X2=0
+ $Y2=0
cc_364 N_A_828_48#_c_320_n N_VGND_c_876_n 0.00685868f $X=6.49 $Y=0.665 $X2=0
+ $Y2=0
cc_365 N_A_828_48#_M1001_g N_VGND_c_879_n 0.0035414f $X=4.215 $Y=0.74 $X2=0
+ $Y2=0
cc_366 N_A_828_48#_M1002_g N_VGND_c_879_n 0.00354087f $X=4.645 $Y=0.74 $X2=0
+ $Y2=0
cc_367 N_A_828_48#_M1004_g N_VGND_c_879_n 0.00354743f $X=5.145 $Y=0.74 $X2=0
+ $Y2=0
cc_368 N_A_828_48#_M1011_g N_VGND_c_879_n 0.00359085f $X=5.645 $Y=0.74 $X2=0
+ $Y2=0
cc_369 N_A_828_48#_c_320_n N_VGND_c_879_n 0.00829701f $X=6.49 $Y=0.665 $X2=0
+ $Y2=0
cc_370 N_B1_N_c_433_n N_VPWR_c_555_n 0.0058365f $X=6.245 $Y=2.045 $X2=0 $Y2=0
cc_371 N_B1_N_c_433_n N_VPWR_c_557_n 6.93274e-19 $X=6.245 $Y=2.045 $X2=0 $Y2=0
cc_372 N_B1_N_c_436_n N_VPWR_c_557_n 0.0183312f $X=6.695 $Y=2.045 $X2=0 $Y2=0
cc_373 B1_N N_VPWR_c_557_n 0.0179834f $X=6.875 $Y=1.58 $X2=0 $Y2=0
cc_374 N_B1_N_c_433_n N_VPWR_c_563_n 0.00445602f $X=6.245 $Y=2.045 $X2=0 $Y2=0
cc_375 N_B1_N_c_436_n N_VPWR_c_563_n 0.00413917f $X=6.695 $Y=2.045 $X2=0 $Y2=0
cc_376 N_B1_N_c_433_n N_VPWR_c_551_n 0.00862391f $X=6.245 $Y=2.045 $X2=0 $Y2=0
cc_377 N_B1_N_c_436_n N_VPWR_c_551_n 0.00817726f $X=6.695 $Y=2.045 $X2=0 $Y2=0
cc_378 N_B1_N_c_430_n N_Y_c_647_n 4.3083e-19 $X=6.695 $Y=1.78 $X2=0 $Y2=0
cc_379 N_B1_N_c_433_n N_Y_c_648_n 0.00536313f $X=6.245 $Y=2.045 $X2=0 $Y2=0
cc_380 N_B1_N_M1007_g N_A_27_74#_c_760_n 5.88438e-19 $X=6.705 $Y=0.89 $X2=0
+ $Y2=0
cc_381 N_B1_N_M1007_g N_A_27_74#_c_761_n 0.00195452f $X=6.705 $Y=0.89 $X2=0
+ $Y2=0
cc_382 N_B1_N_M1007_g N_VGND_c_869_n 0.0160442f $X=6.705 $Y=0.89 $X2=0 $Y2=0
cc_383 B1_N N_VGND_c_869_n 0.0279913f $X=6.875 $Y=1.58 $X2=0 $Y2=0
cc_384 N_B1_N_M1007_g N_VGND_c_876_n 0.00394901f $X=6.705 $Y=0.89 $X2=0 $Y2=0
cc_385 N_B1_N_M1007_g N_VGND_c_879_n 0.00419525f $X=6.705 $Y=0.89 $X2=0 $Y2=0
cc_386 N_A_28_368#_c_481_n N_VPWR_M1008_s 0.00384138f $X=1.02 $Y=2.035 $X2=-0.19
+ $Y2=1.66
cc_387 N_A_28_368#_c_488_n N_VPWR_M1010_s 0.00383853f $X=2 $Y=2.035 $X2=0 $Y2=0
cc_388 N_A_28_368#_c_471_n N_VPWR_c_552_n 0.0453479f $X=0.285 $Y=2.44 $X2=0
+ $Y2=0
cc_389 N_A_28_368#_c_481_n N_VPWR_c_552_n 0.0154248f $X=1.02 $Y=2.035 $X2=0
+ $Y2=0
cc_390 N_A_28_368#_c_472_n N_VPWR_c_552_n 0.0453479f $X=1.185 $Y=2.44 $X2=0
+ $Y2=0
cc_391 N_A_28_368#_c_472_n N_VPWR_c_553_n 0.0462948f $X=1.185 $Y=2.44 $X2=0
+ $Y2=0
cc_392 N_A_28_368#_c_488_n N_VPWR_c_553_n 0.0171814f $X=2 $Y=2.035 $X2=0 $Y2=0
cc_393 N_A_28_368#_c_493_n N_VPWR_c_553_n 0.040027f $X=2.085 $Y=2.4 $X2=0 $Y2=0
cc_394 N_A_28_368#_c_475_n N_VPWR_c_553_n 0.0125885f $X=2.17 $Y=2.99 $X2=0 $Y2=0
cc_395 N_A_28_368#_c_474_n N_VPWR_c_558_n 0.0409869f $X=2.82 $Y=2.99 $X2=0 $Y2=0
cc_396 N_A_28_368#_c_475_n N_VPWR_c_558_n 0.0121867f $X=2.17 $Y=2.99 $X2=0 $Y2=0
cc_397 N_A_28_368#_c_476_n N_VPWR_c_558_n 0.0659319f $X=3.82 $Y=2.99 $X2=0 $Y2=0
cc_398 N_A_28_368#_c_478_n N_VPWR_c_558_n 0.0235512f $X=2.985 $Y=2.99 $X2=0
+ $Y2=0
cc_399 N_A_28_368#_c_471_n N_VPWR_c_560_n 0.011066f $X=0.285 $Y=2.44 $X2=0 $Y2=0
cc_400 N_A_28_368#_c_472_n N_VPWR_c_561_n 0.0110241f $X=1.185 $Y=2.44 $X2=0
+ $Y2=0
cc_401 N_A_28_368#_c_471_n N_VPWR_c_551_n 0.00915947f $X=0.285 $Y=2.44 $X2=0
+ $Y2=0
cc_402 N_A_28_368#_c_472_n N_VPWR_c_551_n 0.00909194f $X=1.185 $Y=2.44 $X2=0
+ $Y2=0
cc_403 N_A_28_368#_c_474_n N_VPWR_c_551_n 0.0231342f $X=2.82 $Y=2.99 $X2=0 $Y2=0
cc_404 N_A_28_368#_c_475_n N_VPWR_c_551_n 0.00660921f $X=2.17 $Y=2.99 $X2=0
+ $Y2=0
cc_405 N_A_28_368#_c_476_n N_VPWR_c_551_n 0.0367158f $X=3.82 $Y=2.99 $X2=0 $Y2=0
cc_406 N_A_28_368#_c_478_n N_VPWR_c_551_n 0.0126924f $X=2.985 $Y=2.99 $X2=0
+ $Y2=0
cc_407 N_A_28_368#_c_474_n N_Y_M1014_d 0.00222494f $X=2.82 $Y=2.99 $X2=0 $Y2=0
cc_408 N_A_28_368#_c_476_n N_Y_M1020_d 0.00250873f $X=3.82 $Y=2.99 $X2=0 $Y2=0
cc_409 N_A_28_368#_c_473_n N_Y_c_652_n 0.013092f $X=2.085 $Y=2.12 $X2=0 $Y2=0
cc_410 N_A_28_368#_c_493_n N_Y_c_655_n 0.0391515f $X=2.085 $Y=2.4 $X2=0 $Y2=0
cc_411 N_A_28_368#_c_474_n N_Y_c_655_n 0.0144323f $X=2.82 $Y=2.99 $X2=0 $Y2=0
cc_412 N_A_28_368#_c_502_n N_Y_c_655_n 0.0298377f $X=2.985 $Y=2.455 $X2=0 $Y2=0
cc_413 N_A_28_368#_M1017_s N_Y_c_657_n 0.00359365f $X=2.835 $Y=1.84 $X2=0 $Y2=0
cc_414 N_A_28_368#_c_502_n N_Y_c_657_n 0.0171813f $X=2.985 $Y=2.455 $X2=0 $Y2=0
cc_415 N_A_28_368#_c_476_n N_Y_c_661_n 0.018923f $X=3.82 $Y=2.99 $X2=0 $Y2=0
cc_416 N_A_28_368#_M1021_s N_Y_c_662_n 0.00595186f $X=3.785 $Y=1.84 $X2=0 $Y2=0
cc_417 N_A_28_368#_c_477_n N_Y_c_662_n 0.00997062f $X=3.985 $Y=2.375 $X2=0 $Y2=0
cc_418 N_A_28_368#_c_476_n N_Y_c_646_n 0.00536548f $X=3.82 $Y=2.99 $X2=0 $Y2=0
cc_419 N_A_28_368#_c_477_n N_Y_c_646_n 0.041429f $X=3.985 $Y=2.375 $X2=0 $Y2=0
cc_420 N_A_28_368#_M1021_s N_Y_c_649_n 0.00336744f $X=3.785 $Y=1.84 $X2=0 $Y2=0
cc_421 N_A_28_368#_c_477_n N_Y_c_649_n 0.0166119f $X=3.985 $Y=2.375 $X2=0 $Y2=0
cc_422 N_A_28_368#_M1021_s Y 0.0021281f $X=3.785 $Y=1.84 $X2=0 $Y2=0
cc_423 N_A_28_368#_c_473_n N_A_27_74#_c_756_n 0.00115483f $X=2.085 $Y=2.12 $X2=0
+ $Y2=0
cc_424 N_A_28_368#_c_473_n N_A_27_74#_c_763_n 0.00499031f $X=2.085 $Y=2.12 $X2=0
+ $Y2=0
cc_425 N_VPWR_c_554_n N_Y_c_646_n 0.0514855f $X=4.995 $Y=2.355 $X2=0 $Y2=0
cc_426 N_VPWR_c_558_n N_Y_c_646_n 0.0145938f $X=4.91 $Y=3.33 $X2=0 $Y2=0
cc_427 N_VPWR_c_551_n N_Y_c_646_n 0.0120466f $X=6.96 $Y=3.33 $X2=0 $Y2=0
cc_428 N_VPWR_M1000_d N_Y_c_691_n 0.0047272f $X=4.845 $Y=1.84 $X2=0 $Y2=0
cc_429 N_VPWR_c_554_n N_Y_c_691_n 0.0136682f $X=4.995 $Y=2.355 $X2=0 $Y2=0
cc_430 N_VPWR_c_554_n N_Y_c_648_n 0.0487067f $X=4.995 $Y=2.355 $X2=0 $Y2=0
cc_431 N_VPWR_c_555_n N_Y_c_648_n 0.0455614f $X=6.02 $Y=2.455 $X2=0 $Y2=0
cc_432 N_VPWR_c_562_n N_Y_c_648_n 0.0145938f $X=5.855 $Y=3.33 $X2=0 $Y2=0
cc_433 N_VPWR_c_551_n N_Y_c_648_n 0.0120466f $X=6.96 $Y=3.33 $X2=0 $Y2=0
cc_434 N_Y_c_643_n N_A_27_74#_M1023_d 0.00261553f $X=4.595 $Y=1.095 $X2=0 $Y2=0
cc_435 N_Y_c_642_n N_A_27_74#_M1002_s 0.00250873f $X=5.265 $Y=1.095 $X2=0 $Y2=0
cc_436 N_Y_c_643_n N_A_27_74#_c_793_n 0.00948342f $X=4.595 $Y=1.095 $X2=0 $Y2=0
cc_437 N_Y_M1001_d N_A_27_74#_c_758_n 0.00176461f $X=4.29 $Y=0.37 $X2=0 $Y2=0
cc_438 N_Y_c_664_n N_A_27_74#_c_758_n 0.0154609f $X=4.43 $Y=0.82 $X2=0 $Y2=0
cc_439 N_Y_c_643_n N_A_27_74#_c_758_n 0.00614817f $X=4.595 $Y=1.095 $X2=0 $Y2=0
cc_440 N_Y_c_642_n N_A_27_74#_c_804_n 0.0207721f $X=5.265 $Y=1.095 $X2=0 $Y2=0
cc_441 N_Y_M1004_d N_A_27_74#_c_760_n 0.00250873f $X=5.22 $Y=0.37 $X2=0 $Y2=0
cc_442 N_Y_c_642_n N_A_27_74#_c_760_n 0.00304353f $X=5.265 $Y=1.095 $X2=0 $Y2=0
cc_443 N_Y_c_695_n N_A_27_74#_c_760_n 0.019446f $X=5.43 $Y=0.86 $X2=0 $Y2=0
cc_444 N_A_27_74#_c_751_n N_VGND_M1006_d 0.00229612f $X=1.105 $Y=1.095 $X2=-0.19
+ $Y2=-0.245
cc_445 N_A_27_74#_c_754_n N_VGND_M1019_d 0.00176461f $X=1.965 $Y=1.095 $X2=0
+ $Y2=0
cc_446 N_A_27_74#_c_756_n N_VGND_M1003_s 0.00176461f $X=2.825 $Y=1.095 $X2=0
+ $Y2=0
cc_447 N_A_27_74#_c_793_n N_VGND_M1013_s 0.00931318f $X=3.765 $Y=0.755 $X2=0
+ $Y2=0
cc_448 N_A_27_74#_c_750_n N_VGND_c_864_n 0.0182902f $X=0.28 $Y=0.515 $X2=0 $Y2=0
cc_449 N_A_27_74#_c_751_n N_VGND_c_864_n 0.0193595f $X=1.105 $Y=1.095 $X2=0
+ $Y2=0
cc_450 N_A_27_74#_c_753_n N_VGND_c_864_n 0.00121793f $X=1.19 $Y=0.515 $X2=0
+ $Y2=0
cc_451 N_A_27_74#_c_753_n N_VGND_c_865_n 0.0182488f $X=1.19 $Y=0.515 $X2=0 $Y2=0
cc_452 N_A_27_74#_c_754_n N_VGND_c_865_n 0.0170777f $X=1.965 $Y=1.095 $X2=0
+ $Y2=0
cc_453 N_A_27_74#_c_755_n N_VGND_c_865_n 0.0182488f $X=2.05 $Y=0.515 $X2=0 $Y2=0
cc_454 N_A_27_74#_c_755_n N_VGND_c_866_n 0.0182488f $X=2.05 $Y=0.515 $X2=0 $Y2=0
cc_455 N_A_27_74#_c_756_n N_VGND_c_866_n 0.0170777f $X=2.825 $Y=1.095 $X2=0
+ $Y2=0
cc_456 N_A_27_74#_c_757_n N_VGND_c_866_n 0.0121972f $X=2.91 $Y=0.515 $X2=0 $Y2=0
cc_457 N_A_27_74#_c_757_n N_VGND_c_867_n 0.00591149f $X=2.91 $Y=0.515 $X2=0
+ $Y2=0
cc_458 N_A_27_74#_c_793_n N_VGND_c_867_n 0.0251188f $X=3.765 $Y=0.755 $X2=0
+ $Y2=0
cc_459 N_A_27_74#_c_759_n N_VGND_c_867_n 0.0114117f $X=4.095 $Y=0.34 $X2=0 $Y2=0
cc_460 N_A_27_74#_c_760_n N_VGND_c_869_n 0.00567334f $X=5.765 $Y=0.34 $X2=0
+ $Y2=0
cc_461 N_A_27_74#_c_761_n N_VGND_c_869_n 0.0020999f $X=5.93 $Y=0.515 $X2=0 $Y2=0
cc_462 N_A_27_74#_c_755_n N_VGND_c_870_n 0.00749631f $X=2.05 $Y=0.515 $X2=0
+ $Y2=0
cc_463 N_A_27_74#_c_757_n N_VGND_c_872_n 0.0109942f $X=2.91 $Y=0.515 $X2=0 $Y2=0
cc_464 N_A_27_74#_c_793_n N_VGND_c_872_n 0.00236055f $X=3.765 $Y=0.755 $X2=0
+ $Y2=0
cc_465 N_A_27_74#_c_750_n N_VGND_c_874_n 0.011066f $X=0.28 $Y=0.515 $X2=0 $Y2=0
cc_466 N_A_27_74#_c_753_n N_VGND_c_875_n 0.00749631f $X=1.19 $Y=0.515 $X2=0
+ $Y2=0
cc_467 N_A_27_74#_c_793_n N_VGND_c_876_n 0.00236055f $X=3.765 $Y=0.755 $X2=0
+ $Y2=0
cc_468 N_A_27_74#_c_758_n N_VGND_c_876_n 0.0422287f $X=4.765 $Y=0.34 $X2=0 $Y2=0
cc_469 N_A_27_74#_c_759_n N_VGND_c_876_n 0.0233032f $X=4.095 $Y=0.34 $X2=0 $Y2=0
cc_470 N_A_27_74#_c_760_n N_VGND_c_876_n 0.0659741f $X=5.765 $Y=0.34 $X2=0 $Y2=0
cc_471 N_A_27_74#_c_764_n N_VGND_c_876_n 0.0233048f $X=4.93 $Y=0.34 $X2=0 $Y2=0
cc_472 N_A_27_74#_c_750_n N_VGND_c_879_n 0.00915947f $X=0.28 $Y=0.515 $X2=0
+ $Y2=0
cc_473 N_A_27_74#_c_753_n N_VGND_c_879_n 0.0062048f $X=1.19 $Y=0.515 $X2=0 $Y2=0
cc_474 N_A_27_74#_c_755_n N_VGND_c_879_n 0.0062048f $X=2.05 $Y=0.515 $X2=0 $Y2=0
cc_475 N_A_27_74#_c_757_n N_VGND_c_879_n 0.00904371f $X=2.91 $Y=0.515 $X2=0
+ $Y2=0
cc_476 N_A_27_74#_c_793_n N_VGND_c_879_n 0.0102106f $X=3.765 $Y=0.755 $X2=0
+ $Y2=0
cc_477 N_A_27_74#_c_758_n N_VGND_c_879_n 0.0238173f $X=4.765 $Y=0.34 $X2=0 $Y2=0
cc_478 N_A_27_74#_c_759_n N_VGND_c_879_n 0.012665f $X=4.095 $Y=0.34 $X2=0 $Y2=0
cc_479 N_A_27_74#_c_760_n N_VGND_c_879_n 0.0367637f $X=5.765 $Y=0.34 $X2=0 $Y2=0
cc_480 N_A_27_74#_c_764_n N_VGND_c_879_n 0.0126653f $X=4.93 $Y=0.34 $X2=0 $Y2=0
