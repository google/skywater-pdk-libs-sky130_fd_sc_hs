* File: sky130_fd_sc_hs__o22ai_2.spice
* Created: Tue Sep  1 20:16:28 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hs__o22ai_2.pex.spice"
.subckt sky130_fd_sc_hs__o22ai_2  VNB VPB B1 B2 A2 A1 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A1	A1
* A2	A2
* B2	B2
* B1	B1
* VPB	VPB
* VNB	VNB
MM1009 N_A_27_74#_M1009_d N_B1_M1009_g N_Y_M1009_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.1406 PD=2.05 PS=1.12 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75000.2
+ SB=75004 A=0.111 P=1.78 MULT=1
MM1012 N_A_27_74#_M1012_d N_B1_M1012_g N_Y_M1009_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1184 AS=0.1406 PD=1.06 PS=1.12 NRD=6.48 NRS=4.86 M=1 R=4.93333 SA=75000.7
+ SB=75003.5 A=0.111 P=1.78 MULT=1
MM1003 N_A_27_74#_M1012_d N_B2_M1003_g N_Y_M1003_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1184 AS=0.1295 PD=1.06 PS=1.09 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75001.2
+ SB=75003 A=0.111 P=1.78 MULT=1
MM1007 N_A_27_74#_M1007_d N_B2_M1007_g N_Y_M1003_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.2812 AS=0.1295 PD=1.5 PS=1.09 NRD=77.832 NRS=0 M=1 R=4.93333 SA=75001.7
+ SB=75002.5 A=0.111 P=1.78 MULT=1
MM1010 N_A_27_74#_M1007_d N_A2_M1010_g N_VGND_M1010_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.2812 AS=0.1184 PD=1.5 PS=1.06 NRD=0 NRS=0 M=1 R=4.93333 SA=75002.6
+ SB=75001.6 A=0.111 P=1.78 MULT=1
MM1014 N_A_27_74#_M1014_d N_A2_M1014_g N_VGND_M1010_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1184 PD=1.02 PS=1.06 NRD=0 NRS=6.48 M=1 R=4.93333 SA=75003.1
+ SB=75001.1 A=0.111 P=1.78 MULT=1
MM1001 N_A_27_74#_M1014_d N_A1_M1001_g N_VGND_M1001_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1295 PD=1.02 PS=1.09 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75003.5
+ SB=75000.7 A=0.111 P=1.78 MULT=1
MM1004 N_A_27_74#_M1004_d N_A1_M1004_g N_VGND_M1001_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.1295 PD=2.05 PS=1.09 NRD=0 NRS=0 M=1 R=4.93333 SA=75004
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1002 N_A_28_368#_M1002_d N_B1_M1002_g N_VPWR_M1002_s VPB PSHORT L=0.15 W=1.12
+ AD=0.3304 AS=0.196 PD=2.83 PS=1.47 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75001.6 A=0.168 P=2.54 MULT=1
MM1006 N_A_28_368#_M1006_d N_B1_M1006_g N_VPWR_M1002_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.196 PD=1.42 PS=1.47 NRD=1.7533 NRS=10.5395 M=1 R=7.46667
+ SA=75000.7 SB=75001.1 A=0.168 P=2.54 MULT=1
MM1005 N_Y_M1005_d N_B2_M1005_g N_A_28_368#_M1006_d VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.2 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1008 N_Y_M1005_d N_B2_M1008_g N_A_28_368#_M1008_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.3304 PD=1.42 PS=2.83 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.6 SB=75000.2 A=0.168 P=2.54 MULT=1
MM1011 N_Y_M1011_d N_A2_M1011_g N_A_510_368#_M1011_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.3304 PD=1.42 PS=2.83 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75001.6 A=0.168 P=2.54 MULT=1
MM1013 N_Y_M1011_d N_A2_M1013_g N_A_510_368#_M1013_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.7 SB=75001.1 A=0.168 P=2.54 MULT=1
MM1000 N_A_510_368#_M1013_s N_A1_M1000_g N_VPWR_M1000_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.1 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1015 N_A_510_368#_M1015_d N_A1_M1015_g N_VPWR_M1000_s VPB PSHORT L=0.15 W=1.12
+ AD=0.3304 AS=0.168 PD=2.83 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.6 SB=75000.2 A=0.168 P=2.54 MULT=1
DX16_noxref VNB VPB NWDIODE A=9.6348 P=14.08
*
.include "sky130_fd_sc_hs__o22ai_2.pxi.spice"
*
.ends
*
*
