* File: sky130_fd_sc_hs__xnor3_1.pex.spice
* Created: Tue Sep  1 20:25:29 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HS__XNOR3_1%A_81_268# 1 2 7 9 10 12 16 17 18 19 20 22 23
+ 24 26 27 28 31 34 36 39
r100 39 41 6.80989 $w=3.28e-07 $l=1.95e-07 $layer=LI1_cond $X=2.49 $Y=2.795
+ $X2=2.49 $Y2=2.99
r101 34 37 8.51103 $w=3.58e-07 $l=1.65e-07 $layer=LI1_cond $X=0.605 $Y=1.505
+ $X2=0.605 $Y2=1.67
r102 34 36 8.51103 $w=3.58e-07 $l=1.65e-07 $layer=LI1_cond $X=0.605 $Y=1.505
+ $X2=0.605 $Y2=1.34
r103 34 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.59
+ $Y=1.505 $X2=0.59 $Y2=1.505
r104 29 31 4.1907 $w=3.28e-07 $l=1.2e-07 $layer=LI1_cond $X=2.5 $Y=0.425 $X2=2.5
+ $Y2=0.545
r105 27 29 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.335 $Y=0.34
+ $X2=2.5 $Y2=0.425
r106 27 28 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.335 $Y=0.34
+ $X2=1.665 $Y2=0.34
r107 25 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.58 $Y=0.425
+ $X2=1.665 $Y2=0.34
r108 25 26 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=1.58 $Y=0.425
+ $X2=1.58 $Y2=0.66
r109 23 41 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.325 $Y=2.99
+ $X2=2.49 $Y2=2.99
r110 23 24 76.984 $w=1.68e-07 $l=1.18e-06 $layer=LI1_cond $X=2.325 $Y=2.99
+ $X2=1.145 $Y2=2.99
r111 22 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.06 $Y=2.905
+ $X2=1.145 $Y2=2.99
r112 21 22 51.2139 $w=1.68e-07 $l=7.85e-07 $layer=LI1_cond $X=1.06 $Y=2.12
+ $X2=1.06 $Y2=2.905
r113 19 21 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.975 $Y=2.035
+ $X2=1.06 $Y2=2.12
r114 19 20 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=0.975 $Y=2.035
+ $X2=0.785 $Y2=2.035
r115 17 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.495 $Y=0.745
+ $X2=1.58 $Y2=0.66
r116 17 18 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=1.495 $Y=0.745
+ $X2=0.785 $Y2=0.745
r117 16 20 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.7 $Y=1.95
+ $X2=0.785 $Y2=2.035
r118 16 37 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=0.7 $Y=1.95 $X2=0.7
+ $Y2=1.67
r119 13 18 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.7 $Y=0.83
+ $X2=0.785 $Y2=0.745
r120 13 36 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=0.7 $Y=0.83 $X2=0.7
+ $Y2=1.34
r121 10 35 53.2088 $w=3.12e-07 $l=2.995e-07 $layer=POLY_cond $X=0.495 $Y=1.765
+ $X2=0.58 $Y2=1.505
r122 10 12 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.495 $Y=1.765
+ $X2=0.495 $Y2=2.4
r123 7 35 38.5325 $w=3.12e-07 $l=2.03101e-07 $layer=POLY_cond $X=0.495 $Y=1.34
+ $X2=0.58 $Y2=1.505
r124 7 9 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=0.495 $Y=1.34
+ $X2=0.495 $Y2=0.86
r125 2 39 600 $w=1.7e-07 $l=9.32939e-07 $layer=licon1_PDIFF $count=1 $X=2.26
+ $Y=1.97 $X2=2.49 $Y2=2.795
r126 1 31 91 $w=1.7e-07 $l=2.84341e-07 $layer=licon1_NDIFF $count=2 $X=2.29
+ $Y=0.37 $X2=2.5 $Y2=0.545
.ends

.subckt PM_SKY130_FD_SC_HS__XNOR3_1%C 1 3 4 6 7 9 10 11 13 14 16 18 23
c77 4 0 1.73622e-19 $X=1.175 $Y=1.765
c78 1 0 1.63453e-19 $X=1.085 $Y=1.35
r79 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.16
+ $Y=1.515 $X2=1.16 $Y2=1.515
r80 20 22 14.5084 $w=2.99e-07 $l=9e-08 $layer=POLY_cond $X=1.16 $Y=1.425
+ $X2=1.16 $Y2=1.515
r81 18 23 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=1.16 $Y=1.665
+ $X2=1.16 $Y2=1.515
r82 14 17 98.2126 $w=1.68e-07 $l=3.51312e-07 $layer=POLY_cond $X=2.215 $Y=1.085
+ $X2=2.192 $Y2=1.425
r83 14 16 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=2.215 $Y=1.085
+ $X2=2.215 $Y2=0.69
r84 11 13 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=2.185 $Y=1.895
+ $X2=2.185 $Y2=2.39
r85 10 11 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=2.185 $Y=1.805
+ $X2=2.185 $Y2=1.895
r86 9 17 44.4659 $w=1.8e-07 $l=1.68464e-07 $layer=POLY_cond $X=2.185 $Y=1.59
+ $X2=2.192 $Y2=1.425
r87 9 10 83.5726 $w=1.8e-07 $l=2.15e-07 $layer=POLY_cond $X=2.185 $Y=1.59
+ $X2=2.185 $Y2=1.805
r88 8 20 18.89 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.325 $Y=1.425
+ $X2=1.16 $Y2=1.425
r89 7 17 5.52526 $w=1.5e-07 $l=9.7e-08 $layer=POLY_cond $X=2.095 $Y=1.425
+ $X2=2.192 $Y2=1.425
r90 7 8 394.83 $w=1.5e-07 $l=7.7e-07 $layer=POLY_cond $X=2.095 $Y=1.425
+ $X2=1.325 $Y2=1.425
r91 4 22 52.2586 $w=2.99e-07 $l=2.57391e-07 $layer=POLY_cond $X=1.175 $Y=1.765
+ $X2=1.16 $Y2=1.515
r92 4 6 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=1.175 $Y=1.765
+ $X2=1.175 $Y2=2.16
r93 1 20 24.0479 $w=2.99e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.085 $Y=1.35
+ $X2=1.16 $Y2=1.425
r94 1 3 106.04 $w=1.5e-07 $l=3.3e-07 $layer=POLY_cond $X=1.085 $Y=1.35 $X2=1.085
+ $Y2=1.02
.ends

.subckt PM_SKY130_FD_SC_HS__XNOR3_1%A_232_162# 1 2 9 11 13 14 18 22 27 28 30 32
r88 30 32 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=2.68 $Y=1.645
+ $X2=2.515 $Y2=1.645
r89 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.68
+ $Y=1.645 $X2=2.68 $Y2=1.645
r90 26 28 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.665 $Y=1.665
+ $X2=1.58 $Y2=1.665
r91 26 32 55.4545 $w=1.68e-07 $l=8.5e-07 $layer=LI1_cond $X=1.665 $Y=1.665
+ $X2=2.515 $Y2=1.665
r92 23 28 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.58 $Y=1.75 $X2=1.58
+ $Y2=1.665
r93 23 27 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=1.58 $Y=1.75 $X2=1.58
+ $Y2=1.95
r94 22 28 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.58 $Y=1.58 $X2=1.58
+ $Y2=1.665
r95 21 22 26.7487 $w=1.68e-07 $l=4.1e-07 $layer=LI1_cond $X=1.58 $Y=1.17
+ $X2=1.58 $Y2=1.58
r96 18 27 8.81775 $w=3.48e-07 $l=1.75e-07 $layer=LI1_cond $X=1.49 $Y=2.125
+ $X2=1.49 $Y2=1.95
r97 18 20 3.48571 $w=3.5e-07 $l=1e-07 $layer=LI1_cond $X=1.49 $Y=2.125 $X2=1.49
+ $Y2=2.225
r98 14 21 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.495 $Y=1.085
+ $X2=1.58 $Y2=1.17
r99 14 16 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=1.495 $Y=1.085
+ $X2=1.3 $Y2=1.085
r100 11 31 51.1109 $w=3.27e-07 $l=2.92831e-07 $layer=POLY_cond $X=2.79 $Y=1.895
+ $X2=2.697 $Y2=1.645
r101 11 13 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=2.79 $Y=1.895
+ $X2=2.79 $Y2=2.39
r102 7 31 38.5818 $w=3.27e-07 $l=1.73767e-07 $layer=POLY_cond $X=2.715 $Y=1.48
+ $X2=2.697 $Y2=1.645
r103 7 9 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.715 $Y=1.48
+ $X2=2.715 $Y2=0.69
r104 2 20 600 $w=1.7e-07 $l=4.53845e-07 $layer=licon1_PDIFF $count=1 $X=1.25
+ $Y=1.84 $X2=1.4 $Y2=2.225
r105 1 16 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=1.16
+ $Y=0.81 $X2=1.3 $Y2=1.085
.ends

.subckt PM_SKY130_FD_SC_HS__XNOR3_1%A_786_100# 1 2 7 9 13 14 15 17 18 20 24 27
+ 29 33 38 40 44
c125 38 0 3.96032e-20 $X=4.63 $Y=1.355
c126 27 0 1.45365e-19 $X=6.095 $Y=1.395
c127 24 0 1.34101e-19 $X=6.095 $Y=1.035
c128 13 0 1.3366e-19 $X=4.97 $Y=0.925
r129 44 45 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.88
+ $Y=1.52 $X2=4.88 $Y2=1.52
r130 41 44 8.73063 $w=3.28e-07 $l=2.5e-07 $layer=LI1_cond $X=4.63 $Y=1.52
+ $X2=4.88 $Y2=1.52
r131 39 41 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.63 $Y=1.685
+ $X2=4.63 $Y2=1.52
r132 39 40 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=4.63 $Y=1.685
+ $X2=4.63 $Y2=1.95
r133 38 41 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.63 $Y=1.355
+ $X2=4.63 $Y2=1.52
r134 37 38 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=4.63 $Y=1.18
+ $X2=4.63 $Y2=1.355
r135 33 40 7.14316 $w=2.5e-07 $l=1.62019e-07 $layer=LI1_cond $X=4.545 $Y=2.075
+ $X2=4.63 $Y2=1.95
r136 33 35 21.205 $w=2.48e-07 $l=4.6e-07 $layer=LI1_cond $X=4.545 $Y=2.075
+ $X2=4.085 $Y2=2.075
r137 29 37 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.545 $Y=1.095
+ $X2=4.63 $Y2=1.18
r138 29 31 30.9893 $w=1.68e-07 $l=4.75e-07 $layer=LI1_cond $X=4.545 $Y=1.095
+ $X2=4.07 $Y2=1.095
r139 22 27 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.095 $Y=1.32
+ $X2=6.095 $Y2=1.395
r140 22 24 146.138 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=6.095 $Y=1.32
+ $X2=6.095 $Y2=1.035
r141 21 24 394.83 $w=1.5e-07 $l=7.7e-07 $layer=POLY_cond $X=6.095 $Y=0.265
+ $X2=6.095 $Y2=1.035
r142 18 20 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=5.94 $Y=1.84
+ $X2=5.94 $Y2=2.235
r143 17 18 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=5.94 $Y=1.75 $X2=5.94
+ $Y2=1.84
r144 16 27 79.4787 $w=1.5e-07 $l=1.55e-07 $layer=POLY_cond $X=5.94 $Y=1.395
+ $X2=6.095 $Y2=1.395
r145 16 17 108.839 $w=1.8e-07 $l=2.8e-07 $layer=POLY_cond $X=5.94 $Y=1.47
+ $X2=5.94 $Y2=1.75
r146 14 21 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=6.02 $Y=0.19
+ $X2=6.095 $Y2=0.265
r147 14 15 499.947 $w=1.5e-07 $l=9.75e-07 $layer=POLY_cond $X=6.02 $Y=0.19
+ $X2=5.045 $Y2=0.19
r148 11 45 38.5916 $w=2.93e-07 $l=2.05122e-07 $layer=POLY_cond $X=4.97 $Y=1.355
+ $X2=4.88 $Y2=1.52
r149 11 13 220.489 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=4.97 $Y=1.355
+ $X2=4.97 $Y2=0.925
r150 10 15 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.97 $Y=0.265
+ $X2=5.045 $Y2=0.19
r151 10 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.97 $Y=0.265
+ $X2=4.97 $Y2=0.925
r152 7 45 55.8646 $w=2.93e-07 $l=3.05205e-07 $layer=POLY_cond $X=4.955 $Y=1.79
+ $X2=4.88 $Y2=1.52
r153 7 9 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=4.955 $Y=1.79
+ $X2=4.955 $Y2=2.285
r154 2 35 600 $w=1.7e-07 $l=3.4187e-07 $layer=licon1_PDIFF $count=1 $X=3.935
+ $Y=1.84 $X2=4.085 $Y2=2.115
r155 1 31 182 $w=1.7e-07 $l=6.61306e-07 $layer=licon1_NDIFF $count=1 $X=3.93
+ $Y=0.5 $X2=4.07 $Y2=1.095
.ends

.subckt PM_SKY130_FD_SC_HS__XNOR3_1%B 1 3 4 6 8 9 10 11 12 16 19 21 23 24 25 28
+ 31 34 35 37 38 40 44
c144 35 0 1.73263e-19 $X=4.295 $Y=1.515
c145 34 0 1.66544e-19 $X=3.705 $Y=1.35
c146 23 0 1.42592e-19 $X=6.575 $Y=2.92
r147 43 44 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.21
+ $Y=1.515 $X2=4.21 $Y2=1.515
r148 40 44 2.67779 $w=6.68e-07 $l=1.5e-07 $layer=LI1_cond $X=4.04 $Y=1.665
+ $X2=4.04 $Y2=1.515
r149 36 37 47.3682 $w=2.1e-07 $l=1.5e-07 $layer=POLY_cond $X=5.505 $Y=1.69
+ $X2=5.505 $Y2=1.84
r150 35 43 14.8632 $w=3.3e-07 $l=8.5e-08 $layer=POLY_cond $X=4.295 $Y=1.515
+ $X2=4.21 $Y2=1.515
r151 33 43 45.4639 $w=3.3e-07 $l=2.6e-07 $layer=POLY_cond $X=3.95 $Y=1.515
+ $X2=4.21 $Y2=1.515
r152 33 34 5.03009 $w=3.3e-07 $l=3.16938e-07 $layer=POLY_cond $X=3.95 $Y=1.515
+ $X2=3.705 $Y2=1.35
r153 31 39 392.266 $w=1.5e-07 $l=7.65e-07 $layer=POLY_cond $X=6.59 $Y=0.925
+ $X2=6.59 $Y2=1.69
r154 26 28 253.819 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=6.575 $Y=2.83
+ $X2=6.575 $Y2=2.335
r155 25 39 58.3064 $w=1.8e-07 $l=1.5e-07 $layer=POLY_cond $X=6.575 $Y=1.84
+ $X2=6.575 $Y2=1.69
r156 25 28 253.819 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=6.575 $Y=1.84
+ $X2=6.575 $Y2=2.335
r157 23 26 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=6.575 $Y=2.92
+ $X2=6.575 $Y2=2.83
r158 23 24 60.25 $w=1.8e-07 $l=1.55e-07 $layer=POLY_cond $X=6.575 $Y=2.92
+ $X2=6.575 $Y2=3.075
r159 22 38 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=5.58 $Y=3.15 $X2=5.49
+ $Y2=3.15
r160 21 24 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=6.485 $Y=3.15
+ $X2=6.575 $Y2=3.075
r161 21 22 464.053 $w=1.5e-07 $l=9.05e-07 $layer=POLY_cond $X=6.485 $Y=3.15
+ $X2=5.58 $Y2=3.15
r162 19 36 392.266 $w=1.5e-07 $l=7.65e-07 $layer=POLY_cond $X=5.535 $Y=0.925
+ $X2=5.535 $Y2=1.69
r163 16 37 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=5.49 $Y=2.235
+ $X2=5.49 $Y2=1.84
r164 14 16 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=5.49 $Y=2.63
+ $X2=5.49 $Y2=2.235
r165 12 38 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=5.49 $Y=3.075
+ $X2=5.49 $Y2=3.15
r166 11 14 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=5.49 $Y=2.72 $X2=5.49
+ $Y2=2.63
r167 11 12 137.992 $w=1.8e-07 $l=3.55e-07 $layer=POLY_cond $X=5.49 $Y=2.72
+ $X2=5.49 $Y2=3.075
r168 9 38 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=5.4 $Y=3.15 $X2=5.49
+ $Y2=3.15
r169 9 10 489.691 $w=1.5e-07 $l=9.55e-07 $layer=POLY_cond $X=5.4 $Y=3.15
+ $X2=4.445 $Y2=3.15
r170 8 10 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.37 $Y=3.075
+ $X2=4.445 $Y2=3.15
r171 7 35 32.1775 $w=3.3e-07 $l=1.98997e-07 $layer=POLY_cond $X=4.37 $Y=1.68
+ $X2=4.295 $Y2=1.515
r172 7 8 715.309 $w=1.5e-07 $l=1.395e-06 $layer=POLY_cond $X=4.37 $Y=1.68
+ $X2=4.37 $Y2=3.075
r173 4 34 37.0704 $w=1.5e-07 $l=4.86364e-07 $layer=POLY_cond $X=3.86 $Y=1.765
+ $X2=3.705 $Y2=1.35
r174 4 6 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.86 $Y=1.765
+ $X2=3.86 $Y2=2.4
r175 1 34 37.0704 $w=1.5e-07 $l=1.5e-07 $layer=POLY_cond $X=3.855 $Y=1.35
+ $X2=3.705 $Y2=1.35
r176 1 3 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=3.855 $Y=1.35
+ $X2=3.855 $Y2=0.87
.ends

.subckt PM_SKY130_FD_SC_HS__XNOR3_1%A 3 5 7 8
c43 5 0 1.78665e-19 $X=7.115 $Y=1.84
c44 3 0 4.37781e-20 $X=7.085 $Y=0.925
r45 8 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.04
+ $Y=1.59 $X2=7.04 $Y2=1.59
r46 5 11 52.2586 $w=2.99e-07 $l=2.85044e-07 $layer=POLY_cond $X=7.115 $Y=1.84
+ $X2=7.04 $Y2=1.59
r47 5 7 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=7.115 $Y=1.84
+ $X2=7.115 $Y2=2.415
r48 1 11 38.5562 $w=2.99e-07 $l=1.86145e-07 $layer=POLY_cond $X=7.085 $Y=1.425
+ $X2=7.04 $Y2=1.59
r49 1 3 256.383 $w=1.5e-07 $l=5e-07 $layer=POLY_cond $X=7.085 $Y=1.425 $X2=7.085
+ $Y2=0.925
.ends

.subckt PM_SKY130_FD_SC_HS__XNOR3_1%A_897_54# 1 2 3 4 13 15 18 20 22 27 28 29 30
+ 31 32 37 41 43 50 52
c124 13 0 1.54564e-19 $X=7.65 $Y=1.84
r125 50 53 8.01359 $w=2.48e-07 $l=1.65e-07 $layer=LI1_cond $X=7.54 $Y=1.59
+ $X2=7.54 $Y2=1.755
r126 50 52 8.01359 $w=2.48e-07 $l=1.65e-07 $layer=LI1_cond $X=7.54 $Y=1.59
+ $X2=7.54 $Y2=1.425
r127 50 51 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.58
+ $Y=1.59 $X2=7.58 $Y2=1.59
r128 43 45 6.80989 $w=3.28e-07 $l=1.95e-07 $layer=LI1_cond $X=4.655 $Y=2.795
+ $X2=4.655 $Y2=2.99
r129 39 41 10.0285 $w=2.43e-07 $l=1.9e-07 $layer=LI1_cond $X=4.65 $Y=0.377
+ $X2=4.84 $Y2=0.377
r130 37 53 10.5499 $w=2.03e-07 $l=1.95e-07 $layer=LI1_cond $X=7.517 $Y=1.95
+ $X2=7.517 $Y2=1.755
r131 34 52 9.19734 $w=2.03e-07 $l=1.7e-07 $layer=LI1_cond $X=7.517 $Y=1.255
+ $X2=7.517 $Y2=1.425
r132 33 48 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.09 $Y=2.035
+ $X2=6.925 $Y2=2.035
r133 32 37 6.89401 $w=1.7e-07 $l=1.38109e-07 $layer=LI1_cond $X=7.415 $Y=2.035
+ $X2=7.517 $Y2=1.95
r134 32 33 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=7.415 $Y=2.035
+ $X2=7.09 $Y2=2.035
r135 30 34 6.89401 $w=1.7e-07 $l=1.38109e-07 $layer=LI1_cond $X=7.415 $Y=1.17
+ $X2=7.517 $Y2=1.255
r136 30 31 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=7.415 $Y=1.17
+ $X2=7.035 $Y2=1.17
r137 28 48 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.925 $Y=2.12
+ $X2=6.925 $Y2=2.035
r138 28 29 27.4142 $w=3.28e-07 $l=7.85e-07 $layer=LI1_cond $X=6.925 $Y=2.12
+ $X2=6.925 $Y2=2.905
r139 25 31 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=6.87 $Y=1.085
+ $X2=7.035 $Y2=1.17
r140 25 27 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=6.87 $Y=1.085
+ $X2=6.87 $Y2=0.75
r141 24 27 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=6.87 $Y=0.425
+ $X2=6.87 $Y2=0.75
r142 22 24 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=6.705 $Y=0.34
+ $X2=6.87 $Y2=0.425
r143 22 41 121.674 $w=1.68e-07 $l=1.865e-06 $layer=LI1_cond $X=6.705 $Y=0.34
+ $X2=4.84 $Y2=0.34
r144 21 45 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.82 $Y=2.99
+ $X2=4.655 $Y2=2.99
r145 20 29 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=6.76 $Y=2.99
+ $X2=6.925 $Y2=2.905
r146 20 21 126.567 $w=1.68e-07 $l=1.94e-06 $layer=LI1_cond $X=6.76 $Y=2.99
+ $X2=4.82 $Y2=2.99
r147 16 51 38.5562 $w=2.99e-07 $l=2.03101e-07 $layer=POLY_cond $X=7.665 $Y=1.425
+ $X2=7.58 $Y2=1.59
r148 16 18 256.383 $w=1.5e-07 $l=5e-07 $layer=POLY_cond $X=7.665 $Y=1.425
+ $X2=7.665 $Y2=0.925
r149 13 51 52.2586 $w=2.99e-07 $l=2.82843e-07 $layer=POLY_cond $X=7.65 $Y=1.84
+ $X2=7.58 $Y2=1.59
r150 13 15 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=7.65 $Y=1.84
+ $X2=7.65 $Y2=2.415
r151 4 48 300 $w=1.7e-07 $l=3.19726e-07 $layer=licon1_PDIFF $count=2 $X=6.65
+ $Y=1.915 $X2=6.885 $Y2=2.115
r152 3 43 600 $w=1.7e-07 $l=9.95214e-07 $layer=licon1_PDIFF $count=1 $X=4.52
+ $Y=1.865 $X2=4.655 $Y2=2.795
r153 2 27 91 $w=1.7e-07 $l=2.67862e-07 $layer=licon1_NDIFF $count=2 $X=6.665
+ $Y=0.605 $X2=6.87 $Y2=0.75
r154 1 39 182 $w=1.7e-07 $l=2.26164e-07 $layer=licon1_NDIFF $count=1 $X=4.485
+ $Y=0.27 $X2=4.65 $Y2=0.415
.ends

.subckt PM_SKY130_FD_SC_HS__XNOR3_1%X 1 2 9 11 15 16 17 28
c22 16 0 1.63453e-19 $X=0.24 $Y=0.555
r23 21 28 2.0808 $w=3.58e-07 $l=6.5e-08 $layer=LI1_cond $X=0.265 $Y=0.99
+ $X2=0.265 $Y2=0.925
r24 17 30 8.67109 $w=3.58e-07 $l=1.7e-07 $layer=LI1_cond $X=0.265 $Y=1 $X2=0.265
+ $Y2=1.17
r25 17 21 0.320123 $w=3.58e-07 $l=1e-08 $layer=LI1_cond $X=0.265 $Y=1 $X2=0.265
+ $Y2=0.99
r26 17 28 0.320123 $w=3.58e-07 $l=1e-08 $layer=LI1_cond $X=0.265 $Y=0.915
+ $X2=0.265 $Y2=0.925
r27 16 17 11.5244 $w=3.58e-07 $l=3.6e-07 $layer=LI1_cond $X=0.265 $Y=0.555
+ $X2=0.265 $Y2=0.915
r28 15 30 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=0.17 $Y=1.84
+ $X2=0.17 $Y2=1.17
r29 11 13 34.5733 $w=2.68e-07 $l=8.1e-07 $layer=LI1_cond $X=0.22 $Y=2.005
+ $X2=0.22 $Y2=2.815
r30 9 15 7.33542 $w=2.68e-07 $l=1.35e-07 $layer=LI1_cond $X=0.22 $Y=1.975
+ $X2=0.22 $Y2=1.84
r31 9 11 1.28049 $w=2.68e-07 $l=3e-08 $layer=LI1_cond $X=0.22 $Y=1.975 $X2=0.22
+ $Y2=2.005
r32 2 13 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.27 $Y2=2.815
r33 2 11 400 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.27 $Y2=2.005
r34 1 16 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.49 $X2=0.28 $Y2=0.635
.ends

.subckt PM_SKY130_FD_SC_HS__XNOR3_1%VPWR 1 2 3 12 16 20 22 24 29 37 47 48 51 54
+ 57
c74 29 0 1.73622e-19 $X=3.395 $Y=3.33
c75 20 0 1.42592e-19 $X=7.425 $Y=2.375
r76 57 58 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r77 54 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r78 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r79 48 58 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=3.33
+ $X2=7.44 $Y2=3.33
r80 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r81 45 57 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.59 $Y=3.33
+ $X2=7.425 $Y2=3.33
r82 45 47 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=7.59 $Y=3.33
+ $X2=7.92 $Y2=3.33
r83 44 58 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=7.44 $Y2=3.33
r84 43 44 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r85 40 43 187.893 $w=1.68e-07 $l=2.88e-06 $layer=LI1_cond $X=4.08 $Y=3.33
+ $X2=6.96 $Y2=3.33
r86 38 54 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.725 $Y=3.33
+ $X2=3.56 $Y2=3.33
r87 38 40 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=3.725 $Y=3.33
+ $X2=4.08 $Y2=3.33
r88 37 57 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.26 $Y=3.33
+ $X2=7.425 $Y2=3.33
r89 37 43 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=7.26 $Y=3.33 $X2=6.96
+ $Y2=3.33
r90 36 55 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=3.6 $Y2=3.33
r91 35 36 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r92 33 36 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=3.12 $Y2=3.33
r93 33 52 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r94 32 35 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=1.2 $Y=3.33
+ $X2=3.12 $Y2=3.33
r95 32 33 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r96 30 51 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.805 $Y=3.33
+ $X2=0.68 $Y2=3.33
r97 30 32 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=0.805 $Y=3.33
+ $X2=1.2 $Y2=3.33
r98 29 54 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.395 $Y=3.33
+ $X2=3.56 $Y2=3.33
r99 29 35 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=3.395 $Y=3.33
+ $X2=3.12 $Y2=3.33
r100 27 52 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r101 26 27 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r102 24 51 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.555 $Y=3.33
+ $X2=0.68 $Y2=3.33
r103 24 26 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=0.555 $Y=3.33
+ $X2=0.24 $Y2=3.33
r104 22 44 0.802756 $w=4.9e-07 $l=2.88e-06 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=6.96 $Y2=3.33
r105 22 55 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=3.6 $Y2=3.33
r106 22 40 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r107 18 57 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.425 $Y=3.245
+ $X2=7.425 $Y2=3.33
r108 18 20 30.3826 $w=3.28e-07 $l=8.7e-07 $layer=LI1_cond $X=7.425 $Y=3.245
+ $X2=7.425 $Y2=2.375
r109 14 54 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.56 $Y=3.245
+ $X2=3.56 $Y2=3.33
r110 14 16 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=3.56 $Y=3.245
+ $X2=3.56 $Y2=2.875
r111 10 51 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=3.245
+ $X2=0.68 $Y2=3.33
r112 10 12 36.4172 $w=2.48e-07 $l=7.9e-07 $layer=LI1_cond $X=0.68 $Y=3.245
+ $X2=0.68 $Y2=2.455
r113 3 20 300 $w=1.7e-07 $l=5.6542e-07 $layer=licon1_PDIFF $count=2 $X=7.19
+ $Y=1.915 $X2=7.425 $Y2=2.375
r114 2 16 600 $w=1.7e-07 $l=1.10043e-06 $layer=licon1_PDIFF $count=1 $X=3.425
+ $Y=1.84 $X2=3.56 $Y2=2.875
r115 1 12 300 $w=1.7e-07 $l=6.85912e-07 $layer=licon1_PDIFF $count=2 $X=0.57
+ $Y=1.84 $X2=0.72 $Y2=2.455
.ends

.subckt PM_SKY130_FD_SC_HS__XNOR3_1%A_363_394# 1 2 3 4 15 17 18 20 22 23 27 29
+ 33 38 39 40
c130 29 0 4.37781e-20 $X=6.255 $Y=0.68
c131 23 0 1.66544e-19 $X=5.015 $Y=2.455
r132 39 40 7.99654 $w=2.43e-07 $l=1.7e-07 $layer=LI1_cond $X=5.01 $Y=0.717
+ $X2=5.18 $Y2=0.717
r133 36 37 13.7351 $w=4.53e-07 $l=5.1e-07 $layer=LI1_cond $X=2.93 $Y=0.67
+ $X2=3.44 $Y2=0.67
r134 31 33 11.5244 $w=2.78e-07 $l=2.8e-07 $layer=LI1_cond $X=6.395 $Y=0.765
+ $X2=6.395 $Y2=1.045
r135 29 31 7.36005 $w=1.7e-07 $l=1.77482e-07 $layer=LI1_cond $X=6.255 $Y=0.68
+ $X2=6.395 $Y2=0.765
r136 29 40 70.1337 $w=1.68e-07 $l=1.075e-06 $layer=LI1_cond $X=6.255 $Y=0.68
+ $X2=5.18 $Y2=0.68
r137 25 27 16.1342 $w=2.48e-07 $l=3.5e-07 $layer=LI1_cond $X=5.14 $Y=2.37
+ $X2=5.14 $Y2=2.02
r138 24 38 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.525 $Y=2.455
+ $X2=3.44 $Y2=2.455
r139 23 25 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=5.015 $Y=2.455
+ $X2=5.14 $Y2=2.37
r140 23 24 97.2086 $w=1.68e-07 $l=1.49e-06 $layer=LI1_cond $X=5.015 $Y=2.455
+ $X2=3.525 $Y2=2.455
r141 22 37 7.27104 $w=4.53e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.525 $Y=0.755
+ $X2=3.44 $Y2=0.67
r142 22 39 96.8824 $w=1.68e-07 $l=1.485e-06 $layer=LI1_cond $X=3.525 $Y=0.755
+ $X2=5.01 $Y2=0.755
r143 20 38 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.44 $Y=2.37
+ $X2=3.44 $Y2=2.455
r144 19 37 6.54142 $w=1.7e-07 $l=3e-07 $layer=LI1_cond $X=3.44 $Y=0.97 $X2=3.44
+ $Y2=0.67
r145 19 20 91.3369 $w=1.68e-07 $l=1.4e-06 $layer=LI1_cond $X=3.44 $Y=0.97
+ $X2=3.44 $Y2=2.37
r146 17 38 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.355 $Y=2.455
+ $X2=3.44 $Y2=2.455
r147 17 18 80.246 $w=1.68e-07 $l=1.23e-06 $layer=LI1_cond $X=3.355 $Y=2.455
+ $X2=2.125 $Y2=2.455
r148 13 18 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=2 $Y=2.37
+ $X2=2.125 $Y2=2.455
r149 13 15 11.7549 $w=2.48e-07 $l=2.55e-07 $layer=LI1_cond $X=2 $Y=2.37 $X2=2
+ $Y2=2.115
r150 4 27 300 $w=1.7e-07 $l=2.17428e-07 $layer=licon1_PDIFF $count=2 $X=5.03
+ $Y=1.865 $X2=5.18 $Y2=2.02
r151 3 15 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=1.815
+ $Y=1.97 $X2=1.96 $Y2=2.115
r152 2 33 182 $w=1.7e-07 $l=3.05778e-07 $layer=licon1_NDIFF $count=1 $X=6.17
+ $Y=0.825 $X2=6.375 $Y2=1.045
r153 1 36 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.79
+ $Y=0.37 $X2=2.93 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__XNOR3_1%A_371_74# 1 2 3 4 15 17 20 21 25 26 27 28 31
+ 34 37 38 44 47
c128 25 0 2.79465e-19 $X=5.52 $Y=1.41
r129 47 48 2.97244 $w=4.38e-07 $l=8.5e-08 $layer=LI1_cond $X=2.055 $Y=1.225
+ $X2=2.055 $Y2=1.14
r130 45 51 9.95397 $w=2.39e-07 $l=1.95e-07 $layer=LI1_cond $X=5.46 $Y=1.295
+ $X2=5.46 $Y2=1.1
r131 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=1.295
+ $X2=5.52 $Y2=1.295
r132 41 47 1.83343 $w=4.38e-07 $l=7e-08 $layer=LI1_cond $X=2.055 $Y=1.295
+ $X2=2.055 $Y2=1.225
r133 40 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=1.295
+ $X2=2.16 $Y2=1.295
r134 38 40 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.305 $Y=1.295
+ $X2=2.16 $Y2=1.295
r135 37 44 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.375 $Y=1.295
+ $X2=5.52 $Y2=1.295
r136 37 38 3.7995 $w=1.4e-07 $l=3.07e-06 $layer=MET1_cond $X=5.375 $Y=1.295
+ $X2=2.305 $Y2=1.295
r137 29 31 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=6.165 $Y=1.935
+ $X2=6.165 $Y2=2.195
r138 27 29 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.08 $Y=1.85
+ $X2=6.165 $Y2=1.935
r139 27 28 30.9893 $w=1.68e-07 $l=4.75e-07 $layer=LI1_cond $X=6.08 $Y=1.85
+ $X2=5.605 $Y2=1.85
r140 26 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.52 $Y=1.765
+ $X2=5.605 $Y2=1.85
r141 25 45 6.90437 $w=2.39e-07 $l=1.41863e-07 $layer=LI1_cond $X=5.52 $Y=1.41
+ $X2=5.46 $Y2=1.295
r142 25 26 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=5.52 $Y=1.41
+ $X2=5.52 $Y2=1.765
r143 21 51 2.73298 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=5.315 $Y=1.1
+ $X2=5.46 $Y2=1.1
r144 21 23 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=5.315 $Y=1.1
+ $X2=5.25 $Y2=1.1
r145 20 34 0.716491 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.1 $Y=2.03
+ $X2=3.015 $Y2=2.115
r146 19 20 46.9733 $w=1.68e-07 $l=7.2e-07 $layer=LI1_cond $X=3.1 $Y=1.31 $X2=3.1
+ $Y2=2.03
r147 18 47 6.36164 $w=1.7e-07 $l=2.2e-07 $layer=LI1_cond $X=2.275 $Y=1.225
+ $X2=2.055 $Y2=1.225
r148 17 19 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.015 $Y=1.225
+ $X2=3.1 $Y2=1.31
r149 17 18 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=3.015 $Y=1.225
+ $X2=2.275 $Y2=1.225
r150 15 48 11.5244 $w=3.28e-07 $l=3.3e-07 $layer=LI1_cond $X=2 $Y=0.81 $X2=2
+ $Y2=1.14
r151 4 31 600 $w=1.7e-07 $l=3.46987e-07 $layer=licon1_PDIFF $count=1 $X=6.015
+ $Y=1.915 $X2=6.165 $Y2=2.195
r152 3 34 600 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=2.865
+ $Y=1.97 $X2=3.015 $Y2=2.115
r153 2 23 182 $w=1.7e-07 $l=5.88643e-07 $layer=licon1_NDIFF $count=1 $X=5.045
+ $Y=0.605 $X2=5.25 $Y2=1.1
r154 1 15 182 $w=1.7e-07 $l=5.07346e-07 $layer=licon1_NDIFF $count=1 $X=1.855
+ $Y=0.37 $X2=2 $Y2=0.81
.ends

.subckt PM_SKY130_FD_SC_HS__XNOR3_1%A_1113_383# 1 2 3 4 15 17 18 19 20 22 23 25
+ 29 35 36 37 43 44 47
c118 36 0 1.54564e-19 $X=7.775 $Y=1.295
c119 19 0 1.78665e-19 $X=6.42 $Y=1.51
r120 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=1.295
+ $X2=7.92 $Y2=1.295
r121 40 47 7.24924 $w=3.08e-07 $l=1.95e-07 $layer=LI1_cond $X=5.93 $Y=1.295
+ $X2=5.93 $Y2=1.1
r122 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=1.295 $X2=6
+ $Y2=1.295
r123 37 39 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.145 $Y=1.295
+ $X2=6 $Y2=1.295
r124 36 43 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=7.775 $Y=1.295
+ $X2=7.92 $Y2=1.295
r125 36 37 2.01732 $w=1.4e-07 $l=1.63e-06 $layer=MET1_cond $X=7.775 $Y=1.295
+ $X2=6.145 $Y2=1.295
r126 35 44 1.92074 $w=2.38e-07 $l=4e-08 $layer=LI1_cond $X=7.955 $Y=1.255
+ $X2=7.955 $Y2=1.295
r127 33 44 42.9765 $w=2.38e-07 $l=8.95e-07 $layer=LI1_cond $X=7.955 $Y=2.19
+ $X2=7.955 $Y2=1.295
r128 31 40 4.83283 $w=3.08e-07 $l=1.3e-07 $layer=LI1_cond $X=5.93 $Y=1.425
+ $X2=5.93 $Y2=1.295
r129 27 35 6.02978 $w=2.78e-07 $l=1.4e-07 $layer=LI1_cond $X=7.935 $Y=1.115
+ $X2=7.935 $Y2=1.255
r130 27 29 15.0229 $w=2.78e-07 $l=3.65e-07 $layer=LI1_cond $X=7.935 $Y=1.115
+ $X2=7.935 $Y2=0.75
r131 23 33 6.0629 $w=2.83e-07 $l=1.42e-07 $layer=LI1_cond $X=7.932 $Y=2.332
+ $X2=7.932 $Y2=2.19
r132 23 25 0.930042 $w=2.83e-07 $l=2.3e-08 $layer=LI1_cond $X=7.932 $Y=2.332
+ $X2=7.932 $Y2=2.355
r133 21 22 63.2834 $w=1.68e-07 $l=9.7e-07 $layer=LI1_cond $X=6.505 $Y=1.595
+ $X2=6.505 $Y2=2.565
r134 20 31 7.59919 $w=1.7e-07 $l=1.92873e-07 $layer=LI1_cond $X=6.085 $Y=1.51
+ $X2=5.93 $Y2=1.425
r135 19 21 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.42 $Y=1.51
+ $X2=6.505 $Y2=1.595
r136 19 20 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=6.42 $Y=1.51
+ $X2=6.085 $Y2=1.51
r137 17 22 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.42 $Y=2.65
+ $X2=6.505 $Y2=2.565
r138 17 18 35.2299 $w=1.68e-07 $l=5.4e-07 $layer=LI1_cond $X=6.42 $Y=2.65
+ $X2=5.88 $Y2=2.65
r139 13 18 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=5.715 $Y=2.565
+ $X2=5.88 $Y2=2.65
r140 13 15 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=5.715 $Y=2.565
+ $X2=5.715 $Y2=2.27
r141 4 25 300 $w=1.7e-07 $l=5.0951e-07 $layer=licon1_PDIFF $count=2 $X=7.725
+ $Y=1.915 $X2=7.875 $Y2=2.355
r142 3 15 600 $w=1.7e-07 $l=4.23409e-07 $layer=licon1_PDIFF $count=1 $X=5.565
+ $Y=1.915 $X2=5.715 $Y2=2.27
r143 2 29 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=7.74
+ $Y=0.605 $X2=7.88 $Y2=0.75
r144 1 47 182 $w=1.7e-07 $l=6.07268e-07 $layer=licon1_NDIFF $count=1 $X=5.61
+ $Y=0.605 $X2=5.86 $Y2=1.1
.ends

.subckt PM_SKY130_FD_SC_HS__XNOR3_1%VGND 1 2 3 12 16 20 22 24 29 37 47 48 51 54
+ 57
r72 57 58 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=0 $X2=7.44
+ $Y2=0
r73 54 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r74 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r75 48 58 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=0 $X2=7.44
+ $Y2=0
r76 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=0 $X2=7.92
+ $Y2=0
r77 45 57 9.97069 $w=1.7e-07 $l=2.05e-07 $layer=LI1_cond $X=7.615 $Y=0 $X2=7.41
+ $Y2=0
r78 45 47 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=7.615 $Y=0 $X2=7.92
+ $Y2=0
r79 44 58 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=0 $X2=7.44
+ $Y2=0
r80 43 44 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=6.96 $Y=0
+ $X2=6.96 $Y2=0
r81 40 43 187.893 $w=1.68e-07 $l=2.88e-06 $layer=LI1_cond $X=4.08 $Y=0 $X2=6.96
+ $Y2=0
r82 38 54 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.725 $Y=0 $X2=3.56
+ $Y2=0
r83 38 40 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=3.725 $Y=0 $X2=4.08
+ $Y2=0
r84 37 57 9.97069 $w=1.7e-07 $l=2.05e-07 $layer=LI1_cond $X=7.205 $Y=0 $X2=7.41
+ $Y2=0
r85 37 43 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=7.205 $Y=0 $X2=6.96
+ $Y2=0
r86 36 55 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=3.6
+ $Y2=0
r87 35 36 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r88 33 36 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=1.2 $Y=0 $X2=3.12
+ $Y2=0
r89 33 52 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r90 32 35 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=1.2 $Y=0 $X2=3.12
+ $Y2=0
r91 32 33 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r92 30 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.955 $Y=0 $X2=0.79
+ $Y2=0
r93 30 32 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=0.955 $Y=0 $X2=1.2
+ $Y2=0
r94 29 54 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.395 $Y=0 $X2=3.56
+ $Y2=0
r95 29 35 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=3.395 $Y=0 $X2=3.12
+ $Y2=0
r96 27 52 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r97 26 27 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r98 24 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.625 $Y=0 $X2=0.79
+ $Y2=0
r99 24 26 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=0.625 $Y=0 $X2=0.24
+ $Y2=0
r100 22 44 0.802756 $w=4.9e-07 $l=2.88e-06 $layer=MET1_cond $X=4.08 $Y=0
+ $X2=6.96 $Y2=0
r101 22 55 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=3.6
+ $Y2=0
r102 22 40 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=4.08 $Y=0
+ $X2=4.08 $Y2=0
r103 18 57 1.53834 $w=4.1e-07 $l=8.5e-08 $layer=LI1_cond $X=7.41 $Y=0.085
+ $X2=7.41 $Y2=0
r104 18 20 18.6921 $w=4.08e-07 $l=6.65e-07 $layer=LI1_cond $X=7.41 $Y=0.085
+ $X2=7.41 $Y2=0.75
r105 14 54 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.56 $Y=0.085
+ $X2=3.56 $Y2=0
r106 14 16 8.73063 $w=3.28e-07 $l=2.5e-07 $layer=LI1_cond $X=3.56 $Y=0.085
+ $X2=3.56 $Y2=0.335
r107 10 51 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.79 $Y=0.085
+ $X2=0.79 $Y2=0
r108 10 12 8.3814 $w=3.28e-07 $l=2.4e-07 $layer=LI1_cond $X=0.79 $Y=0.085
+ $X2=0.79 $Y2=0.325
r109 3 20 182 $w=1.7e-07 $l=3.14245e-07 $layer=licon1_NDIFF $count=1 $X=7.16
+ $Y=0.605 $X2=7.41 $Y2=0.75
r110 2 16 182 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=1 $X=3.415
+ $Y=0.19 $X2=3.56 $Y2=0.335
r111 1 12 182 $w=1.7e-07 $l=2.91033e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.49 $X2=0.79 $Y2=0.325
.ends

