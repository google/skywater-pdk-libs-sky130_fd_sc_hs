* File: sky130_fd_sc_hs__a221oi_4.pxi.spice
* Created: Thu Aug 27 20:26:11 2020
* 
x_PM_SKY130_FD_SC_HS__A221OI_4%C1 N_C1_c_158_n N_C1_M1002_g N_C1_M1015_g
+ N_C1_c_159_n N_C1_M1003_g N_C1_M1022_g N_C1_c_160_n N_C1_M1005_g N_C1_M1027_g
+ N_C1_c_161_n N_C1_M1009_g N_C1_M1039_g C1 C1 C1 N_C1_c_162_n N_C1_c_157_n
+ PM_SKY130_FD_SC_HS__A221OI_4%C1
x_PM_SKY130_FD_SC_HS__A221OI_4%A2 N_A2_c_241_n N_A2_M1016_g N_A2_M1004_g
+ N_A2_M1007_g N_A2_c_242_n N_A2_M1017_g N_A2_M1018_g N_A2_c_243_n N_A2_M1021_g
+ N_A2_M1019_g N_A2_c_244_n N_A2_M1025_g A2 A2 A2 A2 A2 N_A2_c_239_n
+ N_A2_c_240_n PM_SKY130_FD_SC_HS__A221OI_4%A2
x_PM_SKY130_FD_SC_HS__A221OI_4%A1 N_A1_M1012_g N_A1_c_325_n N_A1_M1000_g
+ N_A1_M1024_g N_A1_c_326_n N_A1_M1026_g N_A1_M1033_g N_A1_c_327_n N_A1_M1029_g
+ N_A1_M1034_g N_A1_c_328_n N_A1_M1037_g A1 A1 A1 A1 N_A1_c_324_n
+ PM_SKY130_FD_SC_HS__A221OI_4%A1
x_PM_SKY130_FD_SC_HS__A221OI_4%B1 N_B1_c_424_n N_B1_M1030_g N_B1_M1011_g
+ N_B1_c_425_n N_B1_M1031_g N_B1_M1014_g N_B1_c_426_n N_B1_M1032_g N_B1_M1028_g
+ N_B1_c_427_n N_B1_M1035_g N_B1_M1036_g B1 B1 B1 B1 N_B1_c_428_n N_B1_c_421_n
+ N_B1_c_422_n B1 N_B1_c_423_n PM_SKY130_FD_SC_HS__A221OI_4%B1
x_PM_SKY130_FD_SC_HS__A221OI_4%B2 N_B2_c_511_n N_B2_M1001_g N_B2_M1006_g
+ N_B2_c_512_n N_B2_M1010_g N_B2_M1008_g N_B2_c_513_n N_B2_M1013_g N_B2_M1020_g
+ N_B2_M1023_g N_B2_c_514_n N_B2_M1038_g B2 B2 B2 B2 N_B2_c_510_n
+ PM_SKY130_FD_SC_HS__A221OI_4%B2
x_PM_SKY130_FD_SC_HS__A221OI_4%Y N_Y_M1015_s N_Y_M1022_s N_Y_M1039_s N_Y_M1012_s
+ N_Y_M1033_s N_Y_M1011_s N_Y_M1028_s N_Y_M1002_s N_Y_M1003_s N_Y_M1009_s
+ N_Y_c_599_n N_Y_c_600_n N_Y_c_582_n N_Y_c_611_n N_Y_c_583_n N_Y_c_601_n
+ N_Y_c_584_n N_Y_c_602_n N_Y_c_585_n N_Y_c_586_n N_Y_c_724_p N_Y_c_587_n
+ N_Y_c_729_p N_Y_c_603_n N_Y_c_588_n N_Y_c_589_n N_Y_c_590_n N_Y_c_591_n
+ N_Y_c_592_n N_Y_c_593_n N_Y_c_594_n N_Y_c_595_n Y Y Y Y Y Y Y N_Y_c_597_n
+ N_Y_c_598_n PM_SKY130_FD_SC_HS__A221OI_4%Y
x_PM_SKY130_FD_SC_HS__A221OI_4%A_114_368# N_A_114_368#_M1002_d
+ N_A_114_368#_M1005_d N_A_114_368#_M1030_d N_A_114_368#_M1032_d
+ N_A_114_368#_M1001_s N_A_114_368#_M1013_s N_A_114_368#_c_745_n
+ N_A_114_368#_c_748_n N_A_114_368#_c_749_n N_A_114_368#_c_813_n
+ N_A_114_368#_c_744_n N_A_114_368#_c_773_n N_A_114_368#_c_777_n
+ N_A_114_368#_c_791_n N_A_114_368#_c_756_n N_A_114_368#_c_770_n
+ N_A_114_368#_c_783_n N_A_114_368#_c_788_n N_A_114_368#_c_801_n
+ PM_SKY130_FD_SC_HS__A221OI_4%A_114_368#
x_PM_SKY130_FD_SC_HS__A221OI_4%A_531_368# N_A_531_368#_M1016_s
+ N_A_531_368#_M1017_s N_A_531_368#_M1025_s N_A_531_368#_M1026_s
+ N_A_531_368#_M1037_s N_A_531_368#_M1031_s N_A_531_368#_M1035_s
+ N_A_531_368#_M1010_d N_A_531_368#_M1038_d N_A_531_368#_c_863_n
+ N_A_531_368#_c_865_n N_A_531_368#_c_875_n N_A_531_368#_c_877_n
+ N_A_531_368#_c_879_n N_A_531_368#_c_880_n N_A_531_368#_c_849_n
+ N_A_531_368#_c_850_n N_A_531_368#_c_915_n N_A_531_368#_c_851_n
+ N_A_531_368#_c_918_n N_A_531_368#_c_852_n N_A_531_368#_c_921_n
+ N_A_531_368#_c_853_n N_A_531_368#_c_854_n N_A_531_368#_c_855_n
+ N_A_531_368#_c_856_n N_A_531_368#_c_857_n N_A_531_368#_c_858_n
+ N_A_531_368#_c_859_n N_A_531_368#_c_860_n N_A_531_368#_c_861_n
+ PM_SKY130_FD_SC_HS__A221OI_4%A_531_368#
x_PM_SKY130_FD_SC_HS__A221OI_4%VPWR N_VPWR_M1016_d N_VPWR_M1021_d N_VPWR_M1000_d
+ N_VPWR_M1029_d N_VPWR_c_971_n N_VPWR_c_972_n N_VPWR_c_973_n N_VPWR_c_974_n
+ N_VPWR_c_975_n N_VPWR_c_976_n N_VPWR_c_977_n N_VPWR_c_978_n N_VPWR_c_979_n
+ VPWR N_VPWR_c_980_n N_VPWR_c_981_n N_VPWR_c_970_n N_VPWR_c_983_n
+ N_VPWR_c_984_n PM_SKY130_FD_SC_HS__A221OI_4%VPWR
x_PM_SKY130_FD_SC_HS__A221OI_4%VGND N_VGND_M1015_d N_VGND_M1027_d N_VGND_M1004_d
+ N_VGND_M1018_d N_VGND_M1006_s N_VGND_M1020_s N_VGND_c_1085_n N_VGND_c_1086_n
+ N_VGND_c_1087_n N_VGND_c_1088_n N_VGND_c_1089_n N_VGND_c_1090_n VGND
+ N_VGND_c_1091_n N_VGND_c_1092_n N_VGND_c_1093_n N_VGND_c_1094_n
+ N_VGND_c_1095_n N_VGND_c_1096_n N_VGND_c_1097_n N_VGND_c_1098_n
+ N_VGND_c_1099_n N_VGND_c_1100_n N_VGND_c_1101_n N_VGND_c_1102_n
+ N_VGND_c_1103_n PM_SKY130_FD_SC_HS__A221OI_4%VGND
x_PM_SKY130_FD_SC_HS__A221OI_4%A_534_74# N_A_534_74#_M1004_s N_A_534_74#_M1007_s
+ N_A_534_74#_M1019_s N_A_534_74#_M1024_d N_A_534_74#_M1034_d
+ N_A_534_74#_c_1225_n N_A_534_74#_c_1234_n N_A_534_74#_c_1226_n
+ N_A_534_74#_c_1227_n N_A_534_74#_c_1238_n N_A_534_74#_c_1241_n
+ N_A_534_74#_c_1242_n N_A_534_74#_c_1228_n N_A_534_74#_c_1229_n
+ N_A_534_74#_c_1247_n N_A_534_74#_c_1230_n N_A_534_74#_c_1279_n
+ N_A_534_74#_c_1231_n N_A_534_74#_c_1232_n
+ PM_SKY130_FD_SC_HS__A221OI_4%A_534_74#
x_PM_SKY130_FD_SC_HS__A221OI_4%A_1326_74# N_A_1326_74#_M1011_d
+ N_A_1326_74#_M1014_d N_A_1326_74#_M1036_d N_A_1326_74#_M1008_d
+ N_A_1326_74#_M1023_d N_A_1326_74#_c_1311_n N_A_1326_74#_c_1312_n
+ N_A_1326_74#_c_1313_n N_A_1326_74#_c_1314_n N_A_1326_74#_c_1315_n
+ N_A_1326_74#_c_1316_n N_A_1326_74#_c_1317_n N_A_1326_74#_c_1318_n
+ N_A_1326_74#_c_1319_n N_A_1326_74#_c_1320_n N_A_1326_74#_c_1321_n
+ PM_SKY130_FD_SC_HS__A221OI_4%A_1326_74#
cc_1 VNB N_C1_M1015_g 0.0260102f $X=-0.19 $Y=-0.245 $X2=0.625 $Y2=0.74
cc_2 VNB N_C1_M1022_g 0.0209446f $X=-0.19 $Y=-0.245 $X2=1.055 $Y2=0.74
cc_3 VNB N_C1_M1027_g 0.0209433f $X=-0.19 $Y=-0.245 $X2=1.485 $Y2=0.74
cc_4 VNB N_C1_M1039_g 0.0273441f $X=-0.19 $Y=-0.245 $X2=1.915 $Y2=0.74
cc_5 VNB N_C1_c_157_n 0.0892611f $X=-0.19 $Y=-0.245 $X2=1.845 $Y2=1.542
cc_6 VNB N_A2_M1004_g 0.0300605f $X=-0.19 $Y=-0.245 $X2=0.625 $Y2=0.74
cc_7 VNB N_A2_M1007_g 0.021821f $X=-0.19 $Y=-0.245 $X2=0.945 $Y2=2.4
cc_8 VNB N_A2_M1018_g 0.021821f $X=-0.19 $Y=-0.245 $X2=1.395 $Y2=2.4
cc_9 VNB N_A2_M1019_g 0.0221891f $X=-0.19 $Y=-0.245 $X2=1.845 $Y2=2.4
cc_10 VNB N_A2_c_239_n 0.0152156f $X=-0.19 $Y=-0.245 $X2=1.2 $Y2=1.565
cc_11 VNB N_A2_c_240_n 0.074481f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A1_M1012_g 0.0205994f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.4
cc_13 VNB N_A1_M1024_g 0.0203905f $X=-0.19 $Y=-0.245 $X2=0.945 $Y2=2.4
cc_14 VNB N_A1_M1033_g 0.0203905f $X=-0.19 $Y=-0.245 $X2=1.395 $Y2=2.4
cc_15 VNB N_A1_M1034_g 0.0272298f $X=-0.19 $Y=-0.245 $X2=1.845 $Y2=2.4
cc_16 VNB A1 0.00357027f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A1_c_324_n 0.091885f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.565
cc_18 VNB N_B1_M1011_g 0.0292211f $X=-0.19 $Y=-0.245 $X2=0.625 $Y2=0.74
cc_19 VNB N_B1_M1014_g 0.0230075f $X=-0.19 $Y=-0.245 $X2=1.055 $Y2=0.74
cc_20 VNB N_B1_M1028_g 0.0230075f $X=-0.19 $Y=-0.245 $X2=1.485 $Y2=0.74
cc_21 VNB N_B1_M1036_g 0.0238795f $X=-0.19 $Y=-0.245 $X2=1.915 $Y2=0.74
cc_22 VNB N_B1_c_421_n 0.0728395f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_B1_c_422_n 0.00109917f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_B1_c_423_n 0.0026459f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_B2_M1006_g 0.0230056f $X=-0.19 $Y=-0.245 $X2=0.625 $Y2=0.74
cc_26 VNB N_B2_M1008_g 0.0224899f $X=-0.19 $Y=-0.245 $X2=1.055 $Y2=0.74
cc_27 VNB N_B2_M1020_g 0.0224899f $X=-0.19 $Y=-0.245 $X2=1.485 $Y2=0.74
cc_28 VNB N_B2_M1023_g 0.0318708f $X=-0.19 $Y=-0.245 $X2=1.845 $Y2=2.4
cc_29 VNB B2 0.00453471f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_B2_c_510_n 0.0794465f $X=-0.19 $Y=-0.245 $X2=0.69 $Y2=1.565
cc_31 VNB N_Y_c_582_n 0.00316432f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_Y_c_583_n 0.00178908f $X=-0.19 $Y=-0.245 $X2=1.055 $Y2=1.542
cc_33 VNB N_Y_c_584_n 0.00459798f $X=-0.19 $Y=-0.245 $X2=1.71 $Y2=1.515
cc_34 VNB N_Y_c_585_n 0.0102558f $X=-0.19 $Y=-0.245 $X2=1.2 $Y2=1.565
cc_35 VNB N_Y_c_586_n 0.0305363f $X=-0.19 $Y=-0.245 $X2=1.68 $Y2=1.565
cc_36 VNB N_Y_c_587_n 0.00304134f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_Y_c_588_n 0.00126364f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_Y_c_589_n 0.00542103f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_Y_c_590_n 0.00141635f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_Y_c_591_n 0.00141635f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_Y_c_592_n 0.00317705f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_Y_c_593_n 0.00766831f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_Y_c_594_n 0.00480063f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_Y_c_595_n 0.0106677f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB Y 0.0250032f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_Y_c_597_n 0.0330268f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_Y_c_598_n 0.0113079f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_VPWR_c_970_n 0.442315f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_VGND_c_1085_n 0.00323505f $X=-0.19 $Y=-0.245 $X2=1.845 $Y2=2.4
cc_50 VNB N_VGND_c_1086_n 0.00323505f $X=-0.19 $Y=-0.245 $X2=1.915 $Y2=0.74
cc_51 VNB N_VGND_c_1087_n 0.00323505f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=1.58
cc_52 VNB N_VGND_c_1088_n 0.00323505f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.542
cc_53 VNB N_VGND_c_1089_n 0.00323505f $X=-0.19 $Y=-0.245 $X2=0.69 $Y2=1.515
cc_54 VNB N_VGND_c_1090_n 0.00323505f $X=-0.19 $Y=-0.245 $X2=1.485 $Y2=1.542
cc_55 VNB N_VGND_c_1091_n 0.0151736f $X=-0.19 $Y=-0.245 $X2=1.845 $Y2=1.542
cc_56 VNB N_VGND_c_1092_n 0.0331279f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_VGND_c_1093_n 0.0138836f $X=-0.19 $Y=-0.245 $X2=1.71 $Y2=1.565
cc_58 VNB N_VGND_c_1094_n 0.109557f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_VGND_c_1095_n 0.0151736f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_VGND_c_1096_n 0.0200958f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_VGND_c_1097_n 0.562213f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_VGND_c_1098_n 0.0264764f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_VGND_c_1099_n 0.00604233f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_VGND_c_1100_n 0.00601569f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_VGND_c_1101_n 0.00601569f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_VGND_c_1102_n 0.00604233f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_VGND_c_1103_n 0.00604233f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_A_534_74#_c_1225_n 0.00687082f $X=-0.19 $Y=-0.245 $X2=1.485 $Y2=1.32
cc_69 VNB N_A_534_74#_c_1226_n 0.00231144f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_A_534_74#_c_1227_n 0.00178442f $X=-0.19 $Y=-0.245 $X2=1.845 $Y2=2.4
cc_71 VNB N_A_534_74#_c_1228_n 0.00215453f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_A_534_74#_c_1229_n 0.00230059f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_A_534_74#_c_1230_n 0.00215453f $X=-0.19 $Y=-0.245 $X2=0.69 $Y2=1.515
cc_74 VNB N_A_534_74#_c_1231_n 0.00220113f $X=-0.19 $Y=-0.245 $X2=1.485
+ $Y2=1.542
cc_75 VNB N_A_534_74#_c_1232_n 0.0065966f $X=-0.19 $Y=-0.245 $X2=1.71 $Y2=1.542
cc_76 VNB N_A_1326_74#_c_1311_n 0.00289325f $X=-0.19 $Y=-0.245 $X2=1.485
+ $Y2=1.32
cc_77 VNB N_A_1326_74#_c_1312_n 0.0016059f $X=-0.19 $Y=-0.245 $X2=1.485 $Y2=0.74
cc_78 VNB N_A_1326_74#_c_1313_n 0.00307486f $X=-0.19 $Y=-0.245 $X2=1.845 $Y2=2.4
cc_79 VNB N_A_1326_74#_c_1314_n 0.00205775f $X=-0.19 $Y=-0.245 $X2=1.915
+ $Y2=1.32
cc_80 VNB N_A_1326_74#_c_1315_n 0.00178908f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_81 VNB N_A_1326_74#_c_1316_n 0.0165052f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.58
cc_82 VNB N_A_1326_74#_c_1317_n 0.0270834f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_83 VNB N_A_1326_74#_c_1318_n 0.00597701f $X=-0.19 $Y=-0.245 $X2=0.69
+ $Y2=1.515
cc_84 VNB N_A_1326_74#_c_1319_n 0.00236184f $X=-0.19 $Y=-0.245 $X2=1.395
+ $Y2=1.542
cc_85 VNB N_A_1326_74#_c_1320_n 0.00228921f $X=-0.19 $Y=-0.245 $X2=1.485
+ $Y2=1.542
cc_86 VNB N_A_1326_74#_c_1321_n 0.00127131f $X=-0.19 $Y=-0.245 $X2=1.71
+ $Y2=1.515
cc_87 VPB N_C1_c_158_n 0.0170004f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.765
cc_88 VPB N_C1_c_159_n 0.0146573f $X=-0.19 $Y=1.66 $X2=0.945 $Y2=1.765
cc_89 VPB N_C1_c_160_n 0.0146598f $X=-0.19 $Y=1.66 $X2=1.395 $Y2=1.765
cc_90 VPB N_C1_c_161_n 0.0185593f $X=-0.19 $Y=1.66 $X2=1.845 $Y2=1.765
cc_91 VPB N_C1_c_162_n 0.00839222f $X=-0.19 $Y=1.66 $X2=1.71 $Y2=1.515
cc_92 VPB N_C1_c_157_n 0.0479059f $X=-0.19 $Y=1.66 $X2=1.845 $Y2=1.542
cc_93 VPB N_A2_c_241_n 0.0194207f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.765
cc_94 VPB N_A2_c_242_n 0.0155127f $X=-0.19 $Y=1.66 $X2=1.055 $Y2=0.74
cc_95 VPB N_A2_c_243_n 0.0155127f $X=-0.19 $Y=1.66 $X2=1.485 $Y2=0.74
cc_96 VPB N_A2_c_244_n 0.0159072f $X=-0.19 $Y=1.66 $X2=1.915 $Y2=0.74
cc_97 VPB N_A2_c_239_n 0.0202406f $X=-0.19 $Y=1.66 $X2=1.2 $Y2=1.565
cc_98 VPB N_A2_c_240_n 0.0476542f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_99 VPB N_A1_c_325_n 0.0157881f $X=-0.19 $Y=1.66 $X2=0.625 $Y2=0.74
cc_100 VPB N_A1_c_326_n 0.0155117f $X=-0.19 $Y=1.66 $X2=1.055 $Y2=0.74
cc_101 VPB N_A1_c_327_n 0.017015f $X=-0.19 $Y=1.66 $X2=1.485 $Y2=0.74
cc_102 VPB N_A1_c_328_n 0.0168058f $X=-0.19 $Y=1.66 $X2=1.915 $Y2=0.74
cc_103 VPB A1 0.0126664f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_104 VPB N_A1_c_324_n 0.055793f $X=-0.19 $Y=1.66 $X2=0.72 $Y2=1.565
cc_105 VPB N_B1_c_424_n 0.0147905f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.765
cc_106 VPB N_B1_c_425_n 0.014664f $X=-0.19 $Y=1.66 $X2=0.945 $Y2=1.765
cc_107 VPB N_B1_c_426_n 0.014664f $X=-0.19 $Y=1.66 $X2=1.395 $Y2=1.765
cc_108 VPB N_B1_c_427_n 0.0149102f $X=-0.19 $Y=1.66 $X2=1.845 $Y2=1.765
cc_109 VPB N_B1_c_428_n 0.00800034f $X=-0.19 $Y=1.66 $X2=0.69 $Y2=1.565
cc_110 VPB N_B1_c_421_n 0.046084f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_111 VPB N_B1_c_422_n 6.06119e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_112 VPB N_B1_c_423_n 0.00246497f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_113 VPB N_B2_c_511_n 0.0147911f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.765
cc_114 VPB N_B2_c_512_n 0.014664f $X=-0.19 $Y=1.66 $X2=0.945 $Y2=1.765
cc_115 VPB N_B2_c_513_n 0.0146632f $X=-0.19 $Y=1.66 $X2=1.395 $Y2=1.765
cc_116 VPB N_B2_c_514_n 0.0183915f $X=-0.19 $Y=1.66 $X2=1.915 $Y2=0.74
cc_117 VPB B2 0.0119499f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_118 VPB N_B2_c_510_n 0.0489233f $X=-0.19 $Y=1.66 $X2=0.69 $Y2=1.565
cc_119 VPB N_Y_c_599_n 0.00259172f $X=-0.19 $Y=1.66 $X2=1.595 $Y2=1.58
cc_120 VPB N_Y_c_600_n 0.00938462f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_121 VPB N_Y_c_601_n 0.00759038f $X=-0.19 $Y=1.66 $X2=1.485 $Y2=1.542
cc_122 VPB N_Y_c_602_n 0.00776005f $X=-0.19 $Y=1.66 $X2=0.69 $Y2=1.565
cc_123 VPB N_Y_c_603_n 0.0021839f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_124 VPB Y 0.049211f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_125 VPB N_A_114_368#_c_744_n 0.0208972f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_126 VPB N_A_531_368#_c_849_n 0.0026202f $X=-0.19 $Y=1.66 $X2=1.71 $Y2=1.515
cc_127 VPB N_A_531_368#_c_850_n 0.00192911f $X=-0.19 $Y=1.66 $X2=1.845 $Y2=1.542
cc_128 VPB N_A_531_368#_c_851_n 0.0026202f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_129 VPB N_A_531_368#_c_852_n 0.0026202f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_130 VPB N_A_531_368#_c_853_n 0.012233f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_131 VPB N_A_531_368#_c_854_n 0.0454805f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_132 VPB N_A_531_368#_c_855_n 0.0114591f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_133 VPB N_A_531_368#_c_856_n 0.00257417f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_134 VPB N_A_531_368#_c_857_n 0.00257417f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_135 VPB N_A_531_368#_c_858_n 0.00257417f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_136 VPB N_A_531_368#_c_859_n 0.00167433f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_137 VPB N_A_531_368#_c_860_n 0.00167433f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_138 VPB N_A_531_368#_c_861_n 0.00167433f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_139 VPB N_VPWR_c_971_n 0.00799266f $X=-0.19 $Y=1.66 $X2=1.395 $Y2=1.765
cc_140 VPB N_VPWR_c_972_n 0.0206041f $X=-0.19 $Y=1.66 $X2=1.395 $Y2=2.4
cc_141 VPB N_VPWR_c_973_n 0.00799266f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_142 VPB N_VPWR_c_974_n 0.00799266f $X=-0.19 $Y=1.66 $X2=1.915 $Y2=1.32
cc_143 VPB N_VPWR_c_975_n 0.0107095f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_144 VPB N_VPWR_c_976_n 0.0790487f $X=-0.19 $Y=1.66 $X2=1.595 $Y2=1.58
cc_145 VPB N_VPWR_c_977_n 0.00324402f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_146 VPB N_VPWR_c_978_n 0.0206041f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_147 VPB N_VPWR_c_979_n 0.00324402f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.542
cc_148 VPB N_VPWR_c_980_n 0.0196495f $X=-0.19 $Y=1.66 $X2=0.69 $Y2=1.565
cc_149 VPB N_VPWR_c_981_n 0.100392f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_150 VPB N_VPWR_c_970_n 0.122953f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_151 VPB N_VPWR_c_983_n 0.00324402f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_152 VPB N_VPWR_c_984_n 0.0088184f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_153 N_C1_c_161_n N_A2_c_239_n 2.77359e-19 $X=1.845 $Y=1.765 $X2=0 $Y2=0
cc_154 N_C1_c_162_n N_A2_c_239_n 0.0309808f $X=1.71 $Y=1.515 $X2=0 $Y2=0
cc_155 N_C1_c_157_n N_A2_c_239_n 0.00925123f $X=1.845 $Y=1.542 $X2=0 $Y2=0
cc_156 N_C1_c_158_n N_Y_c_599_n 0.0137046f $X=0.495 $Y=1.765 $X2=0 $Y2=0
cc_157 N_C1_c_159_n N_Y_c_599_n 0.0108414f $X=0.945 $Y=1.765 $X2=0 $Y2=0
cc_158 N_C1_M1015_g N_Y_c_582_n 0.0137752f $X=0.625 $Y=0.74 $X2=0 $Y2=0
cc_159 N_C1_M1022_g N_Y_c_582_n 0.0130918f $X=1.055 $Y=0.74 $X2=0 $Y2=0
cc_160 N_C1_c_162_n N_Y_c_582_n 0.0494694f $X=1.71 $Y=1.515 $X2=0 $Y2=0
cc_161 N_C1_c_157_n N_Y_c_582_n 0.00440402f $X=1.845 $Y=1.542 $X2=0 $Y2=0
cc_162 N_C1_c_158_n N_Y_c_611_n 6.04854e-19 $X=0.495 $Y=1.765 $X2=0 $Y2=0
cc_163 N_C1_c_159_n N_Y_c_611_n 0.00774844f $X=0.945 $Y=1.765 $X2=0 $Y2=0
cc_164 N_C1_c_160_n N_Y_c_611_n 0.00754637f $X=1.395 $Y=1.765 $X2=0 $Y2=0
cc_165 N_C1_c_161_n N_Y_c_611_n 5.52094e-19 $X=1.845 $Y=1.765 $X2=0 $Y2=0
cc_166 N_C1_M1022_g N_Y_c_583_n 3.92313e-19 $X=1.055 $Y=0.74 $X2=0 $Y2=0
cc_167 N_C1_M1027_g N_Y_c_583_n 3.92313e-19 $X=1.485 $Y=0.74 $X2=0 $Y2=0
cc_168 N_C1_c_160_n N_Y_c_601_n 0.0108414f $X=1.395 $Y=1.765 $X2=0 $Y2=0
cc_169 N_C1_c_161_n N_Y_c_601_n 0.0134708f $X=1.845 $Y=1.765 $X2=0 $Y2=0
cc_170 N_C1_M1027_g N_Y_c_584_n 0.0130918f $X=1.485 $Y=0.74 $X2=0 $Y2=0
cc_171 N_C1_M1039_g N_Y_c_584_n 0.0171665f $X=1.915 $Y=0.74 $X2=0 $Y2=0
cc_172 N_C1_c_162_n N_Y_c_584_n 0.039161f $X=1.71 $Y=1.515 $X2=0 $Y2=0
cc_173 N_C1_c_157_n N_Y_c_584_n 0.00236438f $X=1.845 $Y=1.542 $X2=0 $Y2=0
cc_174 N_C1_c_160_n N_Y_c_602_n 5.52094e-19 $X=1.395 $Y=1.765 $X2=0 $Y2=0
cc_175 N_C1_c_161_n N_Y_c_602_n 0.00766159f $X=1.845 $Y=1.765 $X2=0 $Y2=0
cc_176 N_C1_M1039_g N_Y_c_585_n 0.00159319f $X=1.915 $Y=0.74 $X2=0 $Y2=0
cc_177 N_C1_c_159_n N_Y_c_603_n 0.00175197f $X=0.945 $Y=1.765 $X2=0 $Y2=0
cc_178 N_C1_c_160_n N_Y_c_603_n 0.00175197f $X=1.395 $Y=1.765 $X2=0 $Y2=0
cc_179 N_C1_c_162_n N_Y_c_588_n 0.0146025f $X=1.71 $Y=1.515 $X2=0 $Y2=0
cc_180 N_C1_c_157_n N_Y_c_588_n 0.00247319f $X=1.845 $Y=1.542 $X2=0 $Y2=0
cc_181 N_C1_M1039_g N_Y_c_589_n 0.00372818f $X=1.915 $Y=0.74 $X2=0 $Y2=0
cc_182 N_C1_c_158_n Y 0.0102907f $X=0.495 $Y=1.765 $X2=0 $Y2=0
cc_183 N_C1_M1015_g Y 0.00485031f $X=0.625 $Y=0.74 $X2=0 $Y2=0
cc_184 N_C1_c_162_n Y 0.0351326f $X=1.71 $Y=1.515 $X2=0 $Y2=0
cc_185 N_C1_c_157_n Y 0.0135571f $X=1.845 $Y=1.542 $X2=0 $Y2=0
cc_186 N_C1_M1015_g N_Y_c_597_n 0.00159973f $X=0.625 $Y=0.74 $X2=0 $Y2=0
cc_187 N_C1_c_157_n N_Y_c_598_n 0.00445958f $X=1.845 $Y=1.542 $X2=0 $Y2=0
cc_188 N_C1_c_158_n N_A_114_368#_c_745_n 0.00203651f $X=0.495 $Y=1.765 $X2=0
+ $Y2=0
cc_189 N_C1_c_162_n N_A_114_368#_c_745_n 0.0210582f $X=1.71 $Y=1.515 $X2=0 $Y2=0
cc_190 N_C1_c_157_n N_A_114_368#_c_745_n 0.00136566f $X=1.845 $Y=1.542 $X2=0
+ $Y2=0
cc_191 N_C1_c_158_n N_A_114_368#_c_748_n 0.00828329f $X=0.495 $Y=1.765 $X2=0
+ $Y2=0
cc_192 N_C1_c_159_n N_A_114_368#_c_749_n 0.0126853f $X=0.945 $Y=1.765 $X2=0
+ $Y2=0
cc_193 N_C1_c_160_n N_A_114_368#_c_749_n 0.0126853f $X=1.395 $Y=1.765 $X2=0
+ $Y2=0
cc_194 N_C1_c_162_n N_A_114_368#_c_749_n 0.0446098f $X=1.71 $Y=1.515 $X2=0 $Y2=0
cc_195 N_C1_c_157_n N_A_114_368#_c_749_n 0.00130686f $X=1.845 $Y=1.542 $X2=0
+ $Y2=0
cc_196 N_C1_c_161_n N_A_114_368#_c_744_n 0.0159802f $X=1.845 $Y=1.765 $X2=0
+ $Y2=0
cc_197 N_C1_c_162_n N_A_114_368#_c_744_n 0.00914396f $X=1.71 $Y=1.515 $X2=0
+ $Y2=0
cc_198 N_C1_c_157_n N_A_114_368#_c_744_n 0.00112245f $X=1.845 $Y=1.542 $X2=0
+ $Y2=0
cc_199 N_C1_c_162_n N_A_114_368#_c_756_n 0.0183565f $X=1.71 $Y=1.515 $X2=0 $Y2=0
cc_200 N_C1_c_157_n N_A_114_368#_c_756_n 0.00129647f $X=1.845 $Y=1.542 $X2=0
+ $Y2=0
cc_201 N_C1_c_161_n N_A_531_368#_c_855_n 0.00115969f $X=1.845 $Y=1.765 $X2=0
+ $Y2=0
cc_202 N_C1_c_158_n N_VPWR_c_976_n 0.00278271f $X=0.495 $Y=1.765 $X2=0 $Y2=0
cc_203 N_C1_c_159_n N_VPWR_c_976_n 0.00278257f $X=0.945 $Y=1.765 $X2=0 $Y2=0
cc_204 N_C1_c_160_n N_VPWR_c_976_n 0.00278257f $X=1.395 $Y=1.765 $X2=0 $Y2=0
cc_205 N_C1_c_161_n N_VPWR_c_976_n 0.00278257f $X=1.845 $Y=1.765 $X2=0 $Y2=0
cc_206 N_C1_c_158_n N_VPWR_c_970_n 0.00357283f $X=0.495 $Y=1.765 $X2=0 $Y2=0
cc_207 N_C1_c_159_n N_VPWR_c_970_n 0.00353822f $X=0.945 $Y=1.765 $X2=0 $Y2=0
cc_208 N_C1_c_160_n N_VPWR_c_970_n 0.00353822f $X=1.395 $Y=1.765 $X2=0 $Y2=0
cc_209 N_C1_c_161_n N_VPWR_c_970_n 0.00358623f $X=1.845 $Y=1.765 $X2=0 $Y2=0
cc_210 N_C1_M1015_g N_VGND_c_1085_n 0.0137191f $X=0.625 $Y=0.74 $X2=0 $Y2=0
cc_211 N_C1_M1022_g N_VGND_c_1085_n 0.0106755f $X=1.055 $Y=0.74 $X2=0 $Y2=0
cc_212 N_C1_M1027_g N_VGND_c_1085_n 4.71636e-19 $X=1.485 $Y=0.74 $X2=0 $Y2=0
cc_213 N_C1_M1022_g N_VGND_c_1086_n 4.71636e-19 $X=1.055 $Y=0.74 $X2=0 $Y2=0
cc_214 N_C1_M1027_g N_VGND_c_1086_n 0.0106755f $X=1.485 $Y=0.74 $X2=0 $Y2=0
cc_215 N_C1_M1039_g N_VGND_c_1086_n 0.0137191f $X=1.915 $Y=0.74 $X2=0 $Y2=0
cc_216 N_C1_M1022_g N_VGND_c_1091_n 0.00383152f $X=1.055 $Y=0.74 $X2=0 $Y2=0
cc_217 N_C1_M1027_g N_VGND_c_1091_n 0.00383152f $X=1.485 $Y=0.74 $X2=0 $Y2=0
cc_218 N_C1_M1039_g N_VGND_c_1092_n 0.00383152f $X=1.915 $Y=0.74 $X2=0 $Y2=0
cc_219 N_C1_M1015_g N_VGND_c_1097_n 0.00761566f $X=0.625 $Y=0.74 $X2=0 $Y2=0
cc_220 N_C1_M1022_g N_VGND_c_1097_n 0.0075754f $X=1.055 $Y=0.74 $X2=0 $Y2=0
cc_221 N_C1_M1027_g N_VGND_c_1097_n 0.0075754f $X=1.485 $Y=0.74 $X2=0 $Y2=0
cc_222 N_C1_M1039_g N_VGND_c_1097_n 0.00762539f $X=1.915 $Y=0.74 $X2=0 $Y2=0
cc_223 N_C1_M1015_g N_VGND_c_1098_n 0.00383152f $X=0.625 $Y=0.74 $X2=0 $Y2=0
cc_224 N_A2_M1019_g N_A1_M1012_g 0.0207253f $X=4.3 $Y=0.74 $X2=0 $Y2=0
cc_225 N_A2_c_244_n N_A1_c_325_n 0.0258812f $X=4.355 $Y=1.765 $X2=0 $Y2=0
cc_226 N_A2_c_239_n A1 0.0297641f $X=4.1 $Y=1.515 $X2=0 $Y2=0
cc_227 N_A2_c_240_n A1 0.00334761f $X=4.3 $Y=1.557 $X2=0 $Y2=0
cc_228 N_A2_c_239_n N_A1_c_324_n 2.30583e-19 $X=4.1 $Y=1.515 $X2=0 $Y2=0
cc_229 N_A2_c_240_n N_A1_c_324_n 0.023069f $X=4.3 $Y=1.557 $X2=0 $Y2=0
cc_230 N_A2_c_241_n N_Y_c_601_n 0.00250071f $X=3.005 $Y=1.765 $X2=0 $Y2=0
cc_231 N_A2_c_241_n N_Y_c_602_n 0.00134372f $X=3.005 $Y=1.765 $X2=0 $Y2=0
cc_232 N_A2_M1004_g N_Y_c_585_n 0.00247408f $X=3.01 $Y=0.74 $X2=0 $Y2=0
cc_233 N_A2_M1004_g N_Y_c_586_n 0.0125331f $X=3.01 $Y=0.74 $X2=0 $Y2=0
cc_234 N_A2_M1007_g N_Y_c_586_n 0.0104926f $X=3.44 $Y=0.74 $X2=0 $Y2=0
cc_235 N_A2_M1018_g N_Y_c_586_n 0.0104926f $X=3.87 $Y=0.74 $X2=0 $Y2=0
cc_236 N_A2_M1019_g N_Y_c_586_n 0.0137692f $X=4.3 $Y=0.74 $X2=0 $Y2=0
cc_237 N_A2_c_239_n N_Y_c_586_n 0.149442f $X=4.1 $Y=1.515 $X2=0 $Y2=0
cc_238 N_A2_c_240_n N_Y_c_586_n 0.0102156f $X=4.3 $Y=1.557 $X2=0 $Y2=0
cc_239 N_A2_M1004_g N_Y_c_589_n 0.00202289f $X=3.01 $Y=0.74 $X2=0 $Y2=0
cc_240 N_A2_c_239_n N_Y_c_589_n 0.0222088f $X=4.1 $Y=1.515 $X2=0 $Y2=0
cc_241 N_A2_c_241_n N_A_114_368#_c_744_n 0.0126525f $X=3.005 $Y=1.765 $X2=0
+ $Y2=0
cc_242 N_A2_c_242_n N_A_114_368#_c_744_n 0.0107319f $X=3.455 $Y=1.765 $X2=0
+ $Y2=0
cc_243 N_A2_c_243_n N_A_114_368#_c_744_n 0.0107319f $X=3.905 $Y=1.765 $X2=0
+ $Y2=0
cc_244 N_A2_c_244_n N_A_114_368#_c_744_n 0.0151242f $X=4.355 $Y=1.765 $X2=0
+ $Y2=0
cc_245 N_A2_c_239_n N_A_114_368#_c_744_n 0.157589f $X=4.1 $Y=1.515 $X2=0 $Y2=0
cc_246 N_A2_c_240_n N_A_114_368#_c_744_n 0.00392578f $X=4.3 $Y=1.557 $X2=0 $Y2=0
cc_247 N_A2_c_241_n N_A_531_368#_c_863_n 0.011796f $X=3.005 $Y=1.765 $X2=0 $Y2=0
cc_248 N_A2_c_242_n N_A_531_368#_c_863_n 0.011796f $X=3.455 $Y=1.765 $X2=0 $Y2=0
cc_249 N_A2_c_243_n N_A_531_368#_c_865_n 0.011796f $X=3.905 $Y=1.765 $X2=0 $Y2=0
cc_250 N_A2_c_244_n N_A_531_368#_c_865_n 0.011796f $X=4.355 $Y=1.765 $X2=0 $Y2=0
cc_251 N_A2_c_241_n N_A_531_368#_c_855_n 0.0079623f $X=3.005 $Y=1.765 $X2=0
+ $Y2=0
cc_252 N_A2_c_242_n N_A_531_368#_c_855_n 5.64076e-19 $X=3.455 $Y=1.765 $X2=0
+ $Y2=0
cc_253 N_A2_c_241_n N_A_531_368#_c_856_n 5.64076e-19 $X=3.005 $Y=1.765 $X2=0
+ $Y2=0
cc_254 N_A2_c_242_n N_A_531_368#_c_856_n 0.00762432f $X=3.455 $Y=1.765 $X2=0
+ $Y2=0
cc_255 N_A2_c_243_n N_A_531_368#_c_856_n 0.00762432f $X=3.905 $Y=1.765 $X2=0
+ $Y2=0
cc_256 N_A2_c_244_n N_A_531_368#_c_856_n 5.64076e-19 $X=4.355 $Y=1.765 $X2=0
+ $Y2=0
cc_257 N_A2_c_243_n N_A_531_368#_c_857_n 5.64076e-19 $X=3.905 $Y=1.765 $X2=0
+ $Y2=0
cc_258 N_A2_c_244_n N_A_531_368#_c_857_n 0.00761095f $X=4.355 $Y=1.765 $X2=0
+ $Y2=0
cc_259 N_A2_c_241_n N_VPWR_c_971_n 0.00379374f $X=3.005 $Y=1.765 $X2=0 $Y2=0
cc_260 N_A2_c_242_n N_VPWR_c_971_n 0.00379374f $X=3.455 $Y=1.765 $X2=0 $Y2=0
cc_261 N_A2_c_242_n N_VPWR_c_972_n 0.00445602f $X=3.455 $Y=1.765 $X2=0 $Y2=0
cc_262 N_A2_c_243_n N_VPWR_c_972_n 0.00445602f $X=3.905 $Y=1.765 $X2=0 $Y2=0
cc_263 N_A2_c_243_n N_VPWR_c_973_n 0.00379374f $X=3.905 $Y=1.765 $X2=0 $Y2=0
cc_264 N_A2_c_244_n N_VPWR_c_973_n 0.00379374f $X=4.355 $Y=1.765 $X2=0 $Y2=0
cc_265 N_A2_c_241_n N_VPWR_c_976_n 0.00445602f $X=3.005 $Y=1.765 $X2=0 $Y2=0
cc_266 N_A2_c_244_n N_VPWR_c_978_n 0.00445602f $X=4.355 $Y=1.765 $X2=0 $Y2=0
cc_267 N_A2_c_241_n N_VPWR_c_970_n 0.00862391f $X=3.005 $Y=1.765 $X2=0 $Y2=0
cc_268 N_A2_c_242_n N_VPWR_c_970_n 0.00857589f $X=3.455 $Y=1.765 $X2=0 $Y2=0
cc_269 N_A2_c_243_n N_VPWR_c_970_n 0.00857589f $X=3.905 $Y=1.765 $X2=0 $Y2=0
cc_270 N_A2_c_244_n N_VPWR_c_970_n 0.00857673f $X=4.355 $Y=1.765 $X2=0 $Y2=0
cc_271 N_A2_M1004_g N_VGND_c_1087_n 0.0095457f $X=3.01 $Y=0.74 $X2=0 $Y2=0
cc_272 N_A2_M1007_g N_VGND_c_1087_n 0.0066521f $X=3.44 $Y=0.74 $X2=0 $Y2=0
cc_273 N_A2_M1018_g N_VGND_c_1087_n 3.94048e-19 $X=3.87 $Y=0.74 $X2=0 $Y2=0
cc_274 N_A2_M1007_g N_VGND_c_1088_n 3.94048e-19 $X=3.44 $Y=0.74 $X2=0 $Y2=0
cc_275 N_A2_M1018_g N_VGND_c_1088_n 0.0066521f $X=3.87 $Y=0.74 $X2=0 $Y2=0
cc_276 N_A2_M1019_g N_VGND_c_1088_n 0.00637998f $X=4.3 $Y=0.74 $X2=0 $Y2=0
cc_277 N_A2_M1004_g N_VGND_c_1092_n 0.00281141f $X=3.01 $Y=0.74 $X2=0 $Y2=0
cc_278 N_A2_M1007_g N_VGND_c_1093_n 0.00281141f $X=3.44 $Y=0.74 $X2=0 $Y2=0
cc_279 N_A2_M1018_g N_VGND_c_1093_n 0.00281141f $X=3.87 $Y=0.74 $X2=0 $Y2=0
cc_280 N_A2_M1019_g N_VGND_c_1094_n 0.00281141f $X=4.3 $Y=0.74 $X2=0 $Y2=0
cc_281 N_A2_M1004_g N_VGND_c_1097_n 0.00370065f $X=3.01 $Y=0.74 $X2=0 $Y2=0
cc_282 N_A2_M1007_g N_VGND_c_1097_n 0.00365066f $X=3.44 $Y=0.74 $X2=0 $Y2=0
cc_283 N_A2_M1018_g N_VGND_c_1097_n 0.00365066f $X=3.87 $Y=0.74 $X2=0 $Y2=0
cc_284 N_A2_M1019_g N_VGND_c_1097_n 0.00365164f $X=4.3 $Y=0.74 $X2=0 $Y2=0
cc_285 N_A2_M1004_g N_A_534_74#_c_1225_n 0.00178474f $X=3.01 $Y=0.74 $X2=0 $Y2=0
cc_286 N_A2_M1004_g N_A_534_74#_c_1234_n 0.011651f $X=3.01 $Y=0.74 $X2=0 $Y2=0
cc_287 N_A2_M1007_g N_A_534_74#_c_1234_n 0.010916f $X=3.44 $Y=0.74 $X2=0 $Y2=0
cc_288 N_A2_M1007_g N_A_534_74#_c_1227_n 4.34399e-19 $X=3.44 $Y=0.74 $X2=0 $Y2=0
cc_289 N_A2_M1018_g N_A_534_74#_c_1227_n 4.34399e-19 $X=3.87 $Y=0.74 $X2=0 $Y2=0
cc_290 N_A2_M1018_g N_A_534_74#_c_1238_n 0.010916f $X=3.87 $Y=0.74 $X2=0 $Y2=0
cc_291 N_A2_M1019_g N_A_534_74#_c_1238_n 0.00983086f $X=4.3 $Y=0.74 $X2=0 $Y2=0
cc_292 N_A2_M1019_g N_A_534_74#_c_1229_n 5.7591e-19 $X=4.3 $Y=0.74 $X2=0 $Y2=0
cc_293 N_A1_c_328_n N_B1_c_424_n 0.0270824f $X=6.385 $Y=1.765 $X2=-0.19
+ $Y2=-0.245
cc_294 N_A1_c_324_n N_B1_M1011_g 0.00117899f $X=6.02 $Y=1.542 $X2=0 $Y2=0
cc_295 N_A1_c_324_n N_B1_c_421_n 0.0199411f $X=6.02 $Y=1.542 $X2=0 $Y2=0
cc_296 N_A1_c_324_n N_B1_c_422_n 0.00205551f $X=6.02 $Y=1.542 $X2=0 $Y2=0
cc_297 N_A1_c_328_n N_B1_c_423_n 0.00172528f $X=6.385 $Y=1.765 $X2=0 $Y2=0
cc_298 A1 N_B1_c_423_n 0.0218713f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_299 N_A1_c_324_n N_B1_c_423_n 0.0139002f $X=6.02 $Y=1.542 $X2=0 $Y2=0
cc_300 N_A1_M1012_g N_Y_c_586_n 0.012204f $X=4.73 $Y=0.74 $X2=0 $Y2=0
cc_301 A1 N_Y_c_586_n 0.0308513f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_302 N_A1_M1024_g N_Y_c_587_n 0.0122369f $X=5.16 $Y=0.74 $X2=0 $Y2=0
cc_303 N_A1_M1033_g N_Y_c_587_n 0.0122369f $X=5.59 $Y=0.74 $X2=0 $Y2=0
cc_304 A1 N_Y_c_587_n 0.0493873f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_305 N_A1_c_324_n N_Y_c_587_n 0.00263824f $X=6.02 $Y=1.542 $X2=0 $Y2=0
cc_306 A1 N_Y_c_590_n 0.0159678f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_307 N_A1_c_324_n N_Y_c_590_n 0.00269777f $X=6.02 $Y=1.542 $X2=0 $Y2=0
cc_308 A1 N_Y_c_591_n 0.0159678f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_309 N_A1_c_324_n N_Y_c_591_n 0.00284055f $X=6.02 $Y=1.542 $X2=0 $Y2=0
cc_310 N_A1_M1034_g N_Y_c_592_n 0.0143078f $X=6.02 $Y=0.74 $X2=0 $Y2=0
cc_311 A1 N_Y_c_592_n 0.0156329f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_312 N_A1_c_324_n N_Y_c_592_n 0.014872f $X=6.02 $Y=1.542 $X2=0 $Y2=0
cc_313 N_A1_M1034_g N_Y_c_593_n 0.00512693f $X=6.02 $Y=0.74 $X2=0 $Y2=0
cc_314 N_A1_c_325_n N_A_114_368#_c_744_n 0.0106809f $X=4.805 $Y=1.765 $X2=0
+ $Y2=0
cc_315 N_A1_c_326_n N_A_114_368#_c_744_n 0.0107319f $X=5.255 $Y=1.765 $X2=0
+ $Y2=0
cc_316 N_A1_c_327_n N_A_114_368#_c_744_n 0.011734f $X=5.705 $Y=1.765 $X2=0 $Y2=0
cc_317 N_A1_c_328_n N_A_114_368#_c_744_n 0.013276f $X=6.385 $Y=1.765 $X2=0 $Y2=0
cc_318 A1 N_A_114_368#_c_744_n 0.113897f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_319 N_A1_c_324_n N_A_114_368#_c_744_n 0.0103625f $X=6.02 $Y=1.542 $X2=0 $Y2=0
cc_320 N_A1_c_328_n N_A_114_368#_c_770_n 7.3898e-19 $X=6.385 $Y=1.765 $X2=0
+ $Y2=0
cc_321 N_A1_c_325_n N_A_531_368#_c_875_n 0.011796f $X=4.805 $Y=1.765 $X2=0 $Y2=0
cc_322 N_A1_c_326_n N_A_531_368#_c_875_n 0.011796f $X=5.255 $Y=1.765 $X2=0 $Y2=0
cc_323 N_A1_c_327_n N_A_531_368#_c_877_n 0.0127981f $X=5.705 $Y=1.765 $X2=0
+ $Y2=0
cc_324 N_A1_c_328_n N_A_531_368#_c_877_n 0.0127981f $X=6.385 $Y=1.765 $X2=0
+ $Y2=0
cc_325 N_A1_c_328_n N_A_531_368#_c_879_n 4.27055e-19 $X=6.385 $Y=1.765 $X2=0
+ $Y2=0
cc_326 N_A1_c_327_n N_A_531_368#_c_880_n 7.59588e-19 $X=5.705 $Y=1.765 $X2=0
+ $Y2=0
cc_327 N_A1_c_328_n N_A_531_368#_c_880_n 0.00620238f $X=6.385 $Y=1.765 $X2=0
+ $Y2=0
cc_328 N_A1_c_328_n N_A_531_368#_c_850_n 0.00315682f $X=6.385 $Y=1.765 $X2=0
+ $Y2=0
cc_329 N_A1_c_325_n N_A_531_368#_c_857_n 0.00761095f $X=4.805 $Y=1.765 $X2=0
+ $Y2=0
cc_330 N_A1_c_326_n N_A_531_368#_c_857_n 5.64076e-19 $X=5.255 $Y=1.765 $X2=0
+ $Y2=0
cc_331 N_A1_c_325_n N_A_531_368#_c_858_n 5.64076e-19 $X=4.805 $Y=1.765 $X2=0
+ $Y2=0
cc_332 N_A1_c_326_n N_A_531_368#_c_858_n 0.00762432f $X=5.255 $Y=1.765 $X2=0
+ $Y2=0
cc_333 N_A1_c_327_n N_A_531_368#_c_858_n 0.00811901f $X=5.705 $Y=1.765 $X2=0
+ $Y2=0
cc_334 N_A1_c_328_n N_A_531_368#_c_858_n 7.69726e-19 $X=6.385 $Y=1.765 $X2=0
+ $Y2=0
cc_335 N_A1_c_325_n N_VPWR_c_974_n 0.00379374f $X=4.805 $Y=1.765 $X2=0 $Y2=0
cc_336 N_A1_c_326_n N_VPWR_c_974_n 0.00379374f $X=5.255 $Y=1.765 $X2=0 $Y2=0
cc_337 N_A1_c_327_n N_VPWR_c_975_n 0.00624962f $X=5.705 $Y=1.765 $X2=0 $Y2=0
cc_338 N_A1_c_328_n N_VPWR_c_975_n 0.00419392f $X=6.385 $Y=1.765 $X2=0 $Y2=0
cc_339 N_A1_c_325_n N_VPWR_c_978_n 0.00445602f $X=4.805 $Y=1.765 $X2=0 $Y2=0
cc_340 N_A1_c_326_n N_VPWR_c_980_n 0.00445602f $X=5.255 $Y=1.765 $X2=0 $Y2=0
cc_341 N_A1_c_327_n N_VPWR_c_980_n 0.00445602f $X=5.705 $Y=1.765 $X2=0 $Y2=0
cc_342 N_A1_c_328_n N_VPWR_c_981_n 0.0044313f $X=6.385 $Y=1.765 $X2=0 $Y2=0
cc_343 N_A1_c_325_n N_VPWR_c_970_n 0.00857673f $X=4.805 $Y=1.765 $X2=0 $Y2=0
cc_344 N_A1_c_326_n N_VPWR_c_970_n 0.00857589f $X=5.255 $Y=1.765 $X2=0 $Y2=0
cc_345 N_A1_c_327_n N_VPWR_c_970_n 0.00858715f $X=5.705 $Y=1.765 $X2=0 $Y2=0
cc_346 N_A1_c_328_n N_VPWR_c_970_n 0.0085457f $X=6.385 $Y=1.765 $X2=0 $Y2=0
cc_347 N_A1_M1012_g N_VGND_c_1088_n 4.21834e-19 $X=4.73 $Y=0.74 $X2=0 $Y2=0
cc_348 N_A1_M1012_g N_VGND_c_1094_n 0.00284711f $X=4.73 $Y=0.74 $X2=0 $Y2=0
cc_349 N_A1_M1024_g N_VGND_c_1094_n 0.00284711f $X=5.16 $Y=0.74 $X2=0 $Y2=0
cc_350 N_A1_M1033_g N_VGND_c_1094_n 0.00284711f $X=5.59 $Y=0.74 $X2=0 $Y2=0
cc_351 N_A1_M1034_g N_VGND_c_1094_n 0.0028589f $X=6.02 $Y=0.74 $X2=0 $Y2=0
cc_352 N_A1_M1012_g N_VGND_c_1097_n 0.00355092f $X=4.73 $Y=0.74 $X2=0 $Y2=0
cc_353 N_A1_M1024_g N_VGND_c_1097_n 0.00354995f $X=5.16 $Y=0.74 $X2=0 $Y2=0
cc_354 N_A1_M1033_g N_VGND_c_1097_n 0.00354995f $X=5.59 $Y=0.74 $X2=0 $Y2=0
cc_355 N_A1_M1034_g N_VGND_c_1097_n 0.00359075f $X=6.02 $Y=0.74 $X2=0 $Y2=0
cc_356 N_A1_M1012_g N_A_534_74#_c_1241_n 0.00207208f $X=4.73 $Y=0.74 $X2=0 $Y2=0
cc_357 N_A1_M1012_g N_A_534_74#_c_1242_n 0.00405013f $X=4.73 $Y=0.74 $X2=0 $Y2=0
cc_358 N_A1_M1024_g N_A_534_74#_c_1242_n 4.66834e-19 $X=5.16 $Y=0.74 $X2=0 $Y2=0
cc_359 N_A1_M1012_g N_A_534_74#_c_1228_n 0.00832673f $X=4.73 $Y=0.74 $X2=0 $Y2=0
cc_360 N_A1_M1024_g N_A_534_74#_c_1228_n 0.00828016f $X=5.16 $Y=0.74 $X2=0 $Y2=0
cc_361 N_A1_M1012_g N_A_534_74#_c_1229_n 0.0012003f $X=4.73 $Y=0.74 $X2=0 $Y2=0
cc_362 N_A1_M1012_g N_A_534_74#_c_1247_n 5.14064e-19 $X=4.73 $Y=0.74 $X2=0 $Y2=0
cc_363 N_A1_M1024_g N_A_534_74#_c_1247_n 0.00611013f $X=5.16 $Y=0.74 $X2=0 $Y2=0
cc_364 N_A1_M1033_g N_A_534_74#_c_1247_n 0.00611013f $X=5.59 $Y=0.74 $X2=0 $Y2=0
cc_365 N_A1_M1034_g N_A_534_74#_c_1247_n 5.14064e-19 $X=6.02 $Y=0.74 $X2=0 $Y2=0
cc_366 N_A1_M1033_g N_A_534_74#_c_1230_n 0.00832673f $X=5.59 $Y=0.74 $X2=0 $Y2=0
cc_367 N_A1_M1034_g N_A_534_74#_c_1230_n 0.00890733f $X=6.02 $Y=0.74 $X2=0 $Y2=0
cc_368 N_A1_M1024_g N_A_534_74#_c_1231_n 0.001391f $X=5.16 $Y=0.74 $X2=0 $Y2=0
cc_369 N_A1_M1033_g N_A_534_74#_c_1231_n 0.001391f $X=5.59 $Y=0.74 $X2=0 $Y2=0
cc_370 N_A1_M1033_g N_A_534_74#_c_1232_n 5.28405e-19 $X=5.59 $Y=0.74 $X2=0 $Y2=0
cc_371 N_A1_M1034_g N_A_534_74#_c_1232_n 0.00635002f $X=6.02 $Y=0.74 $X2=0 $Y2=0
cc_372 N_A1_M1034_g N_A_1326_74#_c_1318_n 6.29126e-19 $X=6.02 $Y=0.74 $X2=0
+ $Y2=0
cc_373 N_B1_c_427_n N_B2_c_511_n 0.0263546f $X=8.185 $Y=1.765 $X2=-0.19
+ $Y2=-0.245
cc_374 N_B1_M1036_g N_B2_M1006_g 0.019323f $X=8.26 $Y=0.74 $X2=0 $Y2=0
cc_375 N_B1_c_428_n B2 0.0344451f $X=7.93 $Y=1.515 $X2=0 $Y2=0
cc_376 N_B1_c_421_n B2 0.0105978f $X=8.185 $Y=1.557 $X2=0 $Y2=0
cc_377 N_B1_c_428_n N_B2_c_510_n 2.57635e-19 $X=7.93 $Y=1.515 $X2=0 $Y2=0
cc_378 N_B1_c_421_n N_B2_c_510_n 0.0219308f $X=8.185 $Y=1.557 $X2=0 $Y2=0
cc_379 N_B1_M1011_g N_Y_c_593_n 0.00263991f $X=6.97 $Y=0.74 $X2=0 $Y2=0
cc_380 N_B1_c_423_n N_Y_c_593_n 0.0135709f $X=6.73 $Y=1.565 $X2=0 $Y2=0
cc_381 N_B1_M1036_g N_Y_c_594_n 0.00660558f $X=8.26 $Y=0.74 $X2=0 $Y2=0
cc_382 N_B1_c_428_n N_Y_c_594_n 0.0542704f $X=7.93 $Y=1.515 $X2=0 $Y2=0
cc_383 N_B1_c_421_n N_Y_c_594_n 0.00229127f $X=8.185 $Y=1.557 $X2=0 $Y2=0
cc_384 N_B1_M1011_g N_Y_c_595_n 0.0176197f $X=6.97 $Y=0.74 $X2=0 $Y2=0
cc_385 N_B1_M1014_g N_Y_c_595_n 0.0139412f $X=7.4 $Y=0.74 $X2=0 $Y2=0
cc_386 N_B1_M1028_g N_Y_c_595_n 0.014021f $X=7.83 $Y=0.74 $X2=0 $Y2=0
cc_387 N_B1_c_421_n N_Y_c_595_n 0.00867274f $X=8.185 $Y=1.557 $X2=0 $Y2=0
cc_388 N_B1_c_422_n N_Y_c_595_n 0.0542704f $X=6.945 $Y=1.565 $X2=0 $Y2=0
cc_389 N_B1_c_423_n N_Y_c_595_n 0.0127232f $X=6.73 $Y=1.565 $X2=0 $Y2=0
cc_390 N_B1_c_424_n N_A_114_368#_c_744_n 0.0119563f $X=6.835 $Y=1.765 $X2=0
+ $Y2=0
cc_391 N_B1_c_423_n N_A_114_368#_c_744_n 0.0359874f $X=6.73 $Y=1.565 $X2=0 $Y2=0
cc_392 N_B1_c_425_n N_A_114_368#_c_773_n 0.0120074f $X=7.285 $Y=1.765 $X2=0
+ $Y2=0
cc_393 N_B1_c_426_n N_A_114_368#_c_773_n 0.0120074f $X=7.735 $Y=1.765 $X2=0
+ $Y2=0
cc_394 N_B1_c_428_n N_A_114_368#_c_773_n 0.0393875f $X=7.93 $Y=1.515 $X2=0 $Y2=0
cc_395 N_B1_c_421_n N_A_114_368#_c_773_n 0.00130718f $X=8.185 $Y=1.557 $X2=0
+ $Y2=0
cc_396 N_B1_c_427_n N_A_114_368#_c_777_n 0.0160489f $X=8.185 $Y=1.765 $X2=0
+ $Y2=0
cc_397 N_B1_c_424_n N_A_114_368#_c_770_n 0.0103124f $X=6.835 $Y=1.765 $X2=0
+ $Y2=0
cc_398 N_B1_c_425_n N_A_114_368#_c_770_n 0.010266f $X=7.285 $Y=1.765 $X2=0 $Y2=0
cc_399 N_B1_c_426_n N_A_114_368#_c_770_n 5.52094e-19 $X=7.735 $Y=1.765 $X2=0
+ $Y2=0
cc_400 N_B1_c_421_n N_A_114_368#_c_770_n 0.00145694f $X=8.185 $Y=1.557 $X2=0
+ $Y2=0
cc_401 N_B1_c_422_n N_A_114_368#_c_770_n 0.0237163f $X=6.945 $Y=1.565 $X2=0
+ $Y2=0
cc_402 N_B1_c_425_n N_A_114_368#_c_783_n 5.52094e-19 $X=7.285 $Y=1.765 $X2=0
+ $Y2=0
cc_403 N_B1_c_426_n N_A_114_368#_c_783_n 0.010266f $X=7.735 $Y=1.765 $X2=0 $Y2=0
cc_404 N_B1_c_427_n N_A_114_368#_c_783_n 0.0107899f $X=8.185 $Y=1.765 $X2=0
+ $Y2=0
cc_405 N_B1_c_428_n N_A_114_368#_c_783_n 0.0219285f $X=7.93 $Y=1.515 $X2=0 $Y2=0
cc_406 N_B1_c_421_n N_A_114_368#_c_783_n 0.00144162f $X=8.185 $Y=1.557 $X2=0
+ $Y2=0
cc_407 N_B1_c_427_n N_A_114_368#_c_788_n 5.52094e-19 $X=8.185 $Y=1.765 $X2=0
+ $Y2=0
cc_408 N_B1_c_424_n N_A_531_368#_c_849_n 0.0128006f $X=6.835 $Y=1.765 $X2=0
+ $Y2=0
cc_409 N_B1_c_425_n N_A_531_368#_c_849_n 0.0128349f $X=7.285 $Y=1.765 $X2=0
+ $Y2=0
cc_410 N_B1_c_426_n N_A_531_368#_c_851_n 0.0128349f $X=7.735 $Y=1.765 $X2=0
+ $Y2=0
cc_411 N_B1_c_427_n N_A_531_368#_c_851_n 0.0128006f $X=8.185 $Y=1.765 $X2=0
+ $Y2=0
cc_412 N_B1_c_424_n N_VPWR_c_981_n 0.00278271f $X=6.835 $Y=1.765 $X2=0 $Y2=0
cc_413 N_B1_c_425_n N_VPWR_c_981_n 0.00278271f $X=7.285 $Y=1.765 $X2=0 $Y2=0
cc_414 N_B1_c_426_n N_VPWR_c_981_n 0.00278271f $X=7.735 $Y=1.765 $X2=0 $Y2=0
cc_415 N_B1_c_427_n N_VPWR_c_981_n 0.00278271f $X=8.185 $Y=1.765 $X2=0 $Y2=0
cc_416 N_B1_c_424_n N_VPWR_c_970_n 0.00353907f $X=6.835 $Y=1.765 $X2=0 $Y2=0
cc_417 N_B1_c_425_n N_VPWR_c_970_n 0.00353823f $X=7.285 $Y=1.765 $X2=0 $Y2=0
cc_418 N_B1_c_426_n N_VPWR_c_970_n 0.00353823f $X=7.735 $Y=1.765 $X2=0 $Y2=0
cc_419 N_B1_c_427_n N_VPWR_c_970_n 0.00353907f $X=8.185 $Y=1.765 $X2=0 $Y2=0
cc_420 N_B1_M1036_g N_VGND_c_1089_n 6.35276e-19 $X=8.26 $Y=0.74 $X2=0 $Y2=0
cc_421 N_B1_M1011_g N_VGND_c_1094_n 0.00291649f $X=6.97 $Y=0.74 $X2=0 $Y2=0
cc_422 N_B1_M1014_g N_VGND_c_1094_n 0.00291649f $X=7.4 $Y=0.74 $X2=0 $Y2=0
cc_423 N_B1_M1028_g N_VGND_c_1094_n 0.00291649f $X=7.83 $Y=0.74 $X2=0 $Y2=0
cc_424 N_B1_M1036_g N_VGND_c_1094_n 0.00291649f $X=8.26 $Y=0.74 $X2=0 $Y2=0
cc_425 N_B1_M1011_g N_VGND_c_1097_n 0.0036412f $X=6.97 $Y=0.74 $X2=0 $Y2=0
cc_426 N_B1_M1014_g N_VGND_c_1097_n 0.00359121f $X=7.4 $Y=0.74 $X2=0 $Y2=0
cc_427 N_B1_M1028_g N_VGND_c_1097_n 0.00359121f $X=7.83 $Y=0.74 $X2=0 $Y2=0
cc_428 N_B1_M1036_g N_VGND_c_1097_n 0.00359219f $X=8.26 $Y=0.74 $X2=0 $Y2=0
cc_429 N_B1_M1011_g N_A_534_74#_c_1232_n 0.00189749f $X=6.97 $Y=0.74 $X2=0 $Y2=0
cc_430 N_B1_M1028_g N_A_1326_74#_c_1311_n 0.0106239f $X=7.83 $Y=0.74 $X2=0 $Y2=0
cc_431 N_B1_M1036_g N_A_1326_74#_c_1311_n 0.014175f $X=8.26 $Y=0.74 $X2=0 $Y2=0
cc_432 N_B1_M1036_g N_A_1326_74#_c_1314_n 5.97859e-19 $X=8.26 $Y=0.74 $X2=0
+ $Y2=0
cc_433 N_B1_M1011_g N_A_1326_74#_c_1318_n 0.00289501f $X=6.97 $Y=0.74 $X2=0
+ $Y2=0
cc_434 N_B1_M1014_g N_A_1326_74#_c_1318_n 2.3282e-19 $X=7.4 $Y=0.74 $X2=0 $Y2=0
cc_435 N_B1_M1011_g N_A_1326_74#_c_1319_n 0.00920696f $X=6.97 $Y=0.74 $X2=0
+ $Y2=0
cc_436 N_B1_M1014_g N_A_1326_74#_c_1319_n 0.00920696f $X=7.4 $Y=0.74 $X2=0 $Y2=0
cc_437 N_B1_M1011_g N_A_1326_74#_c_1320_n 2.32994e-19 $X=6.97 $Y=0.74 $X2=0
+ $Y2=0
cc_438 N_B1_M1014_g N_A_1326_74#_c_1320_n 0.00274634f $X=7.4 $Y=0.74 $X2=0 $Y2=0
cc_439 N_B2_c_511_n N_A_114_368#_c_777_n 0.0119563f $X=8.635 $Y=1.765 $X2=0
+ $Y2=0
cc_440 B2 N_A_114_368#_c_777_n 0.0284881f $X=9.755 $Y=1.58 $X2=0 $Y2=0
cc_441 N_B2_c_512_n N_A_114_368#_c_791_n 0.0120074f $X=9.085 $Y=1.765 $X2=0
+ $Y2=0
cc_442 N_B2_c_513_n N_A_114_368#_c_791_n 0.0120074f $X=9.535 $Y=1.765 $X2=0
+ $Y2=0
cc_443 B2 N_A_114_368#_c_791_n 0.0393875f $X=9.755 $Y=1.58 $X2=0 $Y2=0
cc_444 N_B2_c_510_n N_A_114_368#_c_791_n 0.00130859f $X=9.98 $Y=1.557 $X2=0
+ $Y2=0
cc_445 N_B2_c_511_n N_A_114_368#_c_783_n 5.52094e-19 $X=8.635 $Y=1.765 $X2=0
+ $Y2=0
cc_446 N_B2_c_511_n N_A_114_368#_c_788_n 0.010266f $X=8.635 $Y=1.765 $X2=0 $Y2=0
cc_447 N_B2_c_512_n N_A_114_368#_c_788_n 0.010266f $X=9.085 $Y=1.765 $X2=0 $Y2=0
cc_448 N_B2_c_513_n N_A_114_368#_c_788_n 5.52094e-19 $X=9.535 $Y=1.765 $X2=0
+ $Y2=0
cc_449 B2 N_A_114_368#_c_788_n 0.0237598f $X=9.755 $Y=1.58 $X2=0 $Y2=0
cc_450 N_B2_c_510_n N_A_114_368#_c_788_n 0.00144162f $X=9.98 $Y=1.557 $X2=0
+ $Y2=0
cc_451 N_B2_c_512_n N_A_114_368#_c_801_n 5.52094e-19 $X=9.085 $Y=1.765 $X2=0
+ $Y2=0
cc_452 N_B2_c_513_n N_A_114_368#_c_801_n 0.010266f $X=9.535 $Y=1.765 $X2=0 $Y2=0
cc_453 N_B2_c_514_n N_A_114_368#_c_801_n 0.0113048f $X=9.985 $Y=1.765 $X2=0
+ $Y2=0
cc_454 B2 N_A_114_368#_c_801_n 0.0237598f $X=9.755 $Y=1.58 $X2=0 $Y2=0
cc_455 N_B2_c_510_n N_A_114_368#_c_801_n 0.00144162f $X=9.98 $Y=1.557 $X2=0
+ $Y2=0
cc_456 N_B2_c_511_n N_A_531_368#_c_852_n 0.0128006f $X=8.635 $Y=1.765 $X2=0
+ $Y2=0
cc_457 N_B2_c_512_n N_A_531_368#_c_852_n 0.0128349f $X=9.085 $Y=1.765 $X2=0
+ $Y2=0
cc_458 N_B2_c_513_n N_A_531_368#_c_853_n 0.0128349f $X=9.535 $Y=1.765 $X2=0
+ $Y2=0
cc_459 N_B2_c_514_n N_A_531_368#_c_853_n 0.0137046f $X=9.985 $Y=1.765 $X2=0
+ $Y2=0
cc_460 N_B2_c_514_n N_A_531_368#_c_854_n 0.010383f $X=9.985 $Y=1.765 $X2=0 $Y2=0
cc_461 N_B2_c_511_n N_VPWR_c_981_n 0.00278271f $X=8.635 $Y=1.765 $X2=0 $Y2=0
cc_462 N_B2_c_512_n N_VPWR_c_981_n 0.00278271f $X=9.085 $Y=1.765 $X2=0 $Y2=0
cc_463 N_B2_c_513_n N_VPWR_c_981_n 0.00278271f $X=9.535 $Y=1.765 $X2=0 $Y2=0
cc_464 N_B2_c_514_n N_VPWR_c_981_n 0.00278271f $X=9.985 $Y=1.765 $X2=0 $Y2=0
cc_465 N_B2_c_511_n N_VPWR_c_970_n 0.00353907f $X=8.635 $Y=1.765 $X2=0 $Y2=0
cc_466 N_B2_c_512_n N_VPWR_c_970_n 0.00353823f $X=9.085 $Y=1.765 $X2=0 $Y2=0
cc_467 N_B2_c_513_n N_VPWR_c_970_n 0.00353823f $X=9.535 $Y=1.765 $X2=0 $Y2=0
cc_468 N_B2_c_514_n N_VPWR_c_970_n 0.00357527f $X=9.985 $Y=1.765 $X2=0 $Y2=0
cc_469 N_B2_M1006_g N_VGND_c_1089_n 0.010782f $X=8.69 $Y=0.74 $X2=0 $Y2=0
cc_470 N_B2_M1008_g N_VGND_c_1089_n 0.0106755f $X=9.12 $Y=0.74 $X2=0 $Y2=0
cc_471 N_B2_M1020_g N_VGND_c_1089_n 4.71636e-19 $X=9.55 $Y=0.74 $X2=0 $Y2=0
cc_472 N_B2_M1008_g N_VGND_c_1090_n 4.71636e-19 $X=9.12 $Y=0.74 $X2=0 $Y2=0
cc_473 N_B2_M1020_g N_VGND_c_1090_n 0.0106755f $X=9.55 $Y=0.74 $X2=0 $Y2=0
cc_474 N_B2_M1023_g N_VGND_c_1090_n 0.0137191f $X=9.98 $Y=0.74 $X2=0 $Y2=0
cc_475 N_B2_M1006_g N_VGND_c_1094_n 0.00383152f $X=8.69 $Y=0.74 $X2=0 $Y2=0
cc_476 N_B2_M1008_g N_VGND_c_1095_n 0.00383152f $X=9.12 $Y=0.74 $X2=0 $Y2=0
cc_477 N_B2_M1020_g N_VGND_c_1095_n 0.00383152f $X=9.55 $Y=0.74 $X2=0 $Y2=0
cc_478 N_B2_M1023_g N_VGND_c_1096_n 0.00383152f $X=9.98 $Y=0.74 $X2=0 $Y2=0
cc_479 N_B2_M1006_g N_VGND_c_1097_n 0.00757637f $X=8.69 $Y=0.74 $X2=0 $Y2=0
cc_480 N_B2_M1008_g N_VGND_c_1097_n 0.0075754f $X=9.12 $Y=0.74 $X2=0 $Y2=0
cc_481 N_B2_M1020_g N_VGND_c_1097_n 0.0075754f $X=9.55 $Y=0.74 $X2=0 $Y2=0
cc_482 N_B2_M1023_g N_VGND_c_1097_n 0.00761455f $X=9.98 $Y=0.74 $X2=0 $Y2=0
cc_483 N_B2_M1006_g N_A_1326_74#_c_1313_n 0.0128967f $X=8.69 $Y=0.74 $X2=0 $Y2=0
cc_484 N_B2_M1008_g N_A_1326_74#_c_1313_n 0.0130453f $X=9.12 $Y=0.74 $X2=0 $Y2=0
cc_485 B2 N_A_1326_74#_c_1313_n 0.0517333f $X=9.755 $Y=1.58 $X2=0 $Y2=0
cc_486 N_B2_c_510_n N_A_1326_74#_c_1313_n 0.00368969f $X=9.98 $Y=1.557 $X2=0
+ $Y2=0
cc_487 B2 N_A_1326_74#_c_1314_n 0.0152645f $X=9.755 $Y=1.58 $X2=0 $Y2=0
cc_488 N_B2_c_510_n N_A_1326_74#_c_1314_n 3.65737e-19 $X=9.98 $Y=1.557 $X2=0
+ $Y2=0
cc_489 N_B2_M1008_g N_A_1326_74#_c_1315_n 3.92313e-19 $X=9.12 $Y=0.74 $X2=0
+ $Y2=0
cc_490 N_B2_M1020_g N_A_1326_74#_c_1315_n 3.92313e-19 $X=9.55 $Y=0.74 $X2=0
+ $Y2=0
cc_491 N_B2_M1020_g N_A_1326_74#_c_1316_n 0.0130918f $X=9.55 $Y=0.74 $X2=0 $Y2=0
cc_492 N_B2_M1023_g N_A_1326_74#_c_1316_n 0.0167076f $X=9.98 $Y=0.74 $X2=0 $Y2=0
cc_493 B2 N_A_1326_74#_c_1316_n 0.0402557f $X=9.755 $Y=1.58 $X2=0 $Y2=0
cc_494 N_B2_c_510_n N_A_1326_74#_c_1316_n 0.00238888f $X=9.98 $Y=1.557 $X2=0
+ $Y2=0
cc_495 N_B2_M1023_g N_A_1326_74#_c_1317_n 0.00159319f $X=9.98 $Y=0.74 $X2=0
+ $Y2=0
cc_496 B2 N_A_1326_74#_c_1321_n 0.0146029f $X=9.755 $Y=1.58 $X2=0 $Y2=0
cc_497 N_B2_c_510_n N_A_1326_74#_c_1321_n 0.00232957f $X=9.98 $Y=1.557 $X2=0
+ $Y2=0
cc_498 N_Y_c_599_n N_A_114_368#_M1002_d 0.00197722f $X=1.005 $Y=2.99 $X2=-0.19
+ $Y2=-0.245
cc_499 N_Y_c_601_n N_A_114_368#_M1005_d 0.00197722f $X=1.905 $Y=2.99 $X2=0 $Y2=0
cc_500 Y N_A_114_368#_c_745_n 0.0121024f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_501 N_Y_c_599_n N_A_114_368#_c_748_n 0.0151173f $X=1.005 $Y=2.99 $X2=0 $Y2=0
cc_502 Y N_A_114_368#_c_748_n 0.0407007f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_503 N_Y_M1003_s N_A_114_368#_c_749_n 0.00359365f $X=1.02 $Y=1.84 $X2=0 $Y2=0
cc_504 N_Y_c_611_n N_A_114_368#_c_749_n 0.0171813f $X=1.17 $Y=2.41 $X2=0 $Y2=0
cc_505 N_Y_c_601_n N_A_114_368#_c_813_n 0.014157f $X=1.905 $Y=2.99 $X2=0 $Y2=0
cc_506 N_Y_M1009_s N_A_114_368#_c_744_n 0.0070945f $X=1.92 $Y=1.84 $X2=0 $Y2=0
cc_507 N_Y_c_602_n N_A_114_368#_c_744_n 0.0220544f $X=2.07 $Y=2.41 $X2=0 $Y2=0
cc_508 N_Y_c_601_n N_A_531_368#_c_855_n 0.00379666f $X=1.905 $Y=2.99 $X2=0 $Y2=0
cc_509 N_Y_c_602_n N_A_531_368#_c_855_n 0.0298129f $X=2.07 $Y=2.41 $X2=0 $Y2=0
cc_510 N_Y_c_599_n N_VPWR_c_976_n 0.0409869f $X=1.005 $Y=2.99 $X2=0 $Y2=0
cc_511 N_Y_c_600_n N_VPWR_c_976_n 0.0178493f $X=0.355 $Y=2.99 $X2=0 $Y2=0
cc_512 N_Y_c_601_n N_VPWR_c_976_n 0.0594839f $X=1.905 $Y=2.99 $X2=0 $Y2=0
cc_513 N_Y_c_603_n N_VPWR_c_976_n 0.0235512f $X=1.17 $Y=2.99 $X2=0 $Y2=0
cc_514 N_Y_c_599_n N_VPWR_c_970_n 0.0231342f $X=1.005 $Y=2.99 $X2=0 $Y2=0
cc_515 N_Y_c_600_n N_VPWR_c_970_n 0.00970886f $X=0.355 $Y=2.99 $X2=0 $Y2=0
cc_516 N_Y_c_601_n N_VPWR_c_970_n 0.0329562f $X=1.905 $Y=2.99 $X2=0 $Y2=0
cc_517 N_Y_c_603_n N_VPWR_c_970_n 0.0126924f $X=1.17 $Y=2.99 $X2=0 $Y2=0
cc_518 N_Y_c_582_n N_VGND_M1015_d 0.00176461f $X=1.185 $Y=1.095 $X2=-0.19
+ $Y2=-0.245
cc_519 N_Y_c_584_n N_VGND_M1027_d 0.00176461f $X=2.045 $Y=1.095 $X2=0 $Y2=0
cc_520 N_Y_c_586_n N_VGND_M1004_d 0.00176891f $X=4.85 $Y=1.175 $X2=0 $Y2=0
cc_521 N_Y_c_586_n N_VGND_M1018_d 0.00176891f $X=4.85 $Y=1.175 $X2=0 $Y2=0
cc_522 N_Y_c_582_n N_VGND_c_1085_n 0.0170777f $X=1.185 $Y=1.095 $X2=0 $Y2=0
cc_523 N_Y_c_583_n N_VGND_c_1085_n 0.0182488f $X=1.27 $Y=0.515 $X2=0 $Y2=0
cc_524 N_Y_c_597_n N_VGND_c_1085_n 0.0183409f $X=0.41 $Y=0.515 $X2=0 $Y2=0
cc_525 N_Y_c_583_n N_VGND_c_1086_n 0.0182488f $X=1.27 $Y=0.515 $X2=0 $Y2=0
cc_526 N_Y_c_584_n N_VGND_c_1086_n 0.0170777f $X=2.045 $Y=1.095 $X2=0 $Y2=0
cc_527 N_Y_c_585_n N_VGND_c_1086_n 0.0182902f $X=2.13 $Y=0.515 $X2=0 $Y2=0
cc_528 N_Y_c_583_n N_VGND_c_1091_n 0.00749631f $X=1.27 $Y=0.515 $X2=0 $Y2=0
cc_529 N_Y_c_585_n N_VGND_c_1092_n 0.011066f $X=2.13 $Y=0.515 $X2=0 $Y2=0
cc_530 N_Y_c_583_n N_VGND_c_1097_n 0.0062048f $X=1.27 $Y=0.515 $X2=0 $Y2=0
cc_531 N_Y_c_585_n N_VGND_c_1097_n 0.00915947f $X=2.13 $Y=0.515 $X2=0 $Y2=0
cc_532 N_Y_c_593_n N_VGND_c_1097_n 0.00945588f $X=6.53 $Y=1.055 $X2=0 $Y2=0
cc_533 N_Y_c_597_n N_VGND_c_1097_n 0.0143301f $X=0.41 $Y=0.515 $X2=0 $Y2=0
cc_534 N_Y_c_597_n N_VGND_c_1098_n 0.0173129f $X=0.41 $Y=0.515 $X2=0 $Y2=0
cc_535 N_Y_c_586_n N_A_534_74#_M1004_s 0.00230047f $X=4.85 $Y=1.175 $X2=-0.19
+ $Y2=-0.245
cc_536 N_Y_c_586_n N_A_534_74#_M1007_s 0.00176461f $X=4.85 $Y=1.175 $X2=0 $Y2=0
cc_537 N_Y_c_586_n N_A_534_74#_M1019_s 0.00176461f $X=4.85 $Y=1.175 $X2=0 $Y2=0
cc_538 N_Y_c_587_n N_A_534_74#_M1024_d 0.00176461f $X=5.71 $Y=1.175 $X2=0 $Y2=0
cc_539 N_Y_c_592_n N_A_534_74#_M1034_d 0.00344852f $X=6.36 $Y=1.055 $X2=0 $Y2=0
cc_540 N_Y_c_593_n N_A_534_74#_M1034_d 0.00287935f $X=6.53 $Y=1.055 $X2=0 $Y2=0
cc_541 N_Y_c_585_n N_A_534_74#_c_1225_n 0.0199479f $X=2.13 $Y=0.515 $X2=0 $Y2=0
cc_542 N_Y_c_586_n N_A_534_74#_c_1234_n 0.0323912f $X=4.85 $Y=1.175 $X2=0 $Y2=0
cc_543 N_Y_c_585_n N_A_534_74#_c_1226_n 0.00920235f $X=2.13 $Y=0.515 $X2=0 $Y2=0
cc_544 N_Y_c_586_n N_A_534_74#_c_1226_n 0.0200122f $X=4.85 $Y=1.175 $X2=0 $Y2=0
cc_545 N_Y_c_586_n N_A_534_74#_c_1238_n 0.0323573f $X=4.85 $Y=1.175 $X2=0 $Y2=0
cc_546 N_Y_c_586_n N_A_534_74#_c_1241_n 0.0152523f $X=4.85 $Y=1.175 $X2=0 $Y2=0
cc_547 N_Y_M1012_s N_A_534_74#_c_1228_n 0.00176461f $X=4.805 $Y=0.37 $X2=0 $Y2=0
cc_548 N_Y_c_586_n N_A_534_74#_c_1228_n 0.00288482f $X=4.85 $Y=1.175 $X2=0 $Y2=0
cc_549 N_Y_c_724_p N_A_534_74#_c_1228_n 0.012662f $X=4.945 $Y=0.805 $X2=0 $Y2=0
cc_550 N_Y_c_587_n N_A_534_74#_c_1228_n 0.00288482f $X=5.71 $Y=1.175 $X2=0 $Y2=0
cc_551 N_Y_c_587_n N_A_534_74#_c_1247_n 0.0169492f $X=5.71 $Y=1.175 $X2=0 $Y2=0
cc_552 N_Y_M1033_s N_A_534_74#_c_1230_n 0.00176461f $X=5.665 $Y=0.37 $X2=0 $Y2=0
cc_553 N_Y_c_587_n N_A_534_74#_c_1230_n 0.00288482f $X=5.71 $Y=1.175 $X2=0 $Y2=0
cc_554 N_Y_c_729_p N_A_534_74#_c_1230_n 0.012662f $X=5.805 $Y=0.805 $X2=0 $Y2=0
cc_555 N_Y_c_592_n N_A_534_74#_c_1230_n 0.0028964f $X=6.36 $Y=1.055 $X2=0 $Y2=0
cc_556 N_Y_c_586_n N_A_534_74#_c_1279_n 0.0133131f $X=4.85 $Y=1.175 $X2=0 $Y2=0
cc_557 N_Y_c_592_n N_A_534_74#_c_1232_n 0.00924091f $X=6.36 $Y=1.055 $X2=0 $Y2=0
cc_558 N_Y_c_593_n N_A_534_74#_c_1232_n 0.00327272f $X=6.53 $Y=1.055 $X2=0 $Y2=0
cc_559 N_Y_c_595_n N_A_1326_74#_M1011_d 0.0034516f $X=7.915 $Y=0.975 $X2=-0.19
+ $Y2=-0.245
cc_560 N_Y_c_595_n N_A_1326_74#_M1014_d 0.00178215f $X=7.915 $Y=0.975 $X2=0
+ $Y2=0
cc_561 N_Y_M1028_s N_A_1326_74#_c_1311_n 0.00179007f $X=7.905 $Y=0.37 $X2=0
+ $Y2=0
cc_562 N_Y_c_594_n N_A_1326_74#_c_1311_n 0.014589f $X=8.045 $Y=0.95 $X2=0 $Y2=0
cc_563 N_Y_c_595_n N_A_1326_74#_c_1311_n 0.00752936f $X=7.915 $Y=0.975 $X2=0
+ $Y2=0
cc_564 N_Y_c_594_n N_A_1326_74#_c_1314_n 0.00988477f $X=8.045 $Y=0.95 $X2=0
+ $Y2=0
cc_565 N_Y_c_595_n N_A_1326_74#_c_1318_n 0.0213291f $X=7.915 $Y=0.975 $X2=0
+ $Y2=0
cc_566 N_Y_M1011_s N_A_1326_74#_c_1319_n 0.00212678f $X=7.045 $Y=0.37 $X2=0
+ $Y2=0
cc_567 N_Y_c_595_n N_A_1326_74#_c_1319_n 0.0217197f $X=7.915 $Y=0.975 $X2=0
+ $Y2=0
cc_568 N_Y_c_595_n N_A_1326_74#_c_1320_n 0.0147899f $X=7.915 $Y=0.975 $X2=0
+ $Y2=0
cc_569 N_A_114_368#_c_744_n N_A_531_368#_M1016_s 0.0055238f $X=6.895 $Y=2.035
+ $X2=-0.19 $Y2=1.66
cc_570 N_A_114_368#_c_744_n N_A_531_368#_M1017_s 0.00359365f $X=6.895 $Y=2.035
+ $X2=0 $Y2=0
cc_571 N_A_114_368#_c_744_n N_A_531_368#_M1025_s 0.00392387f $X=6.895 $Y=2.035
+ $X2=0 $Y2=0
cc_572 N_A_114_368#_c_744_n N_A_531_368#_M1026_s 0.00359365f $X=6.895 $Y=2.035
+ $X2=0 $Y2=0
cc_573 N_A_114_368#_c_744_n N_A_531_368#_M1037_s 0.00395925f $X=6.895 $Y=2.035
+ $X2=0 $Y2=0
cc_574 N_A_114_368#_c_773_n N_A_531_368#_M1031_s 0.00359365f $X=7.795 $Y=2.035
+ $X2=0 $Y2=0
cc_575 N_A_114_368#_c_777_n N_A_531_368#_M1035_s 0.00393511f $X=8.695 $Y=2.035
+ $X2=0 $Y2=0
cc_576 N_A_114_368#_c_791_n N_A_531_368#_M1010_d 0.00359365f $X=9.595 $Y=2.035
+ $X2=0 $Y2=0
cc_577 N_A_114_368#_c_744_n N_A_531_368#_c_863_n 0.0317427f $X=6.895 $Y=2.035
+ $X2=0 $Y2=0
cc_578 N_A_114_368#_c_744_n N_A_531_368#_c_865_n 0.0317427f $X=6.895 $Y=2.035
+ $X2=0 $Y2=0
cc_579 N_A_114_368#_c_744_n N_A_531_368#_c_875_n 0.0317427f $X=6.895 $Y=2.035
+ $X2=0 $Y2=0
cc_580 N_A_114_368#_c_744_n N_A_531_368#_c_877_n 0.0484484f $X=6.895 $Y=2.035
+ $X2=0 $Y2=0
cc_581 N_A_114_368#_c_744_n N_A_531_368#_c_879_n 0.0162332f $X=6.895 $Y=2.035
+ $X2=0 $Y2=0
cc_582 N_A_114_368#_M1030_d N_A_531_368#_c_849_n 0.00197722f $X=6.91 $Y=1.84
+ $X2=0 $Y2=0
cc_583 N_A_114_368#_c_770_n N_A_531_368#_c_849_n 0.0160777f $X=7.06 $Y=2.035
+ $X2=0 $Y2=0
cc_584 N_A_114_368#_c_773_n N_A_531_368#_c_915_n 0.0151327f $X=7.795 $Y=2.035
+ $X2=0 $Y2=0
cc_585 N_A_114_368#_M1032_d N_A_531_368#_c_851_n 0.00197722f $X=7.81 $Y=1.84
+ $X2=0 $Y2=0
cc_586 N_A_114_368#_c_783_n N_A_531_368#_c_851_n 0.0160777f $X=7.96 $Y=2.035
+ $X2=0 $Y2=0
cc_587 N_A_114_368#_c_777_n N_A_531_368#_c_918_n 0.0151327f $X=8.695 $Y=2.035
+ $X2=0 $Y2=0
cc_588 N_A_114_368#_M1001_s N_A_531_368#_c_852_n 0.00197722f $X=8.71 $Y=1.84
+ $X2=0 $Y2=0
cc_589 N_A_114_368#_c_788_n N_A_531_368#_c_852_n 0.0160777f $X=8.86 $Y=2.035
+ $X2=0 $Y2=0
cc_590 N_A_114_368#_c_791_n N_A_531_368#_c_921_n 0.0151327f $X=9.595 $Y=2.035
+ $X2=0 $Y2=0
cc_591 N_A_114_368#_M1013_s N_A_531_368#_c_853_n 0.00197722f $X=9.61 $Y=1.84
+ $X2=0 $Y2=0
cc_592 N_A_114_368#_c_801_n N_A_531_368#_c_853_n 0.0160777f $X=9.76 $Y=2.035
+ $X2=0 $Y2=0
cc_593 N_A_114_368#_c_801_n N_A_531_368#_c_854_n 0.0533059f $X=9.76 $Y=2.035
+ $X2=0 $Y2=0
cc_594 N_A_114_368#_c_744_n N_A_531_368#_c_855_n 0.0222415f $X=6.895 $Y=2.035
+ $X2=0 $Y2=0
cc_595 N_A_114_368#_c_744_n N_A_531_368#_c_856_n 0.0173542f $X=6.895 $Y=2.035
+ $X2=0 $Y2=0
cc_596 N_A_114_368#_c_744_n N_A_531_368#_c_857_n 0.0173542f $X=6.895 $Y=2.035
+ $X2=0 $Y2=0
cc_597 N_A_114_368#_c_744_n N_A_531_368#_c_858_n 0.0173542f $X=6.895 $Y=2.035
+ $X2=0 $Y2=0
cc_598 N_A_114_368#_c_744_n N_VPWR_M1016_d 0.00359847f $X=6.895 $Y=2.035
+ $X2=-0.19 $Y2=1.66
cc_599 N_A_114_368#_c_744_n N_VPWR_M1021_d 0.00359847f $X=6.895 $Y=2.035 $X2=0
+ $Y2=0
cc_600 N_A_114_368#_c_744_n N_VPWR_M1000_d 0.00359847f $X=6.895 $Y=2.035 $X2=0
+ $Y2=0
cc_601 N_A_114_368#_c_744_n N_VPWR_M1029_d 0.0100873f $X=6.895 $Y=2.035 $X2=0
+ $Y2=0
cc_602 N_A_531_368#_c_863_n N_VPWR_M1016_d 0.00428955f $X=3.515 $Y=2.375
+ $X2=-0.19 $Y2=1.66
cc_603 N_A_531_368#_c_865_n N_VPWR_M1021_d 0.00428955f $X=4.415 $Y=2.375 $X2=0
+ $Y2=0
cc_604 N_A_531_368#_c_875_n N_VPWR_M1000_d 0.00428955f $X=5.315 $Y=2.375 $X2=0
+ $Y2=0
cc_605 N_A_531_368#_c_877_n N_VPWR_M1029_d 0.0100354f $X=6.445 $Y=2.375 $X2=0
+ $Y2=0
cc_606 N_A_531_368#_c_863_n N_VPWR_c_971_n 0.0136682f $X=3.515 $Y=2.375 $X2=0
+ $Y2=0
cc_607 N_A_531_368#_c_855_n N_VPWR_c_971_n 0.0228252f $X=2.78 $Y=2.4 $X2=0 $Y2=0
cc_608 N_A_531_368#_c_856_n N_VPWR_c_971_n 0.0228252f $X=3.68 $Y=2.4 $X2=0 $Y2=0
cc_609 N_A_531_368#_c_856_n N_VPWR_c_972_n 0.0145674f $X=3.68 $Y=2.4 $X2=0 $Y2=0
cc_610 N_A_531_368#_c_865_n N_VPWR_c_973_n 0.0136682f $X=4.415 $Y=2.375 $X2=0
+ $Y2=0
cc_611 N_A_531_368#_c_856_n N_VPWR_c_973_n 0.0228252f $X=3.68 $Y=2.4 $X2=0 $Y2=0
cc_612 N_A_531_368#_c_857_n N_VPWR_c_973_n 0.0228252f $X=4.58 $Y=2.4 $X2=0 $Y2=0
cc_613 N_A_531_368#_c_875_n N_VPWR_c_974_n 0.0136682f $X=5.315 $Y=2.375 $X2=0
+ $Y2=0
cc_614 N_A_531_368#_c_857_n N_VPWR_c_974_n 0.0228252f $X=4.58 $Y=2.4 $X2=0 $Y2=0
cc_615 N_A_531_368#_c_858_n N_VPWR_c_974_n 0.0228252f $X=5.48 $Y=2.4 $X2=0 $Y2=0
cc_616 N_A_531_368#_c_877_n N_VPWR_c_975_n 0.0338452f $X=6.445 $Y=2.375 $X2=0
+ $Y2=0
cc_617 N_A_531_368#_c_850_n N_VPWR_c_975_n 0.0121691f $X=6.725 $Y=2.99 $X2=0
+ $Y2=0
cc_618 N_A_531_368#_c_858_n N_VPWR_c_975_n 0.013964f $X=5.48 $Y=2.4 $X2=0 $Y2=0
cc_619 N_A_531_368#_c_855_n N_VPWR_c_976_n 0.0146094f $X=2.78 $Y=2.4 $X2=0 $Y2=0
cc_620 N_A_531_368#_c_857_n N_VPWR_c_978_n 0.0145674f $X=4.58 $Y=2.4 $X2=0 $Y2=0
cc_621 N_A_531_368#_c_858_n N_VPWR_c_980_n 0.0145674f $X=5.48 $Y=2.4 $X2=0 $Y2=0
cc_622 N_A_531_368#_c_849_n N_VPWR_c_981_n 0.0422287f $X=7.395 $Y=2.99 $X2=0
+ $Y2=0
cc_623 N_A_531_368#_c_850_n N_VPWR_c_981_n 0.0200196f $X=6.725 $Y=2.99 $X2=0
+ $Y2=0
cc_624 N_A_531_368#_c_851_n N_VPWR_c_981_n 0.0422287f $X=8.295 $Y=2.99 $X2=0
+ $Y2=0
cc_625 N_A_531_368#_c_852_n N_VPWR_c_981_n 0.0422287f $X=9.195 $Y=2.99 $X2=0
+ $Y2=0
cc_626 N_A_531_368#_c_853_n N_VPWR_c_981_n 0.0620829f $X=10.125 $Y=2.99 $X2=0
+ $Y2=0
cc_627 N_A_531_368#_c_859_n N_VPWR_c_981_n 0.016488f $X=7.51 $Y=2.99 $X2=0 $Y2=0
cc_628 N_A_531_368#_c_860_n N_VPWR_c_981_n 0.016488f $X=8.41 $Y=2.99 $X2=0 $Y2=0
cc_629 N_A_531_368#_c_861_n N_VPWR_c_981_n 0.016488f $X=9.31 $Y=2.99 $X2=0 $Y2=0
cc_630 N_A_531_368#_c_849_n N_VPWR_c_970_n 0.0238173f $X=7.395 $Y=2.99 $X2=0
+ $Y2=0
cc_631 N_A_531_368#_c_850_n N_VPWR_c_970_n 0.0108171f $X=6.725 $Y=2.99 $X2=0
+ $Y2=0
cc_632 N_A_531_368#_c_851_n N_VPWR_c_970_n 0.0238173f $X=8.295 $Y=2.99 $X2=0
+ $Y2=0
cc_633 N_A_531_368#_c_852_n N_VPWR_c_970_n 0.0238173f $X=9.195 $Y=2.99 $X2=0
+ $Y2=0
cc_634 N_A_531_368#_c_853_n N_VPWR_c_970_n 0.0346647f $X=10.125 $Y=2.99 $X2=0
+ $Y2=0
cc_635 N_A_531_368#_c_855_n N_VPWR_c_970_n 0.0120527f $X=2.78 $Y=2.4 $X2=0 $Y2=0
cc_636 N_A_531_368#_c_856_n N_VPWR_c_970_n 0.0119851f $X=3.68 $Y=2.4 $X2=0 $Y2=0
cc_637 N_A_531_368#_c_857_n N_VPWR_c_970_n 0.0119851f $X=4.58 $Y=2.4 $X2=0 $Y2=0
cc_638 N_A_531_368#_c_858_n N_VPWR_c_970_n 0.0119851f $X=5.48 $Y=2.4 $X2=0 $Y2=0
cc_639 N_A_531_368#_c_859_n N_VPWR_c_970_n 0.00894187f $X=7.51 $Y=2.99 $X2=0
+ $Y2=0
cc_640 N_A_531_368#_c_860_n N_VPWR_c_970_n 0.00894187f $X=8.41 $Y=2.99 $X2=0
+ $Y2=0
cc_641 N_A_531_368#_c_861_n N_VPWR_c_970_n 0.00894187f $X=9.31 $Y=2.99 $X2=0
+ $Y2=0
cc_642 N_A_531_368#_c_854_n N_A_1326_74#_c_1316_n 0.00864987f $X=10.21 $Y=1.985
+ $X2=0 $Y2=0
cc_643 N_VGND_c_1087_n N_A_534_74#_c_1225_n 0.00897147f $X=3.225 $Y=0.495 $X2=0
+ $Y2=0
cc_644 N_VGND_c_1092_n N_A_534_74#_c_1225_n 0.0109251f $X=3.06 $Y=0 $X2=0 $Y2=0
cc_645 N_VGND_c_1097_n N_A_534_74#_c_1225_n 0.00910508f $X=10.32 $Y=0 $X2=0
+ $Y2=0
cc_646 N_VGND_M1004_d N_A_534_74#_c_1234_n 0.0033542f $X=3.085 $Y=0.37 $X2=0
+ $Y2=0
cc_647 N_VGND_c_1087_n N_A_534_74#_c_1234_n 0.0165203f $X=3.225 $Y=0.495 $X2=0
+ $Y2=0
cc_648 N_VGND_c_1092_n N_A_534_74#_c_1234_n 0.00197156f $X=3.06 $Y=0 $X2=0 $Y2=0
cc_649 N_VGND_c_1093_n N_A_534_74#_c_1234_n 0.00197156f $X=3.92 $Y=0 $X2=0 $Y2=0
cc_650 N_VGND_c_1097_n N_A_534_74#_c_1234_n 0.00938221f $X=10.32 $Y=0 $X2=0
+ $Y2=0
cc_651 N_VGND_c_1087_n N_A_534_74#_c_1227_n 0.00893007f $X=3.225 $Y=0.495 $X2=0
+ $Y2=0
cc_652 N_VGND_c_1088_n N_A_534_74#_c_1227_n 0.00893007f $X=4.085 $Y=0.495 $X2=0
+ $Y2=0
cc_653 N_VGND_c_1093_n N_A_534_74#_c_1227_n 0.00740085f $X=3.92 $Y=0 $X2=0 $Y2=0
cc_654 N_VGND_c_1097_n N_A_534_74#_c_1227_n 0.00616796f $X=10.32 $Y=0 $X2=0
+ $Y2=0
cc_655 N_VGND_M1018_d N_A_534_74#_c_1238_n 0.0033542f $X=3.945 $Y=0.37 $X2=0
+ $Y2=0
cc_656 N_VGND_c_1088_n N_A_534_74#_c_1238_n 0.0165203f $X=4.085 $Y=0.495 $X2=0
+ $Y2=0
cc_657 N_VGND_c_1093_n N_A_534_74#_c_1238_n 0.00197156f $X=3.92 $Y=0 $X2=0 $Y2=0
cc_658 N_VGND_c_1094_n N_A_534_74#_c_1238_n 0.00197156f $X=8.74 $Y=0 $X2=0 $Y2=0
cc_659 N_VGND_c_1097_n N_A_534_74#_c_1238_n 0.00938221f $X=10.32 $Y=0 $X2=0
+ $Y2=0
cc_660 N_VGND_c_1094_n N_A_534_74#_c_1228_n 0.025931f $X=8.74 $Y=0 $X2=0 $Y2=0
cc_661 N_VGND_c_1097_n N_A_534_74#_c_1228_n 0.0182041f $X=10.32 $Y=0 $X2=0 $Y2=0
cc_662 N_VGND_c_1088_n N_A_534_74#_c_1229_n 0.009209f $X=4.085 $Y=0.495 $X2=0
+ $Y2=0
cc_663 N_VGND_c_1094_n N_A_534_74#_c_1229_n 0.0137625f $X=8.74 $Y=0 $X2=0 $Y2=0
cc_664 N_VGND_c_1097_n N_A_534_74#_c_1229_n 0.009357f $X=10.32 $Y=0 $X2=0 $Y2=0
cc_665 N_VGND_c_1094_n N_A_534_74#_c_1230_n 0.0259505f $X=8.74 $Y=0 $X2=0 $Y2=0
cc_666 N_VGND_c_1097_n N_A_534_74#_c_1230_n 0.018208f $X=10.32 $Y=0 $X2=0 $Y2=0
cc_667 N_VGND_c_1094_n N_A_534_74#_c_1231_n 0.0181125f $X=8.74 $Y=0 $X2=0 $Y2=0
cc_668 N_VGND_c_1097_n N_A_534_74#_c_1231_n 0.0122715f $X=10.32 $Y=0 $X2=0 $Y2=0
cc_669 N_VGND_c_1094_n N_A_534_74#_c_1232_n 0.0174556f $X=8.74 $Y=0 $X2=0 $Y2=0
cc_670 N_VGND_c_1097_n N_A_534_74#_c_1232_n 0.0121438f $X=10.32 $Y=0 $X2=0 $Y2=0
cc_671 N_VGND_c_1089_n N_A_1326_74#_c_1312_n 0.00985092f $X=8.905 $Y=0.675 $X2=0
+ $Y2=0
cc_672 N_VGND_c_1094_n N_A_1326_74#_c_1312_n 0.00758556f $X=8.74 $Y=0 $X2=0
+ $Y2=0
cc_673 N_VGND_c_1097_n N_A_1326_74#_c_1312_n 0.00627867f $X=10.32 $Y=0 $X2=0
+ $Y2=0
cc_674 N_VGND_M1006_s N_A_1326_74#_c_1313_n 0.00176461f $X=8.765 $Y=0.37 $X2=0
+ $Y2=0
cc_675 N_VGND_c_1089_n N_A_1326_74#_c_1313_n 0.0170777f $X=8.905 $Y=0.675 $X2=0
+ $Y2=0
cc_676 N_VGND_c_1089_n N_A_1326_74#_c_1315_n 0.0182488f $X=8.905 $Y=0.675 $X2=0
+ $Y2=0
cc_677 N_VGND_c_1090_n N_A_1326_74#_c_1315_n 0.0182488f $X=9.765 $Y=0.675 $X2=0
+ $Y2=0
cc_678 N_VGND_c_1095_n N_A_1326_74#_c_1315_n 0.00749631f $X=9.6 $Y=0 $X2=0 $Y2=0
cc_679 N_VGND_c_1097_n N_A_1326_74#_c_1315_n 0.0062048f $X=10.32 $Y=0 $X2=0
+ $Y2=0
cc_680 N_VGND_M1020_s N_A_1326_74#_c_1316_n 0.00176461f $X=9.625 $Y=0.37 $X2=0
+ $Y2=0
cc_681 N_VGND_c_1090_n N_A_1326_74#_c_1316_n 0.0170777f $X=9.765 $Y=0.675 $X2=0
+ $Y2=0
cc_682 N_VGND_c_1090_n N_A_1326_74#_c_1317_n 0.0182902f $X=9.765 $Y=0.675 $X2=0
+ $Y2=0
cc_683 N_VGND_c_1096_n N_A_1326_74#_c_1317_n 0.011066f $X=10.32 $Y=0 $X2=0 $Y2=0
cc_684 N_VGND_c_1097_n N_A_1326_74#_c_1317_n 0.00915947f $X=10.32 $Y=0 $X2=0
+ $Y2=0
cc_685 N_VGND_c_1094_n N_A_1326_74#_c_1318_n 0.073391f $X=8.74 $Y=0 $X2=0 $Y2=0
cc_686 N_VGND_c_1097_n N_A_1326_74#_c_1318_n 0.0616471f $X=10.32 $Y=0 $X2=0
+ $Y2=0
cc_687 N_A_534_74#_c_1232_n N_A_1326_74#_c_1318_n 0.0264679f $X=6.235 $Y=0.385
+ $X2=0 $Y2=0
