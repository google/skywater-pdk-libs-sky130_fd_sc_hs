* File: sky130_fd_sc_hs__dfrtp_4.pex.spice
* Created: Thu Aug 27 20:38:53 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HS__DFRTP_4%D 2 4 5 7 10 12 13 14 19 20 23
r32 23 25 35.4289 $w=4e-07 $l=1.65e-07 $layer=POLY_cond $X=0.42 $Y=1.845
+ $X2=0.42 $Y2=2.01
r33 23 24 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=0.385
+ $Y=1.845 $X2=0.385 $Y2=1.845
r34 19 21 45.6753 $w=4e-07 $l=1.65e-07 $layer=POLY_cond $X=0.42 $Y=1.165
+ $X2=0.42 $Y2=1
r35 19 20 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=0.385
+ $Y=1.165 $X2=0.385 $Y2=1.165
r36 14 24 5.61447 $w=3.88e-07 $l=1.9e-07 $layer=LI1_cond $X=0.32 $Y=2.035
+ $X2=0.32 $Y2=1.845
r37 13 24 5.31897 $w=3.88e-07 $l=1.8e-07 $layer=LI1_cond $X=0.32 $Y=1.665
+ $X2=0.32 $Y2=1.845
r38 12 13 10.9334 $w=3.88e-07 $l=3.7e-07 $layer=LI1_cond $X=0.32 $Y=1.295
+ $X2=0.32 $Y2=1.665
r39 12 20 3.84148 $w=3.88e-07 $l=1.3e-07 $layer=LI1_cond $X=0.32 $Y=1.295
+ $X2=0.32 $Y2=1.165
r40 10 21 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=0.545 $Y=0.6 $X2=0.545
+ $Y2=1
r41 5 7 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=0.5 $Y=2.465 $X2=0.5
+ $Y2=2.75
r42 4 5 54.6598 $w=1.94e-07 $l=2.27376e-07 $layer=POLY_cond $X=0.515 $Y=2.245
+ $X2=0.5 $Y2=2.465
r43 4 25 74.2101 $w=2.1e-07 $l=2.35e-07 $layer=POLY_cond $X=0.515 $Y=2.245
+ $X2=0.515 $Y2=2.01
r44 2 23 4.86635 $w=4e-07 $l=3.5e-08 $layer=POLY_cond $X=0.42 $Y=1.81 $X2=0.42
+ $Y2=1.845
r45 1 19 4.86635 $w=4e-07 $l=3.5e-08 $layer=POLY_cond $X=0.42 $Y=1.2 $X2=0.42
+ $Y2=1.165
r46 1 2 84.8135 $w=4e-07 $l=6.1e-07 $layer=POLY_cond $X=0.42 $Y=1.2 $X2=0.42
+ $Y2=1.81
.ends

.subckt PM_SKY130_FD_SC_HS__DFRTP_4%RESET_B 3 6 8 9 11 12 14 16 17 19 21 22 24
+ 27 31 34 35 36 37 38 41 43 44 46 49 53 54 57
c214 54 0 1.353e-19 $X=1.155 $Y=1.295
c215 53 0 1.12283e-19 $X=1.155 $Y=1.295
c216 49 0 1.66354e-20 $X=5.25 $Y=1.835
c217 41 0 1.36553e-19 $X=5.52 $Y=2.035
c218 38 0 1.63054e-19 $X=5.665 $Y=2.035
c219 34 0 1.42958e-20 $X=4.87 $Y=1.835
c220 17 0 1.20728e-19 $X=4.87 $Y=2.24
c221 12 0 1.07817e-19 $X=4.765 $Y=1.185
r222 57 59 41.3282 $w=4.6e-07 $l=1.65e-07 $layer=POLY_cond $X=1.09 $Y=1.975
+ $X2=1.09 $Y2=2.14
r223 57 58 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.155
+ $Y=1.975 $X2=1.155 $Y2=1.975
r224 54 58 30.1408 $w=2.58e-07 $l=6.8e-07 $layer=LI1_cond $X=1.155 $Y=1.295
+ $X2=1.155 $Y2=1.975
r225 53 55 47.2161 $w=4.6e-07 $l=1.65e-07 $layer=POLY_cond $X=1.09 $Y=1.295
+ $X2=1.09 $Y2=1.13
r226 53 54 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.155
+ $Y=1.295 $X2=1.155 $Y2=1.295
r227 49 50 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.25
+ $Y=1.835 $X2=5.25 $Y2=1.835
r228 46 58 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=2.035
+ $X2=1.2 $Y2=2.035
r229 44 61 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.975
+ $Y=2.11 $X2=8.975 $Y2=2.11
r230 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=2.035
+ $X2=8.88 $Y2=2.035
r231 41 50 7.17647 $w=4.48e-07 $l=2.7e-07 $layer=LI1_cond $X=5.52 $Y=1.895
+ $X2=5.25 $Y2=1.895
r232 40 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=2.035
+ $X2=5.52 $Y2=2.035
r233 38 40 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.665 $Y=2.035
+ $X2=5.52 $Y2=2.035
r234 37 43 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=8.735 $Y=2.035
+ $X2=8.88 $Y2=2.035
r235 37 38 3.7995 $w=1.4e-07 $l=3.07e-06 $layer=MET1_cond $X=8.735 $Y=2.035
+ $X2=5.665 $Y2=2.035
r236 36 46 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.345 $Y=2.035
+ $X2=1.2 $Y2=2.035
r237 35 40 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.375 $Y=2.035
+ $X2=5.52 $Y2=2.035
r238 35 36 4.98761 $w=1.4e-07 $l=4.03e-06 $layer=MET1_cond $X=5.375 $Y=2.035
+ $X2=1.345 $Y2=2.035
r239 33 49 50.7098 $w=3.3e-07 $l=2.9e-07 $layer=POLY_cond $X=4.96 $Y=1.835
+ $X2=5.25 $Y2=1.835
r240 33 34 3.90195 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=4.96 $Y=1.835
+ $X2=4.87 $Y2=1.835
r241 29 31 61.5319 $w=1.5e-07 $l=1.2e-07 $layer=POLY_cond $X=4.765 $Y=1.26
+ $X2=4.885 $Y2=1.26
r242 25 61 38.6072 $w=2.91e-07 $l=2.03101e-07 $layer=POLY_cond $X=9.06 $Y=1.945
+ $X2=8.975 $Y2=2.11
r243 25 27 681.979 $w=1.5e-07 $l=1.33e-06 $layer=POLY_cond $X=9.06 $Y=1.945
+ $X2=9.06 $Y2=0.615
r244 22 61 57.6553 $w=2.91e-07 $l=3.01662e-07 $layer=POLY_cond $X=9.02 $Y=2.39
+ $X2=8.975 $Y2=2.11
r245 22 24 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=9.02 $Y=2.39
+ $X2=9.02 $Y2=2.675
r246 21 34 34.7346 $w=1.65e-07 $l=1.72337e-07 $layer=POLY_cond $X=4.885 $Y=1.67
+ $X2=4.87 $Y2=1.835
r247 20 31 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.885 $Y=1.335
+ $X2=4.885 $Y2=1.26
r248 20 21 171.777 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=4.885 $Y=1.335
+ $X2=4.885 $Y2=1.67
r249 17 19 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=4.87 $Y=2.24
+ $X2=4.87 $Y2=2.525
r250 16 17 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=4.87 $Y=2.15 $X2=4.87
+ $Y2=2.24
r251 15 34 34.7346 $w=1.65e-07 $l=1.65e-07 $layer=POLY_cond $X=4.87 $Y=2
+ $X2=4.87 $Y2=1.835
r252 15 16 58.3064 $w=1.8e-07 $l=1.5e-07 $layer=POLY_cond $X=4.87 $Y=2 $X2=4.87
+ $Y2=2.15
r253 12 29 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.765 $Y=1.185
+ $X2=4.765 $Y2=1.26
r254 12 14 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=4.765 $Y=1.185
+ $X2=4.765 $Y2=0.9
r255 9 11 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=0.95 $Y=2.465
+ $X2=0.95 $Y2=2.75
r256 8 9 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=0.95 $Y=2.375 $X2=0.95
+ $Y2=2.465
r257 8 59 91.3468 $w=1.8e-07 $l=2.35e-07 $layer=POLY_cond $X=0.95 $Y=2.375
+ $X2=0.95 $Y2=2.14
r258 6 57 7.8587 $w=4.6e-07 $l=6.5e-08 $layer=POLY_cond $X=1.09 $Y=1.91 $X2=1.09
+ $Y2=1.975
r259 5 53 7.8587 $w=4.6e-07 $l=6.5e-08 $layer=POLY_cond $X=1.09 $Y=1.36 $X2=1.09
+ $Y2=1.295
r260 5 6 66.4967 $w=4.6e-07 $l=5.5e-07 $layer=POLY_cond $X=1.09 $Y=1.36 $X2=1.09
+ $Y2=1.91
r261 3 55 271.766 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=0.935 $Y=0.6
+ $X2=0.935 $Y2=1.13
.ends

.subckt PM_SKY130_FD_SC_HS__DFRTP_4%CLK 3 5 7 8
c44 8 0 1.89442e-19 $X=2.16 $Y=1.665
c45 5 0 3.02652e-19 $X=1.945 $Y=1.755
c46 3 0 7.30529e-21 $X=1.925 $Y=0.74
r47 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.93
+ $Y=1.475 $X2=1.93 $Y2=1.475
r48 8 12 7.06801 $w=3.97e-07 $l=2.3e-07 $layer=LI1_cond $X=2.16 $Y=1.545
+ $X2=1.93 $Y2=1.545
r49 5 11 57.6553 $w=2.91e-07 $l=2.87402e-07 $layer=POLY_cond $X=1.945 $Y=1.755
+ $X2=1.93 $Y2=1.475
r50 5 7 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.945 $Y=1.755
+ $X2=1.945 $Y2=2.39
r51 1 11 38.6072 $w=2.91e-07 $l=1.67481e-07 $layer=POLY_cond $X=1.925 $Y=1.31
+ $X2=1.93 $Y2=1.475
r52 1 3 292.277 $w=1.5e-07 $l=5.7e-07 $layer=POLY_cond $X=1.925 $Y=1.31
+ $X2=1.925 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HS__DFRTP_4%A_494_366# 1 2 8 9 11 12 14 16 18 20 21 22
+ 23 25 28 29 31 32 33 35 39 43 47 53 58 62 68 71 73
c201 58 0 1.07817e-19 $X=4.39 $Y=0.415
c202 39 0 9.26151e-20 $X=7.905 $Y=2.14
c203 29 0 1.27872e-19 $X=4.305 $Y=0.415
c204 16 0 1.85309e-19 $X=3.985 $Y=0.9
c205 14 0 1.35567e-19 $X=3.985 $Y=1.385
r206 70 71 9.95292 $w=3.28e-07 $l=2.85e-07 $layer=LI1_cond $X=7.905 $Y=1.18
+ $X2=8.19 $Y2=1.18
r207 68 79 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=7.71 $Y=1.18 $X2=7.71
+ $Y2=1.27
r208 67 70 6.80989 $w=3.28e-07 $l=1.95e-07 $layer=LI1_cond $X=7.71 $Y=1.18
+ $X2=7.905 $Y2=1.18
r209 67 68 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.71
+ $Y=1.18 $X2=7.71 $Y2=1.18
r210 62 64 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=5.48 $Y=0.34
+ $X2=5.48 $Y2=0.625
r211 58 60 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=4.39 $Y=0.415
+ $X2=4.39 $Y2=0.625
r212 54 76 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.355 $Y=1.725
+ $X2=3.355 $Y2=1.89
r213 54 73 10.4917 $w=3.3e-07 $l=6e-08 $layer=POLY_cond $X=3.355 $Y=1.725
+ $X2=3.355 $Y2=1.665
r214 53 54 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.355
+ $Y=1.725 $X2=3.355 $Y2=1.725
r215 50 51 10.8645 $w=4.68e-07 $l=2.25e-07 $layer=LI1_cond $X=2.78 $Y=0.575
+ $X2=2.78 $Y2=0.8
r216 47 50 4.07176 $w=4.68e-07 $l=1.6e-07 $layer=LI1_cond $X=2.78 $Y=0.415
+ $X2=2.78 $Y2=0.575
r217 43 71 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.19 $Y=1.015
+ $X2=8.19 $Y2=1.18
r218 42 43 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=8.19 $Y=0.425
+ $X2=8.19 $Y2=1.015
r219 39 40 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.905
+ $Y=2.14 $X2=7.905 $Y2=2.14
r220 37 70 0.716491 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=7.905 $Y=1.345
+ $X2=7.905 $Y2=1.18
r221 37 39 27.7634 $w=3.28e-07 $l=7.95e-07 $layer=LI1_cond $X=7.905 $Y=1.345
+ $X2=7.905 $Y2=2.14
r222 36 62 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.565 $Y=0.34
+ $X2=5.48 $Y2=0.34
r223 35 42 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.105 $Y=0.34
+ $X2=8.19 $Y2=0.425
r224 35 36 165.711 $w=1.68e-07 $l=2.54e-06 $layer=LI1_cond $X=8.105 $Y=0.34
+ $X2=5.565 $Y2=0.34
r225 34 60 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.475 $Y=0.625
+ $X2=4.39 $Y2=0.625
r226 33 64 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.395 $Y=0.625
+ $X2=5.48 $Y2=0.625
r227 33 34 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=5.395 $Y=0.625
+ $X2=4.475 $Y2=0.625
r228 31 53 3.47907 $w=2.63e-07 $l=8e-08 $layer=LI1_cond $X=3.322 $Y=1.805
+ $X2=3.322 $Y2=1.725
r229 31 32 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=3.19 $Y=1.805
+ $X2=3.015 $Y2=1.805
r230 30 47 6.76998 $w=1.7e-07 $l=2.35e-07 $layer=LI1_cond $X=3.015 $Y=0.415
+ $X2=2.78 $Y2=0.415
r231 29 58 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.305 $Y=0.415
+ $X2=4.39 $Y2=0.415
r232 29 30 84.1604 $w=1.68e-07 $l=1.29e-06 $layer=LI1_cond $X=4.305 $Y=0.415
+ $X2=3.015 $Y2=0.415
r233 28 32 6.35003 $w=3.65e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.93 $Y=1.72
+ $X2=3.015 $Y2=1.805
r234 28 45 10.3616 $w=3.65e-07 $l=4.07247e-07 $layer=LI1_cond $X=2.93 $Y=1.72
+ $X2=2.62 $Y2=1.945
r235 28 51 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=2.93 $Y=1.72
+ $X2=2.93 $Y2=0.8
r236 23 40 50.2556 $w=3.62e-07 $l=3.02076e-07 $layer=POLY_cond $X=8.06 $Y=2.39
+ $X2=7.945 $Y2=2.14
r237 23 25 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=8.06 $Y=2.39
+ $X2=8.06 $Y2=2.675
r238 21 79 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.545 $Y=1.27
+ $X2=7.71 $Y2=1.27
r239 21 22 184.596 $w=1.5e-07 $l=3.6e-07 $layer=POLY_cond $X=7.545 $Y=1.27
+ $X2=7.185 $Y2=1.27
r240 18 22 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=7.11 $Y=1.195
+ $X2=7.185 $Y2=1.27
r241 18 20 146.207 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=7.11 $Y=1.195
+ $X2=7.11 $Y2=0.74
r242 14 26 71.6325 $w=1.96e-07 $l=3.06268e-07 $layer=POLY_cond $X=3.985 $Y=1.385
+ $X2=3.93 $Y2=1.665
r243 14 16 248.691 $w=1.5e-07 $l=4.85e-07 $layer=POLY_cond $X=3.985 $Y=1.385
+ $X2=3.985 $Y2=0.9
r244 13 73 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.52 $Y=1.665
+ $X2=3.355 $Y2=1.665
r245 12 26 9.11062 $w=1.5e-07 $l=1.3e-07 $layer=POLY_cond $X=3.8 $Y=1.665
+ $X2=3.93 $Y2=1.665
r246 12 13 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=3.8 $Y=1.665
+ $X2=3.52 $Y2=1.665
r247 9 11 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=3.42 $Y=2.24 $X2=3.42
+ $Y2=2.525
r248 8 9 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=3.42 $Y=2.15 $X2=3.42
+ $Y2=2.24
r249 8 76 101.065 $w=1.8e-07 $l=2.6e-07 $layer=POLY_cond $X=3.42 $Y=2.15
+ $X2=3.42 $Y2=1.89
r250 2 45 600 $w=1.7e-07 $l=2.22711e-07 $layer=licon1_PDIFF $count=1 $X=2.47
+ $Y=1.83 $X2=2.62 $Y2=1.99
r251 1 50 182 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_NDIFF $count=1 $X=2.57
+ $Y=0.37 $X2=2.71 $Y2=0.575
.ends

.subckt PM_SKY130_FD_SC_HS__DFRTP_4%A_834_355# 1 2 7 9 12 16 20 22 23 25 29 34
c88 34 0 1.52817e-19 $X=6.45 $Y=2.125
c89 29 0 1.42958e-20 $X=5.735 $Y=0.885
c90 23 0 5.12321e-20 $X=6.325 $Y=0.885
c91 20 0 1.85309e-19 $X=4.57 $Y=0.965
c92 12 0 3.01223e-20 $X=4.375 $Y=0.9
r93 28 30 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=5.9 $Y=0.885
+ $X2=6.24 $Y2=0.885
r94 28 29 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=5.9 $Y=0.885
+ $X2=5.735 $Y2=0.885
r95 23 30 2.96841 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=6.325 $Y=0.885
+ $X2=6.24 $Y2=0.885
r96 23 25 17.4613 $w=3.28e-07 $l=5e-07 $layer=LI1_cond $X=6.325 $Y=0.885
+ $X2=6.825 $Y2=0.885
r97 22 34 8.20383 $w=2.93e-07 $l=2.1e-07 $layer=LI1_cond $X=6.24 $Y=2.087
+ $X2=6.45 $Y2=2.087
r98 21 30 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.24 $Y=1.05
+ $X2=6.24 $Y2=0.885
r99 21 22 58.0642 $w=1.68e-07 $l=8.9e-07 $layer=LI1_cond $X=6.24 $Y=1.05
+ $X2=6.24 $Y2=1.94
r100 20 29 76.0053 $w=1.68e-07 $l=1.165e-06 $layer=LI1_cond $X=4.57 $Y=0.965
+ $X2=5.735 $Y2=0.965
r101 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.405
+ $Y=1.94 $X2=4.405 $Y2=1.94
r102 14 20 7.24806 $w=1.7e-07 $l=1.70276e-07 $layer=LI1_cond $X=4.437 $Y=1.05
+ $X2=4.57 $Y2=0.965
r103 14 16 38.7047 $w=2.63e-07 $l=8.9e-07 $layer=LI1_cond $X=4.437 $Y=1.05
+ $X2=4.437 $Y2=1.94
r104 10 17 38.6446 $w=3.36e-07 $l=1.67481e-07 $layer=POLY_cond $X=4.375 $Y=1.775
+ $X2=4.37 $Y2=1.94
r105 10 12 448.67 $w=1.5e-07 $l=8.75e-07 $layer=POLY_cond $X=4.375 $Y=1.775
+ $X2=4.375 $Y2=0.9
r106 7 17 58.0107 $w=3.36e-07 $l=3.50714e-07 $layer=POLY_cond $X=4.26 $Y=2.24
+ $X2=4.37 $Y2=1.94
r107 7 9 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=4.26 $Y=2.24 $X2=4.26
+ $Y2=2.525
r108 2 34 600 $w=1.7e-07 $l=2.2798e-07 $layer=licon1_PDIFF $count=1 $X=6.3
+ $Y=1.96 $X2=6.45 $Y2=2.125
r109 1 28 182 $w=1.7e-07 $l=5.80797e-07 $layer=licon1_NDIFF $count=1 $X=5.76
+ $Y=0.37 $X2=5.9 $Y2=0.885
r110 1 25 91 $w=1.7e-07 $l=1.29719e-06 $layer=licon1_NDIFF $count=2 $X=5.76
+ $Y=0.37 $X2=6.825 $Y2=0.885
.ends

.subckt PM_SKY130_FD_SC_HS__DFRTP_4%A_313_74# 1 2 7 9 10 12 13 16 17 18 19 21 22
+ 23 24 26 27 30 31 33 34 38 41 44 46 49 52 53 57 58 60 63 64 68 71 72 80
c227 72 0 1.76168e-19 $X=5.56 $Y=2.375
c228 71 0 2.76281e-19 $X=5.56 $Y=2.375
c229 64 0 1.12283e-19 $X=1.665 $Y=1.055
c230 63 0 1.35587e-19 $X=6.87 $Y=2.405
c231 57 0 1.74657e-19 $X=2.56 $Y=1.385
c232 13 0 1.05803e-19 $X=3.41 $Y=1.275
c233 10 0 1.27872e-19 $X=2.495 $Y=1.2
c234 7 0 1.89442e-19 $X=2.395 $Y=1.755
r235 78 88 41.4908 $w=2.73e-07 $l=2.35e-07 $layer=POLY_cond $X=6.66 $Y=1.425
+ $X2=6.66 $Y2=1.66
r236 77 80 7.33373 $w=3.28e-07 $l=2.1e-07 $layer=LI1_cond $X=6.66 $Y=1.425
+ $X2=6.87 $Y2=1.425
r237 77 78 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.66
+ $Y=1.425 $X2=6.66 $Y2=1.425
r238 72 83 30.6007 $w=3.3e-07 $l=1.75e-07 $layer=POLY_cond $X=5.56 $Y=2.375
+ $X2=5.385 $Y2=2.375
r239 71 74 4.01609 $w=3.28e-07 $l=1.15e-07 $layer=LI1_cond $X=5.56 $Y=2.375
+ $X2=5.56 $Y2=2.49
r240 71 72 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.56
+ $Y=2.375 $X2=5.56 $Y2=2.375
r241 65 68 6.28605 $w=3.28e-07 $l=1.8e-07 $layer=LI1_cond $X=1.54 $Y=1.975
+ $X2=1.72 $Y2=1.975
r242 62 80 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.87 $Y=1.59
+ $X2=6.87 $Y2=1.425
r243 62 63 53.1711 $w=1.68e-07 $l=8.15e-07 $layer=LI1_cond $X=6.87 $Y=1.59
+ $X2=6.87 $Y2=2.405
r244 61 74 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.725 $Y=2.49
+ $X2=5.56 $Y2=2.49
r245 60 63 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.785 $Y=2.49
+ $X2=6.87 $Y2=2.405
r246 60 61 69.1551 $w=1.68e-07 $l=1.06e-06 $layer=LI1_cond $X=6.785 $Y=2.49
+ $X2=5.725 $Y2=2.49
r247 57 58 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.56
+ $Y=1.385 $X2=2.56 $Y2=1.385
r248 55 57 12.276 $w=2.28e-07 $l=2.45e-07 $layer=LI1_cond $X=2.56 $Y=1.14
+ $X2=2.56 $Y2=1.385
r249 54 64 3.3845 $w=1.7e-07 $l=2.1e-07 $layer=LI1_cond $X=1.875 $Y=1.055
+ $X2=1.665 $Y2=1.055
r250 53 55 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=2.445 $Y=1.055
+ $X2=2.56 $Y2=1.14
r251 53 54 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=2.445 $Y=1.055
+ $X2=1.875 $Y2=1.055
r252 52 65 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.54 $Y=1.81
+ $X2=1.54 $Y2=1.975
r253 51 64 3.19717 $w=2.95e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.54 $Y=1.14
+ $X2=1.665 $Y2=1.055
r254 51 52 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.54 $Y=1.14
+ $X2=1.54 $Y2=1.81
r255 47 64 3.19717 $w=2.95e-07 $l=8.5e-08 $layer=LI1_cond $X=1.665 $Y=0.97
+ $X2=1.665 $Y2=1.055
r256 47 49 12.4848 $w=4.18e-07 $l=4.55e-07 $layer=LI1_cond $X=1.665 $Y=0.97
+ $X2=1.665 $Y2=0.515
r257 44 58 27.1456 $w=4.2e-07 $l=2.05e-07 $layer=POLY_cond $X=2.515 $Y=1.59
+ $X2=2.515 $Y2=1.385
r258 42 44 37.5584 $w=1.54e-07 $l=1.2e-07 $layer=POLY_cond $X=2.395 $Y=1.672
+ $X2=2.515 $Y2=1.672
r259 40 58 4.63462 $w=4.2e-07 $l=3.5e-08 $layer=POLY_cond $X=2.515 $Y=1.35
+ $X2=2.515 $Y2=1.385
r260 40 41 11.6336 $w=2.85e-07 $l=7.5e-08 $layer=POLY_cond $X=2.515 $Y=1.35
+ $X2=2.515 $Y2=1.275
r261 36 38 497.383 $w=1.5e-07 $l=9.7e-07 $layer=POLY_cond $X=8.16 $Y=1.585
+ $X2=8.16 $Y2=0.615
r262 35 88 16.7618 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.825 $Y=1.66
+ $X2=6.66 $Y2=1.66
r263 34 36 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=8.085 $Y=1.66
+ $X2=8.16 $Y2=1.585
r264 34 35 646.085 $w=1.5e-07 $l=1.26e-06 $layer=POLY_cond $X=8.085 $Y=1.66
+ $X2=6.825 $Y2=1.66
r265 31 88 49.4375 $w=2.73e-07 $l=2.32379e-07 $layer=POLY_cond $X=6.675 $Y=1.885
+ $X2=6.66 $Y2=1.66
r266 31 33 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=6.675 $Y=1.885
+ $X2=6.675 $Y2=2.46
r267 29 83 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.385 $Y=2.54
+ $X2=5.385 $Y2=2.375
r268 29 30 274.33 $w=1.5e-07 $l=5.35e-07 $layer=POLY_cond $X=5.385 $Y=2.54
+ $X2=5.385 $Y2=3.075
r269 28 46 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=3.96 $Y=3.15 $X2=3.87
+ $Y2=3.15
r270 27 30 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.31 $Y=3.15
+ $X2=5.385 $Y2=3.075
r271 27 28 692.234 $w=1.5e-07 $l=1.35e-06 $layer=POLY_cond $X=5.31 $Y=3.15
+ $X2=3.96 $Y2=3.15
r272 24 26 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=3.87 $Y=2.81
+ $X2=3.87 $Y2=2.525
r273 23 46 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=3.87 $Y=3.075
+ $X2=3.87 $Y2=3.15
r274 22 24 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=3.87 $Y=2.9 $X2=3.87
+ $Y2=2.81
r275 22 23 68.0242 $w=1.8e-07 $l=1.75e-07 $layer=POLY_cond $X=3.87 $Y=2.9
+ $X2=3.87 $Y2=3.075
r276 19 21 96.4 $w=1.5e-07 $l=3e-07 $layer=POLY_cond $X=3.485 $Y=1.2 $X2=3.485
+ $Y2=0.9
r277 17 46 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=3.78 $Y=3.15 $X2=3.87
+ $Y2=3.15
r278 17 18 410.213 $w=1.5e-07 $l=8e-07 $layer=POLY_cond $X=3.78 $Y=3.15 $X2=2.98
+ $Y2=3.15
r279 16 18 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.905 $Y=3.075
+ $X2=2.98 $Y2=3.15
r280 15 44 122.065 $w=1.54e-07 $l=3.9e-07 $layer=POLY_cond $X=2.905 $Y=1.672
+ $X2=2.515 $Y2=1.672
r281 15 16 684.543 $w=1.5e-07 $l=1.335e-06 $layer=POLY_cond $X=2.905 $Y=1.74
+ $X2=2.905 $Y2=3.075
r282 14 41 14.7291 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=2.725 $Y=1.275
+ $X2=2.515 $Y2=1.275
r283 13 19 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.41 $Y=1.275
+ $X2=3.485 $Y2=1.2
r284 13 14 351.245 $w=1.5e-07 $l=6.85e-07 $layer=POLY_cond $X=3.41 $Y=1.275
+ $X2=2.725 $Y2=1.275
r285 10 41 11.6336 $w=2.85e-07 $l=8.44097e-08 $layer=POLY_cond $X=2.495 $Y=1.2
+ $X2=2.515 $Y2=1.275
r286 10 12 147.813 $w=1.5e-07 $l=4.6e-07 $layer=POLY_cond $X=2.495 $Y=1.2
+ $X2=2.495 $Y2=0.74
r287 7 42 3.46277 $w=1.5e-07 $l=8.3e-08 $layer=POLY_cond $X=2.395 $Y=1.755
+ $X2=2.395 $Y2=1.672
r288 7 9 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.395 $Y=1.755
+ $X2=2.395 $Y2=2.39
r289 2 68 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.58
+ $Y=1.83 $X2=1.72 $Y2=1.975
r290 1 49 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=1.565
+ $Y=0.37 $X2=1.71 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__DFRTP_4%A_699_463# 1 2 3 10 12 15 17 18 19 20 22 23
+ 24 26 27 29 36 38
c133 26 0 1.38917e-19 $X=4.83 $Y=2.295
c134 23 0 1.50343e-19 $X=4.745 $Y=2.485
c135 22 0 1.05803e-19 $X=4.05 $Y=2.4
c136 20 0 1.30745e-19 $X=6.225 $Y=1.73
c137 18 0 2.99607e-19 $X=5.76 $Y=1.385
c138 15 0 5.6074e-20 $X=6.225 $Y=1.885
r139 38 40 8.354 $w=3.87e-07 $l=2.65e-07 $layer=LI1_cond $X=4.83 $Y=2.525
+ $X2=5.095 $Y2=2.525
r140 33 34 19.764 $w=2.5e-07 $l=4.05e-07 $layer=LI1_cond $X=3.645 $Y=2.57
+ $X2=4.05 $Y2=2.57
r141 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.82
+ $Y=1.385 $X2=5.82 $Y2=1.385
r142 27 29 37.2486 $w=2.78e-07 $l=9.05e-07 $layer=LI1_cond $X=4.915 $Y=1.36
+ $X2=5.82 $Y2=1.36
r143 26 38 5.57805 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=4.83 $Y=2.295
+ $X2=4.83 $Y2=2.525
r144 25 27 7.36005 $w=2.8e-07 $l=1.77482e-07 $layer=LI1_cond $X=4.83 $Y=1.5
+ $X2=4.915 $Y2=1.36
r145 25 26 51.8663 $w=1.68e-07 $l=7.95e-07 $layer=LI1_cond $X=4.83 $Y=1.5
+ $X2=4.83 $Y2=2.295
r146 24 34 5.40474 $w=2.5e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.135 $Y=2.485
+ $X2=4.05 $Y2=2.57
r147 23 38 6.57826 $w=3.87e-07 $l=1.03078e-07 $layer=LI1_cond $X=4.745 $Y=2.485
+ $X2=4.83 $Y2=2.525
r148 23 24 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=4.745 $Y=2.485
+ $X2=4.135 $Y2=2.485
r149 22 34 2.99516 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=4.05 $Y=2.4 $X2=4.05
+ $Y2=2.57
r150 21 36 11.3867 $w=3e-07 $l=3.62767e-07 $layer=LI1_cond $X=4.05 $Y=1.05
+ $X2=3.77 $Y2=0.86
r151 21 22 88.0749 $w=1.68e-07 $l=1.35e-06 $layer=LI1_cond $X=4.05 $Y=1.05
+ $X2=4.05 $Y2=2.4
r152 19 30 55.0813 $w=3.3e-07 $l=3.15e-07 $layer=POLY_cond $X=6.135 $Y=1.385
+ $X2=5.82 $Y2=1.385
r153 18 30 10.4917 $w=3.3e-07 $l=6e-08 $layer=POLY_cond $X=5.76 $Y=1.385
+ $X2=5.82 $Y2=1.385
r154 15 20 60.25 $w=1.8e-07 $l=1.55e-07 $layer=POLY_cond $X=6.225 $Y=1.885
+ $X2=6.225 $Y2=1.73
r155 15 17 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=6.225 $Y=1.885
+ $X2=6.225 $Y2=2.46
r156 13 19 32.1775 $w=3.3e-07 $l=1.98997e-07 $layer=POLY_cond $X=6.21 $Y=1.55
+ $X2=6.135 $Y2=1.385
r157 13 20 92.2979 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=6.21 $Y=1.55
+ $X2=6.21 $Y2=1.73
r158 10 18 17.4878 $w=4.41e-07 $l=1.98997e-07 $layer=POLY_cond $X=5.685 $Y=1.22
+ $X2=5.76 $Y2=1.385
r159 10 12 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=5.685 $Y=1.22
+ $X2=5.685 $Y2=0.74
r160 3 40 600 $w=1.7e-07 $l=2.74955e-07 $layer=licon1_PDIFF $count=1 $X=4.945
+ $Y=2.315 $X2=5.095 $Y2=2.525
r161 2 33 600 $w=1.7e-07 $l=3.26497e-07 $layer=licon1_PDIFF $count=1 $X=3.495
+ $Y=2.315 $X2=3.645 $Y2=2.575
r162 1 36 182 $w=1.7e-07 $l=2.82489e-07 $layer=licon1_NDIFF $count=1 $X=3.56
+ $Y=0.69 $X2=3.77 $Y2=0.86
.ends

.subckt PM_SKY130_FD_SC_HS__DFRTP_4%A_1678_395# 1 2 8 9 11 16 18 19 20 23 24 25
+ 28 31 32 36 41 43
c124 31 0 1.27304e-19 $X=9.86 $Y=1.875
c125 24 0 1.26505e-19 $X=9.775 $Y=1.96
c126 18 0 9.26151e-20 $X=8.492 $Y=1.975
r127 39 41 3.90026 $w=4.58e-07 $l=1.5e-07 $layer=LI1_cond $X=9.245 $Y=2.675
+ $X2=9.395 $Y2=2.675
r128 36 46 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=8.61 $Y=1.2
+ $X2=8.61 $Y2=1.365
r129 36 45 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=8.61 $Y=1.2
+ $X2=8.61 $Y2=1.035
r130 35 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.61
+ $Y=1.2 $X2=8.61 $Y2=1.2
r131 32 35 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=8.61 $Y=1.12 $X2=8.61
+ $Y2=1.2
r132 30 43 3.70735 $w=2.5e-07 $l=1.75425e-07 $layer=LI1_cond $X=9.86 $Y=1.205
+ $X2=9.722 $Y2=1.12
r133 30 31 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=9.86 $Y=1.205
+ $X2=9.86 $Y2=1.875
r134 26 43 3.70735 $w=2.5e-07 $l=1.09864e-07 $layer=LI1_cond $X=9.665 $Y=1.035
+ $X2=9.722 $Y2=1.12
r135 26 28 14.6675 $w=3.28e-07 $l=4.2e-07 $layer=LI1_cond $X=9.665 $Y=1.035
+ $X2=9.665 $Y2=0.615
r136 24 31 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.775 $Y=1.96
+ $X2=9.86 $Y2=1.875
r137 24 25 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=9.775 $Y=1.96
+ $X2=9.48 $Y2=1.96
r138 23 41 6.6364 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=9.395 $Y=2.445
+ $X2=9.395 $Y2=2.675
r139 22 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.395 $Y=2.045
+ $X2=9.48 $Y2=1.96
r140 22 23 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=9.395 $Y=2.045
+ $X2=9.395 $Y2=2.445
r141 21 32 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.775 $Y=1.12
+ $X2=8.61 $Y2=1.12
r142 20 43 2.76166 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=9.5 $Y=1.12
+ $X2=9.722 $Y2=1.12
r143 20 21 47.2995 $w=1.68e-07 $l=7.25e-07 $layer=LI1_cond $X=9.5 $Y=1.12
+ $X2=8.775 $Y2=1.12
r144 18 19 60.4563 $w=1.8e-07 $l=1.5e-07 $layer=POLY_cond $X=8.492 $Y=1.975
+ $X2=8.492 $Y2=2.125
r145 18 46 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=8.52 $Y=1.975
+ $X2=8.52 $Y2=1.365
r146 16 45 215.362 $w=1.5e-07 $l=4.2e-07 $layer=POLY_cond $X=8.55 $Y=0.615
+ $X2=8.55 $Y2=1.035
r147 9 11 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=8.48 $Y=2.39 $X2=8.48
+ $Y2=2.675
r148 8 9 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=8.48 $Y=2.3 $X2=8.48
+ $Y2=2.39
r149 8 19 68.0242 $w=1.8e-07 $l=1.75e-07 $layer=POLY_cond $X=8.48 $Y=2.3
+ $X2=8.48 $Y2=2.125
r150 2 39 600 $w=1.7e-07 $l=2.74955e-07 $layer=licon1_PDIFF $count=1 $X=9.095
+ $Y=2.465 $X2=9.245 $Y2=2.675
r151 1 28 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=9.525
+ $Y=0.405 $X2=9.665 $Y2=0.615
.ends

.subckt PM_SKY130_FD_SC_HS__DFRTP_4%A_1350_392# 1 2 9 12 13 15 16 19 20 22 23 26
+ 27 29 31 34 35 36 37 38 39 40 43 45 50 51 52 58 59
c166 50 0 1.00633e-19 $X=8.325 $Y=2.475
c167 38 0 1.07146e-19 $X=10.475 $Y=1.335
c168 27 0 5.64102e-20 $X=10.425 $Y=1.97
c169 26 0 1.97399e-19 $X=10.425 $Y=1.88
r170 65 66 24.9528 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=9.51 $Y=1.63
+ $X2=9.51 $Y2=1.705
r171 59 65 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=9.51 $Y=1.54 $X2=9.51
+ $Y2=1.63
r172 59 64 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=9.51 $Y=1.54
+ $X2=9.51 $Y2=1.375
r173 58 61 3.54598 $w=2.58e-07 $l=8e-08 $layer=LI1_cond $X=9.475 $Y=1.54
+ $X2=9.475 $Y2=1.62
r174 58 59 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.51
+ $Y=1.54 $X2=9.51 $Y2=1.54
r175 51 61 3.22376 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=9.345 $Y=1.62
+ $X2=9.475 $Y2=1.62
r176 51 52 61 $w=1.68e-07 $l=9.35e-07 $layer=LI1_cond $X=9.345 $Y=1.62 $X2=8.41
+ $Y2=1.62
r177 49 52 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.325 $Y=1.705
+ $X2=8.41 $Y2=1.62
r178 49 50 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=8.325 $Y=1.705
+ $X2=8.325 $Y2=2.475
r179 46 54 2.79691 $w=3.3e-07 $l=1.03e-07 $layer=LI1_cond $X=7.33 $Y=2.64
+ $X2=7.227 $Y2=2.64
r180 46 48 17.6359 $w=3.28e-07 $l=5.05e-07 $layer=LI1_cond $X=7.33 $Y=2.64
+ $X2=7.835 $Y2=2.64
r181 45 50 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=8.24 $Y=2.64
+ $X2=8.325 $Y2=2.475
r182 45 48 14.1436 $w=3.28e-07 $l=4.05e-07 $layer=LI1_cond $X=8.24 $Y=2.64
+ $X2=7.835 $Y2=2.64
r183 41 56 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=7.33 $Y=0.72
+ $X2=7.245 $Y2=0.72
r184 41 43 20.283 $w=2.48e-07 $l=4.4e-07 $layer=LI1_cond $X=7.33 $Y=0.72
+ $X2=7.77 $Y2=0.72
r185 40 54 4.96927 $w=1.7e-07 $l=1.73767e-07 $layer=LI1_cond $X=7.245 $Y=2.475
+ $X2=7.227 $Y2=2.64
r186 39 56 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.245 $Y=0.845
+ $X2=7.245 $Y2=0.72
r187 39 40 106.342 $w=1.68e-07 $l=1.63e-06 $layer=LI1_cond $X=7.245 $Y=0.845
+ $X2=7.245 $Y2=2.475
r188 37 38 43.7534 $w=2.2e-07 $l=1.5e-07 $layer=POLY_cond $X=10.475 $Y=1.185
+ $X2=10.475 $Y2=1.335
r189 34 37 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=10.51 $Y=0.74
+ $X2=10.51 $Y2=1.185
r190 31 36 18.8402 $w=1.65e-07 $l=8.21584e-08 $layer=POLY_cond $X=10.44 $Y=1.555
+ $X2=10.425 $Y2=1.63
r191 31 38 112.809 $w=1.5e-07 $l=2.2e-07 $layer=POLY_cond $X=10.44 $Y=1.555
+ $X2=10.44 $Y2=1.335
r192 27 29 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=10.425 $Y=1.97
+ $X2=10.425 $Y2=2.465
r193 26 27 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=10.425 $Y=1.88
+ $X2=10.425 $Y2=1.97
r194 25 36 18.8402 $w=1.65e-07 $l=7.5e-08 $layer=POLY_cond $X=10.425 $Y=1.705
+ $X2=10.425 $Y2=1.63
r195 25 26 68.0242 $w=1.8e-07 $l=1.75e-07 $layer=POLY_cond $X=10.425 $Y=1.705
+ $X2=10.425 $Y2=1.88
r196 24 35 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=10.065 $Y=1.63
+ $X2=9.975 $Y2=1.63
r197 23 36 6.66866 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=10.335 $Y=1.63
+ $X2=10.425 $Y2=1.63
r198 23 24 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=10.335 $Y=1.63
+ $X2=10.065 $Y2=1.63
r199 20 22 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=9.975 $Y=1.97
+ $X2=9.975 $Y2=2.465
r200 19 20 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=9.975 $Y=1.88
+ $X2=9.975 $Y2=1.97
r201 18 35 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=9.975 $Y=1.705
+ $X2=9.975 $Y2=1.63
r202 18 19 68.0242 $w=1.8e-07 $l=1.75e-07 $layer=POLY_cond $X=9.975 $Y=1.705
+ $X2=9.975 $Y2=1.88
r203 17 65 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.675 $Y=1.63
+ $X2=9.51 $Y2=1.63
r204 16 35 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=9.885 $Y=1.63
+ $X2=9.975 $Y2=1.63
r205 16 17 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=9.885 $Y=1.63
+ $X2=9.675 $Y2=1.63
r206 13 15 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=9.47 $Y=2.39
+ $X2=9.47 $Y2=2.675
r207 12 13 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=9.47 $Y=2.3 $X2=9.47
+ $Y2=2.39
r208 12 66 231.282 $w=1.8e-07 $l=5.95e-07 $layer=POLY_cond $X=9.47 $Y=2.3
+ $X2=9.47 $Y2=1.705
r209 9 64 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=9.45 $Y=0.615
+ $X2=9.45 $Y2=1.375
r210 2 54 600 $w=1.7e-07 $l=8.93868e-07 $layer=licon1_PDIFF $count=1 $X=6.75
+ $Y=1.96 $X2=7.245 $Y2=2.64
r211 2 48 600 $w=1.7e-07 $l=1.38384e-06 $layer=licon1_PDIFF $count=1 $X=6.75
+ $Y=1.96 $X2=7.835 $Y2=2.64
r212 1 56 182 $w=1.7e-07 $l=3.73497e-07 $layer=licon1_NDIFF $count=1 $X=7.185
+ $Y=0.37 $X2=7.325 $Y2=0.68
r213 1 43 182 $w=1.7e-07 $l=7.23585e-07 $layer=licon1_NDIFF $count=1 $X=7.185
+ $Y=0.37 $X2=7.77 $Y2=0.68
.ends

.subckt PM_SKY130_FD_SC_HS__DFRTP_4%A_2010_409# 1 2 7 9 10 12 14 17 19 20 23 25
+ 27 30 32 34 37 39 43 45 46 49 56 59 67
c131 23 0 1.38275e-19 $X=12.025 $Y=0.74
r132 61 62 9.0375 $w=4e-07 $l=7.5e-08 $layer=POLY_cond $X=11.425 $Y=1.532
+ $X2=11.5 $Y2=1.532
r133 57 65 54.5473 $w=2.43e-07 $l=2.75e-07 $layer=POLY_cond $X=12.075 $Y=1.532
+ $X2=12.35 $Y2=1.532
r134 57 63 9.9177 $w=2.43e-07 $l=5e-08 $layer=POLY_cond $X=12.075 $Y=1.532
+ $X2=12.025 $Y2=1.532
r135 56 57 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=12.075
+ $Y=1.465 $X2=12.075 $Y2=1.465
r136 54 61 3.615 $w=4e-07 $l=3e-08 $layer=POLY_cond $X=11.395 $Y=1.532
+ $X2=11.425 $Y2=1.532
r137 53 56 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=11.395 $Y=1.465
+ $X2=12.075 $Y2=1.465
r138 53 54 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=11.395
+ $Y=1.465 $X2=11.395 $Y2=1.465
r139 51 59 6.46576 $w=2.5e-07 $l=1.65e-07 $layer=LI1_cond $X=10.89 $Y=1.465
+ $X2=10.725 $Y2=1.465
r140 51 53 17.6359 $w=3.28e-07 $l=5.05e-07 $layer=LI1_cond $X=10.89 $Y=1.465
+ $X2=11.395 $Y2=1.465
r141 47 59 0.364692 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=10.725 $Y=1.3
+ $X2=10.725 $Y2=1.465
r142 47 49 27.4142 $w=3.28e-07 $l=7.85e-07 $layer=LI1_cond $X=10.725 $Y=1.3
+ $X2=10.725 $Y2=0.515
r143 45 59 6.46576 $w=2.5e-07 $l=2.0106e-07 $layer=LI1_cond $X=10.56 $Y=1.545
+ $X2=10.725 $Y2=1.465
r144 45 46 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=10.56 $Y=1.545
+ $X2=10.365 $Y2=1.545
r145 41 46 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=10.24 $Y=1.63
+ $X2=10.365 $Y2=1.545
r146 41 43 25.8147 $w=2.48e-07 $l=5.6e-07 $layer=LI1_cond $X=10.24 $Y=1.63
+ $X2=10.24 $Y2=2.19
r147 35 67 30.7449 $w=2.43e-07 $l=1.55e-07 $layer=POLY_cond $X=12.955 $Y=1.532
+ $X2=12.8 $Y2=1.532
r148 35 37 379.447 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=12.955 $Y=1.48
+ $X2=12.955 $Y2=0.74
r149 32 67 14.0634 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=12.8 $Y=1.765
+ $X2=12.8 $Y2=1.532
r150 32 34 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=12.8 $Y=1.765
+ $X2=12.8 $Y2=2.4
r151 28 67 54.5473 $w=2.43e-07 $l=2.75e-07 $layer=POLY_cond $X=12.525 $Y=1.532
+ $X2=12.8 $Y2=1.532
r152 28 65 34.7119 $w=2.43e-07 $l=1.75e-07 $layer=POLY_cond $X=12.525 $Y=1.532
+ $X2=12.35 $Y2=1.532
r153 28 30 379.447 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=12.525 $Y=1.48
+ $X2=12.525 $Y2=0.74
r154 25 65 14.0634 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=12.35 $Y=1.765
+ $X2=12.35 $Y2=1.532
r155 25 27 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=12.35 $Y=1.765
+ $X2=12.35 $Y2=2.4
r156 21 63 14.0634 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=12.025 $Y=1.3
+ $X2=12.025 $Y2=1.532
r157 21 23 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=12.025 $Y=1.3
+ $X2=12.025 $Y2=0.74
r158 20 62 10.6563 $w=4e-07 $l=1.03199e-07 $layer=POLY_cond $X=11.575 $Y=1.465
+ $X2=11.5 $Y2=1.532
r159 19 63 14.4 $w=3.3e-07 $l=1.03199e-07 $layer=POLY_cond $X=11.95 $Y=1.465
+ $X2=12.025 $Y2=1.532
r160 19 20 65.573 $w=3.3e-07 $l=3.75e-07 $layer=POLY_cond $X=11.95 $Y=1.465
+ $X2=11.575 $Y2=1.465
r161 15 62 25.8619 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=11.5 $Y=1.3
+ $X2=11.5 $Y2=1.532
r162 15 17 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=11.5 $Y=1.3
+ $X2=11.5 $Y2=0.74
r163 12 61 25.8619 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=11.425 $Y=1.765
+ $X2=11.425 $Y2=1.532
r164 12 14 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=11.425 $Y=1.765
+ $X2=11.425 $Y2=2.4
r165 11 39 7.1379 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=11.02 $Y=1.555
+ $X2=10.93 $Y2=1.555
r166 10 54 39.5853 $w=4e-07 $l=1.76125e-07 $layer=POLY_cond $X=11.23 $Y=1.555
+ $X2=11.395 $Y2=1.532
r167 10 11 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=11.23 $Y=1.555
+ $X2=11.02 $Y2=1.555
r168 7 39 83.7788 $w=1.8e-07 $l=2.1e-07 $layer=POLY_cond $X=10.93 $Y=1.765
+ $X2=10.93 $Y2=1.555
r169 7 9 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=10.93 $Y=1.765
+ $X2=10.93 $Y2=2.4
r170 2 43 300 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=2 $X=10.05
+ $Y=2.045 $X2=10.2 $Y2=2.19
r171 1 49 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=10.585
+ $Y=0.37 $X2=10.725 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__DFRTP_4%VPWR 1 2 3 4 5 6 7 8 9 10 31 33 37 41 45 49
+ 53 57 61 65 67 69 74 75 77 78 80 81 82 84 89 94 102 120 124 133 136 139 142
+ 145 149
c165 149 0 2.33512e-20 $X=13.2 $Y=3.33
c166 102 0 1.50343e-19 $X=5.83 $Y=3.33
c167 61 0 1.07146e-19 $X=10.7 $Y=2.19
r168 148 149 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.2 $Y=3.33
+ $X2=13.2 $Y2=3.33
r169 145 146 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.76 $Y=3.33
+ $X2=11.76 $Y2=3.33
r170 142 143 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r171 139 140 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r172 136 137 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r173 133 134 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r174 130 131 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r175 128 149 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.72 $Y=3.33
+ $X2=13.2 $Y2=3.33
r176 128 146 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=12.72 $Y=3.33
+ $X2=11.76 $Y2=3.33
r177 127 128 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=12.72 $Y=3.33
+ $X2=12.72 $Y2=3.33
r178 125 145 13.7128 $w=1.7e-07 $l=3.53e-07 $layer=LI1_cond $X=12.24 $Y=3.33
+ $X2=11.887 $Y2=3.33
r179 125 127 31.3155 $w=1.68e-07 $l=4.8e-07 $layer=LI1_cond $X=12.24 $Y=3.33
+ $X2=12.72 $Y2=3.33
r180 124 148 4.57341 $w=1.7e-07 $l=2.65e-07 $layer=LI1_cond $X=12.91 $Y=3.33
+ $X2=13.175 $Y2=3.33
r181 124 127 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=12.91 $Y=3.33
+ $X2=12.72 $Y2=3.33
r182 123 146 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.28 $Y=3.33
+ $X2=11.76 $Y2=3.33
r183 122 123 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=11.28 $Y=3.33
+ $X2=11.28 $Y2=3.33
r184 120 145 13.7128 $w=1.7e-07 $l=3.52e-07 $layer=LI1_cond $X=11.535 $Y=3.33
+ $X2=11.887 $Y2=3.33
r185 120 122 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=11.535 $Y=3.33
+ $X2=11.28 $Y2=3.33
r186 119 123 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=10.32 $Y=3.33
+ $X2=11.28 $Y2=3.33
r187 118 119 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.32 $Y=3.33
+ $X2=10.32 $Y2=3.33
r188 116 119 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=9.36 $Y=3.33
+ $X2=10.32 $Y2=3.33
r189 115 116 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.36 $Y=3.33
+ $X2=9.36 $Y2=3.33
r190 113 116 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=8.4 $Y=3.33
+ $X2=9.36 $Y2=3.33
r191 112 113 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=8.4 $Y=3.33
+ $X2=8.4 $Y2=3.33
r192 110 143 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=6 $Y2=3.33
r193 109 112 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=6.48 $Y=3.33
+ $X2=8.4 $Y2=3.33
r194 109 110 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r195 107 142 8.70163 $w=1.7e-07 $l=1.68e-07 $layer=LI1_cond $X=6.165 $Y=3.33
+ $X2=5.997 $Y2=3.33
r196 107 109 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=6.165 $Y=3.33
+ $X2=6.48 $Y2=3.33
r197 106 143 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=6 $Y2=3.33
r198 106 140 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=4.56 $Y2=3.33
r199 105 106 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r200 103 139 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.73 $Y=3.33
+ $X2=4.565 $Y2=3.33
r201 103 105 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=4.73 $Y=3.33
+ $X2=5.52 $Y2=3.33
r202 102 142 8.70163 $w=1.7e-07 $l=1.67e-07 $layer=LI1_cond $X=5.83 $Y=3.33
+ $X2=5.997 $Y2=3.33
r203 102 105 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=5.83 $Y=3.33
+ $X2=5.52 $Y2=3.33
r204 101 140 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=4.56 $Y2=3.33
r205 100 101 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r206 98 101 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=4.08 $Y2=3.33
r207 98 137 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=2.16 $Y2=3.33
r208 97 100 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=2.64 $Y=3.33
+ $X2=4.08 $Y2=3.33
r209 97 98 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r210 95 136 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.335 $Y=3.33
+ $X2=2.17 $Y2=3.33
r211 95 97 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=2.335 $Y=3.33
+ $X2=2.64 $Y2=3.33
r212 94 139 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.4 $Y=3.33
+ $X2=4.565 $Y2=3.33
r213 94 100 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=4.4 $Y=3.33
+ $X2=4.08 $Y2=3.33
r214 93 137 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r215 93 134 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r216 92 93 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r217 90 133 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.34 $Y=3.33
+ $X2=1.215 $Y2=3.33
r218 90 92 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=1.34 $Y=3.33
+ $X2=1.68 $Y2=3.33
r219 89 136 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.005 $Y=3.33
+ $X2=2.17 $Y2=3.33
r220 89 92 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=2.005 $Y=3.33
+ $X2=1.68 $Y2=3.33
r221 88 134 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r222 88 131 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r223 87 88 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r224 85 130 4.01803 $w=1.7e-07 $l=1.8e-07 $layer=LI1_cond $X=0.36 $Y=3.33
+ $X2=0.18 $Y2=3.33
r225 85 87 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=0.36 $Y=3.33
+ $X2=0.72 $Y2=3.33
r226 84 133 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.09 $Y=3.33
+ $X2=1.215 $Y2=3.33
r227 84 87 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=1.09 $Y=3.33
+ $X2=0.72 $Y2=3.33
r228 82 113 0.468274 $w=4.9e-07 $l=1.68e-06 $layer=MET1_cond $X=6.72 $Y=3.33
+ $X2=8.4 $Y2=3.33
r229 82 110 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=6.72 $Y=3.33
+ $X2=6.48 $Y2=3.33
r230 80 118 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=10.535 $Y=3.33
+ $X2=10.32 $Y2=3.33
r231 80 81 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.535 $Y=3.33
+ $X2=10.7 $Y2=3.33
r232 79 122 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=10.865 $Y=3.33
+ $X2=11.28 $Y2=3.33
r233 79 81 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.865 $Y=3.33
+ $X2=10.7 $Y2=3.33
r234 77 115 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=9.65 $Y=3.33
+ $X2=9.36 $Y2=3.33
r235 77 78 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=9.65 $Y=3.33
+ $X2=9.775 $Y2=3.33
r236 76 118 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=9.9 $Y=3.33
+ $X2=10.32 $Y2=3.33
r237 76 78 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=9.9 $Y=3.33
+ $X2=9.775 $Y2=3.33
r238 74 112 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=8.58 $Y=3.33
+ $X2=8.4 $Y2=3.33
r239 74 75 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.58 $Y=3.33
+ $X2=8.745 $Y2=3.33
r240 73 115 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=8.91 $Y=3.33
+ $X2=9.36 $Y2=3.33
r241 73 75 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.91 $Y=3.33
+ $X2=8.745 $Y2=3.33
r242 69 72 24.4458 $w=3.28e-07 $l=7e-07 $layer=LI1_cond $X=13.075 $Y=2.115
+ $X2=13.075 $Y2=2.815
r243 67 148 3.19276 $w=3.3e-07 $l=1.36015e-07 $layer=LI1_cond $X=13.075 $Y=3.245
+ $X2=13.175 $Y2=3.33
r244 67 72 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=13.075 $Y=3.245
+ $X2=13.075 $Y2=2.815
r245 63 145 2.87722 $w=7.05e-07 $l=8.5e-08 $layer=LI1_cond $X=11.887 $Y=3.245
+ $X2=11.887 $Y2=3.33
r246 63 65 15.9477 $w=7.03e-07 $l=9.4e-07 $layer=LI1_cond $X=11.887 $Y=3.245
+ $X2=11.887 $Y2=2.305
r247 59 81 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=10.7 $Y=3.245
+ $X2=10.7 $Y2=3.33
r248 59 61 36.8433 $w=3.28e-07 $l=1.055e-06 $layer=LI1_cond $X=10.7 $Y=3.245
+ $X2=10.7 $Y2=2.19
r249 55 78 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=9.775 $Y=3.245
+ $X2=9.775 $Y2=3.33
r250 55 57 26.2757 $w=2.48e-07 $l=5.7e-07 $layer=LI1_cond $X=9.775 $Y=3.245
+ $X2=9.775 $Y2=2.675
r251 51 75 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.745 $Y=3.245
+ $X2=8.745 $Y2=3.33
r252 51 53 19.9058 $w=3.28e-07 $l=5.7e-07 $layer=LI1_cond $X=8.745 $Y=3.245
+ $X2=8.745 $Y2=2.675
r253 47 142 0.942324 $w=3.35e-07 $l=8.5e-08 $layer=LI1_cond $X=5.997 $Y=3.245
+ $X2=5.997 $Y2=3.33
r254 47 49 14.2765 $w=3.33e-07 $l=4.15e-07 $layer=LI1_cond $X=5.997 $Y=3.245
+ $X2=5.997 $Y2=2.83
r255 43 139 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.565 $Y=3.245
+ $X2=4.565 $Y2=3.33
r256 43 45 14.6675 $w=3.28e-07 $l=4.2e-07 $layer=LI1_cond $X=4.565 $Y=3.245
+ $X2=4.565 $Y2=2.825
r257 39 136 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.17 $Y=3.245
+ $X2=2.17 $Y2=3.33
r258 39 41 16.0644 $w=3.28e-07 $l=4.6e-07 $layer=LI1_cond $X=2.17 $Y=3.245
+ $X2=2.17 $Y2=2.785
r259 35 133 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.215 $Y=3.245
+ $X2=1.215 $Y2=3.33
r260 35 37 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=1.215 $Y=3.245
+ $X2=1.215 $Y2=2.815
r261 31 130 3.12513 $w=2.5e-07 $l=1.09087e-07 $layer=LI1_cond $X=0.235 $Y=3.245
+ $X2=0.18 $Y2=3.33
r262 31 33 22.8184 $w=2.48e-07 $l=4.95e-07 $layer=LI1_cond $X=0.235 $Y=3.245
+ $X2=0.235 $Y2=2.75
r263 10 72 400 $w=1.7e-07 $l=1.07034e-06 $layer=licon1_PDIFF $count=1 $X=12.875
+ $Y=1.84 $X2=13.075 $Y2=2.815
r264 10 69 400 $w=1.7e-07 $l=3.61421e-07 $layer=licon1_PDIFF $count=1 $X=12.875
+ $Y=1.84 $X2=13.075 $Y2=2.115
r265 9 65 150 $w=1.7e-07 $l=8.20183e-07 $layer=licon1_PDIFF $count=4 $X=11.5
+ $Y=1.84 $X2=12.12 $Y2=2.305
r266 8 61 300 $w=1.7e-07 $l=2.62678e-07 $layer=licon1_PDIFF $count=2 $X=10.5
+ $Y=2.045 $X2=10.7 $Y2=2.19
r267 7 57 600 $w=1.7e-07 $l=2.89828e-07 $layer=licon1_PDIFF $count=1 $X=9.545
+ $Y=2.465 $X2=9.735 $Y2=2.675
r268 6 53 600 $w=1.7e-07 $l=2.89828e-07 $layer=licon1_PDIFF $count=1 $X=8.555
+ $Y=2.465 $X2=8.745 $Y2=2.675
r269 5 49 600 $w=1.7e-07 $l=2.41402e-07 $layer=licon1_PDIFF $count=1 $X=5.81
+ $Y=2.7 $X2=5.995 $Y2=2.83
r270 4 45 600 $w=1.7e-07 $l=6.14329e-07 $layer=licon1_PDIFF $count=1 $X=4.335
+ $Y=2.315 $X2=4.565 $Y2=2.825
r271 3 41 600 $w=1.7e-07 $l=1.02727e-06 $layer=licon1_PDIFF $count=1 $X=2.02
+ $Y=1.83 $X2=2.17 $Y2=2.785
r272 2 37 600 $w=1.7e-07 $l=3.4187e-07 $layer=licon1_PDIFF $count=1 $X=1.025
+ $Y=2.54 $X2=1.175 $Y2=2.815
r273 1 33 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.54 $X2=0.275 $Y2=2.75
.ends

.subckt PM_SKY130_FD_SC_HS__DFRTP_4%A_37_78# 1 2 3 4 13 16 19 23 25 27 28 30 32
+ 36 39 40 41
c124 27 0 1.35567e-19 $X=3.625 $Y=1.305
r125 43 45 3.49225 $w=3.28e-07 $l=1e-07 $layer=LI1_cond $X=3.195 $Y=2.425
+ $X2=3.195 $Y2=2.525
r126 41 43 9.7783 $w=3.28e-07 $l=2.8e-07 $layer=LI1_cond $X=3.195 $Y=2.145
+ $X2=3.195 $Y2=2.425
r127 39 40 9.42727 $w=1.98e-07 $l=1.7e-07 $layer=LI1_cond $X=1.51 $Y=2.41
+ $X2=1.68 $Y2=2.41
r128 36 38 14.9345 $w=2.9e-07 $l=3.55e-07 $layer=LI1_cond $X=0.725 $Y=2.395
+ $X2=0.725 $Y2=2.75
r129 32 34 5.06376 $w=3.28e-07 $l=1.45e-07 $layer=LI1_cond $X=0.33 $Y=0.6
+ $X2=0.33 $Y2=0.745
r130 29 30 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.71 $Y=1.39
+ $X2=3.71 $Y2=2.06
r131 27 29 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.625 $Y=1.305
+ $X2=3.71 $Y2=1.39
r132 27 28 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=3.625 $Y=1.305
+ $X2=3.435 $Y2=1.305
r133 26 41 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.36 $Y=2.145
+ $X2=3.195 $Y2=2.145
r134 25 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.625 $Y=2.145
+ $X2=3.71 $Y2=2.06
r135 25 26 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=3.625 $Y=2.145
+ $X2=3.36 $Y2=2.145
r136 21 28 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=3.31 $Y=1.22
+ $X2=3.435 $Y2=1.305
r137 21 23 14.7513 $w=2.48e-07 $l=3.2e-07 $layer=LI1_cond $X=3.31 $Y=1.22
+ $X2=3.31 $Y2=0.9
r138 19 43 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.03 $Y=2.425
+ $X2=3.195 $Y2=2.425
r139 19 40 88.0749 $w=1.68e-07 $l=1.35e-06 $layer=LI1_cond $X=3.03 $Y=2.425
+ $X2=1.68 $Y2=2.425
r140 18 36 3.86198 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.89 $Y=2.395
+ $X2=0.725 $Y2=2.395
r141 18 39 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=0.89 $Y=2.395
+ $X2=1.51 $Y2=2.395
r142 16 36 5.64745 $w=2.9e-07 $l=1.05119e-07 $layer=LI1_cond $X=0.77 $Y=2.31
+ $X2=0.725 $Y2=2.395
r143 15 16 96.5562 $w=1.68e-07 $l=1.48e-06 $layer=LI1_cond $X=0.77 $Y=0.83
+ $X2=0.77 $Y2=2.31
r144 14 34 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.495 $Y=0.745
+ $X2=0.33 $Y2=0.745
r145 13 15 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.685 $Y=0.745
+ $X2=0.77 $Y2=0.83
r146 13 14 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=0.685 $Y=0.745
+ $X2=0.495 $Y2=0.745
r147 4 45 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=3.055
+ $Y=2.315 $X2=3.195 $Y2=2.525
r148 3 38 600 $w=1.7e-07 $l=2.74955e-07 $layer=licon1_PDIFF $count=1 $X=0.575
+ $Y=2.54 $X2=0.725 $Y2=2.75
r149 2 23 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=3.125
+ $Y=0.69 $X2=3.27 $Y2=0.9
r150 1 32 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=0.185
+ $Y=0.39 $X2=0.33 $Y2=0.6
.ends

.subckt PM_SKY130_FD_SC_HS__DFRTP_4%Q 1 2 3 4 15 19 20 21 23 25 29 35 38 41 42
c73 42 0 1.38275e-19 $X=13.2 $Y=1.665
r74 44 45 2.94971 $w=5.17e-07 $l=1.25e-07 $layer=LI1_cond $X=12.575 $Y=1.62
+ $X2=12.7 $Y2=1.62
r75 42 45 11.7988 $w=5.17e-07 $l=5e-07 $layer=LI1_cond $X=13.2 $Y=1.62 $X2=12.7
+ $Y2=1.62
r76 38 45 5.00057 $w=2.5e-07 $l=3.5e-07 $layer=LI1_cond $X=12.7 $Y=1.27 $X2=12.7
+ $Y2=1.62
r77 37 41 5.16603 $w=2.5e-07 $l=1.25e-07 $layer=LI1_cond $X=12.7 $Y=1.13
+ $X2=12.7 $Y2=1.005
r78 37 38 6.45368 $w=2.48e-07 $l=1.4e-07 $layer=LI1_cond $X=12.7 $Y=1.13
+ $X2=12.7 $Y2=1.27
r79 33 41 5.16603 $w=2.5e-07 $l=1.25e-07 $layer=LI1_cond $X=12.7 $Y=0.88
+ $X2=12.7 $Y2=1.005
r80 33 35 16.8257 $w=2.48e-07 $l=3.65e-07 $layer=LI1_cond $X=12.7 $Y=0.88
+ $X2=12.7 $Y2=0.515
r81 29 31 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=12.575 $Y=1.985
+ $X2=12.575 $Y2=2.815
r82 27 44 3.36414 $w=3.3e-07 $l=3.5e-07 $layer=LI1_cond $X=12.575 $Y=1.97
+ $X2=12.575 $Y2=1.62
r83 27 29 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=12.575 $Y=1.97
+ $X2=12.575 $Y2=1.985
r84 26 40 3.87155 $w=2.5e-07 $l=1.58e-07 $layer=LI1_cond $X=11.91 $Y=1.005
+ $X2=11.752 $Y2=1.005
r85 25 41 1.34256 $w=2.5e-07 $l=1.25e-07 $layer=LI1_cond $X=12.575 $Y=1.005
+ $X2=12.7 $Y2=1.005
r86 25 26 30.655 $w=2.48e-07 $l=6.65e-07 $layer=LI1_cond $X=12.575 $Y=1.005
+ $X2=11.91 $Y2=1.005
r87 21 40 3.06294 $w=3.15e-07 $l=1.25e-07 $layer=LI1_cond $X=11.752 $Y=0.88
+ $X2=11.752 $Y2=1.005
r88 21 23 12.8049 $w=3.13e-07 $l=3.5e-07 $layer=LI1_cond $X=11.752 $Y=0.88
+ $X2=11.752 $Y2=0.53
r89 19 44 9.81494 $w=5.17e-07 $l=3.37565e-07 $layer=LI1_cond $X=12.41 $Y=1.885
+ $X2=12.575 $Y2=1.62
r90 19 20 68.1765 $w=1.68e-07 $l=1.045e-06 $layer=LI1_cond $X=12.41 $Y=1.885
+ $X2=11.365 $Y2=1.885
r91 15 17 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=11.2 $Y=1.985
+ $X2=11.2 $Y2=2.815
r92 13 20 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=11.2 $Y=1.97
+ $X2=11.365 $Y2=1.885
r93 13 15 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=11.2 $Y=1.97
+ $X2=11.2 $Y2=1.985
r94 4 31 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=12.425
+ $Y=1.84 $X2=12.575 $Y2=2.815
r95 4 29 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=12.425
+ $Y=1.84 $X2=12.575 $Y2=1.985
r96 3 17 400 $w=1.7e-07 $l=1.06806e-06 $layer=licon1_PDIFF $count=1 $X=11.005
+ $Y=1.84 $X2=11.2 $Y2=2.815
r97 3 15 400 $w=1.7e-07 $l=2.57488e-07 $layer=licon1_PDIFF $count=1 $X=11.005
+ $Y=1.84 $X2=11.2 $Y2=1.985
r98 2 35 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=12.6
+ $Y=0.37 $X2=12.74 $Y2=0.515
r99 1 40 182 $w=1.7e-07 $l=6.81249e-07 $layer=licon1_NDIFF $count=1 $X=11.575
+ $Y=0.37 $X2=11.76 $Y2=0.965
r100 1 23 182 $w=1.7e-07 $l=2.52636e-07 $layer=licon1_NDIFF $count=1 $X=11.575
+ $Y=0.37 $X2=11.76 $Y2=0.53
.ends

.subckt PM_SKY130_FD_SC_HS__DFRTP_4%VGND 1 2 3 4 5 6 7 8 27 31 35 39 43 47 49 51
+ 54 55 57 58 59 65 69 77 89 93 98 104 108 114 117 120 124
c138 124 0 3.01223e-20 $X=13.2 $Y=0
r139 123 124 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.2 $Y=0
+ $X2=13.2 $Y2=0
r140 120 121 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.24 $Y=0
+ $X2=12.24 $Y2=0
r141 117 118 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.28 $Y=0
+ $X2=11.28 $Y2=0
r142 114 115 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=8.88 $Y=0
+ $X2=8.88 $Y2=0
r143 108 111 9.95292 $w=3.28e-07 $l=2.85e-07 $layer=LI1_cond $X=5.06 $Y=0
+ $X2=5.06 $Y2=0.285
r144 108 109 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=0
+ $X2=5.04 $Y2=0
r145 104 105 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0
+ $X2=2.16 $Y2=0
r146 102 124 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.72 $Y=0
+ $X2=13.2 $Y2=0
r147 102 121 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.72 $Y=0
+ $X2=12.24 $Y2=0
r148 101 102 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.72 $Y=0
+ $X2=12.72 $Y2=0
r149 99 120 8.5188 $w=1.7e-07 $l=1.63e-07 $layer=LI1_cond $X=12.405 $Y=0
+ $X2=12.242 $Y2=0
r150 99 101 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=12.405 $Y=0
+ $X2=12.72 $Y2=0
r151 98 123 4.76062 $w=1.7e-07 $l=2.17e-07 $layer=LI1_cond $X=13.005 $Y=0
+ $X2=13.222 $Y2=0
r152 98 101 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=13.005 $Y=0
+ $X2=12.72 $Y2=0
r153 97 121 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.76 $Y=0
+ $X2=12.24 $Y2=0
r154 97 118 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.76 $Y=0
+ $X2=11.28 $Y2=0
r155 96 97 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.76 $Y=0
+ $X2=11.76 $Y2=0
r156 94 117 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=11.41 $Y=0
+ $X2=11.265 $Y2=0
r157 94 96 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=11.41 $Y=0
+ $X2=11.76 $Y2=0
r158 93 120 8.5188 $w=1.7e-07 $l=1.62e-07 $layer=LI1_cond $X=12.08 $Y=0
+ $X2=12.242 $Y2=0
r159 93 96 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=12.08 $Y=0 $X2=11.76
+ $Y2=0
r160 92 118 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.8 $Y=0
+ $X2=11.28 $Y2=0
r161 91 92 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.8 $Y=0 $X2=10.8
+ $Y2=0
r162 89 117 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=11.12 $Y=0
+ $X2=11.265 $Y2=0
r163 89 91 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=11.12 $Y=0 $X2=10.8
+ $Y2=0
r164 88 92 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=9.84 $Y=0 $X2=10.8
+ $Y2=0
r165 88 115 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=9.84 $Y=0
+ $X2=8.88 $Y2=0
r166 87 88 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=9.84 $Y=0 $X2=9.84
+ $Y2=0
r167 85 114 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.955 $Y=0
+ $X2=8.79 $Y2=0
r168 85 87 57.738 $w=1.68e-07 $l=8.85e-07 $layer=LI1_cond $X=8.955 $Y=0 $X2=9.84
+ $Y2=0
r169 84 115 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=0 $X2=8.88
+ $Y2=0
r170 83 84 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=8.4 $Y=0
+ $X2=8.4 $Y2=0
r171 81 109 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=0
+ $X2=5.04 $Y2=0
r172 80 83 187.893 $w=1.68e-07 $l=2.88e-06 $layer=LI1_cond $X=5.52 $Y=0 $X2=8.4
+ $Y2=0
r173 80 81 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=5.52 $Y=0
+ $X2=5.52 $Y2=0
r174 78 108 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.225 $Y=0
+ $X2=5.06 $Y2=0
r175 78 80 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=5.225 $Y=0 $X2=5.52
+ $Y2=0
r176 77 114 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.625 $Y=0
+ $X2=8.79 $Y2=0
r177 77 83 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=8.625 $Y=0 $X2=8.4
+ $Y2=0
r178 76 109 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0
+ $X2=5.04 $Y2=0
r179 75 76 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.56 $Y=0
+ $X2=4.56 $Y2=0
r180 73 76 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=2.64 $Y=0
+ $X2=4.56 $Y2=0
r181 73 105 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0
+ $X2=2.16 $Y2=0
r182 72 75 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=2.64 $Y=0 $X2=4.56
+ $Y2=0
r183 72 73 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.64 $Y=0
+ $X2=2.64 $Y2=0
r184 70 104 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.375 $Y=0
+ $X2=2.21 $Y2=0
r185 70 72 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=2.375 $Y=0
+ $X2=2.64 $Y2=0
r186 69 108 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.895 $Y=0
+ $X2=5.06 $Y2=0
r187 69 75 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=4.895 $Y=0
+ $X2=4.56 $Y2=0
r188 68 105 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0
+ $X2=2.16 $Y2=0
r189 67 68 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r190 65 104 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.045 $Y=0
+ $X2=2.21 $Y2=0
r191 65 67 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=2.045 $Y=0
+ $X2=1.68 $Y2=0
r192 63 68 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r193 62 63 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r194 59 84 0.468274 $w=4.9e-07 $l=1.68e-06 $layer=MET1_cond $X=6.72 $Y=0 $X2=8.4
+ $Y2=0
r195 59 81 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=6.72 $Y=0 $X2=5.52
+ $Y2=0
r196 57 87 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=10.115 $Y=0
+ $X2=9.84 $Y2=0
r197 57 58 7.54988 $w=1.7e-07 $l=1.37e-07 $layer=LI1_cond $X=10.115 $Y=0
+ $X2=10.252 $Y2=0
r198 56 91 26.7487 $w=1.68e-07 $l=4.1e-07 $layer=LI1_cond $X=10.39 $Y=0 $X2=10.8
+ $Y2=0
r199 56 58 7.54988 $w=1.7e-07 $l=1.38e-07 $layer=LI1_cond $X=10.39 $Y=0
+ $X2=10.252 $Y2=0
r200 54 62 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.065 $Y=0 $X2=0.72
+ $Y2=0
r201 54 55 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.065 $Y=0 $X2=1.15
+ $Y2=0
r202 53 67 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=1.235 $Y=0
+ $X2=1.68 $Y2=0
r203 53 55 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.235 $Y=0 $X2=1.15
+ $Y2=0
r204 49 123 3.00555 $w=3.3e-07 $l=1.07912e-07 $layer=LI1_cond $X=13.17 $Y=0.085
+ $X2=13.222 $Y2=0
r205 49 51 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=13.17 $Y=0.085
+ $X2=13.17 $Y2=0.515
r206 45 120 0.848899 $w=3.25e-07 $l=8.5e-08 $layer=LI1_cond $X=12.242 $Y=0.085
+ $X2=12.242 $Y2=0
r207 45 47 15.7796 $w=3.23e-07 $l=4.45e-07 $layer=LI1_cond $X=12.242 $Y=0.085
+ $X2=12.242 $Y2=0.53
r208 41 117 0.489042 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=11.265 $Y=0.085
+ $X2=11.265 $Y2=0
r209 41 43 17.684 $w=2.88e-07 $l=4.45e-07 $layer=LI1_cond $X=11.265 $Y=0.085
+ $X2=11.265 $Y2=0.53
r210 37 58 0.316938 $w=2.75e-07 $l=8.5e-08 $layer=LI1_cond $X=10.252 $Y=0.085
+ $X2=10.252 $Y2=0
r211 37 39 18.02 $w=2.73e-07 $l=4.3e-07 $layer=LI1_cond $X=10.252 $Y=0.085
+ $X2=10.252 $Y2=0.515
r212 33 114 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.79 $Y=0.085
+ $X2=8.79 $Y2=0
r213 33 35 18.5089 $w=3.28e-07 $l=5.3e-07 $layer=LI1_cond $X=8.79 $Y=0.085
+ $X2=8.79 $Y2=0.615
r214 29 104 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.21 $Y=0.085
+ $X2=2.21 $Y2=0
r215 29 31 17.112 $w=3.28e-07 $l=4.9e-07 $layer=LI1_cond $X=2.21 $Y=0.085
+ $X2=2.21 $Y2=0.575
r216 25 55 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.15 $Y=0.085
+ $X2=1.15 $Y2=0
r217 25 27 33.5989 $w=1.68e-07 $l=5.15e-07 $layer=LI1_cond $X=1.15 $Y=0.085
+ $X2=1.15 $Y2=0.6
r218 8 51 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=13.03
+ $Y=0.37 $X2=13.17 $Y2=0.515
r219 7 47 182 $w=1.7e-07 $l=2.19089e-07 $layer=licon1_NDIFF $count=1 $X=12.1
+ $Y=0.37 $X2=12.24 $Y2=0.53
r220 6 43 91 $w=1.7e-07 $l=2.20907e-07 $layer=licon1_NDIFF $count=2 $X=11.14
+ $Y=0.37 $X2=11.285 $Y2=0.53
r221 5 39 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=10.08
+ $Y=0.37 $X2=10.225 $Y2=0.515
r222 4 35 182 $w=1.7e-07 $l=2.80624e-07 $layer=licon1_NDIFF $count=1 $X=8.625
+ $Y=0.405 $X2=8.79 $Y2=0.615
r223 3 111 182 $w=1.7e-07 $l=5.03115e-07 $layer=licon1_NDIFF $count=1 $X=4.84
+ $Y=0.69 $X2=5.06 $Y2=0.285
r224 2 31 182 $w=1.7e-07 $l=2.95212e-07 $layer=licon1_NDIFF $count=1 $X=2
+ $Y=0.37 $X2=2.21 $Y2=0.575
r225 1 27 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.01
+ $Y=0.39 $X2=1.15 $Y2=0.6
.ends

