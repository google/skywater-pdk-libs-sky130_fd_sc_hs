* File: sky130_fd_sc_hs__o2bb2a_4.pex.spice
* Created: Tue Sep  1 20:16:53 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HS__O2BB2A_4%B1 3 6 7 9 11 12 14 17 19 20 30 31
c58 12 0 4.75553e-20 $X=1.025 $Y=1.885
c59 11 0 5.33865e-20 $X=1.025 $Y=1.795
c60 3 0 1.72779e-19 $X=0.495 $Y=0.69
r61 31 32 5.93231 $w=3.25e-07 $l=4e-08 $layer=POLY_cond $X=1.025 $Y=1.425
+ $X2=1.065 $Y2=1.425
r62 29 31 11.1231 $w=3.25e-07 $l=7.5e-08 $layer=POLY_cond $X=0.95 $Y=1.425
+ $X2=1.025 $Y2=1.425
r63 29 30 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.95
+ $Y=1.425 $X2=0.95 $Y2=1.425
r64 27 29 55.6154 $w=3.25e-07 $l=3.75e-07 $layer=POLY_cond $X=0.575 $Y=1.425
+ $X2=0.95 $Y2=1.425
r65 26 27 11.8646 $w=3.25e-07 $l=8e-08 $layer=POLY_cond $X=0.495 $Y=1.425
+ $X2=0.575 $Y2=1.425
r66 24 26 33.3692 $w=3.25e-07 $l=2.25e-07 $layer=POLY_cond $X=0.27 $Y=1.425
+ $X2=0.495 $Y2=1.425
r67 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.27
+ $Y=1.425 $X2=0.27 $Y2=1.425
r68 20 30 5.39408 $w=5.08e-07 $l=2.3e-07 $layer=LI1_cond $X=0.72 $Y=1.515
+ $X2=0.95 $Y2=1.515
r69 20 25 10.5536 $w=5.08e-07 $l=4.5e-07 $layer=LI1_cond $X=0.72 $Y=1.515
+ $X2=0.27 $Y2=1.515
r70 19 25 0.703576 $w=5.08e-07 $l=3e-08 $layer=LI1_cond $X=0.24 $Y=1.515
+ $X2=0.27 $Y2=1.515
r71 15 32 20.86 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.065 $Y=1.26
+ $X2=1.065 $Y2=1.425
r72 15 17 292.277 $w=1.5e-07 $l=5.7e-07 $layer=POLY_cond $X=1.065 $Y=1.26
+ $X2=1.065 $Y2=0.69
r73 12 14 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=1.025 $Y=1.885
+ $X2=1.025 $Y2=2.46
r74 11 12 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=1.025 $Y=1.795
+ $X2=1.025 $Y2=1.885
r75 10 31 16.5763 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.025 $Y=1.59
+ $X2=1.025 $Y2=1.425
r76 10 11 79.6855 $w=1.8e-07 $l=2.05e-07 $layer=POLY_cond $X=1.025 $Y=1.59
+ $X2=1.025 $Y2=1.795
r77 7 9 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=0.575 $Y=1.885
+ $X2=0.575 $Y2=2.46
r78 6 7 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=0.575 $Y=1.795 $X2=0.575
+ $Y2=1.885
r79 5 27 16.5763 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=0.575 $Y=1.59
+ $X2=0.575 $Y2=1.425
r80 5 6 79.6855 $w=1.8e-07 $l=2.05e-07 $layer=POLY_cond $X=0.575 $Y=1.59
+ $X2=0.575 $Y2=1.795
r81 1 26 20.86 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.495 $Y=1.26
+ $X2=0.495 $Y2=1.425
r82 1 3 292.277 $w=1.5e-07 $l=5.7e-07 $layer=POLY_cond $X=0.495 $Y=1.26
+ $X2=0.495 $Y2=0.69
.ends

.subckt PM_SKY130_FD_SC_HS__O2BB2A_4%B2 1 3 6 8 10 13 15 16 23
c58 23 0 3.43014e-19 $X=1.975 $Y=1.615
c59 16 0 5.33865e-20 $X=2.16 $Y=1.665
c60 8 0 5.37684e-20 $X=1.925 $Y=1.885
r61 23 25 2.53684 $w=3.8e-07 $l=2e-08 $layer=POLY_cond $X=1.975 $Y=1.667
+ $X2=1.995 $Y2=1.667
r62 23 24 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.975
+ $Y=1.615 $X2=1.975 $Y2=1.615
r63 21 23 6.34211 $w=3.8e-07 $l=5e-08 $layer=POLY_cond $X=1.925 $Y=1.667
+ $X2=1.975 $Y2=1.667
r64 20 21 54.5421 $w=3.8e-07 $l=4.3e-07 $layer=POLY_cond $X=1.495 $Y=1.667
+ $X2=1.925 $Y2=1.667
r65 19 20 2.53684 $w=3.8e-07 $l=2e-08 $layer=POLY_cond $X=1.475 $Y=1.667
+ $X2=1.495 $Y2=1.667
r66 16 24 6.46067 $w=3.28e-07 $l=1.85e-07 $layer=LI1_cond $X=2.16 $Y=1.615
+ $X2=1.975 $Y2=1.615
r67 15 24 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=1.68 $Y=1.615
+ $X2=1.975 $Y2=1.615
r68 11 25 24.6126 $w=1.5e-07 $l=2.17e-07 $layer=POLY_cond $X=1.995 $Y=1.45
+ $X2=1.995 $Y2=1.667
r69 11 13 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=1.995 $Y=1.45
+ $X2=1.995 $Y2=0.69
r70 8 21 24.6126 $w=1.5e-07 $l=2.18e-07 $layer=POLY_cond $X=1.925 $Y=1.885
+ $X2=1.925 $Y2=1.667
r71 8 10 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=1.925 $Y=1.885
+ $X2=1.925 $Y2=2.46
r72 4 20 24.6126 $w=1.5e-07 $l=2.17e-07 $layer=POLY_cond $X=1.495 $Y=1.45
+ $X2=1.495 $Y2=1.667
r73 4 6 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=1.495 $Y=1.45
+ $X2=1.495 $Y2=0.69
r74 1 19 24.6126 $w=1.5e-07 $l=2.18e-07 $layer=POLY_cond $X=1.475 $Y=1.885
+ $X2=1.475 $Y2=1.667
r75 1 3 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=1.475 $Y=1.885
+ $X2=1.475 $Y2=2.46
.ends

.subckt PM_SKY130_FD_SC_HS__O2BB2A_4%A_476_48# 1 2 9 13 15 17 18 20 21 22 30 31
+ 33 34 36 41 42
c83 33 0 1.74227e-19 $X=3.59 $Y=1.95
c84 22 0 1.82144e-19 $X=3.505 $Y=1.465
c85 15 0 1.6087e-19 $X=2.935 $Y=1.765
c86 9 0 7.85372e-20 $X=2.455 $Y=0.69
r87 46 47 2.15179 $w=3.36e-07 $l=1.5e-08 $layer=POLY_cond $X=2.92 $Y=1.532
+ $X2=2.935 $Y2=1.532
r88 42 47 12.9107 $w=3.36e-07 $l=1.1887e-07 $layer=POLY_cond $X=3.025 $Y=1.465
+ $X2=2.935 $Y2=1.532
r89 34 36 21.8266 $w=3.28e-07 $l=6.25e-07 $layer=LI1_cond $X=3.675 $Y=2.115
+ $X2=4.3 $Y2=2.115
r90 33 34 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.59 $Y=1.95
+ $X2=3.675 $Y2=2.115
r91 32 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.59 $Y=1.63
+ $X2=3.59 $Y2=1.465
r92 32 33 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=3.59 $Y=1.63 $X2=3.59
+ $Y2=1.95
r93 31 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.59 $Y=1.3 $X2=3.59
+ $Y2=1.465
r94 30 40 9.62299 $w=3.74e-07 $l=4.00231e-07 $layer=LI1_cond $X=3.59 $Y=1.13
+ $X2=3.885 $Y2=0.882
r95 30 31 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=3.59 $Y=1.13
+ $X2=3.59 $Y2=1.3
r96 29 42 56.8299 $w=3.3e-07 $l=3.25e-07 $layer=POLY_cond $X=3.35 $Y=1.465
+ $X2=3.025 $Y2=1.465
r97 28 29 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=3.35
+ $Y=1.465 $X2=3.35 $Y2=1.465
r98 25 46 38.0149 $w=3.36e-07 $l=2.65e-07 $layer=POLY_cond $X=2.655 $Y=1.532
+ $X2=2.92 $Y2=1.532
r99 24 28 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=2.655 $Y=1.465
+ $X2=3.35 $Y2=1.465
r100 24 25 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=2.655
+ $Y=1.465 $X2=2.655 $Y2=1.465
r101 22 41 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.505 $Y=1.465
+ $X2=3.59 $Y2=1.465
r102 22 28 5.41299 $w=3.28e-07 $l=1.55e-07 $layer=LI1_cond $X=3.505 $Y=1.465
+ $X2=3.35 $Y2=1.465
r103 21 29 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=3.365 $Y=1.465
+ $X2=3.35 $Y2=1.465
r104 18 21 12.2053 $w=6.32e-07 $l=3.42053e-07 $layer=POLY_cond $X=3.455 $Y=1.765
+ $X2=3.365 $Y2=1.465
r105 18 20 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=3.455 $Y=1.765
+ $X2=3.455 $Y2=2.26
r106 15 47 21.6522 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=2.935 $Y=1.765
+ $X2=2.935 $Y2=1.532
r107 15 17 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=2.935 $Y=1.765
+ $X2=2.935 $Y2=2.26
r108 11 46 21.6522 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=2.92 $Y=1.3
+ $X2=2.92 $Y2=1.532
r109 11 13 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.92 $Y=1.3
+ $X2=2.92 $Y2=0.69
r110 7 25 28.6905 $w=3.36e-07 $l=3.16582e-07 $layer=POLY_cond $X=2.455 $Y=1.3
+ $X2=2.655 $Y2=1.532
r111 7 9 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.455 $Y=1.3
+ $X2=2.455 $Y2=0.69
r112 2 36 600 $w=1.7e-07 $l=3.4187e-07 $layer=licon1_PDIFF $count=1 $X=4.15
+ $Y=1.84 $X2=4.3 $Y2=2.115
r113 1 40 182 $w=1.7e-07 $l=4.04166e-07 $layer=licon1_NDIFF $count=1 $X=3.72
+ $Y=0.47 $X2=3.885 $Y2=0.8
.ends

.subckt PM_SKY130_FD_SC_HS__O2BB2A_4%A2_N 1 3 6 8 12
c34 6 0 1.762e-19 $X=4.1 $Y=0.79
r35 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.01
+ $Y=1.515 $X2=4.01 $Y2=1.515
r36 8 12 4.93904 $w=3.48e-07 $l=1.5e-07 $layer=LI1_cond $X=4.02 $Y=1.665
+ $X2=4.02 $Y2=1.515
r37 4 11 38.5562 $w=2.99e-07 $l=2.05122e-07 $layer=POLY_cond $X=4.1 $Y=1.35
+ $X2=4.01 $Y2=1.515
r38 4 6 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=4.1 $Y=1.35 $X2=4.1
+ $Y2=0.79
r39 1 11 52.2586 $w=2.99e-07 $l=2.80624e-07 $layer=POLY_cond $X=4.075 $Y=1.765
+ $X2=4.01 $Y2=1.515
r40 1 3 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=4.075 $Y=1.765
+ $X2=4.075 $Y2=2.26
.ends

.subckt PM_SKY130_FD_SC_HS__O2BB2A_4%A1_N 3 5 7 8 12
c34 12 0 4.1037e-20 $X=4.58 $Y=1.515
r35 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.58
+ $Y=1.515 $X2=4.58 $Y2=1.515
r36 8 12 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=4.58 $Y=1.665
+ $X2=4.58 $Y2=1.515
r37 5 11 52.2586 $w=2.99e-07 $l=2.76134e-07 $layer=POLY_cond $X=4.525 $Y=1.765
+ $X2=4.58 $Y2=1.515
r38 5 7 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=4.525 $Y=1.765
+ $X2=4.525 $Y2=2.26
r39 1 11 38.5562 $w=2.99e-07 $l=2.05122e-07 $layer=POLY_cond $X=4.49 $Y=1.35
+ $X2=4.58 $Y2=1.515
r40 1 3 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=4.49 $Y=1.35 $X2=4.49
+ $Y2=0.79
.ends

.subckt PM_SKY130_FD_SC_HS__O2BB2A_4%A_310_392# 1 2 3 12 13 15 16 18 20 21 23 24
+ 26 27 29 30 31 32 34 36 37 39 40 45 48 49 50 52 53 54 56 60 62 66 67 74 75 77
+ 81
c182 54 0 2.65681e-20 $X=4.37 $Y=1.035
c183 45 0 7.85372e-20 $X=4.2 $Y=0.34
c184 13 0 4.1037e-20 $X=5.145 $Y=1.765
r185 85 86 1.08804 $w=4.43e-07 $l=1e-08 $layer=POLY_cond $X=6.195 $Y=1.492
+ $X2=6.205 $Y2=1.492
r186 82 83 1.08804 $w=4.43e-07 $l=1e-08 $layer=POLY_cond $X=5.695 $Y=1.492
+ $X2=5.705 $Y2=1.492
r187 73 75 2.96841 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=3.165 $Y=1.985
+ $X2=3.25 $Y2=1.985
r188 73 74 8.63679 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=3.165 $Y=1.985
+ $X2=2.995 $Y2=1.985
r189 67 70 6.28605 $w=3.28e-07 $l=1.8e-07 $layer=LI1_cond $X=2.67 $Y=0.34
+ $X2=2.67 $Y2=0.52
r190 63 85 32.0971 $w=4.43e-07 $l=2.95e-07 $layer=POLY_cond $X=5.9 $Y=1.492
+ $X2=6.195 $Y2=1.492
r191 63 83 21.2167 $w=4.43e-07 $l=1.95e-07 $layer=POLY_cond $X=5.9 $Y=1.492
+ $X2=5.705 $Y2=1.492
r192 62 63 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=5.9
+ $Y=1.385 $X2=5.9 $Y2=1.385
r193 60 81 66.2869 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=5.145 $Y=1.385
+ $X2=5.145 $Y2=1.22
r194 59 62 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=5.22 $Y=1.385
+ $X2=5.9 $Y2=1.385
r195 59 60 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=5.22
+ $Y=1.385 $X2=5.22 $Y2=1.385
r196 57 77 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=5 $Y=1.385 $X2=5
+ $Y2=1.035
r197 57 59 4.71454 $w=3.28e-07 $l=1.35e-07 $layer=LI1_cond $X=5.085 $Y=1.385
+ $X2=5.22 $Y2=1.385
r198 55 57 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=5 $Y=1.55 $X2=5
+ $Y2=1.385
r199 55 56 58.7166 $w=1.68e-07 $l=9e-07 $layer=LI1_cond $X=5 $Y=1.55 $X2=5
+ $Y2=2.45
r200 53 77 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.915 $Y=1.035
+ $X2=5 $Y2=1.035
r201 53 54 35.5561 $w=1.68e-07 $l=5.45e-07 $layer=LI1_cond $X=4.915 $Y=1.035
+ $X2=4.37 $Y2=1.035
r202 52 54 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.285 $Y=0.95
+ $X2=4.37 $Y2=1.035
r203 51 52 34.2513 $w=1.68e-07 $l=5.25e-07 $layer=LI1_cond $X=4.285 $Y=0.425
+ $X2=4.285 $Y2=0.95
r204 49 56 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.915 $Y=2.535
+ $X2=5 $Y2=2.45
r205 49 50 103.08 $w=1.68e-07 $l=1.58e-06 $layer=LI1_cond $X=4.915 $Y=2.535
+ $X2=3.335 $Y2=2.535
r206 48 50 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.25 $Y=2.45
+ $X2=3.335 $Y2=2.535
r207 47 75 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.25 $Y=2.15
+ $X2=3.25 $Y2=1.985
r208 47 48 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=3.25 $Y=2.15 $X2=3.25
+ $Y2=2.45
r209 46 67 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.835 $Y=0.34
+ $X2=2.67 $Y2=0.34
r210 45 51 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.2 $Y=0.34
+ $X2=4.285 $Y2=0.425
r211 45 46 89.0535 $w=1.68e-07 $l=1.365e-06 $layer=LI1_cond $X=4.2 $Y=0.34
+ $X2=2.835 $Y2=0.34
r212 44 66 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.785 $Y=2.035
+ $X2=1.7 $Y2=2.035
r213 44 74 78.9412 $w=1.68e-07 $l=1.21e-06 $layer=LI1_cond $X=1.785 $Y=2.035
+ $X2=2.995 $Y2=2.035
r214 37 39 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=6.65 $Y=1.765
+ $X2=6.65 $Y2=2.4
r215 36 37 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=6.65 $Y=1.675
+ $X2=6.65 $Y2=1.765
r216 35 40 18.8402 $w=1.65e-07 $l=7.5e-08 $layer=POLY_cond $X=6.65 $Y=1.37
+ $X2=6.65 $Y2=1.295
r217 35 36 118.556 $w=1.8e-07 $l=3.05e-07 $layer=POLY_cond $X=6.65 $Y=1.37
+ $X2=6.65 $Y2=1.675
r218 32 40 18.8402 $w=1.65e-07 $l=8.21584e-08 $layer=POLY_cond $X=6.635 $Y=1.22
+ $X2=6.65 $Y2=1.295
r219 32 34 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=6.635 $Y=1.22
+ $X2=6.635 $Y2=0.74
r220 31 86 31.2673 $w=4.43e-07 $l=2.336e-07 $layer=POLY_cond $X=6.285 $Y=1.295
+ $X2=6.205 $Y2=1.492
r221 30 40 6.66866 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=6.56 $Y=1.295
+ $X2=6.65 $Y2=1.295
r222 30 31 141.011 $w=1.5e-07 $l=2.75e-07 $layer=POLY_cond $X=6.56 $Y=1.295
+ $X2=6.285 $Y2=1.295
r223 27 86 28.3771 $w=1.5e-07 $l=2.72e-07 $layer=POLY_cond $X=6.205 $Y=1.22
+ $X2=6.205 $Y2=1.492
r224 27 29 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=6.205 $Y=1.22
+ $X2=6.205 $Y2=0.74
r225 24 85 28.3771 $w=1.5e-07 $l=2.73e-07 $layer=POLY_cond $X=6.195 $Y=1.765
+ $X2=6.195 $Y2=1.492
r226 24 26 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=6.195 $Y=1.765
+ $X2=6.195 $Y2=2.4
r227 21 83 28.3771 $w=1.5e-07 $l=2.72e-07 $layer=POLY_cond $X=5.705 $Y=1.22
+ $X2=5.705 $Y2=1.492
r228 21 23 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=5.705 $Y=1.22
+ $X2=5.705 $Y2=0.74
r229 18 82 28.3771 $w=1.5e-07 $l=2.73e-07 $layer=POLY_cond $X=5.695 $Y=1.765
+ $X2=5.695 $Y2=1.492
r230 18 20 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=5.695 $Y=1.765
+ $X2=5.695 $Y2=2.4
r231 16 82 13.032 $w=4.43e-07 $l=1.45186e-07 $layer=POLY_cond $X=5.605 $Y=1.385
+ $X2=5.695 $Y2=1.492
r232 16 60 64.6987 $w=3.3e-07 $l=3.7e-07 $layer=POLY_cond $X=5.605 $Y=1.385
+ $X2=5.235 $Y2=1.385
r233 13 60 149.859 $w=1.8e-07 $l=3.8e-07 $layer=POLY_cond $X=5.145 $Y=1.765
+ $X2=5.145 $Y2=1.385
r234 13 15 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=5.145 $Y=1.765
+ $X2=5.145 $Y2=2.4
r235 12 81 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=5.13 $Y=0.74
+ $X2=5.13 $Y2=1.22
r236 3 73 600 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_PDIFF $count=1 $X=3.01
+ $Y=1.84 $X2=3.165 $Y2=1.985
r237 2 66 300 $w=1.7e-07 $l=2.17428e-07 $layer=licon1_PDIFF $count=2 $X=1.55
+ $Y=1.96 $X2=1.7 $Y2=2.115
r238 1 70 182 $w=1.7e-07 $l=2.08567e-07 $layer=licon1_NDIFF $count=1 $X=2.53
+ $Y=0.37 $X2=2.67 $Y2=0.52
.ends

.subckt PM_SKY130_FD_SC_HS__O2BB2A_4%A_41_392# 1 2 3 10 12 14 16 19 20 21 24
c52 16 0 5.37684e-20 $X=1.25 $Y=2.12
c53 10 0 4.75553e-20 $X=0.35 $Y=2.12
r54 22 24 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=2.15 $Y=2.905
+ $X2=2.15 $Y2=2.455
r55 20 22 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.985 $Y=2.99
+ $X2=2.15 $Y2=2.905
r56 20 21 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=1.985 $Y=2.99
+ $X2=1.415 $Y2=2.99
r57 17 21 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.25 $Y=2.905
+ $X2=1.415 $Y2=2.99
r58 17 19 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=1.25 $Y=2.905 $X2=1.25
+ $Y2=2.815
r59 16 29 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.25 $Y=2.12 $X2=1.25
+ $Y2=2.035
r60 16 19 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=1.25 $Y=2.12
+ $X2=1.25 $Y2=2.815
r61 15 27 5.07788 $w=1.7e-07 $l=1.67481e-07 $layer=LI1_cond $X=0.515 $Y=2.035
+ $X2=0.35 $Y2=2.03
r62 14 29 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.085 $Y=2.035
+ $X2=1.25 $Y2=2.035
r63 14 15 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=1.085 $Y=2.035
+ $X2=0.515 $Y2=2.035
r64 10 27 2.68829 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=0.35 $Y=2.12 $X2=0.35
+ $Y2=2.03
r65 10 12 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=0.35 $Y=2.12
+ $X2=0.35 $Y2=2.815
r66 3 24 300 $w=1.7e-07 $l=5.65044e-07 $layer=licon1_PDIFF $count=2 $X=2 $Y=1.96
+ $X2=2.15 $Y2=2.455
r67 2 29 400 $w=1.7e-07 $l=2.17428e-07 $layer=licon1_PDIFF $count=1 $X=1.1
+ $Y=1.96 $X2=1.25 $Y2=2.115
r68 2 19 400 $w=1.7e-07 $l=9.26971e-07 $layer=licon1_PDIFF $count=1 $X=1.1
+ $Y=1.96 $X2=1.25 $Y2=2.815
r69 1 27 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.205
+ $Y=1.96 $X2=0.35 $Y2=2.105
r70 1 12 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=0.205
+ $Y=1.96 $X2=0.35 $Y2=2.815
.ends

.subckt PM_SKY130_FD_SC_HS__O2BB2A_4%VPWR 1 2 3 4 5 6 23 27 29 33 37 41 45 47 52
+ 53 54 56 68 72 78 81 84 87 91
r98 90 91 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r99 87 88 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r100 81 82 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r101 78 79 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r102 76 91 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=6.96 $Y2=3.33
r103 76 88 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=3.33 $X2=6
+ $Y2=3.33
r104 75 76 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r105 73 87 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.085 $Y=3.33
+ $X2=5.92 $Y2=3.33
r106 73 75 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=6.085 $Y=3.33
+ $X2=6.48 $Y2=3.33
r107 72 90 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=6.755 $Y=3.33
+ $X2=6.977 $Y2=3.33
r108 72 75 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=6.755 $Y=3.33
+ $X2=6.48 $Y2=3.33
r109 71 88 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=3.33 $X2=6
+ $Y2=3.33
r110 70 71 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r111 68 87 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.755 $Y=3.33
+ $X2=5.92 $Y2=3.33
r112 68 70 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=5.755 $Y=3.33
+ $X2=5.52 $Y2=3.33
r113 67 71 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=5.52 $Y2=3.33
r114 66 67 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r115 64 84 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.93 $Y=3.33
+ $X2=3.765 $Y2=3.33
r116 64 66 41.1016 $w=1.68e-07 $l=6.3e-07 $layer=LI1_cond $X=3.93 $Y=3.33
+ $X2=4.56 $Y2=3.33
r117 63 82 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r118 62 63 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r119 60 63 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.16 $Y2=3.33
r120 60 79 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r121 59 62 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.2 $Y=3.33 $X2=2.16
+ $Y2=3.33
r122 59 60 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r123 57 78 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.885 $Y=3.33
+ $X2=0.8 $Y2=3.33
r124 57 59 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=0.885 $Y=3.33
+ $X2=1.2 $Y2=3.33
r125 56 81 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.545 $Y=3.33
+ $X2=2.71 $Y2=3.33
r126 56 62 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=2.545 $Y=3.33
+ $X2=2.16 $Y2=3.33
r127 54 67 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.56 $Y2=3.33
r128 54 82 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=2.64 $Y2=3.33
r129 54 84 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r130 52 66 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=4.67 $Y=3.33
+ $X2=4.56 $Y2=3.33
r131 52 53 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.67 $Y=3.33
+ $X2=4.835 $Y2=3.33
r132 51 70 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=5 $Y=3.33 $X2=5.52
+ $Y2=3.33
r133 51 53 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5 $Y=3.33 $X2=4.835
+ $Y2=3.33
r134 47 50 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=6.92 $Y=1.985
+ $X2=6.92 $Y2=2.815
r135 45 90 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=6.92 $Y=3.245
+ $X2=6.977 $Y2=3.33
r136 45 50 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=6.92 $Y=3.245
+ $X2=6.92 $Y2=2.815
r137 41 44 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=5.92 $Y=2.145
+ $X2=5.92 $Y2=2.825
r138 39 87 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.92 $Y=3.245
+ $X2=5.92 $Y2=3.33
r139 39 44 14.6675 $w=3.28e-07 $l=4.2e-07 $layer=LI1_cond $X=5.92 $Y=3.245
+ $X2=5.92 $Y2=2.825
r140 35 53 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.835 $Y=3.245
+ $X2=4.835 $Y2=3.33
r141 35 37 10.1275 $w=3.28e-07 $l=2.9e-07 $layer=LI1_cond $X=4.835 $Y=3.245
+ $X2=4.835 $Y2=2.955
r142 31 84 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.765 $Y=3.245
+ $X2=3.765 $Y2=3.33
r143 31 33 10.1275 $w=3.28e-07 $l=2.9e-07 $layer=LI1_cond $X=3.765 $Y=3.245
+ $X2=3.765 $Y2=2.955
r144 30 81 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.875 $Y=3.33
+ $X2=2.71 $Y2=3.33
r145 29 84 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.6 $Y=3.33
+ $X2=3.765 $Y2=3.33
r146 29 30 47.2995 $w=1.68e-07 $l=7.25e-07 $layer=LI1_cond $X=3.6 $Y=3.33
+ $X2=2.875 $Y2=3.33
r147 25 81 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.71 $Y=3.245
+ $X2=2.71 $Y2=3.33
r148 25 27 25.668 $w=3.28e-07 $l=7.35e-07 $layer=LI1_cond $X=2.71 $Y=3.245
+ $X2=2.71 $Y2=2.51
r149 21 78 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.8 $Y=3.245 $X2=0.8
+ $Y2=3.33
r150 21 23 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=0.8 $Y=3.245
+ $X2=0.8 $Y2=2.455
r151 6 50 400 $w=1.7e-07 $l=1.06806e-06 $layer=licon1_PDIFF $count=1 $X=6.725
+ $Y=1.84 $X2=6.92 $Y2=2.815
r152 6 47 400 $w=1.7e-07 $l=2.57488e-07 $layer=licon1_PDIFF $count=1 $X=6.725
+ $Y=1.84 $X2=6.92 $Y2=1.985
r153 5 44 400 $w=1.7e-07 $l=1.05734e-06 $layer=licon1_PDIFF $count=1 $X=5.77
+ $Y=1.84 $X2=5.92 $Y2=2.825
r154 5 41 400 $w=1.7e-07 $l=3.72525e-07 $layer=licon1_PDIFF $count=1 $X=5.77
+ $Y=1.84 $X2=5.92 $Y2=2.145
r155 4 37 600 $w=1.7e-07 $l=1.22689e-06 $layer=licon1_PDIFF $count=1 $X=4.6
+ $Y=1.84 $X2=4.835 $Y2=2.955
r156 3 33 600 $w=1.7e-07 $l=1.22689e-06 $layer=licon1_PDIFF $count=1 $X=3.53
+ $Y=1.84 $X2=3.765 $Y2=2.955
r157 2 27 600 $w=1.7e-07 $l=7.38952e-07 $layer=licon1_PDIFF $count=1 $X=2.565
+ $Y=1.84 $X2=2.71 $Y2=2.51
r158 1 23 300 $w=1.7e-07 $l=5.65044e-07 $layer=licon1_PDIFF $count=2 $X=0.65
+ $Y=1.96 $X2=0.8 $Y2=2.455
.ends

.subckt PM_SKY130_FD_SC_HS__O2BB2A_4%X 1 2 3 4 13 15 19 23 24 27 30 33 37 38 39
+ 40 41
r68 40 45 4.07572 $w=2.4e-07 $l=1.65e-07 $layer=LI1_cond $X=5.42 $Y=0.93
+ $X2=5.585 $Y2=0.93
r69 40 41 19.4475 $w=2.38e-07 $l=4.05e-07 $layer=LI1_cond $X=5.595 $Y=0.93 $X2=6
+ $Y2=0.93
r70 40 45 0.480185 $w=2.38e-07 $l=1e-08 $layer=LI1_cond $X=5.595 $Y=0.93
+ $X2=5.585 $Y2=0.93
r71 37 41 12.2447 $w=2.38e-07 $l=2.55e-07 $layer=LI1_cond $X=6.255 $Y=0.93 $X2=6
+ $Y2=0.93
r72 37 38 2.51069 $w=2.4e-07 $l=1.65e-07 $layer=LI1_cond $X=6.255 $Y=0.93
+ $X2=6.42 $Y2=0.93
r73 33 35 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=6.42 $Y=1.985
+ $X2=6.42 $Y2=2.815
r74 31 39 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.42 $Y=1.89 $X2=6.42
+ $Y2=1.805
r75 31 33 3.31764 $w=3.28e-07 $l=9.5e-08 $layer=LI1_cond $X=6.42 $Y=1.89
+ $X2=6.42 $Y2=1.985
r76 30 39 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.42 $Y=1.72 $X2=6.42
+ $Y2=1.805
r77 29 38 3.93362 $w=3.3e-07 $l=1.2e-07 $layer=LI1_cond $X=6.42 $Y=1.05 $X2=6.42
+ $Y2=0.93
r78 29 30 23.3981 $w=3.28e-07 $l=6.7e-07 $layer=LI1_cond $X=6.42 $Y=1.05
+ $X2=6.42 $Y2=1.72
r79 25 38 3.93362 $w=3.3e-07 $l=1.2e-07 $layer=LI1_cond $X=6.42 $Y=0.81 $X2=6.42
+ $Y2=0.93
r80 25 27 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=6.42 $Y=0.81
+ $X2=6.42 $Y2=0.515
r81 23 39 3.80956 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.255 $Y=1.805
+ $X2=6.42 $Y2=1.805
r82 23 24 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=6.255 $Y=1.805
+ $X2=5.585 $Y2=1.805
r83 19 21 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=5.42 $Y=1.985
+ $X2=5.42 $Y2=2.815
r84 17 24 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=5.42 $Y=1.89
+ $X2=5.585 $Y2=1.805
r85 17 19 3.31764 $w=3.28e-07 $l=9.5e-08 $layer=LI1_cond $X=5.42 $Y=1.89
+ $X2=5.42 $Y2=1.985
r86 13 40 2.96416 $w=3.3e-07 $l=1.2e-07 $layer=LI1_cond $X=5.42 $Y=0.81 $X2=5.42
+ $Y2=0.93
r87 13 15 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=5.42 $Y=0.81
+ $X2=5.42 $Y2=0.515
r88 4 35 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=6.27
+ $Y=1.84 $X2=6.42 $Y2=2.815
r89 4 33 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=6.27
+ $Y=1.84 $X2=6.42 $Y2=1.985
r90 3 21 400 $w=1.7e-07 $l=1.07034e-06 $layer=licon1_PDIFF $count=1 $X=5.22
+ $Y=1.84 $X2=5.42 $Y2=2.815
r91 3 19 400 $w=1.7e-07 $l=2.62678e-07 $layer=licon1_PDIFF $count=1 $X=5.22
+ $Y=1.84 $X2=5.42 $Y2=1.985
r92 2 27 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=6.28
+ $Y=0.37 $X2=6.42 $Y2=0.515
r93 1 15 91 $w=1.7e-07 $l=2.78209e-07 $layer=licon1_NDIFF $count=2 $X=5.205
+ $Y=0.37 $X2=5.42 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__O2BB2A_4%A_27_74# 1 2 3 4 15 17 18 21 23 27 29
c53 21 0 1.72779e-19 $X=1.28 $Y=0.515
r54 29 31 4.36531 $w=3.28e-07 $l=1.25e-07 $layer=LI1_cond $X=3.17 $Y=0.81
+ $X2=3.17 $Y2=0.935
r55 24 27 6.67463 $w=2.4e-07 $l=1.65e-07 $layer=LI1_cond $X=1.445 $Y=0.935
+ $X2=1.28 $Y2=0.935
r56 24 26 28.997 $w=3.08e-07 $l=7.8e-07 $layer=LI1_cond $X=1.445 $Y=0.935
+ $X2=2.225 $Y2=0.935
r57 23 31 1.09485 $w=3.1e-07 $l=1.65e-07 $layer=LI1_cond $X=3.005 $Y=0.935
+ $X2=3.17 $Y2=0.935
r58 23 26 28.997 $w=3.08e-07 $l=7.8e-07 $layer=LI1_cond $X=3.005 $Y=0.935
+ $X2=2.225 $Y2=0.935
r59 19 27 0.225187 $w=3.3e-07 $l=1.55e-07 $layer=LI1_cond $X=1.28 $Y=0.78
+ $X2=1.28 $Y2=0.935
r60 19 21 9.25447 $w=3.28e-07 $l=2.65e-07 $layer=LI1_cond $X=1.28 $Y=0.78
+ $X2=1.28 $Y2=0.515
r61 17 27 6.67463 $w=2.4e-07 $l=1.96914e-07 $layer=LI1_cond $X=1.115 $Y=1.005
+ $X2=1.28 $Y2=0.935
r62 17 18 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.115 $Y=1.005
+ $X2=0.445 $Y2=1.005
r63 13 18 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.28 $Y=0.92
+ $X2=0.445 $Y2=1.005
r64 13 15 14.1436 $w=3.28e-07 $l=4.05e-07 $layer=LI1_cond $X=0.28 $Y=0.92
+ $X2=0.28 $Y2=0.515
r65 4 29 182 $w=1.7e-07 $l=5.20192e-07 $layer=licon1_NDIFF $count=1 $X=2.995
+ $Y=0.37 $X2=3.17 $Y2=0.81
r66 3 26 182 $w=1.7e-07 $l=5.6723e-07 $layer=licon1_NDIFF $count=1 $X=2.07
+ $Y=0.37 $X2=2.225 $Y2=0.865
r67 2 21 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.14
+ $Y=0.37 $X2=1.28 $Y2=0.515
r68 1 15 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__O2BB2A_4%VGND 1 2 3 4 5 18 20 24 28 32 34 36 38 40
+ 45 50 55 61 64 67 70 74
c86 28 0 1.762e-19 $X=4.81 $Y=0.64
r87 73 74 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=0 $X2=6.96
+ $Y2=0
r88 70 71 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=0 $X2=6 $Y2=0
r89 67 68 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r90 64 65 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r91 62 65 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r92 61 62 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r93 59 74 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=0 $X2=6.96
+ $Y2=0
r94 59 71 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=0 $X2=6
+ $Y2=0
r95 58 59 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=0 $X2=6.48
+ $Y2=0
r96 56 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.085 $Y=0 $X2=5.92
+ $Y2=0
r97 56 58 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=6.085 $Y=0 $X2=6.48
+ $Y2=0
r98 55 73 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=6.755 $Y=0 $X2=6.977
+ $Y2=0
r99 55 58 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=6.755 $Y=0 $X2=6.48
+ $Y2=0
r100 54 71 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=6
+ $Y2=0
r101 54 68 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=4.56
+ $Y2=0
r102 53 54 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r103 51 67 11.8214 $w=1.7e-07 $l=2.7e-07 $layer=LI1_cond $X=5.08 $Y=0 $X2=4.81
+ $Y2=0
r104 51 53 28.7059 $w=1.68e-07 $l=4.4e-07 $layer=LI1_cond $X=5.08 $Y=0 $X2=5.52
+ $Y2=0
r105 50 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.755 $Y=0 $X2=5.92
+ $Y2=0
r106 50 53 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=5.755 $Y=0
+ $X2=5.52 $Y2=0
r107 49 65 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.68
+ $Y2=0
r108 48 49 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r109 46 64 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.945 $Y=0 $X2=1.78
+ $Y2=0
r110 46 48 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=1.945 $Y=0
+ $X2=2.16 $Y2=0
r111 45 67 11.8214 $w=1.7e-07 $l=2.7e-07 $layer=LI1_cond $X=4.54 $Y=0 $X2=4.81
+ $Y2=0
r112 45 48 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=4.54 $Y=0 $X2=2.16
+ $Y2=0
r113 43 62 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r114 42 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r115 40 61 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.615 $Y=0 $X2=0.78
+ $Y2=0
r116 40 42 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=0.615 $Y=0
+ $X2=0.24 $Y2=0
r117 38 68 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.56
+ $Y2=0
r118 38 49 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=3.6 $Y=0 $X2=2.16
+ $Y2=0
r119 34 73 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=6.92 $Y=0.085
+ $X2=6.977 $Y2=0
r120 34 36 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=6.92 $Y=0.085
+ $X2=6.92 $Y2=0.515
r121 30 70 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.92 $Y=0.085
+ $X2=5.92 $Y2=0
r122 30 32 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=5.92 $Y=0.085
+ $X2=5.92 $Y2=0.535
r123 26 67 2.26835 $w=5.4e-07 $l=8.5e-08 $layer=LI1_cond $X=4.81 $Y=0.085
+ $X2=4.81 $Y2=0
r124 26 28 12.293 $w=5.38e-07 $l=5.55e-07 $layer=LI1_cond $X=4.81 $Y=0.085
+ $X2=4.81 $Y2=0.64
r125 22 64 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.78 $Y=0.085
+ $X2=1.78 $Y2=0
r126 22 24 15.1913 $w=3.28e-07 $l=4.35e-07 $layer=LI1_cond $X=1.78 $Y=0.085
+ $X2=1.78 $Y2=0.52
r127 21 61 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.945 $Y=0 $X2=0.78
+ $Y2=0
r128 20 64 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.615 $Y=0 $X2=1.78
+ $Y2=0
r129 20 21 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.615 $Y=0
+ $X2=0.945 $Y2=0
r130 16 61 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.78 $Y=0.085
+ $X2=0.78 $Y2=0
r131 16 18 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=0.78 $Y=0.085
+ $X2=0.78 $Y2=0.55
r132 5 36 91 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=2 $X=6.71
+ $Y=0.37 $X2=6.92 $Y2=0.515
r133 4 32 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=5.78
+ $Y=0.37 $X2=5.92 $Y2=0.535
r134 3 28 182 $w=1.7e-07 $l=3.18865e-07 $layer=licon1_NDIFF $count=1 $X=4.565
+ $Y=0.47 $X2=4.81 $Y2=0.64
r135 2 24 182 $w=1.7e-07 $l=2.74955e-07 $layer=licon1_NDIFF $count=1 $X=1.57
+ $Y=0.37 $X2=1.78 $Y2=0.52
r136 1 18 182 $w=1.7e-07 $l=2.86182e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.37 $X2=0.78 $Y2=0.55
.ends

