# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_hs__fah_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  14.40000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.565000 1.290000 2.045000 1.780000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.723000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.555000 1.355000 2.895000 2.150000 ;
        RECT 2.725000 0.595000 5.435000 0.765000 ;
        RECT 2.725000 0.765000 2.895000 1.355000 ;
        RECT 3.440000 1.630000 3.770000 1.960000 ;
        RECT 3.565000 0.765000 3.735000 1.630000 ;
        RECT 4.405000 0.765000 4.595000 1.605000 ;
        RECT 5.265000 0.765000 5.435000 0.920000 ;
        RECT 5.265000 0.920000 6.205000 1.090000 ;
        RECT 5.875000 1.090000 6.205000 1.185000 ;
    END
  END B
  PIN CI
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 11.450000 1.450000 11.875000 1.780000 ;
    END
  END CI
  PIN COUT
    ANTENNADIFFAREA  0.543200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 12.585000 0.350000 12.835000 1.550000 ;
        RECT 12.585000 1.550000 12.920000 2.200000 ;
    END
  END COUT
  PIN SUM
    ANTENNADIFFAREA  0.561800 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 13.515000 0.355000 13.785000 0.800000 ;
        RECT 13.515000 0.800000 14.275000 1.130000 ;
        RECT 13.570000 1.820000 13.875000 2.980000 ;
        RECT 13.705000 1.130000 14.275000 1.505000 ;
        RECT 13.705000 1.505000 13.875000 1.820000 ;
    END
  END SUM
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 14.400000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 14.400000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 14.400000 0.085000 ;
      RECT  0.000000  3.245000 14.400000 3.415000 ;
      RECT  0.105000  2.160000  0.360000 3.245000 ;
      RECT  0.125000  1.180000  0.650000 1.470000 ;
      RECT  0.170000  0.085000  0.535000 0.790000 ;
      RECT  0.335000  1.470000  0.650000 1.820000 ;
      RECT  0.335000  1.820000  0.885000 1.990000 ;
      RECT  0.480000  0.960000  0.965000 1.130000 ;
      RECT  0.480000  1.130000  0.650000 1.180000 ;
      RECT  0.555000  1.990000  0.885000 2.980000 ;
      RECT  0.705000  0.350000  0.965000 0.960000 ;
      RECT  0.820000  1.300000  1.395000 1.630000 ;
      RECT  1.090000  1.630000  1.340000 2.980000 ;
      RECT  1.225000  0.505000  1.705000 1.120000 ;
      RECT  1.225000  1.120000  1.395000 1.300000 ;
      RECT  1.540000  1.950000  1.870000 3.245000 ;
      RECT  1.875000  0.085000  2.125000 0.845000 ;
      RECT  2.055000  2.015000  2.385000 2.890000 ;
      RECT  2.055000  2.890000  6.055000 3.060000 ;
      RECT  2.215000  1.015000  2.555000 1.185000 ;
      RECT  2.215000  1.185000  2.385000 2.015000 ;
      RECT  2.305000  0.255000  5.935000 0.425000 ;
      RECT  2.305000  0.425000  2.555000 1.015000 ;
      RECT  2.555000  2.390000  3.450000 2.550000 ;
      RECT  2.555000  2.550000  5.555000 2.720000 ;
      RECT  3.065000  0.935000  3.395000 1.185000 ;
      RECT  3.065000  1.185000  3.235000 2.390000 ;
      RECT  3.620000  2.130000  4.110000 2.380000 ;
      RECT  3.905000  0.935000  4.235000 1.185000 ;
      RECT  3.940000  1.185000  4.235000 1.410000 ;
      RECT  3.940000  1.410000  4.110000 2.130000 ;
      RECT  4.280000  2.100000  5.215000 2.350000 ;
      RECT  4.765000  0.935000  5.095000 1.260000 ;
      RECT  4.765000  1.260000  5.705000 1.355000 ;
      RECT  4.765000  1.355000  6.545000 1.430000 ;
      RECT  4.765000  1.430000  4.935000 2.100000 ;
      RECT  5.105000  1.600000  5.365000 1.760000 ;
      RECT  5.105000  1.760000  7.045000 1.930000 ;
      RECT  5.385000  2.100000  6.395000 2.240000 ;
      RECT  5.385000  2.240000  7.385000 2.270000 ;
      RECT  5.385000  2.270000  5.555000 2.550000 ;
      RECT  5.535000  1.430000  6.545000 1.525000 ;
      RECT  5.605000  0.425000  5.935000 0.750000 ;
      RECT  5.725000  2.440000  6.055000 2.890000 ;
      RECT  6.225000  2.270000  7.385000 2.410000 ;
      RECT  6.265000  2.580000  6.595000 3.245000 ;
      RECT  6.335000  0.085000  6.665000 0.680000 ;
      RECT  6.375000  0.850000  7.005000 1.020000 ;
      RECT  6.375000  1.020000  6.545000 1.355000 ;
      RECT  6.715000  1.190000  7.505000 1.360000 ;
      RECT  6.715000  1.360000  7.045000 1.760000 ;
      RECT  6.715000  1.930000  7.045000 2.070000 ;
      RECT  6.835000  0.255000  7.845000 0.425000 ;
      RECT  6.835000  0.425000  7.005000 0.850000 ;
      RECT  7.175000  0.630000  7.505000 1.190000 ;
      RECT  7.215000  1.630000  7.505000 1.960000 ;
      RECT  7.215000  1.960000  7.385000 2.240000 ;
      RECT  7.215000  2.410000  7.385000 2.905000 ;
      RECT  7.215000  2.905000  9.575000 3.075000 ;
      RECT  7.555000  2.130000  8.310000 2.735000 ;
      RECT  7.675000  0.425000  7.845000 1.275000 ;
      RECT  7.675000  1.275000  7.970000 1.945000 ;
      RECT  8.015000  0.390000  8.555000 0.640000 ;
      RECT  8.140000  0.640000  8.555000 1.040000 ;
      RECT  8.140000  1.040000  8.310000 2.130000 ;
      RECT  8.480000  1.225000  8.735000 2.905000 ;
      RECT  8.745000  0.255000 10.935000 0.425000 ;
      RECT  8.745000  0.425000  9.075000 1.055000 ;
      RECT  8.905000  1.055000  9.075000 2.130000 ;
      RECT  8.905000  2.130000  9.235000 2.735000 ;
      RECT  9.245000  0.595000 10.255000 0.765000 ;
      RECT  9.245000  0.765000  9.415000 1.630000 ;
      RECT  9.245000  1.630000  9.575000 1.960000 ;
      RECT  9.405000  1.960000  9.575000 2.905000 ;
      RECT  9.585000  0.935000  9.915000 1.185000 ;
      RECT  9.745000  1.185000  9.915000 2.100000 ;
      RECT  9.745000  2.100000 10.075000 2.600000 ;
      RECT  9.745000  2.600000 11.970000 2.770000 ;
      RECT  9.745000  2.770000 10.075000 2.980000 ;
      RECT 10.085000  0.765000 10.255000 1.355000 ;
      RECT 10.085000  1.355000 10.470000 1.685000 ;
      RECT 10.310000  2.130000 10.810000 2.430000 ;
      RECT 10.425000  0.595000 10.595000 1.015000 ;
      RECT 10.425000  1.015000 10.810000 1.185000 ;
      RECT 10.640000  1.185000 10.810000 2.130000 ;
      RECT 10.765000  0.425000 10.935000 0.675000 ;
      RECT 10.765000  0.675000 11.865000 0.845000 ;
      RECT 10.980000  0.845000 11.865000 1.055000 ;
      RECT 10.980000  1.055000 11.240000 1.950000 ;
      RECT 10.980000  1.950000 11.930000 2.200000 ;
      RECT 11.015000  2.940000 11.395000 3.245000 ;
      RECT 11.105000  0.085000 11.355000 0.505000 ;
      RECT 11.535000  0.375000 11.865000 0.675000 ;
      RECT 11.800000  2.370000 13.400000 2.540000 ;
      RECT 11.800000  2.540000 11.970000 2.600000 ;
      RECT 12.075000  0.085000 12.405000 0.640000 ;
      RECT 12.085000  0.810000 12.415000 1.550000 ;
      RECT 12.140000  2.710000 12.470000 3.245000 ;
      RECT 13.015000  0.085000 13.345000 1.130000 ;
      RECT 13.040000  2.710000 13.370000 3.245000 ;
      RECT 13.230000  1.300000 13.535000 1.630000 ;
      RECT 13.230000  1.630000 13.400000 2.370000 ;
      RECT 13.955000  0.085000 14.285000 0.630000 ;
      RECT 14.045000  1.820000 14.295000 3.245000 ;
    LAYER mcon ;
      RECT  0.155000 -0.085000  0.325000 0.085000 ;
      RECT  0.155000  1.210000  0.325000 1.380000 ;
      RECT  0.155000  3.245000  0.325000 3.415000 ;
      RECT  0.635000 -0.085000  0.805000 0.085000 ;
      RECT  0.635000  3.245000  0.805000 3.415000 ;
      RECT  1.115000 -0.085000  1.285000 0.085000 ;
      RECT  1.115000  3.245000  1.285000 3.415000 ;
      RECT  1.595000 -0.085000  1.765000 0.085000 ;
      RECT  1.595000  3.245000  1.765000 3.415000 ;
      RECT  2.075000 -0.085000  2.245000 0.085000 ;
      RECT  2.075000  3.245000  2.245000 3.415000 ;
      RECT  2.555000 -0.085000  2.725000 0.085000 ;
      RECT  2.555000  3.245000  2.725000 3.415000 ;
      RECT  3.035000 -0.085000  3.205000 0.085000 ;
      RECT  3.035000  3.245000  3.205000 3.415000 ;
      RECT  3.515000 -0.085000  3.685000 0.085000 ;
      RECT  3.515000  3.245000  3.685000 3.415000 ;
      RECT  3.995000 -0.085000  4.165000 0.085000 ;
      RECT  3.995000  1.210000  4.165000 1.380000 ;
      RECT  3.995000  3.245000  4.165000 3.415000 ;
      RECT  4.475000 -0.085000  4.645000 0.085000 ;
      RECT  4.475000  3.245000  4.645000 3.415000 ;
      RECT  4.955000 -0.085000  5.125000 0.085000 ;
      RECT  4.955000  3.245000  5.125000 3.415000 ;
      RECT  5.435000 -0.085000  5.605000 0.085000 ;
      RECT  5.435000  3.245000  5.605000 3.415000 ;
      RECT  5.915000 -0.085000  6.085000 0.085000 ;
      RECT  5.915000  3.245000  6.085000 3.415000 ;
      RECT  6.395000 -0.085000  6.565000 0.085000 ;
      RECT  6.395000  3.245000  6.565000 3.415000 ;
      RECT  6.875000 -0.085000  7.045000 0.085000 ;
      RECT  6.875000  3.245000  7.045000 3.415000 ;
      RECT  7.355000 -0.085000  7.525000 0.085000 ;
      RECT  7.355000  3.245000  7.525000 3.415000 ;
      RECT  7.835000 -0.085000  8.005000 0.085000 ;
      RECT  7.835000  3.245000  8.005000 3.415000 ;
      RECT  8.315000 -0.085000  8.485000 0.085000 ;
      RECT  8.315000  0.840000  8.485000 1.010000 ;
      RECT  8.315000  3.245000  8.485000 3.415000 ;
      RECT  8.795000 -0.085000  8.965000 0.085000 ;
      RECT  8.795000  3.245000  8.965000 3.415000 ;
      RECT  9.275000 -0.085000  9.445000 0.085000 ;
      RECT  9.275000  3.245000  9.445000 3.415000 ;
      RECT  9.755000 -0.085000  9.925000 0.085000 ;
      RECT  9.755000  3.245000  9.925000 3.415000 ;
      RECT 10.235000 -0.085000 10.405000 0.085000 ;
      RECT 10.235000  3.245000 10.405000 3.415000 ;
      RECT 10.715000 -0.085000 10.885000 0.085000 ;
      RECT 10.715000  3.245000 10.885000 3.415000 ;
      RECT 11.195000 -0.085000 11.365000 0.085000 ;
      RECT 11.195000  3.245000 11.365000 3.415000 ;
      RECT 11.675000 -0.085000 11.845000 0.085000 ;
      RECT 11.675000  3.245000 11.845000 3.415000 ;
      RECT 12.155000 -0.085000 12.325000 0.085000 ;
      RECT 12.155000  0.840000 12.325000 1.010000 ;
      RECT 12.155000  3.245000 12.325000 3.415000 ;
      RECT 12.635000 -0.085000 12.805000 0.085000 ;
      RECT 12.635000  3.245000 12.805000 3.415000 ;
      RECT 13.115000 -0.085000 13.285000 0.085000 ;
      RECT 13.115000  3.245000 13.285000 3.415000 ;
      RECT 13.595000 -0.085000 13.765000 0.085000 ;
      RECT 13.595000  3.245000 13.765000 3.415000 ;
      RECT 14.075000 -0.085000 14.245000 0.085000 ;
      RECT 14.075000  3.245000 14.245000 3.415000 ;
    LAYER met1 ;
      RECT  0.095000 1.180000  0.385000 1.225000 ;
      RECT  0.095000 1.225000  4.225000 1.365000 ;
      RECT  0.095000 1.365000  0.385000 1.410000 ;
      RECT  3.935000 1.180000  4.225000 1.225000 ;
      RECT  3.935000 1.365000  4.225000 1.410000 ;
      RECT  8.255000 0.810000  8.545000 0.855000 ;
      RECT  8.255000 0.855000 12.385000 0.995000 ;
      RECT  8.255000 0.995000  8.545000 1.040000 ;
      RECT 12.095000 0.810000 12.385000 0.855000 ;
      RECT 12.095000 0.995000 12.385000 1.040000 ;
  END
END sky130_fd_sc_hs__fah_2
END LIBRARY
