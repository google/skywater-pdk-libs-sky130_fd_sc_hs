# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_hs__a41o_4
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_hs__a41o_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  8.160000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.522000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.485000 1.450000 4.195000 1.780000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.522000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.900000 1.450000 5.635000 1.780000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.522000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.885000 1.450000 7.075000 1.780000 ;
    END
  END A3
  PIN A4
    ANTENNAGATEAREA  0.522000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.325000 1.450000 8.035000 1.780000 ;
    END
  END A4
  PIN B1
    ANTENNAGATEAREA  0.522000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.450000 0.550000 1.780000 ;
    END
  END B1
  PIN X
    ANTENNADIFFAREA  1.086400 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.550000 1.000000 3.305000 1.170000 ;
        RECT 2.075000 1.840000 3.305000 2.120000 ;
        RECT 2.555000 1.170000 3.305000 1.840000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 8.160000 0.085000 ;
        RECT 0.110000  0.085000 0.360000 1.250000 ;
        RECT 1.045000  0.085000 1.375000 0.490000 ;
        RECT 2.055000  0.085000 2.385000 0.490000 ;
        RECT 3.055000  0.085000 3.305000 0.490000 ;
        RECT 7.290000  0.085000 7.620000 0.940000 ;
      LAYER mcon ;
        RECT 0.155000 -0.085000 0.325000 0.085000 ;
        RECT 0.635000 -0.085000 0.805000 0.085000 ;
        RECT 1.115000 -0.085000 1.285000 0.085000 ;
        RECT 1.595000 -0.085000 1.765000 0.085000 ;
        RECT 2.075000 -0.085000 2.245000 0.085000 ;
        RECT 2.555000 -0.085000 2.725000 0.085000 ;
        RECT 3.035000 -0.085000 3.205000 0.085000 ;
        RECT 3.515000 -0.085000 3.685000 0.085000 ;
        RECT 3.995000 -0.085000 4.165000 0.085000 ;
        RECT 4.475000 -0.085000 4.645000 0.085000 ;
        RECT 4.955000 -0.085000 5.125000 0.085000 ;
        RECT 5.435000 -0.085000 5.605000 0.085000 ;
        RECT 5.915000 -0.085000 6.085000 0.085000 ;
        RECT 6.395000 -0.085000 6.565000 0.085000 ;
        RECT 6.875000 -0.085000 7.045000 0.085000 ;
        RECT 7.355000 -0.085000 7.525000 0.085000 ;
        RECT 7.835000 -0.085000 8.005000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.245000 8.160000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 3.245000 8.160000 3.415000 ;
        RECT 1.625000 2.630000 1.955000 3.245000 ;
        RECT 2.525000 2.630000 2.855000 3.245000 ;
        RECT 3.425000 2.650000 3.775000 3.245000 ;
        RECT 4.635000 2.290000 5.095000 3.245000 ;
        RECT 5.765000 2.290000 6.095000 3.245000 ;
        RECT 6.765000 2.290000 7.095000 3.245000 ;
        RECT 7.795000 1.950000 8.045000 3.245000 ;
      LAYER mcon ;
        RECT 0.155000 3.245000 0.325000 3.415000 ;
        RECT 0.635000 3.245000 0.805000 3.415000 ;
        RECT 1.115000 3.245000 1.285000 3.415000 ;
        RECT 1.595000 3.245000 1.765000 3.415000 ;
        RECT 2.075000 3.245000 2.245000 3.415000 ;
        RECT 2.555000 3.245000 2.725000 3.415000 ;
        RECT 3.035000 3.245000 3.205000 3.415000 ;
        RECT 3.515000 3.245000 3.685000 3.415000 ;
        RECT 3.995000 3.245000 4.165000 3.415000 ;
        RECT 4.475000 3.245000 4.645000 3.415000 ;
        RECT 4.955000 3.245000 5.125000 3.415000 ;
        RECT 5.435000 3.245000 5.605000 3.415000 ;
        RECT 5.915000 3.245000 6.085000 3.415000 ;
        RECT 6.395000 3.245000 6.565000 3.415000 ;
        RECT 6.875000 3.245000 7.045000 3.415000 ;
        RECT 7.355000 3.245000 7.525000 3.415000 ;
        RECT 7.835000 3.245000 8.005000 3.415000 ;
      LAYER met1 ;
        RECT 0.000000 3.085000 8.160000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.115000 1.950000 0.445000 2.905000 ;
      RECT 0.115000 2.905000 1.395000 3.075000 ;
      RECT 0.540000 0.470000 0.870000 0.660000 ;
      RECT 0.540000 0.660000 3.645000 0.830000 ;
      RECT 0.540000 0.830000 1.225000 1.250000 ;
      RECT 0.615000 1.950000 0.890000 2.735000 ;
      RECT 0.720000 1.250000 1.225000 1.340000 ;
      RECT 0.720000 1.340000 2.385000 1.670000 ;
      RECT 0.720000 1.670000 0.890000 1.950000 ;
      RECT 1.065000 1.940000 1.395000 2.290000 ;
      RECT 1.065000 2.290000 4.375000 2.460000 ;
      RECT 1.065000 2.460000 1.395000 2.905000 ;
      RECT 3.475000 0.255000 4.495000 0.425000 ;
      RECT 3.475000 0.425000 3.645000 0.660000 ;
      RECT 3.815000 0.700000 3.985000 0.770000 ;
      RECT 3.815000 0.770000 4.845000 1.150000 ;
      RECT 4.045000 1.950000 7.595000 2.120000 ;
      RECT 4.045000 2.120000 4.375000 2.290000 ;
      RECT 4.045000 2.460000 4.375000 2.980000 ;
      RECT 4.165000 0.425000 4.495000 0.600000 ;
      RECT 4.675000 0.330000 5.785000 0.600000 ;
      RECT 4.675000 0.600000 4.845000 0.770000 ;
      RECT 5.025000 0.770000 5.285000 1.110000 ;
      RECT 5.025000 1.110000 6.680000 1.280000 ;
      RECT 5.265000 2.120000 5.595000 2.980000 ;
      RECT 5.455000 0.600000 5.785000 0.940000 ;
      RECT 6.000000 0.255000 7.110000 0.425000 ;
      RECT 6.000000 0.425000 6.330000 0.940000 ;
      RECT 6.265000 2.120000 6.595000 2.980000 ;
      RECT 6.510000 0.595000 6.680000 1.110000 ;
      RECT 6.860000 0.425000 7.110000 1.110000 ;
      RECT 6.860000 1.110000 8.050000 1.280000 ;
      RECT 7.265000 2.120000 7.595000 2.980000 ;
      RECT 7.790000 0.350000 8.050000 1.110000 ;
  END
END sky130_fd_sc_hs__a41o_4
