* File: sky130_fd_sc_hs__nand4_4.pxi.spice
* Created: Thu Aug 27 20:51:59 2020
* 
x_PM_SKY130_FD_SC_HS__NAND4_4%D N_D_M1008_g N_D_M1010_g N_D_c_109_n N_D_M1014_g
+ N_D_c_118_n N_D_M1016_g N_D_M1020_g N_D_c_119_n N_D_M1017_g N_D_c_112_n
+ N_D_c_113_n N_D_c_114_n D D D D D N_D_c_116_n PM_SKY130_FD_SC_HS__NAND4_4%D
x_PM_SKY130_FD_SC_HS__NAND4_4%C N_C_M1002_g N_C_c_187_n N_C_M1000_g N_C_M1011_g
+ N_C_c_188_n N_C_M1019_g N_C_M1012_g N_C_M1021_g C C C C N_C_c_186_n
+ PM_SKY130_FD_SC_HS__NAND4_4%C
x_PM_SKY130_FD_SC_HS__NAND4_4%B N_B_c_245_n N_B_M1001_g N_B_M1006_g N_B_c_246_n
+ N_B_M1009_g N_B_M1007_g N_B_M1018_g N_B_M1022_g B B B B N_B_c_244_n
+ PM_SKY130_FD_SC_HS__NAND4_4%B
x_PM_SKY130_FD_SC_HS__NAND4_4%A N_A_M1005_g N_A_M1013_g N_A_c_311_n N_A_M1003_g
+ N_A_M1015_g N_A_c_312_n N_A_M1004_g N_A_M1023_g N_A_c_308_n N_A_c_309_n A A A
+ N_A_c_310_n PM_SKY130_FD_SC_HS__NAND4_4%A
x_PM_SKY130_FD_SC_HS__NAND4_4%VPWR N_VPWR_M1016_d N_VPWR_M1017_d N_VPWR_M1019_d
+ N_VPWR_M1009_s N_VPWR_M1004_s N_VPWR_c_373_n N_VPWR_c_374_n N_VPWR_c_375_n
+ N_VPWR_c_376_n N_VPWR_c_377_n VPWR N_VPWR_c_378_n N_VPWR_c_379_n
+ N_VPWR_c_380_n N_VPWR_c_381_n N_VPWR_c_382_n N_VPWR_c_383_n N_VPWR_c_384_n
+ N_VPWR_c_372_n PM_SKY130_FD_SC_HS__NAND4_4%VPWR
x_PM_SKY130_FD_SC_HS__NAND4_4%Y N_Y_M1005_d N_Y_M1015_d N_Y_M1016_s N_Y_M1000_s
+ N_Y_M1001_d N_Y_M1003_d N_Y_c_449_n N_Y_c_443_n N_Y_c_454_n N_Y_c_444_n
+ N_Y_c_460_n N_Y_c_445_n N_Y_c_469_n N_Y_c_438_n N_Y_c_446_n N_Y_c_439_n
+ N_Y_c_447_n N_Y_c_463_n N_Y_c_473_n N_Y_c_486_n N_Y_c_440_n N_Y_c_441_n Y Y
+ PM_SKY130_FD_SC_HS__NAND4_4%Y
x_PM_SKY130_FD_SC_HS__NAND4_4%A_27_74# N_A_27_74#_M1008_s N_A_27_74#_M1010_s
+ N_A_27_74#_M1020_s N_A_27_74#_M1011_s N_A_27_74#_M1021_s N_A_27_74#_c_535_n
+ N_A_27_74#_c_536_n N_A_27_74#_c_537_n N_A_27_74#_c_538_n N_A_27_74#_c_539_n
+ N_A_27_74#_c_540_n N_A_27_74#_c_559_n N_A_27_74#_c_541_n N_A_27_74#_c_542_n
+ PM_SKY130_FD_SC_HS__NAND4_4%A_27_74#
x_PM_SKY130_FD_SC_HS__NAND4_4%VGND N_VGND_M1008_d N_VGND_M1014_d N_VGND_c_597_n
+ N_VGND_c_598_n N_VGND_c_599_n VGND N_VGND_c_600_n N_VGND_c_601_n
+ N_VGND_c_602_n N_VGND_c_603_n N_VGND_c_604_n PM_SKY130_FD_SC_HS__NAND4_4%VGND
x_PM_SKY130_FD_SC_HS__NAND4_4%A_554_74# N_A_554_74#_M1002_d N_A_554_74#_M1012_d
+ N_A_554_74#_M1006_s N_A_554_74#_M1018_s N_A_554_74#_c_665_n
+ N_A_554_74#_c_666_n N_A_554_74#_c_667_n N_A_554_74#_c_668_n
+ N_A_554_74#_c_669_n PM_SKY130_FD_SC_HS__NAND4_4%A_554_74#
x_PM_SKY130_FD_SC_HS__NAND4_4%A_923_74# N_A_923_74#_M1006_d N_A_923_74#_M1007_d
+ N_A_923_74#_M1022_d N_A_923_74#_M1013_s N_A_923_74#_M1023_s
+ N_A_923_74#_c_705_n N_A_923_74#_c_706_n N_A_923_74#_c_707_n
+ N_A_923_74#_c_708_n N_A_923_74#_c_709_n N_A_923_74#_c_710_n
+ N_A_923_74#_c_711_n N_A_923_74#_c_712_n N_A_923_74#_c_713_n
+ PM_SKY130_FD_SC_HS__NAND4_4%A_923_74#
cc_1 VNB N_D_M1008_g 0.0336211f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_2 VNB N_D_M1010_g 0.024496f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=0.74
cc_3 VNB N_D_c_109_n 0.0155552f $X=-0.19 $Y=-0.245 $X2=1.42 $Y2=1.515
cc_4 VNB N_D_M1014_g 0.0272963f $X=-0.19 $Y=-0.245 $X2=1.495 $Y2=0.74
cc_5 VNB N_D_M1020_g 0.0277516f $X=-0.19 $Y=-0.245 $X2=2.195 $Y2=0.74
cc_6 VNB N_D_c_112_n 0.0137535f $X=-0.19 $Y=-0.245 $X2=0.57 $Y2=1.515
cc_7 VNB N_D_c_113_n 0.0155576f $X=-0.19 $Y=-0.245 $X2=0.92 $Y2=1.515
cc_8 VNB N_D_c_114_n 0.004935f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=1.515
cc_9 VNB D 0.0166475f $X=-0.19 $Y=-0.245 $X2=2.075 $Y2=1.58
cc_10 VNB N_D_c_116_n 0.0479201f $X=-0.19 $Y=-0.245 $X2=2.195 $Y2=1.557
cc_11 VNB N_C_M1002_g 0.0250243f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_12 VNB N_C_M1011_g 0.0234232f $X=-0.19 $Y=-0.245 $X2=1.07 $Y2=1.515
cc_13 VNB N_C_M1012_g 0.0234256f $X=-0.19 $Y=-0.245 $X2=1.76 $Y2=2.4
cc_14 VNB N_C_M1021_g 0.0337355f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB C 0.00704574f $X=-0.19 $Y=-0.245 $X2=0.92 $Y2=1.515
cc_16 VNB N_C_c_186_n 0.0643418f $X=-0.19 $Y=-0.245 $X2=1.425 $Y2=1.515
cc_17 VNB N_B_M1006_g 0.0336884f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=0.74
cc_18 VNB N_B_M1007_g 0.0234256f $X=-0.19 $Y=-0.245 $X2=1.495 $Y2=0.74
cc_19 VNB N_B_M1018_g 0.0234256f $X=-0.19 $Y=-0.245 $X2=1.76 $Y2=2.4
cc_20 VNB N_B_M1022_g 0.0241156f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB B 0.00267486f $X=-0.19 $Y=-0.245 $X2=0.92 $Y2=1.515
cc_22 VNB N_B_c_244_n 0.0917203f $X=-0.19 $Y=-0.245 $X2=1.425 $Y2=1.515
cc_23 VNB N_A_M1005_g 0.0241156f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_24 VNB N_A_M1013_g 0.0234256f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=0.74
cc_25 VNB N_A_M1015_g 0.0255586f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_M1023_g 0.0301963f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_c_308_n 0.0199044f $X=-0.19 $Y=-0.245 $X2=2.26 $Y2=2.4
cc_28 VNB N_A_c_309_n 0.0136818f $X=-0.19 $Y=-0.245 $X2=2.26 $Y2=2.4
cc_29 VNB N_A_c_310_n 0.0443906f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=1.58
cc_30 VNB N_VPWR_c_372_n 0.362705f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_Y_c_438_n 0.00204539f $X=-0.19 $Y=-0.245 $X2=0.745 $Y2=1.515
cc_32 VNB N_Y_c_439_n 0.0145179f $X=-0.19 $Y=-0.245 $X2=1.425 $Y2=1.515
cc_33 VNB N_Y_c_440_n 0.00408444f $X=-0.19 $Y=-0.245 $X2=1.425 $Y2=1.565
cc_34 VNB N_Y_c_441_n 0.00133991f $X=-0.19 $Y=-0.245 $X2=1.68 $Y2=1.565
cc_35 VNB Y 0.0265321f $X=-0.19 $Y=-0.245 $X2=2.16 $Y2=1.565
cc_36 VNB N_A_27_74#_c_535_n 0.0277086f $X=-0.19 $Y=-0.245 $X2=2.195 $Y2=1.35
cc_37 VNB N_A_27_74#_c_536_n 0.00307912f $X=-0.19 $Y=-0.245 $X2=2.195 $Y2=0.74
cc_38 VNB N_A_27_74#_c_537_n 0.0104987f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_27_74#_c_538_n 0.00280455f $X=-0.19 $Y=-0.245 $X2=2.26 $Y2=2.4
cc_40 VNB N_A_27_74#_c_539_n 0.0136988f $X=-0.19 $Y=-0.245 $X2=0.92 $Y2=1.515
cc_41 VNB N_A_27_74#_c_540_n 0.00261637f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_42 VNB N_A_27_74#_c_541_n 0.0136639f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_27_74#_c_542_n 0.00231148f $X=-0.19 $Y=-0.245 $X2=0.745 $Y2=1.515
cc_44 VNB N_VGND_c_597_n 0.00586453f $X=-0.19 $Y=-0.245 $X2=1.42 $Y2=1.515
cc_45 VNB N_VGND_c_598_n 0.0185368f $X=-0.19 $Y=-0.245 $X2=1.495 $Y2=1.35
cc_46 VNB N_VGND_c_599_n 0.00916033f $X=-0.19 $Y=-0.245 $X2=1.76 $Y2=1.765
cc_47 VNB N_VGND_c_600_n 0.0191515f $X=-0.19 $Y=-0.245 $X2=2.195 $Y2=0.74
cc_48 VNB N_VGND_c_601_n 0.168013f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_49 VNB N_VGND_c_602_n 0.467293f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.58
cc_50 VNB N_VGND_c_603_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_VGND_c_604_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_A_554_74#_c_665_n 0.00641753f $X=-0.19 $Y=-0.245 $X2=1.495 $Y2=0.74
cc_53 VNB N_A_554_74#_c_666_n 0.0062129f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_A_554_74#_c_667_n 0.00108276f $X=-0.19 $Y=-0.245 $X2=2.26 $Y2=2.4
cc_55 VNB N_A_554_74#_c_668_n 0.0265392f $X=-0.19 $Y=-0.245 $X2=0.92 $Y2=1.515
cc_56 VNB N_A_554_74#_c_669_n 0.00159267f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=1.515
cc_57 VNB N_A_923_74#_c_705_n 0.00374122f $X=-0.19 $Y=-0.245 $X2=2.26 $Y2=1.765
cc_58 VNB N_A_923_74#_c_706_n 0.00643668f $X=-0.19 $Y=-0.245 $X2=2.26 $Y2=2.4
cc_59 VNB N_A_923_74#_c_707_n 0.002345f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=1.58
cc_60 VNB N_A_923_74#_c_708_n 0.00237781f $X=-0.19 $Y=-0.245 $X2=2.075 $Y2=1.58
cc_61 VNB N_A_923_74#_c_709_n 0.002345f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_A_923_74#_c_710_n 0.00237781f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_A_923_74#_c_711_n 0.002345f $X=-0.19 $Y=-0.245 $X2=0.745 $Y2=1.515
cc_64 VNB N_A_923_74#_c_712_n 0.00237781f $X=-0.19 $Y=-0.245 $X2=0.745 $Y2=1.515
cc_65 VNB N_A_923_74#_c_713_n 0.0171072f $X=-0.19 $Y=-0.245 $X2=1.425 $Y2=1.557
cc_66 VPB N_D_c_109_n 0.0106787f $X=-0.19 $Y=1.66 $X2=1.42 $Y2=1.515
cc_67 VPB N_D_c_118_n 0.0183534f $X=-0.19 $Y=1.66 $X2=1.76 $Y2=1.765
cc_68 VPB N_D_c_119_n 0.0155708f $X=-0.19 $Y=1.66 $X2=2.26 $Y2=1.765
cc_69 VPB N_D_c_112_n 0.00517001f $X=-0.19 $Y=1.66 $X2=0.57 $Y2=1.515
cc_70 VPB N_D_c_113_n 0.0106787f $X=-0.19 $Y=1.66 $X2=0.92 $Y2=1.515
cc_71 VPB N_D_c_114_n 0.00459923f $X=-0.19 $Y=1.66 $X2=0.995 $Y2=1.515
cc_72 VPB D 0.024169f $X=-0.19 $Y=1.66 $X2=2.075 $Y2=1.58
cc_73 VPB N_D_c_116_n 0.0300924f $X=-0.19 $Y=1.66 $X2=2.195 $Y2=1.557
cc_74 VPB N_C_c_187_n 0.0174895f $X=-0.19 $Y=1.66 $X2=0.995 $Y2=1.35
cc_75 VPB N_C_c_188_n 0.0212023f $X=-0.19 $Y=1.66 $X2=1.495 $Y2=0.74
cc_76 VPB C 0.0144832f $X=-0.19 $Y=1.66 $X2=0.92 $Y2=1.515
cc_77 VPB N_C_c_186_n 0.0469223f $X=-0.19 $Y=1.66 $X2=1.425 $Y2=1.515
cc_78 VPB N_B_c_245_n 0.0212023f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.35
cc_79 VPB N_B_c_246_n 0.0212309f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_80 VPB B 0.0160103f $X=-0.19 $Y=1.66 $X2=0.92 $Y2=1.515
cc_81 VPB N_B_c_244_n 0.0614899f $X=-0.19 $Y=1.66 $X2=1.425 $Y2=1.515
cc_82 VPB N_A_c_311_n 0.0239877f $X=-0.19 $Y=1.66 $X2=1.42 $Y2=1.515
cc_83 VPB N_A_c_312_n 0.0222993f $X=-0.19 $Y=1.66 $X2=1.76 $Y2=2.4
cc_84 VPB N_A_c_308_n 0.0125229f $X=-0.19 $Y=1.66 $X2=2.26 $Y2=2.4
cc_85 VPB N_A_c_309_n 0.00761063f $X=-0.19 $Y=1.66 $X2=2.26 $Y2=2.4
cc_86 VPB A 0.0124939f $X=-0.19 $Y=1.66 $X2=0.995 $Y2=1.515
cc_87 VPB N_A_c_310_n 0.0335201f $X=-0.19 $Y=1.66 $X2=1.595 $Y2=1.58
cc_88 VPB N_VPWR_c_373_n 0.00341267f $X=-0.19 $Y=1.66 $X2=2.195 $Y2=1.35
cc_89 VPB N_VPWR_c_374_n 0.0251016f $X=-0.19 $Y=1.66 $X2=2.195 $Y2=0.74
cc_90 VPB N_VPWR_c_375_n 0.00934483f $X=-0.19 $Y=1.66 $X2=2.26 $Y2=2.4
cc_91 VPB N_VPWR_c_376_n 0.0121701f $X=-0.19 $Y=1.66 $X2=0.92 $Y2=1.515
cc_92 VPB N_VPWR_c_377_n 0.0356672f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_93 VPB N_VPWR_c_378_n 0.0185368f $X=-0.19 $Y=1.66 $X2=2.075 $Y2=1.58
cc_94 VPB N_VPWR_c_379_n 0.103552f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_95 VPB N_VPWR_c_380_n 0.027658f $X=-0.19 $Y=1.66 $X2=1.425 $Y2=1.515
cc_96 VPB N_VPWR_c_381_n 0.00601644f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_97 VPB N_VPWR_c_382_n 0.0169248f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_98 VPB N_VPWR_c_383_n 0.0251007f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_99 VPB N_VPWR_c_384_n 0.0498007f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_100 VPB N_VPWR_c_372_n 0.076164f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_101 VPB N_Y_c_443_n 0.00289722f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_102 VPB N_Y_c_444_n 0.00587674f $X=-0.19 $Y=1.66 $X2=0.995 $Y2=1.515
cc_103 VPB N_Y_c_445_n 0.00587584f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_104 VPB N_Y_c_446_n 0.00663864f $X=-0.19 $Y=1.66 $X2=1.425 $Y2=1.557
cc_105 VPB N_Y_c_447_n 0.00714919f $X=-0.19 $Y=1.66 $X2=1.76 $Y2=1.557
cc_106 VPB Y 0.0129336f $X=-0.19 $Y=1.66 $X2=2.16 $Y2=1.565
cc_107 N_D_M1020_g N_C_M1002_g 0.0255149f $X=2.195 $Y=0.74 $X2=0 $Y2=0
cc_108 N_D_c_119_n N_C_c_187_n 0.0263918f $X=2.26 $Y=1.765 $X2=0 $Y2=0
cc_109 D C 0.0285068f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_110 N_D_c_116_n C 0.00356538f $X=2.195 $Y=1.557 $X2=0 $Y2=0
cc_111 D N_C_c_186_n 4.01904e-19 $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_112 N_D_c_116_n N_C_c_186_n 0.0195606f $X=2.195 $Y=1.557 $X2=0 $Y2=0
cc_113 N_D_c_118_n N_VPWR_c_373_n 5.12099e-19 $X=1.76 $Y=1.765 $X2=0 $Y2=0
cc_114 N_D_c_119_n N_VPWR_c_373_n 0.0107539f $X=2.26 $Y=1.765 $X2=0 $Y2=0
cc_115 N_D_c_118_n N_VPWR_c_378_n 0.00445602f $X=1.76 $Y=1.765 $X2=0 $Y2=0
cc_116 N_D_c_119_n N_VPWR_c_378_n 0.00413917f $X=2.26 $Y=1.765 $X2=0 $Y2=0
cc_117 N_D_c_118_n N_VPWR_c_379_n 0.00400188f $X=1.76 $Y=1.765 $X2=0 $Y2=0
cc_118 N_D_c_112_n N_VPWR_c_379_n 0.00744949f $X=0.57 $Y=1.515 $X2=0 $Y2=0
cc_119 D N_VPWR_c_379_n 0.133836f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_120 N_D_c_118_n N_VPWR_c_372_n 0.00862158f $X=1.76 $Y=1.765 $X2=0 $Y2=0
cc_121 N_D_c_119_n N_VPWR_c_372_n 0.00818187f $X=2.26 $Y=1.765 $X2=0 $Y2=0
cc_122 N_D_c_118_n N_Y_c_449_n 0.00189972f $X=1.76 $Y=1.765 $X2=0 $Y2=0
cc_123 D N_Y_c_449_n 0.025478f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_124 N_D_c_116_n N_Y_c_449_n 0.00168024f $X=2.195 $Y=1.557 $X2=0 $Y2=0
cc_125 N_D_c_118_n N_Y_c_443_n 0.00902981f $X=1.76 $Y=1.765 $X2=0 $Y2=0
cc_126 N_D_c_119_n N_Y_c_443_n 0.00464047f $X=2.26 $Y=1.765 $X2=0 $Y2=0
cc_127 N_D_c_119_n N_Y_c_454_n 0.0168344f $X=2.26 $Y=1.765 $X2=0 $Y2=0
cc_128 D N_Y_c_454_n 0.0080834f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_129 N_D_M1008_g N_A_27_74#_c_535_n 0.0102216f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_130 N_D_M1010_g N_A_27_74#_c_535_n 6.38603e-19 $X=0.995 $Y=0.74 $X2=0 $Y2=0
cc_131 N_D_M1008_g N_A_27_74#_c_536_n 0.0115433f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_132 N_D_M1010_g N_A_27_74#_c_536_n 0.0151263f $X=0.995 $Y=0.74 $X2=0 $Y2=0
cc_133 N_D_c_113_n N_A_27_74#_c_536_n 0.00381149f $X=0.92 $Y=1.515 $X2=0 $Y2=0
cc_134 D N_A_27_74#_c_536_n 0.0501792f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_135 N_D_M1008_g N_A_27_74#_c_537_n 0.00214722f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_136 D N_A_27_74#_c_537_n 0.0286342f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_137 N_D_M1010_g N_A_27_74#_c_538_n 0.00350341f $X=0.995 $Y=0.74 $X2=0 $Y2=0
cc_138 N_D_M1014_g N_A_27_74#_c_538_n 0.010082f $X=1.495 $Y=0.74 $X2=0 $Y2=0
cc_139 N_D_M1020_g N_A_27_74#_c_538_n 7.91979e-19 $X=2.195 $Y=0.74 $X2=0 $Y2=0
cc_140 N_D_M1014_g N_A_27_74#_c_539_n 0.0123334f $X=1.495 $Y=0.74 $X2=0 $Y2=0
cc_141 N_D_M1020_g N_A_27_74#_c_539_n 0.013916f $X=2.195 $Y=0.74 $X2=0 $Y2=0
cc_142 D N_A_27_74#_c_539_n 0.062829f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_143 N_D_c_116_n N_A_27_74#_c_539_n 0.0126414f $X=2.195 $Y=1.557 $X2=0 $Y2=0
cc_144 N_D_M1020_g N_A_27_74#_c_540_n 0.00502264f $X=2.195 $Y=0.74 $X2=0 $Y2=0
cc_145 N_D_M1014_g N_A_27_74#_c_559_n 7.59304e-19 $X=1.495 $Y=0.74 $X2=0 $Y2=0
cc_146 N_D_M1020_g N_A_27_74#_c_559_n 0.00666311f $X=2.195 $Y=0.74 $X2=0 $Y2=0
cc_147 N_D_c_109_n N_A_27_74#_c_542_n 0.00396026f $X=1.42 $Y=1.515 $X2=0 $Y2=0
cc_148 N_D_M1014_g N_A_27_74#_c_542_n 0.00173883f $X=1.495 $Y=0.74 $X2=0 $Y2=0
cc_149 D N_A_27_74#_c_542_n 0.0281948f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_150 N_D_M1008_g N_VGND_c_597_n 0.00571035f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_151 N_D_M1010_g N_VGND_c_597_n 0.0109084f $X=0.995 $Y=0.74 $X2=0 $Y2=0
cc_152 N_D_M1014_g N_VGND_c_597_n 4.99121e-19 $X=1.495 $Y=0.74 $X2=0 $Y2=0
cc_153 N_D_M1010_g N_VGND_c_598_n 0.00383152f $X=0.995 $Y=0.74 $X2=0 $Y2=0
cc_154 N_D_M1014_g N_VGND_c_598_n 0.00434272f $X=1.495 $Y=0.74 $X2=0 $Y2=0
cc_155 N_D_M1014_g N_VGND_c_599_n 0.00572004f $X=1.495 $Y=0.74 $X2=0 $Y2=0
cc_156 N_D_M1020_g N_VGND_c_599_n 0.00777206f $X=2.195 $Y=0.74 $X2=0 $Y2=0
cc_157 N_D_M1008_g N_VGND_c_600_n 0.00434272f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_158 N_D_M1020_g N_VGND_c_601_n 0.00433139f $X=2.195 $Y=0.74 $X2=0 $Y2=0
cc_159 N_D_M1008_g N_VGND_c_602_n 0.00824376f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_160 N_D_M1010_g N_VGND_c_602_n 0.00758198f $X=0.995 $Y=0.74 $X2=0 $Y2=0
cc_161 N_D_M1014_g N_VGND_c_602_n 0.00822835f $X=1.495 $Y=0.74 $X2=0 $Y2=0
cc_162 N_D_M1020_g N_VGND_c_602_n 0.0082043f $X=2.195 $Y=0.74 $X2=0 $Y2=0
cc_163 C B 0.0305568f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_164 N_C_c_186_n B 0.00116481f $X=3.805 $Y=1.515 $X2=0 $Y2=0
cc_165 C N_B_c_244_n 0.00207029f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_166 N_C_c_186_n N_B_c_244_n 0.00895304f $X=3.805 $Y=1.515 $X2=0 $Y2=0
cc_167 N_C_c_187_n N_VPWR_c_373_n 0.013525f $X=2.71 $Y=1.765 $X2=0 $Y2=0
cc_168 N_C_c_187_n N_VPWR_c_374_n 0.00413917f $X=2.71 $Y=1.765 $X2=0 $Y2=0
cc_169 N_C_c_188_n N_VPWR_c_374_n 0.00413917f $X=3.54 $Y=1.765 $X2=0 $Y2=0
cc_170 N_C_c_188_n N_VPWR_c_375_n 0.0156654f $X=3.54 $Y=1.765 $X2=0 $Y2=0
cc_171 N_C_c_187_n N_VPWR_c_372_n 0.00820334f $X=2.71 $Y=1.765 $X2=0 $Y2=0
cc_172 N_C_c_188_n N_VPWR_c_372_n 0.00820334f $X=3.54 $Y=1.765 $X2=0 $Y2=0
cc_173 N_C_c_187_n N_Y_c_454_n 0.0126342f $X=2.71 $Y=1.765 $X2=0 $Y2=0
cc_174 C N_Y_c_454_n 0.0191189f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_175 N_C_c_187_n N_Y_c_444_n 3.44078e-19 $X=2.71 $Y=1.765 $X2=0 $Y2=0
cc_176 N_C_c_188_n N_Y_c_444_n 3.44078e-19 $X=3.54 $Y=1.765 $X2=0 $Y2=0
cc_177 N_C_c_188_n N_Y_c_460_n 0.0146058f $X=3.54 $Y=1.765 $X2=0 $Y2=0
cc_178 C N_Y_c_460_n 0.0565548f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_179 N_C_c_186_n N_Y_c_460_n 0.00224564f $X=3.805 $Y=1.515 $X2=0 $Y2=0
cc_180 C N_Y_c_463_n 0.0519473f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_181 N_C_c_186_n N_Y_c_463_n 0.0036208f $X=3.805 $Y=1.515 $X2=0 $Y2=0
cc_182 N_C_M1002_g N_A_27_74#_c_539_n 0.00237285f $X=2.695 $Y=0.74 $X2=0 $Y2=0
cc_183 C N_A_27_74#_c_539_n 0.00450841f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_184 N_C_M1002_g N_A_27_74#_c_541_n 0.0186789f $X=2.695 $Y=0.74 $X2=0 $Y2=0
cc_185 N_C_M1011_g N_A_27_74#_c_541_n 0.0123211f $X=3.125 $Y=0.74 $X2=0 $Y2=0
cc_186 N_C_M1012_g N_A_27_74#_c_541_n 0.0123211f $X=3.555 $Y=0.74 $X2=0 $Y2=0
cc_187 N_C_M1021_g N_A_27_74#_c_541_n 0.0126246f $X=3.985 $Y=0.74 $X2=0 $Y2=0
cc_188 C N_A_27_74#_c_541_n 0.00379054f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_189 N_C_M1002_g N_VGND_c_601_n 0.00291649f $X=2.695 $Y=0.74 $X2=0 $Y2=0
cc_190 N_C_M1011_g N_VGND_c_601_n 0.00291649f $X=3.125 $Y=0.74 $X2=0 $Y2=0
cc_191 N_C_M1012_g N_VGND_c_601_n 0.00291649f $X=3.555 $Y=0.74 $X2=0 $Y2=0
cc_192 N_C_M1021_g N_VGND_c_601_n 0.00291649f $X=3.985 $Y=0.74 $X2=0 $Y2=0
cc_193 N_C_M1002_g N_VGND_c_602_n 0.00359833f $X=2.695 $Y=0.74 $X2=0 $Y2=0
cc_194 N_C_M1011_g N_VGND_c_602_n 0.00359121f $X=3.125 $Y=0.74 $X2=0 $Y2=0
cc_195 N_C_M1012_g N_VGND_c_602_n 0.00359121f $X=3.555 $Y=0.74 $X2=0 $Y2=0
cc_196 N_C_M1021_g N_VGND_c_602_n 0.0036412f $X=3.985 $Y=0.74 $X2=0 $Y2=0
cc_197 N_C_M1002_g N_A_554_74#_c_665_n 0.00380276f $X=2.695 $Y=0.74 $X2=0 $Y2=0
cc_198 N_C_M1011_g N_A_554_74#_c_665_n 0.0119209f $X=3.125 $Y=0.74 $X2=0 $Y2=0
cc_199 N_C_M1012_g N_A_554_74#_c_665_n 0.0119209f $X=3.555 $Y=0.74 $X2=0 $Y2=0
cc_200 C N_A_554_74#_c_665_n 0.0936883f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_201 N_C_c_186_n N_A_554_74#_c_665_n 0.00659531f $X=3.805 $Y=1.515 $X2=0 $Y2=0
cc_202 N_C_M1021_g N_A_554_74#_c_667_n 0.00288027f $X=3.985 $Y=0.74 $X2=0 $Y2=0
cc_203 N_C_M1021_g N_A_554_74#_c_668_n 0.0127268f $X=3.985 $Y=0.74 $X2=0 $Y2=0
cc_204 N_C_M1021_g N_A_923_74#_c_706_n 6.08634e-19 $X=3.985 $Y=0.74 $X2=0 $Y2=0
cc_205 N_B_M1022_g N_A_M1005_g 0.0255996f $X=6.265 $Y=0.74 $X2=0 $Y2=0
cc_206 B A 0.0140912f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_207 N_B_c_244_n A 0.00131406f $X=5.995 $Y=1.515 $X2=0 $Y2=0
cc_208 B N_A_c_310_n 0.00116053f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_209 N_B_c_244_n N_A_c_310_n 0.0255996f $X=5.995 $Y=1.515 $X2=0 $Y2=0
cc_210 N_B_c_245_n N_VPWR_c_375_n 0.0156654f $X=4.56 $Y=1.765 $X2=0 $Y2=0
cc_211 N_B_c_245_n N_VPWR_c_383_n 0.00413917f $X=4.56 $Y=1.765 $X2=0 $Y2=0
cc_212 N_B_c_246_n N_VPWR_c_383_n 0.00413917f $X=5.39 $Y=1.765 $X2=0 $Y2=0
cc_213 N_B_c_246_n N_VPWR_c_384_n 0.0157296f $X=5.39 $Y=1.765 $X2=0 $Y2=0
cc_214 N_B_c_245_n N_VPWR_c_372_n 0.00820334f $X=4.56 $Y=1.765 $X2=0 $Y2=0
cc_215 N_B_c_246_n N_VPWR_c_372_n 0.00815719f $X=5.39 $Y=1.765 $X2=0 $Y2=0
cc_216 N_B_c_245_n N_Y_c_460_n 0.0146058f $X=4.56 $Y=1.765 $X2=0 $Y2=0
cc_217 B N_Y_c_460_n 0.0141607f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_218 N_B_c_245_n N_Y_c_445_n 3.44078e-19 $X=4.56 $Y=1.765 $X2=0 $Y2=0
cc_219 N_B_c_246_n N_Y_c_445_n 3.43681e-19 $X=5.39 $Y=1.765 $X2=0 $Y2=0
cc_220 N_B_c_246_n N_Y_c_469_n 0.0145759f $X=5.39 $Y=1.765 $X2=0 $Y2=0
cc_221 B N_Y_c_469_n 0.0657145f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_222 N_B_c_244_n N_Y_c_469_n 0.0103104f $X=5.995 $Y=1.515 $X2=0 $Y2=0
cc_223 N_B_M1022_g N_Y_c_438_n 7.32989e-19 $X=6.265 $Y=0.74 $X2=0 $Y2=0
cc_224 B N_Y_c_473_n 0.0519473f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_225 N_B_c_244_n N_Y_c_473_n 0.00362999f $X=5.995 $Y=1.515 $X2=0 $Y2=0
cc_226 N_B_M1006_g N_A_27_74#_c_541_n 7.21241e-19 $X=4.975 $Y=0.74 $X2=0 $Y2=0
cc_227 N_B_M1006_g N_VGND_c_601_n 0.00292759f $X=4.975 $Y=0.74 $X2=0 $Y2=0
cc_228 N_B_M1007_g N_VGND_c_601_n 0.00291649f $X=5.405 $Y=0.74 $X2=0 $Y2=0
cc_229 N_B_M1018_g N_VGND_c_601_n 0.00291649f $X=5.835 $Y=0.74 $X2=0 $Y2=0
cc_230 N_B_M1022_g N_VGND_c_601_n 0.00291649f $X=6.265 $Y=0.74 $X2=0 $Y2=0
cc_231 N_B_M1006_g N_VGND_c_602_n 0.00363156f $X=4.975 $Y=0.74 $X2=0 $Y2=0
cc_232 N_B_M1007_g N_VGND_c_602_n 0.00359121f $X=5.405 $Y=0.74 $X2=0 $Y2=0
cc_233 N_B_M1018_g N_VGND_c_602_n 0.00359121f $X=5.835 $Y=0.74 $X2=0 $Y2=0
cc_234 N_B_M1022_g N_VGND_c_602_n 0.00359219f $X=6.265 $Y=0.74 $X2=0 $Y2=0
cc_235 N_B_M1007_g N_A_554_74#_c_666_n 0.0120015f $X=5.405 $Y=0.74 $X2=0 $Y2=0
cc_236 N_B_M1018_g N_A_554_74#_c_666_n 0.0131801f $X=5.835 $Y=0.74 $X2=0 $Y2=0
cc_237 N_B_M1022_g N_A_554_74#_c_666_n 0.00620273f $X=6.265 $Y=0.74 $X2=0 $Y2=0
cc_238 B N_A_554_74#_c_666_n 0.0136738f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_239 N_B_c_244_n N_A_554_74#_c_666_n 0.00440417f $X=5.995 $Y=1.515 $X2=0 $Y2=0
cc_240 N_B_M1006_g N_A_554_74#_c_668_n 0.0149988f $X=4.975 $Y=0.74 $X2=0 $Y2=0
cc_241 B N_A_554_74#_c_668_n 0.0967792f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_242 N_B_c_244_n N_A_554_74#_c_668_n 0.010017f $X=5.995 $Y=1.515 $X2=0 $Y2=0
cc_243 N_B_c_244_n N_A_554_74#_c_669_n 0.00221025f $X=5.995 $Y=1.515 $X2=0 $Y2=0
cc_244 N_B_M1006_g N_A_923_74#_c_706_n 0.00509819f $X=4.975 $Y=0.74 $X2=0 $Y2=0
cc_245 N_B_M1007_g N_A_923_74#_c_706_n 6.42481e-19 $X=5.405 $Y=0.74 $X2=0 $Y2=0
cc_246 N_B_M1006_g N_A_923_74#_c_707_n 0.00833016f $X=4.975 $Y=0.74 $X2=0 $Y2=0
cc_247 N_B_M1007_g N_A_923_74#_c_707_n 0.00775417f $X=5.405 $Y=0.74 $X2=0 $Y2=0
cc_248 N_B_M1006_g N_A_923_74#_c_708_n 5.57235e-19 $X=4.975 $Y=0.74 $X2=0 $Y2=0
cc_249 N_B_M1007_g N_A_923_74#_c_708_n 0.00449305f $X=5.405 $Y=0.74 $X2=0 $Y2=0
cc_250 N_B_M1018_g N_A_923_74#_c_708_n 0.00448992f $X=5.835 $Y=0.74 $X2=0 $Y2=0
cc_251 N_B_M1022_g N_A_923_74#_c_708_n 5.57001e-19 $X=6.265 $Y=0.74 $X2=0 $Y2=0
cc_252 N_B_M1018_g N_A_923_74#_c_709_n 0.00674334f $X=5.835 $Y=0.74 $X2=0 $Y2=0
cc_253 N_B_M1022_g N_A_923_74#_c_709_n 0.00792254f $X=6.265 $Y=0.74 $X2=0 $Y2=0
cc_254 N_B_M1018_g N_A_923_74#_c_710_n 5.57001e-19 $X=5.835 $Y=0.74 $X2=0 $Y2=0
cc_255 N_B_M1022_g N_A_923_74#_c_710_n 0.00530316f $X=6.265 $Y=0.74 $X2=0 $Y2=0
cc_256 N_A_c_312_n N_VPWR_c_377_n 0.0149378f $X=8.13 $Y=1.765 $X2=0 $Y2=0
cc_257 N_A_c_311_n N_VPWR_c_380_n 0.00413917f $X=7.2 $Y=1.765 $X2=0 $Y2=0
cc_258 N_A_c_312_n N_VPWR_c_380_n 0.00413917f $X=8.13 $Y=1.765 $X2=0 $Y2=0
cc_259 N_A_c_311_n N_VPWR_c_384_n 0.0159076f $X=7.2 $Y=1.765 $X2=0 $Y2=0
cc_260 N_A_c_311_n N_VPWR_c_372_n 0.00817913f $X=7.2 $Y=1.765 $X2=0 $Y2=0
cc_261 N_A_c_312_n N_VPWR_c_372_n 0.00822528f $X=8.13 $Y=1.765 $X2=0 $Y2=0
cc_262 N_A_c_311_n N_Y_c_469_n 0.0145759f $X=7.2 $Y=1.765 $X2=0 $Y2=0
cc_263 A N_Y_c_469_n 0.0418544f $X=7.835 $Y=1.58 $X2=0 $Y2=0
cc_264 N_A_c_310_n N_Y_c_469_n 0.00623792f $X=7.63 $Y=1.515 $X2=0 $Y2=0
cc_265 N_A_M1005_g N_Y_c_438_n 0.00550051f $X=6.695 $Y=0.74 $X2=0 $Y2=0
cc_266 A N_Y_c_438_n 0.0171684f $X=7.835 $Y=1.58 $X2=0 $Y2=0
cc_267 N_A_c_310_n N_Y_c_438_n 0.00221206f $X=7.63 $Y=1.515 $X2=0 $Y2=0
cc_268 N_A_c_311_n N_Y_c_446_n 6.58986e-19 $X=7.2 $Y=1.765 $X2=0 $Y2=0
cc_269 N_A_c_312_n N_Y_c_446_n 6.59382e-19 $X=8.13 $Y=1.765 $X2=0 $Y2=0
cc_270 N_A_M1023_g N_Y_c_439_n 0.022034f $X=8.145 $Y=0.74 $X2=0 $Y2=0
cc_271 N_A_c_312_n N_Y_c_447_n 0.0176306f $X=8.13 $Y=1.765 $X2=0 $Y2=0
cc_272 A N_Y_c_447_n 0.00410506f $X=7.835 $Y=1.58 $X2=0 $Y2=0
cc_273 A N_Y_c_486_n 0.0599167f $X=7.835 $Y=1.58 $X2=0 $Y2=0
cc_274 N_A_c_310_n N_Y_c_486_n 0.00416405f $X=7.63 $Y=1.515 $X2=0 $Y2=0
cc_275 N_A_M1013_g N_Y_c_440_n 0.0131801f $X=7.125 $Y=0.74 $X2=0 $Y2=0
cc_276 N_A_M1015_g N_Y_c_440_n 0.0159744f $X=7.555 $Y=0.74 $X2=0 $Y2=0
cc_277 N_A_c_308_n N_Y_c_440_n 0.00572844f $X=8.04 $Y=1.515 $X2=0 $Y2=0
cc_278 A N_Y_c_440_n 0.0691561f $X=7.835 $Y=1.58 $X2=0 $Y2=0
cc_279 N_A_c_310_n N_Y_c_440_n 0.00219211f $X=7.63 $Y=1.515 $X2=0 $Y2=0
cc_280 N_A_M1015_g N_Y_c_441_n 0.0019074f $X=7.555 $Y=0.74 $X2=0 $Y2=0
cc_281 N_A_M1023_g N_Y_c_441_n 0.0019074f $X=8.145 $Y=0.74 $X2=0 $Y2=0
cc_282 N_A_c_312_n Y 0.00696042f $X=8.13 $Y=1.765 $X2=0 $Y2=0
cc_283 N_A_M1023_g Y 0.0207492f $X=8.145 $Y=0.74 $X2=0 $Y2=0
cc_284 A Y 0.0308719f $X=7.835 $Y=1.58 $X2=0 $Y2=0
cc_285 N_A_M1005_g N_VGND_c_601_n 0.00291649f $X=6.695 $Y=0.74 $X2=0 $Y2=0
cc_286 N_A_M1013_g N_VGND_c_601_n 0.00291649f $X=7.125 $Y=0.74 $X2=0 $Y2=0
cc_287 N_A_M1015_g N_VGND_c_601_n 0.00291649f $X=7.555 $Y=0.74 $X2=0 $Y2=0
cc_288 N_A_M1023_g N_VGND_c_601_n 0.00292759f $X=8.145 $Y=0.74 $X2=0 $Y2=0
cc_289 N_A_M1005_g N_VGND_c_602_n 0.00359219f $X=6.695 $Y=0.74 $X2=0 $Y2=0
cc_290 N_A_M1013_g N_VGND_c_602_n 0.00359121f $X=7.125 $Y=0.74 $X2=0 $Y2=0
cc_291 N_A_M1015_g N_VGND_c_602_n 0.00360505f $X=7.555 $Y=0.74 $X2=0 $Y2=0
cc_292 N_A_M1023_g N_VGND_c_602_n 0.00363199f $X=8.145 $Y=0.74 $X2=0 $Y2=0
cc_293 N_A_M1005_g N_A_554_74#_c_666_n 7.32989e-19 $X=6.695 $Y=0.74 $X2=0 $Y2=0
cc_294 N_A_M1015_g N_A_923_74#_c_705_n 0.00855567f $X=7.555 $Y=0.74 $X2=0 $Y2=0
cc_295 N_A_M1023_g N_A_923_74#_c_705_n 0.00913165f $X=8.145 $Y=0.74 $X2=0 $Y2=0
cc_296 N_A_M1005_g N_A_923_74#_c_710_n 0.00530316f $X=6.695 $Y=0.74 $X2=0 $Y2=0
cc_297 N_A_M1013_g N_A_923_74#_c_710_n 5.57001e-19 $X=7.125 $Y=0.74 $X2=0 $Y2=0
cc_298 N_A_M1005_g N_A_923_74#_c_711_n 0.00792254f $X=6.695 $Y=0.74 $X2=0 $Y2=0
cc_299 N_A_M1013_g N_A_923_74#_c_711_n 0.00674334f $X=7.125 $Y=0.74 $X2=0 $Y2=0
cc_300 N_A_M1005_g N_A_923_74#_c_712_n 5.57001e-19 $X=6.695 $Y=0.74 $X2=0 $Y2=0
cc_301 N_A_M1013_g N_A_923_74#_c_712_n 0.00448992f $X=7.125 $Y=0.74 $X2=0 $Y2=0
cc_302 N_A_M1015_g N_A_923_74#_c_712_n 0.00510671f $X=7.555 $Y=0.74 $X2=0 $Y2=0
cc_303 N_A_M1023_g N_A_923_74#_c_712_n 8.54686e-19 $X=8.145 $Y=0.74 $X2=0 $Y2=0
cc_304 N_A_M1015_g N_A_923_74#_c_713_n 9.39838e-19 $X=7.555 $Y=0.74 $X2=0 $Y2=0
cc_305 N_A_M1023_g N_A_923_74#_c_713_n 0.00577613f $X=8.145 $Y=0.74 $X2=0 $Y2=0
cc_306 N_VPWR_c_373_n N_Y_c_443_n 0.0266809f $X=2.485 $Y=2.455 $X2=0 $Y2=0
cc_307 N_VPWR_c_378_n N_Y_c_443_n 0.0145938f $X=2.32 $Y=3.33 $X2=0 $Y2=0
cc_308 N_VPWR_c_379_n N_Y_c_443_n 0.0332705f $X=1.65 $Y=3.33 $X2=0 $Y2=0
cc_309 N_VPWR_c_372_n N_Y_c_443_n 0.0120466f $X=8.4 $Y=3.33 $X2=0 $Y2=0
cc_310 N_VPWR_M1017_d N_Y_c_454_n 0.00761668f $X=2.335 $Y=1.84 $X2=0 $Y2=0
cc_311 N_VPWR_c_373_n N_Y_c_454_n 0.0171814f $X=2.485 $Y=2.455 $X2=0 $Y2=0
cc_312 N_VPWR_c_373_n N_Y_c_444_n 0.0267578f $X=2.485 $Y=2.455 $X2=0 $Y2=0
cc_313 N_VPWR_c_374_n N_Y_c_444_n 0.0271295f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_314 N_VPWR_c_375_n N_Y_c_444_n 0.0297957f $X=4.335 $Y=2.415 $X2=0 $Y2=0
cc_315 N_VPWR_c_372_n N_Y_c_444_n 0.0224555f $X=8.4 $Y=3.33 $X2=0 $Y2=0
cc_316 N_VPWR_M1019_d N_Y_c_460_n 0.0264796f $X=3.615 $Y=1.84 $X2=0 $Y2=0
cc_317 N_VPWR_c_375_n N_Y_c_460_n 0.0635557f $X=4.335 $Y=2.415 $X2=0 $Y2=0
cc_318 N_VPWR_c_375_n N_Y_c_445_n 0.0297957f $X=4.335 $Y=2.415 $X2=0 $Y2=0
cc_319 N_VPWR_c_383_n N_Y_c_445_n 0.0271295f $X=5.45 $Y=2.852 $X2=0 $Y2=0
cc_320 N_VPWR_c_384_n N_Y_c_445_n 0.0298945f $X=7.14 $Y=2.852 $X2=0 $Y2=0
cc_321 N_VPWR_c_372_n N_Y_c_445_n 0.0224555f $X=8.4 $Y=3.33 $X2=0 $Y2=0
cc_322 N_VPWR_M1009_s N_Y_c_469_n 0.0513808f $X=5.465 $Y=1.84 $X2=0 $Y2=0
cc_323 N_VPWR_c_384_n N_Y_c_469_n 0.127419f $X=7.14 $Y=2.852 $X2=0 $Y2=0
cc_324 N_VPWR_c_377_n N_Y_c_446_n 0.0255792f $X=8.355 $Y=2.415 $X2=0 $Y2=0
cc_325 N_VPWR_c_380_n N_Y_c_446_n 0.0306992f $X=8.19 $Y=3.33 $X2=0 $Y2=0
cc_326 N_VPWR_c_384_n N_Y_c_446_n 0.0285677f $X=7.14 $Y=2.852 $X2=0 $Y2=0
cc_327 N_VPWR_c_372_n N_Y_c_446_n 0.0254101f $X=8.4 $Y=3.33 $X2=0 $Y2=0
cc_328 N_VPWR_M1004_s N_Y_c_447_n 0.00452356f $X=8.205 $Y=1.84 $X2=0 $Y2=0
cc_329 N_VPWR_c_377_n N_Y_c_447_n 0.0235574f $X=8.355 $Y=2.415 $X2=0 $Y2=0
cc_330 N_VPWR_M1004_s Y 0.00194528f $X=8.205 $Y=1.84 $X2=0 $Y2=0
cc_331 N_Y_c_438_n N_A_554_74#_c_666_n 0.00828756f $X=7.005 $Y=1.005 $X2=0 $Y2=0
cc_332 N_Y_c_440_n N_A_923_74#_M1013_s 0.00179007f $X=7.755 $Y=0.965 $X2=0 $Y2=0
cc_333 N_Y_c_439_n N_A_923_74#_M1023_s 0.0030137f $X=8.285 $Y=1.005 $X2=0 $Y2=0
cc_334 N_Y_M1015_d N_A_923_74#_c_705_n 0.00526523f $X=7.63 $Y=0.37 $X2=0 $Y2=0
cc_335 N_Y_c_439_n N_A_923_74#_c_705_n 0.00768836f $X=8.285 $Y=1.005 $X2=0 $Y2=0
cc_336 N_Y_c_440_n N_A_923_74#_c_705_n 0.00766981f $X=7.755 $Y=0.965 $X2=0 $Y2=0
cc_337 N_Y_c_441_n N_A_923_74#_c_705_n 0.0091307f $X=7.945 $Y=0.965 $X2=0 $Y2=0
cc_338 N_Y_M1005_d N_A_923_74#_c_711_n 0.00221561f $X=6.77 $Y=0.37 $X2=0 $Y2=0
cc_339 N_Y_c_438_n N_A_923_74#_c_711_n 0.00894405f $X=7.005 $Y=1.005 $X2=0 $Y2=0
cc_340 N_Y_c_440_n N_A_923_74#_c_711_n 0.0028488f $X=7.755 $Y=0.965 $X2=0 $Y2=0
cc_341 N_Y_c_440_n N_A_923_74#_c_712_n 0.0167547f $X=7.755 $Y=0.965 $X2=0 $Y2=0
cc_342 N_Y_c_439_n N_A_923_74#_c_713_n 0.0222972f $X=8.285 $Y=1.005 $X2=0 $Y2=0
cc_343 N_A_27_74#_c_536_n N_VGND_M1008_d 0.00250873f $X=1.115 $Y=1.095 $X2=-0.19
+ $Y2=-0.245
cc_344 N_A_27_74#_c_539_n N_VGND_M1014_d 0.00895142f $X=2.245 $Y=1.095 $X2=0
+ $Y2=0
cc_345 N_A_27_74#_c_535_n N_VGND_c_597_n 0.0191765f $X=0.28 $Y=0.515 $X2=0 $Y2=0
cc_346 N_A_27_74#_c_536_n N_VGND_c_597_n 0.0209867f $X=1.115 $Y=1.095 $X2=0
+ $Y2=0
cc_347 N_A_27_74#_c_538_n N_VGND_c_597_n 0.0191765f $X=1.28 $Y=0.515 $X2=0 $Y2=0
cc_348 N_A_27_74#_c_538_n N_VGND_c_598_n 0.0145639f $X=1.28 $Y=0.515 $X2=0 $Y2=0
cc_349 N_A_27_74#_c_538_n N_VGND_c_599_n 0.0191765f $X=1.28 $Y=0.515 $X2=0 $Y2=0
cc_350 N_A_27_74#_c_539_n N_VGND_c_599_n 0.0257907f $X=2.245 $Y=1.095 $X2=0
+ $Y2=0
cc_351 N_A_27_74#_c_540_n N_VGND_c_599_n 0.0175755f $X=2.41 $Y=0.68 $X2=0 $Y2=0
cc_352 N_A_27_74#_c_559_n N_VGND_c_599_n 0.00801271f $X=2.41 $Y=0.965 $X2=0
+ $Y2=0
cc_353 N_A_27_74#_c_535_n N_VGND_c_600_n 0.0145639f $X=0.28 $Y=0.515 $X2=0 $Y2=0
cc_354 N_A_27_74#_c_540_n N_VGND_c_601_n 0.0146502f $X=2.41 $Y=0.68 $X2=0 $Y2=0
cc_355 N_A_27_74#_c_541_n N_VGND_c_601_n 0.0738988f $X=4.2 $Y=0.515 $X2=0 $Y2=0
cc_356 N_A_27_74#_c_535_n N_VGND_c_602_n 0.0119984f $X=0.28 $Y=0.515 $X2=0 $Y2=0
cc_357 N_A_27_74#_c_538_n N_VGND_c_602_n 0.0119984f $X=1.28 $Y=0.515 $X2=0 $Y2=0
cc_358 N_A_27_74#_c_540_n N_VGND_c_602_n 0.0120674f $X=2.41 $Y=0.68 $X2=0 $Y2=0
cc_359 N_A_27_74#_c_541_n N_VGND_c_602_n 0.0616452f $X=4.2 $Y=0.515 $X2=0 $Y2=0
cc_360 N_A_27_74#_c_541_n N_A_554_74#_M1002_d 0.00172862f $X=4.2 $Y=0.515
+ $X2=-0.19 $Y2=-0.245
cc_361 N_A_27_74#_c_541_n N_A_554_74#_M1012_d 0.00172862f $X=4.2 $Y=0.515 $X2=0
+ $Y2=0
cc_362 N_A_27_74#_M1011_s N_A_554_74#_c_665_n 0.00177318f $X=3.2 $Y=0.37 $X2=0
+ $Y2=0
cc_363 N_A_27_74#_c_539_n N_A_554_74#_c_665_n 0.00587942f $X=2.245 $Y=1.095
+ $X2=0 $Y2=0
cc_364 N_A_27_74#_c_541_n N_A_554_74#_c_665_n 0.0636023f $X=4.2 $Y=0.515 $X2=0
+ $Y2=0
cc_365 N_A_27_74#_M1021_s N_A_554_74#_c_668_n 0.00311853f $X=4.06 $Y=0.37 $X2=0
+ $Y2=0
cc_366 N_A_27_74#_c_541_n N_A_554_74#_c_668_n 0.0254477f $X=4.2 $Y=0.515 $X2=0
+ $Y2=0
cc_367 N_A_27_74#_c_541_n N_A_923_74#_c_706_n 0.0234648f $X=4.2 $Y=0.515 $X2=0
+ $Y2=0
cc_368 N_VGND_c_601_n N_A_923_74#_c_706_n 0.0139208f $X=8.4 $Y=0 $X2=0 $Y2=0
cc_369 N_VGND_c_602_n N_A_923_74#_c_706_n 0.0117508f $X=8.4 $Y=0 $X2=0 $Y2=0
cc_370 N_VGND_c_601_n N_A_923_74#_c_707_n 0.131762f $X=8.4 $Y=0 $X2=0 $Y2=0
cc_371 N_VGND_c_602_n N_A_923_74#_c_707_n 0.111189f $X=8.4 $Y=0 $X2=0 $Y2=0
cc_372 N_VGND_c_601_n N_A_923_74#_c_713_n 0.0139208f $X=8.4 $Y=0 $X2=0 $Y2=0
cc_373 N_VGND_c_602_n N_A_923_74#_c_713_n 0.0117508f $X=8.4 $Y=0 $X2=0 $Y2=0
cc_374 N_A_554_74#_c_668_n N_A_923_74#_M1006_d 0.00296342f $X=5.095 $Y=0.965
+ $X2=-0.19 $Y2=-0.245
cc_375 N_A_554_74#_c_666_n N_A_923_74#_M1007_d 0.00179007f $X=5.955 $Y=1.005
+ $X2=0 $Y2=0
cc_376 N_A_554_74#_c_668_n N_A_923_74#_c_706_n 0.0214875f $X=5.095 $Y=0.965
+ $X2=0 $Y2=0
cc_377 N_A_554_74#_M1006_s N_A_923_74#_c_707_n 0.00221951f $X=5.05 $Y=0.37 $X2=0
+ $Y2=0
cc_378 N_A_554_74#_c_666_n N_A_923_74#_c_707_n 0.00474257f $X=5.955 $Y=1.005
+ $X2=0 $Y2=0
cc_379 N_A_554_74#_c_668_n N_A_923_74#_c_707_n 0.00476112f $X=5.095 $Y=0.965
+ $X2=0 $Y2=0
cc_380 N_A_554_74#_c_669_n N_A_923_74#_c_707_n 0.00797735f $X=5.285 $Y=0.965
+ $X2=0 $Y2=0
cc_381 N_A_554_74#_c_666_n N_A_923_74#_c_708_n 0.0167547f $X=5.955 $Y=1.005
+ $X2=0 $Y2=0
cc_382 N_A_554_74#_M1018_s N_A_923_74#_c_709_n 0.00221561f $X=5.91 $Y=0.37 $X2=0
+ $Y2=0
cc_383 N_A_554_74#_c_666_n N_A_923_74#_c_709_n 0.0117928f $X=5.955 $Y=1.005
+ $X2=0 $Y2=0
