* File: sky130_fd_sc_hs__o221a_4.spice
* Created: Tue Sep  1 20:15:38 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hs__o221a_4.pex.spice"
.subckt sky130_fd_sc_hs__o221a_4  VNB VPB C1 B2 B1 A2 A1 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A1	A1
* A2	A2
* B1	B1
* B2	B2
* C1	C1
* VPB	VPB
* VNB	VNB
MM1016 N_A_27_125#_M1016_d N_C1_M1016_g N_A_114_125#_M1016_s VNB NLOWVT L=0.15
+ W=0.64 AD=0.1824 AS=0.0896 PD=1.85 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75002.5 A=0.096 P=1.58 MULT=1
MM1017 N_A_27_125#_M1017_d N_C1_M1017_g N_A_114_125#_M1016_s VNB NLOWVT L=0.15
+ W=0.64 AD=0.112 AS=0.0896 PD=0.99 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667 SA=75000.6
+ SB=75002.1 A=0.096 P=1.58 MULT=1
MM1002 N_A_27_125#_M1017_d N_B1_M1002_g N_A_300_125#_M1002_s VNB NLOWVT L=0.15
+ W=0.64 AD=0.112 AS=0.1008 PD=0.99 PS=0.955 NRD=13.116 NRS=0 M=1 R=4.26667
+ SA=75001.1 SB=75001.6 A=0.096 P=1.58 MULT=1
MM1007 N_A_300_125#_M1002_s N_B2_M1007_g N_A_27_125#_M1007_s VNB NLOWVT L=0.15
+ W=0.64 AD=0.1008 AS=0.1008 PD=0.955 PS=0.955 NRD=6.552 NRS=6.552 M=1 R=4.26667
+ SA=75001.6 SB=75001.1 A=0.096 P=1.58 MULT=1
MM1023 N_A_300_125#_M1023_d N_B2_M1023_g N_A_27_125#_M1007_s VNB NLOWVT L=0.15
+ W=0.64 AD=0.0912 AS=0.1008 PD=0.925 PS=0.955 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75002.1 SB=75000.6 A=0.096 P=1.58 MULT=1
MM1015 N_A_27_125#_M1015_d N_B1_M1015_g N_A_300_125#_M1023_d VNB NLOWVT L=0.15
+ W=0.64 AD=0.1824 AS=0.0912 PD=1.85 PS=0.925 NRD=0 NRS=0.936 M=1 R=4.26667
+ SA=75002.5 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1012 N_VGND_M1012_d N_A1_M1012_g N_A_300_125#_M1012_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.1824 AS=0.0912 PD=1.85 PS=0.925 NRD=0 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75003.6 A=0.096 P=1.58 MULT=1
MM1013 N_VGND_M1013_d N_A2_M1013_g N_A_300_125#_M1012_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.0896 AS=0.0912 PD=0.92 PS=0.925 NRD=0 NRS=0.936 M=1 R=4.26667 SA=75000.6
+ SB=75003.1 A=0.096 P=1.58 MULT=1
MM1014 N_VGND_M1013_d N_A2_M1014_g N_A_300_125#_M1014_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.0896 AS=0.0896 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667 SA=75001.1
+ SB=75002.7 A=0.096 P=1.58 MULT=1
MM1018 N_VGND_M1018_d N_A1_M1018_g N_A_300_125#_M1014_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.142377 AS=0.0896 PD=1.08058 PS=0.92 NRD=15.468 NRS=0 M=1 R=4.26667
+ SA=75001.5 SB=75002.3 A=0.096 P=1.58 MULT=1
MM1005 N_VGND_M1018_d N_A_114_125#_M1005_g N_X_M1005_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.164623 AS=0.10545 PD=1.24942 PS=1.025 NRD=10.536 NRS=0.804 M=1 R=4.93333
+ SA=75001.8 SB=75001.7 A=0.111 P=1.78 MULT=1
MM1010 N_VGND_M1010_d N_A_114_125#_M1010_g N_X_M1005_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1554 AS=0.10545 PD=1.16 PS=1.025 NRD=5.664 NRS=0 M=1 R=4.93333 SA=75002.3
+ SB=75001.3 A=0.111 P=1.78 MULT=1
MM1021 N_VGND_M1010_d N_A_114_125#_M1021_g N_X_M1021_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1554 AS=0.1036 PD=1.16 PS=1.02 NRD=17.016 NRS=0 M=1 R=4.93333 SA=75002.8
+ SB=75000.7 A=0.111 P=1.78 MULT=1
MM1027 N_VGND_M1027_d N_A_114_125#_M1027_g N_X_M1021_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.2627 AS=0.1036 PD=2.19 PS=1.02 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75003.3
+ SB=75000.3 A=0.111 P=1.78 MULT=1
MM1024 N_A_114_125#_M1024_d N_C1_M1024_g N_VPWR_M1024_s VPB PSHORT L=0.15 W=1
+ AD=0.15 AS=0.295 PD=1.3 PS=2.59 NRD=1.9503 NRS=1.9503 M=1 R=6.66667 SA=75000.2
+ SB=75006.9 A=0.15 P=2.3 MULT=1
MM1025 N_A_114_125#_M1024_d N_C1_M1025_g N_VPWR_M1025_s VPB PSHORT L=0.15 W=1
+ AD=0.15 AS=0.1525 PD=1.3 PS=1.305 NRD=1.9503 NRS=1.9503 M=1 R=6.66667
+ SA=75000.7 SB=75006.4 A=0.15 P=2.3 MULT=1
MM1003 N_VPWR_M1025_s N_B1_M1003_g N_A_297_387#_M1003_s VPB PSHORT L=0.15 W=1
+ AD=0.1525 AS=0.1725 PD=1.305 PS=1.345 NRD=2.9353 NRS=10.8153 M=1 R=6.66667
+ SA=75001.1 SB=75006 A=0.15 P=2.3 MULT=1
MM1000 N_A_114_125#_M1000_d N_B2_M1000_g N_A_297_387#_M1003_s VPB PSHORT L=0.15
+ W=1 AD=0.15 AS=0.1725 PD=1.3 PS=1.345 NRD=1.9503 NRS=1.9503 M=1 R=6.66667
+ SA=75001.6 SB=75005.5 A=0.15 P=2.3 MULT=1
MM1001 N_A_114_125#_M1000_d N_B2_M1001_g N_A_297_387#_M1001_s VPB PSHORT L=0.15
+ W=1 AD=0.15 AS=0.15 PD=1.3 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=6.66667
+ SA=75002.1 SB=75005 A=0.15 P=2.3 MULT=1
MM1019 N_VPWR_M1019_d N_B1_M1019_g N_A_297_387#_M1001_s VPB PSHORT L=0.15 W=1
+ AD=0.3925 AS=0.15 PD=1.785 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=6.66667
+ SA=75002.5 SB=75004.6 A=0.15 P=2.3 MULT=1
MM1004 N_VPWR_M1019_d N_A1_M1004_g N_A_763_387#_M1004_s VPB PSHORT L=0.15 W=1
+ AD=0.3925 AS=0.1625 PD=1.785 PS=1.325 NRD=1.9503 NRS=1.9503 M=1 R=6.66667
+ SA=75003.5 SB=75003.7 A=0.15 P=2.3 MULT=1
MM1020 N_A_114_125#_M1020_d N_A2_M1020_g N_A_763_387#_M1004_s VPB PSHORT L=0.15
+ W=1 AD=0.1625 AS=0.1625 PD=1.325 PS=1.325 NRD=6.8753 NRS=6.8753 M=1 R=6.66667
+ SA=75003.9 SB=75003.2 A=0.15 P=2.3 MULT=1
MM1026 N_A_114_125#_M1020_d N_A2_M1026_g N_A_763_387#_M1026_s VPB PSHORT L=0.15
+ W=1 AD=0.1625 AS=0.175 PD=1.325 PS=1.35 NRD=1.9503 NRS=11.8003 M=1 R=6.66667
+ SA=75004.4 SB=75002.7 A=0.15 P=2.3 MULT=1
MM1022 N_VPWR_M1022_d N_A1_M1022_g N_A_763_387#_M1026_s VPB PSHORT L=0.15 W=1
+ AD=0.182453 AS=0.175 PD=1.39151 PS=1.35 NRD=11.8003 NRS=1.9503 M=1 R=6.66667
+ SA=75004.9 SB=75002.2 A=0.15 P=2.3 MULT=1
MM1006 N_VPWR_M1022_d N_A_114_125#_M1006_g N_X_M1006_s VPB PSHORT L=0.15 W=1.12
+ AD=0.204347 AS=0.21 PD=1.55849 PS=1.495 NRD=2.6201 NRS=14.9326 M=1 R=7.46667
+ SA=75004.9 SB=75001.7 A=0.168 P=2.54 MULT=1
MM1008 N_VPWR_M1008_d N_A_114_125#_M1008_g N_X_M1006_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.21 PD=1.42 PS=1.495 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75005.4 SB=75001.2 A=0.168 P=2.54 MULT=1
MM1009 N_VPWR_M1008_d N_A_114_125#_M1009_g N_X_M1009_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.1988 PD=1.42 PS=1.475 NRD=1.7533 NRS=11.426 M=1 R=7.46667
+ SA=75005.8 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1011 N_VPWR_M1011_d N_A_114_125#_M1011_g N_X_M1009_s VPB PSHORT L=0.15 W=1.12
+ AD=0.3304 AS=0.1988 PD=2.83 PS=1.475 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75006.3 SB=75000.2 A=0.168 P=2.54 MULT=1
DX28_noxref VNB VPB NWDIODE A=14.9916 P=19.84
c_141 VPB 0 1.22796e-19 $X=0 $Y=3.085
*
.include "sky130_fd_sc_hs__o221a_4.pxi.spice"
*
.ends
*
*
