* File: sky130_fd_sc_hs__o41a_1.pxi.spice
* Created: Thu Aug 27 21:04:08 2020
* 
x_PM_SKY130_FD_SC_HS__O41A_1%A_83_270# N_A_83_270#_M1004_s N_A_83_270#_M1006_d
+ N_A_83_270#_M1010_g N_A_83_270#_c_70_n N_A_83_270#_M1005_g N_A_83_270#_c_75_n
+ N_A_83_270#_c_71_n N_A_83_270#_c_72_n N_A_83_270#_c_76_n N_A_83_270#_c_109_p
+ N_A_83_270#_c_73_n N_A_83_270#_c_77_n PM_SKY130_FD_SC_HS__O41A_1%A_83_270#
x_PM_SKY130_FD_SC_HS__O41A_1%B1 N_B1_M1004_g N_B1_c_134_n N_B1_M1006_g B1
+ N_B1_c_135_n PM_SKY130_FD_SC_HS__O41A_1%B1
x_PM_SKY130_FD_SC_HS__O41A_1%A4 N_A4_M1003_g N_A4_c_170_n N_A4_c_171_n
+ N_A4_c_174_n N_A4_M1008_g A4 N_A4_c_172_n PM_SKY130_FD_SC_HS__O41A_1%A4
x_PM_SKY130_FD_SC_HS__O41A_1%A3 N_A3_c_216_n N_A3_M1000_g N_A3_M1011_g A3 A3 A3
+ A3 N_A3_c_218_n PM_SKY130_FD_SC_HS__O41A_1%A3
x_PM_SKY130_FD_SC_HS__O41A_1%A2 N_A2_M1007_g N_A2_c_256_n N_A2_M1002_g A2 A2 A2
+ A2 N_A2_c_257_n PM_SKY130_FD_SC_HS__O41A_1%A2
x_PM_SKY130_FD_SC_HS__O41A_1%A1 N_A1_c_289_n N_A1_M1001_g N_A1_M1009_g A1 A1
+ N_A1_c_291_n PM_SKY130_FD_SC_HS__O41A_1%A1
x_PM_SKY130_FD_SC_HS__O41A_1%X N_X_M1010_s N_X_M1005_s N_X_c_313_n N_X_c_314_n X
+ X N_X_c_315_n X PM_SKY130_FD_SC_HS__O41A_1%X
x_PM_SKY130_FD_SC_HS__O41A_1%VPWR N_VPWR_M1005_d N_VPWR_M1001_d N_VPWR_c_335_n
+ N_VPWR_c_336_n N_VPWR_c_337_n VPWR N_VPWR_c_338_n N_VPWR_c_339_n
+ N_VPWR_c_340_n N_VPWR_c_334_n PM_SKY130_FD_SC_HS__O41A_1%VPWR
x_PM_SKY130_FD_SC_HS__O41A_1%VGND N_VGND_M1010_d N_VGND_M1003_d N_VGND_M1007_d
+ N_VGND_c_379_n N_VGND_c_380_n N_VGND_c_381_n N_VGND_c_382_n N_VGND_c_383_n
+ VGND N_VGND_c_384_n N_VGND_c_385_n N_VGND_c_386_n N_VGND_c_387_n
+ N_VGND_c_388_n N_VGND_c_389_n PM_SKY130_FD_SC_HS__O41A_1%VGND
x_PM_SKY130_FD_SC_HS__O41A_1%A_326_74# N_A_326_74#_M1004_d N_A_326_74#_M1011_d
+ N_A_326_74#_M1009_d N_A_326_74#_c_435_n N_A_326_74#_c_436_n
+ N_A_326_74#_c_437_n N_A_326_74#_c_438_n N_A_326_74#_c_439_n
+ N_A_326_74#_c_440_n N_A_326_74#_c_441_n PM_SKY130_FD_SC_HS__O41A_1%A_326_74#
cc_1 VNB N_A_83_270#_M1010_g 0.0303327f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_2 VNB N_A_83_270#_c_70_n 0.0333324f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.765
cc_3 VNB N_A_83_270#_c_71_n 0.00593596f $X=-0.19 $Y=-0.245 $X2=0.62 $Y2=1.515
cc_4 VNB N_A_83_270#_c_72_n 0.0192328f $X=-0.19 $Y=-0.245 $X2=1.175 $Y2=1.195
cc_5 VNB N_A_83_270#_c_73_n 0.0111398f $X=-0.19 $Y=-0.245 $X2=1.34 $Y2=0.515
cc_6 VNB N_B1_M1004_g 0.042114f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_7 VNB N_B1_c_134_n 0.0229061f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_B1_c_135_n 0.00319006f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_9 VNB N_A4_M1003_g 0.0237112f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A4_c_170_n 0.0332056f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A4_c_171_n 0.0067955f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A4_c_172_n 0.00660497f $X=-0.19 $Y=-0.245 $X2=0.62 $Y2=1.515
cc_13 VNB N_A3_c_216_n 0.0387773f $X=-0.19 $Y=-0.245 $X2=1.195 $Y2=0.37
cc_14 VNB N_A3_M1011_g 0.0253751f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A3_c_218_n 0.00250171f $X=-0.19 $Y=-0.245 $X2=0.62 $Y2=1.515
cc_16 VNB N_A2_M1007_g 0.0309777f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A2_c_256_n 0.032985f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A2_c_257_n 0.00505659f $X=-0.19 $Y=-0.245 $X2=0.62 $Y2=1.515
cc_19 VNB N_A1_c_289_n 0.0305241f $X=-0.19 $Y=-0.245 $X2=1.195 $Y2=0.37
cc_20 VNB N_A1_M1009_g 0.0464113f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A1_c_291_n 0.0184746f $X=-0.19 $Y=-0.245 $X2=0.62 $Y2=1.515
cc_22 VNB N_X_c_313_n 0.0264414f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_23 VNB N_X_c_314_n 0.00871852f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_24 VNB N_X_c_315_n 0.0247491f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_VPWR_c_334_n 0.183584f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_VGND_c_379_n 0.0130175f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_27 VNB N_VGND_c_380_n 0.00900728f $X=-0.19 $Y=-0.245 $X2=0.62 $Y2=1.515
cc_28 VNB N_VGND_c_381_n 0.00814066f $X=-0.19 $Y=-0.245 $X2=0.785 $Y2=1.195
cc_29 VNB N_VGND_c_382_n 0.0339528f $X=-0.19 $Y=-0.245 $X2=1.34 $Y2=1.11
cc_30 VNB N_VGND_c_383_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=1.34 $Y2=0.515
cc_31 VNB N_VGND_c_384_n 0.0173128f $X=-0.19 $Y=-0.245 $X2=1.915 $Y2=2.12
cc_32 VNB N_VGND_c_385_n 0.0185368f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_386_n 0.0191515f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_387_n 0.255913f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_388_n 0.00750435f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_389_n 0.0100141f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_326_74#_c_435_n 0.00280384f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_38 VNB N_A_326_74#_c_436_n 0.00829425f $X=-0.19 $Y=-0.245 $X2=0.62 $Y2=1.515
cc_39 VNB N_A_326_74#_c_437_n 0.00864861f $X=-0.19 $Y=-0.245 $X2=0.62 $Y2=1.95
cc_40 VNB N_A_326_74#_c_438_n 0.00280333f $X=-0.19 $Y=-0.245 $X2=0.62 $Y2=1.515
cc_41 VNB N_A_326_74#_c_439_n 0.0225415f $X=-0.19 $Y=-0.245 $X2=0.785 $Y2=1.195
cc_42 VNB N_A_326_74#_c_440_n 0.0216332f $X=-0.19 $Y=-0.245 $X2=1.34 $Y2=0.515
cc_43 VNB N_A_326_74#_c_441_n 0.00898142f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VPB N_A_83_270#_c_70_n 0.0337329f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.765
cc_45 VPB N_A_83_270#_c_75_n 0.0016796f $X=-0.19 $Y=1.66 $X2=0.62 $Y2=1.95
cc_46 VPB N_A_83_270#_c_76_n 0.0113612f $X=-0.19 $Y=1.66 $X2=1.75 $Y2=2.035
cc_47 VPB N_A_83_270#_c_77_n 3.42873e-19 $X=-0.19 $Y=1.66 $X2=1.915 $Y2=2.13
cc_48 VPB N_B1_c_134_n 0.0527221f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_49 VPB N_B1_c_135_n 0.00256788f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.4
cc_50 VPB N_A4_c_171_n 6.84438e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_51 VPB N_A4_c_174_n 0.0226316f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.35
cc_52 VPB N_A4_c_172_n 0.00584217f $X=-0.19 $Y=1.66 $X2=0.62 $Y2=1.515
cc_53 VPB N_A3_c_216_n 0.0226094f $X=-0.19 $Y=1.66 $X2=1.195 $Y2=0.37
cc_54 VPB N_A3_c_218_n 0.0019602f $X=-0.19 $Y=1.66 $X2=0.62 $Y2=1.515
cc_55 VPB N_A2_c_256_n 0.0236706f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_56 VPB N_A2_c_257_n 0.00255383f $X=-0.19 $Y=1.66 $X2=0.62 $Y2=1.515
cc_57 VPB N_A1_c_289_n 0.0312781f $X=-0.19 $Y=1.66 $X2=1.195 $Y2=0.37
cc_58 VPB N_A1_c_291_n 0.020844f $X=-0.19 $Y=1.66 $X2=0.62 $Y2=1.515
cc_59 VPB X 0.00626527f $X=-0.19 $Y=1.66 $X2=0.62 $Y2=1.515
cc_60 VPB X 0.0226674f $X=-0.19 $Y=1.66 $X2=0.62 $Y2=1.95
cc_61 VPB N_X_c_315_n 0.0240516f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_62 VPB N_VPWR_c_335_n 0.0157896f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.74
cc_63 VPB N_VPWR_c_336_n 0.0142226f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.4
cc_64 VPB N_VPWR_c_337_n 0.0371685f $X=-0.19 $Y=1.66 $X2=0.62 $Y2=1.515
cc_65 VPB N_VPWR_c_338_n 0.0191515f $X=-0.19 $Y=1.66 $X2=0.62 $Y2=1.515
cc_66 VPB N_VPWR_c_339_n 0.0639346f $X=-0.19 $Y=1.66 $X2=1.34 $Y2=1.11
cc_67 VPB N_VPWR_c_340_n 0.0177663f $X=-0.19 $Y=1.66 $X2=0.6 $Y2=1.515
cc_68 VPB N_VPWR_c_334_n 0.0895183f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_69 N_A_83_270#_c_70_n N_B1_M1004_g 0.00112947f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_70 N_A_83_270#_c_71_n N_B1_M1004_g 0.00186326f $X=0.62 $Y=1.515 $X2=0 $Y2=0
cc_71 N_A_83_270#_c_72_n N_B1_M1004_g 0.00743377f $X=1.175 $Y=1.195 $X2=0 $Y2=0
cc_72 N_A_83_270#_c_73_n N_B1_M1004_g 0.0111697f $X=1.34 $Y=0.515 $X2=0 $Y2=0
cc_73 N_A_83_270#_c_70_n N_B1_c_134_n 0.00767667f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_74 N_A_83_270#_c_75_n N_B1_c_134_n 0.00312862f $X=0.62 $Y=1.95 $X2=0 $Y2=0
cc_75 N_A_83_270#_c_72_n N_B1_c_134_n 0.00572457f $X=1.175 $Y=1.195 $X2=0 $Y2=0
cc_76 N_A_83_270#_c_76_n N_B1_c_134_n 0.0286947f $X=1.75 $Y=2.035 $X2=0 $Y2=0
cc_77 N_A_83_270#_c_77_n N_B1_c_134_n 0.00980987f $X=1.915 $Y=2.13 $X2=0 $Y2=0
cc_78 N_A_83_270#_c_70_n N_B1_c_135_n 0.00205993f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_79 N_A_83_270#_c_75_n N_B1_c_135_n 0.0146046f $X=0.62 $Y=1.95 $X2=0 $Y2=0
cc_80 N_A_83_270#_c_71_n N_B1_c_135_n 0.00345372f $X=0.62 $Y=1.515 $X2=0 $Y2=0
cc_81 N_A_83_270#_c_72_n N_B1_c_135_n 0.0351249f $X=1.175 $Y=1.195 $X2=0 $Y2=0
cc_82 N_A_83_270#_c_76_n N_B1_c_135_n 0.0376935f $X=1.75 $Y=2.035 $X2=0 $Y2=0
cc_83 N_A_83_270#_c_72_n N_A4_M1003_g 3.72646e-19 $X=1.175 $Y=1.195 $X2=0 $Y2=0
cc_84 N_A_83_270#_c_73_n N_A4_M1003_g 5.94612e-19 $X=1.34 $Y=0.515 $X2=0 $Y2=0
cc_85 N_A_83_270#_c_72_n N_A4_c_170_n 2.73291e-19 $X=1.175 $Y=1.195 $X2=0 $Y2=0
cc_86 N_A_83_270#_c_76_n N_A4_c_170_n 7.15503e-19 $X=1.75 $Y=2.035 $X2=0 $Y2=0
cc_87 N_A_83_270#_c_76_n N_A4_c_174_n 0.00262338f $X=1.75 $Y=2.035 $X2=0 $Y2=0
cc_88 N_A_83_270#_c_77_n N_A4_c_174_n 0.0125526f $X=1.915 $Y=2.13 $X2=0 $Y2=0
cc_89 N_A_83_270#_c_72_n N_A4_c_172_n 0.00393762f $X=1.175 $Y=1.195 $X2=0 $Y2=0
cc_90 N_A_83_270#_c_76_n N_A4_c_172_n 0.0162867f $X=1.75 $Y=2.035 $X2=0 $Y2=0
cc_91 N_A_83_270#_c_77_n N_A3_c_216_n 7.54461e-19 $X=1.915 $Y=2.13 $X2=-0.19
+ $Y2=-0.245
cc_92 N_A_83_270#_M1010_g N_X_c_313_n 0.00207706f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_93 N_A_83_270#_c_71_n N_X_c_314_n 0.00133215f $X=0.62 $Y=1.515 $X2=0 $Y2=0
cc_94 N_A_83_270#_c_70_n X 0.00231999f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_95 N_A_83_270#_c_70_n X 0.0057471f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_96 N_A_83_270#_M1010_g N_X_c_315_n 0.0047754f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_97 N_A_83_270#_c_70_n N_X_c_315_n 0.022107f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_98 N_A_83_270#_c_75_n N_X_c_315_n 0.0324342f $X=0.62 $Y=1.95 $X2=0 $Y2=0
cc_99 N_A_83_270#_c_71_n N_X_c_315_n 0.0237307f $X=0.62 $Y=1.515 $X2=0 $Y2=0
cc_100 N_A_83_270#_c_109_p N_X_c_315_n 0.0133618f $X=0.785 $Y=2.035 $X2=0 $Y2=0
cc_101 N_A_83_270#_c_75_n N_VPWR_M1005_d 0.00279243f $X=0.62 $Y=1.95 $X2=-0.19
+ $Y2=-0.245
cc_102 N_A_83_270#_c_76_n N_VPWR_M1005_d 0.0127794f $X=1.75 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_103 N_A_83_270#_c_109_p N_VPWR_M1005_d 0.00186198f $X=0.785 $Y=2.035
+ $X2=-0.19 $Y2=-0.245
cc_104 N_A_83_270#_c_70_n N_VPWR_c_335_n 0.0192945f $X=0.505 $Y=1.765 $X2=0
+ $Y2=0
cc_105 N_A_83_270#_c_76_n N_VPWR_c_335_n 0.0565816f $X=1.75 $Y=2.035 $X2=0 $Y2=0
cc_106 N_A_83_270#_c_109_p N_VPWR_c_335_n 0.0132989f $X=0.785 $Y=2.035 $X2=0
+ $Y2=0
cc_107 N_A_83_270#_c_77_n N_VPWR_c_335_n 0.0387143f $X=1.915 $Y=2.13 $X2=0 $Y2=0
cc_108 N_A_83_270#_c_70_n N_VPWR_c_338_n 0.00445602f $X=0.505 $Y=1.765 $X2=0
+ $Y2=0
cc_109 N_A_83_270#_c_77_n N_VPWR_c_339_n 0.00834771f $X=1.915 $Y=2.13 $X2=0
+ $Y2=0
cc_110 N_A_83_270#_c_70_n N_VPWR_c_334_n 0.00865213f $X=0.505 $Y=1.765 $X2=0
+ $Y2=0
cc_111 N_A_83_270#_c_77_n N_VPWR_c_334_n 0.0110052f $X=1.915 $Y=2.13 $X2=0 $Y2=0
cc_112 N_A_83_270#_c_71_n N_VGND_M1010_d 0.00188126f $X=0.62 $Y=1.515 $X2=-0.19
+ $Y2=-0.245
cc_113 N_A_83_270#_M1010_g N_VGND_c_379_n 0.0148187f $X=0.495 $Y=0.74 $X2=0
+ $Y2=0
cc_114 N_A_83_270#_c_70_n N_VGND_c_379_n 7.62615e-19 $X=0.505 $Y=1.765 $X2=0
+ $Y2=0
cc_115 N_A_83_270#_c_71_n N_VGND_c_379_n 0.0166905f $X=0.62 $Y=1.515 $X2=0 $Y2=0
cc_116 N_A_83_270#_c_72_n N_VGND_c_379_n 0.0131435f $X=1.175 $Y=1.195 $X2=0
+ $Y2=0
cc_117 N_A_83_270#_c_73_n N_VGND_c_379_n 0.0403642f $X=1.34 $Y=0.515 $X2=0 $Y2=0
cc_118 N_A_83_270#_c_73_n N_VGND_c_382_n 0.0145639f $X=1.34 $Y=0.515 $X2=0 $Y2=0
cc_119 N_A_83_270#_M1010_g N_VGND_c_384_n 0.00383152f $X=0.495 $Y=0.74 $X2=0
+ $Y2=0
cc_120 N_A_83_270#_M1010_g N_VGND_c_387_n 0.00761198f $X=0.495 $Y=0.74 $X2=0
+ $Y2=0
cc_121 N_A_83_270#_c_73_n N_VGND_c_387_n 0.0119984f $X=1.34 $Y=0.515 $X2=0 $Y2=0
cc_122 N_A_83_270#_c_73_n N_A_326_74#_c_435_n 0.0195517f $X=1.34 $Y=0.515 $X2=0
+ $Y2=0
cc_123 N_A_83_270#_c_73_n N_A_326_74#_c_437_n 0.00682867f $X=1.34 $Y=0.515 $X2=0
+ $Y2=0
cc_124 N_B1_M1004_g N_A4_M1003_g 0.0191404f $X=1.555 $Y=0.69 $X2=0 $Y2=0
cc_125 N_B1_M1004_g N_A4_c_170_n 0.0177663f $X=1.555 $Y=0.69 $X2=0 $Y2=0
cc_126 N_B1_c_135_n N_A4_c_170_n 2.39091e-19 $X=1.415 $Y=1.615 $X2=0 $Y2=0
cc_127 N_B1_c_134_n N_A4_c_171_n 0.00590907f $X=1.605 $Y=1.91 $X2=0 $Y2=0
cc_128 N_B1_c_135_n N_A4_c_171_n 2.2842e-19 $X=1.415 $Y=1.615 $X2=0 $Y2=0
cc_129 N_B1_c_134_n N_A4_c_174_n 0.0233642f $X=1.605 $Y=1.91 $X2=0 $Y2=0
cc_130 N_B1_M1004_g N_A4_c_172_n 0.00168307f $X=1.555 $Y=0.69 $X2=0 $Y2=0
cc_131 N_B1_c_134_n N_A4_c_172_n 0.00235529f $X=1.605 $Y=1.91 $X2=0 $Y2=0
cc_132 N_B1_c_135_n N_A4_c_172_n 0.0180089f $X=1.415 $Y=1.615 $X2=0 $Y2=0
cc_133 N_B1_c_134_n N_VPWR_c_335_n 0.0175164f $X=1.605 $Y=1.91 $X2=0 $Y2=0
cc_134 N_B1_c_134_n N_VPWR_c_339_n 0.00451101f $X=1.605 $Y=1.91 $X2=0 $Y2=0
cc_135 N_B1_c_134_n N_VPWR_c_334_n 0.00473652f $X=1.605 $Y=1.91 $X2=0 $Y2=0
cc_136 N_B1_M1004_g N_VGND_c_379_n 0.00391465f $X=1.555 $Y=0.69 $X2=0 $Y2=0
cc_137 N_B1_M1004_g N_VGND_c_382_n 0.00434272f $X=1.555 $Y=0.69 $X2=0 $Y2=0
cc_138 N_B1_M1004_g N_VGND_c_387_n 0.0082698f $X=1.555 $Y=0.69 $X2=0 $Y2=0
cc_139 N_B1_M1004_g N_A_326_74#_c_435_n 0.00266933f $X=1.555 $Y=0.69 $X2=0 $Y2=0
cc_140 N_B1_M1004_g N_A_326_74#_c_437_n 9.23518e-19 $X=1.555 $Y=0.69 $X2=0 $Y2=0
cc_141 N_A4_c_170_n N_A3_c_216_n 0.0271431f $X=2.14 $Y=1.52 $X2=-0.19 $Y2=-0.245
cc_142 N_A4_c_174_n N_A3_c_216_n 0.0592257f $X=2.14 $Y=1.765 $X2=-0.19
+ $Y2=-0.245
cc_143 N_A4_c_172_n N_A3_c_216_n 0.0033994f $X=2.035 $Y=1.355 $X2=-0.19
+ $Y2=-0.245
cc_144 N_A4_M1003_g N_A3_M1011_g 0.0230092f $X=2.055 $Y=0.69 $X2=0 $Y2=0
cc_145 N_A4_c_170_n N_A3_M1011_g 9.08436e-19 $X=2.14 $Y=1.52 $X2=0 $Y2=0
cc_146 N_A4_c_172_n N_A3_M1011_g 6.6431e-19 $X=2.035 $Y=1.355 $X2=0 $Y2=0
cc_147 N_A4_c_170_n N_A3_c_218_n 6.3137e-19 $X=2.14 $Y=1.52 $X2=0 $Y2=0
cc_148 N_A4_c_174_n N_A3_c_218_n 0.00418263f $X=2.14 $Y=1.765 $X2=0 $Y2=0
cc_149 N_A4_c_172_n N_A3_c_218_n 0.0407164f $X=2.035 $Y=1.355 $X2=0 $Y2=0
cc_150 N_A4_c_174_n N_VPWR_c_335_n 0.00439532f $X=2.14 $Y=1.765 $X2=0 $Y2=0
cc_151 N_A4_c_174_n N_VPWR_c_339_n 0.00447222f $X=2.14 $Y=1.765 $X2=0 $Y2=0
cc_152 N_A4_c_174_n N_VPWR_c_334_n 0.00864918f $X=2.14 $Y=1.765 $X2=0 $Y2=0
cc_153 N_A4_M1003_g N_VGND_c_380_n 0.00525427f $X=2.055 $Y=0.69 $X2=0 $Y2=0
cc_154 N_A4_M1003_g N_VGND_c_382_n 0.00434272f $X=2.055 $Y=0.69 $X2=0 $Y2=0
cc_155 N_A4_M1003_g N_VGND_c_387_n 0.00448875f $X=2.055 $Y=0.69 $X2=0 $Y2=0
cc_156 N_A4_M1003_g N_A_326_74#_c_435_n 0.00731128f $X=2.055 $Y=0.69 $X2=0 $Y2=0
cc_157 N_A4_M1003_g N_A_326_74#_c_436_n 0.00920125f $X=2.055 $Y=0.69 $X2=0 $Y2=0
cc_158 N_A4_c_170_n N_A_326_74#_c_436_n 6.23306e-19 $X=2.14 $Y=1.52 $X2=0 $Y2=0
cc_159 N_A4_c_172_n N_A_326_74#_c_436_n 0.0210835f $X=2.035 $Y=1.355 $X2=0 $Y2=0
cc_160 N_A4_M1003_g N_A_326_74#_c_437_n 8.39937e-19 $X=2.055 $Y=0.69 $X2=0 $Y2=0
cc_161 N_A4_c_170_n N_A_326_74#_c_437_n 8.57327e-19 $X=2.14 $Y=1.52 $X2=0 $Y2=0
cc_162 N_A4_c_172_n N_A_326_74#_c_437_n 0.0116993f $X=2.035 $Y=1.355 $X2=0 $Y2=0
cc_163 N_A4_M1003_g N_A_326_74#_c_438_n 5.97046e-19 $X=2.055 $Y=0.69 $X2=0 $Y2=0
cc_164 N_A3_c_216_n N_A2_M1007_g 0.0177025f $X=2.56 $Y=1.765 $X2=0 $Y2=0
cc_165 N_A3_M1011_g N_A2_M1007_g 0.0222036f $X=2.625 $Y=0.69 $X2=0 $Y2=0
cc_166 N_A3_c_218_n N_A2_M1007_g 5.15832e-19 $X=2.635 $Y=1.385 $X2=0 $Y2=0
cc_167 N_A3_c_216_n N_A2_c_256_n 0.0420633f $X=2.56 $Y=1.765 $X2=0 $Y2=0
cc_168 N_A3_c_218_n N_A2_c_256_n 0.00511818f $X=2.635 $Y=1.385 $X2=0 $Y2=0
cc_169 N_A3_c_216_n N_A2_c_257_n 0.00312103f $X=2.56 $Y=1.765 $X2=0 $Y2=0
cc_170 N_A3_c_218_n N_A2_c_257_n 0.0752933f $X=2.635 $Y=1.385 $X2=0 $Y2=0
cc_171 N_A3_c_216_n N_VPWR_c_339_n 0.00303293f $X=2.56 $Y=1.765 $X2=0 $Y2=0
cc_172 N_A3_c_218_n N_VPWR_c_339_n 0.00909385f $X=2.635 $Y=1.385 $X2=0 $Y2=0
cc_173 N_A3_c_216_n N_VPWR_c_334_n 0.00372936f $X=2.56 $Y=1.765 $X2=0 $Y2=0
cc_174 N_A3_c_218_n N_VPWR_c_334_n 0.0106888f $X=2.635 $Y=1.385 $X2=0 $Y2=0
cc_175 N_A3_c_218_n A_527_368# 0.0114459f $X=2.635 $Y=1.385 $X2=-0.19 $Y2=-0.245
cc_176 N_A3_M1011_g N_VGND_c_380_n 0.00387235f $X=2.625 $Y=0.69 $X2=0 $Y2=0
cc_177 N_A3_M1011_g N_VGND_c_381_n 4.25277e-19 $X=2.625 $Y=0.69 $X2=0 $Y2=0
cc_178 N_A3_M1011_g N_VGND_c_385_n 0.00434272f $X=2.625 $Y=0.69 $X2=0 $Y2=0
cc_179 N_A3_M1011_g N_VGND_c_387_n 0.00448792f $X=2.625 $Y=0.69 $X2=0 $Y2=0
cc_180 N_A3_M1011_g N_A_326_74#_c_435_n 5.97046e-19 $X=2.625 $Y=0.69 $X2=0 $Y2=0
cc_181 N_A3_c_216_n N_A_326_74#_c_436_n 5.31519e-19 $X=2.56 $Y=1.765 $X2=0 $Y2=0
cc_182 N_A3_M1011_g N_A_326_74#_c_436_n 0.00935164f $X=2.625 $Y=0.69 $X2=0 $Y2=0
cc_183 N_A3_c_218_n N_A_326_74#_c_436_n 0.0139058f $X=2.635 $Y=1.385 $X2=0 $Y2=0
cc_184 N_A3_M1011_g N_A_326_74#_c_438_n 0.00730737f $X=2.625 $Y=0.69 $X2=0 $Y2=0
cc_185 N_A3_c_216_n N_A_326_74#_c_441_n 7.62276e-19 $X=2.56 $Y=1.765 $X2=0 $Y2=0
cc_186 N_A3_M1011_g N_A_326_74#_c_441_n 8.85434e-19 $X=2.625 $Y=0.69 $X2=0 $Y2=0
cc_187 N_A3_c_218_n N_A_326_74#_c_441_n 0.00964811f $X=2.635 $Y=1.385 $X2=0
+ $Y2=0
cc_188 N_A2_c_256_n N_A1_c_289_n 0.0511977f $X=3.13 $Y=1.765 $X2=-0.19
+ $Y2=-0.245
cc_189 N_A2_c_257_n N_A1_c_289_n 0.012467f $X=3.205 $Y=1.465 $X2=-0.19
+ $Y2=-0.245
cc_190 N_A2_M1007_g N_A1_M1009_g 0.0200135f $X=3.115 $Y=0.69 $X2=0 $Y2=0
cc_191 N_A2_c_256_n N_A1_M1009_g 0.00172681f $X=3.13 $Y=1.765 $X2=0 $Y2=0
cc_192 N_A2_c_257_n N_A1_M1009_g 2.87867e-19 $X=3.205 $Y=1.465 $X2=0 $Y2=0
cc_193 N_A2_c_256_n N_A1_c_291_n 0.00160884f $X=3.13 $Y=1.765 $X2=0 $Y2=0
cc_194 N_A2_c_257_n N_A1_c_291_n 0.0404044f $X=3.205 $Y=1.465 $X2=0 $Y2=0
cc_195 N_A2_c_256_n N_VPWR_c_337_n 0.0013972f $X=3.13 $Y=1.765 $X2=0 $Y2=0
cc_196 N_A2_c_257_n N_VPWR_c_337_n 0.0240637f $X=3.205 $Y=1.465 $X2=0 $Y2=0
cc_197 N_A2_c_256_n N_VPWR_c_339_n 0.00303293f $X=3.13 $Y=1.765 $X2=0 $Y2=0
cc_198 N_A2_c_257_n N_VPWR_c_339_n 0.00968684f $X=3.205 $Y=1.465 $X2=0 $Y2=0
cc_199 N_A2_c_256_n N_VPWR_c_334_n 0.00374185f $X=3.13 $Y=1.765 $X2=0 $Y2=0
cc_200 N_A2_c_257_n N_VPWR_c_334_n 0.0119091f $X=3.205 $Y=1.465 $X2=0 $Y2=0
cc_201 N_A2_c_257_n A_641_368# 0.0140938f $X=3.205 $Y=1.465 $X2=-0.19 $Y2=-0.245
cc_202 N_A2_M1007_g N_VGND_c_381_n 0.0136443f $X=3.115 $Y=0.69 $X2=0 $Y2=0
cc_203 N_A2_M1007_g N_VGND_c_385_n 0.00413917f $X=3.115 $Y=0.69 $X2=0 $Y2=0
cc_204 N_A2_M1007_g N_VGND_c_387_n 0.00417193f $X=3.115 $Y=0.69 $X2=0 $Y2=0
cc_205 N_A2_M1007_g N_A_326_74#_c_438_n 0.00265992f $X=3.115 $Y=0.69 $X2=0 $Y2=0
cc_206 N_A2_M1007_g N_A_326_74#_c_439_n 0.0138853f $X=3.115 $Y=0.69 $X2=0 $Y2=0
cc_207 N_A2_c_256_n N_A_326_74#_c_439_n 0.00113455f $X=3.13 $Y=1.765 $X2=0 $Y2=0
cc_208 N_A2_c_257_n N_A_326_74#_c_439_n 0.0195066f $X=3.205 $Y=1.465 $X2=0 $Y2=0
cc_209 N_A2_M1007_g N_A_326_74#_c_440_n 9.0724e-19 $X=3.115 $Y=0.69 $X2=0 $Y2=0
cc_210 N_A1_c_291_n N_VPWR_M1001_d 0.00759963f $X=3.775 $Y=1.515 $X2=0 $Y2=0
cc_211 N_A1_c_289_n N_VPWR_c_337_n 0.0165781f $X=3.7 $Y=1.765 $X2=0 $Y2=0
cc_212 N_A1_c_291_n N_VPWR_c_337_n 0.0338132f $X=3.775 $Y=1.515 $X2=0 $Y2=0
cc_213 N_A1_c_289_n N_VPWR_c_339_n 0.00413917f $X=3.7 $Y=1.765 $X2=0 $Y2=0
cc_214 N_A1_c_289_n N_VPWR_c_334_n 0.00818781f $X=3.7 $Y=1.765 $X2=0 $Y2=0
cc_215 N_A1_M1009_g N_VGND_c_381_n 0.00623438f $X=3.825 $Y=0.69 $X2=0 $Y2=0
cc_216 N_A1_M1009_g N_VGND_c_386_n 0.00434272f $X=3.825 $Y=0.69 $X2=0 $Y2=0
cc_217 N_A1_M1009_g N_VGND_c_387_n 0.00452716f $X=3.825 $Y=0.69 $X2=0 $Y2=0
cc_218 N_A1_c_289_n N_A_326_74#_c_439_n 0.00113297f $X=3.7 $Y=1.765 $X2=0 $Y2=0
cc_219 N_A1_M1009_g N_A_326_74#_c_439_n 0.0119089f $X=3.825 $Y=0.69 $X2=0 $Y2=0
cc_220 N_A1_c_291_n N_A_326_74#_c_439_n 0.0310954f $X=3.775 $Y=1.515 $X2=0 $Y2=0
cc_221 N_A1_M1009_g N_A_326_74#_c_440_n 0.00786806f $X=3.825 $Y=0.69 $X2=0 $Y2=0
cc_222 X N_VPWR_c_335_n 0.026735f $X=0.155 $Y=2.32 $X2=0 $Y2=0
cc_223 X N_VPWR_c_338_n 0.0146013f $X=0.155 $Y=2.69 $X2=0 $Y2=0
cc_224 X N_VPWR_c_334_n 0.0120495f $X=0.155 $Y=2.69 $X2=0 $Y2=0
cc_225 N_X_c_313_n N_VGND_c_379_n 0.023562f $X=0.28 $Y=0.515 $X2=0 $Y2=0
cc_226 N_X_c_313_n N_VGND_c_384_n 0.0115122f $X=0.28 $Y=0.515 $X2=0 $Y2=0
cc_227 N_X_c_313_n N_VGND_c_387_n 0.0095288f $X=0.28 $Y=0.515 $X2=0 $Y2=0
cc_228 N_VGND_c_380_n N_A_326_74#_c_435_n 0.0131729f $X=2.34 $Y=0.515 $X2=0
+ $Y2=0
cc_229 N_VGND_c_382_n N_A_326_74#_c_435_n 0.0145482f $X=2.175 $Y=0 $X2=0 $Y2=0
cc_230 N_VGND_c_387_n N_A_326_74#_c_435_n 0.0119922f $X=4.08 $Y=0 $X2=0 $Y2=0
cc_231 N_VGND_M1003_d N_A_326_74#_c_436_n 0.00373913f $X=2.13 $Y=0.37 $X2=0
+ $Y2=0
cc_232 N_VGND_c_380_n N_A_326_74#_c_436_n 0.0243707f $X=2.34 $Y=0.515 $X2=0
+ $Y2=0
cc_233 N_VGND_c_387_n N_A_326_74#_c_436_n 0.0109408f $X=4.08 $Y=0 $X2=0 $Y2=0
cc_234 N_VGND_c_380_n N_A_326_74#_c_438_n 0.0131729f $X=2.34 $Y=0.515 $X2=0
+ $Y2=0
cc_235 N_VGND_c_381_n N_A_326_74#_c_438_n 0.0141032f $X=3.44 $Y=0.515 $X2=0
+ $Y2=0
cc_236 N_VGND_c_385_n N_A_326_74#_c_438_n 0.0145482f $X=3.175 $Y=0 $X2=0 $Y2=0
cc_237 N_VGND_c_387_n N_A_326_74#_c_438_n 0.0119922f $X=4.08 $Y=0 $X2=0 $Y2=0
cc_238 N_VGND_M1007_d N_A_326_74#_c_439_n 0.00644036f $X=3.19 $Y=0.37 $X2=0
+ $Y2=0
cc_239 N_VGND_c_381_n N_A_326_74#_c_439_n 0.0365648f $X=3.44 $Y=0.515 $X2=0
+ $Y2=0
cc_240 N_VGND_c_387_n N_A_326_74#_c_439_n 0.0114864f $X=4.08 $Y=0 $X2=0 $Y2=0
cc_241 N_VGND_c_381_n N_A_326_74#_c_440_n 0.0132315f $X=3.44 $Y=0.515 $X2=0
+ $Y2=0
cc_242 N_VGND_c_386_n N_A_326_74#_c_440_n 0.0145639f $X=4.08 $Y=0 $X2=0 $Y2=0
cc_243 N_VGND_c_387_n N_A_326_74#_c_440_n 0.0119984f $X=4.08 $Y=0 $X2=0 $Y2=0
