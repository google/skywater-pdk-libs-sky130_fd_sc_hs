* NGSPICE file created from sky130_fd_sc_hs__or2_4.ext - technology: sky130A

.subckt sky130_fd_sc_hs__or2_4 A B VGND VNB VPB VPWR X
M1000 VGND B a_83_260# VNB nlowvt w=740000u l=150000u
+  ad=1.6058e+12p pd=1.026e+07u as=2.479e+11p ps=2.15e+06u
M1001 a_83_260# A VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1002 X a_83_260# VGND VNB nlowvt w=740000u l=150000u
+  ad=4.773e+11p pd=4.25e+06u as=0p ps=0u
M1003 VGND a_83_260# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 VPWR a_83_260# X VPB pshort w=1.12e+06u l=150000u
+  ad=1.4068e+12p pd=1.132e+07u as=6.72e+11p ps=5.68e+06u
M1005 X a_83_260# VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 X a_83_260# VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_493_388# A VPWR VPB pshort w=1e+06u l=150000u
+  ad=6.5e+11p pd=5.3e+06u as=0p ps=0u
M1008 VPWR a_83_260# X VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_83_260# B a_493_388# VPB pshort w=1e+06u l=150000u
+  ad=3e+11p pd=2.6e+06u as=0p ps=0u
M1010 VPWR A a_493_388# VPB pshort w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_493_388# B a_83_260# VPB pshort w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 X a_83_260# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VGND a_83_260# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

