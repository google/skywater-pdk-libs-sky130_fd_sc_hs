* File: sky130_fd_sc_hs__or3b_4.spice
* Created: Tue Sep  1 20:20:57 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hs__or3b_4.pex.spice"
.subckt sky130_fd_sc_hs__or3b_4  VNB VPB C_N A B VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* B	B
* A	A
* C_N	C_N
* VPB	VPB
* VNB	VNB
MM1017 N_VGND_M1017_d N_C_N_M1017_g N_A_27_392#_M1017_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.66075 AS=0.1824 PD=3.58 PS=1.85 NRD=183.264 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75000.7 A=0.096 P=1.58 MULT=1
MM1011 N_VGND_M1011_d N_A_27_392#_M1011_g N_A_409_392#_M1011_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1295 AS=0.2072 PD=1.09 PS=2.04 NRD=11.34 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75003 A=0.111 P=1.78 MULT=1
MM1008 N_A_409_392#_M1008_d N_B_M1008_g N_VGND_M1011_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1295 PD=1.02 PS=1.09 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.7
+ SB=75002.5 A=0.111 P=1.78 MULT=1
MM1015 N_VGND_M1015_d N_A_M1015_g N_A_409_392#_M1008_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.1332 AS=0.1036 PD=1.1 PS=1.02 NRD=12.156 NRS=0 M=1 R=4.93333 SA=75001.1
+ SB=75002.1 A=0.111 P=1.78 MULT=1
MM1002 N_X_M1002_d N_A_409_392#_M1002_g N_VGND_M1015_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.11285 AS=0.1332 PD=1.045 PS=1.1 NRD=4.044 NRS=0.804 M=1 R=4.93333
+ SA=75001.6 SB=75001.6 A=0.111 P=1.78 MULT=1
MM1004 N_X_M1002_d N_A_409_392#_M1004_g N_VGND_M1004_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.11285 AS=0.1221 PD=1.045 PS=1.07 NRD=0 NRS=0 M=1 R=4.93333 SA=75002.1
+ SB=75001.1 A=0.111 P=1.78 MULT=1
MM1010 N_X_M1010_d N_A_409_392#_M1010_g N_VGND_M1004_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1221 PD=1.02 PS=1.07 NRD=0 NRS=8.1 M=1 R=4.93333 SA=75002.6
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1018 N_X_M1010_d N_A_409_392#_M1018_g N_VGND_M1018_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.2109 PD=1.02 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333 SA=75003
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1013 N_VPWR_M1013_d N_C_N_M1013_g N_A_27_392#_M1013_s VPB PSHORT L=0.15 W=1
+ AD=0.18 AS=0.29 PD=1.36 PS=2.58 NRD=1.9503 NRS=1.9503 M=1 R=6.66667 SA=75000.2
+ SB=75005 A=0.15 P=2.3 MULT=1
MM1000 N_A_217_392#_M1000_d N_A_M1000_g N_VPWR_M1013_d VPB PSHORT L=0.15 W=1
+ AD=0.15 AS=0.18 PD=1.3 PS=1.36 NRD=1.9503 NRS=13.7703 M=1 R=6.66667 SA=75000.7
+ SB=75004.5 A=0.15 P=2.3 MULT=1
MM1003 N_A_307_392#_M1003_d N_B_M1003_g N_A_217_392#_M1000_d VPB PSHORT L=0.15
+ W=1 AD=0.18 AS=0.15 PD=1.36 PS=1.3 NRD=13.7703 NRS=1.9503 M=1 R=6.66667
+ SA=75001.2 SB=75004 A=0.15 P=2.3 MULT=1
MM1012 N_A_409_392#_M1012_d N_A_27_392#_M1012_g N_A_307_392#_M1003_d VPB PSHORT
+ L=0.15 W=1 AD=0.1625 AS=0.18 PD=1.325 PS=1.36 NRD=3.9203 NRS=1.9503 M=1
+ R=6.66667 SA=75001.7 SB=75003.5 A=0.15 P=2.3 MULT=1
MM1014 N_A_409_392#_M1012_d N_A_27_392#_M1014_g N_A_307_392#_M1014_s VPB PSHORT
+ L=0.15 W=1 AD=0.1625 AS=0.15 PD=1.325 PS=1.3 NRD=4.9053 NRS=1.9503 M=1
+ R=6.66667 SA=75002.2 SB=75003 A=0.15 P=2.3 MULT=1
MM1016 N_A_307_392#_M1014_s N_B_M1016_g N_A_217_392#_M1016_s VPB PSHORT L=0.15
+ W=1 AD=0.15 AS=0.18 PD=1.3 PS=1.36 NRD=1.9503 NRS=11.8003 M=1 R=6.66667
+ SA=75002.6 SB=75002.6 A=0.15 P=2.3 MULT=1
MM1007 N_A_217_392#_M1016_s N_A_M1007_g N_VPWR_M1007_s VPB PSHORT L=0.15 W=1
+ AD=0.18 AS=0.184811 PD=1.36 PS=1.39623 NRD=3.9203 NRS=9.8303 M=1 R=6.66667
+ SA=75003.1 SB=75002.1 A=0.15 P=2.3 MULT=1
MM1001 N_X_M1001_d N_A_409_392#_M1001_g N_VPWR_M1007_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.206989 PD=1.42 PS=1.56377 NRD=1.7533 NRS=5.2599 M=1 R=7.46667
+ SA=75003.3 SB=75001.6 A=0.168 P=2.54 MULT=1
MM1005 N_X_M1001_d N_A_409_392#_M1005_g N_VPWR_M1005_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75003.7 SB=75001.1 A=0.168 P=2.54 MULT=1
MM1006 N_X_M1006_d N_A_409_392#_M1006_g N_VPWR_M1005_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75004.2 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1009 N_X_M1006_d N_A_409_392#_M1009_g N_VPWR_M1009_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.3192 PD=1.42 PS=2.81 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75004.6 SB=75000.2 A=0.168 P=2.54 MULT=1
DX19_noxref VNB VPB NWDIODE A=11.4204 P=16
*
.include "sky130_fd_sc_hs__or3b_4.pxi.spice"
*
.ends
*
*
