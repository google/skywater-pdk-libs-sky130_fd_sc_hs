* File: sky130_fd_sc_hs__a22oi_1.pex.spice
* Created: Tue Sep  1 19:51:23 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HS__A22OI_1%B2 1 3 6 8 9 10 11
c29 1 0 4.6169e-20 $X=0.705 $Y=1.765
r30 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.27
+ $Y=1.385 $X2=0.27 $Y2=1.385
r31 11 16 9.7783 $w=3.28e-07 $l=2.8e-07 $layer=LI1_cond $X=0.27 $Y=1.665
+ $X2=0.27 $Y2=1.385
r32 10 16 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=0.27 $Y=1.295 $X2=0.27
+ $Y2=1.385
r33 8 15 60.3271 $w=3.3e-07 $l=3.45e-07 $layer=POLY_cond $X=0.615 $Y=1.385
+ $X2=0.27 $Y2=1.385
r34 8 9 66.2869 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=0.705 $Y=1.385
+ $X2=0.705 $Y2=1.22
r35 6 9 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=0.72 $Y=0.74 $X2=0.72
+ $Y2=1.22
r36 1 8 149.859 $w=1.8e-07 $l=3.8e-07 $layer=POLY_cond $X=0.705 $Y=1.765
+ $X2=0.705 $Y2=1.385
r37 1 3 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.705 $Y=1.765
+ $X2=0.705 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_HS__A22OI_1%B1 3 5 7 8 12
c33 12 0 4.6169e-20 $X=1.17 $Y=1.515
c34 5 0 4.8353e-20 $X=1.155 $Y=1.765
r35 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.17
+ $Y=1.515 $X2=1.17 $Y2=1.515
r36 8 12 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=1.17 $Y=1.665
+ $X2=1.17 $Y2=1.515
r37 5 11 52.2586 $w=2.99e-07 $l=2.57391e-07 $layer=POLY_cond $X=1.155 $Y=1.765
+ $X2=1.17 $Y2=1.515
r38 5 7 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.155 $Y=1.765
+ $X2=1.155 $Y2=2.4
r39 1 11 38.5562 $w=2.99e-07 $l=2.05122e-07 $layer=POLY_cond $X=1.08 $Y=1.35
+ $X2=1.17 $Y2=1.515
r40 1 3 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.08 $Y=1.35 $X2=1.08
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HS__A22OI_1%A1 3 5 7 8 12
r28 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.71
+ $Y=1.515 $X2=1.71 $Y2=1.515
r29 8 12 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=1.71 $Y=1.665
+ $X2=1.71 $Y2=1.515
r30 5 11 52.2586 $w=2.99e-07 $l=2.85044e-07 $layer=POLY_cond $X=1.635 $Y=1.765
+ $X2=1.71 $Y2=1.515
r31 5 7 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.635 $Y=1.765
+ $X2=1.635 $Y2=2.4
r32 1 11 38.5562 $w=2.99e-07 $l=2.05122e-07 $layer=POLY_cond $X=1.62 $Y=1.35
+ $X2=1.71 $Y2=1.515
r33 1 3 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.62 $Y=1.35 $X2=1.62
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HS__A22OI_1%A2 3 5 7 8 9
r25 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.25
+ $Y=1.515 $X2=2.25 $Y2=1.515
r26 9 14 10.4524 $w=4.28e-07 $l=3.9e-07 $layer=LI1_cond $X=2.64 $Y=1.565
+ $X2=2.25 $Y2=1.565
r27 8 14 2.41209 $w=4.28e-07 $l=9e-08 $layer=LI1_cond $X=2.16 $Y=1.565 $X2=2.25
+ $Y2=1.565
r28 5 13 52.2586 $w=2.99e-07 $l=2.85044e-07 $layer=POLY_cond $X=2.175 $Y=1.765
+ $X2=2.25 $Y2=1.515
r29 5 7 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.175 $Y=1.765
+ $X2=2.175 $Y2=2.4
r30 1 13 38.5562 $w=2.99e-07 $l=2.05122e-07 $layer=POLY_cond $X=2.16 $Y=1.35
+ $X2=2.25 $Y2=1.515
r31 1 3 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.16 $Y=1.35 $X2=2.16
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HS__A22OI_1%A_71_368# 1 2 3 12 14 15 16 19 20 22 24
r39 22 29 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.4 $Y=2.12 $X2=2.4
+ $Y2=2.035
r40 22 24 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=2.4 $Y=2.12 $X2=2.4
+ $Y2=2.815
r41 21 27 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.545 $Y=2.035
+ $X2=1.38 $Y2=2.035
r42 20 29 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.235 $Y=2.035
+ $X2=2.4 $Y2=2.035
r43 20 21 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=2.235 $Y=2.035
+ $X2=1.545 $Y2=2.035
r44 17 19 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=1.38 $Y=2.905 $X2=1.38
+ $Y2=2.815
r45 16 27 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.38 $Y=2.12 $X2=1.38
+ $Y2=2.035
r46 16 19 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=1.38 $Y=2.12
+ $X2=1.38 $Y2=2.815
r47 14 17 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.215 $Y=2.99
+ $X2=1.38 $Y2=2.905
r48 14 15 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=1.215 $Y=2.99
+ $X2=0.645 $Y2=2.99
r49 10 15 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.48 $Y=2.905
+ $X2=0.645 $Y2=2.99
r50 10 12 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=0.48 $Y=2.905
+ $X2=0.48 $Y2=2.455
r51 3 29 400 $w=1.7e-07 $l=3.4187e-07 $layer=licon1_PDIFF $count=1 $X=2.25
+ $Y=1.84 $X2=2.4 $Y2=2.115
r52 3 24 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=2.25
+ $Y=1.84 $X2=2.4 $Y2=2.815
r53 2 27 400 $w=1.7e-07 $l=3.4187e-07 $layer=licon1_PDIFF $count=1 $X=1.23
+ $Y=1.84 $X2=1.38 $Y2=2.115
r54 2 19 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=1.23
+ $Y=1.84 $X2=1.38 $Y2=2.815
r55 1 12 300 $w=1.7e-07 $l=6.74611e-07 $layer=licon1_PDIFF $count=2 $X=0.355
+ $Y=1.84 $X2=0.48 $Y2=2.455
.ends

.subckt PM_SKY130_FD_SC_HS__A22OI_1%Y 1 2 7 8 13 20 22 23
c38 20 0 4.8353e-20 $X=0.93 $Y=2.115
r39 22 23 18.5393 $w=2.28e-07 $l=3.7e-07 $layer=LI1_cond $X=0.72 $Y=1.295
+ $X2=0.72 $Y2=1.665
r40 17 23 14.2803 $w=2.28e-07 $l=2.85e-07 $layer=LI1_cond $X=0.72 $Y=1.95
+ $X2=0.72 $Y2=1.665
r41 17 20 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=0.72 $Y=2.035
+ $X2=0.93 $Y2=2.035
r42 15 22 5.76222 $w=2.28e-07 $l=1.15e-07 $layer=LI1_cond $X=0.72 $Y=1.18
+ $X2=0.72 $Y2=1.295
r43 11 13 12.965 $w=4.38e-07 $l=4.95e-07 $layer=LI1_cond $X=1.35 $Y=1.01
+ $X2=1.35 $Y2=0.515
r44 8 15 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=0.835 $Y=1.095
+ $X2=0.72 $Y2=1.18
r45 7 11 8.71846 $w=1.7e-07 $l=2.59037e-07 $layer=LI1_cond $X=1.13 $Y=1.095
+ $X2=1.35 $Y2=1.01
r46 7 8 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=1.13 $Y=1.095
+ $X2=0.835 $Y2=1.095
r47 2 20 300 $w=1.7e-07 $l=3.4187e-07 $layer=licon1_PDIFF $count=2 $X=0.78
+ $Y=1.84 $X2=0.93 $Y2=2.115
r48 1 13 91 $w=1.7e-07 $l=2.57488e-07 $layer=licon1_NDIFF $count=2 $X=1.155
+ $Y=0.37 $X2=1.35 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__A22OI_1%VPWR 1 6 9 10 11 21 22
r26 21 22 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r27 19 22 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.64 $Y2=3.33
r28 18 19 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r29 14 18 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=0.24 $Y=3.33
+ $X2=1.68 $Y2=3.33
r30 14 15 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r31 11 19 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.44 $Y=3.33
+ $X2=1.68 $Y2=3.33
r32 11 15 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=1.44 $Y=3.33
+ $X2=0.24 $Y2=3.33
r33 9 18 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=1.715 $Y=3.33
+ $X2=1.68 $Y2=3.33
r34 9 10 8.9695 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=1.715 $Y=3.33 $X2=1.89
+ $Y2=3.33
r35 8 21 37.5134 $w=1.68e-07 $l=5.75e-07 $layer=LI1_cond $X=2.065 $Y=3.33
+ $X2=2.64 $Y2=3.33
r36 8 10 8.9695 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=2.065 $Y=3.33 $X2=1.89
+ $Y2=3.33
r37 4 10 1.07557 $w=3.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.89 $Y=3.245 $X2=1.89
+ $Y2=3.33
r38 4 6 26.0123 $w=3.48e-07 $l=7.9e-07 $layer=LI1_cond $X=1.89 $Y=3.245 $X2=1.89
+ $Y2=2.455
r39 1 6 300 $w=1.7e-07 $l=6.99232e-07 $layer=licon1_PDIFF $count=2 $X=1.71
+ $Y=1.84 $X2=1.89 $Y2=2.455
.ends

.subckt PM_SKY130_FD_SC_HS__A22OI_1%VGND 1 2 9 13 16 17 19 20 21 34 35
r30 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r31 32 35 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r32 31 32 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r33 28 31 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=0.72 $Y=0 $X2=2.16
+ $Y2=0
r34 28 29 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r35 25 29 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r36 24 25 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r37 21 32 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.44 $Y=0 $X2=2.16
+ $Y2=0
r38 21 29 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.44 $Y=0 $X2=0.72
+ $Y2=0
r39 19 31 3.26203 $w=1.68e-07 $l=5e-08 $layer=LI1_cond $X=2.21 $Y=0 $X2=2.16
+ $Y2=0
r40 19 20 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.21 $Y=0 $X2=2.375
+ $Y2=0
r41 18 34 6.52406 $w=1.68e-07 $l=1e-07 $layer=LI1_cond $X=2.54 $Y=0 $X2=2.64
+ $Y2=0
r42 18 20 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.54 $Y=0 $X2=2.375
+ $Y2=0
r43 16 24 6.52406 $w=1.68e-07 $l=1e-07 $layer=LI1_cond $X=0.34 $Y=0 $X2=0.24
+ $Y2=0
r44 16 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.34 $Y=0 $X2=0.505
+ $Y2=0
r45 15 28 3.26203 $w=1.68e-07 $l=5e-08 $layer=LI1_cond $X=0.67 $Y=0 $X2=0.72
+ $Y2=0
r46 15 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.67 $Y=0 $X2=0.505
+ $Y2=0
r47 11 20 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.375 $Y=0.085
+ $X2=2.375 $Y2=0
r48 11 13 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=2.375 $Y=0.085
+ $X2=2.375 $Y2=0.515
r49 7 17 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.505 $Y=0.085
+ $X2=0.505 $Y2=0
r50 7 9 20.6043 $w=3.28e-07 $l=5.9e-07 $layer=LI1_cond $X=0.505 $Y=0.085
+ $X2=0.505 $Y2=0.675
r51 2 13 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.235
+ $Y=0.37 $X2=2.375 $Y2=0.515
r52 1 9 182 $w=1.7e-07 $l=3.62146e-07 $layer=licon1_NDIFF $count=1 $X=0.38
+ $Y=0.37 $X2=0.505 $Y2=0.675
.ends

