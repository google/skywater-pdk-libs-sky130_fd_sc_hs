* File: sky130_fd_sc_hs__nor3_4.pex.spice
* Created: Tue Sep  1 20:11:38 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HS__NOR3_4%A 3 5 7 10 12 14 15 17 18 20 21 23 26 28 32
+ 33 37 38 42 43 44 55 58
c138 28 0 1.39786e-19 $X=5.805 $Y=2.105
c139 23 0 1.56752e-19 $X=0.77 $Y=1.515
c140 10 0 7.79871e-20 $X=0.935 $Y=0.74
r141 58 69 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=1.71 $Y=2.045
+ $X2=1.71 $Y2=2.255
r142 55 56 1.92287 $w=3.76e-07 $l=1.5e-08 $layer=POLY_cond $X=0.935 $Y=1.557
+ $X2=0.95 $Y2=1.557
r143 52 53 0.640957 $w=3.76e-07 $l=5e-09 $layer=POLY_cond $X=0.495 $Y=1.557
+ $X2=0.5 $Y2=1.557
r144 44 58 0.652406 $w=1.68e-07 $l=1e-08 $layer=LI1_cond $X=1.71 $Y=2.035
+ $X2=1.71 $Y2=2.045
r145 44 58 0.691466 $w=2.48e-07 $l=1.5e-08 $layer=LI1_cond $X=1.61 $Y=2.045
+ $X2=1.625 $Y2=2.045
r146 43 44 18.9001 $w=2.48e-07 $l=4.1e-07 $layer=LI1_cond $X=1.2 $Y=2.045
+ $X2=1.61 $Y2=2.045
r147 43 59 12.2159 $w=2.48e-07 $l=2.65e-07 $layer=LI1_cond $X=1.2 $Y=2.045
+ $X2=0.935 $Y2=2.045
r148 42 59 3.97509 $w=2.5e-07 $l=1.65e-07 $layer=LI1_cond $X=0.77 $Y=2.045
+ $X2=0.935 $Y2=2.045
r149 38 40 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=3.935 $Y=2.105
+ $X2=3.935 $Y2=2.255
r150 37 49 10.716 $w=5.7e-07 $l=1.2e-07 $layer=POLY_cond $X=6 $Y=1.515 $X2=6
+ $Y2=1.395
r151 36 37 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.97
+ $Y=1.515 $X2=5.97 $Y2=1.515
r152 33 49 84.4783 $w=5.7e-07 $l=9e-07 $layer=POLY_cond $X=6 $Y=0.495 $X2=6
+ $Y2=1.395
r153 32 36 35.621 $w=3.28e-07 $l=1.02e-06 $layer=LI1_cond $X=5.97 $Y=0.495
+ $X2=5.97 $Y2=1.515
r154 32 33 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.97
+ $Y=0.495 $X2=5.97 $Y2=0.495
r155 30 36 17.6359 $w=3.28e-07 $l=5.05e-07 $layer=LI1_cond $X=5.97 $Y=2.02
+ $X2=5.97 $Y2=1.515
r156 29 38 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.02 $Y=2.105
+ $X2=3.935 $Y2=2.105
r157 28 30 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=5.805 $Y=2.105
+ $X2=5.97 $Y2=2.02
r158 28 29 116.455 $w=1.68e-07 $l=1.785e-06 $layer=LI1_cond $X=5.805 $Y=2.105
+ $X2=4.02 $Y2=2.105
r159 27 69 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.795 $Y=2.255
+ $X2=1.71 $Y2=2.255
r160 26 40 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.85 $Y=2.255
+ $X2=3.935 $Y2=2.255
r161 26 27 134.07 $w=1.68e-07 $l=2.055e-06 $layer=LI1_cond $X=3.85 $Y=2.255
+ $X2=1.795 $Y2=2.255
r162 24 55 21.1516 $w=3.76e-07 $l=1.65e-07 $layer=POLY_cond $X=0.77 $Y=1.557
+ $X2=0.935 $Y2=1.557
r163 24 53 34.6117 $w=3.76e-07 $l=2.7e-07 $layer=POLY_cond $X=0.77 $Y=1.557
+ $X2=0.5 $Y2=1.557
r164 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.77
+ $Y=1.515 $X2=0.77 $Y2=1.515
r165 21 42 3.01144 $w=3.3e-07 $l=1.25e-07 $layer=LI1_cond $X=0.77 $Y=1.92
+ $X2=0.77 $Y2=2.045
r166 21 23 14.1436 $w=3.28e-07 $l=4.05e-07 $layer=LI1_cond $X=0.77 $Y=1.92
+ $X2=0.77 $Y2=1.515
r167 18 37 48.6761 $w=2.57e-07 $l=3.44601e-07 $layer=POLY_cond $X=6.225 $Y=1.765
+ $X2=6 $Y2=1.515
r168 18 20 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=6.225 $Y=1.765
+ $X2=6.225 $Y2=2.4
r169 15 37 48.6761 $w=2.57e-07 $l=3.44601e-07 $layer=POLY_cond $X=5.775 $Y=1.765
+ $X2=6 $Y2=1.515
r170 15 17 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=5.775 $Y=1.765
+ $X2=5.775 $Y2=2.4
r171 12 56 24.356 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=0.95 $Y=1.765
+ $X2=0.95 $Y2=1.557
r172 12 14 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.95 $Y=1.765
+ $X2=0.95 $Y2=2.4
r173 8 55 24.356 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.935 $Y=1.35
+ $X2=0.935 $Y2=1.557
r174 8 10 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=0.935 $Y=1.35
+ $X2=0.935 $Y2=0.74
r175 5 53 24.356 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=0.5 $Y=1.765 $X2=0.5
+ $Y2=1.557
r176 5 7 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.5 $Y=1.765 $X2=0.5
+ $Y2=2.4
r177 1 52 24.356 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.495 $Y=1.35
+ $X2=0.495 $Y2=1.557
r178 1 3 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=0.495 $Y=1.35
+ $X2=0.495 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HS__NOR3_4%B 2 3 5 6 8 9 11 13 15 16 18 20 21 23 25 26
+ 28 29 34 37 43 44 54 56 57 61 63 65 67
c126 54 0 1.39786e-19 $X=5.325 $Y=1.345
c127 34 0 1.16344e-19 $X=4.8 $Y=1.345
c128 26 0 9.77441e-20 $X=5.325 $Y=1.765
c129 11 0 4.22428e-20 $X=1.925 $Y=1.185
r130 57 63 1.86425 $w=3.38e-07 $l=5.5e-08 $layer=LI1_cond $X=2.215 $Y=1.35
+ $X2=2.16 $Y2=1.35
r131 56 65 1.86425 $w=3.38e-07 $l=5.5e-08 $layer=LI1_cond $X=2.585 $Y=1.35
+ $X2=2.64 $Y2=1.35
r132 53 54 78.6876 $w=3.3e-07 $l=4.5e-07 $layer=POLY_cond $X=4.875 $Y=1.345
+ $X2=5.325 $Y2=1.345
r133 44 67 3.38954 $w=3.38e-07 $l=1e-07 $layer=LI1_cond $X=2.655 $Y=1.35
+ $X2=2.755 $Y2=1.35
r134 44 65 0.508431 $w=3.38e-07 $l=1.5e-08 $layer=LI1_cond $X=2.655 $Y=1.35
+ $X2=2.64 $Y2=1.35
r135 44 56 0.508431 $w=3.38e-07 $l=1.5e-08 $layer=LI1_cond $X=2.57 $Y=1.35
+ $X2=2.585 $Y2=1.35
r136 43 63 0.508431 $w=3.38e-07 $l=1.5e-08 $layer=LI1_cond $X=2.145 $Y=1.35
+ $X2=2.16 $Y2=1.35
r137 43 61 6.26872 $w=3.38e-07 $l=1e-07 $layer=LI1_cond $X=2.145 $Y=1.35
+ $X2=2.045 $Y2=1.35
r138 43 44 11.5244 $w=3.38e-07 $l=3.4e-07 $layer=LI1_cond $X=2.23 $Y=1.35
+ $X2=2.57 $Y2=1.35
r139 43 57 0.508431 $w=3.38e-07 $l=1.5e-08 $layer=LI1_cond $X=2.23 $Y=1.35
+ $X2=2.215 $Y2=1.35
r140 40 41 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.475
+ $Y=1.515 $X2=1.475 $Y2=1.515
r141 37 40 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=1.475 $Y=1.435
+ $X2=1.475 $Y2=1.515
r142 35 53 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=4.8 $Y=1.345
+ $X2=4.875 $Y2=1.345
r143 35 50 65.573 $w=3.3e-07 $l=3.75e-07 $layer=POLY_cond $X=4.8 $Y=1.345
+ $X2=4.425 $Y2=1.345
r144 34 67 71.4165 $w=3.28e-07 $l=2.045e-06 $layer=LI1_cond $X=4.8 $Y=1.345
+ $X2=2.755 $Y2=1.345
r145 34 35 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.8
+ $Y=1.345 $X2=4.8 $Y2=1.345
r146 31 37 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.64 $Y=1.435
+ $X2=1.475 $Y2=1.435
r147 31 61 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=1.64 $Y=1.435
+ $X2=2.045 $Y2=1.435
r148 26 28 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=5.325 $Y=1.765
+ $X2=5.325 $Y2=2.4
r149 25 26 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=5.325 $Y=1.675
+ $X2=5.325 $Y2=1.765
r150 24 54 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=5.325 $Y=1.51
+ $X2=5.325 $Y2=1.345
r151 24 25 64.1371 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=5.325 $Y=1.51
+ $X2=5.325 $Y2=1.675
r152 21 23 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=4.875 $Y=1.765
+ $X2=4.875 $Y2=2.4
r153 20 21 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=4.875 $Y=1.675
+ $X2=4.875 $Y2=1.765
r154 19 53 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=4.875 $Y=1.51
+ $X2=4.875 $Y2=1.345
r155 19 20 64.1371 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=4.875 $Y=1.51
+ $X2=4.875 $Y2=1.675
r156 16 18 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=4.425 $Y=1.765
+ $X2=4.425 $Y2=2.4
r157 15 16 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=4.425 $Y=1.675
+ $X2=4.425 $Y2=1.765
r158 14 50 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=4.425 $Y=1.51
+ $X2=4.425 $Y2=1.345
r159 14 15 64.1371 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=4.425 $Y=1.51
+ $X2=4.425 $Y2=1.675
r160 11 13 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=1.925 $Y=1.185
+ $X2=1.925 $Y2=0.74
r161 10 29 12.1617 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.64 $Y=1.26
+ $X2=1.475 $Y2=1.26
r162 9 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.85 $Y=1.26
+ $X2=1.925 $Y2=1.185
r163 9 10 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=1.85 $Y=1.26
+ $X2=1.64 $Y2=1.26
r164 6 29 13.5877 $w=2.4e-07 $l=8.44097e-08 $layer=POLY_cond $X=1.495 $Y=1.185
+ $X2=1.475 $Y2=1.26
r165 6 8 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=1.495 $Y=1.185
+ $X2=1.495 $Y2=0.74
r166 3 41 53.429 $w=2.79e-07 $l=2.85044e-07 $layer=POLY_cond $X=1.4 $Y=1.765
+ $X2=1.475 $Y2=1.515
r167 3 5 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.4 $Y=1.765 $X2=1.4
+ $Y2=2.4
r168 2 41 1.29086 $w=3.3e-07 $l=1.75152e-07 $layer=POLY_cond $X=1.475 $Y=1.515
+ $X2=1.475 $Y2=1.515
r169 1 29 13.5877 $w=2.4e-07 $l=7.5e-08 $layer=POLY_cond $X=1.475 $Y=1.335
+ $X2=1.475 $Y2=1.26
r170 1 2 31.475 $w=3.3e-07 $l=1.8e-07 $layer=POLY_cond $X=1.475 $Y=1.335
+ $X2=1.475 $Y2=1.515
.ends

.subckt PM_SKY130_FD_SC_HS__NOR3_4%C 1 3 4 5 8 10 12 13 14 17 19 21 22 23 24 26
+ 33 34 35 36 37 38 39 48
c113 13 0 1.16344e-19 $X=2.85 $Y=1.62
c114 1 0 8.47532e-20 $X=2.005 $Y=1.765
r115 48 49 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=5.31
+ $Y=0.505 $X2=5.31 $Y2=0.505
r116 45 48 237.811 $w=3.3e-07 $l=1.36e-06 $layer=POLY_cond $X=3.95 $Y=0.505
+ $X2=5.31 $Y2=0.505
r117 45 46 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=3.95
+ $Y=0.505 $X2=3.95 $Y2=0.505
r118 39 49 7.33373 $w=3.28e-07 $l=2.1e-07 $layer=LI1_cond $X=5.52 $Y=0.505
+ $X2=5.31 $Y2=0.505
r119 38 49 9.42908 $w=3.28e-07 $l=2.7e-07 $layer=LI1_cond $X=5.04 $Y=0.505
+ $X2=5.31 $Y2=0.505
r120 37 38 16.7628 $w=3.28e-07 $l=4.8e-07 $layer=LI1_cond $X=4.56 $Y=0.505
+ $X2=5.04 $Y2=0.505
r121 36 37 16.7628 $w=3.28e-07 $l=4.8e-07 $layer=LI1_cond $X=4.08 $Y=0.505
+ $X2=4.56 $Y2=0.505
r122 36 46 4.53993 $w=3.28e-07 $l=1.3e-07 $layer=LI1_cond $X=4.08 $Y=0.505
+ $X2=3.95 $Y2=0.505
r123 35 45 7.86876 $w=3.3e-07 $l=4.5e-08 $layer=POLY_cond $X=3.905 $Y=0.505
+ $X2=3.95 $Y2=0.505
r124 33 34 31.303 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=3.815 $Y=1.62
+ $X2=3.815 $Y2=1.545
r125 31 32 78.9717 $w=1.77e-07 $l=2.9e-07 $layer=POLY_cond $X=2.925 $Y=1.655
+ $X2=3.215 $Y2=1.655
r126 29 30 27.1897 $w=1.95e-07 $l=1.1e-07 $layer=POLY_cond $X=2.495 $Y=1.655
+ $X2=2.605 $Y2=1.655
r127 27 35 32.1775 $w=3.3e-07 $l=1.98997e-07 $layer=POLY_cond $X=3.83 $Y=0.67
+ $X2=3.905 $Y2=0.505
r128 27 34 448.67 $w=1.5e-07 $l=8.75e-07 $layer=POLY_cond $X=3.83 $Y=0.67
+ $X2=3.83 $Y2=1.545
r129 24 33 58.5127 $w=1.8e-07 $l=1.45e-07 $layer=POLY_cond $X=3.815 $Y=1.765
+ $X2=3.815 $Y2=1.62
r130 24 26 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.815 $Y=1.765
+ $X2=3.815 $Y2=2.4
r131 23 32 25.7691 $w=1.77e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.305 $Y=1.62
+ $X2=3.215 $Y2=1.655
r132 22 33 7.1379 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=3.725 $Y=1.62
+ $X2=3.815 $Y2=1.62
r133 22 23 215.362 $w=1.5e-07 $l=4.2e-07 $layer=POLY_cond $X=3.725 $Y=1.62
+ $X2=3.305 $Y2=1.62
r134 19 32 6.7465 $w=1.5e-07 $l=1.1e-07 $layer=POLY_cond $X=3.215 $Y=1.765
+ $X2=3.215 $Y2=1.655
r135 19 21 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.215 $Y=1.765
+ $X2=3.215 $Y2=2.4
r136 15 31 6.7465 $w=1.5e-07 $l=1.1e-07 $layer=POLY_cond $X=2.925 $Y=1.545
+ $X2=2.925 $Y2=1.655
r137 15 17 412.777 $w=1.5e-07 $l=8.05e-07 $layer=POLY_cond $X=2.925 $Y=1.545
+ $X2=2.925 $Y2=0.74
r138 14 30 24.9362 $w=1.95e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.695 $Y=1.62
+ $X2=2.605 $Y2=1.655
r139 13 31 21.6843 $w=1.77e-07 $l=9.08295e-08 $layer=POLY_cond $X=2.85 $Y=1.62
+ $X2=2.925 $Y2=1.655
r140 13 14 79.4787 $w=1.5e-07 $l=1.55e-07 $layer=POLY_cond $X=2.85 $Y=1.62
+ $X2=2.695 $Y2=1.62
r141 10 30 8.99251 $w=1.5e-07 $l=1.1e-07 $layer=POLY_cond $X=2.605 $Y=1.765
+ $X2=2.605 $Y2=1.655
r142 10 12 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.605 $Y=1.765
+ $X2=2.605 $Y2=2.4
r143 6 29 8.99251 $w=1.5e-07 $l=1.1e-07 $layer=POLY_cond $X=2.495 $Y=1.545
+ $X2=2.495 $Y2=1.655
r144 6 8 412.777 $w=1.5e-07 $l=8.05e-07 $layer=POLY_cond $X=2.495 $Y=1.545
+ $X2=2.495 $Y2=0.74
r145 4 29 21.2285 $w=1.95e-07 $l=9.08295e-08 $layer=POLY_cond $X=2.42 $Y=1.62
+ $X2=2.495 $Y2=1.655
r146 4 5 166.649 $w=1.5e-07 $l=3.25e-07 $layer=POLY_cond $X=2.42 $Y=1.62
+ $X2=2.095 $Y2=1.62
r147 1 5 26.9307 $w=1.5e-07 $l=1.84594e-07 $layer=POLY_cond $X=2.005 $Y=1.765
+ $X2=2.095 $Y2=1.62
r148 1 3 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.005 $Y=1.765
+ $X2=2.005 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_HS__NOR3_4%A_27_368# 1 2 3 4 5 18 22 24 28 30 32 36 38
+ 42 46 48 51 53 60 61
c88 30 0 4.80254e-20 $X=4.485 $Y=2.595
c89 28 0 8.47532e-20 $X=1.175 $Y=2.815
r90 56 57 2.30489 $w=2.48e-07 $l=5e-08 $layer=LI1_cond $X=4.61 $Y=2.545 $X2=4.61
+ $Y2=2.595
r91 53 56 4.60977 $w=2.48e-07 $l=1e-07 $layer=LI1_cond $X=4.61 $Y=2.445 $X2=4.61
+ $Y2=2.545
r92 51 52 7.83661 $w=2.48e-07 $l=1.7e-07 $layer=LI1_cond $X=1.215 $Y=2.425
+ $X2=1.215 $Y2=2.595
r93 44 61 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.49 $Y=2.53 $X2=6.49
+ $Y2=2.445
r94 44 46 13.1378 $w=2.48e-07 $l=2.85e-07 $layer=LI1_cond $X=6.49 $Y=2.53
+ $X2=6.49 $Y2=2.815
r95 40 61 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.49 $Y=2.36 $X2=6.49
+ $Y2=2.445
r96 40 42 17.2866 $w=2.48e-07 $l=3.75e-07 $layer=LI1_cond $X=6.49 $Y=2.36
+ $X2=6.49 $Y2=1.985
r97 39 60 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.635 $Y=2.445
+ $X2=5.55 $Y2=2.445
r98 38 61 2.76166 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.365 $Y=2.445
+ $X2=6.49 $Y2=2.445
r99 38 39 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=6.365 $Y=2.445
+ $X2=5.635 $Y2=2.445
r100 34 60 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.55 $Y=2.53
+ $X2=5.55 $Y2=2.445
r101 34 36 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=5.55 $Y=2.53
+ $X2=5.55 $Y2=2.835
r102 33 53 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.735 $Y=2.445
+ $X2=4.61 $Y2=2.445
r103 32 60 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.465 $Y=2.445
+ $X2=5.55 $Y2=2.445
r104 32 33 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=5.465 $Y=2.445
+ $X2=4.735 $Y2=2.445
r105 31 52 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.34 $Y=2.595
+ $X2=1.215 $Y2=2.595
r106 30 57 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.485 $Y=2.595
+ $X2=4.61 $Y2=2.595
r107 30 31 205.182 $w=1.68e-07 $l=3.145e-06 $layer=LI1_cond $X=4.485 $Y=2.595
+ $X2=1.34 $Y2=2.595
r108 26 52 3.91831 $w=2.48e-07 $l=8.5e-08 $layer=LI1_cond $X=1.215 $Y=2.68
+ $X2=1.215 $Y2=2.595
r109 26 28 6.22319 $w=2.48e-07 $l=1.35e-07 $layer=LI1_cond $X=1.215 $Y=2.68
+ $X2=1.215 $Y2=2.815
r110 25 48 2.76166 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.36 $Y=2.425
+ $X2=0.235 $Y2=2.425
r111 24 51 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.09 $Y=2.425
+ $X2=1.215 $Y2=2.425
r112 24 25 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=1.09 $Y=2.425
+ $X2=0.36 $Y2=2.425
r113 20 48 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.235 $Y=2.51
+ $X2=0.235 $Y2=2.425
r114 20 22 14.0598 $w=2.48e-07 $l=3.05e-07 $layer=LI1_cond $X=0.235 $Y=2.51
+ $X2=0.235 $Y2=2.815
r115 16 48 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.235 $Y=2.34
+ $X2=0.235 $Y2=2.425
r116 16 18 16.3647 $w=2.48e-07 $l=3.55e-07 $layer=LI1_cond $X=0.235 $Y=2.34
+ $X2=0.235 $Y2=1.985
r117 5 46 600 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=6.3
+ $Y=1.84 $X2=6.45 $Y2=2.815
r118 5 42 300 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=2 $X=6.3
+ $Y=1.84 $X2=6.45 $Y2=1.985
r119 4 60 600 $w=1.7e-07 $l=6.75851e-07 $layer=licon1_PDIFF $count=1 $X=5.4
+ $Y=1.84 $X2=5.55 $Y2=2.445
r120 4 36 600 $w=1.7e-07 $l=1.06737e-06 $layer=licon1_PDIFF $count=1 $X=5.4
+ $Y=1.84 $X2=5.55 $Y2=2.835
r121 3 56 600 $w=1.7e-07 $l=7.76386e-07 $layer=licon1_PDIFF $count=1 $X=4.5
+ $Y=1.84 $X2=4.65 $Y2=2.545
r122 2 51 600 $w=1.7e-07 $l=6.55725e-07 $layer=licon1_PDIFF $count=1 $X=1.025
+ $Y=1.84 $X2=1.175 $Y2=2.425
r123 2 28 600 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=1.025
+ $Y=1.84 $X2=1.175 $Y2=2.815
r124 1 22 600 $w=1.7e-07 $l=1.04265e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.275 $Y2=2.815
r125 1 18 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.84 $X2=0.275 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HS__NOR3_4%VPWR 1 2 9 13 15 17 22 32 33 36 39
c69 1 0 1.56752e-19 $X=0.575 $Y=1.84
r70 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r71 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r72 33 40 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=3.33 $X2=6
+ $Y2=3.33
r73 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r74 30 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.165 $Y=3.33 $X2=6
+ $Y2=3.33
r75 30 32 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=6.165 $Y=3.33
+ $X2=6.48 $Y2=3.33
r76 29 40 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=3.33 $X2=6
+ $Y2=3.33
r77 28 29 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r78 26 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r79 25 28 281.84 $w=1.68e-07 $l=4.32e-06 $layer=LI1_cond $X=1.2 $Y=3.33 $X2=5.52
+ $Y2=3.33
r80 25 26 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r81 23 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.89 $Y=3.33
+ $X2=0.725 $Y2=3.33
r82 23 25 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=0.89 $Y=3.33 $X2=1.2
+ $Y2=3.33
r83 22 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.835 $Y=3.33 $X2=6
+ $Y2=3.33
r84 22 28 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=5.835 $Y=3.33
+ $X2=5.52 $Y2=3.33
r85 20 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r86 19 20 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r87 17 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.56 $Y=3.33
+ $X2=0.725 $Y2=3.33
r88 17 19 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=0.56 $Y=3.33 $X2=0.24
+ $Y2=3.33
r89 15 29 0.602067 $w=4.9e-07 $l=2.16e-06 $layer=MET1_cond $X=3.36 $Y=3.33
+ $X2=5.52 $Y2=3.33
r90 15 26 0.602067 $w=4.9e-07 $l=2.16e-06 $layer=MET1_cond $X=3.36 $Y=3.33
+ $X2=1.2 $Y2=3.33
r91 11 39 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6 $Y=3.245 $X2=6
+ $Y2=3.33
r92 11 13 15.5405 $w=3.28e-07 $l=4.45e-07 $layer=LI1_cond $X=6 $Y=3.245 $X2=6
+ $Y2=2.8
r93 7 36 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.725 $Y=3.245
+ $X2=0.725 $Y2=3.33
r94 7 9 15.8897 $w=3.28e-07 $l=4.55e-07 $layer=LI1_cond $X=0.725 $Y=3.245
+ $X2=0.725 $Y2=2.79
r95 2 13 600 $w=1.7e-07 $l=1.03228e-06 $layer=licon1_PDIFF $count=1 $X=5.85
+ $Y=1.84 $X2=6 $Y2=2.8
r96 1 9 600 $w=1.7e-07 $l=1.02225e-06 $layer=licon1_PDIFF $count=1 $X=0.575
+ $Y=1.84 $X2=0.725 $Y2=2.79
.ends

.subckt PM_SKY130_FD_SC_HS__NOR3_4%A_295_368# 1 2 3 4 13 21 23 25
c46 23 0 1.78868e-19 $X=4.285 $Y=2.962
c47 21 0 7.17547e-20 $X=4.935 $Y=2.99
r48 25 27 6.63528 $w=3.28e-07 $l=1.9e-07 $layer=LI1_cond $X=5.1 $Y=2.8 $X2=5.1
+ $Y2=2.99
r49 21 27 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.935 $Y=2.99
+ $X2=5.1 $Y2=2.99
r50 21 23 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=4.935 $Y=2.99
+ $X2=4.285 $Y2=2.99
r51 18 20 61.9758 $w=2.23e-07 $l=1.21e-06 $layer=LI1_cond $X=2.91 $Y=2.962
+ $X2=4.12 $Y2=2.962
r52 15 18 61.7197 $w=2.23e-07 $l=1.205e-06 $layer=LI1_cond $X=1.705 $Y=2.962
+ $X2=2.91 $Y2=2.962
r53 13 23 6.45221 $w=2.23e-07 $l=1.12e-07 $layer=LI1_cond $X=4.173 $Y=2.962
+ $X2=4.285 $Y2=2.962
r54 13 20 2.71464 $w=2.23e-07 $l=5.3e-08 $layer=LI1_cond $X=4.173 $Y=2.962
+ $X2=4.12 $Y2=2.962
r55 4 25 600 $w=1.7e-07 $l=1.03228e-06 $layer=licon1_PDIFF $count=1 $X=4.95
+ $Y=1.84 $X2=5.1 $Y2=2.8
r56 3 20 600 $w=1.7e-07 $l=1.20452e-06 $layer=licon1_PDIFF $count=1 $X=3.89
+ $Y=1.84 $X2=4.12 $Y2=2.935
r57 2 18 600 $w=1.7e-07 $l=1.20452e-06 $layer=licon1_PDIFF $count=1 $X=2.68
+ $Y=1.84 $X2=2.91 $Y2=2.935
r58 1 15 600 $w=1.7e-07 $l=1.20452e-06 $layer=licon1_PDIFF $count=1 $X=1.475
+ $Y=1.84 $X2=1.705 $Y2=2.935
.ends

.subckt PM_SKY130_FD_SC_HS__NOR3_4%Y 1 2 3 4 5 16 17 20 22 30 32 34 37 39 42 45
+ 46 47
c118 39 0 7.79871e-20 $X=1.71 $Y=0.925
c119 37 0 2.08347e-19 $X=5.22 $Y=1.68
c120 34 0 4.80254e-20 $X=5.135 $Y=1.765
c121 16 0 4.22428e-20 $X=1.545 $Y=1.095
r122 44 46 8.46025 $w=3.18e-07 $l=1.65e-07 $layer=LI1_cond $X=3.515 $Y=1.84
+ $X2=3.68 $Y2=1.84
r123 44 45 6.52497 $w=3.18e-07 $l=1.65e-07 $layer=LI1_cond $X=3.515 $Y=1.84
+ $X2=3.35 $Y2=1.84
r124 39 40 5.93683 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=1.71 $Y=0.925
+ $X2=1.71 $Y2=1.095
r125 38 47 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=0.71 $Y=1.01
+ $X2=0.71 $Y2=0.515
r126 36 37 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.22 $Y=1.01
+ $X2=5.22 $Y2=1.68
r127 34 37 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.135 $Y=1.765
+ $X2=5.22 $Y2=1.68
r128 34 46 94.9251 $w=1.68e-07 $l=1.455e-06 $layer=LI1_cond $X=5.135 $Y=1.765
+ $X2=3.68 $Y2=1.765
r129 33 42 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.875 $Y=0.925
+ $X2=2.71 $Y2=0.925
r130 32 36 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.135 $Y=0.925
+ $X2=5.22 $Y2=1.01
r131 32 33 147.444 $w=1.68e-07 $l=2.26e-06 $layer=LI1_cond $X=5.135 $Y=0.925
+ $X2=2.875 $Y2=0.925
r132 28 42 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.71 $Y=0.84
+ $X2=2.71 $Y2=0.925
r133 28 30 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=2.71 $Y=0.84
+ $X2=2.71 $Y2=0.515
r134 26 45 48.1721 $w=2.48e-07 $l=1.045e-06 $layer=LI1_cond $X=2.305 $Y=1.875
+ $X2=3.35 $Y2=1.875
r135 23 39 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.875 $Y=0.925
+ $X2=1.71 $Y2=0.925
r136 22 42 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.545 $Y=0.925
+ $X2=2.71 $Y2=0.925
r137 22 23 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.545 $Y=0.925
+ $X2=1.875 $Y2=0.925
r138 18 39 2.96841 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=1.71 $Y=0.84
+ $X2=1.71 $Y2=0.925
r139 18 20 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=1.71 $Y=0.84
+ $X2=1.71 $Y2=0.515
r140 17 38 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.875 $Y=1.095
+ $X2=0.71 $Y2=1.01
r141 16 40 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.545 $Y=1.095
+ $X2=1.71 $Y2=1.095
r142 16 17 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.545 $Y=1.095
+ $X2=0.875 $Y2=1.095
r143 5 44 600 $w=1.7e-07 $l=2.59808e-07 $layer=licon1_PDIFF $count=1 $X=3.29
+ $Y=1.84 $X2=3.515 $Y2=1.915
r144 4 26 600 $w=1.7e-07 $l=2.59808e-07 $layer=licon1_PDIFF $count=1 $X=2.08
+ $Y=1.84 $X2=2.305 $Y2=1.915
r145 3 30 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.57
+ $Y=0.37 $X2=2.71 $Y2=0.515
r146 2 20 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.57
+ $Y=0.37 $X2=1.71 $Y2=0.515
r147 1 47 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=0.57
+ $Y=0.37 $X2=0.71 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__NOR3_4%VGND 1 2 3 4 13 15 19 23 25 29 31 33 38 48 49
+ 55 58 61
r62 61 62 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r63 59 62 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=3.12
+ $Y2=0
r64 58 59 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r65 55 56 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r66 52 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r67 48 49 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=6.48 $Y=0
+ $X2=6.48 $Y2=0
r68 46 49 0.802756 $w=4.9e-07 $l=2.88e-06 $layer=MET1_cond $X=3.6 $Y=0 $X2=6.48
+ $Y2=0
r69 45 48 187.893 $w=1.68e-07 $l=2.88e-06 $layer=LI1_cond $X=3.6 $Y=0 $X2=6.48
+ $Y2=0
r70 45 46 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=3.6 $Y=0
+ $X2=3.6 $Y2=0
r71 43 61 8.23795 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=3.365 $Y=0 $X2=3.21
+ $Y2=0
r72 43 45 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=3.365 $Y=0 $X2=3.6
+ $Y2=0
r73 42 59 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r74 42 56 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r75 41 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r76 39 55 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.375 $Y=0 $X2=1.21
+ $Y2=0
r77 39 41 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.375 $Y=0 $X2=1.68
+ $Y2=0
r78 38 58 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.045 $Y=0 $X2=2.21
+ $Y2=0
r79 38 41 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=2.045 $Y=0 $X2=1.68
+ $Y2=0
r80 37 56 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r81 37 53 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r82 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r83 34 52 4.00981 $w=1.7e-07 $l=1.83e-07 $layer=LI1_cond $X=0.365 $Y=0 $X2=0.182
+ $Y2=0
r84 34 36 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=0.365 $Y=0 $X2=0.72
+ $Y2=0
r85 33 55 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.045 $Y=0 $X2=1.21
+ $Y2=0
r86 33 36 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=1.045 $Y=0 $X2=0.72
+ $Y2=0
r87 31 46 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=3.36 $Y=0 $X2=3.6
+ $Y2=0
r88 31 62 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=3.36 $Y=0 $X2=3.12
+ $Y2=0
r89 27 61 0.701276 $w=3.1e-07 $l=8.5e-08 $layer=LI1_cond $X=3.21 $Y=0.085
+ $X2=3.21 $Y2=0
r90 27 29 15.6137 $w=3.08e-07 $l=4.2e-07 $layer=LI1_cond $X=3.21 $Y=0.085
+ $X2=3.21 $Y2=0.505
r91 26 58 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.375 $Y=0 $X2=2.21
+ $Y2=0
r92 25 61 8.23795 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=3.055 $Y=0 $X2=3.21
+ $Y2=0
r93 25 26 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=3.055 $Y=0 $X2=2.375
+ $Y2=0
r94 21 58 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.21 $Y=0.085
+ $X2=2.21 $Y2=0
r95 21 23 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=2.21 $Y=0.085
+ $X2=2.21 $Y2=0.55
r96 17 55 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.21 $Y=0.085
+ $X2=1.21 $Y2=0
r97 17 19 20.6043 $w=3.28e-07 $l=5.9e-07 $layer=LI1_cond $X=1.21 $Y=0.085
+ $X2=1.21 $Y2=0.675
r98 13 52 3.13335 $w=2.5e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.24 $Y=0.085
+ $X2=0.182 $Y2=0
r99 13 15 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=0.24 $Y=0.085
+ $X2=0.24 $Y2=0.515
r100 4 29 182 $w=1.7e-07 $l=1.96214e-07 $layer=licon1_NDIFF $count=1 $X=3
+ $Y=0.37 $X2=3.14 $Y2=0.505
r101 3 23 182 $w=1.7e-07 $l=2.86182e-07 $layer=licon1_NDIFF $count=1 $X=2
+ $Y=0.37 $X2=2.21 $Y2=0.55
r102 2 19 182 $w=1.7e-07 $l=3.9246e-07 $layer=licon1_NDIFF $count=1 $X=1.01
+ $Y=0.37 $X2=1.21 $Y2=0.675
r103 1 15 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.515
.ends

