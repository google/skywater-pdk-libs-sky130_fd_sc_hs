* File: sky130_fd_sc_hs__o2bb2ai_4.pex.spice
* Created: Thu Aug 27 21:01:30 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HS__O2BB2AI_4%A1_N 3 5 7 10 12 14 17 19 21 24 26 28 29
+ 30 31 32 47 48
c83 47 0 9.27533e-20 $X=1.77 $Y=1.515
c84 26 0 1.62199e-20 $X=1.845 $Y=1.765
c85 24 0 8.01953e-20 $X=1.795 $Y=0.74
r86 48 49 6.5847 $w=3.66e-07 $l=5e-08 $layer=POLY_cond $X=1.795 $Y=1.557
+ $X2=1.845 $Y2=1.557
r87 46 48 3.29235 $w=3.66e-07 $l=2.5e-08 $layer=POLY_cond $X=1.77 $Y=1.557
+ $X2=1.795 $Y2=1.557
r88 46 47 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=1.77
+ $Y=1.515 $X2=1.77 $Y2=1.515
r89 44 46 49.3852 $w=3.66e-07 $l=3.75e-07 $layer=POLY_cond $X=1.395 $Y=1.557
+ $X2=1.77 $Y2=1.557
r90 43 44 3.95082 $w=3.66e-07 $l=3e-08 $layer=POLY_cond $X=1.365 $Y=1.557
+ $X2=1.395 $Y2=1.557
r91 42 43 55.3115 $w=3.66e-07 $l=4.2e-07 $layer=POLY_cond $X=0.945 $Y=1.557
+ $X2=1.365 $Y2=1.557
r92 41 42 2.63388 $w=3.66e-07 $l=2e-08 $layer=POLY_cond $X=0.925 $Y=1.557
+ $X2=0.945 $Y2=1.557
r93 40 41 56.6284 $w=3.66e-07 $l=4.3e-07 $layer=POLY_cond $X=0.495 $Y=1.557
+ $X2=0.925 $Y2=1.557
r94 38 40 11.194 $w=3.66e-07 $l=8.5e-08 $layer=POLY_cond $X=0.41 $Y=1.557
+ $X2=0.495 $Y2=1.557
r95 38 39 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=0.41
+ $Y=1.515 $X2=0.41 $Y2=1.515
r96 32 47 2.41209 $w=4.28e-07 $l=9e-08 $layer=LI1_cond $X=1.68 $Y=1.565 $X2=1.77
+ $Y2=1.565
r97 31 32 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=1.2 $Y=1.565
+ $X2=1.68 $Y2=1.565
r98 30 31 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=0.72 $Y=1.565
+ $X2=1.2 $Y2=1.565
r99 30 39 8.30831 $w=4.28e-07 $l=3.1e-07 $layer=LI1_cond $X=0.72 $Y=1.565
+ $X2=0.41 $Y2=1.565
r100 29 39 4.55617 $w=4.28e-07 $l=1.7e-07 $layer=LI1_cond $X=0.24 $Y=1.565
+ $X2=0.41 $Y2=1.565
r101 26 49 23.7042 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=1.845 $Y=1.765
+ $X2=1.845 $Y2=1.557
r102 26 28 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.845 $Y=1.765
+ $X2=1.845 $Y2=2.4
r103 22 48 23.7042 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.795 $Y=1.35
+ $X2=1.795 $Y2=1.557
r104 22 24 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.795 $Y=1.35
+ $X2=1.795 $Y2=0.74
r105 19 44 23.7042 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=1.395 $Y=1.765
+ $X2=1.395 $Y2=1.557
r106 19 21 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.395 $Y=1.765
+ $X2=1.395 $Y2=2.4
r107 15 43 23.7042 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.365 $Y=1.35
+ $X2=1.365 $Y2=1.557
r108 15 17 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.365 $Y=1.35
+ $X2=1.365 $Y2=0.74
r109 12 42 23.7042 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=0.945 $Y=1.765
+ $X2=0.945 $Y2=1.557
r110 12 14 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.945 $Y=1.765
+ $X2=0.945 $Y2=2.4
r111 8 41 23.7042 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.925 $Y=1.35
+ $X2=0.925 $Y2=1.557
r112 8 10 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=0.925 $Y=1.35
+ $X2=0.925 $Y2=0.74
r113 5 40 23.7042 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=0.495 $Y=1.765
+ $X2=0.495 $Y2=1.557
r114 5 7 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.495 $Y=1.765
+ $X2=0.495 $Y2=2.4
r115 1 40 23.7042 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.495 $Y=1.35
+ $X2=0.495 $Y2=1.557
r116 1 3 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=0.495 $Y=1.35
+ $X2=0.495 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HS__O2BB2AI_4%A2_N 3 5 7 10 12 14 17 19 21 22 23 24 26
+ 29 32 33
c95 33 0 1.62199e-20 $X=3.12 $Y=1.665
c96 24 0 1.0348e-19 $X=3.645 $Y=1.765
c97 5 0 9.27533e-20 $X=2.295 $Y=1.765
c98 3 0 1.9142e-19 $X=2.225 $Y=0.74
r99 46 47 1.8075 $w=4e-07 $l=1.5e-08 $layer=POLY_cond $X=3.18 $Y=1.542 $X2=3.195
+ $Y2=1.542
r100 44 46 13.255 $w=4e-07 $l=1.1e-07 $layer=POLY_cond $X=3.07 $Y=1.542 $X2=3.18
+ $Y2=1.542
r101 44 45 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=3.07
+ $Y=1.515 $X2=3.07 $Y2=1.515
r102 42 44 39.1625 $w=4e-07 $l=3.25e-07 $layer=POLY_cond $X=2.745 $Y=1.542
+ $X2=3.07 $Y2=1.542
r103 41 42 10.845 $w=4e-07 $l=9e-08 $layer=POLY_cond $X=2.655 $Y=1.542 $X2=2.745
+ $Y2=1.542
r104 39 41 31.9325 $w=4e-07 $l=2.65e-07 $layer=POLY_cond $X=2.39 $Y=1.542
+ $X2=2.655 $Y2=1.542
r105 39 40 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=2.39
+ $Y=1.515 $X2=2.39 $Y2=1.515
r106 37 39 11.4475 $w=4e-07 $l=9.5e-08 $layer=POLY_cond $X=2.295 $Y=1.542
+ $X2=2.39 $Y2=1.542
r107 36 37 8.435 $w=4e-07 $l=7e-08 $layer=POLY_cond $X=2.225 $Y=1.542 $X2=2.295
+ $Y2=1.542
r108 33 45 1.34005 $w=4.28e-07 $l=5e-08 $layer=LI1_cond $X=3.12 $Y=1.565
+ $X2=3.07 $Y2=1.565
r109 32 45 11.5244 $w=4.28e-07 $l=4.3e-07 $layer=LI1_cond $X=2.64 $Y=1.565
+ $X2=3.07 $Y2=1.565
r110 32 40 6.70025 $w=4.28e-07 $l=2.5e-07 $layer=LI1_cond $X=2.64 $Y=1.565
+ $X2=2.39 $Y2=1.565
r111 27 31 21.642 $w=1.78e-07 $l=7.98436e-08 $layer=POLY_cond $X=3.655 $Y=1.32
+ $X2=3.645 $Y2=1.395
r112 27 29 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=3.655 $Y=1.32
+ $X2=3.655 $Y2=0.74
r113 24 31 101.524 $w=1.78e-07 $l=3.7e-07 $layer=POLY_cond $X=3.645 $Y=1.765
+ $X2=3.645 $Y2=1.395
r114 24 26 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.645 $Y=1.765
+ $X2=3.645 $Y2=2.4
r115 23 47 30.5478 $w=4e-07 $l=1.86652e-07 $layer=POLY_cond $X=3.285 $Y=1.395
+ $X2=3.195 $Y2=1.542
r116 22 31 6.87779 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=3.555 $Y=1.395
+ $X2=3.645 $Y2=1.395
r117 22 23 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=3.555 $Y=1.395
+ $X2=3.285 $Y2=1.395
r118 19 47 25.8619 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=3.195 $Y=1.765
+ $X2=3.195 $Y2=1.542
r119 19 21 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.195 $Y=1.765
+ $X2=3.195 $Y2=2.4
r120 15 46 25.8619 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=3.18 $Y=1.32
+ $X2=3.18 $Y2=1.542
r121 15 17 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=3.18 $Y=1.32
+ $X2=3.18 $Y2=0.74
r122 12 42 25.8619 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=2.745 $Y=1.765
+ $X2=2.745 $Y2=1.542
r123 12 14 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.745 $Y=1.765
+ $X2=2.745 $Y2=2.4
r124 8 41 25.8619 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=2.655 $Y=1.32
+ $X2=2.655 $Y2=1.542
r125 8 10 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=2.655 $Y=1.32
+ $X2=2.655 $Y2=0.74
r126 5 37 25.8619 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=2.295 $Y=1.765
+ $X2=2.295 $Y2=1.542
r127 5 7 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.295 $Y=1.765
+ $X2=2.295 $Y2=2.4
r128 1 36 25.8619 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=2.225 $Y=1.32
+ $X2=2.225 $Y2=1.542
r129 1 3 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=2.225 $Y=1.32
+ $X2=2.225 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HS__O2BB2AI_4%A_114_368# 1 2 3 4 5 6 19 21 22 24 27 29
+ 31 34 36 38 41 43 44 47 49 51 53 57 59 63 67 69 70 71 75 79 81 82 88 94 96 98
c207 82 0 1.74044e-19 $X=3.5 $Y=1.95
c208 70 0 8.01953e-20 $X=2.605 $Y=1.095
c209 47 0 1.9142e-19 $X=5.935 $Y=0.74
c210 44 0 1.50249e-19 $X=5.58 $Y=1.375
r211 108 109 7.57068 $w=3.82e-07 $l=6e-08 $layer=POLY_cond $X=5.445 $Y=1.532
+ $X2=5.505 $Y2=1.532
r212 105 106 10.0942 $w=3.82e-07 $l=8e-08 $layer=POLY_cond $X=4.995 $Y=1.532
+ $X2=5.075 $Y2=1.532
r213 104 105 44.1623 $w=3.82e-07 $l=3.5e-07 $layer=POLY_cond $X=4.645 $Y=1.532
+ $X2=4.995 $Y2=1.532
r214 103 104 12.6178 $w=3.82e-07 $l=1e-07 $layer=POLY_cond $X=4.545 $Y=1.532
+ $X2=4.645 $Y2=1.532
r215 89 108 23.3429 $w=3.82e-07 $l=1.85e-07 $layer=POLY_cond $X=5.26 $Y=1.532
+ $X2=5.445 $Y2=1.532
r216 89 106 23.3429 $w=3.82e-07 $l=1.85e-07 $layer=POLY_cond $X=5.26 $Y=1.532
+ $X2=5.075 $Y2=1.532
r217 88 89 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.26
+ $Y=1.465 $X2=5.26 $Y2=1.465
r218 86 103 38.4843 $w=3.82e-07 $l=3.05e-07 $layer=POLY_cond $X=4.24 $Y=1.532
+ $X2=4.545 $Y2=1.532
r219 86 101 18.2958 $w=3.82e-07 $l=1.45e-07 $layer=POLY_cond $X=4.24 $Y=1.532
+ $X2=4.095 $Y2=1.532
r220 85 88 35.621 $w=3.28e-07 $l=1.02e-06 $layer=LI1_cond $X=4.24 $Y=1.465
+ $X2=5.26 $Y2=1.465
r221 85 86 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.24
+ $Y=1.465 $X2=4.24 $Y2=1.465
r222 83 99 19.7982 $w=2.28e-07 $l=3.7e-07 $layer=LI1_cond $X=3.44 $Y=1.465
+ $X2=3.44 $Y2=1.095
r223 83 85 22.1758 $w=3.28e-07 $l=6.35e-07 $layer=LI1_cond $X=3.605 $Y=1.465
+ $X2=4.24 $Y2=1.465
r224 82 98 3.70735 $w=2.5e-07 $l=1.18427e-07 $layer=LI1_cond $X=3.5 $Y=1.95
+ $X2=3.42 $Y2=2.035
r225 81 83 9.64481 $w=2.28e-07 $l=1.92678e-07 $layer=LI1_cond $X=3.5 $Y=1.63
+ $X2=3.44 $Y2=1.465
r226 81 82 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=3.5 $Y=1.63 $X2=3.5
+ $Y2=1.95
r227 77 99 4.31892 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.44 $Y=1.01
+ $X2=3.44 $Y2=1.095
r228 77 79 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=3.44 $Y=1.01
+ $X2=3.44 $Y2=0.86
r229 73 98 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.42 $Y=2.12
+ $X2=3.42 $Y2=2.035
r230 73 75 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=3.42 $Y=2.12
+ $X2=3.42 $Y2=2.815
r231 72 96 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.685 $Y=2.035
+ $X2=2.52 $Y2=2.035
r232 71 98 2.76166 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.255 $Y=2.035
+ $X2=3.42 $Y2=2.035
r233 71 72 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=3.255 $Y=2.035
+ $X2=2.685 $Y2=2.035
r234 69 99 2.45823 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.275 $Y=1.095
+ $X2=3.44 $Y2=1.095
r235 69 70 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.275 $Y=1.095
+ $X2=2.605 $Y2=1.095
r236 65 96 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.52 $Y=2.12
+ $X2=2.52 $Y2=2.035
r237 65 67 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=2.52 $Y=2.12
+ $X2=2.52 $Y2=2.815
r238 61 70 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.44 $Y=1.01
+ $X2=2.605 $Y2=1.095
r239 61 63 6.63528 $w=3.28e-07 $l=1.9e-07 $layer=LI1_cond $X=2.44 $Y=1.01
+ $X2=2.44 $Y2=0.82
r240 60 94 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.785 $Y=2.035
+ $X2=1.62 $Y2=2.035
r241 59 96 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.355 $Y=2.035
+ $X2=2.52 $Y2=2.035
r242 59 60 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=2.355 $Y=2.035
+ $X2=1.785 $Y2=2.035
r243 55 94 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.62 $Y=2.12
+ $X2=1.62 $Y2=2.035
r244 55 57 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=1.62 $Y=2.12
+ $X2=1.62 $Y2=2.815
r245 54 92 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.885 $Y=2.035
+ $X2=0.72 $Y2=2.035
r246 53 94 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.455 $Y=2.035
+ $X2=1.62 $Y2=2.035
r247 53 54 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=1.455 $Y=2.035
+ $X2=0.885 $Y2=2.035
r248 49 92 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.72 $Y=2.12 $X2=0.72
+ $Y2=2.035
r249 49 51 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=0.72 $Y=2.12
+ $X2=0.72 $Y2=2.815
r250 45 47 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=5.935 $Y=1.3
+ $X2=5.935 $Y2=0.74
r251 44 109 27.8964 $w=3.82e-07 $l=1.90851e-07 $layer=POLY_cond $X=5.58 $Y=1.375
+ $X2=5.505 $Y2=1.532
r252 43 45 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.86 $Y=1.375
+ $X2=5.935 $Y2=1.3
r253 43 44 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=5.86 $Y=1.375
+ $X2=5.58 $Y2=1.375
r254 39 109 24.74 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=5.505 $Y=1.3
+ $X2=5.505 $Y2=1.532
r255 39 41 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=5.505 $Y=1.3
+ $X2=5.505 $Y2=0.74
r256 36 108 24.74 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=5.445 $Y=1.765
+ $X2=5.445 $Y2=1.532
r257 36 38 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=5.445 $Y=1.765
+ $X2=5.445 $Y2=2.4
r258 32 106 24.74 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=5.075 $Y=1.3
+ $X2=5.075 $Y2=1.532
r259 32 34 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=5.075 $Y=1.3
+ $X2=5.075 $Y2=0.74
r260 29 105 24.74 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=4.995 $Y=1.765
+ $X2=4.995 $Y2=1.532
r261 29 31 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=4.995 $Y=1.765
+ $X2=4.995 $Y2=2.4
r262 25 104 24.74 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=4.645 $Y=1.3
+ $X2=4.645 $Y2=1.532
r263 25 27 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=4.645 $Y=1.3
+ $X2=4.645 $Y2=0.74
r264 22 103 24.74 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=4.545 $Y=1.765
+ $X2=4.545 $Y2=1.532
r265 22 24 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=4.545 $Y=1.765
+ $X2=4.545 $Y2=2.4
r266 19 101 24.74 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=4.095 $Y=1.765
+ $X2=4.095 $Y2=1.532
r267 19 21 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=4.095 $Y=1.765
+ $X2=4.095 $Y2=2.4
r268 6 98 400 $w=1.7e-07 $l=2.59374e-07 $layer=licon1_PDIFF $count=1 $X=3.27
+ $Y=1.84 $X2=3.42 $Y2=2.035
r269 6 75 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=3.27
+ $Y=1.84 $X2=3.42 $Y2=2.815
r270 5 96 400 $w=1.7e-07 $l=2.59374e-07 $layer=licon1_PDIFF $count=1 $X=2.37
+ $Y=1.84 $X2=2.52 $Y2=2.035
r271 5 67 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=2.37
+ $Y=1.84 $X2=2.52 $Y2=2.815
r272 4 94 400 $w=1.7e-07 $l=2.59374e-07 $layer=licon1_PDIFF $count=1 $X=1.47
+ $Y=1.84 $X2=1.62 $Y2=2.035
r273 4 57 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=1.47
+ $Y=1.84 $X2=1.62 $Y2=2.815
r274 3 92 400 $w=1.7e-07 $l=2.59374e-07 $layer=licon1_PDIFF $count=1 $X=0.57
+ $Y=1.84 $X2=0.72 $Y2=2.035
r275 3 51 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=0.57
+ $Y=1.84 $X2=0.72 $Y2=2.815
r276 2 79 182 $w=1.7e-07 $l=5.75109e-07 $layer=licon1_NDIFF $count=1 $X=3.255
+ $Y=0.37 $X2=3.44 $Y2=0.86
r277 1 63 182 $w=1.7e-07 $l=5.15267e-07 $layer=licon1_NDIFF $count=1 $X=2.3
+ $Y=0.37 $X2=2.44 $Y2=0.82
.ends

.subckt PM_SKY130_FD_SC_HS__O2BB2AI_4%B2 3 5 7 10 12 14 17 19 21 22 24 27 29 30
+ 31 32 48 49
c91 22 0 3.11558e-19 $X=7.785 $Y=1.765
c92 3 0 2.29387e-19 $X=6.365 $Y=0.74
r93 49 50 1.30978 $w=3.68e-07 $l=1e-08 $layer=POLY_cond $X=7.785 $Y=1.557
+ $X2=7.795 $Y2=1.557
r94 47 49 40.6033 $w=3.68e-07 $l=3.1e-07 $layer=POLY_cond $X=7.475 $Y=1.557
+ $X2=7.785 $Y2=1.557
r95 47 48 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=7.475
+ $Y=1.515 $X2=7.475 $Y2=1.515
r96 45 47 18.337 $w=3.68e-07 $l=1.4e-07 $layer=POLY_cond $X=7.335 $Y=1.557
+ $X2=7.475 $Y2=1.557
r97 44 45 5.23913 $w=3.68e-07 $l=4e-08 $layer=POLY_cond $X=7.295 $Y=1.557
+ $X2=7.335 $Y2=1.557
r98 43 44 53.7011 $w=3.68e-07 $l=4.1e-07 $layer=POLY_cond $X=6.885 $Y=1.557
+ $X2=7.295 $Y2=1.557
r99 42 43 2.61957 $w=3.68e-07 $l=2e-08 $layer=POLY_cond $X=6.865 $Y=1.557
+ $X2=6.885 $Y2=1.557
r100 40 42 53.7011 $w=3.68e-07 $l=4.1e-07 $layer=POLY_cond $X=6.455 $Y=1.557
+ $X2=6.865 $Y2=1.557
r101 40 41 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.455
+ $Y=1.515 $X2=6.455 $Y2=1.515
r102 38 40 2.61957 $w=3.68e-07 $l=2e-08 $layer=POLY_cond $X=6.435 $Y=1.557
+ $X2=6.455 $Y2=1.557
r103 37 38 9.16848 $w=3.68e-07 $l=7e-08 $layer=POLY_cond $X=6.365 $Y=1.557
+ $X2=6.435 $Y2=1.557
r104 32 48 0.938035 $w=4.28e-07 $l=3.5e-08 $layer=LI1_cond $X=7.44 $Y=1.565
+ $X2=7.475 $Y2=1.565
r105 31 32 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=6.96 $Y=1.565
+ $X2=7.44 $Y2=1.565
r106 30 31 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=6.48 $Y=1.565
+ $X2=6.96 $Y2=1.565
r107 30 41 0.670025 $w=4.28e-07 $l=2.5e-08 $layer=LI1_cond $X=6.48 $Y=1.565
+ $X2=6.455 $Y2=1.565
r108 29 41 12.1945 $w=4.28e-07 $l=4.55e-07 $layer=LI1_cond $X=6 $Y=1.565
+ $X2=6.455 $Y2=1.565
r109 25 50 23.8357 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=7.795 $Y=1.35
+ $X2=7.795 $Y2=1.557
r110 25 27 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=7.795 $Y=1.35
+ $X2=7.795 $Y2=0.74
r111 22 49 23.8357 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=7.785 $Y=1.765
+ $X2=7.785 $Y2=1.557
r112 22 24 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=7.785 $Y=1.765
+ $X2=7.785 $Y2=2.4
r113 19 45 23.8357 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=7.335 $Y=1.765
+ $X2=7.335 $Y2=1.557
r114 19 21 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=7.335 $Y=1.765
+ $X2=7.335 $Y2=2.4
r115 15 44 23.8357 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=7.295 $Y=1.35
+ $X2=7.295 $Y2=1.557
r116 15 17 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=7.295 $Y=1.35
+ $X2=7.295 $Y2=0.74
r117 12 43 23.8357 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=6.885 $Y=1.765
+ $X2=6.885 $Y2=1.557
r118 12 14 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=6.885 $Y=1.765
+ $X2=6.885 $Y2=2.4
r119 8 42 23.8357 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=6.865 $Y=1.35
+ $X2=6.865 $Y2=1.557
r120 8 10 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=6.865 $Y=1.35
+ $X2=6.865 $Y2=0.74
r121 5 38 23.8357 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=6.435 $Y=1.765
+ $X2=6.435 $Y2=1.557
r122 5 7 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=6.435 $Y=1.765
+ $X2=6.435 $Y2=2.4
r123 1 37 23.8357 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=6.365 $Y=1.35
+ $X2=6.365 $Y2=1.557
r124 1 3 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=6.365 $Y=1.35
+ $X2=6.365 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HS__O2BB2AI_4%B1 3 5 7 10 12 14 17 19 21 24 26 28 29 30
+ 31 32 46
c81 32 0 1.2677e-19 $X=9.84 $Y=1.665
r82 48 49 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=9.675
+ $Y=1.515 $X2=9.675 $Y2=1.515
r83 46 48 11.8849 $w=3.65e-07 $l=9e-08 $layer=POLY_cond $X=9.585 $Y=1.557
+ $X2=9.675 $Y2=1.557
r84 45 46 59.4247 $w=3.65e-07 $l=4.5e-07 $layer=POLY_cond $X=9.135 $Y=1.557
+ $X2=9.585 $Y2=1.557
r85 44 45 6.60274 $w=3.65e-07 $l=5e-08 $layer=POLY_cond $X=9.085 $Y=1.557
+ $X2=9.135 $Y2=1.557
r86 43 44 52.8219 $w=3.65e-07 $l=4e-07 $layer=POLY_cond $X=8.685 $Y=1.557
+ $X2=9.085 $Y2=1.557
r87 42 43 3.96164 $w=3.65e-07 $l=3e-08 $layer=POLY_cond $X=8.655 $Y=1.557
+ $X2=8.685 $Y2=1.557
r88 40 42 44.8986 $w=3.65e-07 $l=3.4e-07 $layer=POLY_cond $X=8.315 $Y=1.557
+ $X2=8.655 $Y2=1.557
r89 40 41 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=8.315
+ $Y=1.515 $X2=8.315 $Y2=1.515
r90 38 40 10.5644 $w=3.65e-07 $l=8e-08 $layer=POLY_cond $X=8.235 $Y=1.557
+ $X2=8.315 $Y2=1.557
r91 37 38 1.32055 $w=3.65e-07 $l=1e-08 $layer=POLY_cond $X=8.225 $Y=1.557
+ $X2=8.235 $Y2=1.557
r92 32 49 4.42216 $w=4.28e-07 $l=1.65e-07 $layer=LI1_cond $X=9.84 $Y=1.565
+ $X2=9.675 $Y2=1.565
r93 31 49 8.44232 $w=4.28e-07 $l=3.15e-07 $layer=LI1_cond $X=9.36 $Y=1.565
+ $X2=9.675 $Y2=1.565
r94 30 31 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=8.88 $Y=1.565
+ $X2=9.36 $Y2=1.565
r95 29 30 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=8.4 $Y=1.565
+ $X2=8.88 $Y2=1.565
r96 29 41 2.27808 $w=4.28e-07 $l=8.5e-08 $layer=LI1_cond $X=8.4 $Y=1.565
+ $X2=8.315 $Y2=1.565
r97 26 46 23.6381 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=9.585 $Y=1.765
+ $X2=9.585 $Y2=1.557
r98 26 28 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=9.585 $Y=1.765
+ $X2=9.585 $Y2=2.4
r99 22 46 23.6381 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=9.585 $Y=1.35
+ $X2=9.585 $Y2=1.557
r100 22 24 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=9.585 $Y=1.35
+ $X2=9.585 $Y2=0.74
r101 19 45 23.6381 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=9.135 $Y=1.765
+ $X2=9.135 $Y2=1.557
r102 19 21 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=9.135 $Y=1.765
+ $X2=9.135 $Y2=2.4
r103 15 44 23.6381 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=9.085 $Y=1.35
+ $X2=9.085 $Y2=1.557
r104 15 17 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=9.085 $Y=1.35
+ $X2=9.085 $Y2=0.74
r105 12 43 23.6381 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=8.685 $Y=1.765
+ $X2=8.685 $Y2=1.557
r106 12 14 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=8.685 $Y=1.765
+ $X2=8.685 $Y2=2.4
r107 8 42 23.6381 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=8.655 $Y=1.35
+ $X2=8.655 $Y2=1.557
r108 8 10 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=8.655 $Y=1.35
+ $X2=8.655 $Y2=0.74
r109 5 38 23.6381 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=8.235 $Y=1.765
+ $X2=8.235 $Y2=1.557
r110 5 7 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=8.235 $Y=1.765
+ $X2=8.235 $Y2=2.4
r111 1 37 23.6381 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=8.225 $Y=1.35
+ $X2=8.225 $Y2=1.557
r112 1 3 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=8.225 $Y=1.35
+ $X2=8.225 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HS__O2BB2AI_4%VPWR 1 2 3 4 5 6 7 8 9 28 30 36 40 44 48
+ 54 56 60 64 68 71 72 74 75 77 78 80 81 82 83 84 102 110 117 118 124 127 130
c153 64 0 1.84789e-19 $X=8.46 $Y=2.455
r154 130 131 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.36 $Y=3.33
+ $X2=9.36 $Y2=3.33
r155 127 128 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=3.33
+ $X2=8.4 $Y2=3.33
r156 124 125 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r157 121 122 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r158 118 131 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.84 $Y=3.33
+ $X2=9.36 $Y2=3.33
r159 117 118 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.84 $Y=3.33
+ $X2=9.84 $Y2=3.33
r160 115 130 6.01921 $w=1.7e-07 $l=1.03e-07 $layer=LI1_cond $X=9.465 $Y=3.33
+ $X2=9.362 $Y2=3.33
r161 115 117 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=9.465 $Y=3.33
+ $X2=9.84 $Y2=3.33
r162 114 131 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=3.33
+ $X2=9.36 $Y2=3.33
r163 114 128 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=3.33
+ $X2=8.4 $Y2=3.33
r164 113 114 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r165 111 127 7.34436 $w=1.7e-07 $l=1.33e-07 $layer=LI1_cond $X=8.56 $Y=3.33
+ $X2=8.427 $Y2=3.33
r166 111 113 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=8.56 $Y=3.33
+ $X2=8.88 $Y2=3.33
r167 110 130 6.01921 $w=1.7e-07 $l=1.02e-07 $layer=LI1_cond $X=9.26 $Y=3.33
+ $X2=9.362 $Y2=3.33
r168 110 113 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=9.26 $Y=3.33
+ $X2=8.88 $Y2=3.33
r169 109 128 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=3.33
+ $X2=8.4 $Y2=3.33
r170 108 109 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r171 106 109 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=6 $Y=3.33
+ $X2=7.92 $Y2=3.33
r172 106 125 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=3.33
+ $X2=5.52 $Y2=3.33
r173 105 108 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=6 $Y=3.33
+ $X2=7.92 $Y2=3.33
r174 105 106 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r175 103 124 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.835 $Y=3.33
+ $X2=5.67 $Y2=3.33
r176 103 105 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=5.835 $Y=3.33
+ $X2=6 $Y2=3.33
r177 102 127 7.34436 $w=1.7e-07 $l=1.32e-07 $layer=LI1_cond $X=8.295 $Y=3.33
+ $X2=8.427 $Y2=3.33
r178 102 108 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=8.295 $Y=3.33
+ $X2=7.92 $Y2=3.33
r179 100 101 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r180 98 101 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.56 $Y2=3.33
r181 97 98 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r182 95 98 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.6 $Y2=3.33
r183 94 95 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r184 92 95 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.64 $Y2=3.33
r185 91 92 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r186 89 92 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.68 $Y2=3.33
r187 89 122 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r188 88 89 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r189 86 121 4.02368 $w=1.7e-07 $l=1.78e-07 $layer=LI1_cond $X=0.355 $Y=3.33
+ $X2=0.177 $Y2=3.33
r190 86 88 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=0.355 $Y=3.33
+ $X2=0.72 $Y2=3.33
r191 84 125 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=5.52 $Y2=3.33
r192 84 101 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=4.56 $Y2=3.33
r193 82 100 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=4.685 $Y=3.33
+ $X2=4.56 $Y2=3.33
r194 82 83 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.685 $Y=3.33
+ $X2=4.77 $Y2=3.33
r195 80 97 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=3.785 $Y=3.33
+ $X2=3.6 $Y2=3.33
r196 80 81 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.785 $Y=3.33
+ $X2=3.87 $Y2=3.33
r197 79 100 39.4706 $w=1.68e-07 $l=6.05e-07 $layer=LI1_cond $X=3.955 $Y=3.33
+ $X2=4.56 $Y2=3.33
r198 79 81 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.955 $Y=3.33
+ $X2=3.87 $Y2=3.33
r199 77 94 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=2.885 $Y=3.33
+ $X2=2.64 $Y2=3.33
r200 77 78 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.885 $Y=3.33
+ $X2=2.97 $Y2=3.33
r201 76 97 35.5561 $w=1.68e-07 $l=5.45e-07 $layer=LI1_cond $X=3.055 $Y=3.33
+ $X2=3.6 $Y2=3.33
r202 76 78 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.055 $Y=3.33
+ $X2=2.97 $Y2=3.33
r203 74 91 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.985 $Y=3.33
+ $X2=1.68 $Y2=3.33
r204 74 75 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.985 $Y=3.33
+ $X2=2.07 $Y2=3.33
r205 73 94 31.6417 $w=1.68e-07 $l=4.85e-07 $layer=LI1_cond $X=2.155 $Y=3.33
+ $X2=2.64 $Y2=3.33
r206 73 75 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.155 $Y=3.33
+ $X2=2.07 $Y2=3.33
r207 71 88 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=1.085 $Y=3.33
+ $X2=0.72 $Y2=3.33
r208 71 72 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.085 $Y=3.33
+ $X2=1.17 $Y2=3.33
r209 70 91 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=1.255 $Y=3.33
+ $X2=1.68 $Y2=3.33
r210 70 72 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.255 $Y=3.33
+ $X2=1.17 $Y2=3.33
r211 66 130 0.677923 $w=2.05e-07 $l=8.5e-08 $layer=LI1_cond $X=9.362 $Y=3.245
+ $X2=9.362 $Y2=3.33
r212 66 68 42.7406 $w=2.03e-07 $l=7.9e-07 $layer=LI1_cond $X=9.362 $Y=3.245
+ $X2=9.362 $Y2=2.455
r213 62 127 0.195364 $w=2.65e-07 $l=8.5e-08 $layer=LI1_cond $X=8.427 $Y=3.245
+ $X2=8.427 $Y2=3.33
r214 62 64 34.3558 $w=2.63e-07 $l=7.9e-07 $layer=LI1_cond $X=8.427 $Y=3.245
+ $X2=8.427 $Y2=2.455
r215 58 124 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.67 $Y=3.245
+ $X2=5.67 $Y2=3.33
r216 58 60 29.3349 $w=3.28e-07 $l=8.4e-07 $layer=LI1_cond $X=5.67 $Y=3.245
+ $X2=5.67 $Y2=2.405
r217 57 83 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.855 $Y=3.33
+ $X2=4.77 $Y2=3.33
r218 56 124 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.505 $Y=3.33
+ $X2=5.67 $Y2=3.33
r219 56 57 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=5.505 $Y=3.33
+ $X2=4.855 $Y2=3.33
r220 52 83 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.77 $Y=3.245
+ $X2=4.77 $Y2=3.33
r221 52 54 61.3262 $w=1.68e-07 $l=9.4e-07 $layer=LI1_cond $X=4.77 $Y=3.245
+ $X2=4.77 $Y2=2.305
r222 48 51 54.1497 $w=1.68e-07 $l=8.3e-07 $layer=LI1_cond $X=3.87 $Y=1.985
+ $X2=3.87 $Y2=2.815
r223 46 81 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.87 $Y=3.245
+ $X2=3.87 $Y2=3.33
r224 46 51 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=3.87 $Y=3.245
+ $X2=3.87 $Y2=2.815
r225 42 78 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.97 $Y=3.245
+ $X2=2.97 $Y2=3.33
r226 42 44 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=2.97 $Y=3.245
+ $X2=2.97 $Y2=2.455
r227 38 75 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.07 $Y=3.245
+ $X2=2.07 $Y2=3.33
r228 38 40 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=2.07 $Y=3.245
+ $X2=2.07 $Y2=2.455
r229 34 72 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.17 $Y=3.245
+ $X2=1.17 $Y2=3.33
r230 34 36 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=1.17 $Y=3.245
+ $X2=1.17 $Y2=2.455
r231 30 33 32.2684 $w=2.48e-07 $l=7e-07 $layer=LI1_cond $X=0.23 $Y=2.115
+ $X2=0.23 $Y2=2.815
r232 28 121 3.11948 $w=2.5e-07 $l=1.08305e-07 $layer=LI1_cond $X=0.23 $Y=3.245
+ $X2=0.177 $Y2=3.33
r233 28 33 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=0.23 $Y=3.245
+ $X2=0.23 $Y2=2.815
r234 9 68 300 $w=1.7e-07 $l=6.85912e-07 $layer=licon1_PDIFF $count=2 $X=9.21
+ $Y=1.84 $X2=9.36 $Y2=2.455
r235 8 64 300 $w=1.7e-07 $l=6.85912e-07 $layer=licon1_PDIFF $count=2 $X=8.31
+ $Y=1.84 $X2=8.46 $Y2=2.455
r236 7 60 300 $w=1.7e-07 $l=6.3559e-07 $layer=licon1_PDIFF $count=2 $X=5.52
+ $Y=1.84 $X2=5.67 $Y2=2.405
r237 6 54 300 $w=1.7e-07 $l=5.34766e-07 $layer=licon1_PDIFF $count=2 $X=4.62
+ $Y=1.84 $X2=4.77 $Y2=2.305
r238 5 51 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=3.72
+ $Y=1.84 $X2=3.87 $Y2=2.815
r239 5 48 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=3.72
+ $Y=1.84 $X2=3.87 $Y2=1.985
r240 4 44 300 $w=1.7e-07 $l=6.85912e-07 $layer=licon1_PDIFF $count=2 $X=2.82
+ $Y=1.84 $X2=2.97 $Y2=2.455
r241 3 40 300 $w=1.7e-07 $l=6.85912e-07 $layer=licon1_PDIFF $count=2 $X=1.92
+ $Y=1.84 $X2=2.07 $Y2=2.455
r242 2 36 300 $w=1.7e-07 $l=6.85912e-07 $layer=licon1_PDIFF $count=2 $X=1.02
+ $Y=1.84 $X2=1.17 $Y2=2.455
r243 1 33 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.27 $Y2=2.815
r244 1 30 400 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.27 $Y2=2.115
.ends

.subckt PM_SKY130_FD_SC_HS__O2BB2AI_4%Y 1 2 3 4 5 6 21 25 26 29 31 32 35 39 42
+ 43 44 47 51 53 55 56
c111 51 0 4.3658e-20 $X=5.715 $Y=1.045
c112 42 0 1.85729e-19 $X=5.63 $Y=1.8
c113 26 0 1.0348e-19 $X=4.485 $Y=1.885
r114 58 60 1.4104 $w=3.46e-07 $l=4e-08 $layer=LI1_cond $X=5.18 $Y=1.975 $X2=5.22
+ $Y2=1.975
r115 56 63 3.87861 $w=3.46e-07 $l=1.1e-07 $layer=LI1_cond $X=5.52 $Y=1.975
+ $X2=5.63 $Y2=1.975
r116 56 60 10.578 $w=3.46e-07 $l=3e-07 $layer=LI1_cond $X=5.52 $Y=1.975 $X2=5.22
+ $Y2=1.975
r117 48 53 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.825 $Y=2.035
+ $X2=6.66 $Y2=2.035
r118 47 55 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.395 $Y=2.035
+ $X2=7.56 $Y2=2.035
r119 47 48 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=7.395 $Y=2.035
+ $X2=6.825 $Y2=2.035
r120 44 63 6.15745 $w=3.46e-07 $l=1.11018e-07 $layer=LI1_cond $X=5.715 $Y=2.035
+ $X2=5.63 $Y2=1.975
r121 43 53 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.495 $Y=2.035
+ $X2=6.66 $Y2=2.035
r122 43 44 50.8877 $w=1.68e-07 $l=7.8e-07 $layer=LI1_cond $X=6.495 $Y=2.035
+ $X2=5.715 $Y2=2.035
r123 42 63 4.90539 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=5.63 $Y=1.8
+ $X2=5.63 $Y2=1.975
r124 41 51 3.64284 $w=2.55e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.63 $Y=1.13
+ $X2=5.715 $Y2=1.045
r125 41 42 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.63 $Y=1.13
+ $X2=5.63 $Y2=1.8
r126 37 51 3.64284 $w=2.55e-07 $l=8.5e-08 $layer=LI1_cond $X=5.715 $Y=0.96
+ $X2=5.715 $Y2=1.045
r127 37 39 3.38954 $w=3.38e-07 $l=1e-07 $layer=LI1_cond $X=5.715 $Y=0.96
+ $X2=5.715 $Y2=0.86
r128 33 58 2.64155 $w=2.5e-07 $l=1.75e-07 $layer=LI1_cond $X=5.18 $Y=2.15
+ $X2=5.18 $Y2=1.975
r129 33 35 11.5244 $w=2.48e-07 $l=2.5e-07 $layer=LI1_cond $X=5.18 $Y=2.15
+ $X2=5.18 $Y2=2.4
r130 31 51 2.83584 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=5.545 $Y=1.045
+ $X2=5.715 $Y2=1.045
r131 31 32 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=5.545 $Y=1.045
+ $X2=5.025 $Y2=1.045
r132 27 32 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.86 $Y=0.96
+ $X2=5.025 $Y2=1.045
r133 27 29 3.49225 $w=3.28e-07 $l=1e-07 $layer=LI1_cond $X=4.86 $Y=0.96 $X2=4.86
+ $Y2=0.86
r134 25 58 7.56786 $w=3.46e-07 $l=1.63936e-07 $layer=LI1_cond $X=5.055 $Y=1.885
+ $X2=5.18 $Y2=1.975
r135 25 26 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=5.055 $Y=1.885
+ $X2=4.485 $Y2=1.885
r136 21 23 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=4.32 $Y=1.985
+ $X2=4.32 $Y2=2.815
r137 19 26 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.32 $Y=1.97
+ $X2=4.485 $Y2=1.885
r138 19 21 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=4.32 $Y=1.97
+ $X2=4.32 $Y2=1.985
r139 6 55 300 $w=1.7e-07 $l=2.80134e-07 $layer=licon1_PDIFF $count=2 $X=7.41
+ $Y=1.84 $X2=7.56 $Y2=2.055
r140 5 53 300 $w=1.7e-07 $l=2.80134e-07 $layer=licon1_PDIFF $count=2 $X=6.51
+ $Y=1.84 $X2=6.66 $Y2=2.055
r141 4 60 600 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=5.07
+ $Y=1.84 $X2=5.22 $Y2=1.985
r142 4 35 300 $w=1.7e-07 $l=6.30555e-07 $layer=licon1_PDIFF $count=2 $X=5.07
+ $Y=1.84 $X2=5.22 $Y2=2.4
r143 3 23 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=4.17
+ $Y=1.84 $X2=4.32 $Y2=2.815
r144 3 21 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=4.17
+ $Y=1.84 $X2=4.32 $Y2=1.985
r145 2 39 182 $w=1.7e-07 $l=5.55608e-07 $layer=licon1_NDIFF $count=1 $X=5.58
+ $Y=0.37 $X2=5.72 $Y2=0.86
r146 1 29 182 $w=1.7e-07 $l=5.55608e-07 $layer=licon1_NDIFF $count=1 $X=4.72
+ $Y=0.37 $X2=4.86 $Y2=0.86
.ends

.subckt PM_SKY130_FD_SC_HS__O2BB2AI_4%A_1215_368# 1 2 3 4 5 18 20 21 24 26 32 36
+ 38 40 42 44 48
r66 40 50 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.81 $Y=2.12 $X2=9.81
+ $Y2=2.035
r67 40 42 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=9.81 $Y=2.12
+ $X2=9.81 $Y2=2.815
r68 39 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.075 $Y=2.035
+ $X2=8.91 $Y2=2.035
r69 38 50 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.645 $Y=2.035
+ $X2=9.81 $Y2=2.035
r70 38 39 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=9.645 $Y=2.035
+ $X2=9.075 $Y2=2.035
r71 34 48 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.91 $Y=2.12 $X2=8.91
+ $Y2=2.035
r72 34 36 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=8.91 $Y=2.12
+ $X2=8.91 $Y2=2.815
r73 33 46 3.71618 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=8.11 $Y=2.035 $X2=8.01
+ $Y2=2.035
r74 32 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.745 $Y=2.035
+ $X2=8.91 $Y2=2.035
r75 32 33 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=8.745 $Y=2.035
+ $X2=8.11 $Y2=2.035
r76 29 31 4.99091 $w=1.98e-07 $l=9e-08 $layer=LI1_cond $X=8.01 $Y=2.905 $X2=8.01
+ $Y2=2.815
r77 28 46 3.15876 $w=2e-07 $l=8.5e-08 $layer=LI1_cond $X=8.01 $Y=2.12 $X2=8.01
+ $Y2=2.035
r78 28 31 38.5409 $w=1.98e-07 $l=6.95e-07 $layer=LI1_cond $X=8.01 $Y=2.12
+ $X2=8.01 $Y2=2.815
r79 27 44 5.90115 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=7.21 $Y=2.99 $X2=7.11
+ $Y2=2.99
r80 26 29 6.87494 $w=1.7e-07 $l=1.36015e-07 $layer=LI1_cond $X=7.91 $Y=2.99
+ $X2=8.01 $Y2=2.905
r81 26 27 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=7.91 $Y=2.99 $X2=7.21
+ $Y2=2.99
r82 22 44 0.764409 $w=2e-07 $l=8.5e-08 $layer=LI1_cond $X=7.11 $Y=2.905 $X2=7.11
+ $Y2=2.99
r83 22 24 24.9545 $w=1.98e-07 $l=4.5e-07 $layer=LI1_cond $X=7.11 $Y=2.905
+ $X2=7.11 $Y2=2.455
r84 20 44 5.90115 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=7.01 $Y=2.99 $X2=7.11
+ $Y2=2.99
r85 20 21 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=7.01 $Y=2.99 $X2=6.31
+ $Y2=2.99
r86 16 21 7.24806 $w=1.7e-07 $l=1.70276e-07 $layer=LI1_cond $X=6.177 $Y=2.905
+ $X2=6.31 $Y2=2.99
r87 16 18 19.5698 $w=2.63e-07 $l=4.5e-07 $layer=LI1_cond $X=6.177 $Y=2.905
+ $X2=6.177 $Y2=2.455
r88 5 50 400 $w=1.7e-07 $l=2.59374e-07 $layer=licon1_PDIFF $count=1 $X=9.66
+ $Y=1.84 $X2=9.81 $Y2=2.035
r89 5 42 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=9.66
+ $Y=1.84 $X2=9.81 $Y2=2.815
r90 4 48 400 $w=1.7e-07 $l=2.59374e-07 $layer=licon1_PDIFF $count=1 $X=8.76
+ $Y=1.84 $X2=8.91 $Y2=2.035
r91 4 36 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=8.76
+ $Y=1.84 $X2=8.91 $Y2=2.815
r92 3 46 400 $w=1.7e-07 $l=3.4187e-07 $layer=licon1_PDIFF $count=1 $X=7.86
+ $Y=1.84 $X2=8.01 $Y2=2.115
r93 3 31 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=7.86
+ $Y=1.84 $X2=8.01 $Y2=2.815
r94 2 24 300 $w=1.7e-07 $l=6.85912e-07 $layer=licon1_PDIFF $count=2 $X=6.96
+ $Y=1.84 $X2=7.11 $Y2=2.455
r95 1 18 300 $w=1.7e-07 $l=6.79154e-07 $layer=licon1_PDIFF $count=2 $X=6.075
+ $Y=1.84 $X2=6.21 $Y2=2.455
.ends

.subckt PM_SKY130_FD_SC_HS__O2BB2AI_4%A_27_74# 1 2 3 4 5 18 20 21 24 26 32 33 36
+ 38 42 44 45
c68 42 0 1.50249e-19 $X=3.87 $Y=0.515
r69 40 42 4.14879 $w=2.48e-07 $l=9e-08 $layer=LI1_cond $X=3.91 $Y=0.425 $X2=3.91
+ $Y2=0.515
r70 39 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.105 $Y=0.34
+ $X2=2.94 $Y2=0.34
r71 38 40 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=3.785 $Y=0.34
+ $X2=3.91 $Y2=0.425
r72 38 39 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=3.785 $Y=0.34
+ $X2=3.105 $Y2=0.34
r73 34 45 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.94 $Y=0.425
+ $X2=2.94 $Y2=0.34
r74 34 36 5.93683 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=2.94 $Y=0.425
+ $X2=2.94 $Y2=0.595
r75 32 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.775 $Y=0.34
+ $X2=2.94 $Y2=0.34
r76 32 33 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=2.775 $Y=0.34
+ $X2=2.095 $Y2=0.34
r77 29 31 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=2.01 $Y=1.01
+ $X2=2.01 $Y2=0.515
r78 28 33 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.01 $Y=0.425
+ $X2=2.095 $Y2=0.34
r79 28 31 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=2.01 $Y=0.425 $X2=2.01
+ $Y2=0.515
r80 27 44 5.41628 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=1.235 $Y=1.095
+ $X2=1.145 $Y2=1.095
r81 26 29 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.925 $Y=1.095
+ $X2=2.01 $Y2=1.01
r82 26 27 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.925 $Y=1.095
+ $X2=1.235 $Y2=1.095
r83 22 44 1.13756 $w=1.8e-07 $l=8.5e-08 $layer=LI1_cond $X=1.145 $Y=1.01
+ $X2=1.145 $Y2=1.095
r84 22 24 30.5 $w=1.78e-07 $l=4.95e-07 $layer=LI1_cond $X=1.145 $Y=1.01
+ $X2=1.145 $Y2=0.515
r85 20 44 5.41628 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=1.055 $Y=1.095
+ $X2=1.145 $Y2=1.095
r86 20 21 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.055 $Y=1.095
+ $X2=0.365 $Y2=1.095
r87 16 21 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.24 $Y=1.01
+ $X2=0.365 $Y2=1.095
r88 16 18 22.8184 $w=2.48e-07 $l=4.95e-07 $layer=LI1_cond $X=0.24 $Y=1.01
+ $X2=0.24 $Y2=0.515
r89 5 42 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.73
+ $Y=0.37 $X2=3.87 $Y2=0.515
r90 4 36 182 $w=1.7e-07 $l=3.1285e-07 $layer=licon1_NDIFF $count=1 $X=2.73
+ $Y=0.37 $X2=2.94 $Y2=0.595
r91 3 31 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.87
+ $Y=0.37 $X2=2.01 $Y2=0.515
r92 2 24 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=1 $Y=0.37
+ $X2=1.145 $Y2=0.515
r93 1 18 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__O2BB2AI_4%VGND 1 2 3 4 5 6 21 25 27 31 35 39 43 45
+ 47 52 57 62 67 74 75 78 81 84 87 90 93
c129 31 0 1.9142e-19 $X=6.58 $Y=0.65
c130 25 0 1.9142e-19 $X=1.58 $Y=0.595
r131 93 94 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.36 $Y=0 $X2=9.36
+ $Y2=0
r132 90 91 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r133 87 88 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=0 $X2=7.44
+ $Y2=0
r134 84 85 1.69091 $w=1.7e-07 $l=9.35e-07 $layer=mcon $count=5 $X=6.48 $Y=0
+ $X2=6.48 $Y2=0
r135 81 82 1.69091 $w=1.7e-07 $l=9.35e-07 $layer=mcon $count=5 $X=1.68 $Y=0
+ $X2=1.68 $Y2=0
r136 78 79 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r137 75 94 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.84 $Y=0 $X2=9.36
+ $Y2=0
r138 74 75 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.84 $Y=0 $X2=9.84
+ $Y2=0
r139 72 93 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.535 $Y=0 $X2=9.37
+ $Y2=0
r140 72 74 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=9.535 $Y=0
+ $X2=9.84 $Y2=0
r141 71 94 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=0 $X2=9.36
+ $Y2=0
r142 71 91 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=0 $X2=8.4
+ $Y2=0
r143 70 71 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=0 $X2=8.88
+ $Y2=0
r144 68 90 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.605 $Y=0 $X2=8.44
+ $Y2=0
r145 68 70 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=8.605 $Y=0
+ $X2=8.88 $Y2=0
r146 67 93 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.205 $Y=0 $X2=9.37
+ $Y2=0
r147 67 70 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=9.205 $Y=0
+ $X2=8.88 $Y2=0
r148 66 91 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=0 $X2=8.4
+ $Y2=0
r149 66 88 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=0 $X2=7.44
+ $Y2=0
r150 65 66 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=0 $X2=7.92
+ $Y2=0
r151 63 87 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.675 $Y=0 $X2=7.51
+ $Y2=0
r152 63 65 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=7.675 $Y=0 $X2=7.92
+ $Y2=0
r153 62 90 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.275 $Y=0 $X2=8.44
+ $Y2=0
r154 62 65 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=8.275 $Y=0
+ $X2=7.92 $Y2=0
r155 61 88 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=0 $X2=7.44
+ $Y2=0
r156 61 85 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=0 $X2=6.48
+ $Y2=0
r157 60 61 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=0 $X2=6.96
+ $Y2=0
r158 58 84 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.745 $Y=0 $X2=6.58
+ $Y2=0
r159 58 60 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=6.745 $Y=0
+ $X2=6.96 $Y2=0
r160 57 87 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.345 $Y=0 $X2=7.51
+ $Y2=0
r161 57 60 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=7.345 $Y=0
+ $X2=6.96 $Y2=0
r162 56 82 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=1.68
+ $Y2=0
r163 56 79 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r164 55 56 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r165 53 78 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.875 $Y=0 $X2=0.71
+ $Y2=0
r166 53 55 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.875 $Y=0 $X2=1.2
+ $Y2=0
r167 52 81 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.415 $Y=0 $X2=1.58
+ $Y2=0
r168 52 55 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=1.415 $Y=0 $X2=1.2
+ $Y2=0
r169 50 79 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r170 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r171 47 78 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.545 $Y=0 $X2=0.71
+ $Y2=0
r172 47 49 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.545 $Y=0
+ $X2=0.24 $Y2=0
r173 45 85 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=5.04 $Y=0
+ $X2=6.48 $Y2=0
r174 45 82 0.936549 $w=4.9e-07 $l=3.36e-06 $layer=MET1_cond $X=5.04 $Y=0
+ $X2=1.68 $Y2=0
r175 41 93 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.37 $Y=0.085
+ $X2=9.37 $Y2=0
r176 41 43 19.7312 $w=3.28e-07 $l=5.65e-07 $layer=LI1_cond $X=9.37 $Y=0.085
+ $X2=9.37 $Y2=0.65
r177 37 90 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.44 $Y=0.085
+ $X2=8.44 $Y2=0
r178 37 39 19.7312 $w=3.28e-07 $l=5.65e-07 $layer=LI1_cond $X=8.44 $Y=0.085
+ $X2=8.44 $Y2=0.65
r179 33 87 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.51 $Y=0.085
+ $X2=7.51 $Y2=0
r180 33 35 19.7312 $w=3.28e-07 $l=5.65e-07 $layer=LI1_cond $X=7.51 $Y=0.085
+ $X2=7.51 $Y2=0.65
r181 29 84 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.58 $Y=0.085
+ $X2=6.58 $Y2=0
r182 29 31 19.7312 $w=3.28e-07 $l=5.65e-07 $layer=LI1_cond $X=6.58 $Y=0.085
+ $X2=6.58 $Y2=0.65
r183 28 81 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.745 $Y=0 $X2=1.58
+ $Y2=0
r184 27 84 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.415 $Y=0 $X2=6.58
+ $Y2=0
r185 27 28 304.674 $w=1.68e-07 $l=4.67e-06 $layer=LI1_cond $X=6.415 $Y=0
+ $X2=1.745 $Y2=0
r186 23 81 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.58 $Y=0.085
+ $X2=1.58 $Y2=0
r187 23 25 17.8105 $w=3.28e-07 $l=5.1e-07 $layer=LI1_cond $X=1.58 $Y=0.085
+ $X2=1.58 $Y2=0.595
r188 19 78 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.71 $Y=0.085
+ $X2=0.71 $Y2=0
r189 19 21 17.8105 $w=3.28e-07 $l=5.1e-07 $layer=LI1_cond $X=0.71 $Y=0.085
+ $X2=0.71 $Y2=0.595
r190 6 43 182 $w=1.7e-07 $l=3.70405e-07 $layer=licon1_NDIFF $count=1 $X=9.16
+ $Y=0.37 $X2=9.37 $Y2=0.65
r191 5 39 182 $w=1.7e-07 $l=3.42929e-07 $layer=licon1_NDIFF $count=1 $X=8.3
+ $Y=0.37 $X2=8.44 $Y2=0.65
r192 4 35 182 $w=1.7e-07 $l=3.42929e-07 $layer=licon1_NDIFF $count=1 $X=7.37
+ $Y=0.37 $X2=7.51 $Y2=0.65
r193 3 31 182 $w=1.7e-07 $l=3.42929e-07 $layer=licon1_NDIFF $count=1 $X=6.44
+ $Y=0.37 $X2=6.58 $Y2=0.65
r194 2 25 182 $w=1.7e-07 $l=2.86575e-07 $layer=licon1_NDIFF $count=1 $X=1.44
+ $Y=0.37 $X2=1.58 $Y2=0.595
r195 1 21 182 $w=1.7e-07 $l=2.86575e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.37 $X2=0.71 $Y2=0.595
.ends

.subckt PM_SKY130_FD_SC_HS__O2BB2AI_4%A_857_74# 1 2 3 4 5 6 7 24 26 27 30 32 38
+ 39 42 44 48 50 54 56 60 62 63 64 65
r107 58 60 22.8184 $w=2.48e-07 $l=4.95e-07 $layer=LI1_cond $X=9.84 $Y=1.01
+ $X2=9.84 $Y2=0.515
r108 57 65 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=9.035 $Y=1.095
+ $X2=8.91 $Y2=1.095
r109 56 58 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=9.715 $Y=1.095
+ $X2=9.84 $Y2=1.01
r110 56 57 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=9.715 $Y=1.095
+ $X2=9.035 $Y2=1.095
r111 52 65 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=8.91 $Y=1.01
+ $X2=8.91 $Y2=1.095
r112 52 54 22.8184 $w=2.48e-07 $l=4.95e-07 $layer=LI1_cond $X=8.91 $Y=1.01
+ $X2=8.91 $Y2=0.515
r113 51 64 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.095 $Y=1.095
+ $X2=7.97 $Y2=1.095
r114 50 65 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.785 $Y=1.095
+ $X2=8.91 $Y2=1.095
r115 50 51 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=8.785 $Y=1.095
+ $X2=8.095 $Y2=1.095
r116 46 64 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=7.97 $Y=1.01
+ $X2=7.97 $Y2=1.095
r117 46 48 22.8184 $w=2.48e-07 $l=4.95e-07 $layer=LI1_cond $X=7.97 $Y=1.01
+ $X2=7.97 $Y2=0.515
r118 45 63 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.165 $Y=1.095
+ $X2=7.04 $Y2=1.095
r119 44 64 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.845 $Y=1.095
+ $X2=7.97 $Y2=1.095
r120 44 45 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=7.845 $Y=1.095
+ $X2=7.165 $Y2=1.095
r121 40 63 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=7.04 $Y=1.01
+ $X2=7.04 $Y2=1.095
r122 40 42 22.8184 $w=2.48e-07 $l=4.95e-07 $layer=LI1_cond $X=7.04 $Y=1.01
+ $X2=7.04 $Y2=0.515
r123 38 63 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.915 $Y=1.095
+ $X2=7.04 $Y2=1.095
r124 38 39 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=6.915 $Y=1.095
+ $X2=6.235 $Y2=1.095
r125 35 39 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.15 $Y=1.01
+ $X2=6.235 $Y2=1.095
r126 35 37 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=6.15 $Y=1.01
+ $X2=6.15 $Y2=0.515
r127 34 37 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=6.15 $Y=0.425
+ $X2=6.15 $Y2=0.515
r128 33 62 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.375 $Y=0.34
+ $X2=5.29 $Y2=0.34
r129 32 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.065 $Y=0.34
+ $X2=6.15 $Y2=0.425
r130 32 33 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=6.065 $Y=0.34
+ $X2=5.375 $Y2=0.34
r131 28 62 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.29 $Y=0.425
+ $X2=5.29 $Y2=0.34
r132 28 30 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=5.29 $Y=0.425
+ $X2=5.29 $Y2=0.57
r133 26 62 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.205 $Y=0.34
+ $X2=5.29 $Y2=0.34
r134 26 27 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=5.205 $Y=0.34
+ $X2=4.515 $Y2=0.34
r135 22 27 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=4.39 $Y=0.425
+ $X2=4.515 $Y2=0.34
r136 22 24 4.14879 $w=2.48e-07 $l=9e-08 $layer=LI1_cond $X=4.39 $Y=0.425
+ $X2=4.39 $Y2=0.515
r137 7 60 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=9.66
+ $Y=0.37 $X2=9.8 $Y2=0.515
r138 6 54 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=8.73
+ $Y=0.37 $X2=8.87 $Y2=0.515
r139 5 48 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=7.87
+ $Y=0.37 $X2=8.01 $Y2=0.515
r140 4 42 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=6.94
+ $Y=0.37 $X2=7.08 $Y2=0.515
r141 3 37 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=6.01
+ $Y=0.37 $X2=6.15 $Y2=0.515
r142 2 30 182 $w=1.7e-07 $l=2.60768e-07 $layer=licon1_NDIFF $count=1 $X=5.15
+ $Y=0.37 $X2=5.29 $Y2=0.57
r143 1 24 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=4.285
+ $Y=0.37 $X2=4.43 $Y2=0.515
.ends

