* File: sky130_fd_sc_hs__sdfrtp_1.spice
* Created: Tue Sep  1 20:22:38 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hs__sdfrtp_1.pex.spice"
.subckt sky130_fd_sc_hs__sdfrtp_1  VNB VPB SCE D SCD RESET_B CLK VPWR Q VGND
* 
* VGND	VGND
* Q	Q
* VPWR	VPWR
* CLK	CLK
* RESET_B	RESET_B
* SCD	SCD
* D	D
* SCE	SCE
* VPB	VPB
* VNB	VNB
MM1037 N_VGND_M1037_d N_SCE_M1037_g N_A_27_88#_M1037_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.1197 AS=0.1197 PD=1.41 PS=1.41 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1012 noxref_25 N_A_27_88#_M1012_g N_noxref_24_M1012_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.0504 AS=0.1197 PD=0.66 PS=1.41 NRD=18.564 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75002.4 A=0.063 P=1.14 MULT=1
MM1013 N_A_300_464#_M1013_d N_D_M1013_g noxref_25 VNB NLOWVT L=0.15 W=0.42
+ AD=0.13125 AS=0.0504 PD=1.045 PS=0.66 NRD=98.568 NRS=18.564 M=1 R=2.8
+ SA=75000.6 SB=75002 A=0.063 P=1.14 MULT=1
MM1030 noxref_26 N_SCE_M1030_g N_A_300_464#_M1013_d VNB NLOWVT L=0.15 W=0.42
+ AD=0.0504 AS=0.13125 PD=0.66 PS=1.045 NRD=18.564 NRS=0 M=1 R=2.8 SA=75001.4
+ SB=75001.2 A=0.063 P=1.14 MULT=1
MM1021 N_noxref_24_M1021_d N_SCD_M1021_g noxref_26 VNB NLOWVT L=0.15 W=0.42
+ AD=0.09765 AS=0.0504 PD=0.885 PS=0.66 NRD=25.704 NRS=18.564 M=1 R=2.8
+ SA=75001.8 SB=75000.8 A=0.063 P=1.14 MULT=1
MM1016 N_VGND_M1016_d N_RESET_B_M1016_g N_noxref_24_M1021_d VNB NLOWVT L=0.15
+ W=0.42 AD=0.1197 AS=0.09765 PD=1.41 PS=0.885 NRD=0 NRS=27.132 M=1 R=2.8
+ SA=75002.4 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1008 N_VGND_M1008_d N_CLK_M1008_g N_A_855_368#_M1008_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.10545 AS=0.2109 PD=1.025 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75000.6 A=0.111 P=1.78 MULT=1
MM1003 N_A_1034_368#_M1003_d N_A_855_368#_M1003_g N_VGND_M1008_d VNB NLOWVT
+ L=0.15 W=0.74 AD=0.2109 AS=0.10545 PD=2.05 PS=1.025 NRD=0 NRS=0.804 M=1
+ R=4.93333 SA=75000.6 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1009 N_A_1233_118#_M1009_d N_A_855_368#_M1009_g N_A_300_464#_M1009_s VNB
+ NLOWVT L=0.15 W=0.42 AD=0.0588 AS=0.1197 PD=0.7 PS=1.41 NRD=0 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75003.9 A=0.063 P=1.14 MULT=1
MM1000 A_1319_118# N_A_1034_368#_M1000_g N_A_1233_118#_M1009_d VNB NLOWVT L=0.15
+ W=0.42 AD=0.0504 AS=0.0588 PD=0.66 PS=0.7 NRD=18.564 NRS=0 M=1 R=2.8
+ SA=75000.6 SB=75003.4 A=0.063 P=1.14 MULT=1
MM1027 A_1397_118# N_A_1367_92#_M1027_g A_1319_118# VNB NLOWVT L=0.15 W=0.42
+ AD=0.0504 AS=0.0504 PD=0.66 PS=0.66 NRD=18.564 NRS=18.564 M=1 R=2.8 SA=75001
+ SB=75003 A=0.063 P=1.14 MULT=1
MM1019 N_VGND_M1019_d N_RESET_B_M1019_g A_1397_118# VNB NLOWVT L=0.15 W=0.42
+ AD=0.210555 AS=0.0504 PD=1.26792 PS=0.66 NRD=127.512 NRS=18.564 M=1 R=2.8
+ SA=75001.4 SB=75002.6 A=0.063 P=1.14 MULT=1
MM1033 N_A_1367_92#_M1033_d N_A_1233_118#_M1033_g N_VGND_M1019_d VNB NLOWVT
+ L=0.15 W=0.64 AD=0.0896 AS=0.320845 PD=0.92 PS=1.93208 NRD=0 NRS=83.676 M=1
+ R=4.26667 SA=75001.7 SB=75002.1 A=0.096 P=1.58 MULT=1
MM1010 N_A_1745_74#_M1010_d N_A_1034_368#_M1010_g N_A_1367_92#_M1033_d VNB
+ NLOWVT L=0.15 W=0.64 AD=0.282989 AS=0.0896 PD=1.96226 PS=0.92 NRD=132.18 NRS=0
+ M=1 R=4.26667 SA=75002.2 SB=75001.7 A=0.096 P=1.58 MULT=1
MM1007 A_1972_74# N_A_855_368#_M1007_g N_A_1745_74#_M1010_d VNB NLOWVT L=0.15
+ W=0.42 AD=0.0441 AS=0.185711 PD=0.63 PS=1.28774 NRD=14.28 NRS=0 M=1 R=2.8
+ SA=75003 SB=75001.4 A=0.063 P=1.14 MULT=1
MM1005 N_VGND_M1005_d N_A_1997_272#_M1005_g A_1972_74# VNB NLOWVT L=0.15 W=0.42
+ AD=0.06405 AS=0.0441 PD=0.725 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75003.4
+ SB=75001 A=0.063 P=1.14 MULT=1
MM1038 A_2135_74# N_RESET_B_M1038_g N_VGND_M1005_d VNB NLOWVT L=0.15 W=0.42
+ AD=0.0441 AS=0.06405 PD=0.63 PS=0.725 NRD=14.28 NRS=7.14 M=1 R=2.8 SA=75003.8
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1028 N_A_1997_272#_M1028_d N_A_1745_74#_M1028_g A_2135_74# VNB NLOWVT L=0.15
+ W=0.42 AD=0.1197 AS=0.0441 PD=1.41 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8
+ SA=75004.2 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1031 N_A_2399_424#_M1031_d N_A_1745_74#_M1031_g N_VGND_M1031_s VNB NLOWVT
+ L=0.15 W=0.55 AD=0.15675 AS=0.1595 PD=1.67 PS=1.68 NRD=0 NRS=1.08 M=1
+ R=3.66667 SA=75000.2 SB=75000.2 A=0.0825 P=1.4 MULT=1
MM1011 N_Q_M1011_d N_A_2399_424#_M1011_g N_VGND_M1011_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.2109 PD=2.05 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1023 N_VPWR_M1023_d N_SCE_M1023_g N_A_27_88#_M1023_s VPB PSHORT L=0.15 W=0.64
+ AD=0.112 AS=0.1888 PD=0.99 PS=1.87 NRD=18.4589 NRS=3.0732 M=1 R=4.26667
+ SA=75000.2 SB=75003.3 A=0.096 P=1.58 MULT=1
MM1020 A_216_464# N_SCE_M1020_g N_VPWR_M1023_d VPB PSHORT L=0.15 W=0.64
+ AD=0.0864 AS=0.112 PD=0.91 PS=0.99 NRD=24.625 NRS=3.0732 M=1 R=4.26667
+ SA=75000.7 SB=75002.8 A=0.096 P=1.58 MULT=1
MM1036 N_A_300_464#_M1036_d N_D_M1036_g A_216_464# VPB PSHORT L=0.15 W=0.64
+ AD=0.3328 AS=0.0864 PD=1.68 PS=0.91 NRD=3.0732 NRS=24.625 M=1 R=4.26667
+ SA=75001.1 SB=75002.4 A=0.096 P=1.58 MULT=1
MM1024 A_538_464# N_A_27_88#_M1024_g N_A_300_464#_M1036_d VPB PSHORT L=0.15
+ W=0.64 AD=0.0864 AS=0.3328 PD=0.91 PS=1.68 NRD=24.625 NRS=3.0732 M=1 R=4.26667
+ SA=75002.3 SB=75001.2 A=0.096 P=1.58 MULT=1
MM1006 N_VPWR_M1006_d N_SCD_M1006_g A_538_464# VPB PSHORT L=0.15 W=0.64
+ AD=0.1344 AS=0.0864 PD=1.06 PS=0.91 NRD=3.0732 NRS=24.625 M=1 R=4.26667
+ SA=75002.8 SB=75000.8 A=0.096 P=1.58 MULT=1
MM1039 N_A_300_464#_M1039_d N_RESET_B_M1039_g N_VPWR_M1006_d VPB PSHORT L=0.15
+ W=0.64 AD=0.1888 AS=0.1344 PD=1.87 PS=1.06 NRD=3.0732 NRS=40.0107 M=1
+ R=4.26667 SA=75003.3 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1022 N_VPWR_M1022_d N_CLK_M1022_g N_A_855_368#_M1022_s VPB PSHORT L=0.15
+ W=1.12 AD=0.168 AS=0.3304 PD=1.42 PS=2.83 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1029 N_A_1034_368#_M1029_d N_A_855_368#_M1029_g N_VPWR_M1022_d VPB PSHORT
+ L=0.15 W=1.12 AD=0.3304 AS=0.168 PD=2.83 PS=1.42 NRD=1.7533 NRS=1.7533 M=1
+ R=7.46667 SA=75000.7 SB=75000.2 A=0.168 P=2.54 MULT=1
MM1026 N_A_1233_118#_M1026_d N_A_1034_368#_M1026_g N_A_300_464#_M1026_s VPB
+ PSHORT L=0.15 W=0.42 AD=0.0763 AS=0.1239 PD=0.795 PS=1.43 NRD=30.4759
+ NRS=4.6886 M=1 R=2.8 SA=75000.2 SB=75001.7 A=0.063 P=1.14 MULT=1
MM1032 A_1343_461# N_A_855_368#_M1032_g N_A_1233_118#_M1026_d VPB PSHORT L=0.15
+ W=0.42 AD=0.0567 AS=0.0763 PD=0.69 PS=0.795 NRD=37.5088 NRS=4.6886 M=1 R=2.8
+ SA=75000.7 SB=75001.3 A=0.063 P=1.14 MULT=1
MM1002 N_VPWR_M1002_d N_A_1367_92#_M1002_g A_1343_461# VPB PSHORT L=0.15 W=0.42
+ AD=0.135887 AS=0.0567 PD=1.14 PS=0.69 NRD=125.942 NRS=37.5088 M=1 R=2.8
+ SA=75001.1 SB=75000.8 A=0.063 P=1.14 MULT=1
MM1034 N_A_1233_118#_M1034_d N_RESET_B_M1034_g N_VPWR_M1002_d VPB PSHORT L=0.15
+ W=0.42 AD=0.1239 AS=0.135887 PD=1.43 PS=1.14 NRD=4.6886 NRS=125.942 M=1 R=2.8
+ SA=75001.7 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1001 N_A_1367_92#_M1001_d N_A_1233_118#_M1001_g N_VPWR_M1001_s VPB PSHORT
+ L=0.15 W=1 AD=0.15 AS=0.295 PD=1.3 PS=2.59 NRD=1.9503 NRS=1.9503 M=1 R=6.66667
+ SA=75000.2 SB=75001.2 A=0.15 P=2.3 MULT=1
MM1004 N_A_1745_74#_M1004_d N_A_855_368#_M1004_g N_A_1367_92#_M1001_d VPB PSHORT
+ L=0.15 W=1 AD=0.311954 AS=0.15 PD=2.56338 PS=1.3 NRD=40.3653 NRS=1.9503 M=1
+ R=6.66667 SA=75000.7 SB=75000.7 A=0.15 P=2.3 MULT=1
MM1025 A_1993_508# N_A_1034_368#_M1025_g N_A_1745_74#_M1004_d VPB PSHORT L=0.15
+ W=0.42 AD=0.0567 AS=0.131021 PD=0.69 PS=1.07662 NRD=37.5088 NRS=53.9386 M=1
+ R=2.8 SA=75000.9 SB=75002.2 A=0.063 P=1.14 MULT=1
MM1014 N_VPWR_M1014_d N_A_1997_272#_M1014_g A_1993_508# VPB PSHORT L=0.15 W=0.42
+ AD=0.08925 AS=0.0567 PD=0.845 PS=0.69 NRD=21.0987 NRS=37.5088 M=1 R=2.8
+ SA=75001.3 SB=75001.8 A=0.063 P=1.14 MULT=1
MM1015 N_A_1997_272#_M1015_d N_RESET_B_M1015_g N_VPWR_M1014_d VPB PSHORT L=0.15
+ W=0.42 AD=0.063 AS=0.08925 PD=0.72 PS=0.845 NRD=4.6886 NRS=46.886 M=1 R=2.8
+ SA=75001.9 SB=75001.3 A=0.063 P=1.14 MULT=1
MM1018 N_VPWR_M1018_d N_A_1745_74#_M1018_g N_A_1997_272#_M1015_d VPB PSHORT
+ L=0.15 W=0.42 AD=0.1092 AS=0.063 PD=0.85 PS=0.72 NRD=44.5417 NRS=4.6886 M=1
+ R=2.8 SA=75002.3 SB=75000.8 A=0.063 P=1.14 MULT=1
MM1017 N_A_2399_424#_M1017_d N_A_1745_74#_M1017_g N_VPWR_M1018_d VPB PSHORT
+ L=0.15 W=0.84 AD=0.2478 AS=0.2184 PD=2.27 PS=1.7 NRD=2.3443 NRS=14.0658 M=1
+ R=5.6 SA=75001.6 SB=75000.2 A=0.126 P=1.98 MULT=1
MM1035 N_Q_M1035_d N_A_2399_424#_M1035_g N_VPWR_M1035_s VPB PSHORT L=0.15 W=1.12
+ AD=0.3304 AS=0.3304 PD=2.83 PS=2.83 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75000.2 A=0.168 P=2.54 MULT=1
DX40_noxref VNB VPB NWDIODE A=25.8648 P=31.57
c_152 VNB 0 1.07934e-19 $X=0 $Y=0
c_2129 A_1343_461# 0 1.84284e-19 $X=6.715 $Y=2.305
c_2131 A_1993_508# 0 1.05093e-19 $X=9.965 $Y=2.54
*
.include "sky130_fd_sc_hs__sdfrtp_1.pxi.spice"
*
.ends
*
*
