* File: sky130_fd_sc_hs__o211ai_1.spice
* Created: Tue Sep  1 20:13:54 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hs__o211ai_1.pex.spice"
.subckt sky130_fd_sc_hs__o211ai_1  VNB VPB A1 A2 B1 C1 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* C1	C1
* B1	B1
* A2	A2
* A1	A1
* VPB	VPB
* VNB	VNB
MM1006 N_VGND_M1006_d N_A1_M1006_g N_A_31_74#_M1006_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1295 AS=0.2109 PD=1.09 PS=2.05 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75002.1 A=0.111 P=1.78 MULT=1
MM1001 N_A_31_74#_M1001_d N_A2_M1001_g N_VGND_M1006_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.11655 AS=0.1295 PD=1.055 PS=1.09 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.7
+ SB=75001.6 A=0.111 P=1.78 MULT=1
MM1002 A_311_74# N_B1_M1002_g N_A_31_74#_M1001_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.1554 AS=0.11655 PD=1.16 PS=1.055 NRD=25.128 NRS=5.664 M=1 R=4.93333
+ SA=75001.2 SB=75001.1 A=0.111 P=1.78 MULT=1
MM1007 N_Y_M1007_d N_C1_M1007_g A_311_74# VNB NLOWVT L=0.15 W=0.74 AD=0.4588
+ AS=0.1554 PD=2.72 PS=1.16 NRD=0 NRS=25.128 M=1 R=4.93333 SA=75001.7 SB=75000.5
+ A=0.111 P=1.78 MULT=1
MM1005 A_116_368# N_A1_M1005_g N_VPWR_M1005_s VPB PSHORT L=0.15 W=1.12 AD=0.1512
+ AS=0.3304 PD=1.39 PS=2.83 NRD=14.0658 NRS=1.7533 M=1 R=7.46667 SA=75000.2
+ SB=75001.9 A=0.168 P=2.54 MULT=1
MM1000 N_Y_M1000_d N_A2_M1000_g A_116_368# VPB PSHORT L=0.15 W=1.12 AD=0.3192
+ AS=0.1512 PD=1.69 PS=1.39 NRD=26.3783 NRS=14.0658 M=1 R=7.46667 SA=75000.6
+ SB=75001.4 A=0.168 P=2.54 MULT=1
MM1004 N_VPWR_M1004_d N_B1_M1004_g N_Y_M1000_d VPB PSHORT L=0.15 W=1.12 AD=0.196
+ AS=0.3192 PD=1.47 PS=1.69 NRD=1.7533 NRS=24.6053 M=1 R=7.46667 SA=75001.4
+ SB=75000.7 A=0.168 P=2.54 MULT=1
MM1003 N_Y_M1003_d N_C1_M1003_g N_VPWR_M1004_d VPB PSHORT L=0.15 W=1.12
+ AD=0.3304 AS=0.196 PD=2.83 PS=1.47 NRD=1.7533 NRS=10.5395 M=1 R=7.46667
+ SA=75001.9 SB=75000.2 A=0.168 P=2.54 MULT=1
DX8_noxref VNB VPB NWDIODE A=6.0636 P=10.24
*
.include "sky130_fd_sc_hs__o211ai_1.pxi.spice"
*
.ends
*
*
