* File: sky130_fd_sc_hs__dlclkp_1.spice
* Created: Tue Sep  1 20:01:21 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hs__dlclkp_1.pex.spice"
.subckt sky130_fd_sc_hs__dlclkp_1  VNB VPB GATE CLK VPWR GCLK VGND
* 
* VGND	VGND
* GCLK	GCLK
* VPWR	VPWR
* CLK	CLK
* GATE	GATE
* VPB	VPB
* VNB	VNB
MM1017 N_VGND_M1017_d N_A_83_260#_M1017_g N_A_27_74#_M1017_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.235647 AS=0.2109 PD=1.51754 PS=2.05 NRD=13.776 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75002.2 A=0.111 P=1.78 MULT=1
MM1018 A_267_80# N_GATE_M1018_g N_VGND_M1017_d VNB NLOWVT L=0.15 W=0.64
+ AD=0.0768 AS=0.203803 PD=0.88 PS=1.31246 NRD=12.18 NRS=48.744 M=1 R=4.26667
+ SA=75001 SB=75001.7 A=0.096 P=1.58 MULT=1
MM1019 N_A_83_260#_M1019_d N_A_315_54#_M1019_g A_267_80# VNB NLOWVT L=0.15
+ W=0.64 AD=0.162536 AS=0.0768 PD=1.38868 PS=0.88 NRD=21.552 NRS=12.18 M=1
+ R=4.26667 SA=75001.4 SB=75001.3 A=0.096 P=1.58 MULT=1
MM1002 A_477_124# N_A_309_338#_M1002_g N_A_83_260#_M1019_d VNB NLOWVT L=0.15
+ W=0.42 AD=0.0504 AS=0.106664 PD=0.66 PS=0.911321 NRD=18.564 NRS=32.856 M=1
+ R=2.8 SA=75002 SB=75001.2 A=0.063 P=1.14 MULT=1
MM1016 N_VGND_M1016_d N_A_27_74#_M1016_g A_477_124# VNB NLOWVT L=0.15 W=0.42
+ AD=0.102746 AS=0.0504 PD=0.89069 PS=0.66 NRD=28.56 NRS=18.564 M=1 R=2.8
+ SA=75002.4 SB=75000.8 A=0.063 P=1.14 MULT=1
MM1004 N_A_309_338#_M1004_d N_A_315_54#_M1004_g N_VGND_M1016_d VNB NLOWVT L=0.15
+ W=0.74 AD=0.2109 AS=0.181029 PD=2.05 PS=1.56931 NRD=0 NRS=17.016 M=1 R=4.93333
+ SA=75001.8 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1003 N_VGND_M1003_d N_CLK_M1003_g N_A_315_54#_M1003_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.13883 AS=0.2183 PD=1.17971 PS=2.07 NRD=0 NRS=0.804 M=1 R=4.93333
+ SA=75000.2 SB=75001 A=0.111 P=1.78 MULT=1
MM1011 A_984_125# N_CLK_M1011_g N_VGND_M1003_d VNB NLOWVT L=0.15 W=0.64
+ AD=0.0768 AS=0.12007 PD=0.88 PS=1.02029 NRD=12.18 NRS=14.988 M=1 R=4.26667
+ SA=75000.7 SB=75000.6 A=0.096 P=1.58 MULT=1
MM1006 N_A_987_393#_M1006_d N_A_27_74#_M1006_g A_984_125# VNB NLOWVT L=0.15
+ W=0.64 AD=0.1824 AS=0.0768 PD=1.85 PS=0.88 NRD=0 NRS=12.18 M=1 R=4.26667
+ SA=75001.1 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1012 N_GCLK_M1012_d N_A_987_393#_M1012_g N_VGND_M1012_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.2109 AS=0.2109 PD=2.05 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1008 N_VPWR_M1008_d N_A_83_260#_M1008_g N_A_27_74#_M1008_s VPB PSHORT L=0.15
+ W=1.12 AD=0.312649 AS=0.3304 PD=1.77509 PS=2.83 NRD=10.5395 NRS=1.7533 M=1
+ R=7.46667 SA=75000.2 SB=75001.8 A=0.168 P=2.54 MULT=1
MM1005 A_258_392# N_GATE_M1005_g N_VPWR_M1008_d VPB PSHORT L=0.15 W=1 AD=0.135
+ AS=0.279151 PD=1.27 PS=1.58491 NRD=15.7403 NRS=43.3203 M=1 R=6.66667
+ SA=75000.9 SB=75001.3 A=0.15 P=2.3 MULT=1
MM1013 N_A_83_260#_M1013_d N_A_309_338#_M1013_g A_258_392# VPB PSHORT L=0.15 W=1
+ AD=0.273873 AS=0.135 PD=2.19718 PS=1.27 NRD=27.5603 NRS=15.7403 M=1 R=6.66667
+ SA=75001.3 SB=75000.8 A=0.15 P=2.3 MULT=1
MM1009 A_484_508# N_A_315_54#_M1009_g N_A_83_260#_M1013_d VPB PSHORT L=0.15
+ W=0.42 AD=0.0567 AS=0.115027 PD=0.69 PS=0.922817 NRD=37.5088 NRS=65.6601 M=1
+ R=2.8 SA=75002.1 SB=75001 A=0.063 P=1.14 MULT=1
MM1014 N_VPWR_M1014_d N_A_27_74#_M1014_g A_484_508# VPB PSHORT L=0.15 W=0.42
+ AD=0.0999833 AS=0.0567 PD=0.91 PS=0.69 NRD=9.3772 NRS=37.5088 M=1 R=2.8
+ SA=75002.5 SB=75000.6 A=0.063 P=1.14 MULT=1
MM1000 N_A_309_338#_M1000_d N_A_315_54#_M1000_g N_VPWR_M1014_d VPB PSHORT L=0.15
+ W=0.84 AD=0.2478 AS=0.199967 PD=2.27 PS=1.82 NRD=2.3443 NRS=23.443 M=1 R=5.6
+ SA=75001.2 SB=75000.2 A=0.126 P=1.98 MULT=1
MM1010 N_VPWR_M1010_d N_CLK_M1010_g N_A_315_54#_M1010_s VPB PSHORT L=0.15 W=0.84
+ AD=0.1638 AS=0.2478 PD=1.23 PS=2.27 NRD=14.0658 NRS=2.3443 M=1 R=5.6
+ SA=75000.2 SB=75002 A=0.126 P=1.98 MULT=1
MM1001 N_A_987_393#_M1001_d N_CLK_M1001_g N_VPWR_M1010_d VPB PSHORT L=0.15
+ W=0.84 AD=0.1302 AS=0.1638 PD=1.15 PS=1.23 NRD=4.6886 NRS=11.7215 M=1 R=5.6
+ SA=75000.8 SB=75001.5 A=0.126 P=1.98 MULT=1
MM1015 N_VPWR_M1015_d N_A_27_74#_M1015_g N_A_987_393#_M1001_d VPB PSHORT L=0.15
+ W=0.84 AD=0.2844 AS=0.1302 PD=1.53857 PS=1.15 NRD=78.9379 NRS=2.3443 M=1 R=5.6
+ SA=75001.2 SB=75001 A=0.126 P=1.98 MULT=1
MM1007 N_GCLK_M1007_d N_A_987_393#_M1007_g N_VPWR_M1015_d VPB PSHORT L=0.15
+ W=1.12 AD=0.3304 AS=0.3792 PD=2.83 PS=2.05143 NRD=1.7533 NRS=10.5395 M=1
+ R=7.46667 SA=75001.6 SB=75000.2 A=0.168 P=2.54 MULT=1
DX20_noxref VNB VPB NWDIODE A=12.9104 P=18.17
c_120 VPB 0 1.78419e-19 $X=0 $Y=3.085
*
.include "sky130_fd_sc_hs__dlclkp_1.pxi.spice"
*
.ends
*
*
