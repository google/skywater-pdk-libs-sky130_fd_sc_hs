* File: sky130_fd_sc_hs__nand2_4.spice
* Created: Thu Aug 27 20:50:13 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hs__nand2_4.pex.spice"
.subckt sky130_fd_sc_hs__nand2_4  VNB VPB B A VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A	A
* B	B
* VPB	VPB
* VNB	VNB
MM1006 N_VGND_M1006_d N_B_M1006_g N_A_27_74#_M1006_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.2109 PD=1.02 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75003.5 A=0.111 P=1.78 MULT=1
MM1009 N_VGND_M1006_d N_B_M1009_g N_A_27_74#_M1009_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.6
+ SB=75003.1 A=0.111 P=1.78 MULT=1
MM1010 N_VGND_M1010_d N_B_M1010_g N_A_27_74#_M1009_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.1
+ SB=75002.7 A=0.111 P=1.78 MULT=1
MM1011 N_VGND_M1010_d N_B_M1011_g N_A_27_74#_M1011_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1184 PD=1.02 PS=1.06 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.5
+ SB=75002.2 A=0.111 P=1.78 MULT=1
MM1002 N_Y_M1002_d N_A_M1002_g N_A_27_74#_M1011_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1147 AS=0.1184 PD=1.05 PS=1.06 NRD=4.86 NRS=6.48 M=1 R=4.93333 SA=75002
+ SB=75001.8 A=0.111 P=1.78 MULT=1
MM1004 N_Y_M1002_d N_A_M1004_g N_A_27_74#_M1004_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1147 AS=0.1295 PD=1.05 PS=1.09 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75002.4
+ SB=75001.3 A=0.111 P=1.78 MULT=1
MM1007 N_Y_M1007_d N_A_M1007_g N_A_27_74#_M1004_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.15355 AS=0.1295 PD=1.155 PS=1.09 NRD=14.592 NRS=0 M=1 R=4.93333
+ SA=75002.9 SB=75000.8 A=0.111 P=1.78 MULT=1
MM1008 N_Y_M1007_d N_A_M1008_g N_A_27_74#_M1008_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.15355 AS=0.2442 PD=1.155 PS=2.14 NRD=7.296 NRS=7.296 M=1 R=4.93333
+ SA=75003.5 SB=75000.3 A=0.111 P=1.78 MULT=1
MM1001 N_VPWR_M1001_d N_B_M1001_g N_Y_M1001_s VPB PSHORT L=0.15 W=1.12 AD=0.336
+ AS=0.6216 PD=2.84 PS=2.23 NRD=2.6201 NRS=1.7533 M=1 R=7.46667 SA=75000.2
+ SB=75003.5 A=0.168 P=2.54 MULT=1
MM1005 N_VPWR_M1005_d N_B_M1005_g N_Y_M1001_s VPB PSHORT L=0.15 W=1.12 AD=0.196
+ AS=0.6216 PD=1.47 PS=2.23 NRD=1.7533 NRS=1.7533 M=1 R=7.46667 SA=75001.5
+ SB=75002.3 A=0.168 P=2.54 MULT=1
MM1000 N_Y_M1000_d N_A_M1000_g N_VPWR_M1005_d VPB PSHORT L=0.15 W=1.12 AD=0.7532
+ AS=0.196 PD=2.465 PS=1.47 NRD=1.7533 NRS=10.5395 M=1 R=7.46667 SA=75002
+ SB=75001.8 A=0.168 P=2.54 MULT=1
MM1003 N_Y_M1000_d N_A_M1003_g N_VPWR_M1003_s VPB PSHORT L=0.15 W=1.12 AD=0.7532
+ AS=0.3864 PD=2.465 PS=2.93 NRD=1.7533 NRS=10.5395 M=1 R=7.46667 SA=75003.5
+ SB=75000.3 A=0.168 P=2.54 MULT=1
DX12_noxref VNB VPB NWDIODE A=8.742 P=13.12
*
.include "sky130_fd_sc_hs__nand2_4.pxi.spice"
*
.ends
*
*
