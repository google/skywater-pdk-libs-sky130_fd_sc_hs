* File: sky130_fd_sc_hs__nand3_2.pxi.spice
* Created: Tue Sep  1 20:09:18 2020
* 
x_PM_SKY130_FD_SC_HS__NAND3_2%C N_C_c_58_n N_C_M1000_g N_C_c_62_n N_C_M1004_g
+ N_C_c_59_n N_C_M1010_g N_C_c_63_n N_C_M1006_g C N_C_c_60_n N_C_c_61_n
+ PM_SKY130_FD_SC_HS__NAND3_2%C
x_PM_SKY130_FD_SC_HS__NAND3_2%B N_B_M1002_g N_B_c_110_n N_B_M1005_g N_B_c_111_n
+ N_B_M1009_g N_B_M1008_g N_B_c_129_p N_B_c_162_p N_B_c_113_n N_B_c_114_n B
+ N_B_c_115_n B PM_SKY130_FD_SC_HS__NAND3_2%B
x_PM_SKY130_FD_SC_HS__NAND3_2%A N_A_M1001_g N_A_c_204_n N_A_M1003_g N_A_M1011_g
+ N_A_c_205_n N_A_M1007_g A N_A_c_206_n N_A_c_203_n
+ PM_SKY130_FD_SC_HS__NAND3_2%A
x_PM_SKY130_FD_SC_HS__NAND3_2%VPWR N_VPWR_M1004_d N_VPWR_M1006_d N_VPWR_M1003_d
+ N_VPWR_M1009_s N_VPWR_c_259_n N_VPWR_c_260_n N_VPWR_c_261_n N_VPWR_c_262_n
+ N_VPWR_c_263_n N_VPWR_c_264_n VPWR N_VPWR_c_265_n N_VPWR_c_266_n
+ N_VPWR_c_267_n N_VPWR_c_268_n N_VPWR_c_269_n N_VPWR_c_258_n
+ PM_SKY130_FD_SC_HS__NAND3_2%VPWR
x_PM_SKY130_FD_SC_HS__NAND3_2%Y N_Y_M1001_s N_Y_M1004_s N_Y_M1005_d N_Y_M1007_s
+ N_Y_c_318_n N_Y_c_315_n N_Y_c_325_n N_Y_c_329_n N_Y_c_349_n N_Y_c_350_n
+ N_Y_c_319_n N_Y_c_320_n N_Y_c_316_n N_Y_c_317_n Y Y
+ PM_SKY130_FD_SC_HS__NAND3_2%Y
x_PM_SKY130_FD_SC_HS__NAND3_2%A_27_74# N_A_27_74#_M1000_d N_A_27_74#_M1010_d
+ N_A_27_74#_M1008_s N_A_27_74#_c_402_n N_A_27_74#_c_407_n N_A_27_74#_c_415_n
+ N_A_27_74#_c_403_n N_A_27_74#_c_404_n N_A_27_74#_c_405_n
+ PM_SKY130_FD_SC_HS__NAND3_2%A_27_74#
x_PM_SKY130_FD_SC_HS__NAND3_2%VGND N_VGND_M1000_s N_VGND_c_461_n VGND
+ N_VGND_c_462_n N_VGND_c_463_n N_VGND_c_464_n N_VGND_c_465_n
+ PM_SKY130_FD_SC_HS__NAND3_2%VGND
x_PM_SKY130_FD_SC_HS__NAND3_2%A_283_74# N_A_283_74#_M1002_d N_A_283_74#_M1011_d
+ N_A_283_74#_c_501_n PM_SKY130_FD_SC_HS__NAND3_2%A_283_74#
cc_1 VNB N_C_c_58_n 0.0221619f $X=-0.19 $Y=-0.245 $X2=0.48 $Y2=1.22
cc_2 VNB N_C_c_59_n 0.0162301f $X=-0.19 $Y=-0.245 $X2=0.91 $Y2=1.22
cc_3 VNB N_C_c_60_n 0.0251517f $X=-0.19 $Y=-0.245 $X2=0.57 $Y2=1.385
cc_4 VNB N_C_c_61_n 0.0565946f $X=-0.19 $Y=-0.245 $X2=0.91 $Y2=1.492
cc_5 VNB N_B_M1002_g 0.0248915f $X=-0.19 $Y=-0.245 $X2=0.48 $Y2=0.74
cc_6 VNB N_B_c_110_n 0.0232379f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_7 VNB N_B_c_111_n 0.0357817f $X=-0.19 $Y=-0.245 $X2=0.91 $Y2=0.74
cc_8 VNB N_B_M1008_g 0.0280879f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_9 VNB N_B_c_113_n 3.02997e-19 $X=-0.19 $Y=-0.245 $X2=0.57 $Y2=1.385
cc_10 VNB N_B_c_114_n 0.01693f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_B_c_115_n 0.0054119f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_M1001_g 0.0198416f $X=-0.19 $Y=-0.245 $X2=0.48 $Y2=0.74
cc_13 VNB N_A_M1011_g 0.0203106f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=1.765
cc_14 VNB N_A_c_203_n 0.0389124f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.365
cc_15 VNB N_VPWR_c_258_n 0.143779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_Y_c_315_n 0.010102f $X=-0.19 $Y=-0.245 $X2=0.57 $Y2=1.385
cc_17 VNB N_Y_c_316_n 0.00300143f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_Y_c_317_n 0.00225359f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_27_74#_c_402_n 0.0172715f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=2.4
cc_20 VNB N_A_27_74#_c_403_n 0.0110846f $X=-0.19 $Y=-0.245 $X2=0.91 $Y2=1.492
cc_21 VNB N_A_27_74#_c_404_n 0.00213939f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_27_74#_c_405_n 0.0331002f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_VGND_c_461_n 0.00396467f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_24 VNB N_VGND_c_462_n 0.0162587f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=1.765
cc_25 VNB N_VGND_c_463_n 0.0629719f $X=-0.19 $Y=-0.245 $X2=0.91 $Y2=1.492
cc_26 VNB N_VGND_c_464_n 0.205212f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=1.492
cc_27 VNB N_VGND_c_465_n 0.00601569f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_283_74#_c_501_n 0.0141546f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=2.4
cc_29 VPB N_C_c_62_n 0.0176529f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.765
cc_30 VPB N_C_c_63_n 0.0157238f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=1.765
cc_31 VPB N_C_c_61_n 0.0161072f $X=-0.19 $Y=1.66 $X2=0.91 $Y2=1.492
cc_32 VPB N_B_c_110_n 0.0269807f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.4
cc_33 VPB N_B_c_111_n 0.0272659f $X=-0.19 $Y=1.66 $X2=0.91 $Y2=0.74
cc_34 VPB N_B_c_113_n 0.00150792f $X=-0.19 $Y=1.66 $X2=0.57 $Y2=1.385
cc_35 VPB B 0.00120283f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_36 VPB N_B_c_115_n 0.00185734f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_37 VPB N_A_c_204_n 0.0162058f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.4
cc_38 VPB N_A_c_205_n 0.0157504f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=2.4
cc_39 VPB N_A_c_206_n 0.00362397f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=1.492
cc_40 VPB N_A_c_203_n 0.0219875f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=1.365
cc_41 VPB N_VPWR_c_259_n 0.0106521f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.21
cc_42 VPB N_VPWR_c_260_n 0.0575161f $X=-0.19 $Y=1.66 $X2=0.48 $Y2=1.492
cc_43 VPB N_VPWR_c_261_n 0.00886117f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=1.492
cc_44 VPB N_VPWR_c_262_n 0.0059435f $X=-0.19 $Y=1.66 $X2=0.57 $Y2=1.365
cc_45 VPB N_VPWR_c_263_n 0.0106521f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_46 VPB N_VPWR_c_264_n 0.0572108f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_47 VPB N_VPWR_c_265_n 0.0196495f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_48 VPB N_VPWR_c_266_n 0.0196495f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_49 VPB N_VPWR_c_267_n 0.0183691f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_50 VPB N_VPWR_c_268_n 0.0047828f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_51 VPB N_VPWR_c_269_n 0.00614127f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_52 VPB N_VPWR_c_258_n 0.0638197f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_53 VPB N_Y_c_318_n 0.00257348f $X=-0.19 $Y=1.66 $X2=0.48 $Y2=1.492
cc_54 VPB N_Y_c_319_n 0.00234639f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_55 VPB N_Y_c_320_n 0.00597034f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_56 VPB N_Y_c_316_n 0.00122694f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_57 VPB Y 0.00261707f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_58 N_C_c_59_n N_B_M1002_g 0.0140681f $X=0.91 $Y=1.22 $X2=0 $Y2=0
cc_59 N_C_c_61_n N_B_M1002_g 0.0166541f $X=0.91 $Y=1.492 $X2=0 $Y2=0
cc_60 N_C_c_63_n N_B_c_110_n 0.0341021f $X=0.955 $Y=1.765 $X2=0 $Y2=0
cc_61 N_C_c_61_n N_B_c_110_n 0.0109215f $X=0.91 $Y=1.492 $X2=0 $Y2=0
cc_62 N_C_c_63_n B 2.04481e-19 $X=0.955 $Y=1.765 $X2=0 $Y2=0
cc_63 N_C_c_61_n N_B_c_115_n 2.78603e-19 $X=0.91 $Y=1.492 $X2=0 $Y2=0
cc_64 N_C_c_62_n N_VPWR_c_260_n 0.0100916f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_65 N_C_c_60_n N_VPWR_c_260_n 0.0154298f $X=0.57 $Y=1.385 $X2=0 $Y2=0
cc_66 N_C_c_63_n N_VPWR_c_261_n 0.00490136f $X=0.955 $Y=1.765 $X2=0 $Y2=0
cc_67 N_C_c_62_n N_VPWR_c_265_n 0.00445602f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_68 N_C_c_63_n N_VPWR_c_265_n 0.00445602f $X=0.955 $Y=1.765 $X2=0 $Y2=0
cc_69 N_C_c_62_n N_VPWR_c_258_n 0.00861084f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_70 N_C_c_63_n N_VPWR_c_258_n 0.00857432f $X=0.955 $Y=1.765 $X2=0 $Y2=0
cc_71 N_C_c_62_n N_Y_c_318_n 0.00627458f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_72 N_C_c_63_n N_Y_c_318_n 0.00717212f $X=0.955 $Y=1.765 $X2=0 $Y2=0
cc_73 N_C_c_58_n N_Y_c_325_n 5.01846e-19 $X=0.48 $Y=1.22 $X2=0 $Y2=0
cc_74 N_C_c_59_n N_Y_c_325_n 0.0049118f $X=0.91 $Y=1.22 $X2=0 $Y2=0
cc_75 N_C_c_60_n N_Y_c_325_n 0.0061979f $X=0.57 $Y=1.385 $X2=0 $Y2=0
cc_76 N_C_c_61_n N_Y_c_325_n 0.00189162f $X=0.91 $Y=1.492 $X2=0 $Y2=0
cc_77 N_C_c_63_n N_Y_c_329_n 3.73103e-19 $X=0.955 $Y=1.765 $X2=0 $Y2=0
cc_78 N_C_c_62_n N_Y_c_320_n 0.00768381f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_79 N_C_c_63_n N_Y_c_320_n 0.0227034f $X=0.955 $Y=1.765 $X2=0 $Y2=0
cc_80 N_C_c_60_n N_Y_c_320_n 0.0101111f $X=0.57 $Y=1.385 $X2=0 $Y2=0
cc_81 N_C_c_61_n N_Y_c_320_n 0.00412691f $X=0.91 $Y=1.492 $X2=0 $Y2=0
cc_82 N_C_c_62_n N_Y_c_316_n 3.0365e-19 $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_83 N_C_c_63_n N_Y_c_316_n 0.00159392f $X=0.955 $Y=1.765 $X2=0 $Y2=0
cc_84 N_C_c_60_n N_Y_c_316_n 0.0199139f $X=0.57 $Y=1.385 $X2=0 $Y2=0
cc_85 N_C_c_61_n N_Y_c_316_n 0.0164121f $X=0.91 $Y=1.492 $X2=0 $Y2=0
cc_86 N_C_c_63_n Y 6.08775e-19 $X=0.955 $Y=1.765 $X2=0 $Y2=0
cc_87 N_C_c_58_n N_A_27_74#_c_402_n 4.43891e-19 $X=0.48 $Y=1.22 $X2=0 $Y2=0
cc_88 N_C_c_58_n N_A_27_74#_c_407_n 0.00948928f $X=0.48 $Y=1.22 $X2=0 $Y2=0
cc_89 N_C_c_59_n N_A_27_74#_c_407_n 0.0125772f $X=0.91 $Y=1.22 $X2=0 $Y2=0
cc_90 N_C_c_60_n N_A_27_74#_c_407_n 0.0153562f $X=0.57 $Y=1.385 $X2=0 $Y2=0
cc_91 N_C_c_61_n N_A_27_74#_c_407_n 8.56627e-19 $X=0.91 $Y=1.492 $X2=0 $Y2=0
cc_92 N_C_c_58_n N_A_27_74#_c_403_n 0.00343023f $X=0.48 $Y=1.22 $X2=0 $Y2=0
cc_93 N_C_c_59_n N_A_27_74#_c_403_n 5.20319e-19 $X=0.91 $Y=1.22 $X2=0 $Y2=0
cc_94 N_C_c_60_n N_A_27_74#_c_403_n 0.0236506f $X=0.57 $Y=1.385 $X2=0 $Y2=0
cc_95 N_C_c_59_n N_A_27_74#_c_404_n 2.82836e-19 $X=0.91 $Y=1.22 $X2=0 $Y2=0
cc_96 N_C_c_58_n N_VGND_c_461_n 0.0095457f $X=0.48 $Y=1.22 $X2=0 $Y2=0
cc_97 N_C_c_59_n N_VGND_c_461_n 0.00663018f $X=0.91 $Y=1.22 $X2=0 $Y2=0
cc_98 N_C_c_58_n N_VGND_c_462_n 0.00281948f $X=0.48 $Y=1.22 $X2=0 $Y2=0
cc_99 N_C_c_59_n N_VGND_c_463_n 0.00281141f $X=0.91 $Y=1.22 $X2=0 $Y2=0
cc_100 N_C_c_58_n N_VGND_c_464_n 0.00367131f $X=0.48 $Y=1.22 $X2=0 $Y2=0
cc_101 N_C_c_59_n N_VGND_c_464_n 0.00365164f $X=0.91 $Y=1.22 $X2=0 $Y2=0
cc_102 N_B_M1002_g N_A_M1001_g 0.0311226f $X=1.34 $Y=0.74 $X2=0 $Y2=0
cc_103 N_B_c_110_n N_A_c_204_n 0.0234952f $X=1.455 $Y=1.765 $X2=0 $Y2=0
cc_104 N_B_c_129_p N_A_c_204_n 0.0149567f $X=2.655 $Y=2.035 $X2=0 $Y2=0
cc_105 B N_A_c_204_n 0.0023224f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_106 N_B_c_111_n N_A_M1011_g 9.74524e-19 $X=2.855 $Y=1.765 $X2=0 $Y2=0
cc_107 N_B_M1008_g N_A_M1011_g 0.0295756f $X=2.88 $Y=0.795 $X2=0 $Y2=0
cc_108 N_B_c_114_n N_A_M1011_g 6.56671e-19 $X=2.9 $Y=1.485 $X2=0 $Y2=0
cc_109 N_B_c_111_n N_A_c_205_n 0.0232072f $X=2.855 $Y=1.765 $X2=0 $Y2=0
cc_110 N_B_c_129_p N_A_c_205_n 0.015369f $X=2.655 $Y=2.035 $X2=0 $Y2=0
cc_111 N_B_c_113_n N_A_c_205_n 0.00362556f $X=2.74 $Y=1.95 $X2=0 $Y2=0
cc_112 N_B_c_110_n N_A_c_206_n 2.87328e-19 $X=1.455 $Y=1.765 $X2=0 $Y2=0
cc_113 N_B_c_111_n N_A_c_206_n 2.14427e-19 $X=2.855 $Y=1.765 $X2=0 $Y2=0
cc_114 N_B_c_129_p N_A_c_206_n 0.022842f $X=2.655 $Y=2.035 $X2=0 $Y2=0
cc_115 N_B_c_113_n N_A_c_206_n 0.00598821f $X=2.74 $Y=1.95 $X2=0 $Y2=0
cc_116 N_B_c_114_n N_A_c_206_n 0.0101158f $X=2.9 $Y=1.485 $X2=0 $Y2=0
cc_117 B N_A_c_206_n 0.00790544f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_118 N_B_c_115_n N_A_c_206_n 0.015572f $X=1.61 $Y=1.68 $X2=0 $Y2=0
cc_119 N_B_c_110_n N_A_c_203_n 0.0244685f $X=1.455 $Y=1.765 $X2=0 $Y2=0
cc_120 N_B_c_111_n N_A_c_203_n 0.0217358f $X=2.855 $Y=1.765 $X2=0 $Y2=0
cc_121 N_B_c_129_p N_A_c_203_n 0.00147342f $X=2.655 $Y=2.035 $X2=0 $Y2=0
cc_122 N_B_c_113_n N_A_c_203_n 9.35193e-19 $X=2.74 $Y=1.95 $X2=0 $Y2=0
cc_123 N_B_c_114_n N_A_c_203_n 0.00414741f $X=2.9 $Y=1.485 $X2=0 $Y2=0
cc_124 B N_A_c_203_n 6.884e-19 $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_125 N_B_c_115_n N_A_c_203_n 0.00171302f $X=1.61 $Y=1.68 $X2=0 $Y2=0
cc_126 N_B_c_129_p N_VPWR_M1003_d 0.00446461f $X=2.655 $Y=2.035 $X2=0 $Y2=0
cc_127 N_B_c_110_n N_VPWR_c_261_n 0.00417074f $X=1.455 $Y=1.765 $X2=0 $Y2=0
cc_128 N_B_c_111_n N_VPWR_c_262_n 4.41818e-19 $X=2.855 $Y=1.765 $X2=0 $Y2=0
cc_129 N_B_c_111_n N_VPWR_c_264_n 0.0132689f $X=2.855 $Y=1.765 $X2=0 $Y2=0
cc_130 N_B_c_129_p N_VPWR_c_264_n 0.0137304f $X=2.655 $Y=2.035 $X2=0 $Y2=0
cc_131 N_B_c_113_n N_VPWR_c_264_n 0.00940176f $X=2.74 $Y=1.95 $X2=0 $Y2=0
cc_132 N_B_c_114_n N_VPWR_c_264_n 0.005819f $X=2.9 $Y=1.485 $X2=0 $Y2=0
cc_133 N_B_c_110_n N_VPWR_c_266_n 0.00445602f $X=1.455 $Y=1.765 $X2=0 $Y2=0
cc_134 N_B_c_111_n N_VPWR_c_267_n 0.00445602f $X=2.855 $Y=1.765 $X2=0 $Y2=0
cc_135 N_B_c_110_n N_VPWR_c_258_n 0.00858232f $X=1.455 $Y=1.765 $X2=0 $Y2=0
cc_136 N_B_c_111_n N_VPWR_c_258_n 0.00861168f $X=2.855 $Y=1.765 $X2=0 $Y2=0
cc_137 N_B_c_162_p N_Y_M1005_d 0.00210282f $X=1.795 $Y=2.035 $X2=0 $Y2=0
cc_138 N_B_c_129_p N_Y_M1007_s 0.00644106f $X=2.655 $Y=2.035 $X2=0 $Y2=0
cc_139 N_B_c_113_n N_Y_M1007_s 0.00126846f $X=2.74 $Y=1.95 $X2=0 $Y2=0
cc_140 N_B_c_110_n N_Y_c_318_n 5.26453e-19 $X=1.455 $Y=1.765 $X2=0 $Y2=0
cc_141 N_B_M1002_g N_Y_c_315_n 0.0112384f $X=1.34 $Y=0.74 $X2=0 $Y2=0
cc_142 N_B_c_110_n N_Y_c_315_n 0.00494603f $X=1.455 $Y=1.765 $X2=0 $Y2=0
cc_143 N_B_c_115_n N_Y_c_315_n 0.0363457f $X=1.61 $Y=1.68 $X2=0 $Y2=0
cc_144 N_B_c_110_n N_Y_c_329_n 0.0126066f $X=1.455 $Y=1.765 $X2=0 $Y2=0
cc_145 N_B_c_162_p N_Y_c_329_n 0.00678794f $X=1.795 $Y=2.035 $X2=0 $Y2=0
cc_146 N_B_c_115_n N_Y_c_329_n 0.00334286f $X=1.61 $Y=1.68 $X2=0 $Y2=0
cc_147 N_B_c_129_p N_Y_c_349_n 0.0363668f $X=2.655 $Y=2.035 $X2=0 $Y2=0
cc_148 N_B_c_111_n N_Y_c_350_n 0.00202157f $X=2.855 $Y=1.765 $X2=0 $Y2=0
cc_149 N_B_c_129_p N_Y_c_350_n 0.0167008f $X=2.655 $Y=2.035 $X2=0 $Y2=0
cc_150 N_B_c_111_n N_Y_c_319_n 0.00641576f $X=2.855 $Y=1.765 $X2=0 $Y2=0
cc_151 N_B_c_162_p N_Y_c_320_n 0.0087026f $X=1.795 $Y=2.035 $X2=0 $Y2=0
cc_152 N_B_M1002_g N_Y_c_316_n 0.00348765f $X=1.34 $Y=0.74 $X2=0 $Y2=0
cc_153 N_B_c_110_n N_Y_c_316_n 0.00785115f $X=1.455 $Y=1.765 $X2=0 $Y2=0
cc_154 B N_Y_c_316_n 0.0127675f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_155 N_B_c_115_n N_Y_c_316_n 0.0192485f $X=1.61 $Y=1.68 $X2=0 $Y2=0
cc_156 N_B_M1002_g N_Y_c_317_n 7.95487e-19 $X=1.34 $Y=0.74 $X2=0 $Y2=0
cc_157 N_B_M1008_g N_Y_c_317_n 0.00117715f $X=2.88 $Y=0.795 $X2=0 $Y2=0
cc_158 N_B_c_110_n Y 0.00780548f $X=1.455 $Y=1.765 $X2=0 $Y2=0
cc_159 N_B_c_129_p Y 7.20378e-19 $X=2.655 $Y=2.035 $X2=0 $Y2=0
cc_160 N_B_c_162_p Y 0.0182573f $X=1.795 $Y=2.035 $X2=0 $Y2=0
cc_161 N_B_M1002_g N_A_27_74#_c_415_n 0.00503198f $X=1.34 $Y=0.74 $X2=0 $Y2=0
cc_162 N_B_c_111_n N_A_27_74#_c_415_n 0.00106907f $X=2.855 $Y=1.765 $X2=0 $Y2=0
cc_163 N_B_M1008_g N_A_27_74#_c_415_n 0.010205f $X=2.88 $Y=0.795 $X2=0 $Y2=0
cc_164 N_B_c_114_n N_A_27_74#_c_415_n 0.00722399f $X=2.9 $Y=1.485 $X2=0 $Y2=0
cc_165 N_B_M1002_g N_A_27_74#_c_404_n 0.00980692f $X=1.34 $Y=0.74 $X2=0 $Y2=0
cc_166 N_B_c_111_n N_A_27_74#_c_405_n 0.00238884f $X=2.855 $Y=1.765 $X2=0 $Y2=0
cc_167 N_B_M1008_g N_A_27_74#_c_405_n 0.0138289f $X=2.88 $Y=0.795 $X2=0 $Y2=0
cc_168 N_B_c_114_n N_A_27_74#_c_405_n 0.00838142f $X=2.9 $Y=1.485 $X2=0 $Y2=0
cc_169 N_B_M1002_g N_VGND_c_461_n 3.89995e-19 $X=1.34 $Y=0.74 $X2=0 $Y2=0
cc_170 N_B_M1002_g N_VGND_c_463_n 0.00321733f $X=1.34 $Y=0.74 $X2=0 $Y2=0
cc_171 N_B_M1008_g N_VGND_c_463_n 0.00407143f $X=2.88 $Y=0.795 $X2=0 $Y2=0
cc_172 N_B_M1002_g N_VGND_c_464_n 0.00409122f $X=1.34 $Y=0.74 $X2=0 $Y2=0
cc_173 N_B_M1008_g N_VGND_c_464_n 0.00528353f $X=2.88 $Y=0.795 $X2=0 $Y2=0
cc_174 N_B_M1002_g N_A_283_74#_c_501_n 0.00260352f $X=1.34 $Y=0.74 $X2=0 $Y2=0
cc_175 N_B_M1008_g N_A_283_74#_c_501_n 0.00391613f $X=2.88 $Y=0.795 $X2=0 $Y2=0
cc_176 N_A_c_204_n N_VPWR_c_262_n 0.00331824f $X=1.91 $Y=1.765 $X2=0 $Y2=0
cc_177 N_A_c_205_n N_VPWR_c_262_n 0.00746735f $X=2.405 $Y=1.765 $X2=0 $Y2=0
cc_178 N_A_c_204_n N_VPWR_c_266_n 0.00451267f $X=1.91 $Y=1.765 $X2=0 $Y2=0
cc_179 N_A_c_205_n N_VPWR_c_267_n 0.00413917f $X=2.405 $Y=1.765 $X2=0 $Y2=0
cc_180 N_A_c_204_n N_VPWR_c_258_n 0.00875694f $X=1.91 $Y=1.765 $X2=0 $Y2=0
cc_181 N_A_c_205_n N_VPWR_c_258_n 0.0081781f $X=2.405 $Y=1.765 $X2=0 $Y2=0
cc_182 N_A_M1001_g N_Y_c_315_n 0.0134717f $X=1.895 $Y=0.795 $X2=0 $Y2=0
cc_183 N_A_c_204_n N_Y_c_349_n 0.0124044f $X=1.91 $Y=1.765 $X2=0 $Y2=0
cc_184 N_A_c_205_n N_Y_c_349_n 0.0127199f $X=2.405 $Y=1.765 $X2=0 $Y2=0
cc_185 N_A_c_205_n N_Y_c_319_n 3.8272e-19 $X=2.405 $Y=1.765 $X2=0 $Y2=0
cc_186 N_A_M1001_g N_Y_c_317_n 0.00643082f $X=1.895 $Y=0.795 $X2=0 $Y2=0
cc_187 N_A_M1011_g N_Y_c_317_n 0.00830615f $X=2.325 $Y=0.795 $X2=0 $Y2=0
cc_188 N_A_c_206_n N_Y_c_317_n 0.0245791f $X=2.13 $Y=1.515 $X2=0 $Y2=0
cc_189 N_A_c_203_n N_Y_c_317_n 0.00250645f $X=2.325 $Y=1.557 $X2=0 $Y2=0
cc_190 N_A_c_204_n Y 0.00705236f $X=1.91 $Y=1.765 $X2=0 $Y2=0
cc_191 N_A_c_205_n Y 8.03342e-19 $X=2.405 $Y=1.765 $X2=0 $Y2=0
cc_192 N_A_M1001_g N_A_27_74#_c_415_n 0.0117007f $X=1.895 $Y=0.795 $X2=0 $Y2=0
cc_193 N_A_M1011_g N_A_27_74#_c_415_n 0.0145843f $X=2.325 $Y=0.795 $X2=0 $Y2=0
cc_194 N_A_c_206_n N_A_27_74#_c_415_n 4.60142e-19 $X=2.13 $Y=1.515 $X2=0 $Y2=0
cc_195 N_A_c_203_n N_A_27_74#_c_415_n 0.00189149f $X=2.325 $Y=1.557 $X2=0 $Y2=0
cc_196 N_A_M1001_g N_A_27_74#_c_404_n 8.11839e-19 $X=1.895 $Y=0.795 $X2=0 $Y2=0
cc_197 N_A_M1011_g N_A_27_74#_c_405_n 0.00223206f $X=2.325 $Y=0.795 $X2=0 $Y2=0
cc_198 N_A_M1001_g N_VGND_c_463_n 8.63546e-19 $X=1.895 $Y=0.795 $X2=0 $Y2=0
cc_199 N_A_M1011_g N_VGND_c_463_n 8.63546e-19 $X=2.325 $Y=0.795 $X2=0 $Y2=0
cc_200 N_A_M1001_g N_A_283_74#_c_501_n 0.00941316f $X=1.895 $Y=0.795 $X2=0 $Y2=0
cc_201 N_A_M1011_g N_A_283_74#_c_501_n 0.00942684f $X=2.325 $Y=0.795 $X2=0 $Y2=0
cc_202 N_VPWR_c_261_n N_Y_c_318_n 0.0138908f $X=1.23 $Y=2.795 $X2=0 $Y2=0
cc_203 N_VPWR_c_265_n N_Y_c_318_n 0.014552f $X=1.065 $Y=3.33 $X2=0 $Y2=0
cc_204 N_VPWR_c_258_n N_Y_c_318_n 0.0119791f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_205 N_VPWR_M1006_d N_Y_c_329_n 0.01056f $X=1.03 $Y=1.84 $X2=0 $Y2=0
cc_206 N_VPWR_c_261_n N_Y_c_329_n 0.0178175f $X=1.23 $Y=2.795 $X2=0 $Y2=0
cc_207 N_VPWR_M1003_d N_Y_c_349_n 0.00471201f $X=1.985 $Y=1.84 $X2=0 $Y2=0
cc_208 N_VPWR_c_262_n N_Y_c_349_n 0.0198182f $X=2.18 $Y=2.795 $X2=0 $Y2=0
cc_209 N_VPWR_c_264_n N_Y_c_350_n 0.0121024f $X=3.08 $Y=1.985 $X2=0 $Y2=0
cc_210 N_VPWR_c_262_n N_Y_c_319_n 0.013281f $X=2.18 $Y=2.795 $X2=0 $Y2=0
cc_211 N_VPWR_c_264_n N_Y_c_319_n 0.0343455f $X=3.08 $Y=1.985 $X2=0 $Y2=0
cc_212 N_VPWR_c_267_n N_Y_c_319_n 0.0119293f $X=2.995 $Y=3.33 $X2=0 $Y2=0
cc_213 N_VPWR_c_258_n N_Y_c_319_n 0.00983555f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_214 N_VPWR_M1006_d N_Y_c_320_n 0.0063329f $X=1.03 $Y=1.84 $X2=0 $Y2=0
cc_215 N_VPWR_c_260_n N_Y_c_320_n 0.0793896f $X=0.28 $Y=1.985 $X2=0 $Y2=0
cc_216 N_VPWR_c_261_n N_Y_c_320_n 6.31132e-19 $X=1.23 $Y=2.795 $X2=0 $Y2=0
cc_217 N_VPWR_c_261_n Y 0.0234974f $X=1.23 $Y=2.795 $X2=0 $Y2=0
cc_218 N_VPWR_c_262_n Y 0.0139233f $X=2.18 $Y=2.795 $X2=0 $Y2=0
cc_219 N_VPWR_c_266_n Y 0.0145824f $X=2.015 $Y=3.33 $X2=0 $Y2=0
cc_220 N_VPWR_c_258_n Y 0.0120092f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_221 N_VPWR_c_264_n N_A_27_74#_c_405_n 0.00608804f $X=3.08 $Y=1.985 $X2=0
+ $Y2=0
cc_222 N_Y_c_315_n N_A_27_74#_M1010_d 0.00119058f $X=1.945 $Y=1.175 $X2=0 $Y2=0
cc_223 N_Y_c_325_n N_A_27_74#_M1010_d 5.86511e-19 $X=1.095 $Y=1.175 $X2=0 $Y2=0
cc_224 N_Y_c_325_n N_A_27_74#_c_407_n 0.00453647f $X=1.095 $Y=1.175 $X2=0 $Y2=0
cc_225 N_Y_M1001_s N_A_27_74#_c_415_n 0.003356f $X=1.97 $Y=0.425 $X2=0 $Y2=0
cc_226 N_Y_c_315_n N_A_27_74#_c_415_n 0.0199657f $X=1.945 $Y=1.175 $X2=0 $Y2=0
cc_227 N_Y_c_317_n N_A_27_74#_c_415_n 0.0160991f $X=2.11 $Y=1.02 $X2=0 $Y2=0
cc_228 N_Y_c_315_n N_A_27_74#_c_404_n 0.0165421f $X=1.945 $Y=1.175 $X2=0 $Y2=0
cc_229 N_Y_c_325_n N_A_27_74#_c_404_n 0.00472879f $X=1.095 $Y=1.175 $X2=0 $Y2=0
cc_230 N_Y_c_317_n N_A_27_74#_c_405_n 0.00523618f $X=2.11 $Y=1.02 $X2=0 $Y2=0
cc_231 N_Y_c_315_n N_A_283_74#_M1002_d 0.00437664f $X=1.945 $Y=1.175 $X2=-0.19
+ $Y2=-0.245
cc_232 N_A_27_74#_c_407_n N_VGND_M1000_s 0.00447978f $X=1.04 $Y=0.835 $X2=-0.19
+ $Y2=-0.245
cc_233 N_A_27_74#_c_402_n N_VGND_c_461_n 0.00897147f $X=0.265 $Y=0.515 $X2=0
+ $Y2=0
cc_234 N_A_27_74#_c_407_n N_VGND_c_461_n 0.0165203f $X=1.04 $Y=0.835 $X2=0 $Y2=0
cc_235 N_A_27_74#_c_404_n N_VGND_c_461_n 0.0104177f $X=1.205 $Y=0.68 $X2=0 $Y2=0
cc_236 N_A_27_74#_c_402_n N_VGND_c_462_n 0.0110419f $X=0.265 $Y=0.515 $X2=0
+ $Y2=0
cc_237 N_A_27_74#_c_407_n N_VGND_c_462_n 0.00125985f $X=1.04 $Y=0.835 $X2=0
+ $Y2=0
cc_238 N_A_27_74#_c_403_n N_VGND_c_462_n 7.09218e-19 $X=0.265 $Y=0.835 $X2=0
+ $Y2=0
cc_239 N_A_27_74#_c_407_n N_VGND_c_463_n 0.00197156f $X=1.04 $Y=0.835 $X2=0
+ $Y2=0
cc_240 N_A_27_74#_c_415_n N_VGND_c_463_n 0.00390932f $X=2.93 $Y=0.68 $X2=0 $Y2=0
cc_241 N_A_27_74#_c_404_n N_VGND_c_463_n 0.0107219f $X=1.205 $Y=0.68 $X2=0 $Y2=0
cc_242 N_A_27_74#_c_405_n N_VGND_c_463_n 0.0117675f $X=3.095 $Y=0.57 $X2=0 $Y2=0
cc_243 N_A_27_74#_c_402_n N_VGND_c_464_n 0.00915013f $X=0.265 $Y=0.515 $X2=0
+ $Y2=0
cc_244 N_A_27_74#_c_407_n N_VGND_c_464_n 0.00743138f $X=1.04 $Y=0.835 $X2=0
+ $Y2=0
cc_245 N_A_27_74#_c_415_n N_VGND_c_464_n 0.00964348f $X=2.93 $Y=0.68 $X2=0 $Y2=0
cc_246 N_A_27_74#_c_403_n N_VGND_c_464_n 0.00196697f $X=0.265 $Y=0.835 $X2=0
+ $Y2=0
cc_247 N_A_27_74#_c_404_n N_VGND_c_464_n 0.0106167f $X=1.205 $Y=0.68 $X2=0 $Y2=0
cc_248 N_A_27_74#_c_405_n N_VGND_c_464_n 0.0116783f $X=3.095 $Y=0.57 $X2=0 $Y2=0
cc_249 N_A_27_74#_c_415_n N_A_283_74#_M1002_d 0.00737496f $X=2.93 $Y=0.68
+ $X2=-0.19 $Y2=-0.245
cc_250 N_A_27_74#_c_415_n N_A_283_74#_M1011_d 0.0118482f $X=2.93 $Y=0.68 $X2=0
+ $Y2=0
cc_251 N_A_27_74#_c_415_n N_A_283_74#_c_501_n 0.0797775f $X=2.93 $Y=0.68 $X2=0
+ $Y2=0
cc_252 N_A_27_74#_c_404_n N_A_283_74#_c_501_n 0.0025548f $X=1.205 $Y=0.68 $X2=0
+ $Y2=0
cc_253 N_A_27_74#_c_405_n N_A_283_74#_c_501_n 0.00153676f $X=3.095 $Y=0.57 $X2=0
+ $Y2=0
cc_254 N_VGND_c_464_n N_A_283_74#_M1002_d 0.00230295f $X=3.12 $Y=0 $X2=-0.19
+ $Y2=-0.245
cc_255 N_VGND_c_464_n N_A_283_74#_M1011_d 0.00247946f $X=3.12 $Y=0 $X2=0 $Y2=0
cc_256 N_VGND_c_461_n N_A_283_74#_c_501_n 0.00240443f $X=0.695 $Y=0.495 $X2=0
+ $Y2=0
cc_257 N_VGND_c_463_n N_A_283_74#_c_501_n 0.0838614f $X=3.12 $Y=0 $X2=0 $Y2=0
cc_258 N_VGND_c_464_n N_A_283_74#_c_501_n 0.0492532f $X=3.12 $Y=0 $X2=0 $Y2=0
