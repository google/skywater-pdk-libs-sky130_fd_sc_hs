* File: sky130_fd_sc_hs__nand3_4.pxi.spice
* Created: Thu Aug 27 20:51:09 2020
* 
x_PM_SKY130_FD_SC_HS__NAND3_4%A N_A_c_87_n N_A_M1004_g N_A_c_92_n N_A_M1006_g
+ N_A_c_88_n N_A_M1009_g N_A_c_89_n N_A_M1010_g N_A_c_93_n N_A_M1014_g
+ N_A_c_90_n N_A_M1017_g A A N_A_c_94_n N_A_c_91_n PM_SKY130_FD_SC_HS__NAND3_4%A
x_PM_SKY130_FD_SC_HS__NAND3_4%B N_B_c_156_n N_B_M1015_g N_B_M1002_g N_B_c_157_n
+ N_B_M1016_g N_B_M1003_g N_B_M1007_g N_B_M1013_g N_B_c_158_n N_B_c_153_n B B
+ N_B_c_155_n PM_SKY130_FD_SC_HS__NAND3_4%B
x_PM_SKY130_FD_SC_HS__NAND3_4%C N_C_c_221_n N_C_M1011_g N_C_c_222_n N_C_M1012_g
+ N_C_M1000_g N_C_M1001_g N_C_M1005_g N_C_M1008_g N_C_c_223_n N_C_c_227_n C C C
+ N_C_c_220_n PM_SKY130_FD_SC_HS__NAND3_4%C
x_PM_SKY130_FD_SC_HS__NAND3_4%VPWR N_VPWR_M1006_s N_VPWR_M1014_s N_VPWR_M1016_s
+ N_VPWR_M1012_s N_VPWR_c_280_n N_VPWR_c_281_n N_VPWR_c_282_n VPWR
+ N_VPWR_c_283_n N_VPWR_c_284_n N_VPWR_c_285_n N_VPWR_c_279_n N_VPWR_c_287_n
+ N_VPWR_c_288_n N_VPWR_c_289_n N_VPWR_c_290_n PM_SKY130_FD_SC_HS__NAND3_4%VPWR
x_PM_SKY130_FD_SC_HS__NAND3_4%Y N_Y_M1004_d N_Y_M1010_d N_Y_M1006_d N_Y_M1015_d
+ N_Y_M1011_d N_Y_c_333_n N_Y_c_334_n N_Y_c_347_n N_Y_c_338_n N_Y_c_349_n
+ N_Y_c_339_n N_Y_c_335_n N_Y_c_359_n N_Y_c_362_n N_Y_c_340_n N_Y_c_380_n
+ N_Y_c_341_n N_Y_c_342_n N_Y_c_336_n N_Y_c_370_n N_Y_c_343_n Y Y
+ PM_SKY130_FD_SC_HS__NAND3_4%Y
x_PM_SKY130_FD_SC_HS__NAND3_4%A_27_82# N_A_27_82#_M1004_s N_A_27_82#_M1009_s
+ N_A_27_82#_M1017_s N_A_27_82#_M1003_d N_A_27_82#_M1013_d N_A_27_82#_c_430_n
+ N_A_27_82#_c_431_n N_A_27_82#_c_432_n N_A_27_82#_c_460_n N_A_27_82#_c_433_n
+ N_A_27_82#_c_434_n N_A_27_82#_c_435_n N_A_27_82#_c_470_p N_A_27_82#_c_436_n
+ N_A_27_82#_c_437_n N_A_27_82#_c_438_n N_A_27_82#_c_439_n N_A_27_82#_c_440_n
+ PM_SKY130_FD_SC_HS__NAND3_4%A_27_82#
x_PM_SKY130_FD_SC_HS__NAND3_4%A_456_82# N_A_456_82#_M1002_s N_A_456_82#_M1007_s
+ N_A_456_82#_M1000_d N_A_456_82#_M1005_d N_A_456_82#_c_496_n
+ N_A_456_82#_c_497_n N_A_456_82#_c_498_n N_A_456_82#_c_499_n
+ N_A_456_82#_c_500_n N_A_456_82#_c_501_n N_A_456_82#_c_502_n
+ N_A_456_82#_c_503_n N_A_456_82#_c_504_n PM_SKY130_FD_SC_HS__NAND3_4%A_456_82#
x_PM_SKY130_FD_SC_HS__NAND3_4%VGND N_VGND_M1000_s N_VGND_M1001_s N_VGND_M1008_s
+ N_VGND_c_562_n N_VGND_c_563_n N_VGND_c_564_n N_VGND_c_565_n N_VGND_c_566_n
+ N_VGND_c_567_n VGND N_VGND_c_568_n N_VGND_c_569_n N_VGND_c_570_n
+ N_VGND_c_571_n PM_SKY130_FD_SC_HS__NAND3_4%VGND
cc_1 VNB N_A_c_87_n 0.015797f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=1.225
cc_2 VNB N_A_c_88_n 0.0132349f $X=-0.19 $Y=-0.245 $X2=0.915 $Y2=1.225
cc_3 VNB N_A_c_89_n 0.0132368f $X=-0.19 $Y=-0.245 $X2=1.345 $Y2=1.225
cc_4 VNB N_A_c_90_n 0.0135128f $X=-0.19 $Y=-0.245 $X2=1.775 $Y2=1.225
cc_5 VNB N_A_c_91_n 0.0965248f $X=-0.19 $Y=-0.245 $X2=1.475 $Y2=1.495
cc_6 VNB N_B_M1002_g 0.0201101f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_7 VNB N_B_M1003_g 0.0196775f $X=-0.19 $Y=-0.245 $X2=1.475 $Y2=1.765
cc_8 VNB N_B_M1007_g 0.0196642f $X=-0.19 $Y=-0.245 $X2=1.775 $Y2=0.78
cc_9 VNB N_B_M1013_g 0.026969f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_B_c_153_n 0.00319621f $X=-0.19 $Y=-0.245 $X2=1.37 $Y2=1.515
cc_11 VNB B 0.00401758f $X=-0.19 $Y=-0.245 $X2=1.775 $Y2=1.225
cc_12 VNB N_B_c_155_n 0.0756615f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_C_M1000_g 0.0267451f $X=-0.19 $Y=-0.245 $X2=0.915 $Y2=0.78
cc_14 VNB N_C_M1001_g 0.0194534f $X=-0.19 $Y=-0.245 $X2=1.475 $Y2=1.765
cc_15 VNB N_C_M1005_g 0.0194534f $X=-0.19 $Y=-0.245 $X2=1.775 $Y2=0.78
cc_16 VNB N_C_M1008_g 0.0268263f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB C 0.0168872f $X=-0.19 $Y=-0.245 $X2=0.69 $Y2=1.565
cc_18 VNB N_C_c_220_n 0.10532f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_VPWR_c_279_n 0.263193f $X=-0.19 $Y=-0.245 $X2=1.37 $Y2=1.565
cc_20 VNB N_Y_c_333_n 0.00185509f $X=-0.19 $Y=-0.245 $X2=1.775 $Y2=1.225
cc_21 VNB N_Y_c_334_n 0.00754943f $X=-0.19 $Y=-0.245 $X2=1.775 $Y2=0.78
cc_22 VNB N_Y_c_335_n 0.00761155f $X=-0.19 $Y=-0.245 $X2=0.915 $Y2=1.495
cc_23 VNB N_Y_c_336_n 0.0022752f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB Y 0.0235986f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_27_82#_c_430_n 0.0164624f $X=-0.19 $Y=-0.245 $X2=1.775 $Y2=0.78
cc_26 VNB N_A_27_82#_c_431_n 0.00489863f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.58
cc_27 VNB N_A_27_82#_c_432_n 0.00945765f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_27_82#_c_433_n 0.00489863f $X=-0.19 $Y=-0.245 $X2=0.69 $Y2=1.515
cc_29 VNB N_A_27_82#_c_434_n 0.00267069f $X=-0.19 $Y=-0.245 $X2=1.37 $Y2=1.495
cc_30 VNB N_A_27_82#_c_435_n 0.00482743f $X=-0.19 $Y=-0.245 $X2=1.37 $Y2=1.515
cc_31 VNB N_A_27_82#_c_436_n 0.0087562f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_27_82#_c_437_n 0.00308948f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_27_82#_c_438_n 0.00121984f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_27_82#_c_439_n 0.00123754f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_27_82#_c_440_n 0.00136117f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_456_82#_c_496_n 0.00231524f $X=-0.19 $Y=-0.245 $X2=1.475 $Y2=1.765
cc_37 VNB N_A_456_82#_c_497_n 0.0211452f $X=-0.19 $Y=-0.245 $X2=1.475 $Y2=2.4
cc_38 VNB N_A_456_82#_c_498_n 0.00207241f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_39 VNB N_A_456_82#_c_499_n 0.00317575f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_456_82#_c_500_n 0.00140393f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=1.495
cc_41 VNB N_A_456_82#_c_501_n 0.00188975f $X=-0.19 $Y=-0.245 $X2=0.69 $Y2=1.495
cc_42 VNB N_A_456_82#_c_502_n 0.0023444f $X=-0.19 $Y=-0.245 $X2=0.915 $Y2=1.495
cc_43 VNB N_A_456_82#_c_503_n 0.0023444f $X=-0.19 $Y=-0.245 $X2=1.475 $Y2=1.495
cc_44 VNB N_A_456_82#_c_504_n 0.00145912f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_VGND_c_562_n 0.0102622f $X=-0.19 $Y=-0.245 $X2=1.345 $Y2=0.78
cc_46 VNB N_VGND_c_563_n 0.00367233f $X=-0.19 $Y=-0.245 $X2=1.775 $Y2=1.225
cc_47 VNB N_VGND_c_564_n 0.0118978f $X=-0.19 $Y=-0.245 $X2=1.775 $Y2=0.78
cc_48 VNB N_VGND_c_565_n 0.0441986f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.58
cc_49 VNB N_VGND_c_566_n 0.0967194f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=1.495
cc_50 VNB N_VGND_c_567_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.495
cc_51 VNB N_VGND_c_568_n 0.0154442f $X=-0.19 $Y=-0.245 $X2=1.775 $Y2=1.225
cc_52 VNB N_VGND_c_569_n 0.0155887f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_VGND_c_570_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_VGND_c_571_n 0.368708f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VPB N_A_c_92_n 0.0222963f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.765
cc_56 VPB N_A_c_93_n 0.0206882f $X=-0.19 $Y=1.66 $X2=1.475 $Y2=1.765
cc_57 VPB N_A_c_94_n 0.00764076f $X=-0.19 $Y=1.66 $X2=1.37 $Y2=1.515
cc_58 VPB N_A_c_91_n 0.0394357f $X=-0.19 $Y=1.66 $X2=1.475 $Y2=1.495
cc_59 VPB N_B_c_156_n 0.0161908f $X=-0.19 $Y=1.66 $X2=0.485 $Y2=1.225
cc_60 VPB N_B_c_157_n 0.0178234f $X=-0.19 $Y=1.66 $X2=0.915 $Y2=0.78
cc_61 VPB N_B_c_158_n 0.00416485f $X=-0.19 $Y=1.66 $X2=0.915 $Y2=1.495
cc_62 VPB B 0.00805764f $X=-0.19 $Y=1.66 $X2=1.775 $Y2=1.225
cc_63 VPB N_B_c_155_n 0.0559658f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_64 VPB N_C_c_221_n 0.0178273f $X=-0.19 $Y=1.66 $X2=0.485 $Y2=1.225
cc_65 VPB N_C_c_222_n 0.017824f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.765
cc_66 VPB N_C_c_223_n 0.00527478f $X=-0.19 $Y=1.66 $X2=0.915 $Y2=1.495
cc_67 VPB C 0.0265758f $X=-0.19 $Y=1.66 $X2=0.69 $Y2=1.565
cc_68 VPB N_C_c_220_n 0.0617585f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_69 VPB N_VPWR_c_280_n 0.0120106f $X=-0.19 $Y=1.66 $X2=1.475 $Y2=1.765
cc_70 VPB N_VPWR_c_281_n 0.0359868f $X=-0.19 $Y=1.66 $X2=1.475 $Y2=2.4
cc_71 VPB N_VPWR_c_282_n 0.00581763f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_72 VPB N_VPWR_c_283_n 0.028463f $X=-0.19 $Y=1.66 $X2=0.485 $Y2=1.495
cc_73 VPB N_VPWR_c_284_n 0.0187266f $X=-0.19 $Y=1.66 $X2=1.475 $Y2=1.495
cc_74 VPB N_VPWR_c_285_n 0.0172844f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_75 VPB N_VPWR_c_279_n 0.0796344f $X=-0.19 $Y=1.66 $X2=1.37 $Y2=1.565
cc_76 VPB N_VPWR_c_287_n 0.00614127f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_77 VPB N_VPWR_c_288_n 0.0186948f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_78 VPB N_VPWR_c_289_n 0.0421838f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_79 VPB N_VPWR_c_290_n 0.0901606f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_80 VPB N_Y_c_338_n 0.00707089f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_81 VPB N_Y_c_339_n 0.00718169f $X=-0.19 $Y=1.66 $X2=0.69 $Y2=1.515
cc_82 VPB N_Y_c_340_n 0.00257348f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_83 VPB N_Y_c_341_n 0.00249443f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_84 VPB N_Y_c_342_n 0.00257348f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_85 VPB N_Y_c_343_n 0.00437633f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_86 VPB Y 0.0128264f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_87 N_A_c_93_n N_B_c_156_n 0.0297694f $X=1.475 $Y=1.765 $X2=-0.19 $Y2=-0.245
cc_88 N_A_c_90_n N_B_M1002_g 0.0098658f $X=1.775 $Y=1.225 $X2=0 $Y2=0
cc_89 N_A_c_94_n N_B_c_153_n 0.00830118f $X=1.37 $Y=1.515 $X2=0 $Y2=0
cc_90 N_A_c_91_n N_B_c_153_n 0.00136127f $X=1.475 $Y=1.495 $X2=0 $Y2=0
cc_91 N_A_c_94_n N_B_c_155_n 0.00126944f $X=1.37 $Y=1.515 $X2=0 $Y2=0
cc_92 N_A_c_91_n N_B_c_155_n 0.02108f $X=1.475 $Y=1.495 $X2=0 $Y2=0
cc_93 N_A_c_92_n N_VPWR_c_281_n 0.0151681f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_94 N_A_c_93_n N_VPWR_c_282_n 0.0134999f $X=1.475 $Y=1.765 $X2=0 $Y2=0
cc_95 N_A_c_92_n N_VPWR_c_283_n 0.00413917f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_96 N_A_c_93_n N_VPWR_c_283_n 0.00413917f $X=1.475 $Y=1.765 $X2=0 $Y2=0
cc_97 N_A_c_92_n N_VPWR_c_279_n 0.00822528f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_98 N_A_c_93_n N_VPWR_c_279_n 0.00822528f $X=1.475 $Y=1.765 $X2=0 $Y2=0
cc_99 N_A_c_87_n N_Y_c_333_n 0.0138123f $X=0.485 $Y=1.225 $X2=0 $Y2=0
cc_100 N_A_c_94_n N_Y_c_333_n 6.95742e-19 $X=1.37 $Y=1.515 $X2=0 $Y2=0
cc_101 N_A_c_92_n N_Y_c_347_n 0.0168543f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_102 N_A_c_94_n N_Y_c_347_n 0.0054958f $X=1.37 $Y=1.515 $X2=0 $Y2=0
cc_103 N_A_c_87_n N_Y_c_349_n 0.0103239f $X=0.485 $Y=1.225 $X2=0 $Y2=0
cc_104 N_A_c_88_n N_Y_c_349_n 0.00580687f $X=0.915 $Y=1.225 $X2=0 $Y2=0
cc_105 N_A_c_89_n N_Y_c_349_n 5.7278e-19 $X=1.345 $Y=1.225 $X2=0 $Y2=0
cc_106 N_A_c_92_n N_Y_c_339_n 4.68424e-19 $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_107 N_A_c_93_n N_Y_c_339_n 4.68424e-19 $X=1.475 $Y=1.765 $X2=0 $Y2=0
cc_108 N_A_c_88_n N_Y_c_335_n 0.00900535f $X=0.915 $Y=1.225 $X2=0 $Y2=0
cc_109 N_A_c_89_n N_Y_c_335_n 0.0100844f $X=1.345 $Y=1.225 $X2=0 $Y2=0
cc_110 N_A_c_90_n N_Y_c_335_n 0.00328634f $X=1.775 $Y=1.225 $X2=0 $Y2=0
cc_111 N_A_c_94_n N_Y_c_335_n 0.0514236f $X=1.37 $Y=1.515 $X2=0 $Y2=0
cc_112 N_A_c_91_n N_Y_c_335_n 0.00722719f $X=1.475 $Y=1.495 $X2=0 $Y2=0
cc_113 N_A_c_93_n N_Y_c_359_n 0.0133118f $X=1.475 $Y=1.765 $X2=0 $Y2=0
cc_114 N_A_c_94_n N_Y_c_359_n 0.0113329f $X=1.37 $Y=1.515 $X2=0 $Y2=0
cc_115 N_A_c_91_n N_Y_c_359_n 0.00698882f $X=1.475 $Y=1.495 $X2=0 $Y2=0
cc_116 N_A_c_88_n N_Y_c_362_n 5.7278e-19 $X=0.915 $Y=1.225 $X2=0 $Y2=0
cc_117 N_A_c_89_n N_Y_c_362_n 0.00580687f $X=1.345 $Y=1.225 $X2=0 $Y2=0
cc_118 N_A_c_90_n N_Y_c_362_n 0.0046047f $X=1.775 $Y=1.225 $X2=0 $Y2=0
cc_119 N_A_c_93_n N_Y_c_340_n 6.21762e-19 $X=1.475 $Y=1.765 $X2=0 $Y2=0
cc_120 N_A_c_87_n N_Y_c_336_n 0.00107904f $X=0.485 $Y=1.225 $X2=0 $Y2=0
cc_121 N_A_c_88_n N_Y_c_336_n 0.001071f $X=0.915 $Y=1.225 $X2=0 $Y2=0
cc_122 N_A_c_94_n N_Y_c_336_n 0.027783f $X=1.37 $Y=1.515 $X2=0 $Y2=0
cc_123 N_A_c_91_n N_Y_c_336_n 0.00287341f $X=1.475 $Y=1.495 $X2=0 $Y2=0
cc_124 N_A_c_94_n N_Y_c_370_n 0.0643229f $X=1.37 $Y=1.515 $X2=0 $Y2=0
cc_125 N_A_c_91_n N_Y_c_370_n 0.00446803f $X=1.475 $Y=1.495 $X2=0 $Y2=0
cc_126 N_A_c_93_n N_Y_c_343_n 6.04745e-19 $X=1.475 $Y=1.765 $X2=0 $Y2=0
cc_127 N_A_c_87_n Y 0.0178656f $X=0.485 $Y=1.225 $X2=0 $Y2=0
cc_128 N_A_c_92_n Y 0.00699253f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_129 N_A_c_94_n Y 0.0349174f $X=1.37 $Y=1.515 $X2=0 $Y2=0
cc_130 N_A_c_91_n Y 0.00193722f $X=1.475 $Y=1.495 $X2=0 $Y2=0
cc_131 N_A_c_87_n N_A_27_82#_c_431_n 0.0124032f $X=0.485 $Y=1.225 $X2=0 $Y2=0
cc_132 N_A_c_88_n N_A_27_82#_c_431_n 0.0112468f $X=0.915 $Y=1.225 $X2=0 $Y2=0
cc_133 N_A_c_89_n N_A_27_82#_c_433_n 0.0112468f $X=1.345 $Y=1.225 $X2=0 $Y2=0
cc_134 N_A_c_90_n N_A_27_82#_c_433_n 0.0132677f $X=1.775 $Y=1.225 $X2=0 $Y2=0
cc_135 N_A_c_90_n N_A_27_82#_c_434_n 3.92031e-19 $X=1.775 $Y=1.225 $X2=0 $Y2=0
cc_136 N_A_c_87_n N_VGND_c_566_n 9.02242e-19 $X=0.485 $Y=1.225 $X2=0 $Y2=0
cc_137 N_A_c_88_n N_VGND_c_566_n 9.02242e-19 $X=0.915 $Y=1.225 $X2=0 $Y2=0
cc_138 N_A_c_89_n N_VGND_c_566_n 9.02242e-19 $X=1.345 $Y=1.225 $X2=0 $Y2=0
cc_139 N_A_c_90_n N_VGND_c_566_n 9.02242e-19 $X=1.775 $Y=1.225 $X2=0 $Y2=0
cc_140 B N_C_c_221_n 5.9621e-19 $X=3.515 $Y=1.58 $X2=-0.19 $Y2=-0.245
cc_141 B N_C_c_227_n 0.0124198f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_142 N_B_M1013_g N_C_c_220_n 0.0231295f $X=3.495 $Y=0.78 $X2=0 $Y2=0
cc_143 B N_C_c_220_n 0.00766103f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_144 N_B_c_156_n N_VPWR_c_282_n 0.00548019f $X=1.975 $Y=1.765 $X2=0 $Y2=0
cc_145 N_B_c_156_n N_VPWR_c_279_n 0.00857432f $X=1.975 $Y=1.765 $X2=0 $Y2=0
cc_146 N_B_c_157_n N_VPWR_c_279_n 0.00861697f $X=2.425 $Y=1.765 $X2=0 $Y2=0
cc_147 N_B_c_156_n N_VPWR_c_288_n 0.00445602f $X=1.975 $Y=1.765 $X2=0 $Y2=0
cc_148 N_B_c_157_n N_VPWR_c_288_n 0.00445602f $X=2.425 $Y=1.765 $X2=0 $Y2=0
cc_149 N_B_c_157_n N_VPWR_c_289_n 0.00400188f $X=2.425 $Y=1.765 $X2=0 $Y2=0
cc_150 N_B_c_156_n N_Y_c_359_n 0.0157972f $X=1.975 $Y=1.765 $X2=0 $Y2=0
cc_151 N_B_c_156_n N_Y_c_340_n 0.0108556f $X=1.975 $Y=1.765 $X2=0 $Y2=0
cc_152 N_B_c_157_n N_Y_c_340_n 0.0150947f $X=2.425 $Y=1.765 $X2=0 $Y2=0
cc_153 N_B_c_157_n N_Y_c_380_n 0.0141112f $X=2.425 $Y=1.765 $X2=0 $Y2=0
cc_154 N_B_c_158_n N_Y_c_380_n 0.0919525f $X=2.99 $Y=1.565 $X2=0 $Y2=0
cc_155 N_B_c_153_n N_Y_c_380_n 0.00498024f $X=2.56 $Y=1.565 $X2=0 $Y2=0
cc_156 N_B_c_155_n N_Y_c_380_n 0.00820729f $X=3.405 $Y=1.515 $X2=0 $Y2=0
cc_157 N_B_c_156_n N_Y_c_343_n 0.00321262f $X=1.975 $Y=1.765 $X2=0 $Y2=0
cc_158 N_B_c_157_n N_Y_c_343_n 0.00623993f $X=2.425 $Y=1.765 $X2=0 $Y2=0
cc_159 N_B_c_153_n N_Y_c_343_n 0.0179587f $X=2.56 $Y=1.565 $X2=0 $Y2=0
cc_160 N_B_c_155_n N_Y_c_343_n 0.00380406f $X=3.405 $Y=1.515 $X2=0 $Y2=0
cc_161 N_B_M1002_g N_A_27_82#_c_434_n 3.92313e-19 $X=2.205 $Y=0.78 $X2=0 $Y2=0
cc_162 N_B_c_155_n N_A_27_82#_c_434_n 0.00561102f $X=3.405 $Y=1.515 $X2=0 $Y2=0
cc_163 N_B_M1002_g N_A_27_82#_c_435_n 0.0132677f $X=2.205 $Y=0.78 $X2=0 $Y2=0
cc_164 N_B_M1003_g N_A_27_82#_c_435_n 0.0108287f $X=2.635 $Y=0.78 $X2=0 $Y2=0
cc_165 N_B_M1007_g N_A_27_82#_c_436_n 0.0108287f $X=3.065 $Y=0.78 $X2=0 $Y2=0
cc_166 N_B_M1013_g N_A_27_82#_c_436_n 0.0118941f $X=3.495 $Y=0.78 $X2=0 $Y2=0
cc_167 N_B_M1003_g N_A_456_82#_c_496_n 0.0122317f $X=2.635 $Y=0.78 $X2=0 $Y2=0
cc_168 N_B_M1007_g N_A_456_82#_c_496_n 0.0115417f $X=3.065 $Y=0.78 $X2=0 $Y2=0
cc_169 N_B_c_158_n N_A_456_82#_c_496_n 0.0390655f $X=2.99 $Y=1.565 $X2=0 $Y2=0
cc_170 N_B_c_155_n N_A_456_82#_c_496_n 0.00235612f $X=3.405 $Y=1.515 $X2=0 $Y2=0
cc_171 N_B_M1013_g N_A_456_82#_c_497_n 0.014554f $X=3.495 $Y=0.78 $X2=0 $Y2=0
cc_172 B N_A_456_82#_c_497_n 0.0205543f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_173 N_B_M1002_g N_A_456_82#_c_502_n 0.00684098f $X=2.205 $Y=0.78 $X2=0 $Y2=0
cc_174 N_B_M1003_g N_A_456_82#_c_502_n 0.00674834f $X=2.635 $Y=0.78 $X2=0 $Y2=0
cc_175 N_B_M1007_g N_A_456_82#_c_502_n 6.27882e-19 $X=3.065 $Y=0.78 $X2=0 $Y2=0
cc_176 N_B_c_153_n N_A_456_82#_c_502_n 0.0256487f $X=2.56 $Y=1.565 $X2=0 $Y2=0
cc_177 N_B_c_155_n N_A_456_82#_c_502_n 0.00269251f $X=3.405 $Y=1.515 $X2=0 $Y2=0
cc_178 N_B_M1003_g N_A_456_82#_c_503_n 6.27882e-19 $X=2.635 $Y=0.78 $X2=0 $Y2=0
cc_179 N_B_M1007_g N_A_456_82#_c_503_n 0.0067364f $X=3.065 $Y=0.78 $X2=0 $Y2=0
cc_180 N_B_M1013_g N_A_456_82#_c_503_n 0.0112821f $X=3.495 $Y=0.78 $X2=0 $Y2=0
cc_181 B N_A_456_82#_c_503_n 0.0264082f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_182 N_B_c_155_n N_A_456_82#_c_503_n 0.00240984f $X=3.405 $Y=1.515 $X2=0 $Y2=0
cc_183 N_B_M1013_g N_VGND_c_562_n 5.30949e-19 $X=3.495 $Y=0.78 $X2=0 $Y2=0
cc_184 N_B_M1002_g N_VGND_c_566_n 9.02242e-19 $X=2.205 $Y=0.78 $X2=0 $Y2=0
cc_185 N_B_M1003_g N_VGND_c_566_n 9.02242e-19 $X=2.635 $Y=0.78 $X2=0 $Y2=0
cc_186 N_B_M1007_g N_VGND_c_566_n 9.02242e-19 $X=3.065 $Y=0.78 $X2=0 $Y2=0
cc_187 N_B_M1013_g N_VGND_c_566_n 9.02242e-19 $X=3.495 $Y=0.78 $X2=0 $Y2=0
cc_188 N_C_c_221_n N_VPWR_c_284_n 0.00445602f $X=3.9 $Y=1.765 $X2=0 $Y2=0
cc_189 N_C_c_222_n N_VPWR_c_284_n 0.00445602f $X=4.35 $Y=1.765 $X2=0 $Y2=0
cc_190 N_C_c_221_n N_VPWR_c_279_n 0.00861697f $X=3.9 $Y=1.765 $X2=0 $Y2=0
cc_191 N_C_c_222_n N_VPWR_c_279_n 0.00861719f $X=4.35 $Y=1.765 $X2=0 $Y2=0
cc_192 N_C_c_221_n N_VPWR_c_289_n 0.00400188f $X=3.9 $Y=1.765 $X2=0 $Y2=0
cc_193 N_C_c_222_n N_VPWR_c_290_n 0.00399658f $X=4.35 $Y=1.765 $X2=0 $Y2=0
cc_194 N_C_c_223_n N_VPWR_c_290_n 0.112349f $X=4.935 $Y=1.56 $X2=0 $Y2=0
cc_195 N_C_c_227_n N_VPWR_c_290_n 0.00109921f $X=4.495 $Y=1.56 $X2=0 $Y2=0
cc_196 N_C_c_220_n N_VPWR_c_290_n 0.008389f $X=5.665 $Y=1.505 $X2=0 $Y2=0
cc_197 N_C_c_221_n N_Y_c_380_n 0.0160852f $X=3.9 $Y=1.765 $X2=0 $Y2=0
cc_198 N_C_c_221_n N_Y_c_341_n 0.00638955f $X=3.9 $Y=1.765 $X2=0 $Y2=0
cc_199 N_C_c_222_n N_Y_c_341_n 0.00771698f $X=4.35 $Y=1.765 $X2=0 $Y2=0
cc_200 N_C_c_227_n N_Y_c_341_n 0.0114643f $X=4.495 $Y=1.56 $X2=0 $Y2=0
cc_201 N_C_c_220_n N_Y_c_341_n 0.00849236f $X=5.665 $Y=1.505 $X2=0 $Y2=0
cc_202 N_C_c_221_n N_Y_c_342_n 0.0150947f $X=3.9 $Y=1.765 $X2=0 $Y2=0
cc_203 N_C_c_222_n N_Y_c_342_n 0.0095765f $X=4.35 $Y=1.765 $X2=0 $Y2=0
cc_204 N_C_M1000_g N_A_27_82#_c_436_n 5.80377e-19 $X=4.465 $Y=0.78 $X2=0 $Y2=0
cc_205 N_C_M1000_g N_A_456_82#_c_497_n 0.0176619f $X=4.465 $Y=0.78 $X2=0 $Y2=0
cc_206 N_C_c_227_n N_A_456_82#_c_497_n 0.033678f $X=4.495 $Y=1.56 $X2=0 $Y2=0
cc_207 N_C_c_220_n N_A_456_82#_c_497_n 0.0176385f $X=5.665 $Y=1.505 $X2=0 $Y2=0
cc_208 N_C_M1000_g N_A_456_82#_c_498_n 3.99083e-19 $X=4.465 $Y=0.78 $X2=0 $Y2=0
cc_209 N_C_M1001_g N_A_456_82#_c_498_n 3.99083e-19 $X=4.895 $Y=0.78 $X2=0 $Y2=0
cc_210 N_C_M1001_g N_A_456_82#_c_499_n 0.0145809f $X=4.895 $Y=0.78 $X2=0 $Y2=0
cc_211 N_C_M1005_g N_A_456_82#_c_499_n 0.014598f $X=5.325 $Y=0.78 $X2=0 $Y2=0
cc_212 N_C_c_223_n N_A_456_82#_c_499_n 0.0525003f $X=4.935 $Y=1.56 $X2=0 $Y2=0
cc_213 N_C_c_220_n N_A_456_82#_c_499_n 0.00226244f $X=5.665 $Y=1.505 $X2=0 $Y2=0
cc_214 C N_A_456_82#_c_500_n 0.0146264f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_215 N_C_c_220_n N_A_456_82#_c_500_n 0.00232957f $X=5.665 $Y=1.505 $X2=0 $Y2=0
cc_216 N_C_M1005_g N_A_456_82#_c_501_n 3.92313e-19 $X=5.325 $Y=0.78 $X2=0 $Y2=0
cc_217 N_C_M1008_g N_A_456_82#_c_501_n 3.92313e-19 $X=5.755 $Y=0.78 $X2=0 $Y2=0
cc_218 N_C_c_223_n N_A_456_82#_c_504_n 0.0163474f $X=4.935 $Y=1.56 $X2=0 $Y2=0
cc_219 N_C_c_220_n N_A_456_82#_c_504_n 0.00232957f $X=5.665 $Y=1.505 $X2=0 $Y2=0
cc_220 N_C_M1000_g N_VGND_c_562_n 0.00901223f $X=4.465 $Y=0.78 $X2=0 $Y2=0
cc_221 N_C_M1001_g N_VGND_c_562_n 4.25668e-19 $X=4.895 $Y=0.78 $X2=0 $Y2=0
cc_222 N_C_M1000_g N_VGND_c_563_n 4.25668e-19 $X=4.465 $Y=0.78 $X2=0 $Y2=0
cc_223 N_C_M1001_g N_VGND_c_563_n 0.00794874f $X=4.895 $Y=0.78 $X2=0 $Y2=0
cc_224 N_C_M1005_g N_VGND_c_563_n 0.00803145f $X=5.325 $Y=0.78 $X2=0 $Y2=0
cc_225 N_C_M1008_g N_VGND_c_563_n 4.31251e-19 $X=5.755 $Y=0.78 $X2=0 $Y2=0
cc_226 N_C_M1005_g N_VGND_c_565_n 5.64531e-19 $X=5.325 $Y=0.78 $X2=0 $Y2=0
cc_227 N_C_M1008_g N_VGND_c_565_n 0.0150303f $X=5.755 $Y=0.78 $X2=0 $Y2=0
cc_228 C N_VGND_c_565_n 0.0276976f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_229 N_C_M1000_g N_VGND_c_568_n 0.00455951f $X=4.465 $Y=0.78 $X2=0 $Y2=0
cc_230 N_C_M1001_g N_VGND_c_568_n 0.00455951f $X=4.895 $Y=0.78 $X2=0 $Y2=0
cc_231 N_C_M1005_g N_VGND_c_569_n 0.00455951f $X=5.325 $Y=0.78 $X2=0 $Y2=0
cc_232 N_C_M1008_g N_VGND_c_569_n 0.00455951f $X=5.755 $Y=0.78 $X2=0 $Y2=0
cc_233 N_C_M1000_g N_VGND_c_571_n 0.00447788f $X=4.465 $Y=0.78 $X2=0 $Y2=0
cc_234 N_C_M1001_g N_VGND_c_571_n 0.00447788f $X=4.895 $Y=0.78 $X2=0 $Y2=0
cc_235 N_C_M1005_g N_VGND_c_571_n 0.00447788f $X=5.325 $Y=0.78 $X2=0 $Y2=0
cc_236 N_C_M1008_g N_VGND_c_571_n 0.00447788f $X=5.755 $Y=0.78 $X2=0 $Y2=0
cc_237 N_VPWR_M1006_s N_Y_c_347_n 8.29358e-19 $X=0.135 $Y=1.84 $X2=0 $Y2=0
cc_238 N_VPWR_c_281_n N_Y_c_347_n 0.00245231f $X=0.28 $Y=2.395 $X2=0 $Y2=0
cc_239 N_VPWR_M1006_s N_Y_c_338_n 0.00350561f $X=0.135 $Y=1.84 $X2=0 $Y2=0
cc_240 N_VPWR_c_281_n N_Y_c_338_n 0.0206806f $X=0.28 $Y=2.395 $X2=0 $Y2=0
cc_241 N_VPWR_c_281_n N_Y_c_339_n 0.0267725f $X=0.28 $Y=2.395 $X2=0 $Y2=0
cc_242 N_VPWR_c_282_n N_Y_c_339_n 0.0267725f $X=1.7 $Y=2.455 $X2=0 $Y2=0
cc_243 N_VPWR_c_283_n N_Y_c_339_n 0.0333764f $X=1.535 $Y=3.33 $X2=0 $Y2=0
cc_244 N_VPWR_c_279_n N_Y_c_339_n 0.0276261f $X=6 $Y=3.33 $X2=0 $Y2=0
cc_245 N_VPWR_M1014_s N_Y_c_359_n 0.00638497f $X=1.55 $Y=1.84 $X2=0 $Y2=0
cc_246 N_VPWR_c_282_n N_Y_c_359_n 0.0202249f $X=1.7 $Y=2.455 $X2=0 $Y2=0
cc_247 N_VPWR_c_282_n N_Y_c_340_n 0.0266809f $X=1.7 $Y=2.455 $X2=0 $Y2=0
cc_248 N_VPWR_c_279_n N_Y_c_340_n 0.0119791f $X=6 $Y=3.33 $X2=0 $Y2=0
cc_249 N_VPWR_c_288_n N_Y_c_340_n 0.014552f $X=2.535 $Y=2.852 $X2=0 $Y2=0
cc_250 N_VPWR_c_289_n N_Y_c_340_n 0.0268614f $X=3.79 $Y=2.852 $X2=0 $Y2=0
cc_251 N_VPWR_M1016_s N_Y_c_380_n 0.0339419f $X=2.5 $Y=1.84 $X2=0 $Y2=0
cc_252 N_VPWR_c_289_n N_Y_c_380_n 0.0980931f $X=3.79 $Y=2.852 $X2=0 $Y2=0
cc_253 N_VPWR_c_284_n N_Y_c_342_n 0.014552f $X=4.46 $Y=3.33 $X2=0 $Y2=0
cc_254 N_VPWR_c_279_n N_Y_c_342_n 0.0119791f $X=6 $Y=3.33 $X2=0 $Y2=0
cc_255 N_VPWR_c_289_n N_Y_c_342_n 0.0268614f $X=3.79 $Y=2.852 $X2=0 $Y2=0
cc_256 N_VPWR_c_290_n N_Y_c_342_n 0.0331138f $X=4.92 $Y=2.115 $X2=0 $Y2=0
cc_257 N_VPWR_M1006_s Y 0.00194313f $X=0.135 $Y=1.84 $X2=0 $Y2=0
cc_258 N_Y_c_334_n N_A_27_82#_M1004_s 0.00267822f $X=0.355 $Y=1.095 $X2=-0.19
+ $Y2=-0.245
cc_259 N_Y_c_335_n N_A_27_82#_M1009_s 0.00176461f $X=1.395 $Y=1.095 $X2=0 $Y2=0
cc_260 N_Y_c_334_n N_A_27_82#_c_430_n 0.0204519f $X=0.355 $Y=1.095 $X2=0 $Y2=0
cc_261 N_Y_M1004_d N_A_27_82#_c_431_n 0.00176461f $X=0.56 $Y=0.41 $X2=0 $Y2=0
cc_262 N_Y_c_333_n N_A_27_82#_c_431_n 0.0030313f $X=0.535 $Y=1.095 $X2=0 $Y2=0
cc_263 N_Y_c_349_n N_A_27_82#_c_431_n 0.0157965f $X=0.7 $Y=0.68 $X2=0 $Y2=0
cc_264 N_Y_c_335_n N_A_27_82#_c_431_n 0.0030313f $X=1.395 $Y=1.095 $X2=0 $Y2=0
cc_265 N_Y_c_335_n N_A_27_82#_c_460_n 0.0133411f $X=1.395 $Y=1.095 $X2=0 $Y2=0
cc_266 N_Y_M1010_d N_A_27_82#_c_433_n 0.00176461f $X=1.42 $Y=0.41 $X2=0 $Y2=0
cc_267 N_Y_c_335_n N_A_27_82#_c_433_n 0.0030313f $X=1.395 $Y=1.095 $X2=0 $Y2=0
cc_268 N_Y_c_362_n N_A_27_82#_c_433_n 0.0157965f $X=1.56 $Y=0.68 $X2=0 $Y2=0
cc_269 N_Y_c_335_n N_A_27_82#_c_434_n 0.00712541f $X=1.395 $Y=1.095 $X2=0 $Y2=0
cc_270 N_Y_c_343_n N_A_27_82#_c_434_n 0.00135473f $X=2.2 $Y=1.985 $X2=0 $Y2=0
cc_271 N_Y_c_341_n N_A_456_82#_c_497_n 0.00594674f $X=4.125 $Y=2.12 $X2=0 $Y2=0
cc_272 N_A_27_82#_c_435_n N_A_456_82#_M1002_s 0.00176461f $X=2.755 $Y=0.34
+ $X2=-0.19 $Y2=-0.245
cc_273 N_A_27_82#_c_436_n N_A_456_82#_M1007_s 0.00176461f $X=3.615 $Y=0.34 $X2=0
+ $Y2=0
cc_274 N_A_27_82#_M1003_d N_A_456_82#_c_496_n 0.00178571f $X=2.71 $Y=0.41 $X2=0
+ $Y2=0
cc_275 N_A_27_82#_c_435_n N_A_456_82#_c_496_n 0.00364066f $X=2.755 $Y=0.34 $X2=0
+ $Y2=0
cc_276 N_A_27_82#_c_470_p N_A_456_82#_c_496_n 0.0135228f $X=2.85 $Y=0.57 $X2=0
+ $Y2=0
cc_277 N_A_27_82#_c_436_n N_A_456_82#_c_496_n 0.00364066f $X=3.615 $Y=0.34 $X2=0
+ $Y2=0
cc_278 N_A_27_82#_M1013_d N_A_456_82#_c_497_n 0.00296342f $X=3.57 $Y=0.41 $X2=0
+ $Y2=0
cc_279 N_A_27_82#_c_436_n N_A_456_82#_c_497_n 0.00364066f $X=3.615 $Y=0.34 $X2=0
+ $Y2=0
cc_280 N_A_27_82#_c_437_n N_A_456_82#_c_497_n 0.0202474f $X=3.71 $Y=0.57 $X2=0
+ $Y2=0
cc_281 N_A_27_82#_c_434_n N_A_456_82#_c_502_n 0.0212953f $X=1.99 $Y=0.555 $X2=0
+ $Y2=0
cc_282 N_A_27_82#_c_435_n N_A_456_82#_c_502_n 0.0157757f $X=2.755 $Y=0.34 $X2=0
+ $Y2=0
cc_283 N_A_27_82#_c_436_n N_A_456_82#_c_503_n 0.0157757f $X=3.615 $Y=0.34 $X2=0
+ $Y2=0
cc_284 N_A_27_82#_c_436_n N_VGND_c_562_n 0.0129575f $X=3.615 $Y=0.34 $X2=0 $Y2=0
cc_285 N_A_27_82#_c_437_n N_VGND_c_562_n 0.0228893f $X=3.71 $Y=0.57 $X2=0 $Y2=0
cc_286 N_A_27_82#_c_431_n N_VGND_c_566_n 0.0443903f $X=1.045 $Y=0.34 $X2=0 $Y2=0
cc_287 N_A_27_82#_c_432_n N_VGND_c_566_n 0.0177208f $X=0.355 $Y=0.34 $X2=0 $Y2=0
cc_288 N_A_27_82#_c_433_n N_VGND_c_566_n 0.0443903f $X=1.905 $Y=0.34 $X2=0 $Y2=0
cc_289 N_A_27_82#_c_435_n N_VGND_c_566_n 0.0437462f $X=2.755 $Y=0.34 $X2=0 $Y2=0
cc_290 N_A_27_82#_c_436_n N_VGND_c_566_n 0.061305f $X=3.615 $Y=0.34 $X2=0 $Y2=0
cc_291 N_A_27_82#_c_438_n N_VGND_c_566_n 0.0120507f $X=1.13 $Y=0.34 $X2=0 $Y2=0
cc_292 N_A_27_82#_c_439_n N_VGND_c_566_n 0.0121867f $X=1.99 $Y=0.34 $X2=0 $Y2=0
cc_293 N_A_27_82#_c_440_n N_VGND_c_566_n 0.0133031f $X=2.85 $Y=0.34 $X2=0 $Y2=0
cc_294 N_A_27_82#_c_431_n N_VGND_c_571_n 0.0259344f $X=1.045 $Y=0.34 $X2=0 $Y2=0
cc_295 N_A_27_82#_c_432_n N_VGND_c_571_n 0.00968164f $X=0.355 $Y=0.34 $X2=0
+ $Y2=0
cc_296 N_A_27_82#_c_433_n N_VGND_c_571_n 0.0259344f $X=1.905 $Y=0.34 $X2=0 $Y2=0
cc_297 N_A_27_82#_c_435_n N_VGND_c_571_n 0.0255585f $X=2.755 $Y=0.34 $X2=0 $Y2=0
cc_298 N_A_27_82#_c_436_n N_VGND_c_571_n 0.0352091f $X=3.615 $Y=0.34 $X2=0 $Y2=0
cc_299 N_A_27_82#_c_438_n N_VGND_c_571_n 0.00658361f $X=1.13 $Y=0.34 $X2=0 $Y2=0
cc_300 N_A_27_82#_c_439_n N_VGND_c_571_n 0.00660921f $X=1.99 $Y=0.34 $X2=0 $Y2=0
cc_301 N_A_27_82#_c_440_n N_VGND_c_571_n 0.00732729f $X=2.85 $Y=0.34 $X2=0 $Y2=0
cc_302 N_A_456_82#_c_497_n N_VGND_M1000_s 0.00354923f $X=4.585 $Y=1.045
+ $X2=-0.19 $Y2=-0.245
cc_303 N_A_456_82#_c_499_n N_VGND_M1001_s 0.00178571f $X=5.455 $Y=1.045 $X2=0
+ $Y2=0
cc_304 N_A_456_82#_c_497_n N_VGND_c_562_n 0.0225605f $X=4.585 $Y=1.045 $X2=0
+ $Y2=0
cc_305 N_A_456_82#_c_498_n N_VGND_c_562_n 0.0142351f $X=4.68 $Y=0.555 $X2=0
+ $Y2=0
cc_306 N_A_456_82#_c_498_n N_VGND_c_563_n 0.0142351f $X=4.68 $Y=0.555 $X2=0
+ $Y2=0
cc_307 N_A_456_82#_c_499_n N_VGND_c_563_n 0.0175375f $X=5.455 $Y=1.045 $X2=0
+ $Y2=0
cc_308 N_A_456_82#_c_501_n N_VGND_c_563_n 0.0135894f $X=5.54 $Y=0.555 $X2=0
+ $Y2=0
cc_309 N_A_456_82#_c_500_n N_VGND_c_565_n 0.00985092f $X=5.54 $Y=0.92 $X2=0
+ $Y2=0
cc_310 N_A_456_82#_c_501_n N_VGND_c_565_n 0.0196825f $X=5.54 $Y=0.555 $X2=0
+ $Y2=0
cc_311 N_A_456_82#_c_498_n N_VGND_c_568_n 0.00722494f $X=4.68 $Y=0.555 $X2=0
+ $Y2=0
cc_312 N_A_456_82#_c_501_n N_VGND_c_569_n 0.00645633f $X=5.54 $Y=0.555 $X2=0
+ $Y2=0
cc_313 N_A_456_82#_c_498_n N_VGND_c_571_n 0.00677346f $X=4.68 $Y=0.555 $X2=0
+ $Y2=0
cc_314 N_A_456_82#_c_501_n N_VGND_c_571_n 0.00605288f $X=5.54 $Y=0.555 $X2=0
+ $Y2=0
