# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_hs__dfrbp_1
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_hs__dfrbp_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  11.52000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.000000 0.520000 2.195000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.541300 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 11.065000 0.350000 11.435000 1.130000 ;
        RECT 11.075000 1.820000 11.435000 2.980000 ;
        RECT 11.265000 1.130000 11.435000 1.820000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.951500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 9.260000 1.810000 9.950000 2.985000 ;
        RECT 9.560000 0.350000 9.950000 1.810000 ;
    END
  END Q_N
  PIN RESET_B
    ANTENNAGATEAREA  0.378000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.030000 1.130000 1.300000 2.140000 ;
        RECT 5.230000 1.825000 5.610000 2.155000 ;
        RECT 7.835000 1.835000 8.300000 2.165000 ;
      LAYER mcon ;
        RECT 1.115000 1.950000 1.285000 2.120000 ;
        RECT 5.435000 1.950000 5.605000 2.120000 ;
        RECT 7.835000 1.950000 8.005000 2.120000 ;
      LAYER met1 ;
        RECT 1.055000 1.920000 1.345000 1.965000 ;
        RECT 1.055000 1.965000 8.065000 2.105000 ;
        RECT 1.055000 2.105000 1.345000 2.150000 ;
        RECT 5.375000 1.920000 5.665000 1.965000 ;
        RECT 5.375000 2.105000 5.665000 2.150000 ;
        RECT 7.775000 1.920000 8.065000 1.965000 ;
        RECT 7.775000 2.105000 8.065000 2.150000 ;
    END
  END RESET_B
  PIN CLK
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 1.810000 1.310000 2.275000 1.640000 ;
        RECT 2.045000 1.640000 2.275000 1.780000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT  0.000000 -0.085000 11.520000 0.085000 ;
        RECT  1.030000  0.085000  1.280000 0.830000 ;
        RECT  2.090000  0.085000  2.420000 0.800000 ;
        RECT  4.995000  0.085000  5.325000 0.410000 ;
        RECT  7.535000  0.085000  7.995000 0.680000 ;
        RECT  9.140000  0.085000  9.390000 1.130000 ;
        RECT 10.645000  0.085000 10.895000 1.130000 ;
      LAYER mcon ;
        RECT  0.155000 -0.085000  0.325000 0.085000 ;
        RECT  0.635000 -0.085000  0.805000 0.085000 ;
        RECT  1.115000 -0.085000  1.285000 0.085000 ;
        RECT  1.595000 -0.085000  1.765000 0.085000 ;
        RECT  2.075000 -0.085000  2.245000 0.085000 ;
        RECT  2.555000 -0.085000  2.725000 0.085000 ;
        RECT  3.035000 -0.085000  3.205000 0.085000 ;
        RECT  3.515000 -0.085000  3.685000 0.085000 ;
        RECT  3.995000 -0.085000  4.165000 0.085000 ;
        RECT  4.475000 -0.085000  4.645000 0.085000 ;
        RECT  4.955000 -0.085000  5.125000 0.085000 ;
        RECT  5.435000 -0.085000  5.605000 0.085000 ;
        RECT  5.915000 -0.085000  6.085000 0.085000 ;
        RECT  6.395000 -0.085000  6.565000 0.085000 ;
        RECT  6.875000 -0.085000  7.045000 0.085000 ;
        RECT  7.355000 -0.085000  7.525000 0.085000 ;
        RECT  7.835000 -0.085000  8.005000 0.085000 ;
        RECT  8.315000 -0.085000  8.485000 0.085000 ;
        RECT  8.795000 -0.085000  8.965000 0.085000 ;
        RECT  9.275000 -0.085000  9.445000 0.085000 ;
        RECT  9.755000 -0.085000  9.925000 0.085000 ;
        RECT 10.235000 -0.085000 10.405000 0.085000 ;
        RECT 10.715000 -0.085000 10.885000 0.085000 ;
        RECT 11.195000 -0.085000 11.365000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.245000 11.520000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT  0.000000 3.245000 11.520000 3.415000 ;
        RECT  0.115000 2.520000  0.365000 3.245000 ;
        RECT  1.095000 2.650000  1.345000 3.245000 ;
        RECT  2.025000 2.650000  2.355000 3.245000 ;
        RECT  4.440000 2.755000  4.785000 3.245000 ;
        RECT  5.780000 1.740000  6.030000 3.245000 ;
        RECT  7.835000 2.335000  8.060000 3.245000 ;
        RECT  8.810000 2.105000  9.025000 3.245000 ;
        RECT 10.610000 1.820000 10.905000 3.245000 ;
      LAYER mcon ;
        RECT  0.155000 3.245000  0.325000 3.415000 ;
        RECT  0.635000 3.245000  0.805000 3.415000 ;
        RECT  1.115000 3.245000  1.285000 3.415000 ;
        RECT  1.595000 3.245000  1.765000 3.415000 ;
        RECT  2.075000 3.245000  2.245000 3.415000 ;
        RECT  2.555000 3.245000  2.725000 3.415000 ;
        RECT  3.035000 3.245000  3.205000 3.415000 ;
        RECT  3.515000 3.245000  3.685000 3.415000 ;
        RECT  3.995000 3.245000  4.165000 3.415000 ;
        RECT  4.475000 3.245000  4.645000 3.415000 ;
        RECT  4.955000 3.245000  5.125000 3.415000 ;
        RECT  5.435000 3.245000  5.605000 3.415000 ;
        RECT  5.915000 3.245000  6.085000 3.415000 ;
        RECT  6.395000 3.245000  6.565000 3.415000 ;
        RECT  6.875000 3.245000  7.045000 3.415000 ;
        RECT  7.355000 3.245000  7.525000 3.415000 ;
        RECT  7.835000 3.245000  8.005000 3.415000 ;
        RECT  8.315000 3.245000  8.485000 3.415000 ;
        RECT  8.795000 3.245000  8.965000 3.415000 ;
        RECT  9.275000 3.245000  9.445000 3.415000 ;
        RECT  9.755000 3.245000  9.925000 3.415000 ;
        RECT 10.235000 3.245000 10.405000 3.415000 ;
        RECT 10.715000 3.245000 10.885000 3.415000 ;
        RECT 11.195000 3.245000 11.365000 3.415000 ;
      LAYER met1 ;
        RECT 0.000000 3.085000 11.520000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.170000 0.370000  0.500000 0.660000 ;
      RECT  0.170000 0.660000  0.860000 0.830000 ;
      RECT  0.565000 2.520000  0.895000 2.980000 ;
      RECT  0.690000 0.830000  0.860000 2.310000 ;
      RECT  0.690000 2.310000  3.395000 2.480000 ;
      RECT  0.690000 2.480000  0.895000 2.520000 ;
      RECT  1.470000 0.350000  1.920000 0.970000 ;
      RECT  1.470000 0.970000  2.775000 1.140000 ;
      RECT  1.470000 1.140000  1.640000 1.810000 ;
      RECT  1.470000 1.810000  1.825000 2.140000 ;
      RECT  2.445000 1.140000  2.775000 1.550000 ;
      RECT  2.475000 1.735000  3.500000 1.905000 ;
      RECT  2.475000 1.905000  2.805000 2.140000 ;
      RECT  2.590000 0.255000  4.520000 0.425000 ;
      RECT  2.590000 0.425000  3.115000 0.800000 ;
      RECT  2.945000 0.800000  3.115000 1.575000 ;
      RECT  2.945000 1.575000  3.500000 1.735000 ;
      RECT  3.065000 2.075000  3.840000 2.245000 ;
      RECT  3.065000 2.245000  3.395000 2.310000 ;
      RECT  3.065000 2.480000  3.395000 2.755000 ;
      RECT  3.285000 0.595000  3.535000 1.200000 ;
      RECT  3.285000 1.200000  3.840000 1.370000 ;
      RECT  3.595000 2.415000  5.325000 2.585000 ;
      RECT  3.595000 2.585000  3.845000 2.755000 ;
      RECT  3.670000 1.370000  3.840000 2.075000 ;
      RECT  3.705000 0.595000  4.180000 1.030000 ;
      RECT  4.010000 1.030000  4.180000 2.415000 ;
      RECT  4.350000 0.425000  4.520000 0.580000 ;
      RECT  4.350000 0.580000  6.255000 0.750000 ;
      RECT  4.350000 0.920000  5.915000 1.090000 ;
      RECT  4.350000 1.090000  4.630000 2.155000 ;
      RECT  4.890000 1.445000  5.560000 1.615000 ;
      RECT  4.890000 1.615000  5.060000 2.350000 ;
      RECT  4.890000 2.350000  5.325000 2.415000 ;
      RECT  4.990000 2.585000  5.325000 2.680000 ;
      RECT  5.230000 1.285000  5.560000 1.445000 ;
      RECT  5.745000 1.090000  5.915000 1.400000 ;
      RECT  5.745000 1.400000  6.480000 1.570000 ;
      RECT  6.085000 0.750000  6.255000 0.900000 ;
      RECT  6.085000 0.900000  6.820000 1.230000 ;
      RECT  6.230000 1.570000  6.480000 2.755000 ;
      RECT  6.425000 0.400000  7.160000 0.730000 ;
      RECT  6.650000 1.230000  6.820000 1.865000 ;
      RECT  6.650000 1.865000  7.325000 2.195000 ;
      RECT  6.700000 2.365000  7.665000 2.695000 ;
      RECT  6.990000 0.730000  7.160000 1.425000 ;
      RECT  6.990000 1.425000  8.630000 1.595000 ;
      RECT  7.430000 0.900000  8.970000 1.070000 ;
      RECT  7.430000 1.070000  7.760000 1.230000 ;
      RECT  7.495000 1.595000  7.665000 2.365000 ;
      RECT  8.260000 2.335000  8.640000 2.730000 ;
      RECT  8.330000 1.265000  8.630000 1.425000 ;
      RECT  8.470000 1.765000  8.970000 1.935000 ;
      RECT  8.470000 1.935000  8.640000 2.335000 ;
      RECT  8.485000 0.350000  8.970000 0.900000 ;
      RECT  8.800000 1.070000  8.970000 1.765000 ;
      RECT 10.190000 0.350000 10.440000 1.300000 ;
      RECT 10.190000 1.300000 11.095000 1.630000 ;
      RECT 10.190000 1.630000 10.440000 2.975000 ;
  END
END sky130_fd_sc_hs__dfrbp_1
