* NGSPICE file created from sky130_fd_sc_hs__o32ai_1.ext - technology: sky130A

.subckt sky130_fd_sc_hs__o32ai_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
M1000 a_128_368# B1 VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=3.024e+11p pd=2.78e+06u as=7.056e+11p ps=5.74e+06u
M1001 a_342_368# A3 Y VPB pshort w=1.12e+06u l=150000u
+  ad=4.704e+11p pd=3.08e+06u as=5.6e+11p ps=3.24e+06u
M1002 VPWR A1 a_456_368# VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=4.704e+11p ps=3.08e+06u
M1003 VGND A3 a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=5.439e+11p pd=4.43e+06u as=6.771e+11p ps=6.27e+06u
M1004 VGND A1 a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 Y B2 a_128_368# VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_27_74# B2 Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=4.329e+11p ps=2.65e+06u
M1007 a_27_74# A2 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 Y B1 a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_456_368# A2 a_342_368# VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

