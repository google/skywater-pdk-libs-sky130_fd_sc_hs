* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hs__dlxtp_1 D GATE VGND VNB VPB VPWR Q
X0 a_592_149# a_685_59# a_239_85# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X1 VGND a_386_326# a_514_149# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X2 a_229_392# a_562_123# a_592_149# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=150000u
X3 VGND D a_116_424# VNB sky130_fd_pr__nfet_01v8_lvt w=550000u l=150000u
X4 VGND a_386_326# Q VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X5 a_562_123# GATE VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X6 a_239_85# a_116_424# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X7 VPWR a_386_326# Q VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X8 a_386_326# a_592_149# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X9 a_229_392# a_116_424# VPWR VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=150000u
X10 VPWR a_386_326# a_419_392# VPB sky130_fd_pr__pfet_01v8 w=420000u l=150000u
X11 a_592_149# a_685_59# a_419_392# VPB sky130_fd_pr__pfet_01v8 w=420000u l=150000u
X12 a_386_326# a_592_149# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X13 a_514_149# a_562_123# a_592_149# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X14 a_562_123# GATE VPWR VPB sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X15 VPWR D a_116_424# VPB sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X16 VGND a_562_123# a_685_59# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X17 VPWR a_562_123# a_685_59# VPB sky130_fd_pr__pfet_01v8 w=840000u l=150000u
.ends
