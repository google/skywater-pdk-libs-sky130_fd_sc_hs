* File: sky130_fd_sc_hs__nor4b_2.pex.spice
* Created: Tue Sep  1 20:12:27 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HS__NOR4B_2%D_N 1 3 6 8
c32 8 0 1.74586e-19 $X=0.72 $Y=1.665
r33 8 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.7
+ $Y=1.635 $X2=0.7 $Y2=1.635
r34 4 11 39.4698 $w=3.94e-07 $l=1.69926e-07 $layer=POLY_cond $X=0.63 $Y=1.47
+ $X2=0.64 $Y2=1.635
r35 4 6 399.957 $w=1.5e-07 $l=7.8e-07 $layer=POLY_cond $X=0.63 $Y=1.47 $X2=0.63
+ $Y2=0.69
r36 1 11 49.8683 $w=3.94e-07 $l=3.10242e-07 $layer=POLY_cond $X=0.505 $Y=1.885
+ $X2=0.64 $Y2=1.635
r37 1 3 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=0.505 $Y=1.885
+ $X2=0.505 $Y2=2.46
.ends

.subckt PM_SKY130_FD_SC_HS__NOR4B_2%A_27_392# 1 2 7 9 10 12 13 15 16 18 21 25 31
+ 33 35 40
c86 33 0 1.17824e-19 $X=1.61 $Y=1.385
c87 16 0 1.86416e-19 $X=1.965 $Y=1.765
c88 10 0 1.74586e-19 $X=1.515 $Y=1.765
r89 40 41 31.0779 $w=4.11e-07 $l=2.65e-07 $layer=POLY_cond $X=1.7 $Y=1.492
+ $X2=1.965 $Y2=1.492
r90 37 38 36.9416 $w=4.11e-07 $l=3.15e-07 $layer=POLY_cond $X=1.2 $Y=1.492
+ $X2=1.515 $Y2=1.492
r91 34 40 10.5547 $w=4.11e-07 $l=9e-08 $layer=POLY_cond $X=1.61 $Y=1.492 $X2=1.7
+ $Y2=1.492
r92 34 38 11.1411 $w=4.11e-07 $l=9.5e-08 $layer=POLY_cond $X=1.61 $Y=1.492
+ $X2=1.515 $Y2=1.492
r93 33 35 18.0659 $w=4.18e-07 $l=5.05e-07 $layer=LI1_cond $X=1.61 $Y=1.34
+ $X2=1.105 $Y2=1.34
r94 33 34 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.61
+ $Y=1.385 $X2=1.61 $Y2=1.385
r95 30 31 4.11427 $w=1.7e-07 $l=2.33e-07 $layer=LI1_cond $X=0.58 $Y=1.215
+ $X2=0.347 $Y2=1.215
r96 30 35 34.2513 $w=1.68e-07 $l=5.25e-07 $layer=LI1_cond $X=0.58 $Y=1.215
+ $X2=1.105 $Y2=1.215
r97 25 27 32.7294 $w=2.48e-07 $l=7.1e-07 $layer=LI1_cond $X=0.24 $Y=2.105
+ $X2=0.24 $Y2=2.815
r98 23 31 2.68319 $w=3.57e-07 $l=1.43332e-07 $layer=LI1_cond $X=0.24 $Y=1.3
+ $X2=0.347 $Y2=1.215
r99 23 25 37.1087 $w=2.48e-07 $l=8.05e-07 $layer=LI1_cond $X=0.24 $Y=1.3
+ $X2=0.24 $Y2=2.105
r100 19 31 2.68319 $w=3.57e-07 $l=8.5e-08 $layer=LI1_cond $X=0.347 $Y=1.13
+ $X2=0.347 $Y2=1.215
r101 19 21 15.8191 $w=4.63e-07 $l=6.15e-07 $layer=LI1_cond $X=0.347 $Y=1.13
+ $X2=0.347 $Y2=0.515
r102 16 41 26.5265 $w=1.5e-07 $l=2.73e-07 $layer=POLY_cond $X=1.965 $Y=1.765
+ $X2=1.965 $Y2=1.492
r103 16 18 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.965 $Y=1.765
+ $X2=1.965 $Y2=2.4
r104 13 40 26.5265 $w=1.5e-07 $l=2.72e-07 $layer=POLY_cond $X=1.7 $Y=1.22
+ $X2=1.7 $Y2=1.492
r105 13 15 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.7 $Y=1.22 $X2=1.7
+ $Y2=0.74
r106 10 38 26.5265 $w=1.5e-07 $l=2.73e-07 $layer=POLY_cond $X=1.515 $Y=1.765
+ $X2=1.515 $Y2=1.492
r107 10 12 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.515 $Y=1.765
+ $X2=1.515 $Y2=2.4
r108 7 37 26.5265 $w=1.5e-07 $l=2.72e-07 $layer=POLY_cond $X=1.2 $Y=1.22 $X2=1.2
+ $Y2=1.492
r109 7 9 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.2 $Y=1.22 $X2=1.2
+ $Y2=0.74
r110 2 27 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.96 $X2=0.28 $Y2=2.815
r111 2 25 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.96 $X2=0.28 $Y2=2.105
r112 1 21 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.27
+ $Y=0.37 $X2=0.415 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__NOR4B_2%C 3 5 7 10 12 14 15 16 24
c56 24 0 1.53909e-19 $X=2.82 $Y=1.557
c57 12 0 7.48116e-20 $X=2.865 $Y=1.765
c58 5 0 7.17547e-20 $X=2.415 $Y=1.765
r59 24 25 5.75332 $w=3.77e-07 $l=4.5e-08 $layer=POLY_cond $X=2.82 $Y=1.557
+ $X2=2.865 $Y2=1.557
r60 22 24 43.4695 $w=3.77e-07 $l=3.4e-07 $layer=POLY_cond $X=2.48 $Y=1.557
+ $X2=2.82 $Y2=1.557
r61 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.48
+ $Y=1.515 $X2=2.48 $Y2=1.515
r62 20 22 8.31034 $w=3.77e-07 $l=6.5e-08 $layer=POLY_cond $X=2.415 $Y=1.557
+ $X2=2.48 $Y2=1.557
r63 19 20 3.19629 $w=3.77e-07 $l=2.5e-08 $layer=POLY_cond $X=2.39 $Y=1.557
+ $X2=2.415 $Y2=1.557
r64 16 23 4.28816 $w=4.28e-07 $l=1.6e-07 $layer=LI1_cond $X=2.64 $Y=1.565
+ $X2=2.48 $Y2=1.565
r65 15 23 8.57632 $w=4.28e-07 $l=3.2e-07 $layer=LI1_cond $X=2.16 $Y=1.565
+ $X2=2.48 $Y2=1.565
r66 12 25 24.4204 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=2.865 $Y=1.765
+ $X2=2.865 $Y2=1.557
r67 12 14 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.865 $Y=1.765
+ $X2=2.865 $Y2=2.4
r68 8 24 24.4204 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.82 $Y=1.35
+ $X2=2.82 $Y2=1.557
r69 8 10 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.82 $Y=1.35 $X2=2.82
+ $Y2=0.74
r70 5 20 24.4204 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=2.415 $Y=1.765
+ $X2=2.415 $Y2=1.557
r71 5 7 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.415 $Y=1.765
+ $X2=2.415 $Y2=2.4
r72 1 19 24.4204 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.39 $Y=1.35
+ $X2=2.39 $Y2=1.557
r73 1 3 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.39 $Y=1.35 $X2=2.39
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HS__NOR4B_2%B 3 5 6 7 9 12 14 16 18 19 21 22 26
c63 22 0 7.48116e-20 $X=4.08 $Y=1.665
c64 16 0 1.37443e-19 $X=4.325 $Y=1.765
c65 5 0 1.87881e-19 $X=3.785 $Y=1.515
r66 26 27 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.8
+ $Y=1.515 $X2=3.8 $Y2=1.515
r67 22 27 7.50428 $w=4.28e-07 $l=2.8e-07 $layer=LI1_cond $X=4.08 $Y=1.565
+ $X2=3.8 $Y2=1.565
r68 21 27 5.3602 $w=4.28e-07 $l=2e-07 $layer=LI1_cond $X=3.6 $Y=1.565 $X2=3.8
+ $Y2=1.565
r69 16 19 64.3434 $w=1.8e-07 $l=1.6e-07 $layer=POLY_cond $X=4.325 $Y=1.765
+ $X2=4.325 $Y2=1.605
r70 16 18 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=4.325 $Y=1.765
+ $X2=4.325 $Y2=2.4
r71 15 26 6.91837 $w=1.5e-07 $l=1.11445e-07 $layer=POLY_cond $X=3.965 $Y=1.605
+ $X2=3.875 $Y2=1.557
r72 14 19 7.1379 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=4.235 $Y=1.605
+ $X2=4.325 $Y2=1.605
r73 14 15 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=4.235 $Y=1.605
+ $X2=3.965 $Y2=1.605
r74 10 26 18.1359 $w=1.5e-07 $l=2.14369e-07 $layer=POLY_cond $X=3.89 $Y=1.35
+ $X2=3.875 $Y2=1.557
r75 10 12 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=3.89 $Y=1.35
+ $X2=3.89 $Y2=0.74
r76 7 26 18.1359 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=3.875 $Y=1.765
+ $X2=3.875 $Y2=1.557
r77 7 9 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.875 $Y=1.765
+ $X2=3.875 $Y2=2.4
r78 5 26 6.91837 $w=3.3e-07 $l=1.08995e-07 $layer=POLY_cond $X=3.785 $Y=1.515
+ $X2=3.875 $Y2=1.557
r79 5 6 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=3.785 $Y=1.515
+ $X2=3.445 $Y2=1.515
r80 1 6 32.1775 $w=3.3e-07 $l=1.98997e-07 $layer=POLY_cond $X=3.37 $Y=1.35
+ $X2=3.445 $Y2=1.515
r81 1 3 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=3.37 $Y=1.35 $X2=3.37
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HS__NOR4B_2%A 3 5 7 8 10 13 15 16 17 26
c45 17 0 1.37443e-19 $X=5.52 $Y=1.665
r46 26 27 1.928 $w=3.75e-07 $l=1.5e-08 $layer=POLY_cond $X=5.235 $Y=1.557
+ $X2=5.25 $Y2=1.557
r47 24 26 9.64 $w=3.75e-07 $l=7.5e-08 $layer=POLY_cond $X=5.16 $Y=1.557
+ $X2=5.235 $Y2=1.557
r48 24 25 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.16
+ $Y=1.515 $X2=5.16 $Y2=1.515
r49 22 24 49.4853 $w=3.75e-07 $l=3.85e-07 $layer=POLY_cond $X=4.775 $Y=1.557
+ $X2=5.16 $Y2=1.557
r50 21 22 1.28533 $w=3.75e-07 $l=1e-08 $layer=POLY_cond $X=4.765 $Y=1.557
+ $X2=4.775 $Y2=1.557
r51 17 25 9.64836 $w=4.28e-07 $l=3.6e-07 $layer=LI1_cond $X=5.52 $Y=1.565
+ $X2=5.16 $Y2=1.565
r52 16 25 3.21612 $w=4.28e-07 $l=1.2e-07 $layer=LI1_cond $X=5.04 $Y=1.565
+ $X2=5.16 $Y2=1.565
r53 15 16 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=4.56 $Y=1.565
+ $X2=5.04 $Y2=1.565
r54 11 27 24.2915 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=5.25 $Y=1.35
+ $X2=5.25 $Y2=1.557
r55 11 13 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=5.25 $Y=1.35
+ $X2=5.25 $Y2=0.74
r56 8 26 24.2915 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=5.235 $Y=1.765
+ $X2=5.235 $Y2=1.557
r57 8 10 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=5.235 $Y=1.765
+ $X2=5.235 $Y2=2.4
r58 5 22 24.2915 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=4.775 $Y=1.765
+ $X2=4.775 $Y2=1.557
r59 5 7 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=4.775 $Y=1.765
+ $X2=4.775 $Y2=2.4
r60 1 21 24.2915 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.765 $Y=1.35
+ $X2=4.765 $Y2=1.557
r61 1 3 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=4.765 $Y=1.35
+ $X2=4.765 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HS__NOR4B_2%VPWR 1 2 9 15 17 19 24 34 35 38 41
r56 41 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r57 38 39 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r58 35 42 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=5.04 $Y2=3.33
r59 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r60 32 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.165 $Y=3.33 $X2=5
+ $Y2=3.33
r61 32 34 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=5.165 $Y=3.33
+ $X2=5.52 $Y2=3.33
r62 31 42 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=5.04 $Y2=3.33
r63 30 31 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r64 28 39 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r65 27 30 219.209 $w=1.68e-07 $l=3.36e-06 $layer=LI1_cond $X=1.2 $Y=3.33
+ $X2=4.56 $Y2=3.33
r66 27 28 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r67 25 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.895 $Y=3.33
+ $X2=0.73 $Y2=3.33
r68 25 27 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.895 $Y=3.33
+ $X2=1.2 $Y2=3.33
r69 24 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.835 $Y=3.33 $X2=5
+ $Y2=3.33
r70 24 30 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=4.835 $Y=3.33
+ $X2=4.56 $Y2=3.33
r71 22 39 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r72 21 22 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r73 19 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.565 $Y=3.33
+ $X2=0.73 $Y2=3.33
r74 19 21 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.565 $Y=3.33
+ $X2=0.24 $Y2=3.33
r75 17 31 0.468274 $w=4.9e-07 $l=1.68e-06 $layer=MET1_cond $X=2.88 $Y=3.33
+ $X2=4.56 $Y2=3.33
r76 17 28 0.468274 $w=4.9e-07 $l=1.68e-06 $layer=MET1_cond $X=2.88 $Y=3.33
+ $X2=1.2 $Y2=3.33
r77 13 41 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5 $Y=3.245 $X2=5
+ $Y2=3.33
r78 13 15 27.5888 $w=3.28e-07 $l=7.9e-07 $layer=LI1_cond $X=5 $Y=3.245 $X2=5
+ $Y2=2.455
r79 9 12 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=0.73 $Y=2.135
+ $X2=0.73 $Y2=2.815
r80 7 38 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.73 $Y=3.245 $X2=0.73
+ $Y2=3.33
r81 7 12 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=0.73 $Y=3.245
+ $X2=0.73 $Y2=2.815
r82 2 15 300 $w=1.7e-07 $l=6.85912e-07 $layer=licon1_PDIFF $count=2 $X=4.85
+ $Y=1.84 $X2=5 $Y2=2.455
r83 1 12 400 $w=1.7e-07 $l=9.26971e-07 $layer=licon1_PDIFF $count=1 $X=0.58
+ $Y=1.96 $X2=0.73 $Y2=2.815
r84 1 9 400 $w=1.7e-07 $l=2.38485e-07 $layer=licon1_PDIFF $count=1 $X=0.58
+ $Y=1.96 $X2=0.73 $Y2=2.135
.ends

.subckt PM_SKY130_FD_SC_HS__NOR4B_2%A_229_368# 1 2 3 12 16 17 18 19 20 22
r48 22 24 2.44 $w=2.5e-07 $l=5e-08 $layer=LI1_cond $X=3.13 $Y=2.46 $X2=3.13
+ $Y2=2.51
r49 21 26 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.275 $Y=2.375
+ $X2=2.15 $Y2=2.375
r50 20 22 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=3.005 $Y=2.375
+ $X2=3.13 $Y2=2.46
r51 20 21 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=3.005 $Y=2.375
+ $X2=2.275 $Y2=2.375
r52 18 26 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.15 $Y=2.46 $X2=2.15
+ $Y2=2.375
r53 18 19 20.5135 $w=2.48e-07 $l=4.45e-07 $layer=LI1_cond $X=2.15 $Y=2.46
+ $X2=2.15 $Y2=2.905
r54 16 19 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=2.025 $Y=2.99
+ $X2=2.15 $Y2=2.905
r55 16 17 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=2.025 $Y=2.99
+ $X2=1.455 $Y2=2.99
r56 12 15 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=1.29 $Y=1.985
+ $X2=1.29 $Y2=2.815
r57 10 17 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.29 $Y=2.905
+ $X2=1.455 $Y2=2.99
r58 10 15 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=1.29 $Y=2.905 $X2=1.29
+ $Y2=2.815
r59 3 24 600 $w=1.7e-07 $l=7.41215e-07 $layer=licon1_PDIFF $count=1 $X=2.94
+ $Y=1.84 $X2=3.09 $Y2=2.51
r60 2 26 300 $w=1.7e-07 $l=6.85912e-07 $layer=licon1_PDIFF $count=2 $X=2.04
+ $Y=1.84 $X2=2.19 $Y2=2.455
r61 1 15 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=1.145
+ $Y=1.84 $X2=1.29 $Y2=2.815
r62 1 12 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=1.145
+ $Y=1.84 $X2=1.29 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HS__NOR4B_2%Y 1 2 3 4 5 18 20 21 22 24 26 30 33 34 35 36
+ 40 46 47 58
r106 47 58 2.07448 $w=5e-07 $l=8.74643e-08 $layer=LI1_cond $X=3.6 $Y=1.01
+ $X2=3.605 $Y2=1.095
r107 46 47 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=3.605 $Y=0.515
+ $X2=3.605 $Y2=0.925
r108 38 40 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=4.98 $Y=1.01
+ $X2=4.98 $Y2=0.515
r109 37 58 11.2921 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.77 $Y=1.095
+ $X2=3.605 $Y2=1.095
r110 36 38 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.815 $Y=1.095
+ $X2=4.98 $Y2=1.01
r111 36 37 68.1765 $w=1.68e-07 $l=1.045e-06 $layer=LI1_cond $X=4.815 $Y=1.095
+ $X2=3.77 $Y2=1.095
r112 34 58 11.2921 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.44 $Y=1.095
+ $X2=3.605 $Y2=1.095
r113 34 35 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=3.44 $Y=1.095
+ $X2=3.095 $Y2=1.095
r114 32 35 5.57278 $w=2.8e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.01 $Y=1.18
+ $X2=3.095 $Y2=1.095
r115 32 33 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=3.01 $Y=1.18
+ $X2=3.01 $Y2=1.95
r116 28 32 17.6464 $w=2.8e-07 $l=4.9295e-07 $layer=LI1_cond $X=2.605 $Y=0.985
+ $X2=3.01 $Y2=1.18
r117 28 30 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=2.605 $Y=0.79
+ $X2=2.605 $Y2=0.515
r118 27 43 3.40825 $w=1.7e-07 $l=1.12916e-07 $layer=LI1_cond $X=1.825 $Y=2.035
+ $X2=1.74 $Y2=1.97
r119 26 33 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.925 $Y=2.035
+ $X2=3.01 $Y2=1.95
r120 26 27 71.7647 $w=1.68e-07 $l=1.1e-06 $layer=LI1_cond $X=2.925 $Y=2.035
+ $X2=1.825 $Y2=2.035
r121 22 43 3.40825 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=1.74 $Y=2.12
+ $X2=1.74 $Y2=1.97
r122 22 24 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=1.74 $Y=2.12
+ $X2=1.74 $Y2=2.57
r123 20 28 9.0585 $w=2.8e-07 $l=2.13014e-07 $layer=LI1_cond $X=2.44 $Y=0.875
+ $X2=2.605 $Y2=0.985
r124 20 21 56.107 $w=1.68e-07 $l=8.6e-07 $layer=LI1_cond $X=2.44 $Y=0.875
+ $X2=1.58 $Y2=0.875
r125 16 21 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.415 $Y=0.79
+ $X2=1.58 $Y2=0.875
r126 16 18 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=1.415 $Y=0.79
+ $X2=1.415 $Y2=0.495
r127 5 43 600 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=1.59
+ $Y=1.84 $X2=1.74 $Y2=1.985
r128 5 24 600 $w=1.7e-07 $l=8.01499e-07 $layer=licon1_PDIFF $count=1 $X=1.59
+ $Y=1.84 $X2=1.74 $Y2=2.57
r129 4 40 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=4.84
+ $Y=0.37 $X2=4.98 $Y2=0.515
r130 3 46 91 $w=1.7e-07 $l=2.20907e-07 $layer=licon1_NDIFF $count=2 $X=3.445
+ $Y=0.37 $X2=3.605 $Y2=0.515
r131 2 30 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.465
+ $Y=0.37 $X2=2.605 $Y2=0.515
r132 1 18 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=1.275
+ $Y=0.37 $X2=1.415 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_HS__NOR4B_2%A_498_368# 1 2 7 11 14
c31 14 0 1.86416e-19 $X=2.64 $Y=2.805
c32 7 0 7.17547e-20 $X=3.935 $Y=2.99
r33 14 16 6.46067 $w=3.28e-07 $l=1.85e-07 $layer=LI1_cond $X=2.64 $Y=2.805
+ $X2=2.64 $Y2=2.99
r34 9 11 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=4.1 $Y=2.905 $X2=4.1
+ $Y2=2.455
r35 8 16 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.805 $Y=2.99
+ $X2=2.64 $Y2=2.99
r36 7 9 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.935 $Y=2.99
+ $X2=4.1 $Y2=2.905
r37 7 8 73.7219 $w=1.68e-07 $l=1.13e-06 $layer=LI1_cond $X=3.935 $Y=2.99
+ $X2=2.805 $Y2=2.99
r38 2 11 300 $w=1.7e-07 $l=6.85912e-07 $layer=licon1_PDIFF $count=2 $X=3.95
+ $Y=1.84 $X2=4.1 $Y2=2.455
r39 1 14 600 $w=1.7e-07 $l=1.03729e-06 $layer=licon1_PDIFF $count=1 $X=2.49
+ $Y=1.84 $X2=2.64 $Y2=2.805
.ends

.subckt PM_SKY130_FD_SC_HS__NOR4B_2%A_701_368# 1 2 3 10 12 14 18 20 22 24 29
c42 14 0 1.87881e-19 $X=4.465 $Y=2.035
r43 22 31 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.5 $Y=2.12 $X2=5.5
+ $Y2=2.035
r44 22 24 14.0598 $w=2.48e-07 $l=3.05e-07 $layer=LI1_cond $X=5.5 $Y=2.12 $X2=5.5
+ $Y2=2.425
r45 21 29 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.635 $Y=2.035
+ $X2=4.55 $Y2=2.035
r46 20 31 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.375 $Y=2.035
+ $X2=5.5 $Y2=2.035
r47 20 21 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=5.375 $Y=2.035
+ $X2=4.635 $Y2=2.035
r48 16 29 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.55 $Y=2.12 $X2=4.55
+ $Y2=2.035
r49 16 18 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=4.55 $Y=2.12
+ $X2=4.55 $Y2=2.425
r50 15 27 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.735 $Y=2.035
+ $X2=3.61 $Y2=2.035
r51 14 29 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.465 $Y=2.035
+ $X2=4.55 $Y2=2.035
r52 14 15 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=4.465 $Y=2.035
+ $X2=3.735 $Y2=2.035
r53 10 27 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.61 $Y=2.12 $X2=3.61
+ $Y2=2.035
r54 10 12 20.744 $w=2.48e-07 $l=4.5e-07 $layer=LI1_cond $X=3.61 $Y=2.12 $X2=3.61
+ $Y2=2.57
r55 3 31 600 $w=1.7e-07 $l=2.59374e-07 $layer=licon1_PDIFF $count=1 $X=5.31
+ $Y=1.84 $X2=5.46 $Y2=2.035
r56 3 24 300 $w=1.7e-07 $l=6.55725e-07 $layer=licon1_PDIFF $count=2 $X=5.31
+ $Y=1.84 $X2=5.46 $Y2=2.425
r57 2 29 600 $w=1.7e-07 $l=2.59374e-07 $layer=licon1_PDIFF $count=1 $X=4.4
+ $Y=1.84 $X2=4.55 $Y2=2.035
r58 2 18 300 $w=1.7e-07 $l=6.55725e-07 $layer=licon1_PDIFF $count=2 $X=4.4
+ $Y=1.84 $X2=4.55 $Y2=2.425
r59 1 27 600 $w=1.7e-07 $l=2.57488e-07 $layer=licon1_PDIFF $count=1 $X=3.505
+ $Y=1.84 $X2=3.65 $Y2=2.035
r60 1 12 600 $w=1.7e-07 $l=7.99218e-07 $layer=licon1_PDIFF $count=1 $X=3.505
+ $Y=1.84 $X2=3.65 $Y2=2.57
.ends

.subckt PM_SKY130_FD_SC_HS__NOR4B_2%VGND 1 2 3 4 5 18 22 24 26 29 30 31 37 41 46
+ 51 58 64 77
c71 22 0 3.60854e-20 $X=3.105 $Y=0.675
r72 76 77 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r73 69 71 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=4.56
+ $Y2=0
r74 64 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r75 58 61 11.8458 $w=5.18e-07 $l=5.15e-07 $layer=LI1_cond $X=2.01 $Y=0 $X2=2.01
+ $Y2=0.515
r76 58 59 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r77 55 77 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=5.52
+ $Y2=0
r78 55 71 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=4.56
+ $Y2=0
r79 54 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r80 52 54 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=4.645 $Y=0 $X2=5.04
+ $Y2=0
r81 51 76 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=5.315 $Y=0 $X2=5.537
+ $Y2=0
r82 51 54 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=5.315 $Y=0 $X2=5.04
+ $Y2=0
r83 50 69 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.08
+ $Y2=0
r84 50 65 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=3.12
+ $Y2=0
r85 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r86 47 64 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.27 $Y=0 $X2=3.105
+ $Y2=0
r87 47 49 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=3.27 $Y=0 $X2=3.6
+ $Y2=0
r88 46 73 10.6035 $w=7.03e-07 $l=6.25e-07 $layer=LI1_cond $X=4.292 $Y=0
+ $X2=4.292 $Y2=0.625
r89 46 52 9.36843 $w=1.7e-07 $l=3.53e-07 $layer=LI1_cond $X=4.292 $Y=0 $X2=4.645
+ $Y2=0
r90 46 71 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r91 46 69 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r92 46 49 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=3.94 $Y=0 $X2=3.6
+ $Y2=0
r93 45 59 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=2.16
+ $Y2=0
r94 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r95 42 58 7.40362 $w=1.7e-07 $l=2.6e-07 $layer=LI1_cond $X=2.27 $Y=0 $X2=2.01
+ $Y2=0
r96 42 44 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=2.27 $Y=0 $X2=2.64
+ $Y2=0
r97 41 64 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.94 $Y=0 $X2=3.105
+ $Y2=0
r98 41 44 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=2.94 $Y=0 $X2=2.64
+ $Y2=0
r99 40 59 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r100 39 40 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r101 37 58 7.40362 $w=1.7e-07 $l=2.6e-07 $layer=LI1_cond $X=1.75 $Y=0 $X2=2.01
+ $Y2=0
r102 37 39 4.56684 $w=1.68e-07 $l=7e-08 $layer=LI1_cond $X=1.75 $Y=0 $X2=1.68
+ $Y2=0
r103 35 40 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r104 34 35 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r105 31 65 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.88 $Y=0
+ $X2=3.12 $Y2=0
r106 31 45 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.88 $Y=0
+ $X2=2.64 $Y2=0
r107 29 34 1.95722 $w=1.68e-07 $l=3e-08 $layer=LI1_cond $X=0.75 $Y=0 $X2=0.72
+ $Y2=0
r108 29 30 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.75 $Y=0 $X2=0.915
+ $Y2=0
r109 28 39 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=1.08 $Y=0 $X2=1.68
+ $Y2=0
r110 28 30 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.08 $Y=0 $X2=0.915
+ $Y2=0
r111 24 76 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=5.48 $Y=0.085
+ $X2=5.537 $Y2=0
r112 24 26 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=5.48 $Y=0.085
+ $X2=5.48 $Y2=0.515
r113 20 64 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.105 $Y=0.085
+ $X2=3.105 $Y2=0
r114 20 22 20.6043 $w=3.28e-07 $l=5.9e-07 $layer=LI1_cond $X=3.105 $Y=0.085
+ $X2=3.105 $Y2=0.675
r115 16 30 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.915 $Y=0.085
+ $X2=0.915 $Y2=0
r116 16 18 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=0.915 $Y=0.085
+ $X2=0.915 $Y2=0.495
r117 5 26 91 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_NDIFF $count=2 $X=5.325
+ $Y=0.37 $X2=5.48 $Y2=0.515
r118 4 73 91 $w=1.7e-07 $l=7.00999e-07 $layer=licon1_NDIFF $count=2 $X=3.965
+ $Y=0.37 $X2=4.55 $Y2=0.625
r119 3 22 182 $w=1.7e-07 $l=3.96327e-07 $layer=licon1_NDIFF $count=1 $X=2.895
+ $Y=0.37 $X2=3.105 $Y2=0.675
r120 2 61 182 $w=1.7e-07 $l=2.98831e-07 $layer=licon1_NDIFF $count=1 $X=1.775
+ $Y=0.37 $X2=2.01 $Y2=0.515
r121 1 18 91 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=2 $X=0.705
+ $Y=0.37 $X2=0.915 $Y2=0.495
.ends

