* File: sky130_fd_sc_hs__sdfstp_2.pxi.spice
* Created: Tue Sep  1 20:23:17 2020
* 
x_PM_SKY130_FD_SC_HS__SDFSTP_2%SCE N_SCE_c_327_n N_SCE_M1042_g N_SCE_c_328_n
+ N_SCE_M1023_g N_SCE_c_329_n N_SCE_M1024_g N_SCE_M1039_g N_SCE_c_322_n
+ N_SCE_c_323_n N_SCE_c_324_n N_SCE_c_325_n SCE N_SCE_c_326_n
+ PM_SKY130_FD_SC_HS__SDFSTP_2%SCE
x_PM_SKY130_FD_SC_HS__SDFSTP_2%A_27_74# N_A_27_74#_M1042_s N_A_27_74#_M1023_s
+ N_A_27_74#_M1038_g N_A_27_74#_c_402_n N_A_27_74#_M1006_g N_A_27_74#_c_396_n
+ N_A_27_74#_c_397_n N_A_27_74#_c_414_n N_A_27_74#_c_398_n N_A_27_74#_c_399_n
+ N_A_27_74#_c_404_n N_A_27_74#_c_400_n N_A_27_74#_c_405_n N_A_27_74#_c_401_n
+ PM_SKY130_FD_SC_HS__SDFSTP_2%A_27_74#
x_PM_SKY130_FD_SC_HS__SDFSTP_2%D N_D_c_470_n N_D_M1045_g N_D_M1022_g D
+ N_D_c_472_n PM_SKY130_FD_SC_HS__SDFSTP_2%D
x_PM_SKY130_FD_SC_HS__SDFSTP_2%SCD N_SCD_M1035_g N_SCD_c_507_n N_SCD_c_511_n
+ N_SCD_M1041_g SCD SCD SCD N_SCD_c_509_n PM_SKY130_FD_SC_HS__SDFSTP_2%SCD
x_PM_SKY130_FD_SC_HS__SDFSTP_2%CLK N_CLK_c_547_n N_CLK_M1002_g N_CLK_c_548_n
+ N_CLK_M1008_g CLK PM_SKY130_FD_SC_HS__SDFSTP_2%CLK
x_PM_SKY130_FD_SC_HS__SDFSTP_2%A_795_74# N_A_795_74#_M1001_d N_A_795_74#_M1018_d
+ N_A_795_74#_c_604_n N_A_795_74#_c_605_n N_A_795_74#_M1014_g
+ N_A_795_74#_c_582_n N_A_795_74#_c_583_n N_A_795_74#_M1030_g
+ N_A_795_74#_c_585_n N_A_795_74#_c_586_n N_A_795_74#_c_587_n
+ N_A_795_74#_M1000_g N_A_795_74#_c_588_n N_A_795_74#_c_589_n
+ N_A_795_74#_M1036_g N_A_795_74#_c_607_n N_A_795_74#_c_608_n
+ N_A_795_74#_M1044_g N_A_795_74#_c_590_n N_A_795_74#_c_591_n
+ N_A_795_74#_c_609_n N_A_795_74#_c_592_n N_A_795_74#_c_593_n
+ N_A_795_74#_c_610_n N_A_795_74#_c_611_n N_A_795_74#_c_594_n
+ N_A_795_74#_c_595_n N_A_795_74#_c_613_n N_A_795_74#_c_614_n
+ N_A_795_74#_c_615_n N_A_795_74#_c_616_n N_A_795_74#_c_617_n
+ N_A_795_74#_c_618_n N_A_795_74#_c_619_n N_A_795_74#_c_620_n
+ N_A_795_74#_c_596_n N_A_795_74#_c_597_n N_A_795_74#_c_623_n
+ N_A_795_74#_c_624_n N_A_795_74#_c_598_n N_A_795_74#_c_625_n
+ N_A_795_74#_c_599_n N_A_795_74#_c_600_n N_A_795_74#_c_601_n
+ N_A_795_74#_c_602_n N_A_795_74#_c_603_n PM_SKY130_FD_SC_HS__SDFSTP_2%A_795_74#
x_PM_SKY130_FD_SC_HS__SDFSTP_2%A_1185_55# N_A_1185_55#_M1020_s
+ N_A_1185_55#_M1015_d N_A_1185_55#_c_878_n N_A_1185_55#_M1007_g
+ N_A_1185_55#_c_885_n N_A_1185_55#_c_886_n N_A_1185_55#_M1028_g
+ N_A_1185_55#_c_879_n N_A_1185_55#_c_880_n N_A_1185_55#_c_887_n
+ N_A_1185_55#_c_881_n N_A_1185_55#_c_902_n N_A_1185_55#_c_888_n
+ N_A_1185_55#_c_882_n N_A_1185_55#_c_890_n N_A_1185_55#_c_883_n
+ N_A_1185_55#_c_884_n PM_SKY130_FD_SC_HS__SDFSTP_2%A_1185_55#
x_PM_SKY130_FD_SC_HS__SDFSTP_2%A_991_81# N_A_991_81#_M1016_d N_A_991_81#_M1014_d
+ N_A_991_81#_c_979_n N_A_991_81#_c_980_n N_A_991_81#_c_998_n
+ N_A_991_81#_M1015_g N_A_991_81#_c_981_n N_A_991_81#_M1020_g
+ N_A_991_81#_c_982_n N_A_991_81#_c_1000_n N_A_991_81#_M1004_g
+ N_A_991_81#_c_983_n N_A_991_81#_M1025_g N_A_991_81#_c_984_n
+ N_A_991_81#_c_1002_n N_A_991_81#_M1009_g N_A_991_81#_c_985_n
+ N_A_991_81#_M1034_g N_A_991_81#_c_986_n N_A_991_81#_c_1003_n
+ N_A_991_81#_c_1004_n N_A_991_81#_c_987_n N_A_991_81#_c_988_n
+ N_A_991_81#_c_989_n N_A_991_81#_c_1083_n N_A_991_81#_c_990_n
+ N_A_991_81#_c_991_n N_A_991_81#_c_992_n N_A_991_81#_c_993_n
+ N_A_991_81#_c_994_n N_A_991_81#_c_995_n N_A_991_81#_c_996_n
+ PM_SKY130_FD_SC_HS__SDFSTP_2%A_991_81#
x_PM_SKY130_FD_SC_HS__SDFSTP_2%SET_B N_SET_B_c_1174_n N_SET_B_c_1185_n
+ N_SET_B_M1029_g N_SET_B_M1021_g N_SET_B_c_1186_n N_SET_B_c_1187_n
+ N_SET_B_M1019_g N_SET_B_M1017_g N_SET_B_c_1177_n N_SET_B_c_1178_n
+ N_SET_B_c_1179_n SET_B N_SET_B_c_1181_n N_SET_B_c_1182_n N_SET_B_c_1183_n
+ PM_SKY130_FD_SC_HS__SDFSTP_2%SET_B
x_PM_SKY130_FD_SC_HS__SDFSTP_2%A_608_74# N_A_608_74#_M1002_s N_A_608_74#_M1008_s
+ N_A_608_74#_M1001_g N_A_608_74#_c_1331_n N_A_608_74#_M1018_g
+ N_A_608_74#_c_1318_n N_A_608_74#_c_1319_n N_A_608_74#_c_1333_n
+ N_A_608_74#_c_1320_n N_A_608_74#_c_1321_n N_A_608_74#_c_1334_n
+ N_A_608_74#_c_1335_n N_A_608_74#_M1016_g N_A_608_74#_c_1336_n
+ N_A_608_74#_M1027_g N_A_608_74#_c_1337_n N_A_608_74#_c_1323_n
+ N_A_608_74#_c_1339_n N_A_608_74#_M1005_g N_A_608_74#_c_1324_n
+ N_A_608_74#_c_1325_n N_A_608_74#_c_1341_n N_A_608_74#_c_1342_n
+ N_A_608_74#_M1010_g N_A_608_74#_M1043_g N_A_608_74#_c_1343_n
+ N_A_608_74#_c_1344_n N_A_608_74#_c_1345_n N_A_608_74#_c_1346_n
+ N_A_608_74#_c_1327_n N_A_608_74#_c_1328_n N_A_608_74#_c_1348_n
+ N_A_608_74#_c_1349_n N_A_608_74#_c_1329_n N_A_608_74#_c_1330_n
+ PM_SKY130_FD_SC_HS__SDFSTP_2%A_608_74#
x_PM_SKY130_FD_SC_HS__SDFSTP_2%A_2186_367# N_A_2186_367#_M1026_d
+ N_A_2186_367#_M1012_s N_A_2186_367#_c_1532_n N_A_2186_367#_c_1533_n
+ N_A_2186_367#_M1040_g N_A_2186_367#_c_1534_n N_A_2186_367#_M1011_g
+ N_A_2186_367#_c_1524_n N_A_2186_367#_c_1525_n N_A_2186_367#_c_1536_n
+ N_A_2186_367#_c_1537_n N_A_2186_367#_c_1538_n N_A_2186_367#_c_1526_n
+ N_A_2186_367#_c_1527_n N_A_2186_367#_c_1528_n N_A_2186_367#_c_1529_n
+ N_A_2186_367#_c_1530_n N_A_2186_367#_c_1531_n
+ PM_SKY130_FD_SC_HS__SDFSTP_2%A_2186_367#
x_PM_SKY130_FD_SC_HS__SDFSTP_2%A_1804_424# N_A_1804_424#_M1000_d
+ N_A_1804_424#_M1036_d N_A_1804_424#_M1005_s N_A_1804_424#_M1010_s
+ N_A_1804_424#_M1019_d N_A_1804_424#_M1026_g N_A_1804_424#_c_1649_n
+ N_A_1804_424#_c_1650_n N_A_1804_424#_M1012_g N_A_1804_424#_c_1636_n
+ N_A_1804_424#_c_1637_n N_A_1804_424#_M1013_g N_A_1804_424#_c_1638_n
+ N_A_1804_424#_c_1652_n N_A_1804_424#_M1031_g N_A_1804_424#_c_1653_n
+ N_A_1804_424#_c_1639_n N_A_1804_424#_c_1654_n N_A_1804_424#_c_1655_n
+ N_A_1804_424#_c_1656_n N_A_1804_424#_c_1640_n N_A_1804_424#_c_1657_n
+ N_A_1804_424#_c_1725_n N_A_1804_424#_c_1641_n N_A_1804_424#_c_1658_n
+ N_A_1804_424#_c_1642_n N_A_1804_424#_c_1643_n N_A_1804_424#_c_1644_n
+ N_A_1804_424#_c_1660_n N_A_1804_424#_c_1661_n N_A_1804_424#_c_1662_n
+ N_A_1804_424#_c_1645_n N_A_1804_424#_c_1646_n N_A_1804_424#_c_1647_n
+ N_A_1804_424#_c_1709_n N_A_1804_424#_c_1663_n N_A_1804_424#_c_1664_n
+ N_A_1804_424#_c_1648_n PM_SKY130_FD_SC_HS__SDFSTP_2%A_1804_424#
x_PM_SKY130_FD_SC_HS__SDFSTP_2%A_2611_98# N_A_2611_98#_M1013_s
+ N_A_2611_98#_M1031_s N_A_2611_98#_c_1846_n N_A_2611_98#_M1032_g
+ N_A_2611_98#_M1003_g N_A_2611_98#_c_1841_n N_A_2611_98#_M1037_g
+ N_A_2611_98#_c_1847_n N_A_2611_98#_M1033_g N_A_2611_98#_c_1842_n
+ N_A_2611_98#_c_1848_n N_A_2611_98#_c_1843_n N_A_2611_98#_c_1844_n
+ N_A_2611_98#_c_1845_n PM_SKY130_FD_SC_HS__SDFSTP_2%A_2611_98#
x_PM_SKY130_FD_SC_HS__SDFSTP_2%VPWR N_VPWR_M1023_d N_VPWR_M1041_d N_VPWR_M1008_d
+ N_VPWR_M1028_d N_VPWR_M1029_d N_VPWR_M1009_s N_VPWR_M1011_d N_VPWR_M1012_d
+ N_VPWR_M1031_d N_VPWR_M1033_s N_VPWR_c_1921_n N_VPWR_c_1922_n N_VPWR_c_1923_n
+ N_VPWR_c_1924_n N_VPWR_c_1925_n N_VPWR_c_1926_n N_VPWR_c_1927_n
+ N_VPWR_c_1928_n N_VPWR_c_1929_n N_VPWR_c_1930_n N_VPWR_c_1931_n
+ N_VPWR_c_1932_n N_VPWR_c_1933_n N_VPWR_c_1934_n N_VPWR_c_1935_n
+ N_VPWR_c_1936_n N_VPWR_c_1937_n N_VPWR_c_1938_n VPWR N_VPWR_c_1939_n
+ N_VPWR_c_1940_n N_VPWR_c_1941_n N_VPWR_c_1942_n N_VPWR_c_1943_n
+ N_VPWR_c_1944_n N_VPWR_c_1945_n N_VPWR_c_1946_n N_VPWR_c_1947_n
+ N_VPWR_c_1948_n N_VPWR_c_1949_n N_VPWR_c_1950_n N_VPWR_c_1920_n
+ PM_SKY130_FD_SC_HS__SDFSTP_2%VPWR
x_PM_SKY130_FD_SC_HS__SDFSTP_2%A_290_464# N_A_290_464#_M1022_d
+ N_A_290_464#_M1016_s N_A_290_464#_M1045_d N_A_290_464#_M1014_s
+ N_A_290_464#_c_2121_n N_A_290_464#_c_2107_n N_A_290_464#_c_2108_n
+ N_A_290_464#_c_2109_n N_A_290_464#_c_2110_n N_A_290_464#_c_2114_n
+ N_A_290_464#_c_2115_n N_A_290_464#_c_2116_n N_A_290_464#_c_2142_n
+ N_A_290_464#_c_2117_n N_A_290_464#_c_2111_n N_A_290_464#_c_2112_n
+ N_A_290_464#_c_2119_n N_A_290_464#_c_2120_n
+ PM_SKY130_FD_SC_HS__SDFSTP_2%A_290_464#
x_PM_SKY130_FD_SC_HS__SDFSTP_2%A_1584_379# N_A_1584_379#_M1004_d
+ N_A_1584_379#_M1005_d N_A_1584_379#_c_2244_n N_A_1584_379#_c_2241_n
+ N_A_1584_379#_c_2258_n N_A_1584_379#_c_2242_n N_A_1584_379#_c_2243_n
+ PM_SKY130_FD_SC_HS__SDFSTP_2%A_1584_379#
x_PM_SKY130_FD_SC_HS__SDFSTP_2%Q N_Q_M1003_d N_Q_M1032_d N_Q_c_2276_n
+ N_Q_c_2281_n N_Q_c_2277_n N_Q_c_2278_n N_Q_c_2279_n Q Q
+ PM_SKY130_FD_SC_HS__SDFSTP_2%Q
x_PM_SKY130_FD_SC_HS__SDFSTP_2%VGND N_VGND_M1042_d N_VGND_M1035_d N_VGND_M1002_d
+ N_VGND_M1007_d N_VGND_M1021_d N_VGND_M1034_s N_VGND_M1017_d N_VGND_M1013_d
+ N_VGND_M1037_s N_VGND_c_2317_n N_VGND_c_2318_n N_VGND_c_2319_n N_VGND_c_2320_n
+ N_VGND_c_2321_n N_VGND_c_2322_n N_VGND_c_2323_n N_VGND_c_2324_n
+ N_VGND_c_2325_n N_VGND_c_2326_n N_VGND_c_2327_n VGND N_VGND_c_2328_n
+ N_VGND_c_2329_n N_VGND_c_2330_n N_VGND_c_2331_n N_VGND_c_2332_n
+ N_VGND_c_2333_n N_VGND_c_2334_n N_VGND_c_2335_n N_VGND_c_2336_n
+ N_VGND_c_2337_n N_VGND_c_2338_n N_VGND_c_2339_n N_VGND_c_2340_n
+ N_VGND_c_2341_n N_VGND_c_2342_n PM_SKY130_FD_SC_HS__SDFSTP_2%VGND
x_PM_SKY130_FD_SC_HS__SDFSTP_2%A_1641_74# N_A_1641_74#_M1025_d
+ N_A_1641_74#_M1000_s N_A_1641_74#_c_2479_n N_A_1641_74#_c_2480_n
+ N_A_1641_74#_c_2481_n N_A_1641_74#_c_2482_n
+ PM_SKY130_FD_SC_HS__SDFSTP_2%A_1641_74#
cc_1 VNB N_SCE_M1042_g 0.0625566f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.58
cc_2 VNB N_SCE_M1039_g 0.0349556f $X=-0.19 $Y=-0.245 $X2=1.94 $Y2=0.58
cc_3 VNB N_SCE_c_322_n 0.0286809f $X=-0.19 $Y=-0.245 $X2=1.795 $Y2=1.495
cc_4 VNB N_SCE_c_323_n 0.00225026f $X=-0.19 $Y=-0.245 $X2=0.805 $Y2=1.495
cc_5 VNB N_SCE_c_324_n 0.00268133f $X=-0.19 $Y=-0.245 $X2=1.96 $Y2=1.415
cc_6 VNB N_SCE_c_325_n 0.0306519f $X=-0.19 $Y=-0.245 $X2=1.96 $Y2=1.415
cc_7 VNB N_SCE_c_326_n 0.0242481f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.635
cc_8 VNB N_A_27_74#_c_396_n 0.023955f $X=-0.19 $Y=-0.245 $X2=1.94 $Y2=0.58
cc_9 VNB N_A_27_74#_c_397_n 0.0203201f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=2.117
cc_10 VNB N_A_27_74#_c_398_n 0.0100668f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_27_74#_c_399_n 0.0334307f $X=-0.19 $Y=-0.245 $X2=1.92 $Y2=1.495
cc_12 VNB N_A_27_74#_c_400_n 0.0203203f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.635
cc_13 VNB N_A_27_74#_c_401_n 0.0182373f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_D_M1022_g 0.0618257f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_SCD_M1035_g 0.0344632f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.47
cc_16 VNB N_SCD_c_507_n 0.0255215f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB SCD 0.00297672f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=2.245
cc_18 VNB N_SCD_c_509_n 0.0333042f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.117
cc_19 VNB N_CLK_c_547_n 0.0200244f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.665
cc_20 VNB N_CLK_c_548_n 0.0394192f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.58
cc_21 VNB CLK 0.00842451f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.245
cc_22 VNB N_A_795_74#_c_582_n 0.0120986f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=2.64
cc_23 VNB N_A_795_74#_c_583_n 0.00683373f $X=-0.19 $Y=-0.245 $X2=1.94 $Y2=0.58
cc_24 VNB N_A_795_74#_M1030_g 0.0362022f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=2.117
cc_25 VNB N_A_795_74#_c_585_n 0.0279309f $X=-0.19 $Y=-0.245 $X2=1.92 $Y2=1.415
cc_26 VNB N_A_795_74#_c_586_n 0.00949433f $X=-0.19 $Y=-0.245 $X2=1.96 $Y2=1.415
cc_27 VNB N_A_795_74#_c_587_n 0.0175524f $X=-0.19 $Y=-0.245 $X2=1.96 $Y2=1.415
cc_28 VNB N_A_795_74#_c_588_n 0.0168332f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_795_74#_c_589_n 0.0148787f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_795_74#_c_590_n 0.00400906f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_795_74#_c_591_n 0.00168954f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_795_74#_c_592_n 0.0170808f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_795_74#_c_593_n 0.00264685f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_795_74#_c_594_n 0.00341946f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_795_74#_c_595_n 0.00339844f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_795_74#_c_596_n 0.00748821f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_795_74#_c_597_n 0.0169131f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_795_74#_c_598_n 0.0051925f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_795_74#_c_599_n 2.60503e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_795_74#_c_600_n 0.0241397f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_795_74#_c_601_n 0.00785969f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_795_74#_c_602_n 0.0126071f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_795_74#_c_603_n 0.0186057f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_1185_55#_c_878_n 0.0173208f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.245
cc_45 VNB N_A_1185_55#_c_879_n 0.0362711f $X=-0.19 $Y=-0.245 $X2=1.94 $Y2=0.58
cc_46 VNB N_A_1185_55#_c_880_n 0.00116198f $X=-0.19 $Y=-0.245 $X2=0.955
+ $Y2=2.117
cc_47 VNB N_A_1185_55#_c_881_n 0.00722463f $X=-0.19 $Y=-0.245 $X2=1.96 $Y2=1.415
cc_48 VNB N_A_1185_55#_c_882_n 0.00471537f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.635
cc_49 VNB N_A_1185_55#_c_883_n 0.0061097f $X=-0.19 $Y=-0.245 $X2=1.96 $Y2=1.25
cc_50 VNB N_A_1185_55#_c_884_n 0.0204767f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_A_991_81#_c_979_n 0.0149666f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.245
cc_52 VNB N_A_991_81#_c_980_n 0.00584511f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.64
cc_53 VNB N_A_991_81#_c_981_n 0.0180022f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=2.64
cc_54 VNB N_A_991_81#_c_982_n 0.00637895f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_A_991_81#_c_983_n 0.0168452f $X=-0.19 $Y=-0.245 $X2=1.795 $Y2=1.495
cc_56 VNB N_A_991_81#_c_984_n 0.00566411f $X=-0.19 $Y=-0.245 $X2=1.96 $Y2=1.415
cc_57 VNB N_A_991_81#_c_985_n 0.0170434f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_58 VNB N_A_991_81#_c_986_n 0.031795f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.47
cc_59 VNB N_A_991_81#_c_987_n 0.00798345f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_A_991_81#_c_988_n 0.0235266f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_A_991_81#_c_989_n 0.0101867f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_A_991_81#_c_990_n 0.0296742f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_A_991_81#_c_991_n 0.0240823f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_A_991_81#_c_992_n 0.00126724f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_A_991_81#_c_993_n 0.00103134f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_A_991_81#_c_994_n 0.00183906f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_A_991_81#_c_995_n 0.00325464f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_A_991_81#_c_996_n 0.0726615f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_SET_B_c_1174_n 0.00671558f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.99
cc_70 VNB N_SET_B_M1021_g 0.0373019f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.64
cc_71 VNB N_SET_B_M1017_g 0.0515369f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.117
cc_72 VNB N_SET_B_c_1177_n 0.0389494f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=2.117
cc_73 VNB N_SET_B_c_1178_n 0.00220503f $X=-0.19 $Y=-0.245 $X2=1.795 $Y2=1.495
cc_74 VNB N_SET_B_c_1179_n 0.00540182f $X=-0.19 $Y=-0.245 $X2=1.96 $Y2=1.415
cc_75 VNB SET_B 0.0040711f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_SET_B_c_1181_n 0.0378364f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.635
cc_77 VNB N_SET_B_c_1182_n 0.0220211f $X=-0.19 $Y=-0.245 $X2=1.96 $Y2=1.415
cc_78 VNB N_SET_B_c_1183_n 0.00779184f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VNB N_A_608_74#_M1001_g 0.0255853f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.64
cc_80 VNB N_A_608_74#_c_1318_n 0.0103779f $X=-0.19 $Y=-0.245 $X2=1.94 $Y2=0.58
cc_81 VNB N_A_608_74#_c_1319_n 0.0385434f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_82 VNB N_A_608_74#_c_1320_n 0.0292071f $X=-0.19 $Y=-0.245 $X2=1.795 $Y2=1.495
cc_83 VNB N_A_608_74#_c_1321_n 0.0103124f $X=-0.19 $Y=-0.245 $X2=0.805 $Y2=1.495
cc_84 VNB N_A_608_74#_M1016_g 0.0272072f $X=-0.19 $Y=-0.245 $X2=1.92 $Y2=1.495
cc_85 VNB N_A_608_74#_c_1323_n 0.00370714f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.47
cc_86 VNB N_A_608_74#_c_1324_n 0.068993f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_87 VNB N_A_608_74#_c_1325_n 0.00767124f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_88 VNB N_A_608_74#_M1043_g 0.0455489f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_89 VNB N_A_608_74#_c_1327_n 0.00838246f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_90 VNB N_A_608_74#_c_1328_n 0.0120978f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_91 VNB N_A_608_74#_c_1329_n 0.00199494f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_92 VNB N_A_608_74#_c_1330_n 0.00302852f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_93 VNB N_A_2186_367#_c_1524_n 0.0218664f $X=-0.19 $Y=-0.245 $X2=0.505
+ $Y2=2.117
cc_94 VNB N_A_2186_367#_c_1525_n 0.0255406f $X=-0.19 $Y=-0.245 $X2=0.61
+ $Y2=2.117
cc_95 VNB N_A_2186_367#_c_1526_n 0.00775159f $X=-0.19 $Y=-0.245 $X2=0.635
+ $Y2=1.58
cc_96 VNB N_A_2186_367#_c_1527_n 0.00617016f $X=-0.19 $Y=-0.245 $X2=0.61
+ $Y2=1.635
cc_97 VNB N_A_2186_367#_c_1528_n 0.00238188f $X=-0.19 $Y=-0.245 $X2=0.64
+ $Y2=1.635
cc_98 VNB N_A_2186_367#_c_1529_n 0.0330841f $X=-0.19 $Y=-0.245 $X2=1.96 $Y2=1.25
cc_99 VNB N_A_2186_367#_c_1530_n 0.00377829f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_100 VNB N_A_2186_367#_c_1531_n 0.0181222f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_101 VNB N_A_1804_424#_M1026_g 0.0396191f $X=-0.19 $Y=-0.245 $X2=0.61
+ $Y2=2.117
cc_102 VNB N_A_1804_424#_c_1636_n 0.0812455f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_103 VNB N_A_1804_424#_c_1637_n 0.0177817f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_104 VNB N_A_1804_424#_c_1638_n 0.00783058f $X=-0.19 $Y=-0.245 $X2=0.61
+ $Y2=1.635
cc_105 VNB N_A_1804_424#_c_1639_n 0.012429f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_106 VNB N_A_1804_424#_c_1640_n 0.00515896f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_107 VNB N_A_1804_424#_c_1641_n 0.00497081f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_108 VNB N_A_1804_424#_c_1642_n 0.00847186f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_109 VNB N_A_1804_424#_c_1643_n 0.0018227f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_110 VNB N_A_1804_424#_c_1644_n 0.00246574f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_111 VNB N_A_1804_424#_c_1645_n 0.00200957f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_112 VNB N_A_1804_424#_c_1646_n 0.0340509f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_113 VNB N_A_1804_424#_c_1647_n 0.00765385f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_114 VNB N_A_1804_424#_c_1648_n 0.0115341f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_115 VNB N_A_2611_98#_M1003_g 0.0212563f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=2.64
cc_116 VNB N_A_2611_98#_c_1841_n 0.0160455f $X=-0.19 $Y=-0.245 $X2=1.94 $Y2=0.58
cc_117 VNB N_A_2611_98#_c_1842_n 0.00961135f $X=-0.19 $Y=-0.245 $X2=1.92
+ $Y2=1.415
cc_118 VNB N_A_2611_98#_c_1843_n 0.00549082f $X=-0.19 $Y=-0.245 $X2=0.64
+ $Y2=1.635
cc_119 VNB N_A_2611_98#_c_1844_n 0.00102441f $X=-0.19 $Y=-0.245 $X2=1.96
+ $Y2=1.415
cc_120 VNB N_A_2611_98#_c_1845_n 0.0685665f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_121 VNB N_VPWR_c_1920_n 0.621437f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_122 VNB N_A_290_464#_c_2107_n 0.00240191f $X=-0.19 $Y=-0.245 $X2=0.955
+ $Y2=2.117
cc_123 VNB N_A_290_464#_c_2108_n 0.0157325f $X=-0.19 $Y=-0.245 $X2=0.805
+ $Y2=1.495
cc_124 VNB N_A_290_464#_c_2109_n 0.00298819f $X=-0.19 $Y=-0.245 $X2=1.92
+ $Y2=1.415
cc_125 VNB N_A_290_464#_c_2110_n 0.00472436f $X=-0.19 $Y=-0.245 $X2=1.96
+ $Y2=1.415
cc_126 VNB N_A_290_464#_c_2111_n 0.00614445f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_127 VNB N_A_290_464#_c_2112_n 0.00705683f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_128 VNB N_Q_c_2276_n 0.00248472f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.64
cc_129 VNB N_Q_c_2277_n 0.0019936f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.117
cc_130 VNB N_Q_c_2278_n 0.0016018f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=2.117
cc_131 VNB N_Q_c_2279_n 0.0112378f $X=-0.19 $Y=-0.245 $X2=1.795 $Y2=1.495
cc_132 VNB Q 0.00712458f $X=-0.19 $Y=-0.245 $X2=0.805 $Y2=1.495
cc_133 VNB N_VGND_c_2317_n 0.00778079f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.58
cc_134 VNB N_VGND_c_2318_n 0.0101978f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.47
cc_135 VNB N_VGND_c_2319_n 0.0201354f $X=-0.19 $Y=-0.245 $X2=1.96 $Y2=1.25
cc_136 VNB N_VGND_c_2320_n 0.00641543f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_137 VNB N_VGND_c_2321_n 0.00826914f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_138 VNB N_VGND_c_2322_n 0.0130607f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_139 VNB N_VGND_c_2323_n 0.0163952f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_140 VNB N_VGND_c_2324_n 0.010678f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_141 VNB N_VGND_c_2325_n 0.0444854f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_142 VNB N_VGND_c_2326_n 0.0152199f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_143 VNB N_VGND_c_2327_n 0.0590232f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_144 VNB N_VGND_c_2328_n 0.0191515f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_145 VNB N_VGND_c_2329_n 0.0412906f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_146 VNB N_VGND_c_2330_n 0.0293898f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_147 VNB N_VGND_c_2331_n 0.019013f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_148 VNB N_VGND_c_2332_n 0.0345145f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_149 VNB N_VGND_c_2333_n 0.0198784f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_150 VNB N_VGND_c_2334_n 0.00856226f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_151 VNB N_VGND_c_2335_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_152 VNB N_VGND_c_2336_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_153 VNB N_VGND_c_2337_n 0.00942782f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_154 VNB N_VGND_c_2338_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_155 VNB N_VGND_c_2339_n 0.0702539f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_156 VNB N_VGND_c_2340_n 0.0234846f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_157 VNB N_VGND_c_2341_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_158 VNB N_VGND_c_2342_n 0.827876f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_159 VNB N_A_1641_74#_c_2479_n 0.0024035f $X=-0.19 $Y=-0.245 $X2=0.505
+ $Y2=2.64
cc_160 VNB N_A_1641_74#_c_2480_n 0.017548f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=2.64
cc_161 VNB N_A_1641_74#_c_2481_n 0.00262272f $X=-0.19 $Y=-0.245 $X2=0.955
+ $Y2=2.64
cc_162 VNB N_A_1641_74#_c_2482_n 0.00193131f $X=-0.19 $Y=-0.245 $X2=1.94
+ $Y2=0.58
cc_163 VPB N_SCE_c_327_n 0.0740361f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=1.99
cc_164 VPB N_SCE_c_328_n 0.0185154f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.245
cc_165 VPB N_SCE_c_329_n 0.0151606f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=2.245
cc_166 VPB SCE 0.00200129f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_167 VPB N_SCE_c_326_n 4.81492e-19 $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.635
cc_168 VPB N_A_27_74#_c_402_n 0.0538288f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=2.245
cc_169 VPB N_A_27_74#_c_397_n 0.0306448f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=2.117
cc_170 VPB N_A_27_74#_c_404_n 0.00363517f $X=-0.19 $Y=1.66 $X2=0.72 $Y2=1.58
cc_171 VPB N_A_27_74#_c_405_n 0.0311364f $X=-0.19 $Y=1.66 $X2=1.96 $Y2=1.415
cc_172 VPB N_D_c_470_n 0.052443f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=1.665
cc_173 VPB N_D_M1022_g 0.0121448f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_174 VPB N_D_c_472_n 0.00778097f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=2.64
cc_175 VPB N_SCD_c_507_n 0.0251262f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_176 VPB N_SCD_c_511_n 0.0564261f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.245
cc_177 VPB SCD 0.0027614f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=2.245
cc_178 VPB N_CLK_c_548_n 0.0246061f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.58
cc_179 VPB N_A_795_74#_c_604_n 0.0224859f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.64
cc_180 VPB N_A_795_74#_c_605_n 0.0205819f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.64
cc_181 VPB N_A_795_74#_c_582_n 0.00688565f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=2.64
cc_182 VPB N_A_795_74#_c_607_n 0.0143536f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.635
cc_183 VPB N_A_795_74#_c_608_n 0.0228231f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=1.47
cc_184 VPB N_A_795_74#_c_609_n 0.00313813f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_185 VPB N_A_795_74#_c_610_n 0.0227665f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_186 VPB N_A_795_74#_c_611_n 0.00296682f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_187 VPB N_A_795_74#_c_594_n 0.00115773f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_188 VPB N_A_795_74#_c_613_n 0.00574398f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_189 VPB N_A_795_74#_c_614_n 0.0014173f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_190 VPB N_A_795_74#_c_615_n 0.0237345f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_191 VPB N_A_795_74#_c_616_n 0.00244172f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_192 VPB N_A_795_74#_c_617_n 0.0138776f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_193 VPB N_A_795_74#_c_618_n 0.00177503f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_194 VPB N_A_795_74#_c_619_n 0.00543398f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_195 VPB N_A_795_74#_c_620_n 3.46324e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_196 VPB N_A_795_74#_c_596_n 0.0232828f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_197 VPB N_A_795_74#_c_597_n 0.0174517f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_198 VPB N_A_795_74#_c_623_n 0.00570882f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_199 VPB N_A_795_74#_c_624_n 0.0321448f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_200 VPB N_A_795_74#_c_625_n 0.0190886f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_201 VPB N_A_795_74#_c_599_n 0.00413795f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_202 VPB N_A_795_74#_c_600_n 0.00859831f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_203 VPB N_A_795_74#_c_601_n 0.0318194f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_204 VPB N_A_1185_55#_c_885_n 0.0110802f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=2.64
cc_205 VPB N_A_1185_55#_c_886_n 0.021901f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=2.64
cc_206 VPB N_A_1185_55#_c_887_n 0.0155588f $X=-0.19 $Y=1.66 $X2=1.92 $Y2=1.415
cc_207 VPB N_A_1185_55#_c_888_n 0.00762449f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_208 VPB N_A_1185_55#_c_882_n 0.0246878f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.635
cc_209 VPB N_A_1185_55#_c_890_n 0.00167294f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=1.47
cc_210 VPB N_A_991_81#_c_980_n 0.0284432f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.64
cc_211 VPB N_A_991_81#_c_998_n 0.0203615f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.64
cc_212 VPB N_A_991_81#_c_982_n 0.00408855f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_213 VPB N_A_991_81#_c_1000_n 0.0192384f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.117
cc_214 VPB N_A_991_81#_c_984_n 0.00370676f $X=-0.19 $Y=1.66 $X2=1.96 $Y2=1.415
cc_215 VPB N_A_991_81#_c_1002_n 0.0195065f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_216 VPB N_A_991_81#_c_1003_n 0.0040866f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_217 VPB N_A_991_81#_c_1004_n 6.48457e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_218 VPB N_A_991_81#_c_993_n 0.00962356f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_219 VPB N_SET_B_c_1174_n 0.0290969f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=1.99
cc_220 VPB N_SET_B_c_1185_n 0.019778f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.47
cc_221 VPB N_SET_B_c_1186_n 0.0344302f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=2.64
cc_222 VPB N_SET_B_c_1187_n 0.0263253f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=2.64
cc_223 VPB N_SET_B_c_1182_n 0.0169762f $X=-0.19 $Y=1.66 $X2=1.96 $Y2=1.415
cc_224 VPB N_SET_B_c_1183_n 0.00397329f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_225 VPB N_A_608_74#_c_1331_n 0.0151715f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=2.64
cc_226 VPB N_A_608_74#_c_1319_n 0.0178138f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_227 VPB N_A_608_74#_c_1333_n 0.0563946f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=2.117
cc_228 VPB N_A_608_74#_c_1334_n 0.062327f $X=-0.19 $Y=1.66 $X2=1.92 $Y2=1.415
cc_229 VPB N_A_608_74#_c_1335_n 0.0123764f $X=-0.19 $Y=1.66 $X2=1.96 $Y2=1.415
cc_230 VPB N_A_608_74#_c_1336_n 0.0158112f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_231 VPB N_A_608_74#_c_1337_n 0.293738f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=1.635
cc_232 VPB N_A_608_74#_c_1323_n 0.0225218f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=1.47
cc_233 VPB N_A_608_74#_c_1339_n 0.00729337f $X=-0.19 $Y=1.66 $X2=1.96 $Y2=1.415
cc_234 VPB N_A_608_74#_M1005_g 0.00856473f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_235 VPB N_A_608_74#_c_1341_n 0.0359513f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_236 VPB N_A_608_74#_c_1342_n 0.0138501f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_237 VPB N_A_608_74#_c_1343_n 0.0147177f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_238 VPB N_A_608_74#_c_1344_n 0.010113f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_239 VPB N_A_608_74#_c_1345_n 0.0226552f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_240 VPB N_A_608_74#_c_1346_n 0.0122239f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_241 VPB N_A_608_74#_c_1328_n 0.00357202f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_242 VPB N_A_608_74#_c_1348_n 0.0118698f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_243 VPB N_A_608_74#_c_1349_n 0.00459351f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_244 VPB N_A_608_74#_c_1329_n 8.82238e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_245 VPB N_A_2186_367#_c_1532_n 0.00507698f $X=-0.19 $Y=1.66 $X2=0.505
+ $Y2=2.245
cc_246 VPB N_A_2186_367#_c_1533_n 0.0191778f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.64
cc_247 VPB N_A_2186_367#_c_1534_n 0.0196179f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=2.64
cc_248 VPB N_A_2186_367#_c_1524_n 0.0105007f $X=-0.19 $Y=1.66 $X2=0.505
+ $Y2=2.117
cc_249 VPB N_A_2186_367#_c_1536_n 0.00760269f $X=-0.19 $Y=1.66 $X2=1.92
+ $Y2=1.415
cc_250 VPB N_A_2186_367#_c_1537_n 0.00903182f $X=-0.19 $Y=1.66 $X2=1.96
+ $Y2=1.415
cc_251 VPB N_A_2186_367#_c_1538_n 0.0037735f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_252 VPB N_A_2186_367#_c_1527_n 0.0126855f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=1.635
cc_253 VPB N_A_1804_424#_c_1649_n 0.0166506f $X=-0.19 $Y=1.66 $X2=0.805
+ $Y2=1.495
cc_254 VPB N_A_1804_424#_c_1650_n 0.0289592f $X=-0.19 $Y=1.66 $X2=1.92 $Y2=1.415
cc_255 VPB N_A_1804_424#_c_1638_n 0.00921906f $X=-0.19 $Y=1.66 $X2=0.61
+ $Y2=1.635
cc_256 VPB N_A_1804_424#_c_1652_n 0.0259036f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.635
cc_257 VPB N_A_1804_424#_c_1653_n 0.0213273f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_258 VPB N_A_1804_424#_c_1654_n 0.00681579f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_259 VPB N_A_1804_424#_c_1655_n 0.00687114f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_260 VPB N_A_1804_424#_c_1656_n 0.00279745f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_261 VPB N_A_1804_424#_c_1657_n 9.54452e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_262 VPB N_A_1804_424#_c_1658_n 0.0025529f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_263 VPB N_A_1804_424#_c_1644_n 0.00611054f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_264 VPB N_A_1804_424#_c_1660_n 0.00823271f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_265 VPB N_A_1804_424#_c_1661_n 0.0165649f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_266 VPB N_A_1804_424#_c_1662_n 0.00210961f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_267 VPB N_A_1804_424#_c_1663_n 0.0117212f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_268 VPB N_A_1804_424#_c_1664_n 0.0217852f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_269 VPB N_A_1804_424#_c_1648_n 0.0294988f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_270 VPB N_A_2611_98#_c_1846_n 0.0161498f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.245
cc_271 VPB N_A_2611_98#_c_1847_n 0.017582f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.117
cc_272 VPB N_A_2611_98#_c_1848_n 0.0169267f $X=-0.19 $Y=1.66 $X2=1.92 $Y2=1.495
cc_273 VPB N_A_2611_98#_c_1845_n 0.0147442f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_274 VPB N_VPWR_c_1921_n 0.00396467f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.635
cc_275 VPB N_VPWR_c_1922_n 0.00967532f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_276 VPB N_VPWR_c_1923_n 0.0196669f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_277 VPB N_VPWR_c_1924_n 0.00339692f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_278 VPB N_VPWR_c_1925_n 0.00564397f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_279 VPB N_VPWR_c_1926_n 0.0125578f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_280 VPB N_VPWR_c_1927_n 0.0179086f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_281 VPB N_VPWR_c_1928_n 0.00571271f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_282 VPB N_VPWR_c_1929_n 0.0112089f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_283 VPB N_VPWR_c_1930_n 0.0119914f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_284 VPB N_VPWR_c_1931_n 0.0116916f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_285 VPB N_VPWR_c_1932_n 0.0348828f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_286 VPB N_VPWR_c_1933_n 0.0541194f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_287 VPB N_VPWR_c_1934_n 0.00330333f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_288 VPB N_VPWR_c_1935_n 0.027717f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_289 VPB N_VPWR_c_1936_n 0.00223798f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_290 VPB N_VPWR_c_1937_n 0.019428f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_291 VPB N_VPWR_c_1938_n 0.00330333f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_292 VPB N_VPWR_c_1939_n 0.0180274f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_293 VPB N_VPWR_c_1940_n 0.0455708f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_294 VPB N_VPWR_c_1941_n 0.0611503f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_295 VPB N_VPWR_c_1942_n 0.0328287f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_296 VPB N_VPWR_c_1943_n 0.0196104f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_297 VPB N_VPWR_c_1944_n 0.0173363f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_298 VPB N_VPWR_c_1945_n 0.00601644f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_299 VPB N_VPWR_c_1946_n 0.00631651f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_300 VPB N_VPWR_c_1947_n 0.00601644f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_301 VPB N_VPWR_c_1948_n 0.00460249f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_302 VPB N_VPWR_c_1949_n 0.00614127f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_303 VPB N_VPWR_c_1950_n 0.00545601f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_304 VPB N_VPWR_c_1920_n 0.118412f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_305 VPB N_A_290_464#_c_2110_n 0.00529321f $X=-0.19 $Y=1.66 $X2=1.96 $Y2=1.415
cc_306 VPB N_A_290_464#_c_2114_n 0.00531915f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_307 VPB N_A_290_464#_c_2115_n 0.00451248f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_308 VPB N_A_290_464#_c_2116_n 0.00165521f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.635
cc_309 VPB N_A_290_464#_c_2117_n 0.0123642f $X=-0.19 $Y=1.66 $X2=1.96 $Y2=1.25
cc_310 VPB N_A_290_464#_c_2112_n 0.00207118f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_311 VPB N_A_290_464#_c_2119_n 0.00658745f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_312 VPB N_A_290_464#_c_2120_n 0.00497586f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_313 VPB N_A_1584_379#_c_2241_n 0.017113f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=2.64
cc_314 VPB N_A_1584_379#_c_2242_n 0.00244126f $X=-0.19 $Y=1.66 $X2=0.61
+ $Y2=2.117
cc_315 VPB N_A_1584_379#_c_2243_n 0.00694827f $X=-0.19 $Y=1.66 $X2=0.955
+ $Y2=2.117
cc_316 VPB N_Q_c_2281_n 0.00243101f $X=-0.19 $Y=1.66 $X2=1.94 $Y2=1.25
cc_317 VPB Q 0.00758458f $X=-0.19 $Y=1.66 $X2=0.805 $Y2=1.495
cc_318 VPB Q 0.0167374f $X=-0.19 $Y=1.66 $X2=1.92 $Y2=1.415
cc_319 N_SCE_c_324_n N_A_27_74#_c_402_n 3.1694e-19 $X=1.96 $Y=1.415 $X2=0 $Y2=0
cc_320 N_SCE_c_325_n N_A_27_74#_c_402_n 0.0183854f $X=1.96 $Y=1.415 $X2=0 $Y2=0
cc_321 N_SCE_M1042_g N_A_27_74#_c_396_n 0.0115261f $X=0.495 $Y=0.58 $X2=0 $Y2=0
cc_322 N_SCE_M1042_g N_A_27_74#_c_397_n 0.00757393f $X=0.495 $Y=0.58 $X2=0 $Y2=0
cc_323 N_SCE_c_328_n N_A_27_74#_c_397_n 0.00225127f $X=0.505 $Y=2.245 $X2=0
+ $Y2=0
cc_324 N_SCE_c_323_n N_A_27_74#_c_397_n 0.0124456f $X=0.805 $Y=1.495 $X2=0 $Y2=0
cc_325 SCE N_A_27_74#_c_397_n 0.0386025f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_326 N_SCE_c_326_n N_A_27_74#_c_397_n 0.0206346f $X=0.64 $Y=1.635 $X2=0 $Y2=0
cc_327 N_SCE_c_327_n N_A_27_74#_c_414_n 0.00269547f $X=0.61 $Y=1.99 $X2=0 $Y2=0
cc_328 N_SCE_c_328_n N_A_27_74#_c_414_n 0.0112449f $X=0.505 $Y=2.245 $X2=0 $Y2=0
cc_329 N_SCE_c_329_n N_A_27_74#_c_414_n 0.0157821f $X=0.955 $Y=2.245 $X2=0 $Y2=0
cc_330 SCE N_A_27_74#_c_414_n 0.0224122f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_331 N_SCE_M1042_g N_A_27_74#_c_398_n 0.0166195f $X=0.495 $Y=0.58 $X2=0 $Y2=0
cc_332 N_SCE_c_322_n N_A_27_74#_c_398_n 0.030574f $X=1.795 $Y=1.495 $X2=0 $Y2=0
cc_333 N_SCE_c_323_n N_A_27_74#_c_398_n 0.0272015f $X=0.805 $Y=1.495 $X2=0 $Y2=0
cc_334 N_SCE_c_326_n N_A_27_74#_c_398_n 0.00145888f $X=0.64 $Y=1.635 $X2=0 $Y2=0
cc_335 N_SCE_M1042_g N_A_27_74#_c_399_n 0.0123124f $X=0.495 $Y=0.58 $X2=0 $Y2=0
cc_336 N_SCE_c_322_n N_A_27_74#_c_399_n 0.00793591f $X=1.795 $Y=1.495 $X2=0
+ $Y2=0
cc_337 N_SCE_c_324_n N_A_27_74#_c_404_n 0.0145428f $X=1.96 $Y=1.415 $X2=0 $Y2=0
cc_338 N_SCE_c_325_n N_A_27_74#_c_404_n 3.1381e-19 $X=1.96 $Y=1.415 $X2=0 $Y2=0
cc_339 N_SCE_M1042_g N_A_27_74#_c_400_n 0.00874187f $X=0.495 $Y=0.58 $X2=0 $Y2=0
cc_340 N_SCE_c_326_n N_A_27_74#_c_400_n 2.24402e-19 $X=0.64 $Y=1.635 $X2=0 $Y2=0
cc_341 N_SCE_c_328_n N_A_27_74#_c_405_n 0.00545682f $X=0.505 $Y=2.245 $X2=0
+ $Y2=0
cc_342 N_SCE_M1042_g N_A_27_74#_c_401_n 0.0139046f $X=0.495 $Y=0.58 $X2=0 $Y2=0
cc_343 N_SCE_c_327_n N_D_c_470_n 0.0198525f $X=0.61 $Y=1.99 $X2=-0.19 $Y2=-0.245
cc_344 N_SCE_c_329_n N_D_c_470_n 0.0400037f $X=0.955 $Y=2.245 $X2=-0.19
+ $Y2=-0.245
cc_345 N_SCE_c_322_n N_D_c_470_n 0.00435959f $X=1.795 $Y=1.495 $X2=-0.19
+ $Y2=-0.245
cc_346 SCE N_D_c_470_n 2.74008e-19 $X=0.635 $Y=1.58 $X2=-0.19 $Y2=-0.245
cc_347 N_SCE_M1039_g N_D_M1022_g 0.0284734f $X=1.94 $Y=0.58 $X2=0 $Y2=0
cc_348 N_SCE_c_322_n N_D_M1022_g 0.015938f $X=1.795 $Y=1.495 $X2=0 $Y2=0
cc_349 N_SCE_c_324_n N_D_M1022_g 0.00118673f $X=1.96 $Y=1.415 $X2=0 $Y2=0
cc_350 N_SCE_c_325_n N_D_M1022_g 0.0212609f $X=1.96 $Y=1.415 $X2=0 $Y2=0
cc_351 SCE N_D_M1022_g 0.00116396f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_352 N_SCE_c_326_n N_D_M1022_g 0.00639795f $X=0.64 $Y=1.635 $X2=0 $Y2=0
cc_353 N_SCE_c_327_n N_D_c_472_n 0.00328952f $X=0.61 $Y=1.99 $X2=0 $Y2=0
cc_354 N_SCE_c_322_n N_D_c_472_n 0.0291812f $X=1.795 $Y=1.495 $X2=0 $Y2=0
cc_355 SCE N_D_c_472_n 0.0180473f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_356 N_SCE_M1039_g N_SCD_M1035_g 0.0368573f $X=1.94 $Y=0.58 $X2=0 $Y2=0
cc_357 N_SCE_c_324_n N_SCD_c_509_n 2.87119e-19 $X=1.96 $Y=1.415 $X2=0 $Y2=0
cc_358 N_SCE_c_325_n N_SCD_c_509_n 0.0204387f $X=1.96 $Y=1.415 $X2=0 $Y2=0
cc_359 N_SCE_c_328_n N_VPWR_c_1921_n 0.0101271f $X=0.505 $Y=2.245 $X2=0 $Y2=0
cc_360 N_SCE_c_329_n N_VPWR_c_1921_n 0.00946621f $X=0.955 $Y=2.245 $X2=0 $Y2=0
cc_361 N_SCE_c_328_n N_VPWR_c_1939_n 0.00413917f $X=0.505 $Y=2.245 $X2=0 $Y2=0
cc_362 N_SCE_c_329_n N_VPWR_c_1940_n 0.00413917f $X=0.955 $Y=2.245 $X2=0 $Y2=0
cc_363 N_SCE_c_328_n N_VPWR_c_1920_n 0.00417999f $X=0.505 $Y=2.245 $X2=0 $Y2=0
cc_364 N_SCE_c_329_n N_VPWR_c_1920_n 0.00414311f $X=0.955 $Y=2.245 $X2=0 $Y2=0
cc_365 N_SCE_c_329_n N_A_290_464#_c_2121_n 7.12872e-19 $X=0.955 $Y=2.245 $X2=0
+ $Y2=0
cc_366 N_SCE_M1039_g N_A_290_464#_c_2107_n 0.0125369f $X=1.94 $Y=0.58 $X2=0
+ $Y2=0
cc_367 N_SCE_M1039_g N_A_290_464#_c_2108_n 0.0111573f $X=1.94 $Y=0.58 $X2=0
+ $Y2=0
cc_368 N_SCE_c_324_n N_A_290_464#_c_2108_n 0.0111296f $X=1.96 $Y=1.415 $X2=0
+ $Y2=0
cc_369 N_SCE_c_325_n N_A_290_464#_c_2108_n 0.0032473f $X=1.96 $Y=1.415 $X2=0
+ $Y2=0
cc_370 N_SCE_M1039_g N_A_290_464#_c_2109_n 0.00274486f $X=1.94 $Y=0.58 $X2=0
+ $Y2=0
cc_371 N_SCE_c_322_n N_A_290_464#_c_2109_n 0.0123012f $X=1.795 $Y=1.495 $X2=0
+ $Y2=0
cc_372 N_SCE_c_324_n N_A_290_464#_c_2109_n 0.00785342f $X=1.96 $Y=1.415 $X2=0
+ $Y2=0
cc_373 N_SCE_c_325_n N_A_290_464#_c_2109_n 5.46117e-19 $X=1.96 $Y=1.415 $X2=0
+ $Y2=0
cc_374 N_SCE_M1039_g N_A_290_464#_c_2110_n 0.00343685f $X=1.94 $Y=0.58 $X2=0
+ $Y2=0
cc_375 N_SCE_c_324_n N_A_290_464#_c_2110_n 0.0242834f $X=1.96 $Y=1.415 $X2=0
+ $Y2=0
cc_376 N_SCE_c_325_n N_A_290_464#_c_2110_n 0.00204642f $X=1.96 $Y=1.415 $X2=0
+ $Y2=0
cc_377 N_SCE_M1042_g N_VGND_c_2317_n 0.00572943f $X=0.495 $Y=0.58 $X2=0 $Y2=0
cc_378 N_SCE_M1039_g N_VGND_c_2318_n 0.00172001f $X=1.94 $Y=0.58 $X2=0 $Y2=0
cc_379 N_SCE_M1042_g N_VGND_c_2328_n 0.00434272f $X=0.495 $Y=0.58 $X2=0 $Y2=0
cc_380 N_SCE_M1039_g N_VGND_c_2329_n 0.00434272f $X=1.94 $Y=0.58 $X2=0 $Y2=0
cc_381 N_SCE_M1042_g N_VGND_c_2342_n 0.00825349f $X=0.495 $Y=0.58 $X2=0 $Y2=0
cc_382 N_SCE_M1039_g N_VGND_c_2342_n 0.00821825f $X=1.94 $Y=0.58 $X2=0 $Y2=0
cc_383 N_A_27_74#_c_402_n N_D_c_470_n 0.0433856f $X=2.005 $Y=2.245 $X2=-0.19
+ $Y2=-0.245
cc_384 N_A_27_74#_c_414_n N_D_c_470_n 0.0156036f $X=1.795 $Y=2.405 $X2=-0.19
+ $Y2=-0.245
cc_385 N_A_27_74#_c_404_n N_D_c_470_n 0.00360745f $X=1.96 $Y=1.995 $X2=-0.19
+ $Y2=-0.245
cc_386 N_A_27_74#_c_398_n N_D_M1022_g 0.00157925f $X=1.06 $Y=1.065 $X2=0 $Y2=0
cc_387 N_A_27_74#_c_399_n N_D_M1022_g 0.0196496f $X=1.06 $Y=1.065 $X2=0 $Y2=0
cc_388 N_A_27_74#_c_401_n N_D_M1022_g 0.0336314f $X=1.06 $Y=0.9 $X2=0 $Y2=0
cc_389 N_A_27_74#_c_402_n N_D_c_472_n 0.00111057f $X=2.005 $Y=2.245 $X2=0 $Y2=0
cc_390 N_A_27_74#_c_414_n N_D_c_472_n 0.0330418f $X=1.795 $Y=2.405 $X2=0 $Y2=0
cc_391 N_A_27_74#_c_404_n N_D_c_472_n 0.0205429f $X=1.96 $Y=1.995 $X2=0 $Y2=0
cc_392 N_A_27_74#_c_402_n N_SCD_c_507_n 0.0204354f $X=2.005 $Y=2.245 $X2=0 $Y2=0
cc_393 N_A_27_74#_c_404_n N_SCD_c_507_n 3.67751e-19 $X=1.96 $Y=1.995 $X2=0 $Y2=0
cc_394 N_A_27_74#_c_402_n N_SCD_c_511_n 0.0422354f $X=2.005 $Y=2.245 $X2=0 $Y2=0
cc_395 N_A_27_74#_c_414_n N_VPWR_M1023_d 0.00360227f $X=1.795 $Y=2.405 $X2=-0.19
+ $Y2=-0.245
cc_396 N_A_27_74#_c_414_n N_VPWR_c_1921_n 0.0168032f $X=1.795 $Y=2.405 $X2=0
+ $Y2=0
cc_397 N_A_27_74#_c_405_n N_VPWR_c_1921_n 0.0214859f $X=0.28 $Y=2.475 $X2=0
+ $Y2=0
cc_398 N_A_27_74#_c_405_n N_VPWR_c_1939_n 0.0110622f $X=0.28 $Y=2.475 $X2=0
+ $Y2=0
cc_399 N_A_27_74#_c_402_n N_VPWR_c_1940_n 0.00300876f $X=2.005 $Y=2.245 $X2=0
+ $Y2=0
cc_400 N_A_27_74#_c_402_n N_VPWR_c_1920_n 0.00370184f $X=2.005 $Y=2.245 $X2=0
+ $Y2=0
cc_401 N_A_27_74#_c_414_n N_VPWR_c_1920_n 0.0242263f $X=1.795 $Y=2.405 $X2=0
+ $Y2=0
cc_402 N_A_27_74#_c_405_n N_VPWR_c_1920_n 0.00915799f $X=0.28 $Y=2.475 $X2=0
+ $Y2=0
cc_403 N_A_27_74#_c_414_n A_206_464# 0.00479872f $X=1.795 $Y=2.405 $X2=-0.19
+ $Y2=-0.245
cc_404 N_A_27_74#_c_414_n N_A_290_464#_M1045_d 0.0134049f $X=1.795 $Y=2.405
+ $X2=0 $Y2=0
cc_405 N_A_27_74#_c_402_n N_A_290_464#_c_2121_n 0.0149949f $X=2.005 $Y=2.245
+ $X2=0 $Y2=0
cc_406 N_A_27_74#_c_414_n N_A_290_464#_c_2121_n 0.0370379f $X=1.795 $Y=2.405
+ $X2=0 $Y2=0
cc_407 N_A_27_74#_c_398_n N_A_290_464#_c_2107_n 3.9435e-19 $X=1.06 $Y=1.065
+ $X2=0 $Y2=0
cc_408 N_A_27_74#_c_401_n N_A_290_464#_c_2107_n 0.00202258f $X=1.06 $Y=0.9 $X2=0
+ $Y2=0
cc_409 N_A_27_74#_c_398_n N_A_290_464#_c_2109_n 0.00831735f $X=1.06 $Y=1.065
+ $X2=0 $Y2=0
cc_410 N_A_27_74#_c_402_n N_A_290_464#_c_2110_n 0.00762667f $X=2.005 $Y=2.245
+ $X2=0 $Y2=0
cc_411 N_A_27_74#_c_414_n N_A_290_464#_c_2110_n 0.0133253f $X=1.795 $Y=2.405
+ $X2=0 $Y2=0
cc_412 N_A_27_74#_c_404_n N_A_290_464#_c_2110_n 0.0359858f $X=1.96 $Y=1.995
+ $X2=0 $Y2=0
cc_413 N_A_27_74#_c_402_n N_A_290_464#_c_2142_n 2.80564e-19 $X=2.005 $Y=2.245
+ $X2=0 $Y2=0
cc_414 N_A_27_74#_c_396_n N_VGND_c_2317_n 0.0132122f $X=0.28 $Y=0.58 $X2=0 $Y2=0
cc_415 N_A_27_74#_c_398_n N_VGND_c_2317_n 0.0292604f $X=1.06 $Y=1.065 $X2=0
+ $Y2=0
cc_416 N_A_27_74#_c_399_n N_VGND_c_2317_n 0.00320405f $X=1.06 $Y=1.065 $X2=0
+ $Y2=0
cc_417 N_A_27_74#_c_401_n N_VGND_c_2317_n 0.015423f $X=1.06 $Y=0.9 $X2=0 $Y2=0
cc_418 N_A_27_74#_c_396_n N_VGND_c_2328_n 0.0145639f $X=0.28 $Y=0.58 $X2=0 $Y2=0
cc_419 N_A_27_74#_c_401_n N_VGND_c_2329_n 0.00383152f $X=1.06 $Y=0.9 $X2=0 $Y2=0
cc_420 N_A_27_74#_c_396_n N_VGND_c_2342_n 0.0119984f $X=0.28 $Y=0.58 $X2=0 $Y2=0
cc_421 N_A_27_74#_c_401_n N_VGND_c_2342_n 0.0075725f $X=1.06 $Y=0.9 $X2=0 $Y2=0
cc_422 N_D_c_470_n N_VPWR_c_1921_n 0.0016042f $X=1.375 $Y=2.245 $X2=0 $Y2=0
cc_423 N_D_c_470_n N_VPWR_c_1940_n 0.00445405f $X=1.375 $Y=2.245 $X2=0 $Y2=0
cc_424 N_D_c_470_n N_VPWR_c_1920_n 0.00456649f $X=1.375 $Y=2.245 $X2=0 $Y2=0
cc_425 N_D_c_470_n N_A_290_464#_c_2121_n 0.00888514f $X=1.375 $Y=2.245 $X2=0
+ $Y2=0
cc_426 N_D_M1022_g N_A_290_464#_c_2107_n 0.0116998f $X=1.51 $Y=0.58 $X2=0 $Y2=0
cc_427 N_D_M1022_g N_A_290_464#_c_2109_n 0.00483064f $X=1.51 $Y=0.58 $X2=0 $Y2=0
cc_428 N_D_M1022_g N_A_290_464#_c_2110_n 0.00511872f $X=1.51 $Y=0.58 $X2=0 $Y2=0
cc_429 N_D_c_472_n N_A_290_464#_c_2110_n 2.57555e-19 $X=1.42 $Y=1.985 $X2=0
+ $Y2=0
cc_430 N_D_M1022_g N_VGND_c_2317_n 0.00149152f $X=1.51 $Y=0.58 $X2=0 $Y2=0
cc_431 N_D_M1022_g N_VGND_c_2329_n 0.00434272f $X=1.51 $Y=0.58 $X2=0 $Y2=0
cc_432 N_D_M1022_g N_VGND_c_2342_n 0.00821077f $X=1.51 $Y=0.58 $X2=0 $Y2=0
cc_433 N_SCD_c_509_n N_CLK_c_547_n 0.00140608f $X=2.665 $Y=1.305 $X2=-0.19
+ $Y2=-0.245
cc_434 N_SCD_c_507_n N_CLK_c_548_n 0.00682323f $X=2.582 $Y=1.903 $X2=0 $Y2=0
cc_435 N_SCD_c_509_n N_CLK_c_548_n 0.00730373f $X=2.665 $Y=1.305 $X2=0 $Y2=0
cc_436 N_SCD_M1035_g N_A_608_74#_c_1327_n 0.00901831f $X=2.41 $Y=0.58 $X2=0
+ $Y2=0
cc_437 SCD N_A_608_74#_c_1328_n 0.0474887f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_438 N_SCD_c_509_n N_A_608_74#_c_1328_n 0.00688477f $X=2.665 $Y=1.305 $X2=0
+ $Y2=0
cc_439 N_SCD_c_507_n N_A_608_74#_c_1349_n 0.00305508f $X=2.582 $Y=1.903 $X2=0
+ $Y2=0
cc_440 SCD N_A_608_74#_c_1349_n 0.0196463f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_441 N_SCD_c_511_n N_VPWR_c_1922_n 0.00927755f $X=2.425 $Y=2.245 $X2=0 $Y2=0
cc_442 N_SCD_c_511_n N_VPWR_c_1940_n 0.00324189f $X=2.425 $Y=2.245 $X2=0 $Y2=0
cc_443 N_SCD_c_511_n N_VPWR_c_1920_n 0.00412773f $X=2.425 $Y=2.245 $X2=0 $Y2=0
cc_444 N_SCD_c_511_n N_A_290_464#_c_2121_n 2.83395e-19 $X=2.425 $Y=2.245 $X2=0
+ $Y2=0
cc_445 N_SCD_M1035_g N_A_290_464#_c_2107_n 0.00199239f $X=2.41 $Y=0.58 $X2=0
+ $Y2=0
cc_446 N_SCD_M1035_g N_A_290_464#_c_2108_n 0.00850446f $X=2.41 $Y=0.58 $X2=0
+ $Y2=0
cc_447 N_SCD_M1035_g N_A_290_464#_c_2110_n 0.00172798f $X=2.41 $Y=0.58 $X2=0
+ $Y2=0
cc_448 N_SCD_c_507_n N_A_290_464#_c_2110_n 0.0148573f $X=2.582 $Y=1.903 $X2=0
+ $Y2=0
cc_449 N_SCD_c_511_n N_A_290_464#_c_2110_n 0.0173206f $X=2.425 $Y=2.245 $X2=0
+ $Y2=0
cc_450 SCD N_A_290_464#_c_2110_n 0.069827f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_451 N_SCD_c_509_n N_A_290_464#_c_2110_n 0.0060148f $X=2.665 $Y=1.305 $X2=0
+ $Y2=0
cc_452 N_SCD_c_511_n N_A_290_464#_c_2114_n 0.0168177f $X=2.425 $Y=2.245 $X2=0
+ $Y2=0
cc_453 SCD N_A_290_464#_c_2114_n 0.0102308f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_454 N_SCD_c_511_n N_A_290_464#_c_2142_n 0.0122878f $X=2.425 $Y=2.245 $X2=0
+ $Y2=0
cc_455 N_SCD_c_511_n N_A_290_464#_c_2117_n 0.00453491f $X=2.425 $Y=2.245 $X2=0
+ $Y2=0
cc_456 N_SCD_M1035_g N_VGND_c_2318_n 0.0135277f $X=2.41 $Y=0.58 $X2=0 $Y2=0
cc_457 SCD N_VGND_c_2318_n 0.0100559f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_458 N_SCD_c_509_n N_VGND_c_2318_n 0.00355058f $X=2.665 $Y=1.305 $X2=0 $Y2=0
cc_459 N_SCD_M1035_g N_VGND_c_2329_n 0.00383152f $X=2.41 $Y=0.58 $X2=0 $Y2=0
cc_460 N_SCD_M1035_g N_VGND_c_2342_n 0.00757998f $X=2.41 $Y=0.58 $X2=0 $Y2=0
cc_461 N_CLK_c_547_n N_A_608_74#_M1001_g 0.0175799f $X=3.4 $Y=1.22 $X2=0 $Y2=0
cc_462 N_CLK_c_548_n N_A_608_74#_M1001_g 0.0174253f $X=3.485 $Y=1.765 $X2=0
+ $Y2=0
cc_463 CLK N_A_608_74#_M1001_g 0.00597538f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_464 N_CLK_c_548_n N_A_608_74#_c_1331_n 0.0413738f $X=3.485 $Y=1.765 $X2=0
+ $Y2=0
cc_465 N_CLK_c_548_n N_A_608_74#_c_1319_n 0.0112647f $X=3.485 $Y=1.765 $X2=0
+ $Y2=0
cc_466 N_CLK_c_547_n N_A_608_74#_c_1327_n 0.00580215f $X=3.4 $Y=1.22 $X2=0 $Y2=0
cc_467 N_CLK_c_547_n N_A_608_74#_c_1328_n 0.00371193f $X=3.4 $Y=1.22 $X2=0 $Y2=0
cc_468 N_CLK_c_548_n N_A_608_74#_c_1328_n 0.00848825f $X=3.485 $Y=1.765 $X2=0
+ $Y2=0
cc_469 CLK N_A_608_74#_c_1328_n 0.0284508f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_470 N_CLK_c_548_n N_A_608_74#_c_1348_n 0.0166039f $X=3.485 $Y=1.765 $X2=0
+ $Y2=0
cc_471 CLK N_A_608_74#_c_1348_n 0.0229055f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_472 N_CLK_c_548_n N_A_608_74#_c_1329_n 0.00173919f $X=3.485 $Y=1.765 $X2=0
+ $Y2=0
cc_473 CLK N_A_608_74#_c_1329_n 0.0161169f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_474 N_CLK_c_547_n N_A_608_74#_c_1330_n 0.00232554f $X=3.4 $Y=1.22 $X2=0 $Y2=0
cc_475 N_CLK_c_548_n N_A_608_74#_c_1330_n 0.00116809f $X=3.485 $Y=1.765 $X2=0
+ $Y2=0
cc_476 CLK N_A_608_74#_c_1330_n 0.00294872f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_477 N_CLK_c_548_n N_VPWR_c_1922_n 0.00417761f $X=3.485 $Y=1.765 $X2=0 $Y2=0
cc_478 N_CLK_c_548_n N_VPWR_c_1923_n 0.00413917f $X=3.485 $Y=1.765 $X2=0 $Y2=0
cc_479 N_CLK_c_548_n N_VPWR_c_1924_n 0.0161989f $X=3.485 $Y=1.765 $X2=0 $Y2=0
cc_480 N_CLK_c_548_n N_VPWR_c_1920_n 0.00822528f $X=3.485 $Y=1.765 $X2=0 $Y2=0
cc_481 N_CLK_c_548_n N_A_290_464#_c_2115_n 0.0160629f $X=3.485 $Y=1.765 $X2=0
+ $Y2=0
cc_482 N_CLK_c_548_n N_A_290_464#_c_2117_n 0.00725214f $X=3.485 $Y=1.765 $X2=0
+ $Y2=0
cc_483 N_CLK_c_547_n N_VGND_c_2318_n 0.00333233f $X=3.4 $Y=1.22 $X2=0 $Y2=0
cc_484 N_CLK_c_547_n N_VGND_c_2319_n 0.00434272f $X=3.4 $Y=1.22 $X2=0 $Y2=0
cc_485 N_CLK_c_547_n N_VGND_c_2320_n 0.00659657f $X=3.4 $Y=1.22 $X2=0 $Y2=0
cc_486 N_CLK_c_548_n N_VGND_c_2320_n 4.20406e-19 $X=3.485 $Y=1.765 $X2=0 $Y2=0
cc_487 CLK N_VGND_c_2320_n 0.0164658f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_488 N_CLK_c_547_n N_VGND_c_2342_n 0.00825771f $X=3.4 $Y=1.22 $X2=0 $Y2=0
cc_489 N_A_795_74#_M1030_g N_A_1185_55#_c_878_n 0.0474535f $X=5.64 $Y=0.615
+ $X2=0 $Y2=0
cc_490 N_A_795_74#_c_613_n N_A_1185_55#_c_885_n 0.00134246f $X=5.645 $Y=2.255
+ $X2=0 $Y2=0
cc_491 N_A_795_74#_c_615_n N_A_1185_55#_c_885_n 0.00598664f $X=6.515 $Y=2.17
+ $X2=0 $Y2=0
cc_492 N_A_795_74#_c_614_n N_A_1185_55#_c_886_n 0.00719195f $X=5.645 $Y=2.895
+ $X2=0 $Y2=0
cc_493 N_A_795_74#_c_615_n N_A_1185_55#_c_886_n 0.0122739f $X=6.515 $Y=2.17
+ $X2=0 $Y2=0
cc_494 N_A_795_74#_c_616_n N_A_1185_55#_c_886_n 0.00352077f $X=6.6 $Y=2.905
+ $X2=0 $Y2=0
cc_495 N_A_795_74#_M1030_g N_A_1185_55#_c_879_n 0.0118644f $X=5.64 $Y=0.615
+ $X2=0 $Y2=0
cc_496 N_A_795_74#_M1030_g N_A_1185_55#_c_880_n 0.00159877f $X=5.64 $Y=0.615
+ $X2=0 $Y2=0
cc_497 N_A_795_74#_c_615_n N_A_1185_55#_c_887_n 0.0138611f $X=6.515 $Y=2.17
+ $X2=0 $Y2=0
cc_498 N_A_795_74#_c_619_n N_A_1185_55#_c_887_n 0.00157945f $X=7.28 $Y=2.905
+ $X2=0 $Y2=0
cc_499 N_A_795_74#_c_620_n N_A_1185_55#_c_887_n 0.0133719f $X=7.365 $Y=1.81
+ $X2=0 $Y2=0
cc_500 N_A_795_74#_M1030_g N_A_1185_55#_c_902_n 5.16138e-19 $X=5.64 $Y=0.615
+ $X2=0 $Y2=0
cc_501 N_A_795_74#_c_615_n N_A_1185_55#_c_888_n 0.0134997f $X=6.515 $Y=2.17
+ $X2=0 $Y2=0
cc_502 N_A_795_74#_c_616_n N_A_1185_55#_c_888_n 0.0337427f $X=6.6 $Y=2.905 $X2=0
+ $Y2=0
cc_503 N_A_795_74#_c_617_n N_A_1185_55#_c_888_n 0.0130106f $X=7.195 $Y=2.99
+ $X2=0 $Y2=0
cc_504 N_A_795_74#_c_619_n N_A_1185_55#_c_888_n 0.0579875f $X=7.28 $Y=2.905
+ $X2=0 $Y2=0
cc_505 N_A_795_74#_c_613_n N_A_1185_55#_c_882_n 0.00116556f $X=5.645 $Y=2.255
+ $X2=0 $Y2=0
cc_506 N_A_795_74#_c_615_n N_A_1185_55#_c_882_n 0.00367368f $X=6.515 $Y=2.17
+ $X2=0 $Y2=0
cc_507 N_A_795_74#_c_601_n N_A_1185_55#_c_882_n 0.0259356f $X=5.565 $Y=1.655
+ $X2=0 $Y2=0
cc_508 N_A_795_74#_c_613_n N_A_1185_55#_c_890_n 0.0130405f $X=5.645 $Y=2.255
+ $X2=0 $Y2=0
cc_509 N_A_795_74#_c_615_n N_A_1185_55#_c_890_n 0.0415848f $X=6.515 $Y=2.17
+ $X2=0 $Y2=0
cc_510 N_A_795_74#_c_601_n N_A_1185_55#_c_890_n 2.48241e-19 $X=5.565 $Y=1.655
+ $X2=0 $Y2=0
cc_511 N_A_795_74#_c_583_n N_A_1185_55#_c_884_n 0.0118644f $X=5.625 $Y=1.35
+ $X2=0 $Y2=0
cc_512 N_A_795_74#_c_601_n N_A_1185_55#_c_884_n 0.00426508f $X=5.565 $Y=1.655
+ $X2=0 $Y2=0
cc_513 N_A_795_74#_c_592_n N_A_991_81#_M1016_d 2.28826e-19 $X=5 $Y=0.34
+ $X2=-0.19 $Y2=-0.245
cc_514 N_A_795_74#_c_595_n N_A_991_81#_M1016_d 0.00589878f $X=5.085 $Y=1.015
+ $X2=-0.19 $Y2=-0.245
cc_515 N_A_795_74#_c_615_n N_A_991_81#_c_980_n 0.00286592f $X=6.515 $Y=2.17
+ $X2=0 $Y2=0
cc_516 N_A_795_74#_c_620_n N_A_991_81#_c_980_n 2.30351e-19 $X=7.365 $Y=1.81
+ $X2=0 $Y2=0
cc_517 N_A_795_74#_c_615_n N_A_991_81#_c_998_n 0.00360333f $X=6.515 $Y=2.17
+ $X2=0 $Y2=0
cc_518 N_A_795_74#_c_616_n N_A_991_81#_c_998_n 0.01539f $X=6.6 $Y=2.905 $X2=0
+ $Y2=0
cc_519 N_A_795_74#_c_617_n N_A_991_81#_c_998_n 0.00295621f $X=7.195 $Y=2.99
+ $X2=0 $Y2=0
cc_520 N_A_795_74#_c_619_n N_A_991_81#_c_998_n 5.81564e-19 $X=7.28 $Y=2.905
+ $X2=0 $Y2=0
cc_521 N_A_795_74#_c_625_n N_A_991_81#_c_982_n 0.00245883f $X=8.255 $Y=1.685
+ $X2=0 $Y2=0
cc_522 N_A_795_74#_c_599_n N_A_991_81#_c_982_n 9.68097e-19 $X=8.425 $Y=1.685
+ $X2=0 $Y2=0
cc_523 N_A_795_74#_c_619_n N_A_991_81#_c_1000_n 0.00389112f $X=7.28 $Y=2.905
+ $X2=0 $Y2=0
cc_524 N_A_795_74#_c_625_n N_A_991_81#_c_1000_n 0.0138785f $X=8.255 $Y=1.685
+ $X2=0 $Y2=0
cc_525 N_A_795_74#_c_625_n N_A_991_81#_c_984_n 0.00132182f $X=8.255 $Y=1.685
+ $X2=0 $Y2=0
cc_526 N_A_795_74#_c_599_n N_A_991_81#_c_984_n 0.00755698f $X=8.425 $Y=1.685
+ $X2=0 $Y2=0
cc_527 N_A_795_74#_c_625_n N_A_991_81#_c_1002_n 0.00331365f $X=8.255 $Y=1.685
+ $X2=0 $Y2=0
cc_528 N_A_795_74#_c_599_n N_A_991_81#_c_1002_n 0.00628952f $X=8.425 $Y=1.685
+ $X2=0 $Y2=0
cc_529 N_A_795_74#_c_605_n N_A_991_81#_c_1003_n 0.00223259f $X=4.975 $Y=2.21
+ $X2=0 $Y2=0
cc_530 N_A_795_74#_c_614_n N_A_991_81#_c_1003_n 0.0302136f $X=5.645 $Y=2.895
+ $X2=0 $Y2=0
cc_531 N_A_795_74#_c_610_n N_A_991_81#_c_1004_n 0.0191543f $X=5.56 $Y=2.98 $X2=0
+ $Y2=0
cc_532 N_A_795_74#_c_583_n N_A_991_81#_c_987_n 0.00423998f $X=5.625 $Y=1.35
+ $X2=0 $Y2=0
cc_533 N_A_795_74#_M1030_g N_A_991_81#_c_987_n 0.0209349f $X=5.64 $Y=0.615 $X2=0
+ $Y2=0
cc_534 N_A_795_74#_c_592_n N_A_991_81#_c_987_n 0.00340526f $X=5 $Y=0.34 $X2=0
+ $Y2=0
cc_535 N_A_795_74#_c_594_n N_A_991_81#_c_987_n 0.00865059f $X=4.875 $Y=1.565
+ $X2=0 $Y2=0
cc_536 N_A_795_74#_c_595_n N_A_991_81#_c_987_n 0.0446184f $X=5.085 $Y=1.015
+ $X2=0 $Y2=0
cc_537 N_A_795_74#_c_598_n N_A_991_81#_c_987_n 0.0139975f $X=5.085 $Y=1.1 $X2=0
+ $Y2=0
cc_538 N_A_795_74#_c_602_n N_A_991_81#_c_987_n 0.0010998f $X=5.565 $Y=1.58 $X2=0
+ $Y2=0
cc_539 N_A_795_74#_c_615_n N_A_991_81#_c_988_n 0.00708192f $X=6.515 $Y=2.17
+ $X2=0 $Y2=0
cc_540 N_A_795_74#_c_601_n N_A_991_81#_c_988_n 4.23483e-19 $X=5.565 $Y=1.655
+ $X2=0 $Y2=0
cc_541 N_A_795_74#_c_602_n N_A_991_81#_c_988_n 0.011013f $X=5.565 $Y=1.58 $X2=0
+ $Y2=0
cc_542 N_A_795_74#_c_582_n N_A_991_81#_c_989_n 0.0114893f $X=5.4 $Y=1.655 $X2=0
+ $Y2=0
cc_543 N_A_795_74#_c_594_n N_A_991_81#_c_989_n 0.0138133f $X=4.875 $Y=1.565
+ $X2=0 $Y2=0
cc_544 N_A_795_74#_c_613_n N_A_991_81#_c_989_n 0.0192633f $X=5.645 $Y=2.255
+ $X2=0 $Y2=0
cc_545 N_A_795_74#_c_598_n N_A_991_81#_c_989_n 0.00243713f $X=5.085 $Y=1.1 $X2=0
+ $Y2=0
cc_546 N_A_795_74#_c_600_n N_A_991_81#_c_989_n 0.00165075f $X=5.065 $Y=1.565
+ $X2=0 $Y2=0
cc_547 N_A_795_74#_c_602_n N_A_991_81#_c_989_n 0.00452136f $X=5.565 $Y=1.58
+ $X2=0 $Y2=0
cc_548 N_A_795_74#_c_604_n N_A_991_81#_c_993_n 0.00708421f $X=4.975 $Y=2.12
+ $X2=0 $Y2=0
cc_549 N_A_795_74#_c_605_n N_A_991_81#_c_993_n 0.00117893f $X=4.975 $Y=2.21
+ $X2=0 $Y2=0
cc_550 N_A_795_74#_c_582_n N_A_991_81#_c_993_n 0.0132701f $X=5.4 $Y=1.655 $X2=0
+ $Y2=0
cc_551 N_A_795_74#_c_594_n N_A_991_81#_c_993_n 0.0128533f $X=4.875 $Y=1.565
+ $X2=0 $Y2=0
cc_552 N_A_795_74#_c_613_n N_A_991_81#_c_993_n 0.0374763f $X=5.645 $Y=2.255
+ $X2=0 $Y2=0
cc_553 N_A_795_74#_c_614_n N_A_991_81#_c_993_n 5.11009e-19 $X=5.645 $Y=2.895
+ $X2=0 $Y2=0
cc_554 N_A_795_74#_c_600_n N_A_991_81#_c_993_n 3.64028e-19 $X=5.065 $Y=1.565
+ $X2=0 $Y2=0
cc_555 N_A_795_74#_c_601_n N_A_991_81#_c_993_n 0.00251116f $X=5.565 $Y=1.655
+ $X2=0 $Y2=0
cc_556 N_A_795_74#_c_602_n N_A_991_81#_c_993_n 7.34463e-19 $X=5.565 $Y=1.58
+ $X2=0 $Y2=0
cc_557 N_A_795_74#_c_625_n N_A_991_81#_c_994_n 0.0235309f $X=8.255 $Y=1.685
+ $X2=0 $Y2=0
cc_558 N_A_795_74#_c_599_n N_A_991_81#_c_994_n 0.00630615f $X=8.425 $Y=1.685
+ $X2=0 $Y2=0
cc_559 N_A_795_74#_c_586_n N_A_991_81#_c_996_n 0.00756279f $X=9.14 $Y=1.16 $X2=0
+ $Y2=0
cc_560 N_A_795_74#_c_597_n N_A_991_81#_c_996_n 0.00836768f $X=8.975 $Y=1.64
+ $X2=0 $Y2=0
cc_561 N_A_795_74#_c_625_n N_A_991_81#_c_996_n 0.00169988f $X=8.255 $Y=1.685
+ $X2=0 $Y2=0
cc_562 N_A_795_74#_c_599_n N_A_991_81#_c_996_n 0.0106947f $X=8.425 $Y=1.685
+ $X2=0 $Y2=0
cc_563 N_A_795_74#_c_603_n N_A_991_81#_c_996_n 0.00558876f $X=8.975 $Y=1.475
+ $X2=0 $Y2=0
cc_564 N_A_795_74#_c_619_n N_SET_B_c_1174_n 0.00635764f $X=7.28 $Y=2.905 $X2=0
+ $Y2=0
cc_565 N_A_795_74#_c_620_n N_SET_B_c_1174_n 0.00775299f $X=7.365 $Y=1.81 $X2=0
+ $Y2=0
cc_566 N_A_795_74#_c_616_n N_SET_B_c_1185_n 5.25527e-19 $X=6.6 $Y=2.905 $X2=0
+ $Y2=0
cc_567 N_A_795_74#_c_617_n N_SET_B_c_1185_n 0.00184087f $X=7.195 $Y=2.99 $X2=0
+ $Y2=0
cc_568 N_A_795_74#_c_619_n N_SET_B_c_1185_n 0.019399f $X=7.28 $Y=2.905 $X2=0
+ $Y2=0
cc_569 N_A_795_74#_c_585_n N_SET_B_c_1177_n 0.00630186f $X=9.625 $Y=1.16 $X2=0
+ $Y2=0
cc_570 N_A_795_74#_c_586_n N_SET_B_c_1177_n 0.00131559f $X=9.14 $Y=1.16 $X2=0
+ $Y2=0
cc_571 N_A_795_74#_c_588_n N_SET_B_c_1177_n 0.00829517f $X=10.055 $Y=1.16 $X2=0
+ $Y2=0
cc_572 N_A_795_74#_c_590_n N_SET_B_c_1177_n 0.00149277f $X=9.7 $Y=1.16 $X2=0
+ $Y2=0
cc_573 N_A_795_74#_c_596_n N_SET_B_c_1177_n 0.00715649f $X=10 $Y=1.64 $X2=0
+ $Y2=0
cc_574 N_A_795_74#_c_597_n N_SET_B_c_1177_n 0.0045015f $X=8.975 $Y=1.64 $X2=0
+ $Y2=0
cc_575 N_A_795_74#_c_623_n N_SET_B_c_1177_n 0.0100687f $X=10.555 $Y=1.97 $X2=0
+ $Y2=0
cc_576 N_A_795_74#_c_625_n N_SET_B_c_1177_n 0.012825f $X=8.255 $Y=1.685 $X2=0
+ $Y2=0
cc_577 N_A_795_74#_c_599_n N_SET_B_c_1177_n 0.0535919f $X=8.425 $Y=1.685 $X2=0
+ $Y2=0
cc_578 N_A_795_74#_c_603_n N_SET_B_c_1177_n 0.0054977f $X=8.975 $Y=1.475 $X2=0
+ $Y2=0
cc_579 N_A_795_74#_c_620_n N_SET_B_c_1178_n 4.20079e-19 $X=7.365 $Y=1.81 $X2=0
+ $Y2=0
cc_580 N_A_795_74#_c_625_n N_SET_B_c_1178_n 0.0022884f $X=8.255 $Y=1.685 $X2=0
+ $Y2=0
cc_581 N_A_795_74#_c_620_n N_SET_B_c_1179_n 0.0126733f $X=7.365 $Y=1.81 $X2=0
+ $Y2=0
cc_582 N_A_795_74#_c_625_n N_SET_B_c_1179_n 0.0134421f $X=8.255 $Y=1.685 $X2=0
+ $Y2=0
cc_583 N_A_795_74#_c_620_n N_SET_B_c_1181_n 5.14458e-19 $X=7.365 $Y=1.81 $X2=0
+ $Y2=0
cc_584 N_A_795_74#_c_625_n N_SET_B_c_1181_n 0.00118211f $X=8.255 $Y=1.685 $X2=0
+ $Y2=0
cc_585 N_A_795_74#_c_591_n N_A_608_74#_M1001_g 0.00163108f $X=4.115 $Y=0.515
+ $X2=0 $Y2=0
cc_586 N_A_795_74#_c_593_n N_A_608_74#_M1001_g 0.00266901f $X=4.2 $Y=0.34 $X2=0
+ $Y2=0
cc_587 N_A_795_74#_c_609_n N_A_608_74#_c_1331_n 0.00110874f $X=4.16 $Y=2.78
+ $X2=0 $Y2=0
cc_588 N_A_795_74#_c_611_n N_A_608_74#_c_1331_n 0.00129759f $X=4.325 $Y=2.98
+ $X2=0 $Y2=0
cc_589 N_A_795_74#_c_594_n N_A_608_74#_c_1318_n 0.00118998f $X=4.875 $Y=1.565
+ $X2=0 $Y2=0
cc_590 N_A_795_74#_c_591_n N_A_608_74#_c_1319_n 0.00102731f $X=4.115 $Y=0.515
+ $X2=0 $Y2=0
cc_591 N_A_795_74#_c_594_n N_A_608_74#_c_1319_n 3.17258e-19 $X=4.875 $Y=1.565
+ $X2=0 $Y2=0
cc_592 N_A_795_74#_c_600_n N_A_608_74#_c_1319_n 0.021129f $X=5.065 $Y=1.565
+ $X2=0 $Y2=0
cc_593 N_A_795_74#_c_605_n N_A_608_74#_c_1333_n 0.0160432f $X=4.975 $Y=2.21
+ $X2=0 $Y2=0
cc_594 N_A_795_74#_c_609_n N_A_608_74#_c_1333_n 0.00596256f $X=4.16 $Y=2.78
+ $X2=0 $Y2=0
cc_595 N_A_795_74#_c_610_n N_A_608_74#_c_1333_n 0.0135194f $X=5.56 $Y=2.98 $X2=0
+ $Y2=0
cc_596 N_A_795_74#_c_594_n N_A_608_74#_c_1320_n 0.0025543f $X=4.875 $Y=1.565
+ $X2=0 $Y2=0
cc_597 N_A_795_74#_c_598_n N_A_608_74#_c_1320_n 0.007948f $X=5.085 $Y=1.1 $X2=0
+ $Y2=0
cc_598 N_A_795_74#_c_600_n N_A_608_74#_c_1320_n 0.0160256f $X=5.065 $Y=1.565
+ $X2=0 $Y2=0
cc_599 N_A_795_74#_c_591_n N_A_608_74#_c_1321_n 8.15047e-19 $X=4.115 $Y=0.515
+ $X2=0 $Y2=0
cc_600 N_A_795_74#_c_592_n N_A_608_74#_c_1321_n 0.00184816f $X=5 $Y=0.34 $X2=0
+ $Y2=0
cc_601 N_A_795_74#_c_605_n N_A_608_74#_c_1334_n 0.00737233f $X=4.975 $Y=2.21
+ $X2=0 $Y2=0
cc_602 N_A_795_74#_c_610_n N_A_608_74#_c_1334_n 0.0183312f $X=5.56 $Y=2.98 $X2=0
+ $Y2=0
cc_603 N_A_795_74#_M1030_g N_A_608_74#_M1016_g 0.00858665f $X=5.64 $Y=0.615
+ $X2=0 $Y2=0
cc_604 N_A_795_74#_c_591_n N_A_608_74#_M1016_g 0.00311369f $X=4.115 $Y=0.515
+ $X2=0 $Y2=0
cc_605 N_A_795_74#_c_592_n N_A_608_74#_M1016_g 0.0136298f $X=5 $Y=0.34 $X2=0
+ $Y2=0
cc_606 N_A_795_74#_c_595_n N_A_608_74#_M1016_g 0.00592452f $X=5.085 $Y=1.015
+ $X2=0 $Y2=0
cc_607 N_A_795_74#_c_598_n N_A_608_74#_M1016_g 0.00464804f $X=5.085 $Y=1.1 $X2=0
+ $Y2=0
cc_608 N_A_795_74#_c_605_n N_A_608_74#_c_1336_n 0.00896831f $X=4.975 $Y=2.21
+ $X2=0 $Y2=0
cc_609 N_A_795_74#_c_610_n N_A_608_74#_c_1336_n 0.00601296f $X=5.56 $Y=2.98
+ $X2=0 $Y2=0
cc_610 N_A_795_74#_c_613_n N_A_608_74#_c_1336_n 6.45027e-19 $X=5.645 $Y=2.255
+ $X2=0 $Y2=0
cc_611 N_A_795_74#_c_614_n N_A_608_74#_c_1336_n 0.01533f $X=5.645 $Y=2.895 $X2=0
+ $Y2=0
cc_612 N_A_795_74#_c_601_n N_A_608_74#_c_1336_n 0.00908613f $X=5.565 $Y=1.655
+ $X2=0 $Y2=0
cc_613 N_A_795_74#_c_610_n N_A_608_74#_c_1337_n 0.00318219f $X=5.56 $Y=2.98
+ $X2=0 $Y2=0
cc_614 N_A_795_74#_c_617_n N_A_608_74#_c_1337_n 0.0119141f $X=7.195 $Y=2.99
+ $X2=0 $Y2=0
cc_615 N_A_795_74#_c_618_n N_A_608_74#_c_1337_n 0.00345098f $X=6.685 $Y=2.99
+ $X2=0 $Y2=0
cc_616 N_A_795_74#_c_596_n N_A_608_74#_c_1323_n 0.0174119f $X=10 $Y=1.64 $X2=0
+ $Y2=0
cc_617 N_A_795_74#_c_597_n N_A_608_74#_c_1323_n 0.0118f $X=8.975 $Y=1.64 $X2=0
+ $Y2=0
cc_618 N_A_795_74#_c_590_n N_A_608_74#_c_1324_n 0.0283254f $X=9.7 $Y=1.16 $X2=0
+ $Y2=0
cc_619 N_A_795_74#_c_596_n N_A_608_74#_c_1324_n 0.0275131f $X=10 $Y=1.64 $X2=0
+ $Y2=0
cc_620 N_A_795_74#_c_623_n N_A_608_74#_c_1324_n 0.00901037f $X=10.555 $Y=1.97
+ $X2=0 $Y2=0
cc_621 N_A_795_74#_c_624_n N_A_608_74#_c_1324_n 0.0199936f $X=10.555 $Y=1.97
+ $X2=0 $Y2=0
cc_622 N_A_795_74#_c_585_n N_A_608_74#_c_1325_n 0.0283254f $X=9.625 $Y=1.16
+ $X2=0 $Y2=0
cc_623 N_A_795_74#_c_596_n N_A_608_74#_c_1325_n 0.0048077f $X=10 $Y=1.64 $X2=0
+ $Y2=0
cc_624 N_A_795_74#_c_603_n N_A_608_74#_c_1325_n 0.0118f $X=8.975 $Y=1.475 $X2=0
+ $Y2=0
cc_625 N_A_795_74#_c_608_n N_A_608_74#_c_1341_n 9.37481e-19 $X=10.63 $Y=2.465
+ $X2=0 $Y2=0
cc_626 N_A_795_74#_c_607_n N_A_608_74#_c_1342_n 0.0066338f $X=10.63 $Y=2.375
+ $X2=0 $Y2=0
cc_627 N_A_795_74#_c_608_n N_A_608_74#_c_1342_n 0.00656463f $X=10.63 $Y=2.465
+ $X2=0 $Y2=0
cc_628 N_A_795_74#_c_596_n N_A_608_74#_c_1342_n 0.0048641f $X=10 $Y=1.64 $X2=0
+ $Y2=0
cc_629 N_A_795_74#_c_624_n N_A_608_74#_c_1342_n 0.00319597f $X=10.555 $Y=1.97
+ $X2=0 $Y2=0
cc_630 N_A_795_74#_c_589_n N_A_608_74#_M1043_g 0.024414f $X=10.13 $Y=1.085 $X2=0
+ $Y2=0
cc_631 N_A_795_74#_c_604_n N_A_608_74#_c_1343_n 0.00663995f $X=4.975 $Y=2.12
+ $X2=0 $Y2=0
cc_632 N_A_795_74#_c_604_n N_A_608_74#_c_1344_n 0.00365891f $X=4.975 $Y=2.12
+ $X2=0 $Y2=0
cc_633 N_A_795_74#_c_610_n N_A_608_74#_c_1345_n 0.0111526f $X=5.56 $Y=2.98 $X2=0
+ $Y2=0
cc_634 N_A_795_74#_M1018_d N_A_608_74#_c_1348_n 0.00397779f $X=4.01 $Y=1.84
+ $X2=0 $Y2=0
cc_635 N_A_795_74#_c_591_n N_A_608_74#_c_1329_n 0.012379f $X=4.115 $Y=0.515
+ $X2=0 $Y2=0
cc_636 N_A_795_74#_c_624_n N_A_2186_367#_c_1532_n 0.0132478f $X=10.555 $Y=1.97
+ $X2=0 $Y2=0
cc_637 N_A_795_74#_c_607_n N_A_2186_367#_c_1533_n 0.0132478f $X=10.63 $Y=2.375
+ $X2=0 $Y2=0
cc_638 N_A_795_74#_c_608_n N_A_2186_367#_c_1534_n 0.0453641f $X=10.63 $Y=2.465
+ $X2=0 $Y2=0
cc_639 N_A_795_74#_c_624_n N_A_2186_367#_c_1524_n 0.00162157f $X=10.555 $Y=1.97
+ $X2=0 $Y2=0
cc_640 N_A_795_74#_c_596_n N_A_1804_424#_M1010_s 0.00459485f $X=10 $Y=1.64 $X2=0
+ $Y2=0
cc_641 N_A_795_74#_c_623_n N_A_1804_424#_M1010_s 7.16172e-19 $X=10.555 $Y=1.97
+ $X2=0 $Y2=0
cc_642 N_A_795_74#_c_608_n N_A_1804_424#_c_1655_n 0.00296585f $X=10.63 $Y=2.465
+ $X2=0 $Y2=0
cc_643 N_A_795_74#_c_587_n N_A_1804_424#_c_1640_n 0.0109156f $X=9.7 $Y=1.085
+ $X2=0 $Y2=0
cc_644 N_A_795_74#_c_589_n N_A_1804_424#_c_1640_n 0.0133206f $X=10.13 $Y=1.085
+ $X2=0 $Y2=0
cc_645 N_A_795_74#_c_608_n N_A_1804_424#_c_1657_n 0.00885362f $X=10.63 $Y=2.465
+ $X2=0 $Y2=0
cc_646 N_A_795_74#_c_589_n N_A_1804_424#_c_1641_n 0.00571513f $X=10.13 $Y=1.085
+ $X2=0 $Y2=0
cc_647 N_A_795_74#_c_596_n N_A_1804_424#_c_1658_n 0.00575761f $X=10 $Y=1.64
+ $X2=0 $Y2=0
cc_648 N_A_795_74#_c_623_n N_A_1804_424#_c_1658_n 0.0230587f $X=10.555 $Y=1.97
+ $X2=0 $Y2=0
cc_649 N_A_795_74#_c_624_n N_A_1804_424#_c_1658_n 0.0010483f $X=10.555 $Y=1.97
+ $X2=0 $Y2=0
cc_650 N_A_795_74#_c_623_n N_A_1804_424#_c_1642_n 0.00705752f $X=10.555 $Y=1.97
+ $X2=0 $Y2=0
cc_651 N_A_795_74#_c_624_n N_A_1804_424#_c_1642_n 8.56578e-19 $X=10.555 $Y=1.97
+ $X2=0 $Y2=0
cc_652 N_A_795_74#_c_596_n N_A_1804_424#_c_1643_n 0.00546536f $X=10 $Y=1.64
+ $X2=0 $Y2=0
cc_653 N_A_795_74#_c_623_n N_A_1804_424#_c_1643_n 0.00959246f $X=10.555 $Y=1.97
+ $X2=0 $Y2=0
cc_654 N_A_795_74#_c_624_n N_A_1804_424#_c_1643_n 5.88732e-19 $X=10.555 $Y=1.97
+ $X2=0 $Y2=0
cc_655 N_A_795_74#_c_623_n N_A_1804_424#_c_1644_n 0.0128867f $X=10.555 $Y=1.97
+ $X2=0 $Y2=0
cc_656 N_A_795_74#_c_624_n N_A_1804_424#_c_1644_n 4.82162e-19 $X=10.555 $Y=1.97
+ $X2=0 $Y2=0
cc_657 N_A_795_74#_c_587_n N_A_1804_424#_c_1647_n 0.00165289f $X=9.7 $Y=1.085
+ $X2=0 $Y2=0
cc_658 N_A_795_74#_c_607_n N_A_1804_424#_c_1663_n 0.00540489f $X=10.63 $Y=2.375
+ $X2=0 $Y2=0
cc_659 N_A_795_74#_c_608_n N_A_1804_424#_c_1663_n 0.00816299f $X=10.63 $Y=2.465
+ $X2=0 $Y2=0
cc_660 N_A_795_74#_c_623_n N_A_1804_424#_c_1663_n 0.0207081f $X=10.555 $Y=1.97
+ $X2=0 $Y2=0
cc_661 N_A_795_74#_c_624_n N_A_1804_424#_c_1663_n 0.00235196f $X=10.555 $Y=1.97
+ $X2=0 $Y2=0
cc_662 N_A_795_74#_c_623_n N_A_1804_424#_c_1664_n 0.014313f $X=10.555 $Y=1.97
+ $X2=0 $Y2=0
cc_663 N_A_795_74#_c_624_n N_A_1804_424#_c_1664_n 0.00520943f $X=10.555 $Y=1.97
+ $X2=0 $Y2=0
cc_664 N_A_795_74#_c_616_n N_VPWR_M1028_d 0.00440946f $X=6.6 $Y=2.905 $X2=0
+ $Y2=0
cc_665 N_A_795_74#_c_619_n N_VPWR_M1029_d 0.00384943f $X=7.28 $Y=2.905 $X2=0
+ $Y2=0
cc_666 N_A_795_74#_c_609_n N_VPWR_c_1924_n 0.021087f $X=4.16 $Y=2.78 $X2=0 $Y2=0
cc_667 N_A_795_74#_c_611_n N_VPWR_c_1924_n 0.0125705f $X=4.325 $Y=2.98 $X2=0
+ $Y2=0
cc_668 N_A_795_74#_c_610_n N_VPWR_c_1925_n 0.00867487f $X=5.56 $Y=2.98 $X2=0
+ $Y2=0
cc_669 N_A_795_74#_c_614_n N_VPWR_c_1925_n 0.0190646f $X=5.645 $Y=2.895 $X2=0
+ $Y2=0
cc_670 N_A_795_74#_c_615_n N_VPWR_c_1925_n 0.017848f $X=6.515 $Y=2.17 $X2=0
+ $Y2=0
cc_671 N_A_795_74#_c_616_n N_VPWR_c_1925_n 0.0363341f $X=6.6 $Y=2.905 $X2=0
+ $Y2=0
cc_672 N_A_795_74#_c_618_n N_VPWR_c_1925_n 0.0147459f $X=6.685 $Y=2.99 $X2=0
+ $Y2=0
cc_673 N_A_795_74#_c_617_n N_VPWR_c_1926_n 0.0143583f $X=7.195 $Y=2.99 $X2=0
+ $Y2=0
cc_674 N_A_795_74#_c_619_n N_VPWR_c_1926_n 0.0617589f $X=7.28 $Y=2.905 $X2=0
+ $Y2=0
cc_675 N_A_795_74#_c_625_n N_VPWR_c_1926_n 0.0138919f $X=8.255 $Y=1.685 $X2=0
+ $Y2=0
cc_676 N_A_795_74#_c_608_n N_VPWR_c_1928_n 0.00136956f $X=10.63 $Y=2.465 $X2=0
+ $Y2=0
cc_677 N_A_795_74#_c_610_n N_VPWR_c_1933_n 0.0853008f $X=5.56 $Y=2.98 $X2=0
+ $Y2=0
cc_678 N_A_795_74#_c_611_n N_VPWR_c_1933_n 0.0164393f $X=4.325 $Y=2.98 $X2=0
+ $Y2=0
cc_679 N_A_795_74#_c_617_n N_VPWR_c_1935_n 0.0443733f $X=7.195 $Y=2.99 $X2=0
+ $Y2=0
cc_680 N_A_795_74#_c_618_n N_VPWR_c_1935_n 0.0115893f $X=6.685 $Y=2.99 $X2=0
+ $Y2=0
cc_681 N_A_795_74#_c_608_n N_VPWR_c_1941_n 0.00461464f $X=10.63 $Y=2.465 $X2=0
+ $Y2=0
cc_682 N_A_795_74#_c_608_n N_VPWR_c_1920_n 0.00470261f $X=10.63 $Y=2.465 $X2=0
+ $Y2=0
cc_683 N_A_795_74#_c_610_n N_VPWR_c_1920_n 0.0470576f $X=5.56 $Y=2.98 $X2=0
+ $Y2=0
cc_684 N_A_795_74#_c_611_n N_VPWR_c_1920_n 0.00958732f $X=4.325 $Y=2.98 $X2=0
+ $Y2=0
cc_685 N_A_795_74#_c_617_n N_VPWR_c_1920_n 0.0229659f $X=7.195 $Y=2.99 $X2=0
+ $Y2=0
cc_686 N_A_795_74#_c_618_n N_VPWR_c_1920_n 0.00583135f $X=6.685 $Y=2.99 $X2=0
+ $Y2=0
cc_687 N_A_795_74#_c_592_n N_A_290_464#_M1016_s 0.00228614f $X=5 $Y=0.34 $X2=0
+ $Y2=0
cc_688 N_A_795_74#_M1018_d N_A_290_464#_c_2115_n 0.00490079f $X=4.01 $Y=1.84
+ $X2=0 $Y2=0
cc_689 N_A_795_74#_c_609_n N_A_290_464#_c_2115_n 0.019779f $X=4.16 $Y=2.78 $X2=0
+ $Y2=0
cc_690 N_A_795_74#_c_610_n N_A_290_464#_c_2115_n 0.00832556f $X=5.56 $Y=2.98
+ $X2=0 $Y2=0
cc_691 N_A_795_74#_c_604_n N_A_290_464#_c_2116_n 0.00120791f $X=4.975 $Y=2.12
+ $X2=0 $Y2=0
cc_692 N_A_795_74#_c_605_n N_A_290_464#_c_2116_n 0.00327424f $X=4.975 $Y=2.21
+ $X2=0 $Y2=0
cc_693 N_A_795_74#_c_591_n N_A_290_464#_c_2111_n 0.0164119f $X=4.115 $Y=0.515
+ $X2=0 $Y2=0
cc_694 N_A_795_74#_c_592_n N_A_290_464#_c_2111_n 0.0249256f $X=5 $Y=0.34 $X2=0
+ $Y2=0
cc_695 N_A_795_74#_c_595_n N_A_290_464#_c_2111_n 0.0103527f $X=5.085 $Y=1.015
+ $X2=0 $Y2=0
cc_696 N_A_795_74#_c_598_n N_A_290_464#_c_2111_n 0.0052363f $X=5.085 $Y=1.1
+ $X2=0 $Y2=0
cc_697 N_A_795_74#_c_604_n N_A_290_464#_c_2112_n 0.00143241f $X=4.975 $Y=2.12
+ $X2=0 $Y2=0
cc_698 N_A_795_74#_c_591_n N_A_290_464#_c_2112_n 0.0171937f $X=4.115 $Y=0.515
+ $X2=0 $Y2=0
cc_699 N_A_795_74#_c_594_n N_A_290_464#_c_2112_n 0.0403116f $X=4.875 $Y=1.565
+ $X2=0 $Y2=0
cc_700 N_A_795_74#_c_595_n N_A_290_464#_c_2112_n 0.00693452f $X=5.085 $Y=1.015
+ $X2=0 $Y2=0
cc_701 N_A_795_74#_c_598_n N_A_290_464#_c_2112_n 0.0124645f $X=5.085 $Y=1.1
+ $X2=0 $Y2=0
cc_702 N_A_795_74#_c_600_n N_A_290_464#_c_2112_n 0.00203394f $X=5.065 $Y=1.565
+ $X2=0 $Y2=0
cc_703 N_A_795_74#_c_604_n N_A_290_464#_c_2119_n 0.00502684f $X=4.975 $Y=2.12
+ $X2=0 $Y2=0
cc_704 N_A_795_74#_c_594_n N_A_290_464#_c_2119_n 0.0132956f $X=4.875 $Y=1.565
+ $X2=0 $Y2=0
cc_705 N_A_795_74#_c_600_n N_A_290_464#_c_2119_n 0.00324793f $X=5.065 $Y=1.565
+ $X2=0 $Y2=0
cc_706 N_A_795_74#_c_605_n N_A_290_464#_c_2120_n 0.00631852f $X=4.975 $Y=2.21
+ $X2=0 $Y2=0
cc_707 N_A_795_74#_c_609_n N_A_290_464#_c_2120_n 0.00878202f $X=4.16 $Y=2.78
+ $X2=0 $Y2=0
cc_708 N_A_795_74#_c_610_n N_A_290_464#_c_2120_n 0.0259128f $X=5.56 $Y=2.98
+ $X2=0 $Y2=0
cc_709 N_A_795_74#_c_614_n A_1117_483# 0.006138f $X=5.645 $Y=2.895 $X2=-0.19
+ $Y2=-0.245
cc_710 N_A_795_74#_c_596_n N_A_1584_379#_c_2244_n 0.00969718f $X=10 $Y=1.64
+ $X2=0 $Y2=0
cc_711 N_A_795_74#_c_625_n N_A_1584_379#_c_2244_n 0.0120374f $X=8.255 $Y=1.685
+ $X2=0 $Y2=0
cc_712 N_A_795_74#_c_596_n N_A_1584_379#_c_2241_n 0.0948999f $X=10 $Y=1.64 $X2=0
+ $Y2=0
cc_713 N_A_795_74#_c_597_n N_A_1584_379#_c_2241_n 0.00798977f $X=8.975 $Y=1.64
+ $X2=0 $Y2=0
cc_714 N_A_795_74#_c_625_n N_A_1584_379#_c_2242_n 0.0219119f $X=8.255 $Y=1.685
+ $X2=0 $Y2=0
cc_715 N_A_795_74#_c_596_n N_A_1584_379#_c_2243_n 0.0134175f $X=10 $Y=1.64 $X2=0
+ $Y2=0
cc_716 N_A_795_74#_c_593_n N_VGND_c_2320_n 0.0112234f $X=4.2 $Y=0.34 $X2=0 $Y2=0
cc_717 N_A_795_74#_c_587_n N_VGND_c_2322_n 3.14208e-19 $X=9.7 $Y=1.085 $X2=0
+ $Y2=0
cc_718 N_A_795_74#_M1030_g N_VGND_c_2327_n 0.00527282f $X=5.64 $Y=0.615 $X2=0
+ $Y2=0
cc_719 N_A_795_74#_c_592_n N_VGND_c_2327_n 0.0636631f $X=5 $Y=0.34 $X2=0 $Y2=0
cc_720 N_A_795_74#_c_593_n N_VGND_c_2327_n 0.0121867f $X=4.2 $Y=0.34 $X2=0 $Y2=0
cc_721 N_A_795_74#_c_587_n N_VGND_c_2339_n 0.00278271f $X=9.7 $Y=1.085 $X2=0
+ $Y2=0
cc_722 N_A_795_74#_c_589_n N_VGND_c_2339_n 0.00278271f $X=10.13 $Y=1.085 $X2=0
+ $Y2=0
cc_723 N_A_795_74#_M1030_g N_VGND_c_2342_n 0.00534666f $X=5.64 $Y=0.615 $X2=0
+ $Y2=0
cc_724 N_A_795_74#_c_587_n N_VGND_c_2342_n 0.00358427f $X=9.7 $Y=1.085 $X2=0
+ $Y2=0
cc_725 N_A_795_74#_c_589_n N_VGND_c_2342_n 0.0035414f $X=10.13 $Y=1.085 $X2=0
+ $Y2=0
cc_726 N_A_795_74#_c_592_n N_VGND_c_2342_n 0.0366794f $X=5 $Y=0.34 $X2=0 $Y2=0
cc_727 N_A_795_74#_c_593_n N_VGND_c_2342_n 0.00660921f $X=4.2 $Y=0.34 $X2=0
+ $Y2=0
cc_728 N_A_795_74#_c_586_n N_A_1641_74#_c_2480_n 0.0178304f $X=9.14 $Y=1.16
+ $X2=0 $Y2=0
cc_729 N_A_795_74#_c_587_n N_A_1641_74#_c_2480_n 0.0116182f $X=9.7 $Y=1.085
+ $X2=0 $Y2=0
cc_730 N_A_795_74#_c_596_n N_A_1641_74#_c_2480_n 0.0233474f $X=10 $Y=1.64 $X2=0
+ $Y2=0
cc_731 N_A_795_74#_c_597_n N_A_1641_74#_c_2480_n 0.00335664f $X=8.975 $Y=1.64
+ $X2=0 $Y2=0
cc_732 N_A_795_74#_c_625_n N_A_1641_74#_c_2481_n 8.07173e-19 $X=8.255 $Y=1.685
+ $X2=0 $Y2=0
cc_733 N_A_795_74#_c_599_n N_A_1641_74#_c_2481_n 0.00555546f $X=8.425 $Y=1.685
+ $X2=0 $Y2=0
cc_734 N_A_795_74#_c_587_n N_A_1641_74#_c_2482_n 0.0110826f $X=9.7 $Y=1.085
+ $X2=0 $Y2=0
cc_735 N_A_795_74#_c_588_n N_A_1641_74#_c_2482_n 0.0027829f $X=10.055 $Y=1.16
+ $X2=0 $Y2=0
cc_736 N_A_795_74#_c_589_n N_A_1641_74#_c_2482_n 0.00708563f $X=10.13 $Y=1.085
+ $X2=0 $Y2=0
cc_737 N_A_795_74#_c_596_n N_A_1641_74#_c_2482_n 0.00654828f $X=10 $Y=1.64 $X2=0
+ $Y2=0
cc_738 N_A_1185_55#_c_887_n N_A_991_81#_c_979_n 0.00105699f $X=6.855 $Y=1.83
+ $X2=0 $Y2=0
cc_739 N_A_1185_55#_c_885_n N_A_991_81#_c_980_n 0.00305319f $X=6.03 $Y=2.15
+ $X2=0 $Y2=0
cc_740 N_A_1185_55#_c_887_n N_A_991_81#_c_980_n 0.0154198f $X=6.855 $Y=1.83
+ $X2=0 $Y2=0
cc_741 N_A_1185_55#_c_888_n N_A_991_81#_c_980_n 0.00536521f $X=6.94 $Y=2.515
+ $X2=0 $Y2=0
cc_742 N_A_1185_55#_c_882_n N_A_991_81#_c_980_n 0.0120011f $X=6.105 $Y=1.815
+ $X2=0 $Y2=0
cc_743 N_A_1185_55#_c_884_n N_A_991_81#_c_980_n 0.00242176f $X=6.105 $Y=1.65
+ $X2=0 $Y2=0
cc_744 N_A_1185_55#_c_886_n N_A_991_81#_c_998_n 0.0107021f $X=6.03 $Y=2.24 $X2=0
+ $Y2=0
cc_745 N_A_1185_55#_c_888_n N_A_991_81#_c_998_n 0.00186053f $X=6.94 $Y=2.515
+ $X2=0 $Y2=0
cc_746 N_A_1185_55#_c_880_n N_A_991_81#_c_981_n 0.00338254f $X=6.145 $Y=1.1
+ $X2=0 $Y2=0
cc_747 N_A_1185_55#_c_883_n N_A_991_81#_c_981_n 0.00677096f $X=6.855 $Y=0.525
+ $X2=0 $Y2=0
cc_748 N_A_1185_55#_c_878_n N_A_991_81#_c_986_n 0.00146983f $X=6 $Y=0.935 $X2=0
+ $Y2=0
cc_749 N_A_1185_55#_c_879_n N_A_991_81#_c_986_n 0.0177504f $X=6.055 $Y=1.265
+ $X2=0 $Y2=0
cc_750 N_A_1185_55#_c_880_n N_A_991_81#_c_986_n 5.30688e-19 $X=6.145 $Y=1.1
+ $X2=0 $Y2=0
cc_751 N_A_1185_55#_c_881_n N_A_991_81#_c_986_n 0.00370147f $X=6.69 $Y=0.615
+ $X2=0 $Y2=0
cc_752 N_A_1185_55#_c_883_n N_A_991_81#_c_986_n 0.00718643f $X=6.855 $Y=0.525
+ $X2=0 $Y2=0
cc_753 N_A_1185_55#_c_878_n N_A_991_81#_c_987_n 0.00224758f $X=6 $Y=0.935 $X2=0
+ $Y2=0
cc_754 N_A_1185_55#_c_879_n N_A_991_81#_c_987_n 0.00123351f $X=6.055 $Y=1.265
+ $X2=0 $Y2=0
cc_755 N_A_1185_55#_c_880_n N_A_991_81#_c_987_n 0.0189782f $X=6.145 $Y=1.1 $X2=0
+ $Y2=0
cc_756 N_A_1185_55#_c_902_n N_A_991_81#_c_987_n 0.00682346f $X=6.31 $Y=0.615
+ $X2=0 $Y2=0
cc_757 N_A_1185_55#_c_879_n N_A_991_81#_c_988_n 0.00359104f $X=6.055 $Y=1.265
+ $X2=0 $Y2=0
cc_758 N_A_1185_55#_c_880_n N_A_991_81#_c_988_n 0.0256385f $X=6.145 $Y=1.1 $X2=0
+ $Y2=0
cc_759 N_A_1185_55#_c_887_n N_A_991_81#_c_988_n 0.0441129f $X=6.855 $Y=1.83
+ $X2=0 $Y2=0
cc_760 N_A_1185_55#_c_881_n N_A_991_81#_c_988_n 0.0066704f $X=6.69 $Y=0.615
+ $X2=0 $Y2=0
cc_761 N_A_1185_55#_c_882_n N_A_991_81#_c_988_n 0.00167546f $X=6.105 $Y=1.815
+ $X2=0 $Y2=0
cc_762 N_A_1185_55#_c_890_n N_A_991_81#_c_988_n 0.0233235f $X=6.27 $Y=1.815
+ $X2=0 $Y2=0
cc_763 N_A_1185_55#_c_884_n N_A_991_81#_c_988_n 0.0111257f $X=6.105 $Y=1.65
+ $X2=0 $Y2=0
cc_764 N_A_1185_55#_c_879_n N_A_991_81#_c_1083_n 0.00103048f $X=6.055 $Y=1.265
+ $X2=0 $Y2=0
cc_765 N_A_1185_55#_c_880_n N_A_991_81#_c_1083_n 0.00937167f $X=6.145 $Y=1.1
+ $X2=0 $Y2=0
cc_766 N_A_1185_55#_c_884_n N_A_991_81#_c_1083_n 6.17268e-19 $X=6.105 $Y=1.65
+ $X2=0 $Y2=0
cc_767 N_A_1185_55#_c_880_n N_A_991_81#_c_990_n 6.07444e-19 $X=6.145 $Y=1.1
+ $X2=0 $Y2=0
cc_768 N_A_1185_55#_c_884_n N_A_991_81#_c_990_n 0.00843579f $X=6.105 $Y=1.65
+ $X2=0 $Y2=0
cc_769 N_A_1185_55#_c_883_n N_A_991_81#_c_991_n 0.00793363f $X=6.855 $Y=0.525
+ $X2=0 $Y2=0
cc_770 N_A_1185_55#_c_879_n N_A_991_81#_c_992_n 3.96639e-19 $X=6.055 $Y=1.265
+ $X2=0 $Y2=0
cc_771 N_A_1185_55#_c_880_n N_A_991_81#_c_992_n 0.0105303f $X=6.145 $Y=1.1 $X2=0
+ $Y2=0
cc_772 N_A_1185_55#_c_881_n N_A_991_81#_c_992_n 0.0112142f $X=6.69 $Y=0.615
+ $X2=0 $Y2=0
cc_773 N_A_1185_55#_c_883_n N_A_991_81#_c_992_n 0.0157846f $X=6.855 $Y=0.525
+ $X2=0 $Y2=0
cc_774 N_A_1185_55#_c_885_n N_A_991_81#_c_993_n 5.64443e-19 $X=6.03 $Y=2.15
+ $X2=0 $Y2=0
cc_775 N_A_1185_55#_c_882_n N_A_991_81#_c_993_n 2.0933e-19 $X=6.105 $Y=1.815
+ $X2=0 $Y2=0
cc_776 N_A_1185_55#_c_884_n N_A_991_81#_c_993_n 2.07566e-19 $X=6.105 $Y=1.65
+ $X2=0 $Y2=0
cc_777 N_A_1185_55#_c_887_n N_SET_B_c_1174_n 0.00136415f $X=6.855 $Y=1.83 $X2=0
+ $Y2=0
cc_778 N_A_1185_55#_c_888_n N_SET_B_c_1174_n 0.00228039f $X=6.94 $Y=2.515 $X2=0
+ $Y2=0
cc_779 N_A_1185_55#_c_888_n N_SET_B_c_1185_n 0.00169589f $X=6.94 $Y=2.515 $X2=0
+ $Y2=0
cc_780 N_A_1185_55#_c_883_n N_SET_B_M1021_g 0.00103321f $X=6.855 $Y=0.525 $X2=0
+ $Y2=0
cc_781 N_A_1185_55#_c_886_n N_A_608_74#_c_1336_n 0.0161779f $X=6.03 $Y=2.24
+ $X2=0 $Y2=0
cc_782 N_A_1185_55#_c_886_n N_A_608_74#_c_1337_n 0.010379f $X=6.03 $Y=2.24 $X2=0
+ $Y2=0
cc_783 N_A_1185_55#_c_886_n N_VPWR_c_1925_n 0.00802868f $X=6.03 $Y=2.24 $X2=0
+ $Y2=0
cc_784 N_A_1185_55#_c_886_n N_VPWR_c_1920_n 8.82885e-19 $X=6.03 $Y=2.24 $X2=0
+ $Y2=0
cc_785 N_A_1185_55#_c_880_n N_VGND_M1007_d 0.00256846f $X=6.145 $Y=1.1 $X2=0
+ $Y2=0
cc_786 N_A_1185_55#_c_881_n N_VGND_M1007_d 0.00518446f $X=6.69 $Y=0.615 $X2=0
+ $Y2=0
cc_787 N_A_1185_55#_c_902_n N_VGND_M1007_d 0.00235471f $X=6.31 $Y=0.615 $X2=0
+ $Y2=0
cc_788 N_A_1185_55#_c_883_n N_VGND_c_2321_n 0.0107976f $X=6.855 $Y=0.525 $X2=0
+ $Y2=0
cc_789 N_A_1185_55#_c_878_n N_VGND_c_2326_n 0.00357449f $X=6 $Y=0.935 $X2=0
+ $Y2=0
cc_790 N_A_1185_55#_c_879_n N_VGND_c_2326_n 5.89315e-19 $X=6.055 $Y=1.265 $X2=0
+ $Y2=0
cc_791 N_A_1185_55#_c_881_n N_VGND_c_2326_n 0.0109664f $X=6.69 $Y=0.615 $X2=0
+ $Y2=0
cc_792 N_A_1185_55#_c_902_n N_VGND_c_2326_n 0.0144987f $X=6.31 $Y=0.615 $X2=0
+ $Y2=0
cc_793 N_A_1185_55#_c_883_n N_VGND_c_2326_n 6.74191e-19 $X=6.855 $Y=0.525 $X2=0
+ $Y2=0
cc_794 N_A_1185_55#_c_878_n N_VGND_c_2327_n 0.00463637f $X=6 $Y=0.935 $X2=0
+ $Y2=0
cc_795 N_A_1185_55#_c_902_n N_VGND_c_2327_n 0.00291775f $X=6.31 $Y=0.615 $X2=0
+ $Y2=0
cc_796 N_A_1185_55#_c_881_n N_VGND_c_2330_n 0.00533357f $X=6.69 $Y=0.615 $X2=0
+ $Y2=0
cc_797 N_A_1185_55#_c_883_n N_VGND_c_2330_n 0.0138937f $X=6.855 $Y=0.525 $X2=0
+ $Y2=0
cc_798 N_A_1185_55#_c_878_n N_VGND_c_2342_n 0.00534666f $X=6 $Y=0.935 $X2=0
+ $Y2=0
cc_799 N_A_1185_55#_c_881_n N_VGND_c_2342_n 0.00799229f $X=6.69 $Y=0.615 $X2=0
+ $Y2=0
cc_800 N_A_1185_55#_c_902_n N_VGND_c_2342_n 0.00597722f $X=6.31 $Y=0.615 $X2=0
+ $Y2=0
cc_801 N_A_1185_55#_c_883_n N_VGND_c_2342_n 0.0117406f $X=6.855 $Y=0.525 $X2=0
+ $Y2=0
cc_802 N_A_991_81#_c_979_n N_SET_B_c_1174_n 0.00926619f $X=6.715 $Y=1.57 $X2=0
+ $Y2=0
cc_803 N_A_991_81#_c_980_n N_SET_B_c_1174_n 0.0119061f $X=6.715 $Y=2.15 $X2=0
+ $Y2=0
cc_804 N_A_991_81#_c_982_n N_SET_B_c_1174_n 0.00782167f $X=7.845 $Y=1.73 $X2=0
+ $Y2=0
cc_805 N_A_991_81#_c_1000_n N_SET_B_c_1174_n 0.00665068f $X=7.845 $Y=1.82 $X2=0
+ $Y2=0
cc_806 N_A_991_81#_c_998_n N_SET_B_c_1185_n 0.0186157f $X=6.715 $Y=2.24 $X2=0
+ $Y2=0
cc_807 N_A_991_81#_c_1000_n N_SET_B_c_1185_n 0.00730731f $X=7.845 $Y=1.82 $X2=0
+ $Y2=0
cc_808 N_A_991_81#_c_981_n N_SET_B_M1021_g 0.040881f $X=7.07 $Y=0.865 $X2=0
+ $Y2=0
cc_809 N_A_991_81#_c_983_n N_SET_B_M1021_g 0.0171965f $X=8.13 $Y=1.085 $X2=0
+ $Y2=0
cc_810 N_A_991_81#_c_1083_n N_SET_B_M1021_g 8.84629e-19 $X=6.715 $Y=1.065 $X2=0
+ $Y2=0
cc_811 N_A_991_81#_c_990_n N_SET_B_M1021_g 0.00513936f $X=6.715 $Y=1.065 $X2=0
+ $Y2=0
cc_812 N_A_991_81#_c_991_n N_SET_B_M1021_g 0.0146456f $X=7.755 $Y=0.955 $X2=0
+ $Y2=0
cc_813 N_A_991_81#_c_995_n N_SET_B_M1021_g 0.00367161f $X=7.92 $Y=1.225 $X2=0
+ $Y2=0
cc_814 N_A_991_81#_c_991_n N_SET_B_c_1177_n 0.00755992f $X=7.755 $Y=0.955 $X2=0
+ $Y2=0
cc_815 N_A_991_81#_c_994_n N_SET_B_c_1177_n 0.0202042f $X=7.92 $Y=1.39 $X2=0
+ $Y2=0
cc_816 N_A_991_81#_c_996_n N_SET_B_c_1177_n 0.0182276f $X=8.295 $Y=1.32 $X2=0
+ $Y2=0
cc_817 N_A_991_81#_c_988_n N_SET_B_c_1178_n 2.14175e-19 $X=6.55 $Y=1.46 $X2=0
+ $Y2=0
cc_818 N_A_991_81#_c_1083_n N_SET_B_c_1178_n 0.0020303f $X=6.715 $Y=1.065 $X2=0
+ $Y2=0
cc_819 N_A_991_81#_c_990_n N_SET_B_c_1178_n 4.38236e-19 $X=6.715 $Y=1.065 $X2=0
+ $Y2=0
cc_820 N_A_991_81#_c_991_n N_SET_B_c_1178_n 0.00823128f $X=7.755 $Y=0.955 $X2=0
+ $Y2=0
cc_821 N_A_991_81#_c_994_n N_SET_B_c_1178_n 0.00130449f $X=7.92 $Y=1.39 $X2=0
+ $Y2=0
cc_822 N_A_991_81#_c_995_n N_SET_B_c_1178_n 0.00189718f $X=7.92 $Y=1.225 $X2=0
+ $Y2=0
cc_823 N_A_991_81#_c_996_n N_SET_B_c_1178_n 7.09844e-19 $X=8.295 $Y=1.32 $X2=0
+ $Y2=0
cc_824 N_A_991_81#_c_988_n N_SET_B_c_1179_n 0.0082709f $X=6.55 $Y=1.46 $X2=0
+ $Y2=0
cc_825 N_A_991_81#_c_1083_n N_SET_B_c_1179_n 0.00638026f $X=6.715 $Y=1.065 $X2=0
+ $Y2=0
cc_826 N_A_991_81#_c_990_n N_SET_B_c_1179_n 8.13904e-19 $X=6.715 $Y=1.065 $X2=0
+ $Y2=0
cc_827 N_A_991_81#_c_991_n N_SET_B_c_1179_n 0.0233965f $X=7.755 $Y=0.955 $X2=0
+ $Y2=0
cc_828 N_A_991_81#_c_995_n N_SET_B_c_1179_n 0.0216481f $X=7.92 $Y=1.225 $X2=0
+ $Y2=0
cc_829 N_A_991_81#_c_996_n N_SET_B_c_1179_n 0.00178299f $X=8.295 $Y=1.32 $X2=0
+ $Y2=0
cc_830 N_A_991_81#_c_986_n N_SET_B_c_1181_n 0.00166756f $X=7.07 $Y=0.94 $X2=0
+ $Y2=0
cc_831 N_A_991_81#_c_988_n N_SET_B_c_1181_n 8.22009e-19 $X=6.55 $Y=1.46 $X2=0
+ $Y2=0
cc_832 N_A_991_81#_c_1083_n N_SET_B_c_1181_n 6.05847e-19 $X=6.715 $Y=1.065 $X2=0
+ $Y2=0
cc_833 N_A_991_81#_c_990_n N_SET_B_c_1181_n 0.00926619f $X=6.715 $Y=1.065 $X2=0
+ $Y2=0
cc_834 N_A_991_81#_c_991_n N_SET_B_c_1181_n 0.00420665f $X=7.755 $Y=0.955 $X2=0
+ $Y2=0
cc_835 N_A_991_81#_c_994_n N_SET_B_c_1181_n 4.93533e-19 $X=7.92 $Y=1.39 $X2=0
+ $Y2=0
cc_836 N_A_991_81#_c_996_n N_SET_B_c_1181_n 0.0209248f $X=8.295 $Y=1.32 $X2=0
+ $Y2=0
cc_837 N_A_991_81#_c_987_n N_A_608_74#_M1016_g 0.00148512f $X=5.425 $Y=0.615
+ $X2=0 $Y2=0
cc_838 N_A_991_81#_c_1003_n N_A_608_74#_c_1336_n 0.00382716f $X=5.24 $Y=2.39
+ $X2=0 $Y2=0
cc_839 N_A_991_81#_c_998_n N_A_608_74#_c_1337_n 0.00909901f $X=6.715 $Y=2.24
+ $X2=0 $Y2=0
cc_840 N_A_991_81#_c_1000_n N_A_608_74#_c_1337_n 0.0103487f $X=7.845 $Y=1.82
+ $X2=0 $Y2=0
cc_841 N_A_991_81#_c_1002_n N_A_608_74#_c_1337_n 0.0103487f $X=8.295 $Y=1.82
+ $X2=0 $Y2=0
cc_842 N_A_991_81#_c_1002_n N_A_1804_424#_c_1654_n 0.00277632f $X=8.295 $Y=1.82
+ $X2=0 $Y2=0
cc_843 N_A_991_81#_c_998_n N_VPWR_c_1925_n 0.00131022f $X=6.715 $Y=2.24 $X2=0
+ $Y2=0
cc_844 N_A_991_81#_c_1000_n N_VPWR_c_1926_n 0.00516552f $X=7.845 $Y=1.82 $X2=0
+ $Y2=0
cc_845 N_A_991_81#_c_1002_n N_VPWR_c_1927_n 0.00600682f $X=8.295 $Y=1.82 $X2=0
+ $Y2=0
cc_846 N_A_991_81#_c_1000_n N_VPWR_c_1920_n 9.39239e-19 $X=7.845 $Y=1.82 $X2=0
+ $Y2=0
cc_847 N_A_991_81#_c_1002_n N_VPWR_c_1920_n 9.39239e-19 $X=8.295 $Y=1.82 $X2=0
+ $Y2=0
cc_848 N_A_991_81#_c_993_n N_A_290_464#_c_2112_n 0.00564118f $X=5.24 $Y=2.265
+ $X2=0 $Y2=0
cc_849 N_A_991_81#_c_993_n N_A_290_464#_c_2119_n 0.0227835f $X=5.24 $Y=2.265
+ $X2=0 $Y2=0
cc_850 N_A_991_81#_c_1003_n N_A_290_464#_c_2120_n 0.0308684f $X=5.24 $Y=2.39
+ $X2=0 $Y2=0
cc_851 N_A_991_81#_c_1002_n N_A_1584_379#_c_2244_n 0.0128373f $X=8.295 $Y=1.82
+ $X2=0 $Y2=0
cc_852 N_A_991_81#_c_1000_n N_A_1584_379#_c_2242_n 0.00775148f $X=7.845 $Y=1.82
+ $X2=0 $Y2=0
cc_853 N_A_991_81#_c_1002_n N_A_1584_379#_c_2242_n 0.0117861f $X=8.295 $Y=1.82
+ $X2=0 $Y2=0
cc_854 N_A_991_81#_c_1002_n N_A_1584_379#_c_2243_n 0.00364232f $X=8.295 $Y=1.82
+ $X2=0 $Y2=0
cc_855 N_A_991_81#_c_991_n N_VGND_M1021_d 0.00373864f $X=7.755 $Y=0.955 $X2=0
+ $Y2=0
cc_856 N_A_991_81#_c_981_n N_VGND_c_2321_n 0.00149046f $X=7.07 $Y=0.865 $X2=0
+ $Y2=0
cc_857 N_A_991_81#_c_983_n N_VGND_c_2321_n 0.00600886f $X=8.13 $Y=1.085 $X2=0
+ $Y2=0
cc_858 N_A_991_81#_c_991_n N_VGND_c_2321_n 0.0290793f $X=7.755 $Y=0.955 $X2=0
+ $Y2=0
cc_859 N_A_991_81#_c_994_n N_VGND_c_2321_n 0.00136564f $X=7.92 $Y=1.39 $X2=0
+ $Y2=0
cc_860 N_A_991_81#_c_996_n N_VGND_c_2321_n 0.0011328f $X=8.295 $Y=1.32 $X2=0
+ $Y2=0
cc_861 N_A_991_81#_c_985_n N_VGND_c_2322_n 0.011645f $X=8.56 $Y=1.085 $X2=0
+ $Y2=0
cc_862 N_A_991_81#_c_981_n N_VGND_c_2326_n 0.00277351f $X=7.07 $Y=0.865 $X2=0
+ $Y2=0
cc_863 N_A_991_81#_c_987_n N_VGND_c_2327_n 0.00963155f $X=5.425 $Y=0.615 $X2=0
+ $Y2=0
cc_864 N_A_991_81#_c_981_n N_VGND_c_2330_n 0.00434272f $X=7.07 $Y=0.865 $X2=0
+ $Y2=0
cc_865 N_A_991_81#_c_983_n N_VGND_c_2331_n 0.00434272f $X=8.13 $Y=1.085 $X2=0
+ $Y2=0
cc_866 N_A_991_81#_c_985_n N_VGND_c_2331_n 0.00434272f $X=8.56 $Y=1.085 $X2=0
+ $Y2=0
cc_867 N_A_991_81#_c_981_n N_VGND_c_2342_n 0.00825979f $X=7.07 $Y=0.865 $X2=0
+ $Y2=0
cc_868 N_A_991_81#_c_983_n N_VGND_c_2342_n 0.00821975f $X=8.13 $Y=1.085 $X2=0
+ $Y2=0
cc_869 N_A_991_81#_c_985_n N_VGND_c_2342_n 0.00825283f $X=8.56 $Y=1.085 $X2=0
+ $Y2=0
cc_870 N_A_991_81#_c_987_n N_VGND_c_2342_n 0.00894247f $X=5.425 $Y=0.615 $X2=0
+ $Y2=0
cc_871 N_A_991_81#_c_983_n N_A_1641_74#_c_2479_n 0.00822305f $X=8.13 $Y=1.085
+ $X2=0 $Y2=0
cc_872 N_A_991_81#_c_985_n N_A_1641_74#_c_2479_n 0.0117724f $X=8.56 $Y=1.085
+ $X2=0 $Y2=0
cc_873 N_A_991_81#_c_991_n N_A_1641_74#_c_2479_n 8.79632e-19 $X=7.755 $Y=0.955
+ $X2=0 $Y2=0
cc_874 N_A_991_81#_c_985_n N_A_1641_74#_c_2480_n 0.0131495f $X=8.56 $Y=1.085
+ $X2=0 $Y2=0
cc_875 N_A_991_81#_c_983_n N_A_1641_74#_c_2481_n 0.00329746f $X=8.13 $Y=1.085
+ $X2=0 $Y2=0
cc_876 N_A_991_81#_c_985_n N_A_1641_74#_c_2481_n 0.00126919f $X=8.56 $Y=1.085
+ $X2=0 $Y2=0
cc_877 N_A_991_81#_c_991_n N_A_1641_74#_c_2481_n 0.00995113f $X=7.755 $Y=0.955
+ $X2=0 $Y2=0
cc_878 N_A_991_81#_c_995_n N_A_1641_74#_c_2481_n 8.54269e-19 $X=7.92 $Y=1.225
+ $X2=0 $Y2=0
cc_879 N_A_991_81#_c_996_n N_A_1641_74#_c_2481_n 0.00362919f $X=8.295 $Y=1.32
+ $X2=0 $Y2=0
cc_880 N_SET_B_c_1185_n N_A_608_74#_c_1337_n 0.00937227f $X=7.21 $Y=2.24 $X2=0
+ $Y2=0
cc_881 N_SET_B_c_1177_n N_A_608_74#_c_1325_n 0.0158456f $X=11.615 $Y=1.295 $X2=0
+ $Y2=0
cc_882 N_SET_B_c_1177_n N_A_608_74#_M1043_g 0.00705218f $X=11.615 $Y=1.295 $X2=0
+ $Y2=0
cc_883 N_SET_B_c_1186_n N_A_2186_367#_c_1532_n 0.0153072f $X=11.47 $Y=2.375
+ $X2=0 $Y2=0
cc_884 N_SET_B_c_1187_n N_A_2186_367#_c_1533_n 0.0153072f $X=11.47 $Y=2.465
+ $X2=0 $Y2=0
cc_885 N_SET_B_c_1187_n N_A_2186_367#_c_1534_n 0.0111168f $X=11.47 $Y=2.465
+ $X2=0 $Y2=0
cc_886 N_SET_B_M1017_g N_A_2186_367#_c_1524_n 0.00666993f $X=11.59 $Y=0.58 $X2=0
+ $Y2=0
cc_887 N_SET_B_c_1177_n N_A_2186_367#_c_1524_n 0.0036981f $X=11.615 $Y=1.295
+ $X2=0 $Y2=0
cc_888 N_SET_B_c_1182_n N_A_2186_367#_c_1524_n 0.0153072f $X=11.61 $Y=1.635
+ $X2=0 $Y2=0
cc_889 N_SET_B_c_1183_n N_A_2186_367#_c_1524_n 0.00416418f $X=11.76 $Y=1.295
+ $X2=0 $Y2=0
cc_890 N_SET_B_M1017_g N_A_2186_367#_c_1525_n 0.0131197f $X=11.59 $Y=0.58 $X2=0
+ $Y2=0
cc_891 N_SET_B_c_1177_n N_A_2186_367#_c_1525_n 0.00814774f $X=11.615 $Y=1.295
+ $X2=0 $Y2=0
cc_892 SET_B N_A_2186_367#_c_1525_n 0.00328346f $X=11.675 $Y=1.21 $X2=0 $Y2=0
cc_893 N_SET_B_c_1182_n N_A_2186_367#_c_1525_n 0.00258236f $X=11.61 $Y=1.635
+ $X2=0 $Y2=0
cc_894 N_SET_B_c_1183_n N_A_2186_367#_c_1525_n 0.0230245f $X=11.76 $Y=1.295
+ $X2=0 $Y2=0
cc_895 N_SET_B_c_1187_n N_A_2186_367#_c_1536_n 9.87289e-19 $X=11.47 $Y=2.465
+ $X2=0 $Y2=0
cc_896 N_SET_B_c_1186_n N_A_2186_367#_c_1538_n 6.54635e-19 $X=11.47 $Y=2.375
+ $X2=0 $Y2=0
cc_897 N_SET_B_M1017_g N_A_2186_367#_c_1528_n 0.00164729f $X=11.59 $Y=0.58 $X2=0
+ $Y2=0
cc_898 N_SET_B_c_1177_n N_A_2186_367#_c_1528_n 0.0202739f $X=11.615 $Y=1.295
+ $X2=0 $Y2=0
cc_899 SET_B N_A_2186_367#_c_1528_n 2.21379e-19 $X=11.675 $Y=1.21 $X2=0 $Y2=0
cc_900 N_SET_B_c_1183_n N_A_2186_367#_c_1528_n 0.00377693f $X=11.76 $Y=1.295
+ $X2=0 $Y2=0
cc_901 N_SET_B_M1017_g N_A_2186_367#_c_1529_n 0.0182312f $X=11.59 $Y=0.58 $X2=0
+ $Y2=0
cc_902 N_SET_B_c_1177_n N_A_2186_367#_c_1529_n 0.00182071f $X=11.615 $Y=1.295
+ $X2=0 $Y2=0
cc_903 N_SET_B_c_1183_n N_A_2186_367#_c_1529_n 3.01197e-19 $X=11.76 $Y=1.295
+ $X2=0 $Y2=0
cc_904 N_SET_B_M1017_g N_A_2186_367#_c_1531_n 0.0203492f $X=11.59 $Y=0.58 $X2=0
+ $Y2=0
cc_905 N_SET_B_M1017_g N_A_1804_424#_M1026_g 0.00849643f $X=11.59 $Y=0.58 $X2=0
+ $Y2=0
cc_906 N_SET_B_c_1177_n N_A_1804_424#_c_1641_n 0.0226921f $X=11.615 $Y=1.295
+ $X2=0 $Y2=0
cc_907 N_SET_B_c_1177_n N_A_1804_424#_c_1642_n 0.0215392f $X=11.615 $Y=1.295
+ $X2=0 $Y2=0
cc_908 N_SET_B_c_1182_n N_A_1804_424#_c_1642_n 3.78518e-19 $X=11.61 $Y=1.635
+ $X2=0 $Y2=0
cc_909 N_SET_B_c_1183_n N_A_1804_424#_c_1642_n 0.00736758f $X=11.76 $Y=1.295
+ $X2=0 $Y2=0
cc_910 N_SET_B_c_1182_n N_A_1804_424#_c_1644_n 0.00185705f $X=11.61 $Y=1.635
+ $X2=0 $Y2=0
cc_911 N_SET_B_c_1183_n N_A_1804_424#_c_1644_n 0.00867537f $X=11.76 $Y=1.295
+ $X2=0 $Y2=0
cc_912 N_SET_B_c_1187_n N_A_1804_424#_c_1660_n 0.00924537f $X=11.47 $Y=2.465
+ $X2=0 $Y2=0
cc_913 SET_B N_A_1804_424#_c_1661_n 0.00102137f $X=11.675 $Y=1.21 $X2=0 $Y2=0
cc_914 N_SET_B_c_1186_n N_A_1804_424#_c_1645_n 8.79832e-19 $X=11.47 $Y=2.375
+ $X2=0 $Y2=0
cc_915 N_SET_B_M1017_g N_A_1804_424#_c_1645_n 5.52256e-19 $X=11.59 $Y=0.58 $X2=0
+ $Y2=0
cc_916 SET_B N_A_1804_424#_c_1645_n 0.00702776f $X=11.675 $Y=1.21 $X2=0 $Y2=0
cc_917 N_SET_B_c_1182_n N_A_1804_424#_c_1645_n 3.63569e-19 $X=11.61 $Y=1.635
+ $X2=0 $Y2=0
cc_918 N_SET_B_c_1183_n N_A_1804_424#_c_1645_n 0.0327284f $X=11.76 $Y=1.295
+ $X2=0 $Y2=0
cc_919 N_SET_B_M1017_g N_A_1804_424#_c_1646_n 0.00770693f $X=11.59 $Y=0.58 $X2=0
+ $Y2=0
cc_920 SET_B N_A_1804_424#_c_1646_n 0.00460346f $X=11.675 $Y=1.21 $X2=0 $Y2=0
cc_921 N_SET_B_c_1182_n N_A_1804_424#_c_1646_n 0.0104335f $X=11.61 $Y=1.635
+ $X2=0 $Y2=0
cc_922 N_SET_B_c_1183_n N_A_1804_424#_c_1646_n 0.00510479f $X=11.76 $Y=1.295
+ $X2=0 $Y2=0
cc_923 N_SET_B_c_1177_n N_A_1804_424#_c_1709_n 0.00645725f $X=11.615 $Y=1.295
+ $X2=0 $Y2=0
cc_924 N_SET_B_c_1186_n N_A_1804_424#_c_1664_n 0.0226535f $X=11.47 $Y=2.375
+ $X2=0 $Y2=0
cc_925 N_SET_B_c_1187_n N_A_1804_424#_c_1664_n 0.00883221f $X=11.47 $Y=2.465
+ $X2=0 $Y2=0
cc_926 N_SET_B_c_1177_n N_A_1804_424#_c_1664_n 0.0130421f $X=11.615 $Y=1.295
+ $X2=0 $Y2=0
cc_927 SET_B N_A_1804_424#_c_1664_n 9.86625e-19 $X=11.675 $Y=1.21 $X2=0 $Y2=0
cc_928 N_SET_B_c_1182_n N_A_1804_424#_c_1664_n 0.00163909f $X=11.61 $Y=1.635
+ $X2=0 $Y2=0
cc_929 N_SET_B_c_1183_n N_A_1804_424#_c_1664_n 0.0357022f $X=11.76 $Y=1.295
+ $X2=0 $Y2=0
cc_930 N_SET_B_c_1186_n N_A_1804_424#_c_1648_n 0.00647956f $X=11.47 $Y=2.375
+ $X2=0 $Y2=0
cc_931 N_SET_B_c_1174_n N_VPWR_c_1926_n 5.45161e-19 $X=7.21 $Y=2.15 $X2=0 $Y2=0
cc_932 N_SET_B_c_1185_n N_VPWR_c_1926_n 0.00190052f $X=7.21 $Y=2.24 $X2=0 $Y2=0
cc_933 N_SET_B_c_1187_n N_VPWR_c_1928_n 0.0040383f $X=11.47 $Y=2.465 $X2=0 $Y2=0
cc_934 N_SET_B_c_1187_n N_VPWR_c_1942_n 0.00445602f $X=11.47 $Y=2.465 $X2=0
+ $Y2=0
cc_935 N_SET_B_c_1187_n N_VPWR_c_1920_n 0.00462637f $X=11.47 $Y=2.465 $X2=0
+ $Y2=0
cc_936 N_SET_B_M1021_g N_VGND_c_2321_n 0.0159047f $X=7.46 $Y=0.58 $X2=0 $Y2=0
cc_937 N_SET_B_c_1177_n N_VGND_c_2321_n 0.00139039f $X=11.615 $Y=1.295 $X2=0
+ $Y2=0
cc_938 N_SET_B_M1021_g N_VGND_c_2330_n 0.00383152f $X=7.46 $Y=0.58 $X2=0 $Y2=0
cc_939 N_SET_B_M1017_g N_VGND_c_2339_n 0.00383152f $X=11.59 $Y=0.58 $X2=0 $Y2=0
cc_940 N_SET_B_M1017_g N_VGND_c_2340_n 0.0114386f $X=11.59 $Y=0.58 $X2=0 $Y2=0
cc_941 N_SET_B_M1021_g N_VGND_c_2342_n 0.0075725f $X=7.46 $Y=0.58 $X2=0 $Y2=0
cc_942 N_SET_B_M1017_g N_VGND_c_2342_n 0.00373161f $X=11.59 $Y=0.58 $X2=0 $Y2=0
cc_943 N_SET_B_M1021_g N_A_1641_74#_c_2479_n 0.00103176f $X=7.46 $Y=0.58 $X2=0
+ $Y2=0
cc_944 N_SET_B_c_1177_n N_A_1641_74#_c_2480_n 0.0321812f $X=11.615 $Y=1.295
+ $X2=0 $Y2=0
cc_945 N_SET_B_c_1177_n N_A_1641_74#_c_2481_n 0.00922066f $X=11.615 $Y=1.295
+ $X2=0 $Y2=0
cc_946 N_SET_B_c_1177_n N_A_1641_74#_c_2482_n 0.00864504f $X=11.615 $Y=1.295
+ $X2=0 $Y2=0
cc_947 N_A_608_74#_M1043_g N_A_2186_367#_c_1524_n 0.0191919f $X=10.63 $Y=0.58
+ $X2=0 $Y2=0
cc_948 N_A_608_74#_M1043_g N_A_2186_367#_c_1528_n 0.00152879f $X=10.63 $Y=0.58
+ $X2=0 $Y2=0
cc_949 N_A_608_74#_M1043_g N_A_2186_367#_c_1531_n 0.0512761f $X=10.63 $Y=0.58
+ $X2=0 $Y2=0
cc_950 N_A_608_74#_c_1337_n N_A_1804_424#_c_1655_n 4.46185e-19 $X=9.35 $Y=3.15
+ $X2=0 $Y2=0
cc_951 N_A_608_74#_M1005_g N_A_1804_424#_c_1655_n 0.0123295f $X=9.44 $Y=2.54
+ $X2=0 $Y2=0
cc_952 N_A_608_74#_c_1341_n N_A_1804_424#_c_1655_n 0.0101531f $X=9.8 $Y=3.15
+ $X2=0 $Y2=0
cc_953 N_A_608_74#_c_1342_n N_A_1804_424#_c_1655_n 0.0118764f $X=9.89 $Y=3.035
+ $X2=0 $Y2=0
cc_954 N_A_608_74#_c_1346_n N_A_1804_424#_c_1655_n 0.00398289f $X=9.44 $Y=3.13
+ $X2=0 $Y2=0
cc_955 N_A_608_74#_c_1337_n N_A_1804_424#_c_1656_n 0.00815885f $X=9.35 $Y=3.15
+ $X2=0 $Y2=0
cc_956 N_A_608_74#_M1043_g N_A_1804_424#_c_1640_n 0.00520174f $X=10.63 $Y=0.58
+ $X2=0 $Y2=0
cc_957 N_A_608_74#_c_1342_n N_A_1804_424#_c_1657_n 0.00746493f $X=9.89 $Y=3.035
+ $X2=0 $Y2=0
cc_958 N_A_608_74#_M1043_g N_A_1804_424#_c_1725_n 0.00385881f $X=10.63 $Y=0.58
+ $X2=0 $Y2=0
cc_959 N_A_608_74#_M1043_g N_A_1804_424#_c_1641_n 0.0160324f $X=10.63 $Y=0.58
+ $X2=0 $Y2=0
cc_960 N_A_608_74#_c_1342_n N_A_1804_424#_c_1658_n 0.00196063f $X=9.89 $Y=3.035
+ $X2=0 $Y2=0
cc_961 N_A_608_74#_c_1324_n N_A_1804_424#_c_1642_n 0.00361615f $X=10.555 $Y=1.52
+ $X2=0 $Y2=0
cc_962 N_A_608_74#_M1043_g N_A_1804_424#_c_1642_n 0.00274039f $X=10.63 $Y=0.58
+ $X2=0 $Y2=0
cc_963 N_A_608_74#_c_1324_n N_A_1804_424#_c_1643_n 0.00972698f $X=10.555 $Y=1.52
+ $X2=0 $Y2=0
cc_964 N_A_608_74#_M1043_g N_A_1804_424#_c_1643_n 8.62813e-19 $X=10.63 $Y=0.58
+ $X2=0 $Y2=0
cc_965 N_A_608_74#_c_1324_n N_A_1804_424#_c_1644_n 5.16083e-19 $X=10.555 $Y=1.52
+ $X2=0 $Y2=0
cc_966 N_A_608_74#_c_1324_n N_A_1804_424#_c_1709_n 0.00374823f $X=10.555 $Y=1.52
+ $X2=0 $Y2=0
cc_967 N_A_608_74#_M1043_g N_A_1804_424#_c_1709_n 0.00327545f $X=10.63 $Y=0.58
+ $X2=0 $Y2=0
cc_968 N_A_608_74#_c_1348_n N_VPWR_M1008_d 0.00200574f $X=3.885 $Y=1.945 $X2=0
+ $Y2=0
cc_969 N_A_608_74#_c_1331_n N_VPWR_c_1924_n 0.0075987f $X=3.935 $Y=1.765 $X2=0
+ $Y2=0
cc_970 N_A_608_74#_c_1333_n N_VPWR_c_1924_n 3.39122e-19 $X=4.455 $Y=3.075 $X2=0
+ $Y2=0
cc_971 N_A_608_74#_c_1335_n N_VPWR_c_1924_n 0.00232909f $X=4.53 $Y=3.15 $X2=0
+ $Y2=0
cc_972 N_A_608_74#_c_1336_n N_VPWR_c_1925_n 6.16834e-19 $X=5.51 $Y=2.91 $X2=0
+ $Y2=0
cc_973 N_A_608_74#_c_1337_n N_VPWR_c_1925_n 0.0213655f $X=9.35 $Y=3.15 $X2=0
+ $Y2=0
cc_974 N_A_608_74#_c_1345_n N_VPWR_c_1925_n 0.00103172f $X=5.51 $Y=3.15 $X2=0
+ $Y2=0
cc_975 N_A_608_74#_c_1337_n N_VPWR_c_1926_n 0.0170937f $X=9.35 $Y=3.15 $X2=0
+ $Y2=0
cc_976 N_A_608_74#_c_1337_n N_VPWR_c_1927_n 0.0215219f $X=9.35 $Y=3.15 $X2=0
+ $Y2=0
cc_977 N_A_608_74#_M1005_g N_VPWR_c_1927_n 0.00131409f $X=9.44 $Y=2.54 $X2=0
+ $Y2=0
cc_978 N_A_608_74#_c_1331_n N_VPWR_c_1933_n 0.00413917f $X=3.935 $Y=1.765 $X2=0
+ $Y2=0
cc_979 N_A_608_74#_c_1335_n N_VPWR_c_1933_n 0.0413451f $X=4.53 $Y=3.15 $X2=0
+ $Y2=0
cc_980 N_A_608_74#_c_1337_n N_VPWR_c_1935_n 0.0290731f $X=9.35 $Y=3.15 $X2=0
+ $Y2=0
cc_981 N_A_608_74#_c_1337_n N_VPWR_c_1937_n 0.0220248f $X=9.35 $Y=3.15 $X2=0
+ $Y2=0
cc_982 N_A_608_74#_c_1337_n N_VPWR_c_1941_n 0.0319222f $X=9.35 $Y=3.15 $X2=0
+ $Y2=0
cc_983 N_A_608_74#_c_1331_n N_VPWR_c_1920_n 0.0081836f $X=3.935 $Y=1.765 $X2=0
+ $Y2=0
cc_984 N_A_608_74#_c_1334_n N_VPWR_c_1920_n 0.0207008f $X=5.42 $Y=3.15 $X2=0
+ $Y2=0
cc_985 N_A_608_74#_c_1335_n N_VPWR_c_1920_n 0.0060023f $X=4.53 $Y=3.15 $X2=0
+ $Y2=0
cc_986 N_A_608_74#_c_1337_n N_VPWR_c_1920_n 0.106627f $X=9.35 $Y=3.15 $X2=0
+ $Y2=0
cc_987 N_A_608_74#_c_1341_n N_VPWR_c_1920_n 0.0129609f $X=9.8 $Y=3.15 $X2=0
+ $Y2=0
cc_988 N_A_608_74#_c_1345_n N_VPWR_c_1920_n 0.00441434f $X=5.51 $Y=3.15 $X2=0
+ $Y2=0
cc_989 N_A_608_74#_c_1346_n N_VPWR_c_1920_n 0.00440873f $X=9.44 $Y=3.13 $X2=0
+ $Y2=0
cc_990 N_A_608_74#_c_1330_n N_A_290_464#_c_2108_n 0.00556071f $X=3.155 $Y=1.01
+ $X2=0 $Y2=0
cc_991 N_A_608_74#_c_1328_n N_A_290_464#_c_2110_n 0.00168773f $X=3.045 $Y=1.82
+ $X2=0 $Y2=0
cc_992 N_A_608_74#_M1008_s N_A_290_464#_c_2115_n 0.0120356f $X=3.125 $Y=1.84
+ $X2=0 $Y2=0
cc_993 N_A_608_74#_c_1331_n N_A_290_464#_c_2115_n 0.0151245f $X=3.935 $Y=1.765
+ $X2=0 $Y2=0
cc_994 N_A_608_74#_c_1319_n N_A_290_464#_c_2115_n 0.00417303f $X=4.425 $Y=1.68
+ $X2=0 $Y2=0
cc_995 N_A_608_74#_c_1333_n N_A_290_464#_c_2115_n 0.0127413f $X=4.455 $Y=3.075
+ $X2=0 $Y2=0
cc_996 N_A_608_74#_c_1344_n N_A_290_464#_c_2115_n 0.0013146f $X=4.44 $Y=2.12
+ $X2=0 $Y2=0
cc_997 N_A_608_74#_c_1348_n N_A_290_464#_c_2115_n 0.0643262f $X=3.885 $Y=1.945
+ $X2=0 $Y2=0
cc_998 N_A_608_74#_c_1349_n N_A_290_464#_c_2115_n 8.29095e-19 $X=3.13 $Y=1.945
+ $X2=0 $Y2=0
cc_999 N_A_608_74#_c_1344_n N_A_290_464#_c_2116_n 0.00238263f $X=4.44 $Y=2.12
+ $X2=0 $Y2=0
cc_1000 N_A_608_74#_c_1349_n N_A_290_464#_c_2117_n 0.0143305f $X=3.13 $Y=1.945
+ $X2=0 $Y2=0
cc_1001 N_A_608_74#_c_1320_n N_A_290_464#_c_2111_n 0.00627096f $X=4.805 $Y=1.115
+ $X2=0 $Y2=0
cc_1002 N_A_608_74#_c_1321_n N_A_290_464#_c_2111_n 7.52657e-19 $X=4.5 $Y=1.115
+ $X2=0 $Y2=0
cc_1003 N_A_608_74#_M1016_g N_A_290_464#_c_2111_n 0.00370144f $X=4.88 $Y=0.615
+ $X2=0 $Y2=0
cc_1004 N_A_608_74#_M1001_g N_A_290_464#_c_2112_n 0.00116188f $X=3.9 $Y=0.74
+ $X2=0 $Y2=0
cc_1005 N_A_608_74#_c_1331_n N_A_290_464#_c_2112_n 2.64877e-19 $X=3.935 $Y=1.765
+ $X2=0 $Y2=0
cc_1006 N_A_608_74#_c_1318_n N_A_290_464#_c_2112_n 0.00609576f $X=4.425 $Y=1.35
+ $X2=0 $Y2=0
cc_1007 N_A_608_74#_c_1319_n N_A_290_464#_c_2112_n 0.00943493f $X=4.425 $Y=1.68
+ $X2=0 $Y2=0
cc_1008 N_A_608_74#_c_1320_n N_A_290_464#_c_2112_n 0.00700565f $X=4.805 $Y=1.115
+ $X2=0 $Y2=0
cc_1009 N_A_608_74#_c_1321_n N_A_290_464#_c_2112_n 0.00416877f $X=4.5 $Y=1.115
+ $X2=0 $Y2=0
cc_1010 N_A_608_74#_M1016_g N_A_290_464#_c_2112_n 0.0036657f $X=4.88 $Y=0.615
+ $X2=0 $Y2=0
cc_1011 N_A_608_74#_c_1343_n N_A_290_464#_c_2112_n 0.00476159f $X=4.44 $Y=1.97
+ $X2=0 $Y2=0
cc_1012 N_A_608_74#_c_1348_n N_A_290_464#_c_2112_n 0.0179403f $X=3.885 $Y=1.945
+ $X2=0 $Y2=0
cc_1013 N_A_608_74#_c_1329_n N_A_290_464#_c_2112_n 0.0294141f $X=4.05 $Y=1.515
+ $X2=0 $Y2=0
cc_1014 N_A_608_74#_c_1343_n N_A_290_464#_c_2119_n 0.00204773f $X=4.44 $Y=1.97
+ $X2=0 $Y2=0
cc_1015 N_A_608_74#_c_1344_n N_A_290_464#_c_2119_n 0.00520887f $X=4.44 $Y=2.12
+ $X2=0 $Y2=0
cc_1016 N_A_608_74#_c_1333_n N_A_290_464#_c_2120_n 0.00910107f $X=4.455 $Y=3.075
+ $X2=0 $Y2=0
cc_1017 N_A_608_74#_c_1339_n N_A_1584_379#_c_2241_n 0.00680138f $X=9.44 $Y=2.045
+ $X2=0 $Y2=0
cc_1018 N_A_608_74#_M1005_g N_A_1584_379#_c_2241_n 0.0105053f $X=9.44 $Y=2.54
+ $X2=0 $Y2=0
cc_1019 N_A_608_74#_c_1324_n N_A_1584_379#_c_2241_n 0.00145196f $X=10.555
+ $Y=1.52 $X2=0 $Y2=0
cc_1020 N_A_608_74#_c_1342_n N_A_1584_379#_c_2241_n 0.00355999f $X=9.89 $Y=3.035
+ $X2=0 $Y2=0
cc_1021 N_A_608_74#_M1005_g N_A_1584_379#_c_2258_n 0.0115574f $X=9.44 $Y=2.54
+ $X2=0 $Y2=0
cc_1022 N_A_608_74#_c_1342_n N_A_1584_379#_c_2258_n 0.0124025f $X=9.89 $Y=3.035
+ $X2=0 $Y2=0
cc_1023 N_A_608_74#_c_1337_n N_A_1584_379#_c_2242_n 0.00615665f $X=9.35 $Y=3.15
+ $X2=0 $Y2=0
cc_1024 N_A_608_74#_M1005_g N_A_1584_379#_c_2243_n 0.00218712f $X=9.44 $Y=2.54
+ $X2=0 $Y2=0
cc_1025 N_A_608_74#_c_1327_n N_VGND_c_2318_n 0.0328901f $X=3.185 $Y=0.515 $X2=0
+ $Y2=0
cc_1026 N_A_608_74#_c_1327_n N_VGND_c_2319_n 0.0172202f $X=3.185 $Y=0.515 $X2=0
+ $Y2=0
cc_1027 N_A_608_74#_M1001_g N_VGND_c_2320_n 0.0120099f $X=3.9 $Y=0.74 $X2=0
+ $Y2=0
cc_1028 N_A_608_74#_c_1327_n N_VGND_c_2320_n 0.026158f $X=3.185 $Y=0.515 $X2=0
+ $Y2=0
cc_1029 N_A_608_74#_M1001_g N_VGND_c_2327_n 0.00383152f $X=3.9 $Y=0.74 $X2=0
+ $Y2=0
cc_1030 N_A_608_74#_M1016_g N_VGND_c_2327_n 9.15902e-19 $X=4.88 $Y=0.615 $X2=0
+ $Y2=0
cc_1031 N_A_608_74#_M1043_g N_VGND_c_2339_n 0.00430908f $X=10.63 $Y=0.58 $X2=0
+ $Y2=0
cc_1032 N_A_608_74#_M1001_g N_VGND_c_2342_n 0.00762539f $X=3.9 $Y=0.74 $X2=0
+ $Y2=0
cc_1033 N_A_608_74#_M1043_g N_VGND_c_2342_n 0.0081709f $X=10.63 $Y=0.58 $X2=0
+ $Y2=0
cc_1034 N_A_608_74#_c_1327_n N_VGND_c_2342_n 0.0142062f $X=3.185 $Y=0.515 $X2=0
+ $Y2=0
cc_1035 N_A_608_74#_c_1324_n N_A_1641_74#_c_2480_n 2.97622e-19 $X=10.555 $Y=1.52
+ $X2=0 $Y2=0
cc_1036 N_A_608_74#_c_1324_n N_A_1641_74#_c_2482_n 0.00134678f $X=10.555 $Y=1.52
+ $X2=0 $Y2=0
cc_1037 N_A_608_74#_M1043_g N_A_1641_74#_c_2482_n 2.88927e-19 $X=10.63 $Y=0.58
+ $X2=0 $Y2=0
cc_1038 N_A_2186_367#_c_1525_n N_A_1804_424#_M1026_g 0.012172f $X=12.5 $Y=0.875
+ $X2=0 $Y2=0
cc_1039 N_A_2186_367#_c_1526_n N_A_1804_424#_M1026_g 0.0010854f $X=12.64 $Y=0.58
+ $X2=0 $Y2=0
cc_1040 N_A_2186_367#_c_1527_n N_A_1804_424#_M1026_g 0.00600966f $X=12.72
+ $Y=2.31 $X2=0 $Y2=0
cc_1041 N_A_2186_367#_c_1530_n N_A_1804_424#_M1026_g 0.00339418f $X=12.652
+ $Y=0.875 $X2=0 $Y2=0
cc_1042 N_A_2186_367#_c_1537_n N_A_1804_424#_c_1649_n 0.00819862f $X=12.635
+ $Y=2.395 $X2=0 $Y2=0
cc_1043 N_A_2186_367#_c_1536_n N_A_1804_424#_c_1650_n 0.0068126f $X=12.225
+ $Y=2.75 $X2=0 $Y2=0
cc_1044 N_A_2186_367#_c_1537_n N_A_1804_424#_c_1650_n 0.00958888f $X=12.635
+ $Y=2.395 $X2=0 $Y2=0
cc_1045 N_A_2186_367#_c_1527_n N_A_1804_424#_c_1636_n 0.0228379f $X=12.72
+ $Y=2.31 $X2=0 $Y2=0
cc_1046 N_A_2186_367#_c_1530_n N_A_1804_424#_c_1636_n 0.00532238f $X=12.652
+ $Y=0.875 $X2=0 $Y2=0
cc_1047 N_A_2186_367#_c_1526_n N_A_1804_424#_c_1637_n 0.00334701f $X=12.64
+ $Y=0.58 $X2=0 $Y2=0
cc_1048 N_A_2186_367#_c_1527_n N_A_1804_424#_c_1637_n 5.25537e-19 $X=12.72
+ $Y=2.31 $X2=0 $Y2=0
cc_1049 N_A_2186_367#_c_1527_n N_A_1804_424#_c_1638_n 0.00132546f $X=12.72
+ $Y=2.31 $X2=0 $Y2=0
cc_1050 N_A_2186_367#_c_1527_n N_A_1804_424#_c_1652_n 7.74051e-19 $X=12.72
+ $Y=2.31 $X2=0 $Y2=0
cc_1051 N_A_2186_367#_c_1537_n N_A_1804_424#_c_1653_n 3.45584e-19 $X=12.635
+ $Y=2.395 $X2=0 $Y2=0
cc_1052 N_A_2186_367#_c_1538_n N_A_1804_424#_c_1653_n 0.00135996f $X=12.31
+ $Y=2.395 $X2=0 $Y2=0
cc_1053 N_A_2186_367#_c_1527_n N_A_1804_424#_c_1653_n 0.0102395f $X=12.72
+ $Y=2.31 $X2=0 $Y2=0
cc_1054 N_A_2186_367#_c_1531_n N_A_1804_424#_c_1640_n 8.3456e-19 $X=11.11 $Y=0.9
+ $X2=0 $Y2=0
cc_1055 N_A_2186_367#_c_1531_n N_A_1804_424#_c_1725_n 0.00155017f $X=11.11
+ $Y=0.9 $X2=0 $Y2=0
cc_1056 N_A_2186_367#_c_1524_n N_A_1804_424#_c_1641_n 0.00119422f $X=11.02
+ $Y=1.835 $X2=0 $Y2=0
cc_1057 N_A_2186_367#_c_1524_n N_A_1804_424#_c_1642_n 0.00658133f $X=11.02
+ $Y=1.835 $X2=0 $Y2=0
cc_1058 N_A_2186_367#_c_1528_n N_A_1804_424#_c_1642_n 0.00748906f $X=11.11
+ $Y=0.875 $X2=0 $Y2=0
cc_1059 N_A_2186_367#_c_1532_n N_A_1804_424#_c_1644_n 0.00310124f $X=11.02
+ $Y=1.925 $X2=0 $Y2=0
cc_1060 N_A_2186_367#_c_1533_n N_A_1804_424#_c_1644_n 0.00164141f $X=11.02
+ $Y=2.375 $X2=0 $Y2=0
cc_1061 N_A_2186_367#_c_1524_n N_A_1804_424#_c_1644_n 0.00880034f $X=11.02
+ $Y=1.835 $X2=0 $Y2=0
cc_1062 N_A_2186_367#_c_1534_n N_A_1804_424#_c_1660_n 8.52312e-19 $X=11.02
+ $Y=2.465 $X2=0 $Y2=0
cc_1063 N_A_2186_367#_c_1536_n N_A_1804_424#_c_1660_n 0.0363451f $X=12.225
+ $Y=2.75 $X2=0 $Y2=0
cc_1064 N_A_2186_367#_c_1538_n N_A_1804_424#_c_1660_n 3.94351e-19 $X=12.31
+ $Y=2.395 $X2=0 $Y2=0
cc_1065 N_A_2186_367#_c_1538_n N_A_1804_424#_c_1661_n 0.00628904f $X=12.31
+ $Y=2.395 $X2=0 $Y2=0
cc_1066 N_A_2186_367#_c_1537_n N_A_1804_424#_c_1662_n 0.0119564f $X=12.635
+ $Y=2.395 $X2=0 $Y2=0
cc_1067 N_A_2186_367#_c_1538_n N_A_1804_424#_c_1662_n 0.0155839f $X=12.31
+ $Y=2.395 $X2=0 $Y2=0
cc_1068 N_A_2186_367#_c_1527_n N_A_1804_424#_c_1662_n 0.0135424f $X=12.72
+ $Y=2.31 $X2=0 $Y2=0
cc_1069 N_A_2186_367#_c_1525_n N_A_1804_424#_c_1645_n 0.025786f $X=12.5 $Y=0.875
+ $X2=0 $Y2=0
cc_1070 N_A_2186_367#_c_1527_n N_A_1804_424#_c_1645_n 0.0618561f $X=12.72
+ $Y=2.31 $X2=0 $Y2=0
cc_1071 N_A_2186_367#_c_1525_n N_A_1804_424#_c_1646_n 0.00148844f $X=12.5
+ $Y=0.875 $X2=0 $Y2=0
cc_1072 N_A_2186_367#_c_1527_n N_A_1804_424#_c_1646_n 0.00182018f $X=12.72
+ $Y=2.31 $X2=0 $Y2=0
cc_1073 N_A_2186_367#_c_1530_n N_A_1804_424#_c_1646_n 4.75774e-19 $X=12.652
+ $Y=0.875 $X2=0 $Y2=0
cc_1074 N_A_2186_367#_c_1528_n N_A_1804_424#_c_1709_n 0.016946f $X=11.11
+ $Y=0.875 $X2=0 $Y2=0
cc_1075 N_A_2186_367#_c_1529_n N_A_1804_424#_c_1709_n 0.00155017f $X=11.11
+ $Y=1.065 $X2=0 $Y2=0
cc_1076 N_A_2186_367#_c_1533_n N_A_1804_424#_c_1664_n 0.0146624f $X=11.02
+ $Y=2.375 $X2=0 $Y2=0
cc_1077 N_A_2186_367#_c_1534_n N_A_1804_424#_c_1664_n 0.00786238f $X=11.02
+ $Y=2.465 $X2=0 $Y2=0
cc_1078 N_A_2186_367#_c_1538_n N_A_1804_424#_c_1664_n 0.0136908f $X=12.31
+ $Y=2.395 $X2=0 $Y2=0
cc_1079 N_A_2186_367#_c_1527_n N_A_1804_424#_c_1648_n 0.0112411f $X=12.72
+ $Y=2.31 $X2=0 $Y2=0
cc_1080 N_A_2186_367#_c_1526_n N_A_2611_98#_c_1842_n 0.0214128f $X=12.64 $Y=0.58
+ $X2=0 $Y2=0
cc_1081 N_A_2186_367#_c_1527_n N_A_2611_98#_c_1842_n 0.0221171f $X=12.72 $Y=2.31
+ $X2=0 $Y2=0
cc_1082 N_A_2186_367#_c_1530_n N_A_2611_98#_c_1842_n 0.0121616f $X=12.652
+ $Y=0.875 $X2=0 $Y2=0
cc_1083 N_A_2186_367#_c_1537_n N_A_2611_98#_c_1848_n 0.0121747f $X=12.635
+ $Y=2.395 $X2=0 $Y2=0
cc_1084 N_A_2186_367#_c_1527_n N_A_2611_98#_c_1848_n 0.0423532f $X=12.72 $Y=2.31
+ $X2=0 $Y2=0
cc_1085 N_A_2186_367#_c_1527_n N_A_2611_98#_c_1844_n 0.0207869f $X=12.72 $Y=2.31
+ $X2=0 $Y2=0
cc_1086 N_A_2186_367#_c_1534_n N_VPWR_c_1928_n 0.00986158f $X=11.02 $Y=2.465
+ $X2=0 $Y2=0
cc_1087 N_A_2186_367#_c_1536_n N_VPWR_c_1929_n 0.0221564f $X=12.225 $Y=2.75
+ $X2=0 $Y2=0
cc_1088 N_A_2186_367#_c_1537_n N_VPWR_c_1929_n 0.0224772f $X=12.635 $Y=2.395
+ $X2=0 $Y2=0
cc_1089 N_A_2186_367#_c_1534_n N_VPWR_c_1941_n 0.00413917f $X=11.02 $Y=2.465
+ $X2=0 $Y2=0
cc_1090 N_A_2186_367#_c_1536_n N_VPWR_c_1942_n 0.011054f $X=12.225 $Y=2.75 $X2=0
+ $Y2=0
cc_1091 N_A_2186_367#_c_1534_n N_VPWR_c_1920_n 0.00417401f $X=11.02 $Y=2.465
+ $X2=0 $Y2=0
cc_1092 N_A_2186_367#_c_1536_n N_VPWR_c_1920_n 0.00915483f $X=12.225 $Y=2.75
+ $X2=0 $Y2=0
cc_1093 N_A_2186_367#_c_1537_n N_VPWR_c_1920_n 0.00689018f $X=12.635 $Y=2.395
+ $X2=0 $Y2=0
cc_1094 N_A_2186_367#_c_1526_n N_VGND_c_2332_n 0.013473f $X=12.64 $Y=0.58 $X2=0
+ $Y2=0
cc_1095 N_A_2186_367#_c_1531_n N_VGND_c_2339_n 0.00461464f $X=11.11 $Y=0.9 $X2=0
+ $Y2=0
cc_1096 N_A_2186_367#_c_1525_n N_VGND_c_2340_n 0.0458287f $X=12.5 $Y=0.875 $X2=0
+ $Y2=0
cc_1097 N_A_2186_367#_c_1526_n N_VGND_c_2340_n 0.0105067f $X=12.64 $Y=0.58 $X2=0
+ $Y2=0
cc_1098 N_A_2186_367#_c_1531_n N_VGND_c_2340_n 0.00163793f $X=11.11 $Y=0.9 $X2=0
+ $Y2=0
cc_1099 N_A_2186_367#_c_1525_n N_VGND_c_2342_n 0.0198116f $X=12.5 $Y=0.875 $X2=0
+ $Y2=0
cc_1100 N_A_2186_367#_c_1526_n N_VGND_c_2342_n 0.0111726f $X=12.64 $Y=0.58 $X2=0
+ $Y2=0
cc_1101 N_A_2186_367#_c_1528_n N_VGND_c_2342_n 0.0118158f $X=11.11 $Y=0.875
+ $X2=0 $Y2=0
cc_1102 N_A_2186_367#_c_1531_n N_VGND_c_2342_n 0.00451245f $X=11.11 $Y=0.9 $X2=0
+ $Y2=0
cc_1103 N_A_2186_367#_c_1528_n A_2219_74# 0.00386116f $X=11.11 $Y=0.875
+ $X2=-0.19 $Y2=-0.245
cc_1104 N_A_1804_424#_c_1638_n N_A_2611_98#_c_1846_n 0.003789f $X=13.43 $Y=1.795
+ $X2=0 $Y2=0
cc_1105 N_A_1804_424#_c_1652_n N_A_2611_98#_c_1846_n 0.0165135f $X=13.43
+ $Y=1.885 $X2=0 $Y2=0
cc_1106 N_A_1804_424#_c_1637_n N_A_2611_98#_M1003_g 0.0118486f $X=13.415
+ $Y=1.205 $X2=0 $Y2=0
cc_1107 N_A_1804_424#_c_1639_n N_A_2611_98#_M1003_g 0.00434128f $X=13.43
+ $Y=1.365 $X2=0 $Y2=0
cc_1108 N_A_1804_424#_M1026_g N_A_2611_98#_c_1842_n 6.58111e-19 $X=12.425
+ $Y=0.58 $X2=0 $Y2=0
cc_1109 N_A_1804_424#_c_1636_n N_A_2611_98#_c_1842_n 0.0126378f $X=13.34
+ $Y=1.365 $X2=0 $Y2=0
cc_1110 N_A_1804_424#_c_1637_n N_A_2611_98#_c_1842_n 0.0105297f $X=13.415
+ $Y=1.205 $X2=0 $Y2=0
cc_1111 N_A_1804_424#_c_1639_n N_A_2611_98#_c_1842_n 0.00227239f $X=13.43
+ $Y=1.365 $X2=0 $Y2=0
cc_1112 N_A_1804_424#_c_1649_n N_A_2611_98#_c_1848_n 0.00125383f $X=12.45
+ $Y=2.375 $X2=0 $Y2=0
cc_1113 N_A_1804_424#_c_1650_n N_A_2611_98#_c_1848_n 0.00469864f $X=12.45
+ $Y=2.465 $X2=0 $Y2=0
cc_1114 N_A_1804_424#_c_1638_n N_A_2611_98#_c_1848_n 0.00575768f $X=13.43
+ $Y=1.795 $X2=0 $Y2=0
cc_1115 N_A_1804_424#_c_1652_n N_A_2611_98#_c_1848_n 0.0158843f $X=13.43
+ $Y=1.885 $X2=0 $Y2=0
cc_1116 N_A_1804_424#_c_1638_n N_A_2611_98#_c_1843_n 0.00986726f $X=13.43
+ $Y=1.795 $X2=0 $Y2=0
cc_1117 N_A_1804_424#_c_1639_n N_A_2611_98#_c_1843_n 0.0116487f $X=13.43
+ $Y=1.365 $X2=0 $Y2=0
cc_1118 N_A_1804_424#_c_1636_n N_A_2611_98#_c_1844_n 0.0146471f $X=13.34
+ $Y=1.365 $X2=0 $Y2=0
cc_1119 N_A_1804_424#_c_1638_n N_A_2611_98#_c_1844_n 0.00285552f $X=13.43
+ $Y=1.795 $X2=0 $Y2=0
cc_1120 N_A_1804_424#_c_1639_n N_A_2611_98#_c_1844_n 8.38687e-19 $X=13.43
+ $Y=1.365 $X2=0 $Y2=0
cc_1121 N_A_1804_424#_c_1638_n N_A_2611_98#_c_1845_n 0.00465427f $X=13.43
+ $Y=1.795 $X2=0 $Y2=0
cc_1122 N_A_1804_424#_c_1639_n N_A_2611_98#_c_1845_n 0.0215239f $X=13.43
+ $Y=1.365 $X2=0 $Y2=0
cc_1123 N_A_1804_424#_c_1654_n N_VPWR_c_1927_n 0.026573f $X=9.165 $Y=2.4 $X2=0
+ $Y2=0
cc_1124 N_A_1804_424#_c_1656_n N_VPWR_c_1927_n 0.00960002f $X=9.33 $Y=2.99 $X2=0
+ $Y2=0
cc_1125 N_A_1804_424#_c_1655_n N_VPWR_c_1928_n 0.00498298f $X=10.105 $Y=2.99
+ $X2=0 $Y2=0
cc_1126 N_A_1804_424#_c_1657_n N_VPWR_c_1928_n 0.0068533f $X=10.27 $Y=2.745
+ $X2=0 $Y2=0
cc_1127 N_A_1804_424#_c_1660_n N_VPWR_c_1928_n 0.0224916f $X=11.695 $Y=2.75
+ $X2=0 $Y2=0
cc_1128 N_A_1804_424#_c_1664_n N_VPWR_c_1928_n 0.0189806f $X=11.86 $Y=2.222
+ $X2=0 $Y2=0
cc_1129 N_A_1804_424#_c_1650_n N_VPWR_c_1929_n 0.0112254f $X=12.45 $Y=2.465
+ $X2=0 $Y2=0
cc_1130 N_A_1804_424#_c_1652_n N_VPWR_c_1929_n 0.00334463f $X=13.43 $Y=1.885
+ $X2=0 $Y2=0
cc_1131 N_A_1804_424#_c_1652_n N_VPWR_c_1930_n 0.0098356f $X=13.43 $Y=1.885
+ $X2=0 $Y2=0
cc_1132 N_A_1804_424#_c_1655_n N_VPWR_c_1941_n 0.0724392f $X=10.105 $Y=2.99
+ $X2=0 $Y2=0
cc_1133 N_A_1804_424#_c_1656_n N_VPWR_c_1941_n 0.0224969f $X=9.33 $Y=2.99 $X2=0
+ $Y2=0
cc_1134 N_A_1804_424#_c_1650_n N_VPWR_c_1942_n 0.00413917f $X=12.45 $Y=2.465
+ $X2=0 $Y2=0
cc_1135 N_A_1804_424#_c_1660_n N_VPWR_c_1942_n 0.0142841f $X=11.695 $Y=2.75
+ $X2=0 $Y2=0
cc_1136 N_A_1804_424#_c_1652_n N_VPWR_c_1943_n 0.00445602f $X=13.43 $Y=1.885
+ $X2=0 $Y2=0
cc_1137 N_A_1804_424#_c_1650_n N_VPWR_c_1920_n 0.00421563f $X=12.45 $Y=2.465
+ $X2=0 $Y2=0
cc_1138 N_A_1804_424#_c_1652_n N_VPWR_c_1920_n 0.00862274f $X=13.43 $Y=1.885
+ $X2=0 $Y2=0
cc_1139 N_A_1804_424#_c_1655_n N_VPWR_c_1920_n 0.0390733f $X=10.105 $Y=2.99
+ $X2=0 $Y2=0
cc_1140 N_A_1804_424#_c_1656_n N_VPWR_c_1920_n 0.0113197f $X=9.33 $Y=2.99 $X2=0
+ $Y2=0
cc_1141 N_A_1804_424#_c_1660_n N_VPWR_c_1920_n 0.0119269f $X=11.695 $Y=2.75
+ $X2=0 $Y2=0
cc_1142 N_A_1804_424#_c_1663_n N_VPWR_c_1920_n 0.0205786f $X=10.89 $Y=2.222
+ $X2=0 $Y2=0
cc_1143 N_A_1804_424#_c_1664_n N_VPWR_c_1920_n 0.00749032f $X=11.86 $Y=2.222
+ $X2=0 $Y2=0
cc_1144 N_A_1804_424#_c_1655_n N_A_1584_379#_M1005_d 0.00197722f $X=10.105
+ $Y=2.99 $X2=0 $Y2=0
cc_1145 N_A_1804_424#_M1005_s N_A_1584_379#_c_2241_n 0.00326076f $X=9.02 $Y=2.12
+ $X2=0 $Y2=0
cc_1146 N_A_1804_424#_c_1654_n N_A_1584_379#_c_2241_n 0.025036f $X=9.165 $Y=2.4
+ $X2=0 $Y2=0
cc_1147 N_A_1804_424#_c_1655_n N_A_1584_379#_c_2258_n 0.0160776f $X=10.105
+ $Y=2.99 $X2=0 $Y2=0
cc_1148 N_A_1804_424#_c_1657_n N_A_1584_379#_c_2258_n 0.0139312f $X=10.27
+ $Y=2.745 $X2=0 $Y2=0
cc_1149 N_A_1804_424#_c_1658_n N_A_1584_379#_c_2258_n 0.00970046f $X=10.435
+ $Y=2.39 $X2=0 $Y2=0
cc_1150 N_A_1804_424#_c_1647_n N_VGND_c_2322_n 0.0310131f $X=9.415 $Y=0.34 $X2=0
+ $Y2=0
cc_1151 N_A_1804_424#_c_1637_n N_VGND_c_2323_n 0.00876736f $X=13.415 $Y=1.205
+ $X2=0 $Y2=0
cc_1152 N_A_1804_424#_M1026_g N_VGND_c_2332_n 0.00461464f $X=12.425 $Y=0.58
+ $X2=0 $Y2=0
cc_1153 N_A_1804_424#_c_1637_n N_VGND_c_2332_n 0.00473385f $X=13.415 $Y=1.205
+ $X2=0 $Y2=0
cc_1154 N_A_1804_424#_c_1640_n N_VGND_c_2339_n 0.0656534f $X=10.25 $Y=0.34 $X2=0
+ $Y2=0
cc_1155 N_A_1804_424#_c_1647_n N_VGND_c_2339_n 0.0228355f $X=9.415 $Y=0.34 $X2=0
+ $Y2=0
cc_1156 N_A_1804_424#_M1026_g N_VGND_c_2340_n 0.00435671f $X=12.425 $Y=0.58
+ $X2=0 $Y2=0
cc_1157 N_A_1804_424#_M1026_g N_VGND_c_2342_n 0.0045808f $X=12.425 $Y=0.58 $X2=0
+ $Y2=0
cc_1158 N_A_1804_424#_c_1637_n N_VGND_c_2342_n 0.00508379f $X=13.415 $Y=1.205
+ $X2=0 $Y2=0
cc_1159 N_A_1804_424#_c_1640_n N_VGND_c_2342_n 0.0365041f $X=10.25 $Y=0.34 $X2=0
+ $Y2=0
cc_1160 N_A_1804_424#_c_1647_n N_VGND_c_2342_n 0.0126251f $X=9.415 $Y=0.34 $X2=0
+ $Y2=0
cc_1161 N_A_1804_424#_c_1640_n N_A_1641_74#_M1000_s 0.00168754f $X=10.25 $Y=0.34
+ $X2=0 $Y2=0
cc_1162 N_A_1804_424#_M1000_d N_A_1641_74#_c_2480_n 0.0043689f $X=9.27 $Y=0.37
+ $X2=0 $Y2=0
cc_1163 N_A_1804_424#_c_1640_n N_A_1641_74#_c_2480_n 0.0037786f $X=10.25 $Y=0.34
+ $X2=0 $Y2=0
cc_1164 N_A_1804_424#_c_1647_n N_A_1641_74#_c_2480_n 0.024138f $X=9.415 $Y=0.34
+ $X2=0 $Y2=0
cc_1165 N_A_1804_424#_c_1640_n N_A_1641_74#_c_2482_n 0.0155812f $X=10.25 $Y=0.34
+ $X2=0 $Y2=0
cc_1166 N_A_1804_424#_c_1641_n N_A_1641_74#_c_2482_n 0.0109089f $X=10.495 $Y=1.4
+ $X2=0 $Y2=0
cc_1167 N_A_2611_98#_c_1848_n N_VPWR_c_1929_n 0.0249816f $X=13.205 $Y=2.105
+ $X2=0 $Y2=0
cc_1168 N_A_2611_98#_c_1846_n N_VPWR_c_1930_n 0.00226778f $X=13.935 $Y=1.765
+ $X2=0 $Y2=0
cc_1169 N_A_2611_98#_c_1848_n N_VPWR_c_1930_n 0.0500179f $X=13.205 $Y=2.105
+ $X2=0 $Y2=0
cc_1170 N_A_2611_98#_c_1843_n N_VPWR_c_1930_n 0.0246466f $X=13.895 $Y=1.485
+ $X2=0 $Y2=0
cc_1171 N_A_2611_98#_c_1845_n N_VPWR_c_1930_n 0.00218979f $X=14.37 $Y=1.485
+ $X2=0 $Y2=0
cc_1172 N_A_2611_98#_c_1846_n N_VPWR_c_1932_n 5.20717e-19 $X=13.935 $Y=1.765
+ $X2=0 $Y2=0
cc_1173 N_A_2611_98#_c_1847_n N_VPWR_c_1932_n 0.0117458f $X=14.385 $Y=1.765
+ $X2=0 $Y2=0
cc_1174 N_A_2611_98#_c_1848_n N_VPWR_c_1943_n 0.0148169f $X=13.205 $Y=2.105
+ $X2=0 $Y2=0
cc_1175 N_A_2611_98#_c_1846_n N_VPWR_c_1944_n 0.00445602f $X=13.935 $Y=1.765
+ $X2=0 $Y2=0
cc_1176 N_A_2611_98#_c_1847_n N_VPWR_c_1944_n 0.00413917f $X=14.385 $Y=1.765
+ $X2=0 $Y2=0
cc_1177 N_A_2611_98#_c_1846_n N_VPWR_c_1920_n 0.00857473f $X=13.935 $Y=1.765
+ $X2=0 $Y2=0
cc_1178 N_A_2611_98#_c_1847_n N_VPWR_c_1920_n 0.00817726f $X=14.385 $Y=1.765
+ $X2=0 $Y2=0
cc_1179 N_A_2611_98#_c_1848_n N_VPWR_c_1920_n 0.0122313f $X=13.205 $Y=2.105
+ $X2=0 $Y2=0
cc_1180 N_A_2611_98#_M1003_g N_Q_c_2276_n 0.00758611f $X=13.94 $Y=0.76 $X2=0
+ $Y2=0
cc_1181 N_A_2611_98#_c_1841_n N_Q_c_2276_n 0.00889128f $X=14.37 $Y=1.205 $X2=0
+ $Y2=0
cc_1182 N_A_2611_98#_c_1846_n N_Q_c_2281_n 0.00879818f $X=13.935 $Y=1.765 $X2=0
+ $Y2=0
cc_1183 N_A_2611_98#_c_1847_n N_Q_c_2281_n 3.88029e-19 $X=14.385 $Y=1.765 $X2=0
+ $Y2=0
cc_1184 N_A_2611_98#_M1003_g N_Q_c_2277_n 0.00252751f $X=13.94 $Y=0.76 $X2=0
+ $Y2=0
cc_1185 N_A_2611_98#_c_1841_n N_Q_c_2277_n 0.0024145f $X=14.37 $Y=1.205 $X2=0
+ $Y2=0
cc_1186 N_A_2611_98#_c_1843_n N_Q_c_2277_n 0.00111755f $X=13.895 $Y=1.485 $X2=0
+ $Y2=0
cc_1187 N_A_2611_98#_c_1845_n N_Q_c_2277_n 0.00211234f $X=14.37 $Y=1.485 $X2=0
+ $Y2=0
cc_1188 N_A_2611_98#_M1003_g N_Q_c_2278_n 0.00352031f $X=13.94 $Y=0.76 $X2=0
+ $Y2=0
cc_1189 N_A_2611_98#_c_1841_n N_Q_c_2278_n 0.0025985f $X=14.37 $Y=1.205 $X2=0
+ $Y2=0
cc_1190 N_A_2611_98#_c_1845_n N_Q_c_2278_n 0.0056321f $X=14.37 $Y=1.485 $X2=0
+ $Y2=0
cc_1191 N_A_2611_98#_c_1843_n N_Q_c_2279_n 0.0140641f $X=13.895 $Y=1.485 $X2=0
+ $Y2=0
cc_1192 N_A_2611_98#_c_1845_n N_Q_c_2279_n 0.0196468f $X=14.37 $Y=1.485 $X2=0
+ $Y2=0
cc_1193 N_A_2611_98#_c_1846_n Q 3.21813e-19 $X=13.935 $Y=1.765 $X2=0 $Y2=0
cc_1194 N_A_2611_98#_c_1847_n Q 0.0029826f $X=14.385 $Y=1.765 $X2=0 $Y2=0
cc_1195 N_A_2611_98#_c_1843_n Q 0.00775819f $X=13.895 $Y=1.485 $X2=0 $Y2=0
cc_1196 N_A_2611_98#_c_1845_n Q 0.015043f $X=14.37 $Y=1.485 $X2=0 $Y2=0
cc_1197 N_A_2611_98#_c_1846_n Q 0.0036957f $X=13.935 $Y=1.765 $X2=0 $Y2=0
cc_1198 N_A_2611_98#_c_1847_n Q 0.0187908f $X=14.385 $Y=1.765 $X2=0 $Y2=0
cc_1199 N_A_2611_98#_c_1843_n Q 7.50447e-19 $X=13.895 $Y=1.485 $X2=0 $Y2=0
cc_1200 N_A_2611_98#_c_1845_n Q 0.00913763f $X=14.37 $Y=1.485 $X2=0 $Y2=0
cc_1201 N_A_2611_98#_M1003_g N_VGND_c_2323_n 0.00737663f $X=13.94 $Y=0.76 $X2=0
+ $Y2=0
cc_1202 N_A_2611_98#_c_1842_n N_VGND_c_2323_n 0.0474865f $X=13.2 $Y=0.635 $X2=0
+ $Y2=0
cc_1203 N_A_2611_98#_c_1843_n N_VGND_c_2323_n 0.021633f $X=13.895 $Y=1.485 $X2=0
+ $Y2=0
cc_1204 N_A_2611_98#_c_1845_n N_VGND_c_2323_n 0.00172388f $X=14.37 $Y=1.485
+ $X2=0 $Y2=0
cc_1205 N_A_2611_98#_c_1841_n N_VGND_c_2325_n 0.00876453f $X=14.37 $Y=1.205
+ $X2=0 $Y2=0
cc_1206 N_A_2611_98#_c_1842_n N_VGND_c_2332_n 0.00977247f $X=13.2 $Y=0.635 $X2=0
+ $Y2=0
cc_1207 N_A_2611_98#_M1003_g N_VGND_c_2333_n 0.00537471f $X=13.94 $Y=0.76 $X2=0
+ $Y2=0
cc_1208 N_A_2611_98#_c_1841_n N_VGND_c_2333_n 0.0051044f $X=14.37 $Y=1.205 $X2=0
+ $Y2=0
cc_1209 N_A_2611_98#_M1003_g N_VGND_c_2342_n 0.00539454f $X=13.94 $Y=0.76 $X2=0
+ $Y2=0
cc_1210 N_A_2611_98#_c_1841_n N_VGND_c_2342_n 0.00539454f $X=14.37 $Y=1.205
+ $X2=0 $Y2=0
cc_1211 N_A_2611_98#_c_1842_n N_VGND_c_2342_n 0.0111804f $X=13.2 $Y=0.635 $X2=0
+ $Y2=0
cc_1212 N_VPWR_c_1921_n N_A_290_464#_c_2121_n 0.00764771f $X=0.73 $Y=2.78 $X2=0
+ $Y2=0
cc_1213 N_VPWR_c_1940_n N_A_290_464#_c_2121_n 0.021965f $X=2.56 $Y=3.33 $X2=0
+ $Y2=0
cc_1214 N_VPWR_c_1920_n N_A_290_464#_c_2121_n 0.025762f $X=14.64 $Y=3.33 $X2=0
+ $Y2=0
cc_1215 N_VPWR_M1041_d N_A_290_464#_c_2114_n 0.00893529f $X=2.5 $Y=2.32 $X2=0
+ $Y2=0
cc_1216 N_VPWR_c_1922_n N_A_290_464#_c_2114_n 0.0253725f $X=2.725 $Y=2.995 $X2=0
+ $Y2=0
cc_1217 N_VPWR_c_1923_n N_A_290_464#_c_2114_n 0.00100823f $X=3.545 $Y=3.33 $X2=0
+ $Y2=0
cc_1218 N_VPWR_c_1940_n N_A_290_464#_c_2114_n 0.00228238f $X=2.56 $Y=3.33 $X2=0
+ $Y2=0
cc_1219 N_VPWR_c_1920_n N_A_290_464#_c_2114_n 0.0074193f $X=14.64 $Y=3.33 $X2=0
+ $Y2=0
cc_1220 N_VPWR_M1008_d N_A_290_464#_c_2115_n 0.00395925f $X=3.56 $Y=1.84 $X2=0
+ $Y2=0
cc_1221 N_VPWR_c_1924_n N_A_290_464#_c_2115_n 0.0172656f $X=3.71 $Y=2.78 $X2=0
+ $Y2=0
cc_1222 N_VPWR_c_1922_n N_A_290_464#_c_2142_n 0.00578856f $X=2.725 $Y=2.995
+ $X2=0 $Y2=0
cc_1223 N_VPWR_c_1940_n N_A_290_464#_c_2142_n 0.00471211f $X=2.56 $Y=3.33 $X2=0
+ $Y2=0
cc_1224 N_VPWR_c_1920_n N_A_290_464#_c_2142_n 0.00576777f $X=14.64 $Y=3.33 $X2=0
+ $Y2=0
cc_1225 N_VPWR_c_1923_n N_A_290_464#_c_2117_n 0.00305321f $X=3.545 $Y=3.33 $X2=0
+ $Y2=0
cc_1226 N_VPWR_c_1924_n N_A_290_464#_c_2117_n 0.00302728f $X=3.71 $Y=2.78 $X2=0
+ $Y2=0
cc_1227 N_VPWR_c_1920_n N_A_290_464#_c_2117_n 0.00485809f $X=14.64 $Y=3.33 $X2=0
+ $Y2=0
cc_1228 N_VPWR_M1009_s N_A_1584_379#_c_2244_n 0.00511543f $X=8.37 $Y=1.895 $X2=0
+ $Y2=0
cc_1229 N_VPWR_c_1927_n N_A_1584_379#_c_2244_n 0.012936f $X=8.52 $Y=2.58 $X2=0
+ $Y2=0
cc_1230 N_VPWR_c_1926_n N_A_1584_379#_c_2242_n 0.0456552f $X=7.62 $Y=2.23 $X2=0
+ $Y2=0
cc_1231 N_VPWR_c_1927_n N_A_1584_379#_c_2242_n 0.0234974f $X=8.52 $Y=2.58 $X2=0
+ $Y2=0
cc_1232 N_VPWR_c_1937_n N_A_1584_379#_c_2242_n 0.00749334f $X=8.435 $Y=3.33
+ $X2=0 $Y2=0
cc_1233 N_VPWR_c_1920_n N_A_1584_379#_c_2242_n 0.00907476f $X=14.64 $Y=3.33
+ $X2=0 $Y2=0
cc_1234 N_VPWR_M1009_s N_A_1584_379#_c_2243_n 0.00342191f $X=8.37 $Y=1.895 $X2=0
+ $Y2=0
cc_1235 N_VPWR_c_1927_n N_A_1584_379#_c_2243_n 0.00751656f $X=8.52 $Y=2.58 $X2=0
+ $Y2=0
cc_1236 N_VPWR_c_1930_n N_Q_c_2281_n 0.0311427f $X=13.705 $Y=2.085 $X2=0 $Y2=0
cc_1237 N_VPWR_c_1932_n N_Q_c_2281_n 0.0255358f $X=14.61 $Y=2.405 $X2=0 $Y2=0
cc_1238 N_VPWR_c_1944_n N_Q_c_2281_n 0.0123628f $X=14.445 $Y=3.33 $X2=0 $Y2=0
cc_1239 N_VPWR_c_1920_n N_Q_c_2281_n 0.0101999f $X=14.64 $Y=3.33 $X2=0 $Y2=0
cc_1240 N_VPWR_M1033_s Q 0.00418233f $X=14.46 $Y=1.84 $X2=0 $Y2=0
cc_1241 N_VPWR_c_1930_n Q 0.0145522f $X=13.705 $Y=2.085 $X2=0 $Y2=0
cc_1242 N_VPWR_c_1932_n Q 0.0213356f $X=14.61 $Y=2.405 $X2=0 $Y2=0
cc_1243 N_A_290_464#_c_2121_n A_416_464# 0.00472776f $X=2.215 $Y=2.785 $X2=-0.19
+ $Y2=-0.245
cc_1244 N_A_290_464#_c_2110_n A_416_464# 0.0013959f $X=2.3 $Y=2.49 $X2=-0.19
+ $Y2=-0.245
cc_1245 N_A_290_464#_c_2142_n A_416_464# 0.00356936f $X=2.3 $Y=2.575 $X2=-0.19
+ $Y2=-0.245
cc_1246 N_A_290_464#_c_2107_n N_VGND_c_2317_n 0.0107179f $X=1.725 $Y=0.58 $X2=0
+ $Y2=0
cc_1247 N_A_290_464#_c_2107_n N_VGND_c_2318_n 0.0108035f $X=1.725 $Y=0.58 $X2=0
+ $Y2=0
cc_1248 N_A_290_464#_c_2107_n N_VGND_c_2329_n 0.0144922f $X=1.725 $Y=0.58 $X2=0
+ $Y2=0
cc_1249 N_A_290_464#_c_2107_n N_VGND_c_2342_n 0.0118826f $X=1.725 $Y=0.58 $X2=0
+ $Y2=0
cc_1250 N_Q_c_2276_n N_VGND_c_2323_n 0.0558612f $X=14.155 $Y=0.535 $X2=0 $Y2=0
cc_1251 N_Q_c_2276_n N_VGND_c_2325_n 0.0596245f $X=14.155 $Y=0.535 $X2=0 $Y2=0
cc_1252 N_Q_c_2279_n N_VGND_c_2325_n 0.0217963f $X=14.465 $Y=1.49 $X2=0 $Y2=0
cc_1253 N_Q_c_2276_n N_VGND_c_2333_n 0.0143678f $X=14.155 $Y=0.535 $X2=0 $Y2=0
cc_1254 N_Q_c_2276_n N_VGND_c_2342_n 0.0128169f $X=14.155 $Y=0.535 $X2=0 $Y2=0
cc_1255 N_VGND_c_2321_n N_A_1641_74#_c_2479_n 0.0132241f $X=7.76 $Y=0.515 $X2=0
+ $Y2=0
cc_1256 N_VGND_c_2322_n N_A_1641_74#_c_2479_n 0.0138413f $X=8.855 $Y=0.53 $X2=0
+ $Y2=0
cc_1257 N_VGND_c_2331_n N_A_1641_74#_c_2479_n 0.0145302f $X=8.69 $Y=0 $X2=0
+ $Y2=0
cc_1258 N_VGND_c_2342_n N_A_1641_74#_c_2479_n 0.0118976f $X=14.64 $Y=0 $X2=0
+ $Y2=0
cc_1259 N_VGND_M1034_s N_A_1641_74#_c_2480_n 0.00454384f $X=8.635 $Y=0.37 $X2=0
+ $Y2=0
cc_1260 N_VGND_c_2322_n N_A_1641_74#_c_2480_n 0.0256711f $X=8.855 $Y=0.53 $X2=0
+ $Y2=0
