* File: sky130_fd_sc_hs__or3b_1.pex.spice
* Created: Tue Sep  1 20:20:44 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HS__OR3B_1%C_N 2 4 5 7 10 12 13 14 18 19
c34 5 0 1.5681e-19 $X=0.545 $Y=2.045
r35 18 20 46.5827 $w=3.6e-07 $l=1.65e-07 $layer=POLY_cond $X=0.455 $Y=1.275
+ $X2=0.455 $Y2=1.11
r36 18 19 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.44
+ $Y=1.275 $X2=0.44 $Y2=1.275
r37 13 14 9.21977 $w=4.78e-07 $l=3.7e-07 $layer=LI1_cond $X=0.365 $Y=1.295
+ $X2=0.365 $Y2=1.665
r38 13 19 0.498366 $w=4.78e-07 $l=2e-08 $layer=LI1_cond $X=0.365 $Y=1.295
+ $X2=0.365 $Y2=1.275
r39 10 20 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=0.56 $Y=0.645
+ $X2=0.56 $Y2=1.11
r40 5 7 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=0.545 $Y=2.045
+ $X2=0.545 $Y2=2.54
r41 4 5 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=0.545 $Y=1.955 $X2=0.545
+ $Y2=2.045
r42 4 12 68.0242 $w=1.8e-07 $l=1.75e-07 $layer=POLY_cond $X=0.545 $Y=1.955
+ $X2=0.545 $Y2=1.78
r43 2 12 43.2685 $w=3.6e-07 $l=1.8e-07 $layer=POLY_cond $X=0.455 $Y=1.6
+ $X2=0.455 $Y2=1.78
r44 1 18 2.40434 $w=3.6e-07 $l=1.5e-08 $layer=POLY_cond $X=0.455 $Y=1.29
+ $X2=0.455 $Y2=1.275
r45 1 2 49.6898 $w=3.6e-07 $l=3.1e-07 $layer=POLY_cond $X=0.455 $Y=1.29
+ $X2=0.455 $Y2=1.6
.ends

.subckt PM_SKY130_FD_SC_HS__OR3B_1%A_124_424# 1 2 7 8 9 10 13 15 17 22 26 31 34
+ 35 37 38 39 40
c62 35 0 1.5681e-19 $X=0.78 $Y=2.1
c63 13 0 1.89825e-19 $X=1.555 $Y=0.645
r64 37 39 8.78489 $w=4.28e-07 $l=1.65e-07 $layer=LI1_cond $X=0.99 $Y=1.375
+ $X2=0.99 $Y2=1.21
r65 37 38 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.04
+ $Y=1.375 $X2=1.04 $Y2=1.375
r66 35 40 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=0.86 $Y=2.1 $X2=0.86
+ $Y2=1.88
r67 34 39 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=0.86 $Y=0.94 $X2=0.86
+ $Y2=1.21
r68 31 40 10.1249 $w=4.28e-07 $l=2.15e-07 $layer=LI1_cond $X=0.99 $Y=1.665
+ $X2=0.99 $Y2=1.88
r69 30 37 1.34005 $w=4.28e-07 $l=5e-08 $layer=LI1_cond $X=0.99 $Y=1.425 $X2=0.99
+ $Y2=1.375
r70 30 31 6.43224 $w=4.28e-07 $l=2.4e-07 $layer=LI1_cond $X=0.99 $Y=1.425
+ $X2=0.99 $Y2=1.665
r71 26 35 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=0.78 $Y=2.265
+ $X2=0.78 $Y2=2.1
r72 20 34 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=0.78 $Y=0.775
+ $X2=0.78 $Y2=0.94
r73 20 22 4.53993 $w=3.28e-07 $l=1.3e-07 $layer=LI1_cond $X=0.78 $Y=0.775
+ $X2=0.78 $Y2=0.645
r74 19 38 62.0758 $w=3.3e-07 $l=3.55e-07 $layer=POLY_cond $X=1.04 $Y=1.73
+ $X2=1.04 $Y2=1.375
r75 18 38 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=1.04 $Y=1.36
+ $X2=1.04 $Y2=1.375
r76 15 17 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=1.765 $Y=1.88
+ $X2=1.765 $Y2=2.455
r77 11 13 289.713 $w=1.5e-07 $l=5.65e-07 $layer=POLY_cond $X=1.555 $Y=1.21
+ $X2=1.555 $Y2=0.645
r78 10 19 32.1775 $w=1.5e-07 $l=1.98997e-07 $layer=POLY_cond $X=1.205 $Y=1.805
+ $X2=1.04 $Y2=1.73
r79 9 15 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.69 $Y=1.805
+ $X2=1.765 $Y2=1.88
r80 9 10 248.691 $w=1.5e-07 $l=4.85e-07 $layer=POLY_cond $X=1.69 $Y=1.805
+ $X2=1.205 $Y2=1.805
r81 8 18 32.1775 $w=1.5e-07 $l=1.98997e-07 $layer=POLY_cond $X=1.205 $Y=1.285
+ $X2=1.04 $Y2=1.36
r82 7 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.48 $Y=1.285
+ $X2=1.555 $Y2=1.21
r83 7 8 141.011 $w=1.5e-07 $l=2.75e-07 $layer=POLY_cond $X=1.48 $Y=1.285
+ $X2=1.205 $Y2=1.285
r84 2 26 300 $w=1.7e-07 $l=2.20907e-07 $layer=licon1_PDIFF $count=2 $X=0.62
+ $Y=2.12 $X2=0.78 $Y2=2.265
r85 1 22 182 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_NDIFF $count=1 $X=0.635
+ $Y=0.37 $X2=0.78 $Y2=0.645
.ends

.subckt PM_SKY130_FD_SC_HS__OR3B_1%B 3 5 6 7 9 10 11 12 13 20
c45 20 0 1.89825e-19 $X=2.08 $Y=1.355
c46 6 0 1.14684e-19 $X=2.185 $Y=1.79
r47 19 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.08
+ $Y=1.355 $X2=2.08 $Y2=1.355
r48 12 13 11.8446 $w=3.58e-07 $l=3.7e-07 $layer=LI1_cond $X=2.095 $Y=2.405
+ $X2=2.095 $Y2=2.775
r49 11 12 11.8446 $w=3.58e-07 $l=3.7e-07 $layer=LI1_cond $X=2.095 $Y=2.035
+ $X2=2.095 $Y2=2.405
r50 10 11 11.8446 $w=3.58e-07 $l=3.7e-07 $layer=LI1_cond $X=2.095 $Y=1.665
+ $X2=2.095 $Y2=2.035
r51 10 20 9.92381 $w=3.58e-07 $l=3.1e-07 $layer=LI1_cond $X=2.095 $Y=1.665
+ $X2=2.095 $Y2=1.355
r52 7 9 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=2.185 $Y=1.88
+ $X2=2.185 $Y2=2.455
r53 6 7 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=2.185 $Y=1.79 $X2=2.185
+ $Y2=1.88
r54 5 19 48.8089 $w=2.97e-07 $l=2.96606e-07 $layer=POLY_cond $X=2.185 $Y=1.61
+ $X2=2.095 $Y2=1.355
r55 5 6 69.9677 $w=1.8e-07 $l=1.8e-07 $layer=POLY_cond $X=2.185 $Y=1.61
+ $X2=2.185 $Y2=1.79
r56 1 19 38.5662 $w=2.97e-07 $l=1.79374e-07 $layer=POLY_cond $X=2.125 $Y=1.19
+ $X2=2.095 $Y2=1.355
r57 1 3 279.457 $w=1.5e-07 $l=5.45e-07 $layer=POLY_cond $X=2.125 $Y=1.19
+ $X2=2.125 $Y2=0.645
.ends

.subckt PM_SKY130_FD_SC_HS__OR3B_1%A 3 6 7 9 10 13 14
r38 13 16 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.68 $Y=1.465
+ $X2=2.68 $Y2=1.63
r39 13 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.68 $Y=1.465
+ $X2=2.68 $Y2=1.3
r40 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.68
+ $Y=1.465 $X2=2.68 $Y2=1.465
r41 10 14 6.9845 $w=3.28e-07 $l=2e-07 $layer=LI1_cond $X=2.68 $Y=1.665 $X2=2.68
+ $Y2=1.465
r42 7 9 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=2.605 $Y=1.88
+ $X2=2.605 $Y2=2.455
r43 6 7 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=2.605 $Y=1.79 $X2=2.605
+ $Y2=1.88
r44 6 16 62.1936 $w=1.8e-07 $l=1.6e-07 $layer=POLY_cond $X=2.605 $Y=1.79
+ $X2=2.605 $Y2=1.63
r45 3 15 335.862 $w=1.5e-07 $l=6.55e-07 $layer=POLY_cond $X=2.59 $Y=0.645
+ $X2=2.59 $Y2=1.3
.ends

.subckt PM_SKY130_FD_SC_HS__OR3B_1%A_239_74# 1 2 3 10 12 15 19 23 27 31 33 36 37
+ 38 42
c91 37 0 1.96631e-19 $X=1.44 $Y=0.935
c92 23 0 1.14684e-19 $X=1.54 $Y=2.1
r93 42 43 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.25
+ $Y=1.465 $X2=3.25 $Y2=1.465
r94 39 42 3.84148 $w=3.28e-07 $l=1.1e-07 $layer=LI1_cond $X=3.14 $Y=1.465
+ $X2=3.25 $Y2=1.465
r95 36 39 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.14 $Y=1.3 $X2=3.14
+ $Y2=1.465
r96 35 36 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=3.14 $Y=1.02
+ $X2=3.14 $Y2=1.3
r97 34 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.505 $Y=0.935
+ $X2=2.34 $Y2=0.935
r98 33 35 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.055 $Y=0.935
+ $X2=3.14 $Y2=1.02
r99 33 34 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=3.055 $Y=0.935
+ $X2=2.505 $Y2=0.935
r100 29 38 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.34 $Y=0.85
+ $X2=2.34 $Y2=0.935
r101 29 31 7.15912 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=2.34 $Y=0.85
+ $X2=2.34 $Y2=0.645
r102 28 37 3.80956 $w=1.7e-07 $l=2.65e-07 $layer=LI1_cond $X=1.705 $Y=0.935
+ $X2=1.44 $Y2=0.935
r103 27 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.175 $Y=0.935
+ $X2=2.34 $Y2=0.935
r104 27 28 30.6631 $w=1.68e-07 $l=4.7e-07 $layer=LI1_cond $X=2.175 $Y=0.935
+ $X2=1.705 $Y2=0.935
r105 23 25 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=1.54 $Y=2.1 $X2=1.54
+ $Y2=2.81
r106 21 37 2.88756 $w=3.3e-07 $l=1.36015e-07 $layer=LI1_cond $X=1.54 $Y=1.02
+ $X2=1.44 $Y2=0.935
r107 21 23 37.7163 $w=3.28e-07 $l=1.08e-06 $layer=LI1_cond $X=1.54 $Y=1.02
+ $X2=1.54 $Y2=2.1
r108 17 37 2.88756 $w=3.3e-07 $l=1.36015e-07 $layer=LI1_cond $X=1.34 $Y=0.85
+ $X2=1.44 $Y2=0.935
r109 17 19 7.15912 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=1.34 $Y=0.85
+ $X2=1.34 $Y2=0.645
r110 13 43 38.6157 $w=2.9e-07 $l=2.06325e-07 $layer=POLY_cond $X=3.345 $Y=1.3
+ $X2=3.252 $Y2=1.465
r111 13 15 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=3.345 $Y=1.3
+ $X2=3.345 $Y2=0.74
r112 10 43 61.0536 $w=2.9e-07 $l=3.29545e-07 $layer=POLY_cond $X=3.19 $Y=1.765
+ $X2=3.252 $Y2=1.465
r113 10 12 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.19 $Y=1.765
+ $X2=3.19 $Y2=2.4
r114 3 25 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=1.395
+ $Y=1.955 $X2=1.54 $Y2=2.81
r115 3 23 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=1.395
+ $Y=1.955 $X2=1.54 $Y2=2.1
r116 2 31 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=2.2
+ $Y=0.37 $X2=2.34 $Y2=0.645
r117 1 19 182 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_NDIFF $count=1 $X=1.195
+ $Y=0.37 $X2=1.34 $Y2=0.645
.ends

.subckt PM_SKY130_FD_SC_HS__OR3B_1%VPWR 1 2 7 9 13 18 19 20 30 31
r37 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r38 30 31 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r39 28 31 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.6 $Y2=3.33
r40 27 28 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r41 25 35 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r42 24 27 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=0.72 $Y=3.33
+ $X2=2.64 $Y2=3.33
r43 24 25 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r44 22 34 4.73185 $w=1.7e-07 $l=2.23e-07 $layer=LI1_cond $X=0.445 $Y=3.33
+ $X2=0.222 $Y2=3.33
r45 22 24 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=0.445 $Y=3.33
+ $X2=0.72 $Y2=3.33
r46 20 28 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=2.64 $Y2=3.33
r47 20 25 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=0.72 $Y2=3.33
r48 18 27 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=2.75 $Y=3.33
+ $X2=2.64 $Y2=3.33
r49 18 19 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.75 $Y=3.33
+ $X2=2.915 $Y2=3.33
r50 17 30 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=3.08 $Y=3.33 $X2=3.6
+ $Y2=3.33
r51 17 19 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.08 $Y=3.33
+ $X2=2.915 $Y2=3.33
r52 13 16 24.4458 $w=3.28e-07 $l=7e-07 $layer=LI1_cond $X=2.915 $Y=2.115
+ $X2=2.915 $Y2=2.815
r53 11 19 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.915 $Y=3.245
+ $X2=2.915 $Y2=3.33
r54 11 16 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=2.915 $Y=3.245
+ $X2=2.915 $Y2=2.815
r55 7 34 3.03433 $w=3.3e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.28 $Y=3.245
+ $X2=0.222 $Y2=3.33
r56 7 9 34.2241 $w=3.28e-07 $l=9.8e-07 $layer=LI1_cond $X=0.28 $Y=3.245 $X2=0.28
+ $Y2=2.265
r57 2 16 400 $w=1.7e-07 $l=9.70412e-07 $layer=licon1_PDIFF $count=1 $X=2.68
+ $Y=1.955 $X2=2.915 $Y2=2.815
r58 2 13 400 $w=1.7e-07 $l=3.04672e-07 $layer=licon1_PDIFF $count=1 $X=2.68
+ $Y=1.955 $X2=2.915 $Y2=2.115
r59 1 9 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=2.12 $X2=0.28 $Y2=2.265
.ends

.subckt PM_SKY130_FD_SC_HS__OR3B_1%X 1 2 9 14 15 16 17 28
r24 21 28 0.800308 $w=3.58e-07 $l=2.5e-08 $layer=LI1_cond $X=3.575 $Y=0.95
+ $X2=3.575 $Y2=0.925
r25 17 30 8.03084 $w=3.58e-07 $l=1.5e-07 $layer=LI1_cond $X=3.575 $Y=0.98
+ $X2=3.575 $Y2=1.13
r26 17 21 0.960369 $w=3.58e-07 $l=3e-08 $layer=LI1_cond $X=3.575 $Y=0.98
+ $X2=3.575 $Y2=0.95
r27 17 28 0.960369 $w=3.58e-07 $l=3e-08 $layer=LI1_cond $X=3.575 $Y=0.895
+ $X2=3.575 $Y2=0.925
r28 16 17 12.1647 $w=3.58e-07 $l=3.8e-07 $layer=LI1_cond $X=3.575 $Y=0.515
+ $X2=3.575 $Y2=0.895
r29 15 30 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=3.67 $Y=1.82 $X2=3.67
+ $Y2=1.13
r30 14 15 9.54788 $w=5.03e-07 $l=1.65e-07 $layer=LI1_cond $X=3.502 $Y=1.985
+ $X2=3.502 $Y2=1.82
r31 7 14 2.06057 $w=5.03e-07 $l=8.7e-08 $layer=LI1_cond $X=3.502 $Y=2.072
+ $X2=3.502 $Y2=1.985
r32 7 9 17.5977 $w=5.03e-07 $l=7.43e-07 $layer=LI1_cond $X=3.502 $Y=2.072
+ $X2=3.502 $Y2=2.815
r33 2 14 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=3.265
+ $Y=1.84 $X2=3.415 $Y2=1.985
r34 2 9 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=3.265
+ $Y=1.84 $X2=3.415 $Y2=2.815
r35 1 16 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.42
+ $Y=0.37 $X2=3.56 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__OR3B_1%VGND 1 2 3 10 12 16 20 22 24 29 36 37 43 46
c50 2 0 1.96631e-19 $X=1.63 $Y=0.37
r51 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r52 43 44 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r53 40 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r54 37 47 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=3.12
+ $Y2=0
r55 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r56 34 46 11.9488 $w=1.7e-07 $l=2.75e-07 $layer=LI1_cond $X=3.225 $Y=0 $X2=2.95
+ $Y2=0
r57 34 36 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=3.225 $Y=0 $X2=3.6
+ $Y2=0
r58 33 47 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r59 32 33 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r60 30 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.005 $Y=0 $X2=1.84
+ $Y2=0
r61 30 32 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=2.005 $Y=0 $X2=2.64
+ $Y2=0
r62 29 46 11.9488 $w=1.7e-07 $l=2.75e-07 $layer=LI1_cond $X=2.675 $Y=0 $X2=2.95
+ $Y2=0
r63 29 32 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=2.675 $Y=0 $X2=2.64
+ $Y2=0
r64 28 44 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r65 28 41 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r66 27 28 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r67 25 40 4.73185 $w=1.7e-07 $l=2.23e-07 $layer=LI1_cond $X=0.445 $Y=0 $X2=0.222
+ $Y2=0
r68 25 27 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=0.445 $Y=0 $X2=0.72
+ $Y2=0
r69 24 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.675 $Y=0 $X2=1.84
+ $Y2=0
r70 24 27 62.3048 $w=1.68e-07 $l=9.55e-07 $layer=LI1_cond $X=1.675 $Y=0 $X2=0.72
+ $Y2=0
r71 22 33 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=2.64
+ $Y2=0
r72 22 44 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=1.68
+ $Y2=0
r73 18 46 2.31338 $w=5.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.95 $Y=0.085
+ $X2=2.95 $Y2=0
r74 18 20 9.35116 $w=5.48e-07 $l=4.3e-07 $layer=LI1_cond $X=2.95 $Y=0.085
+ $X2=2.95 $Y2=0.515
r75 14 43 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.84 $Y=0.085
+ $X2=1.84 $Y2=0
r76 14 16 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=1.84 $Y=0.085
+ $X2=1.84 $Y2=0.515
r77 10 40 3.03433 $w=3.3e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.28 $Y=0.085
+ $X2=0.222 $Y2=0
r78 10 12 19.5566 $w=3.28e-07 $l=5.6e-07 $layer=LI1_cond $X=0.28 $Y=0.085
+ $X2=0.28 $Y2=0.645
r79 3 20 182 $w=1.7e-07 $l=3.50071e-07 $layer=licon1_NDIFF $count=1 $X=2.665
+ $Y=0.37 $X2=2.95 $Y2=0.515
r80 2 16 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=1.63
+ $Y=0.37 $X2=1.84 $Y2=0.515
r81 1 12 182 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.645
.ends

