# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_hs__a41o_1
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_hs__a41o_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.320000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.261000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.025000 1.450000 2.355000 1.780000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.261000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.525000 0.440000 2.895000 1.550000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.261000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.135000 1.180000 3.715000 1.550000 ;
    END
  END A3
  PIN A4
    ANTENNAGATEAREA  0.261000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.885000 1.180000 4.215000 1.550000 ;
    END
  END A4
  PIN B1
    ANTENNAGATEAREA  0.261000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.485000 1.450000 1.815000 1.780000 ;
    END
  END B1
  PIN X
    ANTENNADIFFAREA  1.040800 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.115000 0.290000 1.120000 0.940000 ;
        RECT 0.115000 0.940000 0.355000 1.820000 ;
        RECT 0.115000 1.820000 0.445000 2.980000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 4.320000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 4.320000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.320000 0.085000 ;
      RECT 0.000000  3.245000 4.320000 3.415000 ;
      RECT 0.575000  1.110000 2.120000 1.280000 ;
      RECT 0.575000  1.280000 1.315000 1.550000 ;
      RECT 0.645000  1.820000 0.895000 3.245000 ;
      RECT 1.145000  1.550000 1.315000 1.950000 ;
      RECT 1.145000  1.950000 1.635000 2.980000 ;
      RECT 1.290000  0.085000 1.620000 0.940000 ;
      RECT 1.790000  0.350000 2.120000 1.110000 ;
      RECT 1.805000  1.950000 3.165000 2.120000 ;
      RECT 1.805000  2.120000 2.135000 2.980000 ;
      RECT 2.305000  2.290000 2.635000 3.245000 ;
      RECT 2.835000  1.720000 4.185000 1.890000 ;
      RECT 2.835000  1.890000 3.165000 1.950000 ;
      RECT 2.835000  2.120000 3.165000 2.980000 ;
      RECT 3.335000  2.060000 3.665000 3.245000 ;
      RECT 3.830000  0.085000 4.160000 1.010000 ;
      RECT 3.855000  1.890000 4.185000 2.980000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
  END
END sky130_fd_sc_hs__a41o_1
END LIBRARY
