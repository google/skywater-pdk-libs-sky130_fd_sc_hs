* File: sky130_fd_sc_hs__bufinv_16.pxi.spice
* Created: Tue Sep  1 19:57:18 2020
* 
x_PM_SKY130_FD_SC_HS__BUFINV_16%A N_A_M1002_g N_A_c_218_n N_A_M1015_g
+ N_A_c_219_n N_A_M1017_g N_A_M1030_g N_A_c_220_n N_A_M1022_g N_A_M1043_g A A A
+ N_A_c_216_n N_A_c_217_n PM_SKY130_FD_SC_HS__BUFINV_16%A
x_PM_SKY130_FD_SC_HS__BUFINV_16%A_27_74# N_A_27_74#_M1002_d N_A_27_74#_M1030_d
+ N_A_27_74#_M1015_d N_A_27_74#_M1017_d N_A_27_74#_M1010_g N_A_27_74#_c_298_n
+ N_A_27_74#_M1000_g N_A_27_74#_M1014_g N_A_27_74#_c_299_n N_A_27_74#_M1004_g
+ N_A_27_74#_M1016_g N_A_27_74#_c_300_n N_A_27_74#_M1009_g N_A_27_74#_M1024_g
+ N_A_27_74#_c_301_n N_A_27_74#_M1026_g N_A_27_74#_M1046_g N_A_27_74#_c_302_n
+ N_A_27_74#_M1044_g N_A_27_74#_c_284_n N_A_27_74#_c_285_n N_A_27_74#_M1049_g
+ N_A_27_74#_c_287_n N_A_27_74#_c_305_n N_A_27_74#_M1047_g N_A_27_74#_c_288_n
+ N_A_27_74#_c_289_n N_A_27_74#_c_306_n N_A_27_74#_c_307_n N_A_27_74#_c_290_n
+ N_A_27_74#_c_291_n N_A_27_74#_c_323_n N_A_27_74#_c_308_n N_A_27_74#_c_292_n
+ N_A_27_74#_c_293_n N_A_27_74#_c_335_n N_A_27_74#_c_294_n N_A_27_74#_c_295_n
+ N_A_27_74#_c_338_n N_A_27_74#_c_296_n N_A_27_74#_c_297_n
+ PM_SKY130_FD_SC_HS__BUFINV_16%A_27_74#
x_PM_SKY130_FD_SC_HS__BUFINV_16%A_384_74# N_A_384_74#_M1010_d
+ N_A_384_74#_M1016_d N_A_384_74#_M1046_d N_A_384_74#_M1000_s
+ N_A_384_74#_M1009_s N_A_384_74#_M1044_s N_A_384_74#_M1003_g
+ N_A_384_74#_c_513_n N_A_384_74#_M1001_g N_A_384_74#_M1006_g
+ N_A_384_74#_c_514_n N_A_384_74#_M1005_g N_A_384_74#_M1012_g
+ N_A_384_74#_c_515_n N_A_384_74#_M1007_g N_A_384_74#_M1018_g
+ N_A_384_74#_c_516_n N_A_384_74#_M1008_g N_A_384_74#_M1020_g
+ N_A_384_74#_c_517_n N_A_384_74#_M1011_g N_A_384_74#_M1021_g
+ N_A_384_74#_c_518_n N_A_384_74#_M1013_g N_A_384_74#_c_519_n
+ N_A_384_74#_M1019_g N_A_384_74#_M1025_g N_A_384_74#_M1027_g
+ N_A_384_74#_c_520_n N_A_384_74#_M1023_g N_A_384_74#_c_521_n
+ N_A_384_74#_M1029_g N_A_384_74#_M1028_g N_A_384_74#_c_522_n
+ N_A_384_74#_M1032_g N_A_384_74#_M1031_g N_A_384_74#_c_523_n
+ N_A_384_74#_M1037_g N_A_384_74#_M1033_g N_A_384_74#_M1034_g
+ N_A_384_74#_c_524_n N_A_384_74#_M1039_g N_A_384_74#_M1035_g
+ N_A_384_74#_c_525_n N_A_384_74#_M1040_g N_A_384_74#_M1036_g
+ N_A_384_74#_c_526_n N_A_384_74#_M1041_g N_A_384_74#_c_527_n
+ N_A_384_74#_M1045_g N_A_384_74#_M1038_g N_A_384_74#_M1042_g
+ N_A_384_74#_c_528_n N_A_384_74#_M1048_g N_A_384_74#_c_529_n
+ N_A_384_74#_c_496_n N_A_384_74#_c_497_n N_A_384_74#_c_498_n
+ N_A_384_74#_c_530_n N_A_384_74#_c_531_n N_A_384_74#_c_499_n
+ N_A_384_74#_c_532_n N_A_384_74#_c_500_n N_A_384_74#_c_533_n
+ N_A_384_74#_c_501_n N_A_384_74#_c_502_n N_A_384_74#_c_535_n
+ N_A_384_74#_c_503_n N_A_384_74#_c_536_n N_A_384_74#_c_504_n
+ N_A_384_74#_c_505_n N_A_384_74#_c_506_n N_A_384_74#_c_507_n
+ N_A_384_74#_c_508_n N_A_384_74#_c_509_n N_A_384_74#_c_510_n
+ N_A_384_74#_c_511_n N_A_384_74#_c_512_n
+ PM_SKY130_FD_SC_HS__BUFINV_16%A_384_74#
x_PM_SKY130_FD_SC_HS__BUFINV_16%VPWR N_VPWR_M1015_s N_VPWR_M1022_s
+ N_VPWR_M1004_d N_VPWR_M1026_d N_VPWR_M1047_d N_VPWR_M1005_d N_VPWR_M1008_d
+ N_VPWR_M1013_d N_VPWR_M1023_d N_VPWR_M1032_d N_VPWR_M1039_d N_VPWR_M1041_d
+ N_VPWR_M1048_d N_VPWR_c_937_n N_VPWR_c_938_n N_VPWR_c_939_n N_VPWR_c_940_n
+ N_VPWR_c_941_n N_VPWR_c_942_n N_VPWR_c_943_n N_VPWR_c_944_n N_VPWR_c_945_n
+ N_VPWR_c_946_n N_VPWR_c_947_n N_VPWR_c_948_n N_VPWR_c_949_n N_VPWR_c_950_n
+ N_VPWR_c_951_n N_VPWR_c_952_n N_VPWR_c_953_n N_VPWR_c_954_n N_VPWR_c_955_n
+ N_VPWR_c_956_n N_VPWR_c_957_n N_VPWR_c_958_n N_VPWR_c_959_n N_VPWR_c_960_n
+ N_VPWR_c_961_n N_VPWR_c_962_n N_VPWR_c_963_n N_VPWR_c_964_n N_VPWR_c_965_n
+ VPWR N_VPWR_c_966_n N_VPWR_c_967_n N_VPWR_c_968_n N_VPWR_c_969_n
+ N_VPWR_c_970_n N_VPWR_c_971_n N_VPWR_c_972_n N_VPWR_c_973_n N_VPWR_c_974_n
+ N_VPWR_c_936_n PM_SKY130_FD_SC_HS__BUFINV_16%VPWR
x_PM_SKY130_FD_SC_HS__BUFINV_16%Y N_Y_M1003_s N_Y_M1012_s N_Y_M1020_s
+ N_Y_M1025_s N_Y_M1028_s N_Y_M1033_s N_Y_M1035_s N_Y_M1038_s N_Y_M1001_s
+ N_Y_M1007_s N_Y_M1011_s N_Y_M1019_s N_Y_M1029_s N_Y_M1037_s N_Y_M1040_s
+ N_Y_M1045_s N_Y_c_1159_n N_Y_c_1160_n N_Y_c_1161_n N_Y_c_1162_n N_Y_c_1171_n
+ N_Y_c_1226_n N_Y_c_1172_n N_Y_c_1163_n N_Y_c_1241_n N_Y_c_1174_n N_Y_c_1164_n
+ N_Y_c_1165_n N_Y_c_1166_n N_Y_c_1276_n N_Y_c_1280_n N_Y_c_1284_n N_Y_c_1288_n
+ N_Y_c_1178_n Y N_Y_c_1179_n N_Y_c_1180_n N_Y_c_1181_n N_Y_c_1182_n
+ N_Y_c_1183_n N_Y_c_1305_n N_Y_c_1328_n PM_SKY130_FD_SC_HS__BUFINV_16%Y
x_PM_SKY130_FD_SC_HS__BUFINV_16%VGND N_VGND_M1002_s N_VGND_M1043_s
+ N_VGND_M1014_s N_VGND_M1024_s N_VGND_M1049_s N_VGND_M1006_d N_VGND_M1018_d
+ N_VGND_M1021_d N_VGND_M1027_d N_VGND_M1031_d N_VGND_M1034_d N_VGND_M1036_d
+ N_VGND_M1042_d N_VGND_c_1421_n N_VGND_c_1422_n N_VGND_c_1423_n N_VGND_c_1424_n
+ N_VGND_c_1425_n N_VGND_c_1426_n N_VGND_c_1427_n N_VGND_c_1428_n
+ N_VGND_c_1429_n N_VGND_c_1430_n N_VGND_c_1431_n N_VGND_c_1432_n
+ N_VGND_c_1433_n N_VGND_c_1434_n N_VGND_c_1435_n N_VGND_c_1436_n
+ N_VGND_c_1437_n N_VGND_c_1438_n N_VGND_c_1439_n N_VGND_c_1440_n
+ N_VGND_c_1441_n N_VGND_c_1442_n VGND N_VGND_c_1443_n N_VGND_c_1444_n
+ N_VGND_c_1445_n N_VGND_c_1446_n N_VGND_c_1447_n N_VGND_c_1448_n
+ N_VGND_c_1449_n N_VGND_c_1450_n N_VGND_c_1451_n N_VGND_c_1452_n
+ N_VGND_c_1453_n N_VGND_c_1454_n N_VGND_c_1455_n N_VGND_c_1456_n
+ N_VGND_c_1457_n N_VGND_c_1458_n N_VGND_c_1459_n N_VGND_c_1460_n
+ PM_SKY130_FD_SC_HS__BUFINV_16%VGND
cc_1 VNB N_A_M1002_g 0.0327337f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_2 VNB N_A_M1030_g 0.0240034f $X=-0.19 $Y=-0.245 $X2=0.985 $Y2=0.74
cc_3 VNB N_A_M1043_g 0.0227235f $X=-0.19 $Y=-0.245 $X2=1.415 $Y2=0.74
cc_4 VNB N_A_c_216_n 0.0166485f $X=-0.19 $Y=-0.245 $X2=1.265 $Y2=1.515
cc_5 VNB N_A_c_217_n 0.0568731f $X=-0.19 $Y=-0.245 $X2=1.41 $Y2=1.557
cc_6 VNB N_A_27_74#_M1010_g 0.0208043f $X=-0.19 $Y=-0.245 $X2=1.41 $Y2=1.765
cc_7 VNB N_A_27_74#_M1014_g 0.0203546f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_8 VNB N_A_27_74#_M1016_g 0.0209331f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=1.557
cc_9 VNB N_A_27_74#_M1024_g 0.0211968f $X=-0.19 $Y=-0.245 $X2=1.265 $Y2=1.515
cc_10 VNB N_A_27_74#_M1046_g 0.0210803f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.565
cc_11 VNB N_A_27_74#_c_284_n 0.00890084f $X=-0.19 $Y=-0.245 $X2=1.265 $Y2=1.565
cc_12 VNB N_A_27_74#_c_285_n 0.123798f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_27_74#_M1049_g 0.0215143f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_27_74#_c_287_n 0.00937171f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_27_74#_c_288_n 0.00787792f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_27_74#_c_289_n 0.0266107f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_27_74#_c_290_n 0.00360698f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_27_74#_c_291_n 0.00998227f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_27_74#_c_292_n 0.00179995f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_27_74#_c_293_n 0.00415915f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_27_74#_c_294_n 4.30857e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_27_74#_c_295_n 6.65696e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_27_74#_c_296_n 0.00127131f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_27_74#_c_297_n 0.00563641f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_384_74#_M1003_g 0.0216367f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_384_74#_M1006_g 0.0204987f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.557
cc_27 VNB N_A_384_74#_M1012_g 0.021162f $X=-0.19 $Y=-0.245 $X2=1.265 $Y2=1.557
cc_28 VNB N_A_384_74#_M1018_g 0.021363f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_384_74#_M1020_g 0.0211843f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_384_74#_M1021_g 0.0213617f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_384_74#_M1025_g 0.0211822f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_384_74#_M1027_g 0.0213612f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_384_74#_M1028_g 0.0211812f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_384_74#_M1031_g 0.0213612f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_384_74#_M1033_g 0.0211812f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_384_74#_M1034_g 0.0213612f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_384_74#_M1035_g 0.0211812f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_384_74#_M1036_g 0.0213612f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_384_74#_M1038_g 0.021184f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_384_74#_M1042_g 0.0260277f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_384_74#_c_496_n 0.00178908f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_384_74#_c_497_n 0.00275044f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_384_74#_c_498_n 0.00140873f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_384_74#_c_499_n 0.00206666f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_A_384_74#_c_500_n 0.00374208f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_A_384_74#_c_501_n 0.00206666f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_384_74#_c_502_n 0.00686392f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_384_74#_c_503_n 0.00178779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A_384_74#_c_504_n 0.00180003f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_A_384_74#_c_505_n 0.00109754f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_A_384_74#_c_506_n 0.00177315f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_A_384_74#_c_507_n 0.00176232f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_A_384_74#_c_508_n 0.00176506f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_A_384_74#_c_509_n 0.00176778f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_A_384_74#_c_510_n 0.00176778f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_A_384_74#_c_511_n 0.00183757f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_A_384_74#_c_512_n 0.476765f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_VPWR_c_936_n 0.502022f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_Y_c_1159_n 0.00378061f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_Y_c_1160_n 0.00574953f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_Y_c_1161_n 0.00397969f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_Y_c_1162_n 0.00398355f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_Y_c_1163_n 0.00398531f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_Y_c_1164_n 0.00398531f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_Y_c_1165_n 0.00398531f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_Y_c_1166_n 0.00269539f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_VGND_c_1421_n 0.00563075f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_VGND_c_1422_n 0.00258815f $X=-0.19 $Y=-0.245 $X2=1.2 $Y2=1.565
cc_69 VNB N_VGND_c_1423_n 0.0040939f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_VGND_c_1424_n 0.00495983f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_VGND_c_1425_n 0.00754943f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_VGND_c_1426_n 0.00419598f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_VGND_c_1427_n 0.00502158f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_VGND_c_1428_n 0.00498499f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_VGND_c_1429_n 0.00494723f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_VGND_c_1430_n 0.00494723f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_VGND_c_1431_n 0.00494723f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_VGND_c_1432_n 0.00508214f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VNB N_VGND_c_1433_n 0.0122168f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_VGND_c_1434_n 0.0547214f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_81 VNB N_VGND_c_1435_n 0.0151736f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_82 VNB N_VGND_c_1436_n 0.00461913f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_83 VNB N_VGND_c_1437_n 0.0172524f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_84 VNB N_VGND_c_1438_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_85 VNB N_VGND_c_1439_n 0.0169342f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_86 VNB N_VGND_c_1440_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_87 VNB N_VGND_c_1441_n 0.0169342f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_88 VNB N_VGND_c_1442_n 0.00461913f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_89 VNB N_VGND_c_1443_n 0.0173909f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_90 VNB N_VGND_c_1444_n 0.0172409f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_91 VNB N_VGND_c_1445_n 0.0175258f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_92 VNB N_VGND_c_1446_n 0.0170514f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_93 VNB N_VGND_c_1447_n 0.0169733f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_94 VNB N_VGND_c_1448_n 0.0169342f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_95 VNB N_VGND_c_1449_n 0.0169342f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_96 VNB N_VGND_c_1450_n 0.0169342f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_97 VNB N_VGND_c_1451_n 0.0186948f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_98 VNB N_VGND_c_1452_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_99 VNB N_VGND_c_1453_n 0.00604233f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_100 VNB N_VGND_c_1454_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_101 VNB N_VGND_c_1455_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_102 VNB N_VGND_c_1456_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_103 VNB N_VGND_c_1457_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_104 VNB N_VGND_c_1458_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_105 VNB N_VGND_c_1459_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_106 VNB N_VGND_c_1460_n 0.623946f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_107 VPB N_A_c_218_n 0.0208611f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=1.765
cc_108 VPB N_A_c_219_n 0.0155109f $X=-0.19 $Y=1.66 $X2=0.96 $Y2=1.765
cc_109 VPB N_A_c_220_n 0.0158647f $X=-0.19 $Y=1.66 $X2=1.41 $Y2=1.765
cc_110 VPB N_A_c_216_n 0.0138362f $X=-0.19 $Y=1.66 $X2=1.265 $Y2=1.515
cc_111 VPB N_A_c_217_n 0.0344244f $X=-0.19 $Y=1.66 $X2=1.41 $Y2=1.557
cc_112 VPB N_A_27_74#_c_298_n 0.0161509f $X=-0.19 $Y=1.66 $X2=1.41 $Y2=2.4
cc_113 VPB N_A_27_74#_c_299_n 0.015404f $X=-0.19 $Y=1.66 $X2=1.115 $Y2=1.58
cc_114 VPB N_A_27_74#_c_300_n 0.015247f $X=-0.19 $Y=1.66 $X2=0.585 $Y2=1.515
cc_115 VPB N_A_27_74#_c_301_n 0.0152262f $X=-0.19 $Y=1.66 $X2=1.41 $Y2=1.557
cc_116 VPB N_A_27_74#_c_302_n 0.0151048f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_117 VPB N_A_27_74#_c_285_n 0.0321912f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_118 VPB N_A_27_74#_c_287_n 6.28632e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_119 VPB N_A_27_74#_c_305_n 0.0205263f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_120 VPB N_A_27_74#_c_306_n 0.00739392f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_121 VPB N_A_27_74#_c_307_n 0.0353617f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_122 VPB N_A_27_74#_c_308_n 0.00257348f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_123 VPB N_A_27_74#_c_294_n 0.00286675f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_124 VPB N_A_384_74#_c_513_n 0.0155385f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_125 VPB N_A_384_74#_c_514_n 0.0154822f $X=-0.19 $Y=1.66 $X2=0.585 $Y2=1.557
cc_126 VPB N_A_384_74#_c_515_n 0.0152343f $X=-0.19 $Y=1.66 $X2=1.265 $Y2=1.515
cc_127 VPB N_A_384_74#_c_516_n 0.0154843f $X=-0.19 $Y=1.66 $X2=0.72 $Y2=1.565
cc_128 VPB N_A_384_74#_c_517_n 0.0152359f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_129 VPB N_A_384_74#_c_518_n 0.0154835f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_130 VPB N_A_384_74#_c_519_n 0.0152376f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_131 VPB N_A_384_74#_c_520_n 0.0154831f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_132 VPB N_A_384_74#_c_521_n 0.0154832f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_133 VPB N_A_384_74#_c_522_n 0.0158611f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_134 VPB N_A_384_74#_c_523_n 0.0156162f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_135 VPB N_A_384_74#_c_524_n 0.0158608f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_136 VPB N_A_384_74#_c_525_n 0.0156138f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_137 VPB N_A_384_74#_c_526_n 0.0155607f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_138 VPB N_A_384_74#_c_527_n 0.0157582f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_139 VPB N_A_384_74#_c_528_n 0.0178344f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_140 VPB N_A_384_74#_c_529_n 0.00291084f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_141 VPB N_A_384_74#_c_530_n 0.00179527f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_142 VPB N_A_384_74#_c_531_n 0.00231059f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_143 VPB N_A_384_74#_c_532_n 0.00257348f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_144 VPB N_A_384_74#_c_533_n 0.00222134f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_145 VPB N_A_384_74#_c_502_n 0.00165499f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_146 VPB N_A_384_74#_c_535_n 0.00257348f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_147 VPB N_A_384_74#_c_536_n 0.00183475f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_148 VPB N_A_384_74#_c_504_n 0.0190681f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_149 VPB N_A_384_74#_c_505_n 0.00147325f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_150 VPB N_A_384_74#_c_506_n 0.00153481f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_151 VPB N_A_384_74#_c_507_n 0.00192338f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_152 VPB N_A_384_74#_c_508_n 0.00218971f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_153 VPB N_A_384_74#_c_509_n 0.0019973f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_154 VPB N_A_384_74#_c_510_n 0.00173921f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_155 VPB N_A_384_74#_c_511_n 0.00195978f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_156 VPB N_A_384_74#_c_512_n 0.0971517f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_157 VPB N_VPWR_c_937_n 0.00799266f $X=-0.19 $Y=1.66 $X2=0.72 $Y2=1.565
cc_158 VPB N_VPWR_c_938_n 0.00799648f $X=-0.19 $Y=1.66 $X2=1.265 $Y2=1.565
cc_159 VPB N_VPWR_c_939_n 0.00799266f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_160 VPB N_VPWR_c_940_n 0.00799266f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_161 VPB N_VPWR_c_941_n 0.00799266f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_162 VPB N_VPWR_c_942_n 0.00799266f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_163 VPB N_VPWR_c_943_n 0.00799266f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_164 VPB N_VPWR_c_944_n 0.00799266f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_165 VPB N_VPWR_c_945_n 0.0206041f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_166 VPB N_VPWR_c_946_n 0.00799266f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_167 VPB N_VPWR_c_947_n 0.00864533f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_168 VPB N_VPWR_c_948_n 0.00875168f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_169 VPB N_VPWR_c_949_n 0.00851573f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_170 VPB N_VPWR_c_950_n 0.0111306f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_171 VPB N_VPWR_c_951_n 0.0645756f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_172 VPB N_VPWR_c_952_n 0.0206041f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_173 VPB N_VPWR_c_953_n 0.00324402f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_174 VPB N_VPWR_c_954_n 0.0212406f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_175 VPB N_VPWR_c_955_n 0.00324402f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_176 VPB N_VPWR_c_956_n 0.0206041f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_177 VPB N_VPWR_c_957_n 0.00324402f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_178 VPB N_VPWR_c_958_n 0.0206041f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_179 VPB N_VPWR_c_959_n 0.00319223f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_180 VPB N_VPWR_c_960_n 0.0206041f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_181 VPB N_VPWR_c_961_n 0.00324402f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_182 VPB N_VPWR_c_962_n 0.0206041f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_183 VPB N_VPWR_c_963_n 0.00324402f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_184 VPB N_VPWR_c_964_n 0.0206041f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_185 VPB N_VPWR_c_965_n 0.00324402f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_186 VPB N_VPWR_c_966_n 0.0206041f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_187 VPB N_VPWR_c_967_n 0.020445f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_188 VPB N_VPWR_c_968_n 0.0201268f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_189 VPB N_VPWR_c_969_n 0.0207632f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_190 VPB N_VPWR_c_970_n 0.0234893f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_191 VPB N_VPWR_c_971_n 0.00324402f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_192 VPB N_VPWR_c_972_n 0.00430193f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_193 VPB N_VPWR_c_973_n 0.00449427f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_194 VPB N_VPWR_c_974_n 0.00410958f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_195 VPB N_VPWR_c_936_n 0.141449f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_196 VPB N_Y_c_1159_n 0.00109191f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_197 VPB N_Y_c_1160_n 0.00127905f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_198 VPB N_Y_c_1161_n 0.00129336f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_199 VPB N_Y_c_1162_n 0.0012737f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_200 VPB N_Y_c_1171_n 0.00257348f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_201 VPB N_Y_c_1172_n 0.00257348f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_202 VPB N_Y_c_1163_n 0.00200376f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_203 VPB N_Y_c_1174_n 0.00257348f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_204 VPB N_Y_c_1164_n 0.00126528f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_205 VPB N_Y_c_1165_n 0.00126894f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_206 VPB N_Y_c_1166_n 0.00126218f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_207 VPB N_Y_c_1178_n 2.17058e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_208 VPB N_Y_c_1179_n 0.00257348f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_209 VPB N_Y_c_1180_n 0.00257348f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_210 VPB N_Y_c_1181_n 0.00257348f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_211 VPB N_Y_c_1182_n 0.00257348f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_212 VPB N_Y_c_1183_n 0.00290896f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_213 N_A_M1043_g N_A_27_74#_M1010_g 0.0296537f $X=1.415 $Y=0.74 $X2=0 $Y2=0
cc_214 N_A_c_220_n N_A_27_74#_c_298_n 0.021493f $X=1.41 $Y=1.765 $X2=0 $Y2=0
cc_215 N_A_c_217_n N_A_27_74#_c_285_n 0.0186443f $X=1.41 $Y=1.557 $X2=0 $Y2=0
cc_216 N_A_M1002_g N_A_27_74#_c_289_n 0.00159319f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_217 N_A_c_218_n N_A_27_74#_c_306_n 4.27055e-19 $X=0.51 $Y=1.765 $X2=0 $Y2=0
cc_218 N_A_c_216_n N_A_27_74#_c_306_n 0.0260502f $X=1.265 $Y=1.515 $X2=0 $Y2=0
cc_219 N_A_c_218_n N_A_27_74#_c_307_n 0.0104891f $X=0.51 $Y=1.765 $X2=0 $Y2=0
cc_220 N_A_c_219_n N_A_27_74#_c_307_n 6.45594e-19 $X=0.96 $Y=1.765 $X2=0 $Y2=0
cc_221 N_A_M1002_g N_A_27_74#_c_290_n 0.013995f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_222 N_A_M1030_g N_A_27_74#_c_290_n 0.0141485f $X=0.985 $Y=0.74 $X2=0 $Y2=0
cc_223 N_A_c_216_n N_A_27_74#_c_290_n 0.056571f $X=1.265 $Y=1.515 $X2=0 $Y2=0
cc_224 N_A_c_217_n N_A_27_74#_c_290_n 0.00358729f $X=1.41 $Y=1.557 $X2=0 $Y2=0
cc_225 N_A_c_216_n N_A_27_74#_c_291_n 0.0216404f $X=1.265 $Y=1.515 $X2=0 $Y2=0
cc_226 N_A_c_218_n N_A_27_74#_c_323_n 0.0120074f $X=0.51 $Y=1.765 $X2=0 $Y2=0
cc_227 N_A_c_219_n N_A_27_74#_c_323_n 0.0120074f $X=0.96 $Y=1.765 $X2=0 $Y2=0
cc_228 N_A_c_216_n N_A_27_74#_c_323_n 0.0393875f $X=1.265 $Y=1.515 $X2=0 $Y2=0
cc_229 N_A_c_217_n N_A_27_74#_c_323_n 0.00131283f $X=1.41 $Y=1.557 $X2=0 $Y2=0
cc_230 N_A_c_218_n N_A_27_74#_c_308_n 6.45594e-19 $X=0.51 $Y=1.765 $X2=0 $Y2=0
cc_231 N_A_c_219_n N_A_27_74#_c_308_n 0.0103431f $X=0.96 $Y=1.765 $X2=0 $Y2=0
cc_232 N_A_c_220_n N_A_27_74#_c_308_n 0.0103958f $X=1.41 $Y=1.765 $X2=0 $Y2=0
cc_233 N_A_M1030_g N_A_27_74#_c_292_n 4.0877e-19 $X=0.985 $Y=0.74 $X2=0 $Y2=0
cc_234 N_A_M1043_g N_A_27_74#_c_292_n 3.92313e-19 $X=1.415 $Y=0.74 $X2=0 $Y2=0
cc_235 N_A_M1043_g N_A_27_74#_c_293_n 0.0139804f $X=1.415 $Y=0.74 $X2=0 $Y2=0
cc_236 N_A_c_216_n N_A_27_74#_c_293_n 0.0107488f $X=1.265 $Y=1.515 $X2=0 $Y2=0
cc_237 N_A_c_217_n N_A_27_74#_c_293_n 3.86519e-19 $X=1.41 $Y=1.557 $X2=0 $Y2=0
cc_238 N_A_c_220_n N_A_27_74#_c_335_n 0.0133449f $X=1.41 $Y=1.765 $X2=0 $Y2=0
cc_239 N_A_c_216_n N_A_27_74#_c_335_n 0.00580317f $X=1.265 $Y=1.515 $X2=0 $Y2=0
cc_240 N_A_c_220_n N_A_27_74#_c_294_n 0.00389155f $X=1.41 $Y=1.765 $X2=0 $Y2=0
cc_241 N_A_c_219_n N_A_27_74#_c_338_n 4.27055e-19 $X=0.96 $Y=1.765 $X2=0 $Y2=0
cc_242 N_A_c_220_n N_A_27_74#_c_338_n 4.27055e-19 $X=1.41 $Y=1.765 $X2=0 $Y2=0
cc_243 N_A_c_216_n N_A_27_74#_c_338_n 0.0237598f $X=1.265 $Y=1.515 $X2=0 $Y2=0
cc_244 N_A_c_217_n N_A_27_74#_c_338_n 0.00144162f $X=1.41 $Y=1.557 $X2=0 $Y2=0
cc_245 N_A_c_216_n N_A_27_74#_c_296_n 0.0146029f $X=1.265 $Y=1.515 $X2=0 $Y2=0
cc_246 N_A_c_217_n N_A_27_74#_c_296_n 0.00232957f $X=1.41 $Y=1.557 $X2=0 $Y2=0
cc_247 N_A_M1043_g N_A_27_74#_c_297_n 0.0040282f $X=1.415 $Y=0.74 $X2=0 $Y2=0
cc_248 N_A_c_216_n N_A_27_74#_c_297_n 0.0341212f $X=1.265 $Y=1.515 $X2=0 $Y2=0
cc_249 N_A_c_217_n N_A_27_74#_c_297_n 0.00314078f $X=1.41 $Y=1.557 $X2=0 $Y2=0
cc_250 N_A_c_218_n N_VPWR_c_937_n 0.00486623f $X=0.51 $Y=1.765 $X2=0 $Y2=0
cc_251 N_A_c_219_n N_VPWR_c_937_n 0.00486623f $X=0.96 $Y=1.765 $X2=0 $Y2=0
cc_252 N_A_c_220_n N_VPWR_c_938_n 0.00486623f $X=1.41 $Y=1.765 $X2=0 $Y2=0
cc_253 N_A_c_219_n N_VPWR_c_952_n 0.00445602f $X=0.96 $Y=1.765 $X2=0 $Y2=0
cc_254 N_A_c_220_n N_VPWR_c_952_n 0.00445602f $X=1.41 $Y=1.765 $X2=0 $Y2=0
cc_255 N_A_c_218_n N_VPWR_c_970_n 0.00445602f $X=0.51 $Y=1.765 $X2=0 $Y2=0
cc_256 N_A_c_218_n N_VPWR_c_936_n 0.008611f $X=0.51 $Y=1.765 $X2=0 $Y2=0
cc_257 N_A_c_219_n N_VPWR_c_936_n 0.00857589f $X=0.96 $Y=1.765 $X2=0 $Y2=0
cc_258 N_A_c_220_n N_VPWR_c_936_n 0.00857673f $X=1.41 $Y=1.765 $X2=0 $Y2=0
cc_259 N_A_M1002_g N_VGND_c_1421_n 0.0136841f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_260 N_A_M1030_g N_VGND_c_1421_n 0.00425844f $X=0.985 $Y=0.74 $X2=0 $Y2=0
cc_261 N_A_M1030_g N_VGND_c_1422_n 4.80113e-19 $X=0.985 $Y=0.74 $X2=0 $Y2=0
cc_262 N_A_M1043_g N_VGND_c_1422_n 0.0107133f $X=1.415 $Y=0.74 $X2=0 $Y2=0
cc_263 N_A_M1002_g N_VGND_c_1443_n 0.00383152f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_264 N_A_M1030_g N_VGND_c_1444_n 0.00461464f $X=0.985 $Y=0.74 $X2=0 $Y2=0
cc_265 N_A_M1043_g N_VGND_c_1444_n 0.00383152f $X=1.415 $Y=0.74 $X2=0 $Y2=0
cc_266 N_A_M1002_g N_VGND_c_1460_n 0.00761198f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_267 N_A_M1030_g N_VGND_c_1460_n 0.00908454f $X=0.985 $Y=0.74 $X2=0 $Y2=0
cc_268 N_A_M1043_g N_VGND_c_1460_n 0.0075754f $X=1.415 $Y=0.74 $X2=0 $Y2=0
cc_269 N_A_27_74#_M1049_g N_A_384_74#_M1003_g 0.020096f $X=4.065 $Y=0.74 $X2=0
+ $Y2=0
cc_270 N_A_27_74#_c_305_n N_A_384_74#_c_513_n 0.00894101f $X=4.13 $Y=1.765 $X2=0
+ $Y2=0
cc_271 N_A_27_74#_c_298_n N_A_384_74#_c_529_n 4.53719e-19 $X=1.86 $Y=1.765 $X2=0
+ $Y2=0
cc_272 N_A_27_74#_c_299_n N_A_384_74#_c_529_n 0.0124249f $X=2.33 $Y=1.765 $X2=0
+ $Y2=0
cc_273 N_A_27_74#_c_300_n N_A_384_74#_c_529_n 6.9119e-19 $X=2.78 $Y=1.765 $X2=0
+ $Y2=0
cc_274 N_A_27_74#_M1010_g N_A_384_74#_c_496_n 3.92313e-19 $X=1.845 $Y=0.74 $X2=0
+ $Y2=0
cc_275 N_A_27_74#_M1014_g N_A_384_74#_c_496_n 3.92313e-19 $X=2.275 $Y=0.74 $X2=0
+ $Y2=0
cc_276 N_A_27_74#_M1014_g N_A_384_74#_c_497_n 0.0124383f $X=2.275 $Y=0.74 $X2=0
+ $Y2=0
cc_277 N_A_27_74#_M1016_g N_A_384_74#_c_497_n 0.0111034f $X=2.705 $Y=0.74 $X2=0
+ $Y2=0
cc_278 N_A_27_74#_c_285_n N_A_384_74#_c_497_n 0.00224206f $X=3.77 $Y=1.375 $X2=0
+ $Y2=0
cc_279 N_A_27_74#_c_295_n N_A_384_74#_c_497_n 0.0447482f $X=3.295 $Y=1.465 $X2=0
+ $Y2=0
cc_280 N_A_27_74#_c_285_n N_A_384_74#_c_498_n 0.00232957f $X=3.77 $Y=1.375 $X2=0
+ $Y2=0
cc_281 N_A_27_74#_c_295_n N_A_384_74#_c_498_n 0.0143381f $X=3.295 $Y=1.465 $X2=0
+ $Y2=0
cc_282 N_A_27_74#_c_297_n N_A_384_74#_c_498_n 0.00140469f $X=1.685 $Y=1.095
+ $X2=0 $Y2=0
cc_283 N_A_27_74#_c_299_n N_A_384_74#_c_530_n 0.0120074f $X=2.33 $Y=1.765 $X2=0
+ $Y2=0
cc_284 N_A_27_74#_c_300_n N_A_384_74#_c_530_n 0.0120074f $X=2.78 $Y=1.765 $X2=0
+ $Y2=0
cc_285 N_A_27_74#_c_285_n N_A_384_74#_c_530_n 0.00765052f $X=3.77 $Y=1.375 $X2=0
+ $Y2=0
cc_286 N_A_27_74#_c_295_n N_A_384_74#_c_530_n 0.0417603f $X=3.295 $Y=1.465 $X2=0
+ $Y2=0
cc_287 N_A_27_74#_c_298_n N_A_384_74#_c_531_n 3.7798e-19 $X=1.86 $Y=1.765 $X2=0
+ $Y2=0
cc_288 N_A_27_74#_c_299_n N_A_384_74#_c_531_n 8.95482e-19 $X=2.33 $Y=1.765 $X2=0
+ $Y2=0
cc_289 N_A_27_74#_c_285_n N_A_384_74#_c_531_n 0.00830678f $X=3.77 $Y=1.375 $X2=0
+ $Y2=0
cc_290 N_A_27_74#_c_294_n N_A_384_74#_c_531_n 0.00329154f $X=1.685 $Y=1.95 $X2=0
+ $Y2=0
cc_291 N_A_27_74#_c_295_n N_A_384_74#_c_531_n 0.027762f $X=3.295 $Y=1.465 $X2=0
+ $Y2=0
cc_292 N_A_27_74#_M1014_g N_A_384_74#_c_499_n 6.20738e-19 $X=2.275 $Y=0.74 $X2=0
+ $Y2=0
cc_293 N_A_27_74#_M1016_g N_A_384_74#_c_499_n 0.00866629f $X=2.705 $Y=0.74 $X2=0
+ $Y2=0
cc_294 N_A_27_74#_M1024_g N_A_384_74#_c_499_n 3.97481e-19 $X=3.135 $Y=0.74 $X2=0
+ $Y2=0
cc_295 N_A_27_74#_c_299_n N_A_384_74#_c_532_n 6.9119e-19 $X=2.33 $Y=1.765 $X2=0
+ $Y2=0
cc_296 N_A_27_74#_c_300_n N_A_384_74#_c_532_n 0.0125029f $X=2.78 $Y=1.765 $X2=0
+ $Y2=0
cc_297 N_A_27_74#_c_301_n N_A_384_74#_c_532_n 0.0125029f $X=3.23 $Y=1.765 $X2=0
+ $Y2=0
cc_298 N_A_27_74#_c_302_n N_A_384_74#_c_532_n 6.9119e-19 $X=3.68 $Y=1.765 $X2=0
+ $Y2=0
cc_299 N_A_27_74#_M1024_g N_A_384_74#_c_500_n 0.0128832f $X=3.135 $Y=0.74 $X2=0
+ $Y2=0
cc_300 N_A_27_74#_M1046_g N_A_384_74#_c_500_n 0.0132728f $X=3.635 $Y=0.74 $X2=0
+ $Y2=0
cc_301 N_A_27_74#_c_285_n N_A_384_74#_c_500_n 0.00390513f $X=3.77 $Y=1.375 $X2=0
+ $Y2=0
cc_302 N_A_27_74#_c_295_n N_A_384_74#_c_500_n 0.0335994f $X=3.295 $Y=1.465 $X2=0
+ $Y2=0
cc_303 N_A_27_74#_c_301_n N_A_384_74#_c_533_n 0.0120074f $X=3.23 $Y=1.765 $X2=0
+ $Y2=0
cc_304 N_A_27_74#_c_302_n N_A_384_74#_c_533_n 0.0137394f $X=3.68 $Y=1.765 $X2=0
+ $Y2=0
cc_305 N_A_27_74#_c_285_n N_A_384_74#_c_533_n 0.00814778f $X=3.77 $Y=1.375 $X2=0
+ $Y2=0
cc_306 N_A_27_74#_c_295_n N_A_384_74#_c_533_n 0.0212559f $X=3.295 $Y=1.465 $X2=0
+ $Y2=0
cc_307 N_A_27_74#_M1024_g N_A_384_74#_c_501_n 8.7513e-19 $X=3.135 $Y=0.74 $X2=0
+ $Y2=0
cc_308 N_A_27_74#_M1046_g N_A_384_74#_c_501_n 0.00862472f $X=3.635 $Y=0.74 $X2=0
+ $Y2=0
cc_309 N_A_27_74#_M1049_g N_A_384_74#_c_501_n 3.97481e-19 $X=4.065 $Y=0.74 $X2=0
+ $Y2=0
cc_310 N_A_27_74#_M1024_g N_A_384_74#_c_502_n 8.02787e-19 $X=3.135 $Y=0.74 $X2=0
+ $Y2=0
cc_311 N_A_27_74#_M1046_g N_A_384_74#_c_502_n 0.00529244f $X=3.635 $Y=0.74 $X2=0
+ $Y2=0
cc_312 N_A_27_74#_c_302_n N_A_384_74#_c_502_n 0.00176384f $X=3.68 $Y=1.765 $X2=0
+ $Y2=0
cc_313 N_A_27_74#_c_284_n N_A_384_74#_c_502_n 0.0105749f $X=3.99 $Y=1.375 $X2=0
+ $Y2=0
cc_314 N_A_27_74#_c_285_n N_A_384_74#_c_502_n 0.0158909f $X=3.77 $Y=1.375 $X2=0
+ $Y2=0
cc_315 N_A_27_74#_M1049_g N_A_384_74#_c_502_n 0.00453721f $X=4.065 $Y=0.74 $X2=0
+ $Y2=0
cc_316 N_A_27_74#_c_287_n N_A_384_74#_c_502_n 0.00827465f $X=4.13 $Y=1.675 $X2=0
+ $Y2=0
cc_317 N_A_27_74#_c_305_n N_A_384_74#_c_502_n 0.0133061f $X=4.13 $Y=1.765 $X2=0
+ $Y2=0
cc_318 N_A_27_74#_c_288_n N_A_384_74#_c_502_n 0.0113158f $X=4.105 $Y=1.375 $X2=0
+ $Y2=0
cc_319 N_A_27_74#_c_295_n N_A_384_74#_c_502_n 0.0185957f $X=3.295 $Y=1.465 $X2=0
+ $Y2=0
cc_320 N_A_27_74#_c_301_n N_A_384_74#_c_535_n 6.9119e-19 $X=3.23 $Y=1.765 $X2=0
+ $Y2=0
cc_321 N_A_27_74#_c_302_n N_A_384_74#_c_535_n 0.0125029f $X=3.68 $Y=1.765 $X2=0
+ $Y2=0
cc_322 N_A_27_74#_c_305_n N_A_384_74#_c_535_n 0.0112516f $X=4.13 $Y=1.765 $X2=0
+ $Y2=0
cc_323 N_A_27_74#_M1016_g N_A_384_74#_c_503_n 9.7541e-19 $X=2.705 $Y=0.74 $X2=0
+ $Y2=0
cc_324 N_A_27_74#_c_285_n N_A_384_74#_c_503_n 0.00232957f $X=3.77 $Y=1.375 $X2=0
+ $Y2=0
cc_325 N_A_27_74#_c_295_n N_A_384_74#_c_503_n 0.0209731f $X=3.295 $Y=1.465 $X2=0
+ $Y2=0
cc_326 N_A_27_74#_c_300_n N_A_384_74#_c_536_n 9.3899e-19 $X=2.78 $Y=1.765 $X2=0
+ $Y2=0
cc_327 N_A_27_74#_c_301_n N_A_384_74#_c_536_n 9.3899e-19 $X=3.23 $Y=1.765 $X2=0
+ $Y2=0
cc_328 N_A_27_74#_c_285_n N_A_384_74#_c_536_n 0.00792231f $X=3.77 $Y=1.375 $X2=0
+ $Y2=0
cc_329 N_A_27_74#_c_295_n N_A_384_74#_c_536_n 0.0276943f $X=3.295 $Y=1.465 $X2=0
+ $Y2=0
cc_330 N_A_27_74#_c_305_n N_A_384_74#_c_504_n 0.00269092f $X=4.13 $Y=1.765 $X2=0
+ $Y2=0
cc_331 N_A_27_74#_c_288_n N_A_384_74#_c_512_n 0.0226086f $X=4.105 $Y=1.375 $X2=0
+ $Y2=0
cc_332 N_A_27_74#_c_323_n N_VPWR_M1015_s 0.00408911f $X=1.02 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_333 N_A_27_74#_c_335_n N_VPWR_M1022_s 0.00533313f $X=1.6 $Y=2.035 $X2=0 $Y2=0
cc_334 N_A_27_74#_c_294_n N_VPWR_M1022_s 0.00160462f $X=1.685 $Y=1.95 $X2=0
+ $Y2=0
cc_335 N_A_27_74#_c_307_n N_VPWR_c_937_n 0.0449718f $X=0.285 $Y=2.815 $X2=0
+ $Y2=0
cc_336 N_A_27_74#_c_323_n N_VPWR_c_937_n 0.0136682f $X=1.02 $Y=2.035 $X2=0 $Y2=0
cc_337 N_A_27_74#_c_308_n N_VPWR_c_937_n 0.0449718f $X=1.185 $Y=2.815 $X2=0
+ $Y2=0
cc_338 N_A_27_74#_c_298_n N_VPWR_c_938_n 0.0050615f $X=1.86 $Y=1.765 $X2=0 $Y2=0
cc_339 N_A_27_74#_c_308_n N_VPWR_c_938_n 0.0449718f $X=1.185 $Y=2.815 $X2=0
+ $Y2=0
cc_340 N_A_27_74#_c_335_n N_VPWR_c_938_n 0.0146343f $X=1.6 $Y=2.035 $X2=0 $Y2=0
cc_341 N_A_27_74#_c_299_n N_VPWR_c_939_n 0.00586501f $X=2.33 $Y=1.765 $X2=0
+ $Y2=0
cc_342 N_A_27_74#_c_300_n N_VPWR_c_939_n 0.00586501f $X=2.78 $Y=1.765 $X2=0
+ $Y2=0
cc_343 N_A_27_74#_c_301_n N_VPWR_c_940_n 0.00586501f $X=3.23 $Y=1.765 $X2=0
+ $Y2=0
cc_344 N_A_27_74#_c_302_n N_VPWR_c_940_n 0.00586501f $X=3.68 $Y=1.765 $X2=0
+ $Y2=0
cc_345 N_A_27_74#_c_305_n N_VPWR_c_941_n 0.00603265f $X=4.13 $Y=1.765 $X2=0
+ $Y2=0
cc_346 N_A_27_74#_c_308_n N_VPWR_c_952_n 0.014552f $X=1.185 $Y=2.815 $X2=0 $Y2=0
cc_347 N_A_27_74#_c_298_n N_VPWR_c_954_n 0.00461464f $X=1.86 $Y=1.765 $X2=0
+ $Y2=0
cc_348 N_A_27_74#_c_299_n N_VPWR_c_954_n 0.00445602f $X=2.33 $Y=1.765 $X2=0
+ $Y2=0
cc_349 N_A_27_74#_c_300_n N_VPWR_c_956_n 0.00445602f $X=2.78 $Y=1.765 $X2=0
+ $Y2=0
cc_350 N_A_27_74#_c_301_n N_VPWR_c_956_n 0.00445602f $X=3.23 $Y=1.765 $X2=0
+ $Y2=0
cc_351 N_A_27_74#_c_302_n N_VPWR_c_958_n 0.00445602f $X=3.68 $Y=1.765 $X2=0
+ $Y2=0
cc_352 N_A_27_74#_c_305_n N_VPWR_c_958_n 0.00445602f $X=4.13 $Y=1.765 $X2=0
+ $Y2=0
cc_353 N_A_27_74#_c_307_n N_VPWR_c_970_n 0.0145938f $X=0.285 $Y=2.815 $X2=0
+ $Y2=0
cc_354 N_A_27_74#_c_298_n N_VPWR_c_936_n 0.00909224f $X=1.86 $Y=1.765 $X2=0
+ $Y2=0
cc_355 N_A_27_74#_c_299_n N_VPWR_c_936_n 0.00857779f $X=2.33 $Y=1.765 $X2=0
+ $Y2=0
cc_356 N_A_27_74#_c_300_n N_VPWR_c_936_n 0.00857589f $X=2.78 $Y=1.765 $X2=0
+ $Y2=0
cc_357 N_A_27_74#_c_301_n N_VPWR_c_936_n 0.00857589f $X=3.23 $Y=1.765 $X2=0
+ $Y2=0
cc_358 N_A_27_74#_c_302_n N_VPWR_c_936_n 0.00857589f $X=3.68 $Y=1.765 $X2=0
+ $Y2=0
cc_359 N_A_27_74#_c_305_n N_VPWR_c_936_n 0.00857673f $X=4.13 $Y=1.765 $X2=0
+ $Y2=0
cc_360 N_A_27_74#_c_307_n N_VPWR_c_936_n 0.0120466f $X=0.285 $Y=2.815 $X2=0
+ $Y2=0
cc_361 N_A_27_74#_c_308_n N_VPWR_c_936_n 0.0119791f $X=1.185 $Y=2.815 $X2=0
+ $Y2=0
cc_362 N_A_27_74#_M1049_g N_Y_c_1159_n 0.0010331f $X=4.065 $Y=0.74 $X2=0 $Y2=0
cc_363 N_A_27_74#_c_305_n N_Y_c_1159_n 4.88979e-19 $X=4.13 $Y=1.765 $X2=0 $Y2=0
cc_364 N_A_27_74#_c_288_n N_Y_c_1159_n 4.12512e-19 $X=4.105 $Y=1.375 $X2=0 $Y2=0
cc_365 N_A_27_74#_c_290_n N_VGND_M1002_s 0.00240242f $X=1.115 $Y=1.095 $X2=-0.19
+ $Y2=-0.245
cc_366 N_A_27_74#_c_293_n N_VGND_M1043_s 8.02634e-19 $X=1.6 $Y=1.095 $X2=0 $Y2=0
cc_367 N_A_27_74#_c_297_n N_VGND_M1043_s 0.00168914f $X=1.685 $Y=1.095 $X2=0
+ $Y2=0
cc_368 N_A_27_74#_c_289_n N_VGND_c_1421_n 0.0182902f $X=0.28 $Y=0.515 $X2=0
+ $Y2=0
cc_369 N_A_27_74#_c_290_n N_VGND_c_1421_n 0.0201731f $X=1.115 $Y=1.095 $X2=0
+ $Y2=0
cc_370 N_A_27_74#_c_292_n N_VGND_c_1421_n 0.00118247f $X=1.2 $Y=0.515 $X2=0
+ $Y2=0
cc_371 N_A_27_74#_M1010_g N_VGND_c_1422_n 0.0108544f $X=1.845 $Y=0.74 $X2=0
+ $Y2=0
cc_372 N_A_27_74#_M1014_g N_VGND_c_1422_n 4.71636e-19 $X=2.275 $Y=0.74 $X2=0
+ $Y2=0
cc_373 N_A_27_74#_c_292_n N_VGND_c_1422_n 0.0182488f $X=1.2 $Y=0.515 $X2=0 $Y2=0
cc_374 N_A_27_74#_c_293_n N_VGND_c_1422_n 0.00609809f $X=1.6 $Y=1.095 $X2=0
+ $Y2=0
cc_375 N_A_27_74#_c_295_n N_VGND_c_1422_n 8.33225e-19 $X=3.295 $Y=1.465 $X2=0
+ $Y2=0
cc_376 N_A_27_74#_c_297_n N_VGND_c_1422_n 0.0100981f $X=1.685 $Y=1.095 $X2=0
+ $Y2=0
cc_377 N_A_27_74#_M1010_g N_VGND_c_1423_n 4.57991e-19 $X=1.845 $Y=0.74 $X2=0
+ $Y2=0
cc_378 N_A_27_74#_M1014_g N_VGND_c_1423_n 0.00900784f $X=2.275 $Y=0.74 $X2=0
+ $Y2=0
cc_379 N_A_27_74#_M1016_g N_VGND_c_1423_n 0.00183835f $X=2.705 $Y=0.74 $X2=0
+ $Y2=0
cc_380 N_A_27_74#_M1016_g N_VGND_c_1424_n 5.04273e-19 $X=2.705 $Y=0.74 $X2=0
+ $Y2=0
cc_381 N_A_27_74#_M1024_g N_VGND_c_1424_n 0.0097054f $X=3.135 $Y=0.74 $X2=0
+ $Y2=0
cc_382 N_A_27_74#_M1046_g N_VGND_c_1424_n 0.00397833f $X=3.635 $Y=0.74 $X2=0
+ $Y2=0
cc_383 N_A_27_74#_M1046_g N_VGND_c_1425_n 6.13182e-19 $X=3.635 $Y=0.74 $X2=0
+ $Y2=0
cc_384 N_A_27_74#_M1049_g N_VGND_c_1425_n 0.0134222f $X=4.065 $Y=0.74 $X2=0
+ $Y2=0
cc_385 N_A_27_74#_c_288_n N_VGND_c_1425_n 6.26412e-19 $X=4.105 $Y=1.375 $X2=0
+ $Y2=0
cc_386 N_A_27_74#_M1010_g N_VGND_c_1435_n 0.00383152f $X=1.845 $Y=0.74 $X2=0
+ $Y2=0
cc_387 N_A_27_74#_M1014_g N_VGND_c_1435_n 0.00383152f $X=2.275 $Y=0.74 $X2=0
+ $Y2=0
cc_388 N_A_27_74#_M1016_g N_VGND_c_1437_n 0.00434272f $X=2.705 $Y=0.74 $X2=0
+ $Y2=0
cc_389 N_A_27_74#_M1024_g N_VGND_c_1437_n 0.00383152f $X=3.135 $Y=0.74 $X2=0
+ $Y2=0
cc_390 N_A_27_74#_M1046_g N_VGND_c_1439_n 0.00434272f $X=3.635 $Y=0.74 $X2=0
+ $Y2=0
cc_391 N_A_27_74#_M1049_g N_VGND_c_1439_n 0.00383152f $X=4.065 $Y=0.74 $X2=0
+ $Y2=0
cc_392 N_A_27_74#_c_289_n N_VGND_c_1443_n 0.011066f $X=0.28 $Y=0.515 $X2=0 $Y2=0
cc_393 N_A_27_74#_c_292_n N_VGND_c_1444_n 0.00749631f $X=1.2 $Y=0.515 $X2=0
+ $Y2=0
cc_394 N_A_27_74#_M1010_g N_VGND_c_1460_n 0.0075754f $X=1.845 $Y=0.74 $X2=0
+ $Y2=0
cc_395 N_A_27_74#_M1014_g N_VGND_c_1460_n 0.0075754f $X=2.275 $Y=0.74 $X2=0
+ $Y2=0
cc_396 N_A_27_74#_M1016_g N_VGND_c_1460_n 0.00820284f $X=2.705 $Y=0.74 $X2=0
+ $Y2=0
cc_397 N_A_27_74#_M1024_g N_VGND_c_1460_n 0.0075754f $X=3.135 $Y=0.74 $X2=0
+ $Y2=0
cc_398 N_A_27_74#_M1046_g N_VGND_c_1460_n 0.00820718f $X=3.635 $Y=0.74 $X2=0
+ $Y2=0
cc_399 N_A_27_74#_M1049_g N_VGND_c_1460_n 0.0075754f $X=4.065 $Y=0.74 $X2=0
+ $Y2=0
cc_400 N_A_27_74#_c_289_n N_VGND_c_1460_n 0.00915947f $X=0.28 $Y=0.515 $X2=0
+ $Y2=0
cc_401 N_A_27_74#_c_292_n N_VGND_c_1460_n 0.0062048f $X=1.2 $Y=0.515 $X2=0 $Y2=0
cc_402 N_A_384_74#_c_530_n N_VPWR_M1004_d 0.00247267f $X=2.84 $Y=1.885 $X2=0
+ $Y2=0
cc_403 N_A_384_74#_c_533_n N_VPWR_M1026_d 0.00247267f $X=3.74 $Y=1.885 $X2=0
+ $Y2=0
cc_404 N_A_384_74#_c_529_n N_VPWR_c_938_n 0.0213938f $X=2.105 $Y=1.985 $X2=0
+ $Y2=0
cc_405 N_A_384_74#_c_529_n N_VPWR_c_939_n 0.0547423f $X=2.105 $Y=1.985 $X2=0
+ $Y2=0
cc_406 N_A_384_74#_c_530_n N_VPWR_c_939_n 0.0136682f $X=2.84 $Y=1.885 $X2=0
+ $Y2=0
cc_407 N_A_384_74#_c_532_n N_VPWR_c_939_n 0.0547423f $X=3.005 $Y=1.985 $X2=0
+ $Y2=0
cc_408 N_A_384_74#_c_532_n N_VPWR_c_940_n 0.0547423f $X=3.005 $Y=1.985 $X2=0
+ $Y2=0
cc_409 N_A_384_74#_c_533_n N_VPWR_c_940_n 0.0136682f $X=3.74 $Y=1.885 $X2=0
+ $Y2=0
cc_410 N_A_384_74#_c_535_n N_VPWR_c_940_n 0.0547423f $X=3.905 $Y=1.985 $X2=0
+ $Y2=0
cc_411 N_A_384_74#_c_513_n N_VPWR_c_941_n 0.00599728f $X=4.58 $Y=1.765 $X2=0
+ $Y2=0
cc_412 N_A_384_74#_c_502_n N_VPWR_c_941_n 0.0152961f $X=3.905 $Y=1.97 $X2=0
+ $Y2=0
cc_413 N_A_384_74#_c_535_n N_VPWR_c_941_n 0.0653172f $X=3.905 $Y=1.985 $X2=0
+ $Y2=0
cc_414 N_A_384_74#_c_504_n N_VPWR_c_941_n 0.00504465f $X=10.71 $Y=1.665 $X2=0
+ $Y2=0
cc_415 N_A_384_74#_c_514_n N_VPWR_c_942_n 0.00592051f $X=5.03 $Y=1.765 $X2=0
+ $Y2=0
cc_416 N_A_384_74#_c_515_n N_VPWR_c_942_n 0.00588387f $X=5.48 $Y=1.765 $X2=0
+ $Y2=0
cc_417 N_A_384_74#_c_504_n N_VPWR_c_942_n 7.18372e-19 $X=10.71 $Y=1.665 $X2=0
+ $Y2=0
cc_418 N_A_384_74#_c_505_n N_VPWR_c_942_n 0.00965197f $X=5.175 $Y=1.465 $X2=0
+ $Y2=0
cc_419 N_A_384_74#_c_512_n N_VPWR_c_942_n 0.00158493f $X=11.435 $Y=1.532 $X2=0
+ $Y2=0
cc_420 N_A_384_74#_c_516_n N_VPWR_c_943_n 0.00592051f $X=5.93 $Y=1.765 $X2=0
+ $Y2=0
cc_421 N_A_384_74#_c_517_n N_VPWR_c_943_n 0.00589619f $X=6.38 $Y=1.765 $X2=0
+ $Y2=0
cc_422 N_A_384_74#_c_504_n N_VPWR_c_943_n 6.09205e-19 $X=10.71 $Y=1.665 $X2=0
+ $Y2=0
cc_423 N_A_384_74#_c_506_n N_VPWR_c_943_n 0.0114663f $X=6.065 $Y=1.465 $X2=0
+ $Y2=0
cc_424 N_A_384_74#_c_512_n N_VPWR_c_943_n 0.00104811f $X=11.435 $Y=1.532 $X2=0
+ $Y2=0
cc_425 N_A_384_74#_c_518_n N_VPWR_c_944_n 0.00592051f $X=6.83 $Y=1.765 $X2=0
+ $Y2=0
cc_426 N_A_384_74#_c_519_n N_VPWR_c_944_n 0.00592051f $X=7.28 $Y=1.765 $X2=0
+ $Y2=0
cc_427 N_A_384_74#_c_504_n N_VPWR_c_944_n 5.65539e-19 $X=10.71 $Y=1.665 $X2=0
+ $Y2=0
cc_428 N_A_384_74#_c_507_n N_VPWR_c_944_n 0.012192f $X=7.005 $Y=1.465 $X2=0
+ $Y2=0
cc_429 N_A_384_74#_c_512_n N_VPWR_c_944_n 8.34596e-19 $X=11.435 $Y=1.532 $X2=0
+ $Y2=0
cc_430 N_A_384_74#_c_519_n N_VPWR_c_945_n 0.00445602f $X=7.28 $Y=1.765 $X2=0
+ $Y2=0
cc_431 N_A_384_74#_c_520_n N_VPWR_c_945_n 0.00445602f $X=7.73 $Y=1.765 $X2=0
+ $Y2=0
cc_432 N_A_384_74#_c_520_n N_VPWR_c_946_n 0.00592051f $X=7.73 $Y=1.765 $X2=0
+ $Y2=0
cc_433 N_A_384_74#_c_521_n N_VPWR_c_946_n 0.00594707f $X=8.18 $Y=1.765 $X2=0
+ $Y2=0
cc_434 N_A_384_74#_c_504_n N_VPWR_c_946_n 5.65539e-19 $X=10.71 $Y=1.665 $X2=0
+ $Y2=0
cc_435 N_A_384_74#_c_508_n N_VPWR_c_946_n 0.012192f $X=7.925 $Y=1.465 $X2=0
+ $Y2=0
cc_436 N_A_384_74#_c_512_n N_VPWR_c_946_n 8.3527e-19 $X=11.435 $Y=1.532 $X2=0
+ $Y2=0
cc_437 N_A_384_74#_c_522_n N_VPWR_c_947_n 0.00633341f $X=8.63 $Y=1.765 $X2=0
+ $Y2=0
cc_438 N_A_384_74#_c_523_n N_VPWR_c_947_n 0.011411f $X=9.13 $Y=1.765 $X2=0 $Y2=0
cc_439 N_A_384_74#_c_504_n N_VPWR_c_947_n 7.50685e-19 $X=10.71 $Y=1.665 $X2=0
+ $Y2=0
cc_440 N_A_384_74#_c_509_n N_VPWR_c_947_n 0.0161834f $X=8.85 $Y=1.465 $X2=0
+ $Y2=0
cc_441 N_A_384_74#_c_512_n N_VPWR_c_947_n 0.00110596f $X=11.435 $Y=1.532 $X2=0
+ $Y2=0
cc_442 N_A_384_74#_c_524_n N_VPWR_c_948_n 0.00638726f $X=9.58 $Y=1.765 $X2=0
+ $Y2=0
cc_443 N_A_384_74#_c_525_n N_VPWR_c_948_n 0.0085568f $X=10.08 $Y=1.765 $X2=0
+ $Y2=0
cc_444 N_A_384_74#_c_504_n N_VPWR_c_948_n 8.28015e-19 $X=10.71 $Y=1.665 $X2=0
+ $Y2=0
cc_445 N_A_384_74#_c_510_n N_VPWR_c_948_n 0.0161834f $X=9.78 $Y=1.465 $X2=0
+ $Y2=0
cc_446 N_A_384_74#_c_512_n N_VPWR_c_948_n 0.00133088f $X=11.435 $Y=1.532 $X2=0
+ $Y2=0
cc_447 N_A_384_74#_c_526_n N_VPWR_c_949_n 0.00621672f $X=10.53 $Y=1.765 $X2=0
+ $Y2=0
cc_448 N_A_384_74#_c_527_n N_VPWR_c_949_n 0.00335732f $X=10.99 $Y=1.765 $X2=0
+ $Y2=0
cc_449 N_A_384_74#_c_504_n N_VPWR_c_949_n 6.194e-19 $X=10.71 $Y=1.665 $X2=0
+ $Y2=0
cc_450 N_A_384_74#_c_511_n N_VPWR_c_949_n 0.0144397f $X=10.71 $Y=1.465 $X2=0
+ $Y2=0
cc_451 N_A_384_74#_c_512_n N_VPWR_c_949_n 0.00127472f $X=11.435 $Y=1.532 $X2=0
+ $Y2=0
cc_452 N_A_384_74#_c_528_n N_VPWR_c_951_n 0.0100916f $X=11.48 $Y=1.765 $X2=0
+ $Y2=0
cc_453 N_A_384_74#_c_529_n N_VPWR_c_954_n 0.0145938f $X=2.105 $Y=1.985 $X2=0
+ $Y2=0
cc_454 N_A_384_74#_c_532_n N_VPWR_c_956_n 0.014552f $X=3.005 $Y=1.985 $X2=0
+ $Y2=0
cc_455 N_A_384_74#_c_535_n N_VPWR_c_958_n 0.014552f $X=3.905 $Y=1.985 $X2=0
+ $Y2=0
cc_456 N_A_384_74#_c_513_n N_VPWR_c_960_n 0.00445602f $X=4.58 $Y=1.765 $X2=0
+ $Y2=0
cc_457 N_A_384_74#_c_514_n N_VPWR_c_960_n 0.00445602f $X=5.03 $Y=1.765 $X2=0
+ $Y2=0
cc_458 N_A_384_74#_c_515_n N_VPWR_c_962_n 0.00445602f $X=5.48 $Y=1.765 $X2=0
+ $Y2=0
cc_459 N_A_384_74#_c_516_n N_VPWR_c_962_n 0.00445602f $X=5.93 $Y=1.765 $X2=0
+ $Y2=0
cc_460 N_A_384_74#_c_517_n N_VPWR_c_964_n 0.00445602f $X=6.38 $Y=1.765 $X2=0
+ $Y2=0
cc_461 N_A_384_74#_c_518_n N_VPWR_c_964_n 0.00445602f $X=6.83 $Y=1.765 $X2=0
+ $Y2=0
cc_462 N_A_384_74#_c_521_n N_VPWR_c_966_n 0.00445602f $X=8.18 $Y=1.765 $X2=0
+ $Y2=0
cc_463 N_A_384_74#_c_522_n N_VPWR_c_966_n 0.00445602f $X=8.63 $Y=1.765 $X2=0
+ $Y2=0
cc_464 N_A_384_74#_c_523_n N_VPWR_c_967_n 0.00445602f $X=9.13 $Y=1.765 $X2=0
+ $Y2=0
cc_465 N_A_384_74#_c_524_n N_VPWR_c_967_n 0.00445602f $X=9.58 $Y=1.765 $X2=0
+ $Y2=0
cc_466 N_A_384_74#_c_525_n N_VPWR_c_968_n 0.00445602f $X=10.08 $Y=1.765 $X2=0
+ $Y2=0
cc_467 N_A_384_74#_c_526_n N_VPWR_c_968_n 0.00445602f $X=10.53 $Y=1.765 $X2=0
+ $Y2=0
cc_468 N_A_384_74#_c_527_n N_VPWR_c_969_n 0.00461464f $X=10.99 $Y=1.765 $X2=0
+ $Y2=0
cc_469 N_A_384_74#_c_528_n N_VPWR_c_969_n 0.00445602f $X=11.48 $Y=1.765 $X2=0
+ $Y2=0
cc_470 N_A_384_74#_c_513_n N_VPWR_c_936_n 0.00857673f $X=4.58 $Y=1.765 $X2=0
+ $Y2=0
cc_471 N_A_384_74#_c_514_n N_VPWR_c_936_n 0.00857589f $X=5.03 $Y=1.765 $X2=0
+ $Y2=0
cc_472 N_A_384_74#_c_515_n N_VPWR_c_936_n 0.00857589f $X=5.48 $Y=1.765 $X2=0
+ $Y2=0
cc_473 N_A_384_74#_c_516_n N_VPWR_c_936_n 0.00857589f $X=5.93 $Y=1.765 $X2=0
+ $Y2=0
cc_474 N_A_384_74#_c_517_n N_VPWR_c_936_n 0.00857589f $X=6.38 $Y=1.765 $X2=0
+ $Y2=0
cc_475 N_A_384_74#_c_518_n N_VPWR_c_936_n 0.00857589f $X=6.83 $Y=1.765 $X2=0
+ $Y2=0
cc_476 N_A_384_74#_c_519_n N_VPWR_c_936_n 0.00857589f $X=7.28 $Y=1.765 $X2=0
+ $Y2=0
cc_477 N_A_384_74#_c_520_n N_VPWR_c_936_n 0.00857589f $X=7.73 $Y=1.765 $X2=0
+ $Y2=0
cc_478 N_A_384_74#_c_521_n N_VPWR_c_936_n 0.00857589f $X=8.18 $Y=1.765 $X2=0
+ $Y2=0
cc_479 N_A_384_74#_c_522_n N_VPWR_c_936_n 0.0085805f $X=8.63 $Y=1.765 $X2=0
+ $Y2=0
cc_480 N_A_384_74#_c_523_n N_VPWR_c_936_n 0.00857938f $X=9.13 $Y=1.765 $X2=0
+ $Y2=0
cc_481 N_A_384_74#_c_524_n N_VPWR_c_936_n 0.0085805f $X=9.58 $Y=1.765 $X2=0
+ $Y2=0
cc_482 N_A_384_74#_c_525_n N_VPWR_c_936_n 0.00857714f $X=10.08 $Y=1.765 $X2=0
+ $Y2=0
cc_483 N_A_384_74#_c_526_n N_VPWR_c_936_n 0.00857685f $X=10.53 $Y=1.765 $X2=0
+ $Y2=0
cc_484 N_A_384_74#_c_527_n N_VPWR_c_936_n 0.00908635f $X=10.99 $Y=1.765 $X2=0
+ $Y2=0
cc_485 N_A_384_74#_c_528_n N_VPWR_c_936_n 0.00861505f $X=11.48 $Y=1.765 $X2=0
+ $Y2=0
cc_486 N_A_384_74#_c_529_n N_VPWR_c_936_n 0.0120466f $X=2.105 $Y=1.985 $X2=0
+ $Y2=0
cc_487 N_A_384_74#_c_532_n N_VPWR_c_936_n 0.0119791f $X=3.005 $Y=1.985 $X2=0
+ $Y2=0
cc_488 N_A_384_74#_c_535_n N_VPWR_c_936_n 0.0119791f $X=3.905 $Y=1.985 $X2=0
+ $Y2=0
cc_489 N_A_384_74#_M1003_g N_Y_c_1159_n 0.0138189f $X=4.565 $Y=0.74 $X2=0 $Y2=0
cc_490 N_A_384_74#_c_513_n N_Y_c_1159_n 0.00349092f $X=4.58 $Y=1.765 $X2=0 $Y2=0
cc_491 N_A_384_74#_M1006_g N_Y_c_1159_n 0.00296452f $X=4.995 $Y=0.74 $X2=0 $Y2=0
cc_492 N_A_384_74#_c_514_n N_Y_c_1159_n 0.0016226f $X=5.03 $Y=1.765 $X2=0 $Y2=0
cc_493 N_A_384_74#_c_502_n N_Y_c_1159_n 0.0375164f $X=3.905 $Y=1.97 $X2=0 $Y2=0
cc_494 N_A_384_74#_c_504_n N_Y_c_1159_n 0.0303937f $X=10.71 $Y=1.665 $X2=0 $Y2=0
cc_495 N_A_384_74#_c_505_n N_Y_c_1159_n 0.0314892f $X=5.175 $Y=1.465 $X2=0 $Y2=0
cc_496 N_A_384_74#_c_512_n N_Y_c_1159_n 0.0252626f $X=11.435 $Y=1.532 $X2=0
+ $Y2=0
cc_497 N_A_384_74#_c_514_n N_Y_c_1160_n 5.01468e-19 $X=5.03 $Y=1.765 $X2=0 $Y2=0
cc_498 N_A_384_74#_M1012_g N_Y_c_1160_n 0.00318673f $X=5.425 $Y=0.74 $X2=0 $Y2=0
cc_499 N_A_384_74#_c_515_n N_Y_c_1160_n 0.00371382f $X=5.48 $Y=1.765 $X2=0 $Y2=0
cc_500 N_A_384_74#_M1018_g N_Y_c_1160_n 0.00511263f $X=5.855 $Y=0.74 $X2=0 $Y2=0
cc_501 N_A_384_74#_c_516_n N_Y_c_1160_n 0.00315768f $X=5.93 $Y=1.765 $X2=0 $Y2=0
cc_502 N_A_384_74#_c_504_n N_Y_c_1160_n 0.0260421f $X=10.71 $Y=1.665 $X2=0 $Y2=0
cc_503 N_A_384_74#_c_505_n N_Y_c_1160_n 0.0263634f $X=5.175 $Y=1.465 $X2=0 $Y2=0
cc_504 N_A_384_74#_c_506_n N_Y_c_1160_n 0.0307253f $X=6.065 $Y=1.465 $X2=0 $Y2=0
cc_505 N_A_384_74#_c_512_n N_Y_c_1160_n 0.0255828f $X=11.435 $Y=1.532 $X2=0
+ $Y2=0
cc_506 N_A_384_74#_M1018_g N_Y_c_1161_n 0.00109749f $X=5.855 $Y=0.74 $X2=0 $Y2=0
cc_507 N_A_384_74#_c_516_n N_Y_c_1161_n 8.03241e-19 $X=5.93 $Y=1.765 $X2=0 $Y2=0
cc_508 N_A_384_74#_M1020_g N_Y_c_1161_n 0.0131322f $X=6.355 $Y=0.74 $X2=0 $Y2=0
cc_509 N_A_384_74#_c_517_n N_Y_c_1161_n 0.00357057f $X=6.38 $Y=1.765 $X2=0 $Y2=0
cc_510 N_A_384_74#_M1021_g N_Y_c_1161_n 0.00519497f $X=6.785 $Y=0.74 $X2=0 $Y2=0
cc_511 N_A_384_74#_c_518_n N_Y_c_1161_n 0.00333565f $X=6.83 $Y=1.765 $X2=0 $Y2=0
cc_512 N_A_384_74#_c_504_n N_Y_c_1161_n 0.0280018f $X=10.71 $Y=1.665 $X2=0 $Y2=0
cc_513 N_A_384_74#_c_506_n N_Y_c_1161_n 0.028655f $X=6.065 $Y=1.465 $X2=0 $Y2=0
cc_514 N_A_384_74#_c_507_n N_Y_c_1161_n 0.0293279f $X=7.005 $Y=1.465 $X2=0 $Y2=0
cc_515 N_A_384_74#_c_512_n N_Y_c_1161_n 0.0271425f $X=11.435 $Y=1.532 $X2=0
+ $Y2=0
cc_516 N_A_384_74#_M1021_g N_Y_c_1162_n 0.00110789f $X=6.785 $Y=0.74 $X2=0 $Y2=0
cc_517 N_A_384_74#_c_518_n N_Y_c_1162_n 0.0011223f $X=6.83 $Y=1.765 $X2=0 $Y2=0
cc_518 N_A_384_74#_c_519_n N_Y_c_1162_n 0.00339593f $X=7.28 $Y=1.765 $X2=0 $Y2=0
cc_519 N_A_384_74#_M1025_g N_Y_c_1162_n 0.0137331f $X=7.285 $Y=0.74 $X2=0 $Y2=0
cc_520 N_A_384_74#_M1027_g N_Y_c_1162_n 0.0052341f $X=7.715 $Y=0.74 $X2=0 $Y2=0
cc_521 N_A_384_74#_c_520_n N_Y_c_1162_n 0.00349095f $X=7.73 $Y=1.765 $X2=0 $Y2=0
cc_522 N_A_384_74#_c_504_n N_Y_c_1162_n 0.0286501f $X=10.71 $Y=1.665 $X2=0 $Y2=0
cc_523 N_A_384_74#_c_507_n N_Y_c_1162_n 0.0317837f $X=7.005 $Y=1.465 $X2=0 $Y2=0
cc_524 N_A_384_74#_c_508_n N_Y_c_1162_n 0.0309189f $X=7.925 $Y=1.465 $X2=0 $Y2=0
cc_525 N_A_384_74#_c_512_n N_Y_c_1162_n 0.0277215f $X=11.435 $Y=1.532 $X2=0
+ $Y2=0
cc_526 N_A_384_74#_c_519_n N_Y_c_1171_n 0.00961693f $X=7.28 $Y=1.765 $X2=0 $Y2=0
cc_527 N_A_384_74#_c_520_n N_Y_c_1171_n 0.00961693f $X=7.73 $Y=1.765 $X2=0 $Y2=0
cc_528 N_A_384_74#_c_521_n N_Y_c_1226_n 0.00163606f $X=8.18 $Y=1.765 $X2=0 $Y2=0
cc_529 N_A_384_74#_c_522_n N_Y_c_1226_n 0.00231761f $X=8.63 $Y=1.765 $X2=0 $Y2=0
cc_530 N_A_384_74#_c_504_n N_Y_c_1226_n 8.5796e-19 $X=10.71 $Y=1.665 $X2=0 $Y2=0
cc_531 N_A_384_74#_c_512_n N_Y_c_1226_n 0.0011003f $X=11.435 $Y=1.532 $X2=0
+ $Y2=0
cc_532 N_A_384_74#_c_521_n N_Y_c_1172_n 0.00899891f $X=8.18 $Y=1.765 $X2=0 $Y2=0
cc_533 N_A_384_74#_c_522_n N_Y_c_1172_n 0.00907095f $X=8.63 $Y=1.765 $X2=0 $Y2=0
cc_534 N_A_384_74#_M1027_g N_Y_c_1163_n 0.00111312f $X=7.715 $Y=0.74 $X2=0 $Y2=0
cc_535 N_A_384_74#_c_521_n N_Y_c_1163_n 0.00197231f $X=8.18 $Y=1.765 $X2=0 $Y2=0
cc_536 N_A_384_74#_M1028_g N_Y_c_1163_n 0.0140323f $X=8.215 $Y=0.74 $X2=0 $Y2=0
cc_537 N_A_384_74#_c_522_n N_Y_c_1163_n 0.00189142f $X=8.63 $Y=1.765 $X2=0 $Y2=0
cc_538 N_A_384_74#_M1031_g N_Y_c_1163_n 0.0052532f $X=8.645 $Y=0.74 $X2=0 $Y2=0
cc_539 N_A_384_74#_c_504_n N_Y_c_1163_n 0.0292669f $X=10.71 $Y=1.665 $X2=0 $Y2=0
cc_540 N_A_384_74#_c_508_n N_Y_c_1163_n 0.0309769f $X=7.925 $Y=1.465 $X2=0 $Y2=0
cc_541 N_A_384_74#_c_509_n N_Y_c_1163_n 0.0317841f $X=8.85 $Y=1.465 $X2=0 $Y2=0
cc_542 N_A_384_74#_c_512_n N_Y_c_1163_n 0.0281939f $X=11.435 $Y=1.532 $X2=0
+ $Y2=0
cc_543 N_A_384_74#_c_523_n N_Y_c_1241_n 0.00205728f $X=9.13 $Y=1.765 $X2=0 $Y2=0
cc_544 N_A_384_74#_c_524_n N_Y_c_1241_n 0.00231761f $X=9.58 $Y=1.765 $X2=0 $Y2=0
cc_545 N_A_384_74#_c_504_n N_Y_c_1241_n 8.08016e-19 $X=10.71 $Y=1.665 $X2=0
+ $Y2=0
cc_546 N_A_384_74#_c_512_n N_Y_c_1241_n 0.00129895f $X=11.435 $Y=1.532 $X2=0
+ $Y2=0
cc_547 N_A_384_74#_c_523_n N_Y_c_1174_n 0.00897724f $X=9.13 $Y=1.765 $X2=0 $Y2=0
cc_548 N_A_384_74#_c_524_n N_Y_c_1174_n 0.00907095f $X=9.58 $Y=1.765 $X2=0 $Y2=0
cc_549 N_A_384_74#_c_522_n N_Y_c_1164_n 6.77785e-19 $X=8.63 $Y=1.765 $X2=0 $Y2=0
cc_550 N_A_384_74#_M1031_g N_Y_c_1164_n 0.00111312f $X=8.645 $Y=0.74 $X2=0 $Y2=0
cc_551 N_A_384_74#_c_523_n N_Y_c_1164_n 0.00345862f $X=9.13 $Y=1.765 $X2=0 $Y2=0
cc_552 N_A_384_74#_M1033_g N_Y_c_1164_n 0.0140323f $X=9.145 $Y=0.74 $X2=0 $Y2=0
cc_553 N_A_384_74#_M1034_g N_Y_c_1164_n 0.0052532f $X=9.575 $Y=0.74 $X2=0 $Y2=0
cc_554 N_A_384_74#_c_524_n N_Y_c_1164_n 0.00354903f $X=9.58 $Y=1.765 $X2=0 $Y2=0
cc_555 N_A_384_74#_c_504_n N_Y_c_1164_n 0.0291792f $X=10.71 $Y=1.665 $X2=0 $Y2=0
cc_556 N_A_384_74#_c_509_n N_Y_c_1164_n 0.0301883f $X=8.85 $Y=1.465 $X2=0 $Y2=0
cc_557 N_A_384_74#_c_510_n N_Y_c_1164_n 0.0317841f $X=9.78 $Y=1.465 $X2=0 $Y2=0
cc_558 N_A_384_74#_c_512_n N_Y_c_1164_n 0.0282137f $X=11.435 $Y=1.532 $X2=0
+ $Y2=0
cc_559 N_A_384_74#_M1034_g N_Y_c_1165_n 0.00111312f $X=9.575 $Y=0.74 $X2=0 $Y2=0
cc_560 N_A_384_74#_c_524_n N_Y_c_1165_n 7.57715e-19 $X=9.58 $Y=1.765 $X2=0 $Y2=0
cc_561 N_A_384_74#_M1035_g N_Y_c_1165_n 0.0140323f $X=10.075 $Y=0.74 $X2=0 $Y2=0
cc_562 N_A_384_74#_c_525_n N_Y_c_1165_n 0.00365835f $X=10.08 $Y=1.765 $X2=0
+ $Y2=0
cc_563 N_A_384_74#_M1036_g N_Y_c_1165_n 0.0052532f $X=10.505 $Y=0.74 $X2=0 $Y2=0
cc_564 N_A_384_74#_c_526_n N_Y_c_1165_n 0.00346205f $X=10.53 $Y=1.765 $X2=0
+ $Y2=0
cc_565 N_A_384_74#_c_504_n N_Y_c_1165_n 0.0291297f $X=10.71 $Y=1.665 $X2=0 $Y2=0
cc_566 N_A_384_74#_c_510_n N_Y_c_1165_n 0.0301883f $X=9.78 $Y=1.465 $X2=0 $Y2=0
cc_567 N_A_384_74#_c_511_n N_Y_c_1165_n 0.0317841f $X=10.71 $Y=1.465 $X2=0 $Y2=0
cc_568 N_A_384_74#_c_512_n N_Y_c_1165_n 0.0277872f $X=11.435 $Y=1.532 $X2=0
+ $Y2=0
cc_569 N_A_384_74#_M1036_g N_Y_c_1166_n 0.00110862f $X=10.505 $Y=0.74 $X2=0
+ $Y2=0
cc_570 N_A_384_74#_c_526_n N_Y_c_1166_n 7.00472e-19 $X=10.53 $Y=1.765 $X2=0
+ $Y2=0
cc_571 N_A_384_74#_c_527_n N_Y_c_1166_n 5.13991e-19 $X=10.99 $Y=1.765 $X2=0
+ $Y2=0
cc_572 N_A_384_74#_M1038_g N_Y_c_1166_n 0.01491f $X=11.005 $Y=0.74 $X2=0 $Y2=0
cc_573 N_A_384_74#_M1042_g N_Y_c_1166_n 0.0190845f $X=11.435 $Y=0.74 $X2=0 $Y2=0
cc_574 N_A_384_74#_c_528_n N_Y_c_1166_n 6.99718e-19 $X=11.48 $Y=1.765 $X2=0
+ $Y2=0
cc_575 N_A_384_74#_c_504_n N_Y_c_1166_n 0.00286257f $X=10.71 $Y=1.665 $X2=0
+ $Y2=0
cc_576 N_A_384_74#_c_511_n N_Y_c_1166_n 0.0313503f $X=10.71 $Y=1.465 $X2=0 $Y2=0
cc_577 N_A_384_74#_c_512_n N_Y_c_1166_n 0.0461404f $X=11.435 $Y=1.532 $X2=0
+ $Y2=0
cc_578 N_A_384_74#_c_513_n N_Y_c_1276_n 0.00237354f $X=4.58 $Y=1.765 $X2=0 $Y2=0
cc_579 N_A_384_74#_c_514_n N_Y_c_1276_n 9.83579e-19 $X=5.03 $Y=1.765 $X2=0 $Y2=0
cc_580 N_A_384_74#_c_504_n N_Y_c_1276_n 9.42848e-19 $X=10.71 $Y=1.665 $X2=0
+ $Y2=0
cc_581 N_A_384_74#_c_512_n N_Y_c_1276_n 0.0020928f $X=11.435 $Y=1.532 $X2=0
+ $Y2=0
cc_582 N_A_384_74#_c_515_n N_Y_c_1280_n 0.00150203f $X=5.48 $Y=1.765 $X2=0 $Y2=0
cc_583 N_A_384_74#_c_516_n N_Y_c_1280_n 9.83579e-19 $X=5.93 $Y=1.765 $X2=0 $Y2=0
cc_584 N_A_384_74#_c_504_n N_Y_c_1280_n 0.00125217f $X=10.71 $Y=1.665 $X2=0
+ $Y2=0
cc_585 N_A_384_74#_c_512_n N_Y_c_1280_n 0.00315126f $X=11.435 $Y=1.532 $X2=0
+ $Y2=0
cc_586 N_A_384_74#_c_517_n N_Y_c_1284_n 0.0012181f $X=6.38 $Y=1.765 $X2=0 $Y2=0
cc_587 N_A_384_74#_c_518_n N_Y_c_1284_n 9.83579e-19 $X=6.83 $Y=1.765 $X2=0 $Y2=0
cc_588 N_A_384_74#_c_504_n N_Y_c_1284_n 0.00102018f $X=10.71 $Y=1.665 $X2=0
+ $Y2=0
cc_589 N_A_384_74#_c_512_n N_Y_c_1284_n 0.00235741f $X=11.435 $Y=1.532 $X2=0
+ $Y2=0
cc_590 N_A_384_74#_c_525_n N_Y_c_1288_n 0.0010526f $X=10.08 $Y=1.765 $X2=0 $Y2=0
cc_591 N_A_384_74#_c_526_n N_Y_c_1288_n 9.83579e-19 $X=10.53 $Y=1.765 $X2=0
+ $Y2=0
cc_592 N_A_384_74#_c_504_n N_Y_c_1288_n 8.65518e-19 $X=10.71 $Y=1.665 $X2=0
+ $Y2=0
cc_593 N_A_384_74#_c_512_n N_Y_c_1288_n 0.00182818f $X=11.435 $Y=1.532 $X2=0
+ $Y2=0
cc_594 N_A_384_74#_c_527_n N_Y_c_1178_n 0.0037886f $X=10.99 $Y=1.765 $X2=0 $Y2=0
cc_595 N_A_384_74#_c_528_n N_Y_c_1178_n 0.00485542f $X=11.48 $Y=1.765 $X2=0
+ $Y2=0
cc_596 N_A_384_74#_c_512_n N_Y_c_1178_n 0.00109503f $X=11.435 $Y=1.532 $X2=0
+ $Y2=0
cc_597 N_A_384_74#_c_513_n N_Y_c_1179_n 0.0104948f $X=4.58 $Y=1.765 $X2=0 $Y2=0
cc_598 N_A_384_74#_c_514_n N_Y_c_1179_n 0.0100549f $X=5.03 $Y=1.765 $X2=0 $Y2=0
cc_599 N_A_384_74#_c_515_n N_Y_c_1180_n 0.0100549f $X=5.48 $Y=1.765 $X2=0 $Y2=0
cc_600 N_A_384_74#_c_516_n N_Y_c_1180_n 0.0100549f $X=5.93 $Y=1.765 $X2=0 $Y2=0
cc_601 N_A_384_74#_c_517_n N_Y_c_1181_n 0.0100549f $X=6.38 $Y=1.765 $X2=0 $Y2=0
cc_602 N_A_384_74#_c_518_n N_Y_c_1181_n 0.0100549f $X=6.83 $Y=1.765 $X2=0 $Y2=0
cc_603 N_A_384_74#_c_525_n N_Y_c_1182_n 0.00980516f $X=10.08 $Y=1.765 $X2=0
+ $Y2=0
cc_604 N_A_384_74#_c_526_n N_Y_c_1182_n 0.0100706f $X=10.53 $Y=1.765 $X2=0 $Y2=0
cc_605 N_A_384_74#_c_527_n N_Y_c_1183_n 6.61845e-19 $X=10.99 $Y=1.765 $X2=0
+ $Y2=0
cc_606 N_A_384_74#_c_528_n N_Y_c_1183_n 0.0112715f $X=11.48 $Y=1.765 $X2=0 $Y2=0
cc_607 N_A_384_74#_c_514_n N_Y_c_1305_n 0.00689819f $X=5.03 $Y=1.765 $X2=0 $Y2=0
cc_608 N_A_384_74#_c_515_n N_Y_c_1305_n 0.0067316f $X=5.48 $Y=1.765 $X2=0 $Y2=0
cc_609 N_A_384_74#_c_516_n N_Y_c_1305_n 0.00677868f $X=5.93 $Y=1.765 $X2=0 $Y2=0
cc_610 N_A_384_74#_c_517_n N_Y_c_1305_n 0.00681955f $X=6.38 $Y=1.765 $X2=0 $Y2=0
cc_611 N_A_384_74#_c_518_n N_Y_c_1305_n 0.00691526f $X=6.83 $Y=1.765 $X2=0 $Y2=0
cc_612 N_A_384_74#_c_519_n N_Y_c_1305_n 0.00701605f $X=7.28 $Y=1.765 $X2=0 $Y2=0
cc_613 N_A_384_74#_c_520_n N_Y_c_1305_n 0.00698355f $X=7.73 $Y=1.765 $X2=0 $Y2=0
cc_614 N_A_384_74#_c_521_n N_Y_c_1305_n 0.00706675f $X=8.18 $Y=1.765 $X2=0 $Y2=0
cc_615 N_A_384_74#_c_522_n N_Y_c_1305_n 0.00700528f $X=8.63 $Y=1.765 $X2=0 $Y2=0
cc_616 N_A_384_74#_c_523_n N_Y_c_1305_n 0.00874967f $X=9.13 $Y=1.765 $X2=0 $Y2=0
cc_617 N_A_384_74#_c_524_n N_Y_c_1305_n 0.00693699f $X=9.58 $Y=1.765 $X2=0 $Y2=0
cc_618 N_A_384_74#_c_525_n N_Y_c_1305_n 0.0086256f $X=10.08 $Y=1.765 $X2=0 $Y2=0
cc_619 N_A_384_74#_c_526_n N_Y_c_1305_n 0.00693233f $X=10.53 $Y=1.765 $X2=0
+ $Y2=0
cc_620 N_A_384_74#_c_527_n N_Y_c_1305_n 0.0123908f $X=10.99 $Y=1.765 $X2=0 $Y2=0
cc_621 N_A_384_74#_c_504_n N_Y_c_1305_n 0.607041f $X=10.71 $Y=1.665 $X2=0 $Y2=0
cc_622 N_A_384_74#_c_505_n N_Y_c_1305_n 0.00188824f $X=5.175 $Y=1.465 $X2=0
+ $Y2=0
cc_623 N_A_384_74#_c_506_n N_Y_c_1305_n 0.00249084f $X=6.065 $Y=1.465 $X2=0
+ $Y2=0
cc_624 N_A_384_74#_c_507_n N_Y_c_1305_n 0.00205675f $X=7.005 $Y=1.465 $X2=0
+ $Y2=0
cc_625 N_A_384_74#_c_508_n N_Y_c_1305_n 0.00186995f $X=7.925 $Y=1.465 $X2=0
+ $Y2=0
cc_626 N_A_384_74#_c_509_n N_Y_c_1305_n 0.00130386f $X=8.85 $Y=1.465 $X2=0 $Y2=0
cc_627 N_A_384_74#_c_510_n N_Y_c_1305_n 0.00149067f $X=9.78 $Y=1.465 $X2=0 $Y2=0
cc_628 N_A_384_74#_c_511_n N_Y_c_1305_n 0.00193542f $X=10.71 $Y=1.465 $X2=0
+ $Y2=0
cc_629 N_A_384_74#_c_512_n N_Y_c_1305_n 0.00285123f $X=11.435 $Y=1.532 $X2=0
+ $Y2=0
cc_630 N_A_384_74#_c_519_n N_Y_c_1328_n 0.00111176f $X=7.28 $Y=1.765 $X2=0 $Y2=0
cc_631 N_A_384_74#_c_520_n N_Y_c_1328_n 0.00142154f $X=7.73 $Y=1.765 $X2=0 $Y2=0
cc_632 N_A_384_74#_c_504_n N_Y_c_1328_n 7.88189e-19 $X=10.71 $Y=1.665 $X2=0
+ $Y2=0
cc_633 N_A_384_74#_c_512_n N_Y_c_1328_n 0.00156357f $X=11.435 $Y=1.532 $X2=0
+ $Y2=0
cc_634 N_A_384_74#_c_497_n N_VGND_M1014_s 0.00176461f $X=2.755 $Y=1.045 $X2=0
+ $Y2=0
cc_635 N_A_384_74#_c_500_n N_VGND_M1024_s 0.00250873f $X=3.685 $Y=1.045 $X2=0
+ $Y2=0
cc_636 N_A_384_74#_c_496_n N_VGND_c_1422_n 0.0182488f $X=2.06 $Y=0.515 $X2=0
+ $Y2=0
cc_637 N_A_384_74#_c_496_n N_VGND_c_1423_n 0.0157999f $X=2.06 $Y=0.515 $X2=0
+ $Y2=0
cc_638 N_A_384_74#_c_497_n N_VGND_c_1423_n 0.0152916f $X=2.755 $Y=1.045 $X2=0
+ $Y2=0
cc_639 N_A_384_74#_c_499_n N_VGND_c_1423_n 0.0158413f $X=2.92 $Y=0.515 $X2=0
+ $Y2=0
cc_640 N_A_384_74#_c_499_n N_VGND_c_1424_n 0.0164981f $X=2.92 $Y=0.515 $X2=0
+ $Y2=0
cc_641 N_A_384_74#_c_500_n N_VGND_c_1424_n 0.0209867f $X=3.685 $Y=1.045 $X2=0
+ $Y2=0
cc_642 N_A_384_74#_c_501_n N_VGND_c_1424_n 0.0166127f $X=3.85 $Y=0.515 $X2=0
+ $Y2=0
cc_643 N_A_384_74#_M1003_g N_VGND_c_1425_n 0.00581358f $X=4.565 $Y=0.74 $X2=0
+ $Y2=0
cc_644 N_A_384_74#_c_501_n N_VGND_c_1425_n 0.0225912f $X=3.85 $Y=0.515 $X2=0
+ $Y2=0
cc_645 N_A_384_74#_c_502_n N_VGND_c_1425_n 0.0342051f $X=3.905 $Y=1.97 $X2=0
+ $Y2=0
cc_646 N_A_384_74#_c_504_n N_VGND_c_1425_n 0.00177399f $X=10.71 $Y=1.665 $X2=0
+ $Y2=0
cc_647 N_A_384_74#_M1003_g N_VGND_c_1426_n 5.98876e-19 $X=4.565 $Y=0.74 $X2=0
+ $Y2=0
cc_648 N_A_384_74#_M1006_g N_VGND_c_1426_n 0.0121668f $X=4.995 $Y=0.74 $X2=0
+ $Y2=0
cc_649 N_A_384_74#_M1012_g N_VGND_c_1426_n 0.00174374f $X=5.425 $Y=0.74 $X2=0
+ $Y2=0
cc_650 N_A_384_74#_c_504_n N_VGND_c_1426_n 0.00123706f $X=10.71 $Y=1.665 $X2=0
+ $Y2=0
cc_651 N_A_384_74#_c_505_n N_VGND_c_1426_n 0.0155643f $X=5.175 $Y=1.465 $X2=0
+ $Y2=0
cc_652 N_A_384_74#_c_512_n N_VGND_c_1426_n 7.77773e-19 $X=11.435 $Y=1.532 $X2=0
+ $Y2=0
cc_653 N_A_384_74#_M1012_g N_VGND_c_1427_n 5.61948e-19 $X=5.425 $Y=0.74 $X2=0
+ $Y2=0
cc_654 N_A_384_74#_M1018_g N_VGND_c_1427_n 0.0126669f $X=5.855 $Y=0.74 $X2=0
+ $Y2=0
cc_655 N_A_384_74#_M1020_g N_VGND_c_1427_n 0.00562547f $X=6.355 $Y=0.74 $X2=0
+ $Y2=0
cc_656 N_A_384_74#_c_504_n N_VGND_c_1427_n 0.00181192f $X=10.71 $Y=1.665 $X2=0
+ $Y2=0
cc_657 N_A_384_74#_c_506_n N_VGND_c_1427_n 0.0207506f $X=6.065 $Y=1.465 $X2=0
+ $Y2=0
cc_658 N_A_384_74#_c_512_n N_VGND_c_1427_n 0.00132221f $X=11.435 $Y=1.532 $X2=0
+ $Y2=0
cc_659 N_A_384_74#_M1020_g N_VGND_c_1428_n 5.96902e-19 $X=6.355 $Y=0.74 $X2=0
+ $Y2=0
cc_660 N_A_384_74#_M1021_g N_VGND_c_1428_n 0.0126964f $X=6.785 $Y=0.74 $X2=0
+ $Y2=0
cc_661 N_A_384_74#_M1025_g N_VGND_c_1428_n 0.00562212f $X=7.285 $Y=0.74 $X2=0
+ $Y2=0
cc_662 N_A_384_74#_c_504_n N_VGND_c_1428_n 0.00179414f $X=10.71 $Y=1.665 $X2=0
+ $Y2=0
cc_663 N_A_384_74#_c_507_n N_VGND_c_1428_n 0.020583f $X=7.005 $Y=1.465 $X2=0
+ $Y2=0
cc_664 N_A_384_74#_c_512_n N_VGND_c_1428_n 0.00132221f $X=11.435 $Y=1.532 $X2=0
+ $Y2=0
cc_665 N_A_384_74#_M1025_g N_VGND_c_1429_n 5.96902e-19 $X=7.285 $Y=0.74 $X2=0
+ $Y2=0
cc_666 N_A_384_74#_M1027_g N_VGND_c_1429_n 0.0126506f $X=7.715 $Y=0.74 $X2=0
+ $Y2=0
cc_667 N_A_384_74#_M1028_g N_VGND_c_1429_n 0.00562044f $X=8.215 $Y=0.74 $X2=0
+ $Y2=0
cc_668 N_A_384_74#_c_504_n N_VGND_c_1429_n 0.00181192f $X=10.71 $Y=1.665 $X2=0
+ $Y2=0
cc_669 N_A_384_74#_c_508_n N_VGND_c_1429_n 0.0207506f $X=7.925 $Y=1.465 $X2=0
+ $Y2=0
cc_670 N_A_384_74#_c_512_n N_VGND_c_1429_n 0.00132221f $X=11.435 $Y=1.532 $X2=0
+ $Y2=0
cc_671 N_A_384_74#_M1028_g N_VGND_c_1430_n 5.96902e-19 $X=8.215 $Y=0.74 $X2=0
+ $Y2=0
cc_672 N_A_384_74#_M1031_g N_VGND_c_1430_n 0.0126506f $X=8.645 $Y=0.74 $X2=0
+ $Y2=0
cc_673 N_A_384_74#_M1033_g N_VGND_c_1430_n 0.00562044f $X=9.145 $Y=0.74 $X2=0
+ $Y2=0
cc_674 N_A_384_74#_c_504_n N_VGND_c_1430_n 0.00197911f $X=10.71 $Y=1.665 $X2=0
+ $Y2=0
cc_675 N_A_384_74#_c_509_n N_VGND_c_1430_n 0.0205727f $X=8.85 $Y=1.465 $X2=0
+ $Y2=0
cc_676 N_A_384_74#_c_512_n N_VGND_c_1430_n 0.00132221f $X=11.435 $Y=1.532 $X2=0
+ $Y2=0
cc_677 N_A_384_74#_M1033_g N_VGND_c_1431_n 5.96902e-19 $X=9.145 $Y=0.74 $X2=0
+ $Y2=0
cc_678 N_A_384_74#_M1034_g N_VGND_c_1431_n 0.0126506f $X=9.575 $Y=0.74 $X2=0
+ $Y2=0
cc_679 N_A_384_74#_M1035_g N_VGND_c_1431_n 0.00562044f $X=10.075 $Y=0.74 $X2=0
+ $Y2=0
cc_680 N_A_384_74#_c_504_n N_VGND_c_1431_n 0.00197911f $X=10.71 $Y=1.665 $X2=0
+ $Y2=0
cc_681 N_A_384_74#_c_510_n N_VGND_c_1431_n 0.0205727f $X=9.78 $Y=1.465 $X2=0
+ $Y2=0
cc_682 N_A_384_74#_c_512_n N_VGND_c_1431_n 0.00132221f $X=11.435 $Y=1.532 $X2=0
+ $Y2=0
cc_683 N_A_384_74#_M1035_g N_VGND_c_1432_n 5.96902e-19 $X=10.075 $Y=0.74 $X2=0
+ $Y2=0
cc_684 N_A_384_74#_M1036_g N_VGND_c_1432_n 0.0126506f $X=10.505 $Y=0.74 $X2=0
+ $Y2=0
cc_685 N_A_384_74#_M1038_g N_VGND_c_1432_n 0.00570988f $X=11.005 $Y=0.74 $X2=0
+ $Y2=0
cc_686 N_A_384_74#_c_504_n N_VGND_c_1432_n 0.00149791f $X=10.71 $Y=1.665 $X2=0
+ $Y2=0
cc_687 N_A_384_74#_c_511_n N_VGND_c_1432_n 0.0206571f $X=10.71 $Y=1.465 $X2=0
+ $Y2=0
cc_688 N_A_384_74#_c_512_n N_VGND_c_1432_n 0.00132221f $X=11.435 $Y=1.532 $X2=0
+ $Y2=0
cc_689 N_A_384_74#_M1042_g N_VGND_c_1434_n 0.0184907f $X=11.435 $Y=0.74 $X2=0
+ $Y2=0
cc_690 N_A_384_74#_c_512_n N_VGND_c_1434_n 6.45246e-19 $X=11.435 $Y=1.532 $X2=0
+ $Y2=0
cc_691 N_A_384_74#_c_496_n N_VGND_c_1435_n 0.00749631f $X=2.06 $Y=0.515 $X2=0
+ $Y2=0
cc_692 N_A_384_74#_c_499_n N_VGND_c_1437_n 0.0109942f $X=2.92 $Y=0.515 $X2=0
+ $Y2=0
cc_693 N_A_384_74#_c_501_n N_VGND_c_1439_n 0.0109942f $X=3.85 $Y=0.515 $X2=0
+ $Y2=0
cc_694 N_A_384_74#_M1003_g N_VGND_c_1441_n 0.00434272f $X=4.565 $Y=0.74 $X2=0
+ $Y2=0
cc_695 N_A_384_74#_M1006_g N_VGND_c_1441_n 0.00383152f $X=4.995 $Y=0.74 $X2=0
+ $Y2=0
cc_696 N_A_384_74#_M1012_g N_VGND_c_1445_n 0.00461464f $X=5.425 $Y=0.74 $X2=0
+ $Y2=0
cc_697 N_A_384_74#_M1018_g N_VGND_c_1445_n 0.00383152f $X=5.855 $Y=0.74 $X2=0
+ $Y2=0
cc_698 N_A_384_74#_M1020_g N_VGND_c_1446_n 0.00451267f $X=6.355 $Y=0.74 $X2=0
+ $Y2=0
cc_699 N_A_384_74#_M1021_g N_VGND_c_1446_n 0.00383152f $X=6.785 $Y=0.74 $X2=0
+ $Y2=0
cc_700 N_A_384_74#_M1025_g N_VGND_c_1447_n 0.00439937f $X=7.285 $Y=0.74 $X2=0
+ $Y2=0
cc_701 N_A_384_74#_M1027_g N_VGND_c_1447_n 0.00383152f $X=7.715 $Y=0.74 $X2=0
+ $Y2=0
cc_702 N_A_384_74#_M1028_g N_VGND_c_1448_n 0.00434272f $X=8.215 $Y=0.74 $X2=0
+ $Y2=0
cc_703 N_A_384_74#_M1031_g N_VGND_c_1448_n 0.00383152f $X=8.645 $Y=0.74 $X2=0
+ $Y2=0
cc_704 N_A_384_74#_M1033_g N_VGND_c_1449_n 0.00434272f $X=9.145 $Y=0.74 $X2=0
+ $Y2=0
cc_705 N_A_384_74#_M1034_g N_VGND_c_1449_n 0.00383152f $X=9.575 $Y=0.74 $X2=0
+ $Y2=0
cc_706 N_A_384_74#_M1035_g N_VGND_c_1450_n 0.00434272f $X=10.075 $Y=0.74 $X2=0
+ $Y2=0
cc_707 N_A_384_74#_M1036_g N_VGND_c_1450_n 0.00383152f $X=10.505 $Y=0.74 $X2=0
+ $Y2=0
cc_708 N_A_384_74#_M1038_g N_VGND_c_1451_n 0.00434272f $X=11.005 $Y=0.74 $X2=0
+ $Y2=0
cc_709 N_A_384_74#_M1042_g N_VGND_c_1451_n 0.00434272f $X=11.435 $Y=0.74 $X2=0
+ $Y2=0
cc_710 N_A_384_74#_M1003_g N_VGND_c_1460_n 0.00820772f $X=4.565 $Y=0.74 $X2=0
+ $Y2=0
cc_711 N_A_384_74#_M1006_g N_VGND_c_1460_n 0.0075754f $X=4.995 $Y=0.74 $X2=0
+ $Y2=0
cc_712 N_A_384_74#_M1012_g N_VGND_c_1460_n 0.00908333f $X=5.425 $Y=0.74 $X2=0
+ $Y2=0
cc_713 N_A_384_74#_M1018_g N_VGND_c_1460_n 0.0075754f $X=5.855 $Y=0.74 $X2=0
+ $Y2=0
cc_714 N_A_384_74#_M1020_g N_VGND_c_1460_n 0.00875749f $X=6.355 $Y=0.74 $X2=0
+ $Y2=0
cc_715 N_A_384_74#_M1021_g N_VGND_c_1460_n 0.0075754f $X=6.785 $Y=0.74 $X2=0
+ $Y2=0
cc_716 N_A_384_74#_M1025_g N_VGND_c_1460_n 0.00839062f $X=7.285 $Y=0.74 $X2=0
+ $Y2=0
cc_717 N_A_384_74#_M1027_g N_VGND_c_1460_n 0.0075754f $X=7.715 $Y=0.74 $X2=0
+ $Y2=0
cc_718 N_A_384_74#_M1028_g N_VGND_c_1460_n 0.00820718f $X=8.215 $Y=0.74 $X2=0
+ $Y2=0
cc_719 N_A_384_74#_M1031_g N_VGND_c_1460_n 0.0075754f $X=8.645 $Y=0.74 $X2=0
+ $Y2=0
cc_720 N_A_384_74#_M1033_g N_VGND_c_1460_n 0.00820718f $X=9.145 $Y=0.74 $X2=0
+ $Y2=0
cc_721 N_A_384_74#_M1034_g N_VGND_c_1460_n 0.0075754f $X=9.575 $Y=0.74 $X2=0
+ $Y2=0
cc_722 N_A_384_74#_M1035_g N_VGND_c_1460_n 0.00820718f $X=10.075 $Y=0.74 $X2=0
+ $Y2=0
cc_723 N_A_384_74#_M1036_g N_VGND_c_1460_n 0.0075754f $X=10.505 $Y=0.74 $X2=0
+ $Y2=0
cc_724 N_A_384_74#_M1038_g N_VGND_c_1460_n 0.00820718f $X=11.005 $Y=0.74 $X2=0
+ $Y2=0
cc_725 N_A_384_74#_M1042_g N_VGND_c_1460_n 0.00823934f $X=11.435 $Y=0.74 $X2=0
+ $Y2=0
cc_726 N_A_384_74#_c_496_n N_VGND_c_1460_n 0.0062048f $X=2.06 $Y=0.515 $X2=0
+ $Y2=0
cc_727 N_A_384_74#_c_499_n N_VGND_c_1460_n 0.00904371f $X=2.92 $Y=0.515 $X2=0
+ $Y2=0
cc_728 N_A_384_74#_c_501_n N_VGND_c_1460_n 0.00904371f $X=3.85 $Y=0.515 $X2=0
+ $Y2=0
cc_729 N_VPWR_c_945_n N_Y_c_1171_n 0.014552f $X=7.87 $Y=3.33 $X2=0 $Y2=0
cc_730 N_VPWR_c_936_n N_Y_c_1171_n 0.0119791f $X=11.76 $Y=3.33 $X2=0 $Y2=0
cc_731 N_VPWR_c_946_n N_Y_c_1226_n 0.0136173f $X=7.955 $Y=2.085 $X2=0 $Y2=0
cc_732 N_VPWR_c_947_n N_Y_c_1226_n 0.0154019f $X=8.855 $Y=2.085 $X2=0 $Y2=0
cc_733 N_VPWR_c_946_n N_Y_c_1172_n 0.0517782f $X=7.955 $Y=2.085 $X2=0 $Y2=0
cc_734 N_VPWR_c_947_n N_Y_c_1172_n 0.0528776f $X=8.855 $Y=2.085 $X2=0 $Y2=0
cc_735 N_VPWR_c_966_n N_Y_c_1172_n 0.014552f $X=8.77 $Y=3.33 $X2=0 $Y2=0
cc_736 N_VPWR_c_936_n N_Y_c_1172_n 0.0119791f $X=11.76 $Y=3.33 $X2=0 $Y2=0
cc_737 N_VPWR_c_947_n N_Y_c_1241_n 0.0156527f $X=8.855 $Y=2.085 $X2=0 $Y2=0
cc_738 N_VPWR_c_948_n N_Y_c_1241_n 0.0154163f $X=9.805 $Y=2.085 $X2=0 $Y2=0
cc_739 N_VPWR_c_947_n N_Y_c_1174_n 0.0539156f $X=8.855 $Y=2.085 $X2=0 $Y2=0
cc_740 N_VPWR_c_948_n N_Y_c_1174_n 0.0530521f $X=9.805 $Y=2.085 $X2=0 $Y2=0
cc_741 N_VPWR_c_967_n N_Y_c_1174_n 0.014552f $X=9.72 $Y=3.33 $X2=0 $Y2=0
cc_742 N_VPWR_c_936_n N_Y_c_1174_n 0.0119791f $X=11.76 $Y=3.33 $X2=0 $Y2=0
cc_743 N_VPWR_c_941_n N_Y_c_1276_n 0.00662689f $X=4.355 $Y=2.085 $X2=0 $Y2=0
cc_744 N_VPWR_c_942_n N_Y_c_1276_n 0.0670269f $X=5.255 $Y=2.085 $X2=0 $Y2=0
cc_745 N_VPWR_c_942_n N_Y_c_1280_n 0.0067098f $X=5.255 $Y=2.085 $X2=0 $Y2=0
cc_746 N_VPWR_c_943_n N_Y_c_1280_n 0.0670272f $X=6.155 $Y=2.085 $X2=0 $Y2=0
cc_747 N_VPWR_c_943_n N_Y_c_1284_n 0.00630839f $X=6.155 $Y=2.085 $X2=0 $Y2=0
cc_748 N_VPWR_c_944_n N_Y_c_1284_n 0.0670266f $X=7.055 $Y=2.085 $X2=0 $Y2=0
cc_749 N_VPWR_c_948_n N_Y_c_1288_n 0.00504547f $X=9.805 $Y=2.085 $X2=0 $Y2=0
cc_750 N_VPWR_c_949_n N_Y_c_1288_n 0.0680133f $X=10.755 $Y=2.085 $X2=0 $Y2=0
cc_751 N_VPWR_c_949_n N_Y_c_1178_n 0.005042f $X=10.755 $Y=2.085 $X2=0 $Y2=0
cc_752 N_VPWR_c_951_n N_Y_c_1178_n 0.0761753f $X=11.705 $Y=1.985 $X2=0 $Y2=0
cc_753 N_VPWR_c_941_n N_Y_c_1179_n 0.0616015f $X=4.355 $Y=2.085 $X2=0 $Y2=0
cc_754 N_VPWR_c_960_n N_Y_c_1179_n 0.014552f $X=5.17 $Y=3.33 $X2=0 $Y2=0
cc_755 N_VPWR_c_936_n N_Y_c_1179_n 0.0119791f $X=11.76 $Y=3.33 $X2=0 $Y2=0
cc_756 N_VPWR_c_942_n N_Y_c_1180_n 0.0613898f $X=5.255 $Y=2.085 $X2=0 $Y2=0
cc_757 N_VPWR_c_962_n N_Y_c_1180_n 0.014552f $X=6.07 $Y=3.33 $X2=0 $Y2=0
cc_758 N_VPWR_c_936_n N_Y_c_1180_n 0.0119791f $X=11.76 $Y=3.33 $X2=0 $Y2=0
cc_759 N_VPWR_c_943_n N_Y_c_1181_n 0.0613898f $X=6.155 $Y=2.085 $X2=0 $Y2=0
cc_760 N_VPWR_c_964_n N_Y_c_1181_n 0.014552f $X=6.97 $Y=3.33 $X2=0 $Y2=0
cc_761 N_VPWR_c_936_n N_Y_c_1181_n 0.0119791f $X=11.76 $Y=3.33 $X2=0 $Y2=0
cc_762 N_VPWR_c_948_n N_Y_c_1182_n 0.0357709f $X=9.805 $Y=2.085 $X2=0 $Y2=0
cc_763 N_VPWR_c_968_n N_Y_c_1182_n 0.014552f $X=10.67 $Y=3.33 $X2=0 $Y2=0
cc_764 N_VPWR_c_936_n N_Y_c_1182_n 0.0119791f $X=11.76 $Y=3.33 $X2=0 $Y2=0
cc_765 N_VPWR_c_949_n N_Y_c_1183_n 0.00519414f $X=10.755 $Y=2.085 $X2=0 $Y2=0
cc_766 N_VPWR_c_969_n N_Y_c_1183_n 0.0145938f $X=11.62 $Y=3.33 $X2=0 $Y2=0
cc_767 N_VPWR_c_936_n N_Y_c_1183_n 0.0120466f $X=11.76 $Y=3.33 $X2=0 $Y2=0
cc_768 N_VPWR_M1005_d N_Y_c_1305_n 0.00673208f $X=5.105 $Y=1.84 $X2=0 $Y2=0
cc_769 N_VPWR_M1008_d N_Y_c_1305_n 0.00667036f $X=6.005 $Y=1.84 $X2=0 $Y2=0
cc_770 N_VPWR_M1013_d N_Y_c_1305_n 0.00657159f $X=6.905 $Y=1.84 $X2=0 $Y2=0
cc_771 N_VPWR_M1023_d N_Y_c_1305_n 0.00651537f $X=7.805 $Y=1.84 $X2=0 $Y2=0
cc_772 N_VPWR_M1032_d N_Y_c_1305_n 0.00664997f $X=8.705 $Y=1.84 $X2=0 $Y2=0
cc_773 N_VPWR_M1039_d N_Y_c_1305_n 0.00613882f $X=9.655 $Y=1.84 $X2=0 $Y2=0
cc_774 N_VPWR_M1041_d N_Y_c_1305_n 0.00526943f $X=10.605 $Y=1.84 $X2=0 $Y2=0
cc_775 N_VPWR_c_941_n N_Y_c_1305_n 0.00152375f $X=4.355 $Y=2.085 $X2=0 $Y2=0
cc_776 N_VPWR_c_942_n N_Y_c_1305_n 0.0186233f $X=5.255 $Y=2.085 $X2=0 $Y2=0
cc_777 N_VPWR_c_943_n N_Y_c_1305_n 0.0186737f $X=6.155 $Y=2.085 $X2=0 $Y2=0
cc_778 N_VPWR_c_944_n N_Y_c_1305_n 0.0187715f $X=7.055 $Y=2.085 $X2=0 $Y2=0
cc_779 N_VPWR_c_946_n N_Y_c_1305_n 0.0188771f $X=7.955 $Y=2.085 $X2=0 $Y2=0
cc_780 N_VPWR_c_947_n N_Y_c_1305_n 0.0232384f $X=8.855 $Y=2.085 $X2=0 $Y2=0
cc_781 N_VPWR_c_948_n N_Y_c_1305_n 0.0239812f $X=9.805 $Y=2.085 $X2=0 $Y2=0
cc_782 N_VPWR_c_949_n N_Y_c_1305_n 0.022642f $X=10.755 $Y=2.085 $X2=0 $Y2=0
cc_783 N_VPWR_c_951_n N_Y_c_1305_n 0.00161542f $X=11.705 $Y=1.985 $X2=0 $Y2=0
cc_784 N_VPWR_c_944_n N_Y_c_1328_n 0.0670252f $X=7.055 $Y=2.085 $X2=0 $Y2=0
cc_785 N_VPWR_c_946_n N_Y_c_1328_n 0.0670252f $X=7.955 $Y=2.085 $X2=0 $Y2=0
cc_786 N_Y_c_1159_n N_VGND_c_1425_n 0.0296294f $X=4.78 $Y=0.515 $X2=0 $Y2=0
cc_787 N_Y_c_1159_n N_VGND_c_1426_n 0.026661f $X=4.78 $Y=0.515 $X2=0 $Y2=0
cc_788 N_Y_c_1160_n N_VGND_c_1426_n 0.00127089f $X=5.64 $Y=0.515 $X2=0 $Y2=0
cc_789 N_Y_c_1160_n N_VGND_c_1427_n 0.0277717f $X=5.64 $Y=0.515 $X2=0 $Y2=0
cc_790 N_Y_c_1161_n N_VGND_c_1427_n 0.0258753f $X=6.57 $Y=0.515 $X2=0 $Y2=0
cc_791 N_Y_c_1161_n N_VGND_c_1428_n 0.0277814f $X=6.57 $Y=0.515 $X2=0 $Y2=0
cc_792 N_Y_c_1162_n N_VGND_c_1428_n 0.0272176f $X=7.5 $Y=0.515 $X2=0 $Y2=0
cc_793 N_Y_c_1162_n N_VGND_c_1429_n 0.0277859f $X=7.5 $Y=0.515 $X2=0 $Y2=0
cc_794 N_Y_c_1163_n N_VGND_c_1429_n 0.0279399f $X=8.43 $Y=0.515 $X2=0 $Y2=0
cc_795 N_Y_c_1163_n N_VGND_c_1430_n 0.0277882f $X=8.43 $Y=0.515 $X2=0 $Y2=0
cc_796 N_Y_c_1164_n N_VGND_c_1430_n 0.0279399f $X=9.36 $Y=0.515 $X2=0 $Y2=0
cc_797 N_Y_c_1164_n N_VGND_c_1431_n 0.0277882f $X=9.36 $Y=0.515 $X2=0 $Y2=0
cc_798 N_Y_c_1165_n N_VGND_c_1431_n 0.0279399f $X=10.29 $Y=0.515 $X2=0 $Y2=0
cc_799 N_Y_c_1165_n N_VGND_c_1432_n 0.0277882f $X=10.29 $Y=0.515 $X2=0 $Y2=0
cc_800 N_Y_c_1166_n N_VGND_c_1432_n 0.0291199f $X=11.22 $Y=0.515 $X2=0 $Y2=0
cc_801 N_Y_c_1166_n N_VGND_c_1434_n 0.0308485f $X=11.22 $Y=0.515 $X2=0 $Y2=0
cc_802 N_Y_c_1159_n N_VGND_c_1441_n 0.0109942f $X=4.78 $Y=0.515 $X2=0 $Y2=0
cc_803 N_Y_c_1160_n N_VGND_c_1445_n 0.00950426f $X=5.64 $Y=0.515 $X2=0 $Y2=0
cc_804 N_Y_c_1161_n N_VGND_c_1446_n 0.0103698f $X=6.57 $Y=0.515 $X2=0 $Y2=0
cc_805 N_Y_c_1162_n N_VGND_c_1447_n 0.0107861f $X=7.5 $Y=0.515 $X2=0 $Y2=0
cc_806 N_Y_c_1163_n N_VGND_c_1448_n 0.0109942f $X=8.43 $Y=0.515 $X2=0 $Y2=0
cc_807 N_Y_c_1164_n N_VGND_c_1449_n 0.0109942f $X=9.36 $Y=0.515 $X2=0 $Y2=0
cc_808 N_Y_c_1165_n N_VGND_c_1450_n 0.0109942f $X=10.29 $Y=0.515 $X2=0 $Y2=0
cc_809 N_Y_c_1166_n N_VGND_c_1451_n 0.0144922f $X=11.22 $Y=0.515 $X2=0 $Y2=0
cc_810 N_Y_c_1159_n N_VGND_c_1460_n 0.00904371f $X=4.78 $Y=0.515 $X2=0 $Y2=0
cc_811 N_Y_c_1160_n N_VGND_c_1460_n 0.0078668f $X=5.64 $Y=0.515 $X2=0 $Y2=0
cc_812 N_Y_c_1161_n N_VGND_c_1460_n 0.00856206f $X=6.57 $Y=0.515 $X2=0 $Y2=0
cc_813 N_Y_c_1162_n N_VGND_c_1460_n 0.00888316f $X=7.5 $Y=0.515 $X2=0 $Y2=0
cc_814 N_Y_c_1163_n N_VGND_c_1460_n 0.00904371f $X=8.43 $Y=0.515 $X2=0 $Y2=0
cc_815 N_Y_c_1164_n N_VGND_c_1460_n 0.00904371f $X=9.36 $Y=0.515 $X2=0 $Y2=0
cc_816 N_Y_c_1165_n N_VGND_c_1460_n 0.00904371f $X=10.29 $Y=0.515 $X2=0 $Y2=0
cc_817 N_Y_c_1166_n N_VGND_c_1460_n 0.0118826f $X=11.22 $Y=0.515 $X2=0 $Y2=0
