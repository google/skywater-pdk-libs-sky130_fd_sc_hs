* File: sky130_fd_sc_hs__o221ai_1.spice
* Created: Thu Aug 27 20:59:36 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hs__o221ai_1.pex.spice"
.subckt sky130_fd_sc_hs__o221ai_1  VNB VPB C1 B1 B2 A2 A1 Y VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* Y	Y
* A1	A1
* A2	A2
* B2	B2
* B1	B1
* C1	C1
* VPB	VPB
* VNB	VNB
MM1009 N_A_114_74#_M1009_d N_C1_M1009_g N_Y_M1009_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.2627 AS=0.2109 PD=2.19 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75000.3 A=0.111 P=1.78 MULT=1
MM1006 N_A_114_74#_M1006_d N_B1_M1006_g N_A_239_74#_M1006_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1295 AS=0.2109 PD=1.09 PS=2.05 NRD=11.34 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75002 A=0.111 P=1.78 MULT=1
MM1005 N_A_239_74#_M1005_d N_B2_M1005_g N_A_114_74#_M1006_d VNB NLOWVT L=0.15
+ W=0.74 AD=0.1295 AS=0.1295 PD=1.09 PS=1.09 NRD=11.34 NRS=0 M=1 R=4.93333
+ SA=75000.7 SB=75001.5 A=0.111 P=1.78 MULT=1
MM1004 N_VGND_M1004_d N_A2_M1004_g N_A_239_74#_M1005_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.2368 AS=0.1295 PD=1.38 PS=1.09 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.2
+ SB=75001 A=0.111 P=1.78 MULT=1
MM1007 N_A_239_74#_M1007_d N_A1_M1007_g N_VGND_M1004_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.2368 PD=2.05 PS=1.38 NRD=0 NRS=0 M=1 R=4.93333 SA=75002
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1001 N_VPWR_M1001_d N_C1_M1001_g N_Y_M1001_s VPB PSHORT L=0.15 W=1.12
+ AD=0.4256 AS=0.3304 PD=1.88 PS=2.83 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75002.7 A=0.168 P=2.54 MULT=1
MM1008 A_324_368# N_B1_M1008_g N_VPWR_M1001_d VPB PSHORT L=0.15 W=1.12 AD=0.1512
+ AS=0.4256 PD=1.39 PS=1.88 NRD=14.0658 NRS=1.7533 M=1 R=7.46667 SA=75001.1
+ SB=75001.8 A=0.168 P=2.54 MULT=1
MM1000 N_Y_M1000_d N_B2_M1000_g A_324_368# VPB PSHORT L=0.15 W=1.12 AD=0.2352
+ AS=0.1512 PD=1.54 PS=1.39 NRD=1.7533 NRS=14.0658 M=1 R=7.46667 SA=75001.5
+ SB=75001.4 A=0.168 P=2.54 MULT=1
MM1003 A_522_368# N_A2_M1003_g N_Y_M1000_d VPB PSHORT L=0.15 W=1.12 AD=0.2352
+ AS=0.2352 PD=1.54 PS=1.54 NRD=27.2451 NRS=22.852 M=1 R=7.46667 SA=75002.1
+ SB=75000.8 A=0.168 P=2.54 MULT=1
MM1002 N_VPWR_M1002_d N_A1_M1002_g A_522_368# VPB PSHORT L=0.15 W=1.12 AD=0.3304
+ AS=0.2352 PD=2.83 PS=1.54 NRD=1.7533 NRS=27.2451 M=1 R=7.46667 SA=75002.7
+ SB=75000.2 A=0.168 P=2.54 MULT=1
DX10_noxref VNB VPB NWDIODE A=7.8492 P=12.16
*
.include "sky130_fd_sc_hs__o221ai_1.pxi.spice"
*
.ends
*
*
