* File: sky130_fd_sc_hs__clkinv_8.spice
* Created: Thu Aug 27 20:37:19 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hs__clkinv_8.pex.spice"
.subckt sky130_fd_sc_hs__clkinv_8  VNB VPB A VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A	A
* VPB	VPB
* VNB	VNB
MM1000 N_Y_M1000_d N_A_M1000_g N_VGND_M1000_s VNB NLOWVT L=0.15 W=0.42 AD=0.4221
+ AS=0.1281 PD=2.43 PS=1.45 NRD=14.28 NRS=5.712 M=1 R=2.8 SA=75000.2 SB=75005.4
+ A=0.063 P=1.14 MULT=1
MM1001 N_Y_M1000_d N_A_M1001_g N_VGND_M1001_s VNB NLOWVT L=0.15 W=0.42 AD=0.4221
+ AS=0.0882 PD=2.43 PS=0.84 NRD=0 NRS=19.992 M=1 R=2.8 SA=75002.4 SB=75003.3
+ A=0.063 P=1.14 MULT=1
MM1004 N_Y_M1004_d N_A_M1004_g N_VGND_M1001_s VNB NLOWVT L=0.15 W=0.42 AD=0.0588
+ AS=0.0882 PD=0.7 PS=0.84 NRD=0 NRS=19.992 M=1 R=2.8 SA=75003 SB=75002.7
+ A=0.063 P=1.14 MULT=1
MM1005 N_Y_M1004_d N_A_M1005_g N_VGND_M1005_s VNB NLOWVT L=0.15 W=0.42 AD=0.0588
+ AS=0.0882 PD=0.7 PS=0.84 NRD=0 NRS=19.992 M=1 R=2.8 SA=75003.4 SB=75002.3
+ A=0.063 P=1.14 MULT=1
MM1006 N_Y_M1006_d N_A_M1006_g N_VGND_M1005_s VNB NLOWVT L=0.15 W=0.42 AD=0.0588
+ AS=0.0882 PD=0.7 PS=0.84 NRD=0 NRS=19.992 M=1 R=2.8 SA=75004 SB=75001.7
+ A=0.063 P=1.14 MULT=1
MM1016 N_Y_M1006_d N_A_M1016_g N_VGND_M1016_s VNB NLOWVT L=0.15 W=0.42 AD=0.0588
+ AS=0.0882 PD=0.7 PS=0.84 NRD=0 NRS=19.992 M=1 R=2.8 SA=75004.4 SB=75001.3
+ A=0.063 P=1.14 MULT=1
MM1017 N_Y_M1017_d N_A_M1017_g N_VGND_M1016_s VNB NLOWVT L=0.15 W=0.42 AD=0.0735
+ AS=0.0882 PD=0.77 PS=0.84 NRD=0 NRS=19.992 M=1 R=2.8 SA=75005 SB=75000.7
+ A=0.063 P=1.14 MULT=1
MM1019 N_Y_M1017_d N_A_M1019_g N_VGND_M1019_s VNB NLOWVT L=0.15 W=0.42 AD=0.0735
+ AS=0.1197 PD=0.77 PS=1.41 NRD=19.992 NRS=0 M=1 R=2.8 SA=75005.5 SB=75000.2
+ A=0.063 P=1.14 MULT=1
MM1002 N_Y_M1002_d N_A_M1002_g N_VPWR_M1002_s VPB PSHORT L=0.15 W=1.12 AD=0.168
+ AS=0.3584 PD=1.42 PS=2.88 NRD=1.7533 NRS=4.3931 M=1 R=7.46667 SA=75000.2
+ SB=75005.4 A=0.168 P=2.54 MULT=1
MM1003 N_Y_M1002_d N_A_M1003_g N_VPWR_M1003_s VPB PSHORT L=0.15 W=1.12 AD=0.168
+ AS=0.196 PD=1.42 PS=1.47 NRD=1.7533 NRS=1.7533 M=1 R=7.46667 SA=75000.7
+ SB=75005 A=0.168 P=2.54 MULT=1
MM1007 N_Y_M1007_d N_A_M1007_g N_VPWR_M1003_s VPB PSHORT L=0.15 W=1.12 AD=0.168
+ AS=0.196 PD=1.42 PS=1.47 NRD=1.7533 NRS=10.5395 M=1 R=7.46667 SA=75001.2
+ SB=75004.5 A=0.168 P=2.54 MULT=1
MM1008 N_Y_M1007_d N_A_M1008_g N_VPWR_M1008_s VPB PSHORT L=0.15 W=1.12 AD=0.168
+ AS=0.196 PD=1.42 PS=1.47 NRD=1.7533 NRS=1.7533 M=1 R=7.46667 SA=75001.6
+ SB=75004 A=0.168 P=2.54 MULT=1
MM1009 N_Y_M1009_d N_A_M1009_g N_VPWR_M1008_s VPB PSHORT L=0.15 W=1.12 AD=0.168
+ AS=0.196 PD=1.42 PS=1.47 NRD=1.7533 NRS=10.5395 M=1 R=7.46667 SA=75002.1
+ SB=75003.5 A=0.168 P=2.54 MULT=1
MM1010 N_Y_M1009_d N_A_M1010_g N_VPWR_M1010_s VPB PSHORT L=0.15 W=1.12 AD=0.168
+ AS=0.196 PD=1.42 PS=1.47 NRD=1.7533 NRS=1.7533 M=1 R=7.46667 SA=75002.6
+ SB=75003.1 A=0.168 P=2.54 MULT=1
MM1011 N_Y_M1011_d N_A_M1011_g N_VPWR_M1010_s VPB PSHORT L=0.15 W=1.12 AD=0.168
+ AS=0.196 PD=1.42 PS=1.47 NRD=1.7533 NRS=10.5395 M=1 R=7.46667 SA=75003.1
+ SB=75002.6 A=0.168 P=2.54 MULT=1
MM1012 N_Y_M1011_d N_A_M1012_g N_VPWR_M1012_s VPB PSHORT L=0.15 W=1.12 AD=0.168
+ AS=0.196 PD=1.42 PS=1.47 NRD=1.7533 NRS=1.7533 M=1 R=7.46667 SA=75003.5
+ SB=75002.1 A=0.168 P=2.54 MULT=1
MM1013 N_Y_M1013_d N_A_M1013_g N_VPWR_M1012_s VPB PSHORT L=0.15 W=1.12 AD=0.168
+ AS=0.196 PD=1.42 PS=1.47 NRD=1.7533 NRS=10.5395 M=1 R=7.46667 SA=75004
+ SB=75001.6 A=0.168 P=2.54 MULT=1
MM1014 N_Y_M1013_d N_A_M1014_g N_VPWR_M1014_s VPB PSHORT L=0.15 W=1.12 AD=0.168
+ AS=0.196 PD=1.42 PS=1.47 NRD=1.7533 NRS=1.7533 M=1 R=7.46667 SA=75004.5
+ SB=75001.2 A=0.168 P=2.54 MULT=1
MM1015 N_Y_M1015_d N_A_M1015_g N_VPWR_M1014_s VPB PSHORT L=0.15 W=1.12 AD=0.168
+ AS=0.196 PD=1.42 PS=1.47 NRD=1.7533 NRS=10.5395 M=1 R=7.46667 SA=75005
+ SB=75000.7 A=0.168 P=2.54 MULT=1
MM1018 N_Y_M1015_d N_A_M1018_g N_VPWR_M1018_s VPB PSHORT L=0.15 W=1.12 AD=0.168
+ AS=0.3304 PD=1.42 PS=2.83 NRD=1.7533 NRS=1.7533 M=1 R=7.46667 SA=75005.4
+ SB=75000.2 A=0.168 P=2.54 MULT=1
DX20_noxref VNB VPB NWDIODE A=12.3132 P=16.96
*
.include "sky130_fd_sc_hs__clkinv_8.pxi.spice"
*
.ends
*
*
