* NGSPICE file created from sky130_fd_sc_hs__clkinv_16.ext - technology: sky130A

.subckt sky130_fd_sc_hs__clkinv_16 A VGND VNB VPB VPWR Y
M1000 Y A VGND VNB nlowvt w=420000u l=150000u
+  ad=9.408e+11p pd=1.12e+07u as=1.83765e+12p ps=1.762e+07u
M1001 Y A VGND VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1002 Y A VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=4.0992e+12p pd=3.42e+07u as=4.4688e+12p ps=3.71e+07u
M1003 VPWR A Y VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 Y A VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VGND A Y VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 Y A VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VPWR A Y VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 Y A VGND VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VGND A Y VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VPWR A Y VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VPWR A Y VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 Y A VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 Y A VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 Y A VGND VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VPWR A Y VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VGND A Y VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 Y A VGND VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 Y A VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 Y A VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 VPWR A Y VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 VPWR A Y VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 Y A VGND VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 Y A VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 Y A VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 Y A VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 VPWR A Y VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 VGND A Y VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1028 Y A VGND VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1029 VPWR A Y VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1030 VGND A Y VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1031 Y A VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1032 Y A VGND VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1033 VPWR A Y VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1034 Y A VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1035 VPWR A Y VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1036 VGND A Y VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1037 VGND A Y VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1038 VGND A Y VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1039 VPWR A Y VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

