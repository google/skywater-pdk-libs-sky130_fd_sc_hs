* File: sky130_fd_sc_hs__o41a_1.spice
* Created: Thu Aug 27 21:04:08 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hs__o41a_1.pex.spice"
.subckt sky130_fd_sc_hs__o41a_1  VNB VPB B1 A4 A3 A2 A1 X VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* X	X
* A1	A1
* A2	A2
* A3	A3
* A4	A4
* B1	B1
* VPB	VPB
* VNB	VNB
MM1010 N_VGND_M1010_d N_A_83_270#_M1010_g N_X_M1010_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.2627 AS=0.2109 PD=2.19 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75000.3 A=0.111 P=1.78 MULT=1
MM1004 N_A_326_74#_M1004_d N_B1_M1004_g N_A_83_270#_M1004_s VNB NLOWVT L=0.15
+ W=0.64 AD=0.112 AS=0.1824 PD=0.99 PS=1.85 NRD=13.116 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75002.5 A=0.096 P=1.58 MULT=1
MM1003 N_VGND_M1003_d N_A4_M1003_g N_A_326_74#_M1004_d VNB NLOWVT L=0.15 W=0.64
+ AD=0.1344 AS=0.112 PD=1.06 PS=0.99 NRD=13.116 NRS=0 M=1 R=4.26667 SA=75000.7
+ SB=75002 A=0.096 P=1.58 MULT=1
MM1011 N_A_326_74#_M1011_d N_A3_M1011_g N_VGND_M1003_d VNB NLOWVT L=0.15 W=0.64
+ AD=0.1088 AS=0.1344 PD=0.98 PS=1.06 NRD=0 NRS=13.116 M=1 R=4.26667 SA=75001.3
+ SB=75001.4 A=0.096 P=1.58 MULT=1
MM1007 N_VGND_M1007_d N_A2_M1007_g N_A_326_74#_M1011_d VNB NLOWVT L=0.15 W=0.64
+ AD=0.1792 AS=0.1088 PD=1.2 PS=0.98 NRD=20.616 NRS=11.244 M=1 R=4.26667
+ SA=75001.8 SB=75000.9 A=0.096 P=1.58 MULT=1
MM1009 N_A_326_74#_M1009_d N_A1_M1009_g N_VGND_M1007_d VNB NLOWVT L=0.15 W=0.64
+ AD=0.1824 AS=0.1792 PD=1.85 PS=1.2 NRD=0 NRS=31.872 M=1 R=4.26667 SA=75002.5
+ SB=75000.2 A=0.096 P=1.58 MULT=1
MM1005 N_VPWR_M1005_d N_A_83_270#_M1005_g N_X_M1005_s VPB PSHORT L=0.15 W=1.12
+ AD=0.538514 AS=0.3304 PD=2.36571 PS=2.83 NRD=10.5395 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75002.8 A=0.168 P=2.54 MULT=1
MM1006 N_A_83_270#_M1006_d N_B1_M1006_g N_VPWR_M1005_d VPB PSHORT L=0.15 W=0.84
+ AD=0.172136 AS=0.403886 PD=1.29 PS=1.77429 NRD=22.261 NRS=23.443 M=1 R=5.6
+ SA=75001.3 SB=75002.4 A=0.126 P=1.98 MULT=1
MM1008 A_443_368# N_A4_M1008_g N_A_83_270#_M1006_d VPB PSHORT L=0.15 W=1.12
+ AD=0.1512 AS=0.229514 PD=1.39 PS=1.72 NRD=14.0658 NRS=1.7533 M=1 R=7.46667
+ SA=75001.4 SB=75001.9 A=0.168 P=2.54 MULT=1
MM1000 A_527_368# N_A3_M1000_g A_443_368# VPB PSHORT L=0.15 W=1.12 AD=0.2352
+ AS=0.1512 PD=1.54 PS=1.39 NRD=27.2451 NRS=14.0658 M=1 R=7.46667 SA=75001.9
+ SB=75001.5 A=0.168 P=2.54 MULT=1
MM1002 A_641_368# N_A2_M1002_g A_527_368# VPB PSHORT L=0.15 W=1.12 AD=0.2352
+ AS=0.2352 PD=1.54 PS=1.54 NRD=27.2451 NRS=27.2451 M=1 R=7.46667 SA=75002.4
+ SB=75000.9 A=0.168 P=2.54 MULT=1
MM1001 N_VPWR_M1001_d N_A1_M1001_g A_641_368# VPB PSHORT L=0.15 W=1.12 AD=0.4592
+ AS=0.2352 PD=3.06 PS=1.54 NRD=1.7533 NRS=27.2451 M=1 R=7.46667 SA=75003
+ SB=75000.3 A=0.168 P=2.54 MULT=1
DX12_noxref VNB VPB NWDIODE A=8.742 P=13.12
*
.include "sky130_fd_sc_hs__o41a_1.pxi.spice"
*
.ends
*
*
