* File: sky130_fd_sc_hs__nand3b_1.pex.spice
* Created: Thu Aug 27 20:51:17 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HS__NAND3B_1%A_N 3 5 7 8 12
r26 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.61
+ $Y=1.515 $X2=0.61 $Y2=1.515
r27 8 12 4.43247 $w=3.88e-07 $l=1.5e-07 $layer=LI1_cond $X=0.64 $Y=1.665
+ $X2=0.64 $Y2=1.515
r28 5 11 51.3895 $w=3.19e-07 $l=2.79732e-07 $layer=POLY_cond $X=0.66 $Y=1.765
+ $X2=0.597 $Y2=1.515
r29 5 7 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=0.66 $Y=1.765 $X2=0.66
+ $Y2=2.26
r30 1 11 38.5462 $w=3.19e-07 $l=2.09893e-07 $layer=POLY_cond $X=0.495 $Y=1.35
+ $X2=0.597 $Y2=1.515
r31 1 3 253.819 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=0.495 $Y=1.35
+ $X2=0.495 $Y2=0.855
.ends

.subckt PM_SKY130_FD_SC_HS__NAND3B_1%C 1 3 6 8 12
r28 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.18
+ $Y=1.515 $X2=1.18 $Y2=1.515
r29 8 12 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=1.18 $Y=1.665
+ $X2=1.18 $Y2=1.515
r30 4 11 38.5562 $w=2.99e-07 $l=2.05122e-07 $layer=POLY_cond $X=1.27 $Y=1.35
+ $X2=1.18 $Y2=1.515
r31 4 6 302.532 $w=1.5e-07 $l=5.9e-07 $layer=POLY_cond $X=1.27 $Y=1.35 $X2=1.27
+ $Y2=0.76
r32 1 11 52.2586 $w=2.99e-07 $l=2.80624e-07 $layer=POLY_cond $X=1.245 $Y=1.765
+ $X2=1.18 $Y2=1.515
r33 1 3 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.245 $Y=1.765
+ $X2=1.245 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_HS__NAND3B_1%B 3 5 7 8 12
r33 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.75
+ $Y=1.515 $X2=1.75 $Y2=1.515
r34 8 12 4.93904 $w=3.48e-07 $l=1.5e-07 $layer=LI1_cond $X=1.74 $Y=1.665
+ $X2=1.74 $Y2=1.515
r35 5 11 52.2586 $w=2.99e-07 $l=2.76134e-07 $layer=POLY_cond $X=1.695 $Y=1.765
+ $X2=1.75 $Y2=1.515
r36 5 7 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.695 $Y=1.765
+ $X2=1.695 $Y2=2.4
r37 1 11 38.5562 $w=2.99e-07 $l=2.05122e-07 $layer=POLY_cond $X=1.66 $Y=1.35
+ $X2=1.75 $Y2=1.515
r38 1 3 302.532 $w=1.5e-07 $l=5.9e-07 $layer=POLY_cond $X=1.66 $Y=1.35 $X2=1.66
+ $Y2=0.76
.ends

.subckt PM_SKY130_FD_SC_HS__NAND3B_1%A_27_116# 1 2 9 11 13 16 22 25 26 28 29 33
r62 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.29
+ $Y=1.485 $X2=2.29 $Y2=1.485
r63 30 33 4.1907 $w=3.28e-07 $l=1.2e-07 $layer=LI1_cond $X=2.17 $Y=1.485
+ $X2=2.29 $Y2=1.485
r64 28 29 9.48656 $w=4.93e-07 $l=1.65e-07 $layer=LI1_cond $X=0.352 $Y=2.115
+ $X2=0.352 $Y2=1.95
r65 25 30 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.17 $Y=1.32
+ $X2=2.17 $Y2=1.485
r66 24 25 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=2.17 $Y=1.15
+ $X2=2.17 $Y2=1.32
r67 23 26 2.28545 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=0.375 $Y=1.065
+ $X2=0.24 $Y2=1.065
r68 22 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.085 $Y=1.065
+ $X2=2.17 $Y2=1.15
r69 22 23 111.561 $w=1.68e-07 $l=1.71e-06 $layer=LI1_cond $X=2.085 $Y=1.065
+ $X2=0.375 $Y2=1.065
r70 18 26 4.14756 $w=2.2e-07 $l=1.07121e-07 $layer=LI1_cond $X=0.19 $Y=1.15
+ $X2=0.24 $Y2=1.065
r71 18 29 52.1925 $w=1.68e-07 $l=8e-07 $layer=LI1_cond $X=0.19 $Y=1.15 $X2=0.19
+ $Y2=1.95
r72 14 26 4.14756 $w=2.2e-07 $l=8.5e-08 $layer=LI1_cond $X=0.24 $Y=0.98 $X2=0.24
+ $Y2=1.065
r73 14 16 5.33538 $w=2.68e-07 $l=1.25e-07 $layer=LI1_cond $X=0.24 $Y=0.98
+ $X2=0.24 $Y2=0.855
r74 11 34 57.6553 $w=2.91e-07 $l=3.01662e-07 $layer=POLY_cond $X=2.245 $Y=1.765
+ $X2=2.29 $Y2=1.485
r75 11 13 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.245 $Y=1.765
+ $X2=2.245 $Y2=2.4
r76 7 34 38.6072 $w=2.91e-07 $l=2.05122e-07 $layer=POLY_cond $X=2.2 $Y=1.32
+ $X2=2.29 $Y2=1.485
r77 7 9 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=2.2 $Y=1.32 $X2=2.2
+ $Y2=0.76
r78 2 28 300 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_PDIFF $count=2 $X=0.29
+ $Y=1.84 $X2=0.435 $Y2=2.115
r79 1 16 182 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.58 $X2=0.28 $Y2=0.855
.ends

.subckt PM_SKY130_FD_SC_HS__NAND3B_1%VPWR 1 2 9 15 18 19 21 22 23 33 34
r35 33 34 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r36 31 34 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.64 $Y2=3.33
r37 30 31 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r38 26 27 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r39 23 31 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.44 $Y=3.33
+ $X2=1.68 $Y2=3.33
r40 23 27 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.44 $Y=3.33
+ $X2=0.72 $Y2=3.33
r41 21 30 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=1.805 $Y=3.33
+ $X2=1.68 $Y2=3.33
r42 21 22 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.805 $Y=3.33
+ $X2=1.97 $Y2=3.33
r43 20 33 32.9465 $w=1.68e-07 $l=5.05e-07 $layer=LI1_cond $X=2.135 $Y=3.33
+ $X2=2.64 $Y2=3.33
r44 20 22 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.135 $Y=3.33
+ $X2=1.97 $Y2=3.33
r45 18 26 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=0.805 $Y=3.33
+ $X2=0.72 $Y2=3.33
r46 18 19 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.805 $Y=3.33
+ $X2=0.97 $Y2=3.33
r47 17 30 35.5561 $w=1.68e-07 $l=5.45e-07 $layer=LI1_cond $X=1.135 $Y=3.33
+ $X2=1.68 $Y2=3.33
r48 17 19 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.135 $Y=3.33
+ $X2=0.97 $Y2=3.33
r49 13 22 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.97 $Y=3.245
+ $X2=1.97 $Y2=3.33
r50 13 15 27.5888 $w=3.28e-07 $l=7.9e-07 $layer=LI1_cond $X=1.97 $Y=3.245
+ $X2=1.97 $Y2=2.455
r51 9 12 27.2396 $w=3.28e-07 $l=7.8e-07 $layer=LI1_cond $X=0.97 $Y=2.035
+ $X2=0.97 $Y2=2.815
r52 7 19 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.97 $Y=3.245 $X2=0.97
+ $Y2=3.33
r53 7 12 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=0.97 $Y=3.245
+ $X2=0.97 $Y2=2.815
r54 2 15 300 $w=1.7e-07 $l=7.07972e-07 $layer=licon1_PDIFF $count=2 $X=1.77
+ $Y=1.84 $X2=1.97 $Y2=2.455
r55 1 12 600 $w=1.7e-07 $l=1.08616e-06 $layer=licon1_PDIFF $count=1 $X=0.735
+ $Y=1.84 $X2=0.97 $Y2=2.815
r56 1 9 300 $w=1.7e-07 $l=3.17884e-07 $layer=licon1_PDIFF $count=2 $X=0.735
+ $Y=1.84 $X2=0.97 $Y2=2.035
.ends

.subckt PM_SKY130_FD_SC_HS__NAND3B_1%Y 1 2 3 10 12 14 16 24 25 26 41 42
r41 41 42 9.45624 $w=4.88e-07 $l=1.65e-07 $layer=LI1_cond $X=2.55 $Y=1.985
+ $X2=2.55 $Y2=1.82
r42 26 38 0.976391 $w=4.88e-07 $l=4e-08 $layer=LI1_cond $X=2.55 $Y=2.775
+ $X2=2.55 $Y2=2.815
r43 25 26 9.03161 $w=4.88e-07 $l=3.7e-07 $layer=LI1_cond $X=2.55 $Y=2.405
+ $X2=2.55 $Y2=2.775
r44 24 41 1.22049 $w=4.88e-07 $l=5e-08 $layer=LI1_cond $X=2.55 $Y=2.035 $X2=2.55
+ $Y2=1.985
r45 24 25 5.98354 $w=6.58e-07 $l=2.85e-07 $layer=LI1_cond $X=2.55 $Y=2.12
+ $X2=2.55 $Y2=2.405
r46 21 23 11.8319 $w=4.64e-07 $l=4.5e-07 $layer=LI1_cond $X=2.522 $Y=0.535
+ $X2=2.522 $Y2=0.985
r47 16 23 9.48898 $w=4.64e-07 $l=2.57612e-07 $layer=LI1_cond $X=2.71 $Y=1.15
+ $X2=2.522 $Y2=0.985
r48 16 42 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.71 $Y=1.15
+ $X2=2.71 $Y2=1.82
r49 15 19 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.635 $Y=2.035
+ $X2=1.47 $Y2=2.035
r50 14 24 7.03003 $w=1.7e-07 $l=2.45e-07 $layer=LI1_cond $X=2.305 $Y=2.035
+ $X2=2.55 $Y2=2.035
r51 14 15 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.305 $Y=2.035
+ $X2=1.635 $Y2=2.035
r52 10 19 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.47 $Y=2.12 $X2=1.47
+ $Y2=2.035
r53 10 12 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=1.47 $Y=2.12
+ $X2=1.47 $Y2=2.815
r54 3 41 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=2.32
+ $Y=1.84 $X2=2.47 $Y2=1.985
r55 3 38 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=2.32
+ $Y=1.84 $X2=2.47 $Y2=2.815
r56 2 19 400 $w=1.7e-07 $l=3.4187e-07 $layer=licon1_PDIFF $count=1 $X=1.32
+ $Y=1.84 $X2=1.47 $Y2=2.115
r57 2 12 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=1.32
+ $Y=1.84 $X2=1.47 $Y2=2.815
r58 1 23 182 $w=1.7e-07 $l=7.35833e-07 $layer=licon1_NDIFF $count=1 $X=2.275
+ $Y=0.39 $X2=2.59 $Y2=0.985
r59 1 21 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=2.275
+ $Y=0.39 $X2=2.415 $Y2=0.535
.ends

.subckt PM_SKY130_FD_SC_HS__NAND3B_1%VGND 1 6 8 10 17 18 21
r23 22 24 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r24 21 24 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r25 21 22 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r26 17 18 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r27 15 21 13.399 $w=1.7e-07 $l=3.38e-07 $layer=LI1_cond $X=1.22 $Y=0 $X2=0.882
+ $Y2=0
r28 15 17 92.6417 $w=1.68e-07 $l=1.42e-06 $layer=LI1_cond $X=1.22 $Y=0 $X2=2.64
+ $Y2=0
r29 13 24 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r30 12 13 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r31 10 21 13.399 $w=1.7e-07 $l=3.37e-07 $layer=LI1_cond $X=0.545 $Y=0 $X2=0.882
+ $Y2=0
r32 10 12 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.545 $Y=0 $X2=0.24
+ $Y2=0
r33 8 18 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=1.44 $Y=0 $X2=2.64
+ $Y2=0
r34 8 22 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.44 $Y=0 $X2=1.2
+ $Y2=0
r35 4 21 2.78459 $w=6.75e-07 $l=8.5e-08 $layer=LI1_cond $X=0.882 $Y=0.085
+ $X2=0.882 $Y2=0
r36 4 6 11.3406 $w=6.73e-07 $l=6.4e-07 $layer=LI1_cond $X=0.882 $Y=0.085
+ $X2=0.882 $Y2=0.725
r37 1 6 91 $w=1.7e-07 $l=5.52766e-07 $layer=licon1_NDIFF $count=2 $X=0.57
+ $Y=0.58 $X2=1.055 $Y2=0.725
.ends

