* File: sky130_fd_sc_hs__dfbbn_2.spice
* Created: Tue Sep  1 19:59:27 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hs__dfbbn_2.pex.spice"
.subckt sky130_fd_sc_hs__dfbbn_2  VNB VPB CLK_N D SET_B RESET_B VPWR Q_N Q VGND
* 
* VGND	VGND
* Q	Q
* Q_N	Q_N
* VPWR	VPWR
* RESET_B	RESET_B
* SET_B	SET_B
* D	D
* CLK_N	CLK_N
* VPB	VPB
* VNB	VNB
MM1034 N_VGND_M1034_d N_CLK_N_M1034_g N_A_27_74#_M1034_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.2109 PD=1.02 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75000.6 A=0.111 P=1.78 MULT=1
MM1035 N_A_200_74#_M1035_d N_A_27_74#_M1035_g N_VGND_M1034_d VNB NLOWVT L=0.15
+ W=0.74 AD=0.2109 AS=0.1036 PD=2.05 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.6 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1012 N_VGND_M1012_d N_D_M1012_g N_A_311_119#_M1012_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.133562 AS=0.1197 PD=1.08 PS=1.41 NRD=32.856 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75002 A=0.063 P=1.14 MULT=1
MM1033 A_529_119# N_A_473_405#_M1033_g N_VGND_M1012_d VNB NLOWVT L=0.15 W=0.42
+ AD=0.0441 AS=0.133562 PD=0.63 PS=1.08 NRD=14.28 NRS=34.284 M=1 R=2.8
+ SA=75000.9 SB=75001.3 A=0.063 P=1.14 MULT=1
MM1042 N_A_601_119#_M1042_d N_A_27_74#_M1042_g A_529_119# VNB NLOWVT L=0.15
+ W=0.42 AD=0.0588 AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75001.2
+ SB=75001 A=0.063 P=1.14 MULT=1
MM1023 N_A_311_119#_M1023_d N_A_200_74#_M1023_g N_A_601_119#_M1042_d VNB NLOWVT
+ L=0.15 W=0.42 AD=0.38115 AS=0.0588 PD=2.52 PS=0.7 NRD=243.564 NRS=0 M=1 R=2.8
+ SA=75001.7 SB=75000.6 A=0.063 P=1.14 MULT=1
MM1039 N_A_473_405#_M1039_d N_A_601_119#_M1039_g N_A_867_125#_M1039_s VNB NLOWVT
+ L=0.15 W=0.55 AD=0.077 AS=0.15675 PD=0.83 PS=1.67 NRD=0 NRS=0 M=1 R=3.66667
+ SA=75000.2 SB=75004.7 A=0.0825 P=1.4 MULT=1
MM1005 N_A_867_125#_M1005_d N_A_975_322#_M1005_g N_A_473_405#_M1039_d VNB NLOWVT
+ L=0.15 W=0.55 AD=0.09625 AS=0.077 PD=0.9 PS=0.83 NRD=15.264 NRS=0 M=1
+ R=3.66667 SA=75000.6 SB=75004.3 A=0.0825 P=1.4 MULT=1
MM1004 N_VGND_M1004_d N_SET_B_M1004_g N_A_867_125#_M1005_d VNB NLOWVT L=0.15
+ W=0.55 AD=0.09625 AS=0.09625 PD=0.9 PS=0.9 NRD=15.264 NRS=0 M=1 R=3.66667
+ SA=75001.1 SB=75003.8 A=0.0825 P=1.4 MULT=1
MM1002 A_1240_125# N_A_473_405#_M1002_g N_VGND_M1004_d VNB NLOWVT L=0.15 W=0.55
+ AD=0.0950625 AS=0.09625 PD=0.94 PS=0.9 NRD=25.704 NRS=0 M=1 R=3.66667
+ SA=75001.6 SB=75003.3 A=0.0825 P=1.4 MULT=1
MM1037 N_A_1335_112#_M1037_d N_A_27_74#_M1037_g A_1240_125# VNB NLOWVT L=0.15
+ W=0.55 AD=0.345876 AS=0.0950625 PD=2.18299 PS=0.94 NRD=0 NRS=25.704 M=1
+ R=3.66667 SA=75001.9 SB=75002.8 A=0.0825 P=1.4 MULT=1
MM1003 A_1640_138# N_A_200_74#_M1003_g N_A_1335_112#_M1037_d VNB NLOWVT L=0.15
+ W=0.42 AD=0.0504 AS=0.264124 PD=0.66 PS=1.66701 NRD=18.564 NRS=0 M=1 R=2.8
+ SA=75003.6 SB=75002.1 A=0.063 P=1.14 MULT=1
MM1013 N_VGND_M1013_d N_A_1555_410#_M1013_g A_1640_138# VNB NLOWVT L=0.15 W=0.42
+ AD=0.0968897 AS=0.0504 PD=0.84 PS=0.66 NRD=50.196 NRS=18.564 M=1 R=2.8
+ SA=75004 SB=75001.7 A=0.063 P=1.14 MULT=1
MM1008 N_A_1832_74#_M1008_d N_SET_B_M1008_g N_VGND_M1013_d VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.17071 PD=1.02 PS=1.48 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75002.7 SB=75001.2 A=0.111 P=1.78 MULT=1
MM1014 N_A_1555_410#_M1014_d N_A_975_322#_M1014_g N_A_1832_74#_M1008_d VNB
+ NLOWVT L=0.15 W=0.74 AD=0.1184 AS=0.1036 PD=1.06 PS=1.02 NRD=6.48 NRS=0 M=1
+ R=4.93333 SA=75003.1 SB=75000.8 A=0.111 P=1.78 MULT=1
MM1007 N_A_1832_74#_M1007_d N_A_1335_112#_M1007_g N_A_1555_410#_M1014_d VNB
+ NLOWVT L=0.15 W=0.74 AD=0.2907 AS=0.1184 PD=2.39 PS=1.06 NRD=12.972 NRS=0 M=1
+ R=4.93333 SA=75003.6 SB=75000.3 A=0.111 P=1.78 MULT=1
MM1020 N_VGND_M1020_d N_RESET_B_M1020_g N_A_975_322#_M1020_s VNB NLOWVT L=0.15
+ W=0.42 AD=0.171892 AS=0.1176 PD=1.45552 PS=1.4 NRD=101.208 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75001.2 A=0.063 P=1.14 MULT=1
MM1031 N_VGND_M1020_d N_A_1555_410#_M1031_g N_Q_N_M1031_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.302858 AS=0.1036 PD=2.56448 PS=1.02 NRD=57.444 NRS=0 M=1 R=4.93333
+ SA=75000.5 SB=75000.7 A=0.111 P=1.78 MULT=1
MM1043 N_VGND_M1043_d N_A_1555_410#_M1043_g N_Q_N_M1031_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.222 AS=0.1036 PD=2.08 PS=1.02 NRD=2.424 NRS=0 M=1 R=4.93333
+ SA=75000.9 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1028 N_VGND_M1028_d N_A_1555_410#_M1028_g N_A_2516_368#_M1028_s VNB NLOWVT
+ L=0.15 W=0.64 AD=0.108058 AS=0.1824 PD=0.987826 PS=1.85 NRD=5.616 NRS=0 M=1
+ R=4.26667 SA=75000.2 SB=75001.1 A=0.096 P=1.58 MULT=1
MM1006 N_Q_M1006_d N_A_2516_368#_M1006_g N_VGND_M1028_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.124942 PD=1.02 PS=1.14217 NRD=0 NRS=2.424 M=1 R=4.93333
+ SA=75000.6 SB=75000.6 A=0.111 P=1.78 MULT=1
MM1029 N_Q_M1006_d N_A_2516_368#_M1029_g N_VGND_M1029_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1998 PD=1.02 PS=2.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1000 N_VPWR_M1000_d N_CLK_N_M1000_g N_A_27_74#_M1000_s VPB PSHORT L=0.15
+ W=1.12 AD=0.168 AS=0.3192 PD=1.42 PS=2.81 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1001 N_A_200_74#_M1001_d N_A_27_74#_M1001_g N_VPWR_M1000_d VPB PSHORT L=0.15
+ W=1.12 AD=0.3136 AS=0.168 PD=2.8 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.7 SB=75000.2 A=0.168 P=2.54 MULT=1
MM1030 N_VPWR_M1030_d N_D_M1030_g N_A_311_119#_M1030_s VPB PSHORT L=0.15 W=0.42
+ AD=0.09345 AS=0.17805 PD=0.865 PS=1.75 NRD=72.693 NRS=46.886 M=1 R=2.8
+ SA=75000.3 SB=75001.8 A=0.063 P=1.14 MULT=1
MM1026 A_536_503# N_A_473_405#_M1026_g N_VPWR_M1030_d VPB PSHORT L=0.15 W=0.42
+ AD=0.0567 AS=0.09345 PD=0.69 PS=0.865 NRD=37.5088 NRS=4.6886 M=1 R=2.8
+ SA=75000.9 SB=75001.2 A=0.063 P=1.14 MULT=1
MM1010 N_A_601_119#_M1010_d N_A_200_74#_M1010_g A_536_503# VPB PSHORT L=0.15
+ W=0.42 AD=0.0756 AS=0.0567 PD=0.78 PS=0.69 NRD=18.7544 NRS=37.5088 M=1 R=2.8
+ SA=75001.3 SB=75000.8 A=0.063 P=1.14 MULT=1
MM1032 N_A_311_119#_M1032_d N_A_27_74#_M1032_g N_A_601_119#_M1010_d VPB PSHORT
+ L=0.15 W=0.42 AD=0.1653 AS=0.0756 PD=1.7 PS=0.78 NRD=37.5088 NRS=18.7544 M=1
+ R=2.8 SA=75001.8 SB=75000.3 A=0.063 P=1.14 MULT=1
MM1021 A_930_424# N_A_601_119#_M1021_g N_A_473_405#_M1021_s VPB PSHORT L=0.15
+ W=0.84 AD=0.1134 AS=0.2352 PD=1.11 PS=2.24 NRD=18.7544 NRS=2.3443 M=1 R=5.6
+ SA=75000.2 SB=75001.1 A=0.126 P=1.98 MULT=1
MM1040 N_VPWR_M1040_d N_A_975_322#_M1040_g A_930_424# VPB PSHORT L=0.15 W=0.84
+ AD=0.1512 AS=0.1134 PD=1.2 PS=1.11 NRD=2.3443 NRS=18.7544 M=1 R=5.6 SA=75000.6
+ SB=75000.7 A=0.126 P=1.98 MULT=1
MM1022 N_A_473_405#_M1022_d N_SET_B_M1022_g N_VPWR_M1040_d VPB PSHORT L=0.15
+ W=0.84 AD=0.2352 AS=0.1512 PD=2.24 PS=1.2 NRD=2.3443 NRS=16.4101 M=1 R=5.6
+ SA=75001.1 SB=75000.2 A=0.126 P=1.98 MULT=1
MM1015 A_1312_424# N_A_473_405#_M1015_g N_VPWR_M1015_s VPB PSHORT L=0.15 W=0.84
+ AD=0.1134 AS=0.2352 PD=1.11 PS=2.24 NRD=18.7544 NRS=2.3443 M=1 R=5.6
+ SA=75000.2 SB=75001.2 A=0.126 P=1.98 MULT=1
MM1027 N_A_1335_112#_M1027_d N_A_200_74#_M1027_g A_1312_424# VPB PSHORT L=0.15
+ W=0.84 AD=0.1918 AS=0.1134 PD=1.64 PS=1.11 NRD=2.3443 NRS=18.7544 M=1 R=5.6
+ SA=75000.6 SB=75000.7 A=0.126 P=1.98 MULT=1
MM1011 A_1504_508# N_A_27_74#_M1011_g N_A_1335_112#_M1027_d VPB PSHORT L=0.15
+ W=0.42 AD=0.0567 AS=0.0959 PD=0.69 PS=0.82 NRD=37.5088 NRS=46.886 M=1 R=2.8
+ SA=75001.2 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1016 N_VPWR_M1016_d N_A_1555_410#_M1016_g A_1504_508# VPB PSHORT L=0.15 W=0.42
+ AD=0.22775 AS=0.0567 PD=2.07 PS=0.69 NRD=228.54 NRS=37.5088 M=1 R=2.8
+ SA=75001.6 SB=75000.3 A=0.063 P=1.14 MULT=1
MM1038 N_VPWR_M1038_d N_SET_B_M1038_g N_A_1555_410#_M1038_s VPB PSHORT L=0.15
+ W=1 AD=0.269075 AS=0.295 PD=1.705 PS=2.59 NRD=42.158 NRS=1.9503 M=1 R=6.66667
+ SA=75000.2 SB=75001.2 A=0.15 P=2.3 MULT=1
MM1041 A_1931_392# N_A_975_322#_M1041_g N_VPWR_M1038_d VPB PSHORT L=0.15 W=1
+ AD=0.135 AS=0.269075 PD=1.27 PS=1.705 NRD=15.7403 NRS=42.158 M=1 R=6.66667
+ SA=75000.8 SB=75000.6 A=0.15 P=2.3 MULT=1
MM1009 N_A_1555_410#_M1009_d N_A_1335_112#_M1009_g A_1931_392# VPB PSHORT L=0.15
+ W=1 AD=0.28 AS=0.135 PD=2.56 PS=1.27 NRD=1.9503 NRS=15.7403 M=1 R=6.66667
+ SA=75001.3 SB=75000.2 A=0.15 P=2.3 MULT=1
MM1036 N_VPWR_M1036_d N_RESET_B_M1036_g N_A_975_322#_M1036_s VPB PSHORT L=0.15
+ W=0.64 AD=0.137018 AS=0.1792 PD=1.08727 PS=1.84 NRD=48.9545 NRS=3.0732 M=1
+ R=4.26667 SA=75000.2 SB=75001.2 A=0.096 P=1.58 MULT=1
MM1017 N_Q_N_M1017_d N_A_1555_410#_M1017_g N_VPWR_M1036_d VPB PSHORT L=0.15
+ W=1.12 AD=0.168 AS=0.239782 PD=1.42 PS=1.90273 NRD=1.7533 NRS=1.7533 M=1
+ R=7.46667 SA=75000.5 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1024 N_Q_N_M1017_d N_A_1555_410#_M1024_g N_VPWR_M1024_s VPB PSHORT L=0.15
+ W=1.12 AD=0.168 AS=0.3136 PD=1.42 PS=2.8 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001 SB=75000.2 A=0.168 P=2.54 MULT=1
MM1018 N_VPWR_M1018_d N_A_1555_410#_M1018_g N_A_2516_368#_M1018_s VPB PSHORT
+ L=0.15 W=1 AD=0.190377 AS=0.28 PD=1.40566 PS=2.56 NRD=15.7403 NRS=1.9503 M=1
+ R=6.66667 SA=75000.2 SB=75001.2 A=0.15 P=2.3 MULT=1
MM1019 N_Q_M1019_d N_A_2516_368#_M1019_g N_VPWR_M1018_d VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.213223 PD=1.42 PS=1.57434 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.7 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1025 N_Q_M1019_d N_A_2516_368#_M1025_g N_VPWR_M1025_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.3192 PD=1.42 PS=2.81 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.1 SB=75000.2 A=0.168 P=2.54 MULT=1
DX44_noxref VNB VPB NWDIODE A=27.4908 P=33.28
c_291 VPB 0 3.14884e-19 $X=0 $Y=3.085
*
.include "sky130_fd_sc_hs__dfbbn_2.pxi.spice"
*
.ends
*
*
