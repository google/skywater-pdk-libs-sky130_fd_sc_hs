* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hs__a2bb2oi_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
M1000 VPWR B1 a_424_368# VPB pshort w=1.12e+06u l=150000u
+  ad=9.47e+11p pd=8.23e+06u as=1.288e+12p ps=1.126e+07u
M1001 a_424_368# B1 VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1002 a_212_102# A2_N a_209_392# VPB pshort w=1e+06u l=150000u
+  ad=2.75e+11p pd=2.55e+06u as=2.4e+11p ps=2.48e+06u
M1003 Y B2 a_615_74# VNB nlowvt w=740000u l=150000u
+  ad=4.144e+11p pd=4.08e+06u as=5.994e+11p ps=6.06e+06u
M1004 Y a_212_102# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=8.17e+11p ps=8.02e+06u
M1005 a_615_74# B1 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_209_392# A1_N VPWR VPB pshort w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_615_74# B2 Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VGND A2_N a_212_102# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=2.08e+11p ps=1.93e+06u
M1009 Y a_212_102# a_424_368# VPB pshort w=1.12e+06u l=150000u
+  ad=3.36e+11p pd=2.84e+06u as=0p ps=0u
M1010 a_212_102# A1_N VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VGND a_212_102# Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_424_368# a_212_102# Y VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VPWR B2 a_424_368# VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 VGND B1 a_615_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_424_368# B2 VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
