* File: sky130_fd_sc_hs__o21bai_2.pex.spice
* Created: Thu Aug 27 20:58:54 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HS__O21BAI_2%B1_N 3 5 7 8 12
r33 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.625
+ $Y=1.515 $X2=0.625 $Y2=1.515
r34 8 12 4.60977 $w=3.73e-07 $l=1.5e-07 $layer=LI1_cond $X=0.647 $Y=1.665
+ $X2=0.647 $Y2=1.515
r35 5 11 50.9845 $w=3.31e-07 $l=2.93684e-07 $layer=POLY_cond $X=0.7 $Y=1.765
+ $X2=0.605 $Y2=1.515
r36 5 7 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=0.7 $Y=1.765 $X2=0.7
+ $Y2=2.34
r37 1 11 38.6069 $w=3.31e-07 $l=2.13014e-07 $layer=POLY_cond $X=0.495 $Y=1.35
+ $X2=0.605 $Y2=1.515
r38 1 3 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.495 $Y=1.35
+ $X2=0.495 $Y2=0.69
.ends

.subckt PM_SKY130_FD_SC_HS__O21BAI_2%A_27_74# 1 2 7 9 10 12 14 15 17 18 20 21 24
+ 28 34 36 40 43 45 46
c87 18 0 1.40781e-19 $X=1.92 $Y=1.765
r88 45 46 7.85017 $w=5.23e-07 $l=8.5e-08 $layer=LI1_cond $X=0.377 $Y=2.035
+ $X2=0.377 $Y2=1.95
r89 40 41 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.195
+ $Y=1.385 $X2=1.195 $Y2=1.385
r90 38 40 7.15912 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=1.195 $Y=1.18
+ $X2=1.195 $Y2=1.385
r91 37 43 2.11342 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.365 $Y=1.095
+ $X2=0.24 $Y2=1.095
r92 36 38 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.03 $Y=1.095
+ $X2=1.195 $Y2=1.18
r93 36 37 43.385 $w=1.68e-07 $l=6.65e-07 $layer=LI1_cond $X=1.03 $Y=1.095
+ $X2=0.365 $Y2=1.095
r94 32 45 4.03249 $w=5.23e-07 $l=1.77e-07 $layer=LI1_cond $X=0.377 $Y=2.212
+ $X2=0.377 $Y2=2.035
r95 32 34 11.4596 $w=5.23e-07 $l=5.03e-07 $layer=LI1_cond $X=0.377 $Y=2.212
+ $X2=0.377 $Y2=2.715
r96 30 43 4.3182 $w=2.1e-07 $l=1.03078e-07 $layer=LI1_cond $X=0.2 $Y=1.18
+ $X2=0.24 $Y2=1.095
r97 30 46 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=0.2 $Y=1.18 $X2=0.2
+ $Y2=1.95
r98 26 43 4.3182 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=0.24 $Y=1.01 $X2=0.24
+ $Y2=1.095
r99 26 28 22.8184 $w=2.48e-07 $l=4.95e-07 $layer=LI1_cond $X=0.24 $Y=1.01
+ $X2=0.24 $Y2=0.515
r100 23 24 56.3207 $w=3.68e-07 $l=4.3e-07 $layer=POLY_cond $X=1.485 $Y=1.492
+ $X2=1.915 $Y2=1.492
r101 22 23 1.96467 $w=3.68e-07 $l=1.5e-08 $layer=POLY_cond $X=1.47 $Y=1.492
+ $X2=1.485 $Y2=1.492
r102 21 41 32.3493 $w=3.3e-07 $l=1.85e-07 $layer=POLY_cond $X=1.38 $Y=1.385
+ $X2=1.195 $Y2=1.385
r103 21 22 12.4101 $w=3.68e-07 $l=1.45186e-07 $layer=POLY_cond $X=1.38 $Y=1.385
+ $X2=1.47 $Y2=1.492
r104 18 20 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.92 $Y=1.765
+ $X2=1.92 $Y2=2.4
r105 15 24 23.8357 $w=1.5e-07 $l=2.72e-07 $layer=POLY_cond $X=1.915 $Y=1.22
+ $X2=1.915 $Y2=1.492
r106 15 17 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.915 $Y=1.22
+ $X2=1.915 $Y2=0.74
r107 14 18 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=1.92 $Y=1.675
+ $X2=1.92 $Y2=1.765
r108 13 24 0.654891 $w=3.68e-07 $l=5e-09 $layer=POLY_cond $X=1.92 $Y=1.492
+ $X2=1.915 $Y2=1.492
r109 13 14 58.3064 $w=1.8e-07 $l=1.5e-07 $layer=POLY_cond $X=1.92 $Y=1.525
+ $X2=1.92 $Y2=1.675
r110 10 23 23.8357 $w=1.5e-07 $l=2.72e-07 $layer=POLY_cond $X=1.485 $Y=1.22
+ $X2=1.485 $Y2=1.492
r111 10 12 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.485 $Y=1.22
+ $X2=1.485 $Y2=0.74
r112 7 22 23.8357 $w=1.5e-07 $l=2.73e-07 $layer=POLY_cond $X=1.47 $Y=1.765
+ $X2=1.47 $Y2=1.492
r113 7 9 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.47 $Y=1.765
+ $X2=1.47 $Y2=2.4
r114 2 45 400 $w=1.7e-07 $l=2.61247e-07 $layer=licon1_PDIFF $count=1 $X=0.32
+ $Y=1.84 $X2=0.475 $Y2=2.035
r115 2 34 400 $w=1.7e-07 $l=9.49342e-07 $layer=licon1_PDIFF $count=1 $X=0.32
+ $Y=1.84 $X2=0.475 $Y2=2.715
r116 1 28 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__O21BAI_2%A1 3 5 7 10 12 14 17 20 21 23 29 32
c81 5 0 7.17547e-20 $X=2.46 $Y=1.765
c82 3 0 1.9405e-19 $X=2.415 $Y=0.74
r83 30 32 0.751593 $w=2.28e-07 $l=1.5e-08 $layer=LI1_cond $X=3.6 $Y=1.65 $X2=3.6
+ $Y2=1.665
r84 28 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.89
+ $Y=1.485 $X2=3.89 $Y2=1.485
r85 23 29 10.1275 $w=3.28e-07 $l=2.9e-07 $layer=LI1_cond $X=3.6 $Y=1.485
+ $X2=3.89 $Y2=1.485
r86 23 30 2.85155 $w=2.3e-07 $l=1.65e-07 $layer=LI1_cond $X=3.6 $Y=1.485 $X2=3.6
+ $Y2=1.65
r87 23 32 1.75372 $w=2.28e-07 $l=3.5e-08 $layer=LI1_cond $X=3.6 $Y=1.7 $X2=3.6
+ $Y2=1.665
r88 22 23 12.5266 $w=2.28e-07 $l=2.5e-07 $layer=LI1_cond $X=3.6 $Y=1.95 $X2=3.6
+ $Y2=1.7
r89 20 22 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=3.485 $Y=2.035
+ $X2=3.6 $Y2=1.95
r90 20 21 59.0428 $w=1.68e-07 $l=9.05e-07 $layer=LI1_cond $X=3.485 $Y=2.035
+ $X2=2.58 $Y2=2.035
r91 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.415
+ $Y=1.515 $X2=2.415 $Y2=1.515
r92 15 21 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.415 $Y=1.95
+ $X2=2.58 $Y2=2.035
r93 15 17 15.1913 $w=3.28e-07 $l=4.35e-07 $layer=LI1_cond $X=2.415 $Y=1.95
+ $X2=2.415 $Y2=1.515
r94 12 28 57.6553 $w=2.91e-07 $l=3.15278e-07 $layer=POLY_cond $X=3.815 $Y=1.765
+ $X2=3.89 $Y2=1.485
r95 12 14 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.815 $Y=1.765
+ $X2=3.815 $Y2=2.4
r96 8 28 38.6072 $w=2.91e-07 $l=2.03101e-07 $layer=POLY_cond $X=3.805 $Y=1.32
+ $X2=3.89 $Y2=1.485
r97 8 10 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=3.805 $Y=1.32
+ $X2=3.805 $Y2=0.74
r98 5 18 52.2586 $w=2.99e-07 $l=2.7157e-07 $layer=POLY_cond $X=2.46 $Y=1.765
+ $X2=2.415 $Y2=1.515
r99 5 7 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.46 $Y=1.765
+ $X2=2.46 $Y2=2.4
r100 1 18 38.5562 $w=2.99e-07 $l=1.65e-07 $layer=POLY_cond $X=2.415 $Y=1.35
+ $X2=2.415 $Y2=1.515
r101 1 3 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.415 $Y=1.35
+ $X2=2.415 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HS__O21BAI_2%A2 1 3 6 8 10 13 15 21 22
r59 22 23 1.9127 $w=3.78e-07 $l=1.5e-08 $layer=POLY_cond $X=3.36 $Y=1.557
+ $X2=3.375 $Y2=1.557
r60 20 22 42.0794 $w=3.78e-07 $l=3.3e-07 $layer=POLY_cond $X=3.03 $Y=1.557
+ $X2=3.36 $Y2=1.557
r61 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.03
+ $Y=1.515 $X2=3.03 $Y2=1.515
r62 18 20 10.8386 $w=3.78e-07 $l=8.5e-08 $layer=POLY_cond $X=2.945 $Y=1.557
+ $X2=3.03 $Y2=1.557
r63 17 18 4.46296 $w=3.78e-07 $l=3.5e-08 $layer=POLY_cond $X=2.91 $Y=1.557
+ $X2=2.945 $Y2=1.557
r64 15 21 4.16546 $w=4.13e-07 $l=1.5e-07 $layer=LI1_cond $X=3.027 $Y=1.665
+ $X2=3.027 $Y2=1.515
r65 11 23 24.4846 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.375 $Y=1.35
+ $X2=3.375 $Y2=1.557
r66 11 13 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=3.375 $Y=1.35
+ $X2=3.375 $Y2=0.74
r67 8 22 24.4846 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=3.36 $Y=1.765
+ $X2=3.36 $Y2=1.557
r68 8 10 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.36 $Y=1.765
+ $X2=3.36 $Y2=2.4
r69 4 18 24.4846 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.945 $Y=1.35
+ $X2=2.945 $Y2=1.557
r70 4 6 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.945 $Y=1.35
+ $X2=2.945 $Y2=0.74
r71 1 17 24.4846 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=2.91 $Y=1.765
+ $X2=2.91 $Y2=1.557
r72 1 3 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.91 $Y=1.765
+ $X2=2.91 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_HS__O21BAI_2%VPWR 1 2 3 12 18 20 22 26 28 33 38 47 50 54
r56 53 54 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r57 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r58 45 54 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.08 $Y2=3.33
r59 44 45 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r60 42 45 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.6 $Y2=3.33
r61 41 44 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=2.64 $Y=3.33 $X2=3.6
+ $Y2=3.33
r62 41 42 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r63 39 50 9.31531 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=2.35 $Y=3.33
+ $X2=2.165 $Y2=3.33
r64 39 41 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=2.35 $Y=3.33
+ $X2=2.64 $Y2=3.33
r65 38 53 4.01252 $w=1.7e-07 $l=1.82e-07 $layer=LI1_cond $X=3.955 $Y=3.33
+ $X2=4.137 $Y2=3.33
r66 38 44 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=3.955 $Y=3.33
+ $X2=3.6 $Y2=3.33
r67 37 48 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r68 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r69 34 47 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.335 $Y=3.33
+ $X2=1.17 $Y2=3.33
r70 34 36 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.335 $Y=3.33
+ $X2=1.68 $Y2=3.33
r71 33 50 9.31531 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=1.98 $Y=3.33
+ $X2=2.165 $Y2=3.33
r72 33 36 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=1.98 $Y=3.33 $X2=1.68
+ $Y2=3.33
r73 31 48 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r74 30 31 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r75 28 47 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.005 $Y=3.33
+ $X2=1.17 $Y2=3.33
r76 28 30 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=1.005 $Y=3.33
+ $X2=0.72 $Y2=3.33
r77 26 42 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r78 26 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.68 $Y2=3.33
r79 26 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r80 22 25 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=4.08 $Y=1.985
+ $X2=4.08 $Y2=2.815
r81 20 53 3.13065 $w=2.5e-07 $l=1.09864e-07 $layer=LI1_cond $X=4.08 $Y=3.245
+ $X2=4.137 $Y2=3.33
r82 20 25 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=4.08 $Y=3.245
+ $X2=4.08 $Y2=2.815
r83 16 50 1.24149 $w=3.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.165 $Y=3.245
+ $X2=2.165 $Y2=3.33
r84 16 18 13.3933 $w=3.68e-07 $l=4.3e-07 $layer=LI1_cond $X=2.165 $Y=3.245
+ $X2=2.165 $Y2=2.815
r85 12 15 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=1.17 $Y=1.985
+ $X2=1.17 $Y2=2.815
r86 10 47 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.17 $Y=3.245
+ $X2=1.17 $Y2=3.33
r87 10 15 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=1.17 $Y=3.245
+ $X2=1.17 $Y2=2.815
r88 3 25 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=3.89
+ $Y=1.84 $X2=4.04 $Y2=2.815
r89 3 22 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=3.89
+ $Y=1.84 $X2=4.04 $Y2=1.985
r90 2 18 600 $w=1.7e-07 $l=1.05659e-06 $layer=licon1_PDIFF $count=1 $X=1.995
+ $Y=1.84 $X2=2.165 $Y2=2.815
r91 1 15 400 $w=1.7e-07 $l=1.15575e-06 $layer=licon1_PDIFF $count=1 $X=0.775
+ $Y=1.84 $X2=1.17 $Y2=2.815
r92 1 12 400 $w=1.7e-07 $l=4.61844e-07 $layer=licon1_PDIFF $count=1 $X=0.775
+ $Y=1.84 $X2=1.17 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HS__O21BAI_2%Y 1 2 3 14 16 18 23 24 25 26 41
c46 14 0 1.9405e-19 $X=1.7 $Y=0.8
r47 31 41 1.78887 $w=3.33e-07 $l=5.2e-08 $layer=LI1_cond $X=1.697 $Y=1.347
+ $X2=1.697 $Y2=1.295
r48 25 26 11.0084 $w=3.33e-07 $l=3.2e-07 $layer=LI1_cond $X=1.697 $Y=1.665
+ $X2=1.697 $Y2=1.985
r49 24 41 0.584822 $w=3.33e-07 $l=1.7e-08 $layer=LI1_cond $X=1.697 $Y=1.278
+ $X2=1.697 $Y2=1.295
r50 24 39 4.13832 $w=3.33e-07 $l=9.8e-08 $layer=LI1_cond $X=1.697 $Y=1.278
+ $X2=1.697 $Y2=1.18
r51 24 25 10.3892 $w=3.33e-07 $l=3.02e-07 $layer=LI1_cond $X=1.697 $Y=1.363
+ $X2=1.697 $Y2=1.665
r52 24 31 0.550421 $w=3.33e-07 $l=1.6e-08 $layer=LI1_cond $X=1.697 $Y=1.363
+ $X2=1.697 $Y2=1.347
r53 21 26 10.4924 $w=3.33e-07 $l=3.05e-07 $layer=LI1_cond $X=1.697 $Y=2.29
+ $X2=1.697 $Y2=1.985
r54 21 23 3.22182 $w=2.92e-07 $l=8.5e-08 $layer=LI1_cond $X=1.697 $Y=2.29
+ $X2=1.697 $Y2=2.375
r55 18 20 3.58824 $w=1.7e-07 $l=5e-08 $layer=LI1_cond $X=3.135 $Y=2.46 $X2=3.135
+ $Y2=2.51
r56 17 23 3.35233 $w=1.7e-07 $l=1.68e-07 $layer=LI1_cond $X=1.865 $Y=2.375
+ $X2=1.697 $Y2=2.375
r57 16 18 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.05 $Y=2.375
+ $X2=3.135 $Y2=2.46
r58 16 17 77.3102 $w=1.68e-07 $l=1.185e-06 $layer=LI1_cond $X=3.05 $Y=2.375
+ $X2=1.865 $Y2=2.375
r59 14 39 17.5171 $w=2.48e-07 $l=3.8e-07 $layer=LI1_cond $X=1.74 $Y=0.8 $X2=1.74
+ $Y2=1.18
r60 3 20 600 $w=1.7e-07 $l=7.41215e-07 $layer=licon1_PDIFF $count=1 $X=2.985
+ $Y=1.84 $X2=3.135 $Y2=2.51
r61 2 26 600 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=1.545
+ $Y=1.84 $X2=1.695 $Y2=1.985
r62 2 23 300 $w=1.7e-07 $l=6.30555e-07 $layer=licon1_PDIFF $count=2 $X=1.545
+ $Y=1.84 $X2=1.695 $Y2=2.4
r63 1 14 182 $w=1.7e-07 $l=4.95076e-07 $layer=licon1_NDIFF $count=1 $X=1.56
+ $Y=0.37 $X2=1.7 $Y2=0.8
.ends

.subckt PM_SKY130_FD_SC_HS__O21BAI_2%A_507_368# 1 2 7 11 14
c31 14 0 1.40781e-19 $X=2.685 $Y=2.805
c32 7 0 7.17547e-20 $X=3.42 $Y=2.99
r33 14 16 6.46067 $w=3.28e-07 $l=1.85e-07 $layer=LI1_cond $X=2.685 $Y=2.805
+ $X2=2.685 $Y2=2.99
r34 9 11 18.2327 $w=3.33e-07 $l=5.3e-07 $layer=LI1_cond $X=3.587 $Y=2.905
+ $X2=3.587 $Y2=2.375
r35 8 16 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.85 $Y=2.99
+ $X2=2.685 $Y2=2.99
r36 7 9 7.80856 $w=1.7e-07 $l=2.05144e-07 $layer=LI1_cond $X=3.42 $Y=2.99
+ $X2=3.587 $Y2=2.905
r37 7 8 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=3.42 $Y=2.99 $X2=2.85
+ $Y2=2.99
r38 2 11 300 $w=1.7e-07 $l=6.05372e-07 $layer=licon1_PDIFF $count=2 $X=3.435
+ $Y=1.84 $X2=3.585 $Y2=2.375
r39 1 14 600 $w=1.7e-07 $l=1.03729e-06 $layer=licon1_PDIFF $count=1 $X=2.535
+ $Y=1.84 $X2=2.685 $Y2=2.805
.ends

.subckt PM_SKY130_FD_SC_HS__O21BAI_2%VGND 1 2 3 12 16 20 22 24 29 37 44 45 48 51
+ 54
r54 54 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r55 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r56 48 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r57 45 55 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=3.6
+ $Y2=0
r58 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r59 42 54 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.755 $Y=0 $X2=3.59
+ $Y2=0
r60 42 44 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=3.755 $Y=0 $X2=4.08
+ $Y2=0
r61 41 55 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=3.6
+ $Y2=0
r62 41 52 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=2.64
+ $Y2=0
r63 40 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r64 38 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.865 $Y=0 $X2=2.7
+ $Y2=0
r65 38 40 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=2.865 $Y=0 $X2=3.12
+ $Y2=0
r66 37 54 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.425 $Y=0 $X2=3.59
+ $Y2=0
r67 37 40 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=3.425 $Y=0 $X2=3.12
+ $Y2=0
r68 33 49 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r69 32 35 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r70 32 33 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r71 30 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.875 $Y=0 $X2=0.71
+ $Y2=0
r72 30 32 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.875 $Y=0 $X2=1.2
+ $Y2=0
r73 29 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.535 $Y=0 $X2=2.7
+ $Y2=0
r74 29 35 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=2.535 $Y=0 $X2=2.16
+ $Y2=0
r75 27 49 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r76 26 27 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r77 24 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.545 $Y=0 $X2=0.71
+ $Y2=0
r78 24 26 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.545 $Y=0 $X2=0.24
+ $Y2=0
r79 22 52 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r80 22 33 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.2
+ $Y2=0
r81 22 35 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r82 18 54 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.59 $Y=0.085
+ $X2=3.59 $Y2=0
r83 18 20 19.5566 $w=3.28e-07 $l=5.6e-07 $layer=LI1_cond $X=3.59 $Y=0.085
+ $X2=3.59 $Y2=0.645
r84 14 51 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.7 $Y=0.085 $X2=2.7
+ $Y2=0
r85 14 16 20.6043 $w=3.28e-07 $l=5.9e-07 $layer=LI1_cond $X=2.7 $Y=0.085 $X2=2.7
+ $Y2=0.675
r86 10 48 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.71 $Y=0.085
+ $X2=0.71 $Y2=0
r87 10 12 20.6043 $w=3.28e-07 $l=5.9e-07 $layer=LI1_cond $X=0.71 $Y=0.085
+ $X2=0.71 $Y2=0.675
r88 3 20 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=3.45
+ $Y=0.37 $X2=3.59 $Y2=0.645
r89 2 16 182 $w=1.7e-07 $l=3.96327e-07 $layer=licon1_NDIFF $count=1 $X=2.49
+ $Y=0.37 $X2=2.7 $Y2=0.675
r90 1 12 182 $w=1.7e-07 $l=3.68409e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.37 $X2=0.71 $Y2=0.675
.ends

.subckt PM_SKY130_FD_SC_HS__O21BAI_2%A_225_74# 1 2 3 4 15 17 18 22 23 24 27 29
+ 33 35
r64 31 33 21.4354 $w=2.48e-07 $l=4.65e-07 $layer=LI1_cond $X=4.06 $Y=0.98
+ $X2=4.06 $Y2=0.515
r65 30 35 5.16603 $w=1.7e-07 $l=9.21954e-08 $layer=LI1_cond $X=3.245 $Y=1.065
+ $X2=3.16 $Y2=1.08
r66 29 31 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=3.935 $Y=1.065
+ $X2=4.06 $Y2=0.98
r67 29 30 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=3.935 $Y=1.065
+ $X2=3.245 $Y2=1.065
r68 25 35 1.34256 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=3.16 $Y=0.98 $X2=3.16
+ $Y2=1.08
r69 25 27 30.3369 $w=1.68e-07 $l=4.65e-07 $layer=LI1_cond $X=3.16 $Y=0.98
+ $X2=3.16 $Y2=0.515
r70 23 35 5.16603 $w=1.7e-07 $l=9.21954e-08 $layer=LI1_cond $X=3.075 $Y=1.095
+ $X2=3.16 $Y2=1.08
r71 23 24 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=3.075 $Y=1.095
+ $X2=2.365 $Y2=1.095
r72 20 24 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.2 $Y=1.01
+ $X2=2.365 $Y2=1.095
r73 20 22 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=2.2 $Y=1.01 $X2=2.2
+ $Y2=0.515
r74 19 22 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=2.2 $Y=0.425 $X2=2.2
+ $Y2=0.515
r75 17 19 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.035 $Y=0.34
+ $X2=2.2 $Y2=0.425
r76 17 18 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=2.035 $Y=0.34
+ $X2=1.435 $Y2=0.34
r77 13 18 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.27 $Y=0.425
+ $X2=1.435 $Y2=0.34
r78 13 15 8.73063 $w=3.28e-07 $l=2.5e-07 $layer=LI1_cond $X=1.27 $Y=0.425
+ $X2=1.27 $Y2=0.675
r79 4 33 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.88
+ $Y=0.37 $X2=4.02 $Y2=0.515
r80 3 27 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.02
+ $Y=0.37 $X2=3.16 $Y2=0.515
r81 2 22 91 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=2 $X=1.99
+ $Y=0.37 $X2=2.2 $Y2=0.515
r82 1 15 182 $w=1.7e-07 $l=3.70473e-07 $layer=licon1_NDIFF $count=1 $X=1.125
+ $Y=0.37 $X2=1.27 $Y2=0.675
.ends

