* File: sky130_fd_sc_hs__a21bo_4.spice
* Created: Thu Aug 27 20:24:16 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hs__a21bo_4.pex.spice"
.subckt sky130_fd_sc_hs__a21bo_4  VNB VPB B1_N A1 A2 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A2	A2
* A1	A1
* B1_N	B1_N
* VPB	VPB
* VNB	VNB
MM1005 N_VGND_M1005_d N_B1_N_M1005_g N_A_29_392#_M1005_s VNB NLOWVT L=0.15
+ W=0.64 AD=0.149542 AS=0.1696 PD=1.10841 PS=1.81 NRD=15.468 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75005 A=0.096 P=1.58 MULT=1
MM1001 N_X_M1001_d N_A_187_338#_M1001_g N_VGND_M1005_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.172908 PD=1.02 PS=1.28159 NRD=0 NRS=12.972 M=1 R=4.93333
+ SA=75000.7 SB=75004.1 A=0.111 P=1.78 MULT=1
MM1003 N_X_M1001_d N_A_187_338#_M1003_g N_VGND_M1003_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.1
+ SB=75003.6 A=0.111 P=1.78 MULT=1
MM1008 N_X_M1008_d N_A_187_338#_M1008_g N_VGND_M1003_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.6
+ SB=75003.2 A=0.111 P=1.78 MULT=1
MM1010 N_X_M1008_d N_A_187_338#_M1010_g N_VGND_M1010_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.132302 PD=1.02 PS=1.17435 NRD=0 NRS=0 M=1 R=4.93333 SA=75002
+ SB=75002.8 A=0.111 P=1.78 MULT=1
MM1015 N_VGND_M1010_s N_A_29_392#_M1015_g N_A_187_338#_M1015_s VNB NLOWVT L=0.15
+ W=0.64 AD=0.114423 AS=0.0896 PD=1.01565 PS=0.92 NRD=11.244 NRS=0 M=1 R=4.26667
+ SA=75002.5 SB=75002.8 A=0.096 P=1.58 MULT=1
MM1021 N_VGND_M1021_d N_A_29_392#_M1021_g N_A_187_338#_M1015_s VNB NLOWVT L=0.15
+ W=0.64 AD=0.2016 AS=0.0896 PD=1.27 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75002.9 SB=75002.3 A=0.096 P=1.58 MULT=1
MM1009 N_VGND_M1021_d N_A2_M1009_g N_A_864_123#_M1009_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.2016 AS=0.1088 PD=1.27 PS=0.98 NRD=65.616 NRS=11.244 M=1 R=4.26667
+ SA=75003.7 SB=75001.5 A=0.096 P=1.58 MULT=1
MM1006 N_A_864_123#_M1009_s N_A1_M1006_g N_A_187_338#_M1006_s VNB NLOWVT L=0.15
+ W=0.64 AD=0.1088 AS=0.0896 PD=0.98 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75004.2 SB=75001.1 A=0.096 P=1.58 MULT=1
MM1012 N_A_864_123#_M1012_d N_A1_M1012_g N_A_187_338#_M1006_s VNB NLOWVT L=0.15
+ W=0.64 AD=0.0896 AS=0.0896 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75004.6 SB=75000.6 A=0.096 P=1.58 MULT=1
MM1020 N_VGND_M1020_d N_A2_M1020_g N_A_864_123#_M1012_d VNB NLOWVT L=0.15 W=0.64
+ AD=0.1696 AS=0.0896 PD=1.81 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667 SA=75005.1
+ SB=75000.2 A=0.096 P=1.58 MULT=1
MM1018 N_VPWR_M1018_d N_B1_N_M1018_g N_A_29_392#_M1018_s VPB PSHORT L=0.15 W=1
+ AD=0.187736 AS=0.275 PD=1.40094 PS=2.55 NRD=14.7553 NRS=1.9503 M=1 R=6.66667
+ SA=75000.2 SB=75002.1 A=0.15 P=2.3 MULT=1
MM1004 N_X_M1004_d N_A_187_338#_M1004_g N_VPWR_M1018_d VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.210264 PD=1.42 PS=1.56906 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.7 SB=75001.5 A=0.168 P=2.54 MULT=1
MM1007 N_X_M1004_d N_A_187_338#_M1007_g N_VPWR_M1007_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.1 SB=75001.1 A=0.168 P=2.54 MULT=1
MM1011 N_X_M1011_d N_A_187_338#_M1011_g N_VPWR_M1007_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.6 SB=75000.6 A=0.168 P=2.54 MULT=1
MM1013 N_X_M1011_d N_A_187_338#_M1013_g N_VPWR_M1013_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.308 PD=1.42 PS=2.79 NRD=1.7533 NRS=1.7533 M=1 R=7.46667 SA=75002
+ SB=75000.2 A=0.168 P=2.54 MULT=1
MM1014 N_A_187_338#_M1014_d N_A_29_392#_M1014_g N_A_596_392#_M1014_s VPB PSHORT
+ L=0.15 W=1 AD=0.15 AS=0.275 PD=1.3 PS=2.55 NRD=1.9503 NRS=1.9503 M=1 R=6.66667
+ SA=75000.2 SB=75002.4 A=0.15 P=2.3 MULT=1
MM1016 N_A_187_338#_M1014_d N_A_29_392#_M1016_g N_A_596_392#_M1016_s VPB PSHORT
+ L=0.15 W=1 AD=0.15 AS=0.15 PD=1.3 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=6.66667
+ SA=75000.6 SB=75002 A=0.15 P=2.3 MULT=1
MM1002 N_A_596_392#_M1016_s N_A2_M1002_g N_VPWR_M1002_s VPB PSHORT L=0.15 W=1
+ AD=0.15 AS=0.15 PD=1.3 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=6.66667 SA=75001.1
+ SB=75001.5 A=0.15 P=2.3 MULT=1
MM1000 N_VPWR_M1002_s N_A1_M1000_g N_A_596_392#_M1000_s VPB PSHORT L=0.15 W=1
+ AD=0.15 AS=0.15 PD=1.3 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=6.66667 SA=75001.5
+ SB=75001.1 A=0.15 P=2.3 MULT=1
MM1019 N_VPWR_M1019_d N_A1_M1019_g N_A_596_392#_M1000_s VPB PSHORT L=0.15 W=1
+ AD=0.15 AS=0.15 PD=1.3 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=6.66667 SA=75002
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1017 N_A_596_392#_M1017_d N_A2_M1017_g N_VPWR_M1019_d VPB PSHORT L=0.15 W=1
+ AD=0.275 AS=0.15 PD=2.55 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=6.66667 SA=75002.4
+ SB=75000.2 A=0.15 P=2.3 MULT=1
DX22_noxref VNB VPB NWDIODE A=12.3132 P=16.96
*
.include "sky130_fd_sc_hs__a21bo_4.pxi.spice"
*
.ends
*
*
