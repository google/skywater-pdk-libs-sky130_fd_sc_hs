# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_hs__sdlclkp_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__sdlclkp_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  9.600000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN GATE
    ANTENNAGATEAREA  0.208500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.835000 1.455000 1.315000 1.785000 ;
    END
  END GATE
  PIN GCLK
    ANTENNADIFFAREA  1.319400 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.705000 1.800000 8.985000 1.970000 ;
        RECT 7.705000 1.970000 8.035000 2.980000 ;
        RECT 7.865000 0.350000 8.115000 0.960000 ;
        RECT 7.865000 0.960000 9.055000 1.130000 ;
        RECT 8.655000 1.970000 8.985000 2.980000 ;
        RECT 8.725000 0.350000 9.055000 0.960000 ;
        RECT 8.725000 1.130000 9.055000 1.410000 ;
        RECT 8.725000 1.410000 8.985000 1.800000 ;
    END
  END GCLK
  PIN SCE
    ANTENNAGATEAREA  0.208500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.455000 0.550000 1.785000 ;
    END
  END SCE
  PIN CLK
    ANTENNAGATEAREA  0.516000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 5.785000 1.180000 6.115000 1.550000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 9.600000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 9.600000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 9.600000 0.085000 ;
      RECT 0.000000  3.245000 9.600000 3.415000 ;
      RECT 0.115000  0.085000 0.445000 1.285000 ;
      RECT 0.115000  1.955000 0.445000 3.245000 ;
      RECT 0.615000  0.615000 2.635000 0.785000 ;
      RECT 0.615000  0.785000 0.945000 1.285000 ;
      RECT 0.985000  1.955000 1.655000 2.310000 ;
      RECT 0.985000  2.310000 3.255000 2.480000 ;
      RECT 0.985000  2.480000 1.315000 2.835000 ;
      RECT 1.125000  0.085000 1.565000 0.445000 ;
      RECT 1.485000  0.785000 1.655000 1.955000 ;
      RECT 1.545000  2.650000 2.160000 3.245000 ;
      RECT 1.825000  0.955000 2.075000 1.565000 ;
      RECT 1.825000  1.565000 3.255000 1.735000 ;
      RECT 2.245000  1.065000 2.975000 1.235000 ;
      RECT 2.245000  1.235000 2.575000 1.395000 ;
      RECT 2.305000  0.350000 2.635000 0.615000 ;
      RECT 2.305000  0.785000 2.635000 0.895000 ;
      RECT 2.365000  1.735000 2.695000 2.140000 ;
      RECT 2.805000  0.270000 3.935000 0.440000 ;
      RECT 2.805000  0.440000 2.975000 1.065000 ;
      RECT 2.925000  1.405000 3.255000 1.565000 ;
      RECT 2.925000  1.905000 3.255000 2.310000 ;
      RECT 2.925000  2.480000 3.255000 2.755000 ;
      RECT 3.145000  0.610000 3.595000 0.940000 ;
      RECT 3.425000  0.940000 3.595000 1.235000 ;
      RECT 3.425000  1.235000 4.930000 1.405000 ;
      RECT 3.425000  1.405000 3.705000 2.755000 ;
      RECT 3.765000  0.440000 3.935000 0.895000 ;
      RECT 3.765000  0.895000 4.775000 1.065000 ;
      RECT 3.960000  1.575000 4.290000 1.735000 ;
      RECT 3.960000  1.735000 5.270000 1.905000 ;
      RECT 4.105000  0.085000 4.435000 0.725000 ;
      RECT 4.430000  2.075000 4.680000 3.245000 ;
      RECT 4.600000  1.405000 4.930000 1.565000 ;
      RECT 4.605000  0.255000 5.835000 0.425000 ;
      RECT 4.605000  0.425000 4.775000 0.895000 ;
      RECT 4.880000  1.905000 5.270000 2.240000 ;
      RECT 4.880000  2.240000 6.455000 2.410000 ;
      RECT 4.880000  2.410000 5.270000 2.895000 ;
      RECT 4.945000  0.595000 5.275000 1.065000 ;
      RECT 5.100000  1.065000 5.270000 1.735000 ;
      RECT 5.440000  1.820000 5.775000 2.070000 ;
      RECT 5.445000  0.425000 5.835000 1.010000 ;
      RECT 5.445000  1.010000 5.615000 1.820000 ;
      RECT 5.980000  2.580000 6.310000 3.245000 ;
      RECT 6.005000  0.085000 6.335000 1.010000 ;
      RECT 6.285000  1.300000 7.030000 1.630000 ;
      RECT 6.285000  1.630000 6.455000 2.240000 ;
      RECT 6.625000  1.800000 7.535000 1.970000 ;
      RECT 6.625000  1.970000 6.955000 2.980000 ;
      RECT 6.825000  0.350000 7.155000 0.960000 ;
      RECT 6.825000  0.960000 7.535000 1.130000 ;
      RECT 7.125000  2.140000 7.455000 3.245000 ;
      RECT 7.365000  1.130000 7.535000 1.300000 ;
      RECT 7.365000  1.300000 8.435000 1.630000 ;
      RECT 7.365000  1.630000 7.535000 1.800000 ;
      RECT 7.385000  0.085000 7.635000 0.790000 ;
      RECT 8.235000  2.140000 8.485000 3.245000 ;
      RECT 8.295000  0.085000 8.545000 0.790000 ;
      RECT 9.155000  1.820000 9.485000 3.245000 ;
      RECT 9.235000  0.085000 9.485000 1.130000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
      RECT 7.835000 -0.085000 8.005000 0.085000 ;
      RECT 7.835000  3.245000 8.005000 3.415000 ;
      RECT 8.315000 -0.085000 8.485000 0.085000 ;
      RECT 8.315000  3.245000 8.485000 3.415000 ;
      RECT 8.795000 -0.085000 8.965000 0.085000 ;
      RECT 8.795000  3.245000 8.965000 3.415000 ;
      RECT 9.275000 -0.085000 9.445000 0.085000 ;
      RECT 9.275000  3.245000 9.445000 3.415000 ;
  END
END sky130_fd_sc_hs__sdlclkp_4
END LIBRARY
