* File: sky130_fd_sc_hs__nor2_2.pex.spice
* Created: Tue Sep  1 20:10:50 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HS__NOR2_2%B 3 6 7 9 11 13 14 16 17
c40 17 0 6.90346e-20 $X=0.24 $Y=1.295
c41 9 0 1.88367e-19 $X=0.995 $Y=1.765
r42 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.28
+ $Y=1.385 $X2=0.28 $Y2=1.385
r43 17 21 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=0.28 $Y=1.295 $X2=0.28
+ $Y2=1.385
r44 15 16 30.3534 $w=1.85e-07 $l=7.5e-08 $layer=POLY_cond $X=0.547 $Y=1.69
+ $X2=0.547 $Y2=1.765
r45 13 20 30.6007 $w=3.3e-07 $l=1.75e-07 $layer=POLY_cond $X=0.455 $Y=1.385
+ $X2=0.28 $Y2=1.385
r46 13 15 112.674 $w=1.85e-07 $l=3.05e-07 $layer=POLY_cond $X=0.547 $Y=1.385
+ $X2=0.547 $Y2=1.69
r47 13 14 63.6015 $w=1.85e-07 $l=1.65e-07 $layer=POLY_cond $X=0.547 $Y=1.385
+ $X2=0.547 $Y2=1.22
r48 9 11 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.995 $Y=1.765
+ $X2=0.995 $Y2=2.4
r49 8 15 7.77431 $w=1.5e-07 $l=9.3e-08 $layer=POLY_cond $X=0.64 $Y=1.69
+ $X2=0.547 $Y2=1.69
r50 7 9 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.92 $Y=1.69
+ $X2=0.995 $Y2=1.765
r51 7 8 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=0.92 $Y=1.69 $X2=0.64
+ $Y2=1.69
r52 6 14 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=0.565 $Y=0.74
+ $X2=0.565 $Y2=1.22
r53 3 16 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.545 $Y=2.4
+ $X2=0.545 $Y2=1.765
.ends

.subckt PM_SKY130_FD_SC_HS__NOR2_2%A 1 3 4 5 6 8 9 11 12 13 14 20 26 28
c46 6 0 1.24794e-19 $X=1.445 $Y=1.765
c47 5 0 6.90346e-20 $X=1.07 $Y=1.26
r48 26 27 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.97
+ $Y=1.44 $X2=1.97 $Y2=1.44
r49 24 26 7.40779 $w=4.88e-07 $l=7.5e-08 $layer=POLY_cond $X=1.895 $Y=1.475
+ $X2=1.97 $Y2=1.475
r50 23 24 44.4467 $w=4.88e-07 $l=4.5e-07 $layer=POLY_cond $X=1.445 $Y=1.475
+ $X2=1.895 $Y2=1.475
r51 20 21 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.97
+ $Y=0.42 $X2=1.97 $Y2=0.42
r52 18 26 11.9614 $w=3.3e-07 $l=2.9e-07 $layer=POLY_cond $X=1.97 $Y=1.185
+ $X2=1.97 $Y2=1.475
r53 18 20 133.769 $w=3.3e-07 $l=7.65e-07 $layer=POLY_cond $X=1.97 $Y=1.185
+ $X2=1.97 $Y2=0.42
r54 14 27 4.35714 $w=4.06e-07 $l=1.45e-07 $layer=LI1_cond $X=2.04 $Y=1.295
+ $X2=2.04 $Y2=1.44
r55 14 29 3.37457 $w=4.7e-07 $l=1.2e-07 $layer=LI1_cond $X=2.04 $Y=1.295
+ $X2=2.04 $Y2=1.175
r56 13 29 6.36212 $w=4.68e-07 $l=2.5e-07 $layer=LI1_cond $X=2.04 $Y=0.925
+ $X2=2.04 $Y2=1.175
r57 13 28 6.36212 $w=4.68e-07 $l=2.5e-07 $layer=LI1_cond $X=2.04 $Y=0.925
+ $X2=2.04 $Y2=0.675
r58 12 28 3.36005 $w=4.7e-07 $l=1.2e-07 $layer=LI1_cond $X=2.04 $Y=0.555
+ $X2=2.04 $Y2=0.675
r59 12 21 4.03676 $w=4.08e-07 $l=1.35e-07 $layer=LI1_cond $X=2.04 $Y=0.555
+ $X2=2.04 $Y2=0.42
r60 9 24 30.7954 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=1.895 $Y=1.765
+ $X2=1.895 $Y2=1.475
r61 9 11 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.895 $Y=1.765
+ $X2=1.895 $Y2=2.4
r62 6 23 30.7954 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=1.445 $Y=1.765
+ $X2=1.445 $Y2=1.475
r63 6 8 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.445 $Y=1.765
+ $X2=1.445 $Y2=2.4
r64 4 23 34.2102 $w=4.88e-07 $l=2.56076e-07 $layer=POLY_cond $X=1.355 $Y=1.26
+ $X2=1.445 $Y2=1.475
r65 4 5 146.138 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=1.355 $Y=1.26
+ $X2=1.07 $Y2=1.26
r66 1 5 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.995 $Y=1.185
+ $X2=1.07 $Y2=1.26
r67 1 3 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=0.995 $Y=1.185
+ $X2=0.995 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HS__NOR2_2%A_35_368# 1 2 3 12 16 17 21 24 25 28
r41 28 30 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=2.12 $Y=1.985
+ $X2=2.12 $Y2=2.815
r42 26 28 1.3969 $w=3.28e-07 $l=4e-08 $layer=LI1_cond $X=2.12 $Y=1.945 $X2=2.12
+ $Y2=1.985
r43 24 26 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.955 $Y=1.86
+ $X2=2.12 $Y2=1.945
r44 24 25 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=1.955 $Y=1.86
+ $X2=1.305 $Y2=1.86
r45 21 23 54.1497 $w=1.68e-07 $l=8.3e-07 $layer=LI1_cond $X=1.22 $Y=1.985
+ $X2=1.22 $Y2=2.815
r46 19 23 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=1.22 $Y=2.905 $X2=1.22
+ $Y2=2.815
r47 18 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.22 $Y=1.945
+ $X2=1.305 $Y2=1.86
r48 18 21 2.60963 $w=1.68e-07 $l=4e-08 $layer=LI1_cond $X=1.22 $Y=1.945 $X2=1.22
+ $Y2=1.985
r49 16 19 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.135 $Y=2.99
+ $X2=1.22 $Y2=2.905
r50 16 17 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=1.135 $Y=2.99
+ $X2=0.405 $Y2=2.99
r51 12 15 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=0.28 $Y=1.985
+ $X2=0.28 $Y2=2.815
r52 10 17 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.28 $Y=2.905
+ $X2=0.405 $Y2=2.99
r53 10 15 4.14879 $w=2.48e-07 $l=9e-08 $layer=LI1_cond $X=0.28 $Y=2.905 $X2=0.28
+ $Y2=2.815
r54 3 30 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=1.97
+ $Y=1.84 $X2=2.12 $Y2=2.815
r55 3 28 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=1.97
+ $Y=1.84 $X2=2.12 $Y2=1.985
r56 2 23 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=1.07
+ $Y=1.84 $X2=1.22 $Y2=2.815
r57 2 21 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=1.07
+ $Y=1.84 $X2=1.22 $Y2=1.985
r58 1 15 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=0.175
+ $Y=1.84 $X2=0.32 $Y2=2.815
r59 1 12 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.175
+ $Y=1.84 $X2=0.32 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HS__NOR2_2%Y 1 2 9 11 12 18
c23 9 0 1.24794e-19 $X=0.78 $Y=0.515
r24 16 18 1.52529 $w=3.38e-07 $l=4.5e-08 $layer=LI1_cond $X=0.775 $Y=1.99
+ $X2=0.775 $Y2=2.035
r25 11 16 0.677908 $w=3.38e-07 $l=2e-08 $layer=LI1_cond $X=0.775 $Y=1.97
+ $X2=0.775 $Y2=1.99
r26 11 24 5.08431 $w=3.38e-07 $l=1.5e-07 $layer=LI1_cond $X=0.775 $Y=1.97
+ $X2=0.775 $Y2=1.82
r27 11 12 11.8634 $w=3.38e-07 $l=3.5e-07 $layer=LI1_cond $X=0.775 $Y=2.055
+ $X2=0.775 $Y2=2.405
r28 11 18 0.677908 $w=3.38e-07 $l=2e-08 $layer=LI1_cond $X=0.775 $Y=2.055
+ $X2=0.775 $Y2=2.035
r29 9 24 45.5739 $w=3.28e-07 $l=1.305e-06 $layer=LI1_cond $X=0.78 $Y=0.515
+ $X2=0.78 $Y2=1.82
r30 2 11 300 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=2 $X=0.62
+ $Y=1.84 $X2=0.77 $Y2=1.985
r31 1 9 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=0.64
+ $Y=0.37 $X2=0.78 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__NOR2_2%VPWR 1 6 9 10 11 21 22
c27 6 0 1.88367e-19 $X=1.67 $Y=2.28
r28 21 22 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r29 14 18 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.24 $Y=3.33 $X2=1.2
+ $Y2=3.33
r30 14 15 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r31 11 22 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.16 $Y2=3.33
r32 11 15 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.24 $Y2=3.33
r33 11 18 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r34 9 18 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.505 $Y=3.33
+ $X2=1.2 $Y2=3.33
r35 9 10 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.505 $Y=3.33
+ $X2=1.63 $Y2=3.33
r36 8 21 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=1.755 $Y=3.33
+ $X2=2.16 $Y2=3.33
r37 8 10 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.755 $Y=3.33
+ $X2=1.63 $Y2=3.33
r38 4 10 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.63 $Y=3.245
+ $X2=1.63 $Y2=3.33
r39 4 6 44.4843 $w=2.48e-07 $l=9.65e-07 $layer=LI1_cond $X=1.63 $Y=3.245
+ $X2=1.63 $Y2=2.28
r40 1 6 300 $w=1.7e-07 $l=5.0951e-07 $layer=licon1_PDIFF $count=2 $X=1.52
+ $Y=1.84 $X2=1.67 $Y2=2.28
.ends

.subckt PM_SKY130_FD_SC_HS__NOR2_2%VGND 1 2 7 9 13 15 17 24 25 31
r28 28 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r29 24 25 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r30 22 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.445 $Y=0 $X2=1.28
+ $Y2=0
r31 22 24 46.6471 $w=1.68e-07 $l=7.15e-07 $layer=LI1_cond $X=1.445 $Y=0 $X2=2.16
+ $Y2=0
r32 21 29 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r33 20 21 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r34 18 28 4.73185 $w=1.7e-07 $l=2.23e-07 $layer=LI1_cond $X=0.445 $Y=0 $X2=0.222
+ $Y2=0
r35 18 20 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=0.445 $Y=0 $X2=0.72
+ $Y2=0
r36 17 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.115 $Y=0 $X2=1.28
+ $Y2=0
r37 17 20 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=1.115 $Y=0 $X2=0.72
+ $Y2=0
r38 15 25 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r39 15 21 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r40 15 31 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r41 11 31 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.28 $Y=0.085
+ $X2=1.28 $Y2=0
r42 11 13 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=1.28 $Y=0.085
+ $X2=1.28 $Y2=0.515
r43 7 28 3.03433 $w=3.3e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.28 $Y=0.085
+ $X2=0.222 $Y2=0
r44 7 9 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=0.28 $Y=0.085 $X2=0.28
+ $Y2=0.515
r45 2 13 91 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=2 $X=1.07
+ $Y=0.37 $X2=1.28 $Y2=0.515
r46 1 9 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.515
.ends

