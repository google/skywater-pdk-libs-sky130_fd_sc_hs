* File: sky130_fd_sc_hs__a21oi_2.pxi.spice
* Created: Thu Aug 27 20:25:18 2020
* 
x_PM_SKY130_FD_SC_HS__A21OI_2%B1 N_B1_M1010_g N_B1_c_70_n N_B1_c_76_n
+ N_B1_M1007_g N_B1_c_71_n N_B1_c_78_n N_B1_M1008_g N_B1_c_72_n B1 N_B1_c_74_n
+ PM_SKY130_FD_SC_HS__A21OI_2%B1
x_PM_SKY130_FD_SC_HS__A21OI_2%A2 N_A2_c_114_n N_A2_M1002_g N_A2_c_118_n
+ N_A2_M1001_g N_A2_c_119_n N_A2_M1009_g N_A2_M1004_g A2 A2 N_A2_c_117_n
+ PM_SKY130_FD_SC_HS__A21OI_2%A2
x_PM_SKY130_FD_SC_HS__A21OI_2%A1 N_A1_c_174_n N_A1_M1003_g N_A1_M1000_g
+ N_A1_M1006_g N_A1_c_175_n N_A1_M1005_g A1 N_A1_c_172_n N_A1_c_173_n
+ PM_SKY130_FD_SC_HS__A21OI_2%A1
x_PM_SKY130_FD_SC_HS__A21OI_2%A_131_368# N_A_131_368#_M1007_s
+ N_A_131_368#_M1008_s N_A_131_368#_M1009_d N_A_131_368#_M1005_s
+ N_A_131_368#_c_220_n N_A_131_368#_c_221_n N_A_131_368#_c_222_n
+ N_A_131_368#_c_229_n N_A_131_368#_c_230_n N_A_131_368#_c_232_n
+ N_A_131_368#_c_236_n N_A_131_368#_c_223_n N_A_131_368#_c_224_n
+ PM_SKY130_FD_SC_HS__A21OI_2%A_131_368#
x_PM_SKY130_FD_SC_HS__A21OI_2%Y N_Y_M1010_d N_Y_M1000_s N_Y_M1007_d N_Y_c_273_n
+ N_Y_c_274_n N_Y_c_275_n N_Y_c_276_n N_Y_c_280_n N_Y_c_277_n N_Y_c_278_n Y Y
+ PM_SKY130_FD_SC_HS__A21OI_2%Y
x_PM_SKY130_FD_SC_HS__A21OI_2%VPWR N_VPWR_M1001_s N_VPWR_M1003_d N_VPWR_c_330_n
+ N_VPWR_c_331_n N_VPWR_c_332_n N_VPWR_c_333_n VPWR N_VPWR_c_334_n
+ N_VPWR_c_335_n N_VPWR_c_329_n N_VPWR_c_337_n PM_SKY130_FD_SC_HS__A21OI_2%VPWR
x_PM_SKY130_FD_SC_HS__A21OI_2%VGND N_VGND_M1010_s N_VGND_M1002_s N_VGND_c_373_n
+ N_VGND_c_374_n N_VGND_c_375_n VGND N_VGND_c_376_n N_VGND_c_377_n
+ N_VGND_c_378_n N_VGND_c_379_n PM_SKY130_FD_SC_HS__A21OI_2%VGND
x_PM_SKY130_FD_SC_HS__A21OI_2%A_280_107# N_A_280_107#_M1002_d
+ N_A_280_107#_M1004_d N_A_280_107#_M1006_d N_A_280_107#_c_410_n
+ N_A_280_107#_c_411_n N_A_280_107#_c_418_n N_A_280_107#_c_458_n
+ N_A_280_107#_c_412_n N_A_280_107#_c_413_n N_A_280_107#_c_414_n
+ N_A_280_107#_c_415_n N_A_280_107#_c_416_n
+ PM_SKY130_FD_SC_HS__A21OI_2%A_280_107#
cc_1 VNB N_B1_M1010_g 0.0431358f $X=-0.19 $Y=-0.245 $X2=0.48 $Y2=0.74
cc_2 VNB N_B1_c_70_n 0.0133105f $X=-0.19 $Y=-0.245 $X2=0.93 $Y2=1.69
cc_3 VNB N_B1_c_71_n 0.0164254f $X=-0.19 $Y=-0.245 $X2=1.38 $Y2=1.69
cc_4 VNB N_B1_c_72_n 0.00499721f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=1.69
cc_5 VNB B1 0.00347618f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_6 VNB N_B1_c_74_n 0.035519f $X=-0.19 $Y=-0.245 $X2=0.555 $Y2=1.6
cc_7 VNB N_A2_c_114_n 0.0207904f $X=-0.19 $Y=-0.245 $X2=0.48 $Y2=1.435
cc_8 VNB N_A2_M1004_g 0.0247974f $X=-0.19 $Y=-0.245 $X2=1.455 $Y2=1.765
cc_9 VNB A2 0.00987786f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_10 VNB N_A2_c_117_n 0.0503242f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A1_M1000_g 0.0238491f $X=-0.19 $Y=-0.245 $X2=0.555 $Y2=1.69
cc_12 VNB N_A1_M1006_g 0.0278198f $X=-0.19 $Y=-0.245 $X2=1.38 $Y2=1.69
cc_13 VNB N_A1_c_172_n 0.00102029f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A1_c_173_n 0.0380232f $X=-0.19 $Y=-0.245 $X2=0.48 $Y2=1.6
cc_15 VNB N_Y_c_273_n 0.017421f $X=-0.19 $Y=-0.245 $X2=1.455 $Y2=1.765
cc_16 VNB N_Y_c_274_n 0.026508f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=1.69
cc_17 VNB N_Y_c_275_n 0.0173725f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_18 VNB N_Y_c_276_n 0.00925586f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.6
cc_19 VNB N_Y_c_277_n 2.51509e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_Y_c_278_n 0.00349834f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_VPWR_c_329_n 0.163682f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_VGND_c_373_n 0.0115487f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=1.765
cc_23 VNB N_VGND_c_374_n 0.0420835f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=2.4
cc_24 VNB N_VGND_c_375_n 0.0159289f $X=-0.19 $Y=-0.245 $X2=1.455 $Y2=2.4
cc_25 VNB N_VGND_c_376_n 0.043727f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_VGND_c_377_n 0.0399389f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_VGND_c_378_n 0.235811f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_379_n 0.00632082f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_280_107#_c_410_n 0.00342239f $X=-0.19 $Y=-0.245 $X2=1.38 $Y2=1.69
cc_30 VNB N_A_280_107#_c_411_n 0.0100707f $X=-0.19 $Y=-0.245 $X2=1.08 $Y2=1.69
cc_31 VNB N_A_280_107#_c_412_n 0.00456651f $X=-0.19 $Y=-0.245 $X2=1.455 $Y2=2.4
cc_32 VNB N_A_280_107#_c_413_n 0.0132061f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.6
cc_33 VNB N_A_280_107#_c_414_n 0.0148263f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.6
cc_34 VNB N_A_280_107#_c_415_n 0.0249441f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_280_107#_c_416_n 0.0113698f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VPB N_B1_c_70_n 0.0157429f $X=-0.19 $Y=1.66 $X2=0.93 $Y2=1.69
cc_37 VPB N_B1_c_76_n 0.018382f $X=-0.19 $Y=1.66 $X2=1.005 $Y2=1.765
cc_38 VPB N_B1_c_71_n 0.0113288f $X=-0.19 $Y=1.66 $X2=1.38 $Y2=1.69
cc_39 VPB N_B1_c_78_n 0.0145507f $X=-0.19 $Y=1.66 $X2=1.455 $Y2=1.765
cc_40 VPB N_B1_c_72_n 0.00167153f $X=-0.19 $Y=1.66 $X2=1.005 $Y2=1.69
cc_41 VPB B1 0.0129596f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_42 VPB N_B1_c_74_n 0.0268817f $X=-0.19 $Y=1.66 $X2=0.555 $Y2=1.6
cc_43 VPB N_A2_c_118_n 0.0157721f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_44 VPB N_A2_c_119_n 0.0162344f $X=-0.19 $Y=1.66 $X2=1.005 $Y2=1.765
cc_45 VPB A2 0.0067772f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_46 VPB N_A2_c_117_n 0.0236526f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_47 VPB N_A1_c_174_n 0.0159044f $X=-0.19 $Y=1.66 $X2=0.48 $Y2=1.435
cc_48 VPB N_A1_c_175_n 0.0192141f $X=-0.19 $Y=1.66 $X2=1.455 $Y2=1.765
cc_49 VPB N_A1_c_172_n 0.00283601f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_50 VPB N_A1_c_173_n 0.0206495f $X=-0.19 $Y=1.66 $X2=0.48 $Y2=1.6
cc_51 VPB N_A_131_368#_c_220_n 0.0364628f $X=-0.19 $Y=1.66 $X2=1.005 $Y2=1.69
cc_52 VPB N_A_131_368#_c_221_n 0.00454203f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.6
cc_53 VPB N_A_131_368#_c_222_n 0.00961757f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.6
cc_54 VPB N_A_131_368#_c_223_n 0.00257417f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_55 VPB N_A_131_368#_c_224_n 0.030827f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_56 VPB N_Y_c_276_n 0.005226f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.6
cc_57 VPB N_Y_c_280_n 7.3738e-19 $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.6
cc_58 VPB N_VPWR_c_330_n 0.00864185f $X=-0.19 $Y=1.66 $X2=1.005 $Y2=2.4
cc_59 VPB N_VPWR_c_331_n 0.00799266f $X=-0.19 $Y=1.66 $X2=1.455 $Y2=2.4
cc_60 VPB N_VPWR_c_332_n 0.0196495f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_61 VPB N_VPWR_c_333_n 0.00324402f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_62 VPB N_VPWR_c_334_n 0.0552656f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.6
cc_63 VPB N_VPWR_c_335_n 0.0207426f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_64 VPB N_VPWR_c_329_n 0.0877938f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_65 VPB N_VPWR_c_337_n 0.00497514f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_66 VPB N_A_280_107#_c_411_n 0.00325045f $X=-0.19 $Y=1.66 $X2=1.08 $Y2=1.69
cc_67 VPB N_A_280_107#_c_418_n 0.00730579f $X=-0.19 $Y=1.66 $X2=1.455 $Y2=1.765
cc_68 VPB N_A_280_107#_c_415_n 0.0122533f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_69 N_B1_c_78_n N_A2_c_118_n 0.0233621f $X=1.455 $Y=1.765 $X2=0 $Y2=0
cc_70 N_B1_c_71_n N_A2_c_117_n 0.00660562f $X=1.38 $Y=1.69 $X2=0 $Y2=0
cc_71 N_B1_c_70_n N_A_131_368#_c_220_n 0.00207738f $X=0.93 $Y=1.69 $X2=0 $Y2=0
cc_72 N_B1_c_76_n N_A_131_368#_c_221_n 0.0137046f $X=1.005 $Y=1.765 $X2=0 $Y2=0
cc_73 N_B1_c_78_n N_A_131_368#_c_221_n 0.0127563f $X=1.455 $Y=1.765 $X2=0 $Y2=0
cc_74 N_B1_M1010_g N_Y_c_273_n 0.0012158f $X=0.48 $Y=0.74 $X2=0 $Y2=0
cc_75 N_B1_M1010_g N_Y_c_274_n 0.0161196f $X=0.48 $Y=0.74 $X2=0 $Y2=0
cc_76 N_B1_c_70_n N_Y_c_274_n 0.00210831f $X=0.93 $Y=1.69 $X2=0 $Y2=0
cc_77 B1 N_Y_c_274_n 0.00891653f $X=0.155 $Y=1.58 $X2=0 $Y2=0
cc_78 N_B1_c_70_n N_Y_c_275_n 0.0022675f $X=0.93 $Y=1.69 $X2=0 $Y2=0
cc_79 N_B1_c_70_n N_Y_c_276_n 0.0162692f $X=0.93 $Y=1.69 $X2=0 $Y2=0
cc_80 N_B1_c_76_n N_Y_c_276_n 0.00688828f $X=1.005 $Y=1.765 $X2=0 $Y2=0
cc_81 N_B1_c_71_n N_Y_c_276_n 0.0122004f $X=1.38 $Y=1.69 $X2=0 $Y2=0
cc_82 N_B1_c_78_n N_Y_c_276_n 3.15021e-19 $X=1.455 $Y=1.765 $X2=0 $Y2=0
cc_83 N_B1_c_72_n N_Y_c_276_n 0.00442527f $X=1.005 $Y=1.69 $X2=0 $Y2=0
cc_84 B1 N_Y_c_276_n 0.0186087f $X=0.155 $Y=1.58 $X2=0 $Y2=0
cc_85 N_B1_c_74_n N_Y_c_276_n 0.0018352f $X=0.555 $Y=1.6 $X2=0 $Y2=0
cc_86 N_B1_c_76_n N_Y_c_280_n 0.0160332f $X=1.005 $Y=1.765 $X2=0 $Y2=0
cc_87 N_B1_c_71_n N_Y_c_280_n 0.00197838f $X=1.38 $Y=1.69 $X2=0 $Y2=0
cc_88 N_B1_c_78_n N_Y_c_280_n 0.0114063f $X=1.455 $Y=1.765 $X2=0 $Y2=0
cc_89 N_B1_c_76_n N_VPWR_c_334_n 0.00278271f $X=1.005 $Y=1.765 $X2=0 $Y2=0
cc_90 N_B1_c_78_n N_VPWR_c_334_n 0.00278271f $X=1.455 $Y=1.765 $X2=0 $Y2=0
cc_91 N_B1_c_76_n N_VPWR_c_329_n 0.00358624f $X=1.005 $Y=1.765 $X2=0 $Y2=0
cc_92 N_B1_c_78_n N_VPWR_c_329_n 0.00353907f $X=1.455 $Y=1.765 $X2=0 $Y2=0
cc_93 N_B1_M1010_g N_VGND_c_374_n 0.0182521f $X=0.48 $Y=0.74 $X2=0 $Y2=0
cc_94 B1 N_VGND_c_374_n 0.0176252f $X=0.155 $Y=1.58 $X2=0 $Y2=0
cc_95 N_B1_c_74_n N_VGND_c_374_n 0.00220195f $X=0.555 $Y=1.6 $X2=0 $Y2=0
cc_96 N_B1_M1010_g N_VGND_c_376_n 0.00383152f $X=0.48 $Y=0.74 $X2=0 $Y2=0
cc_97 N_B1_M1010_g N_VGND_c_378_n 0.00762539f $X=0.48 $Y=0.74 $X2=0 $Y2=0
cc_98 N_B1_c_71_n N_A_280_107#_c_410_n 0.00521306f $X=1.38 $Y=1.69 $X2=0 $Y2=0
cc_99 N_B1_c_71_n N_A_280_107#_c_411_n 0.00140999f $X=1.38 $Y=1.69 $X2=0 $Y2=0
cc_100 N_B1_c_78_n N_A_280_107#_c_411_n 0.00110062f $X=1.455 $Y=1.765 $X2=0
+ $Y2=0
cc_101 N_A2_c_119_n N_A1_c_174_n 0.027449f $X=2.415 $Y=1.765 $X2=-0.19
+ $Y2=-0.245
cc_102 N_A2_M1004_g N_A1_M1000_g 0.035579f $X=2.45 $Y=0.74 $X2=0 $Y2=0
cc_103 A2 N_A1_M1000_g 0.00536167f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_104 A2 N_A1_c_172_n 0.0277147f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_105 N_A2_c_117_n N_A1_c_172_n 2.21765e-19 $X=2.415 $Y=1.557 $X2=0 $Y2=0
cc_106 A2 N_A1_c_173_n 0.00443437f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_107 N_A2_c_117_n N_A1_c_173_n 0.0250278f $X=2.415 $Y=1.557 $X2=0 $Y2=0
cc_108 N_A2_c_118_n N_A_131_368#_c_221_n 0.00324431f $X=1.905 $Y=1.765 $X2=0
+ $Y2=0
cc_109 N_A2_c_118_n N_A_131_368#_c_229_n 4.27055e-19 $X=1.905 $Y=1.765 $X2=0
+ $Y2=0
cc_110 N_A2_c_118_n N_A_131_368#_c_230_n 0.00598174f $X=1.905 $Y=1.765 $X2=0
+ $Y2=0
cc_111 N_A2_c_119_n N_A_131_368#_c_230_n 5.89453e-19 $X=2.415 $Y=1.765 $X2=0
+ $Y2=0
cc_112 N_A2_c_118_n N_A_131_368#_c_232_n 0.0121197f $X=1.905 $Y=1.765 $X2=0
+ $Y2=0
cc_113 N_A2_c_119_n N_A_131_368#_c_232_n 0.0121197f $X=2.415 $Y=1.765 $X2=0
+ $Y2=0
cc_114 N_A2_c_118_n N_A_131_368#_c_223_n 5.49142e-19 $X=1.905 $Y=1.765 $X2=0
+ $Y2=0
cc_115 N_A2_c_119_n N_A_131_368#_c_223_n 0.00730009f $X=2.415 $Y=1.765 $X2=0
+ $Y2=0
cc_116 N_A2_c_114_n N_Y_c_275_n 0.0179555f $X=1.8 $Y=1.35 $X2=0 $Y2=0
cc_117 N_A2_M1004_g N_Y_c_275_n 0.0134085f $X=2.45 $Y=0.74 $X2=0 $Y2=0
cc_118 A2 N_Y_c_275_n 0.0385111f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_119 N_A2_c_117_n N_Y_c_275_n 0.00344153f $X=2.415 $Y=1.557 $X2=0 $Y2=0
cc_120 N_A2_c_118_n N_Y_c_280_n 9.09552e-19 $X=1.905 $Y=1.765 $X2=0 $Y2=0
cc_121 N_A2_M1004_g N_Y_c_278_n 0.0011095f $X=2.45 $Y=0.74 $X2=0 $Y2=0
cc_122 N_A2_c_118_n N_VPWR_c_330_n 0.00250897f $X=1.905 $Y=1.765 $X2=0 $Y2=0
cc_123 N_A2_c_119_n N_VPWR_c_330_n 0.00498232f $X=2.415 $Y=1.765 $X2=0 $Y2=0
cc_124 N_A2_c_119_n N_VPWR_c_332_n 0.00445602f $X=2.415 $Y=1.765 $X2=0 $Y2=0
cc_125 N_A2_c_118_n N_VPWR_c_334_n 0.0044313f $X=1.905 $Y=1.765 $X2=0 $Y2=0
cc_126 N_A2_c_118_n N_VPWR_c_329_n 0.00853993f $X=1.905 $Y=1.765 $X2=0 $Y2=0
cc_127 N_A2_c_119_n N_VPWR_c_329_n 0.00857549f $X=2.415 $Y=1.765 $X2=0 $Y2=0
cc_128 A2 N_VGND_M1002_s 0.00205137f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_129 N_A2_c_114_n N_VGND_c_375_n 0.00475861f $X=1.8 $Y=1.35 $X2=0 $Y2=0
cc_130 N_A2_M1004_g N_VGND_c_375_n 0.00661466f $X=2.45 $Y=0.74 $X2=0 $Y2=0
cc_131 N_A2_c_114_n N_VGND_c_376_n 0.003666f $X=1.8 $Y=1.35 $X2=0 $Y2=0
cc_132 N_A2_M1004_g N_VGND_c_377_n 0.00329872f $X=2.45 $Y=0.74 $X2=0 $Y2=0
cc_133 N_A2_c_114_n N_VGND_c_378_n 0.00495025f $X=1.8 $Y=1.35 $X2=0 $Y2=0
cc_134 N_A2_M1004_g N_VGND_c_378_n 0.00431825f $X=2.45 $Y=0.74 $X2=0 $Y2=0
cc_135 N_A2_c_114_n N_A_280_107#_c_410_n 0.00768497f $X=1.8 $Y=1.35 $X2=0 $Y2=0
cc_136 N_A2_M1004_g N_A_280_107#_c_410_n 4.66537e-19 $X=2.45 $Y=0.74 $X2=0 $Y2=0
cc_137 A2 N_A_280_107#_c_410_n 0.00461694f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_138 N_A2_c_114_n N_A_280_107#_c_411_n 0.0030154f $X=1.8 $Y=1.35 $X2=0 $Y2=0
cc_139 N_A2_c_118_n N_A_280_107#_c_411_n 0.00212266f $X=1.905 $Y=1.765 $X2=0
+ $Y2=0
cc_140 A2 N_A_280_107#_c_411_n 0.0297027f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_141 N_A2_c_117_n N_A_280_107#_c_411_n 0.0122944f $X=2.415 $Y=1.557 $X2=0
+ $Y2=0
cc_142 N_A2_c_118_n N_A_280_107#_c_418_n 0.0152108f $X=1.905 $Y=1.765 $X2=0
+ $Y2=0
cc_143 N_A2_c_119_n N_A_280_107#_c_418_n 0.0110045f $X=2.415 $Y=1.765 $X2=0
+ $Y2=0
cc_144 A2 N_A_280_107#_c_418_n 0.0521676f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_145 N_A2_c_117_n N_A_280_107#_c_418_n 0.00273128f $X=2.415 $Y=1.557 $X2=0
+ $Y2=0
cc_146 N_A2_M1004_g N_A_280_107#_c_412_n 0.00361295f $X=2.45 $Y=0.74 $X2=0 $Y2=0
cc_147 N_A1_c_174_n N_A_131_368#_c_236_n 0.011796f $X=2.865 $Y=1.765 $X2=0 $Y2=0
cc_148 N_A1_c_175_n N_A_131_368#_c_236_n 0.011796f $X=3.315 $Y=1.765 $X2=0 $Y2=0
cc_149 N_A1_c_174_n N_A_131_368#_c_223_n 0.00729973f $X=2.865 $Y=1.765 $X2=0
+ $Y2=0
cc_150 N_A1_c_175_n N_A_131_368#_c_223_n 5.64076e-19 $X=3.315 $Y=1.765 $X2=0
+ $Y2=0
cc_151 N_A1_c_174_n N_A_131_368#_c_224_n 5.64076e-19 $X=2.865 $Y=1.765 $X2=0
+ $Y2=0
cc_152 N_A1_c_175_n N_A_131_368#_c_224_n 0.00745145f $X=3.315 $Y=1.765 $X2=0
+ $Y2=0
cc_153 N_A1_M1000_g N_Y_c_275_n 0.0116659f $X=2.88 $Y=0.74 $X2=0 $Y2=0
cc_154 N_A1_M1000_g N_Y_c_278_n 0.00625373f $X=2.88 $Y=0.74 $X2=0 $Y2=0
cc_155 N_A1_c_172_n N_Y_c_278_n 0.0117303f $X=3.185 $Y=1.515 $X2=0 $Y2=0
cc_156 N_A1_c_173_n N_Y_c_278_n 7.19315e-19 $X=3.31 $Y=1.557 $X2=0 $Y2=0
cc_157 N_A1_c_174_n N_VPWR_c_331_n 0.00379374f $X=2.865 $Y=1.765 $X2=0 $Y2=0
cc_158 N_A1_c_175_n N_VPWR_c_331_n 0.00379374f $X=3.315 $Y=1.765 $X2=0 $Y2=0
cc_159 N_A1_c_174_n N_VPWR_c_332_n 0.00445602f $X=2.865 $Y=1.765 $X2=0 $Y2=0
cc_160 N_A1_c_175_n N_VPWR_c_335_n 0.00445602f $X=3.315 $Y=1.765 $X2=0 $Y2=0
cc_161 N_A1_c_174_n N_VPWR_c_329_n 0.00857673f $X=2.865 $Y=1.765 $X2=0 $Y2=0
cc_162 N_A1_c_175_n N_VPWR_c_329_n 0.00861148f $X=3.315 $Y=1.765 $X2=0 $Y2=0
cc_163 N_A1_M1000_g N_VGND_c_377_n 0.00288916f $X=2.88 $Y=0.74 $X2=0 $Y2=0
cc_164 N_A1_M1006_g N_VGND_c_377_n 0.00288893f $X=3.31 $Y=0.74 $X2=0 $Y2=0
cc_165 N_A1_M1000_g N_VGND_c_378_n 0.00356354f $X=2.88 $Y=0.74 $X2=0 $Y2=0
cc_166 N_A1_M1006_g N_VGND_c_378_n 0.00360947f $X=3.31 $Y=0.74 $X2=0 $Y2=0
cc_167 N_A1_c_174_n N_A_280_107#_c_418_n 0.0152356f $X=2.865 $Y=1.765 $X2=0
+ $Y2=0
cc_168 N_A1_c_175_n N_A_280_107#_c_418_n 0.0132255f $X=3.315 $Y=1.765 $X2=0
+ $Y2=0
cc_169 N_A1_c_172_n N_A_280_107#_c_418_n 0.0246399f $X=3.185 $Y=1.515 $X2=0
+ $Y2=0
cc_170 N_A1_c_173_n N_A_280_107#_c_418_n 0.00235569f $X=3.31 $Y=1.557 $X2=0
+ $Y2=0
cc_171 N_A1_M1000_g N_A_280_107#_c_412_n 0.0102853f $X=2.88 $Y=0.74 $X2=0 $Y2=0
cc_172 N_A1_M1006_g N_A_280_107#_c_412_n 0.0126982f $X=3.31 $Y=0.74 $X2=0 $Y2=0
cc_173 N_A1_M1006_g N_A_280_107#_c_413_n 0.00157834f $X=3.31 $Y=0.74 $X2=0 $Y2=0
cc_174 N_A1_M1000_g N_A_280_107#_c_414_n 9.37628e-19 $X=2.88 $Y=0.74 $X2=0 $Y2=0
cc_175 N_A1_M1006_g N_A_280_107#_c_414_n 0.00650786f $X=3.31 $Y=0.74 $X2=0 $Y2=0
cc_176 N_A1_M1006_g N_A_280_107#_c_415_n 0.00778767f $X=3.31 $Y=0.74 $X2=0 $Y2=0
cc_177 N_A1_c_175_n N_A_280_107#_c_415_n 0.00634278f $X=3.315 $Y=1.765 $X2=0
+ $Y2=0
cc_178 N_A1_c_172_n N_A_280_107#_c_415_n 0.0323874f $X=3.185 $Y=1.515 $X2=0
+ $Y2=0
cc_179 N_A1_c_173_n N_A_280_107#_c_415_n 0.0108185f $X=3.31 $Y=1.557 $X2=0 $Y2=0
cc_180 N_A1_M1006_g N_A_280_107#_c_416_n 0.00333663f $X=3.31 $Y=0.74 $X2=0 $Y2=0
cc_181 N_A1_c_173_n N_A_280_107#_c_416_n 8.76401e-19 $X=3.31 $Y=1.557 $X2=0
+ $Y2=0
cc_182 N_A_131_368#_c_221_n N_Y_M1007_d 0.00197722f $X=1.565 $Y=2.99 $X2=0 $Y2=0
cc_183 N_A_131_368#_c_220_n N_Y_c_276_n 0.0226071f $X=0.78 $Y=2.115 $X2=0 $Y2=0
cc_184 N_A_131_368#_c_221_n N_Y_c_280_n 0.0160777f $X=1.565 $Y=2.99 $X2=0 $Y2=0
cc_185 N_A_131_368#_c_232_n N_VPWR_M1001_s 0.00526572f $X=2.475 $Y=2.375
+ $X2=-0.19 $Y2=1.66
cc_186 N_A_131_368#_c_236_n N_VPWR_M1003_d 0.00428955f $X=3.375 $Y=2.375 $X2=0
+ $Y2=0
cc_187 N_A_131_368#_c_221_n N_VPWR_c_330_n 0.0123076f $X=1.565 $Y=2.99 $X2=0
+ $Y2=0
cc_188 N_A_131_368#_c_230_n N_VPWR_c_330_n 0.0182369f $X=1.705 $Y=2.905 $X2=0
+ $Y2=0
cc_189 N_A_131_368#_c_232_n N_VPWR_c_330_n 0.019282f $X=2.475 $Y=2.375 $X2=0
+ $Y2=0
cc_190 N_A_131_368#_c_223_n N_VPWR_c_330_n 0.0138953f $X=2.64 $Y=2.455 $X2=0
+ $Y2=0
cc_191 N_A_131_368#_c_236_n N_VPWR_c_331_n 0.0136682f $X=3.375 $Y=2.375 $X2=0
+ $Y2=0
cc_192 N_A_131_368#_c_223_n N_VPWR_c_331_n 0.0228252f $X=2.64 $Y=2.455 $X2=0
+ $Y2=0
cc_193 N_A_131_368#_c_224_n N_VPWR_c_331_n 0.0228252f $X=3.54 $Y=2.455 $X2=0
+ $Y2=0
cc_194 N_A_131_368#_c_223_n N_VPWR_c_332_n 0.0145674f $X=2.64 $Y=2.455 $X2=0
+ $Y2=0
cc_195 N_A_131_368#_c_221_n N_VPWR_c_334_n 0.062212f $X=1.565 $Y=2.99 $X2=0
+ $Y2=0
cc_196 N_A_131_368#_c_222_n N_VPWR_c_334_n 0.0200723f $X=0.895 $Y=2.99 $X2=0
+ $Y2=0
cc_197 N_A_131_368#_c_224_n N_VPWR_c_335_n 0.0146094f $X=3.54 $Y=2.455 $X2=0
+ $Y2=0
cc_198 N_A_131_368#_c_221_n N_VPWR_c_329_n 0.0346291f $X=1.565 $Y=2.99 $X2=0
+ $Y2=0
cc_199 N_A_131_368#_c_222_n N_VPWR_c_329_n 0.0108858f $X=0.895 $Y=2.99 $X2=0
+ $Y2=0
cc_200 N_A_131_368#_c_223_n N_VPWR_c_329_n 0.0119851f $X=2.64 $Y=2.455 $X2=0
+ $Y2=0
cc_201 N_A_131_368#_c_224_n N_VPWR_c_329_n 0.0120527f $X=3.54 $Y=2.455 $X2=0
+ $Y2=0
cc_202 N_A_131_368#_M1008_s N_A_280_107#_c_411_n 3.8009e-19 $X=1.53 $Y=1.84
+ $X2=0 $Y2=0
cc_203 N_A_131_368#_M1009_d N_A_280_107#_c_418_n 0.00392387f $X=2.49 $Y=1.84
+ $X2=0 $Y2=0
cc_204 N_A_131_368#_M1005_s N_A_280_107#_c_418_n 0.00600002f $X=3.39 $Y=1.84
+ $X2=0 $Y2=0
cc_205 N_A_131_368#_c_229_n N_A_280_107#_c_418_n 0.0011005f $X=1.705 $Y=2.46
+ $X2=0 $Y2=0
cc_206 N_A_131_368#_c_232_n N_A_280_107#_c_418_n 0.0361007f $X=2.475 $Y=2.375
+ $X2=0 $Y2=0
cc_207 N_A_131_368#_c_236_n N_A_280_107#_c_418_n 0.0317427f $X=3.375 $Y=2.375
+ $X2=0 $Y2=0
cc_208 N_A_131_368#_c_223_n N_A_280_107#_c_418_n 0.0173542f $X=2.64 $Y=2.455
+ $X2=0 $Y2=0
cc_209 N_A_131_368#_c_224_n N_A_280_107#_c_418_n 0.0223522f $X=3.54 $Y=2.455
+ $X2=0 $Y2=0
cc_210 N_A_131_368#_M1008_s N_A_280_107#_c_458_n 0.00265112f $X=1.53 $Y=1.84
+ $X2=0 $Y2=0
cc_211 N_A_131_368#_c_229_n N_A_280_107#_c_458_n 0.0167701f $X=1.705 $Y=2.46
+ $X2=0 $Y2=0
cc_212 N_A_131_368#_M1005_s N_A_280_107#_c_415_n 0.00180719f $X=3.39 $Y=1.84
+ $X2=0 $Y2=0
cc_213 N_Y_c_275_n N_VGND_M1002_s 0.0114207f $X=2.93 $Y=0.835 $X2=0 $Y2=0
cc_214 N_Y_c_273_n N_VGND_c_374_n 0.0154087f $X=0.695 $Y=0.515 $X2=0 $Y2=0
cc_215 N_Y_c_274_n N_VGND_c_374_n 0.00844336f $X=0.732 $Y=1.55 $X2=0 $Y2=0
cc_216 N_Y_c_275_n N_VGND_c_375_n 0.0249524f $X=2.93 $Y=0.835 $X2=0 $Y2=0
cc_217 N_Y_c_273_n N_VGND_c_376_n 0.0112891f $X=0.695 $Y=0.515 $X2=0 $Y2=0
cc_218 N_Y_c_275_n N_VGND_c_376_n 0.0151647f $X=2.93 $Y=0.835 $X2=0 $Y2=0
cc_219 N_Y_c_275_n N_VGND_c_377_n 0.00190416f $X=2.93 $Y=0.835 $X2=0 $Y2=0
cc_220 N_Y_c_273_n N_VGND_c_378_n 0.00934413f $X=0.695 $Y=0.515 $X2=0 $Y2=0
cc_221 N_Y_c_275_n N_VGND_c_378_n 0.0353693f $X=2.93 $Y=0.835 $X2=0 $Y2=0
cc_222 N_Y_c_275_n N_A_280_107#_M1002_d 0.00936585f $X=2.93 $Y=0.835 $X2=-0.19
+ $Y2=-0.245
cc_223 N_Y_c_275_n N_A_280_107#_M1004_d 0.00387088f $X=2.93 $Y=0.835 $X2=0 $Y2=0
cc_224 N_Y_c_274_n N_A_280_107#_c_410_n 0.00663393f $X=0.732 $Y=1.55 $X2=0 $Y2=0
cc_225 N_Y_c_275_n N_A_280_107#_c_410_n 0.0258668f $X=2.93 $Y=0.835 $X2=0 $Y2=0
cc_226 N_Y_c_276_n N_A_280_107#_c_410_n 0.00186174f $X=1.23 $Y=1.78 $X2=0 $Y2=0
cc_227 N_Y_c_276_n N_A_280_107#_c_411_n 0.0187487f $X=1.23 $Y=1.78 $X2=0 $Y2=0
cc_228 N_Y_c_280_n N_A_280_107#_c_411_n 0.00867101f $X=1.23 $Y=1.97 $X2=0 $Y2=0
cc_229 N_Y_M1000_s N_A_280_107#_c_412_n 0.00178571f $X=2.955 $Y=0.37 $X2=0 $Y2=0
cc_230 N_Y_c_275_n N_A_280_107#_c_412_n 0.0220487f $X=2.93 $Y=0.835 $X2=0 $Y2=0
cc_231 N_Y_c_278_n N_A_280_107#_c_412_n 0.0144731f $X=3.055 $Y=0.835 $X2=0 $Y2=0
cc_232 N_Y_c_278_n N_A_280_107#_c_414_n 0.0143118f $X=3.055 $Y=0.835 $X2=0 $Y2=0
cc_233 N_VPWR_M1001_s N_A_280_107#_c_418_n 0.00478997f $X=1.98 $Y=1.84 $X2=0
+ $Y2=0
cc_234 N_VPWR_M1003_d N_A_280_107#_c_418_n 0.0036296f $X=2.94 $Y=1.84 $X2=0
+ $Y2=0
cc_235 N_VGND_c_375_n N_A_280_107#_c_412_n 0.0120344f $X=2.165 $Y=0.495 $X2=0
+ $Y2=0
cc_236 N_VGND_c_377_n N_A_280_107#_c_412_n 0.0378512f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_237 N_VGND_c_378_n N_A_280_107#_c_412_n 0.0297248f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_238 N_VGND_c_377_n N_A_280_107#_c_413_n 0.0159296f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_239 N_VGND_c_378_n N_A_280_107#_c_413_n 0.0122131f $X=3.6 $Y=0 $X2=0 $Y2=0
