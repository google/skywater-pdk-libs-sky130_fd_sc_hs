* File: sky130_fd_sc_hs__o21ai_4.pxi.spice
* Created: Thu Aug 27 20:58:12 2020
* 
x_PM_SKY130_FD_SC_HS__O21AI_4%A1 N_A1_M1006_g N_A1_c_98_n N_A1_M1008_g
+ N_A1_M1018_g N_A1_c_99_n N_A1_M1009_g N_A1_M1019_g N_A1_c_100_n N_A1_M1010_g
+ N_A1_M1021_g N_A1_c_101_n N_A1_M1012_g A1 A1 N_A1_c_97_n N_A1_c_127_p
+ PM_SKY130_FD_SC_HS__O21AI_4%A1
x_PM_SKY130_FD_SC_HS__O21AI_4%B1 N_B1_c_178_n N_B1_M1003_g N_B1_c_185_n
+ N_B1_M1013_g N_B1_c_179_n N_B1_M1004_g N_B1_c_186_n N_B1_M1014_g N_B1_c_180_n
+ N_B1_M1007_g N_B1_c_181_n N_B1_c_182_n N_B1_c_183_n N_B1_M1016_g B1 B1
+ N_B1_c_184_n PM_SKY130_FD_SC_HS__O21AI_4%B1
x_PM_SKY130_FD_SC_HS__O21AI_4%A2 N_A2_c_256_n N_A2_M1002_g N_A2_M1000_g
+ N_A2_c_257_n N_A2_M1015_g N_A2_M1001_g N_A2_c_258_n N_A2_M1017_g N_A2_M1005_g
+ N_A2_c_259_n N_A2_M1020_g N_A2_M1011_g A2 A2 A2 A2 N_A2_c_255_n
+ PM_SKY130_FD_SC_HS__O21AI_4%A2
x_PM_SKY130_FD_SC_HS__O21AI_4%VPWR N_VPWR_M1008_d N_VPWR_M1009_d N_VPWR_M1012_d
+ N_VPWR_M1014_s N_VPWR_c_330_n N_VPWR_c_331_n N_VPWR_c_332_n N_VPWR_c_333_n
+ N_VPWR_c_334_n N_VPWR_c_335_n N_VPWR_c_336_n VPWR N_VPWR_c_337_n
+ N_VPWR_c_338_n N_VPWR_c_339_n N_VPWR_c_329_n N_VPWR_c_341_n N_VPWR_c_342_n
+ PM_SKY130_FD_SC_HS__O21AI_4%VPWR
x_PM_SKY130_FD_SC_HS__O21AI_4%A_116_368# N_A_116_368#_M1008_s
+ N_A_116_368#_M1010_s N_A_116_368#_M1002_d N_A_116_368#_M1015_d
+ N_A_116_368#_M1020_d N_A_116_368#_c_399_n N_A_116_368#_c_400_n
+ N_A_116_368#_c_418_n N_A_116_368#_c_423_n N_A_116_368#_c_427_n
+ N_A_116_368#_c_401_n N_A_116_368#_c_402_n N_A_116_368#_c_403_n
+ N_A_116_368#_c_404_n N_A_116_368#_c_405_n N_A_116_368#_c_406_n
+ N_A_116_368#_c_484_p N_A_116_368#_c_407_n N_A_116_368#_c_408_n
+ N_A_116_368#_c_433_n N_A_116_368#_c_409_n
+ PM_SKY130_FD_SC_HS__O21AI_4%A_116_368#
x_PM_SKY130_FD_SC_HS__O21AI_4%Y N_Y_M1003_d N_Y_M1007_d N_Y_M1013_d N_Y_M1002_s
+ N_Y_M1017_s N_Y_c_495_n N_Y_c_503_n N_Y_c_520_n N_Y_c_521_n N_Y_c_507_n
+ N_Y_c_510_n N_Y_c_525_n N_Y_c_529_n Y N_Y_c_494_n
+ PM_SKY130_FD_SC_HS__O21AI_4%Y
x_PM_SKY130_FD_SC_HS__O21AI_4%A_27_74# N_A_27_74#_M1006_s N_A_27_74#_M1018_s
+ N_A_27_74#_M1021_s N_A_27_74#_M1004_s N_A_27_74#_M1016_s N_A_27_74#_M1001_s
+ N_A_27_74#_M1011_s N_A_27_74#_c_569_n N_A_27_74#_c_570_n N_A_27_74#_c_571_n
+ N_A_27_74#_c_572_n N_A_27_74#_c_591_n N_A_27_74#_c_573_n N_A_27_74#_c_574_n
+ N_A_27_74#_c_575_n N_A_27_74#_c_604_n N_A_27_74#_c_576_n N_A_27_74#_c_577_n
+ N_A_27_74#_c_578_n N_A_27_74#_c_579_n N_A_27_74#_c_580_n N_A_27_74#_c_581_n
+ N_A_27_74#_c_582_n N_A_27_74#_c_583_n PM_SKY130_FD_SC_HS__O21AI_4%A_27_74#
x_PM_SKY130_FD_SC_HS__O21AI_4%VGND N_VGND_M1006_d N_VGND_M1019_d N_VGND_M1000_d
+ N_VGND_M1005_d N_VGND_c_670_n N_VGND_c_671_n N_VGND_c_672_n N_VGND_c_673_n
+ N_VGND_c_674_n VGND N_VGND_c_675_n N_VGND_c_676_n N_VGND_c_677_n
+ N_VGND_c_678_n N_VGND_c_679_n N_VGND_c_680_n N_VGND_c_681_n N_VGND_c_682_n
+ N_VGND_c_683_n PM_SKY130_FD_SC_HS__O21AI_4%VGND
cc_1 VNB N_A1_M1006_g 0.0301354f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_2 VNB N_A1_M1018_g 0.0212151f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=0.74
cc_3 VNB N_A1_M1019_g 0.0217592f $X=-0.19 $Y=-0.245 $X2=1.355 $Y2=0.74
cc_4 VNB N_A1_M1021_g 0.0222874f $X=-0.19 $Y=-0.245 $X2=1.8 $Y2=0.74
cc_5 VNB N_A1_c_97_n 0.11228f $X=-0.19 $Y=-0.245 $X2=1.8 $Y2=1.542
cc_6 VNB N_B1_c_178_n 0.0144853f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.32
cc_7 VNB N_B1_c_179_n 0.0143176f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_8 VNB N_B1_c_180_n 0.0142846f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=2.4
cc_9 VNB N_B1_c_181_n 0.0246434f $X=-0.19 $Y=-0.245 $X2=1.355 $Y2=0.74
cc_10 VNB N_B1_c_182_n 0.0828277f $X=-0.19 $Y=-0.245 $X2=1.355 $Y2=0.74
cc_11 VNB N_B1_c_183_n 0.0143551f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_B1_c_184_n 0.0170818f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.58
cc_13 VNB N_A2_M1000_g 0.0233837f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_14 VNB N_A2_M1001_g 0.0224899f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=2.4
cc_15 VNB N_A2_M1005_g 0.0224899f $X=-0.19 $Y=-0.245 $X2=1.405 $Y2=2.4
cc_16 VNB N_A2_M1011_g 0.0318708f $X=-0.19 $Y=-0.245 $X2=1.855 $Y2=2.4
cc_17 VNB A2 0.0166485f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.485
cc_18 VNB N_A2_c_255_n 0.0779558f $X=-0.19 $Y=-0.245 $X2=1.63 $Y2=1.485
cc_19 VNB N_VPWR_c_329_n 0.243291f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB Y 0.00850576f $X=-0.19 $Y=-0.245 $X2=1.355 $Y2=1.542
cc_21 VNB N_Y_c_494_n 0.00427957f $X=-0.19 $Y=-0.245 $X2=1.63 $Y2=1.485
cc_22 VNB N_A_27_74#_c_569_n 0.0255089f $X=-0.19 $Y=-0.245 $X2=1.8 $Y2=0.74
cc_23 VNB N_A_27_74#_c_570_n 0.00456647f $X=-0.19 $Y=-0.245 $X2=1.855 $Y2=1.765
cc_24 VNB N_A_27_74#_c_571_n 0.0115038f $X=-0.19 $Y=-0.245 $X2=1.855 $Y2=2.4
cc_25 VNB N_A_27_74#_c_572_n 0.00178908f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.485
cc_26 VNB N_A_27_74#_c_573_n 0.00237811f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.542
cc_27 VNB N_A_27_74#_c_574_n 0.00213254f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.542
cc_28 VNB N_A_27_74#_c_575_n 0.00477762f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.542
cc_29 VNB N_A_27_74#_c_576_n 0.00337922f $X=-0.19 $Y=-0.245 $X2=1.355 $Y2=1.542
cc_30 VNB N_A_27_74#_c_577_n 0.00405692f $X=-0.19 $Y=-0.245 $X2=1.405 $Y2=1.542
cc_31 VNB N_A_27_74#_c_578_n 0.00178908f $X=-0.19 $Y=-0.245 $X2=1.63 $Y2=1.485
cc_32 VNB N_A_27_74#_c_579_n 0.0132288f $X=-0.19 $Y=-0.245 $X2=1.855 $Y2=1.542
cc_33 VNB N_A_27_74#_c_580_n 0.0266107f $X=-0.19 $Y=-0.245 $X2=1.29 $Y2=1.55
cc_34 VNB N_A_27_74#_c_581_n 0.00167779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_27_74#_c_582_n 0.00202117f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_27_74#_c_583_n 0.00127131f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_670_n 0.00323505f $X=-0.19 $Y=-0.245 $X2=1.355 $Y2=1.32
cc_38 VNB N_VGND_c_671_n 0.00323505f $X=-0.19 $Y=-0.245 $X2=1.405 $Y2=1.765
cc_39 VNB N_VGND_c_672_n 0.0539351f $X=-0.19 $Y=-0.245 $X2=1.405 $Y2=2.4
cc_40 VNB N_VGND_c_673_n 0.00323505f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_674_n 0.00323505f $X=-0.19 $Y=-0.245 $X2=1.085 $Y2=1.485
cc_42 VNB N_VGND_c_675_n 0.0173909f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_676_n 0.0151736f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.542
cc_44 VNB N_VGND_c_677_n 0.0151736f $X=-0.19 $Y=-0.245 $X2=1.29 $Y2=1.542
cc_45 VNB N_VGND_c_678_n 0.0173909f $X=-0.19 $Y=-0.245 $X2=1.63 $Y2=1.485
cc_46 VNB N_VGND_c_679_n 0.31955f $X=-0.19 $Y=-0.245 $X2=1.8 $Y2=1.542
cc_47 VNB N_VGND_c_680_n 0.00604233f $X=-0.19 $Y=-0.245 $X2=1.085 $Y2=1.55
cc_48 VNB N_VGND_c_681_n 0.00604233f $X=-0.19 $Y=-0.245 $X2=1.63 $Y2=1.55
cc_49 VNB N_VGND_c_682_n 0.00604233f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_VGND_c_683_n 0.00604233f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VPB N_A1_c_98_n 0.01766f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.765
cc_52 VPB N_A1_c_99_n 0.0155173f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=1.765
cc_53 VPB N_A1_c_100_n 0.0155113f $X=-0.19 $Y=1.66 $X2=1.405 $Y2=1.765
cc_54 VPB N_A1_c_101_n 0.0158896f $X=-0.19 $Y=1.66 $X2=1.855 $Y2=1.765
cc_55 VPB A1 0.00637183f $X=-0.19 $Y=1.66 $X2=1.595 $Y2=1.58
cc_56 VPB N_A1_c_97_n 0.0281574f $X=-0.19 $Y=1.66 $X2=1.8 $Y2=1.542
cc_57 VPB N_B1_c_185_n 0.0151476f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_58 VPB N_B1_c_186_n 0.0168537f $X=-0.19 $Y=1.66 $X2=0.925 $Y2=0.74
cc_59 VPB N_B1_c_182_n 0.0141887f $X=-0.19 $Y=1.66 $X2=1.355 $Y2=0.74
cc_60 VPB N_A2_c_256_n 0.0172331f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.32
cc_61 VPB N_A2_c_257_n 0.0150448f $X=-0.19 $Y=1.66 $X2=0.925 $Y2=1.32
cc_62 VPB N_A2_c_258_n 0.014664f $X=-0.19 $Y=1.66 $X2=1.355 $Y2=1.32
cc_63 VPB N_A2_c_259_n 0.0186669f $X=-0.19 $Y=1.66 $X2=1.8 $Y2=1.32
cc_64 VPB A2 0.0190111f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=1.485
cc_65 VPB N_A2_c_255_n 0.0506704f $X=-0.19 $Y=1.66 $X2=1.63 $Y2=1.485
cc_66 VPB N_VPWR_c_330_n 0.0106521f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=2.4
cc_67 VPB N_VPWR_c_331_n 0.0587411f $X=-0.19 $Y=1.66 $X2=1.355 $Y2=1.32
cc_68 VPB N_VPWR_c_332_n 0.00799266f $X=-0.19 $Y=1.66 $X2=1.405 $Y2=2.4
cc_69 VPB N_VPWR_c_333_n 0.00514935f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_70 VPB N_VPWR_c_334_n 0.0122137f $X=-0.19 $Y=1.66 $X2=1.085 $Y2=1.485
cc_71 VPB N_VPWR_c_335_n 0.0206041f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=1.485
cc_72 VPB N_VPWR_c_336_n 0.00324402f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_73 VPB N_VPWR_c_337_n 0.0206041f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=1.542
cc_74 VPB N_VPWR_c_338_n 0.0206218f $X=-0.19 $Y=1.66 $X2=1.29 $Y2=1.485
cc_75 VPB N_VPWR_c_339_n 0.0615915f $X=-0.19 $Y=1.66 $X2=1.085 $Y2=1.55
cc_76 VPB N_VPWR_c_329_n 0.0965427f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_77 VPB N_VPWR_c_341_n 0.00460249f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_78 VPB N_VPWR_c_342_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_79 VPB N_A_116_368#_c_399_n 0.00183525f $X=-0.19 $Y=1.66 $X2=1.355 $Y2=0.74
cc_80 VPB N_A_116_368#_c_400_n 0.00257348f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_81 VPB N_A_116_368#_c_401_n 0.00257348f $X=-0.19 $Y=1.66 $X2=1.855 $Y2=1.765
cc_82 VPB N_A_116_368#_c_402_n 0.0118988f $X=-0.19 $Y=1.66 $X2=1.855 $Y2=2.4
cc_83 VPB N_A_116_368#_c_403_n 3.13193e-19 $X=-0.19 $Y=1.66 $X2=0.61 $Y2=1.485
cc_84 VPB N_A_116_368#_c_404_n 0.00526935f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=1.485
cc_85 VPB N_A_116_368#_c_405_n 0.00294772f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=1.485
cc_86 VPB N_A_116_368#_c_406_n 0.0043681f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_87 VPB N_A_116_368#_c_407_n 0.0124059f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.542
cc_88 VPB N_A_116_368#_c_408_n 0.0351758f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=1.542
cc_89 VPB N_A_116_368#_c_409_n 0.00123754f $X=-0.19 $Y=1.66 $X2=1.2 $Y2=1.55
cc_90 VPB N_Y_c_495_n 0.0109935f $X=-0.19 $Y=1.66 $X2=1.355 $Y2=0.74
cc_91 VPB Y 0.00938845f $X=-0.19 $Y=1.66 $X2=1.355 $Y2=1.542
cc_92 N_A1_M1021_g N_B1_c_178_n 0.0181168f $X=1.8 $Y=0.74 $X2=-0.19 $Y2=-0.245
cc_93 N_A1_c_101_n N_B1_c_185_n 0.0398459f $X=1.855 $Y=1.765 $X2=0 $Y2=0
cc_94 A1 N_B1_c_182_n 0.00120289f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_95 N_A1_c_97_n N_B1_c_182_n 0.0263219f $X=1.8 $Y=1.542 $X2=0 $Y2=0
cc_96 N_A1_M1021_g N_B1_c_184_n 0.00382458f $X=1.8 $Y=0.74 $X2=0 $Y2=0
cc_97 A1 N_B1_c_184_n 0.0151989f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_98 N_A1_c_97_n N_B1_c_184_n 0.00213182f $X=1.8 $Y=1.542 $X2=0 $Y2=0
cc_99 N_A1_c_98_n N_VPWR_c_331_n 0.0100869f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_100 N_A1_c_99_n N_VPWR_c_332_n 0.00486623f $X=0.955 $Y=1.765 $X2=0 $Y2=0
cc_101 N_A1_c_100_n N_VPWR_c_332_n 0.00486381f $X=1.405 $Y=1.765 $X2=0 $Y2=0
cc_102 N_A1_c_101_n N_VPWR_c_333_n 0.00409001f $X=1.855 $Y=1.765 $X2=0 $Y2=0
cc_103 N_A1_c_98_n N_VPWR_c_335_n 0.00445602f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_104 N_A1_c_99_n N_VPWR_c_335_n 0.00445602f $X=0.955 $Y=1.765 $X2=0 $Y2=0
cc_105 N_A1_c_100_n N_VPWR_c_337_n 0.00445602f $X=1.405 $Y=1.765 $X2=0 $Y2=0
cc_106 N_A1_c_101_n N_VPWR_c_337_n 0.00445602f $X=1.855 $Y=1.765 $X2=0 $Y2=0
cc_107 N_A1_c_98_n N_VPWR_c_329_n 0.00861084f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_108 N_A1_c_99_n N_VPWR_c_329_n 0.00857589f $X=0.955 $Y=1.765 $X2=0 $Y2=0
cc_109 N_A1_c_100_n N_VPWR_c_329_n 0.00857589f $X=1.405 $Y=1.765 $X2=0 $Y2=0
cc_110 N_A1_c_101_n N_VPWR_c_329_n 0.00857673f $X=1.855 $Y=1.765 $X2=0 $Y2=0
cc_111 N_A1_c_98_n N_A_116_368#_c_399_n 0.00369554f $X=0.505 $Y=1.765 $X2=0
+ $Y2=0
cc_112 N_A1_c_99_n N_A_116_368#_c_399_n 0.00301134f $X=0.955 $Y=1.765 $X2=0
+ $Y2=0
cc_113 N_A1_c_100_n N_A_116_368#_c_399_n 6.18219e-19 $X=1.405 $Y=1.765 $X2=0
+ $Y2=0
cc_114 N_A1_c_97_n N_A_116_368#_c_399_n 0.00789892f $X=1.8 $Y=1.542 $X2=0 $Y2=0
cc_115 N_A1_c_127_p N_A_116_368#_c_399_n 0.0276944f $X=1.085 $Y=1.55 $X2=0 $Y2=0
cc_116 N_A1_c_98_n N_A_116_368#_c_400_n 0.0102459f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_117 N_A1_c_99_n N_A_116_368#_c_400_n 0.0109808f $X=0.955 $Y=1.765 $X2=0 $Y2=0
cc_118 N_A1_c_100_n N_A_116_368#_c_400_n 6.45594e-19 $X=1.405 $Y=1.765 $X2=0
+ $Y2=0
cc_119 N_A1_c_99_n N_A_116_368#_c_418_n 0.0126678f $X=0.955 $Y=1.765 $X2=0 $Y2=0
cc_120 N_A1_c_100_n N_A_116_368#_c_418_n 0.0120074f $X=1.405 $Y=1.765 $X2=0
+ $Y2=0
cc_121 A1 N_A_116_368#_c_418_n 0.0273513f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_122 N_A1_c_97_n N_A_116_368#_c_418_n 0.00108932f $X=1.8 $Y=1.542 $X2=0 $Y2=0
cc_123 N_A1_c_127_p N_A_116_368#_c_418_n 0.00738639f $X=1.085 $Y=1.55 $X2=0
+ $Y2=0
cc_124 N_A1_c_100_n N_A_116_368#_c_423_n 4.27055e-19 $X=1.405 $Y=1.765 $X2=0
+ $Y2=0
cc_125 N_A1_c_101_n N_A_116_368#_c_423_n 0.00317113f $X=1.855 $Y=1.765 $X2=0
+ $Y2=0
cc_126 A1 N_A_116_368#_c_423_n 0.0239057f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_127 N_A1_c_97_n N_A_116_368#_c_423_n 0.0013489f $X=1.8 $Y=1.542 $X2=0 $Y2=0
cc_128 N_A1_c_99_n N_A_116_368#_c_427_n 4.35082e-19 $X=0.955 $Y=1.765 $X2=0
+ $Y2=0
cc_129 N_A1_c_100_n N_A_116_368#_c_427_n 0.00294319f $X=1.405 $Y=1.765 $X2=0
+ $Y2=0
cc_130 N_A1_c_101_n N_A_116_368#_c_427_n 0.00299327f $X=1.855 $Y=1.765 $X2=0
+ $Y2=0
cc_131 N_A1_c_100_n N_A_116_368#_c_401_n 0.00564712f $X=1.405 $Y=1.765 $X2=0
+ $Y2=0
cc_132 N_A1_c_101_n N_A_116_368#_c_401_n 0.00694321f $X=1.855 $Y=1.765 $X2=0
+ $Y2=0
cc_133 N_A1_c_101_n N_A_116_368#_c_402_n 0.0158375f $X=1.855 $Y=1.765 $X2=0
+ $Y2=0
cc_134 N_A1_c_100_n N_A_116_368#_c_433_n 0.0017329f $X=1.405 $Y=1.765 $X2=0
+ $Y2=0
cc_135 N_A1_c_101_n N_A_116_368#_c_433_n 2.24111e-19 $X=1.855 $Y=1.765 $X2=0
+ $Y2=0
cc_136 N_A1_c_101_n N_Y_c_495_n 0.00110428f $X=1.855 $Y=1.765 $X2=0 $Y2=0
cc_137 N_A1_M1006_g N_A_27_74#_c_569_n 0.00159319f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_138 N_A1_M1006_g N_A_27_74#_c_570_n 0.0137448f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_139 N_A1_M1018_g N_A_27_74#_c_570_n 0.0124568f $X=0.925 $Y=0.74 $X2=0 $Y2=0
cc_140 N_A1_c_97_n N_A_27_74#_c_570_n 0.00243702f $X=1.8 $Y=1.542 $X2=0 $Y2=0
cc_141 N_A1_c_127_p N_A_27_74#_c_570_n 0.0448197f $X=1.085 $Y=1.55 $X2=0 $Y2=0
cc_142 N_A1_M1018_g N_A_27_74#_c_572_n 3.92313e-19 $X=0.925 $Y=0.74 $X2=0 $Y2=0
cc_143 N_A1_M1019_g N_A_27_74#_c_572_n 3.92313e-19 $X=1.355 $Y=0.74 $X2=0 $Y2=0
cc_144 N_A1_M1019_g N_A_27_74#_c_591_n 0.0104439f $X=1.355 $Y=0.74 $X2=0 $Y2=0
cc_145 N_A1_M1021_g N_A_27_74#_c_591_n 0.0125823f $X=1.8 $Y=0.74 $X2=0 $Y2=0
cc_146 A1 N_A_27_74#_c_591_n 0.0227309f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_147 N_A1_c_97_n N_A_27_74#_c_591_n 0.00288743f $X=1.8 $Y=1.542 $X2=0 $Y2=0
cc_148 N_A1_M1021_g N_A_27_74#_c_574_n 9.83948e-19 $X=1.8 $Y=0.74 $X2=0 $Y2=0
cc_149 N_A1_M1019_g N_A_27_74#_c_581_n 9.34957e-19 $X=1.355 $Y=0.74 $X2=0 $Y2=0
cc_150 N_A1_c_97_n N_A_27_74#_c_581_n 0.00232957f $X=1.8 $Y=1.542 $X2=0 $Y2=0
cc_151 N_A1_c_127_p N_A_27_74#_c_581_n 0.0144048f $X=1.085 $Y=1.55 $X2=0 $Y2=0
cc_152 N_A1_M1006_g N_VGND_c_670_n 0.0127296f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_153 N_A1_M1018_g N_VGND_c_670_n 0.00970341f $X=0.925 $Y=0.74 $X2=0 $Y2=0
cc_154 N_A1_M1019_g N_VGND_c_670_n 4.62684e-19 $X=1.355 $Y=0.74 $X2=0 $Y2=0
cc_155 N_A1_M1018_g N_VGND_c_671_n 4.20905e-19 $X=0.925 $Y=0.74 $X2=0 $Y2=0
cc_156 N_A1_M1019_g N_VGND_c_671_n 0.00765209f $X=1.355 $Y=0.74 $X2=0 $Y2=0
cc_157 N_A1_M1021_g N_VGND_c_671_n 0.00617842f $X=1.8 $Y=0.74 $X2=0 $Y2=0
cc_158 N_A1_M1021_g N_VGND_c_672_n 0.00429299f $X=1.8 $Y=0.74 $X2=0 $Y2=0
cc_159 N_A1_M1006_g N_VGND_c_675_n 0.00383152f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_160 N_A1_M1018_g N_VGND_c_676_n 0.00383152f $X=0.925 $Y=0.74 $X2=0 $Y2=0
cc_161 N_A1_M1019_g N_VGND_c_676_n 0.00383152f $X=1.355 $Y=0.74 $X2=0 $Y2=0
cc_162 N_A1_M1006_g N_VGND_c_679_n 0.00761198f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_163 N_A1_M1018_g N_VGND_c_679_n 0.0075754f $X=0.925 $Y=0.74 $X2=0 $Y2=0
cc_164 N_A1_M1019_g N_VGND_c_679_n 0.00383967f $X=1.355 $Y=0.74 $X2=0 $Y2=0
cc_165 N_A1_M1021_g N_VGND_c_679_n 0.00429576f $X=1.8 $Y=0.74 $X2=0 $Y2=0
cc_166 N_B1_c_183_n N_A2_M1000_g 0.0164408f $X=3.52 $Y=1.185 $X2=0 $Y2=0
cc_167 N_B1_c_185_n N_VPWR_c_333_n 0.0103579f $X=2.305 $Y=1.765 $X2=0 $Y2=0
cc_168 N_B1_c_186_n N_VPWR_c_333_n 0.00140581f $X=2.755 $Y=1.765 $X2=0 $Y2=0
cc_169 N_B1_c_186_n N_VPWR_c_334_n 0.0131598f $X=2.755 $Y=1.765 $X2=0 $Y2=0
cc_170 N_B1_c_185_n N_VPWR_c_338_n 0.00413917f $X=2.305 $Y=1.765 $X2=0 $Y2=0
cc_171 N_B1_c_186_n N_VPWR_c_338_n 0.00461464f $X=2.755 $Y=1.765 $X2=0 $Y2=0
cc_172 N_B1_c_185_n N_VPWR_c_329_n 0.00817726f $X=2.305 $Y=1.765 $X2=0 $Y2=0
cc_173 N_B1_c_186_n N_VPWR_c_329_n 0.00913865f $X=2.755 $Y=1.765 $X2=0 $Y2=0
cc_174 N_B1_c_185_n N_A_116_368#_c_423_n 5.01926e-19 $X=2.305 $Y=1.765 $X2=0
+ $Y2=0
cc_175 N_B1_c_185_n N_A_116_368#_c_427_n 8.01914e-19 $X=2.305 $Y=1.765 $X2=0
+ $Y2=0
cc_176 N_B1_c_185_n N_A_116_368#_c_401_n 8.76141e-19 $X=2.305 $Y=1.765 $X2=0
+ $Y2=0
cc_177 N_B1_c_185_n N_A_116_368#_c_402_n 0.0187431f $X=2.305 $Y=1.765 $X2=0
+ $Y2=0
cc_178 N_B1_c_186_n N_A_116_368#_c_402_n 0.0169977f $X=2.755 $Y=1.765 $X2=0
+ $Y2=0
cc_179 N_B1_c_186_n N_A_116_368#_c_404_n 0.00431194f $X=2.755 $Y=1.765 $X2=0
+ $Y2=0
cc_180 N_B1_c_185_n N_Y_c_495_n 0.00616046f $X=2.305 $Y=1.765 $X2=0 $Y2=0
cc_181 N_B1_c_186_n N_Y_c_495_n 0.0159253f $X=2.755 $Y=1.765 $X2=0 $Y2=0
cc_182 N_B1_c_181_n N_Y_c_495_n 0.00492945f $X=3.445 $Y=1.26 $X2=0 $Y2=0
cc_183 N_B1_c_182_n N_Y_c_495_n 0.011339f $X=3.165 $Y=1.26 $X2=0 $Y2=0
cc_184 N_B1_c_184_n N_Y_c_495_n 0.0442063f $X=3 $Y=1.385 $X2=0 $Y2=0
cc_185 N_B1_c_179_n N_Y_c_503_n 0.00950771f $X=2.66 $Y=1.185 $X2=0 $Y2=0
cc_186 N_B1_c_180_n N_Y_c_503_n 0.00950771f $X=3.09 $Y=1.185 $X2=0 $Y2=0
cc_187 N_B1_c_182_n N_Y_c_503_n 6.93344e-19 $X=3.165 $Y=1.26 $X2=0 $Y2=0
cc_188 N_B1_c_184_n N_Y_c_503_n 0.0418422f $X=3 $Y=1.385 $X2=0 $Y2=0
cc_189 N_B1_c_178_n N_Y_c_507_n 0.00516423f $X=2.23 $Y=1.185 $X2=0 $Y2=0
cc_190 N_B1_c_182_n N_Y_c_507_n 7.37755e-19 $X=3.165 $Y=1.26 $X2=0 $Y2=0
cc_191 N_B1_c_184_n N_Y_c_507_n 0.0183113f $X=3 $Y=1.385 $X2=0 $Y2=0
cc_192 N_B1_c_181_n N_Y_c_510_n 0.00304357f $X=3.445 $Y=1.26 $X2=0 $Y2=0
cc_193 N_B1_c_183_n N_Y_c_510_n 0.00625443f $X=3.52 $Y=1.185 $X2=0 $Y2=0
cc_194 N_B1_c_186_n Y 0.00216582f $X=2.755 $Y=1.765 $X2=0 $Y2=0
cc_195 N_B1_c_181_n Y 0.0040411f $X=3.445 $Y=1.26 $X2=0 $Y2=0
cc_196 N_B1_c_182_n Y 0.00591268f $X=3.165 $Y=1.26 $X2=0 $Y2=0
cc_197 N_B1_c_180_n N_Y_c_494_n 0.00351883f $X=3.09 $Y=1.185 $X2=0 $Y2=0
cc_198 N_B1_c_181_n N_Y_c_494_n 0.0112144f $X=3.445 $Y=1.26 $X2=0 $Y2=0
cc_199 N_B1_c_182_n N_Y_c_494_n 0.00148844f $X=3.165 $Y=1.26 $X2=0 $Y2=0
cc_200 N_B1_c_183_n N_Y_c_494_n 0.00324088f $X=3.52 $Y=1.185 $X2=0 $Y2=0
cc_201 N_B1_c_184_n N_Y_c_494_n 0.0288059f $X=3 $Y=1.385 $X2=0 $Y2=0
cc_202 N_B1_c_184_n N_A_27_74#_c_591_n 0.00471836f $X=3 $Y=1.385 $X2=0 $Y2=0
cc_203 N_B1_c_178_n N_A_27_74#_c_573_n 0.0120041f $X=2.23 $Y=1.185 $X2=0 $Y2=0
cc_204 N_B1_c_179_n N_A_27_74#_c_573_n 0.00785166f $X=2.66 $Y=1.185 $X2=0 $Y2=0
cc_205 N_B1_c_180_n N_A_27_74#_c_575_n 0.00785166f $X=3.09 $Y=1.185 $X2=0 $Y2=0
cc_206 N_B1_c_183_n N_A_27_74#_c_575_n 0.0110523f $X=3.52 $Y=1.185 $X2=0 $Y2=0
cc_207 N_B1_c_183_n N_A_27_74#_c_604_n 0.00271595f $X=3.52 $Y=1.185 $X2=0 $Y2=0
cc_208 N_B1_c_183_n N_A_27_74#_c_577_n 9.24829e-19 $X=3.52 $Y=1.185 $X2=0 $Y2=0
cc_209 N_B1_c_178_n N_A_27_74#_c_582_n 6.25215e-19 $X=2.23 $Y=1.185 $X2=0 $Y2=0
cc_210 N_B1_c_179_n N_A_27_74#_c_582_n 0.00663416f $X=2.66 $Y=1.185 $X2=0 $Y2=0
cc_211 N_B1_c_180_n N_A_27_74#_c_582_n 0.00669566f $X=3.09 $Y=1.185 $X2=0 $Y2=0
cc_212 N_B1_c_183_n N_A_27_74#_c_582_n 6.30166e-19 $X=3.52 $Y=1.185 $X2=0 $Y2=0
cc_213 N_B1_c_178_n N_VGND_c_672_n 0.00278271f $X=2.23 $Y=1.185 $X2=0 $Y2=0
cc_214 N_B1_c_179_n N_VGND_c_672_n 0.00279469f $X=2.66 $Y=1.185 $X2=0 $Y2=0
cc_215 N_B1_c_180_n N_VGND_c_672_n 0.00279469f $X=3.09 $Y=1.185 $X2=0 $Y2=0
cc_216 N_B1_c_183_n N_VGND_c_672_n 0.00278271f $X=3.52 $Y=1.185 $X2=0 $Y2=0
cc_217 N_B1_c_178_n N_VGND_c_679_n 0.00353526f $X=2.23 $Y=1.185 $X2=0 $Y2=0
cc_218 N_B1_c_179_n N_VGND_c_679_n 0.00352518f $X=2.66 $Y=1.185 $X2=0 $Y2=0
cc_219 N_B1_c_180_n N_VGND_c_679_n 0.00352518f $X=3.09 $Y=1.185 $X2=0 $Y2=0
cc_220 N_B1_c_183_n N_VGND_c_679_n 0.00353754f $X=3.52 $Y=1.185 $X2=0 $Y2=0
cc_221 N_A2_c_256_n N_VPWR_c_334_n 0.0013297f $X=3.85 $Y=1.765 $X2=0 $Y2=0
cc_222 N_A2_c_256_n N_VPWR_c_339_n 0.00278257f $X=3.85 $Y=1.765 $X2=0 $Y2=0
cc_223 N_A2_c_257_n N_VPWR_c_339_n 0.00278271f $X=4.35 $Y=1.765 $X2=0 $Y2=0
cc_224 N_A2_c_258_n N_VPWR_c_339_n 0.00278271f $X=4.8 $Y=1.765 $X2=0 $Y2=0
cc_225 N_A2_c_259_n N_VPWR_c_339_n 0.00278271f $X=5.25 $Y=1.765 $X2=0 $Y2=0
cc_226 N_A2_c_256_n N_VPWR_c_329_n 0.00359084f $X=3.85 $Y=1.765 $X2=0 $Y2=0
cc_227 N_A2_c_257_n N_VPWR_c_329_n 0.00354284f $X=4.35 $Y=1.765 $X2=0 $Y2=0
cc_228 N_A2_c_258_n N_VPWR_c_329_n 0.00353823f $X=4.8 $Y=1.765 $X2=0 $Y2=0
cc_229 N_A2_c_259_n N_VPWR_c_329_n 0.00357334f $X=5.25 $Y=1.765 $X2=0 $Y2=0
cc_230 N_A2_c_256_n N_A_116_368#_c_403_n 0.00183099f $X=3.85 $Y=1.765 $X2=0
+ $Y2=0
cc_231 N_A2_c_256_n N_A_116_368#_c_404_n 0.00574879f $X=3.85 $Y=1.765 $X2=0
+ $Y2=0
cc_232 N_A2_c_257_n N_A_116_368#_c_404_n 7.18055e-19 $X=4.35 $Y=1.765 $X2=0
+ $Y2=0
cc_233 N_A2_c_256_n N_A_116_368#_c_405_n 0.0111147f $X=3.85 $Y=1.765 $X2=0 $Y2=0
cc_234 N_A2_c_257_n N_A_116_368#_c_405_n 0.0131082f $X=4.35 $Y=1.765 $X2=0 $Y2=0
cc_235 N_A2_c_256_n N_A_116_368#_c_406_n 0.00262934f $X=3.85 $Y=1.765 $X2=0
+ $Y2=0
cc_236 N_A2_c_258_n N_A_116_368#_c_407_n 0.0128349f $X=4.8 $Y=1.765 $X2=0 $Y2=0
cc_237 N_A2_c_259_n N_A_116_368#_c_407_n 0.0137046f $X=5.25 $Y=1.765 $X2=0 $Y2=0
cc_238 A2 N_A_116_368#_c_408_n 0.0215956f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_239 N_A2_c_256_n N_Y_c_520_n 0.0197147f $X=3.85 $Y=1.765 $X2=0 $Y2=0
cc_240 N_A2_c_257_n N_Y_c_521_n 0.0120074f $X=4.35 $Y=1.765 $X2=0 $Y2=0
cc_241 N_A2_c_258_n N_Y_c_521_n 0.0120074f $X=4.8 $Y=1.765 $X2=0 $Y2=0
cc_242 A2 N_Y_c_521_n 0.0393874f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_243 N_A2_c_255_n N_Y_c_521_n 0.00146022f $X=5.25 $Y=1.557 $X2=0 $Y2=0
cc_244 N_A2_c_257_n N_Y_c_525_n 0.00888566f $X=4.35 $Y=1.765 $X2=0 $Y2=0
cc_245 N_A2_c_258_n N_Y_c_525_n 5.7112e-19 $X=4.8 $Y=1.765 $X2=0 $Y2=0
cc_246 A2 N_Y_c_525_n 0.0252603f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_247 N_A2_c_255_n N_Y_c_525_n 0.0018434f $X=5.25 $Y=1.557 $X2=0 $Y2=0
cc_248 N_A2_c_257_n N_Y_c_529_n 5.7112e-19 $X=4.35 $Y=1.765 $X2=0 $Y2=0
cc_249 N_A2_c_258_n N_Y_c_529_n 0.00891808f $X=4.8 $Y=1.765 $X2=0 $Y2=0
cc_250 N_A2_c_259_n N_Y_c_529_n 0.00964697f $X=5.25 $Y=1.765 $X2=0 $Y2=0
cc_251 A2 N_Y_c_529_n 0.0237597f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_252 N_A2_c_255_n N_Y_c_529_n 0.0016057f $X=5.25 $Y=1.557 $X2=0 $Y2=0
cc_253 N_A2_c_256_n Y 0.00907898f $X=3.85 $Y=1.765 $X2=0 $Y2=0
cc_254 A2 Y 0.0147816f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_255 N_A2_c_255_n Y 0.00656268f $X=5.25 $Y=1.557 $X2=0 $Y2=0
cc_256 N_A2_M1000_g N_Y_c_494_n 0.00579798f $X=3.975 $Y=0.74 $X2=0 $Y2=0
cc_257 A2 N_Y_c_494_n 0.00747454f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_258 N_A2_M1000_g N_A_27_74#_c_575_n 9.86481e-19 $X=3.975 $Y=0.74 $X2=0 $Y2=0
cc_259 N_A2_M1000_g N_A_27_74#_c_576_n 0.0148396f $X=3.975 $Y=0.74 $X2=0 $Y2=0
cc_260 N_A2_M1001_g N_A_27_74#_c_576_n 0.0130453f $X=4.405 $Y=0.74 $X2=0 $Y2=0
cc_261 A2 N_A_27_74#_c_576_n 0.0428095f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_262 N_A2_c_255_n N_A_27_74#_c_576_n 0.00408702f $X=5.25 $Y=1.557 $X2=0 $Y2=0
cc_263 N_A2_c_255_n N_A_27_74#_c_577_n 0.0031656f $X=5.25 $Y=1.557 $X2=0 $Y2=0
cc_264 N_A2_M1001_g N_A_27_74#_c_578_n 3.92313e-19 $X=4.405 $Y=0.74 $X2=0 $Y2=0
cc_265 N_A2_M1005_g N_A_27_74#_c_578_n 3.92313e-19 $X=4.835 $Y=0.74 $X2=0 $Y2=0
cc_266 N_A2_M1005_g N_A_27_74#_c_579_n 0.0130918f $X=4.835 $Y=0.74 $X2=0 $Y2=0
cc_267 N_A2_M1011_g N_A_27_74#_c_579_n 0.0136535f $X=5.265 $Y=0.74 $X2=0 $Y2=0
cc_268 A2 N_A_27_74#_c_579_n 0.073609f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_269 N_A2_c_255_n N_A_27_74#_c_579_n 0.00230191f $X=5.25 $Y=1.557 $X2=0 $Y2=0
cc_270 N_A2_M1011_g N_A_27_74#_c_580_n 0.00159319f $X=5.265 $Y=0.74 $X2=0 $Y2=0
cc_271 A2 N_A_27_74#_c_583_n 0.0146029f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_272 N_A2_c_255_n N_A_27_74#_c_583_n 0.00238948f $X=5.25 $Y=1.557 $X2=0 $Y2=0
cc_273 N_A2_M1000_g N_VGND_c_672_n 0.00383152f $X=3.975 $Y=0.74 $X2=0 $Y2=0
cc_274 N_A2_M1000_g N_VGND_c_673_n 0.00971294f $X=3.975 $Y=0.74 $X2=0 $Y2=0
cc_275 N_A2_M1001_g N_VGND_c_673_n 0.0103289f $X=4.405 $Y=0.74 $X2=0 $Y2=0
cc_276 N_A2_M1005_g N_VGND_c_673_n 4.71636e-19 $X=4.835 $Y=0.74 $X2=0 $Y2=0
cc_277 N_A2_M1001_g N_VGND_c_674_n 4.71636e-19 $X=4.405 $Y=0.74 $X2=0 $Y2=0
cc_278 N_A2_M1005_g N_VGND_c_674_n 0.0103289f $X=4.835 $Y=0.74 $X2=0 $Y2=0
cc_279 N_A2_M1011_g N_VGND_c_674_n 0.0133724f $X=5.265 $Y=0.74 $X2=0 $Y2=0
cc_280 N_A2_M1001_g N_VGND_c_677_n 0.00383152f $X=4.405 $Y=0.74 $X2=0 $Y2=0
cc_281 N_A2_M1005_g N_VGND_c_677_n 0.00383152f $X=4.835 $Y=0.74 $X2=0 $Y2=0
cc_282 N_A2_M1011_g N_VGND_c_678_n 0.00383152f $X=5.265 $Y=0.74 $X2=0 $Y2=0
cc_283 N_A2_M1000_g N_VGND_c_679_n 0.00757866f $X=3.975 $Y=0.74 $X2=0 $Y2=0
cc_284 N_A2_M1001_g N_VGND_c_679_n 0.0075754f $X=4.405 $Y=0.74 $X2=0 $Y2=0
cc_285 N_A2_M1005_g N_VGND_c_679_n 0.0075754f $X=4.835 $Y=0.74 $X2=0 $Y2=0
cc_286 N_A2_M1011_g N_VGND_c_679_n 0.00761198f $X=5.265 $Y=0.74 $X2=0 $Y2=0
cc_287 N_VPWR_c_331_n N_A_116_368#_c_399_n 0.0208862f $X=0.28 $Y=1.985 $X2=0
+ $Y2=0
cc_288 N_VPWR_c_331_n N_A_116_368#_c_400_n 0.0576605f $X=0.28 $Y=1.985 $X2=0
+ $Y2=0
cc_289 N_VPWR_c_332_n N_A_116_368#_c_400_n 0.0449718f $X=1.18 $Y=2.455 $X2=0
+ $Y2=0
cc_290 N_VPWR_c_335_n N_A_116_368#_c_400_n 0.014552f $X=1.095 $Y=3.33 $X2=0
+ $Y2=0
cc_291 N_VPWR_c_329_n N_A_116_368#_c_400_n 0.0119791f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_292 N_VPWR_M1009_d N_A_116_368#_c_418_n 0.00410876f $X=1.03 $Y=1.84 $X2=0
+ $Y2=0
cc_293 N_VPWR_c_332_n N_A_116_368#_c_418_n 0.0136682f $X=1.18 $Y=2.455 $X2=0
+ $Y2=0
cc_294 N_VPWR_c_332_n N_A_116_368#_c_401_n 0.0338656f $X=1.18 $Y=2.455 $X2=0
+ $Y2=0
cc_295 N_VPWR_c_333_n N_A_116_368#_c_401_n 0.0234974f $X=2.08 $Y=2.805 $X2=0
+ $Y2=0
cc_296 N_VPWR_c_337_n N_A_116_368#_c_401_n 0.014552f $X=1.995 $Y=3.33 $X2=0
+ $Y2=0
cc_297 N_VPWR_c_329_n N_A_116_368#_c_401_n 0.0119791f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_298 N_VPWR_M1012_d N_A_116_368#_c_402_n 0.00932188f $X=1.93 $Y=1.84 $X2=0
+ $Y2=0
cc_299 N_VPWR_M1014_s N_A_116_368#_c_402_n 0.0091206f $X=2.83 $Y=1.84 $X2=0
+ $Y2=0
cc_300 N_VPWR_c_333_n N_A_116_368#_c_402_n 0.0154248f $X=2.08 $Y=2.805 $X2=0
+ $Y2=0
cc_301 N_VPWR_c_334_n N_A_116_368#_c_402_n 0.0267445f $X=3.065 $Y=2.805 $X2=0
+ $Y2=0
cc_302 N_VPWR_c_334_n N_A_116_368#_c_404_n 0.0185066f $X=3.065 $Y=2.805 $X2=0
+ $Y2=0
cc_303 N_VPWR_c_339_n N_A_116_368#_c_405_n 0.0442078f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_304 N_VPWR_c_329_n N_A_116_368#_c_405_n 0.0250141f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_305 N_VPWR_c_334_n N_A_116_368#_c_406_n 0.0121618f $X=3.065 $Y=2.805 $X2=0
+ $Y2=0
cc_306 N_VPWR_c_339_n N_A_116_368#_c_406_n 0.0236039f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_307 N_VPWR_c_329_n N_A_116_368#_c_406_n 0.012761f $X=5.52 $Y=3.33 $X2=0 $Y2=0
cc_308 N_VPWR_c_339_n N_A_116_368#_c_407_n 0.0640155f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_309 N_VPWR_c_329_n N_A_116_368#_c_407_n 0.0357926f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_310 N_VPWR_c_332_n N_A_116_368#_c_433_n 0.0117758f $X=1.18 $Y=2.455 $X2=0
+ $Y2=0
cc_311 N_VPWR_c_339_n N_A_116_368#_c_409_n 0.0121867f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_312 N_VPWR_c_329_n N_A_116_368#_c_409_n 0.00660921f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_313 N_VPWR_M1014_s N_Y_c_495_n 0.00659121f $X=2.83 $Y=1.84 $X2=0 $Y2=0
cc_314 N_VPWR_c_331_n N_A_27_74#_c_571_n 0.00886035f $X=0.28 $Y=1.985 $X2=0
+ $Y2=0
cc_315 N_A_116_368#_c_402_n N_Y_M1013_d 0.00907897f $X=3.46 $Y=2.375 $X2=0 $Y2=0
cc_316 N_A_116_368#_c_405_n N_Y_M1002_s 0.00250873f $X=4.49 $Y=2.99 $X2=0 $Y2=0
cc_317 N_A_116_368#_c_407_n N_Y_M1017_s 0.00197722f $X=5.39 $Y=2.99 $X2=0 $Y2=0
cc_318 N_A_116_368#_c_423_n N_Y_c_495_n 0.00524731f $X=1.63 $Y=2.12 $X2=0 $Y2=0
cc_319 N_A_116_368#_c_402_n N_Y_c_495_n 0.0600659f $X=3.46 $Y=2.375 $X2=0 $Y2=0
cc_320 N_A_116_368#_M1002_d N_Y_c_520_n 4.9676e-19 $X=3.48 $Y=1.84 $X2=0 $Y2=0
cc_321 N_A_116_368#_c_403_n N_Y_c_520_n 0.00134458f $X=3.625 $Y=2.46 $X2=0 $Y2=0
cc_322 N_A_116_368#_M1015_d N_Y_c_521_n 0.00406069f $X=4.425 $Y=1.84 $X2=0 $Y2=0
cc_323 N_A_116_368#_c_484_p N_Y_c_521_n 0.0136682f $X=4.575 $Y=2.455 $X2=0 $Y2=0
cc_324 N_A_116_368#_c_405_n N_Y_c_525_n 0.018923f $X=4.49 $Y=2.99 $X2=0 $Y2=0
cc_325 N_A_116_368#_c_484_p N_Y_c_525_n 0.0289859f $X=4.575 $Y=2.455 $X2=0 $Y2=0
cc_326 N_A_116_368#_c_484_p N_Y_c_529_n 0.0289859f $X=4.575 $Y=2.455 $X2=0 $Y2=0
cc_327 N_A_116_368#_c_407_n N_Y_c_529_n 0.0160777f $X=5.39 $Y=2.99 $X2=0 $Y2=0
cc_328 N_A_116_368#_c_408_n N_Y_c_529_n 0.0533059f $X=5.475 $Y=2.115 $X2=0 $Y2=0
cc_329 N_A_116_368#_M1002_d Y 0.00608885f $X=3.48 $Y=1.84 $X2=0 $Y2=0
cc_330 N_A_116_368#_c_402_n Y 0.0104353f $X=3.46 $Y=2.375 $X2=0 $Y2=0
cc_331 N_A_116_368#_c_403_n Y 0.0227284f $X=3.625 $Y=2.46 $X2=0 $Y2=0
cc_332 N_Y_c_503_n N_A_27_74#_M1004_s 0.00328233f $X=3.22 $Y=0.925 $X2=0 $Y2=0
cc_333 N_Y_M1003_d N_A_27_74#_c_573_n 0.00176461f $X=2.305 $Y=0.37 $X2=0 $Y2=0
cc_334 N_Y_c_503_n N_A_27_74#_c_573_n 0.0035136f $X=3.22 $Y=0.925 $X2=0 $Y2=0
cc_335 N_Y_c_507_n N_A_27_74#_c_573_n 0.0138155f $X=2.445 $Y=0.8 $X2=0 $Y2=0
cc_336 N_Y_M1007_d N_A_27_74#_c_575_n 0.00176461f $X=3.165 $Y=0.37 $X2=0 $Y2=0
cc_337 N_Y_c_503_n N_A_27_74#_c_575_n 0.0035136f $X=3.22 $Y=0.925 $X2=0 $Y2=0
cc_338 N_Y_c_510_n N_A_27_74#_c_575_n 0.0165223f $X=3.305 $Y=0.8 $X2=0 $Y2=0
cc_339 N_Y_c_510_n N_A_27_74#_c_604_n 0.03026f $X=3.305 $Y=0.8 $X2=0 $Y2=0
cc_340 Y N_A_27_74#_c_577_n 0.0020972f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_341 N_Y_c_494_n N_A_27_74#_c_577_n 0.0135061f $X=3.525 $Y=1.55 $X2=0 $Y2=0
cc_342 N_Y_c_503_n N_A_27_74#_c_582_n 0.0160355f $X=3.22 $Y=0.925 $X2=0 $Y2=0
cc_343 N_Y_c_503_n N_VGND_c_679_n 0.00146755f $X=3.22 $Y=0.925 $X2=0 $Y2=0
cc_344 N_A_27_74#_c_570_n N_VGND_M1006_d 0.00176461f $X=1.055 $Y=1.065 $X2=-0.19
+ $Y2=-0.245
cc_345 N_A_27_74#_c_591_n N_VGND_M1019_d 0.00412925f $X=1.93 $Y=0.925 $X2=0
+ $Y2=0
cc_346 N_A_27_74#_c_576_n N_VGND_M1000_d 0.00176461f $X=4.535 $Y=1.095 $X2=0
+ $Y2=0
cc_347 N_A_27_74#_c_579_n N_VGND_M1005_d 0.00176461f $X=5.395 $Y=1.095 $X2=0
+ $Y2=0
cc_348 N_A_27_74#_c_569_n N_VGND_c_670_n 0.017215f $X=0.28 $Y=0.515 $X2=0 $Y2=0
cc_349 N_A_27_74#_c_570_n N_VGND_c_670_n 0.0170777f $X=1.055 $Y=1.065 $X2=0
+ $Y2=0
cc_350 N_A_27_74#_c_572_n N_VGND_c_670_n 0.0171736f $X=1.14 $Y=0.515 $X2=0 $Y2=0
cc_351 N_A_27_74#_c_572_n N_VGND_c_671_n 0.0121558f $X=1.14 $Y=0.515 $X2=0 $Y2=0
cc_352 N_A_27_74#_c_591_n N_VGND_c_671_n 0.0167779f $X=1.93 $Y=0.925 $X2=0 $Y2=0
cc_353 N_A_27_74#_c_574_n N_VGND_c_671_n 0.010561f $X=2.1 $Y=0.34 $X2=0 $Y2=0
cc_354 N_A_27_74#_c_573_n N_VGND_c_672_n 0.0384655f $X=2.71 $Y=0.34 $X2=0 $Y2=0
cc_355 N_A_27_74#_c_574_n N_VGND_c_672_n 0.0121867f $X=2.1 $Y=0.34 $X2=0 $Y2=0
cc_356 N_A_27_74#_c_575_n N_VGND_c_672_n 0.0522627f $X=3.675 $Y=0.34 $X2=0 $Y2=0
cc_357 N_A_27_74#_c_582_n N_VGND_c_672_n 0.0225055f $X=2.875 $Y=0.34 $X2=0 $Y2=0
cc_358 N_A_27_74#_c_575_n N_VGND_c_673_n 0.0112234f $X=3.675 $Y=0.34 $X2=0 $Y2=0
cc_359 N_A_27_74#_c_576_n N_VGND_c_673_n 0.0171619f $X=4.535 $Y=1.095 $X2=0
+ $Y2=0
cc_360 N_A_27_74#_c_578_n N_VGND_c_673_n 0.0182488f $X=4.62 $Y=0.515 $X2=0 $Y2=0
cc_361 N_A_27_74#_c_578_n N_VGND_c_674_n 0.0182488f $X=4.62 $Y=0.515 $X2=0 $Y2=0
cc_362 N_A_27_74#_c_579_n N_VGND_c_674_n 0.0171619f $X=5.395 $Y=1.095 $X2=0
+ $Y2=0
cc_363 N_A_27_74#_c_580_n N_VGND_c_674_n 0.0182902f $X=5.48 $Y=0.515 $X2=0 $Y2=0
cc_364 N_A_27_74#_c_569_n N_VGND_c_675_n 0.011066f $X=0.28 $Y=0.515 $X2=0 $Y2=0
cc_365 N_A_27_74#_c_572_n N_VGND_c_676_n 0.00749631f $X=1.14 $Y=0.515 $X2=0
+ $Y2=0
cc_366 N_A_27_74#_c_578_n N_VGND_c_677_n 0.00749631f $X=4.62 $Y=0.515 $X2=0
+ $Y2=0
cc_367 N_A_27_74#_c_580_n N_VGND_c_678_n 0.011066f $X=5.48 $Y=0.515 $X2=0 $Y2=0
cc_368 N_A_27_74#_c_569_n N_VGND_c_679_n 0.00915947f $X=0.28 $Y=0.515 $X2=0
+ $Y2=0
cc_369 N_A_27_74#_c_572_n N_VGND_c_679_n 0.0062048f $X=1.14 $Y=0.515 $X2=0 $Y2=0
cc_370 N_A_27_74#_c_591_n N_VGND_c_679_n 0.0120697f $X=1.93 $Y=0.925 $X2=0 $Y2=0
cc_371 N_A_27_74#_c_573_n N_VGND_c_679_n 0.0216792f $X=2.71 $Y=0.34 $X2=0 $Y2=0
cc_372 N_A_27_74#_c_574_n N_VGND_c_679_n 0.00660921f $X=2.1 $Y=0.34 $X2=0 $Y2=0
cc_373 N_A_27_74#_c_575_n N_VGND_c_679_n 0.0292284f $X=3.675 $Y=0.34 $X2=0 $Y2=0
cc_374 N_A_27_74#_c_578_n N_VGND_c_679_n 0.0062048f $X=4.62 $Y=0.515 $X2=0 $Y2=0
cc_375 N_A_27_74#_c_580_n N_VGND_c_679_n 0.00915947f $X=5.48 $Y=0.515 $X2=0
+ $Y2=0
cc_376 N_A_27_74#_c_582_n N_VGND_c_679_n 0.0123739f $X=2.875 $Y=0.34 $X2=0 $Y2=0
