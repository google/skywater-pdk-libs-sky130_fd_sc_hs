* File: sky130_fd_sc_hs__dfxbp_2.pex.spice
* Created: Tue Sep  1 20:00:51 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HS__DFXBP_2%CLK 1 3 4 6 7 11
c27 11 0 8.40497e-20 $X=0.42 $Y=1.385
r28 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.42
+ $Y=1.385 $X2=0.42 $Y2=1.385
r29 7 11 5.60648 $w=3.68e-07 $l=1.8e-07 $layer=LI1_cond $X=0.24 $Y=1.365
+ $X2=0.42 $Y2=1.365
r30 4 10 76.3385 $w=2.76e-07 $l=4.18091e-07 $layer=POLY_cond $X=0.505 $Y=1.765
+ $X2=0.425 $Y2=1.385
r31 4 6 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.505 $Y=1.765
+ $X2=0.505 $Y2=2.4
r32 1 10 38.7914 $w=2.76e-07 $l=1.96914e-07 $layer=POLY_cond $X=0.495 $Y=1.22
+ $X2=0.425 $Y2=1.385
r33 1 3 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=0.495 $Y=1.22 $X2=0.495
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HS__DFXBP_2%A_27_74# 1 2 7 9 10 12 13 15 17 18 20 21 23
+ 24 27 28 33 36 38 40 43 47 51 52 53 54 56 58 59 62 63 64 66 68 69 72 73 74 76
+ 79 82 84 89 93 94 98 107
c265 84 0 4.88492e-20 $X=0.97 $Y=1.385
c266 79 0 6.69395e-20 $X=6.075 $Y=0.365
c267 58 0 1.39925e-19 $X=0.84 $Y=1.72
c268 53 0 7.7167e-20 $X=0.755 $Y=1.805
c269 36 0 2.47898e-20 $X=3.12 $Y=1.165
c270 28 0 2.58209e-19 $X=6.09 $Y=1.245
c271 18 0 1.22911e-19 $X=3.435 $Y=2.15
c272 10 0 1.50442e-19 $X=1.14 $Y=1.22
r273 99 110 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.68 $Y=1.335
+ $X2=5.68 $Y2=1.5
r274 99 107 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=5.68 $Y=1.335
+ $X2=5.68 $Y2=1.245
r275 98 99 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.68
+ $Y=1.335 $X2=5.68 $Y2=1.335
r276 95 98 6.1738 $w=2.78e-07 $l=1.5e-07 $layer=LI1_cond $X=5.53 $Y=1.31
+ $X2=5.68 $Y2=1.31
r277 89 106 6.025 $w=3.6e-07 $l=4.5e-08 $layer=POLY_cond $X=3.39 $Y=1.942
+ $X2=3.435 $Y2=1.942
r278 89 104 36.15 $w=3.6e-07 $l=2.7e-07 $layer=POLY_cond $X=3.39 $Y=1.942
+ $X2=3.12 $Y2=1.942
r279 88 89 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.39
+ $Y=1.9 $X2=3.39 $Y2=1.9
r280 84 86 8.4794 $w=3.43e-07 $l=1.65e-07 $layer=LI1_cond $X=0.927 $Y=1.385
+ $X2=0.927 $Y2=1.55
r281 84 85 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.97
+ $Y=1.385 $X2=0.97 $Y2=1.385
r282 79 80 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.075
+ $Y=0.365 $X2=6.075 $Y2=0.365
r283 77 94 3.40559 $w=2.75e-07 $l=8.5e-08 $layer=LI1_cond $X=5.615 $Y=0.392
+ $X2=5.53 $Y2=0.392
r284 77 79 19.2772 $w=2.73e-07 $l=4.6e-07 $layer=LI1_cond $X=5.615 $Y=0.392
+ $X2=6.075 $Y2=0.392
r285 76 95 3.65648 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=5.53 $Y=1.17
+ $X2=5.53 $Y2=1.31
r286 75 94 3.11956 $w=1.7e-07 $l=1.38e-07 $layer=LI1_cond $X=5.53 $Y=0.53
+ $X2=5.53 $Y2=0.392
r287 75 76 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=5.53 $Y=0.53
+ $X2=5.53 $Y2=1.17
r288 73 94 3.40559 $w=2.75e-07 $l=8.5e-08 $layer=LI1_cond $X=5.445 $Y=0.392
+ $X2=5.53 $Y2=0.392
r289 73 74 26.4014 $w=2.73e-07 $l=6.3e-07 $layer=LI1_cond $X=5.445 $Y=0.392
+ $X2=4.815 $Y2=0.392
r290 71 74 7.32204 $w=2.75e-07 $l=1.75425e-07 $layer=LI1_cond $X=4.73 $Y=0.53
+ $X2=4.815 $Y2=0.392
r291 71 72 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=4.73 $Y=0.53
+ $X2=4.73 $Y2=0.78
r292 70 93 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.64 $Y=0.865
+ $X2=3.555 $Y2=0.865
r293 69 72 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.645 $Y=0.865
+ $X2=4.73 $Y2=0.78
r294 69 70 65.5668 $w=1.68e-07 $l=1.005e-06 $layer=LI1_cond $X=4.645 $Y=0.865
+ $X2=3.64 $Y2=0.865
r295 68 88 6.03661 $w=3.13e-07 $l=1.65e-07 $layer=LI1_cond $X=3.555 $Y=1.907
+ $X2=3.39 $Y2=1.907
r296 67 93 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.555 $Y=0.95
+ $X2=3.555 $Y2=0.865
r297 67 68 52.1925 $w=1.68e-07 $l=8e-07 $layer=LI1_cond $X=3.555 $Y=0.95
+ $X2=3.555 $Y2=1.75
r298 66 93 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.555 $Y=0.78
+ $X2=3.555 $Y2=0.865
r299 65 66 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=3.555 $Y=0.425
+ $X2=3.555 $Y2=0.78
r300 63 65 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.47 $Y=0.34
+ $X2=3.555 $Y2=0.425
r301 63 64 61.3262 $w=1.68e-07 $l=9.4e-07 $layer=LI1_cond $X=3.47 $Y=0.34
+ $X2=2.53 $Y2=0.34
r302 61 64 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.445 $Y=0.425
+ $X2=2.53 $Y2=0.34
r303 61 62 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=2.445 $Y=0.425
+ $X2=2.445 $Y2=0.73
r304 60 82 7.25401 $w=2.25e-07 $l=1.98605e-07 $layer=LI1_cond $X=1.1 $Y=0.815
+ $X2=0.927 $Y2=0.87
r305 59 62 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.36 $Y=0.815
+ $X2=2.445 $Y2=0.73
r306 59 60 82.2032 $w=1.68e-07 $l=1.26e-06 $layer=LI1_cond $X=2.36 $Y=0.815
+ $X2=1.1 $Y2=0.815
r307 58 86 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=0.84 $Y=1.72
+ $X2=0.84 $Y2=1.55
r308 56 84 0.233829 $w=3.43e-07 $l=7e-09 $layer=LI1_cond $X=0.927 $Y=1.378
+ $X2=0.927 $Y2=1.385
r309 55 82 0.140858 $w=3.45e-07 $l=1.4e-07 $layer=LI1_cond $X=0.927 $Y=1.01
+ $X2=0.927 $Y2=0.87
r310 55 56 12.2927 $w=3.43e-07 $l=3.68e-07 $layer=LI1_cond $X=0.927 $Y=1.01
+ $X2=0.927 $Y2=1.378
r311 53 58 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.755 $Y=1.805
+ $X2=0.84 $Y2=1.72
r312 53 54 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=0.755 $Y=1.805
+ $X2=0.445 $Y2=1.805
r313 51 82 7.25401 $w=2.25e-07 $l=1.72e-07 $layer=LI1_cond $X=0.755 $Y=0.87
+ $X2=0.927 $Y2=0.87
r314 51 52 12.7592 $w=2.78e-07 $l=3.1e-07 $layer=LI1_cond $X=0.755 $Y=0.87
+ $X2=0.445 $Y2=0.87
r315 47 49 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=0.28 $Y=1.985
+ $X2=0.28 $Y2=2.815
r316 45 54 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.28 $Y=1.89
+ $X2=0.445 $Y2=1.805
r317 45 47 3.31764 $w=3.28e-07 $l=9.5e-08 $layer=LI1_cond $X=0.28 $Y=1.89
+ $X2=0.28 $Y2=1.985
r318 41 52 6.87623 $w=2.8e-07 $l=2.24332e-07 $layer=LI1_cond $X=0.28 $Y=0.73
+ $X2=0.445 $Y2=0.87
r319 41 43 7.50834 $w=3.28e-07 $l=2.15e-07 $layer=LI1_cond $X=0.28 $Y=0.73
+ $X2=0.28 $Y2=0.515
r320 40 80 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=6.09 $Y=0.365
+ $X2=6.075 $Y2=0.365
r321 34 36 61.5319 $w=1.5e-07 $l=1.2e-07 $layer=POLY_cond $X=3 $Y=1.165 $X2=3.12
+ $Y2=1.165
r322 31 33 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=6.165 $Y=1.17
+ $X2=6.165 $Y2=0.85
r323 30 40 32.1775 $w=3.3e-07 $l=1.98997e-07 $layer=POLY_cond $X=6.165 $Y=0.53
+ $X2=6.09 $Y2=0.365
r324 30 33 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=6.165 $Y=0.53
+ $X2=6.165 $Y2=0.85
r325 29 107 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.845 $Y=1.245
+ $X2=5.68 $Y2=1.245
r326 28 31 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=6.09 $Y=1.245
+ $X2=6.165 $Y2=1.17
r327 28 29 125.628 $w=1.5e-07 $l=2.45e-07 $layer=POLY_cond $X=6.09 $Y=1.245
+ $X2=5.845 $Y2=1.245
r328 27 110 97.4255 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=5.59 $Y=1.69
+ $X2=5.59 $Y2=1.5
r329 25 38 7.1379 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=5.015 $Y=1.765
+ $X2=4.925 $Y2=1.765
r330 24 27 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.515 $Y=1.765
+ $X2=5.59 $Y2=1.69
r331 24 25 256.383 $w=1.5e-07 $l=5e-07 $layer=POLY_cond $X=5.515 $Y=1.765
+ $X2=5.015 $Y2=1.765
r332 21 38 110.989 $w=1.8e-07 $l=2.8e-07 $layer=POLY_cond $X=4.925 $Y=2.045
+ $X2=4.925 $Y2=1.765
r333 21 23 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=4.925 $Y=2.045
+ $X2=4.925 $Y2=2.54
r334 18 106 23.3057 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=3.435 $Y=2.15
+ $X2=3.435 $Y2=1.942
r335 18 20 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=3.435 $Y=2.15
+ $X2=3.435 $Y2=2.435
r336 17 104 23.3057 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.12 $Y=1.735
+ $X2=3.12 $Y2=1.942
r337 16 36 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.12 $Y=1.24
+ $X2=3.12 $Y2=1.165
r338 16 17 253.819 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=3.12 $Y=1.24
+ $X2=3.12 $Y2=1.735
r339 13 34 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3 $Y=1.09 $X2=3
+ $Y2=1.165
r340 13 15 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=3 $Y=1.09 $X2=3
+ $Y2=0.805
r341 10 85 38.5462 $w=3.19e-07 $l=2.20624e-07 $layer=POLY_cond $X=1.14 $Y=1.22
+ $X2=1.01 $Y2=1.385
r342 10 12 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.14 $Y=1.22
+ $X2=1.14 $Y2=0.74
r343 7 85 71.0321 $w=3.19e-07 $l=4.06571e-07 $layer=POLY_cond $X=0.955 $Y=1.765
+ $X2=1.01 $Y2=1.385
r344 7 9 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.955 $Y=1.765
+ $X2=0.955 $Y2=2.4
r345 2 49 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.815
r346 2 47 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=1.985
r347 1 43 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__DFXBP_2%D 1 3 4 6 10 11 12 14 15 22 31
c57 31 0 6.95252e-20 $X=2.16 $Y=1.665
c58 22 0 3.91626e-20 $X=2.21 $Y=1.29
c59 14 0 4.82751e-20 $X=2.16 $Y=1.295
c60 10 0 2.18369e-19 $X=1.99 $Y=2.19
r61 25 31 2.36399 $w=3.88e-07 $l=8e-08 $layer=LI1_cond $X=2.18 $Y=1.585 $X2=2.18
+ $Y2=1.665
r62 15 33 7.07103 $w=3.88e-07 $l=1.13e-07 $layer=LI1_cond $X=2.18 $Y=1.667
+ $X2=2.18 $Y2=1.78
r63 15 31 0.0590996 $w=3.88e-07 $l=2e-09 $layer=LI1_cond $X=2.18 $Y=1.667
+ $X2=2.18 $Y2=1.665
r64 15 25 0.0886495 $w=3.88e-07 $l=3e-09 $layer=LI1_cond $X=2.18 $Y=1.582
+ $X2=2.18 $Y2=1.585
r65 14 15 8.62855 $w=3.88e-07 $l=2.92e-07 $layer=LI1_cond $X=2.18 $Y=1.29
+ $X2=2.18 $Y2=1.582
r66 14 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.21
+ $Y=1.29 $X2=2.21 $Y2=1.29
r67 12 33 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=2.07 $Y=2.025
+ $X2=2.07 $Y2=1.78
r68 11 20 25.1593 $w=3.64e-07 $l=1.9e-07 $layer=POLY_cond $X=1.99 $Y=2.232
+ $X2=2.18 $Y2=2.232
r69 10 12 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=1.99 $Y=2.19
+ $X2=1.99 $Y2=2.025
r70 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.99
+ $Y=2.19 $X2=1.99 $Y2=2.19
r71 4 22 69.6867 $w=2.49e-07 $l=4.34741e-07 $layer=POLY_cond $X=2.57 $Y=1.125
+ $X2=2.21 $Y2=1.29
r72 4 6 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.57 $Y=1.125 $X2=2.57
+ $Y2=0.805
r73 1 20 23.572 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=2.18 $Y=2.44 $X2=2.18
+ $Y2=2.232
r74 1 3 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=2.18 $Y=2.44 $X2=2.18
+ $Y2=2.725
.ends

.subckt PM_SKY130_FD_SC_HS__DFXBP_2%A_206_368# 1 2 9 10 11 14 15 17 20 24 26 28
+ 30 33 35 38 39 43 49 52 56 57 60 64
c189 52 0 2.65941e-19 $X=1.65 $Y=1.65
c190 43 0 1.39777e-19 $X=6.04 $Y=2.07
c191 15 0 9.58637e-20 $X=2.715 $Y=2.15
c192 14 0 1.22505e-19 $X=2.715 $Y=2.06
r193 60 61 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=5.12 $Y=2.71
+ $X2=5.12 $Y2=2.88
r194 57 67 21.8577 $w=3.3e-07 $l=1.25e-07 $layer=POLY_cond $X=5.14 $Y=1.285
+ $X2=5.015 $Y2=1.285
r195 56 59 8.51388 $w=2.88e-07 $l=1.65e-07 $layer=LI1_cond $X=5.13 $Y=1.285
+ $X2=5.13 $Y2=1.45
r196 56 57 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.14
+ $Y=1.285 $X2=5.14 $Y2=1.285
r197 52 65 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=1.65 $Y=1.65 $X2=1.65
+ $Y2=1.74
r198 52 64 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.65 $Y=1.65
+ $X2=1.65 $Y2=1.485
r199 51 52 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.65
+ $Y=1.65 $X2=1.65 $Y2=1.65
r200 49 51 7.9006 $w=3.32e-07 $l=2.15e-07 $layer=LI1_cond $X=1.435 $Y=1.736
+ $X2=1.65 $Y2=1.736
r201 43 44 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.04
+ $Y=2.07 $X2=6.04 $Y2=2.07
r202 41 43 25.3188 $w=3.28e-07 $l=7.25e-07 $layer=LI1_cond $X=6.04 $Y=2.795
+ $X2=6.04 $Y2=2.07
r203 40 61 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.205 $Y=2.88
+ $X2=5.12 $Y2=2.88
r204 39 41 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=5.875 $Y=2.88
+ $X2=6.04 $Y2=2.795
r205 39 40 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.875 $Y=2.88
+ $X2=5.205 $Y2=2.88
r206 38 60 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=5.12 $Y=2.625
+ $X2=5.12 $Y2=2.71
r207 38 59 76.6578 $w=1.68e-07 $l=1.175e-06 $layer=LI1_cond $X=5.12 $Y=2.625
+ $X2=5.12 $Y2=1.45
r208 36 54 4.73278 $w=1.7e-07 $l=2.14114e-07 $layer=LI1_cond $X=1.44 $Y=2.71
+ $X2=1.267 $Y2=2.802
r209 35 60 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.035 $Y=2.71
+ $X2=5.12 $Y2=2.71
r210 35 36 234.54 $w=1.68e-07 $l=3.595e-06 $layer=LI1_cond $X=5.035 $Y=2.71
+ $X2=1.44 $Y2=2.71
r211 31 49 0.753319 $w=3.3e-07 $l=2.51e-07 $layer=LI1_cond $X=1.435 $Y=1.485
+ $X2=1.435 $Y2=1.736
r212 31 33 11.5244 $w=3.28e-07 $l=3.3e-07 $layer=LI1_cond $X=1.435 $Y=1.485
+ $X2=1.435 $Y2=1.155
r213 30 54 3.16114 $w=3.45e-07 $l=1.77e-07 $layer=LI1_cond $X=1.267 $Y=2.625
+ $X2=1.267 $Y2=2.802
r214 29 49 6.17349 $w=3.32e-07 $l=3.24298e-07 $layer=LI1_cond $X=1.267 $Y=1.987
+ $X2=1.435 $Y2=1.736
r215 29 47 3.19699 $w=3.32e-07 $l=8.79943e-08 $layer=LI1_cond $X=1.267 $Y=1.987
+ $X2=1.18 $Y2=1.985
r216 29 30 21.3118 $w=3.43e-07 $l=6.38e-07 $layer=LI1_cond $X=1.267 $Y=1.987
+ $X2=1.267 $Y2=2.625
r217 26 44 52.2586 $w=2.99e-07 $l=2.85044e-07 $layer=POLY_cond $X=5.965 $Y=2.32
+ $X2=6.04 $Y2=2.07
r218 26 28 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=5.965 $Y=2.32
+ $X2=5.965 $Y2=2.605
r219 22 67 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.015 $Y=1.12
+ $X2=5.015 $Y2=1.285
r220 22 24 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=5.015 $Y=1.12
+ $X2=5.015 $Y2=0.655
r221 18 20 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=3.51 $Y=0.255
+ $X2=3.51 $Y2=0.72
r222 15 17 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=2.715 $Y=2.15
+ $X2=2.715 $Y2=2.435
r223 14 15 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=2.715 $Y=2.06
+ $X2=2.715 $Y2=2.15
r224 13 14 95.2339 $w=1.8e-07 $l=2.45e-07 $layer=POLY_cond $X=2.715 $Y=1.815
+ $X2=2.715 $Y2=2.06
r225 12 65 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.815 $Y=1.74
+ $X2=1.65 $Y2=1.74
r226 11 13 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=2.625 $Y=1.74
+ $X2=2.715 $Y2=1.815
r227 11 12 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=2.625 $Y=1.74
+ $X2=1.815 $Y2=1.74
r228 9 18 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.435 $Y=0.18
+ $X2=3.51 $Y2=0.255
r229 9 10 835.809 $w=1.5e-07 $l=1.63e-06 $layer=POLY_cond $X=3.435 $Y=0.18
+ $X2=1.805 $Y2=0.18
r230 7 10 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.73 $Y=0.255
+ $X2=1.805 $Y2=0.18
r231 7 64 630.702 $w=1.5e-07 $l=1.23e-06 $layer=POLY_cond $X=1.73 $Y=0.255
+ $X2=1.73 $Y2=1.485
r232 2 54 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=1.03
+ $Y=1.84 $X2=1.18 $Y2=2.815
r233 2 47 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=1.03
+ $Y=1.84 $X2=1.18 $Y2=1.985
r234 1 33 182 $w=1.7e-07 $l=8.88214e-07 $layer=licon1_NDIFF $count=1 $X=1.215
+ $Y=0.37 $X2=1.435 $Y2=1.155
.ends

.subckt PM_SKY130_FD_SC_HS__DFXBP_2%A_753_284# 1 2 7 8 9 11 14 16 21 22
c57 14 0 3.89984e-20 $X=3.9 $Y=0.72
r58 22 24 1.25721 $w=2.73e-07 $l=3e-08 $layer=LI1_cond $X=4.73 $Y=2.317 $X2=4.7
+ $Y2=2.317
r59 21 29 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.73 $Y=1.45
+ $X2=4.73 $Y2=1.285
r60 21 22 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=4.73 $Y=1.45
+ $X2=4.73 $Y2=2.18
r61 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.975
+ $Y=1.255 $X2=3.975 $Y2=1.255
r62 16 29 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.645 $Y=1.285
+ $X2=4.73 $Y2=1.285
r63 16 18 23.3981 $w=3.28e-07 $l=6.7e-07 $layer=LI1_cond $X=4.645 $Y=1.285
+ $X2=3.975 $Y2=1.285
r64 12 19 38.532 $w=3.09e-07 $l=1.89222e-07 $layer=POLY_cond $X=3.9 $Y=1.09
+ $X2=3.952 $Y2=1.255
r65 12 14 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=3.9 $Y=1.09 $X2=3.9
+ $Y2=0.72
r66 9 11 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=3.855 $Y=2.15
+ $X2=3.855 $Y2=2.435
r67 8 9 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=3.855 $Y=2.06 $X2=3.855
+ $Y2=2.15
r68 7 19 48.107 $w=3.09e-07 $l=2.996e-07 $layer=POLY_cond $X=3.855 $Y=1.51
+ $X2=3.952 $Y2=1.255
r69 7 8 213.79 $w=1.8e-07 $l=5.5e-07 $layer=POLY_cond $X=3.855 $Y=1.51 $X2=3.855
+ $Y2=2.06
r70 2 24 600 $w=1.7e-07 $l=2.17428e-07 $layer=licon1_PDIFF $count=1 $X=4.55
+ $Y=2.12 $X2=4.7 $Y2=2.275
r71 1 29 182 $w=1.7e-07 $l=1.00902e-06 $layer=licon1_NDIFF $count=1 $X=4.5
+ $Y=0.38 $X2=4.72 $Y2=1.285
.ends

.subckt PM_SKY130_FD_SC_HS__DFXBP_2%A_558_445# 1 2 9 11 13 15 16 18 20 21 25 31
c78 18 0 1.01646e-19 $X=3.215 $Y=0.815
r79 31 34 8.46025 $w=3.18e-07 $l=1.65e-07 $layer=LI1_cond $X=4.315 $Y=1.795
+ $X2=4.315 $Y2=1.96
r80 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.32
+ $Y=1.795 $X2=4.32 $Y2=1.795
r81 25 34 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=4.24 $Y=2.285
+ $X2=4.24 $Y2=1.96
r82 21 23 1.95722 $w=1.68e-07 $l=3e-08 $layer=LI1_cond $X=3.055 $Y=2.37
+ $X2=3.085 $Y2=2.37
r83 20 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.155 $Y=2.37
+ $X2=4.24 $Y2=2.285
r84 20 23 69.8075 $w=1.68e-07 $l=1.07e-06 $layer=LI1_cond $X=4.155 $Y=2.37
+ $X2=3.085 $Y2=2.37
r85 16 26 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=3.175 $Y=1.495
+ $X2=2.97 $Y2=1.495
r86 16 18 27.4281 $w=2.48e-07 $l=5.95e-07 $layer=LI1_cond $X=3.175 $Y=1.41
+ $X2=3.175 $Y2=0.815
r87 15 21 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.97 $Y=2.285
+ $X2=3.055 $Y2=2.37
r88 14 26 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.97 $Y=1.58
+ $X2=2.97 $Y2=1.495
r89 14 15 45.9947 $w=1.68e-07 $l=7.05e-07 $layer=LI1_cond $X=2.97 $Y=1.58
+ $X2=2.97 $Y2=2.285
r90 11 32 50.2556 $w=3.62e-07 $l=3.02076e-07 $layer=POLY_cond $X=4.475 $Y=2.045
+ $X2=4.36 $Y2=1.795
r91 11 13 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=4.475 $Y=2.045
+ $X2=4.475 $Y2=2.54
r92 7 32 38.9379 $w=3.62e-07 $l=1.94808e-07 $layer=POLY_cond $X=4.425 $Y=1.63
+ $X2=4.36 $Y2=1.795
r93 7 9 499.947 $w=1.5e-07 $l=9.75e-07 $layer=POLY_cond $X=4.425 $Y=1.63
+ $X2=4.425 $Y2=0.655
r94 2 23 600 $w=1.7e-07 $l=3.60278e-07 $layer=licon1_PDIFF $count=1 $X=2.79
+ $Y=2.225 $X2=3.085 $Y2=2.37
r95 1 18 182 $w=1.7e-07 $l=2.81425e-07 $layer=licon1_NDIFF $count=1 $X=3.075
+ $Y=0.595 $X2=3.215 $Y2=0.815
.ends

.subckt PM_SKY130_FD_SC_HS__DFXBP_2%A_1290_102# 1 2 7 9 12 13 14 16 19 22 23 25
+ 26 30 32 34 35 37 40 43 44 45 49 50 51 54 60 62 65 66 70 74 77 78
c164 7 0 6.69395e-20 $X=6.525 $Y=1.17
r165 76 77 5.26419 $w=2.78e-07 $l=8.5e-08 $layer=LI1_cond $X=7.84 $Y=2.27
+ $X2=7.925 $Y2=2.27
r166 74 76 21.1967 $w=2.78e-07 $l=5.15e-07 $layer=LI1_cond $X=7.325 $Y=2.27
+ $X2=7.84 $Y2=2.27
r167 70 71 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.85
+ $Y=1.485 $X2=8.85 $Y2=1.485
r168 68 70 26.3665 $w=3.28e-07 $l=7.55e-07 $layer=LI1_cond $X=8.85 $Y=2.24
+ $X2=8.85 $Y2=1.485
r169 66 68 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=8.685 $Y=2.325
+ $X2=8.85 $Y2=2.24
r170 66 77 49.5829 $w=1.68e-07 $l=7.6e-07 $layer=LI1_cond $X=8.685 $Y=2.325
+ $X2=7.925 $Y2=2.325
r171 65 76 3.65648 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=7.84 $Y=2.13
+ $X2=7.84 $Y2=2.27
r172 64 65 41.1016 $w=1.68e-07 $l=6.3e-07 $layer=LI1_cond $X=7.84 $Y=1.5
+ $X2=7.84 $Y2=2.13
r173 63 78 5.16603 $w=2.5e-07 $l=1.60078e-07 $layer=LI1_cond $X=7.465 $Y=1.415
+ $X2=7.34 $Y2=1.335
r174 62 64 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.755 $Y=1.415
+ $X2=7.84 $Y2=1.5
r175 62 63 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=7.755 $Y=1.415
+ $X2=7.465 $Y2=1.415
r176 58 78 1.34256 $w=2.5e-07 $l=1.65e-07 $layer=LI1_cond $X=7.34 $Y=1.17
+ $X2=7.34 $Y2=1.335
r177 58 60 29.2721 $w=2.48e-07 $l=6.35e-07 $layer=LI1_cond $X=7.34 $Y=1.17
+ $X2=7.34 $Y2=0.535
r178 53 54 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.88
+ $Y=1.335 $X2=6.88 $Y2=1.335
r179 51 78 5.16603 $w=2.5e-07 $l=1.25e-07 $layer=LI1_cond $X=7.215 $Y=1.335
+ $X2=7.34 $Y2=1.335
r180 51 53 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=7.215 $Y=1.335
+ $X2=6.88 $Y2=1.335
r181 49 71 105.791 $w=3.3e-07 $l=6.05e-07 $layer=POLY_cond $X=9.455 $Y=1.485
+ $X2=8.85 $Y2=1.485
r182 49 50 5.03009 $w=3.3e-07 $l=1.15022e-07 $layer=POLY_cond $X=9.455 $Y=1.485
+ $X2=9.545 $Y2=1.542
r183 48 71 39.3438 $w=3.3e-07 $l=2.25e-07 $layer=POLY_cond $X=8.625 $Y=1.485
+ $X2=8.85 $Y2=1.485
r184 46 48 22.3608 $w=1.94e-07 $l=9e-08 $layer=POLY_cond $X=8.525 $Y=1.395
+ $X2=8.525 $Y2=1.485
r185 42 54 48.9612 $w=3.3e-07 $l=2.8e-07 $layer=POLY_cond $X=6.6 $Y=1.335
+ $X2=6.88 $Y2=1.335
r186 42 43 5.03009 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=6.6 $Y=1.335
+ $X2=6.525 $Y2=1.335
r187 38 50 37.0704 $w=1.5e-07 $l=2.29377e-07 $layer=POLY_cond $X=9.56 $Y=1.32
+ $X2=9.545 $Y2=1.542
r188 38 40 271.766 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=9.56 $Y=1.32
+ $X2=9.56 $Y2=0.79
r189 35 50 37.0704 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=9.545 $Y=1.765
+ $X2=9.545 $Y2=1.542
r190 35 37 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=9.545 $Y=1.765
+ $X2=9.545 $Y2=2.34
r191 32 48 72.1722 $w=1.94e-07 $l=2.84956e-07 $layer=POLY_cond $X=8.535 $Y=1.765
+ $X2=8.525 $Y2=1.485
r192 32 34 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=8.535 $Y=1.765
+ $X2=8.535 $Y2=2.4
r193 28 46 21.2393 $w=1.94e-07 $l=8.66025e-08 $layer=POLY_cond $X=8.5 $Y=1.32
+ $X2=8.525 $Y2=1.395
r194 28 30 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=8.5 $Y=1.32 $X2=8.5
+ $Y2=0.76
r195 27 45 6.66866 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=8.175 $Y=1.395
+ $X2=8.085 $Y2=1.395
r196 26 46 8.87375 $w=1.5e-07 $l=1e-07 $layer=POLY_cond $X=8.425 $Y=1.395
+ $X2=8.525 $Y2=1.395
r197 26 27 128.191 $w=1.5e-07 $l=2.5e-07 $layer=POLY_cond $X=8.425 $Y=1.395
+ $X2=8.175 $Y2=1.395
r198 23 25 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=8.085 $Y=1.765
+ $X2=8.085 $Y2=2.4
r199 22 23 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=8.085 $Y=1.675
+ $X2=8.085 $Y2=1.765
r200 21 45 18.8402 $w=1.65e-07 $l=7.5e-08 $layer=POLY_cond $X=8.085 $Y=1.47
+ $X2=8.085 $Y2=1.395
r201 21 22 79.6855 $w=1.8e-07 $l=2.05e-07 $layer=POLY_cond $X=8.085 $Y=1.47
+ $X2=8.085 $Y2=1.675
r202 17 45 18.8402 $w=1.65e-07 $l=8.21584e-08 $layer=POLY_cond $X=8.07 $Y=1.32
+ $X2=8.085 $Y2=1.395
r203 17 19 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=8.07 $Y=1.32
+ $X2=8.07 $Y2=0.76
r204 14 16 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=6.54 $Y=2.32
+ $X2=6.54 $Y2=2.605
r205 13 14 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=6.54 $Y=2.23 $X2=6.54
+ $Y2=2.32
r206 12 44 37.1337 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=6.54 $Y=1.83 $X2=6.54
+ $Y2=1.74
r207 12 13 155.484 $w=1.8e-07 $l=4e-07 $layer=POLY_cond $X=6.54 $Y=1.83 $X2=6.54
+ $Y2=2.23
r208 10 43 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.525 $Y=1.5
+ $X2=6.525 $Y2=1.335
r209 10 44 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=6.525 $Y=1.5
+ $X2=6.525 $Y2=1.74
r210 7 43 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.525 $Y=1.17
+ $X2=6.525 $Y2=1.335
r211 7 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=6.525 $Y=1.17
+ $X2=6.525 $Y2=0.85
r212 2 74 300 $w=1.7e-07 $l=2.38485e-07 $layer=licon1_PDIFF $count=2 $X=7.175
+ $Y=2.12 $X2=7.325 $Y2=2.295
r213 1 60 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=7.235
+ $Y=0.39 $X2=7.38 $Y2=0.535
.ends

.subckt PM_SKY130_FD_SC_HS__DFXBP_2%A_1000_424# 1 2 7 9 10 12 15 19 21 22 24 29
+ 35 37 38 39 42
c110 35 0 1.18432e-19 $X=6.1 $Y=0.825
r111 42 43 7.01942 $w=3.09e-07 $l=4.5e-08 $layer=POLY_cond $X=7.55 $Y=1.837
+ $X2=7.595 $Y2=1.837
r112 38 39 8.71257 $w=2.88e-07 $l=1.7e-07 $layer=LI1_cond $X=6.375 $Y=1.79
+ $X2=6.545 $Y2=1.79
r113 33 35 6.91466 $w=2.48e-07 $l=1.5e-07 $layer=LI1_cond $X=5.95 $Y=0.825
+ $X2=6.1 $Y2=0.825
r114 30 42 20.2783 $w=3.09e-07 $l=1.3e-07 $layer=POLY_cond $X=7.42 $Y=1.837
+ $X2=7.55 $Y2=1.837
r115 30 40 49.9159 $w=3.09e-07 $l=3.2e-07 $layer=POLY_cond $X=7.42 $Y=1.837
+ $X2=7.1 $Y2=1.837
r116 29 39 34.772 $w=2.88e-07 $l=8.75e-07 $layer=LI1_cond $X=7.42 $Y=1.815
+ $X2=6.545 $Y2=1.815
r117 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.42
+ $Y=1.795 $X2=7.42 $Y2=1.795
r118 26 37 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.185 $Y=1.705
+ $X2=6.1 $Y2=1.705
r119 26 38 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=6.185 $Y=1.705
+ $X2=6.375 $Y2=1.705
r120 24 37 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.1 $Y=1.62 $X2=6.1
+ $Y2=1.705
r121 23 35 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.1 $Y=0.95 $X2=6.1
+ $Y2=0.825
r122 23 24 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=6.1 $Y=0.95 $X2=6.1
+ $Y2=1.62
r123 21 37 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.015 $Y=1.705
+ $X2=6.1 $Y2=1.705
r124 21 22 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=6.015 $Y=1.705
+ $X2=5.705 $Y2=1.705
r125 17 22 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=5.54 $Y=1.79
+ $X2=5.705 $Y2=1.705
r126 17 19 26.1919 $w=3.28e-07 $l=7.5e-07 $layer=LI1_cond $X=5.54 $Y=1.79
+ $X2=5.54 $Y2=2.54
r127 13 43 19.6649 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=7.595 $Y=1.63
+ $X2=7.595 $Y2=1.837
r128 13 15 446.106 $w=1.5e-07 $l=8.7e-07 $layer=POLY_cond $X=7.595 $Y=1.63
+ $X2=7.595 $Y2=0.76
r129 10 42 19.6649 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=7.55 $Y=2.045
+ $X2=7.55 $Y2=1.837
r130 10 12 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=7.55 $Y=2.045
+ $X2=7.55 $Y2=2.54
r131 7 40 19.6649 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=7.1 $Y=2.045
+ $X2=7.1 $Y2=1.837
r132 7 9 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=7.1 $Y=2.045 $X2=7.1
+ $Y2=2.54
r133 2 19 600 $w=1.7e-07 $l=7.2e-07 $layer=licon1_PDIFF $count=1 $X=5 $Y=2.12
+ $X2=5.54 $Y2=2.54
r134 1 33 182 $w=1.7e-07 $l=1.04302e-06 $layer=licon1_NDIFF $count=1 $X=5.09
+ $Y=0.38 $X2=5.95 $Y2=0.785
.ends

.subckt PM_SKY130_FD_SC_HS__DFXBP_2%A_1835_368# 1 2 7 9 12 14 16 19 23 27 33 36
+ 40
c69 27 0 8.25183e-20 $X=9.32 $Y=1.985
c70 7 0 9.96991e-20 $X=10.08 $Y=1.765
r71 40 41 1.84439 $w=3.92e-07 $l=1.5e-08 $layer=POLY_cond $X=10.53 $Y=1.532
+ $X2=10.545 $Y2=1.532
r72 39 40 51.0281 $w=3.92e-07 $l=4.15e-07 $layer=POLY_cond $X=10.115 $Y=1.532
+ $X2=10.53 $Y2=1.532
r73 38 39 4.30357 $w=3.92e-07 $l=3.5e-08 $layer=POLY_cond $X=10.08 $Y=1.532
+ $X2=10.115 $Y2=1.532
r74 34 38 8.60714 $w=3.92e-07 $l=7e-08 $layer=POLY_cond $X=10.01 $Y=1.532
+ $X2=10.08 $Y2=1.532
r75 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.01
+ $Y=1.465 $X2=10.01 $Y2=1.465
r76 31 36 0.533013 $w=3.3e-07 $l=1.38e-07 $layer=LI1_cond $X=9.51 $Y=1.465
+ $X2=9.372 $Y2=1.465
r77 31 33 17.4613 $w=3.28e-07 $l=5e-07 $layer=LI1_cond $X=9.51 $Y=1.465
+ $X2=10.01 $Y2=1.465
r78 27 29 32.7294 $w=2.48e-07 $l=7.1e-07 $layer=LI1_cond $X=9.36 $Y=1.985
+ $X2=9.36 $Y2=2.695
r79 25 36 6.22203 $w=2.62e-07 $l=1.70895e-07 $layer=LI1_cond $X=9.36 $Y=1.63
+ $X2=9.372 $Y2=1.465
r80 25 27 16.3647 $w=2.48e-07 $l=3.55e-07 $layer=LI1_cond $X=9.36 $Y=1.63
+ $X2=9.36 $Y2=1.985
r81 21 36 6.22203 $w=2.62e-07 $l=1.65e-07 $layer=LI1_cond $X=9.372 $Y=1.3
+ $X2=9.372 $Y2=1.465
r82 21 23 19.4868 $w=2.73e-07 $l=4.65e-07 $layer=LI1_cond $X=9.372 $Y=1.3
+ $X2=9.372 $Y2=0.835
r83 17 41 25.3688 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=10.545 $Y=1.3
+ $X2=10.545 $Y2=1.532
r84 17 19 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=10.545 $Y=1.3
+ $X2=10.545 $Y2=0.74
r85 14 40 25.3688 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=10.53 $Y=1.765
+ $X2=10.53 $Y2=1.532
r86 14 16 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=10.53 $Y=1.765
+ $X2=10.53 $Y2=2.4
r87 10 39 25.3688 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=10.115 $Y=1.3
+ $X2=10.115 $Y2=1.532
r88 10 12 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=10.115 $Y=1.3
+ $X2=10.115 $Y2=0.74
r89 7 38 25.3688 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=10.08 $Y=1.765
+ $X2=10.08 $Y2=1.532
r90 7 9 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=10.08 $Y=1.765
+ $X2=10.08 $Y2=2.4
r91 2 29 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=9.175
+ $Y=1.84 $X2=9.32 $Y2=2.695
r92 2 27 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=9.175
+ $Y=1.84 $X2=9.32 $Y2=1.985
r93 1 23 182 $w=1.7e-07 $l=4.31451e-07 $layer=licon1_NDIFF $count=1 $X=9.2
+ $Y=0.47 $X2=9.345 $Y2=0.835
.ends

.subckt PM_SKY130_FD_SC_HS__DFXBP_2%VPWR 1 2 3 4 5 6 7 8 29 33 37 41 45 49 51 56
+ 57 59 60 61 68 80 88 92 98 103 106 108 115 118 122
r118 121 122 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.8 $Y=3.33
+ $X2=10.8 $Y2=3.33
r119 118 119 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.84 $Y=3.33
+ $X2=9.84 $Y2=3.33
r120 115 116 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r121 111 112 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r122 108 111 9.7783 $w=3.28e-07 $l=2.8e-07 $layer=LI1_cond $X=4.165 $Y=3.05
+ $X2=4.165 $Y2=3.33
r123 105 106 10.9518 $w=4.48e-07 $l=2.3e-07 $layer=LI1_cond $X=1.805 $Y=3.19
+ $X2=2.035 $Y2=3.19
r124 101 105 3.32244 $w=4.48e-07 $l=1.25e-07 $layer=LI1_cond $X=1.68 $Y=3.19
+ $X2=1.805 $Y2=3.19
r125 101 103 7.62935 $w=4.48e-07 $l=1.05e-07 $layer=LI1_cond $X=1.68 $Y=3.19
+ $X2=1.575 $Y2=3.19
r126 101 102 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r127 98 99 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r128 96 122 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.32 $Y=3.33
+ $X2=10.8 $Y2=3.33
r129 96 119 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.32 $Y=3.33
+ $X2=9.84 $Y2=3.33
r130 95 96 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.32 $Y=3.33
+ $X2=10.32 $Y2=3.33
r131 93 118 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=9.94 $Y=3.33
+ $X2=9.815 $Y2=3.33
r132 93 95 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=9.94 $Y=3.33
+ $X2=10.32 $Y2=3.33
r133 92 121 4.01252 $w=1.7e-07 $l=1.82e-07 $layer=LI1_cond $X=10.675 $Y=3.33
+ $X2=10.857 $Y2=3.33
r134 92 95 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=10.675 $Y=3.33
+ $X2=10.32 $Y2=3.33
r135 91 119 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.36 $Y=3.33
+ $X2=9.84 $Y2=3.33
r136 90 91 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.36 $Y=3.33
+ $X2=9.36 $Y2=3.33
r137 88 118 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=9.69 $Y=3.33
+ $X2=9.815 $Y2=3.33
r138 88 90 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=9.69 $Y=3.33
+ $X2=9.36 $Y2=3.33
r139 87 91 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=8.4 $Y=3.33
+ $X2=9.36 $Y2=3.33
r140 87 116 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=3.33
+ $X2=7.92 $Y2=3.33
r141 86 87 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=3.33 $X2=8.4
+ $Y2=3.33
r142 84 115 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.025 $Y=3.33
+ $X2=7.86 $Y2=3.33
r143 84 86 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=8.025 $Y=3.33
+ $X2=8.4 $Y2=3.33
r144 83 116 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=7.92 $Y2=3.33
r145 82 83 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r146 80 115 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.695 $Y=3.33
+ $X2=7.86 $Y2=3.33
r147 80 82 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=7.695 $Y=3.33
+ $X2=7.44 $Y2=3.33
r148 79 83 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=7.44 $Y2=3.33
r149 78 79 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r150 76 112 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=4.08 $Y2=3.33
r151 75 78 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=4.56 $Y=3.33
+ $X2=6.48 $Y2=3.33
r152 75 76 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r153 73 111 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.33 $Y=3.33
+ $X2=4.165 $Y2=3.33
r154 73 75 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=4.33 $Y=3.33
+ $X2=4.56 $Y2=3.33
r155 72 112 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=4.08 $Y2=3.33
r156 72 102 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.68 $Y2=3.33
r157 71 106 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=2.16 $Y=3.33
+ $X2=2.035 $Y2=3.33
r158 71 72 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r159 68 111 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4 $Y=3.33
+ $X2=4.165 $Y2=3.33
r160 68 71 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=4 $Y=3.33 $X2=2.16
+ $Y2=3.33
r161 67 102 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=1.68 $Y2=3.33
r162 67 99 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r163 66 103 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=1.2 $Y=3.33
+ $X2=1.575 $Y2=3.33
r164 66 67 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r165 64 98 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.895 $Y=3.33
+ $X2=0.77 $Y2=3.33
r166 64 66 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.895 $Y=3.33
+ $X2=1.2 $Y2=3.33
r167 61 79 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=6.48 $Y2=3.33
r168 61 76 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=4.56 $Y2=3.33
r169 59 86 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=8.595 $Y=3.33
+ $X2=8.4 $Y2=3.33
r170 59 60 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.595 $Y=3.33
+ $X2=8.76 $Y2=3.33
r171 58 90 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=8.925 $Y=3.33
+ $X2=9.36 $Y2=3.33
r172 58 60 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.925 $Y=3.33
+ $X2=8.76 $Y2=3.33
r173 56 78 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=6.6 $Y=3.33
+ $X2=6.48 $Y2=3.33
r174 56 57 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.6 $Y=3.33
+ $X2=6.765 $Y2=3.33
r175 55 82 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=6.93 $Y=3.33
+ $X2=7.44 $Y2=3.33
r176 55 57 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.93 $Y=3.33
+ $X2=6.765 $Y2=3.33
r177 51 54 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=10.8 $Y=1.985
+ $X2=10.8 $Y2=2.815
r178 49 121 3.13065 $w=2.5e-07 $l=1.09864e-07 $layer=LI1_cond $X=10.8 $Y=3.245
+ $X2=10.857 $Y2=3.33
r179 49 54 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=10.8 $Y=3.245
+ $X2=10.8 $Y2=2.815
r180 45 48 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=9.815 $Y=1.985
+ $X2=9.815 $Y2=2.815
r181 43 118 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=9.815 $Y=3.245
+ $X2=9.815 $Y2=3.33
r182 43 48 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=9.815 $Y=3.245
+ $X2=9.815 $Y2=2.815
r183 39 60 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.76 $Y=3.245
+ $X2=8.76 $Y2=3.33
r184 39 41 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=8.76 $Y=3.245
+ $X2=8.76 $Y2=2.78
r185 35 115 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.86 $Y=3.245
+ $X2=7.86 $Y2=3.33
r186 35 37 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=7.86 $Y=3.245
+ $X2=7.86 $Y2=2.78
r187 31 57 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.765 $Y=3.245
+ $X2=6.765 $Y2=3.33
r188 31 33 22.3504 $w=3.28e-07 $l=6.4e-07 $layer=LI1_cond $X=6.765 $Y=3.245
+ $X2=6.765 $Y2=2.605
r189 27 98 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.77 $Y=3.245
+ $X2=0.77 $Y2=3.33
r190 27 29 47.0197 $w=2.48e-07 $l=1.02e-06 $layer=LI1_cond $X=0.77 $Y=3.245
+ $X2=0.77 $Y2=2.225
r191 8 54 400 $w=1.7e-07 $l=1.04964e-06 $layer=licon1_PDIFF $count=1 $X=10.605
+ $Y=1.84 $X2=10.76 $Y2=2.815
r192 8 51 400 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_PDIFF $count=1 $X=10.605
+ $Y=1.84 $X2=10.76 $Y2=1.985
r193 7 48 600 $w=1.7e-07 $l=1.08616e-06 $layer=licon1_PDIFF $count=1 $X=9.62
+ $Y=1.84 $X2=9.855 $Y2=2.815
r194 7 45 300 $w=1.7e-07 $l=2.98831e-07 $layer=licon1_PDIFF $count=2 $X=9.62
+ $Y=1.84 $X2=9.855 $Y2=1.985
r195 6 41 600 $w=1.7e-07 $l=1.01223e-06 $layer=licon1_PDIFF $count=1 $X=8.61
+ $Y=1.84 $X2=8.76 $Y2=2.78
r196 5 37 600 $w=1.7e-07 $l=7.6857e-07 $layer=licon1_PDIFF $count=1 $X=7.625
+ $Y=2.12 $X2=7.86 $Y2=2.78
r197 4 33 600 $w=1.7e-07 $l=2.74955e-07 $layer=licon1_PDIFF $count=1 $X=6.615
+ $Y=2.395 $X2=6.765 $Y2=2.605
r198 3 108 600 $w=1.7e-07 $l=9.35147e-07 $layer=licon1_PDIFF $count=1 $X=3.93
+ $Y=2.225 $X2=4.165 $Y2=3.05
r199 2 105 600 $w=1.7e-07 $l=6.31328e-07 $layer=licon1_PDIFF $count=1 $X=1.595
+ $Y=2.515 $X2=1.805 $Y2=3.05
r200 1 29 300 $w=1.7e-07 $l=4.53845e-07 $layer=licon1_PDIFF $count=2 $X=0.58
+ $Y=1.84 $X2=0.73 $Y2=2.225
.ends

.subckt PM_SKY130_FD_SC_HS__DFXBP_2%A_451_503# 1 2 8 11 16 20
c37 16 0 1.22911e-19 $X=2.63 $Y=2.33
r38 18 20 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=2.63 $Y=1.155
+ $X2=2.785 $Y2=1.155
r39 14 16 6.45368 $w=2.48e-07 $l=1.4e-07 $layer=LI1_cond $X=2.49 $Y=2.33
+ $X2=2.63 $Y2=2.33
r40 9 20 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.785 $Y=1.07
+ $X2=2.785 $Y2=1.155
r41 9 11 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=2.785 $Y=1.07
+ $X2=2.785 $Y2=0.815
r42 8 16 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.63 $Y=2.205
+ $X2=2.63 $Y2=2.33
r43 7 18 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.63 $Y=1.24 $X2=2.63
+ $Y2=1.155
r44 7 8 62.9572 $w=1.68e-07 $l=9.65e-07 $layer=LI1_cond $X=2.63 $Y=1.24 $X2=2.63
+ $Y2=2.205
r45 2 14 600 $w=1.7e-07 $l=2.98831e-07 $layer=licon1_PDIFF $count=1 $X=2.255
+ $Y=2.515 $X2=2.49 $Y2=2.37
r46 1 11 182 $w=1.7e-07 $l=2.81425e-07 $layer=licon1_NDIFF $count=1 $X=2.645
+ $Y=0.595 $X2=2.785 $Y2=0.815
.ends

.subckt PM_SKY130_FD_SC_HS__DFXBP_2%Q 1 2 9 11
r21 11 17 9.96707 $w=3.68e-07 $l=3.2e-07 $layer=LI1_cond $X=8.33 $Y=1.665
+ $X2=8.33 $Y2=1.985
r22 11 14 3.97169 $w=3.68e-07 $l=1.15e-07 $layer=LI1_cond $X=8.33 $Y=1.665
+ $X2=8.33 $Y2=1.55
r23 9 14 38.3518 $w=3.03e-07 $l=1.015e-06 $layer=LI1_cond $X=8.297 $Y=0.535
+ $X2=8.297 $Y2=1.55
r24 2 17 600 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=8.16
+ $Y=1.84 $X2=8.31 $Y2=1.985
r25 1 9 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=8.145
+ $Y=0.39 $X2=8.285 $Y2=0.535
.ends

.subckt PM_SKY130_FD_SC_HS__DFXBP_2%Q_N 1 2 9 13 14 15 16 23 32
c30 32 0 9.96991e-20 $X=10.322 $Y=1.82
r31 21 23 1.04193 $w=3.63e-07 $l=3.3e-08 $layer=LI1_cond $X=10.322 $Y=2.002
+ $X2=10.322 $Y2=2.035
r32 15 16 11.6823 $w=3.63e-07 $l=3.7e-07 $layer=LI1_cond $X=10.322 $Y=2.405
+ $X2=10.322 $Y2=2.775
r33 14 21 0.820918 $w=3.63e-07 $l=2.6e-08 $layer=LI1_cond $X=10.322 $Y=1.976
+ $X2=10.322 $Y2=2.002
r34 14 32 8.24014 $w=3.63e-07 $l=1.56e-07 $layer=LI1_cond $X=10.322 $Y=1.976
+ $X2=10.322 $Y2=1.82
r35 14 15 10.8614 $w=3.63e-07 $l=3.44e-07 $layer=LI1_cond $X=10.322 $Y=2.061
+ $X2=10.322 $Y2=2.405
r36 14 23 0.820918 $w=3.63e-07 $l=2.6e-08 $layer=LI1_cond $X=10.322 $Y=2.061
+ $X2=10.322 $Y2=2.035
r37 13 32 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=10.42 $Y=1.13
+ $X2=10.42 $Y2=1.82
r38 7 13 8.64139 $w=3.38e-07 $l=1.7e-07 $layer=LI1_cond $X=10.335 $Y=0.96
+ $X2=10.335 $Y2=1.13
r39 7 9 15.0834 $w=3.38e-07 $l=4.45e-07 $layer=LI1_cond $X=10.335 $Y=0.96
+ $X2=10.335 $Y2=0.515
r40 2 14 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=10.155
+ $Y=1.84 $X2=10.305 $Y2=1.985
r41 2 16 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=10.155
+ $Y=1.84 $X2=10.305 $Y2=2.815
r42 1 9 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=10.19
+ $Y=0.37 $X2=10.33 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__DFXBP_2%VGND 1 2 3 4 5 6 7 8 27 31 33 37 41 45 49 53
+ 55 57 60 61 63 64 66 67 68 70 75 93 97 103 106 109 112 116
c141 31 0 6.63922e-20 $X=2.025 $Y=0.475
r142 115 116 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.8 $Y=0
+ $X2=10.8 $Y2=0
r143 112 113 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.84 $Y=0
+ $X2=9.84 $Y2=0
r144 109 110 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.08 $Y=0
+ $X2=4.08 $Y2=0
r145 107 110 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=2.16 $Y=0
+ $X2=4.08 $Y2=0
r146 106 107 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.16 $Y=0
+ $X2=2.16 $Y2=0
r147 103 104 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0
+ $X2=0.72 $Y2=0
r148 101 116 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.32 $Y=0
+ $X2=10.8 $Y2=0
r149 101 113 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.32 $Y=0
+ $X2=9.84 $Y2=0
r150 100 101 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.32 $Y=0
+ $X2=10.32 $Y2=0
r151 98 112 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=9.985 $Y=0
+ $X2=9.86 $Y2=0
r152 98 100 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=9.985 $Y=0
+ $X2=10.32 $Y2=0
r153 97 115 4.01252 $w=1.7e-07 $l=1.82e-07 $layer=LI1_cond $X=10.675 $Y=0
+ $X2=10.857 $Y2=0
r154 97 100 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=10.675 $Y=0
+ $X2=10.32 $Y2=0
r155 96 113 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.36 $Y=0
+ $X2=9.84 $Y2=0
r156 95 96 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.36 $Y=0 $X2=9.36
+ $Y2=0
r157 93 112 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=9.735 $Y=0
+ $X2=9.86 $Y2=0
r158 93 95 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=9.735 $Y=0
+ $X2=9.36 $Y2=0
r159 92 96 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=8.4 $Y=0 $X2=9.36
+ $Y2=0
r160 91 92 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r161 89 92 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=7.44 $Y=0 $X2=8.4
+ $Y2=0
r162 88 89 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.44 $Y=0 $X2=7.44
+ $Y2=0
r163 86 89 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.48 $Y=0 $X2=7.44
+ $Y2=0
r164 85 86 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6.48 $Y=0
+ $X2=6.48 $Y2=0
r165 83 110 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0
+ $X2=4.08 $Y2=0
r166 82 85 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=4.56 $Y=0 $X2=6.48
+ $Y2=0
r167 82 83 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.56 $Y=0
+ $X2=4.56 $Y2=0
r168 80 109 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=4.37 $Y=0 $X2=4.2
+ $Y2=0
r169 80 82 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=4.37 $Y=0 $X2=4.56
+ $Y2=0
r170 79 107 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0
+ $X2=2.16 $Y2=0
r171 79 104 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0
+ $X2=0.72 $Y2=0
r172 78 79 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r173 76 103 9.56655 $w=1.7e-07 $l=1.93e-07 $layer=LI1_cond $X=1.01 $Y=0
+ $X2=0.817 $Y2=0
r174 76 78 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.01 $Y=0 $X2=1.68
+ $Y2=0
r175 75 106 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.86 $Y=0
+ $X2=2.025 $Y2=0
r176 75 78 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=1.86 $Y=0 $X2=1.68
+ $Y2=0
r177 73 104 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0
+ $X2=0.72 $Y2=0
r178 72 73 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r179 70 103 9.56655 $w=1.7e-07 $l=1.92e-07 $layer=LI1_cond $X=0.625 $Y=0
+ $X2=0.817 $Y2=0
r180 70 72 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=0.625 $Y=0
+ $X2=0.24 $Y2=0
r181 68 86 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=6.48
+ $Y2=0
r182 68 83 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=4.56
+ $Y2=0
r183 66 91 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=8.62 $Y=0 $X2=8.4
+ $Y2=0
r184 66 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.62 $Y=0 $X2=8.785
+ $Y2=0
r185 65 95 26.7487 $w=1.68e-07 $l=4.1e-07 $layer=LI1_cond $X=8.95 $Y=0 $X2=9.36
+ $Y2=0
r186 65 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.95 $Y=0 $X2=8.785
+ $Y2=0
r187 63 88 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=7.645 $Y=0
+ $X2=7.44 $Y2=0
r188 63 64 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.645 $Y=0 $X2=7.81
+ $Y2=0
r189 62 91 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=7.975 $Y=0 $X2=8.4
+ $Y2=0
r190 62 64 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.975 $Y=0 $X2=7.81
+ $Y2=0
r191 60 85 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=6.655 $Y=0
+ $X2=6.48 $Y2=0
r192 60 61 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.655 $Y=0 $X2=6.82
+ $Y2=0
r193 59 88 29.6845 $w=1.68e-07 $l=4.55e-07 $layer=LI1_cond $X=6.985 $Y=0
+ $X2=7.44 $Y2=0
r194 59 61 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.985 $Y=0 $X2=6.82
+ $Y2=0
r195 55 115 3.13065 $w=2.5e-07 $l=1.09864e-07 $layer=LI1_cond $X=10.8 $Y=0.085
+ $X2=10.857 $Y2=0
r196 55 57 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=10.8 $Y=0.085
+ $X2=10.8 $Y2=0.515
r197 51 112 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=9.86 $Y=0.085
+ $X2=9.86 $Y2=0
r198 51 53 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=9.86 $Y=0.085
+ $X2=9.86 $Y2=0.515
r199 47 67 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.785 $Y=0.085
+ $X2=8.785 $Y2=0
r200 47 49 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=8.785 $Y=0.085
+ $X2=8.785 $Y2=0.535
r201 43 64 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.81 $Y=0.085
+ $X2=7.81 $Y2=0
r202 43 45 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=7.81 $Y=0.085
+ $X2=7.81 $Y2=0.535
r203 39 61 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.82 $Y=0.085
+ $X2=6.82 $Y2=0
r204 39 41 25.3188 $w=3.28e-07 $l=7.25e-07 $layer=LI1_cond $X=6.82 $Y=0.085
+ $X2=6.82 $Y2=0.81
r205 35 109 0.987631 $w=3.4e-07 $l=8.5e-08 $layer=LI1_cond $X=4.2 $Y=0.085
+ $X2=4.2 $Y2=0
r206 35 37 14.914 $w=3.38e-07 $l=4.4e-07 $layer=LI1_cond $X=4.2 $Y=0.085 $X2=4.2
+ $Y2=0.525
r207 34 106 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.19 $Y=0
+ $X2=2.025 $Y2=0
r208 33 109 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=4.03 $Y=0 $X2=4.2
+ $Y2=0
r209 33 34 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=4.03 $Y=0 $X2=2.19
+ $Y2=0
r210 29 106 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.025 $Y=0.085
+ $X2=2.025 $Y2=0
r211 29 31 13.6198 $w=3.28e-07 $l=3.9e-07 $layer=LI1_cond $X=2.025 $Y=0.085
+ $X2=2.025 $Y2=0.475
r212 25 103 1.35792 $w=3.85e-07 $l=8.5e-08 $layer=LI1_cond $X=0.817 $Y=0.085
+ $X2=0.817 $Y2=0
r213 25 27 9.27941 $w=3.83e-07 $l=3.1e-07 $layer=LI1_cond $X=0.817 $Y=0.085
+ $X2=0.817 $Y2=0.395
r214 8 57 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=10.62
+ $Y=0.37 $X2=10.76 $Y2=0.515
r215 7 53 91 $w=1.7e-07 $l=2.86618e-07 $layer=licon1_NDIFF $count=2 $X=9.635
+ $Y=0.47 $X2=9.9 $Y2=0.515
r216 6 49 91 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=2 $X=8.575
+ $Y=0.39 $X2=8.785 $Y2=0.535
r217 5 45 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=7.67
+ $Y=0.39 $X2=7.81 $Y2=0.535
r218 4 41 182 $w=1.7e-07 $l=2.92916e-07 $layer=licon1_NDIFF $count=1 $X=6.6
+ $Y=0.64 $X2=6.82 $Y2=0.81
r219 3 37 182 $w=1.7e-07 $l=2.32379e-07 $layer=licon1_NDIFF $count=1 $X=3.975
+ $Y=0.51 $X2=4.2 $Y2=0.525
r220 2 31 182 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=1 $X=1.88
+ $Y=0.33 $X2=2.025 $Y2=0.475
r221 1 27 182 $w=1.7e-07 $l=2.57196e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.37 $X2=0.815 $Y2=0.395
.ends

