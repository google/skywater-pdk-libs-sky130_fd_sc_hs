* File: sky130_fd_sc_hs__fah_1.pxi.spice
* Created: Tue Sep  1 20:05:39 2020
* 
x_PM_SKY130_FD_SC_HS__FAH_1%CI N_CI_c_284_n N_CI_M1010_g N_CI_c_285_n
+ N_CI_M1022_g CI N_CI_c_286_n PM_SKY130_FD_SC_HS__FAH_1%CI
x_PM_SKY130_FD_SC_HS__FAH_1%A_83_21# N_A_83_21#_M1001_d N_A_83_21#_M1023_d
+ N_A_83_21#_M1029_g N_A_83_21#_c_325_n N_A_83_21#_c_326_n N_A_83_21#_c_343_n
+ N_A_83_21#_M1021_g N_A_83_21#_c_327_n N_A_83_21#_c_328_n N_A_83_21#_c_329_n
+ N_A_83_21#_c_330_n N_A_83_21#_c_331_n N_A_83_21#_c_345_n N_A_83_21#_c_365_p
+ N_A_83_21#_c_366_p N_A_83_21#_c_346_n N_A_83_21#_c_347_n N_A_83_21#_c_332_n
+ N_A_83_21#_c_333_n N_A_83_21#_c_334_n N_A_83_21#_c_400_p N_A_83_21#_c_335_n
+ N_A_83_21#_c_336_n N_A_83_21#_c_337_n N_A_83_21#_c_338_n N_A_83_21#_c_376_p
+ N_A_83_21#_c_348_n N_A_83_21#_c_339_n N_A_83_21#_c_340_n N_A_83_21#_c_341_n
+ PM_SKY130_FD_SC_HS__FAH_1%A_83_21#
x_PM_SKY130_FD_SC_HS__FAH_1%A_410_58# N_A_410_58#_M1000_d N_A_410_58#_M1017_d
+ N_A_410_58#_M1006_g N_A_410_58#_c_514_n N_A_410_58#_c_515_n
+ N_A_410_58#_c_516_n N_A_410_58#_M1015_g N_A_410_58#_c_517_n
+ N_A_410_58#_c_518_n N_A_410_58#_c_550_n N_A_410_58#_c_519_n
+ N_A_410_58#_c_520_n N_A_410_58#_c_521_n N_A_410_58#_c_554_n
+ N_A_410_58#_c_522_n N_A_410_58#_c_523_n N_A_410_58#_c_524_n
+ N_A_410_58#_c_579_p N_A_410_58#_c_563_p PM_SKY130_FD_SC_HS__FAH_1%A_410_58#
x_PM_SKY130_FD_SC_HS__FAH_1%A_231_132# N_A_231_132#_M1010_d N_A_231_132#_M1012_d
+ N_A_231_132#_M1022_d N_A_231_132#_M1005_d N_A_231_132#_c_650_n
+ N_A_231_132#_M1028_g N_A_231_132#_c_651_n N_A_231_132#_M1024_g
+ N_A_231_132#_c_652_n N_A_231_132#_c_660_n N_A_231_132#_c_661_n
+ N_A_231_132#_c_662_n N_A_231_132#_c_695_n N_A_231_132#_c_663_n
+ N_A_231_132#_c_653_n N_A_231_132#_c_654_n N_A_231_132#_c_665_n
+ N_A_231_132#_c_704_n N_A_231_132#_c_655_n N_A_231_132#_c_667_n
+ N_A_231_132#_c_743_n N_A_231_132#_c_746_n N_A_231_132#_c_668_n
+ N_A_231_132#_c_677_n N_A_231_132#_c_656_n N_A_231_132#_c_713_n
+ N_A_231_132#_c_670_n N_A_231_132#_c_716_n N_A_231_132#_c_657_n
+ N_A_231_132#_c_658_n N_A_231_132#_c_672_n N_A_231_132#_c_724_n
+ N_A_231_132#_c_673_n PM_SKY130_FD_SC_HS__FAH_1%A_231_132#
x_PM_SKY130_FD_SC_HS__FAH_1%A_811_379# N_A_811_379#_M1002_d N_A_811_379#_M1018_d
+ N_A_811_379#_c_905_n N_A_811_379#_M1023_g N_A_811_379#_c_894_n
+ N_A_811_379#_c_895_n N_A_811_379#_c_896_n N_A_811_379#_M1000_g
+ N_A_811_379#_c_898_n N_A_811_379#_c_899_n N_A_811_379#_M1001_g
+ N_A_811_379#_c_908_n N_A_811_379#_c_909_n N_A_811_379#_M1017_g
+ N_A_811_379#_c_901_n N_A_811_379#_c_910_n N_A_811_379#_c_911_n
+ N_A_811_379#_c_902_n N_A_811_379#_c_903_n N_A_811_379#_c_904_n
+ N_A_811_379#_c_1010_p N_A_811_379#_c_914_n N_A_811_379#_c_915_n
+ N_A_811_379#_c_916_n N_A_811_379#_c_1016_p N_A_811_379#_c_1017_p
+ PM_SKY130_FD_SC_HS__FAH_1%A_811_379#
x_PM_SKY130_FD_SC_HS__FAH_1%A_1023_379# N_A_1023_379#_M1004_d
+ N_A_1023_379#_M1013_d N_A_1023_379#_M1005_g N_A_1023_379#_M1012_g
+ N_A_1023_379#_c_1117_n N_A_1023_379#_c_1118_n N_A_1023_379#_c_1100_n
+ N_A_1023_379#_M1020_g N_A_1023_379#_c_1101_n N_A_1023_379#_c_1102_n
+ N_A_1023_379#_c_1103_n N_A_1023_379#_c_1120_n N_A_1023_379#_c_1121_n
+ N_A_1023_379#_c_1122_n N_A_1023_379#_M1003_g N_A_1023_379#_c_1104_n
+ N_A_1023_379#_c_1105_n N_A_1023_379#_c_1106_n N_A_1023_379#_c_1107_n
+ N_A_1023_379#_c_1108_n N_A_1023_379#_c_1109_n N_A_1023_379#_c_1125_n
+ N_A_1023_379#_c_1166_n N_A_1023_379#_c_1110_n N_A_1023_379#_c_1111_n
+ N_A_1023_379#_c_1112_n N_A_1023_379#_c_1113_n N_A_1023_379#_c_1129_n
+ N_A_1023_379#_c_1130_n N_A_1023_379#_c_1114_n N_A_1023_379#_c_1115_n
+ PM_SKY130_FD_SC_HS__FAH_1%A_1023_379#
x_PM_SKY130_FD_SC_HS__FAH_1%A_879_55# N_A_879_55#_M1000_s N_A_879_55#_M1026_s
+ N_A_879_55#_M1003_d N_A_879_55#_c_1314_n N_A_879_55#_M1018_g
+ N_A_879_55#_M1004_g N_A_879_55#_c_1316_n N_A_879_55#_M1002_g
+ N_A_879_55#_c_1317_n N_A_879_55#_c_1334_n N_A_879_55#_M1013_g
+ N_A_879_55#_c_1318_n N_A_879_55#_c_1319_n N_A_879_55#_c_1336_n
+ N_A_879_55#_c_1320_n N_A_879_55#_c_1321_n N_A_879_55#_c_1322_n
+ N_A_879_55#_c_1323_n N_A_879_55#_c_1369_n N_A_879_55#_c_1324_n
+ N_A_879_55#_c_1353_n N_A_879_55#_c_1325_n N_A_879_55#_c_1326_n
+ N_A_879_55#_c_1327_n N_A_879_55#_c_1328_n N_A_879_55#_c_1414_n
+ N_A_879_55#_c_1329_n N_A_879_55#_c_1330_n N_A_879_55#_c_1331_n
+ PM_SKY130_FD_SC_HS__FAH_1%A_879_55#
x_PM_SKY130_FD_SC_HS__FAH_1%B N_B_c_1518_n N_B_M1031_g N_B_M1026_g N_B_c_1509_n
+ N_B_c_1520_n N_B_c_1521_n N_B_c_1522_n N_B_c_1510_n N_B_c_1524_n N_B_c_1525_n
+ N_B_c_1526_n N_B_M1019_g N_B_c_1528_n N_B_c_1511_n N_B_M1030_g N_B_M1027_g
+ N_B_c_1513_n N_B_c_1530_n N_B_c_1531_n N_B_c_1532_n N_B_M1016_g N_B_c_1514_n
+ N_B_c_1535_n N_B_c_1515_n B N_B_c_1517_n PM_SKY130_FD_SC_HS__FAH_1%B
x_PM_SKY130_FD_SC_HS__FAH_1%A_2342_48# N_A_2342_48#_M1011_d N_A_2342_48#_M1008_d
+ N_A_2342_48#_M1025_g N_A_2342_48#_c_1673_n N_A_2342_48#_M1007_g
+ N_A_2342_48#_c_1665_n N_A_2342_48#_c_1666_n N_A_2342_48#_c_1667_n
+ N_A_2342_48#_c_1675_n N_A_2342_48#_c_1668_n N_A_2342_48#_c_1669_n
+ N_A_2342_48#_c_1670_n N_A_2342_48#_c_1678_n N_A_2342_48#_c_1671_n
+ N_A_2342_48#_c_1672_n PM_SKY130_FD_SC_HS__FAH_1%A_2342_48#
x_PM_SKY130_FD_SC_HS__FAH_1%A N_A_M1014_g N_A_c_1750_n N_A_M1009_g N_A_c_1751_n
+ N_A_M1008_g N_A_M1011_g A N_A_c_1748_n N_A_c_1749_n
+ PM_SKY130_FD_SC_HS__FAH_1%A
x_PM_SKY130_FD_SC_HS__FAH_1%SUM N_SUM_M1029_s N_SUM_M1021_s SUM SUM SUM SUM SUM
+ N_SUM_c_1794_n PM_SKY130_FD_SC_HS__FAH_1%SUM
x_PM_SKY130_FD_SC_HS__FAH_1%VPWR N_VPWR_M1021_d N_VPWR_M1015_d N_VPWR_M1031_d
+ N_VPWR_M1007_d N_VPWR_M1009_d N_VPWR_c_1813_n N_VPWR_c_1814_n N_VPWR_c_1815_n
+ N_VPWR_c_1816_n N_VPWR_c_1817_n N_VPWR_c_1818_n N_VPWR_c_1819_n VPWR
+ N_VPWR_c_1820_n N_VPWR_c_1821_n N_VPWR_c_1822_n N_VPWR_c_1823_n
+ N_VPWR_c_1812_n N_VPWR_c_1825_n N_VPWR_c_1826_n N_VPWR_c_1827_n
+ N_VPWR_c_1828_n PM_SKY130_FD_SC_HS__FAH_1%VPWR
x_PM_SKY130_FD_SC_HS__FAH_1%COUT N_COUT_M1006_s N_COUT_M1015_s N_COUT_c_1944_n
+ N_COUT_c_1945_n N_COUT_c_1969_n N_COUT_c_1956_n N_COUT_c_1948_n
+ N_COUT_c_1958_n N_COUT_c_1949_n N_COUT_c_1950_n COUT
+ PM_SKY130_FD_SC_HS__FAH_1%COUT
x_PM_SKY130_FD_SC_HS__FAH_1%A_644_104# N_A_644_104#_M1028_d N_A_644_104#_M1020_d
+ N_A_644_104#_M1024_d N_A_644_104#_c_2019_n N_A_644_104#_c_2020_n
+ N_A_644_104#_c_2021_n N_A_644_104#_c_2022_n N_A_644_104#_c_2023_n
+ N_A_644_104#_c_2024_n N_A_644_104#_c_2025_n N_A_644_104#_c_2026_n
+ PM_SKY130_FD_SC_HS__FAH_1%A_644_104#
x_PM_SKY130_FD_SC_HS__FAH_1%A_1660_374# N_A_1660_374#_M1004_s
+ N_A_1660_374#_M1027_d N_A_1660_374#_M1018_s N_A_1660_374#_M1016_d
+ N_A_1660_374#_c_2122_n N_A_1660_374#_c_2123_n N_A_1660_374#_c_2124_n
+ N_A_1660_374#_c_2117_n N_A_1660_374#_c_2118_n N_A_1660_374#_c_2119_n
+ N_A_1660_374#_c_2120_n N_A_1660_374#_c_2132_n N_A_1660_374#_c_2121_n
+ PM_SKY130_FD_SC_HS__FAH_1%A_1660_374#
x_PM_SKY130_FD_SC_HS__FAH_1%A_1849_374# N_A_1849_374#_M1030_d
+ N_A_1849_374#_M1014_s N_A_1849_374#_M1019_d N_A_1849_374#_M1009_s
+ N_A_1849_374#_c_2208_n N_A_1849_374#_c_2209_n N_A_1849_374#_c_2210_n
+ N_A_1849_374#_c_2308_p N_A_1849_374#_c_2214_n N_A_1849_374#_c_2215_n
+ N_A_1849_374#_c_2211_n N_A_1849_374#_c_2216_n N_A_1849_374#_c_2217_n
+ N_A_1849_374#_c_2224_n N_A_1849_374#_c_2218_n N_A_1849_374#_c_2227_n
+ N_A_1849_374#_c_2219_n N_A_1849_374#_c_2220_n
+ PM_SKY130_FD_SC_HS__FAH_1%A_1849_374#
x_PM_SKY130_FD_SC_HS__FAH_1%VGND N_VGND_M1029_d N_VGND_M1006_d N_VGND_M1026_d
+ N_VGND_M1025_d N_VGND_M1014_d N_VGND_c_2317_n N_VGND_c_2318_n N_VGND_c_2319_n
+ N_VGND_c_2320_n N_VGND_c_2321_n N_VGND_c_2322_n N_VGND_c_2323_n
+ N_VGND_c_2324_n N_VGND_c_2325_n VGND N_VGND_c_2326_n N_VGND_c_2327_n
+ N_VGND_c_2328_n N_VGND_c_2329_n N_VGND_c_2330_n N_VGND_c_2331_n
+ N_VGND_c_2332_n N_VGND_c_2333_n PM_SKY130_FD_SC_HS__FAH_1%VGND
cc_1 VNB N_CI_c_284_n 0.0180743f $X=-0.19 $Y=-0.245 $X2=1.08 $Y2=1.41
cc_2 VNB N_CI_c_285_n 0.0250338f $X=-0.19 $Y=-0.245 $X2=1.185 $Y2=1.825
cc_3 VNB N_CI_c_286_n 0.00166349f $X=-0.19 $Y=-0.245 $X2=1.17 $Y2=1.575
cc_4 VNB N_A_83_21#_M1029_g 0.0303307f $X=-0.19 $Y=-0.245 $X2=1.17 $Y2=1.575
cc_5 VNB N_A_83_21#_c_325_n 0.00798644f $X=-0.19 $Y=-0.245 $X2=1.17 $Y2=1.575
cc_6 VNB N_A_83_21#_c_326_n 0.0137495f $X=-0.19 $Y=-0.245 $X2=1.17 $Y2=1.575
cc_7 VNB N_A_83_21#_c_327_n 0.0806199f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_A_83_21#_c_328_n 0.012806f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A_83_21#_c_329_n 0.0564028f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_83_21#_c_330_n 0.0165371f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_83_21#_c_331_n 0.00488345f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_83_21#_c_332_n 0.0022286f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_83_21#_c_333_n 0.0348622f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_83_21#_c_334_n 0.00357079f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_83_21#_c_335_n 0.0121451f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_83_21#_c_336_n 0.00711333f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_83_21#_c_337_n 0.00379131f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_83_21#_c_338_n 0.00355965f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_83_21#_c_339_n 0.0010811f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_83_21#_c_340_n 4.92773e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_83_21#_c_341_n 0.0157991f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_410_58#_M1006_g 0.0211593f $X=-0.19 $Y=-0.245 $X2=1.17 $Y2=1.575
cc_23 VNB N_A_410_58#_c_514_n 0.0256989f $X=-0.19 $Y=-0.245 $X2=1.17 $Y2=1.575
cc_24 VNB N_A_410_58#_c_515_n 0.00694057f $X=-0.19 $Y=-0.245 $X2=1.17 $Y2=1.575
cc_25 VNB N_A_410_58#_c_516_n 0.0352847f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_410_58#_c_517_n 0.00271393f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_410_58#_c_518_n 0.00898084f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_410_58#_c_519_n 0.0121646f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_410_58#_c_520_n 0.00120094f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_410_58#_c_521_n 0.00683747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_410_58#_c_522_n 0.0179487f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_410_58#_c_523_n 0.00776997f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_410_58#_c_524_n 0.00155485f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_231_132#_c_650_n 0.0203077f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_231_132#_c_651_n 0.0362838f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_231_132#_c_652_n 0.00185524f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_231_132#_c_653_n 0.00358783f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_231_132#_c_654_n 0.00114134f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_231_132#_c_655_n 0.00414548f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_231_132#_c_656_n 0.00336481f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_231_132#_c_657_n 0.0700957f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_231_132#_c_658_n 0.00460848f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_811_379#_c_894_n 0.0103399f $X=-0.19 $Y=-0.245 $X2=1.17 $Y2=1.575
cc_44 VNB N_A_811_379#_c_895_n 0.00119363f $X=-0.19 $Y=-0.245 $X2=1.17 $Y2=1.575
cc_45 VNB N_A_811_379#_c_896_n 0.01425f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_A_811_379#_M1000_g 0.0430538f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_811_379#_c_898_n 0.0639671f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_811_379#_c_899_n 0.012806f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A_811_379#_M1001_g 0.0312274f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_A_811_379#_c_901_n 0.0200101f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_A_811_379#_c_902_n 0.00466562f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_A_811_379#_c_903_n 0.00194757f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_A_811_379#_c_904_n 0.0201513f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_A_1023_379#_M1012_g 0.0427265f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_A_1023_379#_c_1100_n 0.0187336f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_A_1023_379#_c_1101_n 0.0254085f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_A_1023_379#_c_1102_n 0.00716314f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_A_1023_379#_c_1103_n 0.0144175f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_A_1023_379#_c_1104_n 0.00808887f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_A_1023_379#_c_1105_n 0.017736f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_A_1023_379#_c_1106_n 0.00340494f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_A_1023_379#_c_1107_n 0.055002f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_A_1023_379#_c_1108_n 0.00504695f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_A_1023_379#_c_1109_n 0.0408024f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_A_1023_379#_c_1110_n 5.75145e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_A_1023_379#_c_1111_n 0.0119849f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_A_1023_379#_c_1112_n 4.30713e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_A_1023_379#_c_1113_n 2.62982e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_A_1023_379#_c_1114_n 0.00166028f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_A_1023_379#_c_1115_n 0.00954575f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_A_879_55#_c_1314_n 0.0212863f $X=-0.19 $Y=-0.245 $X2=1.17 $Y2=1.575
cc_72 VNB N_A_879_55#_M1004_g 0.0290574f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_A_879_55#_c_1316_n 0.021028f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_A_879_55#_c_1317_n 0.0114151f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_A_879_55#_c_1318_n 0.0132907f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_A_879_55#_c_1319_n 0.0523923f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_A_879_55#_c_1320_n 0.00730213f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_A_879_55#_c_1321_n 0.00111269f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VNB N_A_879_55#_c_1322_n 0.0103511f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_A_879_55#_c_1323_n 0.00237617f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_81 VNB N_A_879_55#_c_1324_n 0.00503122f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_82 VNB N_A_879_55#_c_1325_n 0.00797922f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_83 VNB N_A_879_55#_c_1326_n 0.00328646f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_84 VNB N_A_879_55#_c_1327_n 0.00308636f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_85 VNB N_A_879_55#_c_1328_n 0.00385857f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_86 VNB N_A_879_55#_c_1329_n 0.00593009f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_87 VNB N_A_879_55#_c_1330_n 0.00129798f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_88 VNB N_A_879_55#_c_1331_n 0.035184f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_89 VNB N_B_M1026_g 0.0440237f $X=-0.19 $Y=-0.245 $X2=1.185 $Y2=2.4
cc_90 VNB N_B_c_1509_n 0.0285742f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_91 VNB N_B_c_1510_n 0.00342262f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_92 VNB N_B_c_1511_n 0.0194166f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_93 VNB N_B_M1027_g 0.0257958f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_94 VNB N_B_c_1513_n 0.00168574f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_95 VNB N_B_c_1514_n 0.00386338f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_96 VNB N_B_c_1515_n 0.0109549f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_97 VNB B 0.00591564f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_98 VNB N_B_c_1517_n 0.0481078f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_99 VNB N_A_2342_48#_c_1665_n 0.012362f $X=-0.19 $Y=-0.245 $X2=1.17 $Y2=1.665
cc_100 VNB N_A_2342_48#_c_1666_n 0.0194531f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_101 VNB N_A_2342_48#_c_1667_n 0.0143836f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_102 VNB N_A_2342_48#_c_1668_n 0.0339228f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_103 VNB N_A_2342_48#_c_1669_n 0.00491405f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_104 VNB N_A_2342_48#_c_1670_n 0.0517352f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_105 VNB N_A_2342_48#_c_1671_n 0.016963f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_106 VNB N_A_2342_48#_c_1672_n 0.0102948f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_107 VNB N_A_M1014_g 0.0420241f $X=-0.19 $Y=-0.245 $X2=1.08 $Y2=0.98
cc_108 VNB N_A_M1011_g 0.0451104f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_109 VNB N_A_c_1748_n 0.00503377f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_110 VNB N_A_c_1749_n 0.0275155f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_111 VNB N_SUM_c_1794_n 0.047753f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_112 VNB N_VPWR_c_1812_n 0.581632f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_113 VNB N_COUT_c_1944_n 0.00699039f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_114 VNB N_COUT_c_1945_n 8.00153e-19 $X=-0.19 $Y=-0.245 $X2=1.17 $Y2=1.575
cc_115 VNB COUT 0.00961274f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_116 VNB N_A_644_104#_c_2019_n 0.00268697f $X=-0.19 $Y=-0.245 $X2=1.17
+ $Y2=1.575
cc_117 VNB N_A_644_104#_c_2020_n 0.00308986f $X=-0.19 $Y=-0.245 $X2=1.17
+ $Y2=1.665
cc_118 VNB N_A_644_104#_c_2021_n 0.00386933f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_119 VNB N_A_644_104#_c_2022_n 0.0137142f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_120 VNB N_A_644_104#_c_2023_n 0.00447136f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_121 VNB N_A_644_104#_c_2024_n 0.0022959f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_122 VNB N_A_644_104#_c_2025_n 9.98694e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_123 VNB N_A_644_104#_c_2026_n 0.00348609f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_124 VNB N_A_1660_374#_c_2117_n 0.0028553f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_125 VNB N_A_1660_374#_c_2118_n 0.00256092f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_126 VNB N_A_1660_374#_c_2119_n 0.00376487f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_127 VNB N_A_1660_374#_c_2120_n 0.00976345f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_128 VNB N_A_1660_374#_c_2121_n 0.00859629f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_129 VNB N_A_1849_374#_c_2208_n 0.00915134f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_130 VNB N_A_1849_374#_c_2209_n 0.00213506f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_131 VNB N_A_1849_374#_c_2210_n 0.00741456f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_132 VNB N_A_1849_374#_c_2211_n 0.00833203f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_133 VNB N_VGND_c_2317_n 0.00776012f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_134 VNB N_VGND_c_2318_n 0.00967651f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_135 VNB N_VGND_c_2319_n 0.0121719f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_136 VNB N_VGND_c_2320_n 0.0121422f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_137 VNB N_VGND_c_2321_n 0.00975864f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_138 VNB N_VGND_c_2322_n 0.034344f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_139 VNB N_VGND_c_2323_n 0.00326991f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_140 VNB N_VGND_c_2324_n 0.0945588f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_141 VNB N_VGND_c_2325_n 0.00632279f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_142 VNB N_VGND_c_2326_n 0.0190364f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_143 VNB N_VGND_c_2327_n 0.122293f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_144 VNB N_VGND_c_2328_n 0.0205529f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_145 VNB N_VGND_c_2329_n 0.0189562f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_146 VNB N_VGND_c_2330_n 0.725957f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_147 VNB N_VGND_c_2331_n 0.0043669f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_148 VNB N_VGND_c_2332_n 0.0063135f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_149 VNB N_VGND_c_2333_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_150 VPB N_CI_c_285_n 0.0347055f $X=-0.19 $Y=1.66 $X2=1.185 $Y2=1.825
cc_151 VPB N_CI_c_286_n 0.0033715f $X=-0.19 $Y=1.66 $X2=1.17 $Y2=1.575
cc_152 VPB N_A_83_21#_c_326_n 9.92232e-19 $X=-0.19 $Y=1.66 $X2=1.17 $Y2=1.575
cc_153 VPB N_A_83_21#_c_343_n 0.0288209f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_154 VPB N_A_83_21#_c_331_n 6.18558e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_155 VPB N_A_83_21#_c_345_n 0.0891619f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_156 VPB N_A_83_21#_c_346_n 0.00692288f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_157 VPB N_A_83_21#_c_347_n 0.00309886f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_158 VPB N_A_83_21#_c_348_n 0.00227085f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_159 VPB N_A_83_21#_c_341_n 0.00204612f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_160 VPB N_A_410_58#_c_516_n 0.0345705f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_161 VPB N_A_410_58#_c_521_n 0.0013699f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_162 VPB N_A_231_132#_c_651_n 0.0292779f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_163 VPB N_A_231_132#_c_660_n 0.00634393f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_164 VPB N_A_231_132#_c_661_n 0.0146226f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_165 VPB N_A_231_132#_c_662_n 0.00296466f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_166 VPB N_A_231_132#_c_663_n 0.0117181f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_167 VPB N_A_231_132#_c_654_n 0.00188287f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_168 VPB N_A_231_132#_c_665_n 0.00695165f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_169 VPB N_A_231_132#_c_655_n 0.00104012f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_170 VPB N_A_231_132#_c_667_n 0.0183508f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_171 VPB N_A_231_132#_c_668_n 0.00401567f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_172 VPB N_A_231_132#_c_656_n 0.00196245f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_173 VPB N_A_231_132#_c_670_n 0.00229235f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_174 VPB N_A_231_132#_c_657_n 0.0208437f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_175 VPB N_A_231_132#_c_672_n 0.00195335f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_176 VPB N_A_231_132#_c_673_n 0.00585802f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_177 VPB N_A_811_379#_c_905_n 0.0198336f $X=-0.19 $Y=1.66 $X2=1.115 $Y2=1.58
cc_178 VPB N_A_811_379#_c_894_n 0.0236175f $X=-0.19 $Y=1.66 $X2=1.17 $Y2=1.575
cc_179 VPB N_A_811_379#_c_895_n 0.0087198f $X=-0.19 $Y=1.66 $X2=1.17 $Y2=1.575
cc_180 VPB N_A_811_379#_c_908_n 0.0265058f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_181 VPB N_A_811_379#_c_909_n 0.0174068f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_182 VPB N_A_811_379#_c_910_n 0.0100903f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_183 VPB N_A_811_379#_c_911_n 0.00232225f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_184 VPB N_A_811_379#_c_902_n 0.00354633f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_185 VPB N_A_811_379#_c_904_n 0.0202796f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_186 VPB N_A_811_379#_c_914_n 0.00632497f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_187 VPB N_A_811_379#_c_915_n 0.00127378f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_188 VPB N_A_811_379#_c_916_n 0.00328392f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_189 VPB N_A_1023_379#_M1005_g 0.0102152f $X=-0.19 $Y=1.66 $X2=1.17 $Y2=1.575
cc_190 VPB N_A_1023_379#_c_1117_n 0.130356f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_191 VPB N_A_1023_379#_c_1118_n 0.0181541f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_192 VPB N_A_1023_379#_c_1103_n 0.00564425f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_193 VPB N_A_1023_379#_c_1120_n 0.00712649f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_194 VPB N_A_1023_379#_c_1121_n 0.0144823f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_195 VPB N_A_1023_379#_c_1122_n 0.00652025f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_196 VPB N_A_1023_379#_M1003_g 0.00946396f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_197 VPB N_A_1023_379#_c_1104_n 0.012235f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_198 VPB N_A_1023_379#_c_1125_n 0.00282425f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_199 VPB N_A_1023_379#_c_1111_n 0.0256651f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_200 VPB N_A_1023_379#_c_1112_n 0.00112893f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_201 VPB N_A_1023_379#_c_1113_n 0.0011392f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_202 VPB N_A_1023_379#_c_1129_n 0.00432821f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_203 VPB N_A_1023_379#_c_1130_n 0.00250056f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_204 VPB N_A_1023_379#_c_1115_n 2.52545e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_205 VPB N_A_879_55#_c_1314_n 0.0315244f $X=-0.19 $Y=1.66 $X2=1.17 $Y2=1.575
cc_206 VPB N_A_879_55#_c_1317_n 0.00929566f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_207 VPB N_A_879_55#_c_1334_n 0.0176401f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_208 VPB N_A_879_55#_c_1318_n 0.0152791f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_209 VPB N_A_879_55#_c_1336_n 0.00441106f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_210 VPB N_A_879_55#_c_1325_n 9.38584e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_211 VPB N_A_879_55#_c_1328_n 0.00178762f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_212 VPB N_A_879_55#_c_1329_n 0.00271366f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_213 VPB N_A_879_55#_c_1331_n 0.0140276f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_214 VPB N_B_c_1518_n 0.0156123f $X=-0.19 $Y=1.66 $X2=1.08 $Y2=1.41
cc_215 VPB N_B_c_1509_n 0.0153125f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_216 VPB N_B_c_1520_n 0.0771697f $X=-0.19 $Y=1.66 $X2=1.17 $Y2=1.575
cc_217 VPB N_B_c_1521_n 0.0596925f $X=-0.19 $Y=1.66 $X2=1.17 $Y2=1.575
cc_218 VPB N_B_c_1522_n 0.012503f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_219 VPB N_B_c_1510_n 0.0064434f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_220 VPB N_B_c_1524_n 0.00890144f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_221 VPB N_B_c_1525_n 0.0156571f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_222 VPB N_B_c_1526_n 0.00712965f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_223 VPB N_B_M1019_g 0.009998f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_224 VPB N_B_c_1528_n 0.146828f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_225 VPB N_B_c_1513_n 0.00767391f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_226 VPB N_B_c_1530_n 0.00794125f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_227 VPB N_B_c_1531_n 0.0154667f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_228 VPB N_B_c_1532_n 0.0057433f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_229 VPB N_B_M1016_g 0.00862886f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_230 VPB N_B_c_1514_n 0.00457093f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_231 VPB N_B_c_1535_n 0.00898665f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_232 VPB N_B_c_1517_n 0.00362115f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_233 VPB N_A_2342_48#_c_1673_n 0.0179881f $X=-0.19 $Y=1.66 $X2=1.17 $Y2=1.575
cc_234 VPB N_A_2342_48#_c_1665_n 0.0136717f $X=-0.19 $Y=1.66 $X2=1.17 $Y2=1.665
cc_235 VPB N_A_2342_48#_c_1675_n 0.0356154f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_236 VPB N_A_2342_48#_c_1669_n 0.00166579f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_237 VPB N_A_2342_48#_c_1670_n 0.0165636f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_238 VPB N_A_2342_48#_c_1678_n 0.00707313f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_239 VPB N_A_2342_48#_c_1671_n 0.014684f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_240 VPB N_A_c_1750_n 0.0178278f $X=-0.19 $Y=1.66 $X2=1.185 $Y2=2.4
cc_241 VPB N_A_c_1751_n 0.0206916f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_242 VPB N_A_c_1748_n 0.00317944f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_243 VPB N_A_c_1749_n 0.0405103f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_244 VPB N_SUM_c_1794_n 0.0539442f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_245 VPB N_VPWR_c_1813_n 0.00811871f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_246 VPB N_VPWR_c_1814_n 0.0198489f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_247 VPB N_VPWR_c_1815_n 0.00172518f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_248 VPB N_VPWR_c_1816_n 0.0126508f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_249 VPB N_VPWR_c_1817_n 0.00886117f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_250 VPB N_VPWR_c_1818_n 0.0915399f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_251 VPB N_VPWR_c_1819_n 0.00651392f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_252 VPB N_VPWR_c_1820_n 0.0504123f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_253 VPB N_VPWR_c_1821_n 0.102433f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_254 VPB N_VPWR_c_1822_n 0.0215588f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_255 VPB N_VPWR_c_1823_n 0.0190763f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_256 VPB N_VPWR_c_1812_n 0.120131f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_257 VPB N_VPWR_c_1825_n 0.0233111f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_258 VPB N_VPWR_c_1826_n 0.0142668f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_259 VPB N_VPWR_c_1827_n 0.00631825f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_260 VPB N_VPWR_c_1828_n 0.0047828f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_261 VPB N_COUT_c_1944_n 0.00355802f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_262 VPB N_COUT_c_1948_n 0.00242228f $X=-0.19 $Y=1.66 $X2=1.17 $Y2=1.665
cc_263 VPB N_COUT_c_1949_n 0.00260505f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_264 VPB N_COUT_c_1950_n 0.0242637f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_265 VPB N_A_644_104#_c_2022_n 0.00489558f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_266 VPB N_A_644_104#_c_2023_n 0.00214659f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_267 VPB N_A_644_104#_c_2024_n 0.00166693f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_268 VPB N_A_644_104#_c_2025_n 0.00329977f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_269 VPB N_A_644_104#_c_2026_n 0.00917256f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_270 VPB N_A_1660_374#_c_2122_n 0.00111308f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_271 VPB N_A_1660_374#_c_2123_n 0.0505497f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_272 VPB N_A_1660_374#_c_2124_n 5.85313e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_273 VPB N_A_1660_374#_c_2118_n 0.00527952f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_274 VPB N_A_1660_374#_c_2121_n 0.00204935f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_275 VPB N_A_1849_374#_c_2208_n 0.0103766f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_276 VPB N_A_1849_374#_c_2209_n 0.00677983f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_277 VPB N_A_1849_374#_c_2214_n 0.00545578f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_278 VPB N_A_1849_374#_c_2215_n 0.00135635f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_279 VPB N_A_1849_374#_c_2216_n 0.0145105f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_280 VPB N_A_1849_374#_c_2217_n 0.0105002f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_281 VPB N_A_1849_374#_c_2218_n 0.00381488f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_282 VPB N_A_1849_374#_c_2219_n 0.00251594f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_283 VPB N_A_1849_374#_c_2220_n 0.00828332f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_284 N_CI_c_284_n N_A_83_21#_M1029_g 0.0175596f $X=1.08 $Y=1.41 $X2=0 $Y2=0
cc_285 N_CI_c_284_n N_A_83_21#_c_325_n 0.00393369f $X=1.08 $Y=1.41 $X2=0 $Y2=0
cc_286 N_CI_c_285_n N_A_83_21#_c_326_n 0.00393369f $X=1.185 $Y=1.825 $X2=0 $Y2=0
cc_287 N_CI_c_285_n N_A_83_21#_c_343_n 0.0151046f $X=1.185 $Y=1.825 $X2=0 $Y2=0
cc_288 N_CI_c_284_n N_A_83_21#_c_327_n 0.00721051f $X=1.08 $Y=1.41 $X2=0 $Y2=0
cc_289 N_CI_c_284_n N_A_83_21#_c_329_n 0.0199086f $X=1.08 $Y=1.41 $X2=0 $Y2=0
cc_290 N_CI_c_285_n N_A_83_21#_c_345_n 0.0115737f $X=1.185 $Y=1.825 $X2=0 $Y2=0
cc_291 N_CI_c_284_n N_A_83_21#_c_341_n 4.26869e-19 $X=1.08 $Y=1.41 $X2=0 $Y2=0
cc_292 N_CI_c_285_n N_A_83_21#_c_341_n 0.0115388f $X=1.185 $Y=1.825 $X2=0 $Y2=0
cc_293 N_CI_c_286_n N_A_83_21#_c_341_n 3.30521e-19 $X=1.17 $Y=1.575 $X2=0 $Y2=0
cc_294 N_CI_c_284_n N_A_231_132#_c_652_n 0.00290104f $X=1.08 $Y=1.41 $X2=0 $Y2=0
cc_295 N_CI_c_285_n N_A_231_132#_c_652_n 0.00112718f $X=1.185 $Y=1.825 $X2=0
+ $Y2=0
cc_296 N_CI_c_286_n N_A_231_132#_c_652_n 0.0131004f $X=1.17 $Y=1.575 $X2=0 $Y2=0
cc_297 N_CI_c_285_n N_A_231_132#_c_677_n 0.00246364f $X=1.185 $Y=1.825 $X2=0
+ $Y2=0
cc_298 N_CI_c_286_n N_A_231_132#_c_677_n 7.02654e-19 $X=1.17 $Y=1.575 $X2=0
+ $Y2=0
cc_299 N_CI_c_284_n N_A_231_132#_c_656_n 0.00124432f $X=1.08 $Y=1.41 $X2=0 $Y2=0
cc_300 N_CI_c_285_n N_A_231_132#_c_656_n 0.00396448f $X=1.185 $Y=1.825 $X2=0
+ $Y2=0
cc_301 N_CI_c_286_n N_A_231_132#_c_656_n 0.0279725f $X=1.17 $Y=1.575 $X2=0 $Y2=0
cc_302 N_CI_c_284_n N_SUM_c_1794_n 0.00110666f $X=1.08 $Y=1.41 $X2=0 $Y2=0
cc_303 N_CI_c_285_n N_SUM_c_1794_n 4.03567e-19 $X=1.185 $Y=1.825 $X2=0 $Y2=0
cc_304 N_CI_c_285_n N_VPWR_c_1813_n 0.00208117f $X=1.185 $Y=1.825 $X2=0 $Y2=0
cc_305 N_CI_c_285_n N_VPWR_c_1820_n 8.69849e-19 $X=1.185 $Y=1.825 $X2=0 $Y2=0
cc_306 N_CI_c_284_n N_COUT_c_1944_n 0.00985011f $X=1.08 $Y=1.41 $X2=0 $Y2=0
cc_307 N_CI_c_285_n N_COUT_c_1944_n 0.00194352f $X=1.185 $Y=1.825 $X2=0 $Y2=0
cc_308 N_CI_c_286_n N_COUT_c_1944_n 0.0279727f $X=1.17 $Y=1.575 $X2=0 $Y2=0
cc_309 N_CI_c_284_n N_COUT_c_1945_n 0.0134584f $X=1.08 $Y=1.41 $X2=0 $Y2=0
cc_310 N_CI_c_286_n N_COUT_c_1945_n 0.00365255f $X=1.17 $Y=1.575 $X2=0 $Y2=0
cc_311 N_CI_c_285_n N_COUT_c_1956_n 0.0234422f $X=1.185 $Y=1.825 $X2=0 $Y2=0
cc_312 N_CI_c_285_n N_COUT_c_1948_n 0.00262083f $X=1.185 $Y=1.825 $X2=0 $Y2=0
cc_313 N_CI_c_285_n N_COUT_c_1958_n 0.00603264f $X=1.185 $Y=1.825 $X2=0 $Y2=0
cc_314 N_CI_c_286_n N_COUT_c_1958_n 0.00933956f $X=1.17 $Y=1.575 $X2=0 $Y2=0
cc_315 N_CI_c_285_n N_COUT_c_1950_n 0.0103484f $X=1.185 $Y=1.825 $X2=0 $Y2=0
cc_316 N_CI_c_284_n COUT 0.00403824f $X=1.08 $Y=1.41 $X2=0 $Y2=0
cc_317 N_CI_c_284_n N_VGND_c_2317_n 4.52739e-19 $X=1.08 $Y=1.41 $X2=0 $Y2=0
cc_318 N_CI_c_284_n N_VGND_c_2330_n 9.59665e-19 $X=1.08 $Y=1.41 $X2=0 $Y2=0
cc_319 N_A_83_21#_c_338_n N_A_410_58#_M1000_d 0.00261255f $X=5.885 $Y=0.68
+ $X2=-0.19 $Y2=-0.245
cc_320 N_A_83_21#_c_339_n N_A_410_58#_M1000_d 0.00315942f $X=4.96 $Y=0.68
+ $X2=-0.19 $Y2=-0.245
cc_321 N_A_83_21#_c_329_n N_A_410_58#_M1006_g 0.0250002f $X=1.62 $Y=1.235 $X2=0
+ $Y2=0
cc_322 N_A_83_21#_c_330_n N_A_410_58#_M1006_g 0.00553712f $X=1.735 $Y=1.31 $X2=0
+ $Y2=0
cc_323 N_A_83_21#_c_331_n N_A_410_58#_M1006_g 0.0122745f $X=2.01 $Y=1.86 $X2=0
+ $Y2=0
cc_324 N_A_83_21#_c_365_p N_A_410_58#_M1006_g 0.00625054f $X=2.595 $Y=0.985
+ $X2=0 $Y2=0
cc_325 N_A_83_21#_c_366_p N_A_410_58#_M1006_g 0.00907316f $X=2.175 $Y=0.985
+ $X2=0 $Y2=0
cc_326 N_A_83_21#_c_332_n N_A_410_58#_M1006_g 0.00460897f $X=2.68 $Y=0.9 $X2=0
+ $Y2=0
cc_327 N_A_83_21#_c_365_p N_A_410_58#_c_514_n 0.0086249f $X=2.595 $Y=0.985 $X2=0
+ $Y2=0
cc_328 N_A_83_21#_c_331_n N_A_410_58#_c_515_n 0.0071983f $X=2.01 $Y=1.86 $X2=0
+ $Y2=0
cc_329 N_A_83_21#_c_345_n N_A_410_58#_c_515_n 0.00694652f $X=2.01 $Y=1.86 $X2=0
+ $Y2=0
cc_330 N_A_83_21#_c_341_n N_A_410_58#_c_515_n 0.00553712f $X=1.917 $Y=1.695
+ $X2=0 $Y2=0
cc_331 N_A_83_21#_c_331_n N_A_410_58#_c_516_n 0.00494231f $X=2.01 $Y=1.86 $X2=0
+ $Y2=0
cc_332 N_A_83_21#_c_345_n N_A_410_58#_c_516_n 0.0166513f $X=2.01 $Y=1.86 $X2=0
+ $Y2=0
cc_333 N_A_83_21#_c_365_p N_A_410_58#_c_516_n 0.00167876f $X=2.595 $Y=0.985
+ $X2=0 $Y2=0
cc_334 N_A_83_21#_c_346_n N_A_410_58#_c_516_n 0.0182423f $X=3.155 $Y=2.28 $X2=0
+ $Y2=0
cc_335 N_A_83_21#_c_376_p N_A_410_58#_c_516_n 0.00196271f $X=3.24 $Y=2.28 $X2=0
+ $Y2=0
cc_336 N_A_83_21#_c_341_n N_A_410_58#_c_516_n 0.00222905f $X=1.917 $Y=1.695
+ $X2=0 $Y2=0
cc_337 N_A_83_21#_c_365_p N_A_410_58#_c_517_n 0.0138309f $X=2.595 $Y=0.985 $X2=0
+ $Y2=0
cc_338 N_A_83_21#_c_332_n N_A_410_58#_c_517_n 0.00973281f $X=2.68 $Y=0.9 $X2=0
+ $Y2=0
cc_339 N_A_83_21#_c_333_n N_A_410_58#_c_518_n 0.0577593f $X=4.115 $Y=0.34 $X2=0
+ $Y2=0
cc_340 N_A_83_21#_c_335_n N_A_410_58#_c_518_n 0.0134759f $X=4.2 $Y=0.755 $X2=0
+ $Y2=0
cc_341 N_A_83_21#_c_337_n N_A_410_58#_c_518_n 9.36976e-19 $X=4.285 $Y=0.84 $X2=0
+ $Y2=0
cc_342 N_A_83_21#_c_332_n N_A_410_58#_c_550_n 0.0138309f $X=2.68 $Y=0.9 $X2=0
+ $Y2=0
cc_343 N_A_83_21#_c_333_n N_A_410_58#_c_550_n 0.0106895f $X=4.115 $Y=0.34 $X2=0
+ $Y2=0
cc_344 N_A_83_21#_c_337_n N_A_410_58#_c_519_n 0.0134759f $X=4.285 $Y=0.84 $X2=0
+ $Y2=0
cc_345 N_A_83_21#_M1023_d N_A_410_58#_c_521_n 0.00212057f $X=4.22 $Y=2.12 $X2=0
+ $Y2=0
cc_346 N_A_83_21#_M1023_d N_A_410_58#_c_554_n 0.00222934f $X=4.22 $Y=2.12 $X2=0
+ $Y2=0
cc_347 N_A_83_21#_c_331_n N_A_410_58#_c_522_n 0.0191017f $X=2.01 $Y=1.86 $X2=0
+ $Y2=0
cc_348 N_A_83_21#_c_365_p N_A_410_58#_c_522_n 0.0224262f $X=2.595 $Y=0.985 $X2=0
+ $Y2=0
cc_349 N_A_83_21#_c_346_n N_A_410_58#_c_522_n 0.00861567f $X=3.155 $Y=2.28 $X2=0
+ $Y2=0
cc_350 N_A_83_21#_c_333_n N_A_410_58#_c_523_n 0.00488227f $X=4.115 $Y=0.34 $X2=0
+ $Y2=0
cc_351 N_A_83_21#_c_336_n N_A_410_58#_c_523_n 0.0386802f $X=4.875 $Y=0.84 $X2=0
+ $Y2=0
cc_352 N_A_83_21#_c_337_n N_A_410_58#_c_523_n 0.0143396f $X=4.285 $Y=0.84 $X2=0
+ $Y2=0
cc_353 N_A_83_21#_c_339_n N_A_410_58#_c_523_n 0.0087105f $X=4.96 $Y=0.68 $X2=0
+ $Y2=0
cc_354 N_A_83_21#_c_338_n N_A_410_58#_c_524_n 0.00741596f $X=5.885 $Y=0.68 $X2=0
+ $Y2=0
cc_355 N_A_83_21#_c_338_n N_A_231_132#_M1012_d 0.00175311f $X=5.885 $Y=0.68
+ $X2=0 $Y2=0
cc_356 N_A_83_21#_c_365_p N_A_231_132#_c_650_n 9.82061e-19 $X=2.595 $Y=0.985
+ $X2=0 $Y2=0
cc_357 N_A_83_21#_c_332_n N_A_231_132#_c_650_n 0.0065908f $X=2.68 $Y=0.9 $X2=0
+ $Y2=0
cc_358 N_A_83_21#_c_333_n N_A_231_132#_c_650_n 0.0066613f $X=4.115 $Y=0.34 $X2=0
+ $Y2=0
cc_359 N_A_83_21#_c_400_p N_A_231_132#_c_651_n 0.0114233f $X=4.205 $Y=2.37 $X2=0
+ $Y2=0
cc_360 N_A_83_21#_c_348_n N_A_231_132#_c_651_n 0.00159552f $X=4.37 $Y=2.255
+ $X2=0 $Y2=0
cc_361 N_A_83_21#_c_329_n N_A_231_132#_c_652_n 0.00716755f $X=1.62 $Y=1.235
+ $X2=0 $Y2=0
cc_362 N_A_83_21#_c_331_n N_A_231_132#_c_652_n 0.013814f $X=2.01 $Y=1.86 $X2=0
+ $Y2=0
cc_363 N_A_83_21#_c_345_n N_A_231_132#_c_660_n 0.00718697f $X=2.01 $Y=1.86 $X2=0
+ $Y2=0
cc_364 N_A_83_21#_c_347_n N_A_231_132#_c_660_n 0.0136282f $X=2.175 $Y=2.28 $X2=0
+ $Y2=0
cc_365 N_A_83_21#_c_345_n N_A_231_132#_c_661_n 0.00932304f $X=2.01 $Y=1.86 $X2=0
+ $Y2=0
cc_366 N_A_83_21#_c_346_n N_A_231_132#_c_661_n 0.0422491f $X=3.155 $Y=2.28 $X2=0
+ $Y2=0
cc_367 N_A_83_21#_c_347_n N_A_231_132#_c_661_n 0.0263722f $X=2.175 $Y=2.28 $X2=0
+ $Y2=0
cc_368 N_A_83_21#_c_346_n N_A_231_132#_c_695_n 0.00902987f $X=3.155 $Y=2.28
+ $X2=0 $Y2=0
cc_369 N_A_83_21#_c_400_p N_A_231_132#_c_695_n 0.00677804f $X=4.205 $Y=2.37
+ $X2=0 $Y2=0
cc_370 N_A_83_21#_c_376_p N_A_231_132#_c_695_n 0.0110829f $X=3.24 $Y=2.28 $X2=0
+ $Y2=0
cc_371 N_A_83_21#_M1023_d N_A_231_132#_c_663_n 0.010127f $X=4.22 $Y=2.12 $X2=0
+ $Y2=0
cc_372 N_A_83_21#_c_400_p N_A_231_132#_c_663_n 0.0179855f $X=4.205 $Y=2.37 $X2=0
+ $Y2=0
cc_373 N_A_83_21#_c_348_n N_A_231_132#_c_663_n 0.0204134f $X=4.37 $Y=2.255 $X2=0
+ $Y2=0
cc_374 N_A_83_21#_M1023_d N_A_231_132#_c_654_n 0.0165703f $X=4.22 $Y=2.12 $X2=0
+ $Y2=0
cc_375 N_A_83_21#_c_348_n N_A_231_132#_c_654_n 0.0481667f $X=4.37 $Y=2.255 $X2=0
+ $Y2=0
cc_376 N_A_83_21#_M1023_d N_A_231_132#_c_665_n 0.00821661f $X=4.22 $Y=2.12 $X2=0
+ $Y2=0
cc_377 N_A_83_21#_M1001_d N_A_231_132#_c_704_n 0.00345021f $X=5.84 $Y=0.625
+ $X2=0 $Y2=0
cc_378 N_A_83_21#_c_338_n N_A_231_132#_c_704_n 0.00585443f $X=5.885 $Y=0.68
+ $X2=0 $Y2=0
cc_379 N_A_83_21#_c_340_n N_A_231_132#_c_704_n 0.0203544f $X=6.05 $Y=0.68 $X2=0
+ $Y2=0
cc_380 N_A_83_21#_M1001_d N_A_231_132#_c_655_n 7.06785e-19 $X=5.84 $Y=0.625
+ $X2=0 $Y2=0
cc_381 N_A_83_21#_c_345_n N_A_231_132#_c_677_n 0.00502438f $X=2.01 $Y=1.86 $X2=0
+ $Y2=0
cc_382 N_A_83_21#_c_330_n N_A_231_132#_c_656_n 0.00674676f $X=1.735 $Y=1.31
+ $X2=0 $Y2=0
cc_383 N_A_83_21#_c_331_n N_A_231_132#_c_656_n 0.0708186f $X=2.01 $Y=1.86 $X2=0
+ $Y2=0
cc_384 N_A_83_21#_c_345_n N_A_231_132#_c_656_n 0.00626205f $X=2.01 $Y=1.86 $X2=0
+ $Y2=0
cc_385 N_A_83_21#_c_341_n N_A_231_132#_c_656_n 0.00575716f $X=1.917 $Y=1.695
+ $X2=0 $Y2=0
cc_386 N_A_83_21#_c_346_n N_A_231_132#_c_713_n 0.00812609f $X=3.155 $Y=2.28
+ $X2=0 $Y2=0
cc_387 N_A_83_21#_c_400_p N_A_231_132#_c_670_n 0.00848586f $X=4.205 $Y=2.37
+ $X2=0 $Y2=0
cc_388 N_A_83_21#_c_348_n N_A_231_132#_c_670_n 0.00312083f $X=4.37 $Y=2.255
+ $X2=0 $Y2=0
cc_389 N_A_83_21#_c_400_p N_A_231_132#_c_716_n 0.00167184f $X=4.205 $Y=2.37
+ $X2=0 $Y2=0
cc_390 N_A_83_21#_c_400_p N_A_231_132#_c_657_n 0.00104274f $X=4.205 $Y=2.37
+ $X2=0 $Y2=0
cc_391 N_A_83_21#_c_336_n N_A_231_132#_c_657_n 2.68583e-19 $X=4.875 $Y=0.84
+ $X2=0 $Y2=0
cc_392 N_A_83_21#_c_337_n N_A_231_132#_c_657_n 9.39832e-19 $X=4.285 $Y=0.84
+ $X2=0 $Y2=0
cc_393 N_A_83_21#_c_400_p N_A_231_132#_c_658_n 9.53902e-19 $X=4.205 $Y=2.37
+ $X2=0 $Y2=0
cc_394 N_A_83_21#_c_348_n N_A_231_132#_c_658_n 0.0143188f $X=4.37 $Y=2.255 $X2=0
+ $Y2=0
cc_395 N_A_83_21#_M1023_d N_A_231_132#_c_672_n 0.00526596f $X=4.22 $Y=2.12 $X2=0
+ $Y2=0
cc_396 N_A_83_21#_c_348_n N_A_231_132#_c_672_n 4.25819e-19 $X=4.37 $Y=2.255
+ $X2=0 $Y2=0
cc_397 N_A_83_21#_c_338_n N_A_231_132#_c_724_n 0.0158698f $X=5.885 $Y=0.68 $X2=0
+ $Y2=0
cc_398 N_A_83_21#_c_400_p N_A_811_379#_c_905_n 0.011771f $X=4.205 $Y=2.37 $X2=0
+ $Y2=0
cc_399 N_A_83_21#_c_348_n N_A_811_379#_c_905_n 0.0111326f $X=4.37 $Y=2.255 $X2=0
+ $Y2=0
cc_400 N_A_83_21#_c_348_n N_A_811_379#_c_894_n 0.00815895f $X=4.37 $Y=2.255
+ $X2=0 $Y2=0
cc_401 N_A_83_21#_c_335_n N_A_811_379#_M1000_g 0.00302956f $X=4.2 $Y=0.755 $X2=0
+ $Y2=0
cc_402 N_A_83_21#_c_336_n N_A_811_379#_M1000_g 0.0103248f $X=4.875 $Y=0.84 $X2=0
+ $Y2=0
cc_403 N_A_83_21#_c_338_n N_A_811_379#_M1000_g 2.37377e-19 $X=5.885 $Y=0.68
+ $X2=0 $Y2=0
cc_404 N_A_83_21#_c_339_n N_A_811_379#_M1000_g 0.00807936f $X=4.96 $Y=0.68 $X2=0
+ $Y2=0
cc_405 N_A_83_21#_c_338_n N_A_811_379#_M1001_g 0.00987256f $X=5.885 $Y=0.68
+ $X2=0 $Y2=0
cc_406 N_A_83_21#_c_340_n N_A_811_379#_M1001_g 4.44855e-19 $X=6.05 $Y=0.68 $X2=0
+ $Y2=0
cc_407 N_A_83_21#_c_348_n N_A_1023_379#_M1005_g 2.96235e-19 $X=4.37 $Y=2.255
+ $X2=0 $Y2=0
cc_408 N_A_83_21#_c_338_n N_A_1023_379#_M1012_g 0.0130633f $X=5.885 $Y=0.68
+ $X2=0 $Y2=0
cc_409 N_A_83_21#_c_339_n N_A_1023_379#_M1012_g 0.00343987f $X=4.96 $Y=0.68
+ $X2=0 $Y2=0
cc_410 N_A_83_21#_c_340_n N_A_1023_379#_c_1100_n 0.00595239f $X=6.05 $Y=0.68
+ $X2=0 $Y2=0
cc_411 N_A_83_21#_c_336_n N_A_879_55#_M1000_s 0.00416748f $X=4.875 $Y=0.84
+ $X2=-0.19 $Y2=-0.245
cc_412 N_A_83_21#_c_336_n N_A_879_55#_c_1319_n 0.00626942f $X=4.875 $Y=0.84
+ $X2=0 $Y2=0
cc_413 N_A_83_21#_c_338_n N_A_879_55#_c_1319_n 0.0579576f $X=5.885 $Y=0.68 $X2=0
+ $Y2=0
cc_414 N_A_83_21#_c_339_n N_A_879_55#_c_1319_n 0.0123459f $X=4.96 $Y=0.68 $X2=0
+ $Y2=0
cc_415 N_A_83_21#_c_340_n N_A_879_55#_c_1319_n 0.021661f $X=6.05 $Y=0.68 $X2=0
+ $Y2=0
cc_416 N_A_83_21#_c_333_n N_A_879_55#_c_1324_n 0.0145294f $X=4.115 $Y=0.34 $X2=0
+ $Y2=0
cc_417 N_A_83_21#_c_335_n N_A_879_55#_c_1324_n 0.0121714f $X=4.2 $Y=0.755 $X2=0
+ $Y2=0
cc_418 N_A_83_21#_c_336_n N_A_879_55#_c_1324_n 0.0187088f $X=4.875 $Y=0.84 $X2=0
+ $Y2=0
cc_419 N_A_83_21#_M1029_g N_SUM_c_1794_n 0.0150852f $X=0.49 $Y=0.93 $X2=0 $Y2=0
cc_420 N_A_83_21#_c_325_n N_SUM_c_1794_n 0.00295945f $X=0.505 $Y=1.465 $X2=0
+ $Y2=0
cc_421 N_A_83_21#_c_326_n N_SUM_c_1794_n 0.00683961f $X=0.505 $Y=1.675 $X2=0
+ $Y2=0
cc_422 N_A_83_21#_c_343_n N_SUM_c_1794_n 0.0205359f $X=0.505 $Y=1.765 $X2=0
+ $Y2=0
cc_423 N_A_83_21#_c_346_n N_VPWR_M1015_d 0.00835435f $X=3.155 $Y=2.28 $X2=0
+ $Y2=0
cc_424 N_A_83_21#_c_376_p N_VPWR_M1015_d 0.00504006f $X=3.24 $Y=2.28 $X2=0 $Y2=0
cc_425 N_A_83_21#_c_343_n N_VPWR_c_1813_n 0.0059157f $X=0.505 $Y=1.765 $X2=0
+ $Y2=0
cc_426 N_A_83_21#_c_343_n N_VPWR_c_1812_n 0.00865885f $X=0.505 $Y=1.765 $X2=0
+ $Y2=0
cc_427 N_A_83_21#_c_343_n N_VPWR_c_1825_n 0.00445602f $X=0.505 $Y=1.765 $X2=0
+ $Y2=0
cc_428 N_A_83_21#_c_331_n N_COUT_M1006_s 8.27546e-19 $X=2.01 $Y=1.86 $X2=-0.19
+ $Y2=-0.245
cc_429 N_A_83_21#_c_366_p N_COUT_M1006_s 0.00407098f $X=2.175 $Y=0.985 $X2=-0.19
+ $Y2=-0.245
cc_430 N_A_83_21#_c_346_n N_COUT_M1015_s 0.0138834f $X=3.155 $Y=2.28 $X2=0 $Y2=0
cc_431 N_A_83_21#_M1029_g N_COUT_c_1944_n 0.00419714f $X=0.49 $Y=0.93 $X2=0
+ $Y2=0
cc_432 N_A_83_21#_c_325_n N_COUT_c_1944_n 0.0036427f $X=0.505 $Y=1.465 $X2=0
+ $Y2=0
cc_433 N_A_83_21#_c_343_n N_COUT_c_1944_n 0.00184686f $X=0.505 $Y=1.765 $X2=0
+ $Y2=0
cc_434 N_A_83_21#_c_327_n N_COUT_c_1945_n 0.00548628f $X=1.545 $Y=0.18 $X2=0
+ $Y2=0
cc_435 N_A_83_21#_M1029_g N_COUT_c_1969_n 0.00171966f $X=0.49 $Y=0.93 $X2=0
+ $Y2=0
cc_436 N_A_83_21#_c_327_n N_COUT_c_1969_n 7.06095e-19 $X=1.545 $Y=0.18 $X2=0
+ $Y2=0
cc_437 N_A_83_21#_c_343_n N_COUT_c_1956_n 0.00206873f $X=0.505 $Y=1.765 $X2=0
+ $Y2=0
cc_438 N_A_83_21#_c_343_n N_COUT_c_1958_n 0.00184546f $X=0.505 $Y=1.765 $X2=0
+ $Y2=0
cc_439 N_A_83_21#_c_345_n N_COUT_c_1950_n 2.82837e-19 $X=2.01 $Y=1.86 $X2=0
+ $Y2=0
cc_440 N_A_83_21#_c_329_n COUT 0.0249878f $X=1.62 $Y=1.235 $X2=0 $Y2=0
cc_441 N_A_83_21#_c_330_n COUT 0.00359732f $X=1.735 $Y=1.31 $X2=0 $Y2=0
cc_442 N_A_83_21#_c_366_p COUT 0.0146336f $X=2.175 $Y=0.985 $X2=0 $Y2=0
cc_443 N_A_83_21#_c_400_p N_A_644_104#_M1024_d 0.0134075f $X=4.205 $Y=2.37 $X2=0
+ $Y2=0
cc_444 N_A_83_21#_c_400_p N_A_644_104#_c_2022_n 0.00485635f $X=4.205 $Y=2.37
+ $X2=0 $Y2=0
cc_445 N_A_83_21#_c_376_p N_A_644_104#_c_2022_n 2.5231e-19 $X=3.24 $Y=2.28 $X2=0
+ $Y2=0
cc_446 N_A_83_21#_c_348_n N_A_644_104#_c_2022_n 0.00255557f $X=4.37 $Y=2.255
+ $X2=0 $Y2=0
cc_447 N_A_83_21#_c_346_n N_A_644_104#_c_2023_n 0.00178958f $X=3.155 $Y=2.28
+ $X2=0 $Y2=0
cc_448 N_A_83_21#_c_376_p N_A_644_104#_c_2023_n 4.98742e-19 $X=3.24 $Y=2.28
+ $X2=0 $Y2=0
cc_449 N_A_83_21#_c_346_n N_A_644_104#_c_2026_n 0.0112787f $X=3.155 $Y=2.28
+ $X2=0 $Y2=0
cc_450 N_A_83_21#_c_400_p N_A_644_104#_c_2026_n 0.0393078f $X=4.205 $Y=2.37
+ $X2=0 $Y2=0
cc_451 N_A_83_21#_c_376_p N_A_644_104#_c_2026_n 0.0115313f $X=3.24 $Y=2.28 $X2=0
+ $Y2=0
cc_452 N_A_83_21#_c_348_n N_A_644_104#_c_2026_n 0.00107222f $X=4.37 $Y=2.255
+ $X2=0 $Y2=0
cc_453 N_A_83_21#_c_365_p N_VGND_M1006_d 0.0186673f $X=2.595 $Y=0.985 $X2=0
+ $Y2=0
cc_454 N_A_83_21#_c_332_n N_VGND_M1006_d 0.0114553f $X=2.68 $Y=0.9 $X2=0 $Y2=0
cc_455 N_A_83_21#_M1029_g N_VGND_c_2317_n 0.0120264f $X=0.49 $Y=0.93 $X2=0 $Y2=0
cc_456 N_A_83_21#_c_327_n N_VGND_c_2317_n 0.0236598f $X=1.545 $Y=0.18 $X2=0
+ $Y2=0
cc_457 N_A_83_21#_c_329_n N_VGND_c_2317_n 0.00416665f $X=1.62 $Y=1.235 $X2=0
+ $Y2=0
cc_458 N_A_83_21#_c_327_n N_VGND_c_2318_n 0.00339969f $X=1.545 $Y=0.18 $X2=0
+ $Y2=0
cc_459 N_A_83_21#_c_365_p N_VGND_c_2318_n 0.0135869f $X=2.595 $Y=0.985 $X2=0
+ $Y2=0
cc_460 N_A_83_21#_c_332_n N_VGND_c_2318_n 0.022242f $X=2.68 $Y=0.9 $X2=0 $Y2=0
cc_461 N_A_83_21#_c_334_n N_VGND_c_2318_n 0.0143513f $X=2.765 $Y=0.34 $X2=0
+ $Y2=0
cc_462 N_A_83_21#_c_327_n N_VGND_c_2322_n 0.0192056f $X=1.545 $Y=0.18 $X2=0
+ $Y2=0
cc_463 N_A_83_21#_c_328_n N_VGND_c_2326_n 0.00762267f $X=0.565 $Y=0.18 $X2=0
+ $Y2=0
cc_464 N_A_83_21#_c_333_n N_VGND_c_2327_n 0.0990795f $X=4.115 $Y=0.34 $X2=0
+ $Y2=0
cc_465 N_A_83_21#_c_334_n N_VGND_c_2327_n 0.0121867f $X=2.765 $Y=0.34 $X2=0
+ $Y2=0
cc_466 N_A_83_21#_c_336_n N_VGND_c_2327_n 0.00246371f $X=4.875 $Y=0.84 $X2=0
+ $Y2=0
cc_467 N_A_83_21#_c_327_n N_VGND_c_2330_n 0.0257946f $X=1.545 $Y=0.18 $X2=0
+ $Y2=0
cc_468 N_A_83_21#_c_328_n N_VGND_c_2330_n 0.010022f $X=0.565 $Y=0.18 $X2=0 $Y2=0
cc_469 N_A_83_21#_c_333_n N_VGND_c_2330_n 0.0573556f $X=4.115 $Y=0.34 $X2=0
+ $Y2=0
cc_470 N_A_83_21#_c_334_n N_VGND_c_2330_n 0.00660921f $X=2.765 $Y=0.34 $X2=0
+ $Y2=0
cc_471 N_A_83_21#_c_336_n N_VGND_c_2330_n 0.00530161f $X=4.875 $Y=0.84 $X2=0
+ $Y2=0
cc_472 N_A_410_58#_c_563_p N_A_231_132#_M1005_d 0.0218721f $X=6.33 $Y=2.465
+ $X2=0 $Y2=0
cc_473 N_A_410_58#_c_517_n N_A_231_132#_c_650_n 0.0154343f $X=3.02 $Y=1.24 $X2=0
+ $Y2=0
cc_474 N_A_410_58#_c_518_n N_A_231_132#_c_650_n 0.0122461f $X=3.775 $Y=0.68
+ $X2=0 $Y2=0
cc_475 N_A_410_58#_c_550_n N_A_231_132#_c_650_n 0.00395622f $X=3.105 $Y=0.68
+ $X2=0 $Y2=0
cc_476 N_A_410_58#_c_519_n N_A_231_132#_c_650_n 0.00272086f $X=3.86 $Y=1.095
+ $X2=0 $Y2=0
cc_477 N_A_410_58#_c_516_n N_A_231_132#_c_651_n 0.0383705f $X=2.79 $Y=1.765
+ $X2=0 $Y2=0
cc_478 N_A_410_58#_c_518_n N_A_231_132#_c_651_n 0.00477714f $X=3.775 $Y=0.68
+ $X2=0 $Y2=0
cc_479 N_A_410_58#_c_522_n N_A_231_132#_c_651_n 0.00584835f $X=2.665 $Y=1.47
+ $X2=0 $Y2=0
cc_480 N_A_410_58#_c_516_n N_A_231_132#_c_661_n 0.00963087f $X=2.79 $Y=1.765
+ $X2=0 $Y2=0
cc_481 N_A_410_58#_c_516_n N_A_231_132#_c_695_n 3.45448e-19 $X=2.79 $Y=1.765
+ $X2=0 $Y2=0
cc_482 N_A_410_58#_c_521_n N_A_231_132#_c_653_n 0.0122763f $X=5.13 $Y=2.32 $X2=0
+ $Y2=0
cc_483 N_A_410_58#_c_523_n N_A_231_132#_c_653_n 0.0157863f $X=4.88 $Y=1.26 $X2=0
+ $Y2=0
cc_484 N_A_410_58#_c_521_n N_A_231_132#_c_654_n 0.0405706f $X=5.13 $Y=2.32 $X2=0
+ $Y2=0
cc_485 N_A_410_58#_c_554_n N_A_231_132#_c_654_n 0.0138308f $X=5.215 $Y=2.405
+ $X2=0 $Y2=0
cc_486 N_A_410_58#_c_554_n N_A_231_132#_c_665_n 0.00651968f $X=5.215 $Y=2.405
+ $X2=0 $Y2=0
cc_487 N_A_410_58#_c_563_p N_A_231_132#_c_665_n 0.0463983f $X=6.33 $Y=2.465
+ $X2=0 $Y2=0
cc_488 N_A_410_58#_c_579_p N_A_231_132#_c_667_n 0.0153963f $X=6.495 $Y=2.475
+ $X2=0 $Y2=0
cc_489 N_A_410_58#_c_563_p N_A_231_132#_c_667_n 0.00587208f $X=6.33 $Y=2.465
+ $X2=0 $Y2=0
cc_490 N_A_410_58#_M1017_d N_A_231_132#_c_743_n 0.0172302f $X=6.345 $Y=1.865
+ $X2=0 $Y2=0
cc_491 N_A_410_58#_c_579_p N_A_231_132#_c_743_n 0.0188328f $X=6.495 $Y=2.475
+ $X2=0 $Y2=0
cc_492 N_A_410_58#_c_563_p N_A_231_132#_c_743_n 0.00549887f $X=6.33 $Y=2.465
+ $X2=0 $Y2=0
cc_493 N_A_410_58#_c_563_p N_A_231_132#_c_746_n 0.00711829f $X=6.33 $Y=2.465
+ $X2=0 $Y2=0
cc_494 N_A_410_58#_M1017_d N_A_231_132#_c_668_n 0.00686012f $X=6.345 $Y=1.865
+ $X2=0 $Y2=0
cc_495 N_A_410_58#_c_579_p N_A_231_132#_c_668_n 0.0275002f $X=6.495 $Y=2.475
+ $X2=0 $Y2=0
cc_496 N_A_410_58#_c_516_n N_A_231_132#_c_713_n 0.00948606f $X=2.79 $Y=1.765
+ $X2=0 $Y2=0
cc_497 N_A_410_58#_c_516_n N_A_231_132#_c_670_n 7.9135e-19 $X=2.79 $Y=1.765
+ $X2=0 $Y2=0
cc_498 N_A_410_58#_c_518_n N_A_231_132#_c_716_n 0.0026969f $X=3.775 $Y=0.68
+ $X2=0 $Y2=0
cc_499 N_A_410_58#_c_520_n N_A_231_132#_c_716_n 0.0123985f $X=3.945 $Y=1.18
+ $X2=0 $Y2=0
cc_500 N_A_410_58#_c_523_n N_A_231_132#_c_716_n 0.0261106f $X=4.88 $Y=1.26 $X2=0
+ $Y2=0
cc_501 N_A_410_58#_c_520_n N_A_231_132#_c_657_n 0.00734216f $X=3.945 $Y=1.18
+ $X2=0 $Y2=0
cc_502 N_A_410_58#_c_523_n N_A_231_132#_c_657_n 0.0132553f $X=4.88 $Y=1.26 $X2=0
+ $Y2=0
cc_503 N_A_410_58#_c_524_n N_A_231_132#_c_657_n 8.96166e-19 $X=5.13 $Y=1.26
+ $X2=0 $Y2=0
cc_504 N_A_410_58#_c_521_n N_A_811_379#_c_896_n 8.68652e-19 $X=5.13 $Y=2.32
+ $X2=0 $Y2=0
cc_505 N_A_410_58#_c_521_n N_A_811_379#_M1000_g 0.00429432f $X=5.13 $Y=2.32
+ $X2=0 $Y2=0
cc_506 N_A_410_58#_c_523_n N_A_811_379#_M1000_g 0.00972803f $X=4.88 $Y=1.26
+ $X2=0 $Y2=0
cc_507 N_A_410_58#_c_524_n N_A_811_379#_M1000_g 0.00432634f $X=5.13 $Y=1.26
+ $X2=0 $Y2=0
cc_508 N_A_410_58#_c_563_p N_A_811_379#_c_908_n 4.12289e-19 $X=6.33 $Y=2.465
+ $X2=0 $Y2=0
cc_509 N_A_410_58#_c_579_p N_A_811_379#_c_909_n 0.00816607f $X=6.495 $Y=2.475
+ $X2=0 $Y2=0
cc_510 N_A_410_58#_c_563_p N_A_811_379#_c_909_n 0.0104422f $X=6.33 $Y=2.465
+ $X2=0 $Y2=0
cc_511 N_A_410_58#_c_523_n N_A_811_379#_c_901_n 0.00369479f $X=4.88 $Y=1.26
+ $X2=0 $Y2=0
cc_512 N_A_410_58#_c_521_n N_A_811_379#_c_903_n 0.0187771f $X=5.13 $Y=2.32 $X2=0
+ $Y2=0
cc_513 N_A_410_58#_c_524_n N_A_811_379#_c_903_n 0.00362675f $X=5.13 $Y=1.26
+ $X2=0 $Y2=0
cc_514 N_A_410_58#_c_563_p N_A_811_379#_c_903_n 0.00263211f $X=6.33 $Y=2.465
+ $X2=0 $Y2=0
cc_515 N_A_410_58#_c_563_p N_A_811_379#_c_904_n 0.00910537f $X=6.33 $Y=2.465
+ $X2=0 $Y2=0
cc_516 N_A_410_58#_c_579_p N_A_811_379#_c_914_n 0.00260268f $X=6.495 $Y=2.475
+ $X2=0 $Y2=0
cc_517 N_A_410_58#_c_563_p N_A_811_379#_c_914_n 0.0157919f $X=6.33 $Y=2.465
+ $X2=0 $Y2=0
cc_518 N_A_410_58#_c_521_n N_A_811_379#_c_915_n 0.00675927f $X=5.13 $Y=2.32
+ $X2=0 $Y2=0
cc_519 N_A_410_58#_c_563_p N_A_811_379#_c_915_n 0.00424674f $X=6.33 $Y=2.465
+ $X2=0 $Y2=0
cc_520 N_A_410_58#_c_521_n N_A_811_379#_c_916_n 0.0265109f $X=5.13 $Y=2.32 $X2=0
+ $Y2=0
cc_521 N_A_410_58#_c_563_p N_A_811_379#_c_916_n 0.0147997f $X=6.33 $Y=2.465
+ $X2=0 $Y2=0
cc_522 N_A_410_58#_c_521_n N_A_1023_379#_M1005_g 0.0135317f $X=5.13 $Y=2.32
+ $X2=0 $Y2=0
cc_523 N_A_410_58#_c_554_n N_A_1023_379#_M1005_g 0.00552017f $X=5.215 $Y=2.405
+ $X2=0 $Y2=0
cc_524 N_A_410_58#_c_563_p N_A_1023_379#_M1005_g 0.00756207f $X=6.33 $Y=2.465
+ $X2=0 $Y2=0
cc_525 N_A_410_58#_c_521_n N_A_1023_379#_M1012_g 0.00418577f $X=5.13 $Y=2.32
+ $X2=0 $Y2=0
cc_526 N_A_410_58#_c_524_n N_A_1023_379#_M1012_g 0.00447109f $X=5.13 $Y=1.26
+ $X2=0 $Y2=0
cc_527 N_A_410_58#_c_579_p N_A_1023_379#_M1003_g 0.00119931f $X=6.495 $Y=2.475
+ $X2=0 $Y2=0
cc_528 N_A_410_58#_c_521_n N_A_1023_379#_c_1104_n 0.00713612f $X=5.13 $Y=2.32
+ $X2=0 $Y2=0
cc_529 N_A_410_58#_c_524_n N_A_1023_379#_c_1104_n 2.35663e-19 $X=5.13 $Y=1.26
+ $X2=0 $Y2=0
cc_530 N_A_410_58#_c_563_p N_A_1023_379#_c_1104_n 0.0035313f $X=6.33 $Y=2.465
+ $X2=0 $Y2=0
cc_531 N_A_410_58#_c_523_n N_A_879_55#_M1000_s 0.00474163f $X=4.88 $Y=1.26
+ $X2=-0.19 $Y2=-0.245
cc_532 N_A_410_58#_c_516_n N_VPWR_c_1820_n 0.00322669f $X=2.79 $Y=1.765 $X2=0
+ $Y2=0
cc_533 N_A_410_58#_c_516_n N_VPWR_c_1812_n 0.0041252f $X=2.79 $Y=1.765 $X2=0
+ $Y2=0
cc_534 N_A_410_58#_c_516_n N_VPWR_c_1826_n 0.00262972f $X=2.79 $Y=1.765 $X2=0
+ $Y2=0
cc_535 N_A_410_58#_c_516_n N_COUT_c_1949_n 0.00666765f $X=2.79 $Y=1.765 $X2=0
+ $Y2=0
cc_536 N_A_410_58#_M1006_g COUT 0.00537382f $X=2.125 $Y=0.79 $X2=0 $Y2=0
cc_537 N_A_410_58#_c_518_n N_A_644_104#_M1028_d 0.00773538f $X=3.775 $Y=0.68
+ $X2=-0.19 $Y2=-0.245
cc_538 N_A_410_58#_c_516_n N_A_644_104#_c_2019_n 7.36458e-19 $X=2.79 $Y=1.765
+ $X2=0 $Y2=0
cc_539 N_A_410_58#_c_520_n N_A_644_104#_c_2019_n 0.00402215f $X=3.945 $Y=1.18
+ $X2=0 $Y2=0
cc_540 N_A_410_58#_c_522_n N_A_644_104#_c_2019_n 0.0186029f $X=2.665 $Y=1.47
+ $X2=0 $Y2=0
cc_541 N_A_410_58#_c_517_n N_A_644_104#_c_2021_n 0.0133329f $X=3.02 $Y=1.24
+ $X2=0 $Y2=0
cc_542 N_A_410_58#_c_518_n N_A_644_104#_c_2021_n 0.0256727f $X=3.775 $Y=0.68
+ $X2=0 $Y2=0
cc_543 N_A_410_58#_c_519_n N_A_644_104#_c_2021_n 0.012648f $X=3.86 $Y=1.095
+ $X2=0 $Y2=0
cc_544 N_A_410_58#_c_520_n N_A_644_104#_c_2021_n 0.00796151f $X=3.945 $Y=1.18
+ $X2=0 $Y2=0
cc_545 N_A_410_58#_c_520_n N_A_644_104#_c_2022_n 9.38935e-19 $X=3.945 $Y=1.18
+ $X2=0 $Y2=0
cc_546 N_A_410_58#_c_521_n N_A_644_104#_c_2022_n 0.0137335f $X=5.13 $Y=2.32
+ $X2=0 $Y2=0
cc_547 N_A_410_58#_c_523_n N_A_644_104#_c_2022_n 0.0111599f $X=4.88 $Y=1.26
+ $X2=0 $Y2=0
cc_548 N_A_410_58#_c_524_n N_A_644_104#_c_2022_n 0.0086366f $X=5.13 $Y=1.26
+ $X2=0 $Y2=0
cc_549 N_A_410_58#_c_563_p N_A_644_104#_c_2022_n 0.00433386f $X=6.33 $Y=2.465
+ $X2=0 $Y2=0
cc_550 N_A_410_58#_c_516_n N_A_644_104#_c_2023_n 0.00390716f $X=2.79 $Y=1.765
+ $X2=0 $Y2=0
cc_551 N_A_410_58#_c_522_n N_A_644_104#_c_2023_n 0.00744717f $X=2.665 $Y=1.47
+ $X2=0 $Y2=0
cc_552 N_A_410_58#_c_516_n N_A_644_104#_c_2026_n 0.0114948f $X=2.79 $Y=1.765
+ $X2=0 $Y2=0
cc_553 N_A_410_58#_c_522_n N_A_644_104#_c_2026_n 0.0110293f $X=2.665 $Y=1.47
+ $X2=0 $Y2=0
cc_554 N_A_410_58#_c_517_n N_VGND_M1006_d 0.00666905f $X=3.02 $Y=1.24 $X2=0
+ $Y2=0
cc_555 N_A_410_58#_c_550_n N_VGND_M1006_d 0.00271055f $X=3.105 $Y=0.68 $X2=0
+ $Y2=0
cc_556 N_A_410_58#_M1006_g N_VGND_c_2318_n 0.00470773f $X=2.125 $Y=0.79 $X2=0
+ $Y2=0
cc_557 N_A_410_58#_M1006_g N_VGND_c_2322_n 0.00516294f $X=2.125 $Y=0.79 $X2=0
+ $Y2=0
cc_558 N_A_410_58#_M1006_g N_VGND_c_2330_n 0.00529924f $X=2.125 $Y=0.79 $X2=0
+ $Y2=0
cc_559 N_A_231_132#_c_651_n N_A_811_379#_c_905_n 0.0172587f $X=3.435 $Y=1.81
+ $X2=0 $Y2=0
cc_560 N_A_231_132#_c_663_n N_A_811_379#_c_905_n 0.0136824f $X=4.705 $Y=2.99
+ $X2=0 $Y2=0
cc_561 N_A_231_132#_c_654_n N_A_811_379#_c_905_n 0.00215818f $X=4.79 $Y=2.73
+ $X2=0 $Y2=0
cc_562 N_A_231_132#_c_670_n N_A_811_379#_c_905_n 0.00395126f $X=3.545 $Y=2.71
+ $X2=0 $Y2=0
cc_563 N_A_231_132#_c_672_n N_A_811_379#_c_905_n 0.00416934f $X=4.79 $Y=2.902
+ $X2=0 $Y2=0
cc_564 N_A_231_132#_c_653_n N_A_811_379#_c_894_n 0.00368945f $X=4.705 $Y=1.68
+ $X2=0 $Y2=0
cc_565 N_A_231_132#_c_654_n N_A_811_379#_c_894_n 0.00877383f $X=4.79 $Y=2.73
+ $X2=0 $Y2=0
cc_566 N_A_231_132#_c_651_n N_A_811_379#_c_895_n 0.00240122f $X=3.435 $Y=1.81
+ $X2=0 $Y2=0
cc_567 N_A_231_132#_c_716_n N_A_811_379#_c_895_n 7.44199e-19 $X=4.175 $Y=1.52
+ $X2=0 $Y2=0
cc_568 N_A_231_132#_c_657_n N_A_811_379#_c_895_n 0.0182941f $X=4.175 $Y=1.52
+ $X2=0 $Y2=0
cc_569 N_A_231_132#_c_658_n N_A_811_379#_c_895_n 0.00368945f $X=4.34 $Y=1.6
+ $X2=0 $Y2=0
cc_570 N_A_231_132#_c_653_n N_A_811_379#_c_896_n 0.00790075f $X=4.705 $Y=1.68
+ $X2=0 $Y2=0
cc_571 N_A_231_132#_c_654_n N_A_811_379#_c_896_n 0.00668273f $X=4.79 $Y=2.73
+ $X2=0 $Y2=0
cc_572 N_A_231_132#_c_657_n N_A_811_379#_M1000_g 0.00938688f $X=4.175 $Y=1.52
+ $X2=0 $Y2=0
cc_573 N_A_231_132#_c_658_n N_A_811_379#_M1000_g 6.40607e-19 $X=4.34 $Y=1.6
+ $X2=0 $Y2=0
cc_574 N_A_231_132#_c_724_n N_A_811_379#_M1000_g 6.86076e-19 $X=5.55 $Y=1.03
+ $X2=0 $Y2=0
cc_575 N_A_231_132#_c_704_n N_A_811_379#_M1001_g 0.00869923f $X=6.055 $Y=1.12
+ $X2=0 $Y2=0
cc_576 N_A_231_132#_c_655_n N_A_811_379#_M1001_g 0.00342239f $X=6.14 $Y=1.95
+ $X2=0 $Y2=0
cc_577 N_A_231_132#_c_724_n N_A_811_379#_M1001_g 0.00344766f $X=5.55 $Y=1.03
+ $X2=0 $Y2=0
cc_578 N_A_231_132#_c_704_n N_A_811_379#_c_908_n 0.00224077f $X=6.055 $Y=1.12
+ $X2=0 $Y2=0
cc_579 N_A_231_132#_c_655_n N_A_811_379#_c_908_n 0.0119134f $X=6.14 $Y=1.95
+ $X2=0 $Y2=0
cc_580 N_A_231_132#_c_655_n N_A_811_379#_c_909_n 0.00914765f $X=6.14 $Y=1.95
+ $X2=0 $Y2=0
cc_581 N_A_231_132#_c_667_n N_A_811_379#_c_909_n 0.00161872f $X=6.83 $Y=2.99
+ $X2=0 $Y2=0
cc_582 N_A_231_132#_c_743_n N_A_811_379#_c_909_n 0.00767498f $X=6.83 $Y=2.035
+ $X2=0 $Y2=0
cc_583 N_A_231_132#_c_746_n N_A_811_379#_c_909_n 0.00385306f $X=6.225 $Y=2.035
+ $X2=0 $Y2=0
cc_584 N_A_231_132#_c_668_n N_A_811_379#_c_909_n 0.0057579f $X=6.915 $Y=2.905
+ $X2=0 $Y2=0
cc_585 N_A_231_132#_c_673_n N_A_811_379#_c_909_n 0.00476737f $X=6.125 $Y=2.902
+ $X2=0 $Y2=0
cc_586 N_A_231_132#_c_653_n N_A_811_379#_c_901_n 0.0103911f $X=4.705 $Y=1.68
+ $X2=0 $Y2=0
cc_587 N_A_231_132#_c_657_n N_A_811_379#_c_901_n 0.00738436f $X=4.175 $Y=1.52
+ $X2=0 $Y2=0
cc_588 N_A_231_132#_c_658_n N_A_811_379#_c_901_n 3.11201e-19 $X=4.34 $Y=1.6
+ $X2=0 $Y2=0
cc_589 N_A_231_132#_c_704_n N_A_811_379#_c_903_n 0.0101758f $X=6.055 $Y=1.12
+ $X2=0 $Y2=0
cc_590 N_A_231_132#_c_655_n N_A_811_379#_c_903_n 0.0241515f $X=6.14 $Y=1.95
+ $X2=0 $Y2=0
cc_591 N_A_231_132#_c_724_n N_A_811_379#_c_903_n 0.0192285f $X=5.55 $Y=1.03
+ $X2=0 $Y2=0
cc_592 N_A_231_132#_c_704_n N_A_811_379#_c_904_n 0.00326335f $X=6.055 $Y=1.12
+ $X2=0 $Y2=0
cc_593 N_A_231_132#_c_655_n N_A_811_379#_c_904_n 0.00573579f $X=6.14 $Y=1.95
+ $X2=0 $Y2=0
cc_594 N_A_231_132#_c_724_n N_A_811_379#_c_904_n 0.00152514f $X=5.55 $Y=1.03
+ $X2=0 $Y2=0
cc_595 N_A_231_132#_M1005_d N_A_811_379#_c_914_n 0.00214522f $X=5.28 $Y=2.12
+ $X2=0 $Y2=0
cc_596 N_A_231_132#_c_743_n N_A_811_379#_c_914_n 0.0417874f $X=6.83 $Y=2.035
+ $X2=0 $Y2=0
cc_597 N_A_231_132#_c_746_n N_A_811_379#_c_914_n 0.0101765f $X=6.225 $Y=2.035
+ $X2=0 $Y2=0
cc_598 N_A_231_132#_M1005_d N_A_811_379#_c_915_n 0.00321801f $X=5.28 $Y=2.12
+ $X2=0 $Y2=0
cc_599 N_A_231_132#_c_655_n N_A_811_379#_c_915_n 7.51534e-19 $X=6.14 $Y=1.95
+ $X2=0 $Y2=0
cc_600 N_A_231_132#_c_746_n N_A_811_379#_c_915_n 7.983e-19 $X=6.225 $Y=2.035
+ $X2=0 $Y2=0
cc_601 N_A_231_132#_M1005_d N_A_811_379#_c_916_n 0.00182073f $X=5.28 $Y=2.12
+ $X2=0 $Y2=0
cc_602 N_A_231_132#_c_655_n N_A_811_379#_c_916_n 0.00849516f $X=6.14 $Y=1.95
+ $X2=0 $Y2=0
cc_603 N_A_231_132#_c_746_n N_A_811_379#_c_916_n 0.00463277f $X=6.225 $Y=2.035
+ $X2=0 $Y2=0
cc_604 N_A_231_132#_c_654_n N_A_1023_379#_M1005_g 0.0100373f $X=4.79 $Y=2.73
+ $X2=0 $Y2=0
cc_605 N_A_231_132#_c_665_n N_A_1023_379#_M1005_g 0.0154212f $X=5.953 $Y=2.902
+ $X2=0 $Y2=0
cc_606 N_A_231_132#_c_655_n N_A_1023_379#_M1012_g 7.26554e-19 $X=6.14 $Y=1.95
+ $X2=0 $Y2=0
cc_607 N_A_231_132#_c_724_n N_A_1023_379#_M1012_g 0.00494072f $X=5.55 $Y=1.03
+ $X2=0 $Y2=0
cc_608 N_A_231_132#_c_665_n N_A_1023_379#_c_1117_n 0.0340411f $X=5.953 $Y=2.902
+ $X2=0 $Y2=0
cc_609 N_A_231_132#_c_667_n N_A_1023_379#_c_1117_n 0.00312806f $X=6.83 $Y=2.99
+ $X2=0 $Y2=0
cc_610 N_A_231_132#_c_665_n N_A_1023_379#_c_1118_n 0.00470511f $X=5.953 $Y=2.902
+ $X2=0 $Y2=0
cc_611 N_A_231_132#_c_704_n N_A_1023_379#_c_1100_n 0.00490817f $X=6.055 $Y=1.12
+ $X2=0 $Y2=0
cc_612 N_A_231_132#_c_655_n N_A_1023_379#_c_1100_n 8.42764e-19 $X=6.14 $Y=1.95
+ $X2=0 $Y2=0
cc_613 N_A_231_132#_c_724_n N_A_1023_379#_c_1100_n 4.74488e-19 $X=5.55 $Y=1.03
+ $X2=0 $Y2=0
cc_614 N_A_231_132#_c_743_n N_A_1023_379#_c_1101_n 0.00609153f $X=6.83 $Y=2.035
+ $X2=0 $Y2=0
cc_615 N_A_231_132#_c_655_n N_A_1023_379#_c_1102_n 0.00410097f $X=6.14 $Y=1.95
+ $X2=0 $Y2=0
cc_616 N_A_231_132#_c_743_n N_A_1023_379#_c_1102_n 5.01988e-19 $X=6.83 $Y=2.035
+ $X2=0 $Y2=0
cc_617 N_A_231_132#_c_668_n N_A_1023_379#_c_1120_n 0.00282874f $X=6.915 $Y=2.905
+ $X2=0 $Y2=0
cc_618 N_A_231_132#_c_667_n N_A_1023_379#_c_1121_n 0.00799512f $X=6.83 $Y=2.99
+ $X2=0 $Y2=0
cc_619 N_A_231_132#_c_668_n N_A_1023_379#_c_1121_n 9.96081e-19 $X=6.915 $Y=2.905
+ $X2=0 $Y2=0
cc_620 N_A_231_132#_c_743_n N_A_1023_379#_M1003_g 0.00555204f $X=6.83 $Y=2.035
+ $X2=0 $Y2=0
cc_621 N_A_231_132#_c_668_n N_A_1023_379#_M1003_g 0.015959f $X=6.915 $Y=2.905
+ $X2=0 $Y2=0
cc_622 N_A_231_132#_c_654_n N_A_1023_379#_c_1104_n 4.33207e-19 $X=4.79 $Y=2.73
+ $X2=0 $Y2=0
cc_623 N_A_231_132#_c_746_n N_A_1023_379#_c_1104_n 3.30996e-19 $X=6.225 $Y=2.035
+ $X2=0 $Y2=0
cc_624 N_A_231_132#_c_743_n N_A_1023_379#_c_1105_n 5.96439e-19 $X=6.83 $Y=2.035
+ $X2=0 $Y2=0
cc_625 N_A_231_132#_c_743_n N_A_1023_379#_c_1166_n 0.00225902f $X=6.83 $Y=2.035
+ $X2=0 $Y2=0
cc_626 N_A_231_132#_c_743_n N_A_1023_379#_c_1112_n 0.00107496f $X=6.83 $Y=2.035
+ $X2=0 $Y2=0
cc_627 N_A_231_132#_c_743_n N_A_1023_379#_c_1113_n 0.00892773f $X=6.83 $Y=2.035
+ $X2=0 $Y2=0
cc_628 N_A_231_132#_c_704_n N_A_879_55#_c_1319_n 2.89871e-19 $X=6.055 $Y=1.12
+ $X2=0 $Y2=0
cc_629 N_A_231_132#_c_667_n N_A_879_55#_c_1336_n 0.00167808f $X=6.83 $Y=2.99
+ $X2=0 $Y2=0
cc_630 N_A_231_132#_c_668_n N_A_879_55#_c_1336_n 0.0582492f $X=6.915 $Y=2.905
+ $X2=0 $Y2=0
cc_631 N_A_231_132#_c_743_n N_A_879_55#_c_1353_n 0.0119685f $X=6.83 $Y=2.035
+ $X2=0 $Y2=0
cc_632 N_A_231_132#_c_667_n N_B_c_1518_n 3.64859e-19 $X=6.83 $Y=2.99 $X2=-0.19
+ $Y2=-0.245
cc_633 N_A_231_132#_c_695_n N_VPWR_M1015_d 0.00864632f $X=3.46 $Y=2.71 $X2=0
+ $Y2=0
cc_634 N_A_231_132#_c_713_n N_VPWR_M1015_d 0.00302891f $X=2.9 $Y=2.62 $X2=0
+ $Y2=0
cc_635 N_A_231_132#_c_667_n N_VPWR_c_1814_n 0.00434568f $X=6.83 $Y=2.99 $X2=0
+ $Y2=0
cc_636 N_A_231_132#_c_661_n N_VPWR_c_1820_n 0.00247647f $X=2.815 $Y=2.62 $X2=0
+ $Y2=0
cc_637 N_A_231_132#_c_713_n N_VPWR_c_1820_n 0.0020828f $X=2.9 $Y=2.62 $X2=0
+ $Y2=0
cc_638 N_A_231_132#_c_651_n N_VPWR_c_1821_n 0.00291715f $X=3.435 $Y=1.81 $X2=0
+ $Y2=0
cc_639 N_A_231_132#_c_695_n N_VPWR_c_1821_n 0.00310787f $X=3.46 $Y=2.71 $X2=0
+ $Y2=0
cc_640 N_A_231_132#_c_663_n N_VPWR_c_1821_n 0.0687839f $X=4.705 $Y=2.99 $X2=0
+ $Y2=0
cc_641 N_A_231_132#_c_665_n N_VPWR_c_1821_n 0.12933f $X=5.953 $Y=2.902 $X2=0
+ $Y2=0
cc_642 N_A_231_132#_c_667_n N_VPWR_c_1821_n 0.0115566f $X=6.83 $Y=2.99 $X2=0
+ $Y2=0
cc_643 N_A_231_132#_c_670_n N_VPWR_c_1821_n 0.0116773f $X=3.545 $Y=2.71 $X2=0
+ $Y2=0
cc_644 N_A_231_132#_c_672_n N_VPWR_c_1821_n 0.0121505f $X=4.79 $Y=2.902 $X2=0
+ $Y2=0
cc_645 N_A_231_132#_c_651_n N_VPWR_c_1812_n 0.00351561f $X=3.435 $Y=1.81 $X2=0
+ $Y2=0
cc_646 N_A_231_132#_c_661_n N_VPWR_c_1812_n 0.00654036f $X=2.815 $Y=2.62 $X2=0
+ $Y2=0
cc_647 N_A_231_132#_c_695_n N_VPWR_c_1812_n 0.00685329f $X=3.46 $Y=2.71 $X2=0
+ $Y2=0
cc_648 N_A_231_132#_c_663_n N_VPWR_c_1812_n 0.0397311f $X=4.705 $Y=2.99 $X2=0
+ $Y2=0
cc_649 N_A_231_132#_c_665_n N_VPWR_c_1812_n 0.0672694f $X=5.953 $Y=2.902 $X2=0
+ $Y2=0
cc_650 N_A_231_132#_c_667_n N_VPWR_c_1812_n 0.00579705f $X=6.83 $Y=2.99 $X2=0
+ $Y2=0
cc_651 N_A_231_132#_c_713_n N_VPWR_c_1812_n 0.00380867f $X=2.9 $Y=2.62 $X2=0
+ $Y2=0
cc_652 N_A_231_132#_c_670_n N_VPWR_c_1812_n 0.00646299f $X=3.545 $Y=2.71 $X2=0
+ $Y2=0
cc_653 N_A_231_132#_c_672_n N_VPWR_c_1812_n 0.00660393f $X=4.79 $Y=2.902 $X2=0
+ $Y2=0
cc_654 N_A_231_132#_c_651_n N_VPWR_c_1826_n 4.89596e-19 $X=3.435 $Y=1.81 $X2=0
+ $Y2=0
cc_655 N_A_231_132#_c_695_n N_VPWR_c_1826_n 0.0224053f $X=3.46 $Y=2.71 $X2=0
+ $Y2=0
cc_656 N_A_231_132#_c_713_n N_VPWR_c_1826_n 0.00368286f $X=2.9 $Y=2.62 $X2=0
+ $Y2=0
cc_657 N_A_231_132#_c_670_n N_VPWR_c_1826_n 0.00858282f $X=3.545 $Y=2.71 $X2=0
+ $Y2=0
cc_658 N_A_231_132#_c_661_n N_COUT_M1015_s 0.00868396f $X=2.815 $Y=2.62 $X2=0
+ $Y2=0
cc_659 N_A_231_132#_c_652_n N_COUT_c_1944_n 0.00847167f $X=1.505 $Y=1.155 $X2=0
+ $Y2=0
cc_660 N_A_231_132#_c_656_n N_COUT_c_1944_n 0.00936463f $X=1.5 $Y=1.95 $X2=0
+ $Y2=0
cc_661 N_A_231_132#_M1010_d N_COUT_c_1945_n 0.00699152f $X=1.155 $Y=0.66 $X2=0
+ $Y2=0
cc_662 N_A_231_132#_c_652_n N_COUT_c_1945_n 0.0229602f $X=1.505 $Y=1.155 $X2=0
+ $Y2=0
cc_663 N_A_231_132#_c_662_n N_COUT_c_1956_n 0.0156596f $X=1.675 $Y=2.62 $X2=0
+ $Y2=0
cc_664 N_A_231_132#_c_677_n N_COUT_c_1956_n 0.0307726f $X=1.41 $Y=2.115 $X2=0
+ $Y2=0
cc_665 N_A_231_132#_c_677_n N_COUT_c_1958_n 0.0135591f $X=1.41 $Y=2.115 $X2=0
+ $Y2=0
cc_666 N_A_231_132#_c_661_n N_COUT_c_1949_n 0.0230318f $X=2.815 $Y=2.62 $X2=0
+ $Y2=0
cc_667 N_A_231_132#_c_661_n N_COUT_c_1950_n 0.0397244f $X=2.815 $Y=2.62 $X2=0
+ $Y2=0
cc_668 N_A_231_132#_c_662_n N_COUT_c_1950_n 0.0272931f $X=1.675 $Y=2.62 $X2=0
+ $Y2=0
cc_669 N_A_231_132#_c_652_n COUT 0.0144163f $X=1.505 $Y=1.155 $X2=0 $Y2=0
cc_670 N_A_231_132#_c_663_n N_A_644_104#_M1024_d 0.00380577f $X=4.705 $Y=2.99
+ $X2=0 $Y2=0
cc_671 N_A_231_132#_c_670_n N_A_644_104#_M1024_d 0.00460776f $X=3.545 $Y=2.71
+ $X2=0 $Y2=0
cc_672 N_A_231_132#_c_651_n N_A_644_104#_c_2019_n 0.0232561f $X=3.435 $Y=1.81
+ $X2=0 $Y2=0
cc_673 N_A_231_132#_c_716_n N_A_644_104#_c_2019_n 0.00854576f $X=4.175 $Y=1.52
+ $X2=0 $Y2=0
cc_674 N_A_231_132#_c_704_n N_A_644_104#_c_2020_n 0.00795365f $X=6.055 $Y=1.12
+ $X2=0 $Y2=0
cc_675 N_A_231_132#_c_655_n N_A_644_104#_c_2020_n 0.0399443f $X=6.14 $Y=1.95
+ $X2=0 $Y2=0
cc_676 N_A_231_132#_c_650_n N_A_644_104#_c_2021_n 0.00605086f $X=3.145 $Y=1.24
+ $X2=0 $Y2=0
cc_677 N_A_231_132#_c_651_n N_A_644_104#_c_2021_n 0.00562457f $X=3.435 $Y=1.81
+ $X2=0 $Y2=0
cc_678 N_A_231_132#_c_651_n N_A_644_104#_c_2022_n 0.00232855f $X=3.435 $Y=1.81
+ $X2=0 $Y2=0
cc_679 N_A_231_132#_c_653_n N_A_644_104#_c_2022_n 0.0303408f $X=4.705 $Y=1.68
+ $X2=0 $Y2=0
cc_680 N_A_231_132#_c_704_n N_A_644_104#_c_2022_n 0.00674046f $X=6.055 $Y=1.12
+ $X2=0 $Y2=0
cc_681 N_A_231_132#_c_655_n N_A_644_104#_c_2022_n 0.0163998f $X=6.14 $Y=1.95
+ $X2=0 $Y2=0
cc_682 N_A_231_132#_c_743_n N_A_644_104#_c_2022_n 0.00231019f $X=6.83 $Y=2.035
+ $X2=0 $Y2=0
cc_683 N_A_231_132#_c_716_n N_A_644_104#_c_2022_n 0.0190201f $X=4.175 $Y=1.52
+ $X2=0 $Y2=0
cc_684 N_A_231_132#_c_657_n N_A_644_104#_c_2022_n 0.00800818f $X=4.175 $Y=1.52
+ $X2=0 $Y2=0
cc_685 N_A_231_132#_c_658_n N_A_644_104#_c_2022_n 0.00910703f $X=4.34 $Y=1.6
+ $X2=0 $Y2=0
cc_686 N_A_231_132#_c_724_n N_A_644_104#_c_2022_n 0.00209161f $X=5.55 $Y=1.03
+ $X2=0 $Y2=0
cc_687 N_A_231_132#_c_651_n N_A_644_104#_c_2023_n 0.00446096f $X=3.435 $Y=1.81
+ $X2=0 $Y2=0
cc_688 N_A_231_132#_c_655_n N_A_644_104#_c_2024_n 0.00255563f $X=6.14 $Y=1.95
+ $X2=0 $Y2=0
cc_689 N_A_231_132#_c_743_n N_A_644_104#_c_2024_n 0.00308485f $X=6.83 $Y=2.035
+ $X2=0 $Y2=0
cc_690 N_A_231_132#_c_743_n N_A_644_104#_c_2025_n 0.0129936f $X=6.83 $Y=2.035
+ $X2=0 $Y2=0
cc_691 N_A_231_132#_c_651_n N_A_644_104#_c_2026_n 0.0367049f $X=3.435 $Y=1.81
+ $X2=0 $Y2=0
cc_692 N_A_231_132#_c_716_n N_A_644_104#_c_2026_n 0.0266093f $X=4.175 $Y=1.52
+ $X2=0 $Y2=0
cc_693 N_A_231_132#_c_657_n N_A_644_104#_c_2026_n 0.00998674f $X=4.175 $Y=1.52
+ $X2=0 $Y2=0
cc_694 N_A_231_132#_c_650_n N_VGND_c_2318_n 2.64462e-19 $X=3.145 $Y=1.24 $X2=0
+ $Y2=0
cc_695 N_A_231_132#_c_650_n N_VGND_c_2327_n 6.75092e-19 $X=3.145 $Y=1.24 $X2=0
+ $Y2=0
cc_696 N_A_811_379#_c_915_n N_A_1023_379#_M1005_g 0.00287112f $X=5.665 $Y=2.035
+ $X2=0 $Y2=0
cc_697 N_A_811_379#_c_916_n N_A_1023_379#_M1005_g 0.00208045f $X=5.52 $Y=2.035
+ $X2=0 $Y2=0
cc_698 N_A_811_379#_c_896_n N_A_1023_379#_M1012_g 0.00310657f $X=4.655 $Y=1.895
+ $X2=0 $Y2=0
cc_699 N_A_811_379#_M1000_g N_A_1023_379#_M1012_g 0.0317643f $X=4.83 $Y=1.155
+ $X2=0 $Y2=0
cc_700 N_A_811_379#_c_898_n N_A_1023_379#_M1012_g 0.00737859f $X=5.69 $Y=0.18
+ $X2=0 $Y2=0
cc_701 N_A_811_379#_M1001_g N_A_1023_379#_M1012_g 0.0221992f $X=5.765 $Y=0.945
+ $X2=0 $Y2=0
cc_702 N_A_811_379#_c_903_n N_A_1023_379#_M1012_g 0.00571137f $X=5.785 $Y=1.54
+ $X2=0 $Y2=0
cc_703 N_A_811_379#_c_904_n N_A_1023_379#_M1012_g 0.0268717f $X=5.785 $Y=1.54
+ $X2=0 $Y2=0
cc_704 N_A_811_379#_c_916_n N_A_1023_379#_M1012_g 0.0044339f $X=5.52 $Y=2.035
+ $X2=0 $Y2=0
cc_705 N_A_811_379#_c_909_n N_A_1023_379#_c_1117_n 0.00737859f $X=6.27 $Y=1.79
+ $X2=0 $Y2=0
cc_706 N_A_811_379#_M1001_g N_A_1023_379#_c_1100_n 0.0261262f $X=5.765 $Y=0.945
+ $X2=0 $Y2=0
cc_707 N_A_811_379#_c_908_n N_A_1023_379#_c_1102_n 0.0105351f $X=6.195 $Y=1.715
+ $X2=0 $Y2=0
cc_708 N_A_811_379#_c_904_n N_A_1023_379#_c_1102_n 0.00131035f $X=5.785 $Y=1.54
+ $X2=0 $Y2=0
cc_709 N_A_811_379#_c_908_n N_A_1023_379#_c_1103_n 0.00283994f $X=6.195 $Y=1.715
+ $X2=0 $Y2=0
cc_710 N_A_811_379#_c_909_n N_A_1023_379#_c_1120_n 7.8304e-19 $X=6.27 $Y=1.79
+ $X2=0 $Y2=0
cc_711 N_A_811_379#_c_914_n N_A_1023_379#_c_1122_n 2.62074e-19 $X=8.78 $Y=2.035
+ $X2=0 $Y2=0
cc_712 N_A_811_379#_c_909_n N_A_1023_379#_M1003_g 0.0125183f $X=6.27 $Y=1.79
+ $X2=0 $Y2=0
cc_713 N_A_811_379#_c_914_n N_A_1023_379#_M1003_g 0.00593455f $X=8.78 $Y=2.035
+ $X2=0 $Y2=0
cc_714 N_A_811_379#_c_894_n N_A_1023_379#_c_1104_n 0.00444073f $X=4.58 $Y=1.97
+ $X2=0 $Y2=0
cc_715 N_A_811_379#_c_915_n N_A_1023_379#_c_1104_n 0.00168143f $X=5.665 $Y=2.035
+ $X2=0 $Y2=0
cc_716 N_A_811_379#_c_916_n N_A_1023_379#_c_1104_n 0.00429793f $X=5.52 $Y=2.035
+ $X2=0 $Y2=0
cc_717 N_A_811_379#_c_1010_p N_A_1023_379#_c_1109_n 0.0250371f $X=10.65 $Y=0.82
+ $X2=0 $Y2=0
cc_718 N_A_811_379#_c_910_n N_A_1023_379#_c_1125_n 0.0134336f $X=10.645 $Y=2.65
+ $X2=0 $Y2=0
cc_719 N_A_811_379#_c_914_n N_A_1023_379#_c_1166_n 5.2141e-19 $X=8.78 $Y=2.035
+ $X2=0 $Y2=0
cc_720 N_A_811_379#_c_902_n N_A_1023_379#_c_1111_n 0.0163574f $X=10.73 $Y=2.565
+ $X2=0 $Y2=0
cc_721 N_A_811_379#_c_1010_p N_A_1023_379#_c_1111_n 0.00561237f $X=10.65 $Y=0.82
+ $X2=0 $Y2=0
cc_722 N_A_811_379#_c_914_n N_A_1023_379#_c_1111_n 0.122801f $X=8.78 $Y=2.035
+ $X2=0 $Y2=0
cc_723 N_A_811_379#_c_1016_p N_A_1023_379#_c_1111_n 0.0241866f $X=8.925 $Y=2.035
+ $X2=0 $Y2=0
cc_724 N_A_811_379#_c_1017_p N_A_1023_379#_c_1111_n 0.00653929f $X=8.925
+ $Y=2.035 $X2=0 $Y2=0
cc_725 N_A_811_379#_c_914_n N_A_1023_379#_c_1112_n 0.0235648f $X=8.78 $Y=2.035
+ $X2=0 $Y2=0
cc_726 N_A_811_379#_c_914_n N_A_1023_379#_c_1113_n 0.00153114f $X=8.78 $Y=2.035
+ $X2=0 $Y2=0
cc_727 N_A_811_379#_c_902_n N_A_1023_379#_c_1129_n 0.00261636f $X=10.73 $Y=2.565
+ $X2=0 $Y2=0
cc_728 N_A_811_379#_c_902_n N_A_1023_379#_c_1130_n 0.0705982f $X=10.73 $Y=2.565
+ $X2=0 $Y2=0
cc_729 N_A_811_379#_M1002_d N_A_1023_379#_c_1115_n 0.0158189f $X=10.18 $Y=0.47
+ $X2=0 $Y2=0
cc_730 N_A_811_379#_c_1010_p N_A_1023_379#_c_1115_n 0.0705982f $X=10.65 $Y=0.82
+ $X2=0 $Y2=0
cc_731 N_A_811_379#_c_914_n N_A_879_55#_M1003_d 0.00335095f $X=8.78 $Y=2.035
+ $X2=0 $Y2=0
cc_732 N_A_811_379#_c_911_n N_A_879_55#_c_1314_n 0.00100316f $X=9.11 $Y=2.65
+ $X2=0 $Y2=0
cc_733 N_A_811_379#_c_914_n N_A_879_55#_c_1314_n 0.00754601f $X=8.78 $Y=2.035
+ $X2=0 $Y2=0
cc_734 N_A_811_379#_c_1016_p N_A_879_55#_c_1314_n 0.00156324f $X=8.925 $Y=2.035
+ $X2=0 $Y2=0
cc_735 N_A_811_379#_c_1017_p N_A_879_55#_c_1314_n 0.00494152f $X=8.925 $Y=2.035
+ $X2=0 $Y2=0
cc_736 N_A_811_379#_c_902_n N_A_879_55#_c_1316_n 8.12245e-19 $X=10.73 $Y=2.565
+ $X2=0 $Y2=0
cc_737 N_A_811_379#_c_1010_p N_A_879_55#_c_1316_n 0.00313017f $X=10.65 $Y=0.82
+ $X2=0 $Y2=0
cc_738 N_A_811_379#_c_902_n N_A_879_55#_c_1317_n 0.00878214f $X=10.73 $Y=2.565
+ $X2=0 $Y2=0
cc_739 N_A_811_379#_c_1010_p N_A_879_55#_c_1317_n 0.00508142f $X=10.65 $Y=0.82
+ $X2=0 $Y2=0
cc_740 N_A_811_379#_c_910_n N_A_879_55#_c_1334_n 0.00636176f $X=10.645 $Y=2.65
+ $X2=0 $Y2=0
cc_741 N_A_811_379#_c_902_n N_A_879_55#_c_1334_n 0.0221727f $X=10.73 $Y=2.565
+ $X2=0 $Y2=0
cc_742 N_A_811_379#_c_902_n N_A_879_55#_c_1318_n 0.00977631f $X=10.73 $Y=2.565
+ $X2=0 $Y2=0
cc_743 N_A_811_379#_M1000_g N_A_879_55#_c_1319_n 0.0129893f $X=4.83 $Y=1.155
+ $X2=0 $Y2=0
cc_744 N_A_811_379#_c_898_n N_A_879_55#_c_1319_n 0.0117727f $X=5.69 $Y=0.18
+ $X2=0 $Y2=0
cc_745 N_A_811_379#_M1001_g N_A_879_55#_c_1319_n 0.0136053f $X=5.765 $Y=0.945
+ $X2=0 $Y2=0
cc_746 N_A_811_379#_M1002_d N_A_879_55#_c_1369_n 0.00276274f $X=10.18 $Y=0.47
+ $X2=0 $Y2=0
cc_747 N_A_811_379#_c_1010_p N_A_879_55#_c_1369_n 0.0144778f $X=10.65 $Y=0.82
+ $X2=0 $Y2=0
cc_748 N_A_811_379#_M1000_g N_A_879_55#_c_1324_n 0.00815307f $X=4.83 $Y=1.155
+ $X2=0 $Y2=0
cc_749 N_A_811_379#_c_914_n N_A_879_55#_c_1353_n 0.029438f $X=8.78 $Y=2.035
+ $X2=0 $Y2=0
cc_750 N_A_811_379#_c_914_n N_A_879_55#_c_1328_n 0.00269274f $X=8.78 $Y=2.035
+ $X2=0 $Y2=0
cc_751 N_A_811_379#_c_1016_p N_A_879_55#_c_1328_n 2.61696e-19 $X=8.925 $Y=2.035
+ $X2=0 $Y2=0
cc_752 N_A_811_379#_c_1017_p N_A_879_55#_c_1328_n 0.013066f $X=8.925 $Y=2.035
+ $X2=0 $Y2=0
cc_753 N_A_811_379#_c_902_n N_A_879_55#_c_1329_n 0.0242401f $X=10.73 $Y=2.565
+ $X2=0 $Y2=0
cc_754 N_A_811_379#_M1002_d N_A_879_55#_c_1330_n 0.00363108f $X=10.18 $Y=0.47
+ $X2=0 $Y2=0
cc_755 N_A_811_379#_c_902_n N_A_879_55#_c_1330_n 0.00786375f $X=10.73 $Y=2.565
+ $X2=0 $Y2=0
cc_756 N_A_811_379#_c_1010_p N_A_879_55#_c_1330_n 0.0198333f $X=10.65 $Y=0.82
+ $X2=0 $Y2=0
cc_757 N_A_811_379#_c_902_n N_A_879_55#_c_1331_n 0.00429268f $X=10.73 $Y=2.565
+ $X2=0 $Y2=0
cc_758 N_A_811_379#_c_914_n N_B_c_1518_n 0.0082399f $X=8.78 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_759 N_A_811_379#_c_914_n N_B_c_1520_n 0.00720493f $X=8.78 $Y=2.035 $X2=0
+ $Y2=0
cc_760 N_A_811_379#_c_910_n N_B_c_1524_n 4.11423e-19 $X=10.645 $Y=2.65 $X2=0
+ $Y2=0
cc_761 N_A_811_379#_c_911_n N_B_c_1524_n 4.28224e-19 $X=9.11 $Y=2.65 $X2=0 $Y2=0
cc_762 N_A_811_379#_c_910_n N_B_M1019_g 0.0139f $X=10.645 $Y=2.65 $X2=0 $Y2=0
cc_763 N_A_811_379#_c_911_n N_B_M1019_g 7.32783e-19 $X=9.11 $Y=2.65 $X2=0 $Y2=0
cc_764 N_A_811_379#_c_1017_p N_B_M1019_g 0.0138481f $X=8.925 $Y=2.035 $X2=0
+ $Y2=0
cc_765 N_A_811_379#_c_902_n N_B_c_1513_n 2.09199e-19 $X=10.73 $Y=2.565 $X2=0
+ $Y2=0
cc_766 N_A_811_379#_c_914_n N_VPWR_M1031_d 0.00161776f $X=8.78 $Y=2.035 $X2=0
+ $Y2=0
cc_767 N_A_811_379#_c_914_n N_VPWR_c_1814_n 0.0300046f $X=8.78 $Y=2.035 $X2=0
+ $Y2=0
cc_768 N_A_811_379#_c_905_n N_VPWR_c_1821_n 0.00278271f $X=4.145 $Y=2.045 $X2=0
+ $Y2=0
cc_769 N_A_811_379#_c_905_n N_VPWR_c_1812_n 0.00363426f $X=4.145 $Y=2.045 $X2=0
+ $Y2=0
cc_770 N_A_811_379#_c_895_n N_A_644_104#_c_2022_n 0.00150592f $X=4.22 $Y=1.97
+ $X2=0 $Y2=0
cc_771 N_A_811_379#_c_908_n N_A_644_104#_c_2022_n 0.00204651f $X=6.195 $Y=1.715
+ $X2=0 $Y2=0
cc_772 N_A_811_379#_c_901_n N_A_644_104#_c_2022_n 0.00427488f $X=4.83 $Y=1.625
+ $X2=0 $Y2=0
cc_773 N_A_811_379#_c_903_n N_A_644_104#_c_2022_n 0.0177095f $X=5.785 $Y=1.54
+ $X2=0 $Y2=0
cc_774 N_A_811_379#_c_904_n N_A_644_104#_c_2022_n 0.00266701f $X=5.785 $Y=1.54
+ $X2=0 $Y2=0
cc_775 N_A_811_379#_c_914_n N_A_644_104#_c_2022_n 0.0495107f $X=8.78 $Y=2.035
+ $X2=0 $Y2=0
cc_776 N_A_811_379#_c_915_n N_A_644_104#_c_2022_n 0.023446f $X=5.665 $Y=2.035
+ $X2=0 $Y2=0
cc_777 N_A_811_379#_c_916_n N_A_644_104#_c_2022_n 0.00498335f $X=5.52 $Y=2.035
+ $X2=0 $Y2=0
cc_778 N_A_811_379#_c_908_n N_A_644_104#_c_2024_n 0.00136383f $X=6.195 $Y=1.715
+ $X2=0 $Y2=0
cc_779 N_A_811_379#_c_914_n N_A_644_104#_c_2024_n 0.0233656f $X=8.78 $Y=2.035
+ $X2=0 $Y2=0
cc_780 N_A_811_379#_c_908_n N_A_644_104#_c_2025_n 0.00153346f $X=6.195 $Y=1.715
+ $X2=0 $Y2=0
cc_781 N_A_811_379#_c_914_n N_A_644_104#_c_2025_n 2.27622e-19 $X=8.78 $Y=2.035
+ $X2=0 $Y2=0
cc_782 N_A_811_379#_c_905_n N_A_644_104#_c_2026_n 0.00193294f $X=4.145 $Y=2.045
+ $X2=0 $Y2=0
cc_783 N_A_811_379#_c_895_n N_A_644_104#_c_2026_n 0.00562526f $X=4.22 $Y=1.97
+ $X2=0 $Y2=0
cc_784 N_A_811_379#_c_896_n N_A_644_104#_c_2026_n 0.0010623f $X=4.655 $Y=1.895
+ $X2=0 $Y2=0
cc_785 N_A_811_379#_c_911_n N_A_1660_374#_c_2122_n 0.00781631f $X=9.11 $Y=2.65
+ $X2=0 $Y2=0
cc_786 N_A_811_379#_c_914_n N_A_1660_374#_c_2122_n 0.0236002f $X=8.78 $Y=2.035
+ $X2=0 $Y2=0
cc_787 N_A_811_379#_c_1016_p N_A_1660_374#_c_2122_n 0.00129223f $X=8.925
+ $Y=2.035 $X2=0 $Y2=0
cc_788 N_A_811_379#_c_910_n N_A_1660_374#_c_2123_n 0.120902f $X=10.645 $Y=2.65
+ $X2=0 $Y2=0
cc_789 N_A_811_379#_c_911_n N_A_1660_374#_c_2123_n 0.0258986f $X=9.11 $Y=2.65
+ $X2=0 $Y2=0
cc_790 N_A_811_379#_c_914_n N_A_1660_374#_c_2132_n 0.0146707f $X=8.78 $Y=2.035
+ $X2=0 $Y2=0
cc_791 N_A_811_379#_c_1016_p N_A_1660_374#_c_2132_n 0.00129223f $X=8.925
+ $Y=2.035 $X2=0 $Y2=0
cc_792 N_A_811_379#_c_1017_p N_A_1660_374#_c_2132_n 0.0293895f $X=8.925 $Y=2.035
+ $X2=0 $Y2=0
cc_793 N_A_811_379#_c_910_n N_A_1849_374#_M1019_d 0.024542f $X=10.645 $Y=2.65
+ $X2=0 $Y2=0
cc_794 N_A_811_379#_c_902_n N_A_1849_374#_M1019_d 0.0114591f $X=10.73 $Y=2.565
+ $X2=0 $Y2=0
cc_795 N_A_811_379#_c_902_n N_A_1849_374#_c_2208_n 0.00553169f $X=10.73 $Y=2.565
+ $X2=0 $Y2=0
cc_796 N_A_811_379#_c_910_n N_A_1849_374#_c_2224_n 0.00287247f $X=10.645 $Y=2.65
+ $X2=0 $Y2=0
cc_797 N_A_811_379#_c_910_n N_A_1849_374#_c_2218_n 0.00580459f $X=10.645 $Y=2.65
+ $X2=0 $Y2=0
cc_798 N_A_811_379#_c_902_n N_A_1849_374#_c_2218_n 0.0170813f $X=10.73 $Y=2.565
+ $X2=0 $Y2=0
cc_799 N_A_811_379#_c_902_n N_A_1849_374#_c_2227_n 6.59019e-19 $X=10.73 $Y=2.565
+ $X2=0 $Y2=0
cc_800 N_A_811_379#_c_910_n N_A_1849_374#_c_2220_n 0.0916455f $X=10.645 $Y=2.65
+ $X2=0 $Y2=0
cc_801 N_A_811_379#_c_902_n N_A_1849_374#_c_2220_n 0.044926f $X=10.73 $Y=2.565
+ $X2=0 $Y2=0
cc_802 N_A_811_379#_c_1016_p N_A_1849_374#_c_2220_n 0.00171921f $X=8.925
+ $Y=2.035 $X2=0 $Y2=0
cc_803 N_A_811_379#_c_899_n N_VGND_c_2327_n 0.0235892f $X=4.905 $Y=0.18 $X2=0
+ $Y2=0
cc_804 N_A_811_379#_c_898_n N_VGND_c_2330_n 0.024536f $X=5.69 $Y=0.18 $X2=0
+ $Y2=0
cc_805 N_A_811_379#_c_899_n N_VGND_c_2330_n 0.00603608f $X=4.905 $Y=0.18 $X2=0
+ $Y2=0
cc_806 N_A_1023_379#_c_1111_n N_A_879_55#_c_1314_n 0.00404913f $X=10.955
+ $Y=1.665 $X2=0 $Y2=0
cc_807 N_A_1023_379#_c_1108_n N_A_879_55#_M1004_g 0.00379675f $X=9.288 $Y=0.352
+ $X2=0 $Y2=0
cc_808 N_A_1023_379#_c_1109_n N_A_879_55#_c_1316_n 0.00916091f $X=10.985 $Y=0.34
+ $X2=0 $Y2=0
cc_809 N_A_1023_379#_c_1129_n N_A_879_55#_c_1334_n 2.51903e-19 $X=11.1 $Y=1.665
+ $X2=0 $Y2=0
cc_810 N_A_1023_379#_c_1130_n N_A_879_55#_c_1334_n 0.00394475f $X=11.1 $Y=1.665
+ $X2=0 $Y2=0
cc_811 N_A_1023_379#_c_1111_n N_A_879_55#_c_1318_n 0.00643359f $X=10.955
+ $Y=1.665 $X2=0 $Y2=0
cc_812 N_A_1023_379#_c_1129_n N_A_879_55#_c_1318_n 0.00128038f $X=11.1 $Y=1.665
+ $X2=0 $Y2=0
cc_813 N_A_1023_379#_c_1115_n N_A_879_55#_c_1318_n 0.00265776f $X=11.1 $Y=1.55
+ $X2=0 $Y2=0
cc_814 N_A_1023_379#_M1012_g N_A_879_55#_c_1319_n 0.00116683f $X=5.335 $Y=0.945
+ $X2=0 $Y2=0
cc_815 N_A_1023_379#_c_1100_n N_A_879_55#_c_1319_n 0.00930831f $X=6.265 $Y=1.25
+ $X2=0 $Y2=0
cc_816 N_A_1023_379#_c_1106_n N_A_879_55#_c_1319_n 0.0157559f $X=6.9 $Y=0.875
+ $X2=0 $Y2=0
cc_817 N_A_1023_379#_c_1107_n N_A_879_55#_c_1319_n 0.00282291f $X=6.9 $Y=0.875
+ $X2=0 $Y2=0
cc_818 N_A_1023_379#_c_1120_n N_A_879_55#_c_1336_n 0.00127274f $X=7.025 $Y=2.87
+ $X2=0 $Y2=0
cc_819 N_A_1023_379#_c_1106_n N_A_879_55#_c_1321_n 0.0268234f $X=6.9 $Y=0.875
+ $X2=0 $Y2=0
cc_820 N_A_1023_379#_c_1107_n N_A_879_55#_c_1321_n 0.0030771f $X=6.9 $Y=0.875
+ $X2=0 $Y2=0
cc_821 N_A_1023_379#_M1004_d N_A_879_55#_c_1323_n 0.00508114f $X=8.84 $Y=0.47
+ $X2=0 $Y2=0
cc_822 N_A_1023_379#_c_1111_n N_A_879_55#_c_1323_n 7.13018e-19 $X=10.955
+ $Y=1.665 $X2=0 $Y2=0
cc_823 N_A_1023_379#_M1004_d N_A_879_55#_c_1369_n 0.0144412f $X=8.84 $Y=0.47
+ $X2=0 $Y2=0
cc_824 N_A_1023_379#_c_1108_n N_A_879_55#_c_1369_n 0.0283607f $X=9.288 $Y=0.352
+ $X2=0 $Y2=0
cc_825 N_A_1023_379#_c_1109_n N_A_879_55#_c_1369_n 0.0504843f $X=10.985 $Y=0.34
+ $X2=0 $Y2=0
cc_826 N_A_1023_379#_M1003_g N_A_879_55#_c_1353_n 0.00684412f $X=7.025 $Y=2.285
+ $X2=0 $Y2=0
cc_827 N_A_1023_379#_c_1111_n N_A_879_55#_c_1353_n 0.00515509f $X=10.955
+ $Y=1.665 $X2=0 $Y2=0
cc_828 N_A_1023_379#_M1003_g N_A_879_55#_c_1325_n 0.00321135f $X=7.025 $Y=2.285
+ $X2=0 $Y2=0
cc_829 N_A_1023_379#_c_1105_n N_A_879_55#_c_1325_n 0.0040975f $X=6.925 $Y=1.325
+ $X2=0 $Y2=0
cc_830 N_A_1023_379#_c_1106_n N_A_879_55#_c_1325_n 0.0222312f $X=6.9 $Y=0.875
+ $X2=0 $Y2=0
cc_831 N_A_1023_379#_c_1107_n N_A_879_55#_c_1325_n 9.76449e-19 $X=6.9 $Y=0.875
+ $X2=0 $Y2=0
cc_832 N_A_1023_379#_c_1111_n N_A_879_55#_c_1325_n 0.0196475f $X=10.955 $Y=1.665
+ $X2=0 $Y2=0
cc_833 N_A_1023_379#_c_1112_n N_A_879_55#_c_1325_n 0.00218527f $X=7.105 $Y=1.665
+ $X2=0 $Y2=0
cc_834 N_A_1023_379#_c_1113_n N_A_879_55#_c_1325_n 0.00984568f $X=6.96 $Y=1.665
+ $X2=0 $Y2=0
cc_835 N_A_1023_379#_c_1106_n N_A_879_55#_c_1326_n 0.00674647f $X=6.9 $Y=0.875
+ $X2=0 $Y2=0
cc_836 N_A_1023_379#_c_1107_n N_A_879_55#_c_1326_n 7.6719e-19 $X=6.9 $Y=0.875
+ $X2=0 $Y2=0
cc_837 N_A_1023_379#_c_1111_n N_A_879_55#_c_1327_n 0.00595074f $X=10.955
+ $Y=1.665 $X2=0 $Y2=0
cc_838 N_A_1023_379#_c_1111_n N_A_879_55#_c_1328_n 0.0245964f $X=10.955 $Y=1.665
+ $X2=0 $Y2=0
cc_839 N_A_1023_379#_M1004_d N_A_879_55#_c_1414_n 8.29052e-19 $X=8.84 $Y=0.47
+ $X2=0 $Y2=0
cc_840 N_A_1023_379#_c_1108_n N_A_879_55#_c_1414_n 0.00612936f $X=9.288 $Y=0.352
+ $X2=0 $Y2=0
cc_841 N_A_1023_379#_c_1111_n N_A_879_55#_c_1329_n 0.0102318f $X=10.955 $Y=1.665
+ $X2=0 $Y2=0
cc_842 N_A_1023_379#_c_1111_n N_A_879_55#_c_1331_n 0.00739518f $X=10.955
+ $Y=1.665 $X2=0 $Y2=0
cc_843 N_A_1023_379#_c_1120_n N_B_c_1518_n 0.00530961f $X=7.025 $Y=2.87
+ $X2=-0.19 $Y2=-0.245
cc_844 N_A_1023_379#_c_1122_n N_B_c_1518_n 0.00238331f $X=7.025 $Y=1.79
+ $X2=-0.19 $Y2=-0.245
cc_845 N_A_1023_379#_M1003_g N_B_c_1518_n 0.0127864f $X=7.025 $Y=2.285 $X2=-0.19
+ $Y2=-0.245
cc_846 N_A_1023_379#_c_1111_n N_B_c_1518_n 0.00169461f $X=10.955 $Y=1.665
+ $X2=-0.19 $Y2=-0.245
cc_847 N_A_1023_379#_c_1105_n N_B_M1026_g 0.00640007f $X=6.925 $Y=1.325 $X2=0
+ $Y2=0
cc_848 N_A_1023_379#_c_1107_n N_B_M1026_g 0.00726866f $X=6.9 $Y=0.875 $X2=0
+ $Y2=0
cc_849 N_A_1023_379#_c_1111_n N_B_c_1509_n 0.0208981f $X=10.955 $Y=1.665 $X2=0
+ $Y2=0
cc_850 N_A_1023_379#_c_1111_n N_B_c_1520_n 0.0014599f $X=10.955 $Y=1.665 $X2=0
+ $Y2=0
cc_851 N_A_1023_379#_c_1111_n N_B_c_1510_n 0.00651167f $X=10.955 $Y=1.665 $X2=0
+ $Y2=0
cc_852 N_A_1023_379#_c_1111_n N_B_c_1526_n 0.0072595f $X=10.955 $Y=1.665 $X2=0
+ $Y2=0
cc_853 N_A_1023_379#_c_1109_n N_B_c_1511_n 0.00870518f $X=10.985 $Y=0.34 $X2=0
+ $Y2=0
cc_854 N_A_1023_379#_c_1110_n N_B_c_1511_n 7.92841e-19 $X=9.385 $Y=0.352 $X2=0
+ $Y2=0
cc_855 N_A_1023_379#_c_1109_n N_B_M1027_g 0.00234457f $X=10.985 $Y=0.34 $X2=0
+ $Y2=0
cc_856 N_A_1023_379#_c_1115_n N_B_M1027_g 0.0209695f $X=11.1 $Y=1.55 $X2=0 $Y2=0
cc_857 N_A_1023_379#_c_1129_n N_B_c_1513_n 0.00274997f $X=11.1 $Y=1.665 $X2=0
+ $Y2=0
cc_858 N_A_1023_379#_c_1130_n N_B_c_1513_n 0.00216342f $X=11.1 $Y=1.665 $X2=0
+ $Y2=0
cc_859 N_A_1023_379#_c_1115_n N_B_c_1513_n 3.91215e-19 $X=11.1 $Y=1.55 $X2=0
+ $Y2=0
cc_860 N_A_1023_379#_c_1129_n N_B_c_1532_n 7.9617e-19 $X=11.1 $Y=1.665 $X2=0
+ $Y2=0
cc_861 N_A_1023_379#_c_1130_n N_B_c_1532_n 0.00154056f $X=11.1 $Y=1.665 $X2=0
+ $Y2=0
cc_862 N_A_1023_379#_c_1125_n N_B_M1016_g 0.00464865f $X=11.07 $Y=1.98 $X2=0
+ $Y2=0
cc_863 N_A_1023_379#_c_1129_n N_B_M1016_g 4.03853e-19 $X=11.1 $Y=1.665 $X2=0
+ $Y2=0
cc_864 N_A_1023_379#_c_1103_n N_B_c_1514_n 0.00518782f $X=7.025 $Y=1.7 $X2=0
+ $Y2=0
cc_865 N_A_1023_379#_c_1111_n N_B_c_1514_n 0.00639148f $X=10.955 $Y=1.665 $X2=0
+ $Y2=0
cc_866 N_A_1023_379#_c_1113_n N_B_c_1514_n 2.24991e-19 $X=6.96 $Y=1.665 $X2=0
+ $Y2=0
cc_867 N_A_1023_379#_c_1130_n N_B_c_1515_n 2.25647e-19 $X=11.1 $Y=1.665 $X2=0
+ $Y2=0
cc_868 N_A_1023_379#_c_1111_n B 0.0125374f $X=10.955 $Y=1.665 $X2=0 $Y2=0
cc_869 N_A_1023_379#_c_1111_n N_B_c_1517_n 0.00347971f $X=10.955 $Y=1.665 $X2=0
+ $Y2=0
cc_870 N_A_1023_379#_c_1109_n N_A_2342_48#_c_1666_n 0.00235964f $X=10.985
+ $Y=0.34 $X2=0 $Y2=0
cc_871 N_A_1023_379#_c_1121_n N_VPWR_c_1814_n 0.00338783f $X=7.025 $Y=3.075
+ $X2=0 $Y2=0
cc_872 N_A_1023_379#_c_1111_n N_VPWR_c_1814_n 0.0131007f $X=10.955 $Y=1.665
+ $X2=0 $Y2=0
cc_873 N_A_1023_379#_c_1118_n N_VPWR_c_1821_n 0.0431787f $X=5.295 $Y=3.15 $X2=0
+ $Y2=0
cc_874 N_A_1023_379#_c_1117_n N_VPWR_c_1812_n 0.049114f $X=6.935 $Y=3.15 $X2=0
+ $Y2=0
cc_875 N_A_1023_379#_c_1118_n N_VPWR_c_1812_n 0.00674544f $X=5.295 $Y=3.15 $X2=0
+ $Y2=0
cc_876 N_A_1023_379#_c_1100_n N_A_644_104#_c_2020_n 0.00140926f $X=6.265 $Y=1.25
+ $X2=0 $Y2=0
cc_877 N_A_1023_379#_c_1101_n N_A_644_104#_c_2020_n 0.0131359f $X=6.735 $Y=1.325
+ $X2=0 $Y2=0
cc_878 N_A_1023_379#_c_1103_n N_A_644_104#_c_2020_n 8.05667e-19 $X=7.025 $Y=1.7
+ $X2=0 $Y2=0
cc_879 N_A_1023_379#_c_1106_n N_A_644_104#_c_2020_n 0.0491798f $X=6.9 $Y=0.875
+ $X2=0 $Y2=0
cc_880 N_A_1023_379#_c_1107_n N_A_644_104#_c_2020_n 0.0041353f $X=6.9 $Y=0.875
+ $X2=0 $Y2=0
cc_881 N_A_1023_379#_c_1114_n N_A_644_104#_c_2020_n 0.00899568f $X=6.96 $Y=1.55
+ $X2=0 $Y2=0
cc_882 N_A_1023_379#_M1012_g N_A_644_104#_c_2022_n 0.00831542f $X=5.335 $Y=0.945
+ $X2=0 $Y2=0
cc_883 N_A_1023_379#_c_1102_n N_A_644_104#_c_2022_n 0.00145597f $X=6.34 $Y=1.325
+ $X2=0 $Y2=0
cc_884 N_A_1023_379#_c_1104_n N_A_644_104#_c_2022_n 0.00128901f $X=5.335 $Y=1.97
+ $X2=0 $Y2=0
cc_885 N_A_1023_379#_c_1102_n N_A_644_104#_c_2024_n 0.00219086f $X=6.34 $Y=1.325
+ $X2=0 $Y2=0
cc_886 N_A_1023_379#_c_1112_n N_A_644_104#_c_2024_n 0.0225507f $X=7.105 $Y=1.665
+ $X2=0 $Y2=0
cc_887 N_A_1023_379#_c_1113_n N_A_644_104#_c_2024_n 9.8705e-19 $X=6.96 $Y=1.665
+ $X2=0 $Y2=0
cc_888 N_A_1023_379#_c_1101_n N_A_644_104#_c_2025_n 9.28054e-19 $X=6.735
+ $Y=1.325 $X2=0 $Y2=0
cc_889 N_A_1023_379#_c_1103_n N_A_644_104#_c_2025_n 7.95166e-19 $X=7.025 $Y=1.7
+ $X2=0 $Y2=0
cc_890 N_A_1023_379#_c_1112_n N_A_644_104#_c_2025_n 9.88639e-19 $X=7.105
+ $Y=1.665 $X2=0 $Y2=0
cc_891 N_A_1023_379#_c_1113_n N_A_644_104#_c_2025_n 0.0112038f $X=6.96 $Y=1.665
+ $X2=0 $Y2=0
cc_892 N_A_1023_379#_c_1125_n N_A_1660_374#_c_2123_n 0.0132728f $X=11.07 $Y=1.98
+ $X2=0 $Y2=0
cc_893 N_A_1023_379#_c_1115_n N_A_1660_374#_c_2117_n 0.0270149f $X=11.1 $Y=1.55
+ $X2=0 $Y2=0
cc_894 N_A_1023_379#_c_1125_n N_A_1660_374#_c_2118_n 0.0330572f $X=11.07 $Y=1.98
+ $X2=0 $Y2=0
cc_895 N_A_1023_379#_c_1129_n N_A_1660_374#_c_2118_n 0.00661419f $X=11.1
+ $Y=1.665 $X2=0 $Y2=0
cc_896 N_A_1023_379#_c_1130_n N_A_1660_374#_c_2118_n 0.0152718f $X=11.1 $Y=1.665
+ $X2=0 $Y2=0
cc_897 N_A_1023_379#_c_1109_n N_A_1660_374#_c_2119_n 0.005061f $X=10.985 $Y=0.34
+ $X2=0 $Y2=0
cc_898 N_A_1023_379#_c_1115_n N_A_1660_374#_c_2119_n 0.00375546f $X=11.1 $Y=1.55
+ $X2=0 $Y2=0
cc_899 N_A_1023_379#_c_1111_n N_A_1660_374#_c_2120_n 0.00541281f $X=10.955
+ $Y=1.665 $X2=0 $Y2=0
cc_900 N_A_1023_379#_c_1111_n N_A_1660_374#_c_2132_n 0.00362103f $X=10.955
+ $Y=1.665 $X2=0 $Y2=0
cc_901 N_A_1023_379#_c_1111_n N_A_1660_374#_c_2121_n 0.0133101f $X=10.955
+ $Y=1.665 $X2=0 $Y2=0
cc_902 N_A_1023_379#_c_1111_n N_A_1849_374#_c_2208_n 0.0330113f $X=10.955
+ $Y=1.665 $X2=0 $Y2=0
cc_903 N_A_1023_379#_c_1111_n N_A_1849_374#_c_2224_n 0.053525f $X=10.955
+ $Y=1.665 $X2=0 $Y2=0
cc_904 N_A_1023_379#_M1013_d N_A_1849_374#_c_2218_n 0.00583831f $X=10.92 $Y=1.84
+ $X2=0 $Y2=0
cc_905 N_A_1023_379#_c_1125_n N_A_1849_374#_c_2218_n 0.0172139f $X=11.07 $Y=1.98
+ $X2=0 $Y2=0
cc_906 N_A_1023_379#_c_1111_n N_A_1849_374#_c_2218_n 0.0354957f $X=10.955
+ $Y=1.665 $X2=0 $Y2=0
cc_907 N_A_1023_379#_c_1129_n N_A_1849_374#_c_2218_n 0.0236637f $X=11.1 $Y=1.665
+ $X2=0 $Y2=0
cc_908 N_A_1023_379#_c_1130_n N_A_1849_374#_c_2218_n 4.39572e-19 $X=11.1
+ $Y=1.665 $X2=0 $Y2=0
cc_909 N_A_1023_379#_c_1111_n N_A_1849_374#_c_2220_n 0.0272966f $X=10.955
+ $Y=1.665 $X2=0 $Y2=0
cc_910 N_A_1023_379#_c_1108_n N_VGND_c_2324_n 0.13437f $X=9.288 $Y=0.352 $X2=0
+ $Y2=0
cc_911 N_A_1023_379#_c_1109_n N_VGND_c_2324_n 0.0121867f $X=10.985 $Y=0.34 $X2=0
+ $Y2=0
cc_912 N_A_1023_379#_c_1100_n N_VGND_c_2327_n 6.51701e-19 $X=6.265 $Y=1.25 $X2=0
+ $Y2=0
cc_913 N_A_1023_379#_M1004_d N_VGND_c_2330_n 0.00399728f $X=8.84 $Y=0.47 $X2=0
+ $Y2=0
cc_914 N_A_1023_379#_c_1108_n N_VGND_c_2330_n 0.0786214f $X=9.288 $Y=0.352 $X2=0
+ $Y2=0
cc_915 N_A_1023_379#_c_1109_n N_VGND_c_2330_n 0.00660921f $X=10.985 $Y=0.34
+ $X2=0 $Y2=0
cc_916 N_A_879_55#_c_1336_n N_B_c_1518_n 0.00818511f $X=7.335 $Y=2.76 $X2=-0.19
+ $Y2=-0.245
cc_917 N_A_879_55#_c_1353_n N_B_c_1518_n 0.00111743f $X=7.335 $Y=2.05 $X2=-0.19
+ $Y2=-0.245
cc_918 N_A_879_55#_c_1325_n N_B_c_1518_n 0.00405788f $X=7.335 $Y=1.95 $X2=-0.19
+ $Y2=-0.245
cc_919 N_A_879_55#_c_1319_n N_B_M1026_g 0.00474255f $X=7.235 $Y=0.34 $X2=0 $Y2=0
cc_920 N_A_879_55#_c_1320_n N_B_M1026_g 0.00758638f $X=7.4 $Y=0.515 $X2=0 $Y2=0
cc_921 N_A_879_55#_c_1321_n N_B_M1026_g 0.00737435f $X=7.4 $Y=0.965 $X2=0 $Y2=0
cc_922 N_A_879_55#_c_1322_n N_B_M1026_g 0.0141003f $X=8.805 $Y=0.705 $X2=0 $Y2=0
cc_923 N_A_879_55#_c_1325_n N_B_M1026_g 0.00660393f $X=7.335 $Y=1.95 $X2=0 $Y2=0
cc_924 N_A_879_55#_c_1326_n N_B_M1026_g 0.00122503f $X=7.4 $Y=0.705 $X2=0 $Y2=0
cc_925 N_A_879_55#_c_1327_n N_B_M1026_g 0.00433884f $X=7.4 $Y=1.13 $X2=0 $Y2=0
cc_926 N_A_879_55#_c_1314_n N_B_c_1509_n 0.00613107f $X=8.67 $Y=1.795 $X2=0
+ $Y2=0
cc_927 N_A_879_55#_c_1328_n N_B_c_1509_n 2.06293e-19 $X=8.89 $Y=1.545 $X2=0
+ $Y2=0
cc_928 N_A_879_55#_c_1314_n N_B_c_1520_n 0.0220956f $X=8.67 $Y=1.795 $X2=0 $Y2=0
cc_929 N_A_879_55#_c_1325_n N_B_c_1520_n 4.25576e-19 $X=7.335 $Y=1.95 $X2=0
+ $Y2=0
cc_930 N_A_879_55#_c_1314_n N_B_c_1521_n 0.0076828f $X=8.67 $Y=1.795 $X2=0 $Y2=0
cc_931 N_A_879_55#_c_1314_n N_B_c_1510_n 0.0132713f $X=8.67 $Y=1.795 $X2=0 $Y2=0
cc_932 N_A_879_55#_c_1314_n N_B_c_1524_n 0.00211763f $X=8.67 $Y=1.795 $X2=0
+ $Y2=0
cc_933 N_A_879_55#_c_1314_n N_B_c_1526_n 0.00386809f $X=8.67 $Y=1.795 $X2=0
+ $Y2=0
cc_934 N_A_879_55#_c_1314_n N_B_M1019_g 0.0188135f $X=8.67 $Y=1.795 $X2=0 $Y2=0
cc_935 N_A_879_55#_c_1334_n N_B_c_1528_n 0.00661634f $X=10.845 $Y=1.765 $X2=0
+ $Y2=0
cc_936 N_A_879_55#_M1004_g N_B_c_1511_n 0.0137917f $X=8.765 $Y=0.79 $X2=0 $Y2=0
cc_937 N_A_879_55#_c_1316_n N_B_c_1511_n 0.0145345f $X=10.105 $Y=1.22 $X2=0
+ $Y2=0
cc_938 N_A_879_55#_c_1323_n N_B_c_1511_n 0.00465173f $X=8.89 $Y=1.38 $X2=0 $Y2=0
cc_939 N_A_879_55#_c_1369_n N_B_c_1511_n 0.016389f $X=10.145 $Y=0.705 $X2=0
+ $Y2=0
cc_940 N_A_879_55#_c_1330_n N_B_c_1511_n 8.99371e-19 $X=10.31 $Y=1.22 $X2=0
+ $Y2=0
cc_941 N_A_879_55#_c_1318_n N_B_c_1513_n 0.0122493f $X=10.845 $Y=1.475 $X2=0
+ $Y2=0
cc_942 N_A_879_55#_c_1334_n N_B_c_1530_n 0.00253032f $X=10.845 $Y=1.765 $X2=0
+ $Y2=0
cc_943 N_A_879_55#_c_1334_n N_B_M1016_g 0.0111043f $X=10.845 $Y=1.765 $X2=0
+ $Y2=0
cc_944 N_A_879_55#_c_1325_n N_B_c_1514_n 0.00612962f $X=7.335 $Y=1.95 $X2=0
+ $Y2=0
cc_945 N_A_879_55#_c_1327_n N_B_c_1514_n 0.00147078f $X=7.4 $Y=1.13 $X2=0 $Y2=0
cc_946 N_A_879_55#_c_1318_n N_B_c_1515_n 0.00434234f $X=10.845 $Y=1.475 $X2=0
+ $Y2=0
cc_947 N_A_879_55#_M1004_g B 2.69431e-19 $X=8.765 $Y=0.79 $X2=0 $Y2=0
cc_948 N_A_879_55#_c_1323_n B 0.0151952f $X=8.89 $Y=1.38 $X2=0 $Y2=0
cc_949 N_A_879_55#_c_1369_n B 0.0129757f $X=10.145 $Y=0.705 $X2=0 $Y2=0
cc_950 N_A_879_55#_c_1328_n B 0.0138134f $X=8.89 $Y=1.545 $X2=0 $Y2=0
cc_951 N_A_879_55#_M1004_g N_B_c_1517_n 0.0132713f $X=8.765 $Y=0.79 $X2=0 $Y2=0
cc_952 N_A_879_55#_c_1323_n N_B_c_1517_n 0.00110062f $X=8.89 $Y=1.38 $X2=0 $Y2=0
cc_953 N_A_879_55#_c_1369_n N_B_c_1517_n 0.0035026f $X=10.145 $Y=0.705 $X2=0
+ $Y2=0
cc_954 N_A_879_55#_c_1328_n N_B_c_1517_n 0.00305376f $X=8.89 $Y=1.545 $X2=0
+ $Y2=0
cc_955 N_A_879_55#_c_1331_n N_B_c_1517_n 0.0145345f $X=10.475 $Y=1.385 $X2=0
+ $Y2=0
cc_956 N_A_879_55#_c_1325_n N_VPWR_c_1814_n 0.0461644f $X=7.335 $Y=1.95 $X2=0
+ $Y2=0
cc_957 N_A_879_55#_c_1336_n N_VPWR_c_1821_n 0.0119397f $X=7.335 $Y=2.76 $X2=0
+ $Y2=0
cc_958 N_A_879_55#_c_1336_n N_VPWR_c_1812_n 0.0116912f $X=7.335 $Y=2.76 $X2=0
+ $Y2=0
cc_959 N_A_879_55#_c_1319_n N_A_644_104#_c_2020_n 0.00955123f $X=7.235 $Y=0.34
+ $X2=0 $Y2=0
cc_960 N_A_879_55#_c_1326_n N_A_644_104#_c_2020_n 0.00123143f $X=7.4 $Y=0.705
+ $X2=0 $Y2=0
cc_961 N_A_879_55#_c_1322_n N_A_1660_374#_M1004_s 0.0101563f $X=8.805 $Y=0.705
+ $X2=-0.19 $Y2=-0.245
cc_962 N_A_879_55#_c_1314_n N_A_1660_374#_c_2122_n 0.0120528f $X=8.67 $Y=1.795
+ $X2=0 $Y2=0
cc_963 N_A_879_55#_c_1314_n N_A_1660_374#_c_2123_n 0.00328606f $X=8.67 $Y=1.795
+ $X2=0 $Y2=0
cc_964 N_A_879_55#_c_1334_n N_A_1660_374#_c_2123_n 0.00288846f $X=10.845
+ $Y=1.765 $X2=0 $Y2=0
cc_965 N_A_879_55#_c_1314_n N_A_1660_374#_c_2120_n 0.00300193f $X=8.67 $Y=1.795
+ $X2=0 $Y2=0
cc_966 N_A_879_55#_M1004_g N_A_1660_374#_c_2120_n 0.00509805f $X=8.765 $Y=0.79
+ $X2=0 $Y2=0
cc_967 N_A_879_55#_c_1321_n N_A_1660_374#_c_2120_n 0.00527168f $X=7.4 $Y=0.965
+ $X2=0 $Y2=0
cc_968 N_A_879_55#_c_1322_n N_A_1660_374#_c_2120_n 0.0350598f $X=8.805 $Y=0.705
+ $X2=0 $Y2=0
cc_969 N_A_879_55#_c_1323_n N_A_1660_374#_c_2120_n 0.0127597f $X=8.89 $Y=1.38
+ $X2=0 $Y2=0
cc_970 N_A_879_55#_c_1325_n N_A_1660_374#_c_2120_n 0.00243034f $X=7.335 $Y=1.95
+ $X2=0 $Y2=0
cc_971 N_A_879_55#_c_1328_n N_A_1660_374#_c_2120_n 0.00915244f $X=8.89 $Y=1.545
+ $X2=0 $Y2=0
cc_972 N_A_879_55#_c_1314_n N_A_1660_374#_c_2132_n 0.00294666f $X=8.67 $Y=1.795
+ $X2=0 $Y2=0
cc_973 N_A_879_55#_c_1328_n N_A_1660_374#_c_2132_n 0.00470068f $X=8.89 $Y=1.545
+ $X2=0 $Y2=0
cc_974 N_A_879_55#_c_1314_n N_A_1660_374#_c_2121_n 0.00487614f $X=8.67 $Y=1.795
+ $X2=0 $Y2=0
cc_975 N_A_879_55#_M1004_g N_A_1660_374#_c_2121_n 0.00301106f $X=8.765 $Y=0.79
+ $X2=0 $Y2=0
cc_976 N_A_879_55#_c_1323_n N_A_1660_374#_c_2121_n 0.0057164f $X=8.89 $Y=1.38
+ $X2=0 $Y2=0
cc_977 N_A_879_55#_c_1325_n N_A_1660_374#_c_2121_n 0.0125531f $X=7.335 $Y=1.95
+ $X2=0 $Y2=0
cc_978 N_A_879_55#_c_1328_n N_A_1660_374#_c_2121_n 0.024395f $X=8.89 $Y=1.545
+ $X2=0 $Y2=0
cc_979 N_A_879_55#_c_1369_n N_A_1849_374#_M1030_d 0.00772805f $X=10.145 $Y=0.705
+ $X2=-0.19 $Y2=-0.245
cc_980 N_A_879_55#_c_1316_n N_A_1849_374#_c_2208_n 0.00577593f $X=10.105 $Y=1.22
+ $X2=0 $Y2=0
cc_981 N_A_879_55#_c_1323_n N_A_1849_374#_c_2208_n 0.00402151f $X=8.89 $Y=1.38
+ $X2=0 $Y2=0
cc_982 N_A_879_55#_c_1369_n N_A_1849_374#_c_2208_n 0.0265229f $X=10.145 $Y=0.705
+ $X2=0 $Y2=0
cc_983 N_A_879_55#_c_1328_n N_A_1849_374#_c_2208_n 0.00314532f $X=8.89 $Y=1.545
+ $X2=0 $Y2=0
cc_984 N_A_879_55#_c_1330_n N_A_1849_374#_c_2208_n 0.0394249f $X=10.31 $Y=1.22
+ $X2=0 $Y2=0
cc_985 N_A_879_55#_c_1334_n N_A_1849_374#_c_2218_n 0.00543358f $X=10.845
+ $Y=1.765 $X2=0 $Y2=0
cc_986 N_A_879_55#_c_1318_n N_A_1849_374#_c_2218_n 2.30869e-19 $X=10.845
+ $Y=1.475 $X2=0 $Y2=0
cc_987 N_A_879_55#_c_1334_n N_A_1849_374#_c_2220_n 0.00326114f $X=10.845
+ $Y=1.765 $X2=0 $Y2=0
cc_988 N_A_879_55#_c_1329_n N_A_1849_374#_c_2220_n 0.0132213f $X=10.31 $Y=1.385
+ $X2=0 $Y2=0
cc_989 N_A_879_55#_c_1331_n N_A_1849_374#_c_2220_n 0.00741463f $X=10.475
+ $Y=1.385 $X2=0 $Y2=0
cc_990 N_A_879_55#_c_1322_n N_VGND_M1026_d 0.0166098f $X=8.805 $Y=0.705 $X2=0
+ $Y2=0
cc_991 N_A_879_55#_M1004_g N_VGND_c_2319_n 0.00257286f $X=8.765 $Y=0.79 $X2=0
+ $Y2=0
cc_992 N_A_879_55#_c_1319_n N_VGND_c_2319_n 0.0114117f $X=7.235 $Y=0.34 $X2=0
+ $Y2=0
cc_993 N_A_879_55#_c_1322_n N_VGND_c_2319_n 0.0248636f $X=8.805 $Y=0.705 $X2=0
+ $Y2=0
cc_994 N_A_879_55#_M1004_g N_VGND_c_2324_n 0.00387786f $X=8.765 $Y=0.79 $X2=0
+ $Y2=0
cc_995 N_A_879_55#_c_1316_n N_VGND_c_2324_n 7.64118e-19 $X=10.105 $Y=1.22 $X2=0
+ $Y2=0
cc_996 N_A_879_55#_c_1322_n N_VGND_c_2324_n 0.0127782f $X=8.805 $Y=0.705 $X2=0
+ $Y2=0
cc_997 N_A_879_55#_c_1414_n N_VGND_c_2324_n 0.00121079f $X=8.89 $Y=0.705 $X2=0
+ $Y2=0
cc_998 N_A_879_55#_c_1319_n N_VGND_c_2327_n 0.185632f $X=7.235 $Y=0.34 $X2=0
+ $Y2=0
cc_999 N_A_879_55#_c_1322_n N_VGND_c_2327_n 0.00265735f $X=8.805 $Y=0.705 $X2=0
+ $Y2=0
cc_1000 N_A_879_55#_c_1324_n N_VGND_c_2327_n 0.0168534f $X=4.58 $Y=0.34 $X2=0
+ $Y2=0
cc_1001 N_A_879_55#_M1004_g N_VGND_c_2330_n 0.00514438f $X=8.765 $Y=0.79 $X2=0
+ $Y2=0
cc_1002 N_A_879_55#_c_1319_n N_VGND_c_2330_n 0.103281f $X=7.235 $Y=0.34 $X2=0
+ $Y2=0
cc_1003 N_A_879_55#_c_1322_n N_VGND_c_2330_n 0.0271433f $X=8.805 $Y=0.705 $X2=0
+ $Y2=0
cc_1004 N_A_879_55#_c_1324_n N_VGND_c_2330_n 0.00946983f $X=4.58 $Y=0.34 $X2=0
+ $Y2=0
cc_1005 N_A_879_55#_c_1414_n N_VGND_c_2330_n 0.00293042f $X=8.89 $Y=0.705 $X2=0
+ $Y2=0
cc_1006 N_B_c_1530_n N_A_2342_48#_c_1673_n 0.0122727f $X=11.295 $Y=2.85 $X2=0
+ $Y2=0
cc_1007 N_B_M1016_g N_A_2342_48#_c_1673_n 0.00827926f $X=11.295 $Y=2.26 $X2=0
+ $Y2=0
cc_1008 N_B_c_1515_n N_A_2342_48#_c_1665_n 0.0137157f $X=11.292 $Y=1.5 $X2=0
+ $Y2=0
cc_1009 N_B_M1027_g N_A_2342_48#_c_1666_n 0.0175303f $X=11.275 $Y=0.79 $X2=0
+ $Y2=0
cc_1010 N_B_c_1518_n N_VPWR_c_1814_n 0.00925072f $X=7.56 $Y=1.71 $X2=0 $Y2=0
cc_1011 N_B_c_1509_n N_VPWR_c_1814_n 0.010544f $X=8.055 $Y=1.635 $X2=0 $Y2=0
cc_1012 N_B_c_1520_n N_VPWR_c_1814_n 0.0181734f $X=8.13 $Y=3.075 $X2=0 $Y2=0
cc_1013 N_B_c_1528_n N_VPWR_c_1816_n 0.00171071f $X=11.205 $Y=3.15 $X2=0 $Y2=0
cc_1014 N_B_c_1522_n N_VPWR_c_1818_n 0.0718629f $X=8.205 $Y=3.15 $X2=0 $Y2=0
cc_1015 N_B_c_1518_n N_VPWR_c_1821_n 0.00523995f $X=7.56 $Y=1.71 $X2=0 $Y2=0
cc_1016 N_B_c_1518_n N_VPWR_c_1812_n 0.00528353f $X=7.56 $Y=1.71 $X2=0 $Y2=0
cc_1017 N_B_c_1521_n N_VPWR_c_1812_n 0.0205955f $X=9.08 $Y=3.15 $X2=0 $Y2=0
cc_1018 N_B_c_1522_n N_VPWR_c_1812_n 0.0101867f $X=8.205 $Y=3.15 $X2=0 $Y2=0
cc_1019 N_B_c_1528_n N_VPWR_c_1812_n 0.051961f $X=11.205 $Y=3.15 $X2=0 $Y2=0
cc_1020 N_B_c_1535_n N_VPWR_c_1812_n 0.00441592f $X=9.17 $Y=3.15 $X2=0 $Y2=0
cc_1021 N_B_c_1520_n N_A_1660_374#_c_2122_n 0.0213056f $X=8.13 $Y=3.075 $X2=0
+ $Y2=0
cc_1022 N_B_c_1524_n N_A_1660_374#_c_2122_n 0.0020911f $X=9.17 $Y=2.875 $X2=0
+ $Y2=0
cc_1023 N_B_M1019_g N_A_1660_374#_c_2122_n 2.29061e-19 $X=9.17 $Y=2.29 $X2=0
+ $Y2=0
cc_1024 N_B_c_1521_n N_A_1660_374#_c_2123_n 0.0067189f $X=9.08 $Y=3.15 $X2=0
+ $Y2=0
cc_1025 N_B_c_1525_n N_A_1660_374#_c_2123_n 0.014835f $X=9.17 $Y=3.075 $X2=0
+ $Y2=0
cc_1026 N_B_c_1528_n N_A_1660_374#_c_2123_n 0.039059f $X=11.205 $Y=3.15 $X2=0
+ $Y2=0
cc_1027 N_B_c_1531_n N_A_1660_374#_c_2123_n 0.0184827f $X=11.295 $Y=3.075 $X2=0
+ $Y2=0
cc_1028 N_B_c_1520_n N_A_1660_374#_c_2124_n 0.00596594f $X=8.13 $Y=3.075 $X2=0
+ $Y2=0
cc_1029 N_B_c_1521_n N_A_1660_374#_c_2124_n 0.0108374f $X=9.08 $Y=3.15 $X2=0
+ $Y2=0
cc_1030 N_B_c_1522_n N_A_1660_374#_c_2124_n 2.99808e-19 $X=8.205 $Y=3.15 $X2=0
+ $Y2=0
cc_1031 N_B_M1027_g N_A_1660_374#_c_2117_n 0.00218177f $X=11.275 $Y=0.79 $X2=0
+ $Y2=0
cc_1032 N_B_c_1530_n N_A_1660_374#_c_2118_n 0.00440141f $X=11.295 $Y=2.85 $X2=0
+ $Y2=0
cc_1033 N_B_M1016_g N_A_1660_374#_c_2118_n 0.00330146f $X=11.295 $Y=2.26 $X2=0
+ $Y2=0
cc_1034 N_B_c_1515_n N_A_1660_374#_c_2118_n 0.00408817f $X=11.292 $Y=1.5 $X2=0
+ $Y2=0
cc_1035 N_B_M1027_g N_A_1660_374#_c_2119_n 0.00470921f $X=11.275 $Y=0.79 $X2=0
+ $Y2=0
cc_1036 N_B_M1026_g N_A_1660_374#_c_2120_n 0.00426391f $X=7.615 $Y=0.74 $X2=0
+ $Y2=0
cc_1037 N_B_c_1520_n N_A_1660_374#_c_2132_n 0.00527614f $X=8.13 $Y=3.075 $X2=0
+ $Y2=0
cc_1038 N_B_M1019_g N_A_1660_374#_c_2132_n 2.97965e-19 $X=9.17 $Y=2.29 $X2=0
+ $Y2=0
cc_1039 N_B_c_1518_n N_A_1660_374#_c_2121_n 4.40765e-19 $X=7.56 $Y=1.71 $X2=0
+ $Y2=0
cc_1040 N_B_M1026_g N_A_1660_374#_c_2121_n 0.00571899f $X=7.615 $Y=0.74 $X2=0
+ $Y2=0
cc_1041 N_B_c_1509_n N_A_1660_374#_c_2121_n 0.00564986f $X=8.055 $Y=1.635 $X2=0
+ $Y2=0
cc_1042 N_B_c_1520_n N_A_1660_374#_c_2121_n 0.00382019f $X=8.13 $Y=3.075 $X2=0
+ $Y2=0
cc_1043 N_B_c_1510_n N_A_1849_374#_c_2208_n 0.00466121f $X=9.17 $Y=1.705 $X2=0
+ $Y2=0
cc_1044 N_B_M1019_g N_A_1849_374#_c_2208_n 2.77542e-19 $X=9.17 $Y=2.29 $X2=0
+ $Y2=0
cc_1045 N_B_c_1511_n N_A_1849_374#_c_2208_n 0.00620618f $X=9.515 $Y=1.22 $X2=0
+ $Y2=0
cc_1046 B N_A_1849_374#_c_2208_n 0.0292399f $X=9.275 $Y=1.21 $X2=0 $Y2=0
cc_1047 N_B_c_1532_n N_A_1849_374#_c_2218_n 3.80553e-19 $X=11.295 $Y=1.765 $X2=0
+ $Y2=0
cc_1048 N_B_M1016_g N_A_1849_374#_c_2218_n 0.0116096f $X=11.295 $Y=2.26 $X2=0
+ $Y2=0
cc_1049 N_B_M1019_g N_A_1849_374#_c_2220_n 0.0132933f $X=9.17 $Y=2.29 $X2=0
+ $Y2=0
cc_1050 B N_A_1849_374#_c_2220_n 0.00767772f $X=9.275 $Y=1.21 $X2=0 $Y2=0
cc_1051 N_B_c_1517_n N_A_1849_374#_c_2220_n 0.00642818f $X=9.515 $Y=1.385 $X2=0
+ $Y2=0
cc_1052 N_B_M1026_g N_VGND_c_2319_n 0.00471565f $X=7.615 $Y=0.74 $X2=0 $Y2=0
cc_1053 N_B_c_1511_n N_VGND_c_2324_n 7.64118e-19 $X=9.515 $Y=1.22 $X2=0 $Y2=0
cc_1054 N_B_M1027_g N_VGND_c_2324_n 0.00507111f $X=11.275 $Y=0.79 $X2=0 $Y2=0
cc_1055 N_B_M1026_g N_VGND_c_2327_n 0.0031683f $X=7.615 $Y=0.74 $X2=0 $Y2=0
cc_1056 N_B_M1026_g N_VGND_c_2330_n 0.00409665f $X=7.615 $Y=0.74 $X2=0 $Y2=0
cc_1057 N_B_M1027_g N_VGND_c_2330_n 0.00514438f $X=11.275 $Y=0.79 $X2=0 $Y2=0
cc_1058 N_A_2342_48#_c_1667_n N_A_M1014_g 0.0161142f $X=13.475 $Y=1.215 $X2=0
+ $Y2=0
cc_1059 N_A_2342_48#_c_1668_n N_A_M1014_g 8.02192e-19 $X=13.64 $Y=0.515 $X2=0
+ $Y2=0
cc_1060 N_A_2342_48#_c_1669_n N_A_M1014_g 0.00152361f $X=12.415 $Y=1.215 $X2=0
+ $Y2=0
cc_1061 N_A_2342_48#_c_1670_n N_A_M1014_g 0.0191364f $X=12.415 $Y=1.385 $X2=0
+ $Y2=0
cc_1062 N_A_2342_48#_c_1675_n N_A_c_1751_n 0.00843592f $X=13.635 $Y=2.815 $X2=0
+ $Y2=0
cc_1063 N_A_2342_48#_c_1678_n N_A_c_1751_n 0.00184609f $X=13.635 $Y=2.135 $X2=0
+ $Y2=0
cc_1064 N_A_2342_48#_c_1671_n N_A_c_1751_n 0.00117502f $X=13.65 $Y=1.97 $X2=0
+ $Y2=0
cc_1065 N_A_2342_48#_c_1667_n N_A_M1011_g 0.0116904f $X=13.475 $Y=1.215 $X2=0
+ $Y2=0
cc_1066 N_A_2342_48#_c_1668_n N_A_M1011_g 0.0126893f $X=13.64 $Y=0.515 $X2=0
+ $Y2=0
cc_1067 N_A_2342_48#_c_1671_n N_A_M1011_g 0.0158618f $X=13.65 $Y=1.97 $X2=0
+ $Y2=0
cc_1068 N_A_2342_48#_c_1672_n N_A_M1011_g 0.00438068f $X=13.652 $Y=1.215 $X2=0
+ $Y2=0
cc_1069 N_A_2342_48#_c_1667_n N_A_c_1748_n 0.048167f $X=13.475 $Y=1.215 $X2=0
+ $Y2=0
cc_1070 N_A_2342_48#_c_1669_n N_A_c_1748_n 0.00477495f $X=12.415 $Y=1.215 $X2=0
+ $Y2=0
cc_1071 N_A_2342_48#_c_1670_n N_A_c_1748_n 3.37225e-19 $X=12.415 $Y=1.385 $X2=0
+ $Y2=0
cc_1072 N_A_2342_48#_c_1678_n N_A_c_1748_n 0.00126392f $X=13.635 $Y=2.135 $X2=0
+ $Y2=0
cc_1073 N_A_2342_48#_c_1671_n N_A_c_1748_n 0.026181f $X=13.65 $Y=1.97 $X2=0
+ $Y2=0
cc_1074 N_A_2342_48#_c_1672_n N_A_c_1748_n 0.00119737f $X=13.652 $Y=1.215 $X2=0
+ $Y2=0
cc_1075 N_A_2342_48#_c_1667_n N_A_c_1749_n 0.00448411f $X=13.475 $Y=1.215 $X2=0
+ $Y2=0
cc_1076 N_A_2342_48#_c_1673_n N_VPWR_c_1815_n 0.00874897f $X=11.8 $Y=1.765 $X2=0
+ $Y2=0
cc_1077 N_A_2342_48#_c_1670_n N_VPWR_c_1815_n 6.8217e-19 $X=12.415 $Y=1.385
+ $X2=0 $Y2=0
cc_1078 N_A_2342_48#_c_1673_n N_VPWR_c_1816_n 0.0145305f $X=11.8 $Y=1.765 $X2=0
+ $Y2=0
cc_1079 N_A_2342_48#_c_1678_n N_VPWR_c_1817_n 0.0391256f $X=13.635 $Y=2.135
+ $X2=0 $Y2=0
cc_1080 N_A_2342_48#_c_1673_n N_VPWR_c_1818_n 0.00467264f $X=11.8 $Y=1.765 $X2=0
+ $Y2=0
cc_1081 N_A_2342_48#_c_1675_n N_VPWR_c_1823_n 0.0159324f $X=13.635 $Y=2.815
+ $X2=0 $Y2=0
cc_1082 N_A_2342_48#_c_1673_n N_VPWR_c_1812_n 0.0094358f $X=11.8 $Y=1.765 $X2=0
+ $Y2=0
cc_1083 N_A_2342_48#_c_1675_n N_VPWR_c_1812_n 0.0131546f $X=13.635 $Y=2.815
+ $X2=0 $Y2=0
cc_1084 N_A_2342_48#_c_1673_n N_A_1660_374#_c_2123_n 0.0042922f $X=11.8 $Y=1.765
+ $X2=0 $Y2=0
cc_1085 N_A_2342_48#_c_1665_n N_A_1660_374#_c_2117_n 0.00255579f $X=11.89
+ $Y=1.385 $X2=0 $Y2=0
cc_1086 N_A_2342_48#_c_1666_n N_A_1660_374#_c_2117_n 0.00210051f $X=11.8 $Y=1.22
+ $X2=0 $Y2=0
cc_1087 N_A_2342_48#_c_1673_n N_A_1660_374#_c_2118_n 0.0181236f $X=11.8 $Y=1.765
+ $X2=0 $Y2=0
cc_1088 N_A_2342_48#_c_1665_n N_A_1660_374#_c_2118_n 0.012419f $X=11.89 $Y=1.385
+ $X2=0 $Y2=0
cc_1089 N_A_2342_48#_c_1666_n N_A_1660_374#_c_2119_n 0.0156545f $X=11.8 $Y=1.22
+ $X2=0 $Y2=0
cc_1090 N_A_2342_48#_c_1665_n N_A_1849_374#_c_2209_n 0.00403444f $X=11.89
+ $Y=1.385 $X2=0 $Y2=0
cc_1091 N_A_2342_48#_c_1666_n N_A_1849_374#_c_2209_n 0.00529464f $X=11.8 $Y=1.22
+ $X2=0 $Y2=0
cc_1092 N_A_2342_48#_c_1669_n N_A_1849_374#_c_2209_n 0.0307016f $X=12.415
+ $Y=1.215 $X2=0 $Y2=0
cc_1093 N_A_2342_48#_c_1670_n N_A_1849_374#_c_2209_n 0.0213282f $X=12.415
+ $Y=1.385 $X2=0 $Y2=0
cc_1094 N_A_2342_48#_c_1667_n N_A_1849_374#_c_2210_n 0.0165889f $X=13.475
+ $Y=1.215 $X2=0 $Y2=0
cc_1095 N_A_2342_48#_c_1669_n N_A_1849_374#_c_2210_n 0.0273295f $X=12.415
+ $Y=1.215 $X2=0 $Y2=0
cc_1096 N_A_2342_48#_c_1670_n N_A_1849_374#_c_2210_n 0.00770779f $X=12.415
+ $Y=1.385 $X2=0 $Y2=0
cc_1097 N_A_2342_48#_c_1669_n N_A_1849_374#_c_2214_n 0.0103423f $X=12.415
+ $Y=1.215 $X2=0 $Y2=0
cc_1098 N_A_2342_48#_c_1670_n N_A_1849_374#_c_2214_n 0.00758313f $X=12.415
+ $Y=1.385 $X2=0 $Y2=0
cc_1099 N_A_2342_48#_c_1673_n N_A_1849_374#_c_2215_n 0.00370912f $X=11.8
+ $Y=1.765 $X2=0 $Y2=0
cc_1100 N_A_2342_48#_c_1665_n N_A_1849_374#_c_2215_n 0.00112223f $X=11.89
+ $Y=1.385 $X2=0 $Y2=0
cc_1101 N_A_2342_48#_c_1666_n N_A_1849_374#_c_2211_n 0.00437411f $X=11.8 $Y=1.22
+ $X2=0 $Y2=0
cc_1102 N_A_2342_48#_c_1673_n N_A_1849_374#_c_2216_n 0.00187811f $X=11.8
+ $Y=1.765 $X2=0 $Y2=0
cc_1103 N_A_2342_48#_c_1667_n N_A_1849_374#_c_2216_n 0.00750596f $X=13.475
+ $Y=1.215 $X2=0 $Y2=0
cc_1104 N_A_2342_48#_c_1669_n N_A_1849_374#_c_2216_n 0.0150945f $X=12.415
+ $Y=1.215 $X2=0 $Y2=0
cc_1105 N_A_2342_48#_c_1670_n N_A_1849_374#_c_2216_n 0.00145402f $X=12.415
+ $Y=1.385 $X2=0 $Y2=0
cc_1106 N_A_2342_48#_c_1673_n N_A_1849_374#_c_2218_n 0.0136581f $X=11.8 $Y=1.765
+ $X2=0 $Y2=0
cc_1107 N_A_2342_48#_c_1665_n N_A_1849_374#_c_2218_n 3.89416e-19 $X=11.89
+ $Y=1.385 $X2=0 $Y2=0
cc_1108 N_A_2342_48#_c_1670_n N_A_1849_374#_c_2218_n 4.29838e-19 $X=12.415
+ $Y=1.385 $X2=0 $Y2=0
cc_1109 N_A_2342_48#_c_1673_n N_A_1849_374#_c_2219_n 5.99895e-19 $X=11.8
+ $Y=1.765 $X2=0 $Y2=0
cc_1110 N_A_2342_48#_c_1669_n N_A_1849_374#_c_2219_n 9.70457e-19 $X=12.415
+ $Y=1.215 $X2=0 $Y2=0
cc_1111 N_A_2342_48#_c_1666_n N_VGND_c_2320_n 0.00982366f $X=11.8 $Y=1.22 $X2=0
+ $Y2=0
cc_1112 N_A_2342_48#_c_1670_n N_VGND_c_2320_n 7.81927e-19 $X=12.415 $Y=1.385
+ $X2=0 $Y2=0
cc_1113 N_A_2342_48#_c_1667_n N_VGND_c_2321_n 0.0243395f $X=13.475 $Y=1.215
+ $X2=0 $Y2=0
cc_1114 N_A_2342_48#_c_1668_n N_VGND_c_2321_n 0.0239364f $X=13.64 $Y=0.515 $X2=0
+ $Y2=0
cc_1115 N_A_2342_48#_c_1666_n N_VGND_c_2324_n 0.00428607f $X=11.8 $Y=1.22 $X2=0
+ $Y2=0
cc_1116 N_A_2342_48#_c_1668_n N_VGND_c_2329_n 0.0156794f $X=13.64 $Y=0.515 $X2=0
+ $Y2=0
cc_1117 N_A_2342_48#_c_1666_n N_VGND_c_2330_n 0.00811938f $X=11.8 $Y=1.22 $X2=0
+ $Y2=0
cc_1118 N_A_2342_48#_c_1668_n N_VGND_c_2330_n 0.0129217f $X=13.64 $Y=0.515 $X2=0
+ $Y2=0
cc_1119 N_A_c_1750_n N_VPWR_c_1816_n 0.00358265f $X=12.91 $Y=1.885 $X2=0 $Y2=0
cc_1120 N_A_c_1750_n N_VPWR_c_1817_n 0.0064431f $X=12.91 $Y=1.885 $X2=0 $Y2=0
cc_1121 N_A_c_1751_n N_VPWR_c_1817_n 0.0084134f $X=13.41 $Y=1.885 $X2=0 $Y2=0
cc_1122 N_A_c_1748_n N_VPWR_c_1817_n 0.0195375f $X=13.325 $Y=1.635 $X2=0 $Y2=0
cc_1123 N_A_c_1749_n N_VPWR_c_1817_n 0.00590265f $X=13.41 $Y=1.677 $X2=0 $Y2=0
cc_1124 N_A_c_1750_n N_VPWR_c_1822_n 0.00445602f $X=12.91 $Y=1.885 $X2=0 $Y2=0
cc_1125 N_A_c_1751_n N_VPWR_c_1823_n 0.00445602f $X=13.41 $Y=1.885 $X2=0 $Y2=0
cc_1126 N_A_c_1750_n N_VPWR_c_1812_n 0.00862852f $X=12.91 $Y=1.885 $X2=0 $Y2=0
cc_1127 N_A_c_1751_n N_VPWR_c_1812_n 0.00860889f $X=13.41 $Y=1.885 $X2=0 $Y2=0
cc_1128 N_A_M1014_g N_A_1849_374#_c_2211_n 4.67402e-19 $X=12.895 $Y=0.69 $X2=0
+ $Y2=0
cc_1129 N_A_c_1750_n N_A_1849_374#_c_2216_n 0.00496144f $X=12.91 $Y=1.885 $X2=0
+ $Y2=0
cc_1130 N_A_c_1748_n N_A_1849_374#_c_2216_n 0.00875643f $X=13.325 $Y=1.635 $X2=0
+ $Y2=0
cc_1131 N_A_c_1749_n N_A_1849_374#_c_2216_n 0.00422166f $X=13.41 $Y=1.677 $X2=0
+ $Y2=0
cc_1132 N_A_c_1750_n N_A_1849_374#_c_2217_n 0.00891175f $X=12.91 $Y=1.885 $X2=0
+ $Y2=0
cc_1133 N_A_c_1750_n N_A_1849_374#_c_2219_n 0.00110561f $X=12.91 $Y=1.885 $X2=0
+ $Y2=0
cc_1134 N_A_M1014_g N_VGND_c_2320_n 0.00306313f $X=12.895 $Y=0.69 $X2=0 $Y2=0
cc_1135 N_A_M1014_g N_VGND_c_2321_n 0.00349379f $X=12.895 $Y=0.69 $X2=0 $Y2=0
cc_1136 N_A_M1011_g N_VGND_c_2321_n 0.00660592f $X=13.425 $Y=0.69 $X2=0 $Y2=0
cc_1137 N_A_M1014_g N_VGND_c_2328_n 0.00461464f $X=12.895 $Y=0.69 $X2=0 $Y2=0
cc_1138 N_A_M1011_g N_VGND_c_2329_n 0.00434272f $X=13.425 $Y=0.69 $X2=0 $Y2=0
cc_1139 N_A_M1014_g N_VGND_c_2330_n 0.00913126f $X=12.895 $Y=0.69 $X2=0 $Y2=0
cc_1140 N_A_M1011_g N_VGND_c_2330_n 0.00824632f $X=13.425 $Y=0.69 $X2=0 $Y2=0
cc_1141 N_SUM_c_1794_n N_VPWR_c_1813_n 0.0450242f $X=0.275 $Y=0.705 $X2=0 $Y2=0
cc_1142 N_SUM_c_1794_n N_VPWR_c_1812_n 0.0122313f $X=0.275 $Y=0.705 $X2=0 $Y2=0
cc_1143 N_SUM_c_1794_n N_VPWR_c_1825_n 0.0148169f $X=0.275 $Y=0.705 $X2=0 $Y2=0
cc_1144 N_SUM_c_1794_n N_COUT_c_1944_n 0.0642415f $X=0.275 $Y=0.705 $X2=0 $Y2=0
cc_1145 N_SUM_c_1794_n N_COUT_c_1969_n 0.0115198f $X=0.275 $Y=0.705 $X2=0 $Y2=0
cc_1146 N_SUM_c_1794_n N_COUT_c_1956_n 0.00509141f $X=0.275 $Y=0.705 $X2=0 $Y2=0
cc_1147 N_SUM_c_1794_n N_COUT_c_1958_n 0.011089f $X=0.275 $Y=0.705 $X2=0 $Y2=0
cc_1148 N_SUM_c_1794_n N_VGND_c_2317_n 0.00155012f $X=0.275 $Y=0.705 $X2=0 $Y2=0
cc_1149 N_SUM_c_1794_n N_VGND_c_2326_n 0.00826171f $X=0.275 $Y=0.705 $X2=0 $Y2=0
cc_1150 N_SUM_c_1794_n N_VGND_c_2330_n 0.0106812f $X=0.275 $Y=0.705 $X2=0 $Y2=0
cc_1151 N_VPWR_c_1812_n N_COUT_M1015_s 0.00246676f $X=13.68 $Y=3.33 $X2=0 $Y2=0
cc_1152 N_VPWR_M1021_d N_COUT_c_1944_n 0.00418525f $X=0.58 $Y=1.84 $X2=0 $Y2=0
cc_1153 N_VPWR_M1021_d N_COUT_c_1956_n 0.00834514f $X=0.58 $Y=1.84 $X2=0 $Y2=0
cc_1154 N_VPWR_c_1813_n N_COUT_c_1956_n 0.0446382f $X=0.73 $Y=2.455 $X2=0 $Y2=0
cc_1155 N_VPWR_c_1813_n N_COUT_c_1948_n 0.0142842f $X=0.73 $Y=2.455 $X2=0 $Y2=0
cc_1156 N_VPWR_c_1820_n N_COUT_c_1948_n 0.0121867f $X=2.935 $Y=3.33 $X2=0 $Y2=0
cc_1157 N_VPWR_c_1812_n N_COUT_c_1948_n 0.00660921f $X=13.68 $Y=3.33 $X2=0 $Y2=0
cc_1158 N_VPWR_M1021_d N_COUT_c_1958_n 0.0198149f $X=0.58 $Y=1.84 $X2=0 $Y2=0
cc_1159 N_VPWR_c_1813_n N_COUT_c_1958_n 0.0120859f $X=0.73 $Y=2.455 $X2=0 $Y2=0
cc_1160 N_VPWR_c_1826_n N_COUT_c_1949_n 0.00666314f $X=3.11 $Y=3.05 $X2=0 $Y2=0
cc_1161 N_VPWR_c_1820_n N_COUT_c_1950_n 0.0958558f $X=2.935 $Y=3.33 $X2=0 $Y2=0
cc_1162 N_VPWR_c_1812_n N_COUT_c_1950_n 0.056056f $X=13.68 $Y=3.33 $X2=0 $Y2=0
cc_1163 N_VPWR_M1015_d N_A_644_104#_c_2026_n 0.00729118f $X=2.865 $Y=1.84 $X2=0
+ $Y2=0
cc_1164 N_VPWR_c_1816_n N_A_1660_374#_c_2123_n 0.0121002f $X=12.115 $Y=2.615
+ $X2=0 $Y2=0
cc_1165 N_VPWR_c_1818_n N_A_1660_374#_c_2123_n 0.202938f $X=11.95 $Y=3.33 $X2=0
+ $Y2=0
cc_1166 N_VPWR_c_1812_n N_A_1660_374#_c_2123_n 0.106699f $X=13.68 $Y=3.33 $X2=0
+ $Y2=0
cc_1167 N_VPWR_c_1814_n N_A_1660_374#_c_2124_n 0.0142216f $X=7.835 $Y=1.93 $X2=0
+ $Y2=0
cc_1168 N_VPWR_c_1818_n N_A_1660_374#_c_2124_n 0.0299631f $X=11.95 $Y=3.33 $X2=0
+ $Y2=0
cc_1169 N_VPWR_c_1812_n N_A_1660_374#_c_2124_n 0.0150586f $X=13.68 $Y=3.33 $X2=0
+ $Y2=0
cc_1170 N_VPWR_c_1815_n N_A_1660_374#_c_2118_n 0.0257822f $X=12.12 $Y=2.5 $X2=0
+ $Y2=0
cc_1171 N_VPWR_c_1816_n N_A_1660_374#_c_2118_n 0.0268621f $X=12.115 $Y=2.615
+ $X2=0 $Y2=0
cc_1172 N_VPWR_c_1814_n N_A_1660_374#_c_2121_n 0.0897195f $X=7.835 $Y=1.93 $X2=0
+ $Y2=0
cc_1173 N_VPWR_M1007_d N_A_1849_374#_c_2214_n 0.00301654f $X=11.875 $Y=1.84
+ $X2=0 $Y2=0
cc_1174 N_VPWR_c_1815_n N_A_1849_374#_c_2214_n 0.0106222f $X=12.12 $Y=2.5 $X2=0
+ $Y2=0
cc_1175 N_VPWR_M1007_d N_A_1849_374#_c_2215_n 0.0023405f $X=11.875 $Y=1.84 $X2=0
+ $Y2=0
cc_1176 N_VPWR_c_1815_n N_A_1849_374#_c_2215_n 0.00912309f $X=12.12 $Y=2.5 $X2=0
+ $Y2=0
cc_1177 N_VPWR_c_1815_n N_A_1849_374#_c_2216_n 0.00357964f $X=12.12 $Y=2.5 $X2=0
+ $Y2=0
cc_1178 N_VPWR_c_1817_n N_A_1849_374#_c_2216_n 0.0122221f $X=13.135 $Y=2.135
+ $X2=0 $Y2=0
cc_1179 N_VPWR_c_1815_n N_A_1849_374#_c_2217_n 0.0206571f $X=12.12 $Y=2.5 $X2=0
+ $Y2=0
cc_1180 N_VPWR_c_1816_n N_A_1849_374#_c_2217_n 0.0324006f $X=12.115 $Y=2.615
+ $X2=0 $Y2=0
cc_1181 N_VPWR_c_1817_n N_A_1849_374#_c_2217_n 0.0549785f $X=13.135 $Y=2.135
+ $X2=0 $Y2=0
cc_1182 N_VPWR_c_1822_n N_A_1849_374#_c_2217_n 0.0145938f $X=13.05 $Y=3.33 $X2=0
+ $Y2=0
cc_1183 N_VPWR_c_1812_n N_A_1849_374#_c_2217_n 0.0120466f $X=13.68 $Y=3.33 $X2=0
+ $Y2=0
cc_1184 N_VPWR_M1007_d N_A_1849_374#_c_2218_n 0.00936693f $X=11.875 $Y=1.84
+ $X2=0 $Y2=0
cc_1185 N_VPWR_c_1815_n N_A_1849_374#_c_2218_n 0.0105734f $X=12.12 $Y=2.5 $X2=0
+ $Y2=0
cc_1186 N_VPWR_c_1815_n N_A_1849_374#_c_2219_n 0.00117549f $X=12.12 $Y=2.5 $X2=0
+ $Y2=0
cc_1187 N_VPWR_c_1817_n N_A_1849_374#_c_2219_n 9.00695e-19 $X=13.135 $Y=2.135
+ $X2=0 $Y2=0
cc_1188 N_COUT_c_1944_n N_VGND_M1029_d 0.0118219f $X=0.75 $Y=1.95 $X2=-0.19
+ $Y2=-0.245
cc_1189 N_COUT_c_1945_n N_VGND_M1029_d 0.00529767f $X=1.505 $Y=0.815 $X2=-0.19
+ $Y2=-0.245
cc_1190 N_COUT_c_1969_n N_VGND_M1029_d 0.00473001f $X=0.835 $Y=0.815 $X2=-0.19
+ $Y2=-0.245
cc_1191 N_COUT_c_1945_n N_VGND_c_2317_n 0.00889464f $X=1.505 $Y=0.815 $X2=0
+ $Y2=0
cc_1192 N_COUT_c_1969_n N_VGND_c_2317_n 0.0147103f $X=0.835 $Y=0.815 $X2=0 $Y2=0
cc_1193 COUT N_VGND_c_2317_n 0.0061156f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_1194 COUT N_VGND_c_2318_n 0.0136121f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_1195 N_COUT_c_1945_n N_VGND_c_2322_n 0.00704012f $X=1.505 $Y=0.815 $X2=0
+ $Y2=0
cc_1196 COUT N_VGND_c_2322_n 0.0198339f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_1197 N_COUT_c_1945_n N_VGND_c_2330_n 0.0128744f $X=1.505 $Y=0.815 $X2=0 $Y2=0
cc_1198 N_COUT_c_1969_n N_VGND_c_2330_n 7.33912e-19 $X=0.835 $Y=0.815 $X2=0
+ $Y2=0
cc_1199 COUT N_VGND_c_2330_n 0.0190337f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_1200 N_A_1660_374#_c_2119_n N_A_1849_374#_c_2209_n 0.05031f $X=11.57 $Y=0.515
+ $X2=0 $Y2=0
cc_1201 N_A_1660_374#_c_2118_n N_A_1849_374#_c_2215_n 0.0138969f $X=11.545
+ $Y=1.99 $X2=0 $Y2=0
cc_1202 N_A_1660_374#_c_2118_n N_A_1849_374#_c_2216_n 0.00232959f $X=11.545
+ $Y=1.99 $X2=0 $Y2=0
cc_1203 N_A_1660_374#_M1016_d N_A_1849_374#_c_2218_n 7.0241e-19 $X=11.37 $Y=1.84
+ $X2=0 $Y2=0
cc_1204 N_A_1660_374#_c_2118_n N_A_1849_374#_c_2218_n 0.0479486f $X=11.545
+ $Y=1.99 $X2=0 $Y2=0
cc_1205 N_A_1660_374#_c_2119_n N_VGND_c_2320_n 0.0106954f $X=11.57 $Y=0.515
+ $X2=0 $Y2=0
cc_1206 N_A_1660_374#_c_2119_n N_VGND_c_2324_n 0.0147721f $X=11.57 $Y=0.515
+ $X2=0 $Y2=0
cc_1207 N_A_1660_374#_c_2119_n N_VGND_c_2330_n 0.0121589f $X=11.57 $Y=0.515
+ $X2=0 $Y2=0
cc_1208 N_A_1849_374#_c_2209_n N_VGND_M1025_d 0.00638481f $X=11.995 $Y=1.72
+ $X2=0 $Y2=0
cc_1209 N_A_1849_374#_c_2210_n N_VGND_M1025_d 0.00463151f $X=12.475 $Y=0.875
+ $X2=0 $Y2=0
cc_1210 N_A_1849_374#_c_2308_p N_VGND_M1025_d 0.00328667f $X=12.08 $Y=0.875
+ $X2=0 $Y2=0
cc_1211 N_A_1849_374#_c_2210_n N_VGND_c_2320_n 0.0130525f $X=12.475 $Y=0.875
+ $X2=0 $Y2=0
cc_1212 N_A_1849_374#_c_2308_p N_VGND_c_2320_n 0.0143076f $X=12.08 $Y=0.875
+ $X2=0 $Y2=0
cc_1213 N_A_1849_374#_c_2211_n N_VGND_c_2320_n 0.0182033f $X=12.64 $Y=0.515
+ $X2=0 $Y2=0
cc_1214 N_A_1849_374#_c_2211_n N_VGND_c_2321_n 0.00158095f $X=12.64 $Y=0.515
+ $X2=0 $Y2=0
cc_1215 N_A_1849_374#_c_2211_n N_VGND_c_2328_n 0.0145203f $X=12.64 $Y=0.515
+ $X2=0 $Y2=0
cc_1216 N_A_1849_374#_c_2210_n N_VGND_c_2330_n 0.00889179f $X=12.475 $Y=0.875
+ $X2=0 $Y2=0
cc_1217 N_A_1849_374#_c_2308_p N_VGND_c_2330_n 8.90974e-19 $X=12.08 $Y=0.875
+ $X2=0 $Y2=0
cc_1218 N_A_1849_374#_c_2211_n N_VGND_c_2330_n 0.0120696f $X=12.64 $Y=0.515
+ $X2=0 $Y2=0
