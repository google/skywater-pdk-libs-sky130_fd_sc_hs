* File: sky130_fd_sc_hs__nand2b_1.spice
* Created: Tue Sep  1 20:08:54 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hs__nand2b_1.pex.spice"
.subckt sky130_fd_sc_hs__nand2b_1  VNB VPB A_N B VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* B	B
* A_N	A_N
* VPB	VPB
* VNB	VNB
MM1004 N_VGND_M1004_d N_A_N_M1004_g N_A_27_112#_M1004_s VNB NLOWVT L=0.15 W=0.55
+ AD=0.191114 AS=0.15675 PD=1.16395 PS=1.67 NRD=1.08 NRS=0 M=1 R=3.66667
+ SA=75000.2 SB=75001.5 A=0.0825 P=1.4 MULT=1
MM1001 A_269_74# N_B_M1001_g N_VGND_M1004_d VNB NLOWVT L=0.15 W=0.74 AD=0.0888
+ AS=0.257136 PD=0.98 PS=1.56605 NRD=10.536 NRS=0 M=1 R=4.93333 SA=75000.9
+ SB=75000.7 A=0.111 P=1.78 MULT=1
MM1000 N_Y_M1000_d N_A_27_112#_M1000_g A_269_74# VNB NLOWVT L=0.15 W=0.74
+ AD=0.3182 AS=0.0888 PD=2.34 PS=0.98 NRD=10.536 NRS=10.536 M=1 R=4.93333
+ SA=75001.2 SB=75000.4 A=0.111 P=1.78 MULT=1
MM1005 N_VPWR_M1005_d N_A_N_M1005_g N_A_27_112#_M1005_s VPB PSHORT L=0.15 W=0.84
+ AD=0.2388 AS=0.2478 PD=1.40571 PS=2.27 NRD=23.443 NRS=2.3443 M=1 R=5.6
+ SA=75000.2 SB=75001.4 A=0.126 P=1.98 MULT=1
MM1003 N_Y_M1003_d N_B_M1003_g N_VPWR_M1005_d VPB PSHORT L=0.15 W=1.12 AD=0.196
+ AS=0.3184 PD=1.47 PS=1.87429 NRD=1.7533 NRS=24.625 M=1 R=7.46667 SA=75000.8
+ SB=75000.7 A=0.168 P=2.54 MULT=1
MM1002 N_VPWR_M1002_d N_A_27_112#_M1002_g N_Y_M1003_d VPB PSHORT L=0.15 W=1.12
+ AD=0.336 AS=0.196 PD=2.84 PS=1.47 NRD=1.7533 NRS=10.5395 M=1 R=7.46667
+ SA=75001.3 SB=75000.2 A=0.168 P=2.54 MULT=1
DX6_noxref VNB VPB NWDIODE A=5.1708 P=9.28
c_23 VNB 0 1.74227e-19 $X=0 $Y=0
*
.include "sky130_fd_sc_hs__nand2b_1.pxi.spice"
*
.ends
*
*
