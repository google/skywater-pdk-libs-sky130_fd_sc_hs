# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_hs__a21bo_4
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_hs__a21bo_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  6.240000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.445000 1.450000 5.200000 1.780000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.935000 0.255000 4.265000 0.670000 ;
    END
  END A2
  PIN B1_N
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 0.255000 0.625000 0.505000 ;
        RECT 0.125000 0.505000 0.355000 0.670000 ;
    END
  END B1_N
  PIN X
    ANTENNADIFFAREA  1.086400 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605000 1.510000 1.420000 1.850000 ;
        RECT 0.605000 1.850000 2.300000 2.100000 ;
        RECT 1.250000 0.480000 1.555000 1.010000 ;
        RECT 1.250000 1.010000 2.415000 1.180000 ;
        RECT 1.250000 1.180000 1.420000 1.510000 ;
        RECT 2.165000 0.480000 2.415000 1.010000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 6.240000 0.085000 ;
        RECT 0.795000  0.085000 1.045000 1.275000 ;
        RECT 1.735000  0.085000 1.985000 0.840000 ;
        RECT 2.595000  0.085000 2.845000 0.940000 ;
        RECT 3.595000  0.085000 3.765000 0.940000 ;
        RECT 5.725000  0.085000 5.975000 1.275000 ;
      LAYER mcon ;
        RECT 0.155000 -0.085000 0.325000 0.085000 ;
        RECT 0.635000 -0.085000 0.805000 0.085000 ;
        RECT 1.115000 -0.085000 1.285000 0.085000 ;
        RECT 1.595000 -0.085000 1.765000 0.085000 ;
        RECT 2.075000 -0.085000 2.245000 0.085000 ;
        RECT 2.555000 -0.085000 2.725000 0.085000 ;
        RECT 3.035000 -0.085000 3.205000 0.085000 ;
        RECT 3.515000 -0.085000 3.685000 0.085000 ;
        RECT 3.995000 -0.085000 4.165000 0.085000 ;
        RECT 4.475000 -0.085000 4.645000 0.085000 ;
        RECT 4.955000 -0.085000 5.125000 0.085000 ;
        RECT 5.435000 -0.085000 5.605000 0.085000 ;
        RECT 5.915000 -0.085000 6.085000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.245000 6.240000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 3.245000 6.240000 3.415000 ;
        RECT 0.620000 2.610000 0.950000 3.245000 ;
        RECT 1.520000 2.610000 1.850000 3.245000 ;
        RECT 2.420000 2.610000 2.750000 3.245000 ;
        RECT 4.290000 2.290000 4.540000 3.245000 ;
        RECT 5.270000 2.290000 5.520000 3.245000 ;
      LAYER mcon ;
        RECT 0.155000 3.245000 0.325000 3.415000 ;
        RECT 0.635000 3.245000 0.805000 3.415000 ;
        RECT 1.115000 3.245000 1.285000 3.415000 ;
        RECT 1.595000 3.245000 1.765000 3.415000 ;
        RECT 2.075000 3.245000 2.245000 3.415000 ;
        RECT 2.555000 3.245000 2.725000 3.415000 ;
        RECT 3.035000 3.245000 3.205000 3.415000 ;
        RECT 3.515000 3.245000 3.685000 3.415000 ;
        RECT 3.995000 3.245000 4.165000 3.415000 ;
        RECT 4.475000 3.245000 4.645000 3.415000 ;
        RECT 4.955000 3.245000 5.125000 3.415000 ;
        RECT 5.435000 3.245000 5.605000 3.415000 ;
        RECT 5.915000 3.245000 6.085000 3.415000 ;
      LAYER met1 ;
        RECT 0.000000 3.085000 6.240000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.105000 0.840000 0.615000 1.275000 ;
      RECT 0.105000 1.275000 0.435000 2.270000 ;
      RECT 0.105000 2.270000 2.640000 2.440000 ;
      RECT 0.105000 2.440000 0.435000 2.980000 ;
      RECT 1.590000 1.350000 2.755000 1.680000 ;
      RECT 2.470000 1.850000 3.290000 2.020000 ;
      RECT 2.470000 2.020000 2.640000 2.270000 ;
      RECT 2.585000 1.110000 5.035000 1.280000 ;
      RECT 2.585000 1.280000 2.755000 1.350000 ;
      RECT 2.940000 2.190000 3.270000 2.905000 ;
      RECT 2.940000 2.905000 4.090000 3.075000 ;
      RECT 2.960000 1.450000 3.290000 1.850000 ;
      RECT 3.085000 0.595000 3.415000 1.110000 ;
      RECT 3.470000 1.280000 3.720000 2.735000 ;
      RECT 3.920000 1.940000 4.090000 1.950000 ;
      RECT 3.920000 1.950000 5.970000 2.120000 ;
      RECT 3.920000 2.120000 4.090000 2.905000 ;
      RECT 4.435000 0.255000 5.545000 0.425000 ;
      RECT 4.435000 0.425000 4.605000 0.940000 ;
      RECT 4.740000 2.120000 5.070000 2.980000 ;
      RECT 4.785000 0.595000 5.035000 1.110000 ;
      RECT 5.215000 0.425000 5.545000 1.275000 ;
      RECT 5.720000 1.940000 5.970000 1.950000 ;
      RECT 5.720000 2.120000 5.970000 2.980000 ;
  END
END sky130_fd_sc_hs__a21bo_4
