* File: sky130_fd_sc_hs__a21oi_2.spice
* Created: Thu Aug 27 20:25:18 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hs__a21oi_2.pex.spice"
.subckt sky130_fd_sc_hs__a21oi_2  VNB VPB B1 A2 A1 Y VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* Y	Y
* A1	A1
* A2	A2
* B1	B1
* VPB	VPB
* VNB	VNB
MM1010 N_Y_M1010_d N_B1_M1010_g N_VGND_M1010_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1961 AS=0.1961 PD=2.01 PS=2.01 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1002 N_A_280_107#_M1002_d N_A2_M1002_g N_VGND_M1002_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.25175 AS=0.193662 PD=2.22 PS=1.405 NRD=0.396 NRS=33.516 M=1 R=4.93333
+ SA=75000.2 SB=75001.4 A=0.111 P=1.78 MULT=1
MM1004 N_A_280_107#_M1004_d N_A2_M1004_g N_VGND_M1002_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.193662 PD=1.02 PS=1.405 NRD=0 NRS=11.34 M=1 R=4.93333
+ SA=75000.8 SB=75001.1 A=0.111 P=1.78 MULT=1
MM1000 N_A_280_107#_M1004_d N_A1_M1000_g N_Y_M1000_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.2
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1006 N_A_280_107#_M1006_d N_A1_M1006_g N_Y_M1000_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1961 AS=0.1036 PD=2.01 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.6
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1007 N_Y_M1007_d N_B1_M1007_g N_A_131_368#_M1007_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.308 PD=1.42 PS=2.79 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75002.5 A=0.168 P=2.54 MULT=1
MM1008 N_Y_M1007_d N_B1_M1008_g N_A_131_368#_M1008_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.6 SB=75002.1 A=0.168 P=2.54 MULT=1
MM1001 N_A_131_368#_M1008_s N_A2_M1001_g N_VPWR_M1001_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.2016 PD=1.42 PS=1.48 NRD=1.7533 NRS=2.6201 M=1 R=7.46667
+ SA=75001.1 SB=75001.6 A=0.168 P=2.54 MULT=1
MM1009 N_A_131_368#_M1009_d N_A2_M1009_g N_VPWR_M1001_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.2016 PD=1.42 PS=1.48 NRD=1.7533 NRS=11.426 M=1 R=7.46667
+ SA=75001.6 SB=75001.1 A=0.168 P=2.54 MULT=1
MM1003 N_VPWR_M1003_d N_A1_M1003_g N_A_131_368#_M1009_d VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75002.1 SB=75000.6 A=0.168 P=2.54 MULT=1
MM1005 N_VPWR_M1003_d N_A1_M1005_g N_A_131_368#_M1005_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.308 PD=1.42 PS=2.79 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75002.5 SB=75000.2 A=0.168 P=2.54 MULT=1
DX11_noxref VNB VPB NWDIODE A=7.8492 P=12.16
*
.include "sky130_fd_sc_hs__a21oi_2.pxi.spice"
*
.ends
*
*
