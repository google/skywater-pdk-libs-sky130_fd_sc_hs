* NGSPICE file created from sky130_fd_sc_hs__o2bb2ai_2.ext - technology: sky130A

.subckt sky130_fd_sc_hs__o2bb2ai_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
M1000 Y a_133_387# a_518_74# VNB nlowvt w=740000u l=150000u
+  ad=2.072e+11p pd=2.04e+06u as=8.954e+11p ps=8.34e+06u
M1001 VPWR a_133_387# Y VPB pshort w=1.12e+06u l=150000u
+  ad=2.15495e+12p pd=1.515e+07u as=6.888e+11p ps=5.71e+06u
M1002 VGND B2 a_518_74# VNB nlowvt w=740000u l=150000u
+  ad=8.869e+11p pd=8.09e+06u as=0p ps=0u
M1003 a_133_387# A2_N VPWR VPB pshort w=840000u l=150000u
+  ad=5.96625e+11p pd=4.94e+06u as=0p ps=0u
M1004 a_133_387# A1_N VPWR VPB pshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_518_74# a_133_387# Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_134_74# A1_N VGND VNB nlowvt w=640000u l=150000u
+  ad=3.584e+11p pd=3.68e+06u as=0p ps=0u
M1007 a_133_387# A2_N a_134_74# VNB nlowvt w=640000u l=150000u
+  ad=2.272e+11p pd=1.99e+06u as=0p ps=0u
M1008 a_518_74# B1 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VPWR A2_N a_133_387# VPB pshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_796_368# B1 VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=6.72e+11p pd=5.68e+06u as=0p ps=0u
M1011 Y B2 a_796_368# VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VGND A1_N a_134_74# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_796_368# B2 Y VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 Y a_133_387# VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_518_74# B2 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VGND B1 a_518_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 VPWR B1 a_796_368# VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 VPWR A1_N a_133_387# VPB pshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_134_74# A2_N a_133_387# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

