* File: sky130_fd_sc_hs__a311oi_2.spice
* Created: Tue Sep  1 19:52:38 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hs__a311oi_2.pex.spice"
.subckt sky130_fd_sc_hs__a311oi_2  VNB VPB A3 A2 A1 B1 C1 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* C1	C1
* B1	B1
* A1	A1
* A2	A2
* A3	A3
* VPB	VPB
* VNB	VNB
MM1008 N_A_45_74#_M1008_d N_A3_M1008_g N_VGND_M1008_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1961 AS=0.1036 PD=2.01 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75001.5 A=0.111 P=1.78 MULT=1
MM1009 N_A_45_74#_M1009_d N_A3_M1009_g N_VGND_M1008_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.6
+ SB=75001.1 A=0.111 P=1.78 MULT=1
MM1006 N_A_45_74#_M1009_d N_A2_M1006_g N_A_300_74#_M1006_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75001.1 SB=75000.6 A=0.111 P=1.78 MULT=1
MM1014 N_A_45_74#_M1014_d N_A2_M1014_g N_A_300_74#_M1006_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1961 AS=0.1036 PD=2.01 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75001.5 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1011 N_Y_M1011_d N_A1_M1011_g N_A_300_74#_M1011_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1961 AS=0.1036 PD=2.01 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75001.9 A=0.111 P=1.78 MULT=1
MM1017 N_Y_M1017_d N_A1_M1017_g N_A_300_74#_M1011_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.6
+ SB=75001.5 A=0.111 P=1.78 MULT=1
MM1015 N_VGND_M1015_d N_B1_M1015_g N_Y_M1017_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.2553 AS=0.1036 PD=1.43 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.1
+ SB=75001 A=0.111 P=1.78 MULT=1
MM1000 N_Y_M1000_d N_C1_M1000_g N_VGND_M1015_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.1961 AS=0.2553 PD=2.01 PS=1.43 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.9
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1001 N_A_127_368#_M1001_d N_A3_M1001_g N_VPWR_M1001_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.308 PD=1.42 PS=2.79 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75002.5 A=0.168 P=2.54 MULT=1
MM1002 N_A_127_368#_M1001_d N_A3_M1002_g N_VPWR_M1002_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.6 SB=75002 A=0.168 P=2.54 MULT=1
MM1003 N_A_127_368#_M1003_d N_A2_M1003_g N_VPWR_M1002_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.1 SB=75001.6 A=0.168 P=2.54 MULT=1
MM1005 N_A_127_368#_M1003_d N_A2_M1005_g N_VPWR_M1005_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.1848 PD=1.42 PS=1.45 NRD=1.7533 NRS=4.3931 M=1 R=7.46667
+ SA=75001.5 SB=75001.1 A=0.168 P=2.54 MULT=1
MM1004 N_A_127_368#_M1004_d N_A1_M1004_g N_VPWR_M1005_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.1848 PD=1.42 PS=1.45 NRD=1.7533 NRS=4.3931 M=1 R=7.46667
+ SA=75002 SB=75000.6 A=0.168 P=2.54 MULT=1
MM1007 N_A_127_368#_M1004_d N_A1_M1007_g N_VPWR_M1007_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.308 PD=1.42 PS=2.79 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75002.5 SB=75000.2 A=0.168 P=2.54 MULT=1
MM1010 N_A_127_368#_M1010_d N_B1_M1010_g N_A_692_368#_M1010_s VPB PSHORT L=0.15
+ W=1.12 AD=0.168 AS=0.308 PD=1.42 PS=2.79 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75001.5 A=0.168 P=2.54 MULT=1
MM1012 N_A_127_368#_M1010_d N_B1_M1012_g N_A_692_368#_M1012_s VPB PSHORT L=0.15
+ W=1.12 AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.6 SB=75001.1 A=0.168 P=2.54 MULT=1
MM1013 N_Y_M1013_d N_C1_M1013_g N_A_692_368#_M1012_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.1 SB=75000.6 A=0.168 P=2.54 MULT=1
MM1016 N_Y_M1013_d N_C1_M1016_g N_A_692_368#_M1016_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.308 PD=1.42 PS=2.79 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.5 SB=75000.2 A=0.168 P=2.54 MULT=1
DX18_noxref VNB VPB NWDIODE A=11.4204 P=16
*
.include "sky130_fd_sc_hs__a311oi_2.pxi.spice"
*
.ends
*
*
