* File: sky130_fd_sc_hs__o211ai_2.spice
* Created: Thu Aug 27 20:57:17 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hs__o211ai_2.pex.spice"
.subckt sky130_fd_sc_hs__o211ai_2  VNB VPB C1 B1 A2 A1 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A1	A1
* A2	A2
* B1	B1
* C1	C1
* VPB	VPB
* VNB	VNB
MM1003 N_A_30_84#_M1003_d N_C1_M1003_g N_Y_M1003_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.1036 PD=2.05 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75001.6 A=0.111 P=1.78 MULT=1
MM1004 N_A_30_84#_M1004_d N_C1_M1004_g N_Y_M1003_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1295 AS=0.1036 PD=1.09 PS=1.02 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75000.6
+ SB=75001.2 A=0.111 P=1.78 MULT=1
MM1001 N_A_303_84#_M1001_d N_B1_M1001_g N_A_30_84#_M1004_d VNB NLOWVT L=0.15
+ W=0.74 AD=0.1295 AS=0.1295 PD=1.09 PS=1.09 NRD=11.34 NRS=0 M=1 R=4.93333
+ SA=75001.1 SB=75000.7 A=0.111 P=1.78 MULT=1
MM1015 N_A_303_84#_M1001_d N_B1_M1015_g N_A_30_84#_M1015_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1295 AS=0.2183 PD=1.09 PS=2.07 NRD=0 NRS=0.804 M=1 R=4.93333
+ SA=75001.6 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1007 N_VGND_M1007_d N_A2_M1007_g N_A_303_84#_M1007_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.1036 PD=2.05 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75001.6 A=0.111 P=1.78 MULT=1
MM1013 N_VGND_M1013_d N_A2_M1013_g N_A_303_84#_M1007_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.10545 AS=0.1036 PD=1.025 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.6
+ SB=75001.1 A=0.111 P=1.78 MULT=1
MM1008 N_A_303_84#_M1008_d N_A1_M1008_g N_VGND_M1013_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.12025 AS=0.10545 PD=1.065 PS=1.025 NRD=0 NRS=0.804 M=1 R=4.93333
+ SA=75001.1 SB=75000.7 A=0.111 P=1.78 MULT=1
MM1014 N_A_303_84#_M1008_d N_A1_M1014_g N_VGND_M1014_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.12025 AS=0.2294 PD=1.065 PS=2.1 NRD=7.296 NRS=0 M=1 R=4.93333 SA=75001.6
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1009 N_VPWR_M1009_d N_C1_M1009_g N_Y_M1009_s VPB PSHORT L=0.15 W=1.12
+ AD=0.3304 AS=0.168 PD=2.83 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75001.6 A=0.168 P=2.54 MULT=1
MM1010 N_VPWR_M1010_d N_C1_M1010_g N_Y_M1009_s VPB PSHORT L=0.15 W=1.12 AD=0.168
+ AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667 SA=75000.7
+ SB=75001.1 A=0.168 P=2.54 MULT=1
MM1011 N_Y_M1011_d N_B1_M1011_g N_VPWR_M1010_d VPB PSHORT L=0.15 W=1.12 AD=0.168
+ AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667 SA=75001.1
+ SB=75000.7 A=0.168 P=2.54 MULT=1
MM1012 N_Y_M1011_d N_B1_M1012_g N_VPWR_M1012_s VPB PSHORT L=0.15 W=1.12 AD=0.168
+ AS=0.3304 PD=1.42 PS=2.83 NRD=1.7533 NRS=1.7533 M=1 R=7.46667 SA=75001.6
+ SB=75000.2 A=0.168 P=2.54 MULT=1
MM1000 N_Y_M1000_d N_A2_M1000_g N_A_505_368#_M1000_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.3304 PD=1.42 PS=2.83 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75001.6 A=0.168 P=2.54 MULT=1
MM1002 N_Y_M1000_d N_A2_M1002_g N_A_505_368#_M1002_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.7 SB=75001.2 A=0.168 P=2.54 MULT=1
MM1005 N_VPWR_M1005_d N_A1_M1005_g N_A_505_368#_M1002_s VPB PSHORT L=0.15 W=1.12
+ AD=0.196 AS=0.168 PD=1.47 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.1 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1006 N_VPWR_M1005_d N_A1_M1006_g N_A_505_368#_M1006_s VPB PSHORT L=0.15 W=1.12
+ AD=0.196 AS=0.3304 PD=1.47 PS=2.83 NRD=10.5395 NRS=1.7533 M=1 R=7.46667
+ SA=75001.6 SB=75000.2 A=0.168 P=2.54 MULT=1
DX16_noxref VNB VPB NWDIODE A=9.6348 P=14.08
*
.include "sky130_fd_sc_hs__o211ai_2.pxi.spice"
*
.ends
*
*
