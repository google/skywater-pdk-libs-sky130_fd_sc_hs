* File: sky130_fd_sc_hs__o32ai_1.pxi.spice
* Created: Tue Sep  1 20:18:51 2020
* 
x_PM_SKY130_FD_SC_HS__O32AI_1%B1 N_B1_c_48_n N_B1_M1008_g N_B1_c_49_n
+ N_B1_M1000_g B1 PM_SKY130_FD_SC_HS__O32AI_1%B1
x_PM_SKY130_FD_SC_HS__O32AI_1%B2 N_B2_c_71_n N_B2_M1005_g N_B2_M1006_g B2
+ N_B2_c_73_n PM_SKY130_FD_SC_HS__O32AI_1%B2
x_PM_SKY130_FD_SC_HS__O32AI_1%A3 N_A3_c_98_n N_A3_M1001_g N_A3_M1003_g A3 A3 A3
+ N_A3_c_100_n PM_SKY130_FD_SC_HS__O32AI_1%A3
x_PM_SKY130_FD_SC_HS__O32AI_1%A2 N_A2_c_130_n N_A2_M1009_g N_A2_M1007_g A2 A2 A2
+ A2 N_A2_c_132_n PM_SKY130_FD_SC_HS__O32AI_1%A2
x_PM_SKY130_FD_SC_HS__O32AI_1%A1 N_A1_c_163_n N_A1_M1004_g N_A1_c_164_n
+ N_A1_M1002_g A1 PM_SKY130_FD_SC_HS__O32AI_1%A1
x_PM_SKY130_FD_SC_HS__O32AI_1%VPWR N_VPWR_M1000_s N_VPWR_M1002_d N_VPWR_c_185_n
+ N_VPWR_c_186_n N_VPWR_c_187_n N_VPWR_c_188_n VPWR N_VPWR_c_189_n
+ N_VPWR_c_184_n PM_SKY130_FD_SC_HS__O32AI_1%VPWR
x_PM_SKY130_FD_SC_HS__O32AI_1%Y N_Y_M1008_d N_Y_M1005_d N_Y_c_215_n Y
+ N_Y_c_217_n N_Y_c_216_n PM_SKY130_FD_SC_HS__O32AI_1%Y
x_PM_SKY130_FD_SC_HS__O32AI_1%A_27_74# N_A_27_74#_M1008_s N_A_27_74#_M1006_d
+ N_A_27_74#_M1007_d N_A_27_74#_c_247_n N_A_27_74#_c_248_n N_A_27_74#_c_260_n
+ N_A_27_74#_c_249_n N_A_27_74#_c_250_n N_A_27_74#_c_251_n N_A_27_74#_c_252_n
+ PM_SKY130_FD_SC_HS__O32AI_1%A_27_74#
x_PM_SKY130_FD_SC_HS__O32AI_1%VGND N_VGND_M1003_d N_VGND_M1004_d N_VGND_c_292_n
+ N_VGND_c_293_n N_VGND_c_294_n N_VGND_c_295_n N_VGND_c_296_n VGND
+ N_VGND_c_297_n N_VGND_c_298_n PM_SKY130_FD_SC_HS__O32AI_1%VGND
cc_1 VNB N_B1_c_48_n 0.0254704f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.22
cc_2 VNB N_B1_c_49_n 0.0726862f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=1.765
cc_3 VNB B1 0.0084694f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_4 VNB N_B2_c_71_n 0.0300525f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.22
cc_5 VNB N_B2_M1006_g 0.0290226f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=2.4
cc_6 VNB N_B2_c_73_n 0.00473922f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=1.295
cc_7 VNB N_A3_c_98_n 0.0269882f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.22
cc_8 VNB N_A3_M1003_g 0.0270536f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=2.4
cc_9 VNB N_A3_c_100_n 0.00166948f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A2_c_130_n 0.0251332f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.22
cc_11 VNB N_A2_M1007_g 0.0260977f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=2.4
cc_12 VNB N_A2_c_132_n 0.00421825f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A1_c_163_n 0.0198499f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.22
cc_14 VNB N_A1_c_164_n 0.0649949f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=1.765
cc_15 VNB A1 0.0260696f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_16 VNB N_VPWR_c_184_n 0.143779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_Y_c_215_n 0.00685991f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=1.295
cc_18 VNB N_Y_c_216_n 0.00701282f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_27_74#_c_247_n 0.005426f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=1.295
cc_20 VNB N_A_27_74#_c_248_n 0.00261637f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_27_74#_c_249_n 0.018049f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_27_74#_c_250_n 0.00949292f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_27_74#_c_251_n 0.00240191f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_27_74#_c_252_n 0.0284201f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_VGND_c_292_n 0.00977355f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.385
cc_26 VNB N_VGND_c_293_n 0.0142197f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=1.385
cc_27 VNB N_VGND_c_294_n 0.0361072f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_295_n 0.0488022f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_296_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_297_n 0.0196495f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_298_n 0.211748f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VPB N_B1_c_49_n 0.0268816f $X=-0.19 $Y=1.66 $X2=0.565 $Y2=1.765
cc_33 VPB N_B2_c_71_n 0.0307041f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.22
cc_34 VPB N_B2_c_73_n 0.00319058f $X=-0.19 $Y=1.66 $X2=0.28 $Y2=1.295
cc_35 VPB N_A3_c_98_n 0.0293603f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.22
cc_36 VPB N_A3_c_100_n 0.00193983f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_37 VPB N_A2_c_130_n 0.0281441f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.22
cc_38 VPB N_A2_c_132_n 0.00293465f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_39 VPB N_A1_c_164_n 0.030391f $X=-0.19 $Y=1.66 $X2=0.565 $Y2=1.765
cc_40 VPB N_VPWR_c_185_n 0.0128289f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.21
cc_41 VPB N_VPWR_c_186_n 0.0594635f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.385
cc_42 VPB N_VPWR_c_187_n 0.0145625f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_43 VPB N_VPWR_c_188_n 0.0559582f $X=-0.19 $Y=1.66 $X2=0.28 $Y2=1.385
cc_44 VPB N_VPWR_c_189_n 0.0668059f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_45 VPB N_VPWR_c_184_n 0.0832039f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_46 VPB N_Y_c_217_n 0.00533878f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_47 VPB N_Y_c_216_n 0.00125525f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_48 N_B1_c_49_n N_B2_c_71_n 0.0822961f $X=0.565 $Y=1.765 $X2=-0.19 $Y2=-0.245
cc_49 N_B1_c_48_n N_B2_M1006_g 0.0177514f $X=0.495 $Y=1.22 $X2=0 $Y2=0
cc_50 N_B1_c_49_n N_B2_c_73_n 3.24204e-19 $X=0.565 $Y=1.765 $X2=0 $Y2=0
cc_51 N_B1_c_49_n N_VPWR_c_186_n 0.00983179f $X=0.565 $Y=1.765 $X2=0 $Y2=0
cc_52 B1 N_VPWR_c_186_n 0.0186019f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_53 N_B1_c_49_n N_VPWR_c_189_n 0.00456932f $X=0.565 $Y=1.765 $X2=0 $Y2=0
cc_54 N_B1_c_49_n N_VPWR_c_184_n 0.00893078f $X=0.565 $Y=1.765 $X2=0 $Y2=0
cc_55 N_B1_c_48_n N_Y_c_215_n 0.00369403f $X=0.495 $Y=1.22 $X2=0 $Y2=0
cc_56 N_B1_c_49_n N_Y_c_215_n 9.25606e-19 $X=0.565 $Y=1.765 $X2=0 $Y2=0
cc_57 N_B1_c_49_n N_Y_c_217_n 0.0212918f $X=0.565 $Y=1.765 $X2=0 $Y2=0
cc_58 N_B1_c_48_n N_Y_c_216_n 0.0038858f $X=0.495 $Y=1.22 $X2=0 $Y2=0
cc_59 N_B1_c_49_n N_Y_c_216_n 0.0187954f $X=0.565 $Y=1.765 $X2=0 $Y2=0
cc_60 B1 N_Y_c_216_n 0.0249687f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_61 N_B1_c_48_n N_A_27_74#_c_247_n 0.0118798f $X=0.495 $Y=1.22 $X2=0 $Y2=0
cc_62 N_B1_c_48_n N_A_27_74#_c_252_n 0.0130776f $X=0.495 $Y=1.22 $X2=0 $Y2=0
cc_63 N_B1_c_49_n N_A_27_74#_c_252_n 0.00198538f $X=0.565 $Y=1.765 $X2=0 $Y2=0
cc_64 B1 N_A_27_74#_c_252_n 0.0260103f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_65 N_B1_c_48_n N_VGND_c_295_n 0.00291626f $X=0.495 $Y=1.22 $X2=0 $Y2=0
cc_66 N_B1_c_48_n N_VGND_c_298_n 0.00365046f $X=0.495 $Y=1.22 $X2=0 $Y2=0
cc_67 N_B2_c_71_n N_A3_c_98_n 0.0348973f $X=0.985 $Y=1.765 $X2=-0.19 $Y2=-0.245
cc_68 N_B2_c_73_n N_A3_c_98_n 0.00274949f $X=1.14 $Y=1.515 $X2=-0.19 $Y2=-0.245
cc_69 N_B2_M1006_g N_A3_M1003_g 0.0247403f $X=1.23 $Y=0.74 $X2=0 $Y2=0
cc_70 N_B2_c_71_n N_A3_c_100_n 0.00182653f $X=0.985 $Y=1.765 $X2=0 $Y2=0
cc_71 N_B2_c_73_n N_A3_c_100_n 0.0272873f $X=1.14 $Y=1.515 $X2=0 $Y2=0
cc_72 N_B2_c_71_n N_VPWR_c_189_n 0.00291513f $X=0.985 $Y=1.765 $X2=0 $Y2=0
cc_73 N_B2_c_71_n N_VPWR_c_184_n 0.0036081f $X=0.985 $Y=1.765 $X2=0 $Y2=0
cc_74 N_B2_c_71_n N_Y_c_215_n 0.00462376f $X=0.985 $Y=1.765 $X2=0 $Y2=0
cc_75 N_B2_M1006_g N_Y_c_215_n 0.00351046f $X=1.23 $Y=0.74 $X2=0 $Y2=0
cc_76 N_B2_c_73_n N_Y_c_215_n 0.0111437f $X=1.14 $Y=1.515 $X2=0 $Y2=0
cc_77 N_B2_c_71_n N_Y_c_217_n 0.0336287f $X=0.985 $Y=1.765 $X2=0 $Y2=0
cc_78 N_B2_c_73_n N_Y_c_217_n 0.0268169f $X=1.14 $Y=1.515 $X2=0 $Y2=0
cc_79 N_B2_c_71_n N_Y_c_216_n 0.0067159f $X=0.985 $Y=1.765 $X2=0 $Y2=0
cc_80 N_B2_M1006_g N_Y_c_216_n 0.00364258f $X=1.23 $Y=0.74 $X2=0 $Y2=0
cc_81 N_B2_c_73_n N_Y_c_216_n 0.0323503f $X=1.14 $Y=1.515 $X2=0 $Y2=0
cc_82 N_B2_M1006_g N_A_27_74#_c_247_n 0.0160377f $X=1.23 $Y=0.74 $X2=0 $Y2=0
cc_83 N_B2_M1006_g N_A_27_74#_c_250_n 0.0015383f $X=1.23 $Y=0.74 $X2=0 $Y2=0
cc_84 N_B2_M1006_g N_VGND_c_295_n 0.00291649f $X=1.23 $Y=0.74 $X2=0 $Y2=0
cc_85 N_B2_M1006_g N_VGND_c_298_n 0.00362117f $X=1.23 $Y=0.74 $X2=0 $Y2=0
cc_86 N_A3_c_98_n N_A2_c_130_n 0.0550125f $X=1.635 $Y=1.765 $X2=-0.19 $Y2=-0.245
cc_87 N_A3_c_100_n N_A2_c_130_n 0.00303987f $X=1.71 $Y=1.515 $X2=-0.19
+ $Y2=-0.245
cc_88 N_A3_M1003_g N_A2_M1007_g 0.0239043f $X=1.73 $Y=0.74 $X2=0 $Y2=0
cc_89 N_A3_c_98_n N_A2_c_132_n 0.00802653f $X=1.635 $Y=1.765 $X2=0 $Y2=0
cc_90 N_A3_c_100_n N_A2_c_132_n 0.0953748f $X=1.71 $Y=1.515 $X2=0 $Y2=0
cc_91 N_A3_c_98_n N_VPWR_c_189_n 0.00461464f $X=1.635 $Y=1.765 $X2=0 $Y2=0
cc_92 N_A3_c_98_n N_VPWR_c_184_n 0.00459895f $X=1.635 $Y=1.765 $X2=0 $Y2=0
cc_93 N_A3_c_100_n N_VPWR_c_184_n 0.0121164f $X=1.71 $Y=1.515 $X2=0 $Y2=0
cc_94 N_A3_c_98_n N_Y_c_217_n 0.0107259f $X=1.635 $Y=1.765 $X2=0 $Y2=0
cc_95 N_A3_c_100_n A_342_368# 0.00847117f $X=1.71 $Y=1.515 $X2=-0.19 $Y2=-0.245
cc_96 N_A3_M1003_g N_A_27_74#_c_248_n 0.00227966f $X=1.73 $Y=0.74 $X2=0 $Y2=0
cc_97 N_A3_M1003_g N_A_27_74#_c_260_n 0.00785824f $X=1.73 $Y=0.74 $X2=0 $Y2=0
cc_98 N_A3_c_98_n N_A_27_74#_c_249_n 4.86414e-19 $X=1.635 $Y=1.765 $X2=0 $Y2=0
cc_99 N_A3_M1003_g N_A_27_74#_c_249_n 0.0119119f $X=1.73 $Y=0.74 $X2=0 $Y2=0
cc_100 N_A3_c_100_n N_A_27_74#_c_249_n 0.0150021f $X=1.71 $Y=1.515 $X2=0 $Y2=0
cc_101 N_A3_c_98_n N_A_27_74#_c_250_n 8.5334e-19 $X=1.635 $Y=1.765 $X2=0 $Y2=0
cc_102 N_A3_M1003_g N_A_27_74#_c_250_n 0.00158144f $X=1.73 $Y=0.74 $X2=0 $Y2=0
cc_103 N_A3_c_100_n N_A_27_74#_c_250_n 0.0118341f $X=1.71 $Y=1.515 $X2=0 $Y2=0
cc_104 N_A3_M1003_g N_A_27_74#_c_251_n 9.95504e-19 $X=1.73 $Y=0.74 $X2=0 $Y2=0
cc_105 N_A3_M1003_g N_VGND_c_292_n 0.00624419f $X=1.73 $Y=0.74 $X2=0 $Y2=0
cc_106 N_A3_M1003_g N_VGND_c_295_n 0.00433139f $X=1.73 $Y=0.74 $X2=0 $Y2=0
cc_107 N_A3_M1003_g N_VGND_c_298_n 0.00818567f $X=1.73 $Y=0.74 $X2=0 $Y2=0
cc_108 N_A2_M1007_g N_A1_c_163_n 0.0199226f $X=2.33 $Y=0.74 $X2=-0.19 $Y2=-0.245
cc_109 N_A2_c_130_n N_A1_c_164_n 0.0529184f $X=2.205 $Y=1.765 $X2=0 $Y2=0
cc_110 N_A2_c_132_n N_A1_c_164_n 0.0144814f $X=2.28 $Y=1.515 $X2=0 $Y2=0
cc_111 N_A2_c_130_n A1 5.4813e-19 $X=2.205 $Y=1.765 $X2=0 $Y2=0
cc_112 N_A2_M1007_g A1 5.55987e-19 $X=2.33 $Y=0.74 $X2=0 $Y2=0
cc_113 N_A2_c_132_n A1 0.00716206f $X=2.28 $Y=1.515 $X2=0 $Y2=0
cc_114 N_A2_c_130_n N_VPWR_c_188_n 0.00183539f $X=2.205 $Y=1.765 $X2=0 $Y2=0
cc_115 N_A2_c_132_n N_VPWR_c_188_n 0.044568f $X=2.28 $Y=1.515 $X2=0 $Y2=0
cc_116 N_A2_c_130_n N_VPWR_c_189_n 0.00303293f $X=2.205 $Y=1.765 $X2=0 $Y2=0
cc_117 N_A2_c_132_n N_VPWR_c_189_n 0.0106761f $X=2.28 $Y=1.515 $X2=0 $Y2=0
cc_118 N_A2_c_130_n N_VPWR_c_184_n 0.00374185f $X=2.205 $Y=1.765 $X2=0 $Y2=0
cc_119 N_A2_c_132_n N_VPWR_c_184_n 0.0131295f $X=2.28 $Y=1.515 $X2=0 $Y2=0
cc_120 N_A2_c_132_n N_Y_c_217_n 0.0112454f $X=2.28 $Y=1.515 $X2=0 $Y2=0
cc_121 N_A2_c_132_n A_342_368# 0.0127084f $X=2.28 $Y=1.515 $X2=-0.19 $Y2=-0.245
cc_122 N_A2_c_132_n A_456_368# 0.0147038f $X=2.28 $Y=1.515 $X2=-0.19 $Y2=-0.245
cc_123 N_A2_M1007_g N_A_27_74#_c_260_n 9.49738e-19 $X=2.33 $Y=0.74 $X2=0 $Y2=0
cc_124 N_A2_c_130_n N_A_27_74#_c_249_n 0.00128341f $X=2.205 $Y=1.765 $X2=0 $Y2=0
cc_125 N_A2_M1007_g N_A_27_74#_c_249_n 0.013469f $X=2.33 $Y=0.74 $X2=0 $Y2=0
cc_126 N_A2_c_132_n N_A_27_74#_c_249_n 0.0320971f $X=2.28 $Y=1.515 $X2=0 $Y2=0
cc_127 N_A2_M1007_g N_A_27_74#_c_251_n 0.0104013f $X=2.33 $Y=0.74 $X2=0 $Y2=0
cc_128 N_A2_M1007_g N_VGND_c_292_n 0.00754067f $X=2.33 $Y=0.74 $X2=0 $Y2=0
cc_129 N_A2_M1007_g N_VGND_c_297_n 0.00434272f $X=2.33 $Y=0.74 $X2=0 $Y2=0
cc_130 N_A2_M1007_g N_VGND_c_298_n 0.00822293f $X=2.33 $Y=0.74 $X2=0 $Y2=0
cc_131 N_A1_c_164_n N_VPWR_c_188_n 0.0282242f $X=2.775 $Y=1.765 $X2=0 $Y2=0
cc_132 A1 N_VPWR_c_188_n 0.017092f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_133 N_A1_c_164_n N_VPWR_c_189_n 0.00413917f $X=2.775 $Y=1.765 $X2=0 $Y2=0
cc_134 N_A1_c_164_n N_VPWR_c_184_n 0.00818781f $X=2.775 $Y=1.765 $X2=0 $Y2=0
cc_135 N_A1_c_163_n N_A_27_74#_c_249_n 0.0100751f $X=2.76 $Y=1.22 $X2=0 $Y2=0
cc_136 N_A1_c_163_n N_A_27_74#_c_251_n 0.0081858f $X=2.76 $Y=1.22 $X2=0 $Y2=0
cc_137 N_A1_c_163_n N_VGND_c_294_n 0.00495522f $X=2.76 $Y=1.22 $X2=0 $Y2=0
cc_138 N_A1_c_164_n N_VGND_c_294_n 0.00180116f $X=2.775 $Y=1.765 $X2=0 $Y2=0
cc_139 A1 N_VGND_c_294_n 0.0221981f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_140 N_A1_c_163_n N_VGND_c_297_n 0.00434272f $X=2.76 $Y=1.22 $X2=0 $Y2=0
cc_141 N_A1_c_163_n N_VGND_c_298_n 0.00824124f $X=2.76 $Y=1.22 $X2=0 $Y2=0
cc_142 N_VPWR_c_189_n N_Y_c_217_n 0.0324699f $X=2.835 $Y=3.33 $X2=0 $Y2=0
cc_143 N_VPWR_c_184_n N_Y_c_217_n 0.026514f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_144 N_VPWR_c_186_n N_Y_c_216_n 0.0491356f $X=0.3 $Y=1.985 $X2=0 $Y2=0
cc_145 A_128_368# N_Y_c_217_n 0.0021653f $X=0.64 $Y=1.84 $X2=1.21 $Y2=2.115
cc_146 A_128_368# N_Y_c_216_n 0.00121878f $X=0.64 $Y=1.84 $X2=1.005 $Y2=1.95
cc_147 N_Y_M1008_d N_A_27_74#_c_247_n 0.00723582f $X=0.57 $Y=0.37 $X2=0 $Y2=0
cc_148 N_Y_c_215_n N_A_27_74#_c_247_n 0.0305034f $X=0.895 $Y=0.91 $X2=0 $Y2=0
cc_149 N_Y_c_215_n N_A_27_74#_c_250_n 0.00142263f $X=0.895 $Y=0.91 $X2=0 $Y2=0
cc_150 N_Y_c_216_n N_A_27_74#_c_250_n 0.00186133f $X=1.005 $Y=1.95 $X2=0 $Y2=0
cc_151 N_A_27_74#_c_249_n N_VGND_M1003_d 0.0048312f $X=2.38 $Y=1.095 $X2=-0.19
+ $Y2=-0.245
cc_152 N_A_27_74#_c_248_n N_VGND_c_292_n 0.00795492f $X=1.515 $Y=0.52 $X2=0
+ $Y2=0
cc_153 N_A_27_74#_c_249_n N_VGND_c_292_n 0.0228485f $X=2.38 $Y=1.095 $X2=0 $Y2=0
cc_154 N_A_27_74#_c_251_n N_VGND_c_292_n 0.031539f $X=2.545 $Y=0.515 $X2=0 $Y2=0
cc_155 N_A_27_74#_c_251_n N_VGND_c_294_n 0.0254897f $X=2.545 $Y=0.515 $X2=0
+ $Y2=0
cc_156 N_A_27_74#_c_247_n N_VGND_c_295_n 0.0358046f $X=1.35 $Y=0.435 $X2=0 $Y2=0
cc_157 N_A_27_74#_c_248_n N_VGND_c_295_n 0.0146502f $X=1.515 $Y=0.52 $X2=0 $Y2=0
cc_158 N_A_27_74#_c_252_n N_VGND_c_295_n 0.0146186f $X=0.28 $Y=0.515 $X2=0 $Y2=0
cc_159 N_A_27_74#_c_251_n N_VGND_c_297_n 0.0144922f $X=2.545 $Y=0.515 $X2=0
+ $Y2=0
cc_160 N_A_27_74#_c_247_n N_VGND_c_298_n 0.0306817f $X=1.35 $Y=0.435 $X2=0 $Y2=0
cc_161 N_A_27_74#_c_248_n N_VGND_c_298_n 0.0120674f $X=1.515 $Y=0.52 $X2=0 $Y2=0
cc_162 N_A_27_74#_c_251_n N_VGND_c_298_n 0.0118826f $X=2.545 $Y=0.515 $X2=0
+ $Y2=0
cc_163 N_A_27_74#_c_252_n N_VGND_c_298_n 0.0120551f $X=0.28 $Y=0.515 $X2=0 $Y2=0
