* NGSPICE file created from sky130_fd_sc_hs__fah_4.ext - technology: sky130A

.subckt sky130_fd_sc_hs__fah_4 A B CI VGND VNB VPB VPWR COUT SUM
M1000 a_427_362# a_586_257# a_536_114# VPB pshort w=840000u l=150000u
+  ad=6.202e+11p pd=5.22e+06u as=2.52e+11p ps=2.28e+06u
M1001 SUM a_1278_102# VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=6.832e+11p pd=5.7e+06u as=4.77725e+12p ps=2.973e+07u
M1002 VGND a_1278_102# SUM VNB nlowvt w=740000u l=150000u
+  ad=3.15805e+12p pd=2.382e+07u as=4.144e+11p ps=4.08e+06u
M1003 a_528_362# B a_427_362# VPB pshort w=840000u l=150000u
+  ad=2.562e+11p pd=2.29e+06u as=0p ps=0u
M1004 a_427_362# a_27_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=4.026e+11p pd=3.94e+06u as=0p ps=0u
M1005 COUT a_1265_379# VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=6.72e+11p pd=5.68e+06u as=0p ps=0u
M1006 VPWR a_1265_379# COUT VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 COUT a_1265_379# VGND VNB nlowvt w=740000u l=150000u
+  ad=4.144e+11p pd=4.08e+06u as=0p ps=0u
M1008 VPWR a_1265_379# COUT VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VGND a_1265_379# COUT VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_1265_379# a_528_362# a_586_257# VPB pshort w=840000u l=150000u
+  ad=3.738e+11p pd=2.57e+06u as=4.0435e+11p ps=3.01e+06u
M1011 VPWR A a_27_74# VPB pshort w=1e+06u l=150000u
+  ad=0p pd=0u as=2.95e+11p ps=2.59e+06u
M1012 a_200_74# A VPWR VPB pshort w=1e+06u l=150000u
+  ad=7.739e+11p pd=5.79e+06u as=0p ps=0u
M1013 a_427_362# a_27_74# VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_1378_125# a_536_114# a_1265_379# VPB pshort w=840000u l=150000u
+  ad=7.451e+11p pd=5.69e+06u as=0p ps=0u
M1015 VGND a_1265_379# COUT VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VPWR CI a_1378_125# VPB pshort w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_586_257# B VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 VGND CI a_1378_125# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=3.616e+11p ps=3.69e+06u
M1019 a_1278_102# a_528_362# a_1378_125# VPB pshort w=840000u l=150000u
+  ad=6.72e+11p pd=3.28e+06u as=0p ps=0u
M1020 a_536_114# B a_427_362# VNB nlowvt w=640000u l=150000u
+  ad=1.792e+11p pd=1.84e+06u as=0p ps=0u
M1021 SUM a_1278_102# VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 VPWR a_1278_102# SUM VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 VGND a_1378_125# a_1183_102# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=4.4305e+11p ps=3.95e+06u
M1024 a_1183_102# a_536_114# a_1278_102# VPB pshort w=840000u l=150000u
+  ad=3.90725e+11p pd=3e+06u as=0p ps=0u
M1025 a_1278_102# a_528_362# a_1183_102# VNB nlowvt w=640000u l=150000u
+  ad=2.44125e+11p pd=2.21e+06u as=0p ps=0u
M1026 COUT a_1265_379# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 VPWR a_1278_102# SUM VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1028 a_586_257# B VGND VNB nlowvt w=740000u l=150000u
+  ad=5.59925e+11p pd=5.19e+06u as=0p ps=0u
M1029 a_586_257# a_536_114# a_1265_379# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=2.3685e+11p ps=2.18e+06u
M1030 a_528_362# B a_200_74# VNB nlowvt w=640000u l=150000u
+  ad=2.048e+11p pd=1.92e+06u as=4.268e+11p ps=4.01e+06u
M1031 VPWR a_1378_125# a_1183_102# VPB pshort w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1032 SUM a_1278_102# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1033 a_200_74# a_586_257# a_536_114# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1034 VGND a_1278_102# SUM VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1035 COUT a_1265_379# VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1036 a_427_362# a_586_257# a_528_362# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1037 a_200_74# a_586_257# a_528_362# VPB pshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1038 VGND A a_27_74# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=1.824e+11p ps=1.85e+06u
M1039 a_200_74# A VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1040 a_1378_125# a_536_114# a_1278_102# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1041 a_1265_379# a_528_362# a_1378_125# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1042 a_536_114# B a_200_74# VPB pshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1043 SUM a_1278_102# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

