* NGSPICE file created from sky130_fd_sc_hs__and4bb_1.ext - technology: sky130A

.subckt sky130_fd_sc_hs__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
M1000 VPWR D a_179_48# VPB pshort w=840000u l=150000u
+  ad=1.3426e+12p pd=1.028e+07u as=5.46e+11p ps=4.66e+06u
M1001 a_179_48# a_27_74# VPWR VPB pshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1002 VPWR a_503_48# a_179_48# VPB pshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1003 VGND D a_647_74# VNB nlowvt w=640000u l=150000u
+  ad=5.299e+11p pd=4.38e+06u as=2.304e+11p ps=2e+06u
M1004 X a_179_48# VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=4.816e+11p pd=3.1e+06u as=0p ps=0u
M1005 X a_179_48# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1006 a_455_74# a_27_74# a_179_48# VNB nlowvt w=640000u l=150000u
+  ad=1.536e+11p pd=1.76e+06u as=1.824e+11p ps=1.85e+06u
M1007 a_533_74# a_503_48# a_455_74# VNB nlowvt w=640000u l=150000u
+  ad=2.688e+11p pd=2.12e+06u as=0p ps=0u
M1008 VPWR A_N a_27_74# VPB pshort w=840000u l=150000u
+  ad=0p pd=0u as=2.478e+11p ps=2.27e+06u
M1009 a_503_48# B_N VGND VNB nlowvt w=550000u l=150000u
+  ad=1.5675e+11p pd=1.67e+06u as=0p ps=0u
M1010 a_647_74# C a_533_74# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VGND A_N a_27_74# VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=1.5675e+11p ps=1.67e+06u
M1012 a_503_48# B_N VPWR VPB pshort w=840000u l=150000u
+  ad=2.478e+11p pd=2.27e+06u as=0p ps=0u
M1013 a_179_48# C VPWR VPB pshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

