* File: sky130_fd_sc_hs__einvp_1.pxi.spice
* Created: Tue Sep  1 20:04:57 2020
* 
x_PM_SKY130_FD_SC_HS__EINVP_1%TE N_TE_c_51_n N_TE_M1000_g N_TE_M1003_g
+ N_TE_c_46_n N_TE_c_47_n N_TE_M1001_g TE TE N_TE_c_50_n
+ PM_SKY130_FD_SC_HS__EINVP_1%TE
x_PM_SKY130_FD_SC_HS__EINVP_1%A_44_549# N_A_44_549#_M1003_s N_A_44_549#_M1000_s
+ N_A_44_549#_c_95_n N_A_44_549#_c_96_n N_A_44_549#_M1004_g N_A_44_549#_c_92_n
+ N_A_44_549#_c_93_n N_A_44_549#_c_94_n N_A_44_549#_c_98_n N_A_44_549#_c_99_n
+ N_A_44_549#_c_100_n PM_SKY130_FD_SC_HS__EINVP_1%A_44_549#
x_PM_SKY130_FD_SC_HS__EINVP_1%A N_A_M1005_g N_A_M1002_g N_A_c_140_n N_A_c_144_n
+ A N_A_c_141_n N_A_c_142_n PM_SKY130_FD_SC_HS__EINVP_1%A
x_PM_SKY130_FD_SC_HS__EINVP_1%VPWR N_VPWR_M1000_d N_VPWR_c_168_n VPWR
+ N_VPWR_c_169_n N_VPWR_c_170_n N_VPWR_c_167_n N_VPWR_c_172_n
+ PM_SKY130_FD_SC_HS__EINVP_1%VPWR
x_PM_SKY130_FD_SC_HS__EINVP_1%Z N_Z_M1002_d N_Z_M1005_d N_Z_c_196_n N_Z_c_197_n
+ N_Z_c_205_n N_Z_c_198_n N_Z_c_200_n Z Z PM_SKY130_FD_SC_HS__EINVP_1%Z
x_PM_SKY130_FD_SC_HS__EINVP_1%VGND N_VGND_M1003_d N_VGND_c_230_n VGND
+ N_VGND_c_231_n N_VGND_c_232_n N_VGND_c_233_n N_VGND_c_234_n
+ PM_SKY130_FD_SC_HS__EINVP_1%VGND
cc_1 VNB N_TE_M1003_g 0.0564205f $X=-0.19 $Y=-0.245 $X2=1.025 $Y2=0.58
cc_2 VNB N_TE_c_46_n 0.0273253f $X=-0.19 $Y=-0.245 $X2=1.44 $Y2=1.515
cc_3 VNB N_TE_c_47_n 0.0111253f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.515
cc_4 VNB N_TE_M1001_g 0.0293931f $X=-0.19 $Y=-0.245 $X2=1.515 $Y2=0.74
cc_5 VNB TE 0.00267865f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.58
cc_6 VNB N_TE_c_50_n 0.027005f $X=-0.19 $Y=-0.245 $X2=0.85 $Y2=1.605
cc_7 VNB N_A_44_549#_c_92_n 0.0311176f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.58
cc_8 VNB N_A_44_549#_c_93_n 0.0321729f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A_44_549#_c_94_n 0.0209133f $X=-0.19 $Y=-0.245 $X2=0.85 $Y2=1.605
cc_10 VNB N_A_M1002_g 0.0297146f $X=-0.19 $Y=-0.245 $X2=1.025 $Y2=0.58
cc_11 VNB N_A_c_140_n 0.00216621f $X=-0.19 $Y=-0.245 $X2=1.515 $Y2=1.44
cc_12 VNB N_A_c_141_n 0.0560278f $X=-0.19 $Y=-0.245 $X2=0.85 $Y2=1.605
cc_13 VNB N_A_c_142_n 0.00385705f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.605
cc_14 VNB N_VPWR_c_167_n 0.103974f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.605
cc_15 VNB N_Z_c_196_n 0.0103948f $X=-0.19 $Y=-0.245 $X2=1.44 $Y2=1.515
cc_16 VNB N_Z_c_197_n 0.0111859f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.515
cc_17 VNB N_Z_c_198_n 0.02581f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_VGND_c_230_n 0.0169975f $X=-0.19 $Y=-0.245 $X2=1.025 $Y2=0.58
cc_19 VNB N_VGND_c_231_n 0.032472f $X=-0.19 $Y=-0.245 $X2=1.515 $Y2=0.74
cc_20 VNB N_VGND_c_232_n 0.0307665f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.605
cc_21 VNB N_VGND_c_233_n 0.171006f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.605
cc_22 VNB N_VGND_c_234_n 0.00548191f $X=-0.19 $Y=-0.245 $X2=0.94 $Y2=1.662
cc_23 VPB N_TE_c_51_n 0.0188775f $X=-0.19 $Y=1.66 $X2=0.94 $Y2=1.885
cc_24 VPB N_TE_c_47_n 0.0180469f $X=-0.19 $Y=1.66 $X2=1.115 $Y2=1.515
cc_25 VPB TE 0.0108738f $X=-0.19 $Y=1.66 $X2=1.115 $Y2=1.58
cc_26 VPB N_TE_c_50_n 0.019406f $X=-0.19 $Y=1.66 $X2=0.85 $Y2=1.605
cc_27 VPB N_A_44_549#_c_95_n 0.0474067f $X=-0.19 $Y=1.66 $X2=1.115 $Y2=1.515
cc_28 VPB N_A_44_549#_c_96_n 0.0142212f $X=-0.19 $Y=1.66 $X2=1.515 $Y2=0.74
cc_29 VPB N_A_44_549#_c_92_n 0.0172107f $X=-0.19 $Y=1.66 $X2=1.115 $Y2=1.58
cc_30 VPB N_A_44_549#_c_98_n 0.0541373f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=1.605
cc_31 VPB N_A_44_549#_c_99_n 0.0624106f $X=-0.19 $Y=1.66 $X2=0.95 $Y2=1.662
cc_32 VPB N_A_44_549#_c_100_n 0.0295295f $X=-0.19 $Y=1.66 $X2=0.95 $Y2=1.605
cc_33 VPB N_A_c_140_n 0.013048f $X=-0.19 $Y=1.66 $X2=1.515 $Y2=1.44
cc_34 VPB N_A_c_144_n 0.02646f $X=-0.19 $Y=1.66 $X2=1.515 $Y2=0.74
cc_35 VPB N_A_c_142_n 0.00716996f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=1.605
cc_36 VPB N_VPWR_c_168_n 0.00684504f $X=-0.19 $Y=1.66 $X2=1.025 $Y2=0.58
cc_37 VPB N_VPWR_c_169_n 0.02821f $X=-0.19 $Y=1.66 $X2=1.515 $Y2=0.74
cc_38 VPB N_VPWR_c_170_n 0.0301422f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=1.605
cc_39 VPB N_VPWR_c_167_n 0.0582622f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=1.605
cc_40 VPB N_VPWR_c_172_n 0.00485691f $X=-0.19 $Y=1.66 $X2=0.94 $Y2=1.662
cc_41 VPB N_Z_c_196_n 0.0064074f $X=-0.19 $Y=1.66 $X2=1.44 $Y2=1.515
cc_42 VPB N_Z_c_200_n 0.0181642f $X=-0.19 $Y=1.66 $X2=0.85 $Y2=1.605
cc_43 VPB Z 0.0296006f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=1.605
cc_44 N_TE_c_51_n N_A_44_549#_c_95_n 9.93119e-19 $X=0.94 $Y=1.885 $X2=0 $Y2=0
cc_45 N_TE_c_51_n N_A_44_549#_c_96_n 0.0087198f $X=0.94 $Y=1.885 $X2=0 $Y2=0
cc_46 N_TE_c_46_n N_A_44_549#_c_96_n 0.0109392f $X=1.44 $Y=1.515 $X2=0 $Y2=0
cc_47 N_TE_c_47_n N_A_44_549#_c_96_n 0.00194304f $X=1.115 $Y=1.515 $X2=0 $Y2=0
cc_48 N_TE_c_51_n N_A_44_549#_c_92_n 0.00241632f $X=0.94 $Y=1.885 $X2=0 $Y2=0
cc_49 N_TE_M1003_g N_A_44_549#_c_92_n 0.00771354f $X=1.025 $Y=0.58 $X2=0 $Y2=0
cc_50 N_TE_c_47_n N_A_44_549#_c_92_n 0.0024586f $X=1.115 $Y=1.515 $X2=0 $Y2=0
cc_51 TE N_A_44_549#_c_92_n 0.0270525f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_52 N_TE_c_50_n N_A_44_549#_c_92_n 0.00228985f $X=0.85 $Y=1.605 $X2=0 $Y2=0
cc_53 N_TE_M1003_g N_A_44_549#_c_94_n 0.00711567f $X=1.025 $Y=0.58 $X2=0 $Y2=0
cc_54 TE N_A_44_549#_c_94_n 0.0228364f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_55 N_TE_c_50_n N_A_44_549#_c_94_n 0.0103126f $X=0.85 $Y=1.605 $X2=0 $Y2=0
cc_56 N_TE_c_51_n N_A_44_549#_c_98_n 0.00918669f $X=0.94 $Y=1.885 $X2=0 $Y2=0
cc_57 TE N_A_44_549#_c_98_n 0.0281262f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_58 N_TE_c_50_n N_A_44_549#_c_98_n 0.00287124f $X=0.85 $Y=1.605 $X2=0 $Y2=0
cc_59 N_TE_c_51_n N_A_44_549#_c_100_n 0.00143329f $X=0.94 $Y=1.885 $X2=0 $Y2=0
cc_60 N_TE_M1001_g N_A_M1002_g 0.0329902f $X=1.515 $Y=0.74 $X2=0 $Y2=0
cc_61 N_TE_c_46_n N_A_c_141_n 0.0329902f $X=1.44 $Y=1.515 $X2=0 $Y2=0
cc_62 N_TE_c_47_n N_A_c_141_n 0.00156384f $X=1.115 $Y=1.515 $X2=0 $Y2=0
cc_63 N_TE_c_51_n N_VPWR_c_168_n 0.00444601f $X=0.94 $Y=1.885 $X2=0 $Y2=0
cc_64 N_TE_c_46_n N_VPWR_c_168_n 0.00298784f $X=1.44 $Y=1.515 $X2=0 $Y2=0
cc_65 N_TE_c_47_n N_VPWR_c_168_n 2.13311e-19 $X=1.115 $Y=1.515 $X2=0 $Y2=0
cc_66 TE N_VPWR_c_168_n 0.0155105f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_67 N_TE_c_51_n N_VPWR_c_167_n 0.00168326f $X=0.94 $Y=1.885 $X2=0 $Y2=0
cc_68 N_TE_c_47_n N_Z_c_196_n 0.00182281f $X=1.115 $Y=1.515 $X2=0 $Y2=0
cc_69 N_TE_M1001_g N_Z_c_196_n 0.0091827f $X=1.515 $Y=0.74 $X2=0 $Y2=0
cc_70 TE N_Z_c_196_n 0.0189581f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_71 N_TE_M1001_g N_Z_c_205_n 7.6545e-19 $X=1.515 $Y=0.74 $X2=0 $Y2=0
cc_72 N_TE_M1001_g N_Z_c_198_n 0.00176373f $X=1.515 $Y=0.74 $X2=0 $Y2=0
cc_73 N_TE_M1003_g N_VGND_c_230_n 0.0101098f $X=1.025 $Y=0.58 $X2=0 $Y2=0
cc_74 N_TE_c_46_n N_VGND_c_230_n 0.00356442f $X=1.44 $Y=1.515 $X2=0 $Y2=0
cc_75 N_TE_M1001_g N_VGND_c_230_n 0.00387195f $X=1.515 $Y=0.74 $X2=0 $Y2=0
cc_76 TE N_VGND_c_230_n 0.00967694f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_77 N_TE_M1003_g N_VGND_c_231_n 0.00461464f $X=1.025 $Y=0.58 $X2=0 $Y2=0
cc_78 N_TE_M1001_g N_VGND_c_232_n 0.00461464f $X=1.515 $Y=0.74 $X2=0 $Y2=0
cc_79 N_TE_M1003_g N_VGND_c_233_n 0.00913453f $X=1.025 $Y=0.58 $X2=0 $Y2=0
cc_80 N_TE_M1001_g N_VGND_c_233_n 0.00907828f $X=1.515 $Y=0.74 $X2=0 $Y2=0
cc_81 N_A_44_549#_c_95_n N_A_c_144_n 0.00317858f $X=1.4 $Y=3.11 $X2=0 $Y2=0
cc_82 N_A_44_549#_c_96_n N_A_c_144_n 0.0505365f $X=1.475 $Y=3.035 $X2=0 $Y2=0
cc_83 N_A_44_549#_c_95_n N_VPWR_c_168_n 0.0224682f $X=1.4 $Y=3.11 $X2=0 $Y2=0
cc_84 N_A_44_549#_c_96_n N_VPWR_c_168_n 0.0166701f $X=1.475 $Y=3.035 $X2=0 $Y2=0
cc_85 N_A_44_549#_c_98_n N_VPWR_c_168_n 0.0781368f $X=0.715 $Y=2.175 $X2=0 $Y2=0
cc_86 N_A_44_549#_c_100_n N_VPWR_c_168_n 0.00121067f $X=0.89 $Y=2.965 $X2=0
+ $Y2=0
cc_87 N_A_44_549#_c_98_n N_VPWR_c_169_n 0.0538165f $X=0.715 $Y=2.175 $X2=0 $Y2=0
cc_88 N_A_44_549#_c_99_n N_VPWR_c_169_n 0.0207159f $X=0.725 $Y=2.91 $X2=0 $Y2=0
cc_89 N_A_44_549#_c_95_n N_VPWR_c_170_n 0.00538682f $X=1.4 $Y=3.11 $X2=0 $Y2=0
cc_90 N_A_44_549#_c_95_n N_VPWR_c_167_n 0.0188854f $X=1.4 $Y=3.11 $X2=0 $Y2=0
cc_91 N_A_44_549#_c_98_n N_VPWR_c_167_n 0.0274069f $X=0.715 $Y=2.175 $X2=0 $Y2=0
cc_92 N_A_44_549#_c_99_n N_VPWR_c_167_n 0.011903f $X=0.725 $Y=2.91 $X2=0 $Y2=0
cc_93 N_A_44_549#_c_100_n N_VPWR_c_167_n 0.00526618f $X=0.89 $Y=2.965 $X2=0
+ $Y2=0
cc_94 N_A_44_549#_c_96_n N_Z_c_196_n 0.00284788f $X=1.475 $Y=3.035 $X2=0 $Y2=0
cc_95 N_A_44_549#_c_96_n N_Z_c_200_n 0.00153573f $X=1.475 $Y=3.035 $X2=0 $Y2=0
cc_96 N_A_44_549#_c_96_n Z 0.00203425f $X=1.475 $Y=3.035 $X2=0 $Y2=0
cc_97 N_A_44_549#_c_96_n N_VGND_c_230_n 2.97864e-19 $X=1.475 $Y=3.035 $X2=0
+ $Y2=0
cc_98 N_A_44_549#_c_94_n N_VGND_c_230_n 0.0212724f $X=0.81 $Y=0.575 $X2=0 $Y2=0
cc_99 N_A_44_549#_c_93_n N_VGND_c_231_n 0.00610681f $X=0.275 $Y=0.735 $X2=0
+ $Y2=0
cc_100 N_A_44_549#_c_94_n N_VGND_c_231_n 0.0222861f $X=0.81 $Y=0.575 $X2=0 $Y2=0
cc_101 N_A_44_549#_c_93_n N_VGND_c_233_n 0.00604639f $X=0.275 $Y=0.735 $X2=0
+ $Y2=0
cc_102 N_A_44_549#_c_94_n N_VGND_c_233_n 0.0235867f $X=0.81 $Y=0.575 $X2=0 $Y2=0
cc_103 N_A_c_144_n N_VPWR_c_168_n 0.00276443f $X=1.902 $Y=1.885 $X2=0 $Y2=0
cc_104 N_A_c_144_n N_VPWR_c_170_n 0.00445602f $X=1.902 $Y=1.885 $X2=0 $Y2=0
cc_105 N_A_c_144_n N_VPWR_c_167_n 0.00861507f $X=1.902 $Y=1.885 $X2=0 $Y2=0
cc_106 N_A_M1002_g N_Z_c_196_n 0.0104807f $X=1.905 $Y=0.74 $X2=0 $Y2=0
cc_107 N_A_c_144_n N_Z_c_196_n 0.00288515f $X=1.902 $Y=1.885 $X2=0 $Y2=0
cc_108 N_A_c_142_n N_Z_c_196_n 0.0360328f $X=2.11 $Y=1.465 $X2=0 $Y2=0
cc_109 N_A_M1002_g N_Z_c_197_n 0.0151759f $X=1.905 $Y=0.74 $X2=0 $Y2=0
cc_110 N_A_c_141_n N_Z_c_197_n 0.00232659f $X=2.11 $Y=1.465 $X2=0 $Y2=0
cc_111 N_A_c_142_n N_Z_c_197_n 0.0282627f $X=2.11 $Y=1.465 $X2=0 $Y2=0
cc_112 N_A_M1002_g N_Z_c_198_n 0.0123878f $X=1.905 $Y=0.74 $X2=0 $Y2=0
cc_113 N_A_c_144_n N_Z_c_200_n 0.0207334f $X=1.902 $Y=1.885 $X2=0 $Y2=0
cc_114 N_A_c_141_n N_Z_c_200_n 0.00148544f $X=2.11 $Y=1.465 $X2=0 $Y2=0
cc_115 N_A_c_142_n N_Z_c_200_n 0.0279341f $X=2.11 $Y=1.465 $X2=0 $Y2=0
cc_116 N_A_c_144_n Z 0.0124682f $X=1.902 $Y=1.885 $X2=0 $Y2=0
cc_117 N_A_M1002_g N_VGND_c_232_n 0.00434272f $X=1.905 $Y=0.74 $X2=0 $Y2=0
cc_118 N_A_M1002_g N_VGND_c_233_n 0.00824638f $X=1.905 $Y=0.74 $X2=0 $Y2=0
cc_119 N_VPWR_c_168_n Z 0.0205017f $X=1.25 $Y=2.105 $X2=0 $Y2=0
cc_120 N_VPWR_c_170_n Z 0.0146324f $X=2.16 $Y=3.33 $X2=0 $Y2=0
cc_121 N_VPWR_c_167_n Z 0.0120616f $X=2.16 $Y=3.33 $X2=0 $Y2=0
cc_122 A_310_392# N_Z_c_200_n 0.00701052f $X=1.55 $Y=1.96 $X2=2.12 $Y2=2.115
cc_123 N_Z_c_205_n N_VGND_c_230_n 0.00156525f $X=1.775 $Y=1.045 $X2=0 $Y2=0
cc_124 N_Z_c_198_n N_VGND_c_230_n 0.00927251f $X=2.12 $Y=0.515 $X2=0 $Y2=0
cc_125 N_Z_c_198_n N_VGND_c_232_n 0.0145639f $X=2.12 $Y=0.515 $X2=0 $Y2=0
cc_126 N_Z_c_198_n N_VGND_c_233_n 0.0119984f $X=2.12 $Y=0.515 $X2=0 $Y2=0
cc_127 N_Z_c_205_n A_318_74# 0.00570883f $X=1.775 $Y=1.045 $X2=-0.19 $Y2=-0.245
