* File: sky130_fd_sc_hs__o2bb2a_2.pex.spice
* Created: Tue Sep  1 20:16:47 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HS__O2BB2A_2%B1 3 5 7 8 12
r23 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.405
+ $Y=1.615 $X2=0.405 $Y2=1.615
r24 8 12 5.76222 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=0.24 $Y=1.615
+ $X2=0.405 $Y2=1.615
r25 5 11 55.187 $w=3.04e-07 $l=3.11769e-07 $layer=POLY_cond $X=0.51 $Y=1.885
+ $X2=0.42 $Y2=1.615
r26 5 7 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=0.51 $Y=1.885
+ $X2=0.51 $Y2=2.46
r27 1 11 38.539 $w=3.04e-07 $l=1.98997e-07 $layer=POLY_cond $X=0.495 $Y=1.45
+ $X2=0.42 $Y2=1.615
r28 1 3 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=0.495 $Y=1.45
+ $X2=0.495 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HS__O2BB2A_2%B2 3 5 7 8
r29 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.975
+ $Y=1.615 $X2=0.975 $Y2=1.615
r30 8 12 7.85757 $w=3.28e-07 $l=2.25e-07 $layer=LI1_cond $X=1.2 $Y=1.615
+ $X2=0.975 $Y2=1.615
r31 5 11 55.8646 $w=2.93e-07 $l=2.91633e-07 $layer=POLY_cond $X=0.93 $Y=1.885
+ $X2=0.975 $Y2=1.615
r32 5 7 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=0.93 $Y=1.885
+ $X2=0.93 $Y2=2.46
r33 1 11 38.5916 $w=2.93e-07 $l=1.88348e-07 $layer=POLY_cond $X=0.925 $Y=1.45
+ $X2=0.975 $Y2=1.615
r34 1 3 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=0.925 $Y=1.45
+ $X2=0.925 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HS__O2BB2A_2%A_270_48# 1 2 9 11 13 17 18 19 20 22 26 29
+ 31
c68 29 0 1.41594e-19 $X=1.62 $Y=1.615
r69 29 32 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=1.62 $Y=1.615
+ $X2=1.62 $Y2=1.78
r70 29 31 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=1.62 $Y=1.615
+ $X2=1.62 $Y2=1.45
r71 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.62
+ $Y=1.615 $X2=1.62 $Y2=1.615
r72 24 26 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=2.21 $Y=1.135
+ $X2=2.21 $Y2=0.81
r73 20 22 26.2757 $w=2.48e-07 $l=5.7e-07 $layer=LI1_cond $X=1.785 $Y=2.1
+ $X2=2.355 $Y2=2.1
r74 18 24 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.045 $Y=1.22
+ $X2=2.21 $Y2=1.135
r75 18 19 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=2.045 $Y=1.22
+ $X2=1.785 $Y2=1.22
r76 17 20 7.14316 $w=2.5e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.7 $Y=1.975
+ $X2=1.785 $Y2=2.1
r77 17 32 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=1.7 $Y=1.975
+ $X2=1.7 $Y2=1.78
r78 14 19 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.7 $Y=1.305
+ $X2=1.785 $Y2=1.22
r79 14 31 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=1.7 $Y=1.305
+ $X2=1.7 $Y2=1.45
r80 11 30 52.6712 $w=3.73e-07 $l=3.27399e-07 $layer=POLY_cond $X=1.44 $Y=1.885
+ $X2=1.567 $Y2=1.615
r81 11 13 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=1.44 $Y=1.885
+ $X2=1.44 $Y2=2.46
r82 7 30 39.1028 $w=3.73e-07 $l=2.25067e-07 $layer=POLY_cond $X=1.425 $Y=1.45
+ $X2=1.567 $Y2=1.615
r83 7 9 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=1.425 $Y=1.45
+ $X2=1.425 $Y2=0.74
r84 2 22 600 $w=1.7e-07 $l=2.68608e-07 $layer=licon1_PDIFF $count=1 $X=2.16
+ $Y=1.965 $X2=2.355 $Y2=2.14
r85 1 26 182 $w=1.7e-07 $l=5.07346e-07 $layer=licon1_NDIFF $count=1 $X=2.065
+ $Y=0.37 $X2=2.21 $Y2=0.81
.ends

.subckt PM_SKY130_FD_SC_HS__O2BB2A_2%A2_N 1 3 5 6 8 11 13
c44 5 0 1.41594e-19 $X=2.25 $Y=1.475
r45 13 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.16
+ $Y=1.64 $X2=2.16 $Y2=1.64
r46 9 11 89.734 $w=1.5e-07 $l=1.75e-07 $layer=POLY_cond $X=2.25 $Y=1.16
+ $X2=2.425 $Y2=1.16
r47 6 11 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.425 $Y=1.085
+ $X2=2.425 $Y2=1.16
r48 6 8 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=2.425 $Y=1.085
+ $X2=2.425 $Y2=0.69
r49 5 16 38.5562 $w=2.99e-07 $l=2.05122e-07 $layer=POLY_cond $X=2.25 $Y=1.475
+ $X2=2.16 $Y2=1.64
r50 4 9 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.25 $Y=1.235 $X2=2.25
+ $Y2=1.16
r51 4 5 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=2.25 $Y=1.235 $X2=2.25
+ $Y2=1.475
r52 1 16 52.2586 $w=2.99e-07 $l=2.85044e-07 $layer=POLY_cond $X=2.085 $Y=1.89
+ $X2=2.16 $Y2=1.64
r53 1 3 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=2.085 $Y=1.89
+ $X2=2.085 $Y2=2.385
.ends

.subckt PM_SKY130_FD_SC_HS__O2BB2A_2%A1_N 1 3 6 8
c38 8 0 1.85545e-19 $X=2.64 $Y=1.665
c39 6 0 1.63062e-19 $X=2.815 $Y=0.69
r40 8 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.7 $Y=1.64
+ $X2=2.7 $Y2=1.64
r41 4 11 38.5462 $w=3.19e-07 $l=2.10286e-07 $layer=POLY_cond $X=2.815 $Y=1.475
+ $X2=2.712 $Y2=1.64
r42 4 6 402.521 $w=1.5e-07 $l=7.85e-07 $layer=POLY_cond $X=2.815 $Y=1.475
+ $X2=2.815 $Y2=0.69
r43 1 11 51.3895 $w=3.19e-07 $l=2.90259e-07 $layer=POLY_cond $X=2.625 $Y=1.89
+ $X2=2.712 $Y2=1.64
r44 1 3 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=2.625 $Y=1.89
+ $X2=2.625 $Y2=2.385
.ends

.subckt PM_SKY130_FD_SC_HS__O2BB2A_2%A_201_392# 1 2 7 9 12 16 18 20 23 27 29 33
+ 35 36 38 39 40 41 42 43 51
c121 51 0 1.85545e-19 $X=3.81 $Y=1.535
c122 7 0 3.55965e-20 $X=3.365 $Y=1.765
r123 51 52 0.621134 $w=3.88e-07 $l=5e-09 $layer=POLY_cond $X=3.81 $Y=1.535
+ $X2=3.815 $Y2=1.535
r124 50 51 53.4175 $w=3.88e-07 $l=4.3e-07 $layer=POLY_cond $X=3.38 $Y=1.535
+ $X2=3.81 $Y2=1.535
r125 49 50 1.8634 $w=3.88e-07 $l=1.5e-08 $layer=POLY_cond $X=3.365 $Y=1.535
+ $X2=3.38 $Y2=1.535
r126 47 49 12.4227 $w=3.88e-07 $l=1e-07 $layer=POLY_cond $X=3.265 $Y=1.535
+ $X2=3.365 $Y2=1.535
r127 46 47 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.265
+ $Y=1.47 $X2=3.265 $Y2=1.47
r128 41 46 9.03377 $w=2.85e-07 $l=2.03912e-07 $layer=LI1_cond $X=3.17 $Y=1.635
+ $X2=3.257 $Y2=1.47
r129 41 42 49.5829 $w=1.68e-07 $l=7.6e-07 $layer=LI1_cond $X=3.17 $Y=1.635
+ $X2=3.17 $Y2=2.395
r130 39 46 10.7018 $w=2.85e-07 $l=3.24808e-07 $layer=LI1_cond $X=3.085 $Y=1.22
+ $X2=3.257 $Y2=1.47
r131 39 40 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=3.085 $Y=1.22
+ $X2=2.715 $Y2=1.22
r132 38 40 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.63 $Y=1.135
+ $X2=2.715 $Y2=1.22
r133 37 38 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=2.63 $Y=0.425
+ $X2=2.63 $Y2=1.135
r134 35 37 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.545 $Y=0.34
+ $X2=2.63 $Y2=0.425
r135 35 36 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=2.545 $Y=0.34
+ $X2=1.805 $Y2=0.34
r136 31 36 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.64 $Y=0.425
+ $X2=1.805 $Y2=0.34
r137 31 33 2.44458 $w=3.28e-07 $l=7e-08 $layer=LI1_cond $X=1.64 $Y=0.425
+ $X2=1.64 $Y2=0.495
r138 30 43 3.80956 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.38 $Y=2.48
+ $X2=1.215 $Y2=2.48
r139 29 42 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.085 $Y=2.48
+ $X2=3.17 $Y2=2.395
r140 29 30 111.235 $w=1.68e-07 $l=1.705e-06 $layer=LI1_cond $X=3.085 $Y=2.48
+ $X2=1.38 $Y2=2.48
r141 25 43 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.215 $Y=2.565
+ $X2=1.215 $Y2=2.48
r142 25 27 8.73063 $w=3.28e-07 $l=2.5e-07 $layer=LI1_cond $X=1.215 $Y=2.565
+ $X2=1.215 $Y2=2.815
r143 21 43 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.215 $Y=2.395
+ $X2=1.215 $Y2=2.48
r144 21 23 9.7783 $w=3.28e-07 $l=2.8e-07 $layer=LI1_cond $X=1.215 $Y=2.395
+ $X2=1.215 $Y2=2.115
r145 18 52 25.1189 $w=1.5e-07 $l=2.3e-07 $layer=POLY_cond $X=3.815 $Y=1.765
+ $X2=3.815 $Y2=1.535
r146 18 20 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.815 $Y=1.765
+ $X2=3.815 $Y2=2.4
r147 14 51 25.1189 $w=1.5e-07 $l=2.3e-07 $layer=POLY_cond $X=3.81 $Y=1.305
+ $X2=3.81 $Y2=1.535
r148 14 16 289.713 $w=1.5e-07 $l=5.65e-07 $layer=POLY_cond $X=3.81 $Y=1.305
+ $X2=3.81 $Y2=0.74
r149 10 50 25.1189 $w=1.5e-07 $l=2.3e-07 $layer=POLY_cond $X=3.38 $Y=1.305
+ $X2=3.38 $Y2=1.535
r150 10 12 289.713 $w=1.5e-07 $l=5.65e-07 $layer=POLY_cond $X=3.38 $Y=1.305
+ $X2=3.38 $Y2=0.74
r151 7 49 25.1189 $w=1.5e-07 $l=2.3e-07 $layer=POLY_cond $X=3.365 $Y=1.765
+ $X2=3.365 $Y2=1.535
r152 7 9 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.365 $Y=1.765
+ $X2=3.365 $Y2=2.4
r153 2 27 400 $w=1.7e-07 $l=9.54241e-07 $layer=licon1_PDIFF $count=1 $X=1.005
+ $Y=1.96 $X2=1.215 $Y2=2.815
r154 2 23 400 $w=1.7e-07 $l=2.76857e-07 $layer=licon1_PDIFF $count=1 $X=1.005
+ $Y=1.96 $X2=1.215 $Y2=2.115
r155 1 33 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=1.5
+ $Y=0.37 $X2=1.64 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_HS__O2BB2A_2%VPWR 1 2 3 4 13 15 21 25 27 29 33 35 40 45
+ 54 57 61
c53 15 0 1.42909e-19 $X=0.285 $Y=2.115
r54 60 61 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r55 57 58 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r56 54 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r57 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r58 49 61 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.08 $Y2=3.33
r59 49 58 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=3.12 $Y2=3.33
r60 48 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r61 46 57 10.5822 $w=1.7e-07 $l=2.25e-07 $layer=LI1_cond $X=3.22 $Y=3.33
+ $X2=2.995 $Y2=3.33
r62 46 48 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=3.22 $Y=3.33 $X2=3.6
+ $Y2=3.33
r63 45 60 4.01252 $w=1.7e-07 $l=1.82e-07 $layer=LI1_cond $X=3.955 $Y=3.33
+ $X2=4.137 $Y2=3.33
r64 45 48 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=3.955 $Y=3.33
+ $X2=3.6 $Y2=3.33
r65 44 58 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r66 43 44 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r67 41 54 9.05715 $w=1.7e-07 $l=1.78e-07 $layer=LI1_cond $X=1.94 $Y=3.33
+ $X2=1.762 $Y2=3.33
r68 41 43 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=1.94 $Y=3.33 $X2=2.64
+ $Y2=3.33
r69 40 57 10.5822 $w=1.7e-07 $l=2.25e-07 $layer=LI1_cond $X=2.77 $Y=3.33
+ $X2=2.995 $Y2=3.33
r70 40 43 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=2.77 $Y=3.33
+ $X2=2.64 $Y2=3.33
r71 39 55 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=1.68 $Y2=3.33
r72 39 52 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.24 $Y2=3.33
r73 38 39 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r74 36 51 4.72267 $w=1.7e-07 $l=2.25e-07 $layer=LI1_cond $X=0.45 $Y=3.33
+ $X2=0.225 $Y2=3.33
r75 36 38 48.9305 $w=1.68e-07 $l=7.5e-07 $layer=LI1_cond $X=0.45 $Y=3.33 $X2=1.2
+ $Y2=3.33
r76 35 54 9.05715 $w=1.7e-07 $l=1.77e-07 $layer=LI1_cond $X=1.585 $Y=3.33
+ $X2=1.762 $Y2=3.33
r77 35 38 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=1.585 $Y=3.33
+ $X2=1.2 $Y2=3.33
r78 33 44 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r79 33 55 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.68 $Y2=3.33
r80 29 32 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=4.08 $Y=1.985
+ $X2=4.08 $Y2=2.815
r81 27 60 3.13065 $w=2.5e-07 $l=1.09864e-07 $layer=LI1_cond $X=4.08 $Y=3.245
+ $X2=4.137 $Y2=3.33
r82 27 32 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=4.08 $Y=3.245
+ $X2=4.08 $Y2=2.815
r83 23 57 1.79621 $w=4.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.995 $Y=3.245
+ $X2=2.995 $Y2=3.33
r84 23 25 9.16993 $w=4.48e-07 $l=3.45e-07 $layer=LI1_cond $X=2.995 $Y=3.245
+ $X2=2.995 $Y2=2.9
r85 19 54 1.11826 $w=3.55e-07 $l=8.5e-08 $layer=LI1_cond $X=1.762 $Y=3.245
+ $X2=1.762 $Y2=3.33
r86 19 21 11.1998 $w=3.53e-07 $l=3.45e-07 $layer=LI1_cond $X=1.762 $Y=3.245
+ $X2=1.762 $Y2=2.9
r87 15 18 24.4458 $w=3.28e-07 $l=7e-07 $layer=LI1_cond $X=0.285 $Y=2.115
+ $X2=0.285 $Y2=2.815
r88 13 51 3.0435 $w=3.3e-07 $l=1.11018e-07 $layer=LI1_cond $X=0.285 $Y=3.245
+ $X2=0.225 $Y2=3.33
r89 13 18 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=0.285 $Y=3.245
+ $X2=0.285 $Y2=2.815
r90 4 32 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=3.89
+ $Y=1.84 $X2=4.04 $Y2=2.815
r91 4 29 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=3.89
+ $Y=1.84 $X2=4.04 $Y2=1.985
r92 3 25 600 $w=1.7e-07 $l=1.0724e-06 $layer=licon1_PDIFF $count=1 $X=2.7
+ $Y=1.965 $X2=2.995 $Y2=2.9
r93 2 21 600 $w=1.7e-07 $l=1.05541e-06 $layer=licon1_PDIFF $count=1 $X=1.515
+ $Y=1.96 $X2=1.76 $Y2=2.9
r94 1 18 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=0.14
+ $Y=1.96 $X2=0.285 $Y2=2.815
r95 1 15 400 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_PDIFF $count=1 $X=0.14
+ $Y=1.96 $X2=0.285 $Y2=2.115
.ends

.subckt PM_SKY130_FD_SC_HS__O2BB2A_2%X 1 2 9 13 14 15 16 23 32
c32 32 0 3.55965e-20 $X=3.597 $Y=1.82
c33 9 0 1.63062e-19 $X=3.595 $Y=0.515
r34 21 23 1.43638 $w=3.43e-07 $l=4.3e-08 $layer=LI1_cond $X=3.597 $Y=1.992
+ $X2=3.597 $Y2=2.035
r35 15 16 12.3595 $w=3.43e-07 $l=3.7e-07 $layer=LI1_cond $X=3.597 $Y=2.405
+ $X2=3.597 $Y2=2.775
r36 14 21 0.701487 $w=3.43e-07 $l=2.1e-08 $layer=LI1_cond $X=3.597 $Y=1.971
+ $X2=3.597 $Y2=1.992
r37 14 32 8.01174 $w=3.43e-07 $l=1.51e-07 $layer=LI1_cond $X=3.597 $Y=1.971
+ $X2=3.597 $Y2=1.82
r38 14 15 11.658 $w=3.43e-07 $l=3.49e-07 $layer=LI1_cond $X=3.597 $Y=2.056
+ $X2=3.597 $Y2=2.405
r39 14 23 0.701487 $w=3.43e-07 $l=2.1e-08 $layer=LI1_cond $X=3.597 $Y=2.056
+ $X2=3.597 $Y2=2.035
r40 13 32 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=3.685 $Y=1.13
+ $X2=3.685 $Y2=1.82
r41 7 13 8.64139 $w=3.38e-07 $l=1.7e-07 $layer=LI1_cond $X=3.6 $Y=0.96 $X2=3.6
+ $Y2=1.13
r42 7 9 15.0834 $w=3.38e-07 $l=4.45e-07 $layer=LI1_cond $X=3.6 $Y=0.96 $X2=3.6
+ $Y2=0.515
r43 2 14 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=3.44
+ $Y=1.84 $X2=3.59 $Y2=1.985
r44 2 16 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=3.44
+ $Y=1.84 $X2=3.59 $Y2=2.815
r45 1 9 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.455
+ $Y=0.37 $X2=3.595 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__O2BB2A_2%A_27_74# 1 2 9 11 12 15
c26 12 0 1.42909e-19 $X=0.365 $Y=1.195
r27 13 15 27.4281 $w=2.48e-07 $l=5.95e-07 $layer=LI1_cond $X=1.18 $Y=1.11
+ $X2=1.18 $Y2=0.515
r28 11 13 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.055 $Y=1.195
+ $X2=1.18 $Y2=1.11
r29 11 12 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.055 $Y=1.195
+ $X2=0.365 $Y2=1.195
r30 7 12 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.24 $Y=1.11
+ $X2=0.365 $Y2=1.195
r31 7 9 27.4281 $w=2.48e-07 $l=5.95e-07 $layer=LI1_cond $X=0.24 $Y=1.11 $X2=0.24
+ $Y2=0.515
r32 2 15 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1 $Y=0.37
+ $X2=1.14 $Y2=0.515
r33 1 9 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__O2BB2A_2%VGND 1 2 3 12 16 18 20 22 24 29 37 43 46 50
r51 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r52 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r53 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r54 41 50 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.08
+ $Y2=0
r55 41 47 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=3.12
+ $Y2=0
r56 40 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r57 38 46 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.215 $Y=0 $X2=3.05
+ $Y2=0
r58 38 40 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=3.215 $Y=0 $X2=3.6
+ $Y2=0
r59 37 49 3.99177 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.94 $Y=0 $X2=4.13
+ $Y2=0
r60 37 40 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=3.94 $Y=0 $X2=3.6
+ $Y2=0
r61 36 47 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r62 35 36 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r63 33 44 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r64 32 35 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.2 $Y=0 $X2=2.64
+ $Y2=0
r65 32 33 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r66 30 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.875 $Y=0 $X2=0.71
+ $Y2=0
r67 30 32 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.875 $Y=0 $X2=1.2
+ $Y2=0
r68 29 46 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.885 $Y=0 $X2=3.05
+ $Y2=0
r69 29 35 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=2.885 $Y=0 $X2=2.64
+ $Y2=0
r70 27 44 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r71 26 27 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r72 24 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.545 $Y=0 $X2=0.71
+ $Y2=0
r73 24 26 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.545 $Y=0 $X2=0.24
+ $Y2=0
r74 22 36 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r75 22 33 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.2
+ $Y2=0
r76 18 49 3.1514 $w=2.5e-07 $l=1.12916e-07 $layer=LI1_cond $X=4.065 $Y=0.085
+ $X2=4.13 $Y2=0
r77 18 20 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=4.065 $Y=0.085
+ $X2=4.065 $Y2=0.515
r78 14 46 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.05 $Y=0.085
+ $X2=3.05 $Y2=0
r79 14 16 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=3.05 $Y=0.085
+ $X2=3.05 $Y2=0.495
r80 10 43 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.71 $Y=0.085
+ $X2=0.71 $Y2=0
r81 10 12 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=0.71 $Y=0.085
+ $X2=0.71 $Y2=0.495
r82 3 20 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.885
+ $Y=0.37 $X2=4.025 $Y2=0.515
r83 2 16 91 $w=1.7e-07 $l=2.13542e-07 $layer=licon1_NDIFF $count=2 $X=2.89
+ $Y=0.37 $X2=3.05 $Y2=0.495
r84 1 12 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=0.57
+ $Y=0.37 $X2=0.71 $Y2=0.495
.ends

