* File: sky130_fd_sc_hs__sdfbbn_1.pxi.spice
* Created: Thu Aug 27 21:07:51 2020
* 
x_PM_SKY130_FD_SC_HS__SDFBBN_1%SCD N_SCD_c_375_n N_SCD_c_380_n N_SCD_c_381_n
+ N_SCD_M1020_g N_SCD_M1004_g N_SCD_c_382_n SCD N_SCD_c_377_n N_SCD_c_378_n
+ PM_SKY130_FD_SC_HS__SDFBBN_1%SCD
x_PM_SKY130_FD_SC_HS__SDFBBN_1%D N_D_M1023_g N_D_M1000_g N_D_c_412_n N_D_c_413_n
+ D N_D_c_411_n PM_SKY130_FD_SC_HS__SDFBBN_1%D
x_PM_SKY130_FD_SC_HS__SDFBBN_1%A_353_93# N_A_353_93#_M1018_d N_A_353_93#_M1013_d
+ N_A_353_93#_c_469_n N_A_353_93#_M1034_g N_A_353_93#_c_476_n
+ N_A_353_93#_M1029_g N_A_353_93#_c_470_n N_A_353_93#_c_477_n
+ N_A_353_93#_c_471_n N_A_353_93#_c_478_n N_A_353_93#_c_472_n
+ N_A_353_93#_c_473_n N_A_353_93#_c_474_n N_A_353_93#_c_475_n
+ N_A_353_93#_c_482_n N_A_353_93#_c_483_n PM_SKY130_FD_SC_HS__SDFBBN_1%A_353_93#
x_PM_SKY130_FD_SC_HS__SDFBBN_1%SCE N_SCE_M1033_g N_SCE_c_569_n N_SCE_c_570_n
+ N_SCE_M1014_g N_SCE_c_560_n N_SCE_c_561_n N_SCE_M1018_g N_SCE_c_563_n
+ N_SCE_c_564_n N_SCE_c_571_n N_SCE_M1013_g N_SCE_c_565_n N_SCE_c_566_n
+ N_SCE_c_574_n N_SCE_c_575_n SCE N_SCE_c_568_n PM_SKY130_FD_SC_HS__SDFBBN_1%SCE
x_PM_SKY130_FD_SC_HS__SDFBBN_1%CLK_N N_CLK_N_M1015_g N_CLK_N_c_665_n
+ N_CLK_N_M1040_g CLK_N N_CLK_N_c_666_n PM_SKY130_FD_SC_HS__SDFBBN_1%CLK_N
x_PM_SKY130_FD_SC_HS__SDFBBN_1%A_977_243# N_A_977_243#_M1003_d
+ N_A_977_243#_M1046_s N_A_977_243#_M1026_d N_A_977_243#_c_703_n
+ N_A_977_243#_c_704_n N_A_977_243#_c_712_n N_A_977_243#_M1011_g
+ N_A_977_243#_M1021_g N_A_977_243#_M1043_g N_A_977_243#_c_707_n
+ N_A_977_243#_M1012_g N_A_977_243#_c_714_n N_A_977_243#_c_708_n
+ N_A_977_243#_c_716_n N_A_977_243#_c_717_n N_A_977_243#_c_718_n
+ N_A_977_243#_c_719_n N_A_977_243#_c_777_p N_A_977_243#_c_709_n
+ N_A_977_243#_c_779_p N_A_977_243#_c_751_p N_A_977_243#_c_721_n
+ N_A_977_243#_c_710_n N_A_977_243#_c_723_n N_A_977_243#_c_724_n
+ N_A_977_243#_c_725_n N_A_977_243#_c_726_n N_A_977_243#_c_711_n
+ N_A_977_243#_c_781_p N_A_977_243#_c_727_n
+ PM_SKY130_FD_SC_HS__SDFBBN_1%A_977_243#
x_PM_SKY130_FD_SC_HS__SDFBBN_1%A_867_82# N_A_867_82#_M1016_d N_A_867_82#_M1045_d
+ N_A_867_82#_c_922_n N_A_867_82#_c_923_n N_A_867_82#_M1030_g
+ N_A_867_82#_M1001_g N_A_867_82#_c_904_n N_A_867_82#_M1044_g
+ N_A_867_82#_M1039_g N_A_867_82#_c_906_n N_A_867_82#_c_907_n
+ N_A_867_82#_c_926_n N_A_867_82#_c_908_n N_A_867_82#_c_909_n
+ N_A_867_82#_c_910_n N_A_867_82#_c_911_n N_A_867_82#_c_912_n
+ N_A_867_82#_c_913_n N_A_867_82#_c_914_n N_A_867_82#_c_915_n
+ N_A_867_82#_c_916_n N_A_867_82#_c_917_n N_A_867_82#_c_918_n
+ N_A_867_82#_c_919_n N_A_867_82#_c_920_n N_A_867_82#_c_921_n
+ PM_SKY130_FD_SC_HS__SDFBBN_1%A_867_82#
x_PM_SKY130_FD_SC_HS__SDFBBN_1%A_1159_497# N_A_1159_497#_M1017_d
+ N_A_1159_497#_M1030_d N_A_1159_497#_c_1124_n N_A_1159_497#_c_1125_n
+ N_A_1159_497#_c_1126_n N_A_1159_497#_c_1134_n N_A_1159_497#_M1046_g
+ N_A_1159_497#_c_1127_n N_A_1159_497#_M1003_g N_A_1159_497#_c_1128_n
+ N_A_1159_497#_c_1129_n N_A_1159_497#_c_1135_n N_A_1159_497#_c_1130_n
+ N_A_1159_497#_c_1131_n N_A_1159_497#_c_1136_n N_A_1159_497#_c_1132_n
+ N_A_1159_497#_c_1138_n PM_SKY130_FD_SC_HS__SDFBBN_1%A_1159_497#
x_PM_SKY130_FD_SC_HS__SDFBBN_1%A_1579_258# N_A_1579_258#_M1002_s
+ N_A_1579_258#_M1009_s N_A_1579_258#_c_1221_n N_A_1579_258#_c_1243_n
+ N_A_1579_258#_M1022_g N_A_1579_258#_M1047_g N_A_1579_258#_c_1223_n
+ N_A_1579_258#_M1038_g N_A_1579_258#_c_1224_n N_A_1579_258#_c_1225_n
+ N_A_1579_258#_c_1245_n N_A_1579_258#_M1035_g N_A_1579_258#_c_1226_n
+ N_A_1579_258#_c_1227_n N_A_1579_258#_c_1228_n N_A_1579_258#_c_1229_n
+ N_A_1579_258#_c_1230_n N_A_1579_258#_c_1231_n N_A_1579_258#_c_1232_n
+ N_A_1579_258#_c_1233_n N_A_1579_258#_c_1234_n N_A_1579_258#_c_1235_n
+ N_A_1579_258#_c_1236_n N_A_1579_258#_c_1247_n N_A_1579_258#_c_1248_n
+ N_A_1579_258#_c_1237_n N_A_1579_258#_c_1238_n N_A_1579_258#_c_1239_n
+ N_A_1579_258#_c_1240_n N_A_1579_258#_c_1241_n
+ PM_SKY130_FD_SC_HS__SDFBBN_1%A_1579_258#
x_PM_SKY130_FD_SC_HS__SDFBBN_1%SET_B N_SET_B_c_1429_n N_SET_B_M1026_g
+ N_SET_B_M1025_g N_SET_B_c_1424_n N_SET_B_M1042_g N_SET_B_M1007_g
+ N_SET_B_c_1431_n N_SET_B_c_1432_n N_SET_B_c_1426_n SET_B N_SET_B_c_1427_n
+ N_SET_B_c_1428_n PM_SKY130_FD_SC_HS__SDFBBN_1%SET_B
x_PM_SKY130_FD_SC_HS__SDFBBN_1%A_662_82# N_A_662_82#_M1015_s N_A_662_82#_M1040_s
+ N_A_662_82#_M1016_g N_A_662_82#_c_1559_n N_A_662_82#_M1045_g
+ N_A_662_82#_c_1560_n N_A_662_82#_c_1561_n N_A_662_82#_M1017_g
+ N_A_662_82#_c_1563_n N_A_662_82#_c_1564_n N_A_662_82#_c_1576_n
+ N_A_662_82#_M1031_g N_A_662_82#_M1027_g N_A_662_82#_c_1566_n
+ N_A_662_82#_c_1567_n N_A_662_82#_c_1577_n N_A_662_82#_M1041_g
+ N_A_662_82#_c_1568_n N_A_662_82#_c_1569_n N_A_662_82#_c_1578_n
+ N_A_662_82#_c_1570_n N_A_662_82#_c_1571_n N_A_662_82#_c_1580_n
+ N_A_662_82#_c_1581_n N_A_662_82#_c_1603_n N_A_662_82#_c_1572_n
+ N_A_662_82#_c_1582_n N_A_662_82#_c_1573_n
+ PM_SKY130_FD_SC_HS__SDFBBN_1%A_662_82#
x_PM_SKY130_FD_SC_HS__SDFBBN_1%A_2133_410# N_A_2133_410#_M1038_d
+ N_A_2133_410#_M1042_s N_A_2133_410#_M1008_d N_A_2133_410#_c_1756_n
+ N_A_2133_410#_M1024_g N_A_2133_410#_c_1757_n N_A_2133_410#_M1010_g
+ N_A_2133_410#_c_1743_n N_A_2133_410#_M1006_g N_A_2133_410#_M1005_g
+ N_A_2133_410#_c_1745_n N_A_2133_410#_c_1746_n N_A_2133_410#_c_1762_n
+ N_A_2133_410#_M1028_g N_A_2133_410#_M1019_g N_A_2133_410#_c_1748_n
+ N_A_2133_410#_c_1763_n N_A_2133_410#_c_1894_p N_A_2133_410#_c_1764_n
+ N_A_2133_410#_c_1749_n N_A_2133_410#_c_1765_n N_A_2133_410#_c_1766_n
+ N_A_2133_410#_c_1767_n N_A_2133_410#_c_1750_n N_A_2133_410#_c_1751_n
+ N_A_2133_410#_c_1752_n N_A_2133_410#_c_1753_n N_A_2133_410#_c_1868_p
+ N_A_2133_410#_c_1858_p N_A_2133_410#_c_1768_n N_A_2133_410#_c_1769_n
+ N_A_2133_410#_c_1770_n N_A_2133_410#_c_1794_n N_A_2133_410#_c_1754_n
+ N_A_2133_410#_c_1755_n PM_SKY130_FD_SC_HS__SDFBBN_1%A_2133_410#
x_PM_SKY130_FD_SC_HS__SDFBBN_1%A_1954_119# N_A_1954_119#_M1027_d
+ N_A_1954_119#_M1044_d N_A_1954_119#_M1032_g N_A_1954_119#_c_1977_n
+ N_A_1954_119#_M1008_g N_A_1954_119#_c_1984_n N_A_1954_119#_c_1985_n
+ N_A_1954_119#_c_1986_n N_A_1954_119#_c_1987_n N_A_1954_119#_c_1978_n
+ N_A_1954_119#_c_1979_n N_A_1954_119#_c_1989_n N_A_1954_119#_c_1990_n
+ N_A_1954_119#_c_1991_n N_A_1954_119#_c_1992_n N_A_1954_119#_c_1980_n
+ N_A_1954_119#_c_1981_n N_A_1954_119#_c_1982_n N_A_1954_119#_c_1996_n
+ N_A_1954_119#_c_2016_n N_A_1954_119#_c_2019_n N_A_1954_119#_c_2064_n
+ PM_SKY130_FD_SC_HS__SDFBBN_1%A_1954_119#
x_PM_SKY130_FD_SC_HS__SDFBBN_1%RESET_B N_RESET_B_c_2124_n N_RESET_B_M1009_g
+ N_RESET_B_c_2121_n N_RESET_B_M1002_g N_RESET_B_c_2125_n N_RESET_B_c_2126_n
+ N_RESET_B_c_2127_n RESET_B N_RESET_B_c_2123_n
+ PM_SKY130_FD_SC_HS__SDFBBN_1%RESET_B
x_PM_SKY130_FD_SC_HS__SDFBBN_1%A_3078_384# N_A_3078_384#_M1019_s
+ N_A_3078_384#_M1028_s N_A_3078_384#_c_2174_n N_A_3078_384#_M1037_g
+ N_A_3078_384#_c_2175_n N_A_3078_384#_M1036_g N_A_3078_384#_c_2176_n
+ N_A_3078_384#_c_2177_n N_A_3078_384#_c_2178_n N_A_3078_384#_c_2179_n
+ PM_SKY130_FD_SC_HS__SDFBBN_1%A_3078_384#
x_PM_SKY130_FD_SC_HS__SDFBBN_1%A_27_464# N_A_27_464#_M1020_s N_A_27_464#_M1029_d
+ N_A_27_464#_c_2226_n N_A_27_464#_c_2227_n N_A_27_464#_c_2228_n
+ N_A_27_464#_c_2229_n N_A_27_464#_c_2230_n N_A_27_464#_c_2231_n
+ N_A_27_464#_c_2232_n PM_SKY130_FD_SC_HS__SDFBBN_1%A_27_464#
x_PM_SKY130_FD_SC_HS__SDFBBN_1%VPWR N_VPWR_M1020_d N_VPWR_M1013_s N_VPWR_M1040_d
+ N_VPWR_M1011_s N_VPWR_M1022_d N_VPWR_M1012_s N_VPWR_M1024_d N_VPWR_M1042_d
+ N_VPWR_M1009_d N_VPWR_M1028_d N_VPWR_c_2277_n N_VPWR_c_2278_n N_VPWR_c_2279_n
+ N_VPWR_c_2280_n N_VPWR_c_2281_n N_VPWR_c_2282_n N_VPWR_c_2283_n
+ N_VPWR_c_2284_n N_VPWR_c_2285_n N_VPWR_c_2286_n N_VPWR_c_2287_n
+ N_VPWR_c_2288_n N_VPWR_c_2289_n N_VPWR_c_2290_n N_VPWR_c_2291_n VPWR
+ N_VPWR_c_2292_n N_VPWR_c_2293_n N_VPWR_c_2294_n N_VPWR_c_2295_n
+ N_VPWR_c_2296_n N_VPWR_c_2297_n N_VPWR_c_2298_n N_VPWR_c_2276_n
+ N_VPWR_c_2300_n N_VPWR_c_2301_n N_VPWR_c_2302_n N_VPWR_c_2303_n
+ N_VPWR_c_2304_n N_VPWR_c_2305_n N_VPWR_c_2306_n
+ PM_SKY130_FD_SC_HS__SDFBBN_1%VPWR
x_PM_SKY130_FD_SC_HS__SDFBBN_1%A_197_119# N_A_197_119#_M1033_d
+ N_A_197_119#_M1001_d N_A_197_119#_M1023_d N_A_197_119#_M1031_d
+ N_A_197_119#_c_2467_n N_A_197_119#_c_2489_n N_A_197_119#_c_2503_n
+ N_A_197_119#_c_2468_n N_A_197_119#_c_2490_n N_A_197_119#_c_2491_n
+ N_A_197_119#_c_2469_n N_A_197_119#_c_2470_n N_A_197_119#_c_2471_n
+ N_A_197_119#_c_2472_n N_A_197_119#_c_2473_n N_A_197_119#_c_2474_n
+ N_A_197_119#_c_2475_n N_A_197_119#_c_2476_n N_A_197_119#_c_2477_n
+ N_A_197_119#_c_2478_n N_A_197_119#_c_2479_n N_A_197_119#_c_2480_n
+ N_A_197_119#_c_2481_n N_A_197_119#_c_2482_n N_A_197_119#_c_2483_n
+ N_A_197_119#_c_2493_n N_A_197_119#_c_2484_n N_A_197_119#_c_2485_n
+ N_A_197_119#_c_2486_n N_A_197_119#_c_2487_n N_A_197_119#_c_2495_n
+ N_A_197_119#_c_2488_n N_A_197_119#_c_2543_n N_A_197_119#_c_2496_n
+ PM_SKY130_FD_SC_HS__SDFBBN_1%A_197_119#
x_PM_SKY130_FD_SC_HS__SDFBBN_1%Q_N N_Q_N_M1005_d N_Q_N_M1006_d N_Q_N_c_2701_n
+ N_Q_N_c_2702_n Q_N Q_N Q_N Q_N N_Q_N_c_2703_n PM_SKY130_FD_SC_HS__SDFBBN_1%Q_N
x_PM_SKY130_FD_SC_HS__SDFBBN_1%Q N_Q_M1037_d N_Q_M1036_d N_Q_c_2736_n
+ N_Q_c_2737_n Q Q Q Q N_Q_c_2738_n PM_SKY130_FD_SC_HS__SDFBBN_1%Q
x_PM_SKY130_FD_SC_HS__SDFBBN_1%VGND N_VGND_M1004_s N_VGND_M1034_d N_VGND_M1015_d
+ N_VGND_M1021_s N_VGND_M1025_d N_VGND_M1010_d N_VGND_M1002_d N_VGND_M1019_d
+ N_VGND_c_2759_n N_VGND_c_2760_n N_VGND_c_2761_n N_VGND_c_2762_n
+ N_VGND_c_2763_n N_VGND_c_2764_n N_VGND_c_2765_n N_VGND_c_2766_n
+ N_VGND_c_2767_n N_VGND_c_2768_n N_VGND_c_2769_n VGND N_VGND_c_2770_n
+ N_VGND_c_2771_n N_VGND_c_2772_n N_VGND_c_2773_n N_VGND_c_2774_n
+ N_VGND_c_2775_n N_VGND_c_2776_n N_VGND_c_2777_n N_VGND_c_2778_n
+ N_VGND_c_2779_n N_VGND_c_2780_n N_VGND_c_2781_n
+ PM_SKY130_FD_SC_HS__SDFBBN_1%VGND
x_PM_SKY130_FD_SC_HS__SDFBBN_1%A_1434_78# N_A_1434_78#_M1003_s
+ N_A_1434_78#_M1047_d N_A_1434_78#_c_2931_n N_A_1434_78#_c_2932_n
+ N_A_1434_78#_c_2933_n PM_SKY130_FD_SC_HS__SDFBBN_1%A_1434_78#
x_PM_SKY130_FD_SC_HS__SDFBBN_1%A_2392_74# N_A_2392_74#_M1007_d
+ N_A_2392_74#_M1032_d N_A_2392_74#_c_2967_n N_A_2392_74#_c_2964_n
+ N_A_2392_74#_c_2965_n N_A_2392_74#_c_2966_n
+ PM_SKY130_FD_SC_HS__SDFBBN_1%A_2392_74#
cc_1 VNB N_SCD_c_375_n 0.0227054f $X=-0.19 $Y=-0.245 $X2=0.407 $Y2=1.688
cc_2 VNB N_SCD_M1004_g 0.0273411f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=0.805
cc_3 VNB N_SCD_c_377_n 0.021705f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.37
cc_4 VNB N_SCD_c_378_n 0.0188539f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.37
cc_5 VNB N_D_M1000_g 0.0354137f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=1.205
cc_6 VNB D 0.00112383f $X=-0.19 $Y=-0.245 $X2=0.407 $Y2=1.875
cc_7 VNB N_D_c_411_n 0.0216752f $X=-0.19 $Y=-0.245 $X2=0.407 $Y2=1.205
cc_8 VNB N_A_353_93#_c_469_n 0.0145006f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.64
cc_9 VNB N_A_353_93#_c_470_n 0.0138306f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_353_93#_c_471_n 0.0262529f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.54
cc_11 VNB N_A_353_93#_c_472_n 0.00493697f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_353_93#_c_473_n 0.0128457f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_353_93#_c_474_n 0.0285641f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_353_93#_c_475_n 0.00213819f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_SCE_M1033_g 0.0362506f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.155
cc_16 VNB N_SCE_c_560_n 0.133608f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=0.805
cc_17 VNB N_SCE_c_561_n 0.0125534f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_SCE_M1018_g 0.0297697f $X=-0.19 $Y=-0.245 $X2=0.407 $Y2=1.37
cc_19 VNB N_SCE_c_563_n 0.0339866f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.37
cc_20 VNB N_SCE_c_564_n 0.00851842f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.37
cc_21 VNB N_SCE_c_565_n 0.0208752f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.54
cc_22 VNB N_SCE_c_566_n 0.0161476f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB SCE 0.00821433f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_SCE_c_568_n 0.0148961f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_CLK_N_M1015_g 0.0241624f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.875
cc_26 VNB N_CLK_N_c_665_n 0.0360955f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.245
cc_27 VNB N_CLK_N_c_666_n 0.00169104f $X=-0.19 $Y=-0.245 $X2=0.407 $Y2=1.875
cc_28 VNB N_A_977_243#_c_703_n 0.0419268f $X=-0.19 $Y=-0.245 $X2=0.407 $Y2=1.875
cc_29 VNB N_A_977_243#_c_704_n 0.0110024f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_30 VNB N_A_977_243#_M1021_g 0.0220427f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.54
cc_31 VNB N_A_977_243#_M1043_g 0.0381377f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_977_243#_c_707_n 0.00678187f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_977_243#_c_708_n 0.0213071f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_977_243#_c_709_n 0.00420798f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_977_243#_c_710_n 6.05461e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_977_243#_c_711_n 0.0014623f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_867_82#_M1001_g 0.036728f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_867_82#_c_904_n 0.00703065f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.37
cc_39 VNB N_A_867_82#_M1039_g 0.0304832f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_867_82#_c_906_n 0.00558857f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_867_82#_c_907_n 0.0010045f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_867_82#_c_908_n 0.00746161f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_867_82#_c_909_n 0.00184814f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_867_82#_c_910_n 0.0085399f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_A_867_82#_c_911_n 0.0319986f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_A_867_82#_c_912_n 0.00193806f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_867_82#_c_913_n 0.0148502f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_867_82#_c_914_n 0.00476988f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A_867_82#_c_915_n 0.0187935f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_A_867_82#_c_916_n 0.00209826f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_A_867_82#_c_917_n 0.00113735f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_A_867_82#_c_918_n 0.00165111f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_A_867_82#_c_919_n 0.00886767f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_A_867_82#_c_920_n 0.00552553f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_A_867_82#_c_921_n 0.0014707f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_A_1159_497#_c_1124_n 0.0111865f $X=-0.19 $Y=-0.245 $X2=0.505
+ $Y2=2.64
cc_57 VNB N_A_1159_497#_c_1125_n 0.0179103f $X=-0.19 $Y=-0.245 $X2=0.52
+ $Y2=1.205
cc_58 VNB N_A_1159_497#_c_1126_n 0.0116842f $X=-0.19 $Y=-0.245 $X2=0.52
+ $Y2=0.805
cc_59 VNB N_A_1159_497#_c_1127_n 0.017554f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_A_1159_497#_c_1128_n 0.00887168f $X=-0.19 $Y=-0.245 $X2=0.407
+ $Y2=1.205
cc_61 VNB N_A_1159_497#_c_1129_n 0.00193935f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_A_1159_497#_c_1130_n 0.0111908f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_A_1159_497#_c_1131_n 0.00228138f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_A_1159_497#_c_1132_n 0.0166784f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_A_1579_258#_c_1221_n 0.00209711f $X=-0.19 $Y=-0.245 $X2=0.52
+ $Y2=1.205
cc_66 VNB N_A_1579_258#_M1047_g 0.0197908f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_A_1579_258#_c_1223_n 0.0164382f $X=-0.19 $Y=-0.245 $X2=0.385
+ $Y2=1.37
cc_68 VNB N_A_1579_258#_c_1224_n 0.0336392f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.54
cc_69 VNB N_A_1579_258#_c_1225_n 0.00647592f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_A_1579_258#_c_1226_n 0.0186774f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_A_1579_258#_c_1227_n 0.00354122f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_A_1579_258#_c_1228_n 0.0224474f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_A_1579_258#_c_1229_n 0.00293678f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_A_1579_258#_c_1230_n 0.00432188f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_A_1579_258#_c_1231_n 0.00106807f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_A_1579_258#_c_1232_n 0.0158167f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_A_1579_258#_c_1233_n 0.0066041f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_A_1579_258#_c_1234_n 0.0250737f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VNB N_A_1579_258#_c_1235_n 0.00679517f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_A_1579_258#_c_1236_n 0.00329409f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_81 VNB N_A_1579_258#_c_1237_n 0.00624835f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_82 VNB N_A_1579_258#_c_1238_n 0.046662f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_83 VNB N_A_1579_258#_c_1239_n 0.00553857f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_84 VNB N_A_1579_258#_c_1240_n 0.0110986f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_85 VNB N_A_1579_258#_c_1241_n 0.00755219f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_86 VNB N_SET_B_M1025_g 0.0363875f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.64
cc_87 VNB N_SET_B_c_1424_n 0.0195298f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=1.205
cc_88 VNB N_SET_B_M1007_g 0.0308675f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_89 VNB N_SET_B_c_1426_n 0.00112279f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.54
cc_90 VNB N_SET_B_c_1427_n 0.00715852f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_91 VNB N_SET_B_c_1428_n 0.00167869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_92 VNB N_A_662_82#_M1016_g 0.0257732f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=0.805
cc_93 VNB N_A_662_82#_c_1559_n 0.0264437f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_94 VNB N_A_662_82#_c_1560_n 0.120023f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_95 VNB N_A_662_82#_c_1561_n 0.012503f $X=-0.19 $Y=-0.245 $X2=0.407 $Y2=1.37
cc_96 VNB N_A_662_82#_M1017_g 0.0243939f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.54
cc_97 VNB N_A_662_82#_c_1563_n 0.0250852f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_98 VNB N_A_662_82#_c_1564_n 0.268142f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.54
cc_99 VNB N_A_662_82#_M1027_g 0.0319784f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_100 VNB N_A_662_82#_c_1566_n 0.0368616f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_101 VNB N_A_662_82#_c_1567_n 0.00998153f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_102 VNB N_A_662_82#_c_1568_n 0.00749069f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_103 VNB N_A_662_82#_c_1569_n 0.0102676f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_104 VNB N_A_662_82#_c_1570_n 0.0182949f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_105 VNB N_A_662_82#_c_1571_n 0.0121316f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_106 VNB N_A_662_82#_c_1572_n 0.00363763f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_107 VNB N_A_662_82#_c_1573_n 0.0030213f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_108 VNB N_A_2133_410#_M1010_g 0.0473009f $X=-0.19 $Y=-0.245 $X2=0.385
+ $Y2=1.37
cc_109 VNB N_A_2133_410#_c_1743_n 0.0142932f $X=-0.19 $Y=-0.245 $X2=0.24
+ $Y2=1.54
cc_110 VNB N_A_2133_410#_M1005_g 0.0275425f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_111 VNB N_A_2133_410#_c_1745_n 0.0558622f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_112 VNB N_A_2133_410#_c_1746_n 0.00620589f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_113 VNB N_A_2133_410#_M1019_g 0.0397683f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_114 VNB N_A_2133_410#_c_1748_n 0.00814373f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_115 VNB N_A_2133_410#_c_1749_n 0.0070078f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_116 VNB N_A_2133_410#_c_1750_n 0.00688383f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_117 VNB N_A_2133_410#_c_1751_n 0.0166675f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_118 VNB N_A_2133_410#_c_1752_n 0.00370574f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_119 VNB N_A_2133_410#_c_1753_n 0.00213162f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_120 VNB N_A_2133_410#_c_1754_n 0.00151338f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_121 VNB N_A_2133_410#_c_1755_n 0.00158697f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_122 VNB N_A_1954_119#_M1032_g 0.0360248f $X=-0.19 $Y=-0.245 $X2=0.52
+ $Y2=0.805
cc_123 VNB N_A_1954_119#_c_1977_n 0.00771253f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_124 VNB N_A_1954_119#_c_1978_n 0.00444826f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_125 VNB N_A_1954_119#_c_1979_n 0.00675177f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_126 VNB N_A_1954_119#_c_1980_n 0.00183819f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_127 VNB N_A_1954_119#_c_1981_n 5.83966e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_128 VNB N_A_1954_119#_c_1982_n 0.0217424f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_129 VNB N_RESET_B_c_2121_n 0.0190564f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.155
cc_130 VNB RESET_B 0.00269444f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_131 VNB N_RESET_B_c_2123_n 0.0374009f $X=-0.19 $Y=-0.245 $X2=0.407 $Y2=1.205
cc_132 VNB N_A_3078_384#_c_2174_n 0.0221821f $X=-0.19 $Y=-0.245 $X2=0.505
+ $Y2=2.64
cc_133 VNB N_A_3078_384#_c_2175_n 0.0410143f $X=-0.19 $Y=-0.245 $X2=0.52
+ $Y2=0.805
cc_134 VNB N_A_3078_384#_c_2176_n 0.00512138f $X=-0.19 $Y=-0.245 $X2=0.407
+ $Y2=1.37
cc_135 VNB N_A_3078_384#_c_2177_n 6.69403e-19 $X=-0.19 $Y=-0.245 $X2=0.24
+ $Y2=1.54
cc_136 VNB N_A_3078_384#_c_2178_n 0.00750762f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_137 VNB N_A_3078_384#_c_2179_n 6.16118e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_138 VNB N_VPWR_c_2276_n 0.701046f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_139 VNB N_A_197_119#_c_2467_n 0.00166563f $X=-0.19 $Y=-0.245 $X2=0.155
+ $Y2=1.58
cc_140 VNB N_A_197_119#_c_2468_n 0.00762811f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_141 VNB N_A_197_119#_c_2469_n 0.00306689f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_142 VNB N_A_197_119#_c_2470_n 0.0116365f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_143 VNB N_A_197_119#_c_2471_n 0.005791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_144 VNB N_A_197_119#_c_2472_n 0.0155497f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_145 VNB N_A_197_119#_c_2473_n 0.00175986f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_146 VNB N_A_197_119#_c_2474_n 0.00209615f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_147 VNB N_A_197_119#_c_2475_n 0.0107432f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_148 VNB N_A_197_119#_c_2476_n 0.00432316f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_149 VNB N_A_197_119#_c_2477_n 0.0101445f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_150 VNB N_A_197_119#_c_2478_n 0.0169648f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_151 VNB N_A_197_119#_c_2479_n 7.36253e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_152 VNB N_A_197_119#_c_2480_n 0.00266478f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_153 VNB N_A_197_119#_c_2481_n 0.013783f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_154 VNB N_A_197_119#_c_2482_n 0.00159638f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_155 VNB N_A_197_119#_c_2483_n 0.00796442f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_156 VNB N_A_197_119#_c_2484_n 0.00463588f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_157 VNB N_A_197_119#_c_2485_n 3.77841e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_158 VNB N_A_197_119#_c_2486_n 0.002372f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_159 VNB N_A_197_119#_c_2487_n 0.00549494f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_160 VNB N_A_197_119#_c_2488_n 0.00233877f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_161 VNB N_Q_N_c_2701_n 0.0104326f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=0.805
cc_162 VNB N_Q_N_c_2702_n 0.00486315f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_163 VNB N_Q_N_c_2703_n 0.00217925f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_164 VNB N_Q_c_2736_n 0.0237144f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=0.805
cc_165 VNB N_Q_c_2737_n 0.00768928f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_166 VNB N_Q_c_2738_n 0.0286887f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_167 VNB N_VGND_c_2759_n 0.0130142f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_168 VNB N_VGND_c_2760_n 0.0425426f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_169 VNB N_VGND_c_2761_n 0.0113535f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_170 VNB N_VGND_c_2762_n 0.0211187f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_171 VNB N_VGND_c_2763_n 0.00653047f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_172 VNB N_VGND_c_2764_n 0.0087522f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_173 VNB N_VGND_c_2765_n 0.00994235f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_174 VNB N_VGND_c_2766_n 0.0181999f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_175 VNB N_VGND_c_2767_n 0.0577044f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_176 VNB N_VGND_c_2768_n 0.0320808f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_177 VNB N_VGND_c_2769_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_178 VNB N_VGND_c_2770_n 0.042432f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_179 VNB N_VGND_c_2771_n 0.0375776f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_180 VNB N_VGND_c_2772_n 0.0311959f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_181 VNB N_VGND_c_2773_n 0.0743167f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_182 VNB N_VGND_c_2774_n 0.0651782f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_183 VNB N_VGND_c_2775_n 0.0197156f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_184 VNB N_VGND_c_2776_n 0.828436f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_185 VNB N_VGND_c_2777_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_186 VNB N_VGND_c_2778_n 0.0152596f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_187 VNB N_VGND_c_2779_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_188 VNB N_VGND_c_2780_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_189 VNB N_VGND_c_2781_n 0.00596557f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_190 VNB N_A_1434_78#_c_2931_n 0.0225961f $X=-0.19 $Y=-0.245 $X2=0.505
+ $Y2=2.64
cc_191 VNB N_A_1434_78#_c_2932_n 0.00591938f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_192 VNB N_A_1434_78#_c_2933_n 0.00881632f $X=-0.19 $Y=-0.245 $X2=0.155
+ $Y2=1.58
cc_193 VNB N_A_2392_74#_c_2964_n 0.00350421f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_194 VNB N_A_2392_74#_c_2965_n 0.00203957f $X=-0.19 $Y=-0.245 $X2=0.407
+ $Y2=1.875
cc_195 VNB N_A_2392_74#_c_2966_n 0.00423102f $X=-0.19 $Y=-0.245 $X2=0.155
+ $Y2=1.58
cc_196 VPB N_SCD_c_375_n 0.00229605f $X=-0.19 $Y=1.66 $X2=0.407 $Y2=1.688
cc_197 VPB N_SCD_c_380_n 0.0214913f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.155
cc_198 VPB N_SCD_c_381_n 0.0255701f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.245
cc_199 VPB N_SCD_c_382_n 0.0209206f $X=-0.19 $Y=1.66 $X2=0.407 $Y2=1.875
cc_200 VPB N_SCD_c_378_n 0.00912284f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.37
cc_201 VPB N_D_c_412_n 0.0176873f $X=-0.19 $Y=1.66 $X2=0.52 $Y2=0.805
cc_202 VPB N_D_c_413_n 0.022875f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_203 VPB D 9.35477e-19 $X=-0.19 $Y=1.66 $X2=0.407 $Y2=1.875
cc_204 VPB N_D_c_411_n 0.0195092f $X=-0.19 $Y=1.66 $X2=0.407 $Y2=1.205
cc_205 VPB N_A_353_93#_c_476_n 0.0184888f $X=-0.19 $Y=1.66 $X2=0.52 $Y2=0.805
cc_206 VPB N_A_353_93#_c_477_n 0.0150433f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.37
cc_207 VPB N_A_353_93#_c_478_n 0.0318957f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_208 VPB N_A_353_93#_c_472_n 0.00411221f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_209 VPB N_A_353_93#_c_474_n 0.0359665f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_210 VPB N_A_353_93#_c_475_n 0.00238114f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_211 VPB N_A_353_93#_c_482_n 0.0114266f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_212 VPB N_A_353_93#_c_483_n 0.00793835f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_213 VPB N_SCE_c_569_n 0.014768f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.64
cc_214 VPB N_SCE_c_570_n 0.0219533f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.64
cc_215 VPB N_SCE_c_571_n 0.0218634f $X=-0.19 $Y=1.66 $X2=0.407 $Y2=1.205
cc_216 VPB N_SCE_c_565_n 0.0226382f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.54
cc_217 VPB N_SCE_c_566_n 0.00271324f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_218 VPB N_SCE_c_574_n 0.0129976f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_219 VPB N_SCE_c_575_n 0.0372139f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_220 VPB SCE 0.00720768f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_221 VPB N_CLK_N_c_665_n 0.0354311f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.245
cc_222 VPB N_CLK_N_c_666_n 0.00413642f $X=-0.19 $Y=1.66 $X2=0.407 $Y2=1.875
cc_223 VPB N_A_977_243#_c_712_n 0.0165367f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_224 VPB N_A_977_243#_c_707_n 0.0461885f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_225 VPB N_A_977_243#_c_714_n 0.0166641f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_226 VPB N_A_977_243#_c_708_n 0.00525376f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_227 VPB N_A_977_243#_c_716_n 0.0398948f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_228 VPB N_A_977_243#_c_717_n 0.00569037f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_229 VPB N_A_977_243#_c_718_n 0.0030569f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_230 VPB N_A_977_243#_c_719_n 0.00247443f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_231 VPB N_A_977_243#_c_709_n 0.0025142f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_232 VPB N_A_977_243#_c_721_n 0.010787f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_233 VPB N_A_977_243#_c_710_n 0.0030028f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_234 VPB N_A_977_243#_c_723_n 0.0043973f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_235 VPB N_A_977_243#_c_724_n 0.0189072f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_236 VPB N_A_977_243#_c_725_n 0.0252002f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_237 VPB N_A_977_243#_c_726_n 0.0112772f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_238 VPB N_A_977_243#_c_727_n 0.0105943f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_239 VPB N_A_867_82#_c_922_n 0.0238948f $X=-0.19 $Y=1.66 $X2=0.52 $Y2=1.205
cc_240 VPB N_A_867_82#_c_923_n 0.0203105f $X=-0.19 $Y=1.66 $X2=0.52 $Y2=0.805
cc_241 VPB N_A_867_82#_c_904_n 0.0434226f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.37
cc_242 VPB N_A_867_82#_c_907_n 0.00765999f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_243 VPB N_A_867_82#_c_926_n 0.0140344f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_244 VPB N_A_867_82#_c_912_n 7.37857e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_245 VPB N_A_867_82#_c_913_n 0.0159834f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_246 VPB N_A_867_82#_c_914_n 0.00552797f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_247 VPB N_A_867_82#_c_915_n 0.0133672f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_248 VPB N_A_867_82#_c_916_n 0.00101238f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_249 VPB N_A_867_82#_c_917_n 5.82846e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_250 VPB N_A_867_82#_c_918_n 0.00274445f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_251 VPB N_A_867_82#_c_919_n 0.0232f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_252 VPB N_A_867_82#_c_920_n 0.00616144f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_253 VPB N_A_867_82#_c_921_n 0.00177136f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_254 VPB N_A_1159_497#_c_1126_n 0.0140425f $X=-0.19 $Y=1.66 $X2=0.52 $Y2=0.805
cc_255 VPB N_A_1159_497#_c_1134_n 0.0249579f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_256 VPB N_A_1159_497#_c_1135_n 0.0149639f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_257 VPB N_A_1159_497#_c_1136_n 0.00191448f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_258 VPB N_A_1159_497#_c_1132_n 0.0305631f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_259 VPB N_A_1159_497#_c_1138_n 0.00433033f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_260 VPB N_A_1579_258#_c_1221_n 0.016041f $X=-0.19 $Y=1.66 $X2=0.52 $Y2=1.205
cc_261 VPB N_A_1579_258#_c_1243_n 0.0209614f $X=-0.19 $Y=1.66 $X2=0.52 $Y2=0.805
cc_262 VPB N_A_1579_258#_c_1225_n 0.00795556f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_263 VPB N_A_1579_258#_c_1245_n 0.0235235f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_264 VPB N_A_1579_258#_c_1235_n 0.00628773f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_265 VPB N_A_1579_258#_c_1247_n 2.8453e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_266 VPB N_A_1579_258#_c_1248_n 0.00481227f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_267 VPB N_SET_B_c_1429_n 0.0181442f $X=-0.19 $Y=1.66 $X2=0.407 $Y2=1.392
cc_268 VPB N_SET_B_c_1424_n 0.038771f $X=-0.19 $Y=1.66 $X2=0.52 $Y2=1.205
cc_269 VPB N_SET_B_c_1431_n 0.0372704f $X=-0.19 $Y=1.66 $X2=0.407 $Y2=1.37
cc_270 VPB N_SET_B_c_1432_n 0.00255655f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.37
cc_271 VPB N_SET_B_c_1426_n 0.00864679f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=1.54
cc_272 VPB SET_B 5.17315e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_273 VPB N_SET_B_c_1427_n 0.0540421f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_274 VPB N_SET_B_c_1428_n 0.00297931f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_275 VPB N_A_662_82#_c_1559_n 0.0311895f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_276 VPB N_A_662_82#_c_1563_n 0.0229911f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_277 VPB N_A_662_82#_c_1576_n 0.0181314f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_278 VPB N_A_662_82#_c_1577_n 0.0343037f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_279 VPB N_A_662_82#_c_1578_n 0.0233331f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_280 VPB N_A_662_82#_c_1570_n 0.0315192f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_281 VPB N_A_662_82#_c_1580_n 0.00175877f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_282 VPB N_A_662_82#_c_1581_n 0.0102711f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_283 VPB N_A_662_82#_c_1582_n 0.00311108f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_284 VPB N_A_662_82#_c_1573_n 0.00104023f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_285 VPB N_A_2133_410#_c_1756_n 0.0550011f $X=-0.19 $Y=1.66 $X2=0.52 $Y2=0.805
cc_286 VPB N_A_2133_410#_c_1757_n 0.0259723f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_287 VPB N_A_2133_410#_M1010_g 0.0252797f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.37
cc_288 VPB N_A_2133_410#_c_1743_n 0.0385324f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=1.54
cc_289 VPB N_A_2133_410#_c_1745_n 0.0111245f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_290 VPB N_A_2133_410#_c_1746_n 0.00655454f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_291 VPB N_A_2133_410#_c_1762_n 0.0254045f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_292 VPB N_A_2133_410#_c_1763_n 0.00438288f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_293 VPB N_A_2133_410#_c_1764_n 0.00852783f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_294 VPB N_A_2133_410#_c_1765_n 0.00337273f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_295 VPB N_A_2133_410#_c_1766_n 0.00389272f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_296 VPB N_A_2133_410#_c_1767_n 0.0220235f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_297 VPB N_A_2133_410#_c_1768_n 0.00200072f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_298 VPB N_A_2133_410#_c_1769_n 0.00606369f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_299 VPB N_A_2133_410#_c_1770_n 0.0059083f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_300 VPB N_A_2133_410#_c_1754_n 0.00319302f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_301 VPB N_A_1954_119#_c_1977_n 0.0311806f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_302 VPB N_A_1954_119#_c_1984_n 0.00523752f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_303 VPB N_A_1954_119#_c_1985_n 0.00248991f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_304 VPB N_A_1954_119#_c_1986_n 0.0132221f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_305 VPB N_A_1954_119#_c_1987_n 0.00125324f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_306 VPB N_A_1954_119#_c_1979_n 0.00219863f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_307 VPB N_A_1954_119#_c_1989_n 0.00507504f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_308 VPB N_A_1954_119#_c_1990_n 0.0030807f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_309 VPB N_A_1954_119#_c_1991_n 0.00317473f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_310 VPB N_A_1954_119#_c_1992_n 0.00126464f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_311 VPB N_A_1954_119#_c_1980_n 0.00453832f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_312 VPB N_A_1954_119#_c_1981_n 0.00933214f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_313 VPB N_A_1954_119#_c_1982_n 0.0273115f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_314 VPB N_A_1954_119#_c_1996_n 0.00467045f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_315 VPB N_RESET_B_c_2124_n 0.0207148f $X=-0.19 $Y=1.66 $X2=0.407 $Y2=1.392
cc_316 VPB N_RESET_B_c_2125_n 0.0215196f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.64
cc_317 VPB N_RESET_B_c_2126_n 0.0119542f $X=-0.19 $Y=1.66 $X2=0.52 $Y2=1.205
cc_318 VPB N_RESET_B_c_2127_n 0.0284749f $X=-0.19 $Y=1.66 $X2=0.52 $Y2=0.805
cc_319 VPB RESET_B 0.00188312f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_320 VPB N_RESET_B_c_2123_n 0.0071132f $X=-0.19 $Y=1.66 $X2=0.407 $Y2=1.205
cc_321 VPB N_A_3078_384#_c_2175_n 0.0292569f $X=-0.19 $Y=1.66 $X2=0.52 $Y2=0.805
cc_322 VPB N_A_3078_384#_c_2177_n 0.00519655f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=1.54
cc_323 VPB N_A_27_464#_c_2226_n 0.0323906f $X=-0.19 $Y=1.66 $X2=0.52 $Y2=0.805
cc_324 VPB N_A_27_464#_c_2227_n 0.0138099f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_325 VPB N_A_27_464#_c_2228_n 0.0100121f $X=-0.19 $Y=1.66 $X2=0.407 $Y2=1.875
cc_326 VPB N_A_27_464#_c_2229_n 0.00136174f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_327 VPB N_A_27_464#_c_2230_n 0.00711585f $X=-0.19 $Y=1.66 $X2=0.407 $Y2=1.37
cc_328 VPB N_A_27_464#_c_2231_n 0.00226853f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.37
cc_329 VPB N_A_27_464#_c_2232_n 0.00739969f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=1.54
cc_330 VPB N_VPWR_c_2277_n 0.00619043f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_331 VPB N_VPWR_c_2278_n 0.0178548f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_332 VPB N_VPWR_c_2279_n 0.00571271f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_333 VPB N_VPWR_c_2280_n 0.0235577f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_334 VPB N_VPWR_c_2281_n 0.00953088f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_335 VPB N_VPWR_c_2282_n 0.00806851f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_336 VPB N_VPWR_c_2283_n 0.0115529f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_337 VPB N_VPWR_c_2284_n 0.00713932f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_338 VPB N_VPWR_c_2285_n 0.0147501f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_339 VPB N_VPWR_c_2286_n 0.0688573f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_340 VPB N_VPWR_c_2287_n 0.00324402f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_341 VPB N_VPWR_c_2288_n 0.0144232f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_342 VPB N_VPWR_c_2289_n 0.0443291f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_343 VPB N_VPWR_c_2290_n 0.0341433f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_344 VPB N_VPWR_c_2291_n 0.0047828f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_345 VPB N_VPWR_c_2292_n 0.017793f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_346 VPB N_VPWR_c_2293_n 0.0386695f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_347 VPB N_VPWR_c_2294_n 0.033549f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_348 VPB N_VPWR_c_2295_n 0.0213606f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_349 VPB N_VPWR_c_2296_n 0.0196646f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_350 VPB N_VPWR_c_2297_n 0.0473883f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_351 VPB N_VPWR_c_2298_n 0.0198718f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_352 VPB N_VPWR_c_2276_n 0.223377f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_353 VPB N_VPWR_c_2300_n 0.00614127f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_354 VPB N_VPWR_c_2301_n 0.0047828f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_355 VPB N_VPWR_c_2302_n 0.00460249f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_356 VPB N_VPWR_c_2303_n 0.0047828f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_357 VPB N_VPWR_c_2304_n 0.00614127f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_358 VPB N_VPWR_c_2305_n 0.0139421f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_359 VPB N_VPWR_c_2306_n 0.0128855f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_360 VPB N_A_197_119#_c_2489_n 8.66286e-19 $X=-0.19 $Y=1.66 $X2=0.407 $Y2=1.37
cc_361 VPB N_A_197_119#_c_2490_n 0.00484755f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_362 VPB N_A_197_119#_c_2491_n 0.00267979f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_363 VPB N_A_197_119#_c_2469_n 0.00299681f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_364 VPB N_A_197_119#_c_2493_n 0.00874139f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_365 VPB N_A_197_119#_c_2486_n 0.00318629f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_366 VPB N_A_197_119#_c_2495_n 0.00239124f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_367 VPB N_A_197_119#_c_2496_n 0.00834522f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_368 VPB Q_N 0.00504742f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_369 VPB Q_N 0.0171996f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_370 VPB N_Q_N_c_2703_n 0.00365979f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_371 VPB Q 0.0137079f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_372 VPB Q 0.041687f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_373 VPB N_Q_c_2738_n 0.00777552f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_374 N_SCD_M1004_g N_SCE_M1033_g 0.0380401f $X=0.52 $Y=0.805 $X2=0 $Y2=0
cc_375 N_SCD_c_380_n N_SCE_c_569_n 0.00823444f $X=0.505 $Y=2.155 $X2=0 $Y2=0
cc_376 N_SCD_c_381_n N_SCE_c_570_n 0.0149333f $X=0.505 $Y=2.245 $X2=0 $Y2=0
cc_377 N_SCD_c_375_n N_SCE_c_566_n 0.0141465f $X=0.407 $Y=1.688 $X2=0 $Y2=0
cc_378 N_SCD_c_382_n N_SCE_c_574_n 0.0141465f $X=0.407 $Y=1.875 $X2=0 $Y2=0
cc_379 N_SCD_c_377_n SCE 0.0024538f $X=0.385 $Y=1.37 $X2=0 $Y2=0
cc_380 N_SCD_c_378_n SCE 0.0383728f $X=0.385 $Y=1.37 $X2=0 $Y2=0
cc_381 N_SCD_c_377_n N_SCE_c_568_n 0.0141465f $X=0.385 $Y=1.37 $X2=0 $Y2=0
cc_382 N_SCD_c_378_n N_SCE_c_568_n 7.83271e-19 $X=0.385 $Y=1.37 $X2=0 $Y2=0
cc_383 N_SCD_c_381_n N_A_27_464#_c_2226_n 0.00359266f $X=0.505 $Y=2.245 $X2=0
+ $Y2=0
cc_384 N_SCD_c_380_n N_A_27_464#_c_2227_n 0.00918054f $X=0.505 $Y=2.155 $X2=0
+ $Y2=0
cc_385 N_SCD_c_381_n N_A_27_464#_c_2227_n 0.00976364f $X=0.505 $Y=2.245 $X2=0
+ $Y2=0
cc_386 N_SCD_c_382_n N_A_27_464#_c_2227_n 5.17145e-19 $X=0.407 $Y=1.875 $X2=0
+ $Y2=0
cc_387 N_SCD_c_378_n N_A_27_464#_c_2227_n 0.011771f $X=0.385 $Y=1.37 $X2=0 $Y2=0
cc_388 N_SCD_c_382_n N_A_27_464#_c_2228_n 0.00469803f $X=0.407 $Y=1.875 $X2=0
+ $Y2=0
cc_389 N_SCD_c_378_n N_A_27_464#_c_2228_n 0.0243647f $X=0.385 $Y=1.37 $X2=0
+ $Y2=0
cc_390 N_SCD_c_381_n N_VPWR_c_2277_n 0.0124996f $X=0.505 $Y=2.245 $X2=0 $Y2=0
cc_391 N_SCD_c_381_n N_VPWR_c_2292_n 0.00413917f $X=0.505 $Y=2.245 $X2=0 $Y2=0
cc_392 N_SCD_c_381_n N_VPWR_c_2276_n 0.00821221f $X=0.505 $Y=2.245 $X2=0 $Y2=0
cc_393 N_SCD_M1004_g N_A_197_119#_c_2487_n 0.00130204f $X=0.52 $Y=0.805 $X2=0
+ $Y2=0
cc_394 N_SCD_M1004_g N_VGND_c_2760_n 0.0141223f $X=0.52 $Y=0.805 $X2=0 $Y2=0
cc_395 N_SCD_c_377_n N_VGND_c_2760_n 0.00605214f $X=0.385 $Y=1.37 $X2=0 $Y2=0
cc_396 N_SCD_c_378_n N_VGND_c_2760_n 0.0293252f $X=0.385 $Y=1.37 $X2=0 $Y2=0
cc_397 N_SCD_M1004_g N_VGND_c_2770_n 0.0035863f $X=0.52 $Y=0.805 $X2=0 $Y2=0
cc_398 N_SCD_M1004_g N_VGND_c_2776_n 0.00401353f $X=0.52 $Y=0.805 $X2=0 $Y2=0
cc_399 N_D_M1000_g N_A_353_93#_c_469_n 0.0394323f $X=1.45 $Y=0.805 $X2=0 $Y2=0
cc_400 N_D_c_413_n N_A_353_93#_c_476_n 0.0176124f $X=1.412 $Y=2.245 $X2=0 $Y2=0
cc_401 N_D_M1000_g N_A_353_93#_c_470_n 0.00253719f $X=1.45 $Y=0.805 $X2=0 $Y2=0
cc_402 N_D_c_412_n N_A_353_93#_c_477_n 0.00233085f $X=1.412 $Y=2.115 $X2=0 $Y2=0
cc_403 N_D_c_411_n N_A_353_93#_c_471_n 0.00264551f $X=1.65 $Y=1.645 $X2=0 $Y2=0
cc_404 N_D_c_412_n N_A_353_93#_c_478_n 0.0079207f $X=1.412 $Y=2.115 $X2=0 $Y2=0
cc_405 N_D_c_411_n N_A_353_93#_c_478_n 0.00263996f $X=1.65 $Y=1.645 $X2=0 $Y2=0
cc_406 D N_A_353_93#_c_472_n 3.59433e-19 $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_407 N_D_c_411_n N_A_353_93#_c_472_n 0.0182717f $X=1.65 $Y=1.645 $X2=0 $Y2=0
cc_408 N_D_M1000_g N_SCE_M1033_g 0.0161922f $X=1.45 $Y=0.805 $X2=0 $Y2=0
cc_409 N_D_c_412_n N_SCE_c_569_n 0.0116633f $X=1.412 $Y=2.115 $X2=0 $Y2=0
cc_410 N_D_c_413_n N_SCE_c_569_n 0.00592068f $X=1.412 $Y=2.245 $X2=0 $Y2=0
cc_411 N_D_c_413_n N_SCE_c_570_n 0.0321632f $X=1.412 $Y=2.245 $X2=0 $Y2=0
cc_412 N_D_M1000_g N_SCE_c_560_n 0.0100779f $X=1.45 $Y=0.805 $X2=0 $Y2=0
cc_413 D N_SCE_c_566_n 2.37847e-19 $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_414 N_D_c_411_n N_SCE_c_566_n 0.0123129f $X=1.65 $Y=1.645 $X2=0 $Y2=0
cc_415 N_D_c_412_n N_SCE_c_574_n 0.0123129f $X=1.412 $Y=2.115 $X2=0 $Y2=0
cc_416 N_D_M1000_g SCE 0.00327536f $X=1.45 $Y=0.805 $X2=0 $Y2=0
cc_417 D SCE 0.0271418f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_418 N_D_c_411_n SCE 0.00370314f $X=1.65 $Y=1.645 $X2=0 $Y2=0
cc_419 N_D_M1000_g N_SCE_c_568_n 0.013498f $X=1.45 $Y=0.805 $X2=0 $Y2=0
cc_420 N_D_c_412_n N_A_27_464#_c_2227_n 6.64604e-19 $X=1.412 $Y=2.115 $X2=0
+ $Y2=0
cc_421 N_D_c_413_n N_A_27_464#_c_2227_n 9.74204e-19 $X=1.412 $Y=2.245 $X2=0
+ $Y2=0
cc_422 N_D_c_413_n N_A_27_464#_c_2229_n 0.00759296f $X=1.412 $Y=2.245 $X2=0
+ $Y2=0
cc_423 N_D_c_413_n N_A_27_464#_c_2230_n 0.0130117f $X=1.412 $Y=2.245 $X2=0 $Y2=0
cc_424 N_D_c_413_n N_A_27_464#_c_2232_n 9.41798e-19 $X=1.412 $Y=2.245 $X2=0
+ $Y2=0
cc_425 N_D_c_413_n N_VPWR_c_2293_n 0.00278271f $X=1.412 $Y=2.245 $X2=0 $Y2=0
cc_426 N_D_c_413_n N_VPWR_c_2276_n 0.00353713f $X=1.412 $Y=2.245 $X2=0 $Y2=0
cc_427 N_D_M1000_g N_A_197_119#_c_2467_n 0.010538f $X=1.45 $Y=0.805 $X2=0 $Y2=0
cc_428 N_D_c_411_n N_A_197_119#_c_2467_n 9.31825e-19 $X=1.65 $Y=1.645 $X2=0
+ $Y2=0
cc_429 N_D_c_413_n N_A_197_119#_c_2489_n 0.00284379f $X=1.412 $Y=2.245 $X2=0
+ $Y2=0
cc_430 D N_A_197_119#_c_2489_n 0.00220458f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_431 N_D_c_411_n N_A_197_119#_c_2489_n 0.00100464f $X=1.65 $Y=1.645 $X2=0
+ $Y2=0
cc_432 N_D_c_413_n N_A_197_119#_c_2503_n 0.00377073f $X=1.412 $Y=2.245 $X2=0
+ $Y2=0
cc_433 N_D_M1000_g N_A_197_119#_c_2468_n 5.06211e-19 $X=1.45 $Y=0.805 $X2=0
+ $Y2=0
cc_434 D N_A_197_119#_c_2468_n 0.0120251f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_435 N_D_c_411_n N_A_197_119#_c_2468_n 0.00274991f $X=1.65 $Y=1.645 $X2=0
+ $Y2=0
cc_436 D N_A_197_119#_c_2490_n 0.00747803f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_437 N_D_c_411_n N_A_197_119#_c_2490_n 0.00140249f $X=1.65 $Y=1.645 $X2=0
+ $Y2=0
cc_438 N_D_c_412_n N_A_197_119#_c_2491_n 0.00416101f $X=1.412 $Y=2.115 $X2=0
+ $Y2=0
cc_439 D N_A_197_119#_c_2491_n 0.0143367f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_440 N_D_c_411_n N_A_197_119#_c_2491_n 0.00396026f $X=1.65 $Y=1.645 $X2=0
+ $Y2=0
cc_441 N_D_M1000_g N_A_197_119#_c_2469_n 0.00149161f $X=1.45 $Y=0.805 $X2=0
+ $Y2=0
cc_442 N_D_c_412_n N_A_197_119#_c_2469_n 0.00231823f $X=1.412 $Y=2.115 $X2=0
+ $Y2=0
cc_443 D N_A_197_119#_c_2469_n 0.0247729f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_444 N_D_c_411_n N_A_197_119#_c_2469_n 9.87882e-19 $X=1.65 $Y=1.645 $X2=0
+ $Y2=0
cc_445 N_D_M1000_g N_A_197_119#_c_2487_n 0.00447624f $X=1.45 $Y=0.805 $X2=0
+ $Y2=0
cc_446 N_D_c_413_n N_A_197_119#_c_2495_n 0.00133756f $X=1.412 $Y=2.245 $X2=0
+ $Y2=0
cc_447 N_D_M1000_g N_A_197_119#_c_2488_n 0.010065f $X=1.45 $Y=0.805 $X2=0 $Y2=0
cc_448 D N_A_197_119#_c_2488_n 0.013518f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_449 N_D_c_411_n N_A_197_119#_c_2488_n 0.00296428f $X=1.65 $Y=1.645 $X2=0
+ $Y2=0
cc_450 N_D_M1000_g N_VGND_c_2761_n 0.00150032f $X=1.45 $Y=0.805 $X2=0 $Y2=0
cc_451 N_D_M1000_g N_VGND_c_2776_n 9.39239e-19 $X=1.45 $Y=0.805 $X2=0 $Y2=0
cc_452 N_A_353_93#_c_469_n N_SCE_c_560_n 0.0103107f $X=1.84 $Y=1.09 $X2=0 $Y2=0
cc_453 N_A_353_93#_c_469_n N_SCE_M1018_g 0.00391183f $X=1.84 $Y=1.09 $X2=0 $Y2=0
cc_454 N_A_353_93#_c_473_n N_SCE_M1018_g 0.00771436f $X=2.895 $Y=0.815 $X2=0
+ $Y2=0
cc_455 N_A_353_93#_c_473_n N_SCE_c_563_n 0.0182689f $X=2.895 $Y=0.815 $X2=0
+ $Y2=0
cc_456 N_A_353_93#_c_475_n N_SCE_c_563_n 8.83272e-19 $X=2.975 $Y=1.645 $X2=0
+ $Y2=0
cc_457 N_A_353_93#_c_471_n N_SCE_c_564_n 0.0039383f $X=2.13 $Y=1.165 $X2=0 $Y2=0
cc_458 N_A_353_93#_c_473_n N_SCE_c_564_n 0.00179726f $X=2.895 $Y=0.815 $X2=0
+ $Y2=0
cc_459 N_A_353_93#_c_474_n N_SCE_c_564_n 0.01377f $X=2.675 $Y=1.645 $X2=0 $Y2=0
cc_460 N_A_353_93#_c_475_n N_SCE_c_564_n 0.00102404f $X=2.975 $Y=1.645 $X2=0
+ $Y2=0
cc_461 N_A_353_93#_c_482_n N_SCE_c_571_n 0.00936672f $X=3.085 $Y=2.465 $X2=0
+ $Y2=0
cc_462 N_A_353_93#_c_483_n N_SCE_c_571_n 0.00311577f $X=3.07 $Y=2.3 $X2=0 $Y2=0
cc_463 N_A_353_93#_c_473_n N_SCE_c_565_n 0.00443983f $X=2.895 $Y=0.815 $X2=0
+ $Y2=0
cc_464 N_A_353_93#_c_474_n N_SCE_c_565_n 0.0163192f $X=2.675 $Y=1.645 $X2=0
+ $Y2=0
cc_465 N_A_353_93#_c_475_n N_SCE_c_565_n 0.00460554f $X=2.975 $Y=1.645 $X2=0
+ $Y2=0
cc_466 N_A_353_93#_c_483_n N_SCE_c_565_n 0.00591239f $X=3.07 $Y=2.3 $X2=0 $Y2=0
cc_467 N_A_353_93#_c_478_n N_SCE_c_575_n 0.00334442f $X=1.855 $Y=2.147 $X2=0
+ $Y2=0
cc_468 N_A_353_93#_c_474_n N_SCE_c_575_n 0.00426361f $X=2.675 $Y=1.645 $X2=0
+ $Y2=0
cc_469 N_A_353_93#_c_475_n N_SCE_c_575_n 0.0032851f $X=2.975 $Y=1.645 $X2=0
+ $Y2=0
cc_470 N_A_353_93#_c_482_n N_SCE_c_575_n 0.00866124f $X=3.085 $Y=2.465 $X2=0
+ $Y2=0
cc_471 N_A_353_93#_c_483_n N_SCE_c_575_n 0.0164719f $X=3.07 $Y=2.3 $X2=0 $Y2=0
cc_472 N_A_353_93#_c_473_n N_CLK_N_M1015_g 0.00542055f $X=2.895 $Y=0.815 $X2=0
+ $Y2=0
cc_473 N_A_353_93#_c_473_n N_CLK_N_c_666_n 0.00532473f $X=2.895 $Y=0.815 $X2=0
+ $Y2=0
cc_474 N_A_353_93#_c_475_n N_CLK_N_c_666_n 0.0132306f $X=2.975 $Y=1.645 $X2=0
+ $Y2=0
cc_475 N_A_353_93#_c_473_n N_A_662_82#_c_1571_n 0.0174028f $X=2.895 $Y=0.815
+ $X2=0 $Y2=0
cc_476 N_A_353_93#_c_483_n N_A_662_82#_c_1580_n 0.00736629f $X=3.07 $Y=2.3 $X2=0
+ $Y2=0
cc_477 N_A_353_93#_c_482_n N_A_662_82#_c_1581_n 0.0451706f $X=3.085 $Y=2.465
+ $X2=0 $Y2=0
cc_478 N_A_353_93#_c_483_n N_A_662_82#_c_1581_n 0.00712165f $X=3.07 $Y=2.3 $X2=0
+ $Y2=0
cc_479 N_A_353_93#_c_476_n N_A_27_464#_c_2230_n 0.0134197f $X=1.855 $Y=2.245
+ $X2=0 $Y2=0
cc_480 N_A_353_93#_c_476_n N_A_27_464#_c_2232_n 0.00741093f $X=1.855 $Y=2.245
+ $X2=0 $Y2=0
cc_481 N_A_353_93#_c_478_n N_A_27_464#_c_2232_n 0.00763601f $X=1.855 $Y=2.147
+ $X2=0 $Y2=0
cc_482 N_A_353_93#_c_474_n N_A_27_464#_c_2232_n 0.00119962f $X=2.675 $Y=1.645
+ $X2=0 $Y2=0
cc_483 N_A_353_93#_c_476_n N_VPWR_c_2278_n 0.00223475f $X=1.855 $Y=2.245 $X2=0
+ $Y2=0
cc_484 N_A_353_93#_c_474_n N_VPWR_c_2278_n 0.00518466f $X=2.675 $Y=1.645 $X2=0
+ $Y2=0
cc_485 N_A_353_93#_c_475_n N_VPWR_c_2278_n 0.0079892f $X=2.975 $Y=1.645 $X2=0
+ $Y2=0
cc_486 N_A_353_93#_c_482_n N_VPWR_c_2278_n 0.0520379f $X=3.085 $Y=2.465 $X2=0
+ $Y2=0
cc_487 N_A_353_93#_c_476_n N_VPWR_c_2293_n 0.00278257f $X=1.855 $Y=2.245 $X2=0
+ $Y2=0
cc_488 N_A_353_93#_c_482_n N_VPWR_c_2294_n 0.0158428f $X=3.085 $Y=2.465 $X2=0
+ $Y2=0
cc_489 N_A_353_93#_c_476_n N_VPWR_c_2276_n 0.00358707f $X=1.855 $Y=2.245 $X2=0
+ $Y2=0
cc_490 N_A_353_93#_c_482_n N_VPWR_c_2276_n 0.0130099f $X=3.085 $Y=2.465 $X2=0
+ $Y2=0
cc_491 N_A_353_93#_c_471_n N_A_197_119#_c_2468_n 0.0115758f $X=2.13 $Y=1.165
+ $X2=0 $Y2=0
cc_492 N_A_353_93#_c_477_n N_A_197_119#_c_2490_n 0.00362853f $X=2.13 $Y=2.05
+ $X2=0 $Y2=0
cc_493 N_A_353_93#_c_478_n N_A_197_119#_c_2490_n 0.0192477f $X=1.855 $Y=2.147
+ $X2=0 $Y2=0
cc_494 N_A_353_93#_c_470_n N_A_197_119#_c_2469_n 0.00576352f $X=2.13 $Y=1.48
+ $X2=0 $Y2=0
cc_495 N_A_353_93#_c_477_n N_A_197_119#_c_2469_n 0.00932408f $X=2.13 $Y=2.05
+ $X2=0 $Y2=0
cc_496 N_A_353_93#_c_472_n N_A_197_119#_c_2469_n 0.0111597f $X=2.13 $Y=1.645
+ $X2=0 $Y2=0
cc_497 N_A_353_93#_c_473_n N_A_197_119#_c_2469_n 0.00511938f $X=2.895 $Y=0.815
+ $X2=0 $Y2=0
cc_498 N_A_353_93#_c_475_n N_A_197_119#_c_2469_n 0.0135626f $X=2.975 $Y=1.645
+ $X2=0 $Y2=0
cc_499 N_A_353_93#_c_470_n N_A_197_119#_c_2470_n 0.00390368f $X=2.13 $Y=1.48
+ $X2=0 $Y2=0
cc_500 N_A_353_93#_c_471_n N_A_197_119#_c_2470_n 0.00212655f $X=2.13 $Y=1.165
+ $X2=0 $Y2=0
cc_501 N_A_353_93#_c_473_n N_A_197_119#_c_2470_n 0.0146243f $X=2.895 $Y=0.815
+ $X2=0 $Y2=0
cc_502 N_A_353_93#_c_474_n N_A_197_119#_c_2470_n 0.0134099f $X=2.675 $Y=1.645
+ $X2=0 $Y2=0
cc_503 N_A_353_93#_c_475_n N_A_197_119#_c_2470_n 0.00421666f $X=2.975 $Y=1.645
+ $X2=0 $Y2=0
cc_504 N_A_353_93#_c_469_n N_A_197_119#_c_2471_n 0.00274962f $X=1.84 $Y=1.09
+ $X2=0 $Y2=0
cc_505 N_A_353_93#_c_471_n N_A_197_119#_c_2471_n 0.00111927f $X=2.13 $Y=1.165
+ $X2=0 $Y2=0
cc_506 N_A_353_93#_c_473_n N_A_197_119#_c_2471_n 0.0250399f $X=2.895 $Y=0.815
+ $X2=0 $Y2=0
cc_507 N_A_353_93#_c_473_n N_A_197_119#_c_2472_n 0.0230235f $X=2.895 $Y=0.815
+ $X2=0 $Y2=0
cc_508 N_A_353_93#_c_473_n N_A_197_119#_c_2476_n 0.0137113f $X=2.895 $Y=0.815
+ $X2=0 $Y2=0
cc_509 N_A_353_93#_c_469_n N_A_197_119#_c_2487_n 4.8292e-19 $X=1.84 $Y=1.09
+ $X2=0 $Y2=0
cc_510 N_A_353_93#_c_476_n N_A_197_119#_c_2495_n 0.0033357f $X=1.855 $Y=2.245
+ $X2=0 $Y2=0
cc_511 N_A_353_93#_c_478_n N_A_197_119#_c_2495_n 0.00231432f $X=1.855 $Y=2.147
+ $X2=0 $Y2=0
cc_512 N_A_353_93#_c_469_n N_A_197_119#_c_2488_n 0.00446134f $X=1.84 $Y=1.09
+ $X2=0 $Y2=0
cc_513 N_A_353_93#_c_470_n N_A_197_119#_c_2543_n 6.49734e-19 $X=2.13 $Y=1.48
+ $X2=0 $Y2=0
cc_514 N_A_353_93#_c_471_n N_A_197_119#_c_2543_n 0.00435912f $X=2.13 $Y=1.165
+ $X2=0 $Y2=0
cc_515 N_A_353_93#_c_469_n N_VGND_c_2761_n 0.0112979f $X=1.84 $Y=1.09 $X2=0
+ $Y2=0
cc_516 N_A_353_93#_c_471_n N_VGND_c_2761_n 0.00711376f $X=2.13 $Y=1.165 $X2=0
+ $Y2=0
cc_517 N_A_353_93#_c_469_n N_VGND_c_2776_n 7.88961e-19 $X=1.84 $Y=1.09 $X2=0
+ $Y2=0
cc_518 N_SCE_c_563_n N_CLK_N_M1015_g 0.00859889f $X=3.08 $Y=1.165 $X2=0 $Y2=0
cc_519 N_SCE_c_565_n N_CLK_N_c_665_n 0.024867f $X=3.155 $Y=2.05 $X2=0 $Y2=0
cc_520 N_SCE_c_565_n N_CLK_N_c_666_n 0.00219301f $X=3.155 $Y=2.05 $X2=0 $Y2=0
cc_521 N_SCE_M1018_g N_A_662_82#_c_1571_n 5.23339e-19 $X=2.68 $Y=0.805 $X2=0
+ $Y2=0
cc_522 N_SCE_c_563_n N_A_662_82#_c_1571_n 9.71613e-19 $X=3.08 $Y=1.165 $X2=0
+ $Y2=0
cc_523 N_SCE_c_565_n N_A_662_82#_c_1580_n 0.00217384f $X=3.155 $Y=2.05 $X2=0
+ $Y2=0
cc_524 N_SCE_c_571_n N_A_662_82#_c_1581_n 0.00145252f $X=2.86 $Y=2.245 $X2=0
+ $Y2=0
cc_525 N_SCE_c_575_n N_A_662_82#_c_1581_n 0.0011314f $X=2.86 $Y=2.147 $X2=0
+ $Y2=0
cc_526 N_SCE_c_569_n N_A_27_464#_c_2227_n 0.00638477f $X=0.985 $Y=2.155 $X2=0
+ $Y2=0
cc_527 N_SCE_c_570_n N_A_27_464#_c_2227_n 0.00933743f $X=0.985 $Y=2.245 $X2=0
+ $Y2=0
cc_528 N_SCE_c_574_n N_A_27_464#_c_2227_n 0.00397139f $X=0.97 $Y=1.875 $X2=0
+ $Y2=0
cc_529 SCE N_A_27_464#_c_2227_n 0.0354635f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_530 N_SCE_c_570_n N_A_27_464#_c_2229_n 0.00469834f $X=0.985 $Y=2.245 $X2=0
+ $Y2=0
cc_531 N_SCE_c_570_n N_A_27_464#_c_2231_n 0.00126137f $X=0.985 $Y=2.245 $X2=0
+ $Y2=0
cc_532 N_SCE_c_570_n N_VPWR_c_2277_n 0.00141926f $X=0.985 $Y=2.245 $X2=0 $Y2=0
cc_533 N_SCE_c_571_n N_VPWR_c_2278_n 0.00716702f $X=2.86 $Y=2.245 $X2=0 $Y2=0
cc_534 N_SCE_c_570_n N_VPWR_c_2293_n 0.00461464f $X=0.985 $Y=2.245 $X2=0 $Y2=0
cc_535 N_SCE_c_571_n N_VPWR_c_2294_n 0.00411612f $X=2.86 $Y=2.245 $X2=0 $Y2=0
cc_536 N_SCE_c_570_n N_VPWR_c_2276_n 0.00907984f $X=0.985 $Y=2.245 $X2=0 $Y2=0
cc_537 N_SCE_c_571_n N_VPWR_c_2276_n 0.00757132f $X=2.86 $Y=2.245 $X2=0 $Y2=0
cc_538 N_SCE_c_560_n N_A_197_119#_c_2467_n 0.00155845f $X=2.605 $Y=0.18 $X2=0
+ $Y2=0
cc_539 SCE N_A_197_119#_c_2467_n 0.00209962f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_540 N_SCE_c_575_n N_A_197_119#_c_2490_n 5.52612e-19 $X=2.86 $Y=2.147 $X2=0
+ $Y2=0
cc_541 SCE N_A_197_119#_c_2469_n 0.00733237f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_542 N_SCE_c_564_n N_A_197_119#_c_2470_n 0.00120369f $X=2.755 $Y=1.165 $X2=0
+ $Y2=0
cc_543 N_SCE_M1018_g N_A_197_119#_c_2471_n 0.00860995f $X=2.68 $Y=0.805 $X2=0
+ $Y2=0
cc_544 N_SCE_M1018_g N_A_197_119#_c_2472_n 0.0166548f $X=2.68 $Y=0.805 $X2=0
+ $Y2=0
cc_545 N_SCE_c_563_n N_A_197_119#_c_2472_n 0.00496066f $X=3.08 $Y=1.165 $X2=0
+ $Y2=0
cc_546 N_SCE_c_560_n N_A_197_119#_c_2473_n 0.00446747f $X=2.605 $Y=0.18 $X2=0
+ $Y2=0
cc_547 N_SCE_M1018_g N_A_197_119#_c_2474_n 0.00254464f $X=2.68 $Y=0.805 $X2=0
+ $Y2=0
cc_548 N_SCE_M1018_g N_A_197_119#_c_2476_n 6.01013e-19 $X=2.68 $Y=0.805 $X2=0
+ $Y2=0
cc_549 N_SCE_M1033_g N_A_197_119#_c_2487_n 0.00936054f $X=0.91 $Y=0.805 $X2=0
+ $Y2=0
cc_550 N_SCE_c_560_n N_A_197_119#_c_2487_n 0.00422441f $X=2.605 $Y=0.18 $X2=0
+ $Y2=0
cc_551 SCE N_A_197_119#_c_2487_n 0.0287978f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_552 N_SCE_c_568_n N_A_197_119#_c_2487_n 0.00401793f $X=0.97 $Y=1.37 $X2=0
+ $Y2=0
cc_553 N_SCE_M1033_g N_A_197_119#_c_2488_n 8.13451e-19 $X=0.91 $Y=0.805 $X2=0
+ $Y2=0
cc_554 N_SCE_c_560_n N_A_197_119#_c_2488_n 0.00249063f $X=2.605 $Y=0.18 $X2=0
+ $Y2=0
cc_555 SCE N_A_197_119#_c_2488_n 0.00818462f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_556 N_SCE_M1033_g N_VGND_c_2760_n 0.0018473f $X=0.91 $Y=0.805 $X2=0 $Y2=0
cc_557 N_SCE_c_561_n N_VGND_c_2760_n 0.00977077f $X=0.985 $Y=0.18 $X2=0 $Y2=0
cc_558 N_SCE_c_560_n N_VGND_c_2761_n 0.0255808f $X=2.605 $Y=0.18 $X2=0 $Y2=0
cc_559 N_SCE_M1018_g N_VGND_c_2761_n 0.00171036f $X=2.68 $Y=0.805 $X2=0 $Y2=0
cc_560 N_SCE_c_561_n N_VGND_c_2770_n 0.0343879f $X=0.985 $Y=0.18 $X2=0 $Y2=0
cc_561 N_SCE_c_560_n N_VGND_c_2771_n 0.0142019f $X=2.605 $Y=0.18 $X2=0 $Y2=0
cc_562 N_SCE_c_560_n N_VGND_c_2776_n 0.0514593f $X=2.605 $Y=0.18 $X2=0 $Y2=0
cc_563 N_SCE_c_561_n N_VGND_c_2776_n 0.0107881f $X=0.985 $Y=0.18 $X2=0 $Y2=0
cc_564 N_CLK_N_c_665_n N_A_867_82#_c_926_n 7.34107e-19 $X=3.87 $Y=1.765 $X2=0
+ $Y2=0
cc_565 N_CLK_N_M1015_g N_A_662_82#_M1016_g 0.0261259f $X=3.67 $Y=0.78 $X2=0
+ $Y2=0
cc_566 N_CLK_N_M1015_g N_A_662_82#_c_1559_n 2.31546e-19 $X=3.67 $Y=0.78 $X2=0
+ $Y2=0
cc_567 N_CLK_N_c_665_n N_A_662_82#_c_1559_n 0.0461231f $X=3.87 $Y=1.765 $X2=0
+ $Y2=0
cc_568 N_CLK_N_c_666_n N_A_662_82#_c_1559_n 2.18753e-19 $X=3.635 $Y=1.515 $X2=0
+ $Y2=0
cc_569 N_CLK_N_M1015_g N_A_662_82#_c_1571_n 0.0116247f $X=3.67 $Y=0.78 $X2=0
+ $Y2=0
cc_570 N_CLK_N_c_665_n N_A_662_82#_c_1571_n 0.0081008f $X=3.87 $Y=1.765 $X2=0
+ $Y2=0
cc_571 N_CLK_N_c_666_n N_A_662_82#_c_1571_n 0.0243296f $X=3.635 $Y=1.515 $X2=0
+ $Y2=0
cc_572 N_CLK_N_c_665_n N_A_662_82#_c_1580_n 0.00152805f $X=3.87 $Y=1.765 $X2=0
+ $Y2=0
cc_573 N_CLK_N_c_666_n N_A_662_82#_c_1580_n 0.0222375f $X=3.635 $Y=1.515 $X2=0
+ $Y2=0
cc_574 N_CLK_N_c_665_n N_A_662_82#_c_1581_n 0.0043207f $X=3.87 $Y=1.765 $X2=0
+ $Y2=0
cc_575 N_CLK_N_c_665_n N_A_662_82#_c_1603_n 0.016278f $X=3.87 $Y=1.765 $X2=0
+ $Y2=0
cc_576 N_CLK_N_c_666_n N_A_662_82#_c_1603_n 0.00334513f $X=3.635 $Y=1.515 $X2=0
+ $Y2=0
cc_577 N_CLK_N_M1015_g N_A_662_82#_c_1572_n 0.00351998f $X=3.67 $Y=0.78 $X2=0
+ $Y2=0
cc_578 N_CLK_N_c_665_n N_A_662_82#_c_1582_n 0.0028652f $X=3.87 $Y=1.765 $X2=0
+ $Y2=0
cc_579 N_CLK_N_c_666_n N_A_662_82#_c_1582_n 0.00822842f $X=3.635 $Y=1.515 $X2=0
+ $Y2=0
cc_580 N_CLK_N_M1015_g N_A_662_82#_c_1573_n 2.20897e-19 $X=3.67 $Y=0.78 $X2=0
+ $Y2=0
cc_581 N_CLK_N_c_665_n N_A_662_82#_c_1573_n 0.00272959f $X=3.87 $Y=1.765 $X2=0
+ $Y2=0
cc_582 N_CLK_N_c_666_n N_A_662_82#_c_1573_n 0.0260944f $X=3.635 $Y=1.515 $X2=0
+ $Y2=0
cc_583 N_CLK_N_c_665_n N_VPWR_c_2279_n 0.0135832f $X=3.87 $Y=1.765 $X2=0 $Y2=0
cc_584 N_CLK_N_c_665_n N_VPWR_c_2294_n 0.00413917f $X=3.87 $Y=1.765 $X2=0 $Y2=0
cc_585 N_CLK_N_c_665_n N_VPWR_c_2276_n 0.00822528f $X=3.87 $Y=1.765 $X2=0 $Y2=0
cc_586 N_CLK_N_M1015_g N_A_197_119#_c_2472_n 0.00355259f $X=3.67 $Y=0.78 $X2=0
+ $Y2=0
cc_587 N_CLK_N_M1015_g N_A_197_119#_c_2474_n 0.00513179f $X=3.67 $Y=0.78 $X2=0
+ $Y2=0
cc_588 N_CLK_N_M1015_g N_A_197_119#_c_2475_n 0.0135552f $X=3.67 $Y=0.78 $X2=0
+ $Y2=0
cc_589 N_CLK_N_M1015_g N_VGND_c_2771_n 0.00414982f $X=3.67 $Y=0.78 $X2=0 $Y2=0
cc_590 N_CLK_N_M1015_g N_VGND_c_2776_n 0.00533081f $X=3.67 $Y=0.78 $X2=0 $Y2=0
cc_591 N_CLK_N_M1015_g N_VGND_c_2778_n 0.00169411f $X=3.67 $Y=0.78 $X2=0 $Y2=0
cc_592 N_A_977_243#_c_714_n N_A_867_82#_c_922_n 0.00785719f $X=5.05 $Y=1.92
+ $X2=0 $Y2=0
cc_593 N_A_977_243#_c_716_n N_A_867_82#_c_922_n 0.0149921f $X=5.05 $Y=2.145
+ $X2=0 $Y2=0
cc_594 N_A_977_243#_c_717_n N_A_867_82#_c_922_n 0.00189254f $X=5.44 $Y=2.21
+ $X2=0 $Y2=0
cc_595 N_A_977_243#_c_718_n N_A_867_82#_c_922_n 9.05791e-19 $X=5.525 $Y=2.905
+ $X2=0 $Y2=0
cc_596 N_A_977_243#_c_723_n N_A_867_82#_c_922_n 9.36002e-19 $X=5.05 $Y=2.13
+ $X2=0 $Y2=0
cc_597 N_A_977_243#_c_712_n N_A_867_82#_c_923_n 0.0277489f $X=5.33 $Y=2.41 $X2=0
+ $Y2=0
cc_598 N_A_977_243#_c_718_n N_A_867_82#_c_923_n 0.00219826f $X=5.525 $Y=2.905
+ $X2=0 $Y2=0
cc_599 N_A_977_243#_c_725_n N_A_867_82#_c_923_n 0.0144629f $X=6.925 $Y=2.862
+ $X2=0 $Y2=0
cc_600 N_A_977_243#_M1043_g N_A_867_82#_c_904_n 6.85471e-19 $X=9.305 $Y=0.87
+ $X2=0 $Y2=0
cc_601 N_A_977_243#_c_707_n N_A_867_82#_c_904_n 0.0801441f $X=9.44 $Y=2.045
+ $X2=0 $Y2=0
cc_602 N_A_977_243#_c_710_n N_A_867_82#_c_904_n 0.00263288f $X=9.365 $Y=1.795
+ $X2=0 $Y2=0
cc_603 N_A_977_243#_c_708_n N_A_867_82#_c_907_n 0.0054081f $X=5.05 $Y=1.755
+ $X2=0 $Y2=0
cc_604 N_A_977_243#_c_723_n N_A_867_82#_c_907_n 0.00596281f $X=5.05 $Y=2.13
+ $X2=0 $Y2=0
cc_605 N_A_977_243#_c_712_n N_A_867_82#_c_926_n 0.00232031f $X=5.33 $Y=2.41
+ $X2=0 $Y2=0
cc_606 N_A_977_243#_c_716_n N_A_867_82#_c_926_n 0.00208937f $X=5.05 $Y=2.145
+ $X2=0 $Y2=0
cc_607 N_A_977_243#_c_718_n N_A_867_82#_c_926_n 0.0052334f $X=5.525 $Y=2.905
+ $X2=0 $Y2=0
cc_608 N_A_977_243#_c_723_n N_A_867_82#_c_926_n 0.0200965f $X=5.05 $Y=2.13 $X2=0
+ $Y2=0
cc_609 N_A_977_243#_c_724_n N_A_867_82#_c_926_n 0.00276193f $X=5.05 $Y=2.13
+ $X2=0 $Y2=0
cc_610 N_A_977_243#_c_704_n N_A_867_82#_c_908_n 0.00607421f $X=5.035 $Y=1.29
+ $X2=0 $Y2=0
cc_611 N_A_977_243#_M1043_g N_A_867_82#_c_909_n 0.00376456f $X=9.305 $Y=0.87
+ $X2=0 $Y2=0
cc_612 N_A_977_243#_M1043_g N_A_867_82#_c_915_n 0.00194703f $X=9.305 $Y=0.87
+ $X2=0 $Y2=0
cc_613 N_A_977_243#_c_707_n N_A_867_82#_c_915_n 0.00254955f $X=9.44 $Y=2.045
+ $X2=0 $Y2=0
cc_614 N_A_977_243#_c_709_n N_A_867_82#_c_915_n 0.0252739f $X=7.845 $Y=2.31
+ $X2=0 $Y2=0
cc_615 N_A_977_243#_c_751_p N_A_867_82#_c_915_n 0.00917432f $X=8.495 $Y=2.395
+ $X2=0 $Y2=0
cc_616 N_A_977_243#_c_710_n N_A_867_82#_c_915_n 0.0125354f $X=9.365 $Y=1.795
+ $X2=0 $Y2=0
cc_617 N_A_977_243#_c_711_n N_A_867_82#_c_915_n 0.00517428f $X=7.925 $Y=0.855
+ $X2=0 $Y2=0
cc_618 N_A_977_243#_c_714_n N_A_867_82#_c_916_n 3.82815e-19 $X=5.05 $Y=1.92
+ $X2=0 $Y2=0
cc_619 N_A_977_243#_c_708_n N_A_867_82#_c_916_n 5.77178e-19 $X=5.05 $Y=1.755
+ $X2=0 $Y2=0
cc_620 N_A_977_243#_c_717_n N_A_867_82#_c_916_n 0.00205096f $X=5.44 $Y=2.21
+ $X2=0 $Y2=0
cc_621 N_A_977_243#_M1043_g N_A_867_82#_c_917_n 9.84498e-19 $X=9.305 $Y=0.87
+ $X2=0 $Y2=0
cc_622 N_A_977_243#_c_707_n N_A_867_82#_c_917_n 6.86607e-19 $X=9.44 $Y=2.045
+ $X2=0 $Y2=0
cc_623 N_A_977_243#_c_710_n N_A_867_82#_c_917_n 0.00130845f $X=9.365 $Y=1.795
+ $X2=0 $Y2=0
cc_624 N_A_977_243#_M1043_g N_A_867_82#_c_918_n 0.00155948f $X=9.305 $Y=0.87
+ $X2=0 $Y2=0
cc_625 N_A_977_243#_c_707_n N_A_867_82#_c_918_n 0.00156894f $X=9.44 $Y=2.045
+ $X2=0 $Y2=0
cc_626 N_A_977_243#_c_710_n N_A_867_82#_c_918_n 0.020287f $X=9.365 $Y=1.795
+ $X2=0 $Y2=0
cc_627 N_A_977_243#_c_703_n N_A_867_82#_c_919_n 0.021405f $X=5.605 $Y=1.29 $X2=0
+ $Y2=0
cc_628 N_A_977_243#_c_714_n N_A_867_82#_c_919_n 0.0094248f $X=5.05 $Y=1.92 $X2=0
+ $Y2=0
cc_629 N_A_977_243#_c_708_n N_A_867_82#_c_919_n 0.00511549f $X=5.05 $Y=1.755
+ $X2=0 $Y2=0
cc_630 N_A_977_243#_c_717_n N_A_867_82#_c_919_n 0.0041804f $X=5.44 $Y=2.21 $X2=0
+ $Y2=0
cc_631 N_A_977_243#_c_703_n N_A_867_82#_c_920_n 0.00295526f $X=5.605 $Y=1.29
+ $X2=0 $Y2=0
cc_632 N_A_977_243#_c_714_n N_A_867_82#_c_920_n 0.00214398f $X=5.05 $Y=1.92
+ $X2=0 $Y2=0
cc_633 N_A_977_243#_c_708_n N_A_867_82#_c_920_n 0.0154842f $X=5.05 $Y=1.755
+ $X2=0 $Y2=0
cc_634 N_A_977_243#_c_716_n N_A_867_82#_c_920_n 0.00102646f $X=5.05 $Y=2.145
+ $X2=0 $Y2=0
cc_635 N_A_977_243#_c_717_n N_A_867_82#_c_920_n 0.00740117f $X=5.44 $Y=2.21
+ $X2=0 $Y2=0
cc_636 N_A_977_243#_c_723_n N_A_867_82#_c_920_n 0.014763f $X=5.05 $Y=2.13 $X2=0
+ $Y2=0
cc_637 N_A_977_243#_c_714_n N_A_867_82#_c_921_n 0.00157387f $X=5.05 $Y=1.92
+ $X2=0 $Y2=0
cc_638 N_A_977_243#_c_708_n N_A_867_82#_c_921_n 2.4101e-19 $X=5.05 $Y=1.755
+ $X2=0 $Y2=0
cc_639 N_A_977_243#_c_717_n N_A_867_82#_c_921_n 0.0126363f $X=5.44 $Y=2.21 $X2=0
+ $Y2=0
cc_640 N_A_977_243#_c_709_n N_A_1159_497#_c_1126_n 0.00365232f $X=7.845 $Y=2.31
+ $X2=0 $Y2=0
cc_641 N_A_977_243#_c_777_p N_A_1159_497#_c_1134_n 0.00963777f $X=7.76 $Y=2.735
+ $X2=0 $Y2=0
cc_642 N_A_977_243#_c_709_n N_A_1159_497#_c_1134_n 0.00158303f $X=7.845 $Y=2.31
+ $X2=0 $Y2=0
cc_643 N_A_977_243#_c_779_p N_A_1159_497#_c_1134_n 0.00368225f $X=7.845 $Y=2.65
+ $X2=0 $Y2=0
cc_644 N_A_977_243#_c_726_n N_A_1159_497#_c_1134_n 0.00784164f $X=7.505 $Y=2.862
+ $X2=0 $Y2=0
cc_645 N_A_977_243#_c_781_p N_A_1159_497#_c_1134_n 0.00117798f $X=7.845 $Y=2.395
+ $X2=0 $Y2=0
cc_646 N_A_977_243#_c_711_n N_A_1159_497#_c_1127_n 0.00496598f $X=7.925 $Y=0.855
+ $X2=0 $Y2=0
cc_647 N_A_977_243#_c_709_n N_A_1159_497#_c_1128_n 0.00496598f $X=7.845 $Y=2.31
+ $X2=0 $Y2=0
cc_648 N_A_977_243#_M1046_s N_A_1159_497#_c_1135_n 0.00292388f $X=7.025 $Y=2.12
+ $X2=0 $Y2=0
cc_649 N_A_977_243#_c_717_n N_A_1159_497#_c_1138_n 0.00822198f $X=5.44 $Y=2.21
+ $X2=0 $Y2=0
cc_650 N_A_977_243#_c_718_n N_A_1159_497#_c_1138_n 0.0187803f $X=5.525 $Y=2.905
+ $X2=0 $Y2=0
cc_651 N_A_977_243#_c_725_n N_A_1159_497#_c_1138_n 0.0229036f $X=6.925 $Y=2.862
+ $X2=0 $Y2=0
cc_652 N_A_977_243#_c_709_n N_A_1579_258#_c_1221_n 0.00954358f $X=7.845 $Y=2.31
+ $X2=0 $Y2=0
cc_653 N_A_977_243#_c_777_p N_A_1579_258#_c_1243_n 0.00403181f $X=7.76 $Y=2.735
+ $X2=0 $Y2=0
cc_654 N_A_977_243#_c_709_n N_A_1579_258#_c_1243_n 0.00824718f $X=7.845 $Y=2.31
+ $X2=0 $Y2=0
cc_655 N_A_977_243#_c_779_p N_A_1579_258#_c_1243_n 0.00420583f $X=7.845 $Y=2.65
+ $X2=0 $Y2=0
cc_656 N_A_977_243#_c_751_p N_A_1579_258#_c_1243_n 0.010177f $X=8.495 $Y=2.395
+ $X2=0 $Y2=0
cc_657 N_A_977_243#_c_726_n N_A_1579_258#_c_1243_n 7.54449e-19 $X=7.505 $Y=2.862
+ $X2=0 $Y2=0
cc_658 N_A_977_243#_c_781_p N_A_1579_258#_c_1243_n 0.00154168f $X=7.845 $Y=2.395
+ $X2=0 $Y2=0
cc_659 N_A_977_243#_c_727_n N_A_1579_258#_c_1243_n 5.35128e-19 $X=8.66 $Y=2.475
+ $X2=0 $Y2=0
cc_660 N_A_977_243#_c_709_n N_A_1579_258#_M1047_g 0.00474029f $X=7.845 $Y=2.31
+ $X2=0 $Y2=0
cc_661 N_A_977_243#_c_711_n N_A_1579_258#_M1047_g 0.00700206f $X=7.925 $Y=0.855
+ $X2=0 $Y2=0
cc_662 N_A_977_243#_M1043_g N_A_1579_258#_c_1226_n 0.0157265f $X=9.305 $Y=0.87
+ $X2=0 $Y2=0
cc_663 N_A_977_243#_c_707_n N_A_1579_258#_c_1226_n 0.00136408f $X=9.44 $Y=2.045
+ $X2=0 $Y2=0
cc_664 N_A_977_243#_c_721_n N_A_1579_258#_c_1226_n 0.00191594f $X=9.2 $Y=2.215
+ $X2=0 $Y2=0
cc_665 N_A_977_243#_c_710_n N_A_1579_258#_c_1226_n 0.0213603f $X=9.365 $Y=1.795
+ $X2=0 $Y2=0
cc_666 N_A_977_243#_M1043_g N_A_1579_258#_c_1227_n 0.00631281f $X=9.305 $Y=0.87
+ $X2=0 $Y2=0
cc_667 N_A_977_243#_M1043_g N_A_1579_258#_c_1229_n 7.27055e-19 $X=9.305 $Y=0.87
+ $X2=0 $Y2=0
cc_668 N_A_977_243#_c_709_n N_A_1579_258#_c_1237_n 0.0234076f $X=7.845 $Y=2.31
+ $X2=0 $Y2=0
cc_669 N_A_977_243#_c_709_n N_A_1579_258#_c_1238_n 0.00811935f $X=7.845 $Y=2.31
+ $X2=0 $Y2=0
cc_670 N_A_977_243#_c_751_p N_A_1579_258#_c_1238_n 0.00202692f $X=8.495 $Y=2.395
+ $X2=0 $Y2=0
cc_671 N_A_977_243#_c_711_n N_A_1579_258#_c_1238_n 0.00477998f $X=7.925 $Y=0.855
+ $X2=0 $Y2=0
cc_672 N_A_977_243#_c_709_n N_SET_B_c_1429_n 9.03836e-19 $X=7.845 $Y=2.31
+ $X2=-0.19 $Y2=-0.245
cc_673 N_A_977_243#_c_779_p N_SET_B_c_1429_n 4.40639e-19 $X=7.845 $Y=2.65
+ $X2=-0.19 $Y2=-0.245
cc_674 N_A_977_243#_c_751_p N_SET_B_c_1429_n 0.00891054f $X=8.495 $Y=2.395
+ $X2=-0.19 $Y2=-0.245
cc_675 N_A_977_243#_c_710_n N_SET_B_c_1429_n 0.00109172f $X=9.365 $Y=1.795
+ $X2=-0.19 $Y2=-0.245
cc_676 N_A_977_243#_c_727_n N_SET_B_c_1429_n 0.014f $X=8.66 $Y=2.475 $X2=-0.19
+ $Y2=-0.245
cc_677 N_A_977_243#_M1043_g N_SET_B_M1025_g 0.0261819f $X=9.305 $Y=0.87 $X2=0
+ $Y2=0
cc_678 N_A_977_243#_c_707_n N_SET_B_c_1431_n 4.11658e-19 $X=9.44 $Y=2.045 $X2=0
+ $Y2=0
cc_679 N_A_977_243#_c_721_n N_SET_B_c_1431_n 0.0127763f $X=9.2 $Y=2.215 $X2=0
+ $Y2=0
cc_680 N_A_977_243#_c_710_n N_SET_B_c_1431_n 0.0289342f $X=9.365 $Y=1.795 $X2=0
+ $Y2=0
cc_681 N_A_977_243#_c_727_n N_SET_B_c_1431_n 0.00851502f $X=8.66 $Y=2.475 $X2=0
+ $Y2=0
cc_682 N_A_977_243#_M1026_d N_SET_B_c_1432_n 8.54521e-19 $X=8.51 $Y=2.12 $X2=0
+ $Y2=0
cc_683 N_A_977_243#_c_709_n N_SET_B_c_1432_n 0.00655644f $X=7.845 $Y=2.31 $X2=0
+ $Y2=0
cc_684 N_A_977_243#_c_751_p N_SET_B_c_1432_n 0.0067036f $X=8.495 $Y=2.395 $X2=0
+ $Y2=0
cc_685 N_A_977_243#_c_727_n N_SET_B_c_1432_n 0.00243464f $X=8.66 $Y=2.475 $X2=0
+ $Y2=0
cc_686 N_A_977_243#_c_707_n N_SET_B_c_1426_n 0.00113722f $X=9.44 $Y=2.045 $X2=0
+ $Y2=0
cc_687 N_A_977_243#_c_709_n N_SET_B_c_1426_n 0.0124311f $X=7.845 $Y=2.31 $X2=0
+ $Y2=0
cc_688 N_A_977_243#_c_751_p N_SET_B_c_1426_n 0.0101614f $X=8.495 $Y=2.395 $X2=0
+ $Y2=0
cc_689 N_A_977_243#_c_721_n N_SET_B_c_1426_n 0.00935265f $X=9.2 $Y=2.215 $X2=0
+ $Y2=0
cc_690 N_A_977_243#_c_710_n N_SET_B_c_1426_n 0.0204309f $X=9.365 $Y=1.795 $X2=0
+ $Y2=0
cc_691 N_A_977_243#_c_727_n N_SET_B_c_1426_n 0.0151312f $X=8.66 $Y=2.475 $X2=0
+ $Y2=0
cc_692 N_A_977_243#_c_707_n N_SET_B_c_1427_n 0.0230853f $X=9.44 $Y=2.045 $X2=0
+ $Y2=0
cc_693 N_A_977_243#_c_721_n N_SET_B_c_1427_n 0.00301959f $X=9.2 $Y=2.215 $X2=0
+ $Y2=0
cc_694 N_A_977_243#_c_710_n N_SET_B_c_1427_n 0.00180627f $X=9.365 $Y=1.795 $X2=0
+ $Y2=0
cc_695 N_A_977_243#_c_727_n N_SET_B_c_1427_n 0.00544666f $X=8.66 $Y=2.475 $X2=0
+ $Y2=0
cc_696 N_A_977_243#_c_704_n N_A_662_82#_M1016_g 0.00183589f $X=5.035 $Y=1.29
+ $X2=0 $Y2=0
cc_697 N_A_977_243#_c_704_n N_A_662_82#_c_1559_n 0.00823117f $X=5.035 $Y=1.29
+ $X2=0 $Y2=0
cc_698 N_A_977_243#_c_714_n N_A_662_82#_c_1559_n 0.00530385f $X=5.05 $Y=1.92
+ $X2=0 $Y2=0
cc_699 N_A_977_243#_c_708_n N_A_662_82#_c_1559_n 0.00169862f $X=5.05 $Y=1.755
+ $X2=0 $Y2=0
cc_700 N_A_977_243#_M1021_g N_A_662_82#_c_1560_n 0.0103107f $X=5.68 $Y=0.805
+ $X2=0 $Y2=0
cc_701 N_A_977_243#_M1021_g N_A_662_82#_M1017_g 0.0226239f $X=5.68 $Y=0.805
+ $X2=0 $Y2=0
cc_702 N_A_977_243#_c_703_n N_A_662_82#_c_1563_n 0.00540592f $X=5.605 $Y=1.29
+ $X2=0 $Y2=0
cc_703 N_A_977_243#_M1043_g N_A_662_82#_c_1564_n 0.0104164f $X=9.305 $Y=0.87
+ $X2=0 $Y2=0
cc_704 N_A_977_243#_c_725_n N_A_662_82#_c_1576_n 0.0152404f $X=6.925 $Y=2.862
+ $X2=0 $Y2=0
cc_705 N_A_977_243#_c_726_n N_A_662_82#_c_1576_n 0.00458801f $X=7.505 $Y=2.862
+ $X2=0 $Y2=0
cc_706 N_A_977_243#_M1043_g N_A_662_82#_M1027_g 0.0409189f $X=9.305 $Y=0.87
+ $X2=0 $Y2=0
cc_707 N_A_977_243#_c_703_n N_A_662_82#_c_1569_n 0.0226239f $X=5.605 $Y=1.29
+ $X2=0 $Y2=0
cc_708 N_A_977_243#_c_707_n N_A_1954_119#_c_1984_n 0.00227497f $X=9.44 $Y=2.045
+ $X2=0 $Y2=0
cc_709 N_A_977_243#_c_710_n N_A_1954_119#_c_1996_n 6.17874e-19 $X=9.365 $Y=1.795
+ $X2=0 $Y2=0
cc_710 N_A_977_243#_c_751_p N_VPWR_M1022_d 0.00375655f $X=8.495 $Y=2.395 $X2=0
+ $Y2=0
cc_711 N_A_977_243#_c_721_n N_VPWR_M1012_s 0.00562228f $X=9.2 $Y=2.215 $X2=0
+ $Y2=0
cc_712 N_A_977_243#_c_712_n N_VPWR_c_2281_n 0.00925598f $X=5.33 $Y=2.41 $X2=0
+ $Y2=0
cc_713 N_A_977_243#_c_716_n N_VPWR_c_2281_n 0.00244683f $X=5.05 $Y=2.145 $X2=0
+ $Y2=0
cc_714 N_A_977_243#_c_717_n N_VPWR_c_2281_n 0.00429362f $X=5.44 $Y=2.21 $X2=0
+ $Y2=0
cc_715 N_A_977_243#_c_718_n N_VPWR_c_2281_n 0.016537f $X=5.525 $Y=2.905 $X2=0
+ $Y2=0
cc_716 N_A_977_243#_c_719_n N_VPWR_c_2281_n 0.0141804f $X=5.61 $Y=2.99 $X2=0
+ $Y2=0
cc_717 N_A_977_243#_c_723_n N_VPWR_c_2281_n 0.0163558f $X=5.05 $Y=2.13 $X2=0
+ $Y2=0
cc_718 N_A_977_243#_c_777_p N_VPWR_c_2282_n 0.0120091f $X=7.76 $Y=2.735 $X2=0
+ $Y2=0
cc_719 N_A_977_243#_c_751_p N_VPWR_c_2282_n 0.0132576f $X=8.495 $Y=2.395 $X2=0
+ $Y2=0
cc_720 N_A_977_243#_c_726_n N_VPWR_c_2282_n 0.00724127f $X=7.505 $Y=2.862 $X2=0
+ $Y2=0
cc_721 N_A_977_243#_c_727_n N_VPWR_c_2282_n 0.0215476f $X=8.66 $Y=2.475 $X2=0
+ $Y2=0
cc_722 N_A_977_243#_c_707_n N_VPWR_c_2283_n 0.0164499f $X=9.44 $Y=2.045 $X2=0
+ $Y2=0
cc_723 N_A_977_243#_c_721_n N_VPWR_c_2283_n 0.0216233f $X=9.2 $Y=2.215 $X2=0
+ $Y2=0
cc_724 N_A_977_243#_c_727_n N_VPWR_c_2283_n 0.0355056f $X=8.66 $Y=2.475 $X2=0
+ $Y2=0
cc_725 N_A_977_243#_c_712_n N_VPWR_c_2286_n 0.0048289f $X=5.33 $Y=2.41 $X2=0
+ $Y2=0
cc_726 N_A_977_243#_c_719_n N_VPWR_c_2286_n 0.0121867f $X=5.61 $Y=2.99 $X2=0
+ $Y2=0
cc_727 N_A_977_243#_c_777_p N_VPWR_c_2286_n 0.00893233f $X=7.76 $Y=2.735 $X2=0
+ $Y2=0
cc_728 N_A_977_243#_c_725_n N_VPWR_c_2286_n 0.124483f $X=6.925 $Y=2.862 $X2=0
+ $Y2=0
cc_729 N_A_977_243#_c_707_n N_VPWR_c_2289_n 0.00413917f $X=9.44 $Y=2.045 $X2=0
+ $Y2=0
cc_730 N_A_977_243#_c_727_n N_VPWR_c_2295_n 0.0148091f $X=8.66 $Y=2.475 $X2=0
+ $Y2=0
cc_731 N_A_977_243#_c_712_n N_VPWR_c_2276_n 0.0047904f $X=5.33 $Y=2.41 $X2=0
+ $Y2=0
cc_732 N_A_977_243#_c_707_n N_VPWR_c_2276_n 0.00817239f $X=9.44 $Y=2.045 $X2=0
+ $Y2=0
cc_733 N_A_977_243#_c_719_n N_VPWR_c_2276_n 0.00660921f $X=5.61 $Y=2.99 $X2=0
+ $Y2=0
cc_734 N_A_977_243#_c_777_p N_VPWR_c_2276_n 0.0128749f $X=7.76 $Y=2.735 $X2=0
+ $Y2=0
cc_735 N_A_977_243#_c_751_p N_VPWR_c_2276_n 0.0122122f $X=8.495 $Y=2.395 $X2=0
+ $Y2=0
cc_736 N_A_977_243#_c_725_n N_VPWR_c_2276_n 0.0716319f $X=6.925 $Y=2.862 $X2=0
+ $Y2=0
cc_737 N_A_977_243#_c_727_n N_VPWR_c_2276_n 0.0122282f $X=8.66 $Y=2.475 $X2=0
+ $Y2=0
cc_738 N_A_977_243#_c_704_n N_A_197_119#_c_2475_n 0.00226961f $X=5.035 $Y=1.29
+ $X2=0 $Y2=0
cc_739 N_A_977_243#_M1021_g N_A_197_119#_c_2475_n 3.66969e-19 $X=5.68 $Y=0.805
+ $X2=0 $Y2=0
cc_740 N_A_977_243#_M1021_g N_A_197_119#_c_2477_n 0.00323463f $X=5.68 $Y=0.805
+ $X2=0 $Y2=0
cc_741 N_A_977_243#_c_703_n N_A_197_119#_c_2478_n 0.0205411f $X=5.605 $Y=1.29
+ $X2=0 $Y2=0
cc_742 N_A_977_243#_M1021_g N_A_197_119#_c_2478_n 0.00627334f $X=5.68 $Y=0.805
+ $X2=0 $Y2=0
cc_743 N_A_977_243#_c_703_n N_A_197_119#_c_2479_n 0.00405018f $X=5.605 $Y=1.29
+ $X2=0 $Y2=0
cc_744 N_A_977_243#_c_704_n N_A_197_119#_c_2479_n 0.00383886f $X=5.035 $Y=1.29
+ $X2=0 $Y2=0
cc_745 N_A_977_243#_c_708_n N_A_197_119#_c_2479_n 0.00144422f $X=5.05 $Y=1.755
+ $X2=0 $Y2=0
cc_746 N_A_977_243#_M1021_g N_A_197_119#_c_2480_n 0.00439723f $X=5.68 $Y=0.805
+ $X2=0 $Y2=0
cc_747 N_A_977_243#_M1046_s N_A_197_119#_c_2493_n 0.012268f $X=7.025 $Y=2.12
+ $X2=0 $Y2=0
cc_748 N_A_977_243#_c_725_n N_A_197_119#_c_2493_n 0.00782502f $X=6.925 $Y=2.862
+ $X2=0 $Y2=0
cc_749 N_A_977_243#_c_726_n N_A_197_119#_c_2493_n 0.0464242f $X=7.505 $Y=2.862
+ $X2=0 $Y2=0
cc_750 N_A_977_243#_c_781_p N_A_197_119#_c_2493_n 0.0148586f $X=7.845 $Y=2.395
+ $X2=0 $Y2=0
cc_751 N_A_977_243#_c_711_n N_A_197_119#_c_2484_n 0.0140085f $X=7.925 $Y=0.855
+ $X2=0 $Y2=0
cc_752 N_A_977_243#_M1046_s N_A_197_119#_c_2486_n 0.00666089f $X=7.025 $Y=2.12
+ $X2=0 $Y2=0
cc_753 N_A_977_243#_c_711_n N_A_197_119#_c_2486_n 0.0957029f $X=7.925 $Y=0.855
+ $X2=0 $Y2=0
cc_754 N_A_977_243#_c_725_n N_A_197_119#_c_2496_n 0.023777f $X=6.925 $Y=2.862
+ $X2=0 $Y2=0
cc_755 N_A_977_243#_c_726_n N_A_197_119#_c_2496_n 0.00600942f $X=7.505 $Y=2.862
+ $X2=0 $Y2=0
cc_756 N_A_977_243#_c_718_n A_1081_497# 0.00171032f $X=5.525 $Y=2.905 $X2=-0.19
+ $Y2=-0.245
cc_757 N_A_977_243#_c_777_p A_1528_424# 0.00470748f $X=7.76 $Y=2.735 $X2=-0.19
+ $Y2=-0.245
cc_758 N_A_977_243#_c_709_n A_1528_424# 0.00155805f $X=7.845 $Y=2.31 $X2=-0.19
+ $Y2=-0.245
cc_759 N_A_977_243#_c_779_p A_1528_424# 0.00189206f $X=7.845 $Y=2.65 $X2=-0.19
+ $Y2=-0.245
cc_760 N_A_977_243#_c_781_p A_1528_424# 0.00145568f $X=7.845 $Y=2.395 $X2=-0.19
+ $Y2=-0.245
cc_761 N_A_977_243#_c_703_n N_VGND_c_2762_n 0.00236747f $X=5.605 $Y=1.29 $X2=0
+ $Y2=0
cc_762 N_A_977_243#_M1021_g N_VGND_c_2762_n 0.00988925f $X=5.68 $Y=0.805 $X2=0
+ $Y2=0
cc_763 N_A_977_243#_M1043_g N_VGND_c_2763_n 0.00588057f $X=9.305 $Y=0.87 $X2=0
+ $Y2=0
cc_764 N_A_977_243#_M1021_g N_VGND_c_2776_n 7.88961e-19 $X=5.68 $Y=0.805 $X2=0
+ $Y2=0
cc_765 N_A_977_243#_M1043_g N_VGND_c_2776_n 9.39239e-19 $X=9.305 $Y=0.87 $X2=0
+ $Y2=0
cc_766 N_A_977_243#_c_711_n N_A_1434_78#_c_2931_n 0.0228873f $X=7.925 $Y=0.855
+ $X2=0 $Y2=0
cc_767 N_A_867_82#_c_915_n N_A_1159_497#_c_1124_n 9.42131e-19 $X=9.695 $Y=1.665
+ $X2=0 $Y2=0
cc_768 N_A_867_82#_M1001_g N_A_1159_497#_c_1125_n 0.00763412f $X=6.47 $Y=0.805
+ $X2=0 $Y2=0
cc_769 N_A_867_82#_c_915_n N_A_1159_497#_c_1126_n 0.00613284f $X=9.695 $Y=1.665
+ $X2=0 $Y2=0
cc_770 N_A_867_82#_c_915_n N_A_1159_497#_c_1128_n 8.25895e-19 $X=9.695 $Y=1.665
+ $X2=0 $Y2=0
cc_771 N_A_867_82#_M1001_g N_A_1159_497#_c_1129_n 0.0124832f $X=6.47 $Y=0.805
+ $X2=0 $Y2=0
cc_772 N_A_867_82#_c_913_n N_A_1159_497#_c_1135_n 0.00798977f $X=6.545 $Y=1.635
+ $X2=0 $Y2=0
cc_773 N_A_867_82#_c_914_n N_A_1159_497#_c_1135_n 0.0359077f $X=6.38 $Y=1.635
+ $X2=0 $Y2=0
cc_774 N_A_867_82#_c_915_n N_A_1159_497#_c_1135_n 0.00952883f $X=9.695 $Y=1.665
+ $X2=0 $Y2=0
cc_775 N_A_867_82#_M1001_g N_A_1159_497#_c_1130_n 0.012535f $X=6.47 $Y=0.805
+ $X2=0 $Y2=0
cc_776 N_A_867_82#_c_912_n N_A_1159_497#_c_1130_n 0.0198439f $X=6.545 $Y=1.635
+ $X2=0 $Y2=0
cc_777 N_A_867_82#_c_913_n N_A_1159_497#_c_1130_n 0.00369939f $X=6.545 $Y=1.635
+ $X2=0 $Y2=0
cc_778 N_A_867_82#_c_915_n N_A_1159_497#_c_1130_n 0.00734224f $X=9.695 $Y=1.665
+ $X2=0 $Y2=0
cc_779 N_A_867_82#_M1001_g N_A_1159_497#_c_1131_n 0.00236995f $X=6.47 $Y=0.805
+ $X2=0 $Y2=0
cc_780 N_A_867_82#_c_912_n N_A_1159_497#_c_1131_n 0.00302679f $X=6.545 $Y=1.635
+ $X2=0 $Y2=0
cc_781 N_A_867_82#_c_913_n N_A_1159_497#_c_1131_n 3.49216e-19 $X=6.545 $Y=1.635
+ $X2=0 $Y2=0
cc_782 N_A_867_82#_c_914_n N_A_1159_497#_c_1131_n 0.0119633f $X=6.38 $Y=1.635
+ $X2=0 $Y2=0
cc_783 N_A_867_82#_c_915_n N_A_1159_497#_c_1131_n 0.00187073f $X=9.695 $Y=1.665
+ $X2=0 $Y2=0
cc_784 N_A_867_82#_M1001_g N_A_1159_497#_c_1136_n 9.84843e-19 $X=6.47 $Y=0.805
+ $X2=0 $Y2=0
cc_785 N_A_867_82#_c_912_n N_A_1159_497#_c_1136_n 0.0196546f $X=6.545 $Y=1.635
+ $X2=0 $Y2=0
cc_786 N_A_867_82#_c_913_n N_A_1159_497#_c_1136_n 5.12632e-19 $X=6.545 $Y=1.635
+ $X2=0 $Y2=0
cc_787 N_A_867_82#_c_915_n N_A_1159_497#_c_1136_n 0.0303238f $X=9.695 $Y=1.665
+ $X2=0 $Y2=0
cc_788 N_A_867_82#_c_912_n N_A_1159_497#_c_1132_n 0.00114056f $X=6.545 $Y=1.635
+ $X2=0 $Y2=0
cc_789 N_A_867_82#_c_913_n N_A_1159_497#_c_1132_n 0.0214805f $X=6.545 $Y=1.635
+ $X2=0 $Y2=0
cc_790 N_A_867_82#_c_915_n N_A_1159_497#_c_1132_n 0.00138807f $X=9.695 $Y=1.665
+ $X2=0 $Y2=0
cc_791 N_A_867_82#_c_922_n N_A_1159_497#_c_1138_n 0.00341177f $X=5.72 $Y=2.32
+ $X2=0 $Y2=0
cc_792 N_A_867_82#_c_923_n N_A_1159_497#_c_1138_n 0.00321294f $X=5.72 $Y=2.41
+ $X2=0 $Y2=0
cc_793 N_A_867_82#_c_914_n N_A_1159_497#_c_1138_n 0.0179531f $X=6.38 $Y=1.635
+ $X2=0 $Y2=0
cc_794 N_A_867_82#_c_915_n N_A_1159_497#_c_1138_n 0.00230166f $X=9.695 $Y=1.665
+ $X2=0 $Y2=0
cc_795 N_A_867_82#_c_915_n N_A_1579_258#_c_1221_n 0.00331659f $X=9.695 $Y=1.665
+ $X2=0 $Y2=0
cc_796 N_A_867_82#_c_909_n N_A_1579_258#_c_1226_n 0.0155638f $X=10.07 $Y=1.407
+ $X2=0 $Y2=0
cc_797 N_A_867_82#_c_915_n N_A_1579_258#_c_1226_n 0.0311861f $X=9.695 $Y=1.665
+ $X2=0 $Y2=0
cc_798 N_A_867_82#_c_909_n N_A_1579_258#_c_1227_n 0.00235941f $X=10.07 $Y=1.407
+ $X2=0 $Y2=0
cc_799 N_A_867_82#_M1039_g N_A_1579_258#_c_1228_n 0.00540343f $X=10.745 $Y=0.805
+ $X2=0 $Y2=0
cc_800 N_A_867_82#_M1039_g N_A_1579_258#_c_1230_n 3.18691e-19 $X=10.745 $Y=0.805
+ $X2=0 $Y2=0
cc_801 N_A_867_82#_c_915_n N_A_1579_258#_c_1237_n 0.0158677f $X=9.695 $Y=1.665
+ $X2=0 $Y2=0
cc_802 N_A_867_82#_c_915_n N_A_1579_258#_c_1238_n 0.0053521f $X=9.695 $Y=1.665
+ $X2=0 $Y2=0
cc_803 N_A_867_82#_M1039_g N_A_1579_258#_c_1239_n 0.0133178f $X=10.745 $Y=0.805
+ $X2=0 $Y2=0
cc_804 N_A_867_82#_c_915_n N_SET_B_M1025_g 0.00182015f $X=9.695 $Y=1.665 $X2=0
+ $Y2=0
cc_805 N_A_867_82#_c_904_n N_SET_B_c_1431_n 0.00979312f $X=9.83 $Y=2.045 $X2=0
+ $Y2=0
cc_806 N_A_867_82#_c_910_n N_SET_B_c_1431_n 0.0059316f $X=10.835 $Y=1.41 $X2=0
+ $Y2=0
cc_807 N_A_867_82#_c_915_n N_SET_B_c_1431_n 0.0845048f $X=9.695 $Y=1.665 $X2=0
+ $Y2=0
cc_808 N_A_867_82#_c_917_n N_SET_B_c_1431_n 0.0242419f $X=9.84 $Y=1.665 $X2=0
+ $Y2=0
cc_809 N_A_867_82#_c_918_n N_SET_B_c_1431_n 0.00910799f $X=9.84 $Y=1.665 $X2=0
+ $Y2=0
cc_810 N_A_867_82#_c_915_n N_SET_B_c_1432_n 0.0243554f $X=9.695 $Y=1.665 $X2=0
+ $Y2=0
cc_811 N_A_867_82#_c_915_n N_SET_B_c_1426_n 0.0168952f $X=9.695 $Y=1.665 $X2=0
+ $Y2=0
cc_812 N_A_867_82#_c_915_n N_SET_B_c_1427_n 0.00317885f $X=9.695 $Y=1.665 $X2=0
+ $Y2=0
cc_813 N_A_867_82#_c_906_n N_A_662_82#_M1016_g 0.00876799f $X=4.61 $Y=1.045
+ $X2=0 $Y2=0
cc_814 N_A_867_82#_c_908_n N_A_662_82#_M1016_g 0.00204565f $X=4.7 $Y=1.55 $X2=0
+ $Y2=0
cc_815 N_A_867_82#_c_906_n N_A_662_82#_c_1559_n 0.00430983f $X=4.61 $Y=1.045
+ $X2=0 $Y2=0
cc_816 N_A_867_82#_c_907_n N_A_662_82#_c_1559_n 0.00767334f $X=4.58 $Y=2.04
+ $X2=0 $Y2=0
cc_817 N_A_867_82#_c_926_n N_A_662_82#_c_1559_n 0.012147f $X=4.545 $Y=2.815
+ $X2=0 $Y2=0
cc_818 N_A_867_82#_c_908_n N_A_662_82#_c_1559_n 0.00178499f $X=4.7 $Y=1.55 $X2=0
+ $Y2=0
cc_819 N_A_867_82#_M1001_g N_A_662_82#_M1017_g 0.00955219f $X=6.47 $Y=0.805
+ $X2=0 $Y2=0
cc_820 N_A_867_82#_c_912_n N_A_662_82#_c_1563_n 5.27994e-19 $X=6.545 $Y=1.635
+ $X2=0 $Y2=0
cc_821 N_A_867_82#_c_913_n N_A_662_82#_c_1563_n 0.0209314f $X=6.545 $Y=1.635
+ $X2=0 $Y2=0
cc_822 N_A_867_82#_c_914_n N_A_662_82#_c_1563_n 0.0175879f $X=6.38 $Y=1.635
+ $X2=0 $Y2=0
cc_823 N_A_867_82#_c_919_n N_A_662_82#_c_1563_n 0.0226181f $X=5.59 $Y=1.74 $X2=0
+ $Y2=0
cc_824 N_A_867_82#_c_921_n N_A_662_82#_c_1563_n 6.07496e-19 $X=5.755 $Y=1.727
+ $X2=0 $Y2=0
cc_825 N_A_867_82#_M1001_g N_A_662_82#_c_1564_n 0.00882199f $X=6.47 $Y=0.805
+ $X2=0 $Y2=0
cc_826 N_A_867_82#_c_922_n N_A_662_82#_c_1576_n 0.00425795f $X=5.72 $Y=2.32
+ $X2=0 $Y2=0
cc_827 N_A_867_82#_c_923_n N_A_662_82#_c_1576_n 0.0137548f $X=5.72 $Y=2.41 $X2=0
+ $Y2=0
cc_828 N_A_867_82#_M1039_g N_A_662_82#_c_1566_n 0.0100284f $X=10.745 $Y=0.805
+ $X2=0 $Y2=0
cc_829 N_A_867_82#_c_909_n N_A_662_82#_c_1566_n 0.00793522f $X=10.07 $Y=1.407
+ $X2=0 $Y2=0
cc_830 N_A_867_82#_c_910_n N_A_662_82#_c_1566_n 0.0107459f $X=10.835 $Y=1.41
+ $X2=0 $Y2=0
cc_831 N_A_867_82#_c_904_n N_A_662_82#_c_1567_n 0.018105f $X=9.83 $Y=2.045 $X2=0
+ $Y2=0
cc_832 N_A_867_82#_c_909_n N_A_662_82#_c_1567_n 0.00324447f $X=10.07 $Y=1.407
+ $X2=0 $Y2=0
cc_833 N_A_867_82#_c_915_n N_A_662_82#_c_1567_n 0.00201241f $X=9.695 $Y=1.665
+ $X2=0 $Y2=0
cc_834 N_A_867_82#_c_917_n N_A_662_82#_c_1567_n 8.82569e-19 $X=9.84 $Y=1.665
+ $X2=0 $Y2=0
cc_835 N_A_867_82#_c_904_n N_A_662_82#_c_1577_n 0.0122722f $X=9.83 $Y=2.045
+ $X2=0 $Y2=0
cc_836 N_A_867_82#_M1001_g N_A_662_82#_c_1569_n 0.0223854f $X=6.47 $Y=0.805
+ $X2=0 $Y2=0
cc_837 N_A_867_82#_c_914_n N_A_662_82#_c_1569_n 0.00188221f $X=6.38 $Y=1.635
+ $X2=0 $Y2=0
cc_838 N_A_867_82#_c_922_n N_A_662_82#_c_1578_n 0.0138987f $X=5.72 $Y=2.32 $X2=0
+ $Y2=0
cc_839 N_A_867_82#_c_914_n N_A_662_82#_c_1578_n 0.00106428f $X=6.38 $Y=1.635
+ $X2=0 $Y2=0
cc_840 N_A_867_82#_c_904_n N_A_662_82#_c_1570_n 0.0276602f $X=9.83 $Y=2.045
+ $X2=0 $Y2=0
cc_841 N_A_867_82#_c_910_n N_A_662_82#_c_1570_n 0.0106203f $X=10.835 $Y=1.41
+ $X2=0 $Y2=0
cc_842 N_A_867_82#_c_911_n N_A_662_82#_c_1570_n 0.0100284f $X=10.835 $Y=1.41
+ $X2=0 $Y2=0
cc_843 N_A_867_82#_c_918_n N_A_662_82#_c_1570_n 0.00296359f $X=9.84 $Y=1.665
+ $X2=0 $Y2=0
cc_844 N_A_867_82#_c_906_n N_A_662_82#_c_1571_n 0.0107975f $X=4.61 $Y=1.045
+ $X2=0 $Y2=0
cc_845 N_A_867_82#_c_926_n N_A_662_82#_c_1581_n 0.0044927f $X=4.545 $Y=2.815
+ $X2=0 $Y2=0
cc_846 N_A_867_82#_c_907_n N_A_662_82#_c_1603_n 0.00578301f $X=4.58 $Y=2.04
+ $X2=0 $Y2=0
cc_847 N_A_867_82#_c_926_n N_A_662_82#_c_1603_n 0.0050928f $X=4.545 $Y=2.815
+ $X2=0 $Y2=0
cc_848 N_A_867_82#_c_908_n N_A_662_82#_c_1572_n 0.00628822f $X=4.7 $Y=1.55 $X2=0
+ $Y2=0
cc_849 N_A_867_82#_c_907_n N_A_662_82#_c_1582_n 0.0128442f $X=4.58 $Y=2.04 $X2=0
+ $Y2=0
cc_850 N_A_867_82#_c_906_n N_A_662_82#_c_1573_n 0.0099668f $X=4.61 $Y=1.045
+ $X2=0 $Y2=0
cc_851 N_A_867_82#_c_907_n N_A_662_82#_c_1573_n 0.013185f $X=4.58 $Y=2.04 $X2=0
+ $Y2=0
cc_852 N_A_867_82#_c_908_n N_A_662_82#_c_1573_n 0.0162508f $X=4.7 $Y=1.55 $X2=0
+ $Y2=0
cc_853 N_A_867_82#_c_911_n N_A_2133_410#_c_1756_n 0.00776335f $X=10.835 $Y=1.41
+ $X2=0 $Y2=0
cc_854 N_A_867_82#_M1039_g N_A_2133_410#_M1010_g 0.0219184f $X=10.745 $Y=0.805
+ $X2=0 $Y2=0
cc_855 N_A_867_82#_c_910_n N_A_2133_410#_M1010_g 3.39166e-19 $X=10.835 $Y=1.41
+ $X2=0 $Y2=0
cc_856 N_A_867_82#_c_911_n N_A_2133_410#_M1010_g 0.0212382f $X=10.835 $Y=1.41
+ $X2=0 $Y2=0
cc_857 N_A_867_82#_c_904_n N_A_1954_119#_c_1984_n 0.013795f $X=9.83 $Y=2.045
+ $X2=0 $Y2=0
cc_858 N_A_867_82#_c_904_n N_A_1954_119#_c_1985_n 0.00254351f $X=9.83 $Y=2.045
+ $X2=0 $Y2=0
cc_859 N_A_867_82#_c_918_n N_A_1954_119#_c_1985_n 0.00335594f $X=9.84 $Y=1.665
+ $X2=0 $Y2=0
cc_860 N_A_867_82#_c_910_n N_A_1954_119#_c_1986_n 0.0426269f $X=10.835 $Y=1.41
+ $X2=0 $Y2=0
cc_861 N_A_867_82#_c_911_n N_A_1954_119#_c_1986_n 0.00310603f $X=10.835 $Y=1.41
+ $X2=0 $Y2=0
cc_862 N_A_867_82#_c_904_n N_A_1954_119#_c_1987_n 0.00104254f $X=9.83 $Y=2.045
+ $X2=0 $Y2=0
cc_863 N_A_867_82#_c_910_n N_A_1954_119#_c_1987_n 0.0125858f $X=10.835 $Y=1.41
+ $X2=0 $Y2=0
cc_864 N_A_867_82#_c_917_n N_A_1954_119#_c_1987_n 3.73484e-19 $X=9.84 $Y=1.665
+ $X2=0 $Y2=0
cc_865 N_A_867_82#_c_918_n N_A_1954_119#_c_1987_n 0.013985f $X=9.84 $Y=1.665
+ $X2=0 $Y2=0
cc_866 N_A_867_82#_M1039_g N_A_1954_119#_c_1978_n 0.0136417f $X=10.745 $Y=0.805
+ $X2=0 $Y2=0
cc_867 N_A_867_82#_c_911_n N_A_1954_119#_c_1978_n 0.00410729f $X=10.835 $Y=1.41
+ $X2=0 $Y2=0
cc_868 N_A_867_82#_M1039_g N_A_1954_119#_c_1979_n 0.00269838f $X=10.745 $Y=0.805
+ $X2=0 $Y2=0
cc_869 N_A_867_82#_c_910_n N_A_1954_119#_c_1979_n 0.0234153f $X=10.835 $Y=1.41
+ $X2=0 $Y2=0
cc_870 N_A_867_82#_c_911_n N_A_1954_119#_c_1979_n 0.00161194f $X=10.835 $Y=1.41
+ $X2=0 $Y2=0
cc_871 N_A_867_82#_c_904_n N_A_1954_119#_c_1996_n 0.00399114f $X=9.83 $Y=2.045
+ $X2=0 $Y2=0
cc_872 N_A_867_82#_c_910_n N_A_1954_119#_c_1996_n 0.00262016f $X=10.835 $Y=1.41
+ $X2=0 $Y2=0
cc_873 N_A_867_82#_c_918_n N_A_1954_119#_c_1996_n 0.011063f $X=9.84 $Y=1.665
+ $X2=0 $Y2=0
cc_874 N_A_867_82#_c_909_n N_A_1954_119#_c_2016_n 0.0240272f $X=10.07 $Y=1.407
+ $X2=0 $Y2=0
cc_875 N_A_867_82#_c_910_n N_A_1954_119#_c_2016_n 0.0712937f $X=10.835 $Y=1.41
+ $X2=0 $Y2=0
cc_876 N_A_867_82#_c_917_n N_A_1954_119#_c_2016_n 0.00104303f $X=9.84 $Y=1.665
+ $X2=0 $Y2=0
cc_877 N_A_867_82#_M1039_g N_A_1954_119#_c_2019_n 0.00859352f $X=10.745 $Y=0.805
+ $X2=0 $Y2=0
cc_878 N_A_867_82#_c_926_n N_VPWR_c_2279_n 0.0469739f $X=4.545 $Y=2.815 $X2=0
+ $Y2=0
cc_879 N_A_867_82#_c_926_n N_VPWR_c_2280_n 0.0177173f $X=4.545 $Y=2.815 $X2=0
+ $Y2=0
cc_880 N_A_867_82#_c_923_n N_VPWR_c_2281_n 2.33331e-19 $X=5.72 $Y=2.41 $X2=0
+ $Y2=0
cc_881 N_A_867_82#_c_926_n N_VPWR_c_2281_n 0.0328665f $X=4.545 $Y=2.815 $X2=0
+ $Y2=0
cc_882 N_A_867_82#_c_904_n N_VPWR_c_2283_n 0.00197813f $X=9.83 $Y=2.045 $X2=0
+ $Y2=0
cc_883 N_A_867_82#_c_923_n N_VPWR_c_2286_n 8.63546e-19 $X=5.72 $Y=2.41 $X2=0
+ $Y2=0
cc_884 N_A_867_82#_c_904_n N_VPWR_c_2289_n 0.00445602f $X=9.83 $Y=2.045 $X2=0
+ $Y2=0
cc_885 N_A_867_82#_c_904_n N_VPWR_c_2276_n 0.00858657f $X=9.83 $Y=2.045 $X2=0
+ $Y2=0
cc_886 N_A_867_82#_c_926_n N_VPWR_c_2276_n 0.0146319f $X=4.545 $Y=2.815 $X2=0
+ $Y2=0
cc_887 N_A_867_82#_M1016_d N_A_197_119#_c_2475_n 0.0112193f $X=4.335 $Y=0.41
+ $X2=0 $Y2=0
cc_888 N_A_867_82#_c_906_n N_A_197_119#_c_2475_n 0.0327192f $X=4.61 $Y=1.045
+ $X2=0 $Y2=0
cc_889 N_A_867_82#_c_906_n N_A_197_119#_c_2477_n 0.0205248f $X=4.61 $Y=1.045
+ $X2=0 $Y2=0
cc_890 N_A_867_82#_c_908_n N_A_197_119#_c_2477_n 0.00257141f $X=4.7 $Y=1.55
+ $X2=0 $Y2=0
cc_891 N_A_867_82#_c_914_n N_A_197_119#_c_2478_n 0.0130694f $X=6.38 $Y=1.635
+ $X2=0 $Y2=0
cc_892 N_A_867_82#_c_915_n N_A_197_119#_c_2478_n 0.00223165f $X=9.695 $Y=1.665
+ $X2=0 $Y2=0
cc_893 N_A_867_82#_c_916_n N_A_197_119#_c_2478_n 0.0079506f $X=5.665 $Y=1.665
+ $X2=0 $Y2=0
cc_894 N_A_867_82#_c_919_n N_A_197_119#_c_2478_n 0.00117358f $X=5.59 $Y=1.74
+ $X2=0 $Y2=0
cc_895 N_A_867_82#_c_920_n N_A_197_119#_c_2478_n 0.0462297f $X=5.405 $Y=1.727
+ $X2=0 $Y2=0
cc_896 N_A_867_82#_c_908_n N_A_197_119#_c_2479_n 0.013644f $X=4.7 $Y=1.55 $X2=0
+ $Y2=0
cc_897 N_A_867_82#_c_920_n N_A_197_119#_c_2479_n 0.0134395f $X=5.405 $Y=1.727
+ $X2=0 $Y2=0
cc_898 N_A_867_82#_M1001_g N_A_197_119#_c_2480_n 6.63727e-19 $X=6.47 $Y=0.805
+ $X2=0 $Y2=0
cc_899 N_A_867_82#_M1001_g N_A_197_119#_c_2481_n 0.00330666f $X=6.47 $Y=0.805
+ $X2=0 $Y2=0
cc_900 N_A_867_82#_M1001_g N_A_197_119#_c_2483_n 0.00753099f $X=6.47 $Y=0.805
+ $X2=0 $Y2=0
cc_901 N_A_867_82#_c_915_n N_A_197_119#_c_2493_n 0.00639031f $X=9.695 $Y=1.665
+ $X2=0 $Y2=0
cc_902 N_A_867_82#_c_915_n N_A_197_119#_c_2486_n 0.0232935f $X=9.695 $Y=1.665
+ $X2=0 $Y2=0
cc_903 N_A_867_82#_M1039_g N_VGND_c_2767_n 6.52646e-19 $X=10.745 $Y=0.805 $X2=0
+ $Y2=0
cc_904 N_A_867_82#_c_915_n N_A_1434_78#_c_2932_n 7.99965e-19 $X=9.695 $Y=1.665
+ $X2=0 $Y2=0
cc_905 N_A_1159_497#_c_1134_n N_A_1579_258#_c_1221_n 0.0164598f $X=7.565
+ $Y=2.045 $X2=0 $Y2=0
cc_906 N_A_1159_497#_c_1134_n N_A_1579_258#_c_1243_n 0.0452814f $X=7.565
+ $Y=2.045 $X2=0 $Y2=0
cc_907 N_A_1159_497#_c_1127_n N_A_1579_258#_M1047_g 0.0154495f $X=7.61 $Y=1.255
+ $X2=0 $Y2=0
cc_908 N_A_1159_497#_c_1126_n N_A_1579_258#_c_1238_n 0.0164598f $X=7.565
+ $Y=1.955 $X2=0 $Y2=0
cc_909 N_A_1159_497#_c_1128_n N_A_1579_258#_c_1238_n 0.00755082f $X=7.58 $Y=1.33
+ $X2=0 $Y2=0
cc_910 N_A_1159_497#_c_1129_n N_A_662_82#_M1017_g 6.98225e-19 $X=6.255 $Y=0.815
+ $X2=0 $Y2=0
cc_911 N_A_1159_497#_c_1138_n N_A_662_82#_c_1563_n 0.00563053f $X=6.03 $Y=2.055
+ $X2=0 $Y2=0
cc_912 N_A_1159_497#_c_1127_n N_A_662_82#_c_1564_n 0.00882199f $X=7.61 $Y=1.255
+ $X2=0 $Y2=0
cc_913 N_A_1159_497#_c_1138_n N_A_662_82#_c_1576_n 0.0111644f $X=6.03 $Y=2.055
+ $X2=0 $Y2=0
cc_914 N_A_1159_497#_c_1129_n N_A_662_82#_c_1569_n 3.2163e-19 $X=6.255 $Y=0.815
+ $X2=0 $Y2=0
cc_915 N_A_1159_497#_c_1131_n N_A_662_82#_c_1569_n 0.00154023f $X=6.42 $Y=1.215
+ $X2=0 $Y2=0
cc_916 N_A_1159_497#_c_1135_n N_A_662_82#_c_1578_n 0.0126178f $X=6.92 $Y=2.055
+ $X2=0 $Y2=0
cc_917 N_A_1159_497#_c_1138_n N_A_662_82#_c_1578_n 0.0102663f $X=6.03 $Y=2.055
+ $X2=0 $Y2=0
cc_918 N_A_1159_497#_c_1134_n N_VPWR_c_2286_n 0.00308634f $X=7.565 $Y=2.045
+ $X2=0 $Y2=0
cc_919 N_A_1159_497#_c_1134_n N_VPWR_c_2276_n 0.00387099f $X=7.565 $Y=2.045
+ $X2=0 $Y2=0
cc_920 N_A_1159_497#_c_1131_n N_A_197_119#_c_2478_n 0.00728887f $X=6.42 $Y=1.215
+ $X2=0 $Y2=0
cc_921 N_A_1159_497#_c_1129_n N_A_197_119#_c_2480_n 0.0199104f $X=6.255 $Y=0.815
+ $X2=0 $Y2=0
cc_922 N_A_1159_497#_c_1131_n N_A_197_119#_c_2480_n 0.00498269f $X=6.42 $Y=1.215
+ $X2=0 $Y2=0
cc_923 N_A_1159_497#_c_1129_n N_A_197_119#_c_2481_n 0.0168884f $X=6.255 $Y=0.815
+ $X2=0 $Y2=0
cc_924 N_A_1159_497#_c_1127_n N_A_197_119#_c_2483_n 0.00421599f $X=7.61 $Y=1.255
+ $X2=0 $Y2=0
cc_925 N_A_1159_497#_c_1134_n N_A_197_119#_c_2493_n 0.00811038f $X=7.565
+ $Y=2.045 $X2=0 $Y2=0
cc_926 N_A_1159_497#_c_1135_n N_A_197_119#_c_2493_n 0.0429823f $X=6.92 $Y=2.055
+ $X2=0 $Y2=0
cc_927 N_A_1159_497#_c_1132_n N_A_197_119#_c_2493_n 0.0013866f $X=7.085 $Y=1.42
+ $X2=0 $Y2=0
cc_928 N_A_1159_497#_c_1124_n N_A_197_119#_c_2484_n 0.00585102f $X=7.475 $Y=1.33
+ $X2=0 $Y2=0
cc_929 N_A_1159_497#_c_1125_n N_A_197_119#_c_2484_n 0.00165124f $X=7.25 $Y=1.33
+ $X2=0 $Y2=0
cc_930 N_A_1159_497#_c_1127_n N_A_197_119#_c_2484_n 0.00709647f $X=7.61 $Y=1.255
+ $X2=0 $Y2=0
cc_931 N_A_1159_497#_c_1130_n N_A_197_119#_c_2484_n 0.0271622f $X=6.92 $Y=1.215
+ $X2=0 $Y2=0
cc_932 N_A_1159_497#_c_1130_n N_A_197_119#_c_2485_n 0.0271042f $X=6.92 $Y=1.215
+ $X2=0 $Y2=0
cc_933 N_A_1159_497#_c_1124_n N_A_197_119#_c_2486_n 0.00397634f $X=7.475 $Y=1.33
+ $X2=0 $Y2=0
cc_934 N_A_1159_497#_c_1126_n N_A_197_119#_c_2486_n 0.0109871f $X=7.565 $Y=1.955
+ $X2=0 $Y2=0
cc_935 N_A_1159_497#_c_1134_n N_A_197_119#_c_2486_n 0.0112866f $X=7.565 $Y=2.045
+ $X2=0 $Y2=0
cc_936 N_A_1159_497#_c_1127_n N_A_197_119#_c_2486_n 0.00848228f $X=7.61 $Y=1.255
+ $X2=0 $Y2=0
cc_937 N_A_1159_497#_c_1128_n N_A_197_119#_c_2486_n 0.00391652f $X=7.58 $Y=1.33
+ $X2=0 $Y2=0
cc_938 N_A_1159_497#_c_1135_n N_A_197_119#_c_2486_n 0.0142943f $X=6.92 $Y=2.055
+ $X2=0 $Y2=0
cc_939 N_A_1159_497#_c_1130_n N_A_197_119#_c_2486_n 0.013938f $X=6.92 $Y=1.215
+ $X2=0 $Y2=0
cc_940 N_A_1159_497#_c_1136_n N_A_197_119#_c_2486_n 0.0490141f $X=7.085 $Y=1.42
+ $X2=0 $Y2=0
cc_941 N_A_1159_497#_c_1132_n N_A_197_119#_c_2486_n 0.00265527f $X=7.085 $Y=1.42
+ $X2=0 $Y2=0
cc_942 N_A_1159_497#_c_1135_n N_A_197_119#_c_2496_n 0.0246006f $X=6.92 $Y=2.055
+ $X2=0 $Y2=0
cc_943 N_A_1159_497#_c_1130_n N_A_1434_78#_M1003_s 0.00102398f $X=6.92 $Y=1.215
+ $X2=-0.19 $Y2=-0.245
cc_944 N_A_1159_497#_c_1127_n N_A_1434_78#_c_2931_n 0.00292741f $X=7.61 $Y=1.255
+ $X2=0 $Y2=0
cc_945 N_A_1159_497#_c_1124_n N_A_1434_78#_c_2933_n 3.7478e-19 $X=7.475 $Y=1.33
+ $X2=0 $Y2=0
cc_946 N_A_1159_497#_c_1127_n N_A_1434_78#_c_2933_n 0.00592285f $X=7.61 $Y=1.255
+ $X2=0 $Y2=0
cc_947 N_A_1579_258#_c_1243_n N_SET_B_c_1429_n 0.0266092f $X=7.985 $Y=2.045
+ $X2=-0.19 $Y2=-0.245
cc_948 N_A_1579_258#_M1047_g N_SET_B_M1025_g 0.0171555f $X=8.14 $Y=0.87 $X2=0
+ $Y2=0
cc_949 N_A_1579_258#_c_1226_n N_SET_B_M1025_g 0.0145937f $X=9.385 $Y=1.375 $X2=0
+ $Y2=0
cc_950 N_A_1579_258#_c_1237_n N_SET_B_M1025_g 0.00125218f $X=8.265 $Y=1.375
+ $X2=0 $Y2=0
cc_951 N_A_1579_258#_c_1238_n N_SET_B_M1025_g 0.0187498f $X=8.265 $Y=1.455 $X2=0
+ $Y2=0
cc_952 N_A_1579_258#_c_1225_n N_SET_B_c_1424_n 0.00751925f $X=12.47 $Y=1.795
+ $X2=0 $Y2=0
cc_953 N_A_1579_258#_c_1245_n N_SET_B_c_1424_n 0.0305873f $X=12.47 $Y=1.885
+ $X2=0 $Y2=0
cc_954 N_A_1579_258#_c_1232_n N_SET_B_c_1424_n 9.10537e-19 $X=12.2 $Y=1.215
+ $X2=0 $Y2=0
cc_955 N_A_1579_258#_c_1233_n N_SET_B_c_1424_n 3.87822e-19 $X=11.68 $Y=1.215
+ $X2=0 $Y2=0
cc_956 N_A_1579_258#_c_1223_n N_SET_B_M1007_g 0.0127442f $X=12.315 $Y=1.22 $X2=0
+ $Y2=0
cc_957 N_A_1579_258#_c_1224_n N_SET_B_M1007_g 0.0180591f $X=12.47 $Y=1.55 $X2=0
+ $Y2=0
cc_958 N_A_1579_258#_c_1230_n N_SET_B_M1007_g 0.00173868f $X=11.51 $Y=0.665
+ $X2=0 $Y2=0
cc_959 N_A_1579_258#_c_1231_n N_SET_B_M1007_g 0.00584413f $X=11.595 $Y=1.13
+ $X2=0 $Y2=0
cc_960 N_A_1579_258#_c_1232_n N_SET_B_M1007_g 0.0142422f $X=12.2 $Y=1.215 $X2=0
+ $Y2=0
cc_961 N_A_1579_258#_c_1240_n N_SET_B_M1007_g 0.00151951f $X=12.365 $Y=1.215
+ $X2=0 $Y2=0
cc_962 N_A_1579_258#_c_1221_n N_SET_B_c_1432_n 0.00223403f $X=7.985 $Y=1.955
+ $X2=0 $Y2=0
cc_963 N_A_1579_258#_c_1243_n N_SET_B_c_1432_n 0.00183509f $X=7.985 $Y=2.045
+ $X2=0 $Y2=0
cc_964 N_A_1579_258#_c_1237_n N_SET_B_c_1432_n 6.53774e-19 $X=8.265 $Y=1.375
+ $X2=0 $Y2=0
cc_965 N_A_1579_258#_c_1221_n N_SET_B_c_1426_n 0.00307141f $X=7.985 $Y=1.955
+ $X2=0 $Y2=0
cc_966 N_A_1579_258#_c_1243_n N_SET_B_c_1426_n 5.82953e-19 $X=7.985 $Y=2.045
+ $X2=0 $Y2=0
cc_967 N_A_1579_258#_c_1226_n N_SET_B_c_1426_n 0.0265376f $X=9.385 $Y=1.375
+ $X2=0 $Y2=0
cc_968 N_A_1579_258#_c_1237_n N_SET_B_c_1426_n 0.00953422f $X=8.265 $Y=1.375
+ $X2=0 $Y2=0
cc_969 N_A_1579_258#_c_1238_n N_SET_B_c_1426_n 7.33868e-19 $X=8.265 $Y=1.455
+ $X2=0 $Y2=0
cc_970 N_A_1579_258#_c_1233_n SET_B 7.57557e-19 $X=11.68 $Y=1.215 $X2=0 $Y2=0
cc_971 N_A_1579_258#_c_1221_n N_SET_B_c_1427_n 0.0116522f $X=7.985 $Y=1.955
+ $X2=0 $Y2=0
cc_972 N_A_1579_258#_c_1226_n N_SET_B_c_1427_n 0.00249882f $X=9.385 $Y=1.375
+ $X2=0 $Y2=0
cc_973 N_A_1579_258#_c_1238_n N_SET_B_c_1427_n 0.00469195f $X=8.265 $Y=1.455
+ $X2=0 $Y2=0
cc_974 N_A_1579_258#_c_1224_n N_SET_B_c_1428_n 2.99391e-19 $X=12.47 $Y=1.55
+ $X2=0 $Y2=0
cc_975 N_A_1579_258#_c_1225_n N_SET_B_c_1428_n 0.00130171f $X=12.47 $Y=1.795
+ $X2=0 $Y2=0
cc_976 N_A_1579_258#_c_1245_n N_SET_B_c_1428_n 0.00186247f $X=12.47 $Y=1.885
+ $X2=0 $Y2=0
cc_977 N_A_1579_258#_c_1232_n N_SET_B_c_1428_n 0.021621f $X=12.2 $Y=1.215 $X2=0
+ $Y2=0
cc_978 N_A_1579_258#_c_1233_n N_SET_B_c_1428_n 0.00427291f $X=11.68 $Y=1.215
+ $X2=0 $Y2=0
cc_979 N_A_1579_258#_c_1240_n N_SET_B_c_1428_n 0.00455765f $X=12.365 $Y=1.215
+ $X2=0 $Y2=0
cc_980 N_A_1579_258#_M1047_g N_A_662_82#_c_1564_n 0.00882199f $X=8.14 $Y=0.87
+ $X2=0 $Y2=0
cc_981 N_A_1579_258#_c_1229_n N_A_662_82#_c_1564_n 0.00340203f $X=9.555 $Y=0.45
+ $X2=0 $Y2=0
cc_982 N_A_1579_258#_c_1227_n N_A_662_82#_M1027_g 0.0106737f $X=9.47 $Y=1.29
+ $X2=0 $Y2=0
cc_983 N_A_1579_258#_c_1228_n N_A_662_82#_M1027_g 0.0167521f $X=10.75 $Y=0.45
+ $X2=0 $Y2=0
cc_984 N_A_1579_258#_c_1226_n N_A_662_82#_c_1567_n 7.12737e-19 $X=9.385 $Y=1.375
+ $X2=0 $Y2=0
cc_985 N_A_1579_258#_c_1230_n N_A_2133_410#_M1010_g 0.0118286f $X=11.51 $Y=0.665
+ $X2=0 $Y2=0
cc_986 N_A_1579_258#_c_1231_n N_A_2133_410#_M1010_g 0.00545777f $X=11.595
+ $Y=1.13 $X2=0 $Y2=0
cc_987 N_A_1579_258#_c_1233_n N_A_2133_410#_M1010_g 0.00142517f $X=11.68
+ $Y=1.215 $X2=0 $Y2=0
cc_988 N_A_1579_258#_c_1239_n N_A_2133_410#_M1010_g 0.00232774f $X=10.835
+ $Y=0.45 $X2=0 $Y2=0
cc_989 N_A_1579_258#_c_1248_n N_A_2133_410#_c_1743_n 2.06241e-19 $X=13.87
+ $Y=1.875 $X2=0 $Y2=0
cc_990 N_A_1579_258#_c_1245_n N_A_2133_410#_c_1764_n 0.0126852f $X=12.47
+ $Y=1.885 $X2=0 $Y2=0
cc_991 N_A_1579_258#_c_1234_n N_A_2133_410#_c_1749_n 0.0559136f $X=13.61
+ $Y=1.215 $X2=0 $Y2=0
cc_992 N_A_1579_258#_c_1236_n N_A_2133_410#_c_1749_n 0.0141315f $X=13.82 $Y=0.9
+ $X2=0 $Y2=0
cc_993 N_A_1579_258#_c_1245_n N_A_2133_410#_c_1766_n 8.73249e-19 $X=12.47
+ $Y=1.885 $X2=0 $Y2=0
cc_994 N_A_1579_258#_M1009_s N_A_2133_410#_c_1767_n 0.0104464f $X=13.6 $Y=1.73
+ $X2=0 $Y2=0
cc_995 N_A_1579_258#_c_1247_n N_A_2133_410#_c_1767_n 0.0138325f $X=13.78
+ $Y=1.915 $X2=0 $Y2=0
cc_996 N_A_1579_258#_c_1248_n N_A_2133_410#_c_1767_n 0.0260155f $X=13.87
+ $Y=1.875 $X2=0 $Y2=0
cc_997 N_A_1579_258#_c_1236_n N_A_2133_410#_c_1750_n 0.00886483f $X=13.82 $Y=0.9
+ $X2=0 $Y2=0
cc_998 N_A_1579_258#_c_1234_n N_A_2133_410#_c_1751_n 0.00517046f $X=13.61
+ $Y=1.215 $X2=0 $Y2=0
cc_999 N_A_1579_258#_c_1236_n N_A_2133_410#_c_1751_n 0.0130678f $X=13.82 $Y=0.9
+ $X2=0 $Y2=0
cc_1000 N_A_1579_258#_c_1236_n N_A_2133_410#_c_1753_n 0.0067812f $X=13.82 $Y=0.9
+ $X2=0 $Y2=0
cc_1001 N_A_1579_258#_c_1248_n N_A_2133_410#_c_1768_n 0.0106f $X=13.87 $Y=1.875
+ $X2=0 $Y2=0
cc_1002 N_A_1579_258#_c_1245_n N_A_2133_410#_c_1770_n 7.46086e-19 $X=12.47
+ $Y=1.885 $X2=0 $Y2=0
cc_1003 N_A_1579_258#_c_1223_n N_A_2133_410#_c_1794_n 0.0032332f $X=12.315
+ $Y=1.22 $X2=0 $Y2=0
cc_1004 N_A_1579_258#_c_1224_n N_A_2133_410#_c_1794_n 3.68822e-19 $X=12.47
+ $Y=1.55 $X2=0 $Y2=0
cc_1005 N_A_1579_258#_c_1234_n N_A_2133_410#_c_1794_n 0.0182618f $X=13.61
+ $Y=1.215 $X2=0 $Y2=0
cc_1006 N_A_1579_258#_c_1240_n N_A_2133_410#_c_1794_n 0.00533491f $X=12.365
+ $Y=1.215 $X2=0 $Y2=0
cc_1007 N_A_1579_258#_c_1236_n N_A_2133_410#_c_1755_n 0.00175799f $X=13.82
+ $Y=0.9 $X2=0 $Y2=0
cc_1008 N_A_1579_258#_c_1241_n N_A_2133_410#_c_1755_n 0.00193615f $X=13.82
+ $Y=1.215 $X2=0 $Y2=0
cc_1009 N_A_1579_258#_c_1223_n N_A_1954_119#_M1032_g 0.0234354f $X=12.315
+ $Y=1.22 $X2=0 $Y2=0
cc_1010 N_A_1579_258#_c_1224_n N_A_1954_119#_M1032_g 0.0222622f $X=12.47 $Y=1.55
+ $X2=0 $Y2=0
cc_1011 N_A_1579_258#_c_1234_n N_A_1954_119#_M1032_g 0.0123374f $X=13.61
+ $Y=1.215 $X2=0 $Y2=0
cc_1012 N_A_1579_258#_c_1235_n N_A_1954_119#_M1032_g 0.00339989f $X=13.695
+ $Y=1.79 $X2=0 $Y2=0
cc_1013 N_A_1579_258#_c_1240_n N_A_1954_119#_M1032_g 0.00122541f $X=12.365
+ $Y=1.215 $X2=0 $Y2=0
cc_1014 N_A_1579_258#_c_1225_n N_A_1954_119#_c_1977_n 0.0122908f $X=12.47
+ $Y=1.795 $X2=0 $Y2=0
cc_1015 N_A_1579_258#_c_1245_n N_A_1954_119#_c_1977_n 0.0561407f $X=12.47
+ $Y=1.885 $X2=0 $Y2=0
cc_1016 N_A_1579_258#_c_1234_n N_A_1954_119#_c_1977_n 0.011832f $X=13.61
+ $Y=1.215 $X2=0 $Y2=0
cc_1017 N_A_1579_258#_c_1247_n N_A_1954_119#_c_1977_n 0.0038005f $X=13.78
+ $Y=1.915 $X2=0 $Y2=0
cc_1018 N_A_1579_258#_c_1228_n N_A_1954_119#_c_1978_n 0.00537252f $X=10.75
+ $Y=0.45 $X2=0 $Y2=0
cc_1019 N_A_1579_258#_c_1230_n N_A_1954_119#_c_1978_n 0.0268263f $X=11.51
+ $Y=0.665 $X2=0 $Y2=0
cc_1020 N_A_1579_258#_c_1231_n N_A_1954_119#_c_1978_n 0.0134604f $X=11.595
+ $Y=1.13 $X2=0 $Y2=0
cc_1021 N_A_1579_258#_c_1239_n N_A_1954_119#_c_1978_n 0.00827962f $X=10.835
+ $Y=0.45 $X2=0 $Y2=0
cc_1022 N_A_1579_258#_c_1231_n N_A_1954_119#_c_1979_n 0.00278938f $X=11.595
+ $Y=1.13 $X2=0 $Y2=0
cc_1023 N_A_1579_258#_c_1233_n N_A_1954_119#_c_1979_n 0.0137331f $X=11.68
+ $Y=1.215 $X2=0 $Y2=0
cc_1024 N_A_1579_258#_c_1245_n N_A_1954_119#_c_1990_n 0.0154251f $X=12.47
+ $Y=1.885 $X2=0 $Y2=0
cc_1025 N_A_1579_258#_c_1245_n N_A_1954_119#_c_1992_n 0.00682041f $X=12.47
+ $Y=1.885 $X2=0 $Y2=0
cc_1026 N_A_1579_258#_c_1224_n N_A_1954_119#_c_1980_n 0.00142726f $X=12.47
+ $Y=1.55 $X2=0 $Y2=0
cc_1027 N_A_1579_258#_c_1225_n N_A_1954_119#_c_1980_n 0.00260476f $X=12.47
+ $Y=1.795 $X2=0 $Y2=0
cc_1028 N_A_1579_258#_c_1234_n N_A_1954_119#_c_1980_n 0.00797864f $X=13.61
+ $Y=1.215 $X2=0 $Y2=0
cc_1029 N_A_1579_258#_c_1240_n N_A_1954_119#_c_1980_n 0.00483544f $X=12.365
+ $Y=1.215 $X2=0 $Y2=0
cc_1030 N_A_1579_258#_c_1234_n N_A_1954_119#_c_1981_n 0.0499322f $X=13.61
+ $Y=1.215 $X2=0 $Y2=0
cc_1031 N_A_1579_258#_c_1235_n N_A_1954_119#_c_1981_n 0.0253541f $X=13.695
+ $Y=1.79 $X2=0 $Y2=0
cc_1032 N_A_1579_258#_c_1247_n N_A_1954_119#_c_1981_n 0.00888346f $X=13.78
+ $Y=1.915 $X2=0 $Y2=0
cc_1033 N_A_1579_258#_c_1235_n N_A_1954_119#_c_1982_n 0.00196834f $X=13.695
+ $Y=1.79 $X2=0 $Y2=0
cc_1034 N_A_1579_258#_c_1227_n N_A_1954_119#_c_2016_n 0.0276064f $X=9.47 $Y=1.29
+ $X2=0 $Y2=0
cc_1035 N_A_1579_258#_c_1228_n N_A_1954_119#_c_2016_n 0.0605317f $X=10.75
+ $Y=0.45 $X2=0 $Y2=0
cc_1036 N_A_1579_258#_c_1239_n N_A_1954_119#_c_2019_n 0.00347292f $X=10.835
+ $Y=0.45 $X2=0 $Y2=0
cc_1037 N_A_1579_258#_c_1236_n N_RESET_B_c_2121_n 0.0015566f $X=13.82 $Y=0.9
+ $X2=0 $Y2=0
cc_1038 N_A_1579_258#_c_1241_n N_RESET_B_c_2121_n 0.00474542f $X=13.82 $Y=1.215
+ $X2=0 $Y2=0
cc_1039 N_A_1579_258#_c_1248_n N_RESET_B_c_2126_n 0.00515371f $X=13.87 $Y=1.875
+ $X2=0 $Y2=0
cc_1040 N_A_1579_258#_c_1235_n N_RESET_B_c_2127_n 0.00399132f $X=13.695 $Y=1.79
+ $X2=0 $Y2=0
cc_1041 N_A_1579_258#_c_1248_n N_RESET_B_c_2127_n 0.00580189f $X=13.87 $Y=1.875
+ $X2=0 $Y2=0
cc_1042 N_A_1579_258#_c_1235_n RESET_B 0.0123764f $X=13.695 $Y=1.79 $X2=0 $Y2=0
cc_1043 N_A_1579_258#_c_1248_n RESET_B 0.00321191f $X=13.87 $Y=1.875 $X2=0 $Y2=0
cc_1044 N_A_1579_258#_c_1241_n RESET_B 0.00910445f $X=13.82 $Y=1.215 $X2=0 $Y2=0
cc_1045 N_A_1579_258#_c_1235_n N_RESET_B_c_2123_n 0.00507627f $X=13.695 $Y=1.79
+ $X2=0 $Y2=0
cc_1046 N_A_1579_258#_c_1248_n N_RESET_B_c_2123_n 0.00312216f $X=13.87 $Y=1.875
+ $X2=0 $Y2=0
cc_1047 N_A_1579_258#_c_1243_n N_VPWR_c_2282_n 0.0034565f $X=7.985 $Y=2.045
+ $X2=0 $Y2=0
cc_1048 N_A_1579_258#_c_1243_n N_VPWR_c_2286_n 0.00441521f $X=7.985 $Y=2.045
+ $X2=0 $Y2=0
cc_1049 N_A_1579_258#_c_1245_n N_VPWR_c_2297_n 0.00314375f $X=12.47 $Y=1.885
+ $X2=0 $Y2=0
cc_1050 N_A_1579_258#_c_1243_n N_VPWR_c_2276_n 0.00455667f $X=7.985 $Y=2.045
+ $X2=0 $Y2=0
cc_1051 N_A_1579_258#_c_1245_n N_VPWR_c_2276_n 0.00390476f $X=12.47 $Y=1.885
+ $X2=0 $Y2=0
cc_1052 N_A_1579_258#_c_1245_n N_VPWR_c_2305_n 0.00330333f $X=12.47 $Y=1.885
+ $X2=0 $Y2=0
cc_1053 N_A_1579_258#_c_1243_n N_A_197_119#_c_2486_n 2.45932e-19 $X=7.985
+ $Y=2.045 $X2=0 $Y2=0
cc_1054 N_A_1579_258#_c_1238_n N_A_197_119#_c_2486_n 7.29631e-19 $X=8.265
+ $Y=1.455 $X2=0 $Y2=0
cc_1055 N_A_1579_258#_c_1230_n N_VGND_M1010_d 0.00908674f $X=11.51 $Y=0.665
+ $X2=0 $Y2=0
cc_1056 N_A_1579_258#_c_1231_n N_VGND_M1010_d 0.00876391f $X=11.595 $Y=1.13
+ $X2=0 $Y2=0
cc_1057 N_A_1579_258#_c_1226_n N_VGND_c_2763_n 0.0197746f $X=9.385 $Y=1.375
+ $X2=0 $Y2=0
cc_1058 N_A_1579_258#_c_1227_n N_VGND_c_2763_n 0.0176968f $X=9.47 $Y=1.29 $X2=0
+ $Y2=0
cc_1059 N_A_1579_258#_c_1229_n N_VGND_c_2763_n 0.0111637f $X=9.555 $Y=0.45 $X2=0
+ $Y2=0
cc_1060 N_A_1579_258#_c_1230_n N_VGND_c_2766_n 0.0211619f $X=11.51 $Y=0.665
+ $X2=0 $Y2=0
cc_1061 N_A_1579_258#_c_1239_n N_VGND_c_2766_n 0.00170752f $X=10.835 $Y=0.45
+ $X2=0 $Y2=0
cc_1062 N_A_1579_258#_c_1228_n N_VGND_c_2767_n 0.0451243f $X=10.75 $Y=0.45 $X2=0
+ $Y2=0
cc_1063 N_A_1579_258#_c_1229_n N_VGND_c_2767_n 0.0071486f $X=9.555 $Y=0.45 $X2=0
+ $Y2=0
cc_1064 N_A_1579_258#_c_1230_n N_VGND_c_2767_n 0.00989656f $X=11.51 $Y=0.665
+ $X2=0 $Y2=0
cc_1065 N_A_1579_258#_c_1239_n N_VGND_c_2767_n 0.00678948f $X=10.835 $Y=0.45
+ $X2=0 $Y2=0
cc_1066 N_A_1579_258#_c_1223_n N_VGND_c_2774_n 0.00278247f $X=12.315 $Y=1.22
+ $X2=0 $Y2=0
cc_1067 N_A_1579_258#_c_1223_n N_VGND_c_2776_n 0.00354476f $X=12.315 $Y=1.22
+ $X2=0 $Y2=0
cc_1068 N_A_1579_258#_c_1228_n N_VGND_c_2776_n 0.0408085f $X=10.75 $Y=0.45 $X2=0
+ $Y2=0
cc_1069 N_A_1579_258#_c_1229_n N_VGND_c_2776_n 0.00553982f $X=9.555 $Y=0.45
+ $X2=0 $Y2=0
cc_1070 N_A_1579_258#_c_1230_n N_VGND_c_2776_n 0.0160771f $X=11.51 $Y=0.665
+ $X2=0 $Y2=0
cc_1071 N_A_1579_258#_c_1239_n N_VGND_c_2776_n 0.00603183f $X=10.835 $Y=0.45
+ $X2=0 $Y2=0
cc_1072 N_A_1579_258#_M1047_g N_A_1434_78#_c_2931_n 0.00330666f $X=8.14 $Y=0.87
+ $X2=0 $Y2=0
cc_1073 N_A_1579_258#_M1047_g N_A_1434_78#_c_2932_n 0.00697407f $X=8.14 $Y=0.87
+ $X2=0 $Y2=0
cc_1074 N_A_1579_258#_c_1226_n N_A_1434_78#_c_2932_n 0.010602f $X=9.385 $Y=1.375
+ $X2=0 $Y2=0
cc_1075 N_A_1579_258#_c_1237_n N_A_1434_78#_c_2932_n 0.0107488f $X=8.265
+ $Y=1.375 $X2=0 $Y2=0
cc_1076 N_A_1579_258#_c_1238_n N_A_1434_78#_c_2932_n 0.00125757f $X=8.265
+ $Y=1.455 $X2=0 $Y2=0
cc_1077 N_A_1579_258#_c_1227_n A_1876_119# 0.0076632f $X=9.47 $Y=1.29 $X2=-0.19
+ $Y2=-0.245
cc_1078 N_A_1579_258#_c_1230_n A_2164_119# 0.00300803f $X=11.51 $Y=0.665
+ $X2=-0.19 $Y2=-0.245
cc_1079 N_A_1579_258#_c_1239_n A_2164_119# 7.94081e-19 $X=10.835 $Y=0.45
+ $X2=-0.19 $Y2=-0.245
cc_1080 N_A_1579_258#_c_1223_n N_A_2392_74#_c_2967_n 0.00766753f $X=12.315
+ $Y=1.22 $X2=0 $Y2=0
cc_1081 N_A_1579_258#_c_1230_n N_A_2392_74#_c_2967_n 0.0102777f $X=11.51
+ $Y=0.665 $X2=0 $Y2=0
cc_1082 N_A_1579_258#_c_1231_n N_A_2392_74#_c_2967_n 0.0113279f $X=11.595
+ $Y=1.13 $X2=0 $Y2=0
cc_1083 N_A_1579_258#_c_1232_n N_A_2392_74#_c_2967_n 0.0183216f $X=12.2 $Y=1.215
+ $X2=0 $Y2=0
cc_1084 N_A_1579_258#_c_1240_n N_A_2392_74#_c_2967_n 0.00362226f $X=12.365
+ $Y=1.215 $X2=0 $Y2=0
cc_1085 N_A_1579_258#_c_1223_n N_A_2392_74#_c_2964_n 0.0105461f $X=12.315
+ $Y=1.22 $X2=0 $Y2=0
cc_1086 N_A_1579_258#_c_1223_n N_A_2392_74#_c_2965_n 0.00184341f $X=12.315
+ $Y=1.22 $X2=0 $Y2=0
cc_1087 N_SET_B_M1025_g N_A_662_82#_c_1564_n 0.0103107f $X=8.745 $Y=0.87 $X2=0
+ $Y2=0
cc_1088 N_SET_B_c_1431_n N_A_662_82#_c_1577_n 6.68077e-19 $X=11.615 $Y=2.035
+ $X2=0 $Y2=0
cc_1089 N_SET_B_c_1431_n N_A_662_82#_c_1570_n 0.00269682f $X=11.615 $Y=2.035
+ $X2=0 $Y2=0
cc_1090 N_SET_B_c_1431_n N_A_2133_410#_M1042_s 0.00641195f $X=11.615 $Y=2.035
+ $X2=0 $Y2=0
cc_1091 SET_B N_A_2133_410#_M1042_s 0.00176403f $X=11.675 $Y=1.95 $X2=0 $Y2=0
cc_1092 N_SET_B_c_1428_n N_A_2133_410#_M1042_s 0.00164634f $X=11.795 $Y=1.635
+ $X2=0 $Y2=0
cc_1093 N_SET_B_c_1431_n N_A_2133_410#_c_1756_n 0.0013917f $X=11.615 $Y=2.035
+ $X2=0 $Y2=0
cc_1094 N_SET_B_c_1431_n N_A_2133_410#_c_1757_n 0.00432177f $X=11.615 $Y=2.035
+ $X2=0 $Y2=0
cc_1095 SET_B N_A_2133_410#_c_1757_n 7.53207e-19 $X=11.675 $Y=1.95 $X2=0 $Y2=0
cc_1096 N_SET_B_c_1424_n N_A_2133_410#_M1010_g 0.0252868f $X=11.85 $Y=1.885
+ $X2=0 $Y2=0
cc_1097 N_SET_B_M1007_g N_A_2133_410#_M1010_g 0.0214067f $X=11.885 $Y=0.74 $X2=0
+ $Y2=0
cc_1098 N_SET_B_c_1431_n N_A_2133_410#_M1010_g 0.00158114f $X=11.615 $Y=2.035
+ $X2=0 $Y2=0
cc_1099 SET_B N_A_2133_410#_M1010_g 6.80953e-19 $X=11.675 $Y=1.95 $X2=0 $Y2=0
cc_1100 N_SET_B_c_1428_n N_A_2133_410#_M1010_g 0.0031406f $X=11.795 $Y=1.635
+ $X2=0 $Y2=0
cc_1101 N_SET_B_c_1431_n N_A_2133_410#_c_1763_n 0.0215547f $X=11.615 $Y=2.035
+ $X2=0 $Y2=0
cc_1102 N_SET_B_c_1424_n N_A_2133_410#_c_1764_n 0.00834212f $X=11.85 $Y=1.885
+ $X2=0 $Y2=0
cc_1103 N_SET_B_c_1431_n N_A_2133_410#_c_1769_n 0.00617302f $X=11.615 $Y=2.035
+ $X2=0 $Y2=0
cc_1104 N_SET_B_c_1424_n N_A_2133_410#_c_1770_n 0.00451111f $X=11.85 $Y=1.885
+ $X2=0 $Y2=0
cc_1105 N_SET_B_c_1431_n N_A_1954_119#_c_1985_n 0.0147602f $X=11.615 $Y=2.035
+ $X2=0 $Y2=0
cc_1106 N_SET_B_c_1431_n N_A_1954_119#_c_1986_n 0.030797f $X=11.615 $Y=2.035
+ $X2=0 $Y2=0
cc_1107 N_SET_B_c_1424_n N_A_1954_119#_c_1979_n 9.5198e-19 $X=11.85 $Y=1.885
+ $X2=0 $Y2=0
cc_1108 N_SET_B_M1007_g N_A_1954_119#_c_1979_n 0.00106933f $X=11.885 $Y=0.74
+ $X2=0 $Y2=0
cc_1109 N_SET_B_c_1428_n N_A_1954_119#_c_1979_n 0.0118597f $X=11.795 $Y=1.635
+ $X2=0 $Y2=0
cc_1110 N_SET_B_c_1424_n N_A_1954_119#_c_1989_n 0.00303048f $X=11.85 $Y=1.885
+ $X2=0 $Y2=0
cc_1111 N_SET_B_c_1431_n N_A_1954_119#_c_1989_n 0.0203237f $X=11.615 $Y=2.035
+ $X2=0 $Y2=0
cc_1112 SET_B N_A_1954_119#_c_1989_n 0.00279249f $X=11.675 $Y=1.95 $X2=0 $Y2=0
cc_1113 N_SET_B_c_1428_n N_A_1954_119#_c_1989_n 0.00866192f $X=11.795 $Y=1.635
+ $X2=0 $Y2=0
cc_1114 N_SET_B_c_1424_n N_A_1954_119#_c_1990_n 0.0135639f $X=11.85 $Y=1.885
+ $X2=0 $Y2=0
cc_1115 N_SET_B_c_1431_n N_A_1954_119#_c_1990_n 0.0121834f $X=11.615 $Y=2.035
+ $X2=0 $Y2=0
cc_1116 SET_B N_A_1954_119#_c_1990_n 0.00800669f $X=11.675 $Y=1.95 $X2=0 $Y2=0
cc_1117 N_SET_B_c_1428_n N_A_1954_119#_c_1990_n 0.0160506f $X=11.795 $Y=1.635
+ $X2=0 $Y2=0
cc_1118 N_SET_B_c_1428_n N_A_1954_119#_c_1992_n 0.00421876f $X=11.795 $Y=1.635
+ $X2=0 $Y2=0
cc_1119 N_SET_B_c_1428_n N_A_1954_119#_c_1980_n 0.00548815f $X=11.795 $Y=1.635
+ $X2=0 $Y2=0
cc_1120 N_SET_B_c_1431_n N_A_1954_119#_c_1996_n 0.0181235f $X=11.615 $Y=2.035
+ $X2=0 $Y2=0
cc_1121 N_SET_B_c_1424_n N_A_1954_119#_c_2064_n 3.76455e-19 $X=11.85 $Y=1.885
+ $X2=0 $Y2=0
cc_1122 N_SET_B_c_1428_n N_A_1954_119#_c_2064_n 0.00923927f $X=11.795 $Y=1.635
+ $X2=0 $Y2=0
cc_1123 N_SET_B_c_1432_n N_VPWR_M1022_d 0.00116601f $X=8.545 $Y=2.035 $X2=0
+ $Y2=0
cc_1124 N_SET_B_c_1426_n N_VPWR_M1022_d 2.64782e-19 $X=8.4 $Y=2.035 $X2=0 $Y2=0
cc_1125 N_SET_B_c_1429_n N_VPWR_c_2282_n 0.00373065f $X=8.435 $Y=2.045 $X2=0
+ $Y2=0
cc_1126 N_SET_B_c_1429_n N_VPWR_c_2283_n 0.00360601f $X=8.435 $Y=2.045 $X2=0
+ $Y2=0
cc_1127 N_SET_B_c_1431_n N_VPWR_c_2283_n 0.00140127f $X=11.615 $Y=2.035 $X2=0
+ $Y2=0
cc_1128 N_SET_B_c_1424_n N_VPWR_c_2288_n 0.00276611f $X=11.85 $Y=1.885 $X2=0
+ $Y2=0
cc_1129 N_SET_B_c_1429_n N_VPWR_c_2295_n 0.00445602f $X=8.435 $Y=2.045 $X2=0
+ $Y2=0
cc_1130 N_SET_B_c_1424_n N_VPWR_c_2296_n 0.00361132f $X=11.85 $Y=1.885 $X2=0
+ $Y2=0
cc_1131 N_SET_B_c_1429_n N_VPWR_c_2276_n 0.00459843f $X=8.435 $Y=2.045 $X2=0
+ $Y2=0
cc_1132 N_SET_B_c_1424_n N_VPWR_c_2276_n 0.00565696f $X=11.85 $Y=1.885 $X2=0
+ $Y2=0
cc_1133 N_SET_B_c_1424_n N_VPWR_c_2305_n 0.00326445f $X=11.85 $Y=1.885 $X2=0
+ $Y2=0
cc_1134 N_SET_B_M1025_g N_VGND_c_2763_n 0.0104746f $X=8.745 $Y=0.87 $X2=0 $Y2=0
cc_1135 N_SET_B_M1007_g N_VGND_c_2766_n 0.00395402f $X=11.885 $Y=0.74 $X2=0
+ $Y2=0
cc_1136 N_SET_B_M1007_g N_VGND_c_2774_n 0.00430908f $X=11.885 $Y=0.74 $X2=0
+ $Y2=0
cc_1137 N_SET_B_M1025_g N_VGND_c_2776_n 7.88961e-19 $X=8.745 $Y=0.87 $X2=0 $Y2=0
cc_1138 N_SET_B_M1007_g N_VGND_c_2776_n 0.00820779f $X=11.885 $Y=0.74 $X2=0
+ $Y2=0
cc_1139 N_SET_B_M1025_g N_A_1434_78#_c_2932_n 0.00595932f $X=8.745 $Y=0.87 $X2=0
+ $Y2=0
cc_1140 N_SET_B_M1007_g N_A_2392_74#_c_2967_n 0.00910416f $X=11.885 $Y=0.74
+ $X2=0 $Y2=0
cc_1141 N_SET_B_M1007_g N_A_2392_74#_c_2965_n 0.00386319f $X=11.885 $Y=0.74
+ $X2=0 $Y2=0
cc_1142 N_A_662_82#_c_1577_n N_A_2133_410#_c_1756_n 0.0494629f $X=10.365
+ $Y=2.465 $X2=0 $Y2=0
cc_1143 N_A_662_82#_c_1570_n N_A_2133_410#_c_1756_n 0.00743679f $X=10.365
+ $Y=2.18 $X2=0 $Y2=0
cc_1144 N_A_662_82#_c_1577_n N_A_2133_410#_c_1763_n 0.00184147f $X=10.365
+ $Y=2.465 $X2=0 $Y2=0
cc_1145 N_A_662_82#_c_1570_n N_A_2133_410#_c_1763_n 3.77136e-19 $X=10.365
+ $Y=2.18 $X2=0 $Y2=0
cc_1146 N_A_662_82#_c_1577_n N_A_1954_119#_c_1984_n 0.0116657f $X=10.365
+ $Y=2.465 $X2=0 $Y2=0
cc_1147 N_A_662_82#_c_1570_n N_A_1954_119#_c_1985_n 0.00854899f $X=10.365
+ $Y=2.18 $X2=0 $Y2=0
cc_1148 N_A_662_82#_c_1577_n N_A_1954_119#_c_1986_n 8.5645e-19 $X=10.365
+ $Y=2.465 $X2=0 $Y2=0
cc_1149 N_A_662_82#_c_1570_n N_A_1954_119#_c_1986_n 0.00488341f $X=10.365
+ $Y=2.18 $X2=0 $Y2=0
cc_1150 N_A_662_82#_c_1570_n N_A_1954_119#_c_1987_n 0.004329f $X=10.365 $Y=2.18
+ $X2=0 $Y2=0
cc_1151 N_A_662_82#_c_1577_n N_A_1954_119#_c_1996_n 0.00940235f $X=10.365
+ $Y=2.465 $X2=0 $Y2=0
cc_1152 N_A_662_82#_c_1570_n N_A_1954_119#_c_1996_n 0.00268164f $X=10.365
+ $Y=2.18 $X2=0 $Y2=0
cc_1153 N_A_662_82#_M1027_g N_A_1954_119#_c_2016_n 0.00528769f $X=9.695 $Y=0.87
+ $X2=0 $Y2=0
cc_1154 N_A_662_82#_c_1566_n N_A_1954_119#_c_2016_n 0.0144735f $X=10.28 $Y=1.295
+ $X2=0 $Y2=0
cc_1155 N_A_662_82#_c_1603_n N_VPWR_M1040_d 0.00330227f $X=3.97 $Y=2.035 $X2=0
+ $Y2=0
cc_1156 N_A_662_82#_c_1582_n N_VPWR_M1040_d 0.00110097f $X=4.055 $Y=1.95 $X2=0
+ $Y2=0
cc_1157 N_A_662_82#_c_1559_n N_VPWR_c_2279_n 0.00541579f $X=4.32 $Y=1.765 $X2=0
+ $Y2=0
cc_1158 N_A_662_82#_c_1581_n N_VPWR_c_2279_n 0.0453479f $X=3.645 $Y=2.815 $X2=0
+ $Y2=0
cc_1159 N_A_662_82#_c_1603_n N_VPWR_c_2279_n 0.0130547f $X=3.97 $Y=2.035 $X2=0
+ $Y2=0
cc_1160 N_A_662_82#_c_1573_n N_VPWR_c_2279_n 0.00131952f $X=4.335 $Y=1.505 $X2=0
+ $Y2=0
cc_1161 N_A_662_82#_c_1559_n N_VPWR_c_2280_n 0.00445602f $X=4.32 $Y=1.765 $X2=0
+ $Y2=0
cc_1162 N_A_662_82#_c_1559_n N_VPWR_c_2281_n 0.00323052f $X=4.32 $Y=1.765 $X2=0
+ $Y2=0
cc_1163 N_A_662_82#_c_1576_n N_VPWR_c_2286_n 8.63546e-19 $X=6.255 $Y=2.19 $X2=0
+ $Y2=0
cc_1164 N_A_662_82#_c_1577_n N_VPWR_c_2289_n 0.00461464f $X=10.365 $Y=2.465
+ $X2=0 $Y2=0
cc_1165 N_A_662_82#_c_1581_n N_VPWR_c_2294_n 0.011066f $X=3.645 $Y=2.815 $X2=0
+ $Y2=0
cc_1166 N_A_662_82#_c_1559_n N_VPWR_c_2276_n 0.00862475f $X=4.32 $Y=1.765 $X2=0
+ $Y2=0
cc_1167 N_A_662_82#_c_1577_n N_VPWR_c_2276_n 0.00979025f $X=10.365 $Y=2.465
+ $X2=0 $Y2=0
cc_1168 N_A_662_82#_c_1581_n N_VPWR_c_2276_n 0.00915947f $X=3.645 $Y=2.815 $X2=0
+ $Y2=0
cc_1169 N_A_662_82#_M1015_s N_A_197_119#_c_2472_n 2.83864e-19 $X=3.31 $Y=0.41
+ $X2=0 $Y2=0
cc_1170 N_A_662_82#_M1015_s N_A_197_119#_c_2474_n 0.00255936f $X=3.31 $Y=0.41
+ $X2=0 $Y2=0
cc_1171 N_A_662_82#_M1015_s N_A_197_119#_c_2475_n 0.00375964f $X=3.31 $Y=0.41
+ $X2=0 $Y2=0
cc_1172 N_A_662_82#_M1016_g N_A_197_119#_c_2475_n 0.0160561f $X=4.26 $Y=0.78
+ $X2=0 $Y2=0
cc_1173 N_A_662_82#_c_1560_n N_A_197_119#_c_2475_n 0.0133625f $X=5.965 $Y=0.18
+ $X2=0 $Y2=0
cc_1174 N_A_662_82#_c_1571_n N_A_197_119#_c_2475_n 0.045622f $X=3.97 $Y=1.045
+ $X2=0 $Y2=0
cc_1175 N_A_662_82#_c_1573_n N_A_197_119#_c_2475_n 0.00395718f $X=4.335 $Y=1.505
+ $X2=0 $Y2=0
cc_1176 N_A_662_82#_M1015_s N_A_197_119#_c_2476_n 0.00183565f $X=3.31 $Y=0.41
+ $X2=0 $Y2=0
cc_1177 N_A_662_82#_c_1571_n N_A_197_119#_c_2476_n 0.00902297f $X=3.97 $Y=1.045
+ $X2=0 $Y2=0
cc_1178 N_A_662_82#_M1016_g N_A_197_119#_c_2477_n 0.00438612f $X=4.26 $Y=0.78
+ $X2=0 $Y2=0
cc_1179 N_A_662_82#_c_1563_n N_A_197_119#_c_2478_n 0.0030348f $X=6.095 $Y=2.04
+ $X2=0 $Y2=0
cc_1180 N_A_662_82#_c_1569_n N_A_197_119#_c_2478_n 9.15821e-19 $X=6.067 $Y=1.24
+ $X2=0 $Y2=0
cc_1181 N_A_662_82#_M1017_g N_A_197_119#_c_2480_n 0.0122051f $X=6.04 $Y=0.805
+ $X2=0 $Y2=0
cc_1182 N_A_662_82#_c_1569_n N_A_197_119#_c_2480_n 0.00216694f $X=6.067 $Y=1.24
+ $X2=0 $Y2=0
cc_1183 N_A_662_82#_M1017_g N_A_197_119#_c_2481_n 0.0139343f $X=6.04 $Y=0.805
+ $X2=0 $Y2=0
cc_1184 N_A_662_82#_c_1564_n N_A_197_119#_c_2481_n 0.0148027f $X=9.62 $Y=0.18
+ $X2=0 $Y2=0
cc_1185 N_A_662_82#_c_1569_n N_A_197_119#_c_2481_n 0.00137036f $X=6.067 $Y=1.24
+ $X2=0 $Y2=0
cc_1186 N_A_662_82#_c_1560_n N_A_197_119#_c_2482_n 0.00321157f $X=5.965 $Y=0.18
+ $X2=0 $Y2=0
cc_1187 N_A_662_82#_M1017_g N_A_197_119#_c_2482_n 0.0030674f $X=6.04 $Y=0.805
+ $X2=0 $Y2=0
cc_1188 N_A_662_82#_M1017_g N_A_197_119#_c_2483_n 9.13855e-19 $X=6.04 $Y=0.805
+ $X2=0 $Y2=0
cc_1189 N_A_662_82#_c_1564_n N_A_197_119#_c_2484_n 0.0063797f $X=9.62 $Y=0.18
+ $X2=0 $Y2=0
cc_1190 N_A_662_82#_c_1571_n N_VGND_M1015_d 0.00602497f $X=3.97 $Y=1.045 $X2=0
+ $Y2=0
cc_1191 N_A_662_82#_c_1560_n N_VGND_c_2762_n 0.025796f $X=5.965 $Y=0.18 $X2=0
+ $Y2=0
cc_1192 N_A_662_82#_M1017_g N_VGND_c_2762_n 0.00150729f $X=6.04 $Y=0.805 $X2=0
+ $Y2=0
cc_1193 N_A_662_82#_c_1564_n N_VGND_c_2763_n 0.0257121f $X=9.62 $Y=0.18 $X2=0
+ $Y2=0
cc_1194 N_A_662_82#_M1027_g N_VGND_c_2763_n 0.00336259f $X=9.695 $Y=0.87 $X2=0
+ $Y2=0
cc_1195 N_A_662_82#_c_1564_n N_VGND_c_2767_n 0.0183446f $X=9.62 $Y=0.18 $X2=0
+ $Y2=0
cc_1196 N_A_662_82#_c_1561_n N_VGND_c_2772_n 0.0295884f $X=4.335 $Y=0.18 $X2=0
+ $Y2=0
cc_1197 N_A_662_82#_c_1560_n N_VGND_c_2773_n 0.0739828f $X=5.965 $Y=0.18 $X2=0
+ $Y2=0
cc_1198 N_A_662_82#_c_1560_n N_VGND_c_2776_n 0.0400687f $X=5.965 $Y=0.18 $X2=0
+ $Y2=0
cc_1199 N_A_662_82#_c_1561_n N_VGND_c_2776_n 0.00639767f $X=4.335 $Y=0.18 $X2=0
+ $Y2=0
cc_1200 N_A_662_82#_c_1564_n N_VGND_c_2776_n 0.0897088f $X=9.62 $Y=0.18 $X2=0
+ $Y2=0
cc_1201 N_A_662_82#_c_1568_n N_VGND_c_2776_n 0.00370845f $X=6.04 $Y=0.18 $X2=0
+ $Y2=0
cc_1202 N_A_662_82#_c_1561_n N_VGND_c_2778_n 0.0106531f $X=4.335 $Y=0.18 $X2=0
+ $Y2=0
cc_1203 N_A_662_82#_c_1564_n N_A_1434_78#_c_2931_n 0.0214634f $X=9.62 $Y=0.18
+ $X2=0 $Y2=0
cc_1204 N_A_662_82#_c_1564_n N_A_1434_78#_c_2933_n 0.00790476f $X=9.62 $Y=0.18
+ $X2=0 $Y2=0
cc_1205 N_A_2133_410#_c_1749_n N_A_1954_119#_M1032_g 0.0107193f $X=13.395
+ $Y=0.875 $X2=0 $Y2=0
cc_1206 N_A_2133_410#_c_1750_n N_A_1954_119#_M1032_g 0.00288279f $X=13.48
+ $Y=0.79 $X2=0 $Y2=0
cc_1207 N_A_2133_410#_c_1794_n N_A_1954_119#_M1032_g 0.0053774f $X=12.63
+ $Y=0.775 $X2=0 $Y2=0
cc_1208 N_A_2133_410#_c_1764_n N_A_1954_119#_c_1977_n 0.015744f $X=12.95
+ $Y=2.715 $X2=0 $Y2=0
cc_1209 N_A_2133_410#_c_1765_n N_A_1954_119#_c_1977_n 0.00321529f $X=13.115
+ $Y=2.38 $X2=0 $Y2=0
cc_1210 N_A_2133_410#_c_1766_n N_A_1954_119#_c_1977_n 0.00775623f $X=13.115
+ $Y=2.63 $X2=0 $Y2=0
cc_1211 N_A_2133_410#_c_1763_n N_A_1954_119#_c_1984_n 0.0120553f $X=10.83
+ $Y=2.215 $X2=0 $Y2=0
cc_1212 N_A_2133_410#_c_1756_n N_A_1954_119#_c_1985_n 3.1124e-19 $X=10.755
+ $Y=2.465 $X2=0 $Y2=0
cc_1213 N_A_2133_410#_c_1763_n N_A_1954_119#_c_1985_n 0.00190817f $X=10.83
+ $Y=2.215 $X2=0 $Y2=0
cc_1214 N_A_2133_410#_c_1756_n N_A_1954_119#_c_1986_n 0.0079207f $X=10.755
+ $Y=2.465 $X2=0 $Y2=0
cc_1215 N_A_2133_410#_c_1763_n N_A_1954_119#_c_1986_n 0.0205428f $X=10.83
+ $Y=2.215 $X2=0 $Y2=0
cc_1216 N_A_2133_410#_M1010_g N_A_1954_119#_c_1978_n 0.00738916f $X=11.285
+ $Y=0.805 $X2=0 $Y2=0
cc_1217 N_A_2133_410#_M1010_g N_A_1954_119#_c_1979_n 0.0172882f $X=11.285
+ $Y=0.805 $X2=0 $Y2=0
cc_1218 N_A_2133_410#_c_1756_n N_A_1954_119#_c_1989_n 0.00200916f $X=10.755
+ $Y=2.465 $X2=0 $Y2=0
cc_1219 N_A_2133_410#_c_1757_n N_A_1954_119#_c_1989_n 0.00971252f $X=11.21
+ $Y=2.125 $X2=0 $Y2=0
cc_1220 N_A_2133_410#_M1010_g N_A_1954_119#_c_1989_n 0.00492998f $X=11.285
+ $Y=0.805 $X2=0 $Y2=0
cc_1221 N_A_2133_410#_c_1763_n N_A_1954_119#_c_1989_n 0.0157294f $X=10.83
+ $Y=2.215 $X2=0 $Y2=0
cc_1222 N_A_2133_410#_M1042_s N_A_1954_119#_c_1990_n 0.00612902f $X=11.48
+ $Y=1.96 $X2=0 $Y2=0
cc_1223 N_A_2133_410#_c_1757_n N_A_1954_119#_c_1990_n 8.86672e-19 $X=11.21
+ $Y=2.125 $X2=0 $Y2=0
cc_1224 N_A_2133_410#_c_1764_n N_A_1954_119#_c_1990_n 0.0119962f $X=12.95
+ $Y=2.715 $X2=0 $Y2=0
cc_1225 N_A_2133_410#_c_1769_n N_A_1954_119#_c_1990_n 0.0745666f $X=11.46
+ $Y=2.805 $X2=0 $Y2=0
cc_1226 N_A_2133_410#_c_1756_n N_A_1954_119#_c_1991_n 0.00253841f $X=10.755
+ $Y=2.465 $X2=0 $Y2=0
cc_1227 N_A_2133_410#_c_1763_n N_A_1954_119#_c_1991_n 0.0143582f $X=10.83
+ $Y=2.215 $X2=0 $Y2=0
cc_1228 N_A_2133_410#_c_1769_n N_A_1954_119#_c_1991_n 0.0138529f $X=11.46
+ $Y=2.805 $X2=0 $Y2=0
cc_1229 N_A_2133_410#_c_1765_n N_A_1954_119#_c_1981_n 0.0264498f $X=13.115
+ $Y=2.38 $X2=0 $Y2=0
cc_1230 N_A_2133_410#_c_1767_n N_A_1954_119#_c_1981_n 0.00832042f $X=14.55
+ $Y=2.295 $X2=0 $Y2=0
cc_1231 N_A_2133_410#_c_1765_n N_A_1954_119#_c_1982_n 0.00178065f $X=13.115
+ $Y=2.38 $X2=0 $Y2=0
cc_1232 N_A_2133_410#_c_1767_n N_A_1954_119#_c_1982_n 8.26924e-19 $X=14.55
+ $Y=2.295 $X2=0 $Y2=0
cc_1233 N_A_2133_410#_c_1756_n N_A_1954_119#_c_1996_n 6.12517e-19 $X=10.755
+ $Y=2.465 $X2=0 $Y2=0
cc_1234 N_A_2133_410#_c_1763_n N_A_1954_119#_c_1996_n 0.00945054f $X=10.83
+ $Y=2.215 $X2=0 $Y2=0
cc_1235 N_A_2133_410#_M1010_g N_A_1954_119#_c_2064_n 0.00749195f $X=11.285
+ $Y=0.805 $X2=0 $Y2=0
cc_1236 N_A_2133_410#_c_1743_n N_RESET_B_c_2124_n 0.00633653f $X=14.75 $Y=1.765
+ $X2=-0.19 $Y2=-0.245
cc_1237 N_A_2133_410#_c_1764_n N_RESET_B_c_2124_n 0.00888395f $X=12.95 $Y=2.715
+ $X2=-0.19 $Y2=-0.245
cc_1238 N_A_2133_410#_c_1766_n N_RESET_B_c_2124_n 0.00599781f $X=13.115 $Y=2.63
+ $X2=-0.19 $Y2=-0.245
cc_1239 N_A_2133_410#_c_1767_n N_RESET_B_c_2124_n 0.0139706f $X=14.55 $Y=2.295
+ $X2=-0.19 $Y2=-0.245
cc_1240 N_A_2133_410#_M1005_g N_RESET_B_c_2121_n 0.00795349f $X=14.785 $Y=0.74
+ $X2=0 $Y2=0
cc_1241 N_A_2133_410#_c_1750_n N_RESET_B_c_2121_n 0.00205775f $X=13.48 $Y=0.79
+ $X2=0 $Y2=0
cc_1242 N_A_2133_410#_c_1751_n N_RESET_B_c_2121_n 0.00536183f $X=14.075 $Y=0.415
+ $X2=0 $Y2=0
cc_1243 N_A_2133_410#_c_1753_n N_RESET_B_c_2121_n 0.00849055f $X=14.16 $Y=0.85
+ $X2=0 $Y2=0
cc_1244 N_A_2133_410#_c_1858_p N_RESET_B_c_2121_n 0.0057256f $X=14.245 $Y=0.935
+ $X2=0 $Y2=0
cc_1245 N_A_2133_410#_c_1755_n N_RESET_B_c_2121_n 0.00147532f $X=14.742 $Y=1.3
+ $X2=0 $Y2=0
cc_1246 N_A_2133_410#_c_1767_n N_RESET_B_c_2125_n 0.0131005f $X=14.55 $Y=2.295
+ $X2=0 $Y2=0
cc_1247 N_A_2133_410#_c_1768_n N_RESET_B_c_2125_n 0.00543223f $X=14.635 $Y=2.21
+ $X2=0 $Y2=0
cc_1248 N_A_2133_410#_c_1765_n N_RESET_B_c_2126_n 0.00321144f $X=13.115 $Y=2.38
+ $X2=0 $Y2=0
cc_1249 N_A_2133_410#_c_1767_n N_RESET_B_c_2126_n 0.00297501f $X=14.55 $Y=2.295
+ $X2=0 $Y2=0
cc_1250 N_A_2133_410#_c_1743_n N_RESET_B_c_2127_n 0.0242389f $X=14.75 $Y=1.765
+ $X2=0 $Y2=0
cc_1251 N_A_2133_410#_c_1754_n N_RESET_B_c_2127_n 0.00543223f $X=14.77 $Y=1.465
+ $X2=0 $Y2=0
cc_1252 N_A_2133_410#_c_1743_n RESET_B 2.70011e-19 $X=14.75 $Y=1.765 $X2=0 $Y2=0
cc_1253 N_A_2133_410#_c_1767_n RESET_B 0.00593338f $X=14.55 $Y=2.295 $X2=0 $Y2=0
cc_1254 N_A_2133_410#_c_1868_p RESET_B 0.0105326f $X=14.55 $Y=0.935 $X2=0 $Y2=0
cc_1255 N_A_2133_410#_c_1858_p RESET_B 0.011975f $X=14.245 $Y=0.935 $X2=0 $Y2=0
cc_1256 N_A_2133_410#_c_1755_n RESET_B 0.0282196f $X=14.742 $Y=1.3 $X2=0 $Y2=0
cc_1257 N_A_2133_410#_c_1743_n N_RESET_B_c_2123_n 0.0159788f $X=14.75 $Y=1.765
+ $X2=0 $Y2=0
cc_1258 N_A_2133_410#_M1005_g N_RESET_B_c_2123_n 0.00295361f $X=14.785 $Y=0.74
+ $X2=0 $Y2=0
cc_1259 N_A_2133_410#_c_1767_n N_RESET_B_c_2123_n 6.37448e-19 $X=14.55 $Y=2.295
+ $X2=0 $Y2=0
cc_1260 N_A_2133_410#_c_1868_p N_RESET_B_c_2123_n 0.00143975f $X=14.55 $Y=0.935
+ $X2=0 $Y2=0
cc_1261 N_A_2133_410#_c_1858_p N_RESET_B_c_2123_n 8.10892e-19 $X=14.245 $Y=0.935
+ $X2=0 $Y2=0
cc_1262 N_A_2133_410#_c_1755_n N_RESET_B_c_2123_n 0.00209477f $X=14.742 $Y=1.3
+ $X2=0 $Y2=0
cc_1263 N_A_2133_410#_M1019_g N_A_3078_384#_c_2174_n 0.0164933f $X=15.775
+ $Y=0.645 $X2=0 $Y2=0
cc_1264 N_A_2133_410#_c_1762_n N_A_3078_384#_c_2175_n 0.0145446f $X=15.76
+ $Y=1.845 $X2=0 $Y2=0
cc_1265 N_A_2133_410#_M1019_g N_A_3078_384#_c_2175_n 0.02144f $X=15.775 $Y=0.645
+ $X2=0 $Y2=0
cc_1266 N_A_2133_410#_c_1748_n N_A_3078_384#_c_2175_n 0.00719647f $X=15.76
+ $Y=1.435 $X2=0 $Y2=0
cc_1267 N_A_2133_410#_M1005_g N_A_3078_384#_c_2176_n 0.00156859f $X=14.785
+ $Y=0.74 $X2=0 $Y2=0
cc_1268 N_A_2133_410#_M1019_g N_A_3078_384#_c_2176_n 0.0200735f $X=15.775
+ $Y=0.645 $X2=0 $Y2=0
cc_1269 N_A_2133_410#_c_1743_n N_A_3078_384#_c_2177_n 0.00163064f $X=14.75
+ $Y=1.765 $X2=0 $Y2=0
cc_1270 N_A_2133_410#_c_1745_n N_A_3078_384#_c_2177_n 0.00603351f $X=15.67
+ $Y=1.435 $X2=0 $Y2=0
cc_1271 N_A_2133_410#_c_1746_n N_A_3078_384#_c_2177_n 0.00707001f $X=15.76
+ $Y=1.755 $X2=0 $Y2=0
cc_1272 N_A_2133_410#_c_1762_n N_A_3078_384#_c_2177_n 0.0191242f $X=15.76
+ $Y=1.845 $X2=0 $Y2=0
cc_1273 N_A_2133_410#_c_1748_n N_A_3078_384#_c_2177_n 3.77891e-19 $X=15.76
+ $Y=1.435 $X2=0 $Y2=0
cc_1274 N_A_2133_410#_M1019_g N_A_3078_384#_c_2178_n 0.00753093f $X=15.775
+ $Y=0.645 $X2=0 $Y2=0
cc_1275 N_A_2133_410#_c_1748_n N_A_3078_384#_c_2178_n 0.0110454f $X=15.76
+ $Y=1.435 $X2=0 $Y2=0
cc_1276 N_A_2133_410#_c_1745_n N_A_3078_384#_c_2179_n 0.0127506f $X=15.67
+ $Y=1.435 $X2=0 $Y2=0
cc_1277 N_A_2133_410#_M1019_g N_A_3078_384#_c_2179_n 0.00171099f $X=15.775
+ $Y=0.645 $X2=0 $Y2=0
cc_1278 N_A_2133_410#_c_1748_n N_A_3078_384#_c_2179_n 0.00259264f $X=15.76
+ $Y=1.435 $X2=0 $Y2=0
cc_1279 N_A_2133_410#_c_1763_n N_VPWR_M1024_d 0.00367914f $X=10.83 $Y=2.215
+ $X2=0 $Y2=0
cc_1280 N_A_2133_410#_c_1894_p N_VPWR_M1024_d 0.00117264f $X=10.995 $Y=2.715
+ $X2=0 $Y2=0
cc_1281 N_A_2133_410#_c_1769_n N_VPWR_M1024_d 0.00558167f $X=11.46 $Y=2.805
+ $X2=0 $Y2=0
cc_1282 N_A_2133_410#_c_1764_n N_VPWR_M1042_d 0.00848383f $X=12.95 $Y=2.715
+ $X2=0 $Y2=0
cc_1283 N_A_2133_410#_c_1767_n N_VPWR_M1009_d 0.0111157f $X=14.55 $Y=2.295 $X2=0
+ $Y2=0
cc_1284 N_A_2133_410#_c_1768_n N_VPWR_M1009_d 0.00450577f $X=14.635 $Y=2.21
+ $X2=0 $Y2=0
cc_1285 N_A_2133_410#_c_1743_n N_VPWR_c_2284_n 0.0143083f $X=14.75 $Y=1.765
+ $X2=0 $Y2=0
cc_1286 N_A_2133_410#_c_1767_n N_VPWR_c_2284_n 0.0471058f $X=14.55 $Y=2.295
+ $X2=0 $Y2=0
cc_1287 N_A_2133_410#_c_1762_n N_VPWR_c_2285_n 0.00937234f $X=15.76 $Y=1.845
+ $X2=0 $Y2=0
cc_1288 N_A_2133_410#_c_1756_n N_VPWR_c_2288_n 0.00522599f $X=10.755 $Y=2.465
+ $X2=0 $Y2=0
cc_1289 N_A_2133_410#_c_1894_p N_VPWR_c_2288_n 0.007614f $X=10.995 $Y=2.715
+ $X2=0 $Y2=0
cc_1290 N_A_2133_410#_c_1769_n N_VPWR_c_2288_n 0.0172102f $X=11.46 $Y=2.805
+ $X2=0 $Y2=0
cc_1291 N_A_2133_410#_c_1770_n N_VPWR_c_2288_n 6.08883e-19 $X=11.79 $Y=2.805
+ $X2=0 $Y2=0
cc_1292 N_A_2133_410#_c_1756_n N_VPWR_c_2289_n 0.00314257f $X=10.755 $Y=2.465
+ $X2=0 $Y2=0
cc_1293 N_A_2133_410#_c_1894_p N_VPWR_c_2289_n 0.00473541f $X=10.995 $Y=2.715
+ $X2=0 $Y2=0
cc_1294 N_A_2133_410#_c_1743_n N_VPWR_c_2290_n 0.00413917f $X=14.75 $Y=1.765
+ $X2=0 $Y2=0
cc_1295 N_A_2133_410#_c_1762_n N_VPWR_c_2290_n 0.00435405f $X=15.76 $Y=1.845
+ $X2=0 $Y2=0
cc_1296 N_A_2133_410#_c_1764_n N_VPWR_c_2296_n 0.00283195f $X=12.95 $Y=2.715
+ $X2=0 $Y2=0
cc_1297 N_A_2133_410#_c_1769_n N_VPWR_c_2296_n 0.00532338f $X=11.46 $Y=2.805
+ $X2=0 $Y2=0
cc_1298 N_A_2133_410#_c_1770_n N_VPWR_c_2296_n 0.013942f $X=11.79 $Y=2.805 $X2=0
+ $Y2=0
cc_1299 N_A_2133_410#_c_1764_n N_VPWR_c_2297_n 0.0256637f $X=12.95 $Y=2.715
+ $X2=0 $Y2=0
cc_1300 N_A_2133_410#_c_1756_n N_VPWR_c_2276_n 0.00393368f $X=10.755 $Y=2.465
+ $X2=0 $Y2=0
cc_1301 N_A_2133_410#_c_1743_n N_VPWR_c_2276_n 0.00822528f $X=14.75 $Y=1.765
+ $X2=0 $Y2=0
cc_1302 N_A_2133_410#_c_1762_n N_VPWR_c_2276_n 0.00484898f $X=15.76 $Y=1.845
+ $X2=0 $Y2=0
cc_1303 N_A_2133_410#_c_1894_p N_VPWR_c_2276_n 0.00756382f $X=10.995 $Y=2.715
+ $X2=0 $Y2=0
cc_1304 N_A_2133_410#_c_1764_n N_VPWR_c_2276_n 0.0350447f $X=12.95 $Y=2.715
+ $X2=0 $Y2=0
cc_1305 N_A_2133_410#_c_1769_n N_VPWR_c_2276_n 0.00845594f $X=11.46 $Y=2.805
+ $X2=0 $Y2=0
cc_1306 N_A_2133_410#_c_1770_n N_VPWR_c_2276_n 0.0118463f $X=11.79 $Y=2.805
+ $X2=0 $Y2=0
cc_1307 N_A_2133_410#_c_1764_n N_VPWR_c_2305_n 0.0244485f $X=12.95 $Y=2.715
+ $X2=0 $Y2=0
cc_1308 N_A_2133_410#_c_1770_n N_VPWR_c_2305_n 6.21521e-19 $X=11.79 $Y=2.805
+ $X2=0 $Y2=0
cc_1309 N_A_2133_410#_c_1764_n A_2509_392# 0.0040234f $X=12.95 $Y=2.715
+ $X2=-0.19 $Y2=-0.245
cc_1310 N_A_2133_410#_M1005_g N_Q_N_c_2701_n 0.00205269f $X=14.785 $Y=0.74 $X2=0
+ $Y2=0
cc_1311 N_A_2133_410#_M1019_g N_Q_N_c_2701_n 0.00305526f $X=15.775 $Y=0.645
+ $X2=0 $Y2=0
cc_1312 N_A_2133_410#_c_1745_n N_Q_N_c_2702_n 0.00674797f $X=15.67 $Y=1.435
+ $X2=0 $Y2=0
cc_1313 N_A_2133_410#_c_1754_n N_Q_N_c_2702_n 0.00152576f $X=14.77 $Y=1.465
+ $X2=0 $Y2=0
cc_1314 N_A_2133_410#_c_1755_n N_Q_N_c_2702_n 0.00403687f $X=14.742 $Y=1.3 $X2=0
+ $Y2=0
cc_1315 N_A_2133_410#_c_1743_n Q_N 0.00949462f $X=14.75 $Y=1.765 $X2=0 $Y2=0
cc_1316 N_A_2133_410#_c_1745_n Q_N 0.00683658f $X=15.67 $Y=1.435 $X2=0 $Y2=0
cc_1317 N_A_2133_410#_c_1762_n Q_N 0.00291719f $X=15.76 $Y=1.845 $X2=0 $Y2=0
cc_1318 N_A_2133_410#_c_1768_n Q_N 0.0291769f $X=14.635 $Y=2.21 $X2=0 $Y2=0
cc_1319 N_A_2133_410#_c_1754_n Q_N 0.00335008f $X=14.77 $Y=1.465 $X2=0 $Y2=0
cc_1320 N_A_2133_410#_c_1762_n Q_N 0.00203386f $X=15.76 $Y=1.845 $X2=0 $Y2=0
cc_1321 N_A_2133_410#_c_1767_n Q_N 0.0141678f $X=14.55 $Y=2.295 $X2=0 $Y2=0
cc_1322 N_A_2133_410#_c_1743_n N_Q_N_c_2703_n 0.00408557f $X=14.75 $Y=1.765
+ $X2=0 $Y2=0
cc_1323 N_A_2133_410#_M1005_g N_Q_N_c_2703_n 0.00232922f $X=14.785 $Y=0.74 $X2=0
+ $Y2=0
cc_1324 N_A_2133_410#_c_1745_n N_Q_N_c_2703_n 0.0199186f $X=15.67 $Y=1.435 $X2=0
+ $Y2=0
cc_1325 N_A_2133_410#_c_1746_n N_Q_N_c_2703_n 6.03663e-19 $X=15.76 $Y=1.755
+ $X2=0 $Y2=0
cc_1326 N_A_2133_410#_c_1768_n N_Q_N_c_2703_n 0.00541296f $X=14.635 $Y=2.21
+ $X2=0 $Y2=0
cc_1327 N_A_2133_410#_c_1754_n N_Q_N_c_2703_n 0.0240864f $X=14.77 $Y=1.465 $X2=0
+ $Y2=0
cc_1328 N_A_2133_410#_c_1755_n N_Q_N_c_2703_n 0.00465146f $X=14.742 $Y=1.3 $X2=0
+ $Y2=0
cc_1329 N_A_2133_410#_c_1762_n Q 4.88141e-19 $X=15.76 $Y=1.845 $X2=0 $Y2=0
cc_1330 N_A_2133_410#_c_1753_n N_VGND_M1002_d 0.00271078f $X=14.16 $Y=0.85 $X2=0
+ $Y2=0
cc_1331 N_A_2133_410#_c_1868_p N_VGND_M1002_d 0.0153873f $X=14.55 $Y=0.935 $X2=0
+ $Y2=0
cc_1332 N_A_2133_410#_c_1858_p N_VGND_M1002_d 6.76691e-19 $X=14.245 $Y=0.935
+ $X2=0 $Y2=0
cc_1333 N_A_2133_410#_c_1755_n N_VGND_M1002_d 0.00147664f $X=14.742 $Y=1.3 $X2=0
+ $Y2=0
cc_1334 N_A_2133_410#_c_1743_n N_VGND_c_2764_n 2.59535e-19 $X=14.75 $Y=1.765
+ $X2=0 $Y2=0
cc_1335 N_A_2133_410#_M1005_g N_VGND_c_2764_n 0.0118756f $X=14.785 $Y=0.74 $X2=0
+ $Y2=0
cc_1336 N_A_2133_410#_c_1751_n N_VGND_c_2764_n 0.014808f $X=14.075 $Y=0.415
+ $X2=0 $Y2=0
cc_1337 N_A_2133_410#_c_1753_n N_VGND_c_2764_n 0.0139251f $X=14.16 $Y=0.85 $X2=0
+ $Y2=0
cc_1338 N_A_2133_410#_c_1868_p N_VGND_c_2764_n 0.0204933f $X=14.55 $Y=0.935
+ $X2=0 $Y2=0
cc_1339 N_A_2133_410#_c_1754_n N_VGND_c_2764_n 3.81546e-19 $X=14.77 $Y=1.465
+ $X2=0 $Y2=0
cc_1340 N_A_2133_410#_M1019_g N_VGND_c_2765_n 0.00705068f $X=15.775 $Y=0.645
+ $X2=0 $Y2=0
cc_1341 N_A_2133_410#_M1010_g N_VGND_c_2767_n 0.00329274f $X=11.285 $Y=0.805
+ $X2=0 $Y2=0
cc_1342 N_A_2133_410#_M1005_g N_VGND_c_2768_n 0.00383152f $X=14.785 $Y=0.74
+ $X2=0 $Y2=0
cc_1343 N_A_2133_410#_M1019_g N_VGND_c_2768_n 0.00434272f $X=15.775 $Y=0.645
+ $X2=0 $Y2=0
cc_1344 N_A_2133_410#_c_1751_n N_VGND_c_2774_n 0.030562f $X=14.075 $Y=0.415
+ $X2=0 $Y2=0
cc_1345 N_A_2133_410#_c_1752_n N_VGND_c_2774_n 0.00819987f $X=13.565 $Y=0.415
+ $X2=0 $Y2=0
cc_1346 N_A_2133_410#_M1010_g N_VGND_c_2776_n 0.00477801f $X=11.285 $Y=0.805
+ $X2=0 $Y2=0
cc_1347 N_A_2133_410#_M1005_g N_VGND_c_2776_n 0.00762539f $X=14.785 $Y=0.74
+ $X2=0 $Y2=0
cc_1348 N_A_2133_410#_M1019_g N_VGND_c_2776_n 0.00826076f $X=15.775 $Y=0.645
+ $X2=0 $Y2=0
cc_1349 N_A_2133_410#_c_1749_n N_VGND_c_2776_n 0.00704509f $X=13.395 $Y=0.875
+ $X2=0 $Y2=0
cc_1350 N_A_2133_410#_c_1751_n N_VGND_c_2776_n 0.0246282f $X=14.075 $Y=0.415
+ $X2=0 $Y2=0
cc_1351 N_A_2133_410#_c_1752_n N_VGND_c_2776_n 0.00633735f $X=13.565 $Y=0.415
+ $X2=0 $Y2=0
cc_1352 N_A_2133_410#_c_1868_p N_VGND_c_2776_n 0.00687055f $X=14.55 $Y=0.935
+ $X2=0 $Y2=0
cc_1353 N_A_2133_410#_c_1749_n N_A_2392_74#_M1032_d 0.00839898f $X=13.395
+ $Y=0.875 $X2=0 $Y2=0
cc_1354 N_A_2133_410#_M1010_g N_A_2392_74#_c_2967_n 7.01141e-19 $X=11.285
+ $Y=0.805 $X2=0 $Y2=0
cc_1355 N_A_2133_410#_c_1794_n N_A_2392_74#_c_2967_n 0.0250008f $X=12.63
+ $Y=0.775 $X2=0 $Y2=0
cc_1356 N_A_2133_410#_M1038_d N_A_2392_74#_c_2964_n 0.00341039f $X=12.39 $Y=0.37
+ $X2=0 $Y2=0
cc_1357 N_A_2133_410#_c_1749_n N_A_2392_74#_c_2964_n 0.00397331f $X=13.395
+ $Y=0.875 $X2=0 $Y2=0
cc_1358 N_A_2133_410#_c_1794_n N_A_2392_74#_c_2964_n 0.0195324f $X=12.63
+ $Y=0.775 $X2=0 $Y2=0
cc_1359 N_A_2133_410#_c_1749_n N_A_2392_74#_c_2966_n 0.0185865f $X=13.395
+ $Y=0.875 $X2=0 $Y2=0
cc_1360 N_A_2133_410#_c_1750_n N_A_2392_74#_c_2966_n 0.00909745f $X=13.48
+ $Y=0.79 $X2=0 $Y2=0
cc_1361 N_A_2133_410#_c_1752_n N_A_2392_74#_c_2966_n 0.0145005f $X=13.565
+ $Y=0.415 $X2=0 $Y2=0
cc_1362 N_A_1954_119#_c_1982_n N_RESET_B_c_2123_n 0.00140212f $X=13.275 $Y=1.635
+ $X2=0 $Y2=0
cc_1363 N_A_1954_119#_c_1990_n N_VPWR_M1042_d 0.0183998f $X=12.61 $Y=2.375 $X2=0
+ $Y2=0
cc_1364 N_A_1954_119#_c_1984_n N_VPWR_c_2283_n 0.0156011f $X=10.055 $Y=2.815
+ $X2=0 $Y2=0
cc_1365 N_A_1954_119#_c_1984_n N_VPWR_c_2289_n 0.0146247f $X=10.055 $Y=2.815
+ $X2=0 $Y2=0
cc_1366 N_A_1954_119#_c_1977_n N_VPWR_c_2297_n 0.00361118f $X=12.89 $Y=1.885
+ $X2=0 $Y2=0
cc_1367 N_A_1954_119#_c_1977_n N_VPWR_c_2276_n 0.0056474f $X=12.89 $Y=1.885
+ $X2=0 $Y2=0
cc_1368 N_A_1954_119#_c_1984_n N_VPWR_c_2276_n 0.0120586f $X=10.055 $Y=2.815
+ $X2=0 $Y2=0
cc_1369 N_A_1954_119#_c_1990_n A_2509_392# 0.0022665f $X=12.61 $Y=2.375
+ $X2=-0.19 $Y2=-0.245
cc_1370 N_A_1954_119#_c_1992_n A_2509_392# 0.00483806f $X=12.695 $Y=2.29
+ $X2=-0.19 $Y2=-0.245
cc_1371 N_A_1954_119#_M1032_g N_VGND_c_2774_n 0.00278271f $X=12.845 $Y=0.74
+ $X2=0 $Y2=0
cc_1372 N_A_1954_119#_M1032_g N_VGND_c_2776_n 0.0035847f $X=12.845 $Y=0.74 $X2=0
+ $Y2=0
cc_1373 N_A_1954_119#_c_1978_n A_2164_119# 0.00308543f $X=11.17 $Y=1.005
+ $X2=-0.19 $Y2=-0.245
cc_1374 N_A_1954_119#_M1032_g N_A_2392_74#_c_2967_n 7.53527e-19 $X=12.845
+ $Y=0.74 $X2=0 $Y2=0
cc_1375 N_A_1954_119#_M1032_g N_A_2392_74#_c_2964_n 0.0110746f $X=12.845 $Y=0.74
+ $X2=0 $Y2=0
cc_1376 N_A_1954_119#_M1032_g N_A_2392_74#_c_2966_n 0.00150373f $X=12.845
+ $Y=0.74 $X2=0 $Y2=0
cc_1377 N_RESET_B_c_2124_n N_VPWR_c_2284_n 0.0295777f $X=13.94 $Y=2.245 $X2=0
+ $Y2=0
cc_1378 N_RESET_B_c_2125_n N_VPWR_c_2284_n 0.00168808f $X=14.185 $Y=2.17 $X2=0
+ $Y2=0
cc_1379 N_RESET_B_c_2124_n N_VPWR_c_2297_n 0.00413917f $X=13.94 $Y=2.245 $X2=0
+ $Y2=0
cc_1380 N_RESET_B_c_2124_n N_VPWR_c_2276_n 0.00822528f $X=13.94 $Y=2.245 $X2=0
+ $Y2=0
cc_1381 N_RESET_B_c_2121_n N_VGND_c_2764_n 3.74645e-19 $X=14.035 $Y=1.22 $X2=0
+ $Y2=0
cc_1382 N_RESET_B_c_2121_n N_VGND_c_2774_n 2.6303e-19 $X=14.035 $Y=1.22 $X2=0
+ $Y2=0
cc_1383 N_A_3078_384#_c_2175_n N_VPWR_c_2285_n 0.0104544f $X=16.295 $Y=1.765
+ $X2=0 $Y2=0
cc_1384 N_A_3078_384#_c_2177_n N_VPWR_c_2285_n 0.0567727f $X=15.535 $Y=2.065
+ $X2=0 $Y2=0
cc_1385 N_A_3078_384#_c_2178_n N_VPWR_c_2285_n 0.0124476f $X=16.225 $Y=1.385
+ $X2=0 $Y2=0
cc_1386 N_A_3078_384#_c_2177_n N_VPWR_c_2290_n 0.00602538f $X=15.535 $Y=2.065
+ $X2=0 $Y2=0
cc_1387 N_A_3078_384#_c_2175_n N_VPWR_c_2298_n 0.00445602f $X=16.295 $Y=1.765
+ $X2=0 $Y2=0
cc_1388 N_A_3078_384#_c_2175_n N_VPWR_c_2276_n 0.00865885f $X=16.295 $Y=1.765
+ $X2=0 $Y2=0
cc_1389 N_A_3078_384#_c_2177_n N_VPWR_c_2276_n 0.00799129f $X=15.535 $Y=2.065
+ $X2=0 $Y2=0
cc_1390 N_A_3078_384#_c_2176_n N_Q_N_c_2701_n 0.0695681f $X=15.56 $Y=0.645 $X2=0
+ $Y2=0
cc_1391 N_A_3078_384#_c_2177_n N_Q_N_c_2703_n 0.0970792f $X=15.535 $Y=2.065
+ $X2=0 $Y2=0
cc_1392 N_A_3078_384#_c_2179_n N_Q_N_c_2703_n 0.0252224f $X=15.587 $Y=1.385
+ $X2=0 $Y2=0
cc_1393 N_A_3078_384#_c_2174_n N_Q_c_2736_n 0.00596415f $X=16.285 $Y=1.22 $X2=0
+ $Y2=0
cc_1394 N_A_3078_384#_c_2174_n N_Q_c_2737_n 0.00232286f $X=16.285 $Y=1.22 $X2=0
+ $Y2=0
cc_1395 N_A_3078_384#_c_2178_n N_Q_c_2737_n 0.00244346f $X=16.225 $Y=1.385 $X2=0
+ $Y2=0
cc_1396 N_A_3078_384#_c_2175_n Q 0.00404161f $X=16.295 $Y=1.765 $X2=0 $Y2=0
cc_1397 N_A_3078_384#_c_2177_n Q 0.00190906f $X=15.535 $Y=2.065 $X2=0 $Y2=0
cc_1398 N_A_3078_384#_c_2178_n Q 0.00106936f $X=16.225 $Y=1.385 $X2=0 $Y2=0
cc_1399 N_A_3078_384#_c_2175_n Q 0.0116977f $X=16.295 $Y=1.765 $X2=0 $Y2=0
cc_1400 N_A_3078_384#_c_2174_n N_Q_c_2738_n 0.00402581f $X=16.285 $Y=1.22 $X2=0
+ $Y2=0
cc_1401 N_A_3078_384#_c_2175_n N_Q_c_2738_n 0.0153071f $X=16.295 $Y=1.765 $X2=0
+ $Y2=0
cc_1402 N_A_3078_384#_c_2178_n N_Q_c_2738_n 0.0262119f $X=16.225 $Y=1.385 $X2=0
+ $Y2=0
cc_1403 N_A_3078_384#_c_2174_n N_VGND_c_2765_n 0.00308058f $X=16.285 $Y=1.22
+ $X2=0 $Y2=0
cc_1404 N_A_3078_384#_c_2175_n N_VGND_c_2765_n 0.00218674f $X=16.295 $Y=1.765
+ $X2=0 $Y2=0
cc_1405 N_A_3078_384#_c_2176_n N_VGND_c_2765_n 0.0300684f $X=15.56 $Y=0.645
+ $X2=0 $Y2=0
cc_1406 N_A_3078_384#_c_2178_n N_VGND_c_2765_n 0.0211017f $X=16.225 $Y=1.385
+ $X2=0 $Y2=0
cc_1407 N_A_3078_384#_c_2176_n N_VGND_c_2768_n 0.0121098f $X=15.56 $Y=0.645
+ $X2=0 $Y2=0
cc_1408 N_A_3078_384#_c_2174_n N_VGND_c_2775_n 0.00434272f $X=16.285 $Y=1.22
+ $X2=0 $Y2=0
cc_1409 N_A_3078_384#_c_2174_n N_VGND_c_2776_n 0.00824802f $X=16.285 $Y=1.22
+ $X2=0 $Y2=0
cc_1410 N_A_3078_384#_c_2176_n N_VGND_c_2776_n 0.00996704f $X=15.56 $Y=0.645
+ $X2=0 $Y2=0
cc_1411 N_A_27_464#_c_2226_n N_VPWR_c_2277_n 0.0230969f $X=0.28 $Y=2.465 $X2=0
+ $Y2=0
cc_1412 N_A_27_464#_c_2227_n N_VPWR_c_2277_n 0.0225341f $X=1.065 $Y=2.13 $X2=0
+ $Y2=0
cc_1413 N_A_27_464#_c_2231_n N_VPWR_c_2277_n 0.0100772f $X=1.235 $Y=2.99 $X2=0
+ $Y2=0
cc_1414 N_A_27_464#_c_2230_n N_VPWR_c_2278_n 0.0121087f $X=1.915 $Y=2.99 $X2=0
+ $Y2=0
cc_1415 N_A_27_464#_c_2232_n N_VPWR_c_2278_n 0.0391859f $X=2.08 $Y=2.465 $X2=0
+ $Y2=0
cc_1416 N_A_27_464#_c_2226_n N_VPWR_c_2292_n 0.0124046f $X=0.28 $Y=2.465 $X2=0
+ $Y2=0
cc_1417 N_A_27_464#_c_2230_n N_VPWR_c_2293_n 0.0665233f $X=1.915 $Y=2.99 $X2=0
+ $Y2=0
cc_1418 N_A_27_464#_c_2231_n N_VPWR_c_2293_n 0.0121867f $X=1.235 $Y=2.99 $X2=0
+ $Y2=0
cc_1419 N_A_27_464#_c_2226_n N_VPWR_c_2276_n 0.0102675f $X=0.28 $Y=2.465 $X2=0
+ $Y2=0
cc_1420 N_A_27_464#_c_2230_n N_VPWR_c_2276_n 0.0370231f $X=1.915 $Y=2.99 $X2=0
+ $Y2=0
cc_1421 N_A_27_464#_c_2231_n N_VPWR_c_2276_n 0.00660921f $X=1.235 $Y=2.99 $X2=0
+ $Y2=0
cc_1422 N_A_27_464#_c_2229_n A_212_464# 0.00798279f $X=1.15 $Y=2.905 $X2=-0.19
+ $Y2=1.66
cc_1423 N_A_27_464#_c_2230_n A_212_464# 0.00141176f $X=1.915 $Y=2.99 $X2=-0.19
+ $Y2=1.66
cc_1424 N_A_27_464#_c_2230_n N_A_197_119#_M1023_d 0.00222494f $X=1.915 $Y=2.99
+ $X2=0 $Y2=0
cc_1425 N_A_27_464#_c_2229_n N_A_197_119#_c_2489_n 0.0249199f $X=1.15 $Y=2.905
+ $X2=0 $Y2=0
cc_1426 N_A_27_464#_c_2232_n N_A_197_119#_c_2489_n 0.0277921f $X=2.08 $Y=2.465
+ $X2=0 $Y2=0
cc_1427 N_A_27_464#_c_2230_n N_A_197_119#_c_2503_n 0.014415f $X=1.915 $Y=2.99
+ $X2=0 $Y2=0
cc_1428 N_A_27_464#_c_2232_n N_A_197_119#_c_2490_n 0.0176316f $X=2.08 $Y=2.465
+ $X2=0 $Y2=0
cc_1429 N_A_27_464#_c_2227_n N_A_197_119#_c_2491_n 0.00639283f $X=1.065 $Y=2.13
+ $X2=0 $Y2=0
cc_1430 N_A_27_464#_c_2227_n N_A_197_119#_c_2495_n 0.00357858f $X=1.065 $Y=2.13
+ $X2=0 $Y2=0
cc_1431 N_A_27_464#_c_2229_n N_A_197_119#_c_2495_n 0.00415978f $X=1.15 $Y=2.905
+ $X2=0 $Y2=0
cc_1432 N_VPWR_c_2284_n Q_N 0.031531f $X=14.525 $Y=2.685 $X2=0 $Y2=0
cc_1433 N_VPWR_c_2285_n Q_N 0.00658861f $X=16.07 $Y=2.065 $X2=0 $Y2=0
cc_1434 N_VPWR_c_2290_n Q_N 0.0170898f $X=15.905 $Y=3.33 $X2=0 $Y2=0
cc_1435 N_VPWR_c_2276_n Q_N 0.0141455f $X=16.56 $Y=3.33 $X2=0 $Y2=0
cc_1436 N_VPWR_c_2285_n Q 0.0728884f $X=16.07 $Y=2.065 $X2=0 $Y2=0
cc_1437 N_VPWR_c_2298_n Q 0.0159324f $X=16.56 $Y=3.33 $X2=0 $Y2=0
cc_1438 N_VPWR_c_2276_n Q 0.0131546f $X=16.56 $Y=3.33 $X2=0 $Y2=0
cc_1439 N_A_197_119#_c_2471_n N_VGND_M1034_d 0.00778935f $X=2.475 $Y=1.14 $X2=0
+ $Y2=0
cc_1440 N_A_197_119#_c_2475_n N_VGND_M1015_d 0.00736182f $X=4.96 $Y=0.665 $X2=0
+ $Y2=0
cc_1441 N_A_197_119#_c_2487_n N_VGND_c_2760_n 0.0145731f $X=1.125 $Y=0.805 $X2=0
+ $Y2=0
cc_1442 N_A_197_119#_c_2468_n N_VGND_c_2761_n 0.00476116f $X=1.985 $Y=1.225
+ $X2=0 $Y2=0
cc_1443 N_A_197_119#_c_2470_n N_VGND_c_2761_n 0.00507012f $X=2.39 $Y=1.225 $X2=0
+ $Y2=0
cc_1444 N_A_197_119#_c_2471_n N_VGND_c_2761_n 0.0420985f $X=2.475 $Y=1.14 $X2=0
+ $Y2=0
cc_1445 N_A_197_119#_c_2473_n N_VGND_c_2761_n 0.015038f $X=2.56 $Y=0.34 $X2=0
+ $Y2=0
cc_1446 N_A_197_119#_c_2487_n N_VGND_c_2761_n 0.00835434f $X=1.125 $Y=0.805
+ $X2=0 $Y2=0
cc_1447 N_A_197_119#_c_2488_n N_VGND_c_2761_n 0.00604377f $X=1.57 $Y=0.95 $X2=0
+ $Y2=0
cc_1448 N_A_197_119#_c_2543_n N_VGND_c_2761_n 0.0148586f $X=2.07 $Y=1.225 $X2=0
+ $Y2=0
cc_1449 N_A_197_119#_c_2475_n N_VGND_c_2762_n 0.0150383f $X=4.96 $Y=0.665 $X2=0
+ $Y2=0
cc_1450 N_A_197_119#_c_2477_n N_VGND_c_2762_n 0.0225585f $X=5.045 $Y=1.205 $X2=0
+ $Y2=0
cc_1451 N_A_197_119#_c_2478_n N_VGND_c_2762_n 0.0267213f $X=5.8 $Y=1.29 $X2=0
+ $Y2=0
cc_1452 N_A_197_119#_c_2480_n N_VGND_c_2762_n 0.0300896f $X=5.885 $Y=1.205 $X2=0
+ $Y2=0
cc_1453 N_A_197_119#_c_2482_n N_VGND_c_2762_n 0.0150377f $X=5.97 $Y=0.34 $X2=0
+ $Y2=0
cc_1454 N_A_197_119#_c_2487_n N_VGND_c_2770_n 0.00728556f $X=1.125 $Y=0.805
+ $X2=0 $Y2=0
cc_1455 N_A_197_119#_c_2472_n N_VGND_c_2771_n 0.0545651f $X=3.23 $Y=0.34 $X2=0
+ $Y2=0
cc_1456 N_A_197_119#_c_2473_n N_VGND_c_2771_n 0.0115893f $X=2.56 $Y=0.34 $X2=0
+ $Y2=0
cc_1457 N_A_197_119#_c_2475_n N_VGND_c_2771_n 0.00678815f $X=4.96 $Y=0.665 $X2=0
+ $Y2=0
cc_1458 N_A_197_119#_c_2475_n N_VGND_c_2772_n 0.0193121f $X=4.96 $Y=0.665 $X2=0
+ $Y2=0
cc_1459 N_A_197_119#_c_2481_n N_VGND_c_2773_n 0.0623318f $X=6.595 $Y=0.34 $X2=0
+ $Y2=0
cc_1460 N_A_197_119#_c_2482_n N_VGND_c_2773_n 0.0115566f $X=5.97 $Y=0.34 $X2=0
+ $Y2=0
cc_1461 N_A_197_119#_c_2472_n N_VGND_c_2776_n 0.0308464f $X=3.23 $Y=0.34 $X2=0
+ $Y2=0
cc_1462 N_A_197_119#_c_2473_n N_VGND_c_2776_n 0.00583135f $X=2.56 $Y=0.34 $X2=0
+ $Y2=0
cc_1463 N_A_197_119#_c_2475_n N_VGND_c_2776_n 0.0396781f $X=4.96 $Y=0.665 $X2=0
+ $Y2=0
cc_1464 N_A_197_119#_c_2481_n N_VGND_c_2776_n 0.0322209f $X=6.595 $Y=0.34 $X2=0
+ $Y2=0
cc_1465 N_A_197_119#_c_2482_n N_VGND_c_2776_n 0.00579705f $X=5.97 $Y=0.34 $X2=0
+ $Y2=0
cc_1466 N_A_197_119#_c_2484_n N_VGND_c_2776_n 0.008245f $X=7.42 $Y=0.875 $X2=0
+ $Y2=0
cc_1467 N_A_197_119#_c_2487_n N_VGND_c_2776_n 0.008876f $X=1.125 $Y=0.805 $X2=0
+ $Y2=0
cc_1468 N_A_197_119#_c_2488_n N_VGND_c_2776_n 0.00543829f $X=1.57 $Y=0.95 $X2=0
+ $Y2=0
cc_1469 N_A_197_119#_c_2472_n N_VGND_c_2778_n 0.00754448f $X=3.23 $Y=0.34 $X2=0
+ $Y2=0
cc_1470 N_A_197_119#_c_2475_n N_VGND_c_2778_n 0.0244835f $X=4.96 $Y=0.665 $X2=0
+ $Y2=0
cc_1471 N_A_197_119#_c_2488_n A_305_119# 0.00221924f $X=1.57 $Y=0.95 $X2=-0.19
+ $Y2=-0.245
cc_1472 N_A_197_119#_c_2484_n N_A_1434_78#_M1003_s 0.00748686f $X=7.42 $Y=0.875
+ $X2=-0.19 $Y2=-0.245
cc_1473 N_A_197_119#_c_2486_n N_A_1434_78#_M1003_s 0.00660774f $X=7.505 $Y=2.31
+ $X2=-0.19 $Y2=-0.245
cc_1474 N_A_197_119#_c_2484_n N_A_1434_78#_c_2931_n 0.00335832f $X=7.42 $Y=0.875
+ $X2=0 $Y2=0
cc_1475 N_A_197_119#_c_2481_n N_A_1434_78#_c_2933_n 0.0123493f $X=6.595 $Y=0.34
+ $X2=0 $Y2=0
cc_1476 N_A_197_119#_c_2483_n N_A_1434_78#_c_2933_n 0.0133141f $X=6.76 $Y=0.765
+ $X2=0 $Y2=0
cc_1477 N_A_197_119#_c_2484_n N_A_1434_78#_c_2933_n 0.0251076f $X=7.42 $Y=0.875
+ $X2=0 $Y2=0
cc_1478 N_Q_N_c_2701_n N_VGND_c_2764_n 0.0125413f $X=15 $Y=0.515 $X2=0 $Y2=0
cc_1479 N_Q_N_c_2701_n N_VGND_c_2768_n 0.0159743f $X=15 $Y=0.515 $X2=0 $Y2=0
cc_1480 N_Q_N_c_2701_n N_VGND_c_2776_n 0.0132221f $X=15 $Y=0.515 $X2=0 $Y2=0
cc_1481 N_Q_c_2736_n N_VGND_c_2765_n 0.0263278f $X=16.5 $Y=0.515 $X2=0 $Y2=0
cc_1482 N_Q_c_2736_n N_VGND_c_2775_n 0.0168145f $X=16.5 $Y=0.515 $X2=0 $Y2=0
cc_1483 N_Q_c_2736_n N_VGND_c_2776_n 0.0138527f $X=16.5 $Y=0.515 $X2=0 $Y2=0
cc_1484 N_VGND_c_2763_n N_A_1434_78#_c_2931_n 0.0131781f $X=8.96 $Y=0.845 $X2=0
+ $Y2=0
cc_1485 N_VGND_c_2773_n N_A_1434_78#_c_2931_n 0.0726971f $X=8.795 $Y=0 $X2=0
+ $Y2=0
cc_1486 N_VGND_c_2776_n N_A_1434_78#_c_2931_n 0.0375338f $X=16.56 $Y=0 $X2=0
+ $Y2=0
cc_1487 N_VGND_c_2763_n N_A_1434_78#_c_2932_n 0.0444227f $X=8.96 $Y=0.845 $X2=0
+ $Y2=0
cc_1488 N_VGND_c_2773_n N_A_1434_78#_c_2933_n 0.0213919f $X=8.795 $Y=0 $X2=0
+ $Y2=0
cc_1489 N_VGND_c_2776_n N_A_1434_78#_c_2933_n 0.0110564f $X=16.56 $Y=0 $X2=0
+ $Y2=0
cc_1490 N_VGND_c_2774_n N_A_2392_74#_c_2964_n 0.0449102f $X=14.415 $Y=0 $X2=0
+ $Y2=0
cc_1491 N_VGND_c_2776_n N_A_2392_74#_c_2964_n 0.0254396f $X=16.56 $Y=0 $X2=0
+ $Y2=0
cc_1492 N_VGND_c_2766_n N_A_2392_74#_c_2965_n 0.010829f $X=11.585 $Y=0 $X2=0
+ $Y2=0
cc_1493 N_VGND_c_2774_n N_A_2392_74#_c_2965_n 0.0235447f $X=14.415 $Y=0 $X2=0
+ $Y2=0
cc_1494 N_VGND_c_2776_n N_A_2392_74#_c_2965_n 0.0126131f $X=16.56 $Y=0 $X2=0
+ $Y2=0
cc_1495 N_VGND_c_2774_n N_A_2392_74#_c_2966_n 0.0169764f $X=14.415 $Y=0 $X2=0
+ $Y2=0
cc_1496 N_VGND_c_2776_n N_A_2392_74#_c_2966_n 0.00949237f $X=16.56 $Y=0 $X2=0
+ $Y2=0
