* File: sky130_fd_sc_hs__and2b_4.pex.spice
* Created: Tue Sep  1 19:55:03 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HS__AND2B_4%A_N 1 3 6 8
c33 6 0 8.90662e-20 $X=0.59 $Y=0.69
r34 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.58
+ $Y=1.615 $X2=0.58 $Y2=1.615
r35 8 12 4.88915 $w=3.28e-07 $l=1.4e-07 $layer=LI1_cond $X=0.72 $Y=1.615
+ $X2=0.58 $Y2=1.615
r36 4 11 38.5481 $w=3.01e-07 $l=1.72337e-07 $layer=POLY_cond $X=0.59 $Y=1.45
+ $X2=0.575 $Y2=1.615
r37 4 6 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=0.59 $Y=1.45 $X2=0.59
+ $Y2=0.69
r38 1 11 55.362 $w=3.01e-07 $l=3.07409e-07 $layer=POLY_cond $X=0.495 $Y=1.885
+ $X2=0.575 $Y2=1.615
r39 1 3 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=0.495 $Y=1.885
+ $X2=0.495 $Y2=2.46
.ends

.subckt PM_SKY130_FD_SC_HS__AND2B_4%B 3 5 7 8 9 11 12 14 17 19 20 23 24 28 29 36
c105 36 0 1.88563e-19 $X=2.47 $Y=1.385
c106 28 0 7.7817e-20 $X=2.16 $Y=1.295
c107 23 0 8.90662e-20 $X=1.14 $Y=1.52
r108 36 38 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.47 $Y=1.385
+ $X2=2.47 $Y2=1.55
r109 36 37 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.47
+ $Y=1.385 $X2=2.47 $Y2=1.385
r110 29 45 0.885984 $w=5.38e-07 $l=4e-08 $layer=LI1_cond $X=2.315 $Y=1.665
+ $X2=2.315 $Y2=1.705
r111 29 37 6.20189 $w=5.38e-07 $l=2.8e-07 $layer=LI1_cond $X=2.315 $Y=1.665
+ $X2=2.315 $Y2=1.385
r112 28 37 1.99346 $w=5.38e-07 $l=9e-08 $layer=LI1_cond $X=2.315 $Y=1.295
+ $X2=2.315 $Y2=1.385
r113 24 33 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.14 $Y=1.52
+ $X2=1.14 $Y2=1.355
r114 23 26 6.46067 $w=3.28e-07 $l=1.85e-07 $layer=LI1_cond $X=1.14 $Y=1.52
+ $X2=1.14 $Y2=1.705
r115 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.14
+ $Y=1.52 $X2=1.14 $Y2=1.52
r116 21 26 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.305 $Y=1.705
+ $X2=1.14 $Y2=1.705
r117 20 45 7.6426 $w=1.7e-07 $l=2.7e-07 $layer=LI1_cond $X=2.045 $Y=1.705
+ $X2=2.315 $Y2=1.705
r118 20 21 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=2.045 $Y=1.705
+ $X2=1.305 $Y2=1.705
r119 15 36 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.47 $Y=1.22
+ $X2=2.47 $Y2=1.385
r120 15 17 271.766 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=2.47 $Y=1.22
+ $X2=2.47 $Y2=0.69
r121 12 19 20.4101 $w=1.5e-07 $l=8.44097e-08 $layer=POLY_cond $X=2.435 $Y=2.045
+ $X2=2.415 $Y2=1.97
r122 12 14 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=2.435 $Y=2.045
+ $X2=2.435 $Y2=2.54
r123 11 19 20.4101 $w=1.5e-07 $l=9.08295e-08 $layer=POLY_cond $X=2.38 $Y=1.895
+ $X2=2.415 $Y2=1.97
r124 11 38 176.904 $w=1.5e-07 $l=3.45e-07 $layer=POLY_cond $X=2.38 $Y=1.895
+ $X2=2.38 $Y2=1.55
r125 8 19 5.30422 $w=1.5e-07 $l=1.1e-07 $layer=POLY_cond $X=2.305 $Y=1.97
+ $X2=2.415 $Y2=1.97
r126 8 9 125.628 $w=1.5e-07 $l=2.45e-07 $layer=POLY_cond $X=2.305 $Y=1.97
+ $X2=2.06 $Y2=1.97
r127 5 9 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.985 $Y=2.045
+ $X2=2.06 $Y2=1.97
r128 5 7 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=1.985 $Y=2.045
+ $X2=1.985 $Y2=2.54
r129 3 33 340.989 $w=1.5e-07 $l=6.65e-07 $layer=POLY_cond $X=1.09 $Y=0.69
+ $X2=1.09 $Y2=1.355
.ends

.subckt PM_SKY130_FD_SC_HS__AND2B_4%A_27_392# 1 2 7 9 10 11 12 14 15 17 19 20 22
+ 24 28 32 34 38 40 41 42 46
c96 46 0 2.91552e-20 $X=1.68 $Y=1.285
c97 42 0 1.88563e-19 $X=1.68 $Y=1.18
r98 46 48 17.2143 $w=2.52e-07 $l=9e-08 $layer=POLY_cond $X=1.68 $Y=1.285
+ $X2=1.59 $Y2=1.285
r99 45 46 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.68
+ $Y=1.285 $X2=1.68 $Y2=1.285
r100 42 45 3.66686 $w=3.28e-07 $l=1.05e-07 $layer=LI1_cond $X=1.68 $Y=1.18
+ $X2=1.68 $Y2=1.285
r101 39 40 3.60271 $w=1.7e-07 $l=2.28e-07 $layer=LI1_cond $X=0.54 $Y=1.18
+ $X2=0.312 $Y2=1.18
r102 38 42 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.515 $Y=1.18
+ $X2=1.68 $Y2=1.18
r103 38 39 63.6096 $w=1.68e-07 $l=9.75e-07 $layer=LI1_cond $X=1.515 $Y=1.18
+ $X2=0.54 $Y2=1.18
r104 34 36 29.8782 $w=2.68e-07 $l=7e-07 $layer=LI1_cond $X=0.22 $Y=2.115
+ $X2=0.22 $Y2=2.815
r105 32 41 7.33542 $w=2.68e-07 $l=1.35e-07 $layer=LI1_cond $X=0.22 $Y=2.085
+ $X2=0.22 $Y2=1.95
r106 32 34 1.28049 $w=2.68e-07 $l=3e-08 $layer=LI1_cond $X=0.22 $Y=2.085
+ $X2=0.22 $Y2=2.115
r107 30 40 3.03453 $w=3.12e-07 $l=1.79538e-07 $layer=LI1_cond $X=0.17 $Y=1.265
+ $X2=0.312 $Y2=1.18
r108 30 41 44.6898 $w=1.68e-07 $l=6.85e-07 $layer=LI1_cond $X=0.17 $Y=1.265
+ $X2=0.17 $Y2=1.95
r109 26 40 3.03453 $w=3.12e-07 $l=8.5e-08 $layer=LI1_cond $X=0.312 $Y=1.095
+ $X2=0.312 $Y2=1.18
r110 26 28 15.2467 $w=4.53e-07 $l=5.8e-07 $layer=LI1_cond $X=0.312 $Y=1.095
+ $X2=0.312 $Y2=0.515
r111 23 24 64.0957 $w=1.5e-07 $l=1.25e-07 $layer=POLY_cond $X=1.465 $Y=1.97
+ $X2=1.59 $Y2=1.97
r112 20 46 65.0317 $w=2.52e-07 $l=4.14367e-07 $layer=POLY_cond $X=2.02 $Y=1.12
+ $X2=1.68 $Y2=1.285
r113 20 22 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=2.02 $Y=1.12
+ $X2=2.02 $Y2=0.69
r114 19 24 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.59 $Y=1.895
+ $X2=1.59 $Y2=1.97
r115 18 48 14.904 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.59 $Y=1.45
+ $X2=1.59 $Y2=1.285
r116 18 19 228.181 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=1.59 $Y=1.45
+ $X2=1.59 $Y2=1.895
r117 15 48 14.904 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.59 $Y=1.12
+ $X2=1.59 $Y2=1.285
r118 15 17 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=1.59 $Y=1.12
+ $X2=1.59 $Y2=0.69
r119 12 23 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.465 $Y=2.045
+ $X2=1.465 $Y2=1.97
r120 12 14 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=1.465 $Y=2.045
+ $X2=1.465 $Y2=2.54
r121 10 23 38.4574 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.39 $Y=1.97
+ $X2=1.465 $Y2=1.97
r122 10 11 153.83 $w=1.5e-07 $l=3e-07 $layer=POLY_cond $X=1.39 $Y=1.97 $X2=1.09
+ $Y2=1.97
r123 7 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.015 $Y=2.045
+ $X2=1.09 $Y2=1.97
r124 7 9 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=1.015 $Y=2.045
+ $X2=1.015 $Y2=2.54
r125 2 36 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.96 $X2=0.27 $Y2=2.815
r126 2 34 400 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.96 $X2=0.27 $Y2=2.115
r127 1 28 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.23
+ $Y=0.37 $X2=0.375 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__AND2B_4%A_218_424# 1 2 3 12 14 16 19 21 23 24 26 27
+ 29 30 31 32 34 36 37 39 40 43 45 46 47 53 55 58 60 66 69 70
c176 69 0 2.91552e-20 $X=2.21 $Y=2.045
c177 60 0 5.78711e-20 $X=2.84 $Y=1.96
c178 14 0 7.7817e-20 $X=2.955 $Y=1.765
c179 12 0 7.14761e-20 $X=2.955 $Y=0.74
r180 76 77 0.595062 $w=4.05e-07 $l=5e-09 $layer=POLY_cond $X=3.855 $Y=1.475
+ $X2=3.86 $Y2=1.475
r181 67 76 15.4716 $w=4.05e-07 $l=1.3e-07 $layer=POLY_cond $X=3.725 $Y=1.475
+ $X2=3.855 $Y2=1.475
r182 67 74 38.084 $w=4.05e-07 $l=3.2e-07 $layer=POLY_cond $X=3.725 $Y=1.475
+ $X2=3.405 $Y2=1.475
r183 66 67 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=3.725
+ $Y=1.485 $X2=3.725 $Y2=1.485
r184 63 66 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=3.045 $Y=1.485
+ $X2=3.725 $Y2=1.485
r185 63 64 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=3.045
+ $Y=1.485 $X2=3.045 $Y2=1.485
r186 61 70 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.925 $Y=1.485
+ $X2=2.84 $Y2=1.485
r187 61 63 4.1907 $w=3.28e-07 $l=1.2e-07 $layer=LI1_cond $X=2.925 $Y=1.485
+ $X2=3.045 $Y2=1.485
r188 59 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.84 $Y=1.65
+ $X2=2.84 $Y2=1.485
r189 59 60 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=2.84 $Y=1.65
+ $X2=2.84 $Y2=1.96
r190 58 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.84 $Y=1.32
+ $X2=2.84 $Y2=1.485
r191 57 58 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=2.84 $Y=0.925
+ $X2=2.84 $Y2=1.32
r192 56 69 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.375 $Y=2.045
+ $X2=2.21 $Y2=2.045
r193 55 60 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.755 $Y=2.045
+ $X2=2.84 $Y2=1.96
r194 55 56 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=2.755 $Y=2.045
+ $X2=2.375 $Y2=2.045
r195 51 69 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.21 $Y=2.13
+ $X2=2.21 $Y2=2.045
r196 51 53 4.71454 $w=3.28e-07 $l=1.35e-07 $layer=LI1_cond $X=2.21 $Y=2.13
+ $X2=2.21 $Y2=2.265
r197 47 57 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.755 $Y=0.84
+ $X2=2.84 $Y2=0.925
r198 47 49 61.9786 $w=1.68e-07 $l=9.5e-07 $layer=LI1_cond $X=2.755 $Y=0.84
+ $X2=1.805 $Y2=0.84
r199 45 69 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.045 $Y=2.045
+ $X2=2.21 $Y2=2.045
r200 45 46 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=2.045 $Y=2.045
+ $X2=1.405 $Y2=2.045
r201 41 46 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.24 $Y=2.13
+ $X2=1.405 $Y2=2.045
r202 41 43 4.71454 $w=3.28e-07 $l=1.35e-07 $layer=LI1_cond $X=1.24 $Y=2.13
+ $X2=1.24 $Y2=2.265
r203 37 39 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=4.305 $Y=1.765
+ $X2=4.305 $Y2=2.4
r204 36 37 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=4.305 $Y=1.675
+ $X2=4.305 $Y2=1.765
r205 35 40 18.8402 $w=1.65e-07 $l=2.81425e-07 $layer=POLY_cond $X=4.305 $Y=1.425
+ $X2=4.215 $Y2=1.185
r206 35 36 97.1774 $w=1.8e-07 $l=2.5e-07 $layer=POLY_cond $X=4.305 $Y=1.425
+ $X2=4.305 $Y2=1.675
r207 32 40 18.8402 $w=1.65e-07 $l=7.5e-08 $layer=POLY_cond $X=4.29 $Y=1.185
+ $X2=4.215 $Y2=1.185
r208 32 34 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=4.29 $Y=1.185
+ $X2=4.29 $Y2=0.74
r209 31 77 30.1637 $w=4.05e-07 $l=2.53969e-07 $layer=POLY_cond $X=3.945 $Y=1.26
+ $X2=3.86 $Y2=1.475
r210 30 40 6.66866 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.215 $Y=1.26
+ $X2=4.215 $Y2=1.185
r211 30 31 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=4.215 $Y=1.26
+ $X2=3.945 $Y2=1.26
r212 27 77 26.1659 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=3.86 $Y=1.185
+ $X2=3.86 $Y2=1.475
r213 27 29 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=3.86 $Y=1.185
+ $X2=3.86 $Y2=0.74
r214 24 76 26.1659 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=3.855 $Y=1.765
+ $X2=3.855 $Y2=1.475
r215 24 26 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.855 $Y=1.765
+ $X2=3.855 $Y2=2.4
r216 21 74 26.1659 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=3.405 $Y=1.765
+ $X2=3.405 $Y2=1.475
r217 21 23 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.405 $Y=1.765
+ $X2=3.405 $Y2=2.4
r218 17 74 1.19012 $w=4.05e-07 $l=1e-08 $layer=POLY_cond $X=3.395 $Y=1.475
+ $X2=3.405 $Y2=1.475
r219 17 64 41.6543 $w=4.05e-07 $l=3.5e-07 $layer=POLY_cond $X=3.395 $Y=1.475
+ $X2=3.045 $Y2=1.475
r220 17 19 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=3.395 $Y=1.32
+ $X2=3.395 $Y2=0.74
r221 14 16 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.955 $Y=1.765
+ $X2=2.955 $Y2=2.4
r222 10 64 10.7111 $w=4.05e-07 $l=9e-08 $layer=POLY_cond $X=2.955 $Y=1.475
+ $X2=3.045 $Y2=1.475
r223 10 14 26.1659 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=2.955 $Y=1.475
+ $X2=2.955 $Y2=1.765
r224 10 12 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=2.955 $Y=1.32
+ $X2=2.955 $Y2=0.74
r225 3 53 300 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=2 $X=2.06
+ $Y=2.12 $X2=2.21 $Y2=2.265
r226 2 43 300 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=2 $X=1.09
+ $Y=2.12 $X2=1.24 $Y2=2.265
r227 1 49 182 $w=1.7e-07 $l=5.35444e-07 $layer=licon1_NDIFF $count=1 $X=1.665
+ $Y=0.37 $X2=1.805 $Y2=0.84
.ends

.subckt PM_SKY130_FD_SC_HS__AND2B_4%VPWR 1 2 3 4 5 18 20 24 26 30 34 36 38 42 44
+ 49 54 60 63 66 69 73
r79 72 73 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r80 69 70 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r81 66 67 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r82 63 64 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r83 61 64 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.68 $Y2=3.33
r84 60 61 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r85 58 73 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=4.56 $Y2=3.33
r86 58 70 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=3.6 $Y2=3.33
r87 57 58 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r88 55 69 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.795 $Y=3.33
+ $X2=3.63 $Y2=3.33
r89 55 57 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=3.795 $Y=3.33
+ $X2=4.08 $Y2=3.33
r90 54 72 4.76062 $w=1.7e-07 $l=2.17e-07 $layer=LI1_cond $X=4.365 $Y=3.33
+ $X2=4.582 $Y2=3.33
r91 54 57 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=4.365 $Y=3.33
+ $X2=4.08 $Y2=3.33
r92 53 70 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=3.6 $Y2=3.33
r93 53 67 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=2.64 $Y2=3.33
r94 52 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r95 50 66 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.895 $Y=3.33
+ $X2=2.73 $Y2=3.33
r96 50 52 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=2.895 $Y=3.33
+ $X2=3.12 $Y2=3.33
r97 49 69 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.465 $Y=3.33
+ $X2=3.63 $Y2=3.33
r98 49 52 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=3.465 $Y=3.33
+ $X2=3.12 $Y2=3.33
r99 47 61 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r100 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r101 44 60 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.555 $Y=3.33
+ $X2=0.72 $Y2=3.33
r102 44 46 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=0.555 $Y=3.33
+ $X2=0.24 $Y2=3.33
r103 42 67 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.4 $Y=3.33
+ $X2=2.64 $Y2=3.33
r104 42 64 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=2.4 $Y=3.33
+ $X2=1.68 $Y2=3.33
r105 38 41 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=4.53 $Y=1.985
+ $X2=4.53 $Y2=2.815
r106 36 72 3.00555 $w=3.3e-07 $l=1.07912e-07 $layer=LI1_cond $X=4.53 $Y=3.245
+ $X2=4.582 $Y2=3.33
r107 36 41 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=4.53 $Y=3.245
+ $X2=4.53 $Y2=2.815
r108 32 69 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.63 $Y=3.245
+ $X2=3.63 $Y2=3.33
r109 32 34 32.1287 $w=3.28e-07 $l=9.2e-07 $layer=LI1_cond $X=3.63 $Y=3.245
+ $X2=3.63 $Y2=2.325
r110 28 66 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.73 $Y=3.245
+ $X2=2.73 $Y2=3.33
r111 28 30 27.2396 $w=3.28e-07 $l=7.8e-07 $layer=LI1_cond $X=2.73 $Y=3.245
+ $X2=2.73 $Y2=2.465
r112 27 63 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.855 $Y=3.33
+ $X2=1.73 $Y2=3.33
r113 26 66 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.565 $Y=3.33
+ $X2=2.73 $Y2=3.33
r114 26 27 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=2.565 $Y=3.33
+ $X2=1.855 $Y2=3.33
r115 22 63 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.73 $Y=3.245
+ $X2=1.73 $Y2=3.33
r116 22 24 35.9562 $w=2.48e-07 $l=7.8e-07 $layer=LI1_cond $X=1.73 $Y=3.245
+ $X2=1.73 $Y2=2.465
r117 21 60 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.885 $Y=3.33
+ $X2=0.72 $Y2=3.33
r118 20 63 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.605 $Y=3.33
+ $X2=1.73 $Y2=3.33
r119 20 21 46.9733 $w=1.68e-07 $l=7.2e-07 $layer=LI1_cond $X=1.605 $Y=3.33
+ $X2=0.885 $Y2=3.33
r120 16 60 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.72 $Y=3.245
+ $X2=0.72 $Y2=3.33
r121 16 18 34.2241 $w=3.28e-07 $l=9.8e-07 $layer=LI1_cond $X=0.72 $Y=3.245
+ $X2=0.72 $Y2=2.265
r122 5 41 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=4.38
+ $Y=1.84 $X2=4.53 $Y2=2.815
r123 5 38 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=4.38
+ $Y=1.84 $X2=4.53 $Y2=1.985
r124 4 34 300 $w=1.7e-07 $l=5.54955e-07 $layer=licon1_PDIFF $count=2 $X=3.48
+ $Y=1.84 $X2=3.63 $Y2=2.325
r125 3 30 300 $w=1.7e-07 $l=4.41503e-07 $layer=licon1_PDIFF $count=2 $X=2.51
+ $Y=2.12 $X2=2.73 $Y2=2.465
r126 2 24 300 $w=1.7e-07 $l=4.13249e-07 $layer=licon1_PDIFF $count=2 $X=1.54
+ $Y=2.12 $X2=1.69 $Y2=2.465
r127 1 18 300 $w=1.7e-07 $l=3.72525e-07 $layer=licon1_PDIFF $count=2 $X=0.57
+ $Y=1.96 $X2=0.72 $Y2=2.265
.ends

.subckt PM_SKY130_FD_SC_HS__AND2B_4%X 1 2 3 4 15 17 19 21 22 23 27 30 33 35 37
+ 38 41 43 46
c83 43 0 1.47064e-19 $X=4.08 $Y=1.985
c84 30 0 1.63274e-19 $X=4.08 $Y=1.82
r85 45 46 9.26965 $w=2.28e-07 $l=1.85e-07 $layer=LI1_cond $X=4.56 $Y=1.48
+ $X2=4.56 $Y2=1.295
r86 44 46 7.2654 $w=2.28e-07 $l=1.45e-07 $layer=LI1_cond $X=4.56 $Y=1.15
+ $X2=4.56 $Y2=1.295
r87 37 45 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=4.445 $Y=1.565
+ $X2=4.56 $Y2=1.48
r88 37 38 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=4.445 $Y=1.565
+ $X2=4.165 $Y2=1.565
r89 36 41 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.16 $Y=1.065
+ $X2=4.035 $Y2=1.065
r90 35 44 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=4.445 $Y=1.065
+ $X2=4.56 $Y2=1.15
r91 35 36 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=4.445 $Y=1.065
+ $X2=4.16 $Y2=1.065
r92 31 43 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.08 $Y=1.99 $X2=4.08
+ $Y2=1.905
r93 31 33 53.8235 $w=1.68e-07 $l=8.25e-07 $layer=LI1_cond $X=4.08 $Y=1.99
+ $X2=4.08 $Y2=2.815
r94 30 43 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.08 $Y=1.82 $X2=4.08
+ $Y2=1.905
r95 29 38 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.08 $Y=1.65
+ $X2=4.165 $Y2=1.565
r96 29 30 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=4.08 $Y=1.65
+ $X2=4.08 $Y2=1.82
r97 25 41 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.035 $Y=0.98
+ $X2=4.035 $Y2=1.065
r98 25 27 21.4354 $w=2.48e-07 $l=4.65e-07 $layer=LI1_cond $X=4.035 $Y=0.98
+ $X2=4.035 $Y2=0.515
r99 24 40 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.265 $Y=1.905
+ $X2=3.18 $Y2=1.905
r100 23 43 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.995 $Y=1.905
+ $X2=4.08 $Y2=1.905
r101 23 24 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=3.995 $Y=1.905
+ $X2=3.265 $Y2=1.905
r102 21 41 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.91 $Y=1.065
+ $X2=4.035 $Y2=1.065
r103 21 22 42.0802 $w=1.68e-07 $l=6.45e-07 $layer=LI1_cond $X=3.91 $Y=1.065
+ $X2=3.265 $Y2=1.065
r104 17 40 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.18 $Y=1.99
+ $X2=3.18 $Y2=1.905
r105 17 19 53.8235 $w=1.68e-07 $l=8.25e-07 $layer=LI1_cond $X=3.18 $Y=1.99
+ $X2=3.18 $Y2=2.815
r106 13 22 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.18 $Y=0.98
+ $X2=3.265 $Y2=1.065
r107 13 15 30.3369 $w=1.68e-07 $l=4.65e-07 $layer=LI1_cond $X=3.18 $Y=0.98
+ $X2=3.18 $Y2=0.515
r108 4 43 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=3.93
+ $Y=1.84 $X2=4.08 $Y2=1.985
r109 4 33 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=3.93
+ $Y=1.84 $X2=4.08 $Y2=2.815
r110 3 40 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=3.03
+ $Y=1.84 $X2=3.18 $Y2=1.985
r111 3 19 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=3.03
+ $Y=1.84 $X2=3.18 $Y2=2.815
r112 2 27 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.935
+ $Y=0.37 $X2=4.075 $Y2=0.515
r113 1 15 91 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_NDIFF $count=2 $X=3.03
+ $Y=0.37 $X2=3.18 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__AND2B_4%VGND 1 2 3 4 17 21 25 27 29 31 33 38 43 49
+ 52 55 59
r69 58 59 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r70 55 56 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r71 52 53 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r72 49 50 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r73 47 59 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=4.56
+ $Y2=0
r74 47 56 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=3.6
+ $Y2=0
r75 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r76 44 55 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.695 $Y=0 $X2=3.57
+ $Y2=0
r77 44 46 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=3.695 $Y=0 $X2=4.08
+ $Y2=0
r78 43 58 4.70058 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=4.34 $Y=0 $X2=4.57
+ $Y2=0
r79 43 46 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=4.34 $Y=0 $X2=4.08
+ $Y2=0
r80 42 56 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=3.6
+ $Y2=0
r81 42 53 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=2.64
+ $Y2=0
r82 41 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r83 39 52 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.9 $Y=0 $X2=2.735
+ $Y2=0
r84 39 41 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=2.9 $Y=0 $X2=3.12
+ $Y2=0
r85 38 55 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.445 $Y=0 $X2=3.57
+ $Y2=0
r86 38 41 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=3.445 $Y=0 $X2=3.12
+ $Y2=0
r87 37 50 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r88 36 37 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r89 34 49 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.04 $Y=0 $X2=0.875
+ $Y2=0
r90 34 36 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=1.04 $Y=0 $X2=1.2
+ $Y2=0
r91 33 52 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.57 $Y=0 $X2=2.735
+ $Y2=0
r92 33 36 89.3797 $w=1.68e-07 $l=1.37e-06 $layer=LI1_cond $X=2.57 $Y=0 $X2=1.2
+ $Y2=0
r93 31 53 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.4 $Y=0 $X2=2.64
+ $Y2=0
r94 31 37 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=2.4 $Y=0 $X2=1.2
+ $Y2=0
r95 27 58 3.0656 $w=3.3e-07 $l=1.12916e-07 $layer=LI1_cond $X=4.505 $Y=0.085
+ $X2=4.57 $Y2=0
r96 27 29 19.5566 $w=3.28e-07 $l=5.6e-07 $layer=LI1_cond $X=4.505 $Y=0.085
+ $X2=4.505 $Y2=0.645
r97 23 55 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.57 $Y=0.085
+ $X2=3.57 $Y2=0
r98 23 25 25.8147 $w=2.48e-07 $l=5.6e-07 $layer=LI1_cond $X=3.57 $Y=0.085
+ $X2=3.57 $Y2=0.645
r99 19 52 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.735 $Y=0.085
+ $X2=2.735 $Y2=0
r100 19 21 14.4928 $w=3.28e-07 $l=4.15e-07 $layer=LI1_cond $X=2.735 $Y=0.085
+ $X2=2.735 $Y2=0.5
r101 15 49 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.875 $Y=0.085
+ $X2=0.875 $Y2=0
r102 15 17 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=0.875 $Y=0.085
+ $X2=0.875 $Y2=0.495
r103 4 29 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=4.365
+ $Y=0.37 $X2=4.505 $Y2=0.645
r104 3 25 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=3.47
+ $Y=0.37 $X2=3.61 $Y2=0.645
r105 2 21 182 $w=1.7e-07 $l=2.46577e-07 $layer=licon1_NDIFF $count=1 $X=2.545
+ $Y=0.37 $X2=2.735 $Y2=0.5
r106 1 17 91 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=2 $X=0.665
+ $Y=0.37 $X2=0.875 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_HS__AND2B_4%A_233_74# 1 2 7 10 12
c17 12 0 7.14761e-20 $X=2.235 $Y=0.5
r18 10 12 35.2648 $w=2.48e-07 $l=7.65e-07 $layer=LI1_cond $X=1.47 $Y=0.46
+ $X2=2.235 $Y2=0.46
r19 7 10 6.8199 $w=2.5e-07 $l=1.82071e-07 $layer=LI1_cond $X=1.34 $Y=0.585
+ $X2=1.47 $Y2=0.46
r20 7 9 2.81538 $w=2.6e-07 $l=6e-08 $layer=LI1_cond $X=1.34 $Y=0.585 $X2=1.34
+ $Y2=0.645
r21 2 12 182 $w=1.7e-07 $l=1.94422e-07 $layer=licon1_NDIFF $count=1 $X=2.095
+ $Y=0.37 $X2=2.235 $Y2=0.5
r22 1 9 182 $w=1.7e-07 $l=3.49821e-07 $layer=licon1_NDIFF $count=1 $X=1.165
+ $Y=0.37 $X2=1.335 $Y2=0.645
.ends

