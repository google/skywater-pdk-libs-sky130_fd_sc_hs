* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hs__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
M1000 a_437_74# A1 Y VNB nlowvt w=740000u l=150000u
+  ad=2.368e+11p pd=2.12e+06u as=2.072e+11p ps=2.04e+06u
M1001 VGND B1_N a_29_424# VNB nlowvt w=550000u l=150000u
+  ad=5.5275e+11p pd=4.59e+06u as=1.4575e+11p ps=1.63e+06u
M1002 VPWR B1_N a_29_424# VPB pshort w=840000u l=150000u
+  ad=6.006e+11p pd=5.13e+06u as=2.31e+11p ps=2.23e+06u
M1003 a_348_368# a_29_424# Y VPB pshort w=1.12e+06u l=150000u
+  ad=6.44e+11p pd=5.63e+06u as=3.08e+11p ps=2.79e+06u
M1004 a_348_368# A2 VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 Y a_29_424# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VPWR A1 a_348_368# VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VGND A2 a_437_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
