* File: sky130_fd_sc_hs__ha_2.pxi.spice
* Created: Tue Sep  1 20:06:35 2020
* 
x_PM_SKY130_FD_SC_HS__HA_2%B N_B_M1015_g N_B_M1002_g N_B_c_103_n N_B_M1007_g
+ N_B_c_104_n N_B_M1005_g N_B_c_105_n N_B_c_112_n N_B_c_106_n N_B_c_107_n
+ N_B_c_108_n N_B_c_118_p B B B B PM_SKY130_FD_SC_HS__HA_2%B
x_PM_SKY130_FD_SC_HS__HA_2%A N_A_M1009_g N_A_c_191_n N_A_M1003_g N_A_M1004_g
+ N_A_c_192_n N_A_M1012_g A N_A_c_190_n PM_SKY130_FD_SC_HS__HA_2%A
x_PM_SKY130_FD_SC_HS__HA_2%A_27_74# N_A_27_74#_M1015_s N_A_27_74#_M1002_d
+ N_A_27_74#_M1016_g N_A_27_74#_M1000_g N_A_27_74#_c_259_n N_A_27_74#_M1013_g
+ N_A_27_74#_M1001_g N_A_27_74#_c_260_n N_A_27_74#_M1017_g N_A_27_74#_M1008_g
+ N_A_27_74#_c_246_n N_A_27_74#_c_262_n N_A_27_74#_c_247_n N_A_27_74#_c_248_n
+ N_A_27_74#_c_249_n N_A_27_74#_c_250_n N_A_27_74#_c_251_n N_A_27_74#_c_252_n
+ N_A_27_74#_c_318_p N_A_27_74#_c_253_n N_A_27_74#_c_310_p N_A_27_74#_c_286_n
+ N_A_27_74#_c_254_n N_A_27_74#_c_288_n N_A_27_74#_c_255_n N_A_27_74#_c_256_n
+ N_A_27_74#_c_257_n N_A_27_74#_c_258_n PM_SKY130_FD_SC_HS__HA_2%A_27_74#
x_PM_SKY130_FD_SC_HS__HA_2%A_391_388# N_A_391_388#_M1016_s N_A_391_388#_M1005_d
+ N_A_391_388#_c_412_n N_A_391_388#_M1010_g N_A_391_388#_c_404_n
+ N_A_391_388#_M1006_g N_A_391_388#_c_413_n N_A_391_388#_M1011_g
+ N_A_391_388#_c_405_n N_A_391_388#_M1014_g N_A_391_388#_c_414_n
+ N_A_391_388#_c_483_p N_A_391_388#_c_406_n N_A_391_388#_c_407_n
+ N_A_391_388#_c_408_n N_A_391_388#_c_457_p N_A_391_388#_c_409_n
+ N_A_391_388#_c_410_n N_A_391_388#_c_411_n PM_SKY130_FD_SC_HS__HA_2%A_391_388#
x_PM_SKY130_FD_SC_HS__HA_2%VPWR N_VPWR_M1002_s N_VPWR_M1003_d N_VPWR_M1000_d
+ N_VPWR_M1011_s N_VPWR_M1017_s N_VPWR_c_492_n N_VPWR_c_493_n N_VPWR_c_494_n
+ N_VPWR_c_495_n N_VPWR_c_496_n N_VPWR_c_497_n VPWR N_VPWR_c_498_n
+ N_VPWR_c_499_n N_VPWR_c_500_n N_VPWR_c_501_n N_VPWR_c_502_n N_VPWR_c_503_n
+ N_VPWR_c_504_n N_VPWR_c_491_n PM_SKY130_FD_SC_HS__HA_2%VPWR
x_PM_SKY130_FD_SC_HS__HA_2%SUM N_SUM_M1006_d N_SUM_M1010_d N_SUM_c_563_n
+ N_SUM_c_559_n SUM SUM N_SUM_c_561_n PM_SKY130_FD_SC_HS__HA_2%SUM
x_PM_SKY130_FD_SC_HS__HA_2%COUT N_COUT_M1001_d N_COUT_M1013_d N_COUT_c_594_n
+ N_COUT_c_591_n COUT COUT COUT PM_SKY130_FD_SC_HS__HA_2%COUT
x_PM_SKY130_FD_SC_HS__HA_2%VGND N_VGND_M1009_d N_VGND_M1007_d N_VGND_M1006_s
+ N_VGND_M1014_s N_VGND_M1008_s N_VGND_c_624_n N_VGND_c_625_n N_VGND_c_626_n
+ N_VGND_c_627_n N_VGND_c_628_n N_VGND_c_629_n N_VGND_c_630_n N_VGND_c_631_n
+ N_VGND_c_632_n N_VGND_c_633_n VGND N_VGND_c_634_n N_VGND_c_635_n
+ N_VGND_c_636_n N_VGND_c_637_n N_VGND_c_638_n N_VGND_c_639_n
+ PM_SKY130_FD_SC_HS__HA_2%VGND
x_PM_SKY130_FD_SC_HS__HA_2%A_278_74# N_A_278_74#_M1004_d N_A_278_74#_M1016_d
+ N_A_278_74#_c_697_n N_A_278_74#_c_698_n N_A_278_74#_c_699_n
+ N_A_278_74#_c_700_n N_A_278_74#_c_701_n PM_SKY130_FD_SC_HS__HA_2%A_278_74#
cc_1 VNB N_B_M1015_g 0.0297382f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_2 VNB N_B_c_103_n 0.0173977f $X=-0.19 $Y=-0.245 $X2=1.745 $Y2=1.185
cc_3 VNB N_B_c_104_n 0.0492605f $X=-0.19 $Y=-0.245 $X2=1.88 $Y2=1.865
cc_4 VNB N_B_c_105_n 0.00167339f $X=-0.19 $Y=-0.245 $X2=0.497 $Y2=1.79
cc_5 VNB N_B_c_106_n 0.0016809f $X=-0.19 $Y=-0.245 $X2=1.955 $Y2=1.615
cc_6 VNB N_B_c_107_n 0.0137652f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.465
cc_7 VNB N_B_c_108_n 0.0387746f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.465
cc_8 VNB B 0.00154267f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=2.32
cc_9 VNB N_A_M1009_g 0.0232343f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.3
cc_10 VNB N_A_M1004_g 0.0249069f $X=-0.19 $Y=-0.245 $X2=1.745 $Y2=1.185
cc_11 VNB N_A_c_190_n 0.0340356f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_27_74#_M1016_g 0.0257234f $X=-0.19 $Y=-0.245 $X2=1.745 $Y2=0.74
cc_13 VNB N_A_27_74#_M1001_g 0.0207917f $X=-0.19 $Y=-0.245 $X2=0.21 $Y2=1.465
cc_14 VNB N_A_27_74#_M1008_g 0.026707f $X=-0.19 $Y=-0.245 $X2=1.79 $Y2=2.42
cc_15 VNB N_A_27_74#_c_246_n 0.00327664f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=2.32
cc_16 VNB N_A_27_74#_c_247_n 0.02581f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_27_74#_c_248_n 0.0049904f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_27_74#_c_249_n 0.00942532f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_27_74#_c_250_n 0.0023864f $X=-0.19 $Y=-0.245 $X2=0.395 $Y2=1.465
cc_20 VNB N_A_27_74#_c_251_n 0.0286895f $X=-0.19 $Y=-0.245 $X2=0.395 $Y2=1.3
cc_21 VNB N_A_27_74#_c_252_n 9.06092e-19 $X=-0.19 $Y=-0.245 $X2=0.295 $Y2=2.42
cc_22 VNB N_A_27_74#_c_253_n 0.0748099f $X=-0.19 $Y=-0.245 $X2=1.2 $Y2=2.42
cc_23 VNB N_A_27_74#_c_254_n 0.00120577f $X=-0.19 $Y=-0.245 $X2=0.21 $Y2=2.32
cc_24 VNB N_A_27_74#_c_255_n 0.00146718f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_27_74#_c_256_n 0.00717931f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_27_74#_c_257_n 0.00509894f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_27_74#_c_258_n 0.0809936f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_391_388#_c_404_n 0.0198259f $X=-0.19 $Y=-0.245 $X2=1.745 $Y2=1.185
cc_29 VNB N_A_391_388#_c_405_n 0.017136f $X=-0.19 $Y=-0.245 $X2=0.497 $Y2=1.79
cc_30 VNB N_A_391_388#_c_406_n 0.003372f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.465
cc_31 VNB N_A_391_388#_c_407_n 0.00102048f $X=-0.19 $Y=-0.245 $X2=0.385
+ $Y2=1.465
cc_32 VNB N_A_391_388#_c_408_n 0.00213328f $X=-0.19 $Y=-0.245 $X2=1.79 $Y2=2.42
cc_33 VNB N_A_391_388#_c_409_n 0.0119963f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_391_388#_c_410_n 0.0608476f $X=-0.19 $Y=-0.245 $X2=0.395 $Y2=1.465
cc_35 VNB N_A_391_388#_c_411_n 0.0504091f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=2.42
cc_36 VNB N_VPWR_c_491_n 0.243291f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_SUM_c_559_n 0.00991076f $X=-0.19 $Y=-0.245 $X2=1.745 $Y2=0.74
cc_38 VNB N_COUT_c_591_n 0.00134727f $X=-0.19 $Y=-0.245 $X2=1.745 $Y2=0.74
cc_39 VNB COUT 0.00240191f $X=-0.19 $Y=-0.245 $X2=1.88 $Y2=1.865
cc_40 VNB COUT 0.00417716f $X=-0.19 $Y=-0.245 $X2=1.88 $Y2=2.44
cc_41 VNB N_VGND_c_624_n 0.00323505f $X=-0.19 $Y=-0.245 $X2=1.955 $Y2=2.32
cc_42 VNB N_VGND_c_625_n 0.00851745f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_626_n 0.00938716f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.465
cc_44 VNB N_VGND_c_627_n 0.00493915f $X=-0.19 $Y=-0.245 $X2=1.79 $Y2=2.42
cc_45 VNB N_VGND_c_628_n 0.010678f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=2.32
cc_46 VNB N_VGND_c_629_n 0.0450391f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=2.32
cc_47 VNB N_VGND_c_630_n 0.0291765f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_VGND_c_631_n 0.00601668f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_VGND_c_632_n 0.016486f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_VGND_c_633_n 0.00613227f $X=-0.19 $Y=-0.245 $X2=0.395 $Y2=1.465
cc_51 VNB N_VGND_c_634_n 0.0353722f $X=-0.19 $Y=-0.245 $X2=1.68 $Y2=2.42
cc_52 VNB N_VGND_c_635_n 0.0180771f $X=-0.19 $Y=-0.245 $X2=0.21 $Y2=2.42
cc_53 VNB N_VGND_c_636_n 0.0193312f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_VGND_c_637_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_VGND_c_638_n 0.00461913f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_VGND_c_639_n 0.34251f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_A_278_74#_c_697_n 0.0101103f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.845
cc_58 VNB N_A_278_74#_c_698_n 0.00817638f $X=-0.19 $Y=-0.245 $X2=1.745 $Y2=0.74
cc_59 VNB N_A_278_74#_c_699_n 0.013117f $X=-0.19 $Y=-0.245 $X2=1.88 $Y2=1.865
cc_60 VNB N_A_278_74#_c_700_n 0.00353599f $X=-0.19 $Y=-0.245 $X2=1.88 $Y2=2.44
cc_61 VNB N_A_278_74#_c_701_n 0.00359387f $X=-0.19 $Y=-0.245 $X2=0.497 $Y2=1.845
cc_62 VPB N_B_c_104_n 0.0386617f $X=-0.19 $Y=1.66 $X2=1.88 $Y2=1.865
cc_63 VPB N_B_c_105_n 0.00744368f $X=-0.19 $Y=1.66 $X2=0.497 $Y2=1.79
cc_64 VPB N_B_c_112_n 0.0206483f $X=-0.19 $Y=1.66 $X2=0.497 $Y2=1.845
cc_65 VPB N_B_c_106_n 0.00230962f $X=-0.19 $Y=1.66 $X2=1.955 $Y2=1.615
cc_66 VPB B 0.0338761f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=2.32
cc_67 VPB N_A_c_191_n 0.0144258f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.74
cc_68 VPB N_A_c_192_n 0.0148446f $X=-0.19 $Y=1.66 $X2=1.745 $Y2=0.74
cc_69 VPB A 0.00483519f $X=-0.19 $Y=1.66 $X2=1.88 $Y2=2.44
cc_70 VPB N_A_c_190_n 0.0318734f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_71 VPB N_A_27_74#_c_259_n 0.0150909f $X=-0.19 $Y=1.66 $X2=1.955 $Y2=2.32
cc_72 VPB N_A_27_74#_c_260_n 0.0170327f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_73 VPB N_A_27_74#_c_246_n 0.00862625f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=2.32
cc_74 VPB N_A_27_74#_c_262_n 0.0269171f $X=-0.19 $Y=1.66 $X2=1.115 $Y2=2.32
cc_75 VPB N_A_27_74#_c_250_n 0.00213301f $X=-0.19 $Y=1.66 $X2=0.395 $Y2=1.465
cc_76 VPB N_A_27_74#_c_252_n 0.00605612f $X=-0.19 $Y=1.66 $X2=0.295 $Y2=2.42
cc_77 VPB N_A_27_74#_c_254_n 0.00773266f $X=-0.19 $Y=1.66 $X2=0.21 $Y2=2.32
cc_78 VPB N_A_27_74#_c_258_n 0.0130607f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_79 VPB N_A_391_388#_c_412_n 0.0174024f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.845
cc_80 VPB N_A_391_388#_c_413_n 0.014966f $X=-0.19 $Y=1.66 $X2=1.88 $Y2=1.865
cc_81 VPB N_A_391_388#_c_414_n 0.0111715f $X=-0.19 $Y=1.66 $X2=1.955 $Y2=1.615
cc_82 VPB N_A_391_388#_c_408_n 0.00648012f $X=-0.19 $Y=1.66 $X2=1.79 $Y2=2.42
cc_83 VPB N_A_391_388#_c_411_n 0.0138232f $X=-0.19 $Y=1.66 $X2=0.72 $Y2=2.42
cc_84 VPB N_VPWR_c_492_n 0.0121909f $X=-0.19 $Y=1.66 $X2=0.497 $Y2=1.79
cc_85 VPB N_VPWR_c_493_n 0.0209179f $X=-0.19 $Y=1.66 $X2=1.955 $Y2=2.32
cc_86 VPB N_VPWR_c_494_n 0.00454805f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_87 VPB N_VPWR_c_495_n 0.00261656f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.465
cc_88 VPB N_VPWR_c_496_n 0.0120106f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.465
cc_89 VPB N_VPWR_c_497_n 0.0208276f $X=-0.19 $Y=1.66 $X2=1.79 $Y2=2.42
cc_90 VPB N_VPWR_c_498_n 0.0180749f $X=-0.19 $Y=1.66 $X2=1.595 $Y2=2.32
cc_91 VPB N_VPWR_c_499_n 0.017758f $X=-0.19 $Y=1.66 $X2=1.895 $Y2=1.615
cc_92 VPB N_VPWR_c_500_n 0.0177589f $X=-0.19 $Y=1.66 $X2=1.2 $Y2=2.42
cc_93 VPB N_VPWR_c_501_n 0.00734343f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_94 VPB N_VPWR_c_502_n 0.0533445f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_95 VPB N_VPWR_c_503_n 0.0224214f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_96 VPB N_VPWR_c_504_n 0.00601644f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_97 VPB N_VPWR_c_491_n 0.0888061f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_98 VPB N_SUM_c_559_n 0.00296383f $X=-0.19 $Y=1.66 $X2=1.745 $Y2=0.74
cc_99 VPB N_SUM_c_561_n 0.00438767f $X=-0.19 $Y=1.66 $X2=1.955 $Y2=2.32
cc_100 VPB N_COUT_c_594_n 0.00136846f $X=-0.19 $Y=1.66 $X2=1.745 $Y2=1.185
cc_101 VPB N_COUT_c_591_n 0.00114783f $X=-0.19 $Y=1.66 $X2=1.745 $Y2=0.74
cc_102 N_B_M1015_g N_A_M1009_g 0.0340417f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_103 N_B_c_107_n N_A_M1009_g 2.56105e-19 $X=0.385 $Y=1.465 $X2=0 $Y2=0
cc_104 N_B_c_112_n N_A_c_191_n 0.0352089f $X=0.497 $Y=1.845 $X2=0 $Y2=0
cc_105 N_B_c_118_p N_A_c_191_n 0.0176674f $X=1.79 $Y=2.42 $X2=0 $Y2=0
cc_106 N_B_c_103_n N_A_M1004_g 0.0312814f $X=1.745 $Y=1.185 $X2=0 $Y2=0
cc_107 N_B_c_104_n N_A_M1004_g 0.00903936f $X=1.88 $Y=1.865 $X2=0 $Y2=0
cc_108 N_B_c_104_n N_A_c_192_n 0.0560482f $X=1.88 $Y=1.865 $X2=0 $Y2=0
cc_109 N_B_c_106_n N_A_c_192_n 0.00261121f $X=1.955 $Y=1.615 $X2=0 $Y2=0
cc_110 N_B_c_118_p N_A_c_192_n 0.0177597f $X=1.79 $Y=2.42 $X2=0 $Y2=0
cc_111 N_B_c_104_n A 0.00116553f $X=1.88 $Y=1.865 $X2=0 $Y2=0
cc_112 N_B_c_106_n A 0.0124269f $X=1.955 $Y=1.615 $X2=0 $Y2=0
cc_113 N_B_c_118_p A 0.00992318f $X=1.79 $Y=2.42 $X2=0 $Y2=0
cc_114 N_B_c_104_n N_A_c_190_n 0.014075f $X=1.88 $Y=1.865 $X2=0 $Y2=0
cc_115 N_B_c_112_n N_A_c_190_n 0.00218507f $X=0.497 $Y=1.845 $X2=0 $Y2=0
cc_116 N_B_c_106_n N_A_c_190_n 0.00207072f $X=1.955 $Y=1.615 $X2=0 $Y2=0
cc_117 N_B_c_108_n N_A_c_190_n 0.043321f $X=0.385 $Y=1.465 $X2=0 $Y2=0
cc_118 N_B_c_118_p N_A_c_190_n 0.00139277f $X=1.79 $Y=2.42 $X2=0 $Y2=0
cc_119 N_B_c_118_p N_A_27_74#_M1002_d 0.00570774f $X=1.79 $Y=2.42 $X2=0 $Y2=0
cc_120 N_B_M1015_g N_A_27_74#_c_247_n 0.0123382f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_121 N_B_M1015_g N_A_27_74#_c_248_n 0.0108371f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_122 N_B_c_112_n N_A_27_74#_c_248_n 2.50378e-19 $X=0.497 $Y=1.845 $X2=0 $Y2=0
cc_123 N_B_c_107_n N_A_27_74#_c_248_n 0.00746443f $X=0.385 $Y=1.465 $X2=0 $Y2=0
cc_124 N_B_M1015_g N_A_27_74#_c_249_n 0.00113234f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_125 N_B_c_107_n N_A_27_74#_c_249_n 0.0272661f $X=0.385 $Y=1.465 $X2=0 $Y2=0
cc_126 N_B_c_108_n N_A_27_74#_c_249_n 0.00467141f $X=0.385 $Y=1.465 $X2=0 $Y2=0
cc_127 N_B_c_112_n N_A_27_74#_c_250_n 0.00147639f $X=0.497 $Y=1.845 $X2=0 $Y2=0
cc_128 N_B_c_107_n N_A_27_74#_c_250_n 0.025258f $X=0.385 $Y=1.465 $X2=0 $Y2=0
cc_129 N_B_c_108_n N_A_27_74#_c_250_n 0.00348918f $X=0.385 $Y=1.465 $X2=0 $Y2=0
cc_130 B N_A_27_74#_c_250_n 0.0137455f $X=0.155 $Y=2.32 $X2=0 $Y2=0
cc_131 N_B_c_103_n N_A_27_74#_c_251_n 0.00565175f $X=1.745 $Y=1.185 $X2=0 $Y2=0
cc_132 N_B_c_104_n N_A_27_74#_c_251_n 0.0152616f $X=1.88 $Y=1.865 $X2=0 $Y2=0
cc_133 N_B_c_106_n N_A_27_74#_c_251_n 0.0256551f $X=1.955 $Y=1.615 $X2=0 $Y2=0
cc_134 N_B_c_104_n N_A_27_74#_c_252_n 0.00651386f $X=1.88 $Y=1.865 $X2=0 $Y2=0
cc_135 N_B_c_106_n N_A_27_74#_c_252_n 0.0544241f $X=1.955 $Y=1.615 $X2=0 $Y2=0
cc_136 N_B_c_118_p N_A_27_74#_c_252_n 0.00159069f $X=1.79 $Y=2.42 $X2=0 $Y2=0
cc_137 N_B_c_104_n N_A_27_74#_c_253_n 0.0123225f $X=1.88 $Y=1.865 $X2=0 $Y2=0
cc_138 N_B_c_104_n N_A_27_74#_c_286_n 9.20426e-19 $X=1.88 $Y=1.865 $X2=0 $Y2=0
cc_139 N_B_c_118_p N_A_27_74#_c_286_n 0.0153274f $X=1.79 $Y=2.42 $X2=0 $Y2=0
cc_140 N_B_c_112_n N_A_27_74#_c_288_n 0.00288122f $X=0.497 $Y=1.845 $X2=0 $Y2=0
cc_141 N_B_c_118_p N_A_27_74#_c_288_n 0.0156678f $X=1.79 $Y=2.42 $X2=0 $Y2=0
cc_142 B N_A_27_74#_c_288_n 0.00872351f $X=0.155 $Y=2.32 $X2=0 $Y2=0
cc_143 N_B_M1015_g N_A_27_74#_c_255_n 0.0036485f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_144 N_B_c_104_n N_A_27_74#_c_256_n 0.00506711f $X=1.88 $Y=1.865 $X2=0 $Y2=0
cc_145 N_B_c_106_n N_A_27_74#_c_256_n 0.0134933f $X=1.955 $Y=1.615 $X2=0 $Y2=0
cc_146 N_B_c_106_n N_A_391_388#_M1005_d 0.00412198f $X=1.955 $Y=1.615 $X2=0
+ $Y2=0
cc_147 N_B_c_118_p N_A_391_388#_M1005_d 0.00502998f $X=1.79 $Y=2.42 $X2=0 $Y2=0
cc_148 N_B_c_118_p N_VPWR_M1002_s 0.00222182f $X=1.79 $Y=2.42 $X2=-0.19
+ $Y2=-0.245
cc_149 B N_VPWR_M1002_s 0.01041f $X=0.155 $Y=2.32 $X2=-0.19 $Y2=-0.245
cc_150 N_B_c_118_p N_VPWR_M1003_d 0.0064423f $X=1.79 $Y=2.42 $X2=0 $Y2=0
cc_151 N_B_c_112_n N_VPWR_c_493_n 0.0094261f $X=0.497 $Y=1.845 $X2=0 $Y2=0
cc_152 N_B_c_118_p N_VPWR_c_493_n 0.0072308f $X=1.79 $Y=2.42 $X2=0 $Y2=0
cc_153 B N_VPWR_c_493_n 0.0148608f $X=0.155 $Y=2.32 $X2=0 $Y2=0
cc_154 N_B_c_104_n N_VPWR_c_494_n 0.00182212f $X=1.88 $Y=1.865 $X2=0 $Y2=0
cc_155 N_B_c_112_n N_VPWR_c_494_n 0.00106224f $X=0.497 $Y=1.845 $X2=0 $Y2=0
cc_156 N_B_c_118_p N_VPWR_c_494_n 0.0213502f $X=1.79 $Y=2.42 $X2=0 $Y2=0
cc_157 N_B_c_112_n N_VPWR_c_498_n 0.00492531f $X=0.497 $Y=1.845 $X2=0 $Y2=0
cc_158 N_B_c_104_n N_VPWR_c_502_n 0.00563421f $X=1.88 $Y=1.865 $X2=0 $Y2=0
cc_159 N_B_c_104_n N_VPWR_c_491_n 0.00539454f $X=1.88 $Y=1.865 $X2=0 $Y2=0
cc_160 N_B_c_112_n N_VPWR_c_491_n 0.00483326f $X=0.497 $Y=1.845 $X2=0 $Y2=0
cc_161 N_B_c_118_p N_VPWR_c_491_n 0.0477545f $X=1.79 $Y=2.42 $X2=0 $Y2=0
cc_162 B N_VPWR_c_491_n 6.43314e-19 $X=0.155 $Y=2.32 $X2=0 $Y2=0
cc_163 N_B_c_118_p A_307_388# 0.00918698f $X=1.79 $Y=2.42 $X2=-0.19 $Y2=-0.245
cc_164 N_B_M1015_g N_VGND_c_624_n 0.00126873f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_165 N_B_c_103_n N_VGND_c_624_n 0.00106137f $X=1.745 $Y=1.185 $X2=0 $Y2=0
cc_166 N_B_c_103_n N_VGND_c_625_n 0.00970106f $X=1.745 $Y=1.185 $X2=0 $Y2=0
cc_167 N_B_M1015_g N_VGND_c_630_n 0.00434272f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_168 N_B_c_103_n N_VGND_c_632_n 0.00383152f $X=1.745 $Y=1.185 $X2=0 $Y2=0
cc_169 N_B_M1015_g N_VGND_c_639_n 0.00824638f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_170 N_B_c_103_n N_VGND_c_639_n 0.00369368f $X=1.745 $Y=1.185 $X2=0 $Y2=0
cc_171 N_B_c_103_n N_A_278_74#_c_697_n 0.0113476f $X=1.745 $Y=1.185 $X2=0 $Y2=0
cc_172 N_B_c_104_n N_A_278_74#_c_697_n 5.76956e-19 $X=1.88 $Y=1.865 $X2=0 $Y2=0
cc_173 N_B_c_103_n N_A_278_74#_c_698_n 0.0028624f $X=1.745 $Y=1.185 $X2=0 $Y2=0
cc_174 N_B_c_103_n N_A_278_74#_c_700_n 5.73857e-19 $X=1.745 $Y=1.185 $X2=0 $Y2=0
cc_175 N_A_M1009_g N_A_27_74#_c_247_n 0.00248918f $X=0.885 $Y=0.74 $X2=0 $Y2=0
cc_176 N_A_M1009_g N_A_27_74#_c_248_n 2.23249e-19 $X=0.885 $Y=0.74 $X2=0 $Y2=0
cc_177 N_A_M1009_g N_A_27_74#_c_250_n 0.00308843f $X=0.885 $Y=0.74 $X2=0 $Y2=0
cc_178 N_A_c_191_n N_A_27_74#_c_250_n 0.00289279f $X=0.955 $Y=1.845 $X2=0 $Y2=0
cc_179 N_A_c_192_n N_A_27_74#_c_250_n 5.30451e-19 $X=1.46 $Y=1.865 $X2=0 $Y2=0
cc_180 A N_A_27_74#_c_250_n 0.0236478f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_181 N_A_c_190_n N_A_27_74#_c_250_n 0.0141497f $X=1.315 $Y=1.632 $X2=0 $Y2=0
cc_182 N_A_M1009_g N_A_27_74#_c_251_n 0.00934412f $X=0.885 $Y=0.74 $X2=0 $Y2=0
cc_183 N_A_M1004_g N_A_27_74#_c_251_n 0.0137279f $X=1.315 $Y=0.74 $X2=0 $Y2=0
cc_184 A N_A_27_74#_c_251_n 0.0242166f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_185 N_A_c_190_n N_A_27_74#_c_251_n 0.00813003f $X=1.315 $Y=1.632 $X2=0 $Y2=0
cc_186 N_A_c_191_n N_A_27_74#_c_288_n 0.00362798f $X=0.955 $Y=1.845 $X2=0 $Y2=0
cc_187 N_A_c_192_n N_A_27_74#_c_288_n 7.7971e-19 $X=1.46 $Y=1.865 $X2=0 $Y2=0
cc_188 N_A_M1009_g N_A_27_74#_c_255_n 0.0106214f $X=0.885 $Y=0.74 $X2=0 $Y2=0
cc_189 N_A_M1004_g N_A_27_74#_c_255_n 0.00156882f $X=1.315 $Y=0.74 $X2=0 $Y2=0
cc_190 N_A_c_191_n N_VPWR_c_493_n 0.00106331f $X=0.955 $Y=1.845 $X2=0 $Y2=0
cc_191 N_A_c_191_n N_VPWR_c_494_n 0.0086645f $X=0.955 $Y=1.845 $X2=0 $Y2=0
cc_192 N_A_c_192_n N_VPWR_c_494_n 0.00920258f $X=1.46 $Y=1.865 $X2=0 $Y2=0
cc_193 N_A_c_191_n N_VPWR_c_498_n 0.00492531f $X=0.955 $Y=1.845 $X2=0 $Y2=0
cc_194 N_A_c_192_n N_VPWR_c_502_n 0.00505726f $X=1.46 $Y=1.865 $X2=0 $Y2=0
cc_195 N_A_c_191_n N_VPWR_c_491_n 0.00483326f $X=0.955 $Y=1.845 $X2=0 $Y2=0
cc_196 N_A_c_192_n N_VPWR_c_491_n 0.00489105f $X=1.46 $Y=1.865 $X2=0 $Y2=0
cc_197 N_A_M1009_g N_VGND_c_624_n 0.00876864f $X=0.885 $Y=0.74 $X2=0 $Y2=0
cc_198 N_A_M1004_g N_VGND_c_624_n 0.00891708f $X=1.315 $Y=0.74 $X2=0 $Y2=0
cc_199 N_A_M1004_g N_VGND_c_625_n 0.00106137f $X=1.315 $Y=0.74 $X2=0 $Y2=0
cc_200 N_A_M1009_g N_VGND_c_630_n 0.00383152f $X=0.885 $Y=0.74 $X2=0 $Y2=0
cc_201 N_A_M1004_g N_VGND_c_632_n 0.00383152f $X=1.315 $Y=0.74 $X2=0 $Y2=0
cc_202 N_A_M1009_g N_VGND_c_639_n 0.0075725f $X=0.885 $Y=0.74 $X2=0 $Y2=0
cc_203 N_A_M1004_g N_VGND_c_639_n 0.006806f $X=1.315 $Y=0.74 $X2=0 $Y2=0
cc_204 N_A_M1009_g N_A_278_74#_c_697_n 8.11834e-19 $X=0.885 $Y=0.74 $X2=0 $Y2=0
cc_205 N_A_M1004_g N_A_278_74#_c_697_n 0.00416578f $X=1.315 $Y=0.74 $X2=0 $Y2=0
cc_206 N_A_27_74#_c_252_n N_A_391_388#_M1005_d 0.0119981f $X=2.375 $Y=2.34 $X2=0
+ $Y2=0
cc_207 N_A_27_74#_c_310_p N_A_391_388#_M1005_d 0.0204624f $X=5.385 $Y=2.425
+ $X2=0 $Y2=0
cc_208 N_A_27_74#_c_286_n N_A_391_388#_M1005_d 0.00709606f $X=2.46 $Y=2.425
+ $X2=0 $Y2=0
cc_209 N_A_27_74#_c_310_p N_A_391_388#_c_412_n 0.0179844f $X=5.385 $Y=2.425
+ $X2=0 $Y2=0
cc_210 N_A_27_74#_c_259_n N_A_391_388#_c_413_n 0.0390158f $X=4.805 $Y=1.765
+ $X2=0 $Y2=0
cc_211 N_A_27_74#_c_310_p N_A_391_388#_c_413_n 0.0118981f $X=5.385 $Y=2.425
+ $X2=0 $Y2=0
cc_212 N_A_27_74#_M1001_g N_A_391_388#_c_405_n 0.0282033f $X=4.835 $Y=0.74 $X2=0
+ $Y2=0
cc_213 N_A_27_74#_c_262_n N_A_391_388#_c_414_n 0.016066f $X=3.012 $Y=1.865 $X2=0
+ $Y2=0
cc_214 N_A_27_74#_c_252_n N_A_391_388#_c_414_n 0.0202358f $X=2.375 $Y=2.34 $X2=0
+ $Y2=0
cc_215 N_A_27_74#_c_318_p N_A_391_388#_c_414_n 0.0196613f $X=2.87 $Y=1.445 $X2=0
+ $Y2=0
cc_216 N_A_27_74#_c_253_n N_A_391_388#_c_414_n 0.0063963f $X=2.87 $Y=1.445 $X2=0
+ $Y2=0
cc_217 N_A_27_74#_c_310_p N_A_391_388#_c_414_n 0.0560957f $X=5.385 $Y=2.425
+ $X2=0 $Y2=0
cc_218 N_A_27_74#_M1016_g N_A_391_388#_c_406_n 0.012478f $X=2.935 $Y=0.74 $X2=0
+ $Y2=0
cc_219 N_A_27_74#_c_262_n N_A_391_388#_c_406_n 3.68309e-19 $X=3.012 $Y=1.865
+ $X2=0 $Y2=0
cc_220 N_A_27_74#_c_318_p N_A_391_388#_c_406_n 0.0136762f $X=2.87 $Y=1.445 $X2=0
+ $Y2=0
cc_221 N_A_27_74#_c_253_n N_A_391_388#_c_406_n 0.00191708f $X=2.87 $Y=1.445
+ $X2=0 $Y2=0
cc_222 N_A_27_74#_c_318_p N_A_391_388#_c_407_n 0.0136463f $X=2.87 $Y=1.445 $X2=0
+ $Y2=0
cc_223 N_A_27_74#_c_253_n N_A_391_388#_c_407_n 0.00391672f $X=2.87 $Y=1.445
+ $X2=0 $Y2=0
cc_224 N_A_27_74#_c_262_n N_A_391_388#_c_408_n 0.00418912f $X=3.012 $Y=1.865
+ $X2=0 $Y2=0
cc_225 N_A_27_74#_c_253_n N_A_391_388#_c_408_n 0.00722092f $X=2.87 $Y=1.445
+ $X2=0 $Y2=0
cc_226 N_A_27_74#_M1016_g N_A_391_388#_c_409_n 0.00421066f $X=2.935 $Y=0.74
+ $X2=0 $Y2=0
cc_227 N_A_27_74#_c_318_p N_A_391_388#_c_409_n 0.0167012f $X=2.87 $Y=1.445 $X2=0
+ $Y2=0
cc_228 N_A_27_74#_c_253_n N_A_391_388#_c_409_n 0.00118728f $X=2.87 $Y=1.445
+ $X2=0 $Y2=0
cc_229 N_A_27_74#_M1016_g N_A_391_388#_c_410_n 0.00275209f $X=2.935 $Y=0.74
+ $X2=0 $Y2=0
cc_230 N_A_27_74#_c_318_p N_A_391_388#_c_410_n 0.00106912f $X=2.87 $Y=1.445
+ $X2=0 $Y2=0
cc_231 N_A_27_74#_c_253_n N_A_391_388#_c_410_n 0.0158741f $X=2.87 $Y=1.445 $X2=0
+ $Y2=0
cc_232 N_A_27_74#_c_258_n N_A_391_388#_c_411_n 0.0187183f $X=5.265 $Y=1.532
+ $X2=0 $Y2=0
cc_233 N_A_27_74#_c_310_p N_VPWR_M1000_d 0.0243996f $X=5.385 $Y=2.425 $X2=0
+ $Y2=0
cc_234 N_A_27_74#_c_310_p N_VPWR_M1011_s 0.00392503f $X=5.385 $Y=2.425 $X2=0
+ $Y2=0
cc_235 N_A_27_74#_c_310_p N_VPWR_M1017_s 0.00991231f $X=5.385 $Y=2.425 $X2=0
+ $Y2=0
cc_236 N_A_27_74#_c_254_n N_VPWR_M1017_s 0.0224403f $X=5.47 $Y=2.34 $X2=0 $Y2=0
cc_237 N_A_27_74#_c_259_n N_VPWR_c_495_n 0.00924105f $X=4.805 $Y=1.765 $X2=0
+ $Y2=0
cc_238 N_A_27_74#_c_260_n N_VPWR_c_495_n 0.00121234f $X=5.255 $Y=1.765 $X2=0
+ $Y2=0
cc_239 N_A_27_74#_c_310_p N_VPWR_c_495_n 0.0167733f $X=5.385 $Y=2.425 $X2=0
+ $Y2=0
cc_240 N_A_27_74#_c_259_n N_VPWR_c_497_n 0.00121234f $X=4.805 $Y=1.765 $X2=0
+ $Y2=0
cc_241 N_A_27_74#_c_260_n N_VPWR_c_497_n 0.0102712f $X=5.255 $Y=1.765 $X2=0
+ $Y2=0
cc_242 N_A_27_74#_c_310_p N_VPWR_c_497_n 0.0157096f $X=5.385 $Y=2.425 $X2=0
+ $Y2=0
cc_243 N_A_27_74#_c_259_n N_VPWR_c_500_n 0.00413917f $X=4.805 $Y=1.765 $X2=0
+ $Y2=0
cc_244 N_A_27_74#_c_260_n N_VPWR_c_500_n 0.00413917f $X=5.255 $Y=1.765 $X2=0
+ $Y2=0
cc_245 N_A_27_74#_c_262_n N_VPWR_c_502_n 0.00505726f $X=3.012 $Y=1.865 $X2=0
+ $Y2=0
cc_246 N_A_27_74#_c_262_n N_VPWR_c_503_n 0.0216343f $X=3.012 $Y=1.865 $X2=0
+ $Y2=0
cc_247 N_A_27_74#_c_310_p N_VPWR_c_503_n 0.0512284f $X=5.385 $Y=2.425 $X2=0
+ $Y2=0
cc_248 N_A_27_74#_c_259_n N_VPWR_c_491_n 0.00409982f $X=4.805 $Y=1.765 $X2=0
+ $Y2=0
cc_249 N_A_27_74#_c_260_n N_VPWR_c_491_n 0.00409982f $X=5.255 $Y=1.765 $X2=0
+ $Y2=0
cc_250 N_A_27_74#_c_262_n N_VPWR_c_491_n 0.00485508f $X=3.012 $Y=1.865 $X2=0
+ $Y2=0
cc_251 N_A_27_74#_c_310_p N_VPWR_c_491_n 0.0620685f $X=5.385 $Y=2.425 $X2=0
+ $Y2=0
cc_252 N_A_27_74#_c_286_n N_VPWR_c_491_n 0.00678047f $X=2.46 $Y=2.425 $X2=0
+ $Y2=0
cc_253 N_A_27_74#_c_310_p N_SUM_M1010_d 0.00565759f $X=5.385 $Y=2.425 $X2=0
+ $Y2=0
cc_254 N_A_27_74#_M1001_g N_SUM_c_563_n 0.00141692f $X=4.835 $Y=0.74 $X2=0 $Y2=0
cc_255 N_A_27_74#_c_259_n N_SUM_c_559_n 0.00207233f $X=4.805 $Y=1.765 $X2=0
+ $Y2=0
cc_256 N_A_27_74#_M1001_g N_SUM_c_559_n 0.00177272f $X=4.835 $Y=0.74 $X2=0 $Y2=0
cc_257 N_A_27_74#_c_310_p N_SUM_c_559_n 0.0136682f $X=5.385 $Y=2.425 $X2=0 $Y2=0
cc_258 N_A_27_74#_c_258_n N_SUM_c_559_n 0.00413919f $X=5.265 $Y=1.532 $X2=0
+ $Y2=0
cc_259 N_A_27_74#_c_310_p N_SUM_c_561_n 0.0273851f $X=5.385 $Y=2.425 $X2=0 $Y2=0
cc_260 N_A_27_74#_c_310_p N_COUT_M1013_d 0.00565277f $X=5.385 $Y=2.425 $X2=0
+ $Y2=0
cc_261 N_A_27_74#_c_259_n N_COUT_c_594_n 0.00454405f $X=4.805 $Y=1.765 $X2=0
+ $Y2=0
cc_262 N_A_27_74#_c_260_n N_COUT_c_594_n 0.00476771f $X=5.255 $Y=1.765 $X2=0
+ $Y2=0
cc_263 N_A_27_74#_c_310_p N_COUT_c_594_n 0.0167898f $X=5.385 $Y=2.425 $X2=0
+ $Y2=0
cc_264 N_A_27_74#_c_254_n N_COUT_c_594_n 0.0126742f $X=5.47 $Y=2.34 $X2=0 $Y2=0
cc_265 N_A_27_74#_c_258_n N_COUT_c_594_n 0.00565377f $X=5.265 $Y=1.532 $X2=0
+ $Y2=0
cc_266 N_A_27_74#_c_259_n N_COUT_c_591_n 5.42499e-19 $X=4.805 $Y=1.765 $X2=0
+ $Y2=0
cc_267 N_A_27_74#_M1001_g N_COUT_c_591_n 0.00331881f $X=4.835 $Y=0.74 $X2=0
+ $Y2=0
cc_268 N_A_27_74#_M1008_g N_COUT_c_591_n 0.002587f $X=5.265 $Y=0.74 $X2=0 $Y2=0
cc_269 N_A_27_74#_c_254_n N_COUT_c_591_n 0.0066156f $X=5.47 $Y=2.34 $X2=0 $Y2=0
cc_270 N_A_27_74#_c_257_n N_COUT_c_591_n 0.0235661f $X=5.39 $Y=1.465 $X2=0 $Y2=0
cc_271 N_A_27_74#_c_258_n N_COUT_c_591_n 0.02154f $X=5.265 $Y=1.532 $X2=0 $Y2=0
cc_272 N_A_27_74#_M1001_g COUT 0.00892916f $X=4.835 $Y=0.74 $X2=0 $Y2=0
cc_273 N_A_27_74#_M1008_g COUT 0.00788704f $X=5.265 $Y=0.74 $X2=0 $Y2=0
cc_274 N_A_27_74#_M1001_g COUT 0.00203717f $X=4.835 $Y=0.74 $X2=0 $Y2=0
cc_275 N_A_27_74#_M1008_g COUT 0.00327512f $X=5.265 $Y=0.74 $X2=0 $Y2=0
cc_276 N_A_27_74#_c_258_n COUT 0.00199986f $X=5.265 $Y=1.532 $X2=0 $Y2=0
cc_277 N_A_27_74#_c_248_n A_114_74# 0.0039014f $X=0.72 $Y=1.045 $X2=-0.19
+ $Y2=-0.245
cc_278 N_A_27_74#_c_255_n A_114_74# 0.0018016f $X=0.805 $Y=1.045 $X2=-0.19
+ $Y2=-0.245
cc_279 N_A_27_74#_c_247_n N_VGND_c_624_n 0.00792017f $X=0.28 $Y=0.515 $X2=0
+ $Y2=0
cc_280 N_A_27_74#_c_251_n N_VGND_c_624_n 0.00968283f $X=2.29 $Y=1.195 $X2=0
+ $Y2=0
cc_281 N_A_27_74#_M1016_g N_VGND_c_626_n 0.00144451f $X=2.935 $Y=0.74 $X2=0
+ $Y2=0
cc_282 N_A_27_74#_M1001_g N_VGND_c_627_n 0.00294833f $X=4.835 $Y=0.74 $X2=0
+ $Y2=0
cc_283 N_A_27_74#_M1008_g N_VGND_c_629_n 0.00647412f $X=5.265 $Y=0.74 $X2=0
+ $Y2=0
cc_284 N_A_27_74#_c_257_n N_VGND_c_629_n 0.0140864f $X=5.39 $Y=1.465 $X2=0 $Y2=0
cc_285 N_A_27_74#_c_258_n N_VGND_c_629_n 0.00125053f $X=5.265 $Y=1.532 $X2=0
+ $Y2=0
cc_286 N_A_27_74#_c_247_n N_VGND_c_630_n 0.0145639f $X=0.28 $Y=0.515 $X2=0 $Y2=0
cc_287 N_A_27_74#_M1016_g N_VGND_c_634_n 0.00278247f $X=2.935 $Y=0.74 $X2=0
+ $Y2=0
cc_288 N_A_27_74#_M1001_g N_VGND_c_636_n 0.00434272f $X=4.835 $Y=0.74 $X2=0
+ $Y2=0
cc_289 N_A_27_74#_M1008_g N_VGND_c_636_n 0.00434272f $X=5.265 $Y=0.74 $X2=0
+ $Y2=0
cc_290 N_A_27_74#_M1016_g N_VGND_c_639_n 0.00363424f $X=2.935 $Y=0.74 $X2=0
+ $Y2=0
cc_291 N_A_27_74#_M1001_g N_VGND_c_639_n 0.00820382f $X=4.835 $Y=0.74 $X2=0
+ $Y2=0
cc_292 N_A_27_74#_M1008_g N_VGND_c_639_n 0.00823942f $X=5.265 $Y=0.74 $X2=0
+ $Y2=0
cc_293 N_A_27_74#_c_247_n N_VGND_c_639_n 0.0119984f $X=0.28 $Y=0.515 $X2=0 $Y2=0
cc_294 N_A_27_74#_c_251_n N_A_278_74#_c_697_n 0.0613147f $X=2.29 $Y=1.195 $X2=0
+ $Y2=0
cc_295 N_A_27_74#_c_318_p N_A_278_74#_c_697_n 2.30459e-19 $X=2.87 $Y=1.445 $X2=0
+ $Y2=0
cc_296 N_A_27_74#_c_253_n N_A_278_74#_c_697_n 6.05904e-19 $X=2.87 $Y=1.445 $X2=0
+ $Y2=0
cc_297 N_A_27_74#_c_256_n N_A_278_74#_c_697_n 0.0158527f $X=2.375 $Y=1.36 $X2=0
+ $Y2=0
cc_298 N_A_27_74#_M1016_g N_A_278_74#_c_698_n 0.00317277f $X=2.935 $Y=0.74 $X2=0
+ $Y2=0
cc_299 N_A_27_74#_M1016_g N_A_278_74#_c_699_n 0.0131176f $X=2.935 $Y=0.74 $X2=0
+ $Y2=0
cc_300 N_A_27_74#_M1016_g N_A_278_74#_c_701_n 0.00549447f $X=2.935 $Y=0.74 $X2=0
+ $Y2=0
cc_301 N_A_391_388#_c_414_n N_VPWR_M1000_d 0.0097331f $X=3.32 $Y=2.045 $X2=0
+ $Y2=0
cc_302 N_A_391_388#_c_412_n N_VPWR_c_495_n 0.00121367f $X=3.905 $Y=1.765 $X2=0
+ $Y2=0
cc_303 N_A_391_388#_c_413_n N_VPWR_c_495_n 0.00921829f $X=4.355 $Y=1.765 $X2=0
+ $Y2=0
cc_304 N_A_391_388#_c_412_n N_VPWR_c_499_n 0.00413917f $X=3.905 $Y=1.765 $X2=0
+ $Y2=0
cc_305 N_A_391_388#_c_413_n N_VPWR_c_499_n 0.00413917f $X=4.355 $Y=1.765 $X2=0
+ $Y2=0
cc_306 N_A_391_388#_c_412_n N_VPWR_c_503_n 0.0107942f $X=3.905 $Y=1.765 $X2=0
+ $Y2=0
cc_307 N_A_391_388#_c_413_n N_VPWR_c_503_n 0.00120587f $X=4.355 $Y=1.765 $X2=0
+ $Y2=0
cc_308 N_A_391_388#_c_412_n N_VPWR_c_491_n 0.00408365f $X=3.905 $Y=1.765 $X2=0
+ $Y2=0
cc_309 N_A_391_388#_c_413_n N_VPWR_c_491_n 0.00409982f $X=4.355 $Y=1.765 $X2=0
+ $Y2=0
cc_310 N_A_391_388#_c_404_n N_SUM_c_563_n 0.00614403f $X=3.925 $Y=1.22 $X2=0
+ $Y2=0
cc_311 N_A_391_388#_c_405_n N_SUM_c_563_n 0.015895f $X=4.405 $Y=1.22 $X2=0 $Y2=0
cc_312 N_A_391_388#_c_457_p N_SUM_c_563_n 0.021978f $X=4.165 $Y=1.385 $X2=0
+ $Y2=0
cc_313 N_A_391_388#_c_409_n N_SUM_c_563_n 0.00394508f $X=3.405 $Y=1.025 $X2=0
+ $Y2=0
cc_314 N_A_391_388#_c_411_n N_SUM_c_563_n 0.00361918f $X=4.355 $Y=1.492 $X2=0
+ $Y2=0
cc_315 N_A_391_388#_c_413_n N_SUM_c_559_n 0.00127013f $X=4.355 $Y=1.765 $X2=0
+ $Y2=0
cc_316 N_A_391_388#_c_405_n N_SUM_c_559_n 0.00438312f $X=4.405 $Y=1.22 $X2=0
+ $Y2=0
cc_317 N_A_391_388#_c_457_p N_SUM_c_559_n 0.0256364f $X=4.165 $Y=1.385 $X2=0
+ $Y2=0
cc_318 N_A_391_388#_c_411_n N_SUM_c_559_n 0.0067931f $X=4.355 $Y=1.492 $X2=0
+ $Y2=0
cc_319 N_A_391_388#_c_412_n N_SUM_c_561_n 0.00681625f $X=3.905 $Y=1.765 $X2=0
+ $Y2=0
cc_320 N_A_391_388#_c_413_n N_SUM_c_561_n 0.0163825f $X=4.355 $Y=1.765 $X2=0
+ $Y2=0
cc_321 N_A_391_388#_c_414_n N_SUM_c_561_n 0.00983127f $X=3.32 $Y=2.045 $X2=0
+ $Y2=0
cc_322 N_A_391_388#_c_408_n N_SUM_c_561_n 0.00362727f $X=3.405 $Y=1.92 $X2=0
+ $Y2=0
cc_323 N_A_391_388#_c_457_p N_SUM_c_561_n 0.0202968f $X=4.165 $Y=1.385 $X2=0
+ $Y2=0
cc_324 N_A_391_388#_c_411_n N_SUM_c_561_n 0.00483958f $X=4.355 $Y=1.492 $X2=0
+ $Y2=0
cc_325 N_A_391_388#_c_413_n N_COUT_c_594_n 2.55864e-19 $X=4.355 $Y=1.765 $X2=0
+ $Y2=0
cc_326 N_A_391_388#_c_405_n COUT 0.00104911f $X=4.405 $Y=1.22 $X2=0 $Y2=0
cc_327 N_A_391_388#_c_404_n N_VGND_c_626_n 0.0123991f $X=3.925 $Y=1.22 $X2=0
+ $Y2=0
cc_328 N_A_391_388#_c_405_n N_VGND_c_626_n 0.00143104f $X=4.405 $Y=1.22 $X2=0
+ $Y2=0
cc_329 N_A_391_388#_c_457_p N_VGND_c_626_n 0.0104044f $X=4.165 $Y=1.385 $X2=0
+ $Y2=0
cc_330 N_A_391_388#_c_410_n N_VGND_c_626_n 0.00546815f $X=3.815 $Y=1.385 $X2=0
+ $Y2=0
cc_331 N_A_391_388#_c_404_n N_VGND_c_627_n 0.00143325f $X=3.925 $Y=1.22 $X2=0
+ $Y2=0
cc_332 N_A_391_388#_c_405_n N_VGND_c_627_n 0.0106835f $X=4.405 $Y=1.22 $X2=0
+ $Y2=0
cc_333 N_A_391_388#_c_404_n N_VGND_c_635_n 0.00383152f $X=3.925 $Y=1.22 $X2=0
+ $Y2=0
cc_334 N_A_391_388#_c_405_n N_VGND_c_635_n 0.00383152f $X=4.405 $Y=1.22 $X2=0
+ $Y2=0
cc_335 N_A_391_388#_c_404_n N_VGND_c_639_n 0.00758019f $X=3.925 $Y=1.22 $X2=0
+ $Y2=0
cc_336 N_A_391_388#_c_405_n N_VGND_c_639_n 0.00758019f $X=4.405 $Y=1.22 $X2=0
+ $Y2=0
cc_337 N_A_391_388#_c_406_n N_A_278_74#_M1016_d 0.0091494f $X=3.32 $Y=1.025
+ $X2=0 $Y2=0
cc_338 N_A_391_388#_c_483_p N_A_278_74#_c_697_n 0.0140951f $X=2.72 $Y=0.85 $X2=0
+ $Y2=0
cc_339 N_A_391_388#_c_483_p N_A_278_74#_c_698_n 0.0129062f $X=2.72 $Y=0.85 $X2=0
+ $Y2=0
cc_340 N_A_391_388#_M1016_s N_A_278_74#_c_699_n 0.00297651f $X=2.575 $Y=0.615
+ $X2=0 $Y2=0
cc_341 N_A_391_388#_c_404_n N_A_278_74#_c_699_n 6.04331e-19 $X=3.925 $Y=1.22
+ $X2=0 $Y2=0
cc_342 N_A_391_388#_c_483_p N_A_278_74#_c_699_n 0.0124436f $X=2.72 $Y=0.85 $X2=0
+ $Y2=0
cc_343 N_A_391_388#_c_406_n N_A_278_74#_c_699_n 0.00339819f $X=3.32 $Y=1.025
+ $X2=0 $Y2=0
cc_344 N_A_391_388#_c_404_n N_A_278_74#_c_701_n 0.0013469f $X=3.925 $Y=1.22
+ $X2=0 $Y2=0
cc_345 N_A_391_388#_c_406_n N_A_278_74#_c_701_n 0.0214975f $X=3.32 $Y=1.025
+ $X2=0 $Y2=0
cc_346 N_VPWR_M1011_s N_SUM_c_559_n 0.00298305f $X=4.43 $Y=1.84 $X2=0 $Y2=0
cc_347 N_SUM_c_559_n N_COUT_c_594_n 0.0128877f $X=4.59 $Y=1.82 $X2=0 $Y2=0
cc_348 N_SUM_c_563_n COUT 0.0119219f $X=4.505 $Y=0.965 $X2=0 $Y2=0
cc_349 N_SUM_c_559_n COUT 0.0479339f $X=4.59 $Y=1.82 $X2=0 $Y2=0
cc_350 N_SUM_c_563_n N_VGND_M1014_s 0.00322251f $X=4.505 $Y=0.965 $X2=0 $Y2=0
cc_351 N_SUM_c_559_n N_VGND_M1014_s 5.69077e-19 $X=4.59 $Y=1.82 $X2=0 $Y2=0
cc_352 N_SUM_c_563_n N_VGND_c_627_n 0.0142284f $X=4.505 $Y=0.965 $X2=0 $Y2=0
cc_353 COUT N_VGND_c_627_n 0.0136308f $X=4.955 $Y=0.47 $X2=0 $Y2=0
cc_354 COUT N_VGND_c_629_n 0.0293763f $X=4.955 $Y=0.47 $X2=0 $Y2=0
cc_355 COUT N_VGND_c_636_n 0.0144922f $X=4.955 $Y=0.47 $X2=0 $Y2=0
cc_356 COUT N_VGND_c_639_n 0.0118826f $X=4.955 $Y=0.47 $X2=0 $Y2=0
cc_357 N_VGND_M1007_d N_A_278_74#_c_697_n 0.00443918f $X=1.82 $Y=0.37 $X2=0
+ $Y2=0
cc_358 N_VGND_c_625_n N_A_278_74#_c_697_n 0.0213709f $X=1.96 $Y=0.515 $X2=0
+ $Y2=0
cc_359 N_VGND_c_639_n N_A_278_74#_c_697_n 0.0221192f $X=5.52 $Y=0 $X2=0 $Y2=0
cc_360 N_VGND_c_625_n N_A_278_74#_c_698_n 0.0138372f $X=1.96 $Y=0.515 $X2=0
+ $Y2=0
cc_361 N_VGND_c_626_n N_A_278_74#_c_699_n 0.0121616f $X=3.71 $Y=0.53 $X2=0 $Y2=0
cc_362 N_VGND_c_634_n N_A_278_74#_c_699_n 0.0561641f $X=3.545 $Y=0 $X2=0 $Y2=0
cc_363 N_VGND_c_639_n N_A_278_74#_c_699_n 0.0315987f $X=5.52 $Y=0 $X2=0 $Y2=0
cc_364 N_VGND_c_625_n N_A_278_74#_c_700_n 0.0150383f $X=1.96 $Y=0.515 $X2=0
+ $Y2=0
cc_365 N_VGND_c_634_n N_A_278_74#_c_700_n 0.0121935f $X=3.545 $Y=0 $X2=0 $Y2=0
cc_366 N_VGND_c_639_n N_A_278_74#_c_700_n 0.00661049f $X=5.52 $Y=0 $X2=0 $Y2=0
cc_367 N_VGND_c_626_n N_A_278_74#_c_701_n 0.0191805f $X=3.71 $Y=0.53 $X2=0 $Y2=0
