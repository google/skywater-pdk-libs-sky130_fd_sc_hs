* File: sky130_fd_sc_hs__o2bb2ai_2.pxi.spice
* Created: Thu Aug 27 21:01:22 2020
* 
x_PM_SKY130_FD_SC_HS__O2BB2AI_2%A1_N N_A1_N_c_97_n N_A1_N_M1004_g N_A1_N_M1006_g
+ N_A1_N_c_99_n N_A1_N_M1012_g N_A1_N_c_100_n N_A1_N_M1018_g N_A1_N_c_101_n
+ N_A1_N_c_107_n N_A1_N_c_114_p N_A1_N_c_108_n N_A1_N_c_155_p N_A1_N_c_115_p
+ N_A1_N_c_102_n A1_N N_A1_N_c_103_n A1_N PM_SKY130_FD_SC_HS__O2BB2AI_2%A1_N
x_PM_SKY130_FD_SC_HS__O2BB2AI_2%A2_N N_A2_N_M1007_g N_A2_N_c_193_n
+ N_A2_N_M1003_g N_A2_N_M1019_g N_A2_N_c_194_n N_A2_N_M1009_g A2_N
+ N_A2_N_c_192_n PM_SKY130_FD_SC_HS__O2BB2AI_2%A2_N
x_PM_SKY130_FD_SC_HS__O2BB2AI_2%A_133_387# N_A_133_387#_M1007_d
+ N_A_133_387#_M1004_d N_A_133_387#_M1009_d N_A_133_387#_c_260_n
+ N_A_133_387#_M1001_g N_A_133_387#_M1000_g N_A_133_387#_c_261_n
+ N_A_133_387#_M1014_g N_A_133_387#_M1005_g N_A_133_387#_c_268_n
+ N_A_133_387#_c_254_n N_A_133_387#_c_255_n N_A_133_387#_c_344_p
+ N_A_133_387#_c_256_n N_A_133_387#_c_257_n N_A_133_387#_c_278_n
+ N_A_133_387#_c_282_n N_A_133_387#_c_258_n N_A_133_387#_c_259_n
+ PM_SKY130_FD_SC_HS__O2BB2AI_2%A_133_387#
x_PM_SKY130_FD_SC_HS__O2BB2AI_2%B1 N_B1_M1008_g N_B1_c_353_n N_B1_M1010_g
+ N_B1_c_354_n N_B1_M1017_g N_B1_M1016_g N_B1_c_356_n N_B1_c_361_n N_B1_c_362_n
+ B1 PM_SKY130_FD_SC_HS__O2BB2AI_2%B1
x_PM_SKY130_FD_SC_HS__O2BB2AI_2%B2 N_B2_c_432_n N_B2_M1002_g N_B2_c_436_n
+ N_B2_M1011_g N_B2_c_437_n N_B2_M1013_g N_B2_c_433_n N_B2_M1015_g B2
+ N_B2_c_435_n PM_SKY130_FD_SC_HS__O2BB2AI_2%B2
x_PM_SKY130_FD_SC_HS__O2BB2AI_2%VPWR N_VPWR_M1004_s N_VPWR_M1003_s
+ N_VPWR_M1018_s N_VPWR_M1014_d N_VPWR_M1017_s N_VPWR_c_487_n N_VPWR_c_488_n
+ N_VPWR_c_489_n N_VPWR_c_490_n N_VPWR_c_491_n N_VPWR_c_492_n N_VPWR_c_493_n
+ N_VPWR_c_494_n VPWR N_VPWR_c_495_n N_VPWR_c_496_n N_VPWR_c_497_n
+ N_VPWR_c_498_n N_VPWR_c_499_n N_VPWR_c_500_n N_VPWR_c_486_n
+ PM_SKY130_FD_SC_HS__O2BB2AI_2%VPWR
x_PM_SKY130_FD_SC_HS__O2BB2AI_2%Y N_Y_M1000_d N_Y_M1001_s N_Y_M1011_d
+ N_Y_c_566_n N_Y_c_572_n N_Y_c_586_n Y Y Y Y Y Y
+ PM_SKY130_FD_SC_HS__O2BB2AI_2%Y
x_PM_SKY130_FD_SC_HS__O2BB2AI_2%A_796_368# N_A_796_368#_M1010_d
+ N_A_796_368#_M1013_s N_A_796_368#_c_611_n N_A_796_368#_c_607_n
+ N_A_796_368#_c_608_n N_A_796_368#_c_614_n
+ PM_SKY130_FD_SC_HS__O2BB2AI_2%A_796_368#
x_PM_SKY130_FD_SC_HS__O2BB2AI_2%VGND N_VGND_M1006_s N_VGND_M1012_s
+ N_VGND_M1008_s N_VGND_M1015_d N_VGND_c_636_n N_VGND_c_637_n N_VGND_c_638_n
+ N_VGND_c_639_n N_VGND_c_640_n VGND N_VGND_c_641_n N_VGND_c_642_n
+ N_VGND_c_643_n N_VGND_c_644_n N_VGND_c_645_n N_VGND_c_646_n N_VGND_c_647_n
+ N_VGND_c_648_n PM_SKY130_FD_SC_HS__O2BB2AI_2%VGND
x_PM_SKY130_FD_SC_HS__O2BB2AI_2%A_134_74# N_A_134_74#_M1006_d
+ N_A_134_74#_M1019_s N_A_134_74#_c_710_n N_A_134_74#_c_708_n
+ N_A_134_74#_c_709_n N_A_134_74#_c_713_n
+ PM_SKY130_FD_SC_HS__O2BB2AI_2%A_134_74#
x_PM_SKY130_FD_SC_HS__O2BB2AI_2%A_518_74# N_A_518_74#_M1000_s
+ N_A_518_74#_M1005_s N_A_518_74#_M1002_s N_A_518_74#_M1016_d
+ N_A_518_74#_c_732_n N_A_518_74#_c_733_n N_A_518_74#_c_734_n
+ N_A_518_74#_c_745_n N_A_518_74#_c_746_n N_A_518_74#_c_735_n
+ N_A_518_74#_c_736_n N_A_518_74#_c_752_n N_A_518_74#_c_737_n
+ N_A_518_74#_c_738_n N_A_518_74#_c_766_n
+ PM_SKY130_FD_SC_HS__O2BB2AI_2%A_518_74#
cc_1 VNB N_A1_N_c_97_n 0.0133514f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.86
cc_2 VNB N_A1_N_M1006_g 0.033863f $X=-0.19 $Y=-0.245 $X2=0.595 $Y2=0.69
cc_3 VNB N_A1_N_c_99_n 0.0160204f $X=-0.19 $Y=-0.245 $X2=1.96 $Y2=1.085
cc_4 VNB N_A1_N_c_100_n 0.0468159f $X=-0.19 $Y=-0.245 $X2=2.205 $Y2=1.765
cc_5 VNB N_A1_N_c_101_n 0.0444554f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=1.465
cc_6 VNB N_A1_N_c_102_n 0.00491898f $X=-0.19 $Y=-0.245 $X2=2.25 $Y2=1.515
cc_7 VNB N_A1_N_c_103_n 0.0131935f $X=-0.19 $Y=-0.245 $X2=0.315 $Y2=1.465
cc_8 VNB A1_N 0.00134219f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.665
cc_9 VNB N_A2_N_M1007_g 0.0323868f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=2.355
cc_10 VNB N_A2_N_M1019_g 0.0339291f $X=-0.19 $Y=-0.245 $X2=1.96 $Y2=0.69
cc_11 VNB A2_N 0.00179472f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=1.465
cc_12 VNB N_A2_N_c_192_n 0.0315554f $X=-0.19 $Y=-0.245 $X2=2.25 $Y2=2.45
cc_13 VNB N_A_133_387#_M1000_g 0.0224193f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=1.465
cc_14 VNB N_A_133_387#_M1005_g 0.0209341f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=2.415
cc_15 VNB N_A_133_387#_c_254_n 0.00267999f $X=-0.19 $Y=-0.245 $X2=2.13 $Y2=1.515
cc_16 VNB N_A_133_387#_c_255_n 0.00262414f $X=-0.19 $Y=-0.245 $X2=2.13 $Y2=1.515
cc_17 VNB N_A_133_387#_c_256_n 0.0264071f $X=-0.19 $Y=-0.245 $X2=0.315 $Y2=1.465
cc_18 VNB N_A_133_387#_c_257_n 0.00454919f $X=-0.19 $Y=-0.245 $X2=2.09 $Y2=1.515
cc_19 VNB N_A_133_387#_c_258_n 0.0140213f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.465
cc_20 VNB N_A_133_387#_c_259_n 0.0782959f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_B1_M1008_g 0.0255172f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=2.355
cc_22 VNB N_B1_c_353_n 0.027063f $X=-0.19 $Y=-0.245 $X2=0.595 $Y2=0.69
cc_23 VNB N_B1_c_354_n 0.0288682f $X=-0.19 $Y=-0.245 $X2=1.96 $Y2=1.085
cc_24 VNB N_B1_M1016_g 0.0337117f $X=-0.19 $Y=-0.245 $X2=2.205 $Y2=2.26
cc_25 VNB N_B1_c_356_n 0.00205059f $X=-0.19 $Y=-0.245 $X2=0.355 $Y2=2.5
cc_26 VNB B1 0.0201105f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=2.415
cc_27 VNB N_B2_c_432_n 0.0176191f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.86
cc_28 VNB N_B2_c_433_n 0.0172889f $X=-0.19 $Y=-0.245 $X2=1.96 $Y2=0.69
cc_29 VNB B2 0.00363541f $X=-0.19 $Y=-0.245 $X2=2.205 $Y2=2.26
cc_30 VNB N_B2_c_435_n 0.0539423f $X=-0.19 $Y=-0.245 $X2=2.25 $Y2=1.68
cc_31 VNB N_VPWR_c_486_n 0.243291f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB Y 0.00205679f $X=-0.19 $Y=-0.245 $X2=2.25 $Y2=2.45
cc_33 VNB N_VGND_c_636_n 0.01317f $X=-0.19 $Y=-0.245 $X2=2.205 $Y2=2.26
cc_34 VNB N_VGND_c_637_n 0.0407813f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=1.465
cc_35 VNB N_VGND_c_638_n 0.0126674f $X=-0.19 $Y=-0.245 $X2=0.82 $Y2=2.535
cc_36 VNB N_VGND_c_639_n 0.00533463f $X=-0.19 $Y=-0.245 $X2=0.65 $Y2=2.517
cc_37 VNB N_VGND_c_640_n 0.00330537f $X=-0.19 $Y=-0.245 $X2=2.13 $Y2=1.515
cc_38 VNB N_VGND_c_641_n 0.0385965f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_39 VNB N_VGND_c_642_n 0.0396346f $X=-0.19 $Y=-0.245 $X2=0.315 $Y2=1.465
cc_40 VNB N_VGND_c_643_n 0.0163741f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_644_n 0.0173909f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_645_n 0.322373f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_646_n 0.00499734f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_647_n 0.00615422f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_VGND_c_648_n 0.00629135f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_A_134_74#_c_708_n 0.0045598f $X=-0.19 $Y=-0.245 $X2=2.205 $Y2=1.765
cc_47 VNB N_A_134_74#_c_709_n 0.00203831f $X=-0.19 $Y=-0.245 $X2=2.205 $Y2=2.26
cc_48 VNB N_A_518_74#_c_732_n 0.00365422f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=1.465
cc_49 VNB N_A_518_74#_c_733_n 0.00459841f $X=-0.19 $Y=-0.245 $X2=0.355 $Y2=2.5
cc_50 VNB N_A_518_74#_c_734_n 0.0037722f $X=-0.19 $Y=-0.245 $X2=2.165 $Y2=2.535
cc_51 VNB N_A_518_74#_c_735_n 0.01028f $X=-0.19 $Y=-0.245 $X2=0.82 $Y2=2.517
cc_52 VNB N_A_518_74#_c_736_n 0.00225496f $X=-0.19 $Y=-0.245 $X2=2.13 $Y2=1.515
cc_53 VNB N_A_518_74#_c_737_n 0.0217561f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_54 VNB N_A_518_74#_c_738_n 0.0177969f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VPB N_A1_N_c_97_n 0.0275201f $X=-0.19 $Y=1.66 $X2=0.59 $Y2=1.86
cc_56 VPB N_A1_N_c_100_n 0.0325987f $X=-0.19 $Y=1.66 $X2=2.205 $Y2=1.765
cc_57 VPB N_A1_N_c_107_n 0.00702792f $X=-0.19 $Y=1.66 $X2=0.355 $Y2=2.5
cc_58 VPB N_A1_N_c_108_n 0.00191956f $X=-0.19 $Y=1.66 $X2=2.25 $Y2=2.45
cc_59 VPB N_A1_N_c_102_n 4.59347e-19 $X=-0.19 $Y=1.66 $X2=2.25 $Y2=1.515
cc_60 VPB A1_N 0.030084f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=1.665
cc_61 VPB N_A2_N_c_193_n 0.016156f $X=-0.19 $Y=1.66 $X2=0.595 $Y2=0.69
cc_62 VPB N_A2_N_c_194_n 0.0195287f $X=-0.19 $Y=1.66 $X2=2.205 $Y2=2.26
cc_63 VPB A2_N 0.00320714f $X=-0.19 $Y=1.66 $X2=0.5 $Y2=1.465
cc_64 VPB N_A2_N_c_192_n 0.0362647f $X=-0.19 $Y=1.66 $X2=2.25 $Y2=2.45
cc_65 VPB N_A_133_387#_c_260_n 0.0176316f $X=-0.19 $Y=1.66 $X2=1.96 $Y2=0.69
cc_66 VPB N_A_133_387#_c_261_n 0.0166679f $X=-0.19 $Y=1.66 $X2=0.355 $Y2=2.5
cc_67 VPB N_A_133_387#_c_259_n 0.0142577f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_68 VPB N_B1_c_353_n 0.0259913f $X=-0.19 $Y=1.66 $X2=0.595 $Y2=0.69
cc_69 VPB N_B1_c_354_n 0.0294994f $X=-0.19 $Y=1.66 $X2=1.96 $Y2=1.085
cc_70 VPB N_B1_c_356_n 7.62107e-19 $X=-0.19 $Y=1.66 $X2=0.355 $Y2=2.5
cc_71 VPB N_B1_c_361_n 0.0124295f $X=-0.19 $Y=1.66 $X2=2.25 $Y2=1.68
cc_72 VPB N_B1_c_362_n 0.00104655f $X=-0.19 $Y=1.66 $X2=2.25 $Y2=2.45
cc_73 VPB B1 0.0105354f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=2.415
cc_74 VPB N_B2_c_436_n 0.0141341f $X=-0.19 $Y=1.66 $X2=0.595 $Y2=1.3
cc_75 VPB N_B2_c_437_n 0.0141341f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_76 VPB N_B2_c_435_n 0.0122492f $X=-0.19 $Y=1.66 $X2=2.25 $Y2=1.68
cc_77 VPB N_VPWR_c_487_n 0.0121899f $X=-0.19 $Y=1.66 $X2=0.65 $Y2=2.5
cc_78 VPB N_VPWR_c_488_n 0.0282875f $X=-0.19 $Y=1.66 $X2=2.165 $Y2=2.535
cc_79 VPB N_VPWR_c_489_n 0.0207138f $X=-0.19 $Y=1.66 $X2=2.25 $Y2=1.68
cc_80 VPB N_VPWR_c_490_n 0.0231703f $X=-0.19 $Y=1.66 $X2=0.82 $Y2=2.517
cc_81 VPB N_VPWR_c_491_n 0.0190074f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_82 VPB N_VPWR_c_492_n 0.00862004f $X=-0.19 $Y=1.66 $X2=0.315 $Y2=1.465
cc_83 VPB N_VPWR_c_493_n 0.0106521f $X=-0.19 $Y=1.66 $X2=0.315 $Y2=1.465
cc_84 VPB N_VPWR_c_494_n 0.0498574f $X=-0.19 $Y=1.66 $X2=2.09 $Y2=1.515
cc_85 VPB N_VPWR_c_495_n 0.0283053f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_86 VPB N_VPWR_c_496_n 0.0174435f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_87 VPB N_VPWR_c_497_n 0.0389302f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_88 VPB N_VPWR_c_498_n 0.00631873f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_89 VPB N_VPWR_c_499_n 0.00614589f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_90 VPB N_VPWR_c_500_n 0.00631973f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_91 VPB N_VPWR_c_486_n 0.0866249f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_92 VPB N_Y_c_566_n 0.00284934f $X=-0.19 $Y=1.66 $X2=2.205 $Y2=2.26
cc_93 VPB Y 0.00237843f $X=-0.19 $Y=1.66 $X2=2.25 $Y2=2.45
cc_94 VPB N_A_796_368#_c_607_n 0.00431993f $X=-0.19 $Y=1.66 $X2=2.205 $Y2=1.765
cc_95 VPB N_A_796_368#_c_608_n 0.00218363f $X=-0.19 $Y=1.66 $X2=2.205 $Y2=2.26
cc_96 N_A1_N_M1006_g N_A2_N_M1007_g 0.0169811f $X=0.595 $Y=0.69 $X2=0 $Y2=0
cc_97 N_A1_N_c_103_n N_A2_N_M1007_g 2.01039e-19 $X=0.315 $Y=1.465 $X2=0 $Y2=0
cc_98 N_A1_N_c_97_n N_A2_N_c_193_n 0.0299763f $X=0.59 $Y=1.86 $X2=0 $Y2=0
cc_99 N_A1_N_c_114_p N_A2_N_c_193_n 0.0128604f $X=2.165 $Y=2.535 $X2=0 $Y2=0
cc_100 N_A1_N_c_115_p N_A2_N_c_193_n 9.65396e-19 $X=0.82 $Y=2.517 $X2=0 $Y2=0
cc_101 N_A1_N_c_99_n N_A2_N_M1019_g 0.0276245f $X=1.96 $Y=1.085 $X2=0 $Y2=0
cc_102 N_A1_N_c_100_n N_A2_N_M1019_g 0.00733936f $X=2.205 $Y=1.765 $X2=0 $Y2=0
cc_103 N_A1_N_c_102_n N_A2_N_M1019_g 5.52541e-19 $X=2.25 $Y=1.515 $X2=0 $Y2=0
cc_104 N_A1_N_c_100_n N_A2_N_c_194_n 0.02291f $X=2.205 $Y=1.765 $X2=0 $Y2=0
cc_105 N_A1_N_c_114_p N_A2_N_c_194_n 0.0133281f $X=2.165 $Y=2.535 $X2=0 $Y2=0
cc_106 N_A1_N_c_108_n N_A2_N_c_194_n 0.00128994f $X=2.25 $Y=2.45 $X2=0 $Y2=0
cc_107 N_A1_N_c_100_n A2_N 0.00153088f $X=2.205 $Y=1.765 $X2=0 $Y2=0
cc_108 N_A1_N_c_108_n A2_N 0.00428267f $X=2.25 $Y=2.45 $X2=0 $Y2=0
cc_109 N_A1_N_c_102_n A2_N 0.0191382f $X=2.25 $Y=1.515 $X2=0 $Y2=0
cc_110 N_A1_N_c_97_n N_A2_N_c_192_n 0.0278903f $X=0.59 $Y=1.86 $X2=0 $Y2=0
cc_111 N_A1_N_c_100_n N_A2_N_c_192_n 0.0204669f $X=2.205 $Y=1.765 $X2=0 $Y2=0
cc_112 N_A1_N_c_108_n N_A2_N_c_192_n 5.6482e-19 $X=2.25 $Y=2.45 $X2=0 $Y2=0
cc_113 N_A1_N_c_102_n N_A2_N_c_192_n 2.63377e-19 $X=2.25 $Y=1.515 $X2=0 $Y2=0
cc_114 N_A1_N_c_114_p N_A_133_387#_M1004_d 0.00264577f $X=2.165 $Y=2.535 $X2=0
+ $Y2=0
cc_115 N_A1_N_c_115_p N_A_133_387#_M1004_d 0.00337106f $X=0.82 $Y=2.517 $X2=0
+ $Y2=0
cc_116 N_A1_N_c_114_p N_A_133_387#_M1009_d 0.0107402f $X=2.165 $Y=2.535 $X2=0
+ $Y2=0
cc_117 N_A1_N_c_100_n N_A_133_387#_c_260_n 0.00930117f $X=2.205 $Y=1.765 $X2=0
+ $Y2=0
cc_118 N_A1_N_c_108_n N_A_133_387#_c_260_n 4.60283e-19 $X=2.25 $Y=2.45 $X2=0
+ $Y2=0
cc_119 N_A1_N_c_97_n N_A_133_387#_c_268_n 0.0219178f $X=0.59 $Y=1.86 $X2=0 $Y2=0
cc_120 N_A1_N_M1006_g N_A_133_387#_c_268_n 0.00125799f $X=0.595 $Y=0.69 $X2=0
+ $Y2=0
cc_121 N_A1_N_c_114_p N_A_133_387#_c_268_n 0.00710646f $X=2.165 $Y=2.535 $X2=0
+ $Y2=0
cc_122 N_A1_N_c_115_p N_A_133_387#_c_268_n 0.00911315f $X=0.82 $Y=2.517 $X2=0
+ $Y2=0
cc_123 N_A1_N_c_103_n N_A_133_387#_c_268_n 0.0248813f $X=0.315 $Y=1.465 $X2=0
+ $Y2=0
cc_124 A1_N N_A_133_387#_c_268_n 0.0317183f $X=0.24 $Y=1.665 $X2=0 $Y2=0
cc_125 N_A1_N_M1006_g N_A_133_387#_c_255_n 0.0102229f $X=0.595 $Y=0.69 $X2=0
+ $Y2=0
cc_126 N_A1_N_c_99_n N_A_133_387#_c_256_n 0.00951367f $X=1.96 $Y=1.085 $X2=0
+ $Y2=0
cc_127 N_A1_N_c_100_n N_A_133_387#_c_256_n 0.0162401f $X=2.205 $Y=1.765 $X2=0
+ $Y2=0
cc_128 N_A1_N_c_102_n N_A_133_387#_c_256_n 0.0274115f $X=2.25 $Y=1.515 $X2=0
+ $Y2=0
cc_129 N_A1_N_c_100_n N_A_133_387#_c_278_n 0.00338465f $X=2.205 $Y=1.765 $X2=0
+ $Y2=0
cc_130 N_A1_N_c_114_p N_A_133_387#_c_278_n 0.0165473f $X=2.165 $Y=2.535 $X2=0
+ $Y2=0
cc_131 N_A1_N_c_108_n N_A_133_387#_c_278_n 0.0256975f $X=2.25 $Y=2.45 $X2=0
+ $Y2=0
cc_132 N_A1_N_c_102_n N_A_133_387#_c_278_n 0.00163364f $X=2.25 $Y=1.515 $X2=0
+ $Y2=0
cc_133 N_A1_N_c_114_p N_A_133_387#_c_282_n 0.039865f $X=2.165 $Y=2.535 $X2=0
+ $Y2=0
cc_134 N_A1_N_c_100_n N_A_133_387#_c_258_n 0.00394852f $X=2.205 $Y=1.765 $X2=0
+ $Y2=0
cc_135 N_A1_N_c_102_n N_A_133_387#_c_258_n 0.0225013f $X=2.25 $Y=1.515 $X2=0
+ $Y2=0
cc_136 N_A1_N_c_100_n N_A_133_387#_c_259_n 0.0220839f $X=2.205 $Y=1.765 $X2=0
+ $Y2=0
cc_137 N_A1_N_c_108_n N_A_133_387#_c_259_n 6.48994e-19 $X=2.25 $Y=2.45 $X2=0
+ $Y2=0
cc_138 N_A1_N_c_102_n N_A_133_387#_c_259_n 0.00134539f $X=2.25 $Y=1.515 $X2=0
+ $Y2=0
cc_139 N_A1_N_c_107_n N_VPWR_M1004_s 0.00425083f $X=0.355 $Y=2.5 $X2=-0.19
+ $Y2=-0.245
cc_140 N_A1_N_c_155_p N_VPWR_M1004_s 0.00506041f $X=0.65 $Y=2.517 $X2=-0.19
+ $Y2=-0.245
cc_141 A1_N N_VPWR_M1004_s 0.0108991f $X=0.24 $Y=1.665 $X2=-0.19 $Y2=-0.245
cc_142 N_A1_N_c_114_p N_VPWR_M1003_s 0.00871704f $X=2.165 $Y=2.535 $X2=0 $Y2=0
cc_143 N_A1_N_c_97_n N_VPWR_c_488_n 0.00620477f $X=0.59 $Y=1.86 $X2=0 $Y2=0
cc_144 N_A1_N_c_107_n N_VPWR_c_488_n 0.0199258f $X=0.355 $Y=2.5 $X2=0 $Y2=0
cc_145 N_A1_N_c_155_p N_VPWR_c_488_n 0.00696308f $X=0.65 $Y=2.517 $X2=0 $Y2=0
cc_146 N_A1_N_c_97_n N_VPWR_c_489_n 0.00356885f $X=0.59 $Y=1.86 $X2=0 $Y2=0
cc_147 N_A1_N_c_155_p N_VPWR_c_489_n 0.00231655f $X=0.65 $Y=2.517 $X2=0 $Y2=0
cc_148 N_A1_N_c_115_p N_VPWR_c_489_n 0.00661977f $X=0.82 $Y=2.517 $X2=0 $Y2=0
cc_149 N_A1_N_c_114_p N_VPWR_c_490_n 0.025623f $X=2.165 $Y=2.535 $X2=0 $Y2=0
cc_150 N_A1_N_c_100_n N_VPWR_c_491_n 0.00758522f $X=2.205 $Y=1.765 $X2=0 $Y2=0
cc_151 N_A1_N_c_108_n N_VPWR_c_491_n 0.0260114f $X=2.25 $Y=2.45 $X2=0 $Y2=0
cc_152 N_A1_N_c_100_n N_VPWR_c_495_n 0.00315618f $X=2.205 $Y=1.765 $X2=0 $Y2=0
cc_153 N_A1_N_c_114_p N_VPWR_c_495_n 0.0104808f $X=2.165 $Y=2.535 $X2=0 $Y2=0
cc_154 N_A1_N_c_97_n N_VPWR_c_486_n 0.00489211f $X=0.59 $Y=1.86 $X2=0 $Y2=0
cc_155 N_A1_N_c_100_n N_VPWR_c_486_n 0.00462577f $X=2.205 $Y=1.765 $X2=0 $Y2=0
cc_156 N_A1_N_c_107_n N_VPWR_c_486_n 9.6483e-19 $X=0.355 $Y=2.5 $X2=0 $Y2=0
cc_157 N_A1_N_c_114_p N_VPWR_c_486_n 0.0233602f $X=2.165 $Y=2.535 $X2=0 $Y2=0
cc_158 N_A1_N_c_155_p N_VPWR_c_486_n 0.0055879f $X=0.65 $Y=2.517 $X2=0 $Y2=0
cc_159 N_A1_N_c_115_p N_VPWR_c_486_n 0.0143022f $X=0.82 $Y=2.517 $X2=0 $Y2=0
cc_160 N_A1_N_c_108_n Y 0.00415444f $X=2.25 $Y=2.45 $X2=0 $Y2=0
cc_161 N_A1_N_c_102_n Y 0.0015446f $X=2.25 $Y=1.515 $X2=0 $Y2=0
cc_162 N_A1_N_M1006_g N_VGND_c_637_n 0.0164257f $X=0.595 $Y=0.69 $X2=0 $Y2=0
cc_163 N_A1_N_c_101_n N_VGND_c_637_n 0.00713769f $X=0.5 $Y=1.465 $X2=0 $Y2=0
cc_164 N_A1_N_c_103_n N_VGND_c_637_n 0.0196148f $X=0.315 $Y=1.465 $X2=0 $Y2=0
cc_165 N_A1_N_c_99_n N_VGND_c_638_n 0.00500836f $X=1.96 $Y=1.085 $X2=0 $Y2=0
cc_166 N_A1_N_M1006_g N_VGND_c_641_n 0.00430908f $X=0.595 $Y=0.69 $X2=0 $Y2=0
cc_167 N_A1_N_c_99_n N_VGND_c_641_n 0.00430908f $X=1.96 $Y=1.085 $X2=0 $Y2=0
cc_168 N_A1_N_M1006_g N_VGND_c_645_n 0.0081951f $X=0.595 $Y=0.69 $X2=0 $Y2=0
cc_169 N_A1_N_c_99_n N_VGND_c_645_n 0.00820555f $X=1.96 $Y=1.085 $X2=0 $Y2=0
cc_170 N_A1_N_M1006_g N_A_134_74#_c_710_n 0.00569679f $X=0.595 $Y=0.69 $X2=0
+ $Y2=0
cc_171 N_A1_N_c_99_n N_A_134_74#_c_708_n 0.00393598f $X=1.96 $Y=1.085 $X2=0
+ $Y2=0
cc_172 N_A1_N_M1006_g N_A_134_74#_c_709_n 0.00327745f $X=0.595 $Y=0.69 $X2=0
+ $Y2=0
cc_173 N_A1_N_c_99_n N_A_134_74#_c_713_n 0.00505485f $X=1.96 $Y=1.085 $X2=0
+ $Y2=0
cc_174 N_A2_N_M1007_g N_A_133_387#_c_268_n 0.00529294f $X=1.025 $Y=0.69 $X2=0
+ $Y2=0
cc_175 N_A2_N_c_193_n N_A_133_387#_c_268_n 0.00329947f $X=1.04 $Y=1.86 $X2=0
+ $Y2=0
cc_176 N_A2_N_M1019_g N_A_133_387#_c_268_n 8.01327e-19 $X=1.53 $Y=0.69 $X2=0
+ $Y2=0
cc_177 N_A2_N_c_194_n N_A_133_387#_c_268_n 3.8712e-19 $X=1.66 $Y=1.86 $X2=0
+ $Y2=0
cc_178 A2_N N_A_133_387#_c_268_n 0.0129615f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_179 N_A2_N_c_192_n N_A_133_387#_c_268_n 0.0155547f $X=1.54 $Y=1.61 $X2=0
+ $Y2=0
cc_180 N_A2_N_M1007_g N_A_133_387#_c_254_n 0.0127505f $X=1.025 $Y=0.69 $X2=0
+ $Y2=0
cc_181 N_A2_N_M1007_g N_A_133_387#_c_255_n 0.00312194f $X=1.025 $Y=0.69 $X2=0
+ $Y2=0
cc_182 N_A2_N_M1019_g N_A_133_387#_c_256_n 0.0128475f $X=1.53 $Y=0.69 $X2=0
+ $Y2=0
cc_183 A2_N N_A_133_387#_c_256_n 0.0206507f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_184 N_A2_N_c_192_n N_A_133_387#_c_256_n 0.00352326f $X=1.54 $Y=1.61 $X2=0
+ $Y2=0
cc_185 N_A2_N_M1007_g N_A_133_387#_c_257_n 0.00307017f $X=1.025 $Y=0.69 $X2=0
+ $Y2=0
cc_186 N_A2_N_M1019_g N_A_133_387#_c_257_n 0.00311703f $X=1.53 $Y=0.69 $X2=0
+ $Y2=0
cc_187 A2_N N_A_133_387#_c_257_n 0.00253019f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_188 N_A2_N_c_192_n N_A_133_387#_c_257_n 0.0052622f $X=1.54 $Y=1.61 $X2=0
+ $Y2=0
cc_189 N_A2_N_c_194_n N_A_133_387#_c_278_n 0.00146443f $X=1.66 $Y=1.86 $X2=0
+ $Y2=0
cc_190 N_A2_N_c_193_n N_A_133_387#_c_282_n 0.0146938f $X=1.04 $Y=1.86 $X2=0
+ $Y2=0
cc_191 N_A2_N_c_194_n N_A_133_387#_c_282_n 0.0127473f $X=1.66 $Y=1.86 $X2=0
+ $Y2=0
cc_192 A2_N N_A_133_387#_c_282_n 0.0284068f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_193 N_A2_N_c_192_n N_A_133_387#_c_282_n 0.00812857f $X=1.54 $Y=1.61 $X2=0
+ $Y2=0
cc_194 N_A2_N_c_193_n N_VPWR_c_489_n 0.00354798f $X=1.04 $Y=1.86 $X2=0 $Y2=0
cc_195 N_A2_N_c_193_n N_VPWR_c_490_n 0.00331853f $X=1.04 $Y=1.86 $X2=0 $Y2=0
cc_196 N_A2_N_c_194_n N_VPWR_c_490_n 0.00331853f $X=1.66 $Y=1.86 $X2=0 $Y2=0
cc_197 N_A2_N_c_194_n N_VPWR_c_495_n 0.00354798f $X=1.66 $Y=1.86 $X2=0 $Y2=0
cc_198 N_A2_N_c_193_n N_VPWR_c_486_n 0.00489211f $X=1.04 $Y=1.86 $X2=0 $Y2=0
cc_199 N_A2_N_c_194_n N_VPWR_c_486_n 0.00489211f $X=1.66 $Y=1.86 $X2=0 $Y2=0
cc_200 N_A2_N_M1007_g N_VGND_c_641_n 0.00278247f $X=1.025 $Y=0.69 $X2=0 $Y2=0
cc_201 N_A2_N_M1019_g N_VGND_c_641_n 0.00278247f $X=1.53 $Y=0.69 $X2=0 $Y2=0
cc_202 N_A2_N_M1007_g N_VGND_c_645_n 0.00354226f $X=1.025 $Y=0.69 $X2=0 $Y2=0
cc_203 N_A2_N_M1019_g N_VGND_c_645_n 0.00354226f $X=1.53 $Y=0.69 $X2=0 $Y2=0
cc_204 N_A2_N_M1007_g N_A_134_74#_c_710_n 0.00719216f $X=1.025 $Y=0.69 $X2=0
+ $Y2=0
cc_205 N_A2_N_M1019_g N_A_134_74#_c_710_n 6.34304e-19 $X=1.53 $Y=0.69 $X2=0
+ $Y2=0
cc_206 N_A2_N_M1007_g N_A_134_74#_c_708_n 0.0104897f $X=1.025 $Y=0.69 $X2=0
+ $Y2=0
cc_207 N_A2_N_M1019_g N_A_134_74#_c_708_n 0.010847f $X=1.53 $Y=0.69 $X2=0 $Y2=0
cc_208 N_A2_N_M1007_g N_A_134_74#_c_709_n 0.00184341f $X=1.025 $Y=0.69 $X2=0
+ $Y2=0
cc_209 N_A2_N_M1007_g N_A_134_74#_c_713_n 5.5881e-19 $X=1.025 $Y=0.69 $X2=0
+ $Y2=0
cc_210 N_A2_N_M1019_g N_A_134_74#_c_713_n 0.00648761f $X=1.53 $Y=0.69 $X2=0
+ $Y2=0
cc_211 N_A_133_387#_M1005_g N_B1_M1008_g 0.017351f $X=3.38 $Y=0.74 $X2=0 $Y2=0
cc_212 N_A_133_387#_c_261_n N_B1_c_353_n 0.0259512f $X=3.365 $Y=1.765 $X2=0
+ $Y2=0
cc_213 N_A_133_387#_c_259_n N_B1_c_353_n 0.0208636f $X=3.365 $Y=1.532 $X2=0
+ $Y2=0
cc_214 N_A_133_387#_c_259_n N_B1_c_356_n 0.00180218f $X=3.365 $Y=1.532 $X2=0
+ $Y2=0
cc_215 N_A_133_387#_c_261_n N_B1_c_362_n 0.001178f $X=3.365 $Y=1.765 $X2=0 $Y2=0
cc_216 N_A_133_387#_c_259_n N_B1_c_362_n 4.32563e-19 $X=3.365 $Y=1.532 $X2=0
+ $Y2=0
cc_217 N_A_133_387#_c_282_n N_VPWR_M1003_s 0.0101043f $X=1.72 $Y=2.115 $X2=0
+ $Y2=0
cc_218 N_A_133_387#_c_260_n N_VPWR_c_491_n 0.0165788f $X=2.9 $Y=1.765 $X2=0
+ $Y2=0
cc_219 N_A_133_387#_c_261_n N_VPWR_c_491_n 5.69408e-19 $X=3.365 $Y=1.765 $X2=0
+ $Y2=0
cc_220 N_A_133_387#_c_258_n N_VPWR_c_491_n 0.0261023f $X=2.67 $Y=1.095 $X2=0
+ $Y2=0
cc_221 N_A_133_387#_c_259_n N_VPWR_c_491_n 0.00280814f $X=3.365 $Y=1.532 $X2=0
+ $Y2=0
cc_222 N_A_133_387#_c_261_n N_VPWR_c_492_n 0.00198318f $X=3.365 $Y=1.765 $X2=0
+ $Y2=0
cc_223 N_A_133_387#_c_260_n N_VPWR_c_496_n 0.00429299f $X=2.9 $Y=1.765 $X2=0
+ $Y2=0
cc_224 N_A_133_387#_c_261_n N_VPWR_c_496_n 0.00461464f $X=3.365 $Y=1.765 $X2=0
+ $Y2=0
cc_225 N_A_133_387#_c_260_n N_VPWR_c_486_n 0.00847864f $X=2.9 $Y=1.765 $X2=0
+ $Y2=0
cc_226 N_A_133_387#_c_261_n N_VPWR_c_486_n 0.00908918f $X=3.365 $Y=1.765 $X2=0
+ $Y2=0
cc_227 N_A_133_387#_c_260_n N_Y_c_566_n 2.83791e-19 $X=2.9 $Y=1.765 $X2=0 $Y2=0
cc_228 N_A_133_387#_c_261_n N_Y_c_566_n 2.97145e-19 $X=3.365 $Y=1.765 $X2=0
+ $Y2=0
cc_229 N_A_133_387#_c_261_n N_Y_c_572_n 0.0180642f $X=3.365 $Y=1.765 $X2=0 $Y2=0
cc_230 N_A_133_387#_M1000_g Y 0.0139043f $X=2.95 $Y=0.74 $X2=0 $Y2=0
cc_231 N_A_133_387#_M1005_g Y 0.00541215f $X=3.38 $Y=0.74 $X2=0 $Y2=0
cc_232 N_A_133_387#_c_258_n Y 0.00600767f $X=2.67 $Y=1.095 $X2=0 $Y2=0
cc_233 N_A_133_387#_c_260_n Y 9.99405e-19 $X=2.9 $Y=1.765 $X2=0 $Y2=0
cc_234 N_A_133_387#_M1000_g Y 0.0040844f $X=2.95 $Y=0.74 $X2=0 $Y2=0
cc_235 N_A_133_387#_c_261_n Y 9.35809e-19 $X=3.365 $Y=1.765 $X2=0 $Y2=0
cc_236 N_A_133_387#_c_258_n Y 0.0326778f $X=2.67 $Y=1.095 $X2=0 $Y2=0
cc_237 N_A_133_387#_c_259_n Y 0.0326411f $X=3.365 $Y=1.532 $X2=0 $Y2=0
cc_238 N_A_133_387#_c_261_n Y 2.73912e-19 $X=3.365 $Y=1.765 $X2=0 $Y2=0
cc_239 N_A_133_387#_M1000_g N_VGND_c_638_n 0.00164546f $X=2.95 $Y=0.74 $X2=0
+ $Y2=0
cc_240 N_A_133_387#_c_256_n N_VGND_c_638_n 0.0196286f $X=2.505 $Y=1.095 $X2=0
+ $Y2=0
cc_241 N_A_133_387#_M1000_g N_VGND_c_642_n 0.00278271f $X=2.95 $Y=0.74 $X2=0
+ $Y2=0
cc_242 N_A_133_387#_M1005_g N_VGND_c_642_n 0.00278271f $X=3.38 $Y=0.74 $X2=0
+ $Y2=0
cc_243 N_A_133_387#_M1000_g N_VGND_c_645_n 0.00358427f $X=2.95 $Y=0.74 $X2=0
+ $Y2=0
cc_244 N_A_133_387#_M1005_g N_VGND_c_645_n 0.00353799f $X=3.38 $Y=0.74 $X2=0
+ $Y2=0
cc_245 N_A_133_387#_c_255_n N_A_134_74#_c_710_n 0.0242411f $X=0.98 $Y=1.19 $X2=0
+ $Y2=0
cc_246 N_A_133_387#_M1007_d N_A_134_74#_c_708_n 0.00262408f $X=1.1 $Y=0.37 $X2=0
+ $Y2=0
cc_247 N_A_133_387#_c_344_p N_A_134_74#_c_708_n 0.0174435f $X=1.24 $Y=0.78 $X2=0
+ $Y2=0
cc_248 N_A_133_387#_c_256_n N_A_134_74#_c_708_n 0.00382546f $X=2.505 $Y=1.095
+ $X2=0 $Y2=0
cc_249 N_A_133_387#_c_256_n N_A_134_74#_c_713_n 0.020073f $X=2.505 $Y=1.095
+ $X2=0 $Y2=0
cc_250 N_A_133_387#_c_258_n N_A_518_74#_M1000_s 0.00259532f $X=2.67 $Y=1.095
+ $X2=-0.19 $Y2=-0.245
cc_251 N_A_133_387#_c_258_n N_A_518_74#_c_732_n 0.0139685f $X=2.67 $Y=1.095
+ $X2=0 $Y2=0
cc_252 N_A_133_387#_c_259_n N_A_518_74#_c_732_n 0.00137098f $X=3.365 $Y=1.532
+ $X2=0 $Y2=0
cc_253 N_A_133_387#_M1000_g N_A_518_74#_c_733_n 0.0144222f $X=2.95 $Y=0.74 $X2=0
+ $Y2=0
cc_254 N_A_133_387#_M1005_g N_A_518_74#_c_733_n 0.0131461f $X=3.38 $Y=0.74 $X2=0
+ $Y2=0
cc_255 N_B1_M1008_g N_B2_c_432_n 0.0307135f $X=3.84 $Y=0.74 $X2=-0.19 $Y2=-0.245
cc_256 N_B1_c_353_n N_B2_c_436_n 0.0282343f $X=3.905 $Y=1.765 $X2=0 $Y2=0
cc_257 N_B1_c_361_n N_B2_c_436_n 0.00683396f $X=4.925 $Y=1.805 $X2=0 $Y2=0
cc_258 N_B1_c_354_n N_B2_c_437_n 0.0128674f $X=5.255 $Y=1.765 $X2=0 $Y2=0
cc_259 N_B1_c_361_n N_B2_c_437_n 0.010691f $X=4.925 $Y=1.805 $X2=0 $Y2=0
cc_260 N_B1_M1016_g N_B2_c_433_n 0.0337897f $X=5.265 $Y=0.74 $X2=0 $Y2=0
cc_261 N_B1_M1008_g B2 8.65119e-19 $X=3.84 $Y=0.74 $X2=0 $Y2=0
cc_262 N_B1_c_353_n B2 6.51756e-19 $X=3.905 $Y=1.765 $X2=0 $Y2=0
cc_263 N_B1_M1016_g B2 5.30633e-19 $X=5.265 $Y=0.74 $X2=0 $Y2=0
cc_264 N_B1_c_356_n B2 0.0090454f $X=3.86 $Y=1.515 $X2=0 $Y2=0
cc_265 N_B1_c_361_n B2 0.0246222f $X=4.925 $Y=1.805 $X2=0 $Y2=0
cc_266 B1 B2 0.0124556f $X=4.955 $Y=1.58 $X2=0 $Y2=0
cc_267 N_B1_c_353_n N_B2_c_435_n 0.0222941f $X=3.905 $Y=1.765 $X2=0 $Y2=0
cc_268 N_B1_c_354_n N_B2_c_435_n 0.018678f $X=5.255 $Y=1.765 $X2=0 $Y2=0
cc_269 N_B1_c_356_n N_B2_c_435_n 0.00257546f $X=3.86 $Y=1.515 $X2=0 $Y2=0
cc_270 N_B1_c_361_n N_B2_c_435_n 0.018045f $X=4.925 $Y=1.805 $X2=0 $Y2=0
cc_271 B1 N_B2_c_435_n 0.00759459f $X=4.955 $Y=1.58 $X2=0 $Y2=0
cc_272 N_B1_c_362_n N_VPWR_M1014_d 0.00149864f $X=4.025 $Y=1.805 $X2=0 $Y2=0
cc_273 N_B1_c_353_n N_VPWR_c_492_n 0.00469236f $X=3.905 $Y=1.765 $X2=0 $Y2=0
cc_274 N_B1_c_354_n N_VPWR_c_494_n 0.00919044f $X=5.255 $Y=1.765 $X2=0 $Y2=0
cc_275 B1 N_VPWR_c_494_n 0.00879213f $X=4.955 $Y=1.58 $X2=0 $Y2=0
cc_276 N_B1_c_353_n N_VPWR_c_497_n 0.0044313f $X=3.905 $Y=1.765 $X2=0 $Y2=0
cc_277 N_B1_c_354_n N_VPWR_c_497_n 0.0044313f $X=5.255 $Y=1.765 $X2=0 $Y2=0
cc_278 N_B1_c_353_n N_VPWR_c_486_n 0.00853716f $X=3.905 $Y=1.765 $X2=0 $Y2=0
cc_279 N_B1_c_354_n N_VPWR_c_486_n 0.00856939f $X=5.255 $Y=1.765 $X2=0 $Y2=0
cc_280 N_B1_c_361_n N_Y_M1011_d 0.00197722f $X=4.925 $Y=1.805 $X2=0 $Y2=0
cc_281 N_B1_c_353_n N_Y_c_572_n 0.0156781f $X=3.905 $Y=1.765 $X2=0 $Y2=0
cc_282 N_B1_c_361_n N_Y_c_572_n 0.023643f $X=4.925 $Y=1.805 $X2=0 $Y2=0
cc_283 N_B1_c_362_n N_Y_c_572_n 0.0174383f $X=4.025 $Y=1.805 $X2=0 $Y2=0
cc_284 N_B1_c_361_n N_Y_c_586_n 0.0151236f $X=4.925 $Y=1.805 $X2=0 $Y2=0
cc_285 N_B1_M1008_g Y 2.22458e-19 $X=3.84 $Y=0.74 $X2=0 $Y2=0
cc_286 N_B1_c_353_n Y 0.00102381f $X=3.905 $Y=1.765 $X2=0 $Y2=0
cc_287 N_B1_c_356_n Y 0.013779f $X=3.86 $Y=1.515 $X2=0 $Y2=0
cc_288 N_B1_c_362_n Y 0.00781912f $X=4.025 $Y=1.805 $X2=0 $Y2=0
cc_289 N_B1_c_361_n N_A_796_368#_M1010_d 0.00198204f $X=4.925 $Y=1.805 $X2=-0.19
+ $Y2=-0.245
cc_290 B1 N_A_796_368#_M1013_s 0.0023915f $X=4.955 $Y=1.58 $X2=0 $Y2=0
cc_291 N_B1_c_353_n N_A_796_368#_c_611_n 0.00508076f $X=3.905 $Y=1.765 $X2=0
+ $Y2=0
cc_292 N_B1_c_354_n N_A_796_368#_c_607_n 0.00332677f $X=5.255 $Y=1.765 $X2=0
+ $Y2=0
cc_293 N_B1_c_353_n N_A_796_368#_c_608_n 0.00314614f $X=3.905 $Y=1.765 $X2=0
+ $Y2=0
cc_294 N_B1_c_354_n N_A_796_368#_c_614_n 0.00931336f $X=5.255 $Y=1.765 $X2=0
+ $Y2=0
cc_295 N_B1_c_361_n N_A_796_368#_c_614_n 0.00102433f $X=4.925 $Y=1.805 $X2=0
+ $Y2=0
cc_296 B1 N_A_796_368#_c_614_n 0.0182342f $X=4.955 $Y=1.58 $X2=0 $Y2=0
cc_297 N_B1_M1008_g N_VGND_c_639_n 0.00293683f $X=3.84 $Y=0.74 $X2=0 $Y2=0
cc_298 N_B1_M1016_g N_VGND_c_640_n 0.00981808f $X=5.265 $Y=0.74 $X2=0 $Y2=0
cc_299 N_B1_M1008_g N_VGND_c_642_n 0.00430908f $X=3.84 $Y=0.74 $X2=0 $Y2=0
cc_300 N_B1_M1016_g N_VGND_c_644_n 0.00383152f $X=5.265 $Y=0.74 $X2=0 $Y2=0
cc_301 N_B1_M1008_g N_VGND_c_645_n 0.00445932f $X=3.84 $Y=0.74 $X2=0 $Y2=0
cc_302 N_B1_M1016_g N_VGND_c_645_n 0.00372886f $X=5.265 $Y=0.74 $X2=0 $Y2=0
cc_303 N_B1_M1008_g N_A_518_74#_c_733_n 0.00332495f $X=3.84 $Y=0.74 $X2=0 $Y2=0
cc_304 N_B1_M1008_g N_A_518_74#_c_745_n 0.00642991f $X=3.84 $Y=0.74 $X2=0 $Y2=0
cc_305 N_B1_M1008_g N_A_518_74#_c_746_n 0.00963801f $X=3.84 $Y=0.74 $X2=0 $Y2=0
cc_306 N_B1_c_353_n N_A_518_74#_c_746_n 4.88557e-19 $X=3.905 $Y=1.765 $X2=0
+ $Y2=0
cc_307 N_B1_c_356_n N_A_518_74#_c_746_n 0.00900162f $X=3.86 $Y=1.515 $X2=0 $Y2=0
cc_308 N_B1_M1008_g N_A_518_74#_c_735_n 0.00333924f $X=3.84 $Y=0.74 $X2=0 $Y2=0
cc_309 N_B1_c_353_n N_A_518_74#_c_735_n 5.28989e-19 $X=3.905 $Y=1.765 $X2=0
+ $Y2=0
cc_310 N_B1_c_356_n N_A_518_74#_c_735_n 0.00667011f $X=3.86 $Y=1.515 $X2=0 $Y2=0
cc_311 N_B1_M1016_g N_A_518_74#_c_752_n 0.0107539f $X=5.265 $Y=0.74 $X2=0 $Y2=0
cc_312 B1 N_A_518_74#_c_752_n 0.0167053f $X=4.955 $Y=1.58 $X2=0 $Y2=0
cc_313 N_B1_c_354_n N_A_518_74#_c_737_n 0.00116012f $X=5.255 $Y=1.765 $X2=0
+ $Y2=0
cc_314 N_B1_M1016_g N_A_518_74#_c_737_n 0.00412046f $X=5.265 $Y=0.74 $X2=0 $Y2=0
cc_315 B1 N_A_518_74#_c_737_n 0.0124005f $X=4.955 $Y=1.58 $X2=0 $Y2=0
cc_316 N_B1_M1016_g N_A_518_74#_c_738_n 0.00130587f $X=5.265 $Y=0.74 $X2=0 $Y2=0
cc_317 N_B2_c_436_n N_VPWR_c_497_n 0.00278257f $X=4.355 $Y=1.765 $X2=0 $Y2=0
cc_318 N_B2_c_437_n N_VPWR_c_497_n 0.00278257f $X=4.805 $Y=1.765 $X2=0 $Y2=0
cc_319 N_B2_c_436_n N_VPWR_c_486_n 0.00353905f $X=4.355 $Y=1.765 $X2=0 $Y2=0
cc_320 N_B2_c_437_n N_VPWR_c_486_n 0.00353905f $X=4.805 $Y=1.765 $X2=0 $Y2=0
cc_321 N_B2_c_436_n N_Y_c_572_n 0.0105474f $X=4.355 $Y=1.765 $X2=0 $Y2=0
cc_322 N_B2_c_436_n N_A_796_368#_c_611_n 0.00631535f $X=4.355 $Y=1.765 $X2=0
+ $Y2=0
cc_323 N_B2_c_437_n N_A_796_368#_c_611_n 5.2336e-19 $X=4.805 $Y=1.765 $X2=0
+ $Y2=0
cc_324 N_B2_c_436_n N_A_796_368#_c_607_n 0.00879888f $X=4.355 $Y=1.765 $X2=0
+ $Y2=0
cc_325 N_B2_c_437_n N_A_796_368#_c_607_n 0.0125587f $X=4.805 $Y=1.765 $X2=0
+ $Y2=0
cc_326 N_B2_c_436_n N_A_796_368#_c_608_n 0.00171238f $X=4.355 $Y=1.765 $X2=0
+ $Y2=0
cc_327 N_B2_c_436_n N_A_796_368#_c_614_n 5.68027e-19 $X=4.355 $Y=1.765 $X2=0
+ $Y2=0
cc_328 N_B2_c_437_n N_A_796_368#_c_614_n 0.00950859f $X=4.805 $Y=1.765 $X2=0
+ $Y2=0
cc_329 N_B2_c_432_n N_VGND_c_639_n 0.00773369f $X=4.34 $Y=1.22 $X2=0 $Y2=0
cc_330 N_B2_c_433_n N_VGND_c_639_n 4.19327e-19 $X=4.82 $Y=1.22 $X2=0 $Y2=0
cc_331 N_B2_c_432_n N_VGND_c_640_n 4.00885e-19 $X=4.34 $Y=1.22 $X2=0 $Y2=0
cc_332 N_B2_c_433_n N_VGND_c_640_n 0.00702777f $X=4.82 $Y=1.22 $X2=0 $Y2=0
cc_333 N_B2_c_432_n N_VGND_c_643_n 0.00383152f $X=4.34 $Y=1.22 $X2=0 $Y2=0
cc_334 N_B2_c_433_n N_VGND_c_643_n 0.00383152f $X=4.82 $Y=1.22 $X2=0 $Y2=0
cc_335 N_B2_c_432_n N_VGND_c_645_n 0.00384446f $X=4.34 $Y=1.22 $X2=0 $Y2=0
cc_336 N_B2_c_433_n N_VGND_c_645_n 0.00369749f $X=4.82 $Y=1.22 $X2=0 $Y2=0
cc_337 N_B2_c_432_n N_A_518_74#_c_745_n 6.25243e-19 $X=4.34 $Y=1.22 $X2=0 $Y2=0
cc_338 N_B2_c_432_n N_A_518_74#_c_746_n 0.0124209f $X=4.34 $Y=1.22 $X2=0 $Y2=0
cc_339 B2 N_A_518_74#_c_746_n 0.00730648f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_340 N_B2_c_432_n N_A_518_74#_c_735_n 5.68029e-19 $X=4.34 $Y=1.22 $X2=0 $Y2=0
cc_341 N_B2_c_432_n N_A_518_74#_c_736_n 2.53282e-19 $X=4.34 $Y=1.22 $X2=0 $Y2=0
cc_342 N_B2_c_433_n N_A_518_74#_c_736_n 2.53282e-19 $X=4.82 $Y=1.22 $X2=0 $Y2=0
cc_343 N_B2_c_433_n N_A_518_74#_c_752_n 0.0162195f $X=4.82 $Y=1.22 $X2=0 $Y2=0
cc_344 N_B2_c_433_n N_A_518_74#_c_737_n 5.82428e-19 $X=4.82 $Y=1.22 $X2=0 $Y2=0
cc_345 B2 N_A_518_74#_c_766_n 0.0177874f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_346 N_B2_c_435_n N_A_518_74#_c_766_n 0.00105185f $X=4.805 $Y=1.492 $X2=0
+ $Y2=0
cc_347 N_VPWR_c_491_n N_Y_c_566_n 0.0289149f $X=2.67 $Y=1.985 $X2=0 $Y2=0
cc_348 N_VPWR_c_492_n N_Y_c_566_n 0.0233333f $X=3.625 $Y=2.485 $X2=0 $Y2=0
cc_349 N_VPWR_c_496_n N_Y_c_566_n 0.0126277f $X=3.46 $Y=3.33 $X2=0 $Y2=0
cc_350 N_VPWR_c_486_n N_Y_c_566_n 0.0104521f $X=5.52 $Y=3.33 $X2=0 $Y2=0
cc_351 N_VPWR_M1014_d N_Y_c_572_n 0.0114652f $X=3.44 $Y=1.84 $X2=0 $Y2=0
cc_352 N_VPWR_c_492_n N_Y_c_572_n 0.022455f $X=3.625 $Y=2.485 $X2=0 $Y2=0
cc_353 N_VPWR_c_491_n Y 0.00977851f $X=2.67 $Y=1.985 $X2=0 $Y2=0
cc_354 N_VPWR_c_494_n N_A_796_368#_c_607_n 0.012272f $X=5.48 $Y=2.115 $X2=0
+ $Y2=0
cc_355 N_VPWR_c_497_n N_A_796_368#_c_607_n 0.0594312f $X=5.395 $Y=3.33 $X2=0
+ $Y2=0
cc_356 N_VPWR_c_486_n N_A_796_368#_c_607_n 0.0328875f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_357 N_VPWR_c_492_n N_A_796_368#_c_608_n 0.0116611f $X=3.625 $Y=2.485 $X2=0
+ $Y2=0
cc_358 N_VPWR_c_497_n N_A_796_368#_c_608_n 0.0235381f $X=5.395 $Y=3.33 $X2=0
+ $Y2=0
cc_359 N_VPWR_c_486_n N_A_796_368#_c_608_n 0.0126899f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_360 N_VPWR_c_494_n N_A_796_368#_c_614_n 0.0566253f $X=5.48 $Y=2.115 $X2=0
+ $Y2=0
cc_361 N_Y_c_572_n N_A_796_368#_M1010_d 0.00395925f $X=4.465 $Y=2.145 $X2=-0.19
+ $Y2=-0.245
cc_362 N_Y_c_572_n N_A_796_368#_c_611_n 0.017171f $X=4.465 $Y=2.145 $X2=0 $Y2=0
cc_363 N_Y_M1011_d N_A_796_368#_c_607_n 0.00197722f $X=4.43 $Y=1.84 $X2=0 $Y2=0
cc_364 N_Y_c_572_n N_A_796_368#_c_607_n 0.00286566f $X=4.465 $Y=2.145 $X2=0
+ $Y2=0
cc_365 N_Y_c_586_n N_A_796_368#_c_607_n 0.014149f $X=4.58 $Y=2.225 $X2=0 $Y2=0
cc_366 N_Y_M1000_d N_A_518_74#_c_733_n 0.00176461f $X=3.025 $Y=0.37 $X2=0 $Y2=0
cc_367 Y N_A_518_74#_c_733_n 0.0143448f $X=3.035 $Y=0.84 $X2=0 $Y2=0
cc_368 Y N_A_518_74#_c_735_n 0.00157293f $X=3.035 $Y=0.84 $X2=0 $Y2=0
cc_369 N_VGND_c_638_n N_A_134_74#_c_708_n 0.0117551f $X=2.175 $Y=0.66 $X2=0
+ $Y2=0
cc_370 N_VGND_c_641_n N_A_134_74#_c_708_n 0.0613668f $X=2.08 $Y=0 $X2=0 $Y2=0
cc_371 N_VGND_c_645_n N_A_134_74#_c_708_n 0.0341446f $X=5.52 $Y=0 $X2=0 $Y2=0
cc_372 N_VGND_c_637_n N_A_134_74#_c_709_n 0.011924f $X=0.31 $Y=0.515 $X2=0 $Y2=0
cc_373 N_VGND_c_641_n N_A_134_74#_c_709_n 0.0234809f $X=2.08 $Y=0 $X2=0 $Y2=0
cc_374 N_VGND_c_645_n N_A_134_74#_c_709_n 0.0126009f $X=5.52 $Y=0 $X2=0 $Y2=0
cc_375 N_VGND_c_638_n N_A_518_74#_c_732_n 0.025902f $X=2.175 $Y=0.66 $X2=0 $Y2=0
cc_376 N_VGND_c_639_n N_A_518_74#_c_733_n 0.011924f $X=4.125 $Y=0.55 $X2=0 $Y2=0
cc_377 N_VGND_c_642_n N_A_518_74#_c_733_n 0.0638649f $X=3.96 $Y=0 $X2=0 $Y2=0
cc_378 N_VGND_c_645_n N_A_518_74#_c_733_n 0.0354046f $X=5.52 $Y=0 $X2=0 $Y2=0
cc_379 N_VGND_c_638_n N_A_518_74#_c_734_n 0.0119579f $X=2.175 $Y=0.66 $X2=0
+ $Y2=0
cc_380 N_VGND_c_642_n N_A_518_74#_c_734_n 0.0176866f $X=3.96 $Y=0 $X2=0 $Y2=0
cc_381 N_VGND_c_645_n N_A_518_74#_c_734_n 0.00967523f $X=5.52 $Y=0 $X2=0 $Y2=0
cc_382 N_VGND_M1008_s N_A_518_74#_c_746_n 0.0101164f $X=3.915 $Y=0.37 $X2=0
+ $Y2=0
cc_383 N_VGND_c_639_n N_A_518_74#_c_746_n 0.0205261f $X=4.125 $Y=0.55 $X2=0
+ $Y2=0
cc_384 N_VGND_c_645_n N_A_518_74#_c_746_n 0.0113542f $X=5.52 $Y=0 $X2=0 $Y2=0
cc_385 N_VGND_c_639_n N_A_518_74#_c_736_n 0.0121832f $X=4.125 $Y=0.55 $X2=0
+ $Y2=0
cc_386 N_VGND_c_640_n N_A_518_74#_c_736_n 0.0097355f $X=5.04 $Y=0.515 $X2=0
+ $Y2=0
cc_387 N_VGND_c_643_n N_A_518_74#_c_736_n 0.00970617f $X=4.87 $Y=0 $X2=0 $Y2=0
cc_388 N_VGND_c_645_n N_A_518_74#_c_736_n 0.00804326f $X=5.52 $Y=0 $X2=0 $Y2=0
cc_389 N_VGND_M1015_d N_A_518_74#_c_752_n 0.00460082f $X=4.895 $Y=0.37 $X2=0
+ $Y2=0
cc_390 N_VGND_c_640_n N_A_518_74#_c_752_n 0.0181964f $X=5.04 $Y=0.515 $X2=0
+ $Y2=0
cc_391 N_VGND_c_645_n N_A_518_74#_c_752_n 0.0101909f $X=5.52 $Y=0 $X2=0 $Y2=0
cc_392 N_VGND_c_645_n N_A_518_74#_c_737_n 0.00293094f $X=5.52 $Y=0 $X2=0 $Y2=0
cc_393 N_VGND_c_640_n N_A_518_74#_c_738_n 0.00974948f $X=5.04 $Y=0.515 $X2=0
+ $Y2=0
cc_394 N_VGND_c_644_n N_A_518_74#_c_738_n 0.011066f $X=5.52 $Y=0 $X2=0 $Y2=0
cc_395 N_VGND_c_645_n N_A_518_74#_c_738_n 0.00915947f $X=5.52 $Y=0 $X2=0 $Y2=0
