* File: sky130_fd_sc_hs__nor2b_2.spice
* Created: Thu Aug 27 20:53:35 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hs__nor2b_2.pex.spice"
.subckt sky130_fd_sc_hs__nor2b_2  VNB VPB B_N A VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A	A
* B_N	B_N
* VPB	VPB
* VNB	VNB
MM1005 N_VGND_M1005_d N_B_N_M1005_g N_A_27_392#_M1005_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.151513 AS=0.1824 PD=1.10841 PS=1.85 NRD=20.148 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75002.2 A=0.096 P=1.58 MULT=1
MM1000 N_Y_M1000_d N_A_27_392#_M1000_g N_VGND_M1005_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.1221 AS=0.175187 PD=1.07 PS=1.28159 NRD=0 NRS=11.34 M=1 R=4.93333
+ SA=75000.7 SB=75001.6 A=0.111 P=1.78 MULT=1
MM1006 N_Y_M1000_d N_A_27_392#_M1006_g N_VGND_M1006_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1221 AS=0.111 PD=1.07 PS=1.04 NRD=8.1 NRS=3.24 M=1 R=4.93333 SA=75001.2
+ SB=75001.2 A=0.111 P=1.78 MULT=1
MM1008 N_Y_M1008_d N_A_M1008_g N_VGND_M1006_s VNB NLOWVT L=0.15 W=0.74 AD=0.1221
+ AS=0.111 PD=1.07 PS=1.04 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.7 SB=75000.7
+ A=0.111 P=1.78 MULT=1
MM1009 N_Y_M1008_d N_A_M1009_g N_VGND_M1009_s VNB NLOWVT L=0.15 W=0.74 AD=0.1221
+ AS=0.2257 PD=1.07 PS=2.09 NRD=8.1 NRS=3.24 M=1 R=4.93333 SA=75002.2 SB=75000.2
+ A=0.111 P=1.78 MULT=1
MM1007 N_VPWR_M1007_d N_B_N_M1007_g N_A_27_392#_M1007_s VPB PSHORT L=0.15 W=1
+ AD=0.295 AS=0.29 PD=2.59 PS=2.58 NRD=1.9503 NRS=1.9503 M=1 R=6.66667
+ SA=75000.2 SB=75000.2 A=0.15 P=2.3 MULT=1
MM1001 N_Y_M1001_d N_A_27_392#_M1001_g N_A_228_368#_M1001_s VPB PSHORT L=0.15
+ W=1.12 AD=0.168 AS=0.3304 PD=1.42 PS=2.83 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75001.6 A=0.168 P=2.54 MULT=1
MM1002 N_Y_M1001_d N_A_27_392#_M1002_g N_A_228_368#_M1002_s VPB PSHORT L=0.15
+ W=1.12 AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.7 SB=75001.1 A=0.168 P=2.54 MULT=1
MM1003 N_VPWR_M1003_d N_A_M1003_g N_A_228_368#_M1002_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.1 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1004 N_VPWR_M1003_d N_A_M1004_g N_A_228_368#_M1004_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.3248 PD=1.42 PS=2.82 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.6 SB=75000.2 A=0.168 P=2.54 MULT=1
DX10_noxref VNB VPB NWDIODE A=6.9564 P=11.2
*
.include "sky130_fd_sc_hs__nor2b_2.pxi.spice"
*
.ends
*
*
