* File: sky130_fd_sc_hs__o21a_4.pxi.spice
* Created: Tue Sep  1 20:14:24 2020
* 
x_PM_SKY130_FD_SC_HS__O21A_4%A2 N_A2_M1005_g N_A2_c_104_n N_A2_M1015_g
+ N_A2_M1006_g N_A2_c_105_n N_A2_M1018_g A2 N_A2_c_102_n N_A2_c_103_n
+ PM_SKY130_FD_SC_HS__O21A_4%A2
x_PM_SKY130_FD_SC_HS__O21A_4%A1 N_A1_c_152_n N_A1_c_153_n N_A1_M1010_g
+ N_A1_c_161_n N_A1_M1017_g N_A1_c_155_n N_A1_c_156_n N_A1_c_157_n N_A1_M1019_g
+ N_A1_M1012_g A1 PM_SKY130_FD_SC_HS__O21A_4%A1
x_PM_SKY130_FD_SC_HS__O21A_4%B1 N_B1_M1009_g N_B1_c_221_n N_B1_M1003_g
+ N_B1_M1014_g N_B1_c_222_n N_B1_M1004_g B1 B1 N_B1_c_220_n
+ PM_SKY130_FD_SC_HS__O21A_4%B1
x_PM_SKY130_FD_SC_HS__O21A_4%A_216_387# N_A_216_387#_M1009_s
+ N_A_216_387#_M1015_d N_A_216_387#_M1003_s N_A_216_387#_c_281_n
+ N_A_216_387#_M1000_g N_A_216_387#_c_270_n N_A_216_387#_M1001_g
+ N_A_216_387#_c_282_n N_A_216_387#_M1011_g N_A_216_387#_c_271_n
+ N_A_216_387#_M1002_g N_A_216_387#_c_283_n N_A_216_387#_M1013_g
+ N_A_216_387#_c_272_n N_A_216_387#_M1007_g N_A_216_387#_c_284_n
+ N_A_216_387#_M1016_g N_A_216_387#_c_273_n N_A_216_387#_M1008_g
+ N_A_216_387#_c_288_n N_A_216_387#_c_274_n N_A_216_387#_c_275_n
+ N_A_216_387#_c_276_n N_A_216_387#_c_310_n N_A_216_387#_c_277_n
+ N_A_216_387#_c_278_n N_A_216_387#_c_290_n N_A_216_387#_c_286_n
+ N_A_216_387#_c_279_n N_A_216_387#_c_280_n
+ PM_SKY130_FD_SC_HS__O21A_4%A_216_387#
x_PM_SKY130_FD_SC_HS__O21A_4%VPWR N_VPWR_M1017_d N_VPWR_M1019_d N_VPWR_M1004_d
+ N_VPWR_M1011_d N_VPWR_M1016_d N_VPWR_c_413_n N_VPWR_c_414_n N_VPWR_c_415_n
+ N_VPWR_c_416_n N_VPWR_c_417_n N_VPWR_c_418_n N_VPWR_c_419_n N_VPWR_c_420_n
+ N_VPWR_c_421_n VPWR N_VPWR_c_422_n N_VPWR_c_423_n N_VPWR_c_424_n
+ N_VPWR_c_425_n N_VPWR_c_426_n N_VPWR_c_412_n PM_SKY130_FD_SC_HS__O21A_4%VPWR
x_PM_SKY130_FD_SC_HS__O21A_4%A_116_387# N_A_116_387#_M1017_s
+ N_A_116_387#_M1018_s N_A_116_387#_c_484_n N_A_116_387#_c_482_n
+ N_A_116_387#_c_483_n N_A_116_387#_c_490_n
+ PM_SKY130_FD_SC_HS__O21A_4%A_116_387#
x_PM_SKY130_FD_SC_HS__O21A_4%X N_X_M1001_s N_X_M1007_s N_X_M1000_s N_X_M1013_s
+ N_X_c_507_n N_X_c_517_n N_X_c_503_n N_X_c_508_n N_X_c_509_n N_X_c_531_n
+ N_X_c_510_n N_X_c_504_n N_X_c_505_n N_X_c_544_n X PM_SKY130_FD_SC_HS__O21A_4%X
x_PM_SKY130_FD_SC_HS__O21A_4%A_27_125# N_A_27_125#_M1010_s N_A_27_125#_M1005_d
+ N_A_27_125#_M1012_s N_A_27_125#_M1014_d N_A_27_125#_c_573_n
+ N_A_27_125#_c_574_n N_A_27_125#_c_575_n N_A_27_125#_c_576_n
+ N_A_27_125#_c_577_n N_A_27_125#_c_578_n N_A_27_125#_c_579_n
+ N_A_27_125#_c_580_n N_A_27_125#_c_581_n N_A_27_125#_c_582_n
+ PM_SKY130_FD_SC_HS__O21A_4%A_27_125#
x_PM_SKY130_FD_SC_HS__O21A_4%VGND N_VGND_M1010_d N_VGND_M1006_s N_VGND_M1001_d
+ N_VGND_M1002_d N_VGND_M1008_d N_VGND_c_640_n N_VGND_c_641_n N_VGND_c_642_n
+ N_VGND_c_643_n N_VGND_c_644_n N_VGND_c_645_n VGND N_VGND_c_646_n
+ N_VGND_c_647_n N_VGND_c_648_n N_VGND_c_649_n N_VGND_c_650_n N_VGND_c_651_n
+ N_VGND_c_652_n N_VGND_c_653_n N_VGND_c_654_n N_VGND_c_655_n
+ PM_SKY130_FD_SC_HS__O21A_4%VGND
cc_1 VNB N_A2_M1005_g 0.0186294f $X=-0.19 $Y=-0.245 $X2=1 $Y2=0.945
cc_2 VNB N_A2_M1006_g 0.0202457f $X=-0.19 $Y=-0.245 $X2=1.43 $Y2=0.945
cc_3 VNB N_A2_c_102_n 0.00175162f $X=-0.19 $Y=-0.245 $X2=1.34 $Y2=1.61
cc_4 VNB N_A2_c_103_n 0.0305755f $X=-0.19 $Y=-0.245 $X2=1.43 $Y2=1.652
cc_5 VNB N_A1_c_152_n 0.00867293f $X=-0.19 $Y=-0.245 $X2=1 $Y2=1.445
cc_6 VNB N_A1_c_153_n 0.0194277f $X=-0.19 $Y=-0.245 $X2=1 $Y2=0.945
cc_7 VNB N_A1_M1010_g 0.0364999f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=2.435
cc_8 VNB N_A1_c_155_n 0.108819f $X=-0.19 $Y=-0.245 $X2=1.43 $Y2=0.945
cc_9 VNB N_A1_c_156_n 0.012806f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A1_c_157_n 0.0170588f $X=-0.19 $Y=-0.245 $X2=1.455 $Y2=1.86
cc_11 VNB N_A1_M1012_g 0.0331968f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=1.652
cc_12 VNB A1 0.0046028f $X=-0.19 $Y=-0.245 $X2=1.34 $Y2=1.61
cc_13 VNB N_B1_M1009_g 0.0191682f $X=-0.19 $Y=-0.245 $X2=1 $Y2=0.945
cc_14 VNB N_B1_M1014_g 0.0205347f $X=-0.19 $Y=-0.245 $X2=1.43 $Y2=0.945
cc_15 VNB B1 0.0021003f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_B1_c_220_n 0.0320054f $X=-0.19 $Y=-0.245 $X2=1.455 $Y2=1.652
cc_17 VNB N_A_216_387#_c_270_n 0.0198604f $X=-0.19 $Y=-0.245 $X2=1.455 $Y2=2.435
cc_18 VNB N_A_216_387#_c_271_n 0.0164674f $X=-0.19 $Y=-0.245 $X2=1.34 $Y2=1.652
cc_19 VNB N_A_216_387#_c_272_n 0.0166181f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_216_387#_c_273_n 0.021272f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_216_387#_c_274_n 0.00200913f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_216_387#_c_275_n 0.00762265f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_216_387#_c_276_n 0.00269748f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_216_387#_c_277_n 0.00169712f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_216_387#_c_278_n 0.00982261f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_216_387#_c_279_n 0.00906033f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_216_387#_c_280_n 0.154098f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_VPWR_c_412_n 0.243291f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_X_c_503_n 0.00215307f $X=-0.19 $Y=-0.245 $X2=1.34 $Y2=1.61
cc_30 VNB N_X_c_504_n 0.00178908f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_X_c_505_n 0.00177379f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB X 0.00943489f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_27_125#_c_573_n 0.022896f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.58
cc_34 VNB N_A_27_125#_c_574_n 0.00568431f $X=-0.19 $Y=-0.245 $X2=1 $Y2=1.652
cc_35 VNB N_A_27_125#_c_575_n 0.0125745f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=1.652
cc_36 VNB N_A_27_125#_c_576_n 0.00206719f $X=-0.19 $Y=-0.245 $X2=1.34 $Y2=1.61
cc_37 VNB N_A_27_125#_c_577_n 0.00867474f $X=-0.19 $Y=-0.245 $X2=1.455 $Y2=1.652
cc_38 VNB N_A_27_125#_c_578_n 8.44865e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_27_125#_c_579_n 0.0214365f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_27_125#_c_580_n 0.00249092f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_27_125#_c_581_n 0.00923286f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_27_125#_c_582_n 0.00177457f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_640_n 0.00825723f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=1.652
cc_44 VNB N_VGND_c_641_n 0.00930184f $X=-0.19 $Y=-0.245 $X2=1.43 $Y2=1.652
cc_45 VNB N_VGND_c_642_n 0.0149193f $X=-0.19 $Y=-0.245 $X2=1.17 $Y2=1.665
cc_46 VNB N_VGND_c_643_n 0.0026136f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_VGND_c_644_n 0.0120272f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_VGND_c_645_n 0.0425996f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_VGND_c_646_n 0.0191172f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_VGND_c_647_n 0.0160823f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_VGND_c_648_n 0.0403231f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_VGND_c_649_n 0.017175f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_VGND_c_650_n 0.0151736f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_VGND_c_651_n 0.00446116f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_VGND_c_652_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_VGND_c_653_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_VGND_c_654_n 0.00668318f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_VGND_c_655_n 0.320652f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VPB N_A2_c_104_n 0.0143537f $X=-0.19 $Y=1.66 $X2=1.005 $Y2=1.86
cc_60 VPB N_A2_c_105_n 0.0143554f $X=-0.19 $Y=1.66 $X2=1.455 $Y2=1.86
cc_61 VPB N_A2_c_102_n 0.0047247f $X=-0.19 $Y=1.66 $X2=1.34 $Y2=1.61
cc_62 VPB N_A2_c_103_n 0.0344136f $X=-0.19 $Y=1.66 $X2=1.43 $Y2=1.652
cc_63 VPB N_A1_c_153_n 0.00922335f $X=-0.19 $Y=1.66 $X2=1 $Y2=0.945
cc_64 VPB N_A1_c_161_n 0.0274012f $X=-0.19 $Y=1.66 $X2=1.005 $Y2=2.435
cc_65 VPB N_A1_c_157_n 0.0322356f $X=-0.19 $Y=1.66 $X2=1.455 $Y2=1.86
cc_66 VPB A1 0.00434418f $X=-0.19 $Y=1.66 $X2=1.34 $Y2=1.61
cc_67 VPB N_B1_c_221_n 0.0165277f $X=-0.19 $Y=1.66 $X2=1.005 $Y2=1.86
cc_68 VPB N_B1_c_222_n 0.0175905f $X=-0.19 $Y=1.66 $X2=1.455 $Y2=1.86
cc_69 VPB B1 0.0051867f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_70 VPB N_B1_c_220_n 0.0368644f $X=-0.19 $Y=1.66 $X2=1.455 $Y2=1.652
cc_71 VPB N_A_216_387#_c_281_n 0.0164581f $X=-0.19 $Y=1.66 $X2=1.43 $Y2=0.945
cc_72 VPB N_A_216_387#_c_282_n 0.0156627f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_73 VPB N_A_216_387#_c_283_n 0.0156617f $X=-0.19 $Y=1.66 $X2=1.43 $Y2=1.652
cc_74 VPB N_A_216_387#_c_284_n 0.0176935f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_75 VPB N_A_216_387#_c_277_n 0.00446776f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_76 VPB N_A_216_387#_c_286_n 0.00397148f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_77 VPB N_A_216_387#_c_280_n 0.0355354f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_78 VPB N_VPWR_c_413_n 0.0121909f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_79 VPB N_VPWR_c_414_n 0.0556592f $X=-0.19 $Y=1.66 $X2=1.005 $Y2=1.652
cc_80 VPB N_VPWR_c_415_n 0.0173787f $X=-0.19 $Y=1.66 $X2=1.17 $Y2=1.61
cc_81 VPB N_VPWR_c_416_n 0.0205227f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_82 VPB N_VPWR_c_417_n 0.00900305f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_83 VPB N_VPWR_c_418_n 0.0121909f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_84 VPB N_VPWR_c_419_n 0.0513917f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_85 VPB N_VPWR_c_420_n 0.0216748f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_86 VPB N_VPWR_c_421_n 0.00920679f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_87 VPB N_VPWR_c_422_n 0.039459f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_88 VPB N_VPWR_c_423_n 0.0196495f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_89 VPB N_VPWR_c_424_n 0.0186948f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_90 VPB N_VPWR_c_425_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_91 VPB N_VPWR_c_426_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_92 VPB N_VPWR_c_412_n 0.0881897f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_93 VPB N_A_116_387#_c_482_n 0.00746603f $X=-0.19 $Y=1.66 $X2=1.455 $Y2=2.435
cc_94 VPB N_A_116_387#_c_483_n 0.00332693f $X=-0.19 $Y=1.66 $X2=1.455 $Y2=2.435
cc_95 VPB N_X_c_507_n 0.00257348f $X=-0.19 $Y=1.66 $X2=1.115 $Y2=1.58
cc_96 VPB N_X_c_508_n 0.00283613f $X=-0.19 $Y=1.66 $X2=1.455 $Y2=1.652
cc_97 VPB N_X_c_509_n 0.00224287f $X=-0.19 $Y=1.66 $X2=1.17 $Y2=1.61
cc_98 VPB N_X_c_510_n 0.00257348f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_99 VPB X 0.00977006f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_100 N_A2_M1005_g N_A1_c_152_n 0.00461814f $X=1 $Y=0.945 $X2=-0.19 $Y2=-0.245
cc_101 N_A2_c_102_n N_A1_c_153_n 0.00214824f $X=1.34 $Y=1.61 $X2=0 $Y2=0
cc_102 N_A2_c_103_n N_A1_c_153_n 0.0199616f $X=1.43 $Y=1.652 $X2=0 $Y2=0
cc_103 N_A2_M1005_g N_A1_M1010_g 0.0205891f $X=1 $Y=0.945 $X2=0 $Y2=0
cc_104 N_A2_c_104_n N_A1_c_161_n 0.0194511f $X=1.005 $Y=1.86 $X2=0 $Y2=0
cc_105 N_A2_c_103_n N_A1_c_161_n 0.00387721f $X=1.43 $Y=1.652 $X2=0 $Y2=0
cc_106 N_A2_M1005_g N_A1_c_155_n 0.00894529f $X=1 $Y=0.945 $X2=0 $Y2=0
cc_107 N_A2_M1006_g N_A1_c_155_n 0.00895007f $X=1.43 $Y=0.945 $X2=0 $Y2=0
cc_108 N_A2_c_105_n N_A1_c_157_n 0.0272126f $X=1.455 $Y=1.86 $X2=0 $Y2=0
cc_109 N_A2_c_102_n N_A1_c_157_n 3.92399e-19 $X=1.34 $Y=1.61 $X2=0 $Y2=0
cc_110 N_A2_c_103_n N_A1_c_157_n 0.0216779f $X=1.43 $Y=1.652 $X2=0 $Y2=0
cc_111 N_A2_M1006_g N_A1_M1012_g 0.0222303f $X=1.43 $Y=0.945 $X2=0 $Y2=0
cc_112 N_A2_c_102_n A1 0.0177909f $X=1.34 $Y=1.61 $X2=0 $Y2=0
cc_113 N_A2_c_103_n A1 0.00145483f $X=1.43 $Y=1.652 $X2=0 $Y2=0
cc_114 N_A2_c_105_n N_A_216_387#_c_288_n 0.0125107f $X=1.455 $Y=1.86 $X2=0 $Y2=0
cc_115 N_A2_c_102_n N_A_216_387#_c_288_n 0.00780011f $X=1.34 $Y=1.61 $X2=0 $Y2=0
cc_116 N_A2_c_104_n N_A_216_387#_c_290_n 0.0092516f $X=1.005 $Y=1.86 $X2=0 $Y2=0
cc_117 N_A2_c_105_n N_A_216_387#_c_290_n 0.00881955f $X=1.455 $Y=1.86 $X2=0
+ $Y2=0
cc_118 N_A2_c_102_n N_A_216_387#_c_290_n 0.0232219f $X=1.34 $Y=1.61 $X2=0 $Y2=0
cc_119 N_A2_c_103_n N_A_216_387#_c_290_n 0.00183877f $X=1.43 $Y=1.652 $X2=0
+ $Y2=0
cc_120 N_A2_c_104_n N_VPWR_c_414_n 4.43091e-19 $X=1.005 $Y=1.86 $X2=0 $Y2=0
cc_121 N_A2_c_104_n N_VPWR_c_422_n 9.44495e-19 $X=1.005 $Y=1.86 $X2=0 $Y2=0
cc_122 N_A2_c_105_n N_VPWR_c_422_n 9.44495e-19 $X=1.455 $Y=1.86 $X2=0 $Y2=0
cc_123 N_A2_c_102_n N_A_116_387#_c_484_n 0.00244152f $X=1.34 $Y=1.61 $X2=0 $Y2=0
cc_124 N_A2_c_103_n N_A_116_387#_c_484_n 2.18461e-19 $X=1.43 $Y=1.652 $X2=0
+ $Y2=0
cc_125 N_A2_c_104_n N_A_116_387#_c_482_n 0.0140828f $X=1.005 $Y=1.86 $X2=0 $Y2=0
cc_126 N_A2_c_105_n N_A_116_387#_c_482_n 0.014773f $X=1.455 $Y=1.86 $X2=0 $Y2=0
cc_127 N_A2_M1005_g N_A_27_125#_c_573_n 8.14629e-19 $X=1 $Y=0.945 $X2=0 $Y2=0
cc_128 N_A2_M1005_g N_A_27_125#_c_574_n 0.0125078f $X=1 $Y=0.945 $X2=0 $Y2=0
cc_129 N_A2_c_102_n N_A_27_125#_c_574_n 0.0216324f $X=1.34 $Y=1.61 $X2=0 $Y2=0
cc_130 N_A2_c_103_n N_A_27_125#_c_574_n 6.27125e-19 $X=1.43 $Y=1.652 $X2=0 $Y2=0
cc_131 N_A2_M1006_g N_A_27_125#_c_576_n 0.00735846f $X=1.43 $Y=0.945 $X2=0 $Y2=0
cc_132 N_A2_M1006_g N_A_27_125#_c_577_n 0.0116092f $X=1.43 $Y=0.945 $X2=0 $Y2=0
cc_133 N_A2_c_102_n N_A_27_125#_c_577_n 0.0088782f $X=1.34 $Y=1.61 $X2=0 $Y2=0
cc_134 N_A2_c_103_n N_A_27_125#_c_577_n 0.00121018f $X=1.43 $Y=1.652 $X2=0 $Y2=0
cc_135 N_A2_M1006_g N_A_27_125#_c_578_n 8.55081e-19 $X=1.43 $Y=0.945 $X2=0 $Y2=0
cc_136 N_A2_M1006_g N_A_27_125#_c_582_n 8.39256e-19 $X=1.43 $Y=0.945 $X2=0 $Y2=0
cc_137 N_A2_c_102_n N_A_27_125#_c_582_n 0.0210722f $X=1.34 $Y=1.61 $X2=0 $Y2=0
cc_138 N_A2_c_103_n N_A_27_125#_c_582_n 7.86539e-19 $X=1.43 $Y=1.652 $X2=0 $Y2=0
cc_139 N_A2_M1005_g N_VGND_c_640_n 0.00763474f $X=1 $Y=0.945 $X2=0 $Y2=0
cc_140 N_A2_M1006_g N_VGND_c_640_n 4.4191e-19 $X=1.43 $Y=0.945 $X2=0 $Y2=0
cc_141 N_A2_M1006_g N_VGND_c_641_n 0.00378934f $X=1.43 $Y=0.945 $X2=0 $Y2=0
cc_142 N_A2_M1005_g N_VGND_c_655_n 7.97988e-19 $X=1 $Y=0.945 $X2=0 $Y2=0
cc_143 N_A2_M1006_g N_VGND_c_655_n 9.49986e-19 $X=1.43 $Y=0.945 $X2=0 $Y2=0
cc_144 N_A1_M1012_g N_B1_M1009_g 0.0145764f $X=2.01 $Y=0.945 $X2=0 $Y2=0
cc_145 N_A1_c_157_n N_B1_c_221_n 0.0224802f $X=1.955 $Y=1.86 $X2=0 $Y2=0
cc_146 N_A1_c_157_n B1 2.18718e-19 $X=1.955 $Y=1.86 $X2=0 $Y2=0
cc_147 A1 B1 0.022817f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_148 N_A1_c_157_n N_B1_c_220_n 0.0217423f $X=1.955 $Y=1.86 $X2=0 $Y2=0
cc_149 A1 N_B1_c_220_n 0.00413574f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_150 N_A1_c_157_n N_A_216_387#_c_288_n 0.0163558f $X=1.955 $Y=1.86 $X2=0 $Y2=0
cc_151 A1 N_A_216_387#_c_288_n 0.0322164f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_152 N_A1_c_157_n N_A_216_387#_c_290_n 6.56467e-19 $X=1.955 $Y=1.86 $X2=0
+ $Y2=0
cc_153 N_A1_c_157_n N_A_216_387#_c_286_n 8.62472e-19 $X=1.955 $Y=1.86 $X2=0
+ $Y2=0
cc_154 N_A1_c_161_n N_VPWR_c_414_n 0.0155764f $X=0.505 $Y=1.86 $X2=0 $Y2=0
cc_155 N_A1_c_157_n N_VPWR_c_415_n 0.00715123f $X=1.955 $Y=1.86 $X2=0 $Y2=0
cc_156 N_A1_c_161_n N_VPWR_c_422_n 0.00502391f $X=0.505 $Y=1.86 $X2=0 $Y2=0
cc_157 N_A1_c_157_n N_VPWR_c_422_n 0.00513163f $X=1.955 $Y=1.86 $X2=0 $Y2=0
cc_158 N_A1_c_161_n N_VPWR_c_412_n 0.00487653f $X=0.505 $Y=1.86 $X2=0 $Y2=0
cc_159 N_A1_c_157_n N_VPWR_c_412_n 0.00484068f $X=1.955 $Y=1.86 $X2=0 $Y2=0
cc_160 N_A1_c_157_n N_A_116_387#_c_482_n 0.00361932f $X=1.955 $Y=1.86 $X2=0
+ $Y2=0
cc_161 N_A1_c_161_n N_A_116_387#_c_483_n 0.0013728f $X=0.505 $Y=1.86 $X2=0 $Y2=0
cc_162 N_A1_c_157_n N_A_116_387#_c_490_n 0.00662701f $X=1.955 $Y=1.86 $X2=0
+ $Y2=0
cc_163 N_A1_M1010_g N_A_27_125#_c_573_n 0.00756074f $X=0.495 $Y=0.945 $X2=0
+ $Y2=0
cc_164 N_A1_c_152_n N_A_27_125#_c_574_n 0.00113437f $X=0.505 $Y=1.43 $X2=0 $Y2=0
cc_165 N_A1_M1010_g N_A_27_125#_c_574_n 0.0152942f $X=0.495 $Y=0.945 $X2=0 $Y2=0
cc_166 N_A1_M1010_g N_A_27_125#_c_575_n 0.00163942f $X=0.495 $Y=0.945 $X2=0
+ $Y2=0
cc_167 N_A1_c_155_n N_A_27_125#_c_576_n 0.00449567f $X=1.935 $Y=0.18 $X2=0 $Y2=0
cc_168 N_A1_M1012_g N_A_27_125#_c_576_n 8.40186e-19 $X=2.01 $Y=0.945 $X2=0 $Y2=0
cc_169 N_A1_c_157_n N_A_27_125#_c_577_n 0.00430368f $X=1.955 $Y=1.86 $X2=0 $Y2=0
cc_170 N_A1_M1012_g N_A_27_125#_c_577_n 0.0126915f $X=2.01 $Y=0.945 $X2=0 $Y2=0
cc_171 A1 N_A_27_125#_c_577_n 0.0380956f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_172 N_A1_M1012_g N_A_27_125#_c_578_n 0.0113517f $X=2.01 $Y=0.945 $X2=0 $Y2=0
cc_173 N_A1_M1012_g N_A_27_125#_c_580_n 0.00615508f $X=2.01 $Y=0.945 $X2=0 $Y2=0
cc_174 N_A1_M1010_g N_VGND_c_640_n 0.0151444f $X=0.495 $Y=0.945 $X2=0 $Y2=0
cc_175 N_A1_c_155_n N_VGND_c_640_n 0.0235422f $X=1.935 $Y=0.18 $X2=0 $Y2=0
cc_176 N_A1_c_155_n N_VGND_c_641_n 0.0235859f $X=1.935 $Y=0.18 $X2=0 $Y2=0
cc_177 N_A1_M1012_g N_VGND_c_641_n 0.00876868f $X=2.01 $Y=0.945 $X2=0 $Y2=0
cc_178 N_A1_c_156_n N_VGND_c_646_n 0.00730708f $X=0.57 $Y=0.18 $X2=0 $Y2=0
cc_179 N_A1_c_155_n N_VGND_c_647_n 0.0187698f $X=1.935 $Y=0.18 $X2=0 $Y2=0
cc_180 N_A1_c_155_n N_VGND_c_648_n 0.00719493f $X=1.935 $Y=0.18 $X2=0 $Y2=0
cc_181 N_A1_c_155_n N_VGND_c_655_n 0.0361523f $X=1.935 $Y=0.18 $X2=0 $Y2=0
cc_182 N_A1_c_156_n N_VGND_c_655_n 0.0101958f $X=0.57 $Y=0.18 $X2=0 $Y2=0
cc_183 N_B1_c_222_n N_A_216_387#_c_281_n 0.0147592f $X=3.025 $Y=1.86 $X2=0 $Y2=0
cc_184 N_B1_c_220_n N_A_216_387#_c_281_n 0.00122205f $X=2.95 $Y=1.61 $X2=0 $Y2=0
cc_185 N_B1_c_221_n N_A_216_387#_c_288_n 0.0139083f $X=2.495 $Y=1.86 $X2=0 $Y2=0
cc_186 B1 N_A_216_387#_c_288_n 0.0083868f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_187 N_B1_M1014_g N_A_216_387#_c_274_n 0.011831f $X=2.87 $Y=0.945 $X2=0 $Y2=0
cc_188 N_B1_M1014_g N_A_216_387#_c_275_n 0.012382f $X=2.87 $Y=0.945 $X2=0 $Y2=0
cc_189 B1 N_A_216_387#_c_275_n 0.0306534f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_190 N_B1_c_220_n N_A_216_387#_c_275_n 0.00480134f $X=2.95 $Y=1.61 $X2=0 $Y2=0
cc_191 N_B1_M1009_g N_A_216_387#_c_276_n 0.00229365f $X=2.44 $Y=0.945 $X2=0
+ $Y2=0
cc_192 N_B1_M1014_g N_A_216_387#_c_276_n 0.00147096f $X=2.87 $Y=0.945 $X2=0
+ $Y2=0
cc_193 B1 N_A_216_387#_c_276_n 0.0206608f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_194 N_B1_c_220_n N_A_216_387#_c_276_n 0.00253619f $X=2.95 $Y=1.61 $X2=0 $Y2=0
cc_195 N_B1_c_222_n N_A_216_387#_c_310_n 0.0165967f $X=3.025 $Y=1.86 $X2=0 $Y2=0
cc_196 B1 N_A_216_387#_c_310_n 0.020891f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_197 N_B1_c_222_n N_A_216_387#_c_277_n 0.00176786f $X=3.025 $Y=1.86 $X2=0
+ $Y2=0
cc_198 B1 N_A_216_387#_c_277_n 0.0193018f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_199 N_B1_c_220_n N_A_216_387#_c_277_n 0.00229245f $X=2.95 $Y=1.61 $X2=0 $Y2=0
cc_200 N_B1_c_221_n N_A_216_387#_c_286_n 0.00947928f $X=2.495 $Y=1.86 $X2=0
+ $Y2=0
cc_201 N_B1_c_222_n N_A_216_387#_c_286_n 0.00378026f $X=3.025 $Y=1.86 $X2=0
+ $Y2=0
cc_202 B1 N_A_216_387#_c_286_n 0.0253731f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_203 N_B1_c_220_n N_A_216_387#_c_286_n 0.00227154f $X=2.95 $Y=1.61 $X2=0 $Y2=0
cc_204 N_B1_M1014_g N_A_216_387#_c_279_n 0.0021086f $X=2.87 $Y=0.945 $X2=0 $Y2=0
cc_205 B1 N_A_216_387#_c_279_n 0.00318495f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_206 N_B1_c_220_n N_A_216_387#_c_279_n 0.00192995f $X=2.95 $Y=1.61 $X2=0 $Y2=0
cc_207 N_B1_M1014_g N_A_216_387#_c_280_n 0.0043112f $X=2.87 $Y=0.945 $X2=0 $Y2=0
cc_208 N_B1_c_220_n N_A_216_387#_c_280_n 0.00706187f $X=2.95 $Y=1.61 $X2=0 $Y2=0
cc_209 N_B1_c_221_n N_VPWR_c_415_n 0.00418617f $X=2.495 $Y=1.86 $X2=0 $Y2=0
cc_210 N_B1_c_222_n N_VPWR_c_416_n 0.00774357f $X=3.025 $Y=1.86 $X2=0 $Y2=0
cc_211 N_B1_c_221_n N_VPWR_c_420_n 0.00451198f $X=2.495 $Y=1.86 $X2=0 $Y2=0
cc_212 N_B1_c_222_n N_VPWR_c_420_n 0.00454183f $X=3.025 $Y=1.86 $X2=0 $Y2=0
cc_213 N_B1_c_221_n N_VPWR_c_412_n 0.00489211f $X=2.495 $Y=1.86 $X2=0 $Y2=0
cc_214 N_B1_c_222_n N_VPWR_c_412_n 0.00489211f $X=3.025 $Y=1.86 $X2=0 $Y2=0
cc_215 N_B1_M1009_g N_A_27_125#_c_577_n 0.00248344f $X=2.44 $Y=0.945 $X2=0 $Y2=0
cc_216 N_B1_M1009_g N_A_27_125#_c_578_n 0.00918561f $X=2.44 $Y=0.945 $X2=0 $Y2=0
cc_217 N_B1_M1014_g N_A_27_125#_c_578_n 4.92416e-19 $X=2.87 $Y=0.945 $X2=0 $Y2=0
cc_218 N_B1_M1009_g N_A_27_125#_c_579_n 0.00582977f $X=2.44 $Y=0.945 $X2=0 $Y2=0
cc_219 N_B1_M1014_g N_A_27_125#_c_579_n 0.00661564f $X=2.87 $Y=0.945 $X2=0 $Y2=0
cc_220 N_B1_M1014_g N_A_27_125#_c_581_n 0.0108881f $X=2.87 $Y=0.945 $X2=0 $Y2=0
cc_221 N_B1_M1009_g N_VGND_c_648_n 2.28708e-19 $X=2.44 $Y=0.945 $X2=0 $Y2=0
cc_222 N_A_216_387#_c_288_n N_VPWR_M1019_d 0.00698293f $X=2.565 $Y=2.035 $X2=0
+ $Y2=0
cc_223 N_A_216_387#_c_310_n N_VPWR_M1004_d 0.0130167f $X=3.405 $Y=2.035 $X2=0
+ $Y2=0
cc_224 N_A_216_387#_c_277_n N_VPWR_M1004_d 0.00217152f $X=3.49 $Y=1.95 $X2=0
+ $Y2=0
cc_225 N_A_216_387#_c_288_n N_VPWR_c_415_n 0.022455f $X=2.565 $Y=2.035 $X2=0
+ $Y2=0
cc_226 N_A_216_387#_c_286_n N_VPWR_c_415_n 0.0197393f $X=2.73 $Y=2.115 $X2=0
+ $Y2=0
cc_227 N_A_216_387#_c_281_n N_VPWR_c_416_n 0.0134661f $X=3.755 $Y=1.765 $X2=0
+ $Y2=0
cc_228 N_A_216_387#_c_310_n N_VPWR_c_416_n 0.0338933f $X=3.405 $Y=2.035 $X2=0
+ $Y2=0
cc_229 N_A_216_387#_c_286_n N_VPWR_c_416_n 0.00127808f $X=2.73 $Y=2.115 $X2=0
+ $Y2=0
cc_230 N_A_216_387#_c_282_n N_VPWR_c_417_n 0.00874363f $X=4.205 $Y=1.765 $X2=0
+ $Y2=0
cc_231 N_A_216_387#_c_283_n N_VPWR_c_417_n 0.00735548f $X=4.755 $Y=1.765 $X2=0
+ $Y2=0
cc_232 N_A_216_387#_c_284_n N_VPWR_c_419_n 0.0235387f $X=5.205 $Y=1.765 $X2=0
+ $Y2=0
cc_233 N_A_216_387#_c_286_n N_VPWR_c_420_n 0.0082974f $X=2.73 $Y=2.115 $X2=0
+ $Y2=0
cc_234 N_A_216_387#_c_281_n N_VPWR_c_423_n 0.00445602f $X=3.755 $Y=1.765 $X2=0
+ $Y2=0
cc_235 N_A_216_387#_c_282_n N_VPWR_c_423_n 0.00445602f $X=4.205 $Y=1.765 $X2=0
+ $Y2=0
cc_236 N_A_216_387#_c_283_n N_VPWR_c_424_n 0.00445602f $X=4.755 $Y=1.765 $X2=0
+ $Y2=0
cc_237 N_A_216_387#_c_284_n N_VPWR_c_424_n 0.00445602f $X=5.205 $Y=1.765 $X2=0
+ $Y2=0
cc_238 N_A_216_387#_c_281_n N_VPWR_c_412_n 0.00862391f $X=3.755 $Y=1.765 $X2=0
+ $Y2=0
cc_239 N_A_216_387#_c_282_n N_VPWR_c_412_n 0.00857797f $X=4.205 $Y=1.765 $X2=0
+ $Y2=0
cc_240 N_A_216_387#_c_283_n N_VPWR_c_412_n 0.00857797f $X=4.755 $Y=1.765 $X2=0
+ $Y2=0
cc_241 N_A_216_387#_c_284_n N_VPWR_c_412_n 0.00860566f $X=5.205 $Y=1.765 $X2=0
+ $Y2=0
cc_242 N_A_216_387#_c_286_n N_VPWR_c_412_n 0.0107001f $X=2.73 $Y=2.115 $X2=0
+ $Y2=0
cc_243 N_A_216_387#_c_288_n N_A_116_387#_M1018_s 0.00715037f $X=2.565 $Y=2.035
+ $X2=0 $Y2=0
cc_244 N_A_216_387#_c_290_n N_A_116_387#_c_484_n 0.0533059f $X=1.23 $Y=2.115
+ $X2=0 $Y2=0
cc_245 N_A_216_387#_M1015_d N_A_116_387#_c_482_n 0.00197722f $X=1.08 $Y=1.935
+ $X2=0 $Y2=0
cc_246 N_A_216_387#_c_290_n N_A_116_387#_c_482_n 0.0160777f $X=1.23 $Y=2.115
+ $X2=0 $Y2=0
cc_247 N_A_216_387#_c_288_n N_A_116_387#_c_490_n 0.0202249f $X=2.565 $Y=2.035
+ $X2=0 $Y2=0
cc_248 N_A_216_387#_c_281_n N_X_c_507_n 0.0186729f $X=3.755 $Y=1.765 $X2=0 $Y2=0
cc_249 N_A_216_387#_c_282_n N_X_c_507_n 0.0131597f $X=4.205 $Y=1.765 $X2=0 $Y2=0
cc_250 N_A_216_387#_c_283_n N_X_c_507_n 7.1037e-19 $X=4.755 $Y=1.765 $X2=0 $Y2=0
cc_251 N_A_216_387#_c_310_n N_X_c_507_n 0.0107657f $X=3.405 $Y=2.035 $X2=0 $Y2=0
cc_252 N_A_216_387#_c_277_n N_X_c_507_n 0.00334171f $X=3.49 $Y=1.95 $X2=0 $Y2=0
cc_253 N_A_216_387#_c_270_n N_X_c_517_n 0.00219545f $X=3.94 $Y=1.22 $X2=0 $Y2=0
cc_254 N_A_216_387#_c_278_n N_X_c_517_n 0.0190038f $X=4.63 $Y=1.385 $X2=0 $Y2=0
cc_255 N_A_216_387#_c_280_n N_X_c_517_n 6.90776e-19 $X=5.205 $Y=1.492 $X2=0
+ $Y2=0
cc_256 N_A_216_387#_c_270_n N_X_c_503_n 0.00638907f $X=3.94 $Y=1.22 $X2=0 $Y2=0
cc_257 N_A_216_387#_c_271_n N_X_c_503_n 4.40427e-19 $X=4.37 $Y=1.22 $X2=0 $Y2=0
cc_258 N_A_216_387#_c_282_n N_X_c_508_n 0.00941072f $X=4.205 $Y=1.765 $X2=0
+ $Y2=0
cc_259 N_A_216_387#_c_283_n N_X_c_508_n 0.00941072f $X=4.755 $Y=1.765 $X2=0
+ $Y2=0
cc_260 N_A_216_387#_c_278_n N_X_c_508_n 0.0482544f $X=4.63 $Y=1.385 $X2=0 $Y2=0
cc_261 N_A_216_387#_c_280_n N_X_c_508_n 0.0125578f $X=5.205 $Y=1.492 $X2=0 $Y2=0
cc_262 N_A_216_387#_c_281_n N_X_c_509_n 0.0023714f $X=3.755 $Y=1.765 $X2=0 $Y2=0
cc_263 N_A_216_387#_c_282_n N_X_c_509_n 0.00109449f $X=4.205 $Y=1.765 $X2=0
+ $Y2=0
cc_264 N_A_216_387#_c_277_n N_X_c_509_n 0.0103664f $X=3.49 $Y=1.95 $X2=0 $Y2=0
cc_265 N_A_216_387#_c_278_n N_X_c_509_n 0.0278089f $X=4.63 $Y=1.385 $X2=0 $Y2=0
cc_266 N_A_216_387#_c_280_n N_X_c_509_n 0.00584196f $X=5.205 $Y=1.492 $X2=0
+ $Y2=0
cc_267 N_A_216_387#_c_271_n N_X_c_531_n 0.0097547f $X=4.37 $Y=1.22 $X2=0 $Y2=0
cc_268 N_A_216_387#_c_272_n N_X_c_531_n 0.0132906f $X=4.835 $Y=1.22 $X2=0 $Y2=0
cc_269 N_A_216_387#_c_278_n N_X_c_531_n 0.0363197f $X=4.63 $Y=1.385 $X2=0 $Y2=0
cc_270 N_A_216_387#_c_280_n N_X_c_531_n 8.3386e-19 $X=5.205 $Y=1.492 $X2=0 $Y2=0
cc_271 N_A_216_387#_c_282_n N_X_c_510_n 7.1037e-19 $X=4.205 $Y=1.765 $X2=0 $Y2=0
cc_272 N_A_216_387#_c_283_n N_X_c_510_n 0.0131597f $X=4.755 $Y=1.765 $X2=0 $Y2=0
cc_273 N_A_216_387#_c_284_n N_X_c_510_n 0.0137894f $X=5.205 $Y=1.765 $X2=0 $Y2=0
cc_274 N_A_216_387#_c_272_n N_X_c_504_n 3.92313e-19 $X=4.835 $Y=1.22 $X2=0 $Y2=0
cc_275 N_A_216_387#_c_273_n N_X_c_504_n 3.92313e-19 $X=5.265 $Y=1.22 $X2=0 $Y2=0
cc_276 N_A_216_387#_c_272_n N_X_c_505_n 0.00185803f $X=4.835 $Y=1.22 $X2=0 $Y2=0
cc_277 N_A_216_387#_c_273_n N_X_c_505_n 0.00228347f $X=5.265 $Y=1.22 $X2=0 $Y2=0
cc_278 N_A_216_387#_c_278_n N_X_c_505_n 0.0285354f $X=4.63 $Y=1.385 $X2=0 $Y2=0
cc_279 N_A_216_387#_c_280_n N_X_c_505_n 0.0249419f $X=5.205 $Y=1.492 $X2=0 $Y2=0
cc_280 N_A_216_387#_c_283_n N_X_c_544_n 0.00109449f $X=4.755 $Y=1.765 $X2=0
+ $Y2=0
cc_281 N_A_216_387#_c_284_n N_X_c_544_n 0.00603924f $X=5.205 $Y=1.765 $X2=0
+ $Y2=0
cc_282 N_A_216_387#_c_280_n N_X_c_544_n 0.0245632f $X=5.205 $Y=1.492 $X2=0 $Y2=0
cc_283 N_A_216_387#_c_284_n X 0.00657385f $X=5.205 $Y=1.765 $X2=0 $Y2=0
cc_284 N_A_216_387#_c_280_n X 0.0160575f $X=5.205 $Y=1.492 $X2=0 $Y2=0
cc_285 N_A_216_387#_c_275_n N_A_27_125#_M1014_d 0.00396376f $X=3.405 $Y=1.26
+ $X2=0 $Y2=0
cc_286 N_A_216_387#_c_288_n N_A_27_125#_c_577_n 0.0101635f $X=2.565 $Y=2.035
+ $X2=0 $Y2=0
cc_287 N_A_216_387#_c_276_n N_A_27_125#_c_577_n 0.00444516f $X=2.82 $Y=1.26
+ $X2=0 $Y2=0
cc_288 N_A_216_387#_c_274_n N_A_27_125#_c_578_n 0.0186128f $X=2.655 $Y=0.77
+ $X2=0 $Y2=0
cc_289 N_A_216_387#_c_274_n N_A_27_125#_c_579_n 0.0195392f $X=2.655 $Y=0.77
+ $X2=0 $Y2=0
cc_290 N_A_216_387#_c_274_n N_A_27_125#_c_581_n 0.0144986f $X=2.655 $Y=0.77
+ $X2=0 $Y2=0
cc_291 N_A_216_387#_c_275_n N_A_27_125#_c_581_n 0.0266632f $X=3.405 $Y=1.26
+ $X2=0 $Y2=0
cc_292 N_A_216_387#_c_270_n N_VGND_c_642_n 0.00340257f $X=3.94 $Y=1.22 $X2=0
+ $Y2=0
cc_293 N_A_216_387#_c_278_n N_VGND_c_642_n 0.0203976f $X=4.63 $Y=1.385 $X2=0
+ $Y2=0
cc_294 N_A_216_387#_c_279_n N_VGND_c_642_n 0.00131156f $X=3.49 $Y=1.362 $X2=0
+ $Y2=0
cc_295 N_A_216_387#_c_280_n N_VGND_c_642_n 0.00174316f $X=5.205 $Y=1.492 $X2=0
+ $Y2=0
cc_296 N_A_216_387#_c_270_n N_VGND_c_643_n 3.93623e-19 $X=3.94 $Y=1.22 $X2=0
+ $Y2=0
cc_297 N_A_216_387#_c_271_n N_VGND_c_643_n 0.00765879f $X=4.37 $Y=1.22 $X2=0
+ $Y2=0
cc_298 N_A_216_387#_c_272_n N_VGND_c_643_n 0.00768892f $X=4.835 $Y=1.22 $X2=0
+ $Y2=0
cc_299 N_A_216_387#_c_273_n N_VGND_c_643_n 4.1905e-19 $X=5.265 $Y=1.22 $X2=0
+ $Y2=0
cc_300 N_A_216_387#_c_272_n N_VGND_c_645_n 4.70441e-19 $X=4.835 $Y=1.22 $X2=0
+ $Y2=0
cc_301 N_A_216_387#_c_273_n N_VGND_c_645_n 0.0150633f $X=5.265 $Y=1.22 $X2=0
+ $Y2=0
cc_302 N_A_216_387#_c_270_n N_VGND_c_649_n 0.00433834f $X=3.94 $Y=1.22 $X2=0
+ $Y2=0
cc_303 N_A_216_387#_c_271_n N_VGND_c_649_n 0.00383152f $X=4.37 $Y=1.22 $X2=0
+ $Y2=0
cc_304 N_A_216_387#_c_272_n N_VGND_c_650_n 0.00383152f $X=4.835 $Y=1.22 $X2=0
+ $Y2=0
cc_305 N_A_216_387#_c_273_n N_VGND_c_650_n 0.00383152f $X=5.265 $Y=1.22 $X2=0
+ $Y2=0
cc_306 N_A_216_387#_c_270_n N_VGND_c_655_n 0.00824977f $X=3.94 $Y=1.22 $X2=0
+ $Y2=0
cc_307 N_A_216_387#_c_271_n N_VGND_c_655_n 0.00382921f $X=4.37 $Y=1.22 $X2=0
+ $Y2=0
cc_308 N_A_216_387#_c_272_n N_VGND_c_655_n 0.00382921f $X=4.835 $Y=1.22 $X2=0
+ $Y2=0
cc_309 N_A_216_387#_c_273_n N_VGND_c_655_n 0.0075754f $X=5.265 $Y=1.22 $X2=0
+ $Y2=0
cc_310 N_VPWR_c_415_n N_A_116_387#_c_482_n 0.013014f $X=2.23 $Y=2.455 $X2=0
+ $Y2=0
cc_311 N_VPWR_c_422_n N_A_116_387#_c_482_n 0.0686911f $X=2.065 $Y=3.33 $X2=0
+ $Y2=0
cc_312 N_VPWR_c_412_n N_A_116_387#_c_482_n 0.0391401f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_313 N_VPWR_c_414_n N_A_116_387#_c_483_n 0.0129306f $X=0.28 $Y=2.08 $X2=0
+ $Y2=0
cc_314 N_VPWR_c_422_n N_A_116_387#_c_483_n 0.0179217f $X=2.065 $Y=3.33 $X2=0
+ $Y2=0
cc_315 N_VPWR_c_412_n N_A_116_387#_c_483_n 0.00971942f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_316 N_VPWR_c_416_n N_X_c_507_n 0.0479989f $X=3.36 $Y=2.465 $X2=0 $Y2=0
cc_317 N_VPWR_c_417_n N_X_c_507_n 0.0353111f $X=4.48 $Y=2.145 $X2=0 $Y2=0
cc_318 N_VPWR_c_423_n N_X_c_507_n 0.014552f $X=4.315 $Y=3.33 $X2=0 $Y2=0
cc_319 N_VPWR_c_412_n N_X_c_507_n 0.0119791f $X=5.52 $Y=3.33 $X2=0 $Y2=0
cc_320 N_VPWR_M1011_d N_X_c_508_n 0.00306736f $X=4.28 $Y=1.84 $X2=0 $Y2=0
cc_321 N_VPWR_c_417_n N_X_c_508_n 0.0232685f $X=4.48 $Y=2.145 $X2=0 $Y2=0
cc_322 N_VPWR_c_417_n N_X_c_510_n 0.0353111f $X=4.48 $Y=2.145 $X2=0 $Y2=0
cc_323 N_VPWR_c_419_n N_X_c_510_n 0.0394385f $X=5.48 $Y=2.115 $X2=0 $Y2=0
cc_324 N_VPWR_c_424_n N_X_c_510_n 0.014552f $X=5.315 $Y=3.33 $X2=0 $Y2=0
cc_325 N_VPWR_c_412_n N_X_c_510_n 0.0119791f $X=5.52 $Y=3.33 $X2=0 $Y2=0
cc_326 N_VPWR_c_419_n X 0.0260199f $X=5.48 $Y=2.115 $X2=0 $Y2=0
cc_327 N_VPWR_c_414_n N_A_27_125#_c_575_n 0.0120871f $X=0.28 $Y=2.08 $X2=0 $Y2=0
cc_328 N_A_116_387#_c_484_n N_A_27_125#_c_574_n 0.00631305f $X=0.78 $Y=2.115
+ $X2=0 $Y2=0
cc_329 N_X_c_531_n N_VGND_M1002_d 0.00395842f $X=4.965 $Y=0.92 $X2=0 $Y2=0
cc_330 N_X_c_503_n N_VGND_c_642_n 0.0188059f $X=4.155 $Y=0.495 $X2=0 $Y2=0
cc_331 N_X_c_503_n N_VGND_c_643_n 0.0136878f $X=4.155 $Y=0.495 $X2=0 $Y2=0
cc_332 N_X_c_531_n N_VGND_c_643_n 0.0194786f $X=4.965 $Y=0.92 $X2=0 $Y2=0
cc_333 N_X_c_504_n N_VGND_c_643_n 0.0121521f $X=5.05 $Y=0.515 $X2=0 $Y2=0
cc_334 N_X_c_504_n N_VGND_c_645_n 0.0180696f $X=5.05 $Y=0.515 $X2=0 $Y2=0
cc_335 N_X_c_505_n N_VGND_c_645_n 0.00516673f $X=5.05 $Y=1.55 $X2=0 $Y2=0
cc_336 X N_VGND_c_645_n 0.0145768f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_337 N_X_c_503_n N_VGND_c_649_n 0.0119488f $X=4.155 $Y=0.495 $X2=0 $Y2=0
cc_338 N_X_c_504_n N_VGND_c_650_n 0.00749631f $X=5.05 $Y=0.515 $X2=0 $Y2=0
cc_339 N_X_c_503_n N_VGND_c_655_n 0.00915121f $X=4.155 $Y=0.495 $X2=0 $Y2=0
cc_340 N_X_c_531_n N_VGND_c_655_n 0.0118272f $X=4.965 $Y=0.92 $X2=0 $Y2=0
cc_341 N_X_c_504_n N_VGND_c_655_n 0.0062048f $X=5.05 $Y=0.515 $X2=0 $Y2=0
cc_342 N_A_27_125#_c_574_n N_VGND_M1010_d 0.00256188f $X=1.13 $Y=1.19 $X2=-0.19
+ $Y2=-0.245
cc_343 N_A_27_125#_c_577_n N_VGND_M1006_s 0.00397519f $X=2.06 $Y=1.19 $X2=0
+ $Y2=0
cc_344 N_A_27_125#_c_573_n N_VGND_c_640_n 0.0131747f $X=0.28 $Y=0.77 $X2=0 $Y2=0
cc_345 N_A_27_125#_c_574_n N_VGND_c_640_n 0.0213935f $X=1.13 $Y=1.19 $X2=0 $Y2=0
cc_346 N_A_27_125#_c_576_n N_VGND_c_640_n 0.0125829f $X=1.215 $Y=0.77 $X2=0
+ $Y2=0
cc_347 N_A_27_125#_c_576_n N_VGND_c_641_n 0.0120942f $X=1.215 $Y=0.77 $X2=0
+ $Y2=0
cc_348 N_A_27_125#_c_577_n N_VGND_c_641_n 0.0257093f $X=2.06 $Y=1.19 $X2=0 $Y2=0
cc_349 N_A_27_125#_c_578_n N_VGND_c_641_n 0.0265871f $X=2.225 $Y=0.77 $X2=0
+ $Y2=0
cc_350 N_A_27_125#_c_580_n N_VGND_c_641_n 0.0142636f $X=2.39 $Y=0.35 $X2=0 $Y2=0
cc_351 N_A_27_125#_c_579_n N_VGND_c_642_n 0.0119252f $X=3 $Y=0.35 $X2=0 $Y2=0
cc_352 N_A_27_125#_c_581_n N_VGND_c_642_n 0.0376042f $X=3.165 $Y=0.805 $X2=0
+ $Y2=0
cc_353 N_A_27_125#_c_573_n N_VGND_c_646_n 0.00702137f $X=0.28 $Y=0.77 $X2=0
+ $Y2=0
cc_354 N_A_27_125#_c_576_n N_VGND_c_647_n 0.00528099f $X=1.215 $Y=0.77 $X2=0
+ $Y2=0
cc_355 N_A_27_125#_c_579_n N_VGND_c_648_n 0.0591825f $X=3 $Y=0.35 $X2=0 $Y2=0
cc_356 N_A_27_125#_c_580_n N_VGND_c_648_n 0.0221635f $X=2.39 $Y=0.35 $X2=0 $Y2=0
cc_357 N_A_27_125#_c_573_n N_VGND_c_655_n 0.0100521f $X=0.28 $Y=0.77 $X2=0 $Y2=0
cc_358 N_A_27_125#_c_576_n N_VGND_c_655_n 0.00668051f $X=1.215 $Y=0.77 $X2=0
+ $Y2=0
cc_359 N_A_27_125#_c_579_n N_VGND_c_655_n 0.035558f $X=3 $Y=0.35 $X2=0 $Y2=0
cc_360 N_A_27_125#_c_580_n N_VGND_c_655_n 0.0126536f $X=2.39 $Y=0.35 $X2=0 $Y2=0
