* File: sky130_fd_sc_hs__sdfxbp_1.spice
* Created: Thu Aug 27 21:09:51 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hs__sdfxbp_1.pex.spice"
.subckt sky130_fd_sc_hs__sdfxbp_1  VNB VPB SCE D SCD CLK VPWR Q Q_N VGND
* 
* VGND	VGND
* Q_N	Q_N
* Q	Q
* VPWR	VPWR
* CLK	CLK
* SCD	SCD
* D	D
* SCE	SCE
* VPB	VPB
* VNB	VNB
MM1028 N_VGND_M1028_d N_SCE_M1028_g N_A_31_74#_M1028_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.0735 AS=0.1197 PD=0.77 PS=1.41 NRD=19.992 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75002.7 A=0.063 P=1.14 MULT=1
MM1010 A_218_74# N_A_31_74#_M1010_g N_VGND_M1028_d VNB NLOWVT L=0.15 W=0.42
+ AD=0.0504 AS=0.0735 PD=0.66 PS=0.77 NRD=18.564 NRS=0 M=1 R=2.8 SA=75000.7
+ SB=75002.2 A=0.063 P=1.14 MULT=1
MM1011 N_A_296_74#_M1011_d N_D_M1011_g A_218_74# VNB NLOWVT L=0.15 W=0.42
+ AD=0.1134 AS=0.0504 PD=0.96 PS=0.66 NRD=37.14 NRS=18.564 M=1 R=2.8 SA=75001.1
+ SB=75001.8 A=0.063 P=1.14 MULT=1
MM1003 A_434_74# N_SCE_M1003_g N_A_296_74#_M1011_d VNB NLOWVT L=0.15 W=0.42
+ AD=0.0504 AS=0.1134 PD=0.66 PS=0.96 NRD=18.564 NRS=37.14 M=1 R=2.8 SA=75001.8
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1032 N_VGND_M1032_d N_SCD_M1032_g A_434_74# VNB NLOWVT L=0.15 W=0.42
+ AD=0.0821897 AS=0.0504 PD=0.78931 PS=0.66 NRD=11.424 NRS=18.564 M=1 R=2.8
+ SA=75002.2 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1027 N_A_612_74#_M1027_d N_CLK_M1027_g N_VGND_M1032_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.14481 PD=2.05 PS=1.39069 NRD=0 NRS=4.86 M=1 R=4.93333
+ SA=75001.6 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1017 N_A_828_74#_M1017_d N_A_612_74#_M1017_g N_VGND_M1017_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1998 AS=0.2805 PD=2.02 PS=2.25 NRD=0 NRS=13.776 M=1 R=4.93333
+ SA=75000.3 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1035 N_A_1021_100#_M1035_d N_A_612_74#_M1035_g N_A_296_74#_M1035_s VNB NLOWVT
+ L=0.15 W=0.42 AD=0.1113 AS=0.1155 PD=0.95 PS=1.39 NRD=71.424 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75004 A=0.063 P=1.14 MULT=1
MM1009 A_1157_100# N_A_828_74#_M1009_g N_A_1021_100#_M1035_d VNB NLOWVT L=0.15
+ W=0.42 AD=0.0966 AS=0.1113 PD=0.88 PS=0.95 NRD=49.992 NRS=0 M=1 R=2.8
+ SA=75000.9 SB=75003.4 A=0.063 P=1.14 MULT=1
MM1020 N_VGND_M1020_d N_A_1243_398#_M1020_g A_1157_100# VNB NLOWVT L=0.15 W=0.42
+ AD=0.172849 AS=0.0966 PD=1.19072 PS=0.88 NRD=101.868 NRS=49.992 M=1 R=2.8
+ SA=75001.5 SB=75002.8 A=0.063 P=1.14 MULT=1
MM1015 N_A_1243_398#_M1015_d N_A_1021_100#_M1015_g N_VGND_M1020_d VNB NLOWVT
+ L=0.15 W=0.55 AD=0.078375 AS=0.226351 PD=0.835 PS=1.55928 NRD=1.08 NRS=72 M=1
+ R=3.66667 SA=75001.9 SB=75002.1 A=0.0825 P=1.4 MULT=1
MM1013 N_A_1529_74#_M1013_d N_A_828_74#_M1013_g N_A_1243_398#_M1015_d VNB NLOWVT
+ L=0.15 W=0.55 AD=0.163696 AS=0.078375 PD=1.31546 PS=0.835 NRD=72 NRS=0 M=1
+ R=3.66667 SA=75002.3 SB=75001.6 A=0.0825 P=1.4 MULT=1
MM1021 A_1681_74# N_A_612_74#_M1021_g N_A_1529_74#_M1013_d VNB NLOWVT L=0.15
+ W=0.42 AD=0.0441 AS=0.125004 PD=0.63 PS=1.00454 NRD=14.28 NRS=0 M=1 R=2.8
+ SA=75002.9 SB=75001.3 A=0.063 P=1.14 MULT=1
MM1024 N_VGND_M1024_d N_A_1723_48#_M1024_g A_1681_74# VNB NLOWVT L=0.15 W=0.42
+ AD=0.128793 AS=0.0441 PD=1.0132 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75003.3
+ SB=75001 A=0.063 P=1.14 MULT=1
MM1001 N_A_1723_48#_M1001_d N_A_1529_74#_M1001_g N_VGND_M1024_d VNB NLOWVT
+ L=0.15 W=0.55 AD=0.15675 AS=0.168657 PD=1.67 PS=1.3268 NRD=0 NRS=0 M=1
+ R=3.66667 SA=75003.2 SB=75000.2 A=0.0825 P=1.4 MULT=1
MM1016 N_Q_M1016_d N_A_1723_48#_M1016_g N_VGND_M1016_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.2109 PD=2.05 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1004 N_VGND_M1004_d N_A_1723_48#_M1004_g N_A_2216_94#_M1004_s VNB NLOWVT
+ L=0.15 W=0.64 AD=0.132081 AS=0.1824 PD=1.05275 PS=1.85 NRD=11.244 NRS=0 M=1
+ R=4.26667 SA=75000.2 SB=75000.8 A=0.096 P=1.58 MULT=1
MM1031 N_Q_N_M1031_d N_A_2216_94#_M1031_g N_VGND_M1004_d VNB NLOWVT L=0.15
+ W=0.74 AD=0.2109 AS=0.152719 PD=2.05 PS=1.21725 NRD=0 NRS=9.324 M=1 R=4.93333
+ SA=75000.7 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1033 N_VPWR_M1033_d N_SCE_M1033_g N_A_31_74#_M1033_s VPB PSHORT L=0.15 W=0.64
+ AD=0.112 AS=0.1888 PD=0.99 PS=1.87 NRD=18.4589 NRS=3.0732 M=1 R=4.26667
+ SA=75000.2 SB=75002.8 A=0.096 P=1.58 MULT=1
MM1034 A_233_464# N_SCE_M1034_g N_VPWR_M1033_d VPB PSHORT L=0.15 W=0.64
+ AD=0.0864 AS=0.112 PD=0.91 PS=0.99 NRD=24.625 NRS=3.0732 M=1 R=4.26667
+ SA=75000.7 SB=75002.3 A=0.096 P=1.58 MULT=1
MM1002 N_A_296_74#_M1002_d N_D_M1002_g A_233_464# VPB PSHORT L=0.15 W=0.64
+ AD=0.096 AS=0.0864 PD=0.94 PS=0.91 NRD=3.0732 NRS=24.625 M=1 R=4.26667
+ SA=75001.1 SB=75001.9 A=0.096 P=1.58 MULT=1
MM1006 A_407_464# N_A_31_74#_M1006_g N_A_296_74#_M1002_d VPB PSHORT L=0.15
+ W=0.64 AD=0.1248 AS=0.096 PD=1.03 PS=0.94 NRD=43.0839 NRS=3.0732 M=1 R=4.26667
+ SA=75001.6 SB=75001.5 A=0.096 P=1.58 MULT=1
MM1022 N_VPWR_M1022_d N_SCD_M1022_g A_407_464# VPB PSHORT L=0.15 W=0.64
+ AD=0.176582 AS=0.1248 PD=1.22182 PS=1.03 NRD=43.0839 NRS=43.0839 M=1 R=4.26667
+ SA=75002.1 SB=75000.9 A=0.096 P=1.58 MULT=1
MM1026 N_A_612_74#_M1026_d N_CLK_M1026_g N_VPWR_M1022_d VPB PSHORT L=0.15 W=1.12
+ AD=0.3304 AS=0.309018 PD=2.83 PS=2.13818 NRD=1.7533 NRS=24.625 M=1 R=7.46667
+ SA=75001.7 SB=75000.2 A=0.168 P=2.54 MULT=1
MM1000 N_A_828_74#_M1000_d N_A_612_74#_M1000_g N_VPWR_M1000_s VPB PSHORT L=0.15
+ W=1.12 AD=0.3136 AS=0.5264 PD=2.8 PS=3.18 NRD=1.7533 NRS=17.5724 M=1 R=7.46667
+ SA=75000.4 SB=75000.2 A=0.168 P=2.54 MULT=1
MM1019 N_A_1021_100#_M1019_d N_A_828_74#_M1019_g N_A_296_74#_M1019_s VPB PSHORT
+ L=0.15 W=0.42 AD=0.063 AS=0.1176 PD=0.72 PS=1.4 NRD=4.6886 NRS=4.6886 M=1
+ R=2.8 SA=75000.2 SB=75004.1 A=0.063 P=1.14 MULT=1
MM1023 A_1180_496# N_A_612_74#_M1023_g N_A_1021_100#_M1019_d VPB PSHORT L=0.15
+ W=0.42 AD=0.0693 AS=0.063 PD=0.75 PS=0.72 NRD=51.5943 NRS=4.6886 M=1 R=2.8
+ SA=75000.7 SB=75003.7 A=0.063 P=1.14 MULT=1
MM1007 N_VPWR_M1007_d N_A_1243_398#_M1007_g A_1180_496# VPB PSHORT L=0.15 W=0.42
+ AD=0.1255 AS=0.0693 PD=1.01333 PS=0.75 NRD=114.339 NRS=51.5943 M=1 R=2.8
+ SA=75001.1 SB=75003.2 A=0.063 P=1.14 MULT=1
MM1005 N_A_1243_398#_M1005_d N_A_1021_100#_M1005_g N_VPWR_M1007_d VPB PSHORT
+ L=0.15 W=0.84 AD=0.3234 AS=0.251 PD=1.61 PS=2.02667 NRD=0 NRS=57.1694 M=1
+ R=5.6 SA=75001 SB=75002 A=0.126 P=1.98 MULT=1
MM1012 N_A_1529_74#_M1012_d N_A_612_74#_M1012_g N_A_1243_398#_M1005_d VPB PSHORT
+ L=0.15 W=0.84 AD=0.1904 AS=0.3234 PD=1.63333 PS=1.61 NRD=2.3443 NRS=103.189
+ M=1 R=5.6 SA=75001.9 SB=75001.1 A=0.126 P=1.98 MULT=1
MM1008 A_1691_508# N_A_828_74#_M1008_g N_A_1529_74#_M1012_d VPB PSHORT L=0.15
+ W=0.42 AD=0.0567 AS=0.0952 PD=0.69 PS=0.816667 NRD=37.5088 NRS=44.5417 M=1
+ R=2.8 SA=75003 SB=75001.4 A=0.063 P=1.14 MULT=1
MM1014 N_VPWR_M1014_d N_A_1723_48#_M1014_g A_1691_508# VPB PSHORT L=0.15 W=0.42
+ AD=0.118754 AS=0.0567 PD=0.940563 PS=0.69 NRD=68.0044 NRS=37.5088 M=1 R=2.8
+ SA=75003.4 SB=75000.9 A=0.063 P=1.14 MULT=1
MM1029 N_A_1723_48#_M1029_d N_A_1529_74#_M1029_g N_VPWR_M1014_d VPB PSHORT
+ L=0.15 W=1 AD=0.275 AS=0.282746 PD=2.55 PS=2.23944 NRD=1.9503 NRS=32.4853 M=1
+ R=6.66667 SA=75001.9 SB=75000.2 A=0.15 P=2.3 MULT=1
MM1018 N_Q_M1018_d N_A_1723_48#_M1018_g N_VPWR_M1018_s VPB PSHORT L=0.15 W=1.12
+ AD=0.308 AS=0.308 PD=2.79 PS=2.79 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75000.2 A=0.168 P=2.54 MULT=1
MM1030 N_VPWR_M1030_d N_A_1723_48#_M1030_g N_A_2216_94#_M1030_s VPB PSHORT
+ L=0.15 W=0.84 AD=0.1596 AS=0.231 PD=1.26429 PS=2.23 NRD=2.3443 NRS=2.3443 M=1
+ R=5.6 SA=75000.2 SB=75000.7 A=0.126 P=1.98 MULT=1
MM1025 N_Q_N_M1025_d N_A_2216_94#_M1025_g N_VPWR_M1030_d VPB PSHORT L=0.15
+ W=1.12 AD=0.3192 AS=0.2128 PD=2.81 PS=1.68571 NRD=1.7533 NRS=11.426 M=1
+ R=7.46667 SA=75000.6 SB=75000.2 A=0.168 P=2.54 MULT=1
DX36_noxref VNB VPB NWDIODE A=23.9196 P=29.44
c_139 VNB 0 1.65961e-19 $X=0 $Y=0
c_1894 A_434_74# 0 2.47416e-20 $X=2.17 $Y=0.37
*
.include "sky130_fd_sc_hs__sdfxbp_1.pxi.spice"
*
.ends
*
*
