* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hs__nor4_1 A B C D VGND VNB VPB VPWR Y
M1000 a_342_368# C a_228_368# VPB pshort w=1.12e+06u l=150000u
+  ad=4.704e+11p pd=3.08e+06u as=4.704e+11p ps=3.08e+06u
M1001 Y A VGND VNB nlowvt w=740000u l=150000u
+  ad=4.144e+11p pd=4.08e+06u as=8.7975e+11p ps=6.9e+06u
M1002 VGND B Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1003 Y C VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_144_368# A VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=3.024e+11p pd=2.78e+06u as=3.304e+11p ps=2.83e+06u
M1005 a_228_368# B a_144_368# VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VGND D Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 Y D a_342_368# VPB pshort w=1.12e+06u l=150000u
+  ad=3.304e+11p pd=2.83e+06u as=0p ps=0u
.ends
