* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hs__dlxtn_1 D GATE_N VGND VNB VPB VPWR Q
X0 a_27_115# D VGND VNB sky130_fd_pr__nfet_01v8_lvt w=550000u l=150000u
X1 VPWR a_669_392# a_863_441# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=150000u
X2 a_669_392# a_369_392# a_871_139# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X3 a_655_79# a_217_419# a_669_392# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X4 a_27_115# D VPWR VPB sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X5 a_669_392# a_217_419# a_812_508# VPB sky130_fd_pr__pfet_01v8 w=420000u l=150000u
X6 VGND GATE_N a_217_419# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X7 VGND a_27_115# a_655_79# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X8 a_871_139# a_863_441# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X9 a_812_508# a_863_441# VPWR VPB sky130_fd_pr__pfet_01v8 w=420000u l=150000u
X10 VGND a_669_392# a_863_441# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X11 VPWR GATE_N a_217_419# VPB sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X12 VPWR a_27_115# a_585_392# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=150000u
X13 a_369_392# a_217_419# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X14 VGND a_863_441# Q VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X15 a_585_392# a_369_392# a_669_392# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=150000u
X16 VPWR a_863_441# Q VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X17 a_369_392# a_217_419# VPWR VPB sky130_fd_pr__pfet_01v8 w=840000u l=150000u
.ends
