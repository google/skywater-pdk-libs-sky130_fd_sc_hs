* File: sky130_fd_sc_hs__a2111o_1.pxi.spice
* Created: Tue Sep  1 19:47:49 2020
* 
x_PM_SKY130_FD_SC_HS__A2111O_1%A1 N_A1_c_74_n N_A1_c_75_n N_A1_c_81_n
+ N_A1_M1010_g N_A1_M1001_g A1 A1 N_A1_c_77_n N_A1_c_78_n N_A1_c_79_n
+ PM_SKY130_FD_SC_HS__A2111O_1%A1
x_PM_SKY130_FD_SC_HS__A2111O_1%A2 N_A2_M1003_g N_A2_c_113_n N_A2_M1006_g A2 A2
+ A2 PM_SKY130_FD_SC_HS__A2111O_1%A2
x_PM_SKY130_FD_SC_HS__A2111O_1%B1 N_B1_M1004_g N_B1_c_154_n N_B1_c_159_n
+ N_B1_M1007_g N_B1_c_155_n B1 N_B1_c_157_n PM_SKY130_FD_SC_HS__A2111O_1%B1
x_PM_SKY130_FD_SC_HS__A2111O_1%C1 N_C1_c_197_n N_C1_c_198_n N_C1_c_203_n
+ N_C1_M1000_g N_C1_M1005_g C1 N_C1_c_201_n PM_SKY130_FD_SC_HS__A2111O_1%C1
x_PM_SKY130_FD_SC_HS__A2111O_1%D1 N_D1_c_242_n N_D1_M1009_g N_D1_M1002_g D1
+ PM_SKY130_FD_SC_HS__A2111O_1%D1
x_PM_SKY130_FD_SC_HS__A2111O_1%A_85_136# N_A_85_136#_M1001_s N_A_85_136#_M1004_d
+ N_A_85_136#_M1002_d N_A_85_136#_M1009_d N_A_85_136#_c_283_n
+ N_A_85_136#_M1011_g N_A_85_136#_M1008_g N_A_85_136#_c_273_n
+ N_A_85_136#_c_274_n N_A_85_136#_c_275_n N_A_85_136#_c_276_n
+ N_A_85_136#_c_285_n N_A_85_136#_c_277_n N_A_85_136#_c_278_n
+ N_A_85_136#_c_279_n N_A_85_136#_c_280_n N_A_85_136#_c_281_n
+ N_A_85_136#_c_287_n N_A_85_136#_c_282_n PM_SKY130_FD_SC_HS__A2111O_1%A_85_136#
x_PM_SKY130_FD_SC_HS__A2111O_1%A_80_392# N_A_80_392#_M1010_s N_A_80_392#_M1006_d
+ N_A_80_392#_c_365_n N_A_80_392#_c_366_n N_A_80_392#_c_370_n
+ N_A_80_392#_c_375_n N_A_80_392#_c_367_n PM_SKY130_FD_SC_HS__A2111O_1%A_80_392#
x_PM_SKY130_FD_SC_HS__A2111O_1%VPWR N_VPWR_M1010_d N_VPWR_M1011_s N_VPWR_c_394_n
+ N_VPWR_c_395_n N_VPWR_c_396_n N_VPWR_c_397_n N_VPWR_c_398_n N_VPWR_c_399_n
+ VPWR N_VPWR_c_400_n N_VPWR_c_393_n PM_SKY130_FD_SC_HS__A2111O_1%VPWR
x_PM_SKY130_FD_SC_HS__A2111O_1%X N_X_M1008_d N_X_M1011_d X X X X X X X
+ PM_SKY130_FD_SC_HS__A2111O_1%X
x_PM_SKY130_FD_SC_HS__A2111O_1%VGND N_VGND_M1003_d N_VGND_M1005_d N_VGND_M1008_s
+ N_VGND_c_448_n N_VGND_c_449_n N_VGND_c_450_n N_VGND_c_451_n N_VGND_c_452_n
+ N_VGND_c_453_n N_VGND_c_454_n VGND N_VGND_c_455_n N_VGND_c_456_n
+ N_VGND_c_457_n N_VGND_c_458_n N_VGND_c_459_n N_VGND_c_460_n
+ PM_SKY130_FD_SC_HS__A2111O_1%VGND
cc_1 VNB N_A1_c_74_n 0.00825182f $X=-0.19 $Y=-0.245 $X2=0.75 $Y2=1.485
cc_2 VNB N_A1_c_75_n 0.0145126f $X=-0.19 $Y=-0.245 $X2=0.75 $Y2=1.795
cc_3 VNB N_A1_M1001_g 0.0121632f $X=-0.19 $Y=-0.245 $X2=0.765 $Y2=1
cc_4 VNB N_A1_c_77_n 0.050907f $X=-0.19 $Y=-0.245 $X2=0.675 $Y2=0.405
cc_5 VNB N_A1_c_78_n 0.00194614f $X=-0.19 $Y=-0.245 $X2=0.675 $Y2=0.405
cc_6 VNB N_A1_c_79_n 0.0248033f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=0.555
cc_7 VNB N_A2_M1003_g 0.0188883f $X=-0.19 $Y=-0.245 $X2=0.75 $Y2=1.885
cc_8 VNB N_A2_c_113_n 0.0154997f $X=-0.19 $Y=-0.245 $X2=0.75 $Y2=2.46
cc_9 VNB A2 0.00767832f $X=-0.19 $Y=-0.245 $X2=0.75 $Y2=1.395
cc_10 VNB N_B1_M1004_g 0.0116938f $X=-0.19 $Y=-0.245 $X2=0.75 $Y2=2.46
cc_11 VNB N_B1_c_154_n 0.00455744f $X=-0.19 $Y=-0.245 $X2=0.765 $Y2=0.57
cc_12 VNB N_B1_c_155_n 0.00919437f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.47
cc_13 VNB B1 0.00524134f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.47
cc_14 VNB N_B1_c_157_n 0.040608f $X=-0.19 $Y=-0.245 $X2=0.675 $Y2=0.405
cc_15 VNB N_C1_c_197_n 0.00611396f $X=-0.19 $Y=-0.245 $X2=0.75 $Y2=1.485
cc_16 VNB N_C1_c_198_n 0.0070589f $X=-0.19 $Y=-0.245 $X2=0.75 $Y2=1.795
cc_17 VNB N_C1_M1005_g 0.0115624f $X=-0.19 $Y=-0.245 $X2=0.765 $Y2=1
cc_18 VNB C1 0.0072876f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.47
cc_19 VNB N_C1_c_201_n 0.0416442f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_D1_c_242_n 0.0232231f $X=-0.19 $Y=-0.245 $X2=0.75 $Y2=1.485
cc_21 VNB N_D1_M1002_g 0.0231368f $X=-0.19 $Y=-0.245 $X2=0.765 $Y2=0.57
cc_22 VNB N_A_85_136#_M1008_g 0.0284861f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_85_136#_c_273_n 0.0416098f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=0.555
cc_24 VNB N_A_85_136#_c_274_n 0.0181306f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=0.555
cc_25 VNB N_A_85_136#_c_275_n 0.00644288f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_85_136#_c_276_n 0.00713807f $X=-0.19 $Y=-0.245 $X2=0.675 $Y2=0.405
cc_27 VNB N_A_85_136#_c_277_n 0.00982621f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_85_136#_c_278_n 2.31997e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_85_136#_c_279_n 0.0189635f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_85_136#_c_280_n 0.0244976f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_85_136#_c_281_n 0.00237362f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_85_136#_c_282_n 0.00920471f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_VPWR_c_393_n 0.183584f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB X 0.0544527f $X=-0.19 $Y=-0.245 $X2=0.765 $Y2=1.395
cc_35 VNB N_VGND_c_448_n 0.0110058f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.47
cc_36 VNB N_VGND_c_449_n 0.0193596f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_450_n 0.0287345f $X=-0.19 $Y=-0.245 $X2=0.675 $Y2=0.405
cc_38 VNB N_VGND_c_451_n 0.00222109f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=0.555
cc_39 VNB N_VGND_c_452_n 0.00158873f $X=-0.19 $Y=-0.245 $X2=0.675 $Y2=0.555
cc_40 VNB N_VGND_c_453_n 0.0314356f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_454_n 0.00326621f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_455_n 0.0311326f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_456_n 0.0229859f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_457_n 0.0198489f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_VGND_c_458_n 0.279604f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_VGND_c_459_n 0.00326621f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_VGND_c_460_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VPB N_A1_c_75_n 0.0111748f $X=-0.19 $Y=1.66 $X2=0.75 $Y2=1.795
cc_49 VPB N_A1_c_81_n 0.0298714f $X=-0.19 $Y=1.66 $X2=0.75 $Y2=1.885
cc_50 VPB N_A2_c_113_n 0.0338491f $X=-0.19 $Y=1.66 $X2=0.75 $Y2=2.46
cc_51 VPB A2 0.0160983f $X=-0.19 $Y=1.66 $X2=0.75 $Y2=1.395
cc_52 VPB N_B1_c_154_n 0.00535699f $X=-0.19 $Y=1.66 $X2=0.765 $Y2=0.57
cc_53 VPB N_B1_c_159_n 0.0217288f $X=-0.19 $Y=1.66 $X2=0.765 $Y2=1.395
cc_54 VPB N_C1_c_198_n 0.00529161f $X=-0.19 $Y=1.66 $X2=0.75 $Y2=1.795
cc_55 VPB N_C1_c_203_n 0.0216318f $X=-0.19 $Y=1.66 $X2=0.75 $Y2=1.885
cc_56 VPB N_D1_c_242_n 0.0436163f $X=-0.19 $Y=1.66 $X2=0.75 $Y2=1.485
cc_57 VPB N_A_85_136#_c_283_n 0.0209961f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_58 VPB N_A_85_136#_c_274_n 0.00944798f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=0.555
cc_59 VPB N_A_85_136#_c_285_n 0.0170442f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_60 VPB N_A_85_136#_c_278_n 0.00871481f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_61 VPB N_A_85_136#_c_287_n 0.0145556f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_62 VPB N_A_80_392#_c_365_n 0.0140928f $X=-0.19 $Y=1.66 $X2=0.765 $Y2=1.395
cc_63 VPB N_A_80_392#_c_366_n 0.0352424f $X=-0.19 $Y=1.66 $X2=0.765 $Y2=1
cc_64 VPB N_A_80_392#_c_367_n 0.00257348f $X=-0.19 $Y=1.66 $X2=0.675 $Y2=0.405
cc_65 VPB N_VPWR_c_394_n 0.00847102f $X=-0.19 $Y=1.66 $X2=0.765 $Y2=1
cc_66 VPB N_VPWR_c_395_n 0.0314654f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_67 VPB N_VPWR_c_396_n 0.0279026f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_68 VPB N_VPWR_c_397_n 0.00401341f $X=-0.19 $Y=1.66 $X2=0.675 $Y2=0.57
cc_69 VPB N_VPWR_c_398_n 0.0683206f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=0.555
cc_70 VPB N_VPWR_c_399_n 0.0047828f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_71 VPB N_VPWR_c_400_n 0.0205444f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_72 VPB N_VPWR_c_393_n 0.115904f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_73 VPB X 0.0547727f $X=-0.19 $Y=1.66 $X2=0.765 $Y2=1.395
cc_74 N_A1_c_77_n N_A2_M1003_g 0.0379734f $X=0.675 $Y=0.405 $X2=0 $Y2=0
cc_75 N_A1_c_78_n N_A2_M1003_g 3.79132e-19 $X=0.675 $Y=0.405 $X2=0 $Y2=0
cc_76 N_A1_c_74_n N_A2_c_113_n 0.0379734f $X=0.75 $Y=1.485 $X2=0 $Y2=0
cc_77 N_A1_c_81_n N_A2_c_113_n 0.0214432f $X=0.75 $Y=1.885 $X2=0 $Y2=0
cc_78 N_A1_c_75_n A2 0.00199456f $X=0.75 $Y=1.795 $X2=0 $Y2=0
cc_79 N_A1_c_77_n N_B1_c_157_n 0.00402835f $X=0.675 $Y=0.405 $X2=0 $Y2=0
cc_80 N_A1_M1001_g N_A_85_136#_c_275_n 0.010511f $X=0.765 $Y=1 $X2=0 $Y2=0
cc_81 N_A1_c_78_n N_A_85_136#_c_275_n 0.00381804f $X=0.675 $Y=0.405 $X2=0 $Y2=0
cc_82 N_A1_c_74_n N_A_85_136#_c_280_n 0.00110067f $X=0.75 $Y=1.485 $X2=0 $Y2=0
cc_83 N_A1_M1001_g N_A_85_136#_c_280_n 0.00945732f $X=0.765 $Y=1 $X2=0 $Y2=0
cc_84 N_A1_c_77_n N_A_85_136#_c_280_n 9.34446e-19 $X=0.675 $Y=0.405 $X2=0 $Y2=0
cc_85 N_A1_c_78_n N_A_85_136#_c_280_n 0.0146521f $X=0.675 $Y=0.405 $X2=0 $Y2=0
cc_86 N_A1_c_79_n N_A_85_136#_c_280_n 0.0100266f $X=0.51 $Y=0.555 $X2=0 $Y2=0
cc_87 N_A1_c_81_n N_A_80_392#_c_365_n 0.00208878f $X=0.75 $Y=1.885 $X2=0 $Y2=0
cc_88 N_A1_c_81_n N_A_80_392#_c_366_n 0.0104767f $X=0.75 $Y=1.885 $X2=0 $Y2=0
cc_89 N_A1_c_81_n N_A_80_392#_c_370_n 0.0140828f $X=0.75 $Y=1.885 $X2=0 $Y2=0
cc_90 N_A1_c_81_n N_A_80_392#_c_367_n 6.28237e-19 $X=0.75 $Y=1.885 $X2=0 $Y2=0
cc_91 N_A1_c_81_n N_VPWR_c_394_n 0.00507763f $X=0.75 $Y=1.885 $X2=0 $Y2=0
cc_92 N_A1_c_81_n N_VPWR_c_396_n 0.00445602f $X=0.75 $Y=1.885 $X2=0 $Y2=0
cc_93 N_A1_c_81_n N_VPWR_c_393_n 0.0086209f $X=0.75 $Y=1.885 $X2=0 $Y2=0
cc_94 N_A1_c_77_n N_VGND_c_448_n 0.0035084f $X=0.675 $Y=0.405 $X2=0 $Y2=0
cc_95 N_A1_c_78_n N_VGND_c_448_n 0.0220302f $X=0.675 $Y=0.405 $X2=0 $Y2=0
cc_96 N_A1_M1001_g N_VGND_c_451_n 0.00150526f $X=0.765 $Y=1 $X2=0 $Y2=0
cc_97 N_A1_c_78_n N_VGND_c_451_n 4.9027e-19 $X=0.675 $Y=0.405 $X2=0 $Y2=0
cc_98 N_A1_c_77_n N_VGND_c_455_n 0.00586744f $X=0.675 $Y=0.405 $X2=0 $Y2=0
cc_99 N_A1_c_78_n N_VGND_c_455_n 0.0215843f $X=0.675 $Y=0.405 $X2=0 $Y2=0
cc_100 N_A1_c_79_n N_VGND_c_455_n 0.0116351f $X=0.51 $Y=0.555 $X2=0 $Y2=0
cc_101 N_A1_c_77_n N_VGND_c_458_n 0.00754663f $X=0.675 $Y=0.405 $X2=0 $Y2=0
cc_102 N_A1_c_78_n N_VGND_c_458_n 0.0110944f $X=0.675 $Y=0.405 $X2=0 $Y2=0
cc_103 N_A1_c_79_n N_VGND_c_458_n 0.0128919f $X=0.51 $Y=0.555 $X2=0 $Y2=0
cc_104 N_A2_M1003_g N_B1_M1004_g 0.0221727f $X=1.125 $Y=1 $X2=0 $Y2=0
cc_105 N_A2_c_113_n N_B1_c_154_n 0.0155155f $X=1.24 $Y=1.885 $X2=0 $Y2=0
cc_106 A2 N_B1_c_154_n 0.00876296f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_107 N_A2_c_113_n N_B1_c_159_n 0.0137237f $X=1.24 $Y=1.885 $X2=0 $Y2=0
cc_108 A2 N_B1_c_159_n 0.0073676f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_109 N_A2_c_113_n N_B1_c_155_n 0.00505817f $X=1.24 $Y=1.885 $X2=0 $Y2=0
cc_110 A2 N_B1_c_155_n 0.00417922f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_111 A2 N_C1_c_198_n 0.0112402f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_112 A2 N_C1_c_203_n 0.00835824f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_113 A2 N_D1_c_242_n 0.0021316f $X=2.075 $Y=1.58 $X2=-0.19 $Y2=-0.245
cc_114 A2 D1 0.0252516f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_115 N_A2_M1003_g N_A_85_136#_c_275_n 0.011795f $X=1.125 $Y=1 $X2=0 $Y2=0
cc_116 N_A2_c_113_n N_A_85_136#_c_275_n 0.00466536f $X=1.24 $Y=1.885 $X2=0 $Y2=0
cc_117 A2 N_A_85_136#_c_275_n 0.0494435f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_118 A2 N_A_85_136#_c_276_n 0.017121f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_119 N_A2_M1003_g N_A_85_136#_c_280_n 0.00137574f $X=1.125 $Y=1 $X2=0 $Y2=0
cc_120 N_A2_M1003_g N_A_85_136#_c_281_n 8.00461e-19 $X=1.125 $Y=1 $X2=0 $Y2=0
cc_121 A2 N_A_85_136#_c_281_n 0.0273946f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_122 N_A2_c_113_n N_A_80_392#_c_366_n 6.28237e-19 $X=1.24 $Y=1.885 $X2=0 $Y2=0
cc_123 N_A2_c_113_n N_A_80_392#_c_370_n 0.0147139f $X=1.24 $Y=1.885 $X2=0 $Y2=0
cc_124 A2 N_A_80_392#_c_370_n 0.0158922f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_125 N_A2_c_113_n N_A_80_392#_c_375_n 0.00146386f $X=1.24 $Y=1.885 $X2=0 $Y2=0
cc_126 A2 N_A_80_392#_c_375_n 0.0226807f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_127 N_A2_c_113_n N_A_80_392#_c_367_n 0.010325f $X=1.24 $Y=1.885 $X2=0 $Y2=0
cc_128 N_A2_c_113_n N_VPWR_c_394_n 0.00507763f $X=1.24 $Y=1.885 $X2=0 $Y2=0
cc_129 N_A2_c_113_n N_VPWR_c_398_n 0.00445602f $X=1.24 $Y=1.885 $X2=0 $Y2=0
cc_130 N_A2_c_113_n N_VPWR_c_393_n 0.00858105f $X=1.24 $Y=1.885 $X2=0 $Y2=0
cc_131 N_A2_M1003_g N_VGND_c_448_n 0.00547724f $X=1.125 $Y=1 $X2=0 $Y2=0
cc_132 N_A2_M1003_g N_VGND_c_451_n 0.00908429f $X=1.125 $Y=1 $X2=0 $Y2=0
cc_133 N_A2_M1003_g N_VGND_c_455_n 0.00115433f $X=1.125 $Y=1 $X2=0 $Y2=0
cc_134 N_A2_M1003_g N_VGND_c_458_n 0.00139378f $X=1.125 $Y=1 $X2=0 $Y2=0
cc_135 N_B1_c_155_n N_C1_c_197_n 0.010711f $X=1.685 $Y=1.545 $X2=-0.19
+ $Y2=-0.245
cc_136 N_B1_c_154_n N_C1_c_198_n 0.010711f $X=1.69 $Y=1.795 $X2=0 $Y2=0
cc_137 N_B1_c_159_n N_C1_c_203_n 0.0761177f $X=1.69 $Y=1.885 $X2=0 $Y2=0
cc_138 N_B1_M1004_g N_C1_M1005_g 0.0213181f $X=1.665 $Y=1 $X2=0 $Y2=0
cc_139 B1 N_C1_M1005_g 4.39948e-19 $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_140 N_B1_M1004_g C1 4.14714e-19 $X=1.665 $Y=1 $X2=0 $Y2=0
cc_141 B1 C1 0.0281802f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_142 N_B1_c_157_n C1 3.38136e-19 $X=1.6 $Y=0.37 $X2=0 $Y2=0
cc_143 B1 N_C1_c_201_n 9.98522e-19 $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_144 N_B1_c_157_n N_C1_c_201_n 0.0185027f $X=1.6 $Y=0.37 $X2=0 $Y2=0
cc_145 N_B1_M1004_g N_A_85_136#_c_275_n 0.00979317f $X=1.665 $Y=1 $X2=0 $Y2=0
cc_146 B1 N_A_85_136#_c_275_n 0.00683244f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_147 N_B1_c_157_n N_A_85_136#_c_275_n 0.002282f $X=1.6 $Y=0.37 $X2=0 $Y2=0
cc_148 N_B1_M1004_g N_A_85_136#_c_281_n 0.00810118f $X=1.665 $Y=1 $X2=0 $Y2=0
cc_149 N_B1_c_155_n N_A_85_136#_c_281_n 0.00118931f $X=1.685 $Y=1.545 $X2=0
+ $Y2=0
cc_150 B1 N_A_85_136#_c_281_n 0.0042544f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_151 N_B1_c_159_n N_A_80_392#_c_375_n 0.00333375f $X=1.69 $Y=1.885 $X2=0 $Y2=0
cc_152 N_B1_c_159_n N_A_80_392#_c_367_n 0.0145945f $X=1.69 $Y=1.885 $X2=0 $Y2=0
cc_153 N_B1_c_159_n N_VPWR_c_398_n 0.00445602f $X=1.69 $Y=1.885 $X2=0 $Y2=0
cc_154 N_B1_c_159_n N_VPWR_c_393_n 0.00857948f $X=1.69 $Y=1.885 $X2=0 $Y2=0
cc_155 N_B1_M1004_g N_VGND_c_448_n 9.4076e-19 $X=1.665 $Y=1 $X2=0 $Y2=0
cc_156 B1 N_VGND_c_448_n 0.0253807f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_157 N_B1_c_157_n N_VGND_c_448_n 0.0028006f $X=1.6 $Y=0.37 $X2=0 $Y2=0
cc_158 N_B1_M1004_g N_VGND_c_451_n 0.00558866f $X=1.665 $Y=1 $X2=0 $Y2=0
cc_159 B1 N_VGND_c_451_n 6.94247e-19 $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_160 B1 N_VGND_c_453_n 0.0233865f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_161 N_B1_c_157_n N_VGND_c_453_n 0.00623567f $X=1.6 $Y=0.37 $X2=0 $Y2=0
cc_162 B1 N_VGND_c_458_n 0.0122355f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_163 N_B1_c_157_n N_VGND_c_458_n 0.00873446f $X=1.6 $Y=0.37 $X2=0 $Y2=0
cc_164 N_C1_c_197_n N_D1_c_242_n 0.026715f $X=2.08 $Y=1.485 $X2=-0.19 $Y2=-0.245
cc_165 N_C1_c_203_n N_D1_c_242_n 0.0654165f $X=2.08 $Y=1.885 $X2=-0.19
+ $Y2=-0.245
cc_166 N_C1_M1005_g N_D1_M1002_g 0.0170371f $X=2.095 $Y=1 $X2=0 $Y2=0
cc_167 C1 N_D1_M1002_g 3.54912e-19 $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_168 N_C1_c_198_n D1 2.74575e-19 $X=2.08 $Y=1.795 $X2=0 $Y2=0
cc_169 N_C1_M1005_g N_A_85_136#_c_276_n 0.0100922f $X=2.095 $Y=1 $X2=0 $Y2=0
cc_170 C1 N_A_85_136#_c_276_n 0.0078915f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_171 N_C1_c_201_n N_A_85_136#_c_276_n 0.00161934f $X=2.17 $Y=0.37 $X2=0 $Y2=0
cc_172 N_C1_c_203_n N_A_85_136#_c_285_n 0.00408342f $X=2.08 $Y=1.885 $X2=0 $Y2=0
cc_173 N_C1_c_197_n N_A_85_136#_c_281_n 8.83432e-19 $X=2.08 $Y=1.485 $X2=0 $Y2=0
cc_174 N_C1_M1005_g N_A_85_136#_c_281_n 0.0086072f $X=2.095 $Y=1 $X2=0 $Y2=0
cc_175 C1 N_A_85_136#_c_281_n 0.00251454f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_176 N_C1_c_203_n N_A_85_136#_c_287_n 8.11289e-19 $X=2.08 $Y=1.885 $X2=0 $Y2=0
cc_177 N_C1_c_203_n N_A_80_392#_c_375_n 8.18438e-19 $X=2.08 $Y=1.885 $X2=0 $Y2=0
cc_178 N_C1_c_203_n N_A_80_392#_c_367_n 0.00408054f $X=2.08 $Y=1.885 $X2=0 $Y2=0
cc_179 N_C1_c_203_n N_VPWR_c_398_n 0.00461464f $X=2.08 $Y=1.885 $X2=0 $Y2=0
cc_180 N_C1_c_203_n N_VPWR_c_393_n 0.00908738f $X=2.08 $Y=1.885 $X2=0 $Y2=0
cc_181 N_C1_M1005_g N_VGND_c_449_n 4.35288e-19 $X=2.095 $Y=1 $X2=0 $Y2=0
cc_182 C1 N_VGND_c_449_n 0.0273749f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_183 N_C1_c_201_n N_VGND_c_449_n 0.00422608f $X=2.17 $Y=0.37 $X2=0 $Y2=0
cc_184 N_C1_M1005_g N_VGND_c_452_n 0.00511653f $X=2.095 $Y=1 $X2=0 $Y2=0
cc_185 C1 N_VGND_c_452_n 7.25307e-19 $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_186 C1 N_VGND_c_453_n 0.0214896f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_187 N_C1_c_201_n N_VGND_c_453_n 0.00623567f $X=2.17 $Y=0.37 $X2=0 $Y2=0
cc_188 C1 N_VGND_c_458_n 0.011118f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_189 N_C1_c_201_n N_VGND_c_458_n 0.00876197f $X=2.17 $Y=0.37 $X2=0 $Y2=0
cc_190 N_D1_M1002_g N_A_85_136#_c_273_n 0.00470073f $X=2.715 $Y=1 $X2=0 $Y2=0
cc_191 N_D1_c_242_n N_A_85_136#_c_276_n 0.00769547f $X=2.47 $Y=1.885 $X2=0 $Y2=0
cc_192 N_D1_M1002_g N_A_85_136#_c_276_n 0.0128941f $X=2.715 $Y=1 $X2=0 $Y2=0
cc_193 D1 N_A_85_136#_c_276_n 0.0241162f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_194 N_D1_c_242_n N_A_85_136#_c_285_n 0.0148434f $X=2.47 $Y=1.885 $X2=0 $Y2=0
cc_195 N_D1_M1002_g N_A_85_136#_c_277_n 4.47467e-19 $X=2.715 $Y=1 $X2=0 $Y2=0
cc_196 N_D1_c_242_n N_A_85_136#_c_278_n 0.00809159f $X=2.47 $Y=1.885 $X2=0 $Y2=0
cc_197 D1 N_A_85_136#_c_278_n 0.0112155f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_198 N_D1_M1002_g N_A_85_136#_c_281_n 7.63247e-19 $X=2.715 $Y=1 $X2=0 $Y2=0
cc_199 N_D1_c_242_n N_A_85_136#_c_287_n 0.0090023f $X=2.47 $Y=1.885 $X2=0 $Y2=0
cc_200 D1 N_A_85_136#_c_287_n 0.0158167f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_201 N_D1_M1002_g N_A_85_136#_c_282_n 0.00696805f $X=2.715 $Y=1 $X2=0 $Y2=0
cc_202 D1 N_A_85_136#_c_282_n 0.0126267f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_203 N_D1_c_242_n N_VPWR_c_398_n 0.00445602f $X=2.47 $Y=1.885 $X2=0 $Y2=0
cc_204 N_D1_c_242_n N_VPWR_c_393_n 0.00862666f $X=2.47 $Y=1.885 $X2=0 $Y2=0
cc_205 N_D1_M1002_g N_VGND_c_449_n 0.00661179f $X=2.715 $Y=1 $X2=0 $Y2=0
cc_206 N_D1_M1002_g N_VGND_c_450_n 0.00331675f $X=2.715 $Y=1 $X2=0 $Y2=0
cc_207 N_D1_M1002_g N_VGND_c_452_n 0.0045349f $X=2.715 $Y=1 $X2=0 $Y2=0
cc_208 N_D1_M1002_g N_VGND_c_456_n 0.00296257f $X=2.715 $Y=1 $X2=0 $Y2=0
cc_209 N_D1_M1002_g N_VGND_c_458_n 0.00351476f $X=2.715 $Y=1 $X2=0 $Y2=0
cc_210 N_A_85_136#_c_280_n N_A_80_392#_c_365_n 0.0114345f $X=0.55 $Y=1.09 $X2=0
+ $Y2=0
cc_211 N_A_85_136#_c_275_n N_A_80_392#_c_370_n 0.0080253f $X=1.715 $Y=1.245
+ $X2=0 $Y2=0
cc_212 N_A_85_136#_c_280_n N_A_80_392#_c_370_n 5.86784e-19 $X=0.55 $Y=1.09 $X2=0
+ $Y2=0
cc_213 N_A_85_136#_c_283_n N_VPWR_c_395_n 0.0100916f $X=3.8 $Y=1.765 $X2=0 $Y2=0
cc_214 N_A_85_136#_c_273_n N_VPWR_c_395_n 0.00577732f $X=3.71 $Y=1.485 $X2=0
+ $Y2=0
cc_215 N_A_85_136#_c_285_n N_VPWR_c_395_n 0.0303536f $X=2.695 $Y=2.815 $X2=0
+ $Y2=0
cc_216 N_A_85_136#_c_278_n N_VPWR_c_395_n 0.00793894f $X=3.03 $Y=1.97 $X2=0
+ $Y2=0
cc_217 N_A_85_136#_c_279_n N_VPWR_c_395_n 0.0209147f $X=3.525 $Y=1.485 $X2=0
+ $Y2=0
cc_218 N_A_85_136#_c_287_n N_VPWR_c_395_n 0.00980487f $X=3.03 $Y=2.055 $X2=0
+ $Y2=0
cc_219 N_A_85_136#_c_285_n N_VPWR_c_398_n 0.0145938f $X=2.695 $Y=2.815 $X2=0
+ $Y2=0
cc_220 N_A_85_136#_c_283_n N_VPWR_c_400_n 0.00445602f $X=3.8 $Y=1.765 $X2=0
+ $Y2=0
cc_221 N_A_85_136#_c_283_n N_VPWR_c_393_n 0.00865934f $X=3.8 $Y=1.765 $X2=0
+ $Y2=0
cc_222 N_A_85_136#_c_285_n N_VPWR_c_393_n 0.0120466f $X=2.695 $Y=2.815 $X2=0
+ $Y2=0
cc_223 N_A_85_136#_c_283_n X 0.0178122f $X=3.8 $Y=1.765 $X2=0 $Y2=0
cc_224 N_A_85_136#_M1008_g X 0.0217973f $X=3.815 $Y=0.76 $X2=0 $Y2=0
cc_225 N_A_85_136#_c_274_n X 0.0199666f $X=3.8 $Y=1.542 $X2=0 $Y2=0
cc_226 N_A_85_136#_c_279_n X 0.026211f $X=3.525 $Y=1.485 $X2=0 $Y2=0
cc_227 N_A_85_136#_c_275_n A_168_136# 0.00366293f $X=1.715 $Y=1.245 $X2=-0.19
+ $Y2=-0.245
cc_228 N_A_85_136#_c_275_n N_VGND_M1003_d 0.00421607f $X=1.715 $Y=1.245
+ $X2=-0.19 $Y2=-0.245
cc_229 N_A_85_136#_c_276_n N_VGND_M1005_d 0.00772935f $X=2.845 $Y=1.245 $X2=0
+ $Y2=0
cc_230 N_A_85_136#_M1008_g N_VGND_c_450_n 0.00650419f $X=3.815 $Y=0.76 $X2=0
+ $Y2=0
cc_231 N_A_85_136#_c_273_n N_VGND_c_450_n 0.00577732f $X=3.71 $Y=1.485 $X2=0
+ $Y2=0
cc_232 N_A_85_136#_c_277_n N_VGND_c_450_n 0.0253945f $X=2.93 $Y=0.825 $X2=0
+ $Y2=0
cc_233 N_A_85_136#_c_279_n N_VGND_c_450_n 0.0209147f $X=3.525 $Y=1.485 $X2=0
+ $Y2=0
cc_234 N_A_85_136#_c_275_n N_VGND_c_451_n 0.0202621f $X=1.715 $Y=1.245 $X2=0
+ $Y2=0
cc_235 N_A_85_136#_c_280_n N_VGND_c_451_n 0.00587041f $X=0.55 $Y=1.09 $X2=0
+ $Y2=0
cc_236 N_A_85_136#_c_281_n N_VGND_c_451_n 0.00770511f $X=1.88 $Y=1.085 $X2=0
+ $Y2=0
cc_237 N_A_85_136#_c_276_n N_VGND_c_452_n 0.0152633f $X=2.845 $Y=1.245 $X2=0
+ $Y2=0
cc_238 N_A_85_136#_c_277_n N_VGND_c_452_n 0.0126658f $X=2.93 $Y=0.825 $X2=0
+ $Y2=0
cc_239 N_A_85_136#_c_281_n N_VGND_c_452_n 0.0062632f $X=1.88 $Y=1.085 $X2=0
+ $Y2=0
cc_240 N_A_85_136#_c_277_n N_VGND_c_456_n 0.00515577f $X=2.93 $Y=0.825 $X2=0
+ $Y2=0
cc_241 N_A_85_136#_M1008_g N_VGND_c_457_n 0.00532065f $X=3.815 $Y=0.76 $X2=0
+ $Y2=0
cc_242 N_A_85_136#_M1008_g N_VGND_c_458_n 0.00539454f $X=3.815 $Y=0.76 $X2=0
+ $Y2=0
cc_243 N_A_85_136#_c_277_n N_VGND_c_458_n 0.00798209f $X=2.93 $Y=0.825 $X2=0
+ $Y2=0
cc_244 N_A_85_136#_c_280_n N_VGND_c_458_n 5.92647e-19 $X=0.55 $Y=1.09 $X2=0
+ $Y2=0
cc_245 N_A_85_136#_c_281_n N_VGND_c_458_n 0.00820329f $X=1.88 $Y=1.085 $X2=0
+ $Y2=0
cc_246 N_A_80_392#_c_370_n N_VPWR_M1010_d 0.00684424f $X=1.3 $Y=2.055 $X2=-0.19
+ $Y2=1.66
cc_247 N_A_80_392#_c_366_n N_VPWR_c_394_n 0.0443643f $X=0.525 $Y=2.815 $X2=0
+ $Y2=0
cc_248 N_A_80_392#_c_370_n N_VPWR_c_394_n 0.0169226f $X=1.3 $Y=2.055 $X2=0 $Y2=0
cc_249 N_A_80_392#_c_367_n N_VPWR_c_394_n 0.0443643f $X=1.465 $Y=2.815 $X2=0
+ $Y2=0
cc_250 N_A_80_392#_c_366_n N_VPWR_c_396_n 0.0145938f $X=0.525 $Y=2.815 $X2=0
+ $Y2=0
cc_251 N_A_80_392#_c_367_n N_VPWR_c_398_n 0.014552f $X=1.465 $Y=2.815 $X2=0
+ $Y2=0
cc_252 N_A_80_392#_c_366_n N_VPWR_c_393_n 0.0120466f $X=0.525 $Y=2.815 $X2=0
+ $Y2=0
cc_253 N_A_80_392#_c_367_n N_VPWR_c_393_n 0.0119791f $X=1.465 $Y=2.815 $X2=0
+ $Y2=0
cc_254 N_VPWR_c_395_n X 0.0779264f $X=3.575 $Y=1.985 $X2=0 $Y2=0
cc_255 N_VPWR_c_400_n X 0.0148169f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_256 N_VPWR_c_393_n X 0.0122313f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_257 X N_VGND_c_450_n 0.0301457f $X=3.995 $Y=0.47 $X2=0 $Y2=0
cc_258 X N_VGND_c_457_n 0.0136693f $X=3.995 $Y=0.47 $X2=0 $Y2=0
cc_259 X N_VGND_c_458_n 0.0121248f $X=3.995 $Y=0.47 $X2=0 $Y2=0
