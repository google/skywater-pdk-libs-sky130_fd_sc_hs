* File: sky130_fd_sc_hs__a22o_2.spice
* Created: Tue Sep  1 19:51:12 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hs__a22o_2.pex.spice"
.subckt sky130_fd_sc_hs__a22o_2  VNB VPB A1 B1 B2 A2 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A2	A2
* B2	B2
* B1	B1
* A1	A1
* VPB	VPB
* VNB	VNB
MM1000 N_VGND_M1000_d N_A_81_48#_M1000_g N_X_M1000_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1961 AS=0.1036 PD=2.01 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1010 N_VGND_M1010_d N_A_81_48#_M1010_g N_X_M1000_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1961 AS=0.1036 PD=2.01 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.6
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1009 N_A_81_48#_M1009_d N_A1_M1009_g N_A_304_74#_M1009_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1295 AS=0.2109 PD=1.09 PS=2.05 NRD=11.34 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75001.6 A=0.111 P=1.78 MULT=1
MM1007 A_491_74# N_B1_M1007_g N_A_81_48#_M1009_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.0925 AS=0.1295 PD=0.99 PS=1.09 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75000.7
+ SB=75001.1 A=0.111 P=1.78 MULT=1
MM1011 N_VGND_M1011_d N_B2_M1011_g A_491_74# VNB NLOWVT L=0.15 W=0.74 AD=0.1443
+ AS=0.0925 PD=1.13 PS=0.99 NRD=6.48 NRS=11.34 M=1 R=4.93333 SA=75001.1
+ SB=75000.7 A=0.111 P=1.78 MULT=1
MM1006 N_A_304_74#_M1006_d N_A2_M1006_g N_VGND_M1011_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.1443 PD=2.05 PS=1.13 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75001.6
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1001 N_X_M1001_d N_A_81_48#_M1001_g N_VPWR_M1001_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.308 PD=1.42 PS=2.79 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75002.4 A=0.168 P=2.54 MULT=1
MM1002 N_X_M1001_d N_A_81_48#_M1002_g N_VPWR_M1002_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.222838 PD=1.42 PS=1.59547 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.6 SB=75002 A=0.168 P=2.54 MULT=1
MM1003 N_A_388_368#_M1003_d N_A1_M1003_g N_VPWR_M1002_s VPB PSHORT L=0.15 W=1
+ AD=0.15 AS=0.198962 PD=1.3 PS=1.42453 NRD=1.9503 NRS=19.7 M=1 R=6.66667
+ SA=75001.2 SB=75001.7 A=0.15 P=2.3 MULT=1
MM1004 N_A_81_48#_M1004_d N_B1_M1004_g N_A_388_368#_M1003_d VPB PSHORT L=0.15
+ W=1 AD=0.175 AS=0.15 PD=1.35 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=6.66667
+ SA=75001.6 SB=75001.2 A=0.15 P=2.3 MULT=1
MM1005 N_A_388_368#_M1005_d N_B2_M1005_g N_A_81_48#_M1004_d VPB PSHORT L=0.15
+ W=1 AD=0.185 AS=0.175 PD=1.37 PS=1.35 NRD=3.9203 NRS=11.8003 M=1 R=6.66667
+ SA=75002.1 SB=75000.7 A=0.15 P=2.3 MULT=1
MM1008 N_VPWR_M1008_d N_A2_M1008_g N_A_388_368#_M1005_d VPB PSHORT L=0.15 W=1
+ AD=0.275 AS=0.185 PD=2.55 PS=1.37 NRD=1.9503 NRS=13.7703 M=1 R=6.66667
+ SA=75002.7 SB=75000.2 A=0.15 P=2.3 MULT=1
DX12_noxref VNB VPB NWDIODE A=7.8492 P=12.16
c_453 A_491_74# 0 1.11531e-19 $X=2.455 $Y=0.37
*
.include "sky130_fd_sc_hs__a22o_2.pxi.spice"
*
.ends
*
*
