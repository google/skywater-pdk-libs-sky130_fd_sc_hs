* File: sky130_fd_sc_hs__decap_8.pex.spice
* Created: Thu Aug 27 20:37:42 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HS__DECAP_8%VGND 1 12 17 20 22 25 29 33 36 38 44 49 56
+ 57 63 66
r41 66 67 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r42 63 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r43 60 61 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r44 57 67 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=2.64
+ $Y2=0
r45 56 57 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r46 54 66 13.6613 $w=1.7e-07 $l=3.5e-07 $layer=LI1_cond $X=3.055 $Y=0 $X2=2.705
+ $Y2=0
r47 54 56 35.5561 $w=1.68e-07 $l=5.45e-07 $layer=LI1_cond $X=3.055 $Y=0 $X2=3.6
+ $Y2=0
r48 53 67 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r49 52 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r50 50 63 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.78 $Y=0 $X2=1.615
+ $Y2=0
r51 50 52 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=1.78 $Y=0 $X2=2.16
+ $Y2=0
r52 49 66 13.6613 $w=1.7e-07 $l=3.5e-07 $layer=LI1_cond $X=2.355 $Y=0 $X2=2.705
+ $Y2=0
r53 49 52 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=2.355 $Y=0 $X2=2.16
+ $Y2=0
r54 48 64 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=1.68
+ $Y2=0
r55 48 61 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.24
+ $Y2=0
r56 47 48 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r57 45 60 6.71932 $w=1.7e-07 $l=3.7e-07 $layer=LI1_cond $X=0.74 $Y=0 $X2=0.37
+ $Y2=0
r58 45 47 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=0.74 $Y=0 $X2=1.2
+ $Y2=0
r59 44 63 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.45 $Y=0 $X2=1.615
+ $Y2=0
r60 44 47 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=1.45 $Y=0 $X2=1.2
+ $Y2=0
r61 38 53 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=2.16
+ $Y2=0
r62 38 64 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=1.68
+ $Y2=0
r63 35 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.52
+ $Y=1.42 $X2=2.52 $Y2=1.42
r64 33 35 13.3277 $w=6.98e-07 $l=7.8e-07 $layer=LI1_cond $X=2.705 $Y=0.64
+ $X2=2.705 $Y2=1.42
r65 31 66 2.86223 $w=7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.705 $Y=0.085
+ $X2=2.705 $Y2=0
r66 31 33 9.48319 $w=6.98e-07 $l=5.55e-07 $layer=LI1_cond $X=2.705 $Y=0.085
+ $X2=2.705 $Y2=0.64
r67 27 63 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.615 $Y=0.085
+ $X2=1.615 $Y2=0
r68 27 29 19.382 $w=3.28e-07 $l=5.55e-07 $layer=LI1_cond $X=1.615 $Y=0.085
+ $X2=1.615 $Y2=0.64
r69 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.575
+ $Y=1.42 $X2=0.575 $Y2=1.42
r70 22 24 16.3674 $w=5.68e-07 $l=7.8e-07 $layer=LI1_cond $X=0.455 $Y=0.64
+ $X2=0.455 $Y2=1.42
r71 20 60 3.08726 $w=5.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.455 $Y=0.085
+ $X2=0.37 $Y2=0
r72 20 22 11.646 $w=5.68e-07 $l=5.55e-07 $layer=LI1_cond $X=0.455 $Y=0.085
+ $X2=0.455 $Y2=0.64
r73 18 36 71.6931 $w=3.3e-07 $l=4.1e-07 $layer=POLY_cond $X=2.52 $Y=1.83
+ $X2=2.52 $Y2=1.42
r74 17 18 57.2398 $w=1e-06 $l=6.3e-07 $layer=POLY_cond $X=2.185 $Y=2.46
+ $X2=2.185 $Y2=1.83
r75 13 25 71.6931 $w=3.3e-07 $l=4.1e-07 $layer=POLY_cond $X=0.575 $Y=1.83
+ $X2=0.575 $Y2=1.42
r76 12 13 57.2398 $w=1e-06 $l=6.3e-07 $layer=POLY_cond $X=0.91 $Y=2.46 $X2=0.91
+ $Y2=1.83
r77 1 33 182 $w=1.7e-07 $l=2.7627e-07 $layer=licon1_NDIFF $count=1 $X=2.75
+ $Y=0.425 $X2=2.89 $Y2=0.64
r78 1 29 182 $w=1.7e-07 $l=2.7627e-07 $layer=licon1_NDIFF $count=1 $X=1.475
+ $Y=0.425 $X2=1.615 $Y2=0.64
r79 1 22 182 $w=1.7e-07 $l=2.7037e-07 $layer=licon1_NDIFF $count=1 $X=1.475
+ $Y=0.425 $X2=0.335 $Y2=0.64
.ends

.subckt PM_SKY130_FD_SC_HS__DECAP_8%VPWR 1 10 12 16 20 21 29 34 35 36 39 42 48
+ 49 55
r38 56 58 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r39 55 58 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r40 55 56 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r41 53 58 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=1.2 $Y2=3.33
r42 52 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r43 48 49 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r44 46 49 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.6 $Y2=3.33
r45 45 46 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r46 43 55 15.7884 $w=1.7e-07 $l=4.68e-07 $layer=LI1_cond $X=2.08 $Y=3.33
+ $X2=1.612 $Y2=3.33
r47 43 45 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=2.08 $Y=3.33
+ $X2=2.64 $Y2=3.33
r48 36 46 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=2.64 $Y2=3.33
r49 36 56 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=1.68 $Y2=3.33
r50 34 45 1.30481 $w=1.68e-07 $l=2e-08 $layer=LI1_cond $X=2.66 $Y=3.33 $X2=2.64
+ $Y2=3.33
r51 34 35 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.66 $Y=3.33
+ $X2=2.825 $Y2=3.33
r52 33 48 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=2.99 $Y=3.33 $X2=3.6
+ $Y2=3.33
r53 33 35 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.99 $Y=3.33
+ $X2=2.825 $Y2=3.33
r54 29 32 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=2.825 $Y=2.105
+ $X2=2.825 $Y2=2.815
r55 27 35 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.825 $Y=3.245
+ $X2=2.825 $Y2=3.33
r56 27 32 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=2.825 $Y=3.245
+ $X2=2.825 $Y2=2.815
r57 24 26 9.26417 $w=9.33e-07 $l=7.1e-07 $layer=LI1_cond $X=1.612 $Y=2.105
+ $X2=1.612 $Y2=2.815
r58 21 42 17.6663 $w=9.14e-07 $l=3.35e-07 $layer=POLY_cond $X=1.915 $Y=0.712
+ $X2=2.25 $Y2=0.712
r59 21 39 49.5711 $w=9.14e-07 $l=9.4e-07 $layer=POLY_cond $X=1.915 $Y=0.712
+ $X2=0.975 $Y2=0.712
r60 20 24 9.00321 $w=9.33e-07 $l=6.9e-07 $layer=LI1_cond $X=1.612 $Y=1.415
+ $X2=1.612 $Y2=2.105
r61 20 21 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.915
+ $Y=1.415 $X2=1.915 $Y2=1.415
r62 18 55 3.4167 $w=9.35e-07 $l=8.5e-08 $layer=LI1_cond $X=1.612 $Y=3.245
+ $X2=1.612 $Y2=3.33
r63 18 26 5.6107 $w=9.33e-07 $l=4.3e-07 $layer=LI1_cond $X=1.612 $Y=3.245
+ $X2=1.612 $Y2=2.815
r64 17 52 4.78091 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=0.425 $Y=3.33
+ $X2=0.212 $Y2=3.33
r65 16 55 15.7884 $w=1.7e-07 $l=4.67e-07 $layer=LI1_cond $X=1.145 $Y=3.33
+ $X2=1.612 $Y2=3.33
r66 16 17 46.9733 $w=1.68e-07 $l=7.2e-07 $layer=LI1_cond $X=1.145 $Y=3.33
+ $X2=0.425 $Y2=3.33
r67 12 15 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=0.26 $Y=2.105
+ $X2=0.26 $Y2=2.815
r68 10 52 2.98526 $w=3.3e-07 $l=1.06325e-07 $layer=LI1_cond $X=0.26 $Y=3.245
+ $X2=0.212 $Y2=3.33
r69 10 15 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=0.26 $Y=3.245
+ $X2=0.26 $Y2=2.815
r70 1 32 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=2.685
+ $Y=1.96 $X2=2.825 $Y2=2.815
r71 1 29 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=2.685
+ $Y=1.96 $X2=2.825 $Y2=2.105
r72 1 26 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=1.41
+ $Y=1.96 $X2=1.55 $Y2=2.815
r73 1 24 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.41
+ $Y=1.96 $X2=1.55 $Y2=2.105
r74 1 15 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=1.41
+ $Y=1.96 $X2=0.26 $Y2=2.815
r75 1 12 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=1.41
+ $Y=1.96 $X2=0.26 $Y2=2.105
.ends

