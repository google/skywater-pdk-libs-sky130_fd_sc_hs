# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_hs__a222o_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__a222o_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.280000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.925000 1.350000 3.255000 2.150000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.685000 1.350000 5.155000 1.780000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.465000 1.350000 3.795000 1.780000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.965000 1.350000 4.445000 1.780000 ;
    END
  END B2
  PIN C1
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105000 1.300000 0.435000 1.780000 ;
    END
  END C1
  PIN C2
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605000 1.260000 1.140000 1.780000 ;
    END
  END C2
  PIN X
    ANTENNADIFFAREA  0.543200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.695000 0.920000 2.025000 1.820000 ;
        RECT 1.695000 1.820000 2.440000 2.200000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 5.280000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 5.280000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.280000 0.085000 ;
      RECT 0.000000  3.245000 5.280000 3.415000 ;
      RECT 0.115000  0.390000 0.365000 0.920000 ;
      RECT 0.115000  0.920000 1.525000 1.090000 ;
      RECT 0.115000  1.950000 1.525000 2.200000 ;
      RECT 0.115000  2.200000 0.365000 2.980000 ;
      RECT 0.565000  2.370000 4.165000 2.540000 ;
      RECT 0.565000  2.540000 0.895000 2.980000 ;
      RECT 0.935000  0.085000 1.185000 0.750000 ;
      RECT 1.355000  0.580000 2.400000 0.750000 ;
      RECT 1.355000  0.750000 1.525000 0.920000 ;
      RECT 1.355000  1.090000 1.525000 1.950000 ;
      RECT 1.575000  2.710000 1.905000 3.245000 ;
      RECT 2.205000  0.085000 2.535000 0.410000 ;
      RECT 2.230000  0.750000 2.400000 1.010000 ;
      RECT 2.230000  1.010000 3.750000 1.180000 ;
      RECT 2.230000  1.180000 2.560000 1.590000 ;
      RECT 2.645000  2.710000 2.975000 3.245000 ;
      RECT 2.765000  0.350000 4.090000 0.520000 ;
      RECT 2.765000  0.520000 3.095000 0.840000 ;
      RECT 3.265000  0.700000 3.750000 1.010000 ;
      RECT 3.265000  2.710000 3.630000 2.905000 ;
      RECT 3.265000  2.905000 4.665000 3.075000 ;
      RECT 3.835000  1.950000 4.165000 2.370000 ;
      RECT 3.835000  2.540000 4.165000 2.735000 ;
      RECT 3.920000  0.520000 4.090000 1.010000 ;
      RECT 3.920000  1.010000 5.140000 1.180000 ;
      RECT 4.260000  0.085000 4.590000 0.840000 ;
      RECT 4.335000  1.950000 4.665000 2.905000 ;
      RECT 4.810000  0.350000 5.140000 1.010000 ;
      RECT 4.835000  1.950000 5.165000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
  END
END sky130_fd_sc_hs__a222o_2
END LIBRARY
