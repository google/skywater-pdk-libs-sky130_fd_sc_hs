* File: sky130_fd_sc_hs__o22a_1.spice
* Created: Thu Aug 27 21:00:00 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hs__o22a_1.pex.spice"
.subckt sky130_fd_sc_hs__o22a_1  VNB VPB B1 B2 A2 A1 X VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* X	X
* A1	A1
* A2	A2
* B2	B2
* B1	B1
* VPB	VPB
* VNB	VNB
MM1009 N_VGND_M1009_d N_A_83_260#_M1009_g N_X_M1009_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.2109 PD=2.05 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1001 N_A_83_260#_M1001_d N_B1_M1001_g N_A_299_139#_M1001_s VNB NLOWVT L=0.15
+ W=0.64 AD=0.1024 AS=0.1705 PD=0.96 PS=1.85 NRD=3.744 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75001.7 A=0.096 P=1.58 MULT=1
MM1006 N_A_299_139#_M1006_d N_B2_M1006_g N_A_83_260#_M1001_d VNB NLOWVT L=0.15
+ W=0.64 AD=0.0896 AS=0.1024 PD=0.92 PS=0.96 NRD=0 NRS=3.744 M=1 R=4.26667
+ SA=75000.7 SB=75001.2 A=0.096 P=1.58 MULT=1
MM1004 N_VGND_M1004_d N_A2_M1004_g N_A_299_139#_M1006_d VNB NLOWVT L=0.15 W=0.64
+ AD=0.144737 AS=0.0896 PD=1.125 PS=0.92 NRD=15.936 NRS=0 M=1 R=4.26667
+ SA=75001.1 SB=75000.8 A=0.096 P=1.58 MULT=1
MM1000 N_A_299_139#_M1000_d N_A1_M1000_g N_VGND_M1004_d VNB NLOWVT L=0.15 W=0.64
+ AD=0.18205 AS=0.144737 PD=1.85 PS=1.125 NRD=0 NRS=14.052 M=1 R=4.26667
+ SA=75001.6 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1005 N_VPWR_M1005_d N_A_83_260#_M1005_g N_X_M1005_s VPB PSHORT L=0.15 W=1.12
+ AD=0.68246 AS=0.3304 PD=2.51472 PS=2.83 NRD=2.6201 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75002.7 A=0.168 P=2.54 MULT=1
MM1008 A_398_392# N_B1_M1008_g N_VPWR_M1005_d VPB PSHORT L=0.15 W=1 AD=0.135
+ AS=0.60934 PD=1.27 PS=2.24528 NRD=15.7403 NRS=2.9353 M=1 R=6.66667 SA=75001.6
+ SB=75001.6 A=0.15 P=2.3 MULT=1
MM1002 N_A_83_260#_M1002_d N_B2_M1002_g A_398_392# VPB PSHORT L=0.15 W=1 AD=0.15
+ AS=0.135 PD=1.3 PS=1.27 NRD=1.9503 NRS=15.7403 M=1 R=6.66667 SA=75002
+ SB=75001.2 A=0.15 P=2.3 MULT=1
MM1003 A_572_392# N_A2_M1003_g N_A_83_260#_M1002_d VPB PSHORT L=0.15 W=1
+ AD=0.195 AS=0.15 PD=1.39 PS=1.3 NRD=27.5603 NRS=1.9503 M=1 R=6.66667
+ SA=75002.5 SB=75000.8 A=0.15 P=2.3 MULT=1
MM1007 N_VPWR_M1007_d N_A1_M1007_g A_572_392# VPB PSHORT L=0.15 W=1 AD=0.295
+ AS=0.195 PD=2.59 PS=1.39 NRD=1.9503 NRS=27.5603 M=1 R=6.66667 SA=75003
+ SB=75000.2 A=0.15 P=2.3 MULT=1
DX10_noxref VNB VPB NWDIODE A=7.81875 P=12.19
c_346 A_398_392# 0 1.97013e-19 $X=1.99 $Y=1.96
*
.include "sky130_fd_sc_hs__o22a_1.pxi.spice"
*
.ends
*
*
