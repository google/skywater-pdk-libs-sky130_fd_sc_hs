* File: sky130_fd_sc_hs__inv_1.spice
* Created: Tue Sep  1 20:06:53 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hs__inv_1.pex.spice"
.subckt sky130_fd_sc_hs__inv_1  VNB VPB A VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A	A
* VPB	VPB
* VNB	VNB
MM1001 N_Y_M1001_d N_A_M1001_g N_VGND_M1001_s VNB NLOWVT L=0.15 W=0.74 AD=0.2109
+ AS=0.2627 PD=2.05 PS=2.19 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75000.3 SB=75000.2
+ A=0.111 P=1.78 MULT=1
MM1000 N_Y_M1000_d N_A_M1000_g N_VPWR_M1000_s VPB PSHORT L=0.15 W=1.12 AD=0.3304
+ AS=0.3864 PD=2.83 PS=2.93 NRD=1.7533 NRS=10.5395 M=1 R=7.46667 SA=75000.3
+ SB=75000.2 A=0.168 P=2.54 MULT=1
DX2_noxref VNB VPB NWDIODE A=3.3852 P=7.36
*
.include "sky130_fd_sc_hs__inv_1.pxi.spice"
*
.ends
*
*
