* File: sky130_fd_sc_hs__sdfxtp_2.pex.spice
* Created: Tue Sep  1 20:23:48 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HS__SDFXTP_2%A_27_74# 1 2 9 11 13 14 16 19 21 26 34 36
c82 36 0 6.89189e-20 $X=2.045 $Y=1.94
c83 34 0 1.9954e-19 $X=0.915 $Y=1.827
c84 14 0 1.79254e-19 $X=0.965 $Y=1.635
r85 36 39 5.5876 $w=3.28e-07 $l=1.6e-07 $layer=LI1_cond $X=2.045 $Y=1.94
+ $X2=2.045 $Y2=2.1
r86 36 37 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.045
+ $Y=1.94 $X2=2.045 $Y2=1.94
r87 32 34 10.9011 $w=7.13e-07 $l=1.65e-07 $layer=LI1_cond $X=0.75 $Y=1.827
+ $X2=0.915 $Y2=1.827
r88 32 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.75
+ $Y=1.635 $X2=0.75 $Y2=1.635
r89 30 32 8.11326 $w=7.13e-07 $l=4.85e-07 $layer=LI1_cond $X=0.265 $Y=1.827
+ $X2=0.75 $Y2=1.827
r90 23 26 5.9927 $w=2.48e-07 $l=1.3e-07 $layer=LI1_cond $X=0.17 $Y=0.515 $X2=0.3
+ $Y2=0.515
r91 21 39 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.88 $Y=2.1
+ $X2=2.045 $Y2=2.1
r92 21 34 62.9572 $w=1.68e-07 $l=9.65e-07 $layer=LI1_cond $X=1.88 $Y=2.1
+ $X2=0.915 $Y2=2.1
r93 17 30 4.75969 $w=3.6e-07 $l=3.58e-07 $layer=LI1_cond $X=0.265 $Y=2.185
+ $X2=0.265 $Y2=1.827
r94 17 19 7.20277 $w=3.58e-07 $l=2.25e-07 $layer=LI1_cond $X=0.265 $Y=2.185
+ $X2=0.265 $Y2=2.41
r95 16 30 1.5892 $w=7.13e-07 $l=9.5e-08 $layer=LI1_cond $X=0.17 $Y=1.827
+ $X2=0.265 $Y2=1.827
r96 15 23 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.17 $Y=0.64
+ $X2=0.17 $Y2=0.515
r97 15 16 54.1497 $w=1.68e-07 $l=8.3e-07 $layer=LI1_cond $X=0.17 $Y=0.64
+ $X2=0.17 $Y2=1.47
r98 14 33 37.5952 $w=3.3e-07 $l=2.15e-07 $layer=POLY_cond $X=0.965 $Y=1.635
+ $X2=0.75 $Y2=1.635
r99 11 37 52.2586 $w=2.99e-07 $l=2.85044e-07 $layer=POLY_cond $X=2.12 $Y=2.19
+ $X2=2.045 $Y2=1.94
r100 11 13 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=2.12 $Y=2.19
+ $X2=2.12 $Y2=2.585
r101 7 14 32.1775 $w=3.3e-07 $l=1.98997e-07 $layer=POLY_cond $X=1.04 $Y=1.47
+ $X2=0.965 $Y2=1.635
r102 7 9 456.362 $w=1.5e-07 $l=8.9e-07 $layer=POLY_cond $X=1.04 $Y=1.47 $X2=1.04
+ $Y2=0.58
r103 2 19 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=2.265 $X2=0.28 $Y2=2.41
r104 1 26 182 $w=1.7e-07 $l=2.5446e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.37 $X2=0.3 $Y2=0.555
.ends

.subckt PM_SKY130_FD_SC_HS__SDFXTP_2%SCE 2 3 5 6 8 9 10 11 13 14 16 20 22 28 31
+ 37 43
c83 37 0 1.36067e-19 $X=2.135 $Y=1.065
c84 31 0 3.45016e-20 $X=0.54 $Y=1.065
c85 22 0 4.92605e-20 $X=2.04 $Y=0.935
c86 9 0 3.61584e-20 $X=0.93 $Y=2.115
r87 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.59
+ $Y=1.065 $X2=0.59 $Y2=1.065
r88 31 33 9.41406 $w=2.56e-07 $l=5e-08 $layer=POLY_cond $X=0.54 $Y=1.065
+ $X2=0.59 $Y2=1.065
r89 28 43 7.36464 $w=4.18e-07 $l=1.15e-07 $layer=LI1_cond $X=0.72 $Y=1.02
+ $X2=0.835 $Y2=1.02
r90 28 34 3.56709 $w=4.18e-07 $l=1.3e-07 $layer=LI1_cond $X=0.72 $Y=1.02
+ $X2=0.59 $Y2=1.02
r91 26 37 16.6118 $w=3.3e-07 $l=9.5e-08 $layer=POLY_cond $X=2.04 $Y=1.065
+ $X2=2.135 $Y2=1.065
r92 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.04
+ $Y=1.065 $X2=2.04 $Y2=1.065
r93 22 25 4.53993 $w=3.28e-07 $l=1.3e-07 $layer=LI1_cond $X=2.04 $Y=0.935
+ $X2=2.04 $Y2=1.065
r94 20 22 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.875 $Y=0.935
+ $X2=2.04 $Y2=0.935
r95 20 43 67.8503 $w=1.68e-07 $l=1.04e-06 $layer=LI1_cond $X=1.875 $Y=0.935
+ $X2=0.835 $Y2=0.935
r96 17 19 120.5 $w=1.5e-07 $l=2.35e-07 $layer=POLY_cond $X=0.27 $Y=2.115
+ $X2=0.505 $Y2=2.115
r97 14 37 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.135 $Y=0.9
+ $X2=2.135 $Y2=1.065
r98 14 16 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.135 $Y=0.9
+ $X2=2.135 $Y2=0.58
r99 11 13 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=1.005 $Y=2.19
+ $X2=1.005 $Y2=2.585
r100 10 19 38.4574 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.58 $Y=2.115
+ $X2=0.505 $Y2=2.115
r101 9 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.93 $Y=2.115
+ $X2=1.005 $Y2=2.19
r102 9 10 179.468 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=0.93 $Y=2.115
+ $X2=0.58 $Y2=2.115
r103 6 31 15.2686 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.54 $Y=0.9
+ $X2=0.54 $Y2=1.065
r104 6 8 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.54 $Y=0.9 $X2=0.54
+ $Y2=0.58
r105 3 19 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.505 $Y=2.19
+ $X2=0.505 $Y2=2.115
r106 3 5 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=0.505 $Y=2.19
+ $X2=0.505 $Y2=2.585
r107 2 17 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.27 $Y=2.04
+ $X2=0.27 $Y2=2.115
r108 1 31 50.8359 $w=2.56e-07 $l=3.4271e-07 $layer=POLY_cond $X=0.27 $Y=1.23
+ $X2=0.54 $Y2=1.065
r109 1 2 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=0.27 $Y=1.23 $X2=0.27
+ $Y2=2.04
.ends

.subckt PM_SKY130_FD_SC_HS__SDFXTP_2%D 2 3 5 8 12 13 14 17 18
c46 18 0 2.06727e-19 $X=1.5 $Y=1.355
c47 17 0 4.92605e-20 $X=1.5 $Y=1.355
c48 12 0 1.9954e-19 $X=1.5 $Y=1.695
c49 3 0 2.16829e-19 $X=1.425 $Y=2.19
r50 17 18 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.5
+ $Y=1.355 $X2=1.5 $Y2=1.355
r51 14 18 5.47822 $w=6.53e-07 $l=3e-07 $layer=LI1_cond $X=1.2 $Y=1.517 $X2=1.5
+ $Y2=1.517
r52 12 17 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.5 $Y=1.695 $X2=1.5
+ $Y2=1.355
r53 12 13 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.5 $Y=1.695
+ $X2=1.5 $Y2=1.86
r54 11 17 43.0552 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.5 $Y=1.19 $X2=1.5
+ $Y2=1.355
r55 8 11 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.43 $Y=0.58 $X2=1.43
+ $Y2=1.19
r56 3 5 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=1.425 $Y=2.19
+ $X2=1.425 $Y2=2.585
r57 2 3 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=1.425 $Y=2.1 $X2=1.425
+ $Y2=2.19
r58 2 13 93.2903 $w=1.8e-07 $l=2.4e-07 $layer=POLY_cond $X=1.425 $Y=2.1
+ $X2=1.425 $Y2=1.86
.ends

.subckt PM_SKY130_FD_SC_HS__SDFXTP_2%SCD 3 5 7 10 11 12 16
r43 11 12 15.1913 $w=3.28e-07 $l=4.35e-07 $layer=LI1_cond $X=2.615 $Y=1.6
+ $X2=2.615 $Y2=2.035
r44 11 16 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.615
+ $Y=1.6 $X2=2.615 $Y2=1.6
r45 10 16 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.615 $Y=1.94
+ $X2=2.615 $Y2=1.6
r46 9 16 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.615 $Y=1.435
+ $X2=2.615 $Y2=1.6
r47 5 10 43.19 $w=2.79e-07 $l=2.85044e-07 $layer=POLY_cond $X=2.54 $Y=2.19
+ $X2=2.615 $Y2=1.94
r48 5 7 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=2.54 $Y=2.19 $X2=2.54
+ $Y2=2.585
r49 3 9 438.415 $w=1.5e-07 $l=8.55e-07 $layer=POLY_cond $X=2.525 $Y=0.58
+ $X2=2.525 $Y2=1.435
.ends

.subckt PM_SKY130_FD_SC_HS__SDFXTP_2%CLK 3 5 7 8 11 14
c46 11 0 1.00538e-19 $X=3.28 $Y=1.557
r47 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.455
+ $Y=1.515 $X2=3.455 $Y2=1.515
r48 11 13 23.7606 $w=3.55e-07 $l=1.75e-07 $layer=POLY_cond $X=3.28 $Y=1.557
+ $X2=3.455 $Y2=1.557
r49 10 11 25.1183 $w=3.55e-07 $l=1.85e-07 $layer=POLY_cond $X=3.095 $Y=1.557
+ $X2=3.28 $Y2=1.557
r50 8 14 4.37637 $w=3.93e-07 $l=1.5e-07 $layer=LI1_cond $X=3.487 $Y=1.665
+ $X2=3.487 $Y2=1.515
r51 5 11 22.9692 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=3.28 $Y=1.765
+ $X2=3.28 $Y2=1.557
r52 5 7 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.28 $Y=1.765
+ $X2=3.28 $Y2=2.4
r53 1 10 22.9692 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.095 $Y=1.35
+ $X2=3.095 $Y2=1.557
r54 1 3 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=3.095 $Y=1.35
+ $X2=3.095 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HS__SDFXTP_2%A_846_74# 1 2 7 9 12 15 16 18 20 24 26 27
+ 29 30 33 36 37 39 42 43 44 46 48 52 53 55 56 61 62 67 73 76
c191 67 0 1.91717e-19 $X=8.58 $Y=2.155
c192 61 0 1.80614e-19 $X=8.26 $Y=1.195
c193 53 0 5.96821e-20 $X=5.21 $Y=1.775
c194 52 0 1.28501e-19 $X=5.21 $Y=1.775
c195 36 0 1.59795e-19 $X=6.11 $Y=1.195
c196 20 0 1.74027e-19 $X=5.21 $Y=2.13
r197 67 68 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.58
+ $Y=2.155 $X2=8.58 $Y2=2.155
r198 64 67 7.33373 $w=3.28e-07 $l=2.1e-07 $layer=LI1_cond $X=8.37 $Y=2.155
+ $X2=8.58 $Y2=2.155
r199 61 76 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=8.26 $Y=1.195
+ $X2=8.26 $Y2=1.03
r200 60 62 3.84148 $w=3.28e-07 $l=1.1e-07 $layer=LI1_cond $X=8.26 $Y=1.195
+ $X2=8.37 $Y2=1.195
r201 60 61 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.26
+ $Y=1.195 $X2=8.26 $Y2=1.195
r202 57 60 4.01609 $w=3.28e-07 $l=1.15e-07 $layer=LI1_cond $X=8.145 $Y=1.195
+ $X2=8.26 $Y2=1.195
r203 52 54 1.31655 $w=5.56e-07 $l=6e-08 $layer=LI1_cond $X=5.21 $Y=1.945
+ $X2=5.27 $Y2=1.945
r204 52 53 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.21
+ $Y=1.775 $X2=5.21 $Y2=1.775
r205 50 52 10.3129 $w=5.56e-07 $l=4.7e-07 $layer=LI1_cond $X=4.74 $Y=1.945
+ $X2=5.21 $Y2=1.945
r206 48 64 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.37 $Y=1.99
+ $X2=8.37 $Y2=2.155
r207 47 62 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.37 $Y=1.36
+ $X2=8.37 $Y2=1.195
r208 47 48 41.1016 $w=1.68e-07 $l=6.3e-07 $layer=LI1_cond $X=8.37 $Y=1.36
+ $X2=8.37 $Y2=1.99
r209 46 57 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.145 $Y=1.03
+ $X2=8.145 $Y2=1.195
r210 45 46 39.4706 $w=1.68e-07 $l=6.05e-07 $layer=LI1_cond $X=8.145 $Y=0.425
+ $X2=8.145 $Y2=1.03
r211 43 45 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.06 $Y=0.34
+ $X2=8.145 $Y2=0.425
r212 43 44 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=8.06 $Y=0.34
+ $X2=7.39 $Y2=0.34
r213 41 44 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.305 $Y=0.425
+ $X2=7.39 $Y2=0.34
r214 41 42 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=7.305 $Y=0.425
+ $X2=7.305 $Y2=0.72
r215 40 56 2.76166 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.275 $Y=0.805
+ $X2=6.11 $Y2=0.805
r216 39 42 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.22 $Y=0.805
+ $X2=7.305 $Y2=0.72
r217 39 40 61.6524 $w=1.68e-07 $l=9.45e-07 $layer=LI1_cond $X=7.22 $Y=0.805
+ $X2=6.275 $Y2=0.805
r218 37 73 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.11 $Y=1.195
+ $X2=6.11 $Y2=1.03
r219 36 37 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.11
+ $Y=1.195 $X2=6.11 $Y2=1.195
r220 34 56 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.11 $Y=0.89
+ $X2=6.11 $Y2=0.805
r221 34 36 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=6.11 $Y=0.89
+ $X2=6.11 $Y2=1.195
r222 33 56 3.70735 $w=2.5e-07 $l=1.18427e-07 $layer=LI1_cond $X=6.03 $Y=0.72
+ $X2=6.11 $Y2=0.805
r223 32 33 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=6.03 $Y=0.425
+ $X2=6.03 $Y2=0.72
r224 31 55 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.355 $Y=0.34
+ $X2=5.27 $Y2=0.34
r225 30 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.945 $Y=0.34
+ $X2=6.03 $Y2=0.425
r226 30 31 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=5.945 $Y=0.34
+ $X2=5.355 $Y2=0.34
r227 29 54 7.82841 $w=1.7e-07 $l=3.35e-07 $layer=LI1_cond $X=5.27 $Y=1.61
+ $X2=5.27 $Y2=1.945
r228 28 55 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.27 $Y=0.425
+ $X2=5.27 $Y2=0.34
r229 28 29 77.3102 $w=1.68e-07 $l=1.185e-06 $layer=LI1_cond $X=5.27 $Y=0.425
+ $X2=5.27 $Y2=1.61
r230 26 55 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.185 $Y=0.34
+ $X2=5.27 $Y2=0.34
r231 26 27 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=5.185 $Y=0.34
+ $X2=4.535 $Y2=0.34
r232 22 27 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.37 $Y=0.425
+ $X2=4.535 $Y2=0.34
r233 22 24 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=4.37 $Y=0.425
+ $X2=4.37 $Y2=0.515
r234 20 53 62.0758 $w=3.3e-07 $l=3.55e-07 $layer=POLY_cond $X=5.21 $Y=2.13
+ $X2=5.21 $Y2=1.775
r235 20 21 72.9952 $w=2.08e-07 $l=3.15e-07 $layer=POLY_cond $X=5.21 $Y=2.28
+ $X2=5.525 $Y2=2.28
r236 16 68 50.5804 $w=3.46e-07 $l=2.97909e-07 $layer=POLY_cond $X=8.445 $Y=2.405
+ $X2=8.55 $Y2=2.155
r237 16 18 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=8.445 $Y=2.405
+ $X2=8.445 $Y2=2.69
r238 15 76 123.713 $w=1.5e-07 $l=3.85e-07 $layer=POLY_cond $X=8.35 $Y=0.645
+ $X2=8.35 $Y2=1.03
r239 12 73 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=6.02 $Y=0.71
+ $X2=6.02 $Y2=1.03
r240 7 21 10.4806 $w=1.5e-07 $l=1.85e-07 $layer=POLY_cond $X=5.525 $Y=2.465
+ $X2=5.525 $Y2=2.28
r241 7 9 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=5.525 $Y=2.465
+ $X2=5.525 $Y2=2.75
r242 2 50 600 $w=1.7e-07 $l=2.74955e-07 $layer=licon1_PDIFF $count=1 $X=4.59
+ $Y=1.84 $X2=4.74 $Y2=2.05
r243 1 24 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=4.23
+ $Y=0.37 $X2=4.37 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__SDFXTP_2%A_634_74# 1 2 7 9 10 12 13 14 17 19 22 23
+ 24 25 27 28 30 31 35 37 42 44 46 50 52 55 57 60 61 62 64 68 76
c214 76 0 7.36295e-20 $X=7.95 $Y=1.765
c215 68 0 1.74027e-19 $X=6.06 $Y=2.135
c216 57 0 1.10031e-19 $X=7.005 $Y=2.215
c217 52 0 1.00538e-19 $X=4 $Y=1.445
c218 35 0 1.57288e-19 $X=8.86 $Y=0.58
c219 19 0 2.88296e-19 $X=5.585 $Y=1.295
r220 80 81 39.3469 $w=4.41e-07 $l=3.6e-07 $layer=POLY_cond $X=4.155 $Y=1.492
+ $X2=4.515 $Y2=1.492
r221 77 83 14.9072 $w=2.91e-07 $l=9e-08 $layer=POLY_cond $X=7.95 $Y=1.765
+ $X2=7.95 $Y2=1.675
r222 76 77 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.95
+ $Y=1.765 $X2=7.95 $Y2=1.765
r223 73 76 6.28605 $w=3.28e-07 $l=1.8e-07 $layer=LI1_cond $X=7.77 $Y=1.765
+ $X2=7.95 $Y2=1.765
r224 68 71 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=6.06 $Y=2.135 $X2=6.06
+ $Y2=2.215
r225 68 69 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.06
+ $Y=2.135 $X2=6.06 $Y2=2.135
r226 63 73 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.77 $Y=1.93
+ $X2=7.77 $Y2=1.765
r227 63 64 63.6096 $w=1.68e-07 $l=9.75e-07 $layer=LI1_cond $X=7.77 $Y=1.93
+ $X2=7.77 $Y2=2.905
r228 61 64 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.685 $Y=2.99
+ $X2=7.77 $Y2=2.905
r229 61 62 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=7.685 $Y=2.99
+ $X2=7.175 $Y2=2.99
r230 60 62 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.09 $Y=2.905
+ $X2=7.175 $Y2=2.99
r231 59 60 39.4706 $w=1.68e-07 $l=6.05e-07 $layer=LI1_cond $X=7.09 $Y=2.3
+ $X2=7.09 $Y2=2.905
r232 58 71 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.225 $Y=2.215
+ $X2=6.06 $Y2=2.215
r233 57 59 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.005 $Y=2.215
+ $X2=7.09 $Y2=2.3
r234 57 58 50.8877 $w=1.68e-07 $l=7.8e-07 $layer=LI1_cond $X=7.005 $Y=2.215
+ $X2=6.225 $Y2=2.215
r235 56 80 16.941 $w=4.41e-07 $l=1.55e-07 $layer=POLY_cond $X=4 $Y=1.492
+ $X2=4.155 $Y2=1.492
r236 55 56 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4
+ $Y=1.465 $X2=4 $Y2=1.465
r237 53 55 19.2736 $w=2.88e-07 $l=4.85e-07 $layer=LI1_cond $X=4 $Y=1.95 $X2=4
+ $Y2=1.465
r238 52 66 15.6734 $w=2.9e-07 $l=3.5e-07 $layer=LI1_cond $X=4 $Y=1.445 $X2=4
+ $Y2=1.095
r239 52 55 0.794788 $w=2.88e-07 $l=2e-08 $layer=LI1_cond $X=4 $Y=1.445 $X2=4
+ $Y2=1.465
r240 51 65 2.55969 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.475 $Y=1.095
+ $X2=3.31 $Y2=1.095
r241 50 66 1.9771 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=3.855 $Y=1.095 $X2=4
+ $Y2=1.095
r242 50 51 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=3.855 $Y=1.095
+ $X2=3.475 $Y2=1.095
r243 46 53 6.85346 $w=3.3e-07 $l=2.26164e-07 $layer=LI1_cond $X=3.855 $Y=2.115
+ $X2=4 $Y2=1.95
r244 46 48 12.2229 $w=3.28e-07 $l=3.5e-07 $layer=LI1_cond $X=3.855 $Y=2.115
+ $X2=3.505 $Y2=2.115
r245 42 65 13.6603 $w=3.3e-07 $l=3.4e-07 $layer=LI1_cond $X=3.31 $Y=0.755
+ $X2=3.31 $Y2=1.095
r246 42 44 9.07985 $w=3.28e-07 $l=2.6e-07 $layer=LI1_cond $X=3.31 $Y=0.755
+ $X2=3.31 $Y2=0.495
r247 33 35 523.021 $w=1.5e-07 $l=1.02e-06 $layer=POLY_cond $X=8.86 $Y=1.6
+ $X2=8.86 $Y2=0.58
r248 32 83 18.2534 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.115 $Y=1.675
+ $X2=7.95 $Y2=1.675
r249 31 33 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=8.785 $Y=1.675
+ $X2=8.86 $Y2=1.6
r250 31 32 343.553 $w=1.5e-07 $l=6.7e-07 $layer=POLY_cond $X=8.785 $Y=1.675
+ $X2=8.115 $Y2=1.675
r251 28 77 57.6553 $w=2.91e-07 $l=3.10805e-07 $layer=POLY_cond $X=7.885 $Y=2.045
+ $X2=7.95 $Y2=1.765
r252 28 30 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=7.885 $Y=2.045
+ $X2=7.885 $Y2=2.54
r253 25 69 69.5873 $w=2.61e-07 $l=3.67831e-07 $layer=POLY_cond $X=5.975 $Y=2.465
+ $X2=6.055 $Y2=2.135
r254 25 27 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=5.975 $Y=2.465
+ $X2=5.975 $Y2=2.75
r255 24 69 3.43315 $w=3.4e-07 $l=5e-09 $layer=POLY_cond $X=6.055 $Y=2.13
+ $X2=6.055 $Y2=2.135
r256 23 38 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=6.055 $Y=1.815
+ $X2=5.66 $Y2=1.815
r257 23 24 40.7324 $w=3.4e-07 $l=2.4e-07 $layer=POLY_cond $X=6.055 $Y=1.89
+ $X2=6.055 $Y2=2.13
r258 22 38 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.66 $Y=1.74
+ $X2=5.66 $Y2=1.815
r259 21 22 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=5.66 $Y=1.37
+ $X2=5.66 $Y2=1.74
r260 20 37 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.22 $Y=1.295
+ $X2=5.145 $Y2=1.295
r261 19 21 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.585 $Y=1.295
+ $X2=5.66 $Y2=1.37
r262 19 20 187.16 $w=1.5e-07 $l=3.65e-07 $layer=POLY_cond $X=5.585 $Y=1.295
+ $X2=5.22 $Y2=1.295
r263 15 37 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.145 $Y=1.22
+ $X2=5.145 $Y2=1.295
r264 15 17 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=5.145 $Y=1.22
+ $X2=5.145 $Y2=0.71
r265 14 81 32.2719 $w=4.41e-07 $l=2.37779e-07 $layer=POLY_cond $X=4.605 $Y=1.295
+ $X2=4.515 $Y2=1.492
r266 13 37 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.07 $Y=1.295
+ $X2=5.145 $Y2=1.295
r267 13 14 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=5.07 $Y=1.295
+ $X2=4.605 $Y2=1.295
r268 10 81 28.2648 $w=1.5e-07 $l=2.73e-07 $layer=POLY_cond $X=4.515 $Y=1.765
+ $X2=4.515 $Y2=1.492
r269 10 12 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=4.515 $Y=1.765
+ $X2=4.515 $Y2=2.4
r270 7 80 28.2648 $w=1.5e-07 $l=2.72e-07 $layer=POLY_cond $X=4.155 $Y=1.22
+ $X2=4.155 $Y2=1.492
r271 7 9 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=4.155 $Y=1.22
+ $X2=4.155 $Y2=0.74
r272 2 48 600 $w=1.7e-07 $l=3.4187e-07 $layer=licon1_PDIFF $count=1 $X=3.355
+ $Y=1.84 $X2=3.505 $Y2=2.115
r273 1 44 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=3.17
+ $Y=0.37 $X2=3.31 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_HS__SDFXTP_2%A_1287_320# 1 2 8 9 11 16 18 19 21 22 25 29
+ 33 35
c85 33 0 1.06984e-19 $X=7.725 $Y=0.765
c86 19 0 1.86347e-19 $X=6.535 $Y=1.75
r87 31 35 6.46576 $w=2.5e-07 $l=3.8e-07 $layer=LI1_cond $X=7.725 $Y=1.06
+ $X2=7.345 $Y2=1.06
r88 31 33 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=7.725 $Y=1.06
+ $X2=7.725 $Y2=0.765
r89 27 35 6.46576 $w=2.5e-07 $l=3.70068e-07 $layer=LI1_cond $X=7.43 $Y=1.39
+ $X2=7.345 $Y2=1.06
r90 27 29 66.5455 $w=1.68e-07 $l=1.02e-06 $layer=LI1_cond $X=7.43 $Y=1.39
+ $X2=7.43 $Y2=2.41
r91 24 25 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.99
+ $Y=1.225 $X2=6.99 $Y2=1.225
r92 22 35 0.364692 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=7.345 $Y=1.225
+ $X2=7.345 $Y2=1.06
r93 22 24 12.3975 $w=3.28e-07 $l=3.55e-07 $layer=LI1_cond $X=7.345 $Y=1.225
+ $X2=6.99 $Y2=1.225
r94 20 25 56.8299 $w=3.3e-07 $l=3.25e-07 $layer=POLY_cond $X=6.665 $Y=1.225
+ $X2=6.99 $Y2=1.225
r95 20 21 5.03009 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=6.665 $Y=1.225
+ $X2=6.575 $Y2=1.225
r96 18 19 60.4563 $w=1.8e-07 $l=1.5e-07 $layer=POLY_cond $X=6.535 $Y=1.6
+ $X2=6.535 $Y2=1.75
r97 14 21 37.0704 $w=1.5e-07 $l=1.72337e-07 $layer=POLY_cond $X=6.59 $Y=1.06
+ $X2=6.575 $Y2=1.225
r98 14 16 179.468 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=6.59 $Y=1.06
+ $X2=6.59 $Y2=0.71
r99 12 21 37.0704 $w=1.5e-07 $l=1.72337e-07 $layer=POLY_cond $X=6.56 $Y=1.39
+ $X2=6.575 $Y2=1.225
r100 12 18 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=6.56 $Y=1.39
+ $X2=6.56 $Y2=1.6
r101 9 11 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=6.525 $Y=2.465
+ $X2=6.525 $Y2=2.75
r102 8 9 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=6.525 $Y=2.375
+ $X2=6.525 $Y2=2.465
r103 8 19 242.944 $w=1.8e-07 $l=6.25e-07 $layer=POLY_cond $X=6.525 $Y=2.375
+ $X2=6.525 $Y2=1.75
r104 2 29 600 $w=1.7e-07 $l=3.57211e-07 $layer=licon1_PDIFF $count=1 $X=7.28
+ $Y=2.12 $X2=7.43 $Y2=2.41
r105 1 33 182 $w=1.7e-07 $l=4.59701e-07 $layer=licon1_NDIFF $count=1 $X=7.585
+ $Y=0.37 $X2=7.725 $Y2=0.765
.ends

.subckt PM_SKY130_FD_SC_HS__SDFXTP_2%A_1044_100# 1 2 7 9 11 14 15 16 18 21 24 27
+ 29 30 32 39
c105 32 0 7.63155e-20 $X=7.01 $Y=1.715
c106 27 0 1.87953e-19 $X=5.665 $Y=1.715
c107 18 0 5.96821e-20 $X=5.665 $Y=1.63
r108 39 40 36.3903 $w=3.51e-07 $l=2.65e-07 $layer=POLY_cond $X=7.205 $Y=1.837
+ $X2=7.47 $Y2=1.837
r109 36 39 26.7778 $w=3.51e-07 $l=1.95e-07 $layer=POLY_cond $X=7.01 $Y=1.837
+ $X2=7.205 $Y2=1.837
r110 35 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.01
+ $Y=1.795 $X2=7.01 $Y2=1.795
r111 32 35 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=7.01 $Y=1.715 $X2=7.01
+ $Y2=1.795
r112 29 30 10.5918 $w=3.58e-07 $l=2.3e-07 $layer=LI1_cond $X=5.735 $Y=2.75
+ $X2=5.735 $Y2=2.52
r113 24 26 8.26222 $w=2.48e-07 $l=1.75e-07 $layer=LI1_cond $X=5.65 $Y=0.765
+ $X2=5.65 $Y2=0.94
r114 22 27 1.84097 $w=1.7e-07 $l=1.1e-07 $layer=LI1_cond $X=5.775 $Y=1.715
+ $X2=5.665 $Y2=1.715
r115 21 32 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.845 $Y=1.715
+ $X2=7.01 $Y2=1.715
r116 21 22 69.8075 $w=1.68e-07 $l=1.07e-06 $layer=LI1_cond $X=6.845 $Y=1.715
+ $X2=5.775 $Y2=1.715
r117 19 27 4.60183 $w=1.95e-07 $l=9.66954e-08 $layer=LI1_cond $X=5.64 $Y=1.8
+ $X2=5.665 $Y2=1.715
r118 19 30 46.9733 $w=1.68e-07 $l=7.2e-07 $layer=LI1_cond $X=5.64 $Y=1.8
+ $X2=5.64 $Y2=2.52
r119 18 27 4.60183 $w=1.95e-07 $l=8.5e-08 $layer=LI1_cond $X=5.665 $Y=1.63
+ $X2=5.665 $Y2=1.715
r120 18 26 36.1448 $w=2.18e-07 $l=6.9e-07 $layer=LI1_cond $X=5.665 $Y=1.63
+ $X2=5.665 $Y2=0.94
r121 15 16 53.9552 $w=1.9e-07 $l=1.5e-07 $layer=POLY_cond $X=7.49 $Y=0.995
+ $X2=7.49 $Y2=1.145
r122 14 15 112.467 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=7.51 $Y=0.645
+ $X2=7.51 $Y2=0.995
r123 11 40 22.6971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=7.47 $Y=1.63
+ $X2=7.47 $Y2=1.837
r124 11 16 248.691 $w=1.5e-07 $l=4.85e-07 $layer=POLY_cond $X=7.47 $Y=1.63
+ $X2=7.47 $Y2=1.145
r125 7 39 22.6971 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=7.205 $Y=2.045
+ $X2=7.205 $Y2=1.837
r126 7 9 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=7.205 $Y=2.045
+ $X2=7.205 $Y2=2.54
r127 2 29 600 $w=1.7e-07 $l=2.74955e-07 $layer=licon1_PDIFF $count=1 $X=5.6
+ $Y=2.54 $X2=5.75 $Y2=2.75
r128 1 24 182 $w=1.7e-07 $l=5.05421e-07 $layer=licon1_NDIFF $count=1 $X=5.22
+ $Y=0.5 $X2=5.61 $Y2=0.765
.ends

.subckt PM_SKY130_FD_SC_HS__SDFXTP_2%A_1829_398# 1 2 7 8 9 11 14 16 18 19 21 22
+ 24 25 27 28 31 35 38 39 42 46 48 54 55
c103 39 0 1.57288e-19 $X=9.535 $Y=1.155
c104 28 0 1.40987e-19 $X=10.93 $Y=1.385
c105 19 0 1.10546e-19 $X=11.045 $Y=1.765
c106 14 0 1.58278e-19 $X=9.25 $Y=0.58
c107 8 0 2.29134e-20 $X=9.235 $Y=2.315
c108 7 0 1.68803e-19 $X=9.235 $Y=2.08
r109 54 55 11.2873 $w=3.48e-07 $l=2.5e-07 $layer=LI1_cond $X=10.27 $Y=2.665
+ $X2=10.27 $Y2=2.415
r110 48 49 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=10.88
+ $Y=1.385 $X2=10.88 $Y2=1.385
r111 46 52 3.87119 $w=3.3e-07 $l=1.8262e-07 $layer=LI1_cond $X=10.445 $Y=1.385
+ $X2=10.36 $Y2=1.24
r112 46 48 15.1913 $w=3.28e-07 $l=4.35e-07 $layer=LI1_cond $X=10.445 $Y=1.385
+ $X2=10.88 $Y2=1.385
r113 44 52 3.01842 $w=1.7e-07 $l=3.1e-07 $layer=LI1_cond $X=10.36 $Y=1.55
+ $X2=10.36 $Y2=1.24
r114 44 55 56.4332 $w=1.68e-07 $l=8.65e-07 $layer=LI1_cond $X=10.36 $Y=1.55
+ $X2=10.36 $Y2=2.415
r115 40 52 19.1992 $w=2.51e-07 $l=3.95e-07 $layer=LI1_cond $X=9.965 $Y=1.24
+ $X2=10.36 $Y2=1.24
r116 40 42 19.382 $w=3.28e-07 $l=5.55e-07 $layer=LI1_cond $X=9.965 $Y=1.07
+ $X2=9.965 $Y2=0.515
r117 38 40 9.29704 $w=2.51e-07 $l=2.03101e-07 $layer=LI1_cond $X=9.8 $Y=1.155
+ $X2=9.965 $Y2=1.24
r118 38 39 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=9.8 $Y=1.155
+ $X2=9.535 $Y2=1.155
r119 35 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.37
+ $Y=1.74 $X2=9.37 $Y2=1.74
r120 33 39 7.55824 $w=1.7e-07 $l=1.90825e-07 $layer=LI1_cond $X=9.382 $Y=1.24
+ $X2=9.535 $Y2=1.155
r121 33 35 18.8925 $w=3.03e-07 $l=5e-07 $layer=LI1_cond $X=9.382 $Y=1.24
+ $X2=9.382 $Y2=1.74
r122 31 32 1.61384 $w=4.48e-07 $l=1.5e-08 $layer=POLY_cond $X=11.48 $Y=1.492
+ $X2=11.495 $Y2=1.492
r123 30 31 46.8013 $w=4.48e-07 $l=4.35e-07 $layer=POLY_cond $X=11.045 $Y=1.492
+ $X2=11.48 $Y2=1.492
r124 29 30 4.30357 $w=4.48e-07 $l=4e-08 $layer=POLY_cond $X=11.005 $Y=1.492
+ $X2=11.045 $Y2=1.492
r125 28 49 8.74306 $w=3.3e-07 $l=5e-08 $layer=POLY_cond $X=10.93 $Y=1.385
+ $X2=10.88 $Y2=1.385
r126 28 29 11.5087 $w=4.48e-07 $l=1.39549e-07 $layer=POLY_cond $X=10.93 $Y=1.385
+ $X2=11.005 $Y2=1.492
r127 25 32 28.6558 $w=1.5e-07 $l=2.73e-07 $layer=POLY_cond $X=11.495 $Y=1.765
+ $X2=11.495 $Y2=1.492
r128 25 27 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=11.495 $Y=1.765
+ $X2=11.495 $Y2=2.4
r129 22 31 28.6558 $w=1.5e-07 $l=2.72e-07 $layer=POLY_cond $X=11.48 $Y=1.22
+ $X2=11.48 $Y2=1.492
r130 22 24 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=11.48 $Y=1.22
+ $X2=11.48 $Y2=0.74
r131 19 30 28.6558 $w=1.5e-07 $l=2.73e-07 $layer=POLY_cond $X=11.045 $Y=1.765
+ $X2=11.045 $Y2=1.492
r132 19 21 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=11.045 $Y=1.765
+ $X2=11.045 $Y2=2.4
r133 16 29 28.6558 $w=1.5e-07 $l=2.72e-07 $layer=POLY_cond $X=11.005 $Y=1.22
+ $X2=11.005 $Y2=1.492
r134 16 18 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=11.005 $Y=1.22
+ $X2=11.005 $Y2=0.74
r135 12 36 38.5991 $w=2.92e-07 $l=2.05122e-07 $layer=POLY_cond $X=9.25 $Y=1.575
+ $X2=9.34 $Y2=1.74
r136 12 14 510.202 $w=1.5e-07 $l=9.95e-07 $layer=POLY_cond $X=9.25 $Y=1.575
+ $X2=9.25 $Y2=0.58
r137 9 11 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=9.235 $Y=2.405
+ $X2=9.235 $Y2=2.69
r138 8 9 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=9.235 $Y=2.315
+ $X2=9.235 $Y2=2.405
r139 7 36 63.1688 $w=2.92e-07 $l=3.88973e-07 $layer=POLY_cond $X=9.235 $Y=2.08
+ $X2=9.34 $Y2=1.74
r140 7 8 91.3468 $w=1.8e-07 $l=2.35e-07 $layer=POLY_cond $X=9.235 $Y=2.08
+ $X2=9.235 $Y2=2.315
r141 2 54 600 $w=1.7e-07 $l=8.36645e-07 $layer=licon1_PDIFF $count=1 $X=10.11
+ $Y=1.9 $X2=10.26 $Y2=2.665
r142 1 42 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=9.825
+ $Y=0.37 $X2=9.965 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__SDFXTP_2%A_1592_424# 1 2 7 9 10 12 13 16 18 19 23 26
+ 32 34
c88 23 0 2.99265e-19 $X=9.94 $Y=1.575
r89 26 29 5.9927 $w=2.48e-07 $l=1.3e-07 $layer=LI1_cond $X=8.15 $Y=2.575
+ $X2=8.15 $Y2=2.705
r90 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.94
+ $Y=1.575 $X2=9.94 $Y2=1.575
r91 21 23 17.4613 $w=3.28e-07 $l=5e-07 $layer=LI1_cond $X=9.94 $Y=2.075 $X2=9.94
+ $Y2=1.575
r92 20 34 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.06 $Y=2.16
+ $X2=8.975 $Y2=2.16
r93 19 21 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=9.775 $Y=2.16
+ $X2=9.94 $Y2=2.075
r94 19 20 46.6471 $w=1.68e-07 $l=7.15e-07 $layer=LI1_cond $X=9.775 $Y=2.16
+ $X2=9.06 $Y2=2.16
r95 17 34 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.975 $Y=2.245
+ $X2=8.975 $Y2=2.16
r96 17 18 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=8.975 $Y=2.245
+ $X2=8.975 $Y2=2.49
r97 16 34 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.975 $Y=2.075
+ $X2=8.975 $Y2=2.16
r98 15 32 14.5831 $w=3.43e-07 $l=5.1225e-07 $layer=LI1_cond $X=8.975 $Y=0.81
+ $X2=8.565 $Y2=0.58
r99 15 16 82.5294 $w=1.68e-07 $l=1.265e-06 $layer=LI1_cond $X=8.975 $Y=0.81
+ $X2=8.975 $Y2=2.075
r100 14 26 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.275 $Y=2.575
+ $X2=8.15 $Y2=2.575
r101 13 18 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.89 $Y=2.575
+ $X2=8.975 $Y2=2.49
r102 13 14 40.123 $w=1.68e-07 $l=6.15e-07 $layer=LI1_cond $X=8.89 $Y=2.575
+ $X2=8.275 $Y2=2.575
r103 10 24 53.362 $w=2.8e-07 $l=3.10242e-07 $layer=POLY_cond $X=10.035 $Y=1.825
+ $X2=9.9 $Y2=1.575
r104 10 12 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=10.035 $Y=1.825
+ $X2=10.035 $Y2=2.4
r105 7 24 77.462 $w=2.8e-07 $l=4.58912e-07 $layer=POLY_cond $X=9.75 $Y=1.185
+ $X2=9.9 $Y2=1.575
r106 7 9 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=9.75 $Y=1.185
+ $X2=9.75 $Y2=0.74
r107 2 29 600 $w=1.7e-07 $l=6.55725e-07 $layer=licon1_PDIFF $count=1 $X=7.96
+ $Y=2.12 $X2=8.11 $Y2=2.705
r108 1 32 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=8.425
+ $Y=0.37 $X2=8.565 $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_HS__SDFXTP_2%VPWR 1 2 3 4 5 6 7 24 28 32 36 40 44 46 51
+ 52 54 55 56 58 70 81 85 90 96 99 106 111 115
c137 24 0 1.79254e-19 $X=0.78 $Y=2.44
r138 114 115 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.76 $Y=3.33
+ $X2=11.76 $Y2=3.33
r139 111 112 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.8 $Y=3.33
+ $X2=10.8 $Y2=3.33
r140 107 109 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.84 $Y=3.33
+ $X2=9.36 $Y2=3.33
r141 106 109 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=9.36 $Y=3.33
+ $X2=9.36 $Y2=3.33
r142 106 107 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.84 $Y=3.33
+ $X2=9.84 $Y2=3.33
r143 102 103 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r144 99 102 9.54318 $w=4.68e-07 $l=3.75e-07 $layer=LI1_cond $X=4.135 $Y=2.955
+ $X2=4.135 $Y2=3.33
r145 96 97 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r146 94 115 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.28 $Y=3.33
+ $X2=11.76 $Y2=3.33
r147 94 112 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.28 $Y=3.33
+ $X2=10.8 $Y2=3.33
r148 93 94 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.28 $Y=3.33
+ $X2=11.28 $Y2=3.33
r149 91 111 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=10.905 $Y=3.33
+ $X2=10.78 $Y2=3.33
r150 91 93 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=10.905 $Y=3.33
+ $X2=11.28 $Y2=3.33
r151 90 114 4.01252 $w=1.7e-07 $l=1.82e-07 $layer=LI1_cond $X=11.635 $Y=3.33
+ $X2=11.817 $Y2=3.33
r152 90 93 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=11.635 $Y=3.33
+ $X2=11.28 $Y2=3.33
r153 89 112 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.32 $Y=3.33
+ $X2=10.8 $Y2=3.33
r154 89 107 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.32 $Y=3.33
+ $X2=9.84 $Y2=3.33
r155 88 89 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.32 $Y=3.33
+ $X2=10.32 $Y2=3.33
r156 86 106 12.9051 $w=1.7e-07 $l=3.15e-07 $layer=LI1_cond $X=9.925 $Y=3.33
+ $X2=9.61 $Y2=3.33
r157 86 88 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=9.925 $Y=3.33
+ $X2=10.32 $Y2=3.33
r158 85 111 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=10.655 $Y=3.33
+ $X2=10.78 $Y2=3.33
r159 85 88 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=10.655 $Y=3.33
+ $X2=10.32 $Y2=3.33
r160 84 109 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=9.36 $Y2=3.33
r161 83 84 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r162 81 106 12.9051 $w=1.7e-07 $l=3.15e-07 $layer=LI1_cond $X=9.295 $Y=3.33
+ $X2=9.61 $Y2=3.33
r163 81 83 152.337 $w=1.68e-07 $l=2.335e-06 $layer=LI1_cond $X=9.295 $Y=3.33
+ $X2=6.96 $Y2=3.33
r164 80 84 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=6.96 $Y2=3.33
r165 79 80 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r166 77 103 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=4.08 $Y2=3.33
r167 76 79 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=4.56 $Y=3.33
+ $X2=6.48 $Y2=3.33
r168 76 77 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r169 74 102 6.76998 $w=1.7e-07 $l=2.35e-07 $layer=LI1_cond $X=4.37 $Y=3.33
+ $X2=4.135 $Y2=3.33
r170 74 76 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=4.37 $Y=3.33
+ $X2=4.56 $Y2=3.33
r171 73 103 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.08 $Y2=3.33
r172 72 73 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r173 70 102 6.76998 $w=1.7e-07 $l=2.35e-07 $layer=LI1_cond $X=3.9 $Y=3.33
+ $X2=4.135 $Y2=3.33
r174 70 72 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=3.9 $Y=3.33 $X2=3.6
+ $Y2=3.33
r175 69 73 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.6 $Y2=3.33
r176 68 69 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r177 66 69 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.64 $Y2=3.33
r178 66 97 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r179 65 68 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.2 $Y=3.33
+ $X2=2.64 $Y2=3.33
r180 65 66 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r181 63 96 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.945 $Y=3.33
+ $X2=0.78 $Y2=3.33
r182 63 65 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.945 $Y=3.33
+ $X2=1.2 $Y2=3.33
r183 61 97 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r184 60 61 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r185 58 96 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.615 $Y=3.33
+ $X2=0.78 $Y2=3.33
r186 58 60 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=0.615 $Y=3.33
+ $X2=0.24 $Y2=3.33
r187 56 80 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=3.33 $X2=6.48
+ $Y2=3.33
r188 56 77 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=6 $Y=3.33
+ $X2=4.56 $Y2=3.33
r189 54 79 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=6.585 $Y=3.33
+ $X2=6.48 $Y2=3.33
r190 54 55 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.585 $Y=3.33
+ $X2=6.71 $Y2=3.33
r191 53 83 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=6.835 $Y=3.33
+ $X2=6.96 $Y2=3.33
r192 53 55 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.835 $Y=3.33
+ $X2=6.71 $Y2=3.33
r193 51 68 2.93583 $w=1.68e-07 $l=4.5e-08 $layer=LI1_cond $X=2.685 $Y=3.33
+ $X2=2.64 $Y2=3.33
r194 51 52 10.5822 $w=1.7e-07 $l=2.25e-07 $layer=LI1_cond $X=2.685 $Y=3.33
+ $X2=2.91 $Y2=3.33
r195 50 72 30.3369 $w=1.68e-07 $l=4.65e-07 $layer=LI1_cond $X=3.135 $Y=3.33
+ $X2=3.6 $Y2=3.33
r196 50 52 10.5822 $w=1.7e-07 $l=2.25e-07 $layer=LI1_cond $X=3.135 $Y=3.33
+ $X2=2.91 $Y2=3.33
r197 46 49 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=11.76 $Y=1.985
+ $X2=11.76 $Y2=2.815
r198 44 114 3.13065 $w=2.5e-07 $l=1.09864e-07 $layer=LI1_cond $X=11.76 $Y=3.245
+ $X2=11.817 $Y2=3.33
r199 44 49 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=11.76 $Y=3.245
+ $X2=11.76 $Y2=2.815
r200 40 43 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=10.78 $Y=1.985
+ $X2=10.78 $Y2=2.815
r201 38 111 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=10.78 $Y=3.245
+ $X2=10.78 $Y2=3.33
r202 38 43 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=10.78 $Y=3.245
+ $X2=10.78 $Y2=2.815
r203 34 106 2.6323 $w=6.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.61 $Y=3.245
+ $X2=9.61 $Y2=3.33
r204 34 36 9.30283 $w=6.28e-07 $l=4.9e-07 $layer=LI1_cond $X=9.61 $Y=3.245
+ $X2=9.61 $Y2=2.755
r205 30 55 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.71 $Y=3.245
+ $X2=6.71 $Y2=3.33
r206 30 32 22.8184 $w=2.48e-07 $l=4.95e-07 $layer=LI1_cond $X=6.71 $Y=3.245
+ $X2=6.71 $Y2=2.75
r207 26 52 1.79621 $w=4.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.91 $Y=3.245
+ $X2=2.91 $Y2=3.33
r208 26 28 7.70806 $w=4.48e-07 $l=2.9e-07 $layer=LI1_cond $X=2.91 $Y=3.245
+ $X2=2.91 $Y2=2.955
r209 22 96 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.78 $Y=3.245
+ $X2=0.78 $Y2=3.33
r210 22 24 28.1126 $w=3.28e-07 $l=8.05e-07 $layer=LI1_cond $X=0.78 $Y=3.245
+ $X2=0.78 $Y2=2.44
r211 7 49 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=11.57
+ $Y=1.84 $X2=11.72 $Y2=2.815
r212 7 46 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=11.57
+ $Y=1.84 $X2=11.72 $Y2=1.985
r213 6 43 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=10.675
+ $Y=1.84 $X2=10.82 $Y2=2.815
r214 6 40 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=10.675
+ $Y=1.84 $X2=10.82 $Y2=1.985
r215 5 36 300 $w=1.7e-07 $l=6.22495e-07 $layer=licon1_PDIFF $count=2 $X=9.31
+ $Y=2.48 $X2=9.81 $Y2=2.755
r216 4 32 600 $w=1.7e-07 $l=2.74955e-07 $layer=licon1_PDIFF $count=1 $X=6.6
+ $Y=2.54 $X2=6.75 $Y2=2.75
r217 3 99 600 $w=1.7e-07 $l=1.21776e-06 $layer=licon1_PDIFF $count=1 $X=3.92
+ $Y=1.84 $X2=4.135 $Y2=2.955
r218 2 28 600 $w=1.7e-07 $l=8.24409e-07 $layer=licon1_PDIFF $count=1 $X=2.615
+ $Y=2.265 $X2=2.91 $Y2=2.955
r219 1 24 300 $w=1.7e-07 $l=2.73861e-07 $layer=licon1_PDIFF $count=2 $X=0.58
+ $Y=2.265 $X2=0.78 $Y2=2.44
.ends

.subckt PM_SKY130_FD_SC_HS__SDFXTP_2%A_300_453# 1 2 3 4 13 17 20 21 22 24 25 28
+ 29 30 31 34 37 40 44 45 49
c135 17 0 1.47911e-19 $X=2.95 $Y=2.487
r136 46 49 4.67658 $w=3.43e-07 $l=1.4e-07 $layer=LI1_cond $X=4.79 $Y=0.767
+ $X2=4.93 $Y2=0.767
r137 40 42 0.977664 $w=5.73e-07 $l=4.7e-08 $layer=LI1_cond $X=1.772 $Y=2.44
+ $X2=1.772 $Y2=2.487
r138 35 37 5.9927 $w=2.48e-07 $l=1.3e-07 $layer=LI1_cond $X=5.26 $Y=2.62
+ $X2=5.26 $Y2=2.75
r139 33 46 4.88813 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=4.79 $Y=0.94
+ $X2=4.79 $Y2=0.767
r140 33 34 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=4.79 $Y=0.94
+ $X2=4.79 $Y2=1.3
r141 32 45 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.485 $Y=2.535
+ $X2=4.4 $Y2=2.535
r142 31 35 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=5.135 $Y=2.535
+ $X2=5.26 $Y2=2.62
r143 31 32 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=5.135 $Y=2.535
+ $X2=4.485 $Y2=2.535
r144 29 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.705 $Y=1.385
+ $X2=4.79 $Y2=1.3
r145 29 30 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=4.705 $Y=1.385
+ $X2=4.485 $Y2=1.385
r146 28 45 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.4 $Y=2.45 $X2=4.4
+ $Y2=2.535
r147 27 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.4 $Y=1.47
+ $X2=4.485 $Y2=1.385
r148 27 28 63.9358 $w=1.68e-07 $l=9.8e-07 $layer=LI1_cond $X=4.4 $Y=1.47 $X2=4.4
+ $Y2=2.45
r149 26 44 4.18896 $w=2.17e-07 $l=1.06325e-07 $layer=LI1_cond $X=3.12 $Y=2.535
+ $X2=3.035 $Y2=2.487
r150 25 45 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.315 $Y=2.535
+ $X2=4.4 $Y2=2.535
r151 25 26 77.9626 $w=1.68e-07 $l=1.195e-06 $layer=LI1_cond $X=4.315 $Y=2.535
+ $X2=3.12 $Y2=2.535
r152 24 44 2.24312 $w=1.7e-07 $l=1.32e-07 $layer=LI1_cond $X=3.035 $Y=2.355
+ $X2=3.035 $Y2=2.487
r153 23 24 71.1123 $w=1.68e-07 $l=1.09e-06 $layer=LI1_cond $X=3.035 $Y=1.265
+ $X2=3.035 $Y2=2.355
r154 21 23 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.95 $Y=1.18
+ $X2=3.035 $Y2=1.265
r155 21 22 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=2.95 $Y=1.18
+ $X2=2.545 $Y2=1.18
r156 20 22 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.46 $Y=1.095
+ $X2=2.545 $Y2=1.18
r157 19 20 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=2.46 $Y=0.68
+ $X2=2.46 $Y2=1.095
r158 18 42 5.29924 $w=2.65e-07 $l=2.88e-07 $layer=LI1_cond $X=2.06 $Y=2.487
+ $X2=1.772 $Y2=2.487
r159 17 44 4.18896 $w=2.17e-07 $l=8.5e-08 $layer=LI1_cond $X=2.95 $Y=2.487
+ $X2=3.035 $Y2=2.487
r160 17 18 38.7047 $w=2.63e-07 $l=8.9e-07 $layer=LI1_cond $X=2.95 $Y=2.487
+ $X2=2.06 $Y2=2.487
r161 13 19 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.375 $Y=0.515
+ $X2=2.46 $Y2=0.68
r162 13 15 20.7789 $w=3.28e-07 $l=5.95e-07 $layer=LI1_cond $X=2.375 $Y=0.515
+ $X2=1.78 $Y2=0.515
r163 4 37 600 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_PDIFF $count=1 $X=5.155
+ $Y=2.54 $X2=5.3 $Y2=2.75
r164 3 40 300 $w=1.7e-07 $l=3.46627e-07 $layer=licon1_PDIFF $count=2 $X=1.5
+ $Y=2.265 $X2=1.77 $Y2=2.44
r165 2 49 182 $w=1.7e-07 $l=3.29621e-07 $layer=licon1_NDIFF $count=1 $X=4.785
+ $Y=0.5 $X2=4.93 $Y2=0.765
r166 1 15 182 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_NDIFF $count=1 $X=1.505
+ $Y=0.37 $X2=1.78 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__SDFXTP_2%Q 1 2 9 13 14 15 16 24 33
c23 33 0 1.10546e-19 $X=11.27 $Y=1.82
r24 15 16 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=11.27 $Y=2.405
+ $X2=11.27 $Y2=2.775
r25 14 24 0.628605 $w=3.28e-07 $l=1.8e-08 $layer=LI1_cond $X=11.27 $Y=1.967
+ $X2=11.27 $Y2=1.985
r26 14 33 7.83357 $w=3.28e-07 $l=1.47e-07 $layer=LI1_cond $X=11.27 $Y=1.967
+ $X2=11.27 $Y2=1.82
r27 14 15 12.3276 $w=3.28e-07 $l=3.53e-07 $layer=LI1_cond $X=11.27 $Y=2.052
+ $X2=11.27 $Y2=2.405
r28 14 24 2.33981 $w=3.28e-07 $l=6.7e-08 $layer=LI1_cond $X=11.27 $Y=2.052
+ $X2=11.27 $Y2=1.985
r29 13 33 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=11.3 $Y=1.05
+ $X2=11.3 $Y2=1.82
r30 7 13 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=11.22 $Y=0.885
+ $X2=11.22 $Y2=1.05
r31 7 9 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=11.22 $Y=0.885
+ $X2=11.22 $Y2=0.515
r32 2 16 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=11.12
+ $Y=1.84 $X2=11.27 $Y2=2.815
r33 2 24 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=11.12
+ $Y=1.84 $X2=11.27 $Y2=1.985
r34 1 9 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=11.08
+ $Y=0.37 $X2=11.22 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__SDFXTP_2%VGND 1 2 3 4 5 6 7 26 30 34 38 42 46 48 50
+ 53 54 56 57 58 70 77 82 87 93 96 99 102 106
r135 105 106 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.76 $Y=0
+ $X2=11.76 $Y2=0
r136 102 103 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.8 $Y=0
+ $X2=10.8 $Y2=0
r137 99 100 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=9.36 $Y=0
+ $X2=9.36 $Y2=0
r138 96 97 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=0 $X2=6.96
+ $Y2=0
r139 93 94 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r140 91 106 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.28 $Y=0
+ $X2=11.76 $Y2=0
r141 91 103 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.28 $Y=0
+ $X2=10.8 $Y2=0
r142 90 91 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.28 $Y=0
+ $X2=11.28 $Y2=0
r143 88 102 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=10.885 $Y=0
+ $X2=10.75 $Y2=0
r144 88 90 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=10.885 $Y=0
+ $X2=11.28 $Y2=0
r145 87 105 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=11.555 $Y=0
+ $X2=11.777 $Y2=0
r146 87 90 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=11.555 $Y=0
+ $X2=11.28 $Y2=0
r147 86 103 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.32 $Y=0
+ $X2=10.8 $Y2=0
r148 86 100 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=10.32 $Y=0
+ $X2=9.36 $Y2=0
r149 85 86 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.32 $Y=0
+ $X2=10.32 $Y2=0
r150 83 99 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.63 $Y=0 $X2=9.465
+ $Y2=0
r151 83 85 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=9.63 $Y=0 $X2=10.32
+ $Y2=0
r152 82 102 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=10.615 $Y=0
+ $X2=10.75 $Y2=0
r153 82 85 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=10.615 $Y=0
+ $X2=10.32 $Y2=0
r154 81 100 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=7.44 $Y=0
+ $X2=9.36 $Y2=0
r155 81 97 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=0 $X2=6.96
+ $Y2=0
r156 80 81 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=7.44 $Y=0
+ $X2=7.44 $Y2=0
r157 78 96 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.05 $Y=0 $X2=6.885
+ $Y2=0
r158 78 80 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=7.05 $Y=0 $X2=7.44
+ $Y2=0
r159 77 99 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.3 $Y=0 $X2=9.465
+ $Y2=0
r160 77 80 121.348 $w=1.68e-07 $l=1.86e-06 $layer=LI1_cond $X=9.3 $Y=0 $X2=7.44
+ $Y2=0
r161 76 97 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=0 $X2=6.96
+ $Y2=0
r162 75 76 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=6.48 $Y=0 $X2=6.48
+ $Y2=0
r163 72 75 156.578 $w=1.68e-07 $l=2.4e-06 $layer=LI1_cond $X=4.08 $Y=0 $X2=6.48
+ $Y2=0
r164 72 73 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r165 70 96 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.72 $Y=0 $X2=6.885
+ $Y2=0
r166 70 75 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=6.72 $Y=0 $X2=6.48
+ $Y2=0
r167 69 73 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.08
+ $Y2=0
r168 68 69 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r169 66 69 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.6
+ $Y2=0
r170 65 66 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r171 63 66 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=1.2 $Y=0 $X2=2.64
+ $Y2=0
r172 63 94 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r173 62 65 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.2 $Y=0 $X2=2.64
+ $Y2=0
r174 62 63 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r175 60 93 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.99 $Y=0 $X2=0.825
+ $Y2=0
r176 60 62 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=0.99 $Y=0 $X2=1.2
+ $Y2=0
r177 58 76 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=0 $X2=6.48
+ $Y2=0
r178 58 73 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=6 $Y=0 $X2=4.08
+ $Y2=0
r179 56 68 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=3.705 $Y=0 $X2=3.6
+ $Y2=0
r180 56 57 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.705 $Y=0 $X2=3.87
+ $Y2=0
r181 55 72 2.93583 $w=1.68e-07 $l=4.5e-08 $layer=LI1_cond $X=4.035 $Y=0 $X2=4.08
+ $Y2=0
r182 55 57 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.035 $Y=0 $X2=3.87
+ $Y2=0
r183 53 65 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=2.715 $Y=0 $X2=2.64
+ $Y2=0
r184 53 54 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.715 $Y=0 $X2=2.845
+ $Y2=0
r185 52 68 40.7754 $w=1.68e-07 $l=6.25e-07 $layer=LI1_cond $X=2.975 $Y=0 $X2=3.6
+ $Y2=0
r186 52 54 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.975 $Y=0 $X2=2.845
+ $Y2=0
r187 48 105 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=11.72 $Y=0.085
+ $X2=11.777 $Y2=0
r188 48 50 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=11.72 $Y=0.085
+ $X2=11.72 $Y2=0.515
r189 44 102 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.75 $Y=0.085
+ $X2=10.75 $Y2=0
r190 44 46 18.3537 $w=2.68e-07 $l=4.3e-07 $layer=LI1_cond $X=10.75 $Y=0.085
+ $X2=10.75 $Y2=0.515
r191 40 99 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.465 $Y=0.085
+ $X2=9.465 $Y2=0
r192 40 42 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=9.465 $Y=0.085
+ $X2=9.465 $Y2=0.58
r193 36 96 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.885 $Y=0.085
+ $X2=6.885 $Y2=0
r194 36 38 10.4768 $w=3.28e-07 $l=3e-07 $layer=LI1_cond $X=6.885 $Y=0.085
+ $X2=6.885 $Y2=0.385
r195 32 57 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.87 $Y=0.085
+ $X2=3.87 $Y2=0
r196 32 34 17.8105 $w=3.28e-07 $l=5.1e-07 $layer=LI1_cond $X=3.87 $Y=0.085
+ $X2=3.87 $Y2=0.595
r197 28 54 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=2.845 $Y=0.085
+ $X2=2.845 $Y2=0
r198 28 30 21.9407 $w=2.58e-07 $l=4.95e-07 $layer=LI1_cond $X=2.845 $Y=0.085
+ $X2=2.845 $Y2=0.58
r199 24 93 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.825 $Y=0.085
+ $X2=0.825 $Y2=0
r200 24 26 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=0.825 $Y=0.085
+ $X2=0.825 $Y2=0.535
r201 7 50 91 $w=1.7e-07 $l=2.26164e-07 $layer=licon1_NDIFF $count=2 $X=11.555
+ $Y=0.37 $X2=11.72 $Y2=0.515
r202 6 46 91 $w=1.7e-07 $l=2.78209e-07 $layer=licon1_NDIFF $count=2 $X=10.575
+ $Y=0.37 $X2=10.79 $Y2=0.515
r203 5 42 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=9.325
+ $Y=0.37 $X2=9.465 $Y2=0.58
r204 4 38 182 $w=1.7e-07 $l=2.71477e-07 $layer=licon1_NDIFF $count=1 $X=6.665
+ $Y=0.5 $X2=6.885 $Y2=0.385
r205 3 34 182 $w=1.7e-07 $l=2.88531e-07 $layer=licon1_NDIFF $count=1 $X=3.725
+ $Y=0.37 $X2=3.87 $Y2=0.595
r206 2 30 182 $w=1.7e-07 $l=3.44347e-07 $layer=licon1_NDIFF $count=1 $X=2.6
+ $Y=0.37 $X2=2.855 $Y2=0.58
r207 1 26 182 $w=1.7e-07 $l=2.80624e-07 $layer=licon1_NDIFF $count=1 $X=0.615
+ $Y=0.37 $X2=0.825 $Y2=0.535
.ends

