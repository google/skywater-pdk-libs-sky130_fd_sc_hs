* File: sky130_fd_sc_hs__nand4_4.pex.spice
* Created: Tue Sep  1 20:10:01 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HS__NAND4_4%D 3 7 9 13 15 17 20 22 24 25 26 27 28 29 30
+ 31 32 49
c74 32 0 1.29429e-20 $X=2.16 $Y=1.665
c75 22 0 1.02686e-19 $X=2.26 $Y=1.765
c76 20 0 7.27676e-20 $X=2.195 $Y=0.74
r77 49 50 8.6547 $w=3.62e-07 $l=6.5e-08 $layer=POLY_cond $X=2.195 $Y=1.557
+ $X2=2.26 $Y2=1.557
r78 47 49 11.9834 $w=3.62e-07 $l=9e-08 $layer=POLY_cond $X=2.105 $Y=1.557
+ $X2=2.195 $Y2=1.557
r79 47 48 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.105
+ $Y=1.515 $X2=2.105 $Y2=1.515
r80 45 47 45.9365 $w=3.62e-07 $l=3.45e-07 $layer=POLY_cond $X=1.76 $Y=1.557
+ $X2=2.105 $Y2=1.557
r81 44 45 35.2845 $w=3.62e-07 $l=2.65e-07 $layer=POLY_cond $X=1.495 $Y=1.557
+ $X2=1.76 $Y2=1.557
r82 42 44 9.32044 $w=3.62e-07 $l=7e-08 $layer=POLY_cond $X=1.425 $Y=1.557
+ $X2=1.495 $Y2=1.557
r83 42 43 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.425
+ $Y=1.515 $X2=1.425 $Y2=1.515
r84 39 40 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=0.745
+ $Y=1.515 $X2=0.745 $Y2=1.515
r85 32 48 1.47406 $w=4.28e-07 $l=5.5e-08 $layer=LI1_cond $X=2.16 $Y=1.565
+ $X2=2.105 $Y2=1.565
r86 31 48 11.3904 $w=4.28e-07 $l=4.25e-07 $layer=LI1_cond $X=1.68 $Y=1.565
+ $X2=2.105 $Y2=1.565
r87 31 43 6.83426 $w=4.28e-07 $l=2.55e-07 $layer=LI1_cond $X=1.68 $Y=1.565
+ $X2=1.425 $Y2=1.565
r88 30 43 6.03022 $w=4.28e-07 $l=2.25e-07 $layer=LI1_cond $X=1.2 $Y=1.565
+ $X2=1.425 $Y2=1.565
r89 30 40 12.1945 $w=4.28e-07 $l=4.55e-07 $layer=LI1_cond $X=1.2 $Y=1.565
+ $X2=0.745 $Y2=1.565
r90 29 40 0.670025 $w=4.28e-07 $l=2.5e-08 $layer=LI1_cond $X=0.72 $Y=1.565
+ $X2=0.745 $Y2=1.565
r91 28 29 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=0.24 $Y=1.565
+ $X2=0.72 $Y2=1.565
r92 26 39 30.6007 $w=3.3e-07 $l=1.75e-07 $layer=POLY_cond $X=0.92 $Y=1.515
+ $X2=0.745 $Y2=1.515
r93 26 27 10.1687 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=0.92 $Y=1.515
+ $X2=0.995 $Y2=1.515
r94 25 39 30.6007 $w=3.3e-07 $l=1.75e-07 $layer=POLY_cond $X=0.57 $Y=1.515
+ $X2=0.745 $Y2=1.515
r95 22 50 23.4391 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=2.26 $Y=1.765
+ $X2=2.26 $Y2=1.557
r96 22 24 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.26 $Y=1.765
+ $X2=2.26 $Y2=2.4
r97 18 49 23.4391 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.195 $Y=1.35
+ $X2=2.195 $Y2=1.557
r98 18 20 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.195 $Y=1.35
+ $X2=2.195 $Y2=0.74
r99 15 45 23.4391 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=1.76 $Y=1.765
+ $X2=1.76 $Y2=1.557
r100 15 17 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.76 $Y=1.765
+ $X2=1.76 $Y2=2.4
r101 11 44 23.4391 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.495 $Y=1.35
+ $X2=1.495 $Y2=1.557
r102 11 13 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.495 $Y=1.35
+ $X2=1.495 $Y2=0.74
r103 10 27 10.1687 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=1.07 $Y=1.515
+ $X2=0.995 $Y2=1.515
r104 9 42 1.13569 $w=3.62e-07 $l=4.44297e-08 $layer=POLY_cond $X=1.42 $Y=1.515
+ $X2=1.425 $Y2=1.557
r105 9 10 61.2015 $w=3.3e-07 $l=3.5e-07 $layer=POLY_cond $X=1.42 $Y=1.515
+ $X2=1.07 $Y2=1.515
r106 5 27 16.9349 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.995 $Y=1.35
+ $X2=0.995 $Y2=1.515
r107 5 7 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=0.995 $Y=1.35
+ $X2=0.995 $Y2=0.74
r108 1 25 32.1775 $w=3.3e-07 $l=1.98997e-07 $layer=POLY_cond $X=0.495 $Y=1.35
+ $X2=0.57 $Y2=1.515
r109 1 3 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=0.495 $Y=1.35
+ $X2=0.495 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HS__NAND4_4%C 3 5 7 10 12 14 17 21 23 24 25 26 43
c58 26 0 1.96965e-19 $X=4.08 $Y=1.665
c59 5 0 1.29429e-20 $X=2.71 $Y=1.765
r60 43 45 24.7179 $w=3.51e-07 $l=1.8e-07 $layer=POLY_cond $X=3.805 $Y=1.557
+ $X2=3.985 $Y2=1.557
r61 43 44 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.805
+ $Y=1.515 $X2=3.805 $Y2=1.515
r62 41 43 34.3305 $w=3.51e-07 $l=2.5e-07 $layer=POLY_cond $X=3.555 $Y=1.557
+ $X2=3.805 $Y2=1.557
r63 40 41 2.05983 $w=3.51e-07 $l=1.5e-08 $layer=POLY_cond $X=3.54 $Y=1.557
+ $X2=3.555 $Y2=1.557
r64 38 40 10.2991 $w=3.51e-07 $l=7.5e-08 $layer=POLY_cond $X=3.465 $Y=1.557
+ $X2=3.54 $Y2=1.557
r65 38 39 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=3.465
+ $Y=1.515 $X2=3.465 $Y2=1.515
r66 36 38 46.6895 $w=3.51e-07 $l=3.4e-07 $layer=POLY_cond $X=3.125 $Y=1.557
+ $X2=3.465 $Y2=1.557
r67 34 36 46.6895 $w=3.51e-07 $l=3.4e-07 $layer=POLY_cond $X=2.785 $Y=1.557
+ $X2=3.125 $Y2=1.557
r68 34 35 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=2.785
+ $Y=1.515 $X2=2.785 $Y2=1.515
r69 32 34 10.2991 $w=3.51e-07 $l=7.5e-08 $layer=POLY_cond $X=2.71 $Y=1.557
+ $X2=2.785 $Y2=1.557
r70 31 32 2.05983 $w=3.51e-07 $l=1.5e-08 $layer=POLY_cond $X=2.695 $Y=1.557
+ $X2=2.71 $Y2=1.557
r71 26 44 7.37028 $w=4.28e-07 $l=2.75e-07 $layer=LI1_cond $X=4.08 $Y=1.565
+ $X2=3.805 $Y2=1.565
r72 25 44 5.4942 $w=4.28e-07 $l=2.05e-07 $layer=LI1_cond $X=3.6 $Y=1.565
+ $X2=3.805 $Y2=1.565
r73 25 39 3.61813 $w=4.28e-07 $l=1.35e-07 $layer=LI1_cond $X=3.6 $Y=1.565
+ $X2=3.465 $Y2=1.565
r74 24 39 9.24634 $w=4.28e-07 $l=3.45e-07 $layer=LI1_cond $X=3.12 $Y=1.565
+ $X2=3.465 $Y2=1.565
r75 24 35 8.97834 $w=4.28e-07 $l=3.35e-07 $layer=LI1_cond $X=3.12 $Y=1.565
+ $X2=2.785 $Y2=1.565
r76 23 35 3.88615 $w=4.28e-07 $l=1.45e-07 $layer=LI1_cond $X=2.64 $Y=1.565
+ $X2=2.785 $Y2=1.565
r77 19 45 22.6971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.985 $Y=1.35
+ $X2=3.985 $Y2=1.557
r78 19 21 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=3.985 $Y=1.35
+ $X2=3.985 $Y2=0.74
r79 15 41 22.6971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.555 $Y=1.35
+ $X2=3.555 $Y2=1.557
r80 15 17 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=3.555 $Y=1.35
+ $X2=3.555 $Y2=0.74
r81 12 40 22.6971 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=3.54 $Y=1.765
+ $X2=3.54 $Y2=1.557
r82 12 14 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.54 $Y=1.765
+ $X2=3.54 $Y2=2.4
r83 8 36 22.6971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.125 $Y=1.35
+ $X2=3.125 $Y2=1.557
r84 8 10 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=3.125 $Y=1.35
+ $X2=3.125 $Y2=0.74
r85 5 32 22.6971 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=2.71 $Y=1.765
+ $X2=2.71 $Y2=1.557
r86 5 7 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.71 $Y=1.765
+ $X2=2.71 $Y2=2.4
r87 1 31 22.6971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.695 $Y=1.35
+ $X2=2.695 $Y2=1.557
r88 1 3 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.695 $Y=1.35
+ $X2=2.695 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HS__NAND4_4%B 1 3 6 8 10 13 17 21 23 24 25 26 43
c65 1 0 9.42782e-20 $X=4.56 $Y=1.765
r66 43 45 37.6127 $w=3.46e-07 $l=2.7e-07 $layer=POLY_cond $X=5.995 $Y=1.557
+ $X2=6.265 $Y2=1.557
r67 43 44 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.995
+ $Y=1.515 $X2=5.995 $Y2=1.515
r68 41 43 22.289 $w=3.46e-07 $l=1.6e-07 $layer=POLY_cond $X=5.835 $Y=1.557
+ $X2=5.995 $Y2=1.557
r69 40 41 59.9017 $w=3.46e-07 $l=4.3e-07 $layer=POLY_cond $X=5.405 $Y=1.557
+ $X2=5.835 $Y2=1.557
r70 39 40 2.0896 $w=3.46e-07 $l=1.5e-08 $layer=POLY_cond $X=5.39 $Y=1.557
+ $X2=5.405 $Y2=1.557
r71 37 39 10.448 $w=3.46e-07 $l=7.5e-08 $layer=POLY_cond $X=5.315 $Y=1.557
+ $X2=5.39 $Y2=1.557
r72 37 38 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=5.315
+ $Y=1.515 $X2=5.315 $Y2=1.515
r73 35 37 47.3642 $w=3.46e-07 $l=3.4e-07 $layer=POLY_cond $X=4.975 $Y=1.557
+ $X2=5.315 $Y2=1.557
r74 33 35 47.3642 $w=3.46e-07 $l=3.4e-07 $layer=POLY_cond $X=4.635 $Y=1.557
+ $X2=4.975 $Y2=1.557
r75 33 34 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=4.635
+ $Y=1.515 $X2=4.635 $Y2=1.515
r76 31 33 10.448 $w=3.46e-07 $l=7.5e-08 $layer=POLY_cond $X=4.56 $Y=1.557
+ $X2=4.635 $Y2=1.557
r77 26 44 0.134005 $w=4.28e-07 $l=5e-09 $layer=LI1_cond $X=6 $Y=1.565 $X2=5.995
+ $Y2=1.565
r78 25 44 12.7305 $w=4.28e-07 $l=4.75e-07 $layer=LI1_cond $X=5.52 $Y=1.565
+ $X2=5.995 $Y2=1.565
r79 25 38 5.4942 $w=4.28e-07 $l=2.05e-07 $layer=LI1_cond $X=5.52 $Y=1.565
+ $X2=5.315 $Y2=1.565
r80 24 38 7.37028 $w=4.28e-07 $l=2.75e-07 $layer=LI1_cond $X=5.04 $Y=1.565
+ $X2=5.315 $Y2=1.565
r81 24 34 10.8544 $w=4.28e-07 $l=4.05e-07 $layer=LI1_cond $X=5.04 $Y=1.565
+ $X2=4.635 $Y2=1.565
r82 23 34 2.01008 $w=4.28e-07 $l=7.5e-08 $layer=LI1_cond $X=4.56 $Y=1.565
+ $X2=4.635 $Y2=1.565
r83 19 45 22.3532 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=6.265 $Y=1.35
+ $X2=6.265 $Y2=1.557
r84 19 21 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=6.265 $Y=1.35
+ $X2=6.265 $Y2=0.74
r85 15 41 22.3532 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=5.835 $Y=1.35
+ $X2=5.835 $Y2=1.557
r86 15 17 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=5.835 $Y=1.35
+ $X2=5.835 $Y2=0.74
r87 11 40 22.3532 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=5.405 $Y=1.35
+ $X2=5.405 $Y2=1.557
r88 11 13 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=5.405 $Y=1.35
+ $X2=5.405 $Y2=0.74
r89 8 39 22.3532 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=5.39 $Y=1.765
+ $X2=5.39 $Y2=1.557
r90 8 10 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=5.39 $Y=1.765
+ $X2=5.39 $Y2=2.4
r91 4 35 22.3532 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.975 $Y=1.35
+ $X2=4.975 $Y2=1.557
r92 4 6 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=4.975 $Y=1.35
+ $X2=4.975 $Y2=0.74
r93 1 31 22.3532 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=4.56 $Y=1.765
+ $X2=4.56 $Y2=1.557
r94 1 3 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=4.56 $Y=1.765
+ $X2=4.56 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_HS__NAND4_4%A 3 7 9 11 14 16 18 21 23 24 25 26 27 31
r68 42 44 44.0087 $w=3.45e-07 $l=3.15e-07 $layer=POLY_cond $X=7.24 $Y=1.557
+ $X2=7.555 $Y2=1.557
r69 42 43 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=7.24
+ $Y=1.515 $X2=7.24 $Y2=1.515
r70 40 42 5.58841 $w=3.45e-07 $l=4e-08 $layer=POLY_cond $X=7.2 $Y=1.557 $X2=7.24
+ $Y2=1.557
r71 39 40 10.4783 $w=3.45e-07 $l=7.5e-08 $layer=POLY_cond $X=7.125 $Y=1.557
+ $X2=7.2 $Y2=1.557
r72 37 39 31.4348 $w=3.45e-07 $l=2.25e-07 $layer=POLY_cond $X=6.9 $Y=1.557
+ $X2=7.125 $Y2=1.557
r73 37 38 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.9
+ $Y=1.515 $X2=6.9 $Y2=1.515
r74 35 37 28.6406 $w=3.45e-07 $l=2.05e-07 $layer=POLY_cond $X=6.695 $Y=1.557
+ $X2=6.9 $Y2=1.557
r75 31 44 10.4783 $w=3.45e-07 $l=9.3675e-08 $layer=POLY_cond $X=7.63 $Y=1.515
+ $X2=7.555 $Y2=1.557
r76 31 33 50.7098 $w=3.3e-07 $l=2.9e-07 $layer=POLY_cond $X=7.63 $Y=1.515
+ $X2=7.92 $Y2=1.515
r77 27 33 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=7.92
+ $Y=1.515 $X2=7.92 $Y2=1.515
r78 26 27 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=7.44 $Y=1.565
+ $X2=7.92 $Y2=1.565
r79 26 43 5.3602 $w=4.28e-07 $l=2e-07 $layer=LI1_cond $X=7.44 $Y=1.565 $X2=7.24
+ $Y2=1.565
r80 25 43 7.50428 $w=4.28e-07 $l=2.8e-07 $layer=LI1_cond $X=6.96 $Y=1.565
+ $X2=7.24 $Y2=1.565
r81 25 38 1.60806 $w=4.28e-07 $l=6e-08 $layer=LI1_cond $X=6.96 $Y=1.565 $X2=6.9
+ $Y2=1.565
r82 23 33 20.9834 $w=3.3e-07 $l=1.2e-07 $layer=POLY_cond $X=8.04 $Y=1.515
+ $X2=7.92 $Y2=1.515
r83 23 24 5.03009 $w=3.3e-07 $l=1.08995e-07 $layer=POLY_cond $X=8.04 $Y=1.515
+ $X2=8.13 $Y2=1.557
r84 19 24 37.0704 $w=1.5e-07 $l=2.14369e-07 $layer=POLY_cond $X=8.145 $Y=1.35
+ $X2=8.13 $Y2=1.557
r85 19 21 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=8.145 $Y=1.35
+ $X2=8.145 $Y2=0.74
r86 16 24 37.0704 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=8.13 $Y=1.765
+ $X2=8.13 $Y2=1.557
r87 16 18 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=8.13 $Y=1.765
+ $X2=8.13 $Y2=2.4
r88 12 44 22.2839 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=7.555 $Y=1.35
+ $X2=7.555 $Y2=1.557
r89 12 14 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=7.555 $Y=1.35
+ $X2=7.555 $Y2=0.74
r90 9 40 22.2839 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=7.2 $Y=1.765 $X2=7.2
+ $Y2=1.557
r91 9 11 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=7.2 $Y=1.765 $X2=7.2
+ $Y2=2.4
r92 5 39 22.2839 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=7.125 $Y=1.35
+ $X2=7.125 $Y2=1.557
r93 5 7 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=7.125 $Y=1.35
+ $X2=7.125 $Y2=0.74
r94 1 35 22.2839 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=6.695 $Y=1.35
+ $X2=6.695 $Y2=1.557
r95 1 3 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=6.695 $Y=1.35
+ $X2=6.695 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HS__NAND4_4%VPWR 1 2 3 4 5 18 20 24 26 28 30 32 33 42 61
+ 64 71 82 85
r66 84 85 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=3.33 $X2=8.4
+ $Y2=3.33
r67 81 82 13.5255 $w=1.123e-06 $l=1.65e-07 $layer=LI1_cond $X=6.975 $Y=2.852
+ $X2=7.14 $Y2=2.852
r68 78 81 0.162667 $w=1.123e-06 $l=1.5e-08 $layer=LI1_cond $X=6.96 $Y=2.852
+ $X2=6.975 $Y2=2.852
r69 78 79 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r70 76 79 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6 $Y=3.33 $X2=6.96
+ $Y2=3.33
r71 75 78 10.4107 $w=1.123e-06 $l=9.6e-07 $layer=LI1_cond $X=6 $Y=2.852 $X2=6.96
+ $Y2=2.852
r72 75 76 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r73 73 75 4.17511 $w=1.123e-06 $l=3.85e-07 $layer=LI1_cond $X=5.615 $Y=2.852
+ $X2=6 $Y2=2.852
r74 70 76 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=3.33 $X2=6
+ $Y2=3.33
r75 69 73 1.03022 $w=1.123e-06 $l=9.5e-08 $layer=LI1_cond $X=5.52 $Y=2.852
+ $X2=5.615 $Y2=2.852
r76 69 71 12.4953 $w=1.123e-06 $l=7e-08 $layer=LI1_cond $X=5.52 $Y=2.852
+ $X2=5.45 $Y2=2.852
r77 69 70 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r78 65 67 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=3.6 $Y2=3.33
r79 64 67 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r80 64 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r81 62 67 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.6 $Y2=3.33
r82 61 62 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r83 56 59 2.93013 $w=1.374e-06 $l=3.3e-07 $layer=LI1_cond $X=1.2 $Y=2.682
+ $X2=1.53 $Y2=2.682
r84 56 57 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r85 53 56 4.21761 $w=1.374e-06 $l=4.75e-07 $layer=LI1_cond $X=0.725 $Y=2.682
+ $X2=1.2 $Y2=2.682
r86 51 53 3.55167 $w=1.374e-06 $l=4e-07 $layer=LI1_cond $X=0.325 $Y=2.682
+ $X2=0.725 $Y2=2.682
r87 49 57 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=1.2 $Y2=3.33
r88 48 51 0.754731 $w=1.374e-06 $l=8.5e-08 $layer=LI1_cond $X=0.24 $Y=2.682
+ $X2=0.325 $Y2=2.682
r89 48 49 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r90 46 85 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=3.33
+ $X2=8.4 $Y2=3.33
r91 46 79 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=7.92 $Y=3.33
+ $X2=6.96 $Y2=3.33
r92 45 82 50.8877 $w=1.68e-07 $l=7.8e-07 $layer=LI1_cond $X=7.92 $Y=3.33
+ $X2=7.14 $Y2=3.33
r93 45 46 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r94 42 84 4.72267 $w=1.7e-07 $l=2.25e-07 $layer=LI1_cond $X=8.19 $Y=3.33
+ $X2=8.415 $Y2=3.33
r95 42 45 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=8.19 $Y=3.33 $X2=7.92
+ $Y2=3.33
r96 41 70 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=5.52 $Y2=3.33
r97 40 71 58.0642 $w=1.68e-07 $l=8.9e-07 $layer=LI1_cond $X=4.56 $Y=3.33
+ $X2=5.45 $Y2=3.33
r98 40 41 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r99 38 64 15.5046 $w=1.7e-07 $l=4.5e-07 $layer=LI1_cond $X=4.5 $Y=3.33 $X2=4.05
+ $Y2=3.33
r100 38 40 3.91444 $w=1.68e-07 $l=6e-08 $layer=LI1_cond $X=4.5 $Y=3.33 $X2=4.56
+ $Y2=3.33
r101 36 62 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r102 36 57 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.2 $Y2=3.33
r103 35 36 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r104 33 59 14.335 $w=1.374e-06 $l=7.05453e-07 $layer=LI1_cond $X=1.65 $Y=3.33
+ $X2=1.53 $Y2=2.682
r105 33 35 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=1.65 $Y=3.33
+ $X2=2.16 $Y2=3.33
r106 32 61 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.32 $Y=3.33
+ $X2=2.485 $Y2=3.33
r107 32 35 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=2.32 $Y=3.33
+ $X2=2.16 $Y2=3.33
r108 30 41 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=4.32 $Y=3.33
+ $X2=4.56 $Y2=3.33
r109 30 65 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=4.32 $Y=3.33
+ $X2=4.08 $Y2=3.33
r110 26 84 3.0435 $w=3.3e-07 $l=1.11018e-07 $layer=LI1_cond $X=8.355 $Y=3.245
+ $X2=8.415 $Y2=3.33
r111 26 28 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=8.355 $Y=3.245
+ $X2=8.355 $Y2=2.415
r112 22 64 3.34993 $w=9e-07 $l=8.5e-08 $layer=LI1_cond $X=4.05 $Y=3.245 $X2=4.05
+ $Y2=3.33
r113 22 24 11.2511 $w=8.98e-07 $l=8.3e-07 $layer=LI1_cond $X=4.05 $Y=3.245
+ $X2=4.05 $Y2=2.415
r114 21 61 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.65 $Y=3.33
+ $X2=2.485 $Y2=3.33
r115 20 64 15.5046 $w=1.7e-07 $l=4.5e-07 $layer=LI1_cond $X=3.6 $Y=3.33 $X2=4.05
+ $Y2=3.33
r116 20 21 61.9786 $w=1.68e-07 $l=9.5e-07 $layer=LI1_cond $X=3.6 $Y=3.33
+ $X2=2.65 $Y2=3.33
r117 16 61 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.485 $Y=3.245
+ $X2=2.485 $Y2=3.33
r118 16 18 27.5888 $w=3.28e-07 $l=7.9e-07 $layer=LI1_cond $X=2.485 $Y=3.245
+ $X2=2.485 $Y2=2.455
r119 5 28 300 $w=1.7e-07 $l=6.45659e-07 $layer=licon1_PDIFF $count=2 $X=8.205
+ $Y=1.84 $X2=8.355 $Y2=2.415
r120 4 81 120 $w=1.7e-07 $l=1.77436e-06 $layer=licon1_PDIFF $count=5 $X=5.465
+ $Y=1.84 $X2=6.975 $Y2=2.415
r121 4 73 120 $w=1.7e-07 $l=6.45659e-07 $layer=licon1_PDIFF $count=5 $X=5.465
+ $Y=1.84 $X2=5.615 $Y2=2.415
r122 3 24 150 $w=1.7e-07 $l=9.65609e-07 $layer=licon1_PDIFF $count=4 $X=3.615
+ $Y=1.84 $X2=4.335 $Y2=2.415
r123 2 18 300 $w=1.7e-07 $l=6.85912e-07 $layer=licon1_PDIFF $count=2 $X=2.335
+ $Y=1.84 $X2=2.485 $Y2=2.455
r124 1 59 200 $w=1.7e-07 $l=1.6745e-06 $layer=licon1_PDIFF $count=3 $X=0.135
+ $Y=1.84 $X2=1.53 $Y2=2.455
r125 1 53 200 $w=1.7e-07 $l=1.23526e-06 $layer=licon1_PDIFF $count=3 $X=0.135
+ $Y=1.84 $X2=0.725 $Y2=2.815
r126 1 53 200 $w=1.7e-07 $l=7.14388e-07 $layer=licon1_PDIFF $count=3 $X=0.135
+ $Y=1.84 $X2=0.725 $Y2=2.115
r127 1 51 200 $w=1.7e-07 $l=7.03616e-07 $layer=licon1_PDIFF $count=3 $X=0.135
+ $Y=1.84 $X2=0.325 $Y2=2.455
.ends

.subckt PM_SKY130_FD_SC_HS__NAND4_4%Y 1 2 3 4 5 6 19 21 23 27 29 33 35 38 41 43
+ 45 50 52 56 59 60 63 64
r97 63 64 18.5393 $w=2.28e-07 $l=3.7e-07 $layer=LI1_cond $X=8.4 $Y=1.295 $X2=8.4
+ $Y2=1.665
r98 62 64 14.2803 $w=2.28e-07 $l=2.85e-07 $layer=LI1_cond $X=8.4 $Y=1.95 $X2=8.4
+ $Y2=1.665
r99 61 63 8.26753 $w=2.28e-07 $l=1.65e-07 $layer=LI1_cond $X=8.4 $Y=1.13 $X2=8.4
+ $Y2=1.295
r100 58 60 4.02231 $w=3.28e-07 $l=9.5e-08 $layer=LI1_cond $X=7.85 $Y=0.965
+ $X2=7.945 $Y2=0.965
r101 58 59 4.02231 $w=3.28e-07 $l=9.5e-08 $layer=LI1_cond $X=7.85 $Y=0.965
+ $X2=7.755 $Y2=0.965
r102 46 56 13.5574 $w=1.7e-07 $l=3.45e-07 $layer=LI1_cond $X=8.01 $Y=2.035
+ $X2=7.665 $Y2=2.035
r103 45 62 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=8.285 $Y=2.035
+ $X2=8.4 $Y2=1.95
r104 45 46 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=8.285 $Y=2.035
+ $X2=8.01 $Y2=2.035
r105 43 61 6.8319 $w=2.5e-07 $l=1.73205e-07 $layer=LI1_cond $X=8.285 $Y=1.005
+ $X2=8.4 $Y2=1.13
r106 43 60 15.6732 $w=2.48e-07 $l=3.4e-07 $layer=LI1_cond $X=8.285 $Y=1.005
+ $X2=7.945 $Y2=1.005
r107 39 56 2.83173 $w=6.9e-07 $l=8.5e-08 $layer=LI1_cond $X=7.665 $Y=2.12
+ $X2=7.665 $Y2=2.035
r108 39 41 5.11367 $w=6.88e-07 $l=2.95e-07 $layer=LI1_cond $X=7.665 $Y=2.12
+ $X2=7.665 $Y2=2.415
r109 38 54 4.23145 $w=3.08e-07 $l=1.13248e-07 $layer=LI1_cond $X=7.005 $Y=1.005
+ $X2=6.91 $Y2=0.965
r110 38 59 34.5733 $w=2.48e-07 $l=7.5e-07 $layer=LI1_cond $X=7.005 $Y=1.005
+ $X2=7.755 $Y2=1.005
r111 36 52 12.6759 $w=1.7e-07 $l=3.05e-07 $layer=LI1_cond $X=5.28 $Y=2.035
+ $X2=4.975 $Y2=2.035
r112 35 56 13.5574 $w=1.7e-07 $l=3.45e-07 $layer=LI1_cond $X=7.32 $Y=2.035
+ $X2=7.665 $Y2=2.035
r113 35 36 133.091 $w=1.68e-07 $l=2.04e-06 $layer=LI1_cond $X=7.32 $Y=2.035
+ $X2=5.28 $Y2=2.035
r114 31 52 2.55884 $w=6.1e-07 $l=8.5e-08 $layer=LI1_cond $X=4.975 $Y=2.12
+ $X2=4.975 $Y2=2.035
r115 31 33 5.78431 $w=6.08e-07 $l=2.95e-07 $layer=LI1_cond $X=4.975 $Y=2.12
+ $X2=4.975 $Y2=2.415
r116 30 50 12.6759 $w=1.7e-07 $l=3.05e-07 $layer=LI1_cond $X=3.43 $Y=2.035
+ $X2=3.125 $Y2=2.035
r117 29 52 12.6759 $w=1.7e-07 $l=3.05e-07 $layer=LI1_cond $X=4.67 $Y=2.035
+ $X2=4.975 $Y2=2.035
r118 29 30 80.8984 $w=1.68e-07 $l=1.24e-06 $layer=LI1_cond $X=4.67 $Y=2.035
+ $X2=3.43 $Y2=2.035
r119 25 50 2.55884 $w=6.1e-07 $l=8.5e-08 $layer=LI1_cond $X=3.125 $Y=2.12
+ $X2=3.125 $Y2=2.035
r120 25 27 5.78431 $w=6.08e-07 $l=2.95e-07 $layer=LI1_cond $X=3.125 $Y=2.12
+ $X2=3.125 $Y2=2.415
r121 24 48 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.15 $Y=2.035
+ $X2=1.985 $Y2=2.035
r122 23 50 12.6759 $w=1.7e-07 $l=3.05e-07 $layer=LI1_cond $X=2.82 $Y=2.035
+ $X2=3.125 $Y2=2.035
r123 23 24 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.82 $Y=2.035
+ $X2=2.15 $Y2=2.035
r124 19 48 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.985 $Y=2.12
+ $X2=1.985 $Y2=2.035
r125 19 21 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=1.985 $Y=2.12
+ $X2=1.985 $Y2=2.415
r126 6 56 300 $w=1.7e-07 $l=7.20937e-07 $layer=licon1_PDIFF $count=2 $X=7.275
+ $Y=1.84 $X2=7.905 $Y2=2.035
r127 6 41 150 $w=1.7e-07 $l=8.71292e-07 $layer=licon1_PDIFF $count=4 $X=7.275
+ $Y=1.84 $X2=7.905 $Y2=2.415
r128 5 52 300 $w=1.7e-07 $l=6.19879e-07 $layer=licon1_PDIFF $count=2 $X=4.635
+ $Y=1.84 $X2=5.165 $Y2=2.035
r129 5 33 150 $w=1.7e-07 $l=7.97104e-07 $layer=licon1_PDIFF $count=4 $X=4.635
+ $Y=1.84 $X2=5.165 $Y2=2.415
r130 4 50 300 $w=1.7e-07 $l=6.19879e-07 $layer=licon1_PDIFF $count=2 $X=2.785
+ $Y=1.84 $X2=3.315 $Y2=2.035
r131 4 27 150 $w=1.7e-07 $l=7.97104e-07 $layer=licon1_PDIFF $count=4 $X=2.785
+ $Y=1.84 $X2=3.315 $Y2=2.415
r132 3 48 600 $w=1.7e-07 $l=2.59374e-07 $layer=licon1_PDIFF $count=1 $X=1.835
+ $Y=1.84 $X2=1.985 $Y2=2.035
r133 3 21 300 $w=1.7e-07 $l=6.45659e-07 $layer=licon1_PDIFF $count=2 $X=1.835
+ $Y=1.84 $X2=1.985 $Y2=2.415
r134 2 58 182 $w=1.7e-07 $l=6.96366e-07 $layer=licon1_NDIFF $count=1 $X=7.63
+ $Y=0.37 $X2=7.85 $Y2=0.965
r135 1 54 182 $w=1.7e-07 $l=6.61306e-07 $layer=licon1_NDIFF $count=1 $X=6.77
+ $Y=0.37 $X2=6.91 $Y2=0.965
.ends

.subckt PM_SKY130_FD_SC_HS__NAND4_4%A_27_74# 1 2 3 4 5 18 20 21 24 26 28 31 36
+ 38
r62 34 36 30.0334 $w=3.28e-07 $l=8.6e-07 $layer=LI1_cond $X=3.34 $Y=0.515
+ $X2=4.2 $Y2=0.515
r63 32 40 3.40825 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=2.575 $Y=0.515
+ $X2=2.41 $Y2=0.515
r64 32 34 26.7157 $w=3.28e-07 $l=7.65e-07 $layer=LI1_cond $X=2.575 $Y=0.515
+ $X2=3.34 $Y2=0.515
r65 29 31 1.57151 $w=3.28e-07 $l=4.5e-08 $layer=LI1_cond $X=2.41 $Y=1.01
+ $X2=2.41 $Y2=0.965
r66 28 40 3.40825 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=2.41 $Y=0.68
+ $X2=2.41 $Y2=0.515
r67 28 31 9.95292 $w=3.28e-07 $l=2.85e-07 $layer=LI1_cond $X=2.41 $Y=0.68
+ $X2=2.41 $Y2=0.965
r68 27 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.445 $Y=1.095
+ $X2=1.28 $Y2=1.095
r69 26 29 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.245 $Y=1.095
+ $X2=2.41 $Y2=1.01
r70 26 27 52.1925 $w=1.68e-07 $l=8e-07 $layer=LI1_cond $X=2.245 $Y=1.095
+ $X2=1.445 $Y2=1.095
r71 22 38 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.28 $Y=1.01 $X2=1.28
+ $Y2=1.095
r72 22 24 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=1.28 $Y=1.01
+ $X2=1.28 $Y2=0.515
r73 20 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.115 $Y=1.095
+ $X2=1.28 $Y2=1.095
r74 20 21 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.115 $Y=1.095
+ $X2=0.445 $Y2=1.095
r75 16 21 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.28 $Y=1.01
+ $X2=0.445 $Y2=1.095
r76 16 18 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=0.28 $Y=1.01
+ $X2=0.28 $Y2=0.515
r77 5 36 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=4.06
+ $Y=0.37 $X2=4.2 $Y2=0.515
r78 4 34 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=3.2
+ $Y=0.37 $X2=3.34 $Y2=0.515
r79 3 40 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=2.27
+ $Y=0.37 $X2=2.41 $Y2=0.515
r80 3 31 182 $w=1.7e-07 $l=6.61306e-07 $layer=licon1_NDIFF $count=1 $X=2.27
+ $Y=0.37 $X2=2.41 $Y2=0.965
r81 2 24 91 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=2 $X=1.07
+ $Y=0.37 $X2=1.28 $Y2=0.515
r82 1 18 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__NAND4_4%VGND 1 2 9 11 15 17 19 29 30 33 36
r68 36 37 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r69 34 37 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r70 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r71 29 30 1.32857 $w=1.7e-07 $l=1.19e-06 $layer=mcon $count=7 $X=8.4 $Y=0
+ $X2=8.4 $Y2=0
r72 27 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.68
+ $Y2=0
r73 26 29 407.102 $w=1.68e-07 $l=6.24e-06 $layer=LI1_cond $X=2.16 $Y=0 $X2=8.4
+ $Y2=0
r74 26 27 1.32857 $w=1.7e-07 $l=1.19e-06 $layer=mcon $count=7 $X=2.16 $Y=0
+ $X2=2.16 $Y2=0
r75 24 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.945 $Y=0 $X2=1.78
+ $Y2=0
r76 24 26 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=1.945 $Y=0 $X2=2.16
+ $Y2=0
r77 22 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r78 21 22 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r79 19 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.615 $Y=0 $X2=0.78
+ $Y2=0
r80 19 21 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=0.615 $Y=0 $X2=0.24
+ $Y2=0
r81 17 30 1.13724 $w=4.9e-07 $l=4.08e-06 $layer=MET1_cond $X=4.32 $Y=0 $X2=8.4
+ $Y2=0
r82 17 27 0.602067 $w=4.9e-07 $l=2.16e-06 $layer=MET1_cond $X=4.32 $Y=0 $X2=2.16
+ $Y2=0
r83 13 36 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.78 $Y=0.085
+ $X2=1.78 $Y2=0
r84 13 15 20.6043 $w=3.28e-07 $l=5.9e-07 $layer=LI1_cond $X=1.78 $Y=0.085
+ $X2=1.78 $Y2=0.675
r85 12 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.945 $Y=0 $X2=0.78
+ $Y2=0
r86 11 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.615 $Y=0 $X2=1.78
+ $Y2=0
r87 11 12 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.615 $Y=0 $X2=0.945
+ $Y2=0
r88 7 33 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.78 $Y=0.085 $X2=0.78
+ $Y2=0
r89 7 9 20.6043 $w=3.28e-07 $l=5.9e-07 $layer=LI1_cond $X=0.78 $Y=0.085 $X2=0.78
+ $Y2=0.675
r90 2 15 182 $w=1.7e-07 $l=3.96327e-07 $layer=licon1_NDIFF $count=1 $X=1.57
+ $Y=0.37 $X2=1.78 $Y2=0.675
r91 1 9 182 $w=1.7e-07 $l=3.96327e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.37 $X2=0.78 $Y2=0.675
.ends

.subckt PM_SKY130_FD_SC_HS__NAND4_4%A_554_74# 1 2 3 4 13 21 23 26 27
c40 13 0 7.27676e-20 $X=3.795 $Y=0.99
r41 25 27 4.02231 $w=3.28e-07 $l=9.5e-08 $layer=LI1_cond $X=5.19 $Y=0.965
+ $X2=5.285 $Y2=0.965
r42 25 26 4.02231 $w=3.28e-07 $l=9.5e-08 $layer=LI1_cond $X=5.19 $Y=0.965
+ $X2=5.095 $Y2=0.965
r43 23 26 53.4734 $w=2.48e-07 $l=1.16e-06 $layer=LI1_cond $X=3.935 $Y=1.005
+ $X2=5.095 $Y2=1.005
r44 21 29 4.23145 $w=3.08e-07 $l=1.13248e-07 $layer=LI1_cond $X=5.955 $Y=1.005
+ $X2=6.05 $Y2=0.965
r45 21 27 30.8855 $w=2.48e-07 $l=6.7e-07 $layer=LI1_cond $X=5.955 $Y=1.005
+ $X2=5.285 $Y2=1.005
r46 15 18 35.3965 $w=2.78e-07 $l=8.6e-07 $layer=LI1_cond $X=2.91 $Y=0.99
+ $X2=3.77 $Y2=0.99
r47 13 23 5.9212 $w=2.78e-07 $l=1.4e-07 $layer=LI1_cond $X=3.795 $Y=0.99
+ $X2=3.935 $Y2=0.99
r48 13 18 1.02897 $w=2.78e-07 $l=2.5e-08 $layer=LI1_cond $X=3.795 $Y=0.99
+ $X2=3.77 $Y2=0.99
r49 4 29 182 $w=1.7e-07 $l=6.61306e-07 $layer=licon1_NDIFF $count=1 $X=5.91
+ $Y=0.37 $X2=6.05 $Y2=0.965
r50 3 25 182 $w=1.7e-07 $l=6.61306e-07 $layer=licon1_NDIFF $count=1 $X=5.05
+ $Y=0.37 $X2=5.19 $Y2=0.965
r51 2 18 182 $w=1.7e-07 $l=6.4622e-07 $layer=licon1_NDIFF $count=1 $X=3.63
+ $Y=0.37 $X2=3.77 $Y2=0.95
r52 1 15 182 $w=1.7e-07 $l=6.4622e-07 $layer=licon1_NDIFF $count=1 $X=2.77
+ $Y=0.37 $X2=2.91 $Y2=0.95
.ends

.subckt PM_SKY130_FD_SC_HS__NAND4_4%A_923_74# 1 2 3 4 5 22 24 31 32 35 36 39 40
+ 41
r62 41 44 3.84148 $w=3.28e-07 $l=1.1e-07 $layer=LI1_cond $X=8.36 $Y=0.435
+ $X2=8.36 $Y2=0.545
r63 38 40 8.51103 $w=3.58e-07 $l=1.65e-07 $layer=LI1_cond $X=7.34 $Y=0.53
+ $X2=7.505 $Y2=0.53
r64 38 39 8.51103 $w=3.58e-07 $l=1.65e-07 $layer=LI1_cond $X=7.34 $Y=0.53
+ $X2=7.175 $Y2=0.53
r65 36 39 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=6.645 $Y=0.435
+ $X2=7.175 $Y2=0.435
r66 34 36 8.51103 $w=3.58e-07 $l=1.65e-07 $layer=LI1_cond $X=6.48 $Y=0.53
+ $X2=6.645 $Y2=0.53
r67 34 35 8.51103 $w=3.58e-07 $l=1.65e-07 $layer=LI1_cond $X=6.48 $Y=0.53
+ $X2=6.315 $Y2=0.53
r68 32 35 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=5.785 $Y=0.435
+ $X2=6.315 $Y2=0.435
r69 30 32 8.51103 $w=3.58e-07 $l=1.65e-07 $layer=LI1_cond $X=5.62 $Y=0.53
+ $X2=5.785 $Y2=0.53
r70 30 31 8.51103 $w=3.58e-07 $l=1.65e-07 $layer=LI1_cond $X=5.62 $Y=0.53
+ $X2=5.455 $Y2=0.53
r71 24 27 3.84148 $w=3.28e-07 $l=1.1e-07 $layer=LI1_cond $X=4.76 $Y=0.435
+ $X2=4.76 $Y2=0.545
r72 22 41 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.195 $Y=0.435
+ $X2=8.36 $Y2=0.435
r73 22 40 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=8.195 $Y=0.435
+ $X2=7.505 $Y2=0.435
r74 17 24 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.925 $Y=0.435
+ $X2=4.76 $Y2=0.435
r75 17 31 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=4.925 $Y=0.435
+ $X2=5.455 $Y2=0.435
r76 5 44 182 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_NDIFF $count=1 $X=8.22
+ $Y=0.37 $X2=8.36 $Y2=0.545
r77 4 38 182 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_NDIFF $count=1 $X=7.2
+ $Y=0.37 $X2=7.34 $Y2=0.545
r78 3 34 182 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_NDIFF $count=1 $X=6.34
+ $Y=0.37 $X2=6.48 $Y2=0.545
r79 2 30 182 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_NDIFF $count=1 $X=5.48
+ $Y=0.37 $X2=5.62 $Y2=0.545
r80 1 27 182 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_NDIFF $count=1 $X=4.615
+ $Y=0.37 $X2=4.76 $Y2=0.545
.ends

