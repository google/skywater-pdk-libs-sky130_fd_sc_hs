* File: sky130_fd_sc_hs__sdfrbp_1.pex.spice
* Created: Thu Aug 27 21:08:19 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HS__SDFRBP_1%A_27_74# 1 2 7 9 10 12 15 18 21 22 24 26 31
+ 33
c80 33 0 4.33637e-20 $X=2.53 $Y=1.995
r81 33 36 4.88915 $w=3.28e-07 $l=1.4e-07 $layer=LI1_cond $X=2.53 $Y=1.995
+ $X2=2.53 $Y2=2.135
r82 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.53
+ $Y=1.995 $X2=2.53 $Y2=1.995
r83 30 31 12.4206 $w=9.23e-07 $l=1.65e-07 $layer=LI1_cond $X=0.89 $Y=2.512
+ $X2=1.055 $Y2=2.512
r84 24 36 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.365 $Y=2.135
+ $X2=2.53 $Y2=2.135
r85 24 31 85.4652 $w=1.68e-07 $l=1.31e-06 $layer=LI1_cond $X=2.365 $Y=2.135
+ $X2=1.055 $Y2=2.135
r86 21 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.23
+ $Y=1.145 $X2=1.23 $Y2=1.145
r87 19 26 0.221902 $w=3.3e-07 $l=1.25e-07 $layer=LI1_cond $X=0.365 $Y=1.145
+ $X2=0.24 $Y2=1.145
r88 19 21 30.208 $w=3.28e-07 $l=8.65e-07 $layer=LI1_cond $X=0.365 $Y=1.145
+ $X2=1.23 $Y2=1.145
r89 18 30 9.10054 $w=9.23e-07 $l=6.9e-07 $layer=LI1_cond $X=0.2 $Y=2.512
+ $X2=0.89 $Y2=2.512
r90 17 26 7.38875 $w=2.1e-07 $l=1.83916e-07 $layer=LI1_cond $X=0.2 $Y=1.31
+ $X2=0.24 $Y2=1.145
r91 17 18 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=0.2 $Y=1.31 $X2=0.2
+ $Y2=2.05
r92 13 26 7.38875 $w=2.1e-07 $l=1.65e-07 $layer=LI1_cond $X=0.24 $Y=0.98
+ $X2=0.24 $Y2=1.145
r93 13 15 18.4391 $w=2.48e-07 $l=4e-07 $layer=LI1_cond $X=0.24 $Y=0.98 $X2=0.24
+ $Y2=0.58
r94 10 34 52.2586 $w=2.99e-07 $l=2.7157e-07 $layer=POLY_cond $X=2.485 $Y=2.245
+ $X2=2.53 $Y2=1.995
r95 10 12 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=2.485 $Y=2.245
+ $X2=2.485 $Y2=2.64
r96 7 22 45.5222 $w=2.7e-07 $l=3.27261e-07 $layer=POLY_cond $X=1.485 $Y=0.98
+ $X2=1.23 $Y2=1.145
r97 7 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.485 $Y=0.98
+ $X2=1.485 $Y2=0.66
r98 2 30 150 $w=1.7e-07 $l=8.24318e-07 $layer=licon1_PDIFF $count=4 $X=0.135
+ $Y=2.32 $X2=0.89 $Y2=2.465
r99 1 15 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_HS__SDFRBP_1%SCE 3 6 7 9 11 12 14 17 19 20 23 24 28 29
+ 30 35 43 48 57 59
c89 24 0 1.81012e-19 $X=2.56 $Y=1.425
r90 48 57 2.36399 $w=3.88e-07 $l=8e-08 $layer=LI1_cond $X=1.6 $Y=1.685 $X2=1.68
+ $Y2=1.685
r91 41 43 28.8521 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.45 $Y=1.715
+ $X2=1.615 $Y2=1.715
r92 41 42 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.45
+ $Y=1.715 $X2=1.45 $Y2=1.715
r93 39 41 58.5785 $w=3.3e-07 $l=3.35e-07 $layer=POLY_cond $X=1.115 $Y=1.715
+ $X2=1.45 $Y2=1.715
r94 35 39 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=1.025 $Y=1.715
+ $X2=1.115 $Y2=1.715
r95 35 37 44.5896 $w=3.3e-07 $l=2.55e-07 $layer=POLY_cond $X=1.025 $Y=1.715
+ $X2=0.77 $Y2=1.715
r96 30 59 7.07103 $w=3.88e-07 $l=1.13e-07 $layer=LI1_cond $X=1.682 $Y=1.685
+ $X2=1.795 $Y2=1.685
r97 30 57 0.0590996 $w=3.88e-07 $l=2e-09 $layer=LI1_cond $X=1.682 $Y=1.685
+ $X2=1.68 $Y2=1.685
r98 30 48 0.0886495 $w=3.88e-07 $l=3e-09 $layer=LI1_cond $X=1.597 $Y=1.685
+ $X2=1.6 $Y2=1.685
r99 30 42 4.34382 $w=3.88e-07 $l=1.47e-07 $layer=LI1_cond $X=1.597 $Y=1.685
+ $X2=1.45 $Y2=1.685
r100 29 42 7.38745 $w=3.88e-07 $l=2.5e-07 $layer=LI1_cond $X=1.2 $Y=1.685
+ $X2=1.45 $Y2=1.685
r101 28 29 14.1839 $w=3.88e-07 $l=4.8e-07 $layer=LI1_cond $X=0.72 $Y=1.685
+ $X2=1.2 $Y2=1.685
r102 28 37 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=0.77
+ $Y=1.715 $X2=0.77 $Y2=1.715
r103 24 46 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.56 $Y=1.425
+ $X2=2.56 $Y2=1.26
r104 23 26 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=2.56 $Y=1.425
+ $X2=2.56 $Y2=1.575
r105 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.56
+ $Y=1.425 $X2=2.56 $Y2=1.425
r106 20 26 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.395 $Y=1.575
+ $X2=2.56 $Y2=1.575
r107 20 59 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=2.395 $Y=1.575
+ $X2=1.795 $Y2=1.575
r108 19 37 34.9723 $w=3.3e-07 $l=2e-07 $layer=POLY_cond $X=0.57 $Y=1.715
+ $X2=0.77 $Y2=1.715
r109 17 46 289.713 $w=1.5e-07 $l=5.65e-07 $layer=POLY_cond $X=2.65 $Y=0.695
+ $X2=2.65 $Y2=1.26
r110 12 14 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=1.615 $Y=2.245
+ $X2=1.615 $Y2=2.64
r111 11 12 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=1.615 $Y=2.155
+ $X2=1.615 $Y2=2.245
r112 10 43 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.615 $Y=1.88
+ $X2=1.615 $Y2=1.715
r113 10 11 106.895 $w=1.8e-07 $l=2.75e-07 $layer=POLY_cond $X=1.615 $Y=1.88
+ $X2=1.615 $Y2=2.155
r114 7 9 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=1.115 $Y=2.245
+ $X2=1.115 $Y2=2.64
r115 6 7 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=1.115 $Y=2.155
+ $X2=1.115 $Y2=2.245
r116 5 39 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.115 $Y=1.88
+ $X2=1.115 $Y2=1.715
r117 5 6 106.895 $w=1.8e-07 $l=2.75e-07 $layer=POLY_cond $X=1.115 $Y=1.88
+ $X2=1.115 $Y2=2.155
r118 1 19 32.1775 $w=3.3e-07 $l=1.98997e-07 $layer=POLY_cond $X=0.495 $Y=1.55
+ $X2=0.57 $Y2=1.715
r119 1 3 497.383 $w=1.5e-07 $l=9.7e-07 $layer=POLY_cond $X=0.495 $Y=1.55
+ $X2=0.495 $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_HS__SDFRBP_1%D 3 5 6 8 9 12 13 14
c44 13 0 1.81012e-19 $X=1.935 $Y=1.145
c45 6 0 4.33637e-20 $X=2.035 $Y=2.245
r46 12 15 40.8147 $w=3.55e-07 $l=1.65e-07 $layer=POLY_cond $X=1.947 $Y=1.145
+ $X2=1.947 $Y2=1.31
r47 12 14 46.504 $w=3.55e-07 $l=1.65e-07 $layer=POLY_cond $X=1.947 $Y=1.145
+ $X2=1.947 $Y2=0.98
r48 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.935
+ $Y=1.145 $X2=1.935 $Y2=1.145
r49 9 13 6.1 $w=4.98e-07 $l=2.55e-07 $layer=LI1_cond $X=1.68 $Y=1.06 $X2=1.935
+ $Y2=1.06
r50 6 8 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=2.035 $Y=2.245
+ $X2=2.035 $Y2=2.64
r51 5 6 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=2.035 $Y=2.155 $X2=2.035
+ $Y2=2.245
r52 5 15 328.46 $w=1.8e-07 $l=8.45e-07 $layer=POLY_cond $X=2.035 $Y=2.155
+ $X2=2.035 $Y2=1.31
r53 3 14 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.99 $Y=0.66 $X2=1.99
+ $Y2=0.98
.ends

.subckt PM_SKY130_FD_SC_HS__SDFRBP_1%SCD 1 3 6 10 11 12 16
c44 11 0 1.32707e-19 $X=3.12 $Y=1.665
r45 11 12 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=3.1 $Y=1.605 $X2=3.1
+ $Y2=2.035
r46 11 16 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.1
+ $Y=1.605 $X2=3.1 $Y2=1.605
r47 10 16 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=3.1 $Y=1.945 $X2=3.1
+ $Y2=1.605
r48 9 16 41.8716 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.1 $Y=1.44 $X2=3.1
+ $Y2=1.605
r49 6 9 382.011 $w=1.5e-07 $l=7.45e-07 $layer=POLY_cond $X=3.04 $Y=0.695
+ $X2=3.04 $Y2=1.44
r50 1 10 55.1908 $w=2.62e-07 $l=3.3541e-07 $layer=POLY_cond $X=3.025 $Y=2.245
+ $X2=3.1 $Y2=1.945
r51 1 3 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=3.025 $Y=2.245
+ $X2=3.025 $Y2=2.64
.ends

.subckt PM_SKY130_FD_SC_HS__SDFRBP_1%RESET_B 3 5 7 10 12 14 16 19 23 30 36 38 39
+ 40 41 42 43 51 54 55 58 61 63 64 65
c220 64 0 1.5378e-19 $X=10.9 $Y=1.845
c221 63 0 2.44776e-20 $X=10.9 $Y=1.845
c222 58 0 1.32707e-19 $X=3.595 $Y=2.032
c223 39 0 8.18376e-20 $X=10.81 $Y=2.37
c224 36 0 6.47027e-20 $X=10.81 $Y=1.335
r225 64 76 5.91795 $w=3.68e-07 $l=1.9e-07 $layer=LI1_cond $X=10.88 $Y=1.845
+ $X2=10.88 $Y2=2.035
r226 63 66 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=10.9 $Y=1.845
+ $X2=10.9 $Y2=2.01
r227 63 65 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=10.9 $Y=1.845
+ $X2=10.9 $Y2=1.68
r228 63 64 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.9
+ $Y=1.845 $X2=10.9 $Y2=1.845
r229 60 61 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.95
+ $Y=1.985 $X2=3.95 $Y2=1.985
r230 58 60 47.7961 $w=3.58e-07 $l=3.55e-07 $layer=POLY_cond $X=3.595 $Y=2.032
+ $X2=3.95 $Y2=2.032
r231 57 58 2.01955 $w=3.58e-07 $l=1.5e-08 $layer=POLY_cond $X=3.58 $Y=2.032
+ $X2=3.595 $Y2=2.032
r232 54 55 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.86
+ $Y=1.985 $X2=7.86 $Y2=1.985
r233 51 76 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.8 $Y=2.035
+ $X2=10.8 $Y2=2.035
r234 49 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=2.035
+ $X2=7.92 $Y2=2.035
r235 45 61 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=2.035
+ $X2=4.08 $Y2=2.035
r236 43 49 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=8.065 $Y=2.035
+ $X2=7.92 $Y2=2.035
r237 42 51 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=10.655 $Y=2.035
+ $X2=10.8 $Y2=2.035
r238 42 43 3.20544 $w=1.4e-07 $l=2.59e-06 $layer=MET1_cond $X=10.655 $Y=2.035
+ $X2=8.065 $Y2=2.035
r239 41 45 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.225 $Y=2.035
+ $X2=4.08 $Y2=2.035
r240 40 49 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=7.775 $Y=2.035
+ $X2=7.92 $Y2=2.035
r241 40 41 4.39356 $w=1.4e-07 $l=3.55e-06 $layer=MET1_cond $X=7.775 $Y=2.035
+ $X2=4.225 $Y2=2.035
r242 38 39 47.3682 $w=2.1e-07 $l=1.5e-07 $layer=POLY_cond $X=10.81 $Y=2.22
+ $X2=10.81 $Y2=2.37
r243 38 66 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=10.84 $Y=2.22
+ $X2=10.84 $Y2=2.01
r244 34 36 135.883 $w=1.5e-07 $l=2.65e-07 $layer=POLY_cond $X=10.545 $Y=1.335
+ $X2=10.81 $Y2=1.335
r245 33 54 31.475 $w=3.3e-07 $l=1.8e-07 $layer=POLY_cond $X=7.68 $Y=1.985
+ $X2=7.86 $Y2=1.985
r246 28 30 151.266 $w=1.5e-07 $l=2.95e-07 $layer=POLY_cond $X=7.31 $Y=1.145
+ $X2=7.605 $Y2=1.145
r247 24 36 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=10.81 $Y=1.41
+ $X2=10.81 $Y2=1.335
r248 24 65 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=10.81 $Y=1.41
+ $X2=10.81 $Y2=1.68
r249 23 39 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=10.795 $Y=2.655
+ $X2=10.795 $Y2=2.37
r250 17 34 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=10.545 $Y=1.26
+ $X2=10.545 $Y2=1.335
r251 17 19 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=10.545 $Y=1.26
+ $X2=10.545 $Y2=0.58
r252 16 33 45.8367 $w=1.79e-07 $l=1.80748e-07 $layer=POLY_cond $X=7.605 $Y=1.82
+ $X2=7.572 $Y2=1.985
r253 15 30 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.605 $Y=1.22
+ $X2=7.605 $Y2=1.145
r254 15 16 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=7.605 $Y=1.22
+ $X2=7.605 $Y2=1.82
r255 12 33 70.0713 $w=1.79e-07 $l=2.63363e-07 $layer=POLY_cond $X=7.555 $Y=2.24
+ $X2=7.572 $Y2=1.985
r256 12 14 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=7.555 $Y=2.24
+ $X2=7.555 $Y2=2.525
r257 8 28 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.31 $Y=1.07
+ $X2=7.31 $Y2=1.145
r258 8 10 192.287 $w=1.5e-07 $l=3.75e-07 $layer=POLY_cond $X=7.31 $Y=1.07
+ $X2=7.31 $Y2=0.695
r259 5 58 23.1716 $w=1.5e-07 $l=2.13e-07 $layer=POLY_cond $X=3.595 $Y=2.245
+ $X2=3.595 $Y2=2.032
r260 5 7 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=3.595 $Y=2.245
+ $X2=3.595 $Y2=2.64
r261 1 57 23.1716 $w=1.5e-07 $l=2.12e-07 $layer=POLY_cond $X=3.58 $Y=1.82
+ $X2=3.58 $Y2=2.032
r262 1 3 599.936 $w=1.5e-07 $l=1.17e-06 $layer=POLY_cond $X=3.58 $Y=1.82
+ $X2=3.58 $Y2=0.65
.ends

.subckt PM_SKY130_FD_SC_HS__SDFRBP_1%CLK 1 3 4 6 8 9 13
c48 13 0 1.07514e-19 $X=4.48 $Y=1.385
c49 8 0 1.5551e-19 $X=4.535 $Y=1.385
r50 12 13 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.48
+ $Y=1.385 $X2=4.48 $Y2=1.385
r51 9 13 12.4588 $w=3.68e-07 $l=4e-07 $layer=LI1_cond $X=4.08 $Y=1.365 $X2=4.48
+ $Y2=1.365
r52 8 12 9.61737 $w=3.3e-07 $l=5.5e-08 $layer=POLY_cond $X=4.535 $Y=1.385
+ $X2=4.48 $Y2=1.385
r53 4 8 100.273 $w=1.75e-07 $l=3.64966e-07 $layer=POLY_cond $X=4.645 $Y=1.745
+ $X2=4.635 $Y2=1.385
r54 4 6 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=4.645 $Y=1.745
+ $X2=4.645 $Y2=2.38
r55 1 8 46.5648 $w=1.75e-07 $l=1.77059e-07 $layer=POLY_cond $X=4.61 $Y=1.22
+ $X2=4.635 $Y2=1.385
r56 1 3 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=4.61 $Y=1.22 $X2=4.61
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HS__SDFRBP_1%A_1023_74# 1 2 8 9 11 12 16 18 20 21 22 23
+ 25 29 30 31 33 34 36 40 41 42 44 45 46 48 50 53 61 66 67 71 73
c209 67 0 1.52128e-19 $X=9.27 $Y=1.07
c210 66 0 1.89691e-19 $X=9.27 $Y=1.07
r211 67 79 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=9.27 $Y=1.07 $X2=9.27
+ $Y2=1.16
r212 66 67 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.27
+ $Y=1.07 $X2=9.27 $Y2=1.07
r213 63 66 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=8.865 $Y=0.99
+ $X2=9.27 $Y2=0.99
r214 53 54 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.67
+ $Y=2.065 $X2=9.67 $Y2=2.065
r215 51 71 0.201461 $w=2.5e-07 $l=1.15e-07 $layer=LI1_cond $X=9.63 $Y=1.575
+ $X2=9.63 $Y2=1.46
r216 51 53 22.5879 $w=2.48e-07 $l=4.9e-07 $layer=LI1_cond $X=9.63 $Y=1.575
+ $X2=9.63 $Y2=2.065
r217 50 71 18.0382 $w=2.28e-07 $l=3.6e-07 $layer=LI1_cond $X=9.27 $Y=1.46
+ $X2=9.63 $Y2=1.46
r218 50 66 9.42908 $w=3.28e-07 $l=2.7e-07 $layer=LI1_cond $X=9.27 $Y=1.345
+ $X2=9.27 $Y2=1.075
r219 48 63 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.865 $Y=0.905
+ $X2=8.865 $Y2=0.99
r220 47 48 31.3155 $w=1.68e-07 $l=4.8e-07 $layer=LI1_cond $X=8.865 $Y=0.425
+ $X2=8.865 $Y2=0.905
r221 45 47 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.78 $Y=0.34
+ $X2=8.865 $Y2=0.425
r222 45 46 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=8.78 $Y=0.34
+ $X2=8.11 $Y2=0.34
r223 43 46 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.025 $Y=0.425
+ $X2=8.11 $Y2=0.34
r224 43 44 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=8.025 $Y=0.425
+ $X2=8.025 $Y2=0.595
r225 41 44 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.94 $Y=0.68
+ $X2=8.025 $Y2=0.595
r226 41 42 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=7.94 $Y=0.68
+ $X2=7.185 $Y2=0.68
r227 40 42 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.1 $Y=0.595
+ $X2=7.185 $Y2=0.68
r228 39 40 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=7.1 $Y=0.425
+ $X2=7.1 $Y2=0.595
r229 37 76 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.055 $Y=1.74
+ $X2=6.055 $Y2=1.905
r230 37 73 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=6.055 $Y=1.74
+ $X2=6.055 $Y2=1.65
r231 36 37 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.055
+ $Y=1.74 $X2=6.055 $Y2=1.74
r232 34 58 7.95652 $w=3.45e-07 $l=3.26671e-07 $layer=LI1_cond $X=5.62 $Y=1.74
+ $X2=5.387 $Y2=1.965
r233 34 36 15.1913 $w=3.28e-07 $l=4.35e-07 $layer=LI1_cond $X=5.62 $Y=1.74
+ $X2=6.055 $Y2=1.74
r234 33 34 8.97647 $w=3.45e-07 $l=2.03101e-07 $layer=LI1_cond $X=5.535 $Y=1.575
+ $X2=5.62 $Y2=1.74
r235 32 61 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.535 $Y=1.13
+ $X2=5.535 $Y2=1.045
r236 32 33 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=5.535 $Y=1.13
+ $X2=5.535 $Y2=1.575
r237 30 39 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.015 $Y=0.34
+ $X2=7.1 $Y2=0.425
r238 30 31 104.059 $w=1.68e-07 $l=1.595e-06 $layer=LI1_cond $X=7.015 $Y=0.34
+ $X2=5.42 $Y2=0.34
r239 27 61 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=5.295 $Y=1.045
+ $X2=5.535 $Y2=1.045
r240 27 29 20.5135 $w=2.48e-07 $l=4.45e-07 $layer=LI1_cond $X=5.295 $Y=0.96
+ $X2=5.295 $Y2=0.515
r241 26 31 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=5.295 $Y=0.425
+ $X2=5.42 $Y2=0.34
r242 26 29 4.14879 $w=2.48e-07 $l=9e-08 $layer=LI1_cond $X=5.295 $Y=0.425
+ $X2=5.295 $Y2=0.515
r243 23 54 60.889 $w=3.02e-07 $l=3.46215e-07 $layer=POLY_cond $X=9.77 $Y=2.37
+ $X2=9.682 $Y2=2.065
r244 23 25 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=9.77 $Y=2.37
+ $X2=9.77 $Y2=2.655
r245 21 79 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.105 $Y=1.16
+ $X2=9.27 $Y2=1.16
r246 21 22 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=9.105 $Y=1.16
+ $X2=8.735 $Y2=1.16
r247 18 22 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=8.66 $Y=1.085
+ $X2=8.735 $Y2=1.16
r248 18 20 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=8.66 $Y=1.085
+ $X2=8.66 $Y2=0.69
r249 14 16 451.234 $w=1.5e-07 $l=8.8e-07 $layer=POLY_cond $X=6.53 $Y=1.575
+ $X2=6.53 $Y2=0.695
r250 13 73 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.22 $Y=1.65
+ $X2=6.055 $Y2=1.65
r251 12 14 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=6.455 $Y=1.65
+ $X2=6.53 $Y2=1.575
r252 12 13 120.5 $w=1.5e-07 $l=2.35e-07 $layer=POLY_cond $X=6.455 $Y=1.65
+ $X2=6.22 $Y2=1.65
r253 9 11 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=6.115 $Y=2.24
+ $X2=6.115 $Y2=2.525
r254 8 9 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=6.115 $Y=2.15 $X2=6.115
+ $Y2=2.24
r255 8 76 95.2339 $w=1.8e-07 $l=2.45e-07 $layer=POLY_cond $X=6.115 $Y=2.15
+ $X2=6.115 $Y2=1.905
r256 2 58 600 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=5.17
+ $Y=1.82 $X2=5.32 $Y2=1.965
r257 1 29 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=5.115
+ $Y=0.37 $X2=5.255 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__SDFRBP_1%A_1369_71# 1 2 9 12 13 15 18 19 21 22 25 28
+ 29 31 35
c108 35 0 1.32669e-19 $X=8.445 $Y=1.02
c109 29 0 4.08738e-20 $X=8.81 $Y=1.415
c110 25 0 1.94589e-20 $X=8.445 $Y=0.81
r111 40 42 6.12014 $w=3.3e-07 $l=3.5e-08 $layer=POLY_cond $X=6.92 $Y=1.595
+ $X2=6.955 $Y2=1.595
r112 31 33 32.7294 $w=2.48e-07 $l=7.1e-07 $layer=LI1_cond $X=8.81 $Y=1.88
+ $X2=8.81 $Y2=2.59
r113 29 36 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=8.81 $Y=1.33
+ $X2=8.525 $Y2=1.33
r114 29 31 21.4354 $w=2.48e-07 $l=4.65e-07 $layer=LI1_cond $X=8.81 $Y=1.415
+ $X2=8.81 $Y2=1.88
r115 28 36 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.525 $Y=1.245
+ $X2=8.525 $Y2=1.33
r116 27 35 3.70735 $w=2.5e-07 $l=1.18427e-07 $layer=LI1_cond $X=8.525 $Y=1.105
+ $X2=8.445 $Y2=1.02
r117 27 28 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=8.525 $Y=1.105
+ $X2=8.525 $Y2=1.245
r118 23 35 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=8.445 $Y=0.935
+ $X2=8.445 $Y2=1.02
r119 23 25 4.36531 $w=3.28e-07 $l=1.25e-07 $layer=LI1_cond $X=8.445 $Y=0.935
+ $X2=8.445 $Y2=0.81
r120 21 35 2.76166 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.28 $Y=1.02
+ $X2=8.445 $Y2=1.02
r121 21 22 68.1765 $w=1.68e-07 $l=1.045e-06 $layer=LI1_cond $X=8.28 $Y=1.02
+ $X2=7.235 $Y2=1.02
r122 19 42 29.7264 $w=3.3e-07 $l=1.7e-07 $layer=POLY_cond $X=7.125 $Y=1.595
+ $X2=6.955 $Y2=1.595
r123 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.125
+ $Y=1.595 $X2=7.125 $Y2=1.595
r124 16 22 6.96323 $w=1.7e-07 $l=1.46458e-07 $layer=LI1_cond $X=7.125 $Y=1.105
+ $X2=7.235 $Y2=1.02
r125 16 18 25.668 $w=2.18e-07 $l=4.9e-07 $layer=LI1_cond $X=7.125 $Y=1.105
+ $X2=7.125 $Y2=1.595
r126 13 15 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=6.955 $Y=2.24
+ $X2=6.955 $Y2=2.525
r127 12 13 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=6.955 $Y=2.15
+ $X2=6.955 $Y2=2.24
r128 11 42 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=6.955 $Y=1.76
+ $X2=6.955 $Y2=1.595
r129 11 12 151.597 $w=1.8e-07 $l=3.9e-07 $layer=POLY_cond $X=6.955 $Y=1.76
+ $X2=6.955 $Y2=2.15
r130 7 40 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.92 $Y=1.43
+ $X2=6.92 $Y2=1.595
r131 7 9 376.883 $w=1.5e-07 $l=7.35e-07 $layer=POLY_cond $X=6.92 $Y=1.43
+ $X2=6.92 $Y2=0.695
r132 2 33 400 $w=1.7e-07 $l=9.26971e-07 $layer=licon1_PDIFF $count=1 $X=8.62
+ $Y=1.735 $X2=8.77 $Y2=2.59
r133 2 31 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=8.62
+ $Y=1.735 $X2=8.77 $Y2=1.88
r134 1 25 182 $w=1.7e-07 $l=5.05173e-07 $layer=licon1_NDIFF $count=1 $X=8.305
+ $Y=0.37 $X2=8.445 $Y2=0.81
.ends

.subckt PM_SKY130_FD_SC_HS__SDFRBP_1%A_1221_97# 1 2 3 12 14 16 17 21 26 27 30 31
+ 33 36 41
c115 33 0 2.05564e-20 $X=8.105 $Y=1.41
c116 30 0 1.29256e-19 $X=7.49 $Y=2.32
c117 21 0 1.35224e-19 $X=6.675 $Y=2.585
r118 41 42 56.0258 $w=2.71e-07 $l=3.15e-07 $layer=POLY_cond $X=8.23 $Y=1.452
+ $X2=8.545 $Y2=1.452
r119 34 41 22.2325 $w=2.71e-07 $l=1.25e-07 $layer=POLY_cond $X=8.105 $Y=1.452
+ $X2=8.23 $Y2=1.452
r120 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.105
+ $Y=1.41 $X2=8.105 $Y2=1.41
r121 31 33 22.622 $w=2.68e-07 $l=5.3e-07 $layer=LI1_cond $X=7.575 $Y=1.41
+ $X2=8.105 $Y2=1.41
r122 30 39 10.6888 $w=3.31e-07 $l=3.83445e-07 $layer=LI1_cond $X=7.49 $Y=2.32
+ $X2=7.78 $Y2=2.537
r123 29 31 7.28469 $w=2.7e-07 $l=1.72337e-07 $layer=LI1_cond $X=7.49 $Y=1.545
+ $X2=7.575 $Y2=1.41
r124 29 30 50.5615 $w=1.68e-07 $l=7.75e-07 $layer=LI1_cond $X=7.49 $Y=1.545
+ $X2=7.49 $Y2=2.32
r125 28 36 3.64284 $w=2.55e-07 $l=1.69245e-07 $layer=LI1_cond $X=6.845 $Y=2.405
+ $X2=6.76 $Y2=2.537
r126 27 30 6.01027 $w=3.31e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.405 $Y=2.405
+ $X2=7.49 $Y2=2.32
r127 27 28 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=7.405 $Y=2.405
+ $X2=6.845 $Y2=2.405
r128 26 36 2.83584 $w=1.7e-07 $l=2.17e-07 $layer=LI1_cond $X=6.76 $Y=2.32
+ $X2=6.76 $Y2=2.537
r129 25 26 91.0107 $w=1.68e-07 $l=1.395e-06 $layer=LI1_cond $X=6.76 $Y=0.925
+ $X2=6.76 $Y2=2.32
r130 21 36 3.64284 $w=2.55e-07 $l=1.06325e-07 $layer=LI1_cond $X=6.675 $Y=2.585
+ $X2=6.76 $Y2=2.537
r131 21 23 11.355 $w=3.38e-07 $l=3.35e-07 $layer=LI1_cond $X=6.675 $Y=2.585
+ $X2=6.34 $Y2=2.585
r132 17 25 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=6.675 $Y=0.76
+ $X2=6.76 $Y2=0.925
r133 17 19 12.5721 $w=3.28e-07 $l=3.6e-07 $layer=LI1_cond $X=6.675 $Y=0.76
+ $X2=6.315 $Y2=0.76
r134 14 42 16.5906 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=8.545 $Y=1.66
+ $X2=8.545 $Y2=1.452
r135 14 16 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=8.545 $Y=1.66
+ $X2=8.545 $Y2=2.235
r136 10 41 16.5906 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=8.23 $Y=1.245
+ $X2=8.23 $Y2=1.452
r137 10 12 284.585 $w=1.5e-07 $l=5.55e-07 $layer=POLY_cond $X=8.23 $Y=1.245
+ $X2=8.23 $Y2=0.69
r138 3 39 600 $w=1.7e-07 $l=2.85307e-07 $layer=licon1_PDIFF $count=1 $X=7.63
+ $Y=2.315 $X2=7.78 $Y2=2.535
r139 2 23 600 $w=1.7e-07 $l=3.36749e-07 $layer=licon1_PDIFF $count=1 $X=6.19
+ $Y=2.315 $X2=6.34 $Y2=2.585
r140 1 19 182 $w=1.7e-07 $l=3.65205e-07 $layer=licon1_NDIFF $count=1 $X=6.105
+ $Y=0.485 $X2=6.315 $Y2=0.76
.ends

.subckt PM_SKY130_FD_SC_HS__SDFRBP_1%A_850_74# 1 2 7 9 10 12 13 16 17 19 20 23
+ 25 26 27 29 30 32 33 37 38 39 42 44 45 46 48 50 52 55 57 60 68
c192 68 0 1.36582e-19 $X=5.13 $Y=1.465
c193 42 0 1.87517e-19 $X=9.755 $Y=0.58
c194 39 0 6.14302e-20 $X=9.07 $Y=1.585
c195 38 0 2.17443e-21 $X=9.68 $Y=1.585
c196 17 0 1.69935e-19 $X=5.955 $Y=1.26
c197 16 0 1.35224e-19 $X=5.605 $Y=3.075
c198 7 0 2.4889e-19 $X=5.04 $Y=1.185
r199 69 71 33.0468 $w=2.99e-07 $l=2.05e-07 $layer=POLY_cond $X=5.13 $Y=1.465
+ $X2=5.13 $Y2=1.26
r200 68 69 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.13
+ $Y=1.465 $X2=5.13 $Y2=1.465
r201 65 68 8.03218 $w=3.28e-07 $l=2.3e-07 $layer=LI1_cond $X=4.9 $Y=1.465
+ $X2=5.13 $Y2=1.465
r202 60 63 4.84026 $w=2.48e-07 $l=1.05e-07 $layer=LI1_cond $X=4.46 $Y=1.885
+ $X2=4.46 $Y2=1.99
r203 56 65 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.9 $Y=1.63 $X2=4.9
+ $Y2=1.465
r204 56 57 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=4.9 $Y=1.63 $X2=4.9
+ $Y2=1.8
r205 55 65 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.9 $Y=1.3 $X2=4.9
+ $Y2=1.465
r206 54 55 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=4.9 $Y=1.01 $X2=4.9
+ $Y2=1.3
r207 53 60 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.585 $Y=1.885
+ $X2=4.46 $Y2=1.885
r208 52 57 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.815 $Y=1.885
+ $X2=4.9 $Y2=1.8
r209 52 53 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=4.815 $Y=1.885
+ $X2=4.585 $Y2=1.885
r210 51 59 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.48 $Y=0.925
+ $X2=4.355 $Y2=0.925
r211 50 54 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.815 $Y=0.925
+ $X2=4.9 $Y2=1.01
r212 50 51 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=4.815 $Y=0.925
+ $X2=4.48 $Y2=0.925
r213 46 59 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.355 $Y=0.84
+ $X2=4.355 $Y2=0.925
r214 46 48 14.9818 $w=2.48e-07 $l=3.25e-07 $layer=LI1_cond $X=4.355 $Y=0.84
+ $X2=4.355 $Y2=0.515
r215 40 42 476.872 $w=1.5e-07 $l=9.3e-07 $layer=POLY_cond $X=9.755 $Y=1.51
+ $X2=9.755 $Y2=0.58
r216 38 40 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=9.68 $Y=1.585
+ $X2=9.755 $Y2=1.51
r217 38 39 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=9.68 $Y=1.585
+ $X2=9.07 $Y2=1.585
r218 35 37 294.84 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=8.995 $Y=2.81
+ $X2=8.995 $Y2=2.235
r219 34 39 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=8.995 $Y=1.66
+ $X2=9.07 $Y2=1.585
r220 34 37 294.84 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=8.995 $Y=1.66
+ $X2=8.995 $Y2=2.235
r221 32 35 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=8.995 $Y=2.9
+ $X2=8.995 $Y2=2.81
r222 32 33 68.0242 $w=1.8e-07 $l=1.75e-07 $layer=POLY_cond $X=8.995 $Y=2.9
+ $X2=8.995 $Y2=3.075
r223 31 45 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=6.655 $Y=3.15
+ $X2=6.565 $Y2=3.15
r224 30 33 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=8.905 $Y=3.15
+ $X2=8.995 $Y2=3.075
r225 30 31 1153.72 $w=1.5e-07 $l=2.25e-06 $layer=POLY_cond $X=8.905 $Y=3.15
+ $X2=6.655 $Y2=3.15
r226 27 29 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=6.565 $Y=2.81
+ $X2=6.565 $Y2=2.525
r227 26 45 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=6.565 $Y=3.075
+ $X2=6.565 $Y2=3.15
r228 25 27 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=6.565 $Y=2.9
+ $X2=6.565 $Y2=2.81
r229 25 26 68.0242 $w=1.8e-07 $l=1.75e-07 $layer=POLY_cond $X=6.565 $Y=2.9
+ $X2=6.565 $Y2=3.075
r230 21 23 251.255 $w=1.5e-07 $l=4.9e-07 $layer=POLY_cond $X=6.03 $Y=1.185
+ $X2=6.03 $Y2=0.695
r231 19 45 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=6.475 $Y=3.15
+ $X2=6.565 $Y2=3.15
r232 19 20 407.649 $w=1.5e-07 $l=7.95e-07 $layer=POLY_cond $X=6.475 $Y=3.15
+ $X2=5.68 $Y2=3.15
r233 18 44 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.68 $Y=1.26
+ $X2=5.605 $Y2=1.26
r234 17 21 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.955 $Y=1.26
+ $X2=6.03 $Y2=1.185
r235 17 18 141.011 $w=1.5e-07 $l=2.75e-07 $layer=POLY_cond $X=5.955 $Y=1.26
+ $X2=5.68 $Y2=1.26
r236 16 20 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.605 $Y=3.075
+ $X2=5.68 $Y2=3.15
r237 15 44 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.605 $Y=1.335
+ $X2=5.605 $Y2=1.26
r238 15 16 892.213 $w=1.5e-07 $l=1.74e-06 $layer=POLY_cond $X=5.605 $Y=1.335
+ $X2=5.605 $Y2=3.075
r239 14 71 18.89 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.295 $Y=1.26
+ $X2=5.13 $Y2=1.26
r240 13 44 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.53 $Y=1.26
+ $X2=5.605 $Y2=1.26
r241 13 14 120.5 $w=1.5e-07 $l=2.35e-07 $layer=POLY_cond $X=5.53 $Y=1.26
+ $X2=5.295 $Y2=1.26
r242 10 69 57.0947 $w=2.99e-07 $l=2.96985e-07 $layer=POLY_cond $X=5.095 $Y=1.745
+ $X2=5.13 $Y2=1.465
r243 10 12 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=5.095 $Y=1.745
+ $X2=5.095 $Y2=2.38
r244 7 71 24.0479 $w=2.99e-07 $l=1.21861e-07 $layer=POLY_cond $X=5.04 $Y=1.185
+ $X2=5.13 $Y2=1.26
r245 7 9 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=5.04 $Y=1.185
+ $X2=5.04 $Y2=0.74
r246 2 63 600 $w=1.7e-07 $l=2.31409e-07 $layer=licon1_PDIFF $count=1 $X=4.275
+ $Y=1.82 $X2=4.42 $Y2=1.99
r247 1 59 182 $w=1.7e-07 $l=6.23298e-07 $layer=licon1_NDIFF $count=1 $X=4.25
+ $Y=0.37 $X2=4.395 $Y2=0.925
r248 1 48 182 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=1 $X=4.25
+ $Y=0.37 $X2=4.395 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__SDFRBP_1%A_2008_48# 1 2 9 11 12 13 15 18 21 22 25 28
+ 29 31 32 34 35 37
c136 29 0 1.60243e-20 $X=11.675 $Y=0.665
c137 21 0 2.44776e-20 $X=10.855 $Y=2.405
c138 18 0 6.47027e-20 $X=10.36 $Y=1.815
r139 37 39 4.01609 $w=3.28e-07 $l=1.15e-07 $layer=LI1_cond $X=11.12 $Y=0.55
+ $X2=11.12 $Y2=0.665
r140 33 34 57.4118 $w=1.68e-07 $l=8.8e-07 $layer=LI1_cond $X=11.76 $Y=0.75
+ $X2=11.76 $Y2=1.63
r141 31 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=11.675 $Y=1.715
+ $X2=11.76 $Y2=1.63
r142 31 32 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=11.675 $Y=1.715
+ $X2=11.405 $Y2=1.715
r143 30 39 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.285 $Y=0.665
+ $X2=11.12 $Y2=0.665
r144 29 33 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=11.675 $Y=0.665
+ $X2=11.76 $Y2=0.75
r145 29 30 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=11.675 $Y=0.665
+ $X2=11.285 $Y2=0.665
r146 28 35 3.70735 $w=2.5e-07 $l=2.28583e-07 $layer=LI1_cond $X=11.32 $Y=2.32
+ $X2=11.13 $Y2=2.405
r147 27 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=11.32 $Y=1.8
+ $X2=11.405 $Y2=1.715
r148 27 28 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=11.32 $Y=1.8
+ $X2=11.32 $Y2=2.32
r149 23 35 3.70735 $w=2.5e-07 $l=1.46458e-07 $layer=LI1_cond $X=11.02 $Y=2.49
+ $X2=11.13 $Y2=2.405
r150 23 25 5.76222 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=11.02 $Y=2.49
+ $X2=11.02 $Y2=2.655
r151 21 35 2.76166 $w=1.7e-07 $l=2.75e-07 $layer=LI1_cond $X=10.855 $Y=2.405
+ $X2=11.13 $Y2=2.405
r152 21 22 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=10.855 $Y=2.405
+ $X2=10.525 $Y2=2.405
r153 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.36
+ $Y=1.815 $X2=10.36 $Y2=1.815
r154 16 22 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=10.395 $Y=2.32
+ $X2=10.525 $Y2=2.405
r155 16 18 22.384 $w=2.58e-07 $l=5.05e-07 $layer=LI1_cond $X=10.395 $Y=2.32
+ $X2=10.395 $Y2=1.815
r156 13 15 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=10.16 $Y=2.37
+ $X2=10.16 $Y2=2.655
r157 12 13 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=10.16 $Y=2.28
+ $X2=10.16 $Y2=2.37
r158 11 19 34.2225 $w=3.69e-07 $l=2.17612e-07 $layer=POLY_cond $X=10.16 $Y=1.98
+ $X2=10.282 $Y2=1.815
r159 11 12 116.613 $w=1.8e-07 $l=3e-07 $layer=POLY_cond $X=10.16 $Y=1.98
+ $X2=10.16 $Y2=2.28
r160 7 19 58.6339 $w=3.69e-07 $l=3.89654e-07 $layer=POLY_cond $X=10.115 $Y=1.5
+ $X2=10.282 $Y2=1.815
r161 7 9 471.745 $w=1.5e-07 $l=9.2e-07 $layer=POLY_cond $X=10.115 $Y=1.5
+ $X2=10.115 $Y2=0.58
r162 2 25 600 $w=1.7e-07 $l=2.74955e-07 $layer=licon1_PDIFF $count=1 $X=10.87
+ $Y=2.445 $X2=11.02 $Y2=2.655
r163 1 37 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=10.98
+ $Y=0.37 $X2=11.12 $Y2=0.55
.ends

.subckt PM_SKY130_FD_SC_HS__SDFRBP_1%A_1747_74# 1 2 7 9 10 11 12 14 16 17 19 20
+ 22 23 24 26 27 29 32 40 42 45 47 51 52 56 58 59 61
c180 58 0 8.18376e-20 $X=10.01 $Y=2.425
c181 10 0 1.78926e-19 $X=11.26 $Y=1.02
c182 7 0 1.60243e-20 $X=10.905 $Y=0.87
r183 68 69 4.6235 $w=4.17e-07 $l=4e-08 $layer=POLY_cond $X=11.925 $Y=1.5
+ $X2=11.965 $Y2=1.5
r184 64 65 15.0154 $w=2.6e-07 $l=3.2e-07 $layer=LI1_cond $X=9.69 $Y=1.175
+ $X2=10.01 $Y2=1.175
r185 59 65 4.30428 $w=4.3e-07 $l=1.05119e-07 $layer=LI1_cond $X=10.095 $Y=1.22
+ $X2=10.01 $Y2=1.175
r186 59 61 31.2232 $w=4.28e-07 $l=1.165e-06 $layer=LI1_cond $X=10.095 $Y=1.22
+ $X2=11.26 $Y2=1.22
r187 57 65 3.22376 $w=1.7e-07 $l=2.6e-07 $layer=LI1_cond $X=10.01 $Y=1.435
+ $X2=10.01 $Y2=1.175
r188 57 58 64.5882 $w=1.68e-07 $l=9.9e-07 $layer=LI1_cond $X=10.01 $Y=1.435
+ $X2=10.01 $Y2=2.425
r189 56 64 3.22376 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=9.69 $Y=1.005
+ $X2=9.69 $Y2=1.175
r190 55 56 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=9.69 $Y=0.735
+ $X2=9.69 $Y2=1.005
r191 52 54 7.68295 $w=3.28e-07 $l=2.2e-07 $layer=LI1_cond $X=9.325 $Y=2.59
+ $X2=9.545 $Y2=2.59
r192 51 58 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=9.925 $Y=2.59
+ $X2=10.01 $Y2=2.425
r193 51 54 13.2706 $w=3.28e-07 $l=3.8e-07 $layer=LI1_cond $X=9.925 $Y=2.59
+ $X2=9.545 $Y2=2.59
r194 47 55 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=9.605 $Y=0.57
+ $X2=9.69 $Y2=0.735
r195 47 49 8.20679 $w=3.28e-07 $l=2.35e-07 $layer=LI1_cond $X=9.605 $Y=0.57
+ $X2=9.37 $Y2=0.57
r196 43 52 7.17723 $w=3.3e-07 $l=2.13014e-07 $layer=LI1_cond $X=9.215 $Y=2.425
+ $X2=9.325 $Y2=2.59
r197 43 45 26.4538 $w=2.18e-07 $l=5.05e-07 $layer=LI1_cond $X=9.215 $Y=2.425
+ $X2=9.215 $Y2=1.92
r198 38 40 53.8404 $w=1.5e-07 $l=1.05e-07 $layer=POLY_cond $X=11.245 $Y=2.295
+ $X2=11.35 $Y2=2.295
r199 30 42 34.7346 $w=1.65e-07 $l=1.72337e-07 $layer=POLY_cond $X=12.93 $Y=1.355
+ $X2=12.915 $Y2=1.52
r200 30 32 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=12.93 $Y=1.355
+ $X2=12.93 $Y2=0.645
r201 27 29 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=12.915 $Y=2.045
+ $X2=12.915 $Y2=2.54
r202 26 27 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=12.915 $Y=1.955
+ $X2=12.915 $Y2=2.045
r203 25 42 34.7346 $w=1.65e-07 $l=1.65e-07 $layer=POLY_cond $X=12.915 $Y=1.685
+ $X2=12.915 $Y2=1.52
r204 25 26 104.952 $w=1.8e-07 $l=2.7e-07 $layer=POLY_cond $X=12.915 $Y=1.685
+ $X2=12.915 $Y2=1.955
r205 24 69 10.9026 $w=4.17e-07 $l=8.44097e-08 $layer=POLY_cond $X=12.04 $Y=1.52
+ $X2=11.965 $Y2=1.5
r206 23 42 3.90195 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=12.825 $Y=1.52
+ $X2=12.915 $Y2=1.52
r207 23 24 137.266 $w=3.3e-07 $l=7.85e-07 $layer=POLY_cond $X=12.825 $Y=1.52
+ $X2=12.04 $Y2=1.52
r208 20 69 26.8826 $w=1.5e-07 $l=2.65e-07 $layer=POLY_cond $X=11.965 $Y=1.235
+ $X2=11.965 $Y2=1.5
r209 20 22 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=11.965 $Y=1.235
+ $X2=11.965 $Y2=0.74
r210 17 68 26.8826 $w=1.5e-07 $l=2.65e-07 $layer=POLY_cond $X=11.925 $Y=1.765
+ $X2=11.925 $Y2=1.5
r211 17 19 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=11.925 $Y=1.765
+ $X2=11.925 $Y2=2.4
r212 16 40 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=11.35 $Y=2.22
+ $X2=11.35 $Y2=2.295
r213 15 68 66.4628 $w=4.17e-07 $l=5.75e-07 $layer=POLY_cond $X=11.35 $Y=1.5
+ $X2=11.925 $Y2=1.5
r214 15 16 274.33 $w=1.5e-07 $l=5.35e-07 $layer=POLY_cond $X=11.35 $Y=1.685
+ $X2=11.35 $Y2=2.22
r215 12 38 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=11.245 $Y=2.37
+ $X2=11.245 $Y2=2.295
r216 12 14 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=11.245 $Y=2.37
+ $X2=11.245 $Y2=2.655
r217 11 15 10.4029 $w=4.17e-07 $l=3.06716e-07 $layer=POLY_cond $X=11.26 $Y=1.235
+ $X2=11.35 $Y2=1.5
r218 11 61 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=11.26
+ $Y=1.27 $X2=11.26 $Y2=1.27
r219 10 34 182.032 $w=1.5e-07 $l=3.55e-07 $layer=POLY_cond $X=11.26 $Y=0.945
+ $X2=10.905 $Y2=0.945
r220 10 11 37.5952 $w=3.3e-07 $l=2.15e-07 $layer=POLY_cond $X=11.26 $Y=1.02
+ $X2=11.26 $Y2=1.235
r221 7 34 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=10.905 $Y=0.87
+ $X2=10.905 $Y2=0.945
r222 7 9 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=10.905 $Y=0.87
+ $X2=10.905 $Y2=0.58
r223 2 54 600 $w=1.7e-07 $l=1.06637e-06 $layer=licon1_PDIFF $count=1 $X=9.07
+ $Y=1.735 $X2=9.545 $Y2=2.59
r224 2 45 300 $w=1.7e-07 $l=2.48948e-07 $layer=licon1_PDIFF $count=2 $X=9.07
+ $Y=1.735 $X2=9.22 $Y2=1.92
r225 1 49 182 $w=1.7e-07 $l=7.28166e-07 $layer=licon1_NDIFF $count=1 $X=8.735
+ $Y=0.37 $X2=9.37 $Y2=0.57
.ends

.subckt PM_SKY130_FD_SC_HS__SDFRBP_1%A_2513_424# 1 2 9 11 13 16 20 24 27
r50 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=13.38
+ $Y=1.465 $X2=13.38 $Y2=1.465
r51 22 27 0.820356 $w=3.3e-07 $l=1.43e-07 $layer=LI1_cond $X=12.855 $Y=1.465
+ $X2=12.712 $Y2=1.465
r52 22 24 18.3343 $w=3.28e-07 $l=5.25e-07 $layer=LI1_cond $X=12.855 $Y=1.465
+ $X2=13.38 $Y2=1.465
r53 18 27 5.82594 $w=2.85e-07 $l=1.65e-07 $layer=LI1_cond $X=12.712 $Y=1.63
+ $X2=12.712 $Y2=1.465
r54 18 20 25.6772 $w=2.83e-07 $l=6.35e-07 $layer=LI1_cond $X=12.712 $Y=1.63
+ $X2=12.712 $Y2=2.265
r55 14 27 5.82594 $w=2.85e-07 $l=1.65e-07 $layer=LI1_cond $X=12.712 $Y=1.3
+ $X2=12.712 $Y2=1.465
r56 14 16 26.486 $w=2.83e-07 $l=6.55e-07 $layer=LI1_cond $X=12.712 $Y=1.3
+ $X2=12.712 $Y2=0.645
r57 11 25 61.4066 $w=2.86e-07 $l=3.26343e-07 $layer=POLY_cond $X=13.435 $Y=1.765
+ $X2=13.38 $Y2=1.465
r58 11 13 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=13.435 $Y=1.765
+ $X2=13.435 $Y2=2.4
r59 7 25 38.6549 $w=2.86e-07 $l=1.83916e-07 $layer=POLY_cond $X=13.42 $Y=1.3
+ $X2=13.38 $Y2=1.465
r60 7 9 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=13.42 $Y=1.3 $X2=13.42
+ $Y2=0.74
r61 2 20 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=12.565
+ $Y=2.12 $X2=12.69 $Y2=2.265
r62 1 16 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=12.59
+ $Y=0.37 $X2=12.715 $Y2=0.645
.ends

.subckt PM_SKY130_FD_SC_HS__SDFRBP_1%VPWR 1 2 3 4 5 6 7 8 27 31 35 39 43 49 52
+ 55 59 64 65 67 68 70 71 73 75 84 101 105 110 115 122 123 126 129 132 135 138
c182 4 0 1.29256e-19 $X=7.03 $Y=2.315
c183 2 0 5.02674e-20 $X=3.1 $Y=2.32
r184 138 139 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.2 $Y=3.33
+ $X2=13.2 $Y2=3.33
r185 135 136 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=11.76 $Y=3.33
+ $X2=11.76 $Y2=3.33
r186 132 133 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.32 $Y=3.33
+ $X2=10.32 $Y2=3.33
r187 129 130 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=3.33
+ $X2=8.4 $Y2=3.33
r188 126 127 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r189 123 139 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=13.68 $Y=3.33
+ $X2=13.2 $Y2=3.33
r190 122 123 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.68 $Y=3.33
+ $X2=13.68 $Y2=3.33
r191 120 138 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=13.325 $Y=3.33
+ $X2=13.185 $Y2=3.33
r192 120 122 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=13.325 $Y=3.33
+ $X2=13.68 $Y2=3.33
r193 119 139 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.72 $Y=3.33
+ $X2=13.2 $Y2=3.33
r194 119 136 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=12.72 $Y=3.33
+ $X2=11.76 $Y2=3.33
r195 118 119 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=12.72 $Y=3.33
+ $X2=12.72 $Y2=3.33
r196 116 135 10.508 $w=1.7e-07 $l=2.23e-07 $layer=LI1_cond $X=11.815 $Y=3.33
+ $X2=11.592 $Y2=3.33
r197 116 118 59.0428 $w=1.68e-07 $l=9.05e-07 $layer=LI1_cond $X=11.815 $Y=3.33
+ $X2=12.72 $Y2=3.33
r198 115 138 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=13.045 $Y=3.33
+ $X2=13.185 $Y2=3.33
r199 115 118 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=13.045 $Y=3.33
+ $X2=12.72 $Y2=3.33
r200 114 136 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.28 $Y=3.33
+ $X2=11.76 $Y2=3.33
r201 114 133 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=11.28 $Y=3.33
+ $X2=10.32 $Y2=3.33
r202 113 114 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=11.28 $Y=3.33
+ $X2=11.28 $Y2=3.33
r203 111 132 8.88104 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=10.65 $Y=3.33
+ $X2=10.477 $Y2=3.33
r204 111 113 41.1016 $w=1.68e-07 $l=6.3e-07 $layer=LI1_cond $X=10.65 $Y=3.33
+ $X2=11.28 $Y2=3.33
r205 110 135 10.508 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=11.37 $Y=3.33
+ $X2=11.592 $Y2=3.33
r206 110 113 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=11.37 $Y=3.33
+ $X2=11.28 $Y2=3.33
r207 109 133 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=8.88 $Y=3.33
+ $X2=10.32 $Y2=3.33
r208 109 130 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=3.33
+ $X2=8.4 $Y2=3.33
r209 108 109 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r210 106 129 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.485 $Y=3.33
+ $X2=8.36 $Y2=3.33
r211 106 108 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=8.485 $Y=3.33
+ $X2=8.88 $Y2=3.33
r212 105 132 8.88104 $w=1.7e-07 $l=1.72e-07 $layer=LI1_cond $X=10.305 $Y=3.33
+ $X2=10.477 $Y2=3.33
r213 105 108 92.9679 $w=1.68e-07 $l=1.425e-06 $layer=LI1_cond $X=10.305 $Y=3.33
+ $X2=8.88 $Y2=3.33
r214 104 130 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=3.33
+ $X2=8.4 $Y2=3.33
r215 103 104 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r216 101 129 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.235 $Y=3.33
+ $X2=8.36 $Y2=3.33
r217 101 103 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=8.235 $Y=3.33
+ $X2=7.92 $Y2=3.33
r218 96 99 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=5.04 $Y=3.33
+ $X2=6.96 $Y2=3.33
r219 96 97 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r220 94 97 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=5.04 $Y2=3.33
r221 93 94 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r222 91 94 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.56 $Y2=3.33
r223 91 127 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=3.12 $Y2=3.33
r224 90 93 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=3.6 $Y=3.33 $X2=4.56
+ $Y2=3.33
r225 90 91 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r226 88 126 9.14399 $w=1.7e-07 $l=1.8e-07 $layer=LI1_cond $X=3.445 $Y=3.33
+ $X2=3.265 $Y2=3.33
r227 88 90 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=3.445 $Y=3.33
+ $X2=3.6 $Y2=3.33
r228 87 127 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=3.12 $Y2=3.33
r229 86 87 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r230 84 126 9.14399 $w=1.7e-07 $l=1.8e-07 $layer=LI1_cond $X=3.085 $Y=3.33
+ $X2=3.265 $Y2=3.33
r231 84 86 91.6631 $w=1.68e-07 $l=1.405e-06 $layer=LI1_cond $X=3.085 $Y=3.33
+ $X2=1.68 $Y2=3.33
r232 83 87 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=1.68 $Y2=3.33
r233 82 83 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r234 79 83 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=1.2 $Y2=3.33
r235 78 82 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.24 $Y=3.33 $X2=1.2
+ $Y2=3.33
r236 78 79 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r237 75 104 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=7.92 $Y2=3.33
r238 75 97 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=5.04 $Y2=3.33
r239 75 99 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r240 73 74 5.78802 $w=4.43e-07 $l=1.2e-07 $layer=LI1_cond $X=11.592 $Y=2.815
+ $X2=11.592 $Y2=2.695
r241 70 99 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=7.09 $Y=3.33
+ $X2=6.96 $Y2=3.33
r242 70 71 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.09 $Y=3.33
+ $X2=7.255 $Y2=3.33
r243 69 103 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=7.42 $Y=3.33
+ $X2=7.92 $Y2=3.33
r244 69 71 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.42 $Y=3.33
+ $X2=7.255 $Y2=3.33
r245 67 93 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=4.705 $Y=3.33
+ $X2=4.56 $Y2=3.33
r246 67 68 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.705 $Y=3.33
+ $X2=4.87 $Y2=3.33
r247 66 96 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=5.035 $Y=3.33
+ $X2=5.04 $Y2=3.33
r248 66 68 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.035 $Y=3.33
+ $X2=4.87 $Y2=3.33
r249 64 82 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=1.225 $Y=3.33
+ $X2=1.2 $Y2=3.33
r250 64 65 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.225 $Y=3.33
+ $X2=1.39 $Y2=3.33
r251 63 86 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=1.555 $Y=3.33
+ $X2=1.68 $Y2=3.33
r252 63 65 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.555 $Y=3.33
+ $X2=1.39 $Y2=3.33
r253 59 62 17.0809 $w=2.78e-07 $l=4.15e-07 $layer=LI1_cond $X=13.185 $Y=1.985
+ $X2=13.185 $Y2=2.4
r254 57 138 0.375625 $w=2.8e-07 $l=8.5e-08 $layer=LI1_cond $X=13.185 $Y=3.245
+ $X2=13.185 $Y2=3.33
r255 57 62 34.7791 $w=2.78e-07 $l=8.45e-07 $layer=LI1_cond $X=13.185 $Y=3.245
+ $X2=13.185 $Y2=2.4
r256 55 74 28.0595 $w=2.28e-07 $l=5.6e-07 $layer=LI1_cond $X=11.7 $Y=2.135
+ $X2=11.7 $Y2=2.695
r257 52 135 1.76584 $w=4.45e-07 $l=8.5e-08 $layer=LI1_cond $X=11.592 $Y=3.245
+ $X2=11.592 $Y2=3.33
r258 51 73 2.64155 $w=4.43e-07 $l=1.02e-07 $layer=LI1_cond $X=11.592 $Y=2.917
+ $X2=11.592 $Y2=2.815
r259 51 52 8.49441 $w=4.43e-07 $l=3.28e-07 $layer=LI1_cond $X=11.592 $Y=2.917
+ $X2=11.592 $Y2=3.245
r260 47 132 1.03204 $w=3.45e-07 $l=8.5e-08 $layer=LI1_cond $X=10.477 $Y=3.245
+ $X2=10.477 $Y2=3.33
r261 47 49 14.0297 $w=3.43e-07 $l=4.2e-07 $layer=LI1_cond $X=10.477 $Y=3.245
+ $X2=10.477 $Y2=2.825
r262 43 46 32.7294 $w=2.48e-07 $l=7.1e-07 $layer=LI1_cond $X=8.36 $Y=1.88
+ $X2=8.36 $Y2=2.59
r263 41 129 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=8.36 $Y=3.245
+ $X2=8.36 $Y2=3.33
r264 41 46 30.194 $w=2.48e-07 $l=6.55e-07 $layer=LI1_cond $X=8.36 $Y=3.245
+ $X2=8.36 $Y2=2.59
r265 37 71 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.255 $Y=3.245
+ $X2=7.255 $Y2=3.33
r266 37 39 14.6675 $w=3.28e-07 $l=4.2e-07 $layer=LI1_cond $X=7.255 $Y=3.245
+ $X2=7.255 $Y2=2.825
r267 33 68 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.87 $Y=3.245
+ $X2=4.87 $Y2=3.33
r268 33 35 16.0644 $w=3.28e-07 $l=4.6e-07 $layer=LI1_cond $X=4.87 $Y=3.245
+ $X2=4.87 $Y2=2.785
r269 29 126 1.16013 $w=3.6e-07 $l=8.5e-08 $layer=LI1_cond $X=3.265 $Y=3.245
+ $X2=3.265 $Y2=3.33
r270 29 31 13.7653 $w=3.58e-07 $l=4.3e-07 $layer=LI1_cond $X=3.265 $Y=3.245
+ $X2=3.265 $Y2=2.815
r271 25 65 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.39 $Y=3.245
+ $X2=1.39 $Y2=3.33
r272 25 27 26.8903 $w=3.28e-07 $l=7.7e-07 $layer=LI1_cond $X=1.39 $Y=3.245
+ $X2=1.39 $Y2=2.475
r273 8 62 300 $w=1.7e-07 $l=3.60832e-07 $layer=licon1_PDIFF $count=2 $X=12.99
+ $Y=2.12 $X2=13.175 $Y2=2.4
r274 8 59 600 $w=1.7e-07 $l=2.79464e-07 $layer=licon1_PDIFF $count=1 $X=12.99
+ $Y=2.12 $X2=13.21 $Y2=1.985
r275 7 73 600 $w=1.7e-07 $l=4.65242e-07 $layer=licon1_PDIFF $count=1 $X=11.32
+ $Y=2.445 $X2=11.535 $Y2=2.815
r276 7 55 300 $w=1.7e-07 $l=5.06828e-07 $layer=licon1_PDIFF $count=2 $X=11.32
+ $Y=2.445 $X2=11.695 $Y2=2.135
r277 6 49 600 $w=1.7e-07 $l=4.85386e-07 $layer=licon1_PDIFF $count=1 $X=10.235
+ $Y=2.445 $X2=10.475 $Y2=2.825
r278 5 46 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=8.185
+ $Y=1.735 $X2=8.32 $Y2=2.59
r279 5 43 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=8.185
+ $Y=1.735 $X2=8.32 $Y2=1.88
r280 4 39 600 $w=1.7e-07 $l=6.1225e-07 $layer=licon1_PDIFF $count=1 $X=7.03
+ $Y=2.315 $X2=7.255 $Y2=2.825
r281 3 35 600 $w=1.7e-07 $l=1.03729e-06 $layer=licon1_PDIFF $count=1 $X=4.72
+ $Y=1.82 $X2=4.87 $Y2=2.785
r282 2 31 600 $w=1.7e-07 $l=5.71577e-07 $layer=licon1_PDIFF $count=1 $X=3.1
+ $Y=2.32 $X2=3.265 $Y2=2.815
r283 1 27 300 $w=1.7e-07 $l=2.66458e-07 $layer=licon1_PDIFF $count=2 $X=1.19
+ $Y=2.32 $X2=1.39 $Y2=2.475
.ends

.subckt PM_SKY130_FD_SC_HS__SDFRBP_1%A_413_90# 1 2 3 4 5 20 23 24 26 29 30 32 33
+ 35 37 39 44 47 51 54
c146 51 0 1.69935e-19 $X=5.895 $Y=0.692
c147 33 0 1.41376e-19 $X=5.98 $Y=1.18
c148 23 0 5.02674e-20 $X=3.53 $Y=2.32
r149 54 56 4.92377 $w=2.23e-07 $l=9e-08 $layer=LI1_cond $X=5.85 $Y=2.435
+ $X2=5.85 $Y2=2.525
r150 53 54 15.0448 $w=2.23e-07 $l=2.75e-07 $layer=LI1_cond $X=5.85 $Y=2.16
+ $X2=5.85 $Y2=2.435
r151 49 51 4.55012 $w=1.93e-07 $l=8e-08 $layer=LI1_cond $X=5.815 $Y=0.692
+ $X2=5.895 $Y2=0.692
r152 43 44 5.07737 $w=2.38e-07 $l=8.5e-08 $layer=LI1_cond $X=3.53 $Y=2.44
+ $X2=3.445 $Y2=2.44
r153 39 41 8.55602 $w=3.28e-07 $l=2.45e-07 $layer=LI1_cond $X=2.435 $Y=0.76
+ $X2=2.435 $Y2=1.005
r154 34 35 52.8449 $w=1.68e-07 $l=8.1e-07 $layer=LI1_cond $X=6.42 $Y=1.265
+ $X2=6.42 $Y2=2.075
r155 32 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.335 $Y=1.18
+ $X2=6.42 $Y2=1.265
r156 32 33 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=6.335 $Y=1.18
+ $X2=5.98 $Y2=1.18
r157 31 53 2.32876 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.975 $Y=2.16
+ $X2=5.85 $Y2=2.16
r158 30 35 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.335 $Y=2.16
+ $X2=6.42 $Y2=2.075
r159 30 31 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=6.335 $Y=2.16
+ $X2=5.975 $Y2=2.16
r160 29 33 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.895 $Y=1.095
+ $X2=5.98 $Y2=1.18
r161 28 51 1.54022 $w=1.7e-07 $l=9.8e-08 $layer=LI1_cond $X=5.895 $Y=0.79
+ $X2=5.895 $Y2=0.692
r162 28 29 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=5.895 $Y=0.79
+ $X2=5.895 $Y2=1.095
r163 26 54 2.32876 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.725 $Y=2.435
+ $X2=5.85 $Y2=2.435
r164 26 47 113.519 $w=1.68e-07 $l=1.74e-06 $layer=LI1_cond $X=5.725 $Y=2.435
+ $X2=3.985 $Y2=2.435
r165 24 47 9.87921 $w=2.38e-07 $l=1.85e-07 $layer=LI1_cond $X=3.8 $Y=2.44
+ $X2=3.985 $Y2=2.44
r166 24 43 12.965 $w=2.38e-07 $l=2.7e-07 $layer=LI1_cond $X=3.8 $Y=2.44 $X2=3.53
+ $Y2=2.44
r167 23 43 2.75731 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=3.53 $Y=2.32
+ $X2=3.53 $Y2=2.44
r168 22 23 80.246 $w=1.68e-07 $l=1.23e-06 $layer=LI1_cond $X=3.53 $Y=1.09
+ $X2=3.53 $Y2=2.32
r169 21 41 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.6 $Y=1.005
+ $X2=2.435 $Y2=1.005
r170 20 22 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.445 $Y=1.005
+ $X2=3.53 $Y2=1.09
r171 20 21 55.1283 $w=1.68e-07 $l=8.45e-07 $layer=LI1_cond $X=3.445 $Y=1.005
+ $X2=2.6 $Y2=1.005
r172 19 37 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.425 $Y=2.475
+ $X2=2.26 $Y2=2.475
r173 19 44 66.5455 $w=1.68e-07 $l=1.02e-06 $layer=LI1_cond $X=2.425 $Y=2.475
+ $X2=3.445 $Y2=2.475
r174 5 56 600 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_PDIFF $count=1 $X=5.755
+ $Y=2.315 $X2=5.89 $Y2=2.525
r175 4 24 300 $w=1.7e-07 $l=2.17428e-07 $layer=licon1_PDIFF $count=2 $X=3.67
+ $Y=2.32 $X2=3.82 $Y2=2.475
r176 3 37 300 $w=1.7e-07 $l=2.17428e-07 $layer=licon1_PDIFF $count=2 $X=2.11
+ $Y=2.32 $X2=2.26 $Y2=2.475
r177 2 49 182 $w=1.7e-07 $l=2.67862e-07 $layer=licon1_NDIFF $count=1 $X=5.67
+ $Y=0.485 $X2=5.815 $Y2=0.69
r178 1 39 182 $w=1.7e-07 $l=5.01597e-07 $layer=licon1_NDIFF $count=1 $X=2.065
+ $Y=0.45 $X2=2.435 $Y2=0.76
.ends

.subckt PM_SKY130_FD_SC_HS__SDFRBP_1%Q_N 1 2 7 8 9 10 11 12 13
r21 13 40 1.3969 $w=3.28e-07 $l=4e-08 $layer=LI1_cond $X=12.18 $Y=2.775
+ $X2=12.18 $Y2=2.815
r22 12 13 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=12.18 $Y=2.405
+ $X2=12.18 $Y2=2.775
r23 12 34 12.2229 $w=3.28e-07 $l=3.5e-07 $layer=LI1_cond $X=12.18 $Y=2.405
+ $X2=12.18 $Y2=2.055
r24 11 34 0.69845 $w=3.28e-07 $l=2e-08 $layer=LI1_cond $X=12.18 $Y=2.035
+ $X2=12.18 $Y2=2.055
r25 10 11 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=12.18 $Y=1.665
+ $X2=12.18 $Y2=2.035
r26 9 10 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=12.18 $Y=1.295
+ $X2=12.18 $Y2=1.665
r27 8 9 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=12.18 $Y=0.925
+ $X2=12.18 $Y2=1.295
r28 7 8 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=12.18 $Y=0.515
+ $X2=12.18 $Y2=0.925
r29 2 40 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=12
+ $Y=1.84 $X2=12.15 $Y2=2.815
r30 2 34 400 $w=1.7e-07 $l=2.80134e-07 $layer=licon1_PDIFF $count=1 $X=12
+ $Y=1.84 $X2=12.15 $Y2=2.055
r31 1 7 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=12.04
+ $Y=0.37 $X2=12.18 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__SDFRBP_1%Q 1 2 9 10 11 12 13 28 32 43
r20 41 43 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=13.75 $Y=1.13
+ $X2=13.75 $Y2=1.82
r21 29 32 1.02897 $w=2.78e-07 $l=2.5e-08 $layer=LI1_cond $X=13.695 $Y=1.96
+ $X2=13.695 $Y2=1.985
r22 21 28 0.726197 $w=3.63e-07 $l=2.3e-08 $layer=LI1_cond $X=13.652 $Y=0.948
+ $X2=13.652 $Y2=0.925
r23 12 13 15.2287 $w=2.78e-07 $l=3.7e-07 $layer=LI1_cond $X=13.695 $Y=2.405
+ $X2=13.695 $Y2=2.775
r24 11 29 0.205793 $w=2.78e-07 $l=5e-09 $layer=LI1_cond $X=13.695 $Y=1.955
+ $X2=13.695 $Y2=1.96
r25 11 43 7.32213 $w=2.78e-07 $l=1.35e-07 $layer=LI1_cond $X=13.695 $Y=1.955
+ $X2=13.695 $Y2=1.82
r26 11 12 15.0229 $w=2.78e-07 $l=3.65e-07 $layer=LI1_cond $X=13.695 $Y=2.04
+ $X2=13.695 $Y2=2.405
r27 11 32 2.26373 $w=2.78e-07 $l=5.5e-08 $layer=LI1_cond $X=13.695 $Y=2.04
+ $X2=13.695 $Y2=1.985
r28 10 41 8.08227 $w=3.63e-07 $l=1.51e-07 $layer=LI1_cond $X=13.652 $Y=0.979
+ $X2=13.652 $Y2=1.13
r29 10 21 0.978787 $w=3.63e-07 $l=3.1e-08 $layer=LI1_cond $X=13.652 $Y=0.979
+ $X2=13.652 $Y2=0.948
r30 10 28 0.978787 $w=3.63e-07 $l=3.1e-08 $layer=LI1_cond $X=13.652 $Y=0.894
+ $X2=13.652 $Y2=0.925
r31 9 10 11.9665 $w=3.63e-07 $l=3.79e-07 $layer=LI1_cond $X=13.652 $Y=0.515
+ $X2=13.652 $Y2=0.894
r32 2 13 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=13.51
+ $Y=1.84 $X2=13.66 $Y2=2.815
r33 2 32 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=13.51
+ $Y=1.84 $X2=13.66 $Y2=1.985
r34 1 9 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=13.495
+ $Y=0.37 $X2=13.635 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__SDFRBP_1%VGND 1 2 3 4 5 6 7 24 28 32 36 40 42 46 49
+ 50 52 53 54 56 71 75 83 90 91 94 97 100 104 110
c139 91 0 2.51459e-20 $X=13.68 $Y=0
c140 32 0 1.36582e-19 $X=4.825 $Y=0.55
c141 28 0 1.5551e-19 $X=3.835 $Y=0.585
r142 110 111 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=13.2 $Y=0
+ $X2=13.2 $Y2=0
r143 105 111 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=11.76 $Y=0
+ $X2=13.2 $Y2=0
r144 104 107 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=11.675 $Y=0
+ $X2=11.675 $Y2=0.325
r145 104 105 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=11.76 $Y=0
+ $X2=11.76 $Y2=0
r146 100 101 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.32 $Y=0
+ $X2=10.32 $Y2=0
r147 97 98 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=7.44 $Y=0 $X2=7.44
+ $Y2=0
r148 94 95 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r149 91 111 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=13.68 $Y=0
+ $X2=13.2 $Y2=0
r150 90 91 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.68 $Y=0
+ $X2=13.68 $Y2=0
r151 88 110 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=13.29 $Y=0
+ $X2=13.205 $Y2=0
r152 88 90 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=13.29 $Y=0
+ $X2=13.68 $Y2=0
r153 87 105 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.28 $Y=0
+ $X2=11.76 $Y2=0
r154 87 101 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=11.28 $Y=0
+ $X2=10.32 $Y2=0
r155 86 87 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=11.28 $Y=0
+ $X2=11.28 $Y2=0
r156 84 100 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.495 $Y=0
+ $X2=10.33 $Y2=0
r157 84 86 51.2139 $w=1.68e-07 $l=7.85e-07 $layer=LI1_cond $X=10.495 $Y=0
+ $X2=11.28 $Y2=0
r158 83 104 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.51 $Y=0
+ $X2=11.675 $Y2=0
r159 83 86 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=11.51 $Y=0
+ $X2=11.28 $Y2=0
r160 82 101 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.84 $Y=0
+ $X2=10.32 $Y2=0
r161 81 82 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=9.84 $Y=0
+ $X2=9.84 $Y2=0
r162 79 82 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=7.92 $Y=0
+ $X2=9.84 $Y2=0
r163 79 98 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=0 $X2=7.44
+ $Y2=0
r164 78 81 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=7.92 $Y=0 $X2=9.84
+ $Y2=0
r165 78 79 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=7.92 $Y=0
+ $X2=7.92 $Y2=0
r166 76 97 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.77 $Y=0 $X2=7.605
+ $Y2=0
r167 76 78 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=7.77 $Y=0 $X2=7.92
+ $Y2=0
r168 75 100 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.165 $Y=0
+ $X2=10.33 $Y2=0
r169 75 81 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=10.165 $Y=0
+ $X2=9.84 $Y2=0
r170 73 74 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r171 71 97 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.44 $Y=0 $X2=7.605
+ $Y2=0
r172 71 73 156.578 $w=1.68e-07 $l=2.4e-06 $layer=LI1_cond $X=7.44 $Y=0 $X2=5.04
+ $Y2=0
r173 70 74 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=5.04
+ $Y2=0
r174 69 70 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r175 67 70 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.56
+ $Y2=0
r176 66 67 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r177 64 67 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=1.2 $Y=0 $X2=3.6
+ $Y2=0
r178 64 95 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r179 63 66 156.578 $w=1.68e-07 $l=2.4e-06 $layer=LI1_cond $X=1.2 $Y=0 $X2=3.6
+ $Y2=0
r180 63 64 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r181 61 94 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.875 $Y=0 $X2=0.71
+ $Y2=0
r182 61 63 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.875 $Y=0 $X2=1.2
+ $Y2=0
r183 59 95 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r184 58 59 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r185 56 94 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.545 $Y=0 $X2=0.71
+ $Y2=0
r186 56 58 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.545 $Y=0
+ $X2=0.24 $Y2=0
r187 54 98 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=0 $X2=7.44
+ $Y2=0
r188 54 74 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=6.96 $Y=0
+ $X2=5.04 $Y2=0
r189 52 69 6.52406 $w=1.68e-07 $l=1e-07 $layer=LI1_cond $X=4.66 $Y=0 $X2=4.56
+ $Y2=0
r190 52 53 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.66 $Y=0 $X2=4.825
+ $Y2=0
r191 51 73 3.26203 $w=1.68e-07 $l=5e-08 $layer=LI1_cond $X=4.99 $Y=0 $X2=5.04
+ $Y2=0
r192 51 53 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.99 $Y=0 $X2=4.825
+ $Y2=0
r193 49 66 4.56684 $w=1.68e-07 $l=7e-08 $layer=LI1_cond $X=3.67 $Y=0 $X2=3.6
+ $Y2=0
r194 49 50 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.67 $Y=0 $X2=3.835
+ $Y2=0
r195 48 69 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=4 $Y=0 $X2=4.56
+ $Y2=0
r196 48 50 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4 $Y=0 $X2=3.835
+ $Y2=0
r197 44 110 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=13.205 $Y=0.085
+ $X2=13.205 $Y2=0
r198 44 46 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=13.205 $Y=0.085
+ $X2=13.205 $Y2=0.515
r199 43 104 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.84 $Y=0
+ $X2=11.675 $Y2=0
r200 42 110 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=13.12 $Y=0
+ $X2=13.205 $Y2=0
r201 42 43 83.508 $w=1.68e-07 $l=1.28e-06 $layer=LI1_cond $X=13.12 $Y=0
+ $X2=11.84 $Y2=0
r202 38 100 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=10.33 $Y=0.085
+ $X2=10.33 $Y2=0
r203 38 40 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=10.33 $Y=0.085
+ $X2=10.33 $Y2=0.58
r204 34 97 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.605 $Y=0.085
+ $X2=7.605 $Y2=0
r205 34 36 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=7.605 $Y=0.085
+ $X2=7.605 $Y2=0.34
r206 30 53 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.825 $Y=0.085
+ $X2=4.825 $Y2=0
r207 30 32 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=4.825 $Y=0.085
+ $X2=4.825 $Y2=0.55
r208 26 50 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.835 $Y=0.085
+ $X2=3.835 $Y2=0
r209 26 28 17.4613 $w=3.28e-07 $l=5e-07 $layer=LI1_cond $X=3.835 $Y=0.085
+ $X2=3.835 $Y2=0.585
r210 22 94 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.71 $Y=0.085
+ $X2=0.71 $Y2=0
r211 22 24 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=0.71 $Y=0.085
+ $X2=0.71 $Y2=0.58
r212 7 46 91 $w=1.7e-07 $l=2.62678e-07 $layer=licon1_NDIFF $count=2 $X=13.005
+ $Y=0.37 $X2=13.205 $Y2=0.515
r213 6 107 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=11.535
+ $Y=0.18 $X2=11.675 $Y2=0.325
r214 5 40 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=10.19
+ $Y=0.37 $X2=10.33 $Y2=0.58
r215 4 36 182 $w=1.7e-07 $l=2.83373e-07 $layer=licon1_NDIFF $count=1 $X=7.385
+ $Y=0.485 $X2=7.605 $Y2=0.34
r216 3 32 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=4.685
+ $Y=0.37 $X2=4.825 $Y2=0.55
r217 2 28 182 $w=1.7e-07 $l=2.41868e-07 $layer=licon1_NDIFF $count=1 $X=3.655
+ $Y=0.44 $X2=3.835 $Y2=0.585
r218 1 24 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.37 $X2=0.71 $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_HS__SDFRBP_1%noxref_25 1 2 9 11 12 13
r31 13 16 8.55602 $w=3.28e-07 $l=2.45e-07 $layer=LI1_cond $X=3.335 $Y=0.34
+ $X2=3.335 $Y2=0.585
r32 11 13 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.17 $Y=0.34
+ $X2=3.335 $Y2=0.34
r33 11 12 118.412 $w=1.68e-07 $l=1.815e-06 $layer=LI1_cond $X=3.17 $Y=0.34
+ $X2=1.355 $Y2=0.34
r34 7 12 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.23 $Y=0.425
+ $X2=1.355 $Y2=0.34
r35 7 9 8.98906 $w=2.48e-07 $l=1.95e-07 $layer=LI1_cond $X=1.23 $Y=0.425
+ $X2=1.23 $Y2=0.62
r36 2 16 182 $w=1.7e-07 $l=2.6533e-07 $layer=licon1_NDIFF $count=1 $X=3.115
+ $Y=0.485 $X2=3.335 $Y2=0.585
r37 1 9 182 $w=1.7e-07 $l=2.31409e-07 $layer=licon1_NDIFF $count=1 $X=1.125
+ $Y=0.45 $X2=1.27 $Y2=0.62
.ends

