* File: sky130_fd_sc_hs__o2111a_4.pxi.spice
* Created: Tue Sep  1 20:13:10 2020
* 
x_PM_SKY130_FD_SC_HS__O2111A_4%D1 N_D1_M1019_g N_D1_c_150_n N_D1_M1004_g
+ N_D1_c_151_n N_D1_M1020_g N_D1_c_157_n N_D1_M1011_g N_D1_c_153_n D1
+ N_D1_c_154_n PM_SKY130_FD_SC_HS__O2111A_4%D1
x_PM_SKY130_FD_SC_HS__O2111A_4%C1 N_C1_c_206_n N_C1_M1005_g N_C1_c_210_n
+ N_C1_M1006_g N_C1_c_207_n N_C1_M1017_g N_C1_c_211_n N_C1_M1007_g C1 C1
+ N_C1_c_209_n PM_SKY130_FD_SC_HS__O2111A_4%C1
x_PM_SKY130_FD_SC_HS__O2111A_4%B1 N_B1_c_262_n N_B1_M1008_g N_B1_M1009_g
+ N_B1_c_263_n N_B1_M1012_g N_B1_M1025_g B1 N_B1_c_261_n
+ PM_SKY130_FD_SC_HS__O2111A_4%B1
x_PM_SKY130_FD_SC_HS__O2111A_4%A2 N_A2_c_312_n N_A2_M1015_g N_A2_M1014_g
+ N_A2_c_313_n N_A2_M1016_g N_A2_M1027_g A2 A2 A2 A2 N_A2_c_311_n
+ PM_SKY130_FD_SC_HS__O2111A_4%A2
x_PM_SKY130_FD_SC_HS__O2111A_4%A1 N_A1_M1010_g N_A1_c_363_n N_A1_M1000_g
+ N_A1_M1022_g N_A1_c_364_n N_A1_M1002_g A1 N_A1_c_362_n
+ PM_SKY130_FD_SC_HS__O2111A_4%A1
x_PM_SKY130_FD_SC_HS__O2111A_4%A_27_392# N_A_27_392#_M1019_d N_A_27_392#_M1004_d
+ N_A_27_392#_M1011_d N_A_27_392#_M1007_d N_A_27_392#_M1012_s
+ N_A_27_392#_M1016_d N_A_27_392#_M1013_g N_A_27_392#_c_418_n
+ N_A_27_392#_M1001_g N_A_27_392#_M1018_g N_A_27_392#_c_419_n
+ N_A_27_392#_M1003_g N_A_27_392#_M1021_g N_A_27_392#_c_420_n
+ N_A_27_392#_M1024_g N_A_27_392#_c_410_n N_A_27_392#_c_411_n
+ N_A_27_392#_M1023_g N_A_27_392#_c_413_n N_A_27_392#_c_423_n
+ N_A_27_392#_M1026_g N_A_27_392#_c_414_n N_A_27_392#_c_424_n
+ N_A_27_392#_c_415_n N_A_27_392#_c_426_n N_A_27_392#_c_427_n
+ N_A_27_392#_c_428_n N_A_27_392#_c_429_n N_A_27_392#_c_430_n
+ N_A_27_392#_c_431_n N_A_27_392#_c_432_n N_A_27_392#_c_433_n
+ N_A_27_392#_c_416_n N_A_27_392#_c_568_p N_A_27_392#_c_434_n
+ N_A_27_392#_c_417_n N_A_27_392#_c_507_p N_A_27_392#_c_435_n
+ N_A_27_392#_c_436_n N_A_27_392#_c_437_n N_A_27_392#_c_438_n
+ PM_SKY130_FD_SC_HS__O2111A_4%A_27_392#
x_PM_SKY130_FD_SC_HS__O2111A_4%VPWR N_VPWR_M1004_s N_VPWR_M1006_s N_VPWR_M1008_d
+ N_VPWR_M1000_s N_VPWR_M1002_s N_VPWR_M1003_s N_VPWR_M1026_s N_VPWR_c_631_n
+ N_VPWR_c_632_n N_VPWR_c_633_n N_VPWR_c_634_n N_VPWR_c_635_n N_VPWR_c_636_n
+ N_VPWR_c_637_n N_VPWR_c_638_n N_VPWR_c_639_n N_VPWR_c_640_n N_VPWR_c_641_n
+ N_VPWR_c_642_n N_VPWR_c_643_n VPWR N_VPWR_c_644_n N_VPWR_c_645_n
+ N_VPWR_c_646_n N_VPWR_c_647_n N_VPWR_c_648_n N_VPWR_c_649_n N_VPWR_c_650_n
+ N_VPWR_c_651_n N_VPWR_c_630_n PM_SKY130_FD_SC_HS__O2111A_4%VPWR
x_PM_SKY130_FD_SC_HS__O2111A_4%A_747_392# N_A_747_392#_M1015_s
+ N_A_747_392#_M1000_d N_A_747_392#_c_753_n N_A_747_392#_c_756_n
+ N_A_747_392#_c_754_n PM_SKY130_FD_SC_HS__O2111A_4%A_747_392#
x_PM_SKY130_FD_SC_HS__O2111A_4%X N_X_M1013_d N_X_M1021_d N_X_M1001_d N_X_M1024_d
+ N_X_c_776_n N_X_c_791_n N_X_c_785_n N_X_c_777_n N_X_c_778_n N_X_c_803_n
+ N_X_c_779_n N_X_c_786_n N_X_c_787_n N_X_c_780_n N_X_c_781_n N_X_c_782_n
+ N_X_c_783_n N_X_c_829_n X PM_SKY130_FD_SC_HS__O2111A_4%X
x_PM_SKY130_FD_SC_HS__O2111A_4%A_27_74# N_A_27_74#_M1019_s N_A_27_74#_M1020_s
+ N_A_27_74#_M1017_s N_A_27_74#_c_858_n N_A_27_74#_c_859_n N_A_27_74#_c_860_n
+ N_A_27_74#_c_861_n N_A_27_74#_c_862_n N_A_27_74#_c_863_n N_A_27_74#_c_864_n
+ PM_SKY130_FD_SC_HS__O2111A_4%A_27_74#
x_PM_SKY130_FD_SC_HS__O2111A_4%A_287_74# N_A_287_74#_M1005_d N_A_287_74#_M1009_d
+ N_A_287_74#_c_897_n N_A_287_74#_c_898_n N_A_287_74#_c_899_n
+ PM_SKY130_FD_SC_HS__O2111A_4%A_287_74#
x_PM_SKY130_FD_SC_HS__O2111A_4%A_477_198# N_A_477_198#_M1009_s
+ N_A_477_198#_M1025_s N_A_477_198#_M1027_d N_A_477_198#_M1010_d
+ N_A_477_198#_c_926_n N_A_477_198#_c_936_n N_A_477_198#_c_927_n
+ N_A_477_198#_c_946_n N_A_477_198#_c_928_n N_A_477_198#_c_929_n
+ N_A_477_198#_c_930_n N_A_477_198#_c_931_n N_A_477_198#_c_932_n
+ N_A_477_198#_c_933_n PM_SKY130_FD_SC_HS__O2111A_4%A_477_198#
x_PM_SKY130_FD_SC_HS__O2111A_4%VGND N_VGND_M1014_s N_VGND_M1010_s N_VGND_M1022_s
+ N_VGND_M1018_s N_VGND_M1023_s N_VGND_c_990_n N_VGND_c_991_n N_VGND_c_992_n
+ N_VGND_c_993_n N_VGND_c_994_n N_VGND_c_995_n N_VGND_c_996_n N_VGND_c_997_n
+ N_VGND_c_998_n N_VGND_c_999_n N_VGND_c_1000_n N_VGND_c_1001_n VGND
+ N_VGND_c_1002_n N_VGND_c_1003_n N_VGND_c_1004_n N_VGND_c_1005_n
+ PM_SKY130_FD_SC_HS__O2111A_4%VGND
cc_1 VNB N_D1_M1019_g 0.0398087f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=0.74
cc_2 VNB N_D1_c_150_n 0.0244877f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.885
cc_3 VNB N_D1_c_151_n 0.00812914f $X=-0.19 $Y=-0.245 $X2=0.855 $Y2=1.705
cc_4 VNB N_D1_M1020_g 0.0367314f $X=-0.19 $Y=-0.245 $X2=0.93 $Y2=0.74
cc_5 VNB N_D1_c_153_n 0.00691334f $X=-0.19 $Y=-0.245 $X2=0.93 $Y2=1.757
cc_6 VNB N_D1_c_154_n 0.00919084f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.615
cc_7 VNB N_C1_c_206_n 0.014489f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=1.45
cc_8 VNB N_C1_c_207_n 0.0173034f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.38
cc_9 VNB C1 0.00620616f $X=-0.19 $Y=-0.245 $X2=1.055 $Y2=1.885
cc_10 VNB N_C1_c_209_n 0.0710768f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.615
cc_11 VNB N_B1_M1009_g 0.0254353f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.38
cc_12 VNB N_B1_M1025_g 0.0198802f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB B1 9.27509e-19 $X=-0.19 $Y=-0.245 $X2=1.055 $Y2=2.38
cc_14 VNB N_B1_c_261_n 0.0327986f $X=-0.19 $Y=-0.245 $X2=0.407 $Y2=1.615
cc_15 VNB N_A2_M1014_g 0.0201199f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.38
cc_16 VNB N_A2_M1027_g 0.026686f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB A2 0.0142547f $X=-0.19 $Y=-0.245 $X2=1.055 $Y2=1.757
cc_18 VNB N_A2_c_311_n 0.0284336f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.615
cc_19 VNB N_A1_M1010_g 0.0363489f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=0.74
cc_20 VNB N_A1_M1022_g 0.0297668f $X=-0.19 $Y=-0.245 $X2=0.93 $Y2=1.63
cc_21 VNB A1 9.25683e-19 $X=-0.19 $Y=-0.245 $X2=1.055 $Y2=2.38
cc_22 VNB N_A1_c_362_n 0.0276131f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.615
cc_23 VNB N_A_27_392#_M1013_g 0.024894f $X=-0.19 $Y=-0.245 $X2=0.407 $Y2=1.615
cc_24 VNB N_A_27_392#_M1018_g 0.024924f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.615
cc_25 VNB N_A_27_392#_M1021_g 0.0249207f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_27_392#_c_410_n 0.00880736f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_27_392#_c_411_n 0.0557112f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_27_392#_M1023_g 0.0255042f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_27_392#_c_413_n 0.00983424f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_27_392#_c_414_n 0.00852688f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_27_392#_c_415_n 0.00406729f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_27_392#_c_416_n 0.00516444f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_27_392#_c_417_n 0.00199603f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_VPWR_c_630_n 0.342803f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_X_c_776_n 0.00240191f $X=-0.19 $Y=-0.245 $X2=1.055 $Y2=2.38
cc_36 VNB N_X_c_777_n 0.00323083f $X=-0.19 $Y=-0.245 $X2=0.407 $Y2=1.615
cc_37 VNB N_X_c_778_n 0.00230427f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.615
cc_38 VNB N_X_c_779_n 0.00240191f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_X_c_780_n 0.00997592f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_X_c_781_n 0.0126045f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_X_c_782_n 8.8527e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_X_c_783_n 0.00273044f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB X 0.0155405f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_27_74#_c_858_n 0.0167032f $X=-0.19 $Y=-0.245 $X2=0.93 $Y2=1.63
cc_45 VNB N_A_27_74#_c_859_n 0.0219399f $X=-0.19 $Y=-0.245 $X2=0.93 $Y2=0.74
cc_46 VNB N_A_27_74#_c_860_n 0.00272448f $X=-0.19 $Y=-0.245 $X2=1.055 $Y2=1.885
cc_47 VNB N_A_27_74#_c_861_n 0.00226074f $X=-0.19 $Y=-0.245 $X2=1.055 $Y2=1.757
cc_48 VNB N_A_27_74#_c_862_n 0.00123754f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.615
cc_49 VNB N_A_27_74#_c_863_n 0.00987713f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_A_27_74#_c_864_n 0.0027795f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.615
cc_51 VNB N_A_287_74#_c_897_n 0.0168718f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.38
cc_52 VNB N_A_287_74#_c_898_n 0.00289336f $X=-0.19 $Y=-0.245 $X2=0.93 $Y2=0.74
cc_53 VNB N_A_287_74#_c_899_n 0.00264166f $X=-0.19 $Y=-0.245 $X2=1.055 $Y2=1.885
cc_54 VNB N_A_477_198#_c_926_n 0.0080669f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_A_477_198#_c_927_n 0.00267457f $X=-0.19 $Y=-0.245 $X2=0.407
+ $Y2=1.615
cc_56 VNB N_A_477_198#_c_928_n 0.0101622f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_A_477_198#_c_929_n 0.0252068f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_A_477_198#_c_930_n 0.00178908f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_A_477_198#_c_931_n 0.00108544f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_A_477_198#_c_932_n 0.00230918f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_A_477_198#_c_933_n 0.0025485f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_VGND_c_990_n 0.0206912f $X=-0.19 $Y=-0.245 $X2=1.055 $Y2=1.757
cc_63 VNB N_VGND_c_991_n 0.0166086f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.615
cc_64 VNB N_VGND_c_992_n 0.0154673f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_VGND_c_993_n 0.00830803f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_VGND_c_994_n 0.0131737f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_VGND_c_995_n 0.029666f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_VGND_c_996_n 0.0952344f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_VGND_c_997_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_VGND_c_998_n 0.0151736f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_VGND_c_999_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_VGND_c_1000_n 0.0186948f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_VGND_c_1001_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_VGND_c_1002_n 0.0222872f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_VGND_c_1003_n 0.0186948f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_VGND_c_1004_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_VGND_c_1005_n 0.456094f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VPB N_D1_c_150_n 0.0436497f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.885
cc_79 VPB N_D1_c_151_n 0.00985951f $X=-0.19 $Y=1.66 $X2=0.855 $Y2=1.705
cc_80 VPB N_D1_c_157_n 0.0157133f $X=-0.19 $Y=1.66 $X2=1.055 $Y2=1.885
cc_81 VPB N_D1_c_153_n 0.0150067f $X=-0.19 $Y=1.66 $X2=0.93 $Y2=1.757
cc_82 VPB N_D1_c_154_n 0.0054581f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.615
cc_83 VPB N_C1_c_210_n 0.0154054f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_84 VPB N_C1_c_211_n 0.0161168f $X=-0.19 $Y=1.66 $X2=0.93 $Y2=1.63
cc_85 VPB C1 0.00250401f $X=-0.19 $Y=1.66 $X2=1.055 $Y2=1.885
cc_86 VPB N_C1_c_209_n 0.0356219f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.615
cc_87 VPB N_B1_c_262_n 0.0157358f $X=-0.19 $Y=1.66 $X2=0.5 $Y2=1.45
cc_88 VPB N_B1_c_263_n 0.0154596f $X=-0.19 $Y=1.66 $X2=0.855 $Y2=1.705
cc_89 VPB B1 0.00138027f $X=-0.19 $Y=1.66 $X2=1.055 $Y2=2.38
cc_90 VPB N_B1_c_261_n 0.041099f $X=-0.19 $Y=1.66 $X2=0.407 $Y2=1.615
cc_91 VPB N_A2_c_312_n 0.0173428f $X=-0.19 $Y=1.66 $X2=0.5 $Y2=1.45
cc_92 VPB N_A2_c_313_n 0.018883f $X=-0.19 $Y=1.66 $X2=0.855 $Y2=1.705
cc_93 VPB A2 0.0119806f $X=-0.19 $Y=1.66 $X2=1.055 $Y2=1.757
cc_94 VPB N_A2_c_311_n 0.0384902f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.615
cc_95 VPB N_A1_c_363_n 0.0179782f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.885
cc_96 VPB N_A1_c_364_n 0.0163389f $X=-0.19 $Y=1.66 $X2=0.93 $Y2=0.74
cc_97 VPB A1 0.00235587f $X=-0.19 $Y=1.66 $X2=1.055 $Y2=2.38
cc_98 VPB N_A1_c_362_n 0.038041f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.615
cc_99 VPB N_A_27_392#_c_418_n 0.0157919f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.615
cc_100 VPB N_A_27_392#_c_419_n 0.0154901f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_101 VPB N_A_27_392#_c_420_n 0.0150811f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_102 VPB N_A_27_392#_c_411_n 0.0351244f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_103 VPB N_A_27_392#_c_413_n 0.00111912f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_104 VPB N_A_27_392#_c_423_n 0.0257552f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_105 VPB N_A_27_392#_c_424_n 0.00132673f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_106 VPB N_A_27_392#_c_415_n 0.00313061f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_107 VPB N_A_27_392#_c_426_n 8.4684e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_108 VPB N_A_27_392#_c_427_n 0.00456859f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_109 VPB N_A_27_392#_c_428_n 0.00433366f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_110 VPB N_A_27_392#_c_429_n 7.2018e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_111 VPB N_A_27_392#_c_430_n 0.0208557f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_112 VPB N_A_27_392#_c_431_n 0.00273412f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_113 VPB N_A_27_392#_c_432_n 0.00484195f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_114 VPB N_A_27_392#_c_433_n 0.00136802f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_115 VPB N_A_27_392#_c_434_n 0.0397524f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_116 VPB N_A_27_392#_c_435_n 0.0058322f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_117 VPB N_A_27_392#_c_436_n 0.0151238f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_118 VPB N_A_27_392#_c_437_n 0.00403686f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_119 VPB N_A_27_392#_c_438_n 0.00697293f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_120 VPB N_VPWR_c_631_n 0.0191693f $X=-0.19 $Y=1.66 $X2=0.407 $Y2=1.705
cc_121 VPB N_VPWR_c_632_n 0.0193866f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_122 VPB N_VPWR_c_633_n 0.0158144f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_123 VPB N_VPWR_c_634_n 0.0127873f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_124 VPB N_VPWR_c_635_n 0.0128087f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_125 VPB N_VPWR_c_636_n 0.00599091f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_126 VPB N_VPWR_c_637_n 0.00274649f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_127 VPB N_VPWR_c_638_n 0.0121909f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_128 VPB N_VPWR_c_639_n 0.0594132f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_129 VPB N_VPWR_c_640_n 0.0216142f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_130 VPB N_VPWR_c_641_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_131 VPB N_VPWR_c_642_n 0.0432956f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_132 VPB N_VPWR_c_643_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_133 VPB N_VPWR_c_644_n 0.0198433f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_134 VPB N_VPWR_c_645_n 0.0198086f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_135 VPB N_VPWR_c_646_n 0.0172173f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_136 VPB N_VPWR_c_647_n 0.0175706f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_137 VPB N_VPWR_c_648_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_138 VPB N_VPWR_c_649_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_139 VPB N_VPWR_c_650_n 0.00614127f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_140 VPB N_VPWR_c_651_n 0.00601644f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_141 VPB N_VPWR_c_630_n 0.117049f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_142 VPB N_A_747_392#_c_753_n 0.0124765f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.38
cc_143 VPB N_A_747_392#_c_754_n 0.00257417f $X=-0.19 $Y=1.66 $X2=0.93 $Y2=1.757
cc_144 VPB N_X_c_785_n 0.00275689f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_145 VPB N_X_c_786_n 0.00163506f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_146 VPB N_X_c_787_n 0.00216998f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_147 N_D1_M1020_g N_C1_c_206_n 0.0187348f $X=0.93 $Y=0.74 $X2=-0.19 $Y2=-0.245
cc_148 N_D1_c_157_n N_C1_c_210_n 0.0144223f $X=1.055 $Y=1.885 $X2=0 $Y2=0
cc_149 N_D1_M1020_g C1 0.00173097f $X=0.93 $Y=0.74 $X2=0 $Y2=0
cc_150 N_D1_c_153_n C1 0.00672465f $X=0.93 $Y=1.757 $X2=0 $Y2=0
cc_151 N_D1_M1020_g N_C1_c_209_n 0.00802884f $X=0.93 $Y=0.74 $X2=0 $Y2=0
cc_152 N_D1_c_153_n N_C1_c_209_n 0.0124404f $X=0.93 $Y=1.757 $X2=0 $Y2=0
cc_153 N_D1_c_150_n N_A_27_392#_c_424_n 0.0140774f $X=0.505 $Y=1.885 $X2=0 $Y2=0
cc_154 N_D1_c_151_n N_A_27_392#_c_424_n 0.00424535f $X=0.855 $Y=1.705 $X2=0
+ $Y2=0
cc_155 N_D1_c_154_n N_A_27_392#_c_424_n 0.00746443f $X=0.385 $Y=1.615 $X2=0
+ $Y2=0
cc_156 N_D1_M1019_g N_A_27_392#_c_415_n 0.00680216f $X=0.5 $Y=0.74 $X2=0 $Y2=0
cc_157 N_D1_c_150_n N_A_27_392#_c_415_n 0.00508079f $X=0.505 $Y=1.885 $X2=0
+ $Y2=0
cc_158 N_D1_c_151_n N_A_27_392#_c_415_n 0.00987117f $X=0.855 $Y=1.705 $X2=0
+ $Y2=0
cc_159 N_D1_M1020_g N_A_27_392#_c_415_n 0.0114191f $X=0.93 $Y=0.74 $X2=0 $Y2=0
cc_160 N_D1_c_157_n N_A_27_392#_c_415_n 0.00155171f $X=1.055 $Y=1.885 $X2=0
+ $Y2=0
cc_161 N_D1_c_153_n N_A_27_392#_c_415_n 0.00585164f $X=0.93 $Y=1.757 $X2=0 $Y2=0
cc_162 N_D1_c_154_n N_A_27_392#_c_415_n 0.0247006f $X=0.385 $Y=1.615 $X2=0 $Y2=0
cc_163 N_D1_c_157_n N_A_27_392#_c_426_n 0.0154073f $X=1.055 $Y=1.885 $X2=0 $Y2=0
cc_164 N_D1_c_153_n N_A_27_392#_c_426_n 0.0037937f $X=0.93 $Y=1.757 $X2=0 $Y2=0
cc_165 N_D1_c_150_n N_A_27_392#_c_434_n 0.0178942f $X=0.505 $Y=1.885 $X2=0 $Y2=0
cc_166 N_D1_c_157_n N_A_27_392#_c_434_n 7.02865e-19 $X=1.055 $Y=1.885 $X2=0
+ $Y2=0
cc_167 N_D1_c_154_n N_A_27_392#_c_434_n 0.027311f $X=0.385 $Y=1.615 $X2=0 $Y2=0
cc_168 N_D1_M1019_g N_A_27_392#_c_417_n 0.00603749f $X=0.5 $Y=0.74 $X2=0 $Y2=0
cc_169 N_D1_c_150_n N_A_27_392#_c_417_n 7.30743e-19 $X=0.505 $Y=1.885 $X2=0
+ $Y2=0
cc_170 N_D1_c_151_n N_A_27_392#_c_417_n 0.00331039f $X=0.855 $Y=1.705 $X2=0
+ $Y2=0
cc_171 N_D1_M1020_g N_A_27_392#_c_417_n 0.00453298f $X=0.93 $Y=0.74 $X2=0 $Y2=0
cc_172 N_D1_c_150_n N_A_27_392#_c_435_n 7.02865e-19 $X=0.505 $Y=1.885 $X2=0
+ $Y2=0
cc_173 N_D1_c_157_n N_A_27_392#_c_435_n 0.0114959f $X=1.055 $Y=1.885 $X2=0 $Y2=0
cc_174 N_D1_c_153_n N_A_27_392#_c_435_n 3.77791e-19 $X=0.93 $Y=1.757 $X2=0 $Y2=0
cc_175 N_D1_c_150_n N_VPWR_c_631_n 0.00630009f $X=0.505 $Y=1.885 $X2=0 $Y2=0
cc_176 N_D1_c_151_n N_VPWR_c_631_n 8.20775e-19 $X=0.855 $Y=1.705 $X2=0 $Y2=0
cc_177 N_D1_c_157_n N_VPWR_c_631_n 0.00489938f $X=1.055 $Y=1.885 $X2=0 $Y2=0
cc_178 N_D1_c_157_n N_VPWR_c_632_n 0.00458031f $X=1.055 $Y=1.885 $X2=0 $Y2=0
cc_179 N_D1_c_150_n N_VPWR_c_644_n 0.00458031f $X=0.505 $Y=1.885 $X2=0 $Y2=0
cc_180 N_D1_c_150_n N_VPWR_c_630_n 0.0049649f $X=0.505 $Y=1.885 $X2=0 $Y2=0
cc_181 N_D1_c_157_n N_VPWR_c_630_n 0.0049649f $X=1.055 $Y=1.885 $X2=0 $Y2=0
cc_182 N_D1_M1019_g N_A_27_74#_c_859_n 9.80934e-19 $X=0.5 $Y=0.74 $X2=0 $Y2=0
cc_183 N_D1_c_150_n N_A_27_74#_c_859_n 0.00335778f $X=0.505 $Y=1.885 $X2=0 $Y2=0
cc_184 N_D1_c_154_n N_A_27_74#_c_859_n 0.0133432f $X=0.385 $Y=1.615 $X2=0 $Y2=0
cc_185 N_D1_M1019_g N_A_27_74#_c_860_n 0.0182491f $X=0.5 $Y=0.74 $X2=0 $Y2=0
cc_186 N_D1_M1020_g N_A_27_74#_c_860_n 0.0169848f $X=0.93 $Y=0.74 $X2=0 $Y2=0
cc_187 N_D1_M1020_g N_A_27_74#_c_861_n 3.89484e-19 $X=0.93 $Y=0.74 $X2=0 $Y2=0
cc_188 N_D1_c_153_n N_A_27_74#_c_861_n 0.00113532f $X=0.93 $Y=1.757 $X2=0 $Y2=0
cc_189 N_D1_M1019_g N_VGND_c_996_n 0.00278271f $X=0.5 $Y=0.74 $X2=0 $Y2=0
cc_190 N_D1_M1020_g N_VGND_c_996_n 0.00278271f $X=0.93 $Y=0.74 $X2=0 $Y2=0
cc_191 N_D1_M1019_g N_VGND_c_1005_n 0.00357103f $X=0.5 $Y=0.74 $X2=0 $Y2=0
cc_192 N_D1_M1020_g N_VGND_c_1005_n 0.00353526f $X=0.93 $Y=0.74 $X2=0 $Y2=0
cc_193 N_C1_c_211_n N_B1_c_262_n 0.0191061f $X=2.005 $Y=1.885 $X2=-0.19
+ $Y2=-0.245
cc_194 N_C1_c_209_n N_B1_c_261_n 0.0151976f $X=1.79 $Y=1.535 $X2=0 $Y2=0
cc_195 C1 N_A_27_392#_c_415_n 0.0232485f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_196 N_C1_c_209_n N_A_27_392#_c_415_n 0.00145788f $X=1.79 $Y=1.535 $X2=0 $Y2=0
cc_197 C1 N_A_27_392#_c_426_n 0.00210849f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_198 N_C1_c_210_n N_A_27_392#_c_427_n 0.0122806f $X=1.505 $Y=1.885 $X2=0 $Y2=0
cc_199 N_C1_c_211_n N_A_27_392#_c_427_n 0.0201067f $X=2.005 $Y=1.885 $X2=0 $Y2=0
cc_200 C1 N_A_27_392#_c_427_n 0.0257653f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_201 N_C1_c_209_n N_A_27_392#_c_427_n 0.0117775f $X=1.79 $Y=1.535 $X2=0 $Y2=0
cc_202 N_C1_c_206_n N_A_27_392#_c_417_n 6.23466e-19 $X=1.36 $Y=1.185 $X2=0 $Y2=0
cc_203 N_C1_c_210_n N_A_27_392#_c_435_n 0.0112639f $X=1.505 $Y=1.885 $X2=0 $Y2=0
cc_204 N_C1_c_211_n N_A_27_392#_c_435_n 0.00101598f $X=2.005 $Y=1.885 $X2=0
+ $Y2=0
cc_205 C1 N_A_27_392#_c_435_n 0.028809f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_206 N_C1_c_209_n N_A_27_392#_c_435_n 4.63579e-19 $X=1.79 $Y=1.535 $X2=0 $Y2=0
cc_207 N_C1_c_211_n N_A_27_392#_c_436_n 0.01097f $X=2.005 $Y=1.885 $X2=0 $Y2=0
cc_208 N_C1_c_210_n N_VPWR_c_632_n 0.00458031f $X=1.505 $Y=1.885 $X2=0 $Y2=0
cc_209 N_C1_c_210_n N_VPWR_c_633_n 0.00451095f $X=1.505 $Y=1.885 $X2=0 $Y2=0
cc_210 N_C1_c_211_n N_VPWR_c_633_n 0.0112032f $X=2.005 $Y=1.885 $X2=0 $Y2=0
cc_211 N_C1_c_211_n N_VPWR_c_634_n 5.85107e-19 $X=2.005 $Y=1.885 $X2=0 $Y2=0
cc_212 N_C1_c_211_n N_VPWR_c_640_n 0.00421101f $X=2.005 $Y=1.885 $X2=0 $Y2=0
cc_213 N_C1_c_210_n N_VPWR_c_630_n 0.0049649f $X=1.505 $Y=1.885 $X2=0 $Y2=0
cc_214 N_C1_c_211_n N_VPWR_c_630_n 0.00450151f $X=2.005 $Y=1.885 $X2=0 $Y2=0
cc_215 N_C1_c_206_n N_A_27_74#_c_861_n 4.08775e-19 $X=1.36 $Y=1.185 $X2=0 $Y2=0
cc_216 C1 N_A_27_74#_c_861_n 0.00820373f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_217 N_C1_c_206_n N_A_27_74#_c_864_n 0.0122675f $X=1.36 $Y=1.185 $X2=0 $Y2=0
cc_218 N_C1_c_207_n N_A_27_74#_c_864_n 0.0113109f $X=1.79 $Y=1.185 $X2=0 $Y2=0
cc_219 N_C1_c_207_n N_A_287_74#_c_897_n 0.0127544f $X=1.79 $Y=1.185 $X2=0 $Y2=0
cc_220 C1 N_A_287_74#_c_897_n 0.00143794f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_221 N_C1_c_209_n N_A_287_74#_c_897_n 0.00546102f $X=1.79 $Y=1.535 $X2=0 $Y2=0
cc_222 N_C1_c_206_n N_A_287_74#_c_898_n 0.00805309f $X=1.36 $Y=1.185 $X2=0 $Y2=0
cc_223 N_C1_c_207_n N_A_287_74#_c_898_n 0.0169798f $X=1.79 $Y=1.185 $X2=0 $Y2=0
cc_224 C1 N_A_287_74#_c_898_n 0.0167849f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_225 N_C1_c_209_n N_A_287_74#_c_898_n 0.00333691f $X=1.79 $Y=1.535 $X2=0 $Y2=0
cc_226 N_C1_c_207_n N_A_477_198#_c_926_n 0.00673386f $X=1.79 $Y=1.185 $X2=0
+ $Y2=0
cc_227 N_C1_c_206_n N_VGND_c_996_n 0.00278271f $X=1.36 $Y=1.185 $X2=0 $Y2=0
cc_228 N_C1_c_207_n N_VGND_c_996_n 0.00278271f $X=1.79 $Y=1.185 $X2=0 $Y2=0
cc_229 N_C1_c_206_n N_VGND_c_1005_n 0.00353526f $X=1.36 $Y=1.185 $X2=0 $Y2=0
cc_230 N_C1_c_207_n N_VGND_c_1005_n 0.00358427f $X=1.79 $Y=1.185 $X2=0 $Y2=0
cc_231 N_B1_c_263_n N_A2_c_312_n 0.0209644f $X=3.075 $Y=1.885 $X2=-0.19
+ $Y2=-0.245
cc_232 N_B1_M1025_g N_A2_M1014_g 0.0159516f $X=3.255 $Y=0.91 $X2=0 $Y2=0
cc_233 B1 A2 0.0276607f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_234 N_B1_c_261_n A2 0.00240023f $X=3.15 $Y=1.615 $X2=0 $Y2=0
cc_235 B1 N_A2_c_311_n 3.40273e-19 $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_236 N_B1_c_261_n N_A2_c_311_n 0.0222416f $X=3.15 $Y=1.615 $X2=0 $Y2=0
cc_237 N_B1_c_262_n N_A_27_392#_c_428_n 0.0170851f $X=2.625 $Y=1.885 $X2=0 $Y2=0
cc_238 N_B1_c_263_n N_A_27_392#_c_428_n 0.0154824f $X=3.075 $Y=1.885 $X2=0 $Y2=0
cc_239 B1 N_A_27_392#_c_428_n 0.0170742f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_240 N_B1_c_261_n N_A_27_392#_c_428_n 0.0103291f $X=3.15 $Y=1.615 $X2=0 $Y2=0
cc_241 N_B1_c_263_n N_A_27_392#_c_429_n 0.0112272f $X=3.075 $Y=1.885 $X2=0 $Y2=0
cc_242 N_B1_c_263_n N_A_27_392#_c_432_n 2.59907e-19 $X=3.075 $Y=1.885 $X2=0
+ $Y2=0
cc_243 N_B1_c_262_n N_A_27_392#_c_436_n 0.01097f $X=2.625 $Y=1.885 $X2=0 $Y2=0
cc_244 B1 N_A_27_392#_c_437_n 0.00796601f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_245 N_B1_c_261_n N_A_27_392#_c_437_n 0.00128085f $X=3.15 $Y=1.615 $X2=0 $Y2=0
cc_246 N_B1_c_262_n N_VPWR_c_633_n 5.85107e-19 $X=2.625 $Y=1.885 $X2=0 $Y2=0
cc_247 N_B1_c_262_n N_VPWR_c_634_n 0.0113303f $X=2.625 $Y=1.885 $X2=0 $Y2=0
cc_248 N_B1_c_263_n N_VPWR_c_634_n 0.010209f $X=3.075 $Y=1.885 $X2=0 $Y2=0
cc_249 N_B1_c_262_n N_VPWR_c_640_n 0.00421101f $X=2.625 $Y=1.885 $X2=0 $Y2=0
cc_250 N_B1_c_263_n N_VPWR_c_642_n 0.00421101f $X=3.075 $Y=1.885 $X2=0 $Y2=0
cc_251 N_B1_c_262_n N_VPWR_c_630_n 0.00450151f $X=2.625 $Y=1.885 $X2=0 $Y2=0
cc_252 N_B1_c_263_n N_VPWR_c_630_n 0.00450151f $X=3.075 $Y=1.885 $X2=0 $Y2=0
cc_253 N_B1_M1009_g N_A_27_74#_c_863_n 0.00324596f $X=2.825 $Y=0.91 $X2=0 $Y2=0
cc_254 N_B1_M1009_g N_A_287_74#_c_897_n 0.0109615f $X=2.825 $Y=0.91 $X2=0 $Y2=0
cc_255 N_B1_M1009_g N_A_287_74#_c_899_n 0.00936405f $X=2.825 $Y=0.91 $X2=0 $Y2=0
cc_256 N_B1_c_261_n N_A_477_198#_c_926_n 0.00526284f $X=3.15 $Y=1.615 $X2=0
+ $Y2=0
cc_257 N_B1_M1009_g N_A_477_198#_c_936_n 0.0102868f $X=2.825 $Y=0.91 $X2=0 $Y2=0
cc_258 N_B1_M1025_g N_A_477_198#_c_936_n 0.0125752f $X=3.255 $Y=0.91 $X2=0 $Y2=0
cc_259 B1 N_A_477_198#_c_936_n 0.0216895f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_260 N_B1_c_261_n N_A_477_198#_c_936_n 7.11881e-19 $X=3.15 $Y=1.615 $X2=0
+ $Y2=0
cc_261 N_B1_M1009_g N_A_477_198#_c_927_n 9.14331e-19 $X=2.825 $Y=0.91 $X2=0
+ $Y2=0
cc_262 N_B1_M1025_g N_A_477_198#_c_927_n 0.00758705f $X=3.255 $Y=0.91 $X2=0
+ $Y2=0
cc_263 N_B1_M1009_g N_A_477_198#_c_931_n 0.00222768f $X=2.825 $Y=0.91 $X2=0
+ $Y2=0
cc_264 N_B1_M1025_g N_A_477_198#_c_932_n 0.00103783f $X=3.255 $Y=0.91 $X2=0
+ $Y2=0
cc_265 B1 N_A_477_198#_c_932_n 7.22171e-19 $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_266 N_B1_M1025_g N_VGND_c_990_n 6.8897e-19 $X=3.255 $Y=0.91 $X2=0 $Y2=0
cc_267 N_B1_M1009_g N_VGND_c_996_n 0.00359961f $X=2.825 $Y=0.91 $X2=0 $Y2=0
cc_268 N_B1_M1025_g N_VGND_c_996_n 0.00444543f $X=3.255 $Y=0.91 $X2=0 $Y2=0
cc_269 N_B1_M1009_g N_VGND_c_1005_n 0.00493565f $X=2.825 $Y=0.91 $X2=0 $Y2=0
cc_270 N_B1_M1025_g N_VGND_c_1005_n 0.00493565f $X=3.255 $Y=0.91 $X2=0 $Y2=0
cc_271 A2 A1 0.0261825f $X=4.955 $Y=1.58 $X2=0 $Y2=0
cc_272 A2 N_A1_c_362_n 0.0143298f $X=4.955 $Y=1.58 $X2=0 $Y2=0
cc_273 N_A2_c_312_n N_A_27_392#_c_430_n 0.0157477f $X=3.66 $Y=1.885 $X2=0 $Y2=0
cc_274 N_A2_c_313_n N_A_27_392#_c_430_n 0.0129264f $X=4.16 $Y=1.885 $X2=0 $Y2=0
cc_275 A2 N_A_27_392#_c_430_n 0.123143f $X=4.955 $Y=1.58 $X2=0 $Y2=0
cc_276 N_A2_c_311_n N_A_27_392#_c_430_n 0.00954984f $X=4.16 $Y=1.667 $X2=0 $Y2=0
cc_277 N_A2_c_312_n N_A_27_392#_c_431_n 0.0151061f $X=3.66 $Y=1.885 $X2=0 $Y2=0
cc_278 N_A2_c_313_n N_A_27_392#_c_431_n 0.00887409f $X=4.16 $Y=1.885 $X2=0 $Y2=0
cc_279 A2 N_A_27_392#_c_437_n 0.00575f $X=4.955 $Y=1.58 $X2=0 $Y2=0
cc_280 N_A2_c_312_n N_A_27_392#_c_438_n 6.42635e-19 $X=3.66 $Y=1.885 $X2=0 $Y2=0
cc_281 N_A2_c_313_n N_A_27_392#_c_438_n 0.00758595f $X=4.16 $Y=1.885 $X2=0 $Y2=0
cc_282 N_A2_c_312_n N_VPWR_c_634_n 9.85938e-19 $X=3.66 $Y=1.885 $X2=0 $Y2=0
cc_283 N_A2_c_313_n N_VPWR_c_635_n 0.00133087f $X=4.16 $Y=1.885 $X2=0 $Y2=0
cc_284 N_A2_c_312_n N_VPWR_c_642_n 0.00278271f $X=3.66 $Y=1.885 $X2=0 $Y2=0
cc_285 N_A2_c_313_n N_VPWR_c_642_n 0.00279479f $X=4.16 $Y=1.885 $X2=0 $Y2=0
cc_286 N_A2_c_312_n N_VPWR_c_630_n 0.00359085f $X=3.66 $Y=1.885 $X2=0 $Y2=0
cc_287 N_A2_c_313_n N_VPWR_c_630_n 0.00358175f $X=4.16 $Y=1.885 $X2=0 $Y2=0
cc_288 N_A2_c_313_n N_A_747_392#_c_753_n 0.0127395f $X=4.16 $Y=1.885 $X2=0 $Y2=0
cc_289 N_A2_c_312_n N_A_747_392#_c_756_n 0.00534929f $X=3.66 $Y=1.885 $X2=0
+ $Y2=0
cc_290 N_A2_M1014_g N_A_477_198#_c_927_n 3.13308e-19 $X=3.685 $Y=0.91 $X2=0
+ $Y2=0
cc_291 N_A2_M1014_g N_A_477_198#_c_946_n 0.0125873f $X=3.685 $Y=0.91 $X2=0 $Y2=0
cc_292 N_A2_M1027_g N_A_477_198#_c_946_n 0.0122289f $X=4.175 $Y=0.91 $X2=0 $Y2=0
cc_293 A2 N_A_477_198#_c_946_n 0.0433751f $X=4.955 $Y=1.58 $X2=0 $Y2=0
cc_294 N_A2_c_311_n N_A_477_198#_c_946_n 0.00358729f $X=4.16 $Y=1.667 $X2=0
+ $Y2=0
cc_295 N_A2_M1014_g N_A_477_198#_c_928_n 9.05595e-19 $X=3.685 $Y=0.91 $X2=0
+ $Y2=0
cc_296 N_A2_M1027_g N_A_477_198#_c_928_n 0.00850927f $X=4.175 $Y=0.91 $X2=0
+ $Y2=0
cc_297 A2 N_A_477_198#_c_929_n 0.0465439f $X=4.955 $Y=1.58 $X2=0 $Y2=0
cc_298 A2 N_A_477_198#_c_932_n 0.00597859f $X=4.955 $Y=1.58 $X2=0 $Y2=0
cc_299 N_A2_M1027_g N_A_477_198#_c_933_n 4.27055e-19 $X=4.175 $Y=0.91 $X2=0
+ $Y2=0
cc_300 A2 N_A_477_198#_c_933_n 0.02594f $X=4.955 $Y=1.58 $X2=0 $Y2=0
cc_301 N_A2_M1014_g N_VGND_c_990_n 0.00895009f $X=3.685 $Y=0.91 $X2=0 $Y2=0
cc_302 N_A2_M1027_g N_VGND_c_990_n 0.00539056f $X=4.175 $Y=0.91 $X2=0 $Y2=0
cc_303 N_A2_M1027_g N_VGND_c_991_n 0.00356388f $X=4.175 $Y=0.91 $X2=0 $Y2=0
cc_304 N_A2_M1014_g N_VGND_c_996_n 0.00384833f $X=3.685 $Y=0.91 $X2=0 $Y2=0
cc_305 N_A2_M1027_g N_VGND_c_1002_n 0.00452252f $X=4.175 $Y=0.91 $X2=0 $Y2=0
cc_306 N_A2_M1014_g N_VGND_c_1005_n 0.00414594f $X=3.685 $Y=0.91 $X2=0 $Y2=0
cc_307 N_A2_M1027_g N_VGND_c_1005_n 0.00493565f $X=4.175 $Y=0.91 $X2=0 $Y2=0
cc_308 N_A1_M1022_g N_A_27_392#_M1013_g 0.0259675f $X=5.635 $Y=0.74 $X2=0 $Y2=0
cc_309 N_A1_c_362_n N_A_27_392#_c_418_n 0.0256329f $X=5.635 $Y=1.667 $X2=0 $Y2=0
cc_310 A1 N_A_27_392#_c_411_n 3.03891e-19 $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_311 N_A1_c_362_n N_A_27_392#_c_411_n 0.00961693f $X=5.635 $Y=1.667 $X2=0
+ $Y2=0
cc_312 N_A1_c_363_n N_A_27_392#_c_430_n 0.0147792f $X=5.22 $Y=1.885 $X2=0 $Y2=0
cc_313 N_A1_c_364_n N_A_27_392#_c_430_n 0.0178766f $X=5.67 $Y=1.885 $X2=0 $Y2=0
cc_314 A1 N_A_27_392#_c_430_n 0.0245521f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_315 N_A1_c_362_n N_A_27_392#_c_430_n 0.00370716f $X=5.635 $Y=1.667 $X2=0
+ $Y2=0
cc_316 A1 N_A_27_392#_c_433_n 0.00466348f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_317 N_A1_c_362_n N_A_27_392#_c_433_n 0.00428371f $X=5.635 $Y=1.667 $X2=0
+ $Y2=0
cc_318 N_A1_M1022_g N_A_27_392#_c_416_n 0.00252208f $X=5.635 $Y=0.74 $X2=0 $Y2=0
cc_319 A1 N_A_27_392#_c_416_n 0.0121153f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_320 N_A1_c_362_n N_A_27_392#_c_416_n 0.0022552f $X=5.635 $Y=1.667 $X2=0 $Y2=0
cc_321 N_A1_c_363_n N_VPWR_c_635_n 0.0116111f $X=5.22 $Y=1.885 $X2=0 $Y2=0
cc_322 N_A1_c_364_n N_VPWR_c_636_n 0.0093094f $X=5.67 $Y=1.885 $X2=0 $Y2=0
cc_323 N_A1_c_363_n N_VPWR_c_645_n 0.00445602f $X=5.22 $Y=1.885 $X2=0 $Y2=0
cc_324 N_A1_c_364_n N_VPWR_c_645_n 0.00445602f $X=5.67 $Y=1.885 $X2=0 $Y2=0
cc_325 N_A1_c_363_n N_VPWR_c_630_n 0.00861719f $X=5.22 $Y=1.885 $X2=0 $Y2=0
cc_326 N_A1_c_364_n N_VPWR_c_630_n 0.00858495f $X=5.67 $Y=1.885 $X2=0 $Y2=0
cc_327 N_A1_c_363_n N_A_747_392#_c_753_n 0.0137166f $X=5.22 $Y=1.885 $X2=0 $Y2=0
cc_328 N_A1_c_363_n N_A_747_392#_c_754_n 0.0114674f $X=5.22 $Y=1.885 $X2=0 $Y2=0
cc_329 N_A1_c_364_n N_A_747_392#_c_754_n 0.00775254f $X=5.67 $Y=1.885 $X2=0
+ $Y2=0
cc_330 N_A1_M1010_g N_A_477_198#_c_928_n 0.00293386f $X=5.205 $Y=0.74 $X2=0
+ $Y2=0
cc_331 N_A1_M1010_g N_A_477_198#_c_929_n 0.0177833f $X=5.205 $Y=0.74 $X2=0 $Y2=0
cc_332 N_A1_M1022_g N_A_477_198#_c_929_n 0.00415797f $X=5.635 $Y=0.74 $X2=0
+ $Y2=0
cc_333 A1 N_A_477_198#_c_929_n 0.0150501f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_334 N_A1_c_362_n N_A_477_198#_c_929_n 7.91474e-19 $X=5.635 $Y=1.667 $X2=0
+ $Y2=0
cc_335 N_A1_M1010_g N_A_477_198#_c_930_n 3.92313e-19 $X=5.205 $Y=0.74 $X2=0
+ $Y2=0
cc_336 N_A1_M1022_g N_A_477_198#_c_930_n 3.92313e-19 $X=5.635 $Y=0.74 $X2=0
+ $Y2=0
cc_337 N_A1_M1010_g N_VGND_c_991_n 0.0114363f $X=5.205 $Y=0.74 $X2=0 $Y2=0
cc_338 N_A1_M1022_g N_VGND_c_991_n 5.01478e-19 $X=5.635 $Y=0.74 $X2=0 $Y2=0
cc_339 N_A1_M1010_g N_VGND_c_992_n 5.68935e-19 $X=5.205 $Y=0.74 $X2=0 $Y2=0
cc_340 N_A1_M1022_g N_VGND_c_992_n 0.0142039f $X=5.635 $Y=0.74 $X2=0 $Y2=0
cc_341 N_A1_c_362_n N_VGND_c_992_n 0.0012667f $X=5.635 $Y=1.667 $X2=0 $Y2=0
cc_342 N_A1_M1010_g N_VGND_c_998_n 0.00383152f $X=5.205 $Y=0.74 $X2=0 $Y2=0
cc_343 N_A1_M1022_g N_VGND_c_998_n 0.00383152f $X=5.635 $Y=0.74 $X2=0 $Y2=0
cc_344 N_A1_M1010_g N_VGND_c_1005_n 0.0075754f $X=5.205 $Y=0.74 $X2=0 $Y2=0
cc_345 N_A1_M1022_g N_VGND_c_1005_n 0.0075754f $X=5.635 $Y=0.74 $X2=0 $Y2=0
cc_346 N_A_27_392#_c_424_n N_VPWR_M1004_s 9.24238e-19 $X=0.72 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_347 N_A_27_392#_c_426_n N_VPWR_M1004_s 3.60678e-19 $X=1.115 $Y=2.035
+ $X2=-0.19 $Y2=-0.245
cc_348 N_A_27_392#_c_507_p N_VPWR_M1004_s 0.00235005f $X=0.805 $Y=2.035
+ $X2=-0.19 $Y2=-0.245
cc_349 N_A_27_392#_c_427_n N_VPWR_M1006_s 0.00266f $X=2.15 $Y=2.035 $X2=0 $Y2=0
cc_350 N_A_27_392#_c_428_n N_VPWR_M1008_d 0.00209644f $X=3.22 $Y=2.035 $X2=0
+ $Y2=0
cc_351 N_A_27_392#_c_430_n N_VPWR_M1000_s 0.00452107f $X=5.975 $Y=2.035 $X2=0
+ $Y2=0
cc_352 N_A_27_392#_c_430_n N_VPWR_M1002_s 0.0076786f $X=5.975 $Y=2.035 $X2=0
+ $Y2=0
cc_353 N_A_27_392#_c_433_n N_VPWR_M1002_s 0.00132117f $X=6.06 $Y=1.95 $X2=0
+ $Y2=0
cc_354 N_A_27_392#_c_424_n N_VPWR_c_631_n 0.00606292f $X=0.72 $Y=2.035 $X2=0
+ $Y2=0
cc_355 N_A_27_392#_c_426_n N_VPWR_c_631_n 0.00239072f $X=1.115 $Y=2.035 $X2=0
+ $Y2=0
cc_356 N_A_27_392#_c_434_n N_VPWR_c_631_n 0.0197393f $X=0.28 $Y=2.115 $X2=0
+ $Y2=0
cc_357 N_A_27_392#_c_507_p N_VPWR_c_631_n 0.0138281f $X=0.805 $Y=2.035 $X2=0
+ $Y2=0
cc_358 N_A_27_392#_c_435_n N_VPWR_c_631_n 0.0197393f $X=1.28 $Y=2.115 $X2=0
+ $Y2=0
cc_359 N_A_27_392#_c_435_n N_VPWR_c_632_n 0.00877065f $X=1.28 $Y=2.115 $X2=0
+ $Y2=0
cc_360 N_A_27_392#_c_427_n N_VPWR_c_633_n 0.01825f $X=2.15 $Y=2.035 $X2=0 $Y2=0
cc_361 N_A_27_392#_c_435_n N_VPWR_c_633_n 0.0197393f $X=1.28 $Y=2.115 $X2=0
+ $Y2=0
cc_362 N_A_27_392#_c_436_n N_VPWR_c_633_n 0.0339726f $X=2.315 $Y=2.105 $X2=0
+ $Y2=0
cc_363 N_A_27_392#_c_428_n N_VPWR_c_634_n 0.0154949f $X=3.22 $Y=2.035 $X2=0
+ $Y2=0
cc_364 N_A_27_392#_c_429_n N_VPWR_c_634_n 0.0397821f $X=3.385 $Y=2.815 $X2=0
+ $Y2=0
cc_365 N_A_27_392#_c_432_n N_VPWR_c_634_n 0.0130718f $X=3.55 $Y=2.99 $X2=0 $Y2=0
cc_366 N_A_27_392#_c_436_n N_VPWR_c_634_n 0.0339726f $X=2.315 $Y=2.105 $X2=0
+ $Y2=0
cc_367 N_A_27_392#_c_438_n N_VPWR_c_635_n 0.0300015f $X=4.385 $Y=2.805 $X2=0
+ $Y2=0
cc_368 N_A_27_392#_c_418_n N_VPWR_c_636_n 0.0107376f $X=6.205 $Y=1.765 $X2=0
+ $Y2=0
cc_369 N_A_27_392#_c_419_n N_VPWR_c_636_n 4.93059e-19 $X=6.705 $Y=1.765 $X2=0
+ $Y2=0
cc_370 N_A_27_392#_c_430_n N_VPWR_c_636_n 0.0228331f $X=5.975 $Y=2.035 $X2=0
+ $Y2=0
cc_371 N_A_27_392#_c_418_n N_VPWR_c_637_n 4.83252e-19 $X=6.205 $Y=1.765 $X2=0
+ $Y2=0
cc_372 N_A_27_392#_c_419_n N_VPWR_c_637_n 0.0102165f $X=6.705 $Y=1.765 $X2=0
+ $Y2=0
cc_373 N_A_27_392#_c_420_n N_VPWR_c_637_n 0.0105015f $X=7.155 $Y=1.765 $X2=0
+ $Y2=0
cc_374 N_A_27_392#_c_423_n N_VPWR_c_637_n 5.44284e-19 $X=7.605 $Y=1.765 $X2=0
+ $Y2=0
cc_375 N_A_27_392#_c_423_n N_VPWR_c_639_n 0.0260843f $X=7.605 $Y=1.765 $X2=0
+ $Y2=0
cc_376 N_A_27_392#_c_436_n N_VPWR_c_640_n 0.00884037f $X=2.315 $Y=2.105 $X2=0
+ $Y2=0
cc_377 N_A_27_392#_c_431_n N_VPWR_c_642_n 0.0423015f $X=4.22 $Y=2.99 $X2=0 $Y2=0
cc_378 N_A_27_392#_c_432_n N_VPWR_c_642_n 0.0236566f $X=3.55 $Y=2.99 $X2=0 $Y2=0
cc_379 N_A_27_392#_c_438_n N_VPWR_c_642_n 0.0227333f $X=4.385 $Y=2.805 $X2=0
+ $Y2=0
cc_380 N_A_27_392#_c_434_n N_VPWR_c_644_n 0.00880551f $X=0.28 $Y=2.115 $X2=0
+ $Y2=0
cc_381 N_A_27_392#_c_418_n N_VPWR_c_646_n 0.00413917f $X=6.205 $Y=1.765 $X2=0
+ $Y2=0
cc_382 N_A_27_392#_c_419_n N_VPWR_c_646_n 0.00413917f $X=6.705 $Y=1.765 $X2=0
+ $Y2=0
cc_383 N_A_27_392#_c_420_n N_VPWR_c_647_n 0.00413917f $X=7.155 $Y=1.765 $X2=0
+ $Y2=0
cc_384 N_A_27_392#_c_423_n N_VPWR_c_647_n 0.00445602f $X=7.605 $Y=1.765 $X2=0
+ $Y2=0
cc_385 N_A_27_392#_c_418_n N_VPWR_c_630_n 0.00818187f $X=6.205 $Y=1.765 $X2=0
+ $Y2=0
cc_386 N_A_27_392#_c_419_n N_VPWR_c_630_n 0.00818187f $X=6.705 $Y=1.765 $X2=0
+ $Y2=0
cc_387 N_A_27_392#_c_420_n N_VPWR_c_630_n 0.00817726f $X=7.155 $Y=1.765 $X2=0
+ $Y2=0
cc_388 N_A_27_392#_c_423_n N_VPWR_c_630_n 0.00860566f $X=7.605 $Y=1.765 $X2=0
+ $Y2=0
cc_389 N_A_27_392#_c_431_n N_VPWR_c_630_n 0.0238896f $X=4.22 $Y=2.99 $X2=0 $Y2=0
cc_390 N_A_27_392#_c_432_n N_VPWR_c_630_n 0.0128296f $X=3.55 $Y=2.99 $X2=0 $Y2=0
cc_391 N_A_27_392#_c_434_n N_VPWR_c_630_n 0.0108814f $X=0.28 $Y=2.115 $X2=0
+ $Y2=0
cc_392 N_A_27_392#_c_435_n N_VPWR_c_630_n 0.0108663f $X=1.28 $Y=2.115 $X2=0
+ $Y2=0
cc_393 N_A_27_392#_c_436_n N_VPWR_c_630_n 0.0108964f $X=2.315 $Y=2.105 $X2=0
+ $Y2=0
cc_394 N_A_27_392#_c_438_n N_VPWR_c_630_n 0.0125508f $X=4.385 $Y=2.805 $X2=0
+ $Y2=0
cc_395 N_A_27_392#_c_430_n N_A_747_392#_M1015_s 0.00250873f $X=5.975 $Y=2.035
+ $X2=-0.19 $Y2=-0.245
cc_396 N_A_27_392#_c_431_n N_A_747_392#_M1015_s 0.00250873f $X=4.22 $Y=2.99
+ $X2=-0.19 $Y2=-0.245
cc_397 N_A_27_392#_c_430_n N_A_747_392#_M1000_d 0.00197722f $X=5.975 $Y=2.035
+ $X2=0 $Y2=0
cc_398 N_A_27_392#_M1016_d N_A_747_392#_c_753_n 0.00613551f $X=4.235 $Y=1.96
+ $X2=0 $Y2=0
cc_399 N_A_27_392#_c_430_n N_A_747_392#_c_753_n 0.0778199f $X=5.975 $Y=2.035
+ $X2=0 $Y2=0
cc_400 N_A_27_392#_c_431_n N_A_747_392#_c_753_n 0.00419805f $X=4.22 $Y=2.99
+ $X2=0 $Y2=0
cc_401 N_A_27_392#_c_438_n N_A_747_392#_c_753_n 0.0212524f $X=4.385 $Y=2.805
+ $X2=0 $Y2=0
cc_402 N_A_27_392#_c_430_n N_A_747_392#_c_756_n 0.0195846f $X=5.975 $Y=2.035
+ $X2=0 $Y2=0
cc_403 N_A_27_392#_c_431_n N_A_747_392#_c_756_n 0.0183575f $X=4.22 $Y=2.99 $X2=0
+ $Y2=0
cc_404 N_A_27_392#_c_430_n N_A_747_392#_c_754_n 0.0173542f $X=5.975 $Y=2.035
+ $X2=0 $Y2=0
cc_405 N_A_27_392#_M1013_g N_X_c_776_n 0.00792144f $X=6.135 $Y=0.74 $X2=0 $Y2=0
cc_406 N_A_27_392#_M1018_g N_X_c_776_n 0.00993385f $X=6.565 $Y=0.74 $X2=0 $Y2=0
cc_407 N_A_27_392#_M1021_g N_X_c_776_n 7.02145e-19 $X=7.135 $Y=0.74 $X2=0 $Y2=0
cc_408 N_A_27_392#_c_411_n N_X_c_791_n 0.00703686f $X=7.245 $Y=1.425 $X2=0 $Y2=0
cc_409 N_A_27_392#_c_568_p N_X_c_791_n 0.0209593f $X=6.96 $Y=1.515 $X2=0 $Y2=0
cc_410 N_A_27_392#_c_418_n N_X_c_785_n 0.00431856f $X=6.205 $Y=1.765 $X2=0 $Y2=0
cc_411 N_A_27_392#_c_419_n N_X_c_785_n 2.99529e-19 $X=6.705 $Y=1.765 $X2=0 $Y2=0
cc_412 N_A_27_392#_M1018_g N_X_c_777_n 0.0118691f $X=6.565 $Y=0.74 $X2=0 $Y2=0
cc_413 N_A_27_392#_M1021_g N_X_c_777_n 0.0127389f $X=7.135 $Y=0.74 $X2=0 $Y2=0
cc_414 N_A_27_392#_c_411_n N_X_c_777_n 0.00559421f $X=7.245 $Y=1.425 $X2=0 $Y2=0
cc_415 N_A_27_392#_c_568_p N_X_c_777_n 0.0451032f $X=6.96 $Y=1.515 $X2=0 $Y2=0
cc_416 N_A_27_392#_M1013_g N_X_c_778_n 0.00343246f $X=6.135 $Y=0.74 $X2=0 $Y2=0
cc_417 N_A_27_392#_M1018_g N_X_c_778_n 0.00157732f $X=6.565 $Y=0.74 $X2=0 $Y2=0
cc_418 N_A_27_392#_c_411_n N_X_c_778_n 0.00232957f $X=7.245 $Y=1.425 $X2=0 $Y2=0
cc_419 N_A_27_392#_c_568_p N_X_c_778_n 0.0276081f $X=6.96 $Y=1.515 $X2=0 $Y2=0
cc_420 N_A_27_392#_c_419_n N_X_c_803_n 0.0174967f $X=6.705 $Y=1.765 $X2=0 $Y2=0
cc_421 N_A_27_392#_c_420_n N_X_c_803_n 0.018987f $X=7.155 $Y=1.765 $X2=0 $Y2=0
cc_422 N_A_27_392#_c_411_n N_X_c_803_n 0.00631084f $X=7.245 $Y=1.425 $X2=0 $Y2=0
cc_423 N_A_27_392#_c_568_p N_X_c_803_n 0.0348131f $X=6.96 $Y=1.515 $X2=0 $Y2=0
cc_424 N_A_27_392#_M1018_g N_X_c_779_n 7.02145e-19 $X=6.565 $Y=0.74 $X2=0 $Y2=0
cc_425 N_A_27_392#_M1021_g N_X_c_779_n 0.00993385f $X=7.135 $Y=0.74 $X2=0 $Y2=0
cc_426 N_A_27_392#_M1023_g N_X_c_779_n 0.0145491f $X=7.565 $Y=0.74 $X2=0 $Y2=0
cc_427 N_A_27_392#_c_420_n N_X_c_786_n 0.00210897f $X=7.155 $Y=1.765 $X2=0 $Y2=0
cc_428 N_A_27_392#_c_411_n N_X_c_786_n 0.00248482f $X=7.245 $Y=1.425 $X2=0 $Y2=0
cc_429 N_A_27_392#_c_413_n N_X_c_786_n 0.00118727f $X=7.605 $Y=1.675 $X2=0 $Y2=0
cc_430 N_A_27_392#_c_423_n N_X_c_786_n 0.00820943f $X=7.605 $Y=1.765 $X2=0 $Y2=0
cc_431 N_A_27_392#_c_568_p N_X_c_786_n 0.00234327f $X=6.96 $Y=1.515 $X2=0 $Y2=0
cc_432 N_A_27_392#_c_420_n N_X_c_787_n 0.00606506f $X=7.155 $Y=1.765 $X2=0 $Y2=0
cc_433 N_A_27_392#_c_423_n N_X_c_787_n 0.00876549f $X=7.605 $Y=1.765 $X2=0 $Y2=0
cc_434 N_A_27_392#_M1023_g N_X_c_780_n 0.0131828f $X=7.565 $Y=0.74 $X2=0 $Y2=0
cc_435 N_A_27_392#_c_414_n N_X_c_780_n 0.00148797f $X=7.592 $Y=1.425 $X2=0 $Y2=0
cc_436 N_A_27_392#_c_413_n N_X_c_781_n 0.0116389f $X=7.605 $Y=1.675 $X2=0 $Y2=0
cc_437 N_A_27_392#_c_414_n N_X_c_781_n 0.00293976f $X=7.592 $Y=1.425 $X2=0 $Y2=0
cc_438 N_A_27_392#_c_410_n N_X_c_782_n 0.00565298f $X=7.49 $Y=1.425 $X2=0 $Y2=0
cc_439 N_A_27_392#_c_411_n N_X_c_782_n 0.00146733f $X=7.245 $Y=1.425 $X2=0 $Y2=0
cc_440 N_A_27_392#_c_413_n N_X_c_782_n 0.00172267f $X=7.605 $Y=1.675 $X2=0 $Y2=0
cc_441 N_A_27_392#_c_414_n N_X_c_782_n 0.0010485f $X=7.592 $Y=1.425 $X2=0 $Y2=0
cc_442 N_A_27_392#_c_568_p N_X_c_782_n 0.0150643f $X=6.96 $Y=1.515 $X2=0 $Y2=0
cc_443 N_A_27_392#_M1021_g N_X_c_783_n 0.00192507f $X=7.135 $Y=0.74 $X2=0 $Y2=0
cc_444 N_A_27_392#_c_410_n N_X_c_783_n 0.00245515f $X=7.49 $Y=1.425 $X2=0 $Y2=0
cc_445 N_A_27_392#_M1023_g N_X_c_783_n 0.00164391f $X=7.565 $Y=0.74 $X2=0 $Y2=0
cc_446 N_A_27_392#_c_423_n N_X_c_829_n 0.00330225f $X=7.605 $Y=1.765 $X2=0 $Y2=0
cc_447 N_A_27_392#_M1023_g X 0.00602992f $X=7.565 $Y=0.74 $X2=0 $Y2=0
cc_448 N_A_27_392#_c_414_n X 0.0059128f $X=7.592 $Y=1.425 $X2=0 $Y2=0
cc_449 N_A_27_392#_c_417_n N_A_27_74#_c_859_n 0.0131655f $X=0.715 $Y=0.95 $X2=0
+ $Y2=0
cc_450 N_A_27_392#_M1019_d N_A_27_74#_c_860_n 0.00180346f $X=0.575 $Y=0.37 $X2=0
+ $Y2=0
cc_451 N_A_27_392#_c_417_n N_A_27_74#_c_860_n 0.0176997f $X=0.715 $Y=0.95 $X2=0
+ $Y2=0
cc_452 N_A_27_392#_c_417_n N_A_27_74#_c_861_n 0.0142848f $X=0.715 $Y=0.95 $X2=0
+ $Y2=0
cc_453 N_A_27_392#_c_428_n N_A_477_198#_c_926_n 0.00825032f $X=3.22 $Y=2.035
+ $X2=0 $Y2=0
cc_454 N_A_27_392#_c_436_n N_A_477_198#_c_926_n 0.00394735f $X=2.315 $Y=2.105
+ $X2=0 $Y2=0
cc_455 N_A_27_392#_c_428_n N_A_477_198#_c_936_n 0.00478817f $X=3.22 $Y=2.035
+ $X2=0 $Y2=0
cc_456 N_A_27_392#_c_430_n N_A_477_198#_c_929_n 0.00395758f $X=5.975 $Y=2.035
+ $X2=0 $Y2=0
cc_457 N_A_27_392#_c_437_n N_A_477_198#_c_932_n 0.00481287f $X=3.385 $Y=2.115
+ $X2=0 $Y2=0
cc_458 N_A_27_392#_M1013_g N_VGND_c_992_n 0.00590268f $X=6.135 $Y=0.74 $X2=0
+ $Y2=0
cc_459 N_A_27_392#_c_416_n N_VGND_c_992_n 0.00304495f $X=6.145 $Y=1.515 $X2=0
+ $Y2=0
cc_460 N_A_27_392#_M1018_g N_VGND_c_993_n 0.00469226f $X=6.565 $Y=0.74 $X2=0
+ $Y2=0
cc_461 N_A_27_392#_M1021_g N_VGND_c_993_n 0.00469226f $X=7.135 $Y=0.74 $X2=0
+ $Y2=0
cc_462 N_A_27_392#_M1023_g N_VGND_c_995_n 0.0123273f $X=7.565 $Y=0.74 $X2=0
+ $Y2=0
cc_463 N_A_27_392#_M1013_g N_VGND_c_1000_n 0.00434272f $X=6.135 $Y=0.74 $X2=0
+ $Y2=0
cc_464 N_A_27_392#_M1018_g N_VGND_c_1000_n 0.00434272f $X=6.565 $Y=0.74 $X2=0
+ $Y2=0
cc_465 N_A_27_392#_M1021_g N_VGND_c_1003_n 0.00434272f $X=7.135 $Y=0.74 $X2=0
+ $Y2=0
cc_466 N_A_27_392#_M1023_g N_VGND_c_1003_n 0.00434272f $X=7.565 $Y=0.74 $X2=0
+ $Y2=0
cc_467 N_A_27_392#_M1013_g N_VGND_c_1005_n 0.00820772f $X=6.135 $Y=0.74 $X2=0
+ $Y2=0
cc_468 N_A_27_392#_M1018_g N_VGND_c_1005_n 0.00821294f $X=6.565 $Y=0.74 $X2=0
+ $Y2=0
cc_469 N_A_27_392#_M1021_g N_VGND_c_1005_n 0.00821294f $X=7.135 $Y=0.74 $X2=0
+ $Y2=0
cc_470 N_A_27_392#_M1023_g N_VGND_c_1005_n 0.00824014f $X=7.565 $Y=0.74 $X2=0
+ $Y2=0
cc_471 N_VPWR_M1000_s N_A_747_392#_c_753_n 0.00766476f $X=4.8 $Y=1.96 $X2=0
+ $Y2=0
cc_472 N_VPWR_c_635_n N_A_747_392#_c_753_n 0.025036f $X=4.945 $Y=2.805 $X2=0
+ $Y2=0
cc_473 N_VPWR_c_635_n N_A_747_392#_c_754_n 0.0139233f $X=4.945 $Y=2.805 $X2=0
+ $Y2=0
cc_474 N_VPWR_c_636_n N_A_747_392#_c_754_n 0.047064f $X=5.98 $Y=2.455 $X2=0
+ $Y2=0
cc_475 N_VPWR_c_645_n N_A_747_392#_c_754_n 0.0145674f $X=5.815 $Y=3.33 $X2=0
+ $Y2=0
cc_476 N_VPWR_c_630_n N_A_747_392#_c_754_n 0.0119851f $X=7.92 $Y=3.33 $X2=0
+ $Y2=0
cc_477 N_VPWR_c_636_n N_X_c_785_n 0.0266594f $X=5.98 $Y=2.455 $X2=0 $Y2=0
cc_478 N_VPWR_c_637_n N_X_c_785_n 0.023849f $X=6.93 $Y=2.435 $X2=0 $Y2=0
cc_479 N_VPWR_c_646_n N_X_c_785_n 0.0121815f $X=6.765 $Y=3.33 $X2=0 $Y2=0
cc_480 N_VPWR_c_630_n N_X_c_785_n 0.0100828f $X=7.92 $Y=3.33 $X2=0 $Y2=0
cc_481 N_VPWR_M1003_s N_X_c_803_n 0.00360677f $X=6.78 $Y=1.84 $X2=0 $Y2=0
cc_482 N_VPWR_c_637_n N_X_c_803_n 0.0179913f $X=6.93 $Y=2.435 $X2=0 $Y2=0
cc_483 N_VPWR_c_639_n N_X_c_786_n 0.00183331f $X=7.88 $Y=1.985 $X2=0 $Y2=0
cc_484 N_VPWR_c_637_n N_X_c_787_n 0.0422717f $X=6.93 $Y=2.435 $X2=0 $Y2=0
cc_485 N_VPWR_c_639_n N_X_c_787_n 0.0295221f $X=7.88 $Y=1.985 $X2=0 $Y2=0
cc_486 N_VPWR_c_647_n N_X_c_787_n 0.0110241f $X=7.715 $Y=3.33 $X2=0 $Y2=0
cc_487 N_VPWR_c_630_n N_X_c_787_n 0.00909194f $X=7.92 $Y=3.33 $X2=0 $Y2=0
cc_488 N_VPWR_c_639_n N_X_c_781_n 0.0289318f $X=7.88 $Y=1.985 $X2=0 $Y2=0
cc_489 N_X_c_778_n N_A_477_198#_c_929_n 0.00152173f $X=6.515 $Y=1.095 $X2=0
+ $Y2=0
cc_490 N_X_c_777_n N_VGND_M1018_s 0.00377777f $X=7.185 $Y=1.095 $X2=0 $Y2=0
cc_491 N_X_c_780_n N_VGND_M1023_s 0.0044011f $X=7.805 $Y=1.095 $X2=0 $Y2=0
cc_492 N_X_c_776_n N_VGND_c_992_n 0.0255177f $X=6.35 $Y=0.515 $X2=0 $Y2=0
cc_493 N_X_c_778_n N_VGND_c_992_n 0.00584871f $X=6.515 $Y=1.095 $X2=0 $Y2=0
cc_494 N_X_c_776_n N_VGND_c_993_n 0.0182384f $X=6.35 $Y=0.515 $X2=0 $Y2=0
cc_495 N_X_c_777_n N_VGND_c_993_n 0.0224739f $X=7.185 $Y=1.095 $X2=0 $Y2=0
cc_496 N_X_c_779_n N_VGND_c_993_n 0.0182384f $X=7.35 $Y=0.515 $X2=0 $Y2=0
cc_497 N_X_c_779_n N_VGND_c_995_n 0.0182384f $X=7.35 $Y=0.515 $X2=0 $Y2=0
cc_498 N_X_c_780_n N_VGND_c_995_n 0.0248922f $X=7.805 $Y=1.095 $X2=0 $Y2=0
cc_499 N_X_c_776_n N_VGND_c_1000_n 0.0144922f $X=6.35 $Y=0.515 $X2=0 $Y2=0
cc_500 N_X_c_779_n N_VGND_c_1003_n 0.0144922f $X=7.35 $Y=0.515 $X2=0 $Y2=0
cc_501 N_X_c_776_n N_VGND_c_1005_n 0.0118826f $X=6.35 $Y=0.515 $X2=0 $Y2=0
cc_502 N_X_c_779_n N_VGND_c_1005_n 0.0118826f $X=7.35 $Y=0.515 $X2=0 $Y2=0
cc_503 N_A_27_74#_c_864_n N_A_287_74#_M1005_d 0.00176891f $X=1.92 $Y=0.397
+ $X2=-0.19 $Y2=-0.245
cc_504 N_A_27_74#_M1017_s N_A_287_74#_c_897_n 0.00624487f $X=1.865 $Y=0.37 $X2=0
+ $Y2=0
cc_505 N_A_27_74#_c_863_n N_A_287_74#_c_897_n 0.024192f $X=2.085 $Y=0.375 $X2=0
+ $Y2=0
cc_506 N_A_27_74#_c_864_n N_A_287_74#_c_897_n 0.00497069f $X=1.92 $Y=0.397 $X2=0
+ $Y2=0
cc_507 N_A_27_74#_c_861_n N_A_287_74#_c_898_n 0.0204279f $X=1.145 $Y=0.965 $X2=0
+ $Y2=0
cc_508 N_A_27_74#_c_864_n N_A_287_74#_c_898_n 0.0158153f $X=1.92 $Y=0.397 $X2=0
+ $Y2=0
cc_509 N_A_27_74#_c_863_n N_A_287_74#_c_899_n 5.51636e-19 $X=2.085 $Y=0.375
+ $X2=0 $Y2=0
cc_510 N_A_27_74#_c_858_n N_VGND_c_996_n 0.018997f $X=0.247 $Y=0.6 $X2=0 $Y2=0
cc_511 N_A_27_74#_c_860_n N_VGND_c_996_n 0.0450241f $X=1.06 $Y=0.427 $X2=0 $Y2=0
cc_512 N_A_27_74#_c_862_n N_VGND_c_996_n 0.0121867f $X=1.145 $Y=0.515 $X2=0
+ $Y2=0
cc_513 N_A_27_74#_c_864_n N_VGND_c_996_n 0.0658946f $X=1.92 $Y=0.397 $X2=0 $Y2=0
cc_514 N_A_27_74#_M1017_s N_VGND_c_1005_n 0.00242558f $X=1.865 $Y=0.37 $X2=0
+ $Y2=0
cc_515 N_A_27_74#_c_858_n N_VGND_c_1005_n 0.0103026f $X=0.247 $Y=0.6 $X2=0 $Y2=0
cc_516 N_A_27_74#_c_860_n N_VGND_c_1005_n 0.0245954f $X=1.06 $Y=0.427 $X2=0
+ $Y2=0
cc_517 N_A_27_74#_c_862_n N_VGND_c_1005_n 0.00660921f $X=1.145 $Y=0.515 $X2=0
+ $Y2=0
cc_518 N_A_27_74#_c_864_n N_VGND_c_1005_n 0.0372424f $X=1.92 $Y=0.397 $X2=0
+ $Y2=0
cc_519 N_A_287_74#_c_897_n N_A_477_198#_M1009_s 0.00635284f $X=2.875 $Y=0.795
+ $X2=-0.19 $Y2=-0.245
cc_520 N_A_287_74#_c_897_n N_A_477_198#_c_926_n 0.0333166f $X=2.875 $Y=0.795
+ $X2=0 $Y2=0
cc_521 N_A_287_74#_c_898_n N_A_477_198#_c_926_n 0.00246079f $X=1.74 $Y=0.862
+ $X2=0 $Y2=0
cc_522 N_A_287_74#_M1009_d N_A_477_198#_c_936_n 0.00359685f $X=2.9 $Y=0.54 $X2=0
+ $Y2=0
cc_523 N_A_287_74#_c_899_n N_A_477_198#_c_936_n 0.014851f $X=3.04 $Y=0.7 $X2=0
+ $Y2=0
cc_524 N_A_287_74#_c_899_n N_A_477_198#_c_927_n 0.0130934f $X=3.04 $Y=0.7 $X2=0
+ $Y2=0
cc_525 N_A_287_74#_c_897_n N_VGND_c_996_n 0.0089723f $X=2.875 $Y=0.795 $X2=0
+ $Y2=0
cc_526 N_A_287_74#_c_899_n N_VGND_c_996_n 0.00617201f $X=3.04 $Y=0.7 $X2=0 $Y2=0
cc_527 N_A_287_74#_c_897_n N_VGND_c_1005_n 0.0178492f $X=2.875 $Y=0.795 $X2=0
+ $Y2=0
cc_528 N_A_287_74#_c_899_n N_VGND_c_1005_n 0.00794446f $X=3.04 $Y=0.7 $X2=0
+ $Y2=0
cc_529 N_A_477_198#_c_946_n N_VGND_M1014_s 0.00444479f $X=4.235 $Y=1.195
+ $X2=-0.19 $Y2=-0.245
cc_530 N_A_477_198#_c_927_n N_VGND_c_990_n 0.0157813f $X=3.47 $Y=0.685 $X2=0
+ $Y2=0
cc_531 N_A_477_198#_c_946_n N_VGND_c_990_n 0.0202152f $X=4.235 $Y=1.195 $X2=0
+ $Y2=0
cc_532 N_A_477_198#_c_928_n N_VGND_c_990_n 0.0165499f $X=4.4 $Y=0.685 $X2=0
+ $Y2=0
cc_533 N_A_477_198#_c_928_n N_VGND_c_991_n 0.0260211f $X=4.4 $Y=0.685 $X2=0
+ $Y2=0
cc_534 N_A_477_198#_c_929_n N_VGND_c_991_n 0.0243991f $X=5.335 $Y=1.195 $X2=0
+ $Y2=0
cc_535 N_A_477_198#_c_930_n N_VGND_c_991_n 0.0218329f $X=5.42 $Y=0.515 $X2=0
+ $Y2=0
cc_536 N_A_477_198#_c_929_n N_VGND_c_992_n 0.00157055f $X=5.335 $Y=1.195 $X2=0
+ $Y2=0
cc_537 N_A_477_198#_c_930_n N_VGND_c_992_n 0.027926f $X=5.42 $Y=0.515 $X2=0
+ $Y2=0
cc_538 N_A_477_198#_c_927_n N_VGND_c_996_n 0.00645818f $X=3.47 $Y=0.685 $X2=0
+ $Y2=0
cc_539 N_A_477_198#_c_930_n N_VGND_c_998_n 0.00749631f $X=5.42 $Y=0.515 $X2=0
+ $Y2=0
cc_540 N_A_477_198#_c_928_n N_VGND_c_1002_n 0.00858533f $X=4.4 $Y=0.685 $X2=0
+ $Y2=0
cc_541 N_A_477_198#_c_927_n N_VGND_c_1005_n 0.00815448f $X=3.47 $Y=0.685 $X2=0
+ $Y2=0
cc_542 N_A_477_198#_c_928_n N_VGND_c_1005_n 0.0108043f $X=4.4 $Y=0.685 $X2=0
+ $Y2=0
cc_543 N_A_477_198#_c_930_n N_VGND_c_1005_n 0.0062048f $X=5.42 $Y=0.515 $X2=0
+ $Y2=0
