* File: sky130_fd_sc_hs__a41oi_4.spice
* Created: Tue Sep  1 19:54:28 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hs__a41oi_4.pex.spice"
.subckt sky130_fd_sc_hs__a41oi_4  VNB VPB B1 A1 A2 A3 A4 Y VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* Y	Y
* A4	A4
* A3	A3
* A2	A2
* A1	A1
* B1	B1
* VPB	VPB
* VNB	VNB
MM1016 N_VGND_M1016_d N_B1_M1016_g N_Y_M1016_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.1295 PD=2.05 PS=1.09 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75000.7 A=0.111 P=1.78 MULT=1
MM1035 N_VGND_M1035_d N_B1_M1035_g N_Y_M1016_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.1295 PD=2.05 PS=1.09 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75000.7
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1027 N_Y_M1027_d N_A1_M1027_g N_A_325_74#_M1027_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1295 AS=0.2109 PD=1.09 PS=2.05 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75003.8 A=0.111 P=1.78 MULT=1
MM1029 N_Y_M1027_d N_A1_M1029_g N_A_325_74#_M1029_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1295 AS=0.2294 PD=1.09 PS=1.36 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.7
+ SB=75003.3 A=0.111 P=1.78 MULT=1
MM1032 N_Y_M1032_d N_A1_M1032_g N_A_325_74#_M1029_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.2294 PD=1.02 PS=1.36 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.5
+ SB=75002.5 A=0.111 P=1.78 MULT=1
MM1037 N_Y_M1032_d N_A1_M1037_g N_A_325_74#_M1037_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1295 PD=1.02 PS=1.09 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75001.9
+ SB=75002.1 A=0.111 P=1.78 MULT=1
MM1006 N_A_852_74#_M1006_d N_A2_M1006_g N_A_325_74#_M1037_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1295 AS=0.1295 PD=1.09 PS=1.09 NRD=11.34 NRS=0 M=1 R=4.93333
+ SA=75002.4 SB=75001.6 A=0.111 P=1.78 MULT=1
MM1007 N_A_852_74#_M1006_d N_A2_M1007_g N_A_325_74#_M1007_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1295 AS=0.1036 PD=1.09 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75002.9 SB=75001.1 A=0.111 P=1.78 MULT=1
MM1030 N_A_852_74#_M1030_d N_A2_M1030_g N_A_325_74#_M1007_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75003.3 SB=75000.6 A=0.111 P=1.78 MULT=1
MM1033 N_A_852_74#_M1030_d N_A2_M1033_g N_A_325_74#_M1033_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.2109 PD=1.02 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75003.8 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1010 N_A_1235_74#_M1010_d N_A3_M1010_g N_A_852_74#_M1010_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.2109 AS=0.1036 PD=2.05 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75003.3 A=0.111 P=1.78 MULT=1
MM1024 N_A_1235_74#_M1024_d N_A3_M1024_g N_A_852_74#_M1010_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.6 SB=75002.8 A=0.111 P=1.78 MULT=1
MM1028 N_A_1235_74#_M1024_d N_A3_M1028_g N_A_852_74#_M1028_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75001.1 SB=75002.4 A=0.111 P=1.78 MULT=1
MM1036 N_A_1235_74#_M1036_d N_A3_M1036_g N_A_852_74#_M1028_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75001.5 SB=75002 A=0.111 P=1.78 MULT=1
MM1003 N_A_1235_74#_M1036_d N_A4_M1003_g N_VGND_M1003_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.9
+ SB=75001.5 A=0.111 P=1.78 MULT=1
MM1017 N_A_1235_74#_M1017_d N_A4_M1017_g N_VGND_M1003_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75002.4
+ SB=75001.1 A=0.111 P=1.78 MULT=1
MM1022 N_A_1235_74#_M1017_d N_A4_M1022_g N_VGND_M1022_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1184 PD=1.02 PS=1.06 NRD=0 NRS=0 M=1 R=4.93333 SA=75002.8
+ SB=75000.7 A=0.111 P=1.78 MULT=1
MM1034 N_A_1235_74#_M1034_d N_A4_M1034_g N_VGND_M1022_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.1184 PD=2.05 PS=1.06 NRD=0 NRS=6.48 M=1 R=4.93333 SA=75003.3
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1014 N_Y_M1014_d N_B1_M1014_g N_A_27_368#_M1014_s VPB PSHORT L=0.15 W=1.12
+ AD=0.1932 AS=0.336 PD=1.465 PS=2.84 NRD=9.6727 NRS=2.6201 M=1 R=7.46667
+ SA=75000.2 SB=75009.3 A=0.168 P=2.54 MULT=1
MM1018 N_Y_M1014_d N_B1_M1018_g N_A_27_368#_M1018_s VPB PSHORT L=0.15 W=1.12
+ AD=0.1932 AS=0.196 PD=1.465 PS=1.47 NRD=1.7533 NRS=10.5395 M=1 R=7.46667
+ SA=75000.7 SB=75008.8 A=0.168 P=2.54 MULT=1
MM1019 N_Y_M1019_d N_B1_M1019_g N_A_27_368#_M1018_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.196 PD=1.42 PS=1.47 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.2 SB=75008.3 A=0.168 P=2.54 MULT=1
MM1023 N_Y_M1019_d N_B1_M1023_g N_A_27_368#_M1023_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.7 SB=75007.8 A=0.168 P=2.54 MULT=1
MM1012 N_A_27_368#_M1023_s N_A1_M1012_g N_VPWR_M1012_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.224 PD=1.42 PS=1.52 NRD=1.7533 NRS=10.5395 M=1 R=7.46667
+ SA=75002.1 SB=75007.4 A=0.168 P=2.54 MULT=1
MM1020 N_A_27_368#_M1020_d N_A1_M1020_g N_VPWR_M1012_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.224 PD=1.42 PS=1.52 NRD=1.7533 NRS=10.5395 M=1 R=7.46667
+ SA=75002.7 SB=75006.8 A=0.168 P=2.54 MULT=1
MM1025 N_A_27_368#_M1020_d N_A1_M1025_g N_VPWR_M1025_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.1988 PD=1.42 PS=1.475 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75003.1 SB=75006.4 A=0.168 P=2.54 MULT=1
MM1026 N_A_27_368#_M1026_d N_A1_M1026_g N_VPWR_M1025_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.1988 PD=1.42 PS=1.475 NRD=1.7533 NRS=11.426 M=1 R=7.46667
+ SA=75003.6 SB=75005.9 A=0.168 P=2.54 MULT=1
MM1000 N_VPWR_M1000_d N_A2_M1000_g N_A_27_368#_M1026_d VPB PSHORT L=0.15 W=1.12
+ AD=0.2016 AS=0.168 PD=1.48 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75004.1 SB=75005.4 A=0.168 P=2.54 MULT=1
MM1001 N_VPWR_M1000_d N_A2_M1001_g N_A_27_368#_M1001_s VPB PSHORT L=0.15 W=1.12
+ AD=0.2016 AS=0.168 PD=1.48 PS=1.42 NRD=12.2928 NRS=1.7533 M=1 R=7.46667
+ SA=75004.6 SB=75004.9 A=0.168 P=2.54 MULT=1
MM1015 N_VPWR_M1015_d N_A2_M1015_g N_A_27_368#_M1001_s VPB PSHORT L=0.15 W=1.12
+ AD=0.196 AS=0.168 PD=1.47 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667 SA=75005
+ SB=75004.5 A=0.168 P=2.54 MULT=1
MM1031 N_VPWR_M1015_d N_A2_M1031_g N_A_27_368#_M1031_s VPB PSHORT L=0.15 W=1.12
+ AD=0.196 AS=0.168 PD=1.47 PS=1.42 NRD=10.5395 NRS=1.7533 M=1 R=7.46667
+ SA=75005.5 SB=75004 A=0.168 P=2.54 MULT=1
MM1002 N_A_27_368#_M1031_s N_A3_M1002_g N_VPWR_M1002_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.196 PD=1.42 PS=1.47 NRD=1.7533 NRS=1.7533 M=1 R=7.46667 SA=75006
+ SB=75003.5 A=0.168 P=2.54 MULT=1
MM1004 N_A_27_368#_M1004_d N_A3_M1004_g N_VPWR_M1002_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.196 PD=1.42 PS=1.47 NRD=1.7533 NRS=10.5395 M=1 R=7.46667
+ SA=75006.5 SB=75003 A=0.168 P=2.54 MULT=1
MM1008 N_A_27_368#_M1004_d N_A3_M1008_g N_VPWR_M1008_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.196 PD=1.42 PS=1.47 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75006.9 SB=75002.6 A=0.168 P=2.54 MULT=1
MM1009 N_A_27_368#_M1009_d N_A3_M1009_g N_VPWR_M1008_s VPB PSHORT L=0.15 W=1.12
+ AD=0.196 AS=0.196 PD=1.47 PS=1.47 NRD=1.7533 NRS=10.5395 M=1 R=7.46667
+ SA=75007.4 SB=75002.1 A=0.168 P=2.54 MULT=1
MM1005 N_VPWR_M1005_d N_A4_M1005_g N_A_27_368#_M1009_d VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.196 PD=1.42 PS=1.47 NRD=1.7533 NRS=10.5395 M=1 R=7.46667
+ SA=75007.9 SB=75001.6 A=0.168 P=2.54 MULT=1
MM1011 N_VPWR_M1005_d N_A4_M1011_g N_A_27_368#_M1011_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75008.4 SB=75001.1 A=0.168 P=2.54 MULT=1
MM1013 N_VPWR_M1013_d N_A4_M1013_g N_A_27_368#_M1011_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75008.8 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1021 N_VPWR_M1013_d N_A4_M1021_g N_A_27_368#_M1021_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.3304 PD=1.42 PS=2.83 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75009.3 SB=75000.2 A=0.168 P=2.54 MULT=1
DX38_noxref VNB VPB NWDIODE A=19.4556 P=24.64
c_72 VNB 0 1.1015e-19 $X=0 $Y=0
*
.include "sky130_fd_sc_hs__a41oi_4.pxi.spice"
*
.ends
*
*
