* File: sky130_fd_sc_hs__a31o_2.pxi.spice
* Created: Tue Sep  1 19:52:56 2020
* 
x_PM_SKY130_FD_SC_HS__A31O_2%A_97_296# N_A_97_296#_M1007_d N_A_97_296#_M1001_d
+ N_A_97_296#_M1005_g N_A_97_296#_c_62_n N_A_97_296#_M1008_g N_A_97_296#_M1006_g
+ N_A_97_296#_c_63_n N_A_97_296#_M1009_g N_A_97_296#_c_58_n N_A_97_296#_c_71_p
+ N_A_97_296#_c_140_p N_A_97_296#_c_64_n N_A_97_296#_c_91_p N_A_97_296#_c_59_n
+ N_A_97_296#_c_65_n N_A_97_296#_c_60_n N_A_97_296#_c_61_n
+ PM_SKY130_FD_SC_HS__A31O_2%A_97_296#
x_PM_SKY130_FD_SC_HS__A31O_2%A3 N_A3_c_158_n N_A3_M1010_g N_A3_c_159_n
+ N_A3_M1002_g A3 PM_SKY130_FD_SC_HS__A31O_2%A3
x_PM_SKY130_FD_SC_HS__A31O_2%A2 N_A2_c_189_n N_A2_M1004_g N_A2_c_190_n
+ N_A2_M1011_g A2 N_A2_c_191_n PM_SKY130_FD_SC_HS__A31O_2%A2
x_PM_SKY130_FD_SC_HS__A31O_2%A1 N_A1_c_217_n N_A1_M1007_g N_A1_c_218_n
+ N_A1_M1003_g A1 PM_SKY130_FD_SC_HS__A31O_2%A1
x_PM_SKY130_FD_SC_HS__A31O_2%B1 N_B1_c_248_n N_B1_M1000_g N_B1_c_249_n
+ N_B1_M1001_g B1 PM_SKY130_FD_SC_HS__A31O_2%B1
x_PM_SKY130_FD_SC_HS__A31O_2%VPWR N_VPWR_M1008_s N_VPWR_M1009_s N_VPWR_M1011_d
+ N_VPWR_c_270_n N_VPWR_c_271_n N_VPWR_c_272_n N_VPWR_c_273_n VPWR
+ N_VPWR_c_274_n N_VPWR_c_275_n N_VPWR_c_276_n N_VPWR_c_269_n N_VPWR_c_278_n
+ N_VPWR_c_279_n PM_SKY130_FD_SC_HS__A31O_2%VPWR
x_PM_SKY130_FD_SC_HS__A31O_2%X N_X_M1005_s N_X_M1008_d N_X_c_319_n N_X_c_320_n X
+ X X X N_X_c_321_n PM_SKY130_FD_SC_HS__A31O_2%X
x_PM_SKY130_FD_SC_HS__A31O_2%A_362_368# N_A_362_368#_M1010_d
+ N_A_362_368#_M1003_d N_A_362_368#_c_353_n N_A_362_368#_c_349_n
+ N_A_362_368#_c_350_n PM_SKY130_FD_SC_HS__A31O_2%A_362_368#
x_PM_SKY130_FD_SC_HS__A31O_2%VGND N_VGND_M1005_d N_VGND_M1006_d N_VGND_M1000_d
+ N_VGND_c_375_n N_VGND_c_376_n N_VGND_c_377_n N_VGND_c_378_n VGND
+ N_VGND_c_379_n N_VGND_c_380_n N_VGND_c_381_n N_VGND_c_382_n
+ PM_SKY130_FD_SC_HS__A31O_2%VGND
cc_1 VNB N_A_97_296#_M1005_g 0.0260123f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=0.74
cc_2 VNB N_A_97_296#_M1006_g 0.0235682f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=0.74
cc_3 VNB N_A_97_296#_c_58_n 0.00317249f $X=-0.19 $Y=-0.245 $X2=1.22 $Y2=1.3
cc_4 VNB N_A_97_296#_c_59_n 0.00335352f $X=-0.19 $Y=-0.245 $X2=3.015 $Y2=0.495
cc_5 VNB N_A_97_296#_c_60_n 0.00590395f $X=-0.19 $Y=-0.245 $X2=1.12 $Y2=1.465
cc_6 VNB N_A_97_296#_c_61_n 0.0762146f $X=-0.19 $Y=-0.245 $X2=1.025 $Y2=1.532
cc_7 VNB N_A3_c_158_n 0.0399734f $X=-0.19 $Y=-0.245 $X2=2.815 $Y2=0.37
cc_8 VNB N_A3_c_159_n 0.0188039f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB A3 0.00334701f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=1.3
cc_10 VNB N_A2_c_189_n 0.0183498f $X=-0.19 $Y=-0.245 $X2=2.815 $Y2=0.37
cc_11 VNB N_A2_c_190_n 0.0349366f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A2_c_191_n 0.00752993f $X=-0.19 $Y=-0.245 $X2=0.575 $Y2=1.765
cc_13 VNB N_A1_c_217_n 0.0198831f $X=-0.19 $Y=-0.245 $X2=2.815 $Y2=0.37
cc_14 VNB N_A1_c_218_n 0.0352811f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB A1 0.0109964f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=1.3
cc_16 VNB N_B1_c_248_n 0.0220404f $X=-0.19 $Y=-0.245 $X2=2.815 $Y2=0.37
cc_17 VNB N_B1_c_249_n 0.0676131f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB B1 0.00926001f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=1.3
cc_19 VNB N_VPWR_c_269_n 0.163682f $X=-0.19 $Y=-0.245 $X2=3.015 $Y2=0.925
cc_20 VNB N_X_c_319_n 0.00229096f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=0.74
cc_21 VNB N_X_c_320_n 0.00306343f $X=-0.19 $Y=-0.245 $X2=0.575 $Y2=2.4
cc_22 VNB N_X_c_321_n 0.00113823f $X=-0.19 $Y=-0.245 $X2=3.555 $Y2=1.985
cc_23 VNB N_VGND_c_375_n 0.0122168f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_VGND_c_376_n 0.0550278f $X=-0.19 $Y=-0.245 $X2=0.575 $Y2=2.4
cc_25 VNB N_VGND_c_377_n 0.0131437f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=1.3
cc_26 VNB N_VGND_c_378_n 0.0344105f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=0.74
cc_27 VNB N_VGND_c_379_n 0.0172472f $X=-0.19 $Y=-0.245 $X2=1.025 $Y2=2.4
cc_28 VNB N_VGND_c_380_n 0.0489588f $X=-0.19 $Y=-0.245 $X2=3.385 $Y2=1.805
cc_29 VNB N_VGND_c_381_n 0.0187802f $X=-0.19 $Y=-0.245 $X2=3.555 $Y2=2.695
cc_30 VNB N_VGND_c_382_n 0.228974f $X=-0.19 $Y=-0.245 $X2=0.575 $Y2=1.532
cc_31 VPB N_A_97_296#_c_62_n 0.0173551f $X=-0.19 $Y=1.66 $X2=0.575 $Y2=1.765
cc_32 VPB N_A_97_296#_c_63_n 0.017491f $X=-0.19 $Y=1.66 $X2=1.025 $Y2=1.765
cc_33 VPB N_A_97_296#_c_64_n 0.0376948f $X=-0.19 $Y=1.66 $X2=3.385 $Y2=1.805
cc_34 VPB N_A_97_296#_c_65_n 0.0404069f $X=-0.19 $Y=1.66 $X2=3.555 $Y2=1.985
cc_35 VPB N_A_97_296#_c_60_n 0.00232882f $X=-0.19 $Y=1.66 $X2=1.12 $Y2=1.465
cc_36 VPB N_A_97_296#_c_61_n 0.0173848f $X=-0.19 $Y=1.66 $X2=1.025 $Y2=1.532
cc_37 VPB N_A3_c_158_n 0.0230895f $X=-0.19 $Y=1.66 $X2=2.815 $Y2=0.37
cc_38 VPB N_A2_c_190_n 0.022641f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_39 VPB N_A1_c_218_n 0.0232123f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_40 VPB N_B1_c_249_n 0.0281798f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_41 VPB N_VPWR_c_270_n 0.012885f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_42 VPB N_VPWR_c_271_n 0.0638092f $X=-0.19 $Y=1.66 $X2=0.575 $Y2=2.4
cc_43 VPB N_VPWR_c_272_n 0.0131994f $X=-0.19 $Y=1.66 $X2=1.025 $Y2=1.765
cc_44 VPB N_VPWR_c_273_n 0.0200045f $X=-0.19 $Y=1.66 $X2=1.305 $Y2=0.925
cc_45 VPB N_VPWR_c_274_n 0.0181766f $X=-0.19 $Y=1.66 $X2=3.015 $Y2=0.495
cc_46 VPB N_VPWR_c_275_n 0.0209833f $X=-0.19 $Y=1.66 $X2=3.555 $Y2=1.985
cc_47 VPB N_VPWR_c_276_n 0.034947f $X=-0.19 $Y=1.66 $X2=1.305 $Y2=1.805
cc_48 VPB N_VPWR_c_269_n 0.082478f $X=-0.19 $Y=1.66 $X2=3.015 $Y2=0.925
cc_49 VPB N_VPWR_c_278_n 0.010089f $X=-0.19 $Y=1.66 $X2=1.12 $Y2=1.532
cc_50 VPB N_VPWR_c_279_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_51 VPB X 0.00171795f $X=-0.19 $Y=1.66 $X2=0.995 $Y2=1.3
cc_52 VPB X 0.00247758f $X=-0.19 $Y=1.66 $X2=1.305 $Y2=0.925
cc_53 VPB N_X_c_321_n 8.38373e-19 $X=-0.19 $Y=1.66 $X2=3.555 $Y2=1.985
cc_54 VPB N_A_362_368#_c_349_n 0.003137f $X=-0.19 $Y=1.66 $X2=0.995 $Y2=1.3
cc_55 VPB N_A_362_368#_c_350_n 0.00348704f $X=-0.19 $Y=1.66 $X2=0.995 $Y2=0.74
cc_56 N_A_97_296#_M1006_g N_A3_c_158_n 0.00147268f $X=0.995 $Y=0.74 $X2=-0.19
+ $Y2=-0.245
cc_57 N_A_97_296#_c_63_n N_A3_c_158_n 0.0102934f $X=1.025 $Y=1.765 $X2=-0.19
+ $Y2=-0.245
cc_58 N_A_97_296#_c_58_n N_A3_c_158_n 6.42308e-19 $X=1.22 $Y=1.3 $X2=-0.19
+ $Y2=-0.245
cc_59 N_A_97_296#_c_71_p N_A3_c_158_n 0.00100895f $X=2.85 $Y=0.925 $X2=-0.19
+ $Y2=-0.245
cc_60 N_A_97_296#_c_64_n N_A3_c_158_n 0.0176628f $X=3.385 $Y=1.805 $X2=-0.19
+ $Y2=-0.245
cc_61 N_A_97_296#_c_60_n N_A3_c_158_n 0.00486307f $X=1.12 $Y=1.465 $X2=-0.19
+ $Y2=-0.245
cc_62 N_A_97_296#_c_61_n N_A3_c_158_n 0.0177963f $X=1.025 $Y=1.532 $X2=-0.19
+ $Y2=-0.245
cc_63 N_A_97_296#_M1006_g N_A3_c_159_n 0.00877705f $X=0.995 $Y=0.74 $X2=0 $Y2=0
cc_64 N_A_97_296#_c_58_n N_A3_c_159_n 0.00315986f $X=1.22 $Y=1.3 $X2=0 $Y2=0
cc_65 N_A_97_296#_c_71_p N_A3_c_159_n 0.0126481f $X=2.85 $Y=0.925 $X2=0 $Y2=0
cc_66 N_A_97_296#_c_58_n A3 0.00757247f $X=1.22 $Y=1.3 $X2=0 $Y2=0
cc_67 N_A_97_296#_c_71_p A3 0.0228656f $X=2.85 $Y=0.925 $X2=0 $Y2=0
cc_68 N_A_97_296#_c_64_n A3 0.024317f $X=3.385 $Y=1.805 $X2=0 $Y2=0
cc_69 N_A_97_296#_c_60_n A3 0.0164597f $X=1.12 $Y=1.465 $X2=0 $Y2=0
cc_70 N_A_97_296#_c_61_n A3 3.04404e-19 $X=1.025 $Y=1.532 $X2=0 $Y2=0
cc_71 N_A_97_296#_c_71_p N_A2_c_189_n 0.0122562f $X=2.85 $Y=0.925 $X2=-0.19
+ $Y2=-0.245
cc_72 N_A_97_296#_c_71_p N_A2_c_190_n 0.0010191f $X=2.85 $Y=0.925 $X2=0 $Y2=0
cc_73 N_A_97_296#_c_64_n N_A2_c_190_n 0.0157598f $X=3.385 $Y=1.805 $X2=0 $Y2=0
cc_74 N_A_97_296#_c_71_p N_A2_c_191_n 0.0250213f $X=2.85 $Y=0.925 $X2=0 $Y2=0
cc_75 N_A_97_296#_c_64_n N_A2_c_191_n 0.0283471f $X=3.385 $Y=1.805 $X2=0 $Y2=0
cc_76 N_A_97_296#_c_71_p N_A1_c_217_n 0.012933f $X=2.85 $Y=0.925 $X2=-0.19
+ $Y2=-0.245
cc_77 N_A_97_296#_c_59_n N_A1_c_217_n 0.00348158f $X=3.015 $Y=0.495 $X2=-0.19
+ $Y2=-0.245
cc_78 N_A_97_296#_c_64_n N_A1_c_218_n 0.0163035f $X=3.385 $Y=1.805 $X2=0 $Y2=0
cc_79 N_A_97_296#_c_91_p N_A1_c_218_n 9.58112e-19 $X=3.015 $Y=0.84 $X2=0 $Y2=0
cc_80 N_A_97_296#_c_65_n N_A1_c_218_n 8.4488e-19 $X=3.555 $Y=1.985 $X2=0 $Y2=0
cc_81 N_A_97_296#_c_71_p A1 0.012294f $X=2.85 $Y=0.925 $X2=0 $Y2=0
cc_82 N_A_97_296#_c_64_n A1 0.0435494f $X=3.385 $Y=1.805 $X2=0 $Y2=0
cc_83 N_A_97_296#_c_91_p A1 0.0277108f $X=3.015 $Y=0.84 $X2=0 $Y2=0
cc_84 N_A_97_296#_c_59_n N_B1_c_248_n 0.00298143f $X=3.015 $Y=0.495 $X2=-0.19
+ $Y2=-0.245
cc_85 N_A_97_296#_c_64_n N_B1_c_249_n 0.0239144f $X=3.385 $Y=1.805 $X2=0 $Y2=0
cc_86 N_A_97_296#_c_65_n N_B1_c_249_n 0.011338f $X=3.555 $Y=1.985 $X2=0 $Y2=0
cc_87 N_A_97_296#_c_64_n B1 0.0272055f $X=3.385 $Y=1.805 $X2=0 $Y2=0
cc_88 N_A_97_296#_c_64_n N_VPWR_M1009_s 0.0035884f $X=3.385 $Y=1.805 $X2=0 $Y2=0
cc_89 N_A_97_296#_c_60_n N_VPWR_M1009_s 0.00197987f $X=1.12 $Y=1.465 $X2=0 $Y2=0
cc_90 N_A_97_296#_c_64_n N_VPWR_M1011_d 0.00427791f $X=3.385 $Y=1.805 $X2=0
+ $Y2=0
cc_91 N_A_97_296#_c_62_n N_VPWR_c_271_n 0.00823862f $X=0.575 $Y=1.765 $X2=0
+ $Y2=0
cc_92 N_A_97_296#_c_62_n N_VPWR_c_272_n 5.98333e-19 $X=0.575 $Y=1.765 $X2=0
+ $Y2=0
cc_93 N_A_97_296#_c_63_n N_VPWR_c_272_n 0.0190899f $X=1.025 $Y=1.765 $X2=0 $Y2=0
cc_94 N_A_97_296#_c_64_n N_VPWR_c_272_n 0.0242084f $X=3.385 $Y=1.805 $X2=0 $Y2=0
cc_95 N_A_97_296#_c_60_n N_VPWR_c_272_n 0.0142866f $X=1.12 $Y=1.465 $X2=0 $Y2=0
cc_96 N_A_97_296#_c_61_n N_VPWR_c_272_n 6.27077e-19 $X=1.025 $Y=1.532 $X2=0
+ $Y2=0
cc_97 N_A_97_296#_c_62_n N_VPWR_c_274_n 0.00411612f $X=0.575 $Y=1.765 $X2=0
+ $Y2=0
cc_98 N_A_97_296#_c_63_n N_VPWR_c_274_n 0.00429299f $X=1.025 $Y=1.765 $X2=0
+ $Y2=0
cc_99 N_A_97_296#_c_65_n N_VPWR_c_276_n 0.010098f $X=3.555 $Y=1.985 $X2=0 $Y2=0
cc_100 N_A_97_296#_c_62_n N_VPWR_c_269_n 0.00751233f $X=0.575 $Y=1.765 $X2=0
+ $Y2=0
cc_101 N_A_97_296#_c_63_n N_VPWR_c_269_n 0.00847721f $X=1.025 $Y=1.765 $X2=0
+ $Y2=0
cc_102 N_A_97_296#_c_65_n N_VPWR_c_269_n 0.0115323f $X=3.555 $Y=1.985 $X2=0
+ $Y2=0
cc_103 N_A_97_296#_M1005_g N_X_c_319_n 0.0078359f $X=0.565 $Y=0.74 $X2=0 $Y2=0
cc_104 N_A_97_296#_M1006_g N_X_c_319_n 5.92016e-19 $X=0.995 $Y=0.74 $X2=0 $Y2=0
cc_105 N_A_97_296#_M1005_g N_X_c_320_n 0.00164237f $X=0.565 $Y=0.74 $X2=0 $Y2=0
cc_106 N_A_97_296#_c_58_n N_X_c_320_n 0.00392342f $X=1.22 $Y=1.3 $X2=0 $Y2=0
cc_107 N_A_97_296#_c_61_n N_X_c_320_n 0.00199986f $X=1.025 $Y=1.532 $X2=0 $Y2=0
cc_108 N_A_97_296#_c_62_n X 0.00255173f $X=0.575 $Y=1.765 $X2=0 $Y2=0
cc_109 N_A_97_296#_c_63_n X 5.67061e-19 $X=1.025 $Y=1.765 $X2=0 $Y2=0
cc_110 N_A_97_296#_c_60_n X 0.00141815f $X=1.12 $Y=1.465 $X2=0 $Y2=0
cc_111 N_A_97_296#_c_61_n X 0.00617155f $X=1.025 $Y=1.532 $X2=0 $Y2=0
cc_112 N_A_97_296#_c_62_n X 0.0131908f $X=0.575 $Y=1.765 $X2=0 $Y2=0
cc_113 N_A_97_296#_M1005_g N_X_c_321_n 0.00856132f $X=0.565 $Y=0.74 $X2=0 $Y2=0
cc_114 N_A_97_296#_c_62_n N_X_c_321_n 0.00297978f $X=0.575 $Y=1.765 $X2=0 $Y2=0
cc_115 N_A_97_296#_M1006_g N_X_c_321_n 9.64425e-19 $X=0.995 $Y=0.74 $X2=0 $Y2=0
cc_116 N_A_97_296#_c_58_n N_X_c_321_n 0.00544148f $X=1.22 $Y=1.3 $X2=0 $Y2=0
cc_117 N_A_97_296#_c_60_n N_X_c_321_n 0.0304594f $X=1.12 $Y=1.465 $X2=0 $Y2=0
cc_118 N_A_97_296#_c_61_n N_X_c_321_n 0.0346741f $X=1.025 $Y=1.532 $X2=0 $Y2=0
cc_119 N_A_97_296#_c_64_n N_A_362_368#_M1010_d 0.00197722f $X=3.385 $Y=1.805
+ $X2=-0.19 $Y2=-0.245
cc_120 N_A_97_296#_c_64_n N_A_362_368#_M1003_d 0.00250873f $X=3.385 $Y=1.805
+ $X2=0 $Y2=0
cc_121 N_A_97_296#_c_64_n N_A_362_368#_c_353_n 0.045543f $X=3.385 $Y=1.805 $X2=0
+ $Y2=0
cc_122 N_A_97_296#_c_63_n N_A_362_368#_c_349_n 2.1805e-19 $X=1.025 $Y=1.765
+ $X2=0 $Y2=0
cc_123 N_A_97_296#_c_64_n N_A_362_368#_c_349_n 0.0173337f $X=3.385 $Y=1.805
+ $X2=0 $Y2=0
cc_124 N_A_97_296#_c_64_n N_A_362_368#_c_350_n 0.0203011f $X=3.385 $Y=1.805
+ $X2=0 $Y2=0
cc_125 N_A_97_296#_c_65_n N_A_362_368#_c_350_n 0.0245379f $X=3.555 $Y=1.985
+ $X2=0 $Y2=0
cc_126 N_A_97_296#_c_58_n N_VGND_M1006_d 0.00324595f $X=1.22 $Y=1.3 $X2=0 $Y2=0
cc_127 N_A_97_296#_c_71_p N_VGND_M1006_d 0.0156289f $X=2.85 $Y=0.925 $X2=0 $Y2=0
cc_128 N_A_97_296#_c_140_p N_VGND_M1006_d 0.00542593f $X=1.305 $Y=0.925 $X2=0
+ $Y2=0
cc_129 N_A_97_296#_M1005_g N_VGND_c_376_n 0.0184209f $X=0.565 $Y=0.74 $X2=0
+ $Y2=0
cc_130 N_A_97_296#_c_59_n N_VGND_c_378_n 0.0183215f $X=3.015 $Y=0.495 $X2=0
+ $Y2=0
cc_131 N_A_97_296#_M1005_g N_VGND_c_379_n 0.00434272f $X=0.565 $Y=0.74 $X2=0
+ $Y2=0
cc_132 N_A_97_296#_M1006_g N_VGND_c_379_n 0.004307f $X=0.995 $Y=0.74 $X2=0 $Y2=0
cc_133 N_A_97_296#_c_59_n N_VGND_c_380_n 0.0146038f $X=3.015 $Y=0.495 $X2=0
+ $Y2=0
cc_134 N_A_97_296#_M1005_g N_VGND_c_381_n 4.01823e-19 $X=0.565 $Y=0.74 $X2=0
+ $Y2=0
cc_135 N_A_97_296#_M1006_g N_VGND_c_381_n 0.00736755f $X=0.995 $Y=0.74 $X2=0
+ $Y2=0
cc_136 N_A_97_296#_c_71_p N_VGND_c_381_n 0.021742f $X=2.85 $Y=0.925 $X2=0 $Y2=0
cc_137 N_A_97_296#_c_140_p N_VGND_c_381_n 0.0111679f $X=1.305 $Y=0.925 $X2=0
+ $Y2=0
cc_138 N_A_97_296#_c_61_n N_VGND_c_381_n 7.08877e-19 $X=1.025 $Y=1.532 $X2=0
+ $Y2=0
cc_139 N_A_97_296#_M1005_g N_VGND_c_382_n 0.00823934f $X=0.565 $Y=0.74 $X2=0
+ $Y2=0
cc_140 N_A_97_296#_M1006_g N_VGND_c_382_n 0.00847524f $X=0.995 $Y=0.74 $X2=0
+ $Y2=0
cc_141 N_A_97_296#_c_71_p N_VGND_c_382_n 0.0372445f $X=2.85 $Y=0.925 $X2=0 $Y2=0
cc_142 N_A_97_296#_c_140_p N_VGND_c_382_n 7.38843e-19 $X=1.305 $Y=0.925 $X2=0
+ $Y2=0
cc_143 N_A_97_296#_c_59_n N_VGND_c_382_n 0.0121018f $X=3.015 $Y=0.495 $X2=0
+ $Y2=0
cc_144 N_A_97_296#_c_71_p A_371_74# 0.00734082f $X=2.85 $Y=0.925 $X2=-0.19
+ $Y2=-0.245
cc_145 N_A_97_296#_c_71_p A_449_74# 0.0147367f $X=2.85 $Y=0.925 $X2=-0.19
+ $Y2=-0.245
cc_146 N_A3_c_159_n N_A2_c_189_n 0.0359536f $X=1.78 $Y=1.22 $X2=-0.19 $Y2=-0.245
cc_147 A3 N_A2_c_189_n 4.24429e-19 $X=1.595 $Y=1.21 $X2=-0.19 $Y2=-0.245
cc_148 N_A3_c_158_n N_A2_c_190_n 0.0670278f $X=1.735 $Y=1.765 $X2=0 $Y2=0
cc_149 N_A3_c_159_n N_A2_c_191_n 0.00224187f $X=1.78 $Y=1.22 $X2=0 $Y2=0
cc_150 A3 N_A2_c_191_n 0.0271823f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_151 N_A3_c_158_n N_VPWR_c_272_n 0.00700002f $X=1.735 $Y=1.765 $X2=0 $Y2=0
cc_152 N_A3_c_158_n N_VPWR_c_275_n 0.00481995f $X=1.735 $Y=1.765 $X2=0 $Y2=0
cc_153 N_A3_c_158_n N_VPWR_c_269_n 0.00508379f $X=1.735 $Y=1.765 $X2=0 $Y2=0
cc_154 N_A3_c_158_n N_A_362_368#_c_349_n 0.0102336f $X=1.735 $Y=1.765 $X2=0
+ $Y2=0
cc_155 N_A3_c_159_n N_VGND_c_380_n 0.00384553f $X=1.78 $Y=1.22 $X2=0 $Y2=0
cc_156 N_A3_c_159_n N_VGND_c_381_n 0.0103313f $X=1.78 $Y=1.22 $X2=0 $Y2=0
cc_157 N_A3_c_159_n N_VGND_c_382_n 0.00383677f $X=1.78 $Y=1.22 $X2=0 $Y2=0
cc_158 N_A2_c_189_n N_A1_c_217_n 0.0301845f $X=2.17 $Y=1.22 $X2=-0.19 $Y2=-0.245
cc_159 N_A2_c_190_n N_A1_c_218_n 0.0479837f $X=2.185 $Y=1.765 $X2=0 $Y2=0
cc_160 N_A2_c_191_n N_A1_c_218_n 4.20673e-19 $X=2.26 $Y=1.385 $X2=0 $Y2=0
cc_161 N_A2_c_190_n A1 4.18553e-19 $X=2.185 $Y=1.765 $X2=0 $Y2=0
cc_162 N_A2_c_191_n A1 0.0224075f $X=2.26 $Y=1.385 $X2=0 $Y2=0
cc_163 N_A2_c_190_n N_VPWR_c_273_n 0.00779845f $X=2.185 $Y=1.765 $X2=0 $Y2=0
cc_164 N_A2_c_190_n N_VPWR_c_275_n 0.00481995f $X=2.185 $Y=1.765 $X2=0 $Y2=0
cc_165 N_A2_c_190_n N_VPWR_c_269_n 0.00508379f $X=2.185 $Y=1.765 $X2=0 $Y2=0
cc_166 N_A2_c_190_n N_A_362_368#_c_353_n 0.0127987f $X=2.185 $Y=1.765 $X2=0
+ $Y2=0
cc_167 N_A2_c_190_n N_A_362_368#_c_349_n 0.0112251f $X=2.185 $Y=1.765 $X2=0
+ $Y2=0
cc_168 N_A2_c_190_n N_A_362_368#_c_350_n 8.23919e-19 $X=2.185 $Y=1.765 $X2=0
+ $Y2=0
cc_169 N_A2_c_189_n N_VGND_c_380_n 0.00461464f $X=2.17 $Y=1.22 $X2=0 $Y2=0
cc_170 N_A2_c_189_n N_VGND_c_381_n 0.00178416f $X=2.17 $Y=1.22 $X2=0 $Y2=0
cc_171 N_A2_c_189_n N_VGND_c_382_n 0.00465551f $X=2.17 $Y=1.22 $X2=0 $Y2=0
cc_172 N_A1_c_217_n N_B1_c_248_n 0.0234037f $X=2.74 $Y=1.22 $X2=-0.19 $Y2=-0.245
cc_173 A1 N_B1_c_248_n 0.00355487f $X=3.035 $Y=1.21 $X2=-0.19 $Y2=-0.245
cc_174 N_A1_c_218_n N_B1_c_249_n 0.0535236f $X=2.825 $Y=1.765 $X2=0 $Y2=0
cc_175 N_A1_c_218_n B1 2.16754e-19 $X=2.825 $Y=1.765 $X2=0 $Y2=0
cc_176 A1 B1 0.0290828f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_177 N_A1_c_218_n N_VPWR_c_273_n 0.00792131f $X=2.825 $Y=1.765 $X2=0 $Y2=0
cc_178 N_A1_c_218_n N_VPWR_c_276_n 0.00481995f $X=2.825 $Y=1.765 $X2=0 $Y2=0
cc_179 N_A1_c_218_n N_VPWR_c_269_n 0.00508379f $X=2.825 $Y=1.765 $X2=0 $Y2=0
cc_180 N_A1_c_218_n N_A_362_368#_c_353_n 0.0127987f $X=2.825 $Y=1.765 $X2=0
+ $Y2=0
cc_181 N_A1_c_218_n N_A_362_368#_c_349_n 8.32166e-19 $X=2.825 $Y=1.765 $X2=0
+ $Y2=0
cc_182 N_A1_c_218_n N_A_362_368#_c_350_n 0.0108459f $X=2.825 $Y=1.765 $X2=0
+ $Y2=0
cc_183 N_A1_c_217_n N_VGND_c_378_n 7.29208e-19 $X=2.74 $Y=1.22 $X2=0 $Y2=0
cc_184 N_A1_c_217_n N_VGND_c_380_n 0.00461464f $X=2.74 $Y=1.22 $X2=0 $Y2=0
cc_185 N_A1_c_217_n N_VGND_c_382_n 0.00467093f $X=2.74 $Y=1.22 $X2=0 $Y2=0
cc_186 N_B1_c_249_n N_VPWR_c_276_n 0.00481995f $X=3.325 $Y=1.765 $X2=0 $Y2=0
cc_187 N_B1_c_249_n N_VPWR_c_269_n 0.00508379f $X=3.325 $Y=1.765 $X2=0 $Y2=0
cc_188 N_B1_c_249_n N_A_362_368#_c_350_n 0.00341658f $X=3.325 $Y=1.765 $X2=0
+ $Y2=0
cc_189 N_B1_c_248_n N_VGND_c_378_n 0.0134916f $X=3.31 $Y=1.22 $X2=0 $Y2=0
cc_190 N_B1_c_249_n N_VGND_c_378_n 0.00190818f $X=3.325 $Y=1.765 $X2=0 $Y2=0
cc_191 B1 N_VGND_c_378_n 0.0232669f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_192 N_B1_c_248_n N_VGND_c_380_n 0.00383152f $X=3.31 $Y=1.22 $X2=0 $Y2=0
cc_193 N_B1_c_248_n N_VGND_c_382_n 0.00758792f $X=3.31 $Y=1.22 $X2=0 $Y2=0
cc_194 N_VPWR_c_271_n X 0.0878655f $X=0.35 $Y=1.985 $X2=0 $Y2=0
cc_195 N_VPWR_c_272_n X 0.0379525f $X=1.255 $Y=2.145 $X2=0 $Y2=0
cc_196 N_VPWR_c_274_n X 0.0138348f $X=1.09 $Y=3.33 $X2=0 $Y2=0
cc_197 N_VPWR_c_269_n X 0.0113479f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_198 N_VPWR_M1011_d N_A_362_368#_c_353_n 0.0103765f $X=2.26 $Y=1.84 $X2=0
+ $Y2=0
cc_199 N_VPWR_c_273_n N_A_362_368#_c_353_n 0.0266856f $X=2.515 $Y=2.565 $X2=0
+ $Y2=0
cc_200 N_VPWR_c_272_n N_A_362_368#_c_349_n 0.0244519f $X=1.255 $Y=2.145 $X2=0
+ $Y2=0
cc_201 N_VPWR_c_273_n N_A_362_368#_c_349_n 0.0288223f $X=2.515 $Y=2.565 $X2=0
+ $Y2=0
cc_202 N_VPWR_c_275_n N_A_362_368#_c_349_n 0.00976219f $X=2.35 $Y=3.33 $X2=0
+ $Y2=0
cc_203 N_VPWR_c_269_n N_A_362_368#_c_349_n 0.0111764f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_204 N_VPWR_c_273_n N_A_362_368#_c_350_n 0.0309481f $X=2.515 $Y=2.565 $X2=0
+ $Y2=0
cc_205 N_VPWR_c_276_n N_A_362_368#_c_350_n 0.0097982f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_206 N_VPWR_c_269_n N_A_362_368#_c_350_n 0.0111907f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_207 N_X_c_319_n N_VGND_c_376_n 0.0300058f $X=0.78 $Y=0.515 $X2=0 $Y2=0
cc_208 N_X_c_319_n N_VGND_c_379_n 0.0121098f $X=0.78 $Y=0.515 $X2=0 $Y2=0
cc_209 N_X_c_319_n N_VGND_c_381_n 0.0112219f $X=0.78 $Y=0.515 $X2=0 $Y2=0
cc_210 N_X_c_319_n N_VGND_c_382_n 0.00996704f $X=0.78 $Y=0.515 $X2=0 $Y2=0
