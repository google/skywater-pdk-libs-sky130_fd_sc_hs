* File: sky130_fd_sc_hs__sdfrtp_2.pxi.spice
* Created: Tue Sep  1 20:22:45 2020
* 
x_PM_SKY130_FD_SC_HS__SDFRTP_2%A_27_74# N_A_27_74#_M1039_s N_A_27_74#_M1020_s
+ N_A_27_74#_c_280_n N_A_27_74#_c_281_n N_A_27_74#_M1010_g N_A_27_74#_c_287_n
+ N_A_27_74#_M1036_g N_A_27_74#_c_282_n N_A_27_74#_c_283_n N_A_27_74#_c_289_n
+ N_A_27_74#_c_284_n N_A_27_74#_c_290_n N_A_27_74#_c_285_n N_A_27_74#_c_291_n
+ N_A_27_74#_c_292_n N_A_27_74#_c_286_n PM_SKY130_FD_SC_HS__SDFRTP_2%A_27_74#
x_PM_SKY130_FD_SC_HS__SDFRTP_2%SCE N_SCE_c_369_n N_SCE_M1039_g N_SCE_c_370_n
+ N_SCE_M1020_g N_SCE_c_371_n N_SCE_c_372_n N_SCE_M1017_g N_SCE_M1006_g
+ N_SCE_c_362_n N_SCE_c_363_n N_SCE_c_364_n N_SCE_c_365_n SCE SCE SCE
+ N_SCE_c_366_n N_SCE_c_367_n SCE N_SCE_c_368_n PM_SKY130_FD_SC_HS__SDFRTP_2%SCE
x_PM_SKY130_FD_SC_HS__SDFRTP_2%D N_D_c_444_n N_D_M1011_g N_D_c_445_n N_D_c_449_n
+ N_D_M1033_g D N_D_c_446_n N_D_c_447_n PM_SKY130_FD_SC_HS__SDFRTP_2%D
x_PM_SKY130_FD_SC_HS__SDFRTP_2%SCD N_SCD_c_493_n N_SCD_M1005_g N_SCD_M1038_g
+ N_SCD_c_490_n SCD SCD N_SCD_c_492_n PM_SKY130_FD_SC_HS__SDFRTP_2%SCD
x_PM_SKY130_FD_SC_HS__SDFRTP_2%RESET_B N_RESET_B_M1002_g N_RESET_B_c_544_n
+ N_RESET_B_M1041_g N_RESET_B_c_539_n N_RESET_B_M1021_g N_RESET_B_c_545_n
+ N_RESET_B_M1037_g N_RESET_B_c_540_n N_RESET_B_M1023_g N_RESET_B_c_548_n
+ N_RESET_B_c_549_n N_RESET_B_M1026_g N_RESET_B_c_542_n N_RESET_B_c_550_n
+ N_RESET_B_c_551_n N_RESET_B_c_552_n N_RESET_B_c_553_n N_RESET_B_c_554_n
+ RESET_B N_RESET_B_c_555_n N_RESET_B_c_556_n N_RESET_B_c_557_n
+ N_RESET_B_c_558_n N_RESET_B_c_653_p PM_SKY130_FD_SC_HS__SDFRTP_2%RESET_B
x_PM_SKY130_FD_SC_HS__SDFRTP_2%CLK N_CLK_c_735_n N_CLK_M1018_g N_CLK_M1019_g
+ N_CLK_c_737_n N_CLK_c_748_n CLK N_CLK_c_738_n PM_SKY130_FD_SC_HS__SDFRTP_2%CLK
x_PM_SKY130_FD_SC_HS__SDFRTP_2%A_1034_368# N_A_1034_368#_M1007_d
+ N_A_1034_368#_M1032_d N_A_1034_368#_c_812_n N_A_1034_368#_c_813_n
+ N_A_1034_368#_M1028_g N_A_1034_368#_c_790_n N_A_1034_368#_c_791_n
+ N_A_1034_368#_M1003_g N_A_1034_368#_c_793_n N_A_1034_368#_M1024_g
+ N_A_1034_368#_c_794_n N_A_1034_368#_c_795_n N_A_1034_368#_c_816_n
+ N_A_1034_368#_M1027_g N_A_1034_368#_c_796_n N_A_1034_368#_c_797_n
+ N_A_1034_368#_c_798_n N_A_1034_368#_c_799_n N_A_1034_368#_c_800_n
+ N_A_1034_368#_c_801_n N_A_1034_368#_c_972_p N_A_1034_368#_c_802_n
+ N_A_1034_368#_c_803_n N_A_1034_368#_c_858_p N_A_1034_368#_c_804_n
+ N_A_1034_368#_c_805_n N_A_1034_368#_c_806_n N_A_1034_368#_c_807_n
+ N_A_1034_368#_c_808_n N_A_1034_368#_c_809_n N_A_1034_368#_c_810_n
+ N_A_1034_368#_c_811_n PM_SKY130_FD_SC_HS__SDFRTP_2%A_1034_368#
x_PM_SKY130_FD_SC_HS__SDFRTP_2%A_1383_349# N_A_1383_349#_M1040_d
+ N_A_1383_349#_M1016_d N_A_1383_349#_c_996_n N_A_1383_349#_M1000_g
+ N_A_1383_349#_M1035_g N_A_1383_349#_c_993_n N_A_1383_349#_c_1013_n
+ N_A_1383_349#_c_1030_n N_A_1383_349#_c_999_n N_A_1383_349#_c_994_n
+ N_A_1383_349#_c_1000_n N_A_1383_349#_c_995_n
+ PM_SKY130_FD_SC_HS__SDFRTP_2%A_1383_349#
x_PM_SKY130_FD_SC_HS__SDFRTP_2%A_1242_457# N_A_1242_457#_M1004_d
+ N_A_1242_457#_M1028_d N_A_1242_457#_M1037_d N_A_1242_457#_M1040_g
+ N_A_1242_457#_c_1083_n N_A_1242_457#_M1016_g N_A_1242_457#_c_1084_n
+ N_A_1242_457#_c_1092_n N_A_1242_457#_c_1085_n N_A_1242_457#_c_1105_n
+ N_A_1242_457#_c_1086_n N_A_1242_457#_c_1087_n N_A_1242_457#_c_1088_n
+ N_A_1242_457#_c_1089_n N_A_1242_457#_c_1095_n
+ PM_SKY130_FD_SC_HS__SDFRTP_2%A_1242_457#
x_PM_SKY130_FD_SC_HS__SDFRTP_2%A_855_368# N_A_855_368#_M1019_s
+ N_A_855_368#_M1018_s N_A_855_368#_c_1202_n N_A_855_368#_M1032_g
+ N_A_855_368#_M1007_g N_A_855_368#_c_1204_n N_A_855_368#_c_1205_n
+ N_A_855_368#_c_1206_n N_A_855_368#_c_1219_n N_A_855_368#_c_1220_n
+ N_A_855_368#_M1004_g N_A_855_368#_c_1221_n N_A_855_368#_c_1222_n
+ N_A_855_368#_c_1223_n N_A_855_368#_M1034_g N_A_855_368#_c_1224_n
+ N_A_855_368#_M1025_g N_A_855_368#_c_1208_n N_A_855_368#_c_1227_n
+ N_A_855_368#_c_1209_n N_A_855_368#_M1008_g N_A_855_368#_c_1211_n
+ N_A_855_368#_c_1228_n N_A_855_368#_c_1229_n N_A_855_368#_c_1212_n
+ N_A_855_368#_c_1213_n N_A_855_368#_c_1253_n N_A_855_368#_c_1255_n
+ N_A_855_368#_c_1230_n N_A_855_368#_c_1214_n N_A_855_368#_c_1215_n
+ N_A_855_368#_c_1232_n N_A_855_368#_c_1216_n
+ PM_SKY130_FD_SC_HS__SDFRTP_2%A_855_368#
x_PM_SKY130_FD_SC_HS__SDFRTP_2%A_2082_446# N_A_2082_446#_M1013_d
+ N_A_2082_446#_M1026_d N_A_2082_446#_c_1408_n N_A_2082_446#_M1015_g
+ N_A_2082_446#_M1009_g N_A_2082_446#_c_1409_n N_A_2082_446#_c_1419_n
+ N_A_2082_446#_c_1400_n N_A_2082_446#_c_1401_n N_A_2082_446#_c_1412_n
+ N_A_2082_446#_c_1469_p N_A_2082_446#_c_1413_n N_A_2082_446#_c_1402_n
+ N_A_2082_446#_c_1403_n N_A_2082_446#_c_1404_n N_A_2082_446#_c_1405_n
+ N_A_2082_446#_c_1406_n N_A_2082_446#_c_1407_n
+ PM_SKY130_FD_SC_HS__SDFRTP_2%A_2082_446#
x_PM_SKY130_FD_SC_HS__SDFRTP_2%A_1824_74# N_A_1824_74#_M1024_d
+ N_A_1824_74#_M1025_d N_A_1824_74#_M1013_g N_A_1824_74#_c_1535_n
+ N_A_1824_74#_c_1536_n N_A_1824_74#_c_1537_n N_A_1824_74#_M1029_g
+ N_A_1824_74#_c_1522_n N_A_1824_74#_c_1523_n N_A_1824_74#_c_1524_n
+ N_A_1824_74#_c_1539_n N_A_1824_74#_M1022_g N_A_1824_74#_c_1525_n
+ N_A_1824_74#_M1030_g N_A_1824_74#_c_1526_n N_A_1824_74#_c_1527_n
+ N_A_1824_74#_c_1553_n N_A_1824_74#_c_1528_n N_A_1824_74#_c_1540_n
+ N_A_1824_74#_c_1541_n N_A_1824_74#_c_1529_n N_A_1824_74#_c_1530_n
+ N_A_1824_74#_c_1531_n N_A_1824_74#_c_1532_n N_A_1824_74#_c_1533_n
+ N_A_1824_74#_c_1534_n PM_SKY130_FD_SC_HS__SDFRTP_2%A_1824_74#
x_PM_SKY130_FD_SC_HS__SDFRTP_2%A_2492_392# N_A_2492_392#_M1030_d
+ N_A_2492_392#_M1022_d N_A_2492_392#_c_1672_n N_A_2492_392#_M1012_g
+ N_A_2492_392#_M1001_g N_A_2492_392#_c_1673_n N_A_2492_392#_M1014_g
+ N_A_2492_392#_M1031_g N_A_2492_392#_c_1674_n N_A_2492_392#_c_1675_n
+ N_A_2492_392#_c_1667_n N_A_2492_392#_c_1668_n N_A_2492_392#_c_1669_n
+ N_A_2492_392#_c_1670_n N_A_2492_392#_c_1671_n
+ PM_SKY130_FD_SC_HS__SDFRTP_2%A_2492_392#
x_PM_SKY130_FD_SC_HS__SDFRTP_2%VPWR N_VPWR_M1020_d N_VPWR_M1005_d N_VPWR_M1018_d
+ N_VPWR_M1000_d N_VPWR_M1016_s N_VPWR_M1015_d N_VPWR_M1029_d N_VPWR_M1012_s
+ N_VPWR_M1014_s N_VPWR_c_1728_n N_VPWR_c_1729_n N_VPWR_c_1730_n N_VPWR_c_1731_n
+ N_VPWR_c_1732_n N_VPWR_c_1733_n N_VPWR_c_1734_n N_VPWR_c_1735_n
+ N_VPWR_c_1736_n N_VPWR_c_1737_n N_VPWR_c_1738_n N_VPWR_c_1739_n
+ N_VPWR_c_1740_n N_VPWR_c_1741_n VPWR N_VPWR_c_1742_n N_VPWR_c_1743_n
+ N_VPWR_c_1744_n N_VPWR_c_1745_n N_VPWR_c_1746_n N_VPWR_c_1747_n
+ N_VPWR_c_1748_n N_VPWR_c_1749_n N_VPWR_c_1750_n N_VPWR_c_1751_n
+ N_VPWR_c_1752_n N_VPWR_c_1727_n PM_SKY130_FD_SC_HS__SDFRTP_2%VPWR
x_PM_SKY130_FD_SC_HS__SDFRTP_2%A_390_81# N_A_390_81#_M1011_d N_A_390_81#_M1004_s
+ N_A_390_81#_M1033_d N_A_390_81#_M1041_d N_A_390_81#_M1028_s
+ N_A_390_81#_c_1902_n N_A_390_81#_c_1919_n N_A_390_81#_c_1903_n
+ N_A_390_81#_c_1904_n N_A_390_81#_c_1905_n N_A_390_81#_c_1906_n
+ N_A_390_81#_c_1912_n N_A_390_81#_c_1913_n N_A_390_81#_c_1914_n
+ N_A_390_81#_c_1907_n N_A_390_81#_c_1915_n N_A_390_81#_c_1908_n
+ N_A_390_81#_c_1909_n N_A_390_81#_c_1910_n N_A_390_81#_c_1917_n
+ N_A_390_81#_c_1918_n PM_SKY130_FD_SC_HS__SDFRTP_2%A_390_81#
x_PM_SKY130_FD_SC_HS__SDFRTP_2%Q N_Q_M1001_d N_Q_M1012_d N_Q_c_2057_n Q Q Q Q
+ PM_SKY130_FD_SC_HS__SDFRTP_2%Q
x_PM_SKY130_FD_SC_HS__SDFRTP_2%VGND N_VGND_M1039_d N_VGND_M1002_d N_VGND_M1019_d
+ N_VGND_M1021_d N_VGND_M1009_d N_VGND_M1030_s N_VGND_M1001_s N_VGND_M1031_s
+ N_VGND_c_2078_n N_VGND_c_2079_n N_VGND_c_2080_n N_VGND_c_2081_n
+ N_VGND_c_2082_n N_VGND_c_2083_n N_VGND_c_2084_n N_VGND_c_2085_n
+ N_VGND_c_2086_n N_VGND_c_2087_n VGND N_VGND_c_2088_n N_VGND_c_2089_n
+ N_VGND_c_2090_n N_VGND_c_2091_n N_VGND_c_2092_n N_VGND_c_2093_n
+ N_VGND_c_2094_n N_VGND_c_2095_n N_VGND_c_2096_n N_VGND_c_2097_n
+ N_VGND_c_2098_n N_VGND_c_2099_n N_VGND_c_2100_n
+ PM_SKY130_FD_SC_HS__SDFRTP_2%VGND
x_PM_SKY130_FD_SC_HS__SDFRTP_2%noxref_24 N_noxref_24_M1010_s N_noxref_24_M1038_d
+ N_noxref_24_c_2215_n N_noxref_24_c_2216_n N_noxref_24_c_2217_n
+ PM_SKY130_FD_SC_HS__SDFRTP_2%noxref_24
cc_1 VNB N_A_27_74#_c_280_n 0.0258189f $X=-0.19 $Y=-0.245 $X2=1.41 $Y2=1.01
cc_2 VNB N_A_27_74#_c_281_n 0.0202565f $X=-0.19 $Y=-0.245 $X2=1.485 $Y2=0.935
cc_3 VNB N_A_27_74#_c_282_n 0.0257773f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=0.58
cc_4 VNB N_A_27_74#_c_283_n 0.0190417f $X=-0.19 $Y=-0.245 $X2=0.2 $Y2=2.005
cc_5 VNB N_A_27_74#_c_284_n 0.00987534f $X=-0.19 $Y=-0.245 $X2=0.975 $Y2=1.1
cc_6 VNB N_A_27_74#_c_285_n 0.018224f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.1
cc_7 VNB N_A_27_74#_c_286_n 0.0395906f $X=-0.19 $Y=-0.245 $X2=0.975 $Y2=1.01
cc_8 VNB N_SCE_M1039_g 0.0668709f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_SCE_M1006_g 0.0362271f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=0.58
cc_10 VNB N_SCE_c_362_n 0.00775502f $X=-0.19 $Y=-0.245 $X2=0.2 $Y2=2.005
cc_11 VNB N_SCE_c_363_n 0.0420954f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=2.175
cc_12 VNB N_SCE_c_364_n 0.01245f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=2.465
cc_13 VNB N_SCE_c_365_n 0.00344346f $X=-0.19 $Y=-0.245 $X2=0.365 $Y2=1.1
cc_14 VNB N_SCE_c_366_n 0.0351466f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_SCE_c_367_n 0.0106235f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_SCE_c_368_n 0.00168276f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_D_c_444_n 0.0162211f $X=-0.19 $Y=-0.245 $X2=0.135 $Y2=0.37
cc_18 VNB N_D_c_445_n 0.0275832f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_D_c_446_n 0.00758117f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=0.935
cc_20 VNB N_D_c_447_n 0.0380459f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=0.58
cc_21 VNB N_SCD_M1038_g 0.0431772f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_SCD_c_490_n 0.00107072f $X=-0.19 $Y=-0.245 $X2=1.485 $Y2=0.615
cc_23 VNB SCD 0.00167055f $X=-0.19 $Y=-0.245 $X2=1.485 $Y2=0.615
cc_24 VNB N_SCD_c_492_n 0.0170281f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=0.58
cc_25 VNB N_RESET_B_M1002_g 0.0676013f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_RESET_B_c_539_n 0.0185871f $X=-0.19 $Y=-0.245 $X2=1.14 $Y2=1.01
cc_27 VNB N_RESET_B_c_540_n 0.0189013f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=0.935
cc_28 VNB N_RESET_B_M1023_g 0.0531601f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_RESET_B_c_542_n 0.0224087f $X=-0.19 $Y=-0.245 $X2=0.975 $Y2=1.1
cc_30 VNB N_CLK_c_735_n 0.0212209f $X=-0.19 $Y=-0.245 $X2=0.135 $Y2=0.37
cc_31 VNB N_CLK_M1019_g 0.0236484f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_CLK_c_737_n 0.060774f $X=-0.19 $Y=-0.245 $X2=1.485 $Y2=0.935
cc_33 VNB N_CLK_c_738_n 0.0111142f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=2.465
cc_34 VNB N_A_1034_368#_c_790_n 0.00766157f $X=-0.19 $Y=-0.245 $X2=2.495
+ $Y2=2.245
cc_35 VNB N_A_1034_368#_c_791_n 0.0255078f $X=-0.19 $Y=-0.245 $X2=2.495 $Y2=2.64
cc_36 VNB N_A_1034_368#_M1003_g 0.0226179f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=0.58
cc_37 VNB N_A_1034_368#_c_793_n 0.0171555f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_1034_368#_c_794_n 0.0222225f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=2.175
cc_39 VNB N_A_1034_368#_c_795_n 0.0102361f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=2.465
cc_40 VNB N_A_1034_368#_c_796_n 0.00706325f $X=-0.19 $Y=-0.245 $X2=2.375
+ $Y2=2.09
cc_41 VNB N_A_1034_368#_c_797_n 0.00336558f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.1
cc_42 VNB N_A_1034_368#_c_798_n 0.0412728f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=2.09
cc_43 VNB N_A_1034_368#_c_799_n 0.00390309f $X=-0.19 $Y=-0.245 $X2=2.54
+ $Y2=1.995
cc_44 VNB N_A_1034_368#_c_800_n 0.00190641f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_A_1034_368#_c_801_n 0.00328545f $X=-0.19 $Y=-0.245 $X2=0.975
+ $Y2=1.01
cc_46 VNB N_A_1034_368#_c_802_n 0.00854373f $X=-0.19 $Y=-0.245 $X2=2.54
+ $Y2=1.995
cc_47 VNB N_A_1034_368#_c_803_n 0.00245962f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_1034_368#_c_804_n 0.00595338f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A_1034_368#_c_805_n 0.00363165f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_A_1034_368#_c_806_n 0.0322711f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_A_1034_368#_c_807_n 0.0101868f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_A_1034_368#_c_808_n 2.31855e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_A_1034_368#_c_809_n 0.00412914f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_A_1034_368#_c_810_n 0.0108699f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_A_1034_368#_c_811_n 0.0070601f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_A_1383_349#_M1035_g 0.0373116f $X=-0.19 $Y=-0.245 $X2=2.495
+ $Y2=2.245
cc_57 VNB N_A_1383_349#_c_993_n 0.00395139f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=0.58
cc_58 VNB N_A_1383_349#_c_994_n 0.00239154f $X=-0.19 $Y=-0.245 $X2=0.975 $Y2=1.1
cc_59 VNB N_A_1383_349#_c_995_n 0.0143226f $X=-0.19 $Y=-0.245 $X2=2.54 $Y2=1.995
cc_60 VNB N_A_1242_457#_M1040_g 0.0241865f $X=-0.19 $Y=-0.245 $X2=2.495
+ $Y2=2.245
cc_61 VNB N_A_1242_457#_c_1083_n 0.0171771f $X=-0.19 $Y=-0.245 $X2=2.495
+ $Y2=2.64
cc_62 VNB N_A_1242_457#_c_1084_n 0.0274099f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_A_1242_457#_c_1085_n 0.00406303f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_A_1242_457#_c_1086_n 5.47821e-19 $X=-0.19 $Y=-0.245 $X2=0.975
+ $Y2=1.1
cc_65 VNB N_A_1242_457#_c_1087_n 0.00159936f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_A_1242_457#_c_1088_n 0.00560512f $X=-0.19 $Y=-0.245 $X2=0.445
+ $Y2=2.09
cc_67 VNB N_A_1242_457#_c_1089_n 0.00553892f $X=-0.19 $Y=-0.245 $X2=2.54
+ $Y2=1.995
cc_68 VNB N_A_855_368#_c_1202_n 0.0315269f $X=-0.19 $Y=-0.245 $X2=1.41 $Y2=1.01
cc_69 VNB N_A_855_368#_M1007_g 0.0232873f $X=-0.19 $Y=-0.245 $X2=2.495 $Y2=2.245
cc_70 VNB N_A_855_368#_c_1204_n 0.00980266f $X=-0.19 $Y=-0.245 $X2=2.495
+ $Y2=2.64
cc_71 VNB N_A_855_368#_c_1205_n 0.0122914f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=0.58
cc_72 VNB N_A_855_368#_c_1206_n 0.0333628f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_A_855_368#_M1004_g 0.0210546f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_A_855_368#_c_1208_n 0.012531f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_A_855_368#_c_1209_n 0.0236403f $X=-0.19 $Y=-0.245 $X2=0.975 $Y2=1.01
cc_76 VNB N_A_855_368#_M1008_g 0.027022f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_A_855_368#_c_1211_n 0.00789845f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_A_855_368#_c_1212_n 0.0209137f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VNB N_A_855_368#_c_1213_n 0.00192022f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_A_855_368#_c_1214_n 0.00314875f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_81 VNB N_A_855_368#_c_1215_n 0.00106788f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_82 VNB N_A_855_368#_c_1216_n 0.00438178f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_83 VNB N_A_2082_446#_M1009_g 0.0407896f $X=-0.19 $Y=-0.245 $X2=2.495
+ $Y2=2.245
cc_84 VNB N_A_2082_446#_c_1400_n 0.00604102f $X=-0.19 $Y=-0.245 $X2=0.2
+ $Y2=1.265
cc_85 VNB N_A_2082_446#_c_1401_n 0.00978233f $X=-0.19 $Y=-0.245 $X2=0.2
+ $Y2=2.005
cc_86 VNB N_A_2082_446#_c_1402_n 0.00743589f $X=-0.19 $Y=-0.245 $X2=2.375
+ $Y2=2.09
cc_87 VNB N_A_2082_446#_c_1403_n 0.00688415f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.1
cc_88 VNB N_A_2082_446#_c_1404_n 0.00281201f $X=-0.19 $Y=-0.245 $X2=0.28
+ $Y2=2.09
cc_89 VNB N_A_2082_446#_c_1405_n 0.00528256f $X=-0.19 $Y=-0.245 $X2=2.54
+ $Y2=1.995
cc_90 VNB N_A_2082_446#_c_1406_n 0.00129589f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_91 VNB N_A_2082_446#_c_1407_n 0.0231274f $X=-0.19 $Y=-0.245 $X2=2.54 $Y2=2.09
cc_92 VNB N_A_1824_74#_M1013_g 0.0313995f $X=-0.19 $Y=-0.245 $X2=1.485 $Y2=0.935
cc_93 VNB N_A_1824_74#_c_1522_n 0.0313227f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_94 VNB N_A_1824_74#_c_1523_n 0.0323107f $X=-0.19 $Y=-0.245 $X2=0.2 $Y2=1.265
cc_95 VNB N_A_1824_74#_c_1524_n 0.0156535f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=2.175
cc_96 VNB N_A_1824_74#_c_1525_n 0.0193338f $X=-0.19 $Y=-0.245 $X2=0.365 $Y2=1.1
cc_97 VNB N_A_1824_74#_c_1526_n 0.0143534f $X=-0.19 $Y=-0.245 $X2=0.975 $Y2=1.1
cc_98 VNB N_A_1824_74#_c_1527_n 0.0203145f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_99 VNB N_A_1824_74#_c_1528_n 0.00728448f $X=-0.19 $Y=-0.245 $X2=2.54
+ $Y2=1.995
cc_100 VNB N_A_1824_74#_c_1529_n 0.00580575f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_101 VNB N_A_1824_74#_c_1530_n 0.00783827f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_102 VNB N_A_1824_74#_c_1531_n 0.0103967f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_103 VNB N_A_1824_74#_c_1532_n 4.11765e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_104 VNB N_A_1824_74#_c_1533_n 0.0164314f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_105 VNB N_A_1824_74#_c_1534_n 0.00253069f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_106 VNB N_A_2492_392#_M1001_g 0.0229518f $X=-0.19 $Y=-0.245 $X2=2.495
+ $Y2=2.245
cc_107 VNB N_A_2492_392#_M1031_g 0.0260209f $X=-0.19 $Y=-0.245 $X2=0.2 $Y2=1.265
cc_108 VNB N_A_2492_392#_c_1667_n 0.0162202f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_109 VNB N_A_2492_392#_c_1668_n 0.0113264f $X=-0.19 $Y=-0.245 $X2=2.54
+ $Y2=1.995
cc_110 VNB N_A_2492_392#_c_1669_n 7.87382e-19 $X=-0.19 $Y=-0.245 $X2=2.54
+ $Y2=2.09
cc_111 VNB N_A_2492_392#_c_1670_n 0.00922601f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_112 VNB N_A_2492_392#_c_1671_n 0.0953071f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_113 VNB N_VPWR_c_1727_n 0.601534f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_114 VNB N_A_390_81#_c_1902_n 0.00895762f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_115 VNB N_A_390_81#_c_1903_n 0.00275942f $X=-0.19 $Y=-0.245 $X2=0.365 $Y2=1.1
cc_116 VNB N_A_390_81#_c_1904_n 0.0135173f $X=-0.19 $Y=-0.245 $X2=0.975 $Y2=1.1
cc_117 VNB N_A_390_81#_c_1905_n 0.00472946f $X=-0.19 $Y=-0.245 $X2=0.975 $Y2=1.1
cc_118 VNB N_A_390_81#_c_1906_n 0.00291665f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_119 VNB N_A_390_81#_c_1907_n 0.00721563f $X=-0.19 $Y=-0.245 $X2=2.54
+ $Y2=1.995
cc_120 VNB N_A_390_81#_c_1908_n 0.00546923f $X=-0.19 $Y=-0.245 $X2=0.975
+ $Y2=1.01
cc_121 VNB N_A_390_81#_c_1909_n 0.00265013f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_122 VNB N_A_390_81#_c_1910_n 0.00287507f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_123 VNB N_Q_c_2057_n 2.86109e-19 $X=-0.19 $Y=-0.245 $X2=1.485 $Y2=0.935
cc_124 VNB Q 0.00240191f $X=-0.19 $Y=-0.245 $X2=2.495 $Y2=2.64
cc_125 VNB N_VGND_c_2078_n 0.0110567f $X=-0.19 $Y=-0.245 $X2=0.975 $Y2=1.1
cc_126 VNB N_VGND_c_2079_n 0.0270283f $X=-0.19 $Y=-0.245 $X2=0.445 $Y2=2.09
cc_127 VNB N_VGND_c_2080_n 0.00632134f $X=-0.19 $Y=-0.245 $X2=2.54 $Y2=1.995
cc_128 VNB N_VGND_c_2081_n 0.0067048f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_129 VNB N_VGND_c_2082_n 0.00861345f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_130 VNB N_VGND_c_2083_n 0.0169646f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_131 VNB N_VGND_c_2084_n 0.010678f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_132 VNB N_VGND_c_2085_n 0.0505973f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_133 VNB N_VGND_c_2086_n 0.0673948f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_134 VNB N_VGND_c_2087_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_135 VNB N_VGND_c_2088_n 0.0173909f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_136 VNB N_VGND_c_2089_n 0.0205822f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_137 VNB N_VGND_c_2090_n 0.0833231f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_138 VNB N_VGND_c_2091_n 0.0684884f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_139 VNB N_VGND_c_2092_n 0.0296745f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_140 VNB N_VGND_c_2093_n 0.0187654f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_141 VNB N_VGND_c_2094_n 0.0193312f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_142 VNB N_VGND_c_2095_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_143 VNB N_VGND_c_2096_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_144 VNB N_VGND_c_2097_n 0.00604233f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_145 VNB N_VGND_c_2098_n 0.00613227f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_146 VNB N_VGND_c_2099_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_147 VNB N_VGND_c_2100_n 0.792467f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_148 VNB N_noxref_24_c_2215_n 0.0170004f $X=-0.19 $Y=-0.245 $X2=1.41 $Y2=1.01
cc_149 VNB N_noxref_24_c_2216_n 0.00359395f $X=-0.19 $Y=-0.245 $X2=1.485
+ $Y2=0.615
cc_150 VNB N_noxref_24_c_2217_n 0.00655627f $X=-0.19 $Y=-0.245 $X2=2.495
+ $Y2=2.64
cc_151 VPB N_A_27_74#_c_287_n 0.0530057f $X=-0.19 $Y=1.66 $X2=2.495 $Y2=2.245
cc_152 VPB N_A_27_74#_c_283_n 0.016494f $X=-0.19 $Y=1.66 $X2=0.2 $Y2=2.005
cc_153 VPB N_A_27_74#_c_289_n 0.0338402f $X=-0.19 $Y=1.66 $X2=0.28 $Y2=2.465
cc_154 VPB N_A_27_74#_c_290_n 0.0351167f $X=-0.19 $Y=1.66 $X2=2.375 $Y2=2.09
cc_155 VPB N_A_27_74#_c_291_n 0.0129728f $X=-0.19 $Y=1.66 $X2=0.28 $Y2=2.09
cc_156 VPB N_A_27_74#_c_292_n 0.00362322f $X=-0.19 $Y=1.66 $X2=2.54 $Y2=1.995
cc_157 VPB N_SCE_c_369_n 0.0264922f $X=-0.19 $Y=1.66 $X2=0.135 $Y2=2.32
cc_158 VPB N_SCE_c_370_n 0.0318721f $X=-0.19 $Y=1.66 $X2=1.41 $Y2=1.01
cc_159 VPB N_SCE_c_371_n 0.0231924f $X=-0.19 $Y=1.66 $X2=1.485 $Y2=0.615
cc_160 VPB N_SCE_c_372_n 0.0275749f $X=-0.19 $Y=1.66 $X2=2.495 $Y2=2.245
cc_161 VPB N_SCE_c_362_n 0.00782879f $X=-0.19 $Y=1.66 $X2=0.2 $Y2=2.005
cc_162 VPB N_SCE_c_363_n 0.0410982f $X=-0.19 $Y=1.66 $X2=0.28 $Y2=2.175
cc_163 VPB N_SCE_c_365_n 0.00199215f $X=-0.19 $Y=1.66 $X2=0.365 $Y2=1.1
cc_164 VPB N_SCE_c_368_n 0.00270951f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_165 VPB N_D_c_445_n 0.030204f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_166 VPB N_D_c_449_n 0.0220375f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_167 VPB N_SCD_c_493_n 0.0170214f $X=-0.19 $Y=1.66 $X2=0.135 $Y2=0.37
cc_168 VPB N_SCD_c_490_n 0.0512537f $X=-0.19 $Y=1.66 $X2=1.485 $Y2=0.615
cc_169 VPB SCD 0.00146742f $X=-0.19 $Y=1.66 $X2=1.485 $Y2=0.615
cc_170 VPB N_RESET_B_M1002_g 0.0125098f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_171 VPB N_RESET_B_c_544_n 0.021814f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_172 VPB N_RESET_B_c_545_n 0.0178721f $X=-0.19 $Y=1.66 $X2=1.485 $Y2=0.615
cc_173 VPB N_RESET_B_c_540_n 0.0105327f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=0.935
cc_174 VPB N_RESET_B_M1023_g 0.0132171f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_175 VPB N_RESET_B_c_548_n 0.00850302f $X=-0.19 $Y=1.66 $X2=0.28 $Y2=2.175
cc_176 VPB N_RESET_B_c_549_n 0.0233033f $X=-0.19 $Y=1.66 $X2=0.28 $Y2=2.465
cc_177 VPB N_RESET_B_c_550_n 0.0195989f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_178 VPB N_RESET_B_c_551_n 0.00161953f $X=-0.19 $Y=1.66 $X2=2.375 $Y2=2.09
cc_179 VPB N_RESET_B_c_552_n 0.0135889f $X=-0.19 $Y=1.66 $X2=0.445 $Y2=2.09
cc_180 VPB N_RESET_B_c_553_n 3.23518e-19 $X=-0.19 $Y=1.66 $X2=0.24 $Y2=1.1
cc_181 VPB N_RESET_B_c_554_n 0.0118766f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_182 VPB N_RESET_B_c_555_n 0.0663796f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_183 VPB N_RESET_B_c_556_n 0.00233009f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_184 VPB N_RESET_B_c_557_n 0.0604769f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_185 VPB N_RESET_B_c_558_n 0.035184f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_186 VPB N_CLK_c_735_n 0.029777f $X=-0.19 $Y=1.66 $X2=0.135 $Y2=0.37
cc_187 VPB N_A_1034_368#_c_812_n 0.00944036f $X=-0.19 $Y=1.66 $X2=1.14 $Y2=1.01
cc_188 VPB N_A_1034_368#_c_813_n 0.0193299f $X=-0.19 $Y=1.66 $X2=1.485 $Y2=0.935
cc_189 VPB N_A_1034_368#_c_790_n 0.0111871f $X=-0.19 $Y=1.66 $X2=2.495 $Y2=2.245
cc_190 VPB N_A_1034_368#_c_791_n 0.0079794f $X=-0.19 $Y=1.66 $X2=2.495 $Y2=2.64
cc_191 VPB N_A_1034_368#_c_816_n 0.0670682f $X=-0.19 $Y=1.66 $X2=0.28 $Y2=2.465
cc_192 VPB N_A_1034_368#_c_800_n 0.0016505f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_193 VPB N_A_1034_368#_c_807_n 0.00643236f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_194 VPB N_A_1034_368#_c_808_n 0.00774017f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_195 VPB N_A_1034_368#_c_811_n 0.0242323f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_196 VPB N_A_1383_349#_c_996_n 0.069852f $X=-0.19 $Y=1.66 $X2=1.41 $Y2=1.01
cc_197 VPB N_A_1383_349#_M1035_g 0.00462646f $X=-0.19 $Y=1.66 $X2=2.495
+ $Y2=2.245
cc_198 VPB N_A_1383_349#_c_993_n 0.00156886f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=0.58
cc_199 VPB N_A_1383_349#_c_999_n 5.83952e-19 $X=-0.19 $Y=1.66 $X2=0.365 $Y2=1.1
cc_200 VPB N_A_1383_349#_c_1000_n 0.00552703f $X=-0.19 $Y=1.66 $X2=0.28 $Y2=2.09
cc_201 VPB N_A_1383_349#_c_995_n 0.00449517f $X=-0.19 $Y=1.66 $X2=2.54 $Y2=1.995
cc_202 VPB N_A_1242_457#_c_1083_n 0.0305943f $X=-0.19 $Y=1.66 $X2=2.495 $Y2=2.64
cc_203 VPB N_A_1242_457#_c_1084_n 0.00914718f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_204 VPB N_A_1242_457#_c_1092_n 0.00318329f $X=-0.19 $Y=1.66 $X2=0.2 $Y2=1.265
cc_205 VPB N_A_1242_457#_c_1085_n 0.0102264f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_206 VPB N_A_1242_457#_c_1086_n 0.0107635f $X=-0.19 $Y=1.66 $X2=0.975 $Y2=1.1
cc_207 VPB N_A_1242_457#_c_1095_n 0.00159706f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_208 VPB N_A_855_368#_c_1202_n 0.0225132f $X=-0.19 $Y=1.66 $X2=1.41 $Y2=1.01
cc_209 VPB N_A_855_368#_c_1205_n 0.0769332f $X=-0.19 $Y=1.66 $X2=0.28 $Y2=0.58
cc_210 VPB N_A_855_368#_c_1219_n 0.0560362f $X=-0.19 $Y=1.66 $X2=0.2 $Y2=2.005
cc_211 VPB N_A_855_368#_c_1220_n 0.0123764f $X=-0.19 $Y=1.66 $X2=0.28 $Y2=2.175
cc_212 VPB N_A_855_368#_c_1221_n 0.00717482f $X=-0.19 $Y=1.66 $X2=0.975 $Y2=1.1
cc_213 VPB N_A_855_368#_c_1222_n 0.0193529f $X=-0.19 $Y=1.66 $X2=0.975 $Y2=1.1
cc_214 VPB N_A_855_368#_c_1223_n 0.0133882f $X=-0.19 $Y=1.66 $X2=0.975 $Y2=1.1
cc_215 VPB N_A_855_368#_c_1224_n 0.189544f $X=-0.19 $Y=1.66 $X2=0.445 $Y2=2.09
cc_216 VPB N_A_855_368#_M1025_g 0.010423f $X=-0.19 $Y=1.66 $X2=2.54 $Y2=1.995
cc_217 VPB N_A_855_368#_c_1208_n 0.03645f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_218 VPB N_A_855_368#_c_1227_n 0.0129219f $X=-0.19 $Y=1.66 $X2=2.54 $Y2=2.09
cc_219 VPB N_A_855_368#_c_1228_n 0.0089867f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_220 VPB N_A_855_368#_c_1229_n 0.0289165f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_221 VPB N_A_855_368#_c_1230_n 0.00228081f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_222 VPB N_A_855_368#_c_1215_n 0.00277049f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_223 VPB N_A_855_368#_c_1232_n 0.00185952f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_224 VPB N_A_2082_446#_c_1408_n 0.0165865f $X=-0.19 $Y=1.66 $X2=1.41 $Y2=1.01
cc_225 VPB N_A_2082_446#_c_1409_n 0.0276144f $X=-0.19 $Y=1.66 $X2=2.495 $Y2=2.64
cc_226 VPB N_A_2082_446#_c_1400_n 0.0447354f $X=-0.19 $Y=1.66 $X2=0.2 $Y2=1.265
cc_227 VPB N_A_2082_446#_c_1401_n 0.0137444f $X=-0.19 $Y=1.66 $X2=0.2 $Y2=2.005
cc_228 VPB N_A_2082_446#_c_1412_n 0.00779622f $X=-0.19 $Y=1.66 $X2=0.28
+ $Y2=2.465
cc_229 VPB N_A_2082_446#_c_1413_n 0.00256678f $X=-0.19 $Y=1.66 $X2=0.975 $Y2=1.1
cc_230 VPB N_A_1824_74#_c_1535_n 0.00554553f $X=-0.19 $Y=1.66 $X2=1.485
+ $Y2=0.615
cc_231 VPB N_A_1824_74#_c_1536_n 0.0382574f $X=-0.19 $Y=1.66 $X2=2.495 $Y2=2.245
cc_232 VPB N_A_1824_74#_c_1537_n 0.0224017f $X=-0.19 $Y=1.66 $X2=2.495 $Y2=2.64
cc_233 VPB N_A_1824_74#_c_1524_n 0.00845967f $X=-0.19 $Y=1.66 $X2=0.28 $Y2=2.175
cc_234 VPB N_A_1824_74#_c_1539_n 0.0253471f $X=-0.19 $Y=1.66 $X2=0.28 $Y2=2.465
cc_235 VPB N_A_1824_74#_c_1540_n 0.0061417f $X=-0.19 $Y=1.66 $X2=2.54 $Y2=2.09
cc_236 VPB N_A_1824_74#_c_1541_n 0.00281397f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_237 VPB N_A_1824_74#_c_1530_n 0.0144635f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_238 VPB N_A_2492_392#_c_1672_n 0.0177177f $X=-0.19 $Y=1.66 $X2=1.41 $Y2=1.01
cc_239 VPB N_A_2492_392#_c_1673_n 0.0174134f $X=-0.19 $Y=1.66 $X2=2.495 $Y2=2.64
cc_240 VPB N_A_2492_392#_c_1674_n 0.00506653f $X=-0.19 $Y=1.66 $X2=0.28
+ $Y2=2.465
cc_241 VPB N_A_2492_392#_c_1675_n 0.0105448f $X=-0.19 $Y=1.66 $X2=0.365 $Y2=1.1
cc_242 VPB N_A_2492_392#_c_1669_n 0.00706142f $X=-0.19 $Y=1.66 $X2=2.54 $Y2=2.09
cc_243 VPB N_A_2492_392#_c_1671_n 0.0176866f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_244 VPB N_VPWR_c_1728_n 0.0066125f $X=-0.19 $Y=1.66 $X2=2.375 $Y2=2.09
cc_245 VPB N_VPWR_c_1729_n 0.00396467f $X=-0.19 $Y=1.66 $X2=2.54 $Y2=1.995
cc_246 VPB N_VPWR_c_1730_n 0.0154251f $X=-0.19 $Y=1.66 $X2=2.54 $Y2=2.09
cc_247 VPB N_VPWR_c_1731_n 0.0189554f $X=-0.19 $Y=1.66 $X2=0.975 $Y2=1.1
cc_248 VPB N_VPWR_c_1732_n 0.0194601f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_249 VPB N_VPWR_c_1733_n 0.0187962f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_250 VPB N_VPWR_c_1734_n 0.0121909f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_251 VPB N_VPWR_c_1735_n 0.0688105f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_252 VPB N_VPWR_c_1736_n 0.0375576f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_253 VPB N_VPWR_c_1737_n 0.00601668f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_254 VPB N_VPWR_c_1738_n 0.0616623f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_255 VPB N_VPWR_c_1739_n 0.00443527f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_256 VPB N_VPWR_c_1740_n 0.0198404f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_257 VPB N_VPWR_c_1741_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_258 VPB N_VPWR_c_1742_n 0.0191816f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_259 VPB N_VPWR_c_1743_n 0.0457766f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_260 VPB N_VPWR_c_1744_n 0.0206273f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_261 VPB N_VPWR_c_1745_n 0.0534696f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_262 VPB N_VPWR_c_1746_n 0.0206041f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_263 VPB N_VPWR_c_1747_n 0.0174925f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_264 VPB N_VPWR_c_1748_n 0.0312859f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_265 VPB N_VPWR_c_1749_n 0.00614127f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_266 VPB N_VPWR_c_1750_n 0.00436868f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_267 VPB N_VPWR_c_1751_n 0.0232464f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_268 VPB N_VPWR_c_1752_n 0.00614127f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_269 VPB N_VPWR_c_1727_n 0.117523f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_270 VPB N_A_390_81#_c_1906_n 0.00480127f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_271 VPB N_A_390_81#_c_1912_n 0.00940845f $X=-0.19 $Y=1.66 $X2=2.375 $Y2=2.09
cc_272 VPB N_A_390_81#_c_1913_n 0.0124867f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=1.1
cc_273 VPB N_A_390_81#_c_1914_n 0.00122623f $X=-0.19 $Y=1.66 $X2=0.28 $Y2=2.09
cc_274 VPB N_A_390_81#_c_1915_n 0.00158904f $X=-0.19 $Y=1.66 $X2=2.54 $Y2=2.09
cc_275 VPB N_A_390_81#_c_1910_n 0.00505466f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_276 VPB N_A_390_81#_c_1917_n 0.00257025f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_277 VPB N_A_390_81#_c_1918_n 0.00869982f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_278 VPB N_Q_c_2057_n 0.00395156f $X=-0.19 $Y=1.66 $X2=1.485 $Y2=0.935
cc_279 N_A_27_74#_c_290_n N_SCE_c_369_n 0.0121883f $X=2.375 $Y=2.09 $X2=0 $Y2=0
cc_280 N_A_27_74#_c_291_n N_SCE_c_369_n 0.00496169f $X=0.28 $Y=2.09 $X2=0 $Y2=0
cc_281 N_A_27_74#_c_282_n N_SCE_M1039_g 0.00686809f $X=0.28 $Y=0.58 $X2=0 $Y2=0
cc_282 N_A_27_74#_c_283_n N_SCE_M1039_g 0.00830473f $X=0.2 $Y=2.005 $X2=0 $Y2=0
cc_283 N_A_27_74#_c_284_n N_SCE_M1039_g 0.0281157f $X=0.975 $Y=1.1 $X2=0 $Y2=0
cc_284 N_A_27_74#_c_286_n N_SCE_M1039_g 0.0181297f $X=0.975 $Y=1.01 $X2=0 $Y2=0
cc_285 N_A_27_74#_c_289_n N_SCE_c_370_n 0.0173713f $X=0.28 $Y=2.465 $X2=0 $Y2=0
cc_286 N_A_27_74#_c_290_n N_SCE_c_370_n 0.00721429f $X=2.375 $Y=2.09 $X2=0 $Y2=0
cc_287 N_A_27_74#_c_291_n N_SCE_c_370_n 4.59028e-19 $X=0.28 $Y=2.09 $X2=0 $Y2=0
cc_288 N_A_27_74#_c_290_n N_SCE_c_371_n 0.0100663f $X=2.375 $Y=2.09 $X2=0 $Y2=0
cc_289 N_A_27_74#_c_290_n N_SCE_c_372_n 0.00784761f $X=2.375 $Y=2.09 $X2=0 $Y2=0
cc_290 N_A_27_74#_c_283_n N_SCE_c_362_n 0.0158921f $X=0.2 $Y=2.005 $X2=0 $Y2=0
cc_291 N_A_27_74#_c_284_n N_SCE_c_362_n 0.00162366f $X=0.975 $Y=1.1 $X2=0 $Y2=0
cc_292 N_A_27_74#_c_280_n N_SCE_c_363_n 0.0106974f $X=1.41 $Y=1.01 $X2=0 $Y2=0
cc_293 N_A_27_74#_c_284_n N_SCE_c_363_n 0.00180358f $X=0.975 $Y=1.1 $X2=0 $Y2=0
cc_294 N_A_27_74#_c_290_n N_SCE_c_363_n 0.0170396f $X=2.375 $Y=2.09 $X2=0 $Y2=0
cc_295 N_A_27_74#_c_286_n N_SCE_c_363_n 0.0175645f $X=0.975 $Y=1.01 $X2=0 $Y2=0
cc_296 N_A_27_74#_c_290_n N_SCE_c_364_n 0.0253562f $X=2.375 $Y=2.09 $X2=0 $Y2=0
cc_297 N_A_27_74#_c_287_n N_SCE_c_365_n 0.00114249f $X=2.495 $Y=2.245 $X2=0
+ $Y2=0
cc_298 N_A_27_74#_c_292_n N_SCE_c_365_n 0.0267028f $X=2.54 $Y=1.995 $X2=0 $Y2=0
cc_299 N_A_27_74#_c_287_n N_SCE_c_366_n 0.0182385f $X=2.495 $Y=2.245 $X2=0 $Y2=0
cc_300 N_A_27_74#_c_292_n N_SCE_c_366_n 3.6101e-19 $X=2.54 $Y=1.995 $X2=0 $Y2=0
cc_301 N_A_27_74#_c_280_n N_SCE_c_367_n 0.00818136f $X=1.41 $Y=1.01 $X2=0 $Y2=0
cc_302 N_A_27_74#_c_283_n N_SCE_c_367_n 0.0170838f $X=0.2 $Y=2.005 $X2=0 $Y2=0
cc_303 N_A_27_74#_c_284_n N_SCE_c_367_n 0.0353374f $X=0.975 $Y=1.1 $X2=0 $Y2=0
cc_304 N_A_27_74#_c_290_n N_SCE_c_367_n 0.0893268f $X=2.375 $Y=2.09 $X2=0 $Y2=0
cc_305 N_A_27_74#_c_286_n N_SCE_c_367_n 0.00202099f $X=0.975 $Y=1.01 $X2=0 $Y2=0
cc_306 N_A_27_74#_c_281_n N_D_c_444_n 0.0356736f $X=1.485 $Y=0.935 $X2=-0.19
+ $Y2=-0.245
cc_307 N_A_27_74#_c_287_n N_D_c_445_n 0.0183644f $X=2.495 $Y=2.245 $X2=0 $Y2=0
cc_308 N_A_27_74#_c_290_n N_D_c_445_n 0.00915555f $X=2.375 $Y=2.09 $X2=0 $Y2=0
cc_309 N_A_27_74#_c_292_n N_D_c_445_n 0.00125897f $X=2.54 $Y=1.995 $X2=0 $Y2=0
cc_310 N_A_27_74#_c_287_n N_D_c_449_n 0.0140909f $X=2.495 $Y=2.245 $X2=0 $Y2=0
cc_311 N_A_27_74#_c_290_n N_D_c_449_n 0.00753583f $X=2.375 $Y=2.09 $X2=0 $Y2=0
cc_312 N_A_27_74#_c_281_n N_D_c_446_n 0.00558783f $X=1.485 $Y=0.935 $X2=0 $Y2=0
cc_313 N_A_27_74#_c_284_n N_D_c_446_n 0.0143876f $X=0.975 $Y=1.1 $X2=0 $Y2=0
cc_314 N_A_27_74#_c_286_n N_D_c_446_n 8.79717e-19 $X=0.975 $Y=1.01 $X2=0 $Y2=0
cc_315 N_A_27_74#_c_280_n N_D_c_447_n 0.00979811f $X=1.41 $Y=1.01 $X2=0 $Y2=0
cc_316 N_A_27_74#_c_284_n N_D_c_447_n 2.46751e-19 $X=0.975 $Y=1.1 $X2=0 $Y2=0
cc_317 N_A_27_74#_c_286_n N_D_c_447_n 0.00223479f $X=0.975 $Y=1.01 $X2=0 $Y2=0
cc_318 N_A_27_74#_c_287_n N_SCD_c_493_n 0.0258628f $X=2.495 $Y=2.245 $X2=-0.19
+ $Y2=-0.245
cc_319 N_A_27_74#_c_287_n N_SCD_c_490_n 0.0204601f $X=2.495 $Y=2.245 $X2=0 $Y2=0
cc_320 N_A_27_74#_c_292_n N_SCD_c_490_n 0.001579f $X=2.54 $Y=1.995 $X2=0 $Y2=0
cc_321 N_A_27_74#_c_287_n SCD 0.00117743f $X=2.495 $Y=2.245 $X2=0 $Y2=0
cc_322 N_A_27_74#_c_292_n SCD 0.0182021f $X=2.54 $Y=1.995 $X2=0 $Y2=0
cc_323 N_A_27_74#_c_287_n N_VPWR_c_1728_n 0.00141778f $X=2.495 $Y=2.245 $X2=0
+ $Y2=0
cc_324 N_A_27_74#_c_289_n N_VPWR_c_1742_n 0.0145938f $X=0.28 $Y=2.465 $X2=0
+ $Y2=0
cc_325 N_A_27_74#_c_287_n N_VPWR_c_1743_n 0.00445602f $X=2.495 $Y=2.245 $X2=0
+ $Y2=0
cc_326 N_A_27_74#_c_289_n N_VPWR_c_1748_n 0.0247088f $X=0.28 $Y=2.465 $X2=0
+ $Y2=0
cc_327 N_A_27_74#_c_290_n N_VPWR_c_1748_n 0.0746993f $X=2.375 $Y=2.09 $X2=0
+ $Y2=0
cc_328 N_A_27_74#_c_287_n N_VPWR_c_1727_n 0.00448781f $X=2.495 $Y=2.245 $X2=0
+ $Y2=0
cc_329 N_A_27_74#_c_289_n N_VPWR_c_1727_n 0.0120466f $X=0.28 $Y=2.465 $X2=0
+ $Y2=0
cc_330 N_A_27_74#_c_287_n N_A_390_81#_c_1919_n 0.010208f $X=2.495 $Y=2.245 $X2=0
+ $Y2=0
cc_331 N_A_27_74#_c_292_n N_A_390_81#_c_1919_n 0.0180834f $X=2.54 $Y=1.995 $X2=0
+ $Y2=0
cc_332 N_A_27_74#_c_287_n N_A_390_81#_c_1917_n 0.00974144f $X=2.495 $Y=2.245
+ $X2=0 $Y2=0
cc_333 N_A_27_74#_c_290_n N_A_390_81#_c_1917_n 0.0189432f $X=2.375 $Y=2.09 $X2=0
+ $Y2=0
cc_334 N_A_27_74#_c_292_n N_A_390_81#_c_1917_n 0.00295889f $X=2.54 $Y=1.995
+ $X2=0 $Y2=0
cc_335 N_A_27_74#_c_281_n N_VGND_c_2078_n 0.00287309f $X=1.485 $Y=0.935 $X2=0
+ $Y2=0
cc_336 N_A_27_74#_c_282_n N_VGND_c_2078_n 0.0156021f $X=0.28 $Y=0.58 $X2=0 $Y2=0
cc_337 N_A_27_74#_c_284_n N_VGND_c_2078_n 0.0254818f $X=0.975 $Y=1.1 $X2=0 $Y2=0
cc_338 N_A_27_74#_c_286_n N_VGND_c_2078_n 0.00149092f $X=0.975 $Y=1.01 $X2=0
+ $Y2=0
cc_339 N_A_27_74#_c_281_n N_VGND_c_2086_n 9.09582e-19 $X=1.485 $Y=0.935 $X2=0
+ $Y2=0
cc_340 N_A_27_74#_c_282_n N_VGND_c_2088_n 0.011066f $X=0.28 $Y=0.58 $X2=0 $Y2=0
cc_341 N_A_27_74#_c_282_n N_VGND_c_2100_n 0.00915947f $X=0.28 $Y=0.58 $X2=0
+ $Y2=0
cc_342 N_A_27_74#_c_281_n N_noxref_24_c_2215_n 0.0108727f $X=1.485 $Y=0.935
+ $X2=0 $Y2=0
cc_343 N_A_27_74#_c_281_n N_noxref_24_c_2217_n 0.00859442f $X=1.485 $Y=0.935
+ $X2=0 $Y2=0
cc_344 N_A_27_74#_c_284_n N_noxref_24_c_2217_n 0.00178881f $X=0.975 $Y=1.1 $X2=0
+ $Y2=0
cc_345 N_A_27_74#_c_286_n N_noxref_24_c_2217_n 0.00859402f $X=0.975 $Y=1.01
+ $X2=0 $Y2=0
cc_346 N_SCE_M1006_g N_D_c_444_n 0.00721309f $X=2.66 $Y=0.615 $X2=-0.19
+ $Y2=-0.245
cc_347 N_SCE_c_363_n N_D_c_445_n 0.0203026f $X=1.535 $Y=1.67 $X2=0 $Y2=0
cc_348 N_SCE_c_364_n N_D_c_445_n 0.0144918f $X=2.375 $Y=1.575 $X2=0 $Y2=0
cc_349 N_SCE_c_365_n N_D_c_445_n 3.41462e-19 $X=2.54 $Y=1.425 $X2=0 $Y2=0
cc_350 N_SCE_c_368_n N_D_c_445_n 0.00479409f $X=1.795 $Y=1.662 $X2=0 $Y2=0
cc_351 N_SCE_c_371_n N_D_c_449_n 0.0203026f $X=1.625 $Y=2.155 $X2=0 $Y2=0
cc_352 N_SCE_c_372_n N_D_c_449_n 0.0373591f $X=1.625 $Y=2.245 $X2=0 $Y2=0
cc_353 N_SCE_M1006_g N_D_c_446_n 0.0035822f $X=2.66 $Y=0.615 $X2=0 $Y2=0
cc_354 N_SCE_c_363_n N_D_c_446_n 0.00106377f $X=1.535 $Y=1.67 $X2=0 $Y2=0
cc_355 N_SCE_c_367_n N_D_c_446_n 0.0344941f $X=1.623 $Y=1.662 $X2=0 $Y2=0
cc_356 N_SCE_M1006_g N_D_c_447_n 0.00967695f $X=2.66 $Y=0.615 $X2=0 $Y2=0
cc_357 N_SCE_c_365_n N_D_c_447_n 0.00152136f $X=2.54 $Y=1.425 $X2=0 $Y2=0
cc_358 N_SCE_c_366_n N_D_c_447_n 0.0185773f $X=2.66 $Y=1.425 $X2=0 $Y2=0
cc_359 N_SCE_c_368_n N_D_c_447_n 0.004564f $X=1.795 $Y=1.662 $X2=0 $Y2=0
cc_360 N_SCE_M1006_g N_SCD_M1038_g 0.0638139f $X=2.66 $Y=0.615 $X2=0 $Y2=0
cc_361 N_SCE_c_365_n N_SCD_M1038_g 0.00107576f $X=2.54 $Y=1.425 $X2=0 $Y2=0
cc_362 N_SCE_c_365_n SCD 0.0105222f $X=2.54 $Y=1.425 $X2=0 $Y2=0
cc_363 N_SCE_c_366_n SCD 3.98419e-19 $X=2.66 $Y=1.425 $X2=0 $Y2=0
cc_364 N_SCE_c_365_n N_SCD_c_492_n 0.0018749f $X=2.54 $Y=1.425 $X2=0 $Y2=0
cc_365 N_SCE_c_366_n N_SCD_c_492_n 0.0067837f $X=2.66 $Y=1.425 $X2=0 $Y2=0
cc_366 N_SCE_c_370_n N_VPWR_c_1742_n 0.00445602f $X=0.505 $Y=2.245 $X2=0 $Y2=0
cc_367 N_SCE_c_372_n N_VPWR_c_1743_n 0.00415318f $X=1.625 $Y=2.245 $X2=0 $Y2=0
cc_368 N_SCE_c_370_n N_VPWR_c_1748_n 0.017697f $X=0.505 $Y=2.245 $X2=0 $Y2=0
cc_369 N_SCE_c_372_n N_VPWR_c_1748_n 0.0163904f $X=1.625 $Y=2.245 $X2=0 $Y2=0
cc_370 N_SCE_c_370_n N_VPWR_c_1727_n 0.00865213f $X=0.505 $Y=2.245 $X2=0 $Y2=0
cc_371 N_SCE_c_372_n N_VPWR_c_1727_n 0.00817532f $X=1.625 $Y=2.245 $X2=0 $Y2=0
cc_372 N_SCE_M1006_g N_A_390_81#_c_1902_n 0.0124804f $X=2.66 $Y=0.615 $X2=0
+ $Y2=0
cc_373 N_SCE_c_364_n N_A_390_81#_c_1902_n 0.00321433f $X=2.375 $Y=1.575 $X2=0
+ $Y2=0
cc_374 N_SCE_c_365_n N_A_390_81#_c_1902_n 0.0127797f $X=2.54 $Y=1.425 $X2=0
+ $Y2=0
cc_375 N_SCE_c_366_n N_A_390_81#_c_1902_n 0.00126581f $X=2.66 $Y=1.425 $X2=0
+ $Y2=0
cc_376 N_SCE_M1006_g N_A_390_81#_c_1903_n 0.00615828f $X=2.66 $Y=0.615 $X2=0
+ $Y2=0
cc_377 N_SCE_M1006_g N_A_390_81#_c_1905_n 0.00371736f $X=2.66 $Y=0.615 $X2=0
+ $Y2=0
cc_378 N_SCE_c_365_n N_A_390_81#_c_1905_n 0.00421648f $X=2.54 $Y=1.425 $X2=0
+ $Y2=0
cc_379 N_SCE_c_372_n N_A_390_81#_c_1917_n 0.00182961f $X=1.625 $Y=2.245 $X2=0
+ $Y2=0
cc_380 N_SCE_M1039_g N_VGND_c_2078_n 0.0129468f $X=0.495 $Y=0.58 $X2=0 $Y2=0
cc_381 N_SCE_M1006_g N_VGND_c_2086_n 9.15902e-19 $X=2.66 $Y=0.615 $X2=0 $Y2=0
cc_382 N_SCE_M1039_g N_VGND_c_2088_n 0.00383152f $X=0.495 $Y=0.58 $X2=0 $Y2=0
cc_383 N_SCE_M1039_g N_VGND_c_2100_n 0.00761198f $X=0.495 $Y=0.58 $X2=0 $Y2=0
cc_384 N_SCE_M1006_g N_noxref_24_c_2215_n 0.0107628f $X=2.66 $Y=0.615 $X2=0
+ $Y2=0
cc_385 N_SCE_M1039_g N_noxref_24_c_2217_n 9.19966e-19 $X=0.495 $Y=0.58 $X2=0
+ $Y2=0
cc_386 N_D_c_449_n N_VPWR_c_1743_n 0.00445602f $X=2.045 $Y=2.245 $X2=0 $Y2=0
cc_387 N_D_c_449_n N_VPWR_c_1748_n 0.00236192f $X=2.045 $Y=2.245 $X2=0 $Y2=0
cc_388 N_D_c_449_n N_VPWR_c_1727_n 0.00858241f $X=2.045 $Y=2.245 $X2=0 $Y2=0
cc_389 N_D_c_446_n N_A_390_81#_M1011_d 0.00160203f $X=1.935 $Y=1.1 $X2=-0.19
+ $Y2=-0.245
cc_390 N_D_c_444_n N_A_390_81#_c_1902_n 0.00564096f $X=1.875 $Y=0.935 $X2=0
+ $Y2=0
cc_391 N_D_c_446_n N_A_390_81#_c_1902_n 0.00298881f $X=1.935 $Y=1.1 $X2=0 $Y2=0
cc_392 N_D_c_449_n N_A_390_81#_c_1917_n 0.0112736f $X=2.045 $Y=2.245 $X2=0 $Y2=0
cc_393 N_D_c_444_n N_VGND_c_2086_n 9.15902e-19 $X=1.875 $Y=0.935 $X2=0 $Y2=0
cc_394 N_D_c_444_n N_noxref_24_c_2215_n 0.0119231f $X=1.875 $Y=0.935 $X2=0 $Y2=0
cc_395 N_D_c_446_n N_noxref_24_c_2215_n 0.0128576f $X=1.935 $Y=1.1 $X2=0 $Y2=0
cc_396 N_D_c_447_n N_noxref_24_c_2215_n 0.00157776f $X=2.045 $Y=1.1 $X2=0 $Y2=0
cc_397 N_D_c_444_n N_noxref_24_c_2217_n 0.00113655f $X=1.875 $Y=0.935 $X2=0
+ $Y2=0
cc_398 N_D_c_446_n noxref_25 0.00198619f $X=1.935 $Y=1.1 $X2=-0.19 $Y2=-0.245
cc_399 N_SCD_M1038_g N_RESET_B_M1002_g 0.0276502f $X=3.05 $Y=0.615 $X2=0 $Y2=0
cc_400 SCD N_RESET_B_M1002_g 3.882e-19 $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_401 N_SCD_c_492_n N_RESET_B_M1002_g 0.0178289f $X=3.11 $Y=1.645 $X2=0 $Y2=0
cc_402 N_SCD_c_493_n N_RESET_B_c_544_n 0.0163026f $X=3.035 $Y=2.245 $X2=0 $Y2=0
cc_403 N_SCD_c_490_n N_RESET_B_c_555_n 0.019443f $X=3.11 $Y=1.985 $X2=0 $Y2=0
cc_404 SCD N_RESET_B_c_555_n 3.50716e-19 $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_405 N_SCD_c_493_n N_VPWR_c_1728_n 0.0100582f $X=3.035 $Y=2.245 $X2=0 $Y2=0
cc_406 N_SCD_c_493_n N_VPWR_c_1743_n 0.00413917f $X=3.035 $Y=2.245 $X2=0 $Y2=0
cc_407 N_SCD_c_493_n N_VPWR_c_1727_n 0.00409681f $X=3.035 $Y=2.245 $X2=0 $Y2=0
cc_408 N_SCD_M1038_g N_A_390_81#_c_1902_n 0.00688594f $X=3.05 $Y=0.615 $X2=0
+ $Y2=0
cc_409 N_SCD_c_493_n N_A_390_81#_c_1919_n 0.0130079f $X=3.035 $Y=2.245 $X2=0
+ $Y2=0
cc_410 N_SCD_c_490_n N_A_390_81#_c_1919_n 9.09052e-19 $X=3.11 $Y=1.985 $X2=0
+ $Y2=0
cc_411 SCD N_A_390_81#_c_1919_n 0.02044f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_412 N_SCD_M1038_g N_A_390_81#_c_1903_n 0.00797437f $X=3.05 $Y=0.615 $X2=0
+ $Y2=0
cc_413 N_SCD_M1038_g N_A_390_81#_c_1904_n 0.00837073f $X=3.05 $Y=0.615 $X2=0
+ $Y2=0
cc_414 SCD N_A_390_81#_c_1904_n 0.0179457f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_415 N_SCD_c_492_n N_A_390_81#_c_1904_n 0.00103763f $X=3.11 $Y=1.645 $X2=0
+ $Y2=0
cc_416 N_SCD_M1038_g N_A_390_81#_c_1905_n 0.0030063f $X=3.05 $Y=0.615 $X2=0
+ $Y2=0
cc_417 SCD N_A_390_81#_c_1905_n 0.00853461f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_418 N_SCD_c_492_n N_A_390_81#_c_1905_n 2.26648e-19 $X=3.11 $Y=1.645 $X2=0
+ $Y2=0
cc_419 N_SCD_c_493_n N_A_390_81#_c_1906_n 0.00151656f $X=3.035 $Y=2.245 $X2=0
+ $Y2=0
cc_420 N_SCD_M1038_g N_A_390_81#_c_1906_n 0.00307473f $X=3.05 $Y=0.615 $X2=0
+ $Y2=0
cc_421 N_SCD_c_490_n N_A_390_81#_c_1906_n 0.00173845f $X=3.11 $Y=1.985 $X2=0
+ $Y2=0
cc_422 SCD N_A_390_81#_c_1906_n 0.0502799f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_423 N_SCD_c_492_n N_A_390_81#_c_1906_n 0.00381694f $X=3.11 $Y=1.645 $X2=0
+ $Y2=0
cc_424 N_SCD_c_493_n N_A_390_81#_c_1912_n 4.52461e-19 $X=3.035 $Y=2.245 $X2=0
+ $Y2=0
cc_425 N_SCD_c_493_n N_A_390_81#_c_1914_n 5.56969e-19 $X=3.035 $Y=2.245 $X2=0
+ $Y2=0
cc_426 N_SCD_c_493_n N_A_390_81#_c_1917_n 0.00167919f $X=3.035 $Y=2.245 $X2=0
+ $Y2=0
cc_427 N_SCD_M1038_g N_VGND_c_2086_n 9.15902e-19 $X=3.05 $Y=0.615 $X2=0 $Y2=0
cc_428 N_SCD_M1038_g N_noxref_24_c_2215_n 0.0125096f $X=3.05 $Y=0.615 $X2=0
+ $Y2=0
cc_429 N_SCD_M1038_g N_noxref_24_c_2216_n 0.00668662f $X=3.05 $Y=0.615 $X2=0
+ $Y2=0
cc_430 N_RESET_B_c_550_n N_CLK_c_735_n 0.00217929f $X=8.255 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_431 N_RESET_B_c_555_n N_CLK_c_735_n 0.00390967f $X=3.605 $Y=2.037 $X2=-0.19
+ $Y2=-0.245
cc_432 N_RESET_B_c_556_n N_CLK_c_735_n 4.10166e-19 $X=3.95 $Y=1.995 $X2=-0.19
+ $Y2=-0.245
cc_433 N_RESET_B_M1002_g N_CLK_c_737_n 0.0123949f $X=3.595 $Y=0.615 $X2=0 $Y2=0
cc_434 N_RESET_B_c_550_n N_CLK_c_737_n 0.00236558f $X=8.255 $Y=2.035 $X2=0 $Y2=0
cc_435 N_RESET_B_c_551_n N_CLK_c_737_n 0.00141283f $X=4.225 $Y=2.035 $X2=0 $Y2=0
cc_436 N_RESET_B_c_555_n N_CLK_c_737_n 0.00724732f $X=3.605 $Y=2.037 $X2=0 $Y2=0
cc_437 N_RESET_B_c_556_n N_CLK_c_737_n 0.00160635f $X=3.95 $Y=1.995 $X2=0 $Y2=0
cc_438 N_RESET_B_c_550_n N_CLK_c_748_n 0.00561721f $X=8.255 $Y=2.035 $X2=0 $Y2=0
cc_439 N_RESET_B_M1002_g N_CLK_c_738_n 0.00388719f $X=3.595 $Y=0.615 $X2=0 $Y2=0
cc_440 N_RESET_B_c_551_n N_CLK_c_738_n 0.00358893f $X=4.225 $Y=2.035 $X2=0 $Y2=0
cc_441 N_RESET_B_c_555_n N_CLK_c_738_n 7.34666e-19 $X=3.605 $Y=2.037 $X2=0 $Y2=0
cc_442 N_RESET_B_c_556_n N_CLK_c_738_n 0.0104842f $X=3.95 $Y=1.995 $X2=0 $Y2=0
cc_443 N_RESET_B_c_550_n N_A_1034_368#_c_812_n 0.00524451f $X=8.255 $Y=2.035
+ $X2=0 $Y2=0
cc_444 N_RESET_B_c_550_n N_A_1034_368#_c_790_n 0.0046221f $X=8.255 $Y=2.035
+ $X2=0 $Y2=0
cc_445 N_RESET_B_c_550_n N_A_1034_368#_c_791_n 9.63386e-19 $X=8.255 $Y=2.035
+ $X2=0 $Y2=0
cc_446 N_RESET_B_c_552_n N_A_1034_368#_c_794_n 3.77242e-19 $X=11.135 $Y=2.035
+ $X2=0 $Y2=0
cc_447 N_RESET_B_c_552_n N_A_1034_368#_c_816_n 0.00339815f $X=11.135 $Y=2.035
+ $X2=0 $Y2=0
cc_448 N_RESET_B_c_550_n N_A_1034_368#_c_800_n 0.016155f $X=8.255 $Y=2.035 $X2=0
+ $Y2=0
cc_449 N_RESET_B_c_539_n N_A_1034_368#_c_801_n 0.0116554f $X=7.475 $Y=1.185
+ $X2=0 $Y2=0
cc_450 N_RESET_B_c_552_n N_A_1034_368#_c_807_n 0.0178906f $X=11.135 $Y=2.035
+ $X2=0 $Y2=0
cc_451 N_RESET_B_c_550_n N_A_1034_368#_c_808_n 0.0320515f $X=8.255 $Y=2.035
+ $X2=0 $Y2=0
cc_452 N_RESET_B_c_539_n N_A_1034_368#_c_810_n 5.48446e-19 $X=7.475 $Y=1.185
+ $X2=0 $Y2=0
cc_453 N_RESET_B_c_550_n N_A_1034_368#_c_811_n 0.00546521f $X=8.255 $Y=2.035
+ $X2=0 $Y2=0
cc_454 N_RESET_B_c_552_n N_A_1383_349#_M1016_d 0.00622796f $X=11.135 $Y=2.035
+ $X2=0 $Y2=0
cc_455 N_RESET_B_c_545_n N_A_1383_349#_c_996_n 0.0122885f $X=7.63 $Y=2.21 $X2=0
+ $Y2=0
cc_456 N_RESET_B_c_540_n N_A_1383_349#_c_996_n 0.00263372f $X=7.645 $Y=1.795
+ $X2=0 $Y2=0
cc_457 N_RESET_B_c_550_n N_A_1383_349#_c_996_n 0.0113866f $X=8.255 $Y=2.035
+ $X2=0 $Y2=0
cc_458 N_RESET_B_c_557_n N_A_1383_349#_c_996_n 0.0214958f $X=7.645 $Y=2.002
+ $X2=0 $Y2=0
cc_459 N_RESET_B_c_539_n N_A_1383_349#_M1035_g 0.0418792f $X=7.475 $Y=1.185
+ $X2=0 $Y2=0
cc_460 N_RESET_B_c_540_n N_A_1383_349#_M1035_g 0.0108937f $X=7.645 $Y=1.795
+ $X2=0 $Y2=0
cc_461 N_RESET_B_c_539_n N_A_1383_349#_c_993_n 0.00474717f $X=7.475 $Y=1.185
+ $X2=0 $Y2=0
cc_462 N_RESET_B_c_540_n N_A_1383_349#_c_993_n 0.00131101f $X=7.645 $Y=1.795
+ $X2=0 $Y2=0
cc_463 N_RESET_B_c_550_n N_A_1383_349#_c_993_n 0.0210957f $X=8.255 $Y=2.035
+ $X2=0 $Y2=0
cc_464 N_RESET_B_c_557_n N_A_1383_349#_c_993_n 3.6329e-19 $X=7.645 $Y=2.002
+ $X2=0 $Y2=0
cc_465 N_RESET_B_c_539_n N_A_1383_349#_c_1013_n 0.0144265f $X=7.475 $Y=1.185
+ $X2=0 $Y2=0
cc_466 N_RESET_B_c_542_n N_A_1383_349#_c_1013_n 0.00458767f $X=7.645 $Y=1.26
+ $X2=0 $Y2=0
cc_467 N_RESET_B_c_552_n N_A_1383_349#_c_999_n 0.0436073f $X=11.135 $Y=2.035
+ $X2=0 $Y2=0
cc_468 N_RESET_B_c_553_n N_A_1383_349#_c_999_n 0.00263797f $X=8.545 $Y=2.035
+ $X2=0 $Y2=0
cc_469 N_RESET_B_c_554_n N_A_1383_349#_c_999_n 0.00493501f $X=8.4 $Y=2.035 $X2=0
+ $Y2=0
cc_470 N_RESET_B_c_552_n N_A_1242_457#_c_1083_n 0.0150817f $X=11.135 $Y=2.035
+ $X2=0 $Y2=0
cc_471 N_RESET_B_c_553_n N_A_1242_457#_c_1083_n 0.00261991f $X=8.545 $Y=2.035
+ $X2=0 $Y2=0
cc_472 N_RESET_B_c_554_n N_A_1242_457#_c_1083_n 0.0027848f $X=8.4 $Y=2.035 $X2=0
+ $Y2=0
cc_473 N_RESET_B_c_557_n N_A_1242_457#_c_1083_n 0.00817914f $X=7.645 $Y=2.002
+ $X2=0 $Y2=0
cc_474 N_RESET_B_c_542_n N_A_1242_457#_c_1084_n 0.0105479f $X=7.645 $Y=1.26
+ $X2=0 $Y2=0
cc_475 N_RESET_B_c_554_n N_A_1242_457#_c_1084_n 0.0100815f $X=8.4 $Y=2.035 $X2=0
+ $Y2=0
cc_476 N_RESET_B_c_557_n N_A_1242_457#_c_1084_n 0.00287914f $X=7.645 $Y=2.002
+ $X2=0 $Y2=0
cc_477 N_RESET_B_c_550_n N_A_1242_457#_c_1092_n 0.00732961f $X=8.255 $Y=2.035
+ $X2=0 $Y2=0
cc_478 N_RESET_B_c_550_n N_A_1242_457#_c_1085_n 0.0221124f $X=8.255 $Y=2.035
+ $X2=0 $Y2=0
cc_479 N_RESET_B_c_550_n N_A_1242_457#_c_1105_n 0.0205065f $X=8.255 $Y=2.035
+ $X2=0 $Y2=0
cc_480 N_RESET_B_c_545_n N_A_1242_457#_c_1086_n 0.0185053f $X=7.63 $Y=2.21 $X2=0
+ $Y2=0
cc_481 N_RESET_B_c_540_n N_A_1242_457#_c_1086_n 0.0114947f $X=7.645 $Y=1.795
+ $X2=0 $Y2=0
cc_482 N_RESET_B_c_550_n N_A_1242_457#_c_1086_n 0.0293845f $X=8.255 $Y=2.035
+ $X2=0 $Y2=0
cc_483 N_RESET_B_c_553_n N_A_1242_457#_c_1086_n 2.62119e-19 $X=8.545 $Y=2.035
+ $X2=0 $Y2=0
cc_484 N_RESET_B_c_554_n N_A_1242_457#_c_1086_n 0.0403998f $X=8.4 $Y=2.035 $X2=0
+ $Y2=0
cc_485 N_RESET_B_c_557_n N_A_1242_457#_c_1086_n 0.0179852f $X=7.645 $Y=2.002
+ $X2=0 $Y2=0
cc_486 N_RESET_B_c_540_n N_A_1242_457#_c_1087_n 0.00390473f $X=7.645 $Y=1.795
+ $X2=0 $Y2=0
cc_487 N_RESET_B_c_542_n N_A_1242_457#_c_1087_n 0.00529036f $X=7.645 $Y=1.26
+ $X2=0 $Y2=0
cc_488 N_RESET_B_c_540_n N_A_1242_457#_c_1088_n 0.00623197f $X=7.645 $Y=1.795
+ $X2=0 $Y2=0
cc_489 N_RESET_B_c_542_n N_A_1242_457#_c_1088_n 0.00198801f $X=7.645 $Y=1.26
+ $X2=0 $Y2=0
cc_490 N_RESET_B_c_550_n N_A_1242_457#_c_1088_n 0.0080909f $X=8.255 $Y=2.035
+ $X2=0 $Y2=0
cc_491 N_RESET_B_c_553_n N_A_1242_457#_c_1088_n 8.96068e-19 $X=8.545 $Y=2.035
+ $X2=0 $Y2=0
cc_492 N_RESET_B_c_554_n N_A_1242_457#_c_1088_n 0.0351039f $X=8.4 $Y=2.035 $X2=0
+ $Y2=0
cc_493 N_RESET_B_c_557_n N_A_1242_457#_c_1088_n 0.0100276f $X=7.645 $Y=2.002
+ $X2=0 $Y2=0
cc_494 N_RESET_B_c_550_n N_A_855_368#_M1018_s 0.0011702f $X=8.255 $Y=2.035 $X2=0
+ $Y2=0
cc_495 N_RESET_B_c_550_n N_A_855_368#_c_1202_n 0.00465858f $X=8.255 $Y=2.035
+ $X2=0 $Y2=0
cc_496 N_RESET_B_c_550_n N_A_855_368#_c_1205_n 0.00471468f $X=8.255 $Y=2.035
+ $X2=0 $Y2=0
cc_497 N_RESET_B_c_550_n N_A_855_368#_c_1223_n 0.00215571f $X=8.255 $Y=2.035
+ $X2=0 $Y2=0
cc_498 N_RESET_B_c_545_n N_A_855_368#_c_1224_n 0.00859125f $X=7.63 $Y=2.21 $X2=0
+ $Y2=0
cc_499 N_RESET_B_c_552_n N_A_855_368#_M1025_g 0.00944311f $X=11.135 $Y=2.035
+ $X2=0 $Y2=0
cc_500 N_RESET_B_c_552_n N_A_855_368#_c_1208_n 0.00577012f $X=11.135 $Y=2.035
+ $X2=0 $Y2=0
cc_501 N_RESET_B_c_552_n N_A_855_368#_c_1227_n 3.19444e-19 $X=11.135 $Y=2.035
+ $X2=0 $Y2=0
cc_502 N_RESET_B_c_550_n N_A_855_368#_c_1230_n 0.0152754f $X=8.255 $Y=2.035
+ $X2=0 $Y2=0
cc_503 N_RESET_B_M1002_g N_A_855_368#_c_1232_n 2.05047e-19 $X=3.595 $Y=0.615
+ $X2=0 $Y2=0
cc_504 N_RESET_B_c_550_n N_A_855_368#_c_1232_n 0.014404f $X=8.255 $Y=2.035 $X2=0
+ $Y2=0
cc_505 N_RESET_B_c_551_n N_A_855_368#_c_1232_n 0.00277564f $X=4.225 $Y=2.035
+ $X2=0 $Y2=0
cc_506 N_RESET_B_c_555_n N_A_855_368#_c_1232_n 0.0023658f $X=3.605 $Y=2.037
+ $X2=0 $Y2=0
cc_507 N_RESET_B_c_556_n N_A_855_368#_c_1232_n 0.0240037f $X=3.95 $Y=1.995 $X2=0
+ $Y2=0
cc_508 N_RESET_B_c_550_n N_A_855_368#_c_1216_n 0.00716742f $X=8.255 $Y=2.035
+ $X2=0 $Y2=0
cc_509 N_RESET_B_c_549_n N_A_2082_446#_c_1408_n 0.00549853f $X=11.35 $Y=2.465
+ $X2=0 $Y2=0
cc_510 N_RESET_B_M1023_g N_A_2082_446#_M1009_g 0.0332604f $X=11.135 $Y=0.58
+ $X2=0 $Y2=0
cc_511 N_RESET_B_c_548_n N_A_2082_446#_c_1409_n 0.00482347f $X=11.35 $Y=2.375
+ $X2=0 $Y2=0
cc_512 N_RESET_B_c_549_n N_A_2082_446#_c_1409_n 9.24257e-19 $X=11.35 $Y=2.465
+ $X2=0 $Y2=0
cc_513 N_RESET_B_c_552_n N_A_2082_446#_c_1409_n 7.79989e-19 $X=11.135 $Y=2.035
+ $X2=0 $Y2=0
cc_514 N_RESET_B_c_548_n N_A_2082_446#_c_1419_n 8.40443e-19 $X=11.35 $Y=2.375
+ $X2=0 $Y2=0
cc_515 N_RESET_B_c_552_n N_A_2082_446#_c_1419_n 0.0371304f $X=11.135 $Y=2.035
+ $X2=0 $Y2=0
cc_516 RESET_B N_A_2082_446#_c_1419_n 5.86564e-19 $X=11.195 $Y=1.95 $X2=0 $Y2=0
cc_517 N_RESET_B_c_558_n N_A_2082_446#_c_1419_n 0.00153537f $X=11.275 $Y=2.07
+ $X2=0 $Y2=0
cc_518 N_RESET_B_c_653_p N_A_2082_446#_c_1419_n 0.0134652f $X=11.28 $Y=2.035
+ $X2=0 $Y2=0
cc_519 N_RESET_B_c_552_n N_A_2082_446#_c_1400_n 0.0118555f $X=11.135 $Y=2.035
+ $X2=0 $Y2=0
cc_520 N_RESET_B_c_558_n N_A_2082_446#_c_1400_n 0.031607f $X=11.275 $Y=2.07
+ $X2=0 $Y2=0
cc_521 N_RESET_B_c_653_p N_A_2082_446#_c_1400_n 0.00107974f $X=11.28 $Y=2.035
+ $X2=0 $Y2=0
cc_522 N_RESET_B_M1023_g N_A_2082_446#_c_1401_n 0.0112646f $X=11.135 $Y=0.58
+ $X2=0 $Y2=0
cc_523 N_RESET_B_c_552_n N_A_2082_446#_c_1401_n 0.00766736f $X=11.135 $Y=2.035
+ $X2=0 $Y2=0
cc_524 RESET_B N_A_2082_446#_c_1401_n 0.0021857f $X=11.195 $Y=1.95 $X2=0 $Y2=0
cc_525 N_RESET_B_c_558_n N_A_2082_446#_c_1401_n 0.00565198f $X=11.275 $Y=2.07
+ $X2=0 $Y2=0
cc_526 N_RESET_B_c_653_p N_A_2082_446#_c_1401_n 0.0208148f $X=11.28 $Y=2.035
+ $X2=0 $Y2=0
cc_527 N_RESET_B_c_549_n N_A_2082_446#_c_1412_n 0.0137666f $X=11.35 $Y=2.465
+ $X2=0 $Y2=0
cc_528 N_RESET_B_c_552_n N_A_2082_446#_c_1412_n 0.00726729f $X=11.135 $Y=2.035
+ $X2=0 $Y2=0
cc_529 RESET_B N_A_2082_446#_c_1412_n 0.00176886f $X=11.195 $Y=1.95 $X2=0 $Y2=0
cc_530 N_RESET_B_c_558_n N_A_2082_446#_c_1412_n 0.00469264f $X=11.275 $Y=2.07
+ $X2=0 $Y2=0
cc_531 N_RESET_B_c_653_p N_A_2082_446#_c_1412_n 0.0223172f $X=11.28 $Y=2.035
+ $X2=0 $Y2=0
cc_532 N_RESET_B_c_549_n N_A_2082_446#_c_1413_n 0.0102517f $X=11.35 $Y=2.465
+ $X2=0 $Y2=0
cc_533 N_RESET_B_M1023_g N_A_2082_446#_c_1402_n 0.00114233f $X=11.135 $Y=0.58
+ $X2=0 $Y2=0
cc_534 N_RESET_B_M1023_g N_A_2082_446#_c_1404_n 7.54334e-19 $X=11.135 $Y=0.58
+ $X2=0 $Y2=0
cc_535 N_RESET_B_M1023_g N_A_2082_446#_c_1406_n 0.00211977f $X=11.135 $Y=0.58
+ $X2=0 $Y2=0
cc_536 N_RESET_B_M1023_g N_A_2082_446#_c_1407_n 0.0225188f $X=11.135 $Y=0.58
+ $X2=0 $Y2=0
cc_537 N_RESET_B_c_552_n N_A_1824_74#_M1025_d 6.85563e-19 $X=11.135 $Y=2.035
+ $X2=0 $Y2=0
cc_538 N_RESET_B_M1023_g N_A_1824_74#_M1013_g 0.0603983f $X=11.135 $Y=0.58 $X2=0
+ $Y2=0
cc_539 N_RESET_B_M1023_g N_A_1824_74#_c_1535_n 0.00632307f $X=11.135 $Y=0.58
+ $X2=0 $Y2=0
cc_540 N_RESET_B_c_558_n N_A_1824_74#_c_1536_n 0.013294f $X=11.275 $Y=2.07 $X2=0
+ $Y2=0
cc_541 N_RESET_B_c_653_p N_A_1824_74#_c_1536_n 0.00121903f $X=11.28 $Y=2.035
+ $X2=0 $Y2=0
cc_542 N_RESET_B_c_548_n N_A_1824_74#_c_1537_n 0.013294f $X=11.35 $Y=2.375 $X2=0
+ $Y2=0
cc_543 N_RESET_B_c_549_n N_A_1824_74#_c_1537_n 0.00940262f $X=11.35 $Y=2.465
+ $X2=0 $Y2=0
cc_544 N_RESET_B_M1023_g N_A_1824_74#_c_1523_n 0.00629822f $X=11.135 $Y=0.58
+ $X2=0 $Y2=0
cc_545 N_RESET_B_c_558_n N_A_1824_74#_c_1523_n 2.27226e-19 $X=11.275 $Y=2.07
+ $X2=0 $Y2=0
cc_546 N_RESET_B_M1023_g N_A_1824_74#_c_1526_n 0.00585373f $X=11.135 $Y=0.58
+ $X2=0 $Y2=0
cc_547 N_RESET_B_c_552_n N_A_1824_74#_c_1553_n 0.0283424f $X=11.135 $Y=2.035
+ $X2=0 $Y2=0
cc_548 N_RESET_B_c_552_n N_A_1824_74#_c_1540_n 0.0138963f $X=11.135 $Y=2.035
+ $X2=0 $Y2=0
cc_549 N_RESET_B_c_552_n N_A_1824_74#_c_1530_n 0.023417f $X=11.135 $Y=2.035
+ $X2=0 $Y2=0
cc_550 N_RESET_B_M1023_g N_A_1824_74#_c_1531_n 0.00517953f $X=11.135 $Y=0.58
+ $X2=0 $Y2=0
cc_551 N_RESET_B_M1023_g N_A_1824_74#_c_1534_n 0.0159185f $X=11.135 $Y=0.58
+ $X2=0 $Y2=0
cc_552 N_RESET_B_c_550_n N_VPWR_M1018_d 0.00304398f $X=8.255 $Y=2.035 $X2=0
+ $Y2=0
cc_553 N_RESET_B_c_552_n N_VPWR_M1016_s 4.03369e-19 $X=11.135 $Y=2.035 $X2=0
+ $Y2=0
cc_554 N_RESET_B_c_553_n N_VPWR_M1016_s 0.00325449f $X=8.545 $Y=2.035 $X2=0
+ $Y2=0
cc_555 N_RESET_B_c_554_n N_VPWR_M1016_s 0.00690849f $X=8.4 $Y=2.035 $X2=0 $Y2=0
cc_556 N_RESET_B_c_544_n N_VPWR_c_1728_n 0.00548967f $X=3.605 $Y=2.245 $X2=0
+ $Y2=0
cc_557 N_RESET_B_c_545_n N_VPWR_c_1730_n 0.00384546f $X=7.63 $Y=2.21 $X2=0 $Y2=0
cc_558 N_RESET_B_c_545_n N_VPWR_c_1731_n 0.00350108f $X=7.63 $Y=2.21 $X2=0 $Y2=0
cc_559 N_RESET_B_c_552_n N_VPWR_c_1731_n 0.00158286f $X=11.135 $Y=2.035 $X2=0
+ $Y2=0
cc_560 N_RESET_B_c_553_n N_VPWR_c_1731_n 0.00903602f $X=8.545 $Y=2.035 $X2=0
+ $Y2=0
cc_561 N_RESET_B_c_554_n N_VPWR_c_1731_n 0.0187103f $X=8.4 $Y=2.035 $X2=0 $Y2=0
cc_562 RESET_B N_VPWR_c_1732_n 0.00143958f $X=11.195 $Y=1.95 $X2=0 $Y2=0
cc_563 N_RESET_B_c_653_p N_VPWR_c_1732_n 0.00812957f $X=11.28 $Y=2.035 $X2=0
+ $Y2=0
cc_564 N_RESET_B_c_544_n N_VPWR_c_1736_n 0.00388952f $X=3.605 $Y=2.245 $X2=0
+ $Y2=0
cc_565 N_RESET_B_c_549_n N_VPWR_c_1740_n 0.00445602f $X=11.35 $Y=2.465 $X2=0
+ $Y2=0
cc_566 N_RESET_B_c_549_n N_VPWR_c_1751_n 0.00638397f $X=11.35 $Y=2.465 $X2=0
+ $Y2=0
cc_567 N_RESET_B_c_544_n N_VPWR_c_1727_n 0.00420469f $X=3.605 $Y=2.245 $X2=0
+ $Y2=0
cc_568 N_RESET_B_c_545_n N_VPWR_c_1727_n 9.49986e-19 $X=7.63 $Y=2.21 $X2=0 $Y2=0
cc_569 N_RESET_B_c_549_n N_VPWR_c_1727_n 0.00439026f $X=11.35 $Y=2.465 $X2=0
+ $Y2=0
cc_570 N_RESET_B_M1002_g N_A_390_81#_c_1903_n 0.00147981f $X=3.595 $Y=0.615
+ $X2=0 $Y2=0
cc_571 N_RESET_B_M1002_g N_A_390_81#_c_1904_n 0.0113777f $X=3.595 $Y=0.615 $X2=0
+ $Y2=0
cc_572 N_RESET_B_M1002_g N_A_390_81#_c_1906_n 0.019178f $X=3.595 $Y=0.615 $X2=0
+ $Y2=0
cc_573 N_RESET_B_c_544_n N_A_390_81#_c_1906_n 0.00445911f $X=3.605 $Y=2.245
+ $X2=0 $Y2=0
cc_574 N_RESET_B_c_551_n N_A_390_81#_c_1906_n 0.00108729f $X=4.225 $Y=2.035
+ $X2=0 $Y2=0
cc_575 N_RESET_B_c_555_n N_A_390_81#_c_1906_n 0.0139492f $X=3.605 $Y=2.037 $X2=0
+ $Y2=0
cc_576 N_RESET_B_c_556_n N_A_390_81#_c_1906_n 0.0228135f $X=3.95 $Y=1.995 $X2=0
+ $Y2=0
cc_577 N_RESET_B_c_544_n N_A_390_81#_c_1912_n 0.00791994f $X=3.605 $Y=2.245
+ $X2=0 $Y2=0
cc_578 N_RESET_B_c_550_n N_A_390_81#_c_1913_n 0.0290511f $X=8.255 $Y=2.035 $X2=0
+ $Y2=0
cc_579 N_RESET_B_c_551_n N_A_390_81#_c_1913_n 0.00388056f $X=4.225 $Y=2.035
+ $X2=0 $Y2=0
cc_580 N_RESET_B_c_555_n N_A_390_81#_c_1913_n 0.00258186f $X=3.605 $Y=2.037
+ $X2=0 $Y2=0
cc_581 N_RESET_B_c_556_n N_A_390_81#_c_1913_n 0.00903824f $X=3.95 $Y=1.995 $X2=0
+ $Y2=0
cc_582 N_RESET_B_c_544_n N_A_390_81#_c_1914_n 0.0119634f $X=3.605 $Y=2.245 $X2=0
+ $Y2=0
cc_583 N_RESET_B_c_551_n N_A_390_81#_c_1914_n 4.98701e-19 $X=4.225 $Y=2.035
+ $X2=0 $Y2=0
cc_584 N_RESET_B_c_555_n N_A_390_81#_c_1914_n 0.00783424f $X=3.605 $Y=2.037
+ $X2=0 $Y2=0
cc_585 N_RESET_B_c_556_n N_A_390_81#_c_1914_n 0.0168153f $X=3.95 $Y=1.995 $X2=0
+ $Y2=0
cc_586 N_RESET_B_c_550_n N_A_390_81#_c_1915_n 0.0114008f $X=8.255 $Y=2.035 $X2=0
+ $Y2=0
cc_587 N_RESET_B_c_550_n N_A_390_81#_c_1908_n 0.0036393f $X=8.255 $Y=2.035 $X2=0
+ $Y2=0
cc_588 N_RESET_B_c_550_n N_A_390_81#_c_1910_n 0.0156292f $X=8.255 $Y=2.035 $X2=0
+ $Y2=0
cc_589 N_RESET_B_c_550_n N_A_390_81#_c_1918_n 0.00761582f $X=8.255 $Y=2.035
+ $X2=0 $Y2=0
cc_590 N_RESET_B_M1002_g N_VGND_c_2079_n 0.0115263f $X=3.595 $Y=0.615 $X2=0
+ $Y2=0
cc_591 N_RESET_B_M1023_g N_VGND_c_2081_n 0.0122528f $X=11.135 $Y=0.58 $X2=0
+ $Y2=0
cc_592 N_RESET_B_M1002_g N_VGND_c_2086_n 0.0047553f $X=3.595 $Y=0.615 $X2=0
+ $Y2=0
cc_593 N_RESET_B_c_539_n N_VGND_c_2090_n 0.00294166f $X=7.475 $Y=1.185 $X2=0
+ $Y2=0
cc_594 N_RESET_B_M1023_g N_VGND_c_2092_n 0.00383152f $X=11.135 $Y=0.58 $X2=0
+ $Y2=0
cc_595 N_RESET_B_M1002_g N_VGND_c_2100_n 0.00445555f $X=3.595 $Y=0.615 $X2=0
+ $Y2=0
cc_596 N_RESET_B_c_539_n N_VGND_c_2100_n 0.00451834f $X=7.475 $Y=1.185 $X2=0
+ $Y2=0
cc_597 N_RESET_B_M1023_g N_VGND_c_2100_n 0.0075694f $X=11.135 $Y=0.58 $X2=0
+ $Y2=0
cc_598 N_RESET_B_M1002_g N_noxref_24_c_2215_n 0.00417413f $X=3.595 $Y=0.615
+ $X2=0 $Y2=0
cc_599 N_RESET_B_M1002_g N_noxref_24_c_2216_n 0.00538329f $X=3.595 $Y=0.615
+ $X2=0 $Y2=0
cc_600 N_CLK_M1019_g N_A_1034_368#_c_796_n 9.99563e-19 $X=4.69 $Y=0.74 $X2=0
+ $Y2=0
cc_601 N_CLK_c_735_n N_A_1034_368#_c_808_n 8.48532e-19 $X=4.645 $Y=1.765 $X2=0
+ $Y2=0
cc_602 N_CLK_c_735_n N_A_855_368#_c_1202_n 0.0481718f $X=4.645 $Y=1.765 $X2=0
+ $Y2=0
cc_603 N_CLK_M1019_g N_A_855_368#_c_1202_n 0.0224827f $X=4.69 $Y=0.74 $X2=0
+ $Y2=0
cc_604 N_CLK_c_748_n N_A_855_368#_c_1202_n 2.48882e-19 $X=4.48 $Y=1.425 $X2=0
+ $Y2=0
cc_605 N_CLK_M1019_g N_A_855_368#_M1007_g 0.0230598f $X=4.69 $Y=0.74 $X2=0 $Y2=0
cc_606 N_CLK_M1019_g N_A_855_368#_c_1213_n 8.21824e-19 $X=4.69 $Y=0.74 $X2=0
+ $Y2=0
cc_607 N_CLK_M1019_g N_A_855_368#_c_1253_n 0.015589f $X=4.69 $Y=0.74 $X2=0 $Y2=0
cc_608 N_CLK_c_748_n N_A_855_368#_c_1253_n 0.00417222f $X=4.48 $Y=1.425 $X2=0
+ $Y2=0
cc_609 N_CLK_c_737_n N_A_855_368#_c_1255_n 0.00394119f $X=4.555 $Y=1.425 $X2=0
+ $Y2=0
cc_610 N_CLK_c_748_n N_A_855_368#_c_1255_n 0.0138664f $X=4.48 $Y=1.425 $X2=0
+ $Y2=0
cc_611 N_CLK_c_735_n N_A_855_368#_c_1230_n 0.0125528f $X=4.645 $Y=1.765 $X2=0
+ $Y2=0
cc_612 N_CLK_c_748_n N_A_855_368#_c_1230_n 0.00302347f $X=4.48 $Y=1.425 $X2=0
+ $Y2=0
cc_613 N_CLK_M1019_g N_A_855_368#_c_1214_n 0.00317215f $X=4.69 $Y=0.74 $X2=0
+ $Y2=0
cc_614 N_CLK_c_748_n N_A_855_368#_c_1214_n 0.00271679f $X=4.48 $Y=1.425 $X2=0
+ $Y2=0
cc_615 N_CLK_c_738_n N_A_855_368#_c_1214_n 0.00245197f $X=4.195 $Y=1.385 $X2=0
+ $Y2=0
cc_616 N_CLK_c_735_n N_A_855_368#_c_1215_n 0.00448074f $X=4.645 $Y=1.765 $X2=0
+ $Y2=0
cc_617 N_CLK_c_735_n N_A_855_368#_c_1232_n 0.00541631f $X=4.645 $Y=1.765 $X2=0
+ $Y2=0
cc_618 N_CLK_c_737_n N_A_855_368#_c_1232_n 0.004824f $X=4.555 $Y=1.425 $X2=0
+ $Y2=0
cc_619 N_CLK_c_748_n N_A_855_368#_c_1232_n 0.0144756f $X=4.48 $Y=1.425 $X2=0
+ $Y2=0
cc_620 N_CLK_c_735_n N_A_855_368#_c_1216_n 0.00340618f $X=4.645 $Y=1.765 $X2=0
+ $Y2=0
cc_621 N_CLK_c_748_n N_A_855_368#_c_1216_n 0.0254591f $X=4.48 $Y=1.425 $X2=0
+ $Y2=0
cc_622 N_CLK_c_735_n N_VPWR_c_1729_n 0.0172823f $X=4.645 $Y=1.765 $X2=0 $Y2=0
cc_623 N_CLK_c_735_n N_VPWR_c_1736_n 0.00413917f $X=4.645 $Y=1.765 $X2=0 $Y2=0
cc_624 N_CLK_c_735_n N_VPWR_c_1727_n 0.00403443f $X=4.645 $Y=1.765 $X2=0 $Y2=0
cc_625 N_CLK_c_738_n N_A_390_81#_c_1904_n 0.00635568f $X=4.195 $Y=1.385 $X2=0
+ $Y2=0
cc_626 N_CLK_c_737_n N_A_390_81#_c_1906_n 3.23617e-19 $X=4.555 $Y=1.425 $X2=0
+ $Y2=0
cc_627 N_CLK_c_738_n N_A_390_81#_c_1906_n 0.0131632f $X=4.195 $Y=1.385 $X2=0
+ $Y2=0
cc_628 N_CLK_c_735_n N_A_390_81#_c_1912_n 0.0103912f $X=4.645 $Y=1.765 $X2=0
+ $Y2=0
cc_629 N_CLK_c_735_n N_A_390_81#_c_1913_n 0.0146064f $X=4.645 $Y=1.765 $X2=0
+ $Y2=0
cc_630 N_CLK_c_735_n N_A_390_81#_c_1914_n 0.00160388f $X=4.645 $Y=1.765 $X2=0
+ $Y2=0
cc_631 N_CLK_M1019_g N_VGND_c_2079_n 0.0038126f $X=4.69 $Y=0.74 $X2=0 $Y2=0
cc_632 N_CLK_c_737_n N_VGND_c_2079_n 4.3166e-19 $X=4.555 $Y=1.425 $X2=0 $Y2=0
cc_633 N_CLK_c_738_n N_VGND_c_2079_n 0.00442933f $X=4.195 $Y=1.385 $X2=0 $Y2=0
cc_634 N_CLK_M1019_g N_VGND_c_2080_n 0.0114836f $X=4.69 $Y=0.74 $X2=0 $Y2=0
cc_635 N_CLK_M1019_g N_VGND_c_2089_n 0.00383152f $X=4.69 $Y=0.74 $X2=0 $Y2=0
cc_636 N_CLK_M1019_g N_VGND_c_2100_n 0.00762539f $X=4.69 $Y=0.74 $X2=0 $Y2=0
cc_637 N_A_1034_368#_c_802_n N_A_1383_349#_M1040_d 0.00256188f $X=9.09 $Y=0.34
+ $X2=-0.19 $Y2=-0.245
cc_638 N_A_1034_368#_c_812_n N_A_1383_349#_c_996_n 0.00260777f $X=6.135 $Y=2.12
+ $X2=0 $Y2=0
cc_639 N_A_1034_368#_c_791_n N_A_1383_349#_c_996_n 0.00193915f $X=6.695 $Y=1.355
+ $X2=0 $Y2=0
cc_640 N_A_1034_368#_c_811_n N_A_1383_349#_c_996_n 0.00175484f $X=6.065 $Y=1.71
+ $X2=0 $Y2=0
cc_641 N_A_1034_368#_c_791_n N_A_1383_349#_M1035_g 0.00646846f $X=6.695 $Y=1.355
+ $X2=0 $Y2=0
cc_642 N_A_1034_368#_M1003_g N_A_1383_349#_M1035_g 0.0474823f $X=6.695 $Y=0.9
+ $X2=0 $Y2=0
cc_643 N_A_1034_368#_c_798_n N_A_1383_349#_M1035_g 0.00140384f $X=7.04 $Y=0.415
+ $X2=0 $Y2=0
cc_644 N_A_1034_368#_c_801_n N_A_1383_349#_M1035_g 3.08289e-19 $X=8.25 $Y=0.665
+ $X2=0 $Y2=0
cc_645 N_A_1034_368#_c_810_n N_A_1383_349#_M1035_g 0.00894962f $X=7.125 $Y=0.415
+ $X2=0 $Y2=0
cc_646 N_A_1034_368#_M1003_g N_A_1383_349#_c_993_n 4.19676e-19 $X=6.695 $Y=0.9
+ $X2=0 $Y2=0
cc_647 N_A_1034_368#_c_801_n N_A_1383_349#_c_1013_n 0.0713598f $X=8.25 $Y=0.665
+ $X2=0 $Y2=0
cc_648 N_A_1034_368#_c_802_n N_A_1383_349#_c_1013_n 0.00354657f $X=9.09 $Y=0.34
+ $X2=0 $Y2=0
cc_649 N_A_1034_368#_M1003_g N_A_1383_349#_c_1030_n 2.50187e-19 $X=6.695 $Y=0.9
+ $X2=0 $Y2=0
cc_650 N_A_1034_368#_c_801_n N_A_1383_349#_c_1030_n 0.00797314f $X=8.25 $Y=0.665
+ $X2=0 $Y2=0
cc_651 N_A_1034_368#_c_810_n N_A_1383_349#_c_1030_n 0.00971736f $X=7.125
+ $Y=0.415 $X2=0 $Y2=0
cc_652 N_A_1034_368#_c_793_n N_A_1383_349#_c_994_n 0.00241408f $X=9.045 $Y=1.185
+ $X2=0 $Y2=0
cc_653 N_A_1034_368#_c_802_n N_A_1383_349#_c_994_n 0.0199132f $X=9.09 $Y=0.34
+ $X2=0 $Y2=0
cc_654 N_A_1034_368#_c_805_n N_A_1383_349#_c_994_n 0.0223601f $X=9.26 $Y=1.17
+ $X2=0 $Y2=0
cc_655 N_A_1034_368#_c_795_n N_A_1383_349#_c_1000_n 0.00481612f $X=9.12 $Y=1.26
+ $X2=0 $Y2=0
cc_656 N_A_1034_368#_c_805_n N_A_1383_349#_c_1000_n 0.0011706f $X=9.26 $Y=1.17
+ $X2=0 $Y2=0
cc_657 N_A_1034_368#_c_807_n N_A_1383_349#_c_1000_n 0.00385352f $X=9.95 $Y=2.165
+ $X2=0 $Y2=0
cc_658 N_A_1034_368#_c_795_n N_A_1383_349#_c_995_n 0.00241408f $X=9.12 $Y=1.26
+ $X2=0 $Y2=0
cc_659 N_A_1034_368#_c_793_n N_A_1242_457#_M1040_g 0.0131362f $X=9.045 $Y=1.185
+ $X2=0 $Y2=0
cc_660 N_A_1034_368#_c_802_n N_A_1242_457#_M1040_g 0.0120273f $X=9.09 $Y=0.34
+ $X2=0 $Y2=0
cc_661 N_A_1034_368#_c_858_p N_A_1242_457#_M1040_g 6.7135e-19 $X=9.175 $Y=1.005
+ $X2=0 $Y2=0
cc_662 N_A_1034_368#_c_795_n N_A_1242_457#_c_1083_n 0.0131362f $X=9.12 $Y=1.26
+ $X2=0 $Y2=0
cc_663 N_A_1034_368#_c_813_n N_A_1242_457#_c_1092_n 0.00318252f $X=6.135 $Y=2.21
+ $X2=0 $Y2=0
cc_664 N_A_1034_368#_c_790_n N_A_1242_457#_c_1092_n 4.39571e-19 $X=6.51 $Y=1.71
+ $X2=0 $Y2=0
cc_665 N_A_1034_368#_c_791_n N_A_1242_457#_c_1092_n 5.28117e-19 $X=6.695
+ $Y=1.355 $X2=0 $Y2=0
cc_666 N_A_1034_368#_c_813_n N_A_1242_457#_c_1085_n 2.13752e-19 $X=6.135 $Y=2.21
+ $X2=0 $Y2=0
cc_667 N_A_1034_368#_c_791_n N_A_1242_457#_c_1085_n 0.00803564f $X=6.695
+ $Y=1.355 $X2=0 $Y2=0
cc_668 N_A_1034_368#_M1003_g N_A_1242_457#_c_1085_n 0.00554176f $X=6.695 $Y=0.9
+ $X2=0 $Y2=0
cc_669 N_A_1034_368#_c_790_n N_A_1242_457#_c_1089_n 6.35169e-19 $X=6.51 $Y=1.71
+ $X2=0 $Y2=0
cc_670 N_A_1034_368#_c_791_n N_A_1242_457#_c_1089_n 0.00378246f $X=6.695
+ $Y=1.355 $X2=0 $Y2=0
cc_671 N_A_1034_368#_M1003_g N_A_1242_457#_c_1089_n 0.0149994f $X=6.695 $Y=0.9
+ $X2=0 $Y2=0
cc_672 N_A_1034_368#_c_798_n N_A_1242_457#_c_1089_n 0.0329234f $X=7.04 $Y=0.415
+ $X2=0 $Y2=0
cc_673 N_A_1034_368#_c_810_n N_A_1242_457#_c_1089_n 0.00290442f $X=7.125
+ $Y=0.415 $X2=0 $Y2=0
cc_674 N_A_1034_368#_c_797_n N_A_855_368#_c_1202_n 7.62202e-19 $X=5.56 $Y=1.635
+ $X2=0 $Y2=0
cc_675 N_A_1034_368#_c_808_n N_A_855_368#_c_1202_n 0.0119607f $X=5.4 $Y=1.8
+ $X2=0 $Y2=0
cc_676 N_A_1034_368#_c_796_n N_A_855_368#_M1007_g 0.00707355f $X=5.405 $Y=0.515
+ $X2=0 $Y2=0
cc_677 N_A_1034_368#_c_797_n N_A_855_368#_M1007_g 0.00254048f $X=5.56 $Y=1.635
+ $X2=0 $Y2=0
cc_678 N_A_1034_368#_c_799_n N_A_855_368#_M1007_g 0.00290968f $X=5.645 $Y=0.415
+ $X2=0 $Y2=0
cc_679 N_A_1034_368#_c_809_n N_A_855_368#_M1007_g 0.00309908f $X=5.442 $Y=1.125
+ $X2=0 $Y2=0
cc_680 N_A_1034_368#_c_797_n N_A_855_368#_c_1204_n 0.00504919f $X=5.56 $Y=1.635
+ $X2=0 $Y2=0
cc_681 N_A_1034_368#_c_808_n N_A_855_368#_c_1204_n 0.00105281f $X=5.4 $Y=1.8
+ $X2=0 $Y2=0
cc_682 N_A_1034_368#_c_809_n N_A_855_368#_c_1204_n 0.00394715f $X=5.442 $Y=1.125
+ $X2=0 $Y2=0
cc_683 N_A_1034_368#_c_812_n N_A_855_368#_c_1205_n 0.00852849f $X=6.135 $Y=2.12
+ $X2=0 $Y2=0
cc_684 N_A_1034_368#_c_813_n N_A_855_368#_c_1205_n 0.0127466f $X=6.135 $Y=2.21
+ $X2=0 $Y2=0
cc_685 N_A_1034_368#_c_797_n N_A_855_368#_c_1205_n 0.0106342f $X=5.56 $Y=1.635
+ $X2=0 $Y2=0
cc_686 N_A_1034_368#_c_800_n N_A_855_368#_c_1205_n 0.00715637f $X=6.065 $Y=1.8
+ $X2=0 $Y2=0
cc_687 N_A_1034_368#_c_808_n N_A_855_368#_c_1205_n 0.0134367f $X=5.4 $Y=1.8
+ $X2=0 $Y2=0
cc_688 N_A_1034_368#_c_811_n N_A_855_368#_c_1205_n 0.0213787f $X=6.065 $Y=1.71
+ $X2=0 $Y2=0
cc_689 N_A_1034_368#_c_791_n N_A_855_368#_c_1206_n 0.00220632f $X=6.695 $Y=1.355
+ $X2=0 $Y2=0
cc_690 N_A_1034_368#_c_800_n N_A_855_368#_c_1206_n 0.00513789f $X=6.065 $Y=1.8
+ $X2=0 $Y2=0
cc_691 N_A_1034_368#_c_811_n N_A_855_368#_c_1206_n 0.0198941f $X=6.065 $Y=1.71
+ $X2=0 $Y2=0
cc_692 N_A_1034_368#_c_813_n N_A_855_368#_c_1219_n 0.00899647f $X=6.135 $Y=2.21
+ $X2=0 $Y2=0
cc_693 N_A_1034_368#_M1003_g N_A_855_368#_M1004_g 0.0185497f $X=6.695 $Y=0.9
+ $X2=0 $Y2=0
cc_694 N_A_1034_368#_c_796_n N_A_855_368#_M1004_g 0.00432442f $X=5.405 $Y=0.515
+ $X2=0 $Y2=0
cc_695 N_A_1034_368#_c_798_n N_A_855_368#_M1004_g 0.00661564f $X=7.04 $Y=0.415
+ $X2=0 $Y2=0
cc_696 N_A_1034_368#_c_813_n N_A_855_368#_c_1221_n 0.00278823f $X=6.135 $Y=2.21
+ $X2=0 $Y2=0
cc_697 N_A_1034_368#_c_813_n N_A_855_368#_c_1223_n 0.0120679f $X=6.135 $Y=2.21
+ $X2=0 $Y2=0
cc_698 N_A_1034_368#_c_791_n N_A_855_368#_c_1223_n 0.0058266f $X=6.695 $Y=1.355
+ $X2=0 $Y2=0
cc_699 N_A_1034_368#_c_816_n N_A_855_368#_M1025_g 0.001338f $X=10.11 $Y=2.465
+ $X2=0 $Y2=0
cc_700 N_A_1034_368#_c_807_n N_A_855_368#_M1025_g 0.00134374f $X=9.95 $Y=2.165
+ $X2=0 $Y2=0
cc_701 N_A_1034_368#_c_816_n N_A_855_368#_c_1208_n 0.0207729f $X=10.11 $Y=2.465
+ $X2=0 $Y2=0
cc_702 N_A_1034_368#_c_806_n N_A_855_368#_c_1208_n 0.0169827f $X=9.645 $Y=1.17
+ $X2=0 $Y2=0
cc_703 N_A_1034_368#_c_807_n N_A_855_368#_c_1208_n 0.0202931f $X=9.95 $Y=2.165
+ $X2=0 $Y2=0
cc_704 N_A_1034_368#_c_794_n N_A_855_368#_c_1227_n 0.0169827f $X=9.48 $Y=1.26
+ $X2=0 $Y2=0
cc_705 N_A_1034_368#_c_804_n N_A_855_368#_c_1227_n 0.00271869f $X=9.785 $Y=1.17
+ $X2=0 $Y2=0
cc_706 N_A_1034_368#_c_805_n N_A_855_368#_c_1227_n 6.613e-19 $X=9.26 $Y=1.17
+ $X2=0 $Y2=0
cc_707 N_A_1034_368#_c_807_n N_A_855_368#_c_1227_n 5.48883e-19 $X=9.95 $Y=2.165
+ $X2=0 $Y2=0
cc_708 N_A_1034_368#_c_807_n N_A_855_368#_c_1209_n 0.00569302f $X=9.95 $Y=2.165
+ $X2=0 $Y2=0
cc_709 N_A_1034_368#_c_797_n N_A_855_368#_c_1211_n 0.00611873f $X=5.56 $Y=1.635
+ $X2=0 $Y2=0
cc_710 N_A_1034_368#_c_816_n N_A_855_368#_c_1229_n 0.00415106f $X=10.11 $Y=2.465
+ $X2=0 $Y2=0
cc_711 N_A_1034_368#_c_804_n N_A_855_368#_c_1212_n 0.00289132f $X=9.785 $Y=1.17
+ $X2=0 $Y2=0
cc_712 N_A_1034_368#_c_806_n N_A_855_368#_c_1212_n 0.0181127f $X=9.645 $Y=1.17
+ $X2=0 $Y2=0
cc_713 N_A_1034_368#_c_796_n N_A_855_368#_c_1253_n 0.0102862f $X=5.405 $Y=0.515
+ $X2=0 $Y2=0
cc_714 N_A_1034_368#_c_808_n N_A_855_368#_c_1230_n 0.00824733f $X=5.4 $Y=1.8
+ $X2=0 $Y2=0
cc_715 N_A_1034_368#_c_797_n N_A_855_368#_c_1214_n 0.00572729f $X=5.56 $Y=1.635
+ $X2=0 $Y2=0
cc_716 N_A_1034_368#_c_809_n N_A_855_368#_c_1214_n 0.00191706f $X=5.442 $Y=1.125
+ $X2=0 $Y2=0
cc_717 N_A_1034_368#_c_797_n N_A_855_368#_c_1215_n 3.41517e-19 $X=5.56 $Y=1.635
+ $X2=0 $Y2=0
cc_718 N_A_1034_368#_c_808_n N_A_855_368#_c_1215_n 0.00842419f $X=5.4 $Y=1.8
+ $X2=0 $Y2=0
cc_719 N_A_1034_368#_c_808_n N_A_855_368#_c_1232_n 0.00452944f $X=5.4 $Y=1.8
+ $X2=0 $Y2=0
cc_720 N_A_1034_368#_c_797_n N_A_855_368#_c_1216_n 0.02517f $X=5.56 $Y=1.635
+ $X2=0 $Y2=0
cc_721 N_A_1034_368#_c_808_n N_A_855_368#_c_1216_n 0.0114292f $X=5.4 $Y=1.8
+ $X2=0 $Y2=0
cc_722 N_A_1034_368#_c_809_n N_A_855_368#_c_1216_n 0.00528992f $X=5.442 $Y=1.125
+ $X2=0 $Y2=0
cc_723 N_A_1034_368#_c_816_n N_A_2082_446#_c_1408_n 0.0313578f $X=10.11 $Y=2.465
+ $X2=0 $Y2=0
cc_724 N_A_1034_368#_c_816_n N_A_2082_446#_c_1409_n 0.0134605f $X=10.11 $Y=2.465
+ $X2=0 $Y2=0
cc_725 N_A_1034_368#_c_816_n N_A_2082_446#_c_1400_n 0.0127423f $X=10.11 $Y=2.465
+ $X2=0 $Y2=0
cc_726 N_A_1034_368#_c_802_n N_A_1824_74#_M1024_d 0.00248108f $X=9.09 $Y=0.34
+ $X2=-0.19 $Y2=-0.245
cc_727 N_A_1034_368#_c_858_p N_A_1824_74#_M1024_d 0.0130256f $X=9.175 $Y=1.005
+ $X2=-0.19 $Y2=-0.245
cc_728 N_A_1034_368#_c_804_n N_A_1824_74#_M1024_d 0.00450592f $X=9.785 $Y=1.17
+ $X2=-0.19 $Y2=-0.245
cc_729 N_A_1034_368#_c_816_n N_A_1824_74#_c_1553_n 0.004427f $X=10.11 $Y=2.465
+ $X2=0 $Y2=0
cc_730 N_A_1034_368#_c_804_n N_A_1824_74#_c_1553_n 0.00861974f $X=9.785 $Y=1.17
+ $X2=0 $Y2=0
cc_731 N_A_1034_368#_c_807_n N_A_1824_74#_c_1553_n 0.0339543f $X=9.95 $Y=2.165
+ $X2=0 $Y2=0
cc_732 N_A_1034_368#_c_793_n N_A_1824_74#_c_1528_n 0.0018748f $X=9.045 $Y=1.185
+ $X2=0 $Y2=0
cc_733 N_A_1034_368#_c_794_n N_A_1824_74#_c_1528_n 2.42458e-19 $X=9.48 $Y=1.26
+ $X2=0 $Y2=0
cc_734 N_A_1034_368#_c_858_p N_A_1824_74#_c_1528_n 0.026719f $X=9.175 $Y=1.005
+ $X2=0 $Y2=0
cc_735 N_A_1034_368#_c_804_n N_A_1824_74#_c_1528_n 0.0466861f $X=9.785 $Y=1.17
+ $X2=0 $Y2=0
cc_736 N_A_1034_368#_c_806_n N_A_1824_74#_c_1528_n 0.0070276f $X=9.645 $Y=1.17
+ $X2=0 $Y2=0
cc_737 N_A_1034_368#_c_816_n N_A_1824_74#_c_1540_n 0.0157095f $X=10.11 $Y=2.465
+ $X2=0 $Y2=0
cc_738 N_A_1034_368#_c_807_n N_A_1824_74#_c_1540_n 0.019012f $X=9.95 $Y=2.165
+ $X2=0 $Y2=0
cc_739 N_A_1034_368#_c_804_n N_A_1824_74#_c_1529_n 0.00187033f $X=9.785 $Y=1.17
+ $X2=0 $Y2=0
cc_740 N_A_1034_368#_c_816_n N_A_1824_74#_c_1530_n 0.00479636f $X=10.11 $Y=2.465
+ $X2=0 $Y2=0
cc_741 N_A_1034_368#_c_804_n N_A_1824_74#_c_1530_n 0.0107493f $X=9.785 $Y=1.17
+ $X2=0 $Y2=0
cc_742 N_A_1034_368#_c_807_n N_A_1824_74#_c_1530_n 0.0746733f $X=9.95 $Y=2.165
+ $X2=0 $Y2=0
cc_743 N_A_1034_368#_c_804_n N_A_1824_74#_c_1532_n 0.0146626f $X=9.785 $Y=1.17
+ $X2=0 $Y2=0
cc_744 N_A_1034_368#_c_816_n N_VPWR_c_1745_n 0.00308386f $X=10.11 $Y=2.465 $X2=0
+ $Y2=0
cc_745 N_A_1034_368#_c_816_n N_VPWR_c_1751_n 0.0012612f $X=10.11 $Y=2.465 $X2=0
+ $Y2=0
cc_746 N_A_1034_368#_c_813_n N_VPWR_c_1727_n 9.49986e-19 $X=6.135 $Y=2.21 $X2=0
+ $Y2=0
cc_747 N_A_1034_368#_c_816_n N_VPWR_c_1727_n 0.00381714f $X=10.11 $Y=2.465 $X2=0
+ $Y2=0
cc_748 N_A_1034_368#_M1032_d N_A_390_81#_c_1913_n 0.00696197f $X=5.17 $Y=1.84
+ $X2=0 $Y2=0
cc_749 N_A_1034_368#_c_800_n N_A_390_81#_c_1913_n 0.00189471f $X=6.065 $Y=1.8
+ $X2=0 $Y2=0
cc_750 N_A_1034_368#_c_808_n N_A_390_81#_c_1913_n 0.0233646f $X=5.4 $Y=1.8 $X2=0
+ $Y2=0
cc_751 N_A_1034_368#_M1003_g N_A_390_81#_c_1907_n 6.49857e-19 $X=6.695 $Y=0.9
+ $X2=0 $Y2=0
cc_752 N_A_1034_368#_c_796_n N_A_390_81#_c_1907_n 0.0514496f $X=5.405 $Y=0.515
+ $X2=0 $Y2=0
cc_753 N_A_1034_368#_c_798_n N_A_390_81#_c_1907_n 0.0262076f $X=7.04 $Y=0.415
+ $X2=0 $Y2=0
cc_754 N_A_1034_368#_c_813_n N_A_390_81#_c_1915_n 0.0147311f $X=6.135 $Y=2.21
+ $X2=0 $Y2=0
cc_755 N_A_1034_368#_c_790_n N_A_390_81#_c_1915_n 0.00246862f $X=6.51 $Y=1.71
+ $X2=0 $Y2=0
cc_756 N_A_1034_368#_c_800_n N_A_390_81#_c_1915_n 0.0109321f $X=6.065 $Y=1.8
+ $X2=0 $Y2=0
cc_757 N_A_1034_368#_c_811_n N_A_390_81#_c_1915_n 9.60671e-19 $X=6.065 $Y=1.71
+ $X2=0 $Y2=0
cc_758 N_A_1034_368#_c_791_n N_A_390_81#_c_1908_n 0.00410506f $X=6.695 $Y=1.355
+ $X2=0 $Y2=0
cc_759 N_A_1034_368#_M1003_g N_A_390_81#_c_1908_n 4.96156e-19 $X=6.695 $Y=0.9
+ $X2=0 $Y2=0
cc_760 N_A_1034_368#_c_800_n N_A_390_81#_c_1908_n 0.00322721f $X=6.065 $Y=1.8
+ $X2=0 $Y2=0
cc_761 N_A_1034_368#_c_811_n N_A_390_81#_c_1908_n 0.00328043f $X=6.065 $Y=1.71
+ $X2=0 $Y2=0
cc_762 N_A_1034_368#_c_797_n N_A_390_81#_c_1909_n 0.0132897f $X=5.56 $Y=1.635
+ $X2=0 $Y2=0
cc_763 N_A_1034_368#_c_800_n N_A_390_81#_c_1909_n 0.0271035f $X=6.065 $Y=1.8
+ $X2=0 $Y2=0
cc_764 N_A_1034_368#_c_811_n N_A_390_81#_c_1909_n 0.0016654f $X=6.065 $Y=1.71
+ $X2=0 $Y2=0
cc_765 N_A_1034_368#_c_812_n N_A_390_81#_c_1910_n 0.00365666f $X=6.135 $Y=2.12
+ $X2=0 $Y2=0
cc_766 N_A_1034_368#_c_790_n N_A_390_81#_c_1910_n 0.0104977f $X=6.51 $Y=1.71
+ $X2=0 $Y2=0
cc_767 N_A_1034_368#_c_791_n N_A_390_81#_c_1910_n 0.00657268f $X=6.695 $Y=1.355
+ $X2=0 $Y2=0
cc_768 N_A_1034_368#_c_800_n N_A_390_81#_c_1910_n 0.0257057f $X=6.065 $Y=1.8
+ $X2=0 $Y2=0
cc_769 N_A_1034_368#_c_811_n N_A_390_81#_c_1910_n 0.00207319f $X=6.065 $Y=1.71
+ $X2=0 $Y2=0
cc_770 N_A_1034_368#_c_813_n N_A_390_81#_c_1918_n 0.00510388f $X=6.135 $Y=2.21
+ $X2=0 $Y2=0
cc_771 N_A_1034_368#_c_800_n N_A_390_81#_c_1918_n 0.0165466f $X=6.065 $Y=1.8
+ $X2=0 $Y2=0
cc_772 N_A_1034_368#_c_808_n N_A_390_81#_c_1918_n 0.00516423f $X=5.4 $Y=1.8
+ $X2=0 $Y2=0
cc_773 N_A_1034_368#_c_811_n N_A_390_81#_c_1918_n 0.00166973f $X=6.065 $Y=1.71
+ $X2=0 $Y2=0
cc_774 N_A_1034_368#_c_801_n N_VGND_M1021_d 0.0214581f $X=8.25 $Y=0.665 $X2=0
+ $Y2=0
cc_775 N_A_1034_368#_c_972_p N_VGND_M1021_d 0.00612573f $X=8.335 $Y=0.58 $X2=0
+ $Y2=0
cc_776 N_A_1034_368#_c_803_n N_VGND_M1021_d 0.00122695f $X=8.42 $Y=0.34 $X2=0
+ $Y2=0
cc_777 N_A_1034_368#_c_799_n N_VGND_c_2080_n 0.0087905f $X=5.645 $Y=0.415 $X2=0
+ $Y2=0
cc_778 N_A_1034_368#_c_798_n N_VGND_c_2090_n 0.0611023f $X=7.04 $Y=0.415 $X2=0
+ $Y2=0
cc_779 N_A_1034_368#_c_799_n N_VGND_c_2090_n 0.0195675f $X=5.645 $Y=0.415 $X2=0
+ $Y2=0
cc_780 N_A_1034_368#_c_801_n N_VGND_c_2090_n 0.0432912f $X=8.25 $Y=0.665 $X2=0
+ $Y2=0
cc_781 N_A_1034_368#_c_803_n N_VGND_c_2090_n 0.0139413f $X=8.42 $Y=0.34 $X2=0
+ $Y2=0
cc_782 N_A_1034_368#_c_810_n N_VGND_c_2090_n 0.0115182f $X=7.125 $Y=0.415 $X2=0
+ $Y2=0
cc_783 N_A_1034_368#_c_793_n N_VGND_c_2091_n 0.00278242f $X=9.045 $Y=1.185 $X2=0
+ $Y2=0
cc_784 N_A_1034_368#_c_801_n N_VGND_c_2091_n 0.00335833f $X=8.25 $Y=0.665 $X2=0
+ $Y2=0
cc_785 N_A_1034_368#_c_802_n N_VGND_c_2091_n 0.0544002f $X=9.09 $Y=0.34 $X2=0
+ $Y2=0
cc_786 N_A_1034_368#_c_803_n N_VGND_c_2091_n 0.0118998f $X=8.42 $Y=0.34 $X2=0
+ $Y2=0
cc_787 N_A_1034_368#_c_793_n N_VGND_c_2100_n 0.00359177f $X=9.045 $Y=1.185 $X2=0
+ $Y2=0
cc_788 N_A_1034_368#_c_798_n N_VGND_c_2100_n 0.0500008f $X=7.04 $Y=0.415 $X2=0
+ $Y2=0
cc_789 N_A_1034_368#_c_799_n N_VGND_c_2100_n 0.015016f $X=5.645 $Y=0.415 $X2=0
+ $Y2=0
cc_790 N_A_1034_368#_c_801_n N_VGND_c_2100_n 0.0191252f $X=8.25 $Y=0.665 $X2=0
+ $Y2=0
cc_791 N_A_1034_368#_c_802_n N_VGND_c_2100_n 0.0304263f $X=9.09 $Y=0.34 $X2=0
+ $Y2=0
cc_792 N_A_1034_368#_c_803_n N_VGND_c_2100_n 0.00655543f $X=8.42 $Y=0.34 $X2=0
+ $Y2=0
cc_793 N_A_1034_368#_c_810_n N_VGND_c_2100_n 0.00618366f $X=7.125 $Y=0.415 $X2=0
+ $Y2=0
cc_794 N_A_1034_368#_c_801_n A_1432_138# 0.0013295f $X=8.25 $Y=0.665 $X2=-0.19
+ $Y2=-0.245
cc_795 N_A_1383_349#_c_1013_n N_A_1242_457#_M1040_g 0.0148889f $X=8.59 $Y=1.005
+ $X2=0 $Y2=0
cc_796 N_A_1383_349#_c_994_n N_A_1242_457#_M1040_g 0.0150489f $X=8.755 $Y=0.86
+ $X2=0 $Y2=0
cc_797 N_A_1383_349#_c_995_n N_A_1242_457#_M1040_g 0.00617118f $X=8.932 $Y=1.715
+ $X2=0 $Y2=0
cc_798 N_A_1383_349#_c_994_n N_A_1242_457#_c_1083_n 0.00463727f $X=8.755 $Y=0.86
+ $X2=0 $Y2=0
cc_799 N_A_1383_349#_c_995_n N_A_1242_457#_c_1083_n 0.016456f $X=8.932 $Y=1.715
+ $X2=0 $Y2=0
cc_800 N_A_1383_349#_c_1013_n N_A_1242_457#_c_1084_n 0.00840745f $X=8.59
+ $Y=1.005 $X2=0 $Y2=0
cc_801 N_A_1383_349#_c_996_n N_A_1242_457#_c_1085_n 0.00743747f $X=7.005 $Y=2.21
+ $X2=0 $Y2=0
cc_802 N_A_1383_349#_M1035_g N_A_1242_457#_c_1085_n 0.0036446f $X=7.085 $Y=0.9
+ $X2=0 $Y2=0
cc_803 N_A_1383_349#_c_993_n N_A_1242_457#_c_1085_n 0.0696484f $X=7.165 $Y=1.91
+ $X2=0 $Y2=0
cc_804 N_A_1383_349#_c_996_n N_A_1242_457#_c_1105_n 0.0124345f $X=7.005 $Y=2.21
+ $X2=0 $Y2=0
cc_805 N_A_1383_349#_c_993_n N_A_1242_457#_c_1105_n 0.010168f $X=7.165 $Y=1.91
+ $X2=0 $Y2=0
cc_806 N_A_1383_349#_c_996_n N_A_1242_457#_c_1086_n 0.00433331f $X=7.005 $Y=2.21
+ $X2=0 $Y2=0
cc_807 N_A_1383_349#_M1035_g N_A_1242_457#_c_1086_n 4.10299e-19 $X=7.085 $Y=0.9
+ $X2=0 $Y2=0
cc_808 N_A_1383_349#_c_993_n N_A_1242_457#_c_1086_n 0.0370159f $X=7.165 $Y=1.91
+ $X2=0 $Y2=0
cc_809 N_A_1383_349#_M1035_g N_A_1242_457#_c_1087_n 7.98464e-19 $X=7.085 $Y=0.9
+ $X2=0 $Y2=0
cc_810 N_A_1383_349#_c_993_n N_A_1242_457#_c_1087_n 0.0271618f $X=7.165 $Y=1.91
+ $X2=0 $Y2=0
cc_811 N_A_1383_349#_c_1013_n N_A_1242_457#_c_1087_n 0.0111252f $X=8.59 $Y=1.005
+ $X2=0 $Y2=0
cc_812 N_A_1383_349#_c_1013_n N_A_1242_457#_c_1088_n 0.0573215f $X=8.59 $Y=1.005
+ $X2=0 $Y2=0
cc_813 N_A_1383_349#_c_995_n N_A_1242_457#_c_1088_n 0.0151715f $X=8.932 $Y=1.715
+ $X2=0 $Y2=0
cc_814 N_A_1383_349#_M1035_g N_A_1242_457#_c_1089_n 0.002196f $X=7.085 $Y=0.9
+ $X2=0 $Y2=0
cc_815 N_A_1383_349#_c_993_n N_A_1242_457#_c_1089_n 0.00279586f $X=7.165 $Y=1.91
+ $X2=0 $Y2=0
cc_816 N_A_1383_349#_c_1030_n N_A_1242_457#_c_1089_n 0.0130355f $X=7.315
+ $Y=1.005 $X2=0 $Y2=0
cc_817 N_A_1383_349#_c_996_n N_A_1242_457#_c_1095_n 0.00590261f $X=7.005 $Y=2.21
+ $X2=0 $Y2=0
cc_818 N_A_1383_349#_c_996_n N_A_855_368#_c_1221_n 0.00284772f $X=7.005 $Y=2.21
+ $X2=0 $Y2=0
cc_819 N_A_1383_349#_c_996_n N_A_855_368#_c_1223_n 0.0259599f $X=7.005 $Y=2.21
+ $X2=0 $Y2=0
cc_820 N_A_1383_349#_c_996_n N_A_855_368#_c_1224_n 0.00862445f $X=7.005 $Y=2.21
+ $X2=0 $Y2=0
cc_821 N_A_1383_349#_c_999_n N_A_855_368#_c_1224_n 0.00737375f $X=8.95 $Y=2.235
+ $X2=0 $Y2=0
cc_822 N_A_1383_349#_c_1000_n N_A_855_368#_M1025_g 0.0104192f $X=8.95 $Y=1.88
+ $X2=0 $Y2=0
cc_823 N_A_1383_349#_c_1000_n N_A_855_368#_c_1227_n 7.1022e-19 $X=8.95 $Y=1.88
+ $X2=0 $Y2=0
cc_824 N_A_1383_349#_c_995_n N_A_855_368#_c_1227_n 0.00307401f $X=8.932 $Y=1.715
+ $X2=0 $Y2=0
cc_825 N_A_1383_349#_c_1000_n N_A_1824_74#_c_1553_n 0.0438134f $X=8.95 $Y=1.88
+ $X2=0 $Y2=0
cc_826 N_A_1383_349#_c_999_n N_A_1824_74#_c_1541_n 0.0168727f $X=8.95 $Y=2.235
+ $X2=0 $Y2=0
cc_827 N_A_1383_349#_c_996_n N_VPWR_c_1730_n 0.00392315f $X=7.005 $Y=2.21 $X2=0
+ $Y2=0
cc_828 N_A_1383_349#_c_999_n N_VPWR_c_1731_n 0.0171249f $X=8.95 $Y=2.235 $X2=0
+ $Y2=0
cc_829 N_A_1383_349#_c_999_n N_VPWR_c_1745_n 0.00805754f $X=8.95 $Y=2.235 $X2=0
+ $Y2=0
cc_830 N_A_1383_349#_c_996_n N_VPWR_c_1727_n 9.49986e-19 $X=7.005 $Y=2.21 $X2=0
+ $Y2=0
cc_831 N_A_1383_349#_c_999_n N_VPWR_c_1727_n 0.0100713f $X=8.95 $Y=2.235 $X2=0
+ $Y2=0
cc_832 N_A_1383_349#_c_1013_n N_VGND_M1021_d 0.0209614f $X=8.59 $Y=1.005 $X2=0
+ $Y2=0
cc_833 N_A_1383_349#_M1035_g N_VGND_c_2090_n 4.68109e-19 $X=7.085 $Y=0.9 $X2=0
+ $Y2=0
cc_834 N_A_1383_349#_c_993_n A_1432_138# 2.2331e-19 $X=7.165 $Y=1.91 $X2=-0.19
+ $Y2=-0.245
cc_835 N_A_1383_349#_c_1013_n A_1432_138# 0.00102891f $X=8.59 $Y=1.005 $X2=-0.19
+ $Y2=-0.245
cc_836 N_A_1383_349#_c_1030_n A_1432_138# 0.00108716f $X=7.315 $Y=1.005
+ $X2=-0.19 $Y2=-0.245
cc_837 N_A_1242_457#_c_1092_n N_A_855_368#_c_1219_n 0.00366466f $X=6.7 $Y=2.6
+ $X2=0 $Y2=0
cc_838 N_A_1242_457#_c_1085_n N_A_855_368#_M1004_g 6.17163e-19 $X=6.785 $Y=2.32
+ $X2=0 $Y2=0
cc_839 N_A_1242_457#_c_1089_n N_A_855_368#_M1004_g 0.00249151f $X=6.48 $Y=0.895
+ $X2=0 $Y2=0
cc_840 N_A_1242_457#_c_1092_n N_A_855_368#_c_1221_n 9.75099e-19 $X=6.7 $Y=2.6
+ $X2=0 $Y2=0
cc_841 N_A_1242_457#_c_1092_n N_A_855_368#_c_1223_n 0.0105779f $X=6.7 $Y=2.6
+ $X2=0 $Y2=0
cc_842 N_A_1242_457#_c_1085_n N_A_855_368#_c_1223_n 0.00105048f $X=6.785 $Y=2.32
+ $X2=0 $Y2=0
cc_843 N_A_1242_457#_c_1083_n N_A_855_368#_c_1224_n 0.0103562f $X=8.64 $Y=1.66
+ $X2=0 $Y2=0
cc_844 N_A_1242_457#_c_1092_n N_A_855_368#_c_1224_n 4.45551e-19 $X=6.7 $Y=2.6
+ $X2=0 $Y2=0
cc_845 N_A_1242_457#_c_1105_n N_A_855_368#_c_1224_n 0.00245825f $X=7.485
+ $Y=2.405 $X2=0 $Y2=0
cc_846 N_A_1242_457#_c_1086_n N_A_855_368#_c_1224_n 0.00747767f $X=7.57 $Y=2.32
+ $X2=0 $Y2=0
cc_847 N_A_1242_457#_c_1095_n N_A_855_368#_c_1224_n 0.00336263f $X=6.785
+ $Y=2.522 $X2=0 $Y2=0
cc_848 N_A_1242_457#_c_1083_n N_A_855_368#_M1025_g 0.0199663f $X=8.64 $Y=1.66
+ $X2=0 $Y2=0
cc_849 N_A_1242_457#_c_1083_n N_A_855_368#_c_1227_n 0.00359436f $X=8.64 $Y=1.66
+ $X2=0 $Y2=0
cc_850 N_A_1242_457#_c_1083_n N_A_1824_74#_c_1541_n 4.59845e-19 $X=8.64 $Y=1.66
+ $X2=0 $Y2=0
cc_851 N_A_1242_457#_c_1105_n N_VPWR_M1000_d 0.00807089f $X=7.485 $Y=2.405 $X2=0
+ $Y2=0
cc_852 N_A_1242_457#_c_1086_n N_VPWR_M1000_d 5.12435e-19 $X=7.57 $Y=2.32 $X2=0
+ $Y2=0
cc_853 N_A_1242_457#_c_1105_n N_VPWR_c_1730_n 0.0256457f $X=7.485 $Y=2.405 $X2=0
+ $Y2=0
cc_854 N_A_1242_457#_c_1086_n N_VPWR_c_1730_n 0.00442355f $X=7.57 $Y=2.32 $X2=0
+ $Y2=0
cc_855 N_A_1242_457#_c_1095_n N_VPWR_c_1730_n 0.00389678f $X=6.785 $Y=2.522
+ $X2=0 $Y2=0
cc_856 N_A_1242_457#_c_1083_n N_VPWR_c_1731_n 0.0100186f $X=8.64 $Y=1.66 $X2=0
+ $Y2=0
cc_857 N_A_1242_457#_c_1086_n N_VPWR_c_1731_n 0.0280602f $X=7.57 $Y=2.32 $X2=0
+ $Y2=0
cc_858 N_A_1242_457#_c_1092_n N_VPWR_c_1738_n 0.00974072f $X=6.7 $Y=2.6 $X2=0
+ $Y2=0
cc_859 N_A_1242_457#_c_1095_n N_VPWR_c_1738_n 0.00364053f $X=6.785 $Y=2.522
+ $X2=0 $Y2=0
cc_860 N_A_1242_457#_c_1086_n N_VPWR_c_1744_n 0.00680673f $X=7.57 $Y=2.32 $X2=0
+ $Y2=0
cc_861 N_A_1242_457#_c_1083_n N_VPWR_c_1727_n 8.51577e-19 $X=8.64 $Y=1.66 $X2=0
+ $Y2=0
cc_862 N_A_1242_457#_c_1092_n N_VPWR_c_1727_n 0.0127724f $X=6.7 $Y=2.6 $X2=0
+ $Y2=0
cc_863 N_A_1242_457#_c_1105_n N_VPWR_c_1727_n 0.00916028f $X=7.485 $Y=2.405
+ $X2=0 $Y2=0
cc_864 N_A_1242_457#_c_1086_n N_VPWR_c_1727_n 0.0152918f $X=7.57 $Y=2.32 $X2=0
+ $Y2=0
cc_865 N_A_1242_457#_c_1095_n N_VPWR_c_1727_n 0.00458771f $X=6.785 $Y=2.522
+ $X2=0 $Y2=0
cc_866 N_A_1242_457#_c_1085_n N_A_390_81#_c_1907_n 0.00454965f $X=6.785 $Y=2.32
+ $X2=0 $Y2=0
cc_867 N_A_1242_457#_c_1089_n N_A_390_81#_c_1907_n 0.0185813f $X=6.48 $Y=0.895
+ $X2=0 $Y2=0
cc_868 N_A_1242_457#_M1028_d N_A_390_81#_c_1915_n 0.00201205f $X=6.21 $Y=2.285
+ $X2=0 $Y2=0
cc_869 N_A_1242_457#_c_1092_n N_A_390_81#_c_1915_n 0.0163086f $X=6.7 $Y=2.6
+ $X2=0 $Y2=0
cc_870 N_A_1242_457#_c_1085_n N_A_390_81#_c_1915_n 0.0126252f $X=6.785 $Y=2.32
+ $X2=0 $Y2=0
cc_871 N_A_1242_457#_c_1085_n N_A_390_81#_c_1908_n 0.0132424f $X=6.785 $Y=2.32
+ $X2=0 $Y2=0
cc_872 N_A_1242_457#_c_1089_n N_A_390_81#_c_1908_n 0.0191012f $X=6.48 $Y=0.895
+ $X2=0 $Y2=0
cc_873 N_A_1242_457#_c_1085_n N_A_390_81#_c_1910_n 0.048352f $X=6.785 $Y=2.32
+ $X2=0 $Y2=0
cc_874 N_A_1242_457#_c_1092_n N_A_390_81#_c_1918_n 0.0176736f $X=6.7 $Y=2.6
+ $X2=0 $Y2=0
cc_875 N_A_1242_457#_c_1085_n A_1332_457# 4.63054e-19 $X=6.785 $Y=2.32 $X2=-0.19
+ $Y2=-0.245
cc_876 N_A_1242_457#_c_1095_n A_1332_457# 0.0027348f $X=6.785 $Y=2.522 $X2=-0.19
+ $Y2=-0.245
cc_877 N_A_1242_457#_M1040_g N_VGND_c_2090_n 0.00115066f $X=8.54 $Y=0.74 $X2=0
+ $Y2=0
cc_878 N_A_1242_457#_M1040_g N_VGND_c_2091_n 0.00278271f $X=8.54 $Y=0.74 $X2=0
+ $Y2=0
cc_879 N_A_1242_457#_M1040_g N_VGND_c_2100_n 0.0035918f $X=8.54 $Y=0.74 $X2=0
+ $Y2=0
cc_880 N_A_1242_457#_c_1089_n A_1354_138# 0.0020913f $X=6.48 $Y=0.895 $X2=-0.19
+ $Y2=-0.245
cc_881 N_A_855_368#_c_1209_n N_A_2082_446#_M1009_g 0.00472321f $X=10.125
+ $Y=1.575 $X2=0 $Y2=0
cc_882 N_A_855_368#_M1008_g N_A_2082_446#_M1009_g 0.0465564f $X=10.315 $Y=0.58
+ $X2=0 $Y2=0
cc_883 N_A_855_368#_c_1208_n N_A_2082_446#_c_1400_n 0.00873113f $X=10.05 $Y=1.65
+ $X2=0 $Y2=0
cc_884 N_A_855_368#_c_1209_n N_A_2082_446#_c_1407_n 0.00873113f $X=10.125
+ $Y=1.575 $X2=0 $Y2=0
cc_885 N_A_855_368#_M1025_g N_A_1824_74#_c_1553_n 0.00686632f $X=9.26 $Y=2.33
+ $X2=0 $Y2=0
cc_886 N_A_855_368#_c_1208_n N_A_1824_74#_c_1553_n 0.00627973f $X=10.05 $Y=1.65
+ $X2=0 $Y2=0
cc_887 N_A_855_368#_M1008_g N_A_1824_74#_c_1528_n 0.0085841f $X=10.315 $Y=0.58
+ $X2=0 $Y2=0
cc_888 N_A_855_368#_c_1212_n N_A_1824_74#_c_1528_n 0.0073765f $X=10.315 $Y=1.055
+ $X2=0 $Y2=0
cc_889 N_A_855_368#_M1025_g N_A_1824_74#_c_1541_n 0.00525155f $X=9.26 $Y=2.33
+ $X2=0 $Y2=0
cc_890 N_A_855_368#_c_1229_n N_A_1824_74#_c_1541_n 4.63769e-19 $X=9.26 $Y=3.15
+ $X2=0 $Y2=0
cc_891 N_A_855_368#_M1008_g N_A_1824_74#_c_1529_n 0.00682018f $X=10.315 $Y=0.58
+ $X2=0 $Y2=0
cc_892 N_A_855_368#_c_1212_n N_A_1824_74#_c_1529_n 0.00308052f $X=10.315
+ $Y=1.055 $X2=0 $Y2=0
cc_893 N_A_855_368#_c_1209_n N_A_1824_74#_c_1530_n 0.00432791f $X=10.125
+ $Y=1.575 $X2=0 $Y2=0
cc_894 N_A_855_368#_c_1209_n N_A_1824_74#_c_1532_n 7.4004e-19 $X=10.125 $Y=1.575
+ $X2=0 $Y2=0
cc_895 N_A_855_368#_c_1212_n N_A_1824_74#_c_1532_n 0.00823777f $X=10.315
+ $Y=1.055 $X2=0 $Y2=0
cc_896 N_A_855_368#_c_1230_n N_VPWR_M1018_d 0.00232663f $X=4.815 $Y=1.905 $X2=0
+ $Y2=0
cc_897 N_A_855_368#_c_1202_n N_VPWR_c_1729_n 0.00888208f $X=5.095 $Y=1.765 $X2=0
+ $Y2=0
cc_898 N_A_855_368#_c_1205_n N_VPWR_c_1729_n 0.0017658f $X=5.615 $Y=3.075 $X2=0
+ $Y2=0
cc_899 N_A_855_368#_c_1220_n N_VPWR_c_1729_n 0.00232909f $X=5.69 $Y=3.15 $X2=0
+ $Y2=0
cc_900 N_A_855_368#_c_1221_n N_VPWR_c_1730_n 0.0066733f $X=6.585 $Y=2.87 $X2=0
+ $Y2=0
cc_901 N_A_855_368#_c_1224_n N_VPWR_c_1730_n 0.025635f $X=9.17 $Y=3.15 $X2=0
+ $Y2=0
cc_902 N_A_855_368#_c_1224_n N_VPWR_c_1731_n 0.0259473f $X=9.17 $Y=3.15 $X2=0
+ $Y2=0
cc_903 N_A_855_368#_M1025_g N_VPWR_c_1731_n 0.00149031f $X=9.26 $Y=2.33 $X2=0
+ $Y2=0
cc_904 N_A_855_368#_c_1229_n N_VPWR_c_1731_n 0.00415487f $X=9.26 $Y=3.15 $X2=0
+ $Y2=0
cc_905 N_A_855_368#_c_1202_n N_VPWR_c_1738_n 0.00413917f $X=5.095 $Y=1.765 $X2=0
+ $Y2=0
cc_906 N_A_855_368#_c_1220_n N_VPWR_c_1738_n 0.0484733f $X=5.69 $Y=3.15 $X2=0
+ $Y2=0
cc_907 N_A_855_368#_c_1224_n N_VPWR_c_1744_n 0.0233394f $X=9.17 $Y=3.15 $X2=0
+ $Y2=0
cc_908 N_A_855_368#_c_1224_n N_VPWR_c_1745_n 0.0232816f $X=9.17 $Y=3.15 $X2=0
+ $Y2=0
cc_909 N_A_855_368#_c_1202_n N_VPWR_c_1727_n 0.00399275f $X=5.095 $Y=1.765 $X2=0
+ $Y2=0
cc_910 N_A_855_368#_c_1219_n N_VPWR_c_1727_n 0.0243437f $X=6.495 $Y=3.15 $X2=0
+ $Y2=0
cc_911 N_A_855_368#_c_1220_n N_VPWR_c_1727_n 0.00693725f $X=5.69 $Y=3.15 $X2=0
+ $Y2=0
cc_912 N_A_855_368#_c_1224_n N_VPWR_c_1727_n 0.0584197f $X=9.17 $Y=3.15 $X2=0
+ $Y2=0
cc_913 N_A_855_368#_c_1228_n N_VPWR_c_1727_n 0.00504011f $X=6.585 $Y=3.15 $X2=0
+ $Y2=0
cc_914 N_A_855_368#_c_1229_n N_VPWR_c_1727_n 0.0122553f $X=9.26 $Y=3.15 $X2=0
+ $Y2=0
cc_915 N_A_855_368#_M1018_s N_A_390_81#_c_1913_n 0.0082239f $X=4.275 $Y=1.84
+ $X2=0 $Y2=0
cc_916 N_A_855_368#_c_1202_n N_A_390_81#_c_1913_n 0.0125758f $X=5.095 $Y=1.765
+ $X2=0 $Y2=0
cc_917 N_A_855_368#_c_1205_n N_A_390_81#_c_1913_n 0.0124767f $X=5.615 $Y=3.075
+ $X2=0 $Y2=0
cc_918 N_A_855_368#_c_1230_n N_A_390_81#_c_1913_n 0.00796999f $X=4.815 $Y=1.905
+ $X2=0 $Y2=0
cc_919 N_A_855_368#_c_1232_n N_A_390_81#_c_1913_n 0.013838f $X=4.46 $Y=1.905
+ $X2=0 $Y2=0
cc_920 N_A_855_368#_M1007_g N_A_390_81#_c_1907_n 7.30108e-19 $X=5.19 $Y=0.74
+ $X2=0 $Y2=0
cc_921 N_A_855_368#_c_1206_n N_A_390_81#_c_1907_n 0.00792986f $X=6.12 $Y=1.32
+ $X2=0 $Y2=0
cc_922 N_A_855_368#_M1004_g N_A_390_81#_c_1907_n 0.0107286f $X=6.195 $Y=0.9
+ $X2=0 $Y2=0
cc_923 N_A_855_368#_c_1223_n N_A_390_81#_c_1915_n 0.0038729f $X=6.585 $Y=2.78
+ $X2=0 $Y2=0
cc_924 N_A_855_368#_c_1206_n N_A_390_81#_c_1908_n 0.00824418f $X=6.12 $Y=1.32
+ $X2=0 $Y2=0
cc_925 N_A_855_368#_c_1206_n N_A_390_81#_c_1909_n 0.00689048f $X=6.12 $Y=1.32
+ $X2=0 $Y2=0
cc_926 N_A_855_368#_c_1205_n N_A_390_81#_c_1910_n 0.00311796f $X=5.615 $Y=3.075
+ $X2=0 $Y2=0
cc_927 N_A_855_368#_c_1205_n N_A_390_81#_c_1918_n 0.0102854f $X=5.615 $Y=3.075
+ $X2=0 $Y2=0
cc_928 N_A_855_368#_c_1219_n N_A_390_81#_c_1918_n 0.00419186f $X=6.495 $Y=3.15
+ $X2=0 $Y2=0
cc_929 N_A_855_368#_c_1253_n N_VGND_M1019_d 0.00379589f $X=4.815 $Y=1.005 $X2=0
+ $Y2=0
cc_930 N_A_855_368#_c_1213_n N_VGND_c_2079_n 0.0233464f $X=4.475 $Y=0.515 $X2=0
+ $Y2=0
cc_931 N_A_855_368#_c_1202_n N_VGND_c_2080_n 0.00178148f $X=5.095 $Y=1.765 $X2=0
+ $Y2=0
cc_932 N_A_855_368#_M1007_g N_VGND_c_2080_n 0.00484359f $X=5.19 $Y=0.74 $X2=0
+ $Y2=0
cc_933 N_A_855_368#_c_1213_n N_VGND_c_2080_n 0.0150231f $X=4.475 $Y=0.515 $X2=0
+ $Y2=0
cc_934 N_A_855_368#_c_1253_n N_VGND_c_2080_n 0.0159075f $X=4.815 $Y=1.005 $X2=0
+ $Y2=0
cc_935 N_A_855_368#_c_1216_n N_VGND_c_2080_n 0.00262017f $X=5.14 $Y=1.46 $X2=0
+ $Y2=0
cc_936 N_A_855_368#_M1008_g N_VGND_c_2081_n 0.00155929f $X=10.315 $Y=0.58 $X2=0
+ $Y2=0
cc_937 N_A_855_368#_c_1213_n N_VGND_c_2089_n 0.00749631f $X=4.475 $Y=0.515 $X2=0
+ $Y2=0
cc_938 N_A_855_368#_M1007_g N_VGND_c_2090_n 0.00432683f $X=5.19 $Y=0.74 $X2=0
+ $Y2=0
cc_939 N_A_855_368#_M1008_g N_VGND_c_2091_n 0.00308264f $X=10.315 $Y=0.58 $X2=0
+ $Y2=0
cc_940 N_A_855_368#_M1007_g N_VGND_c_2100_n 0.00821783f $X=5.19 $Y=0.74 $X2=0
+ $Y2=0
cc_941 N_A_855_368#_M1008_g N_VGND_c_2100_n 0.00383744f $X=10.315 $Y=0.58 $X2=0
+ $Y2=0
cc_942 N_A_855_368#_c_1213_n N_VGND_c_2100_n 0.0062048f $X=4.475 $Y=0.515 $X2=0
+ $Y2=0
cc_943 N_A_2082_446#_c_1402_n N_A_1824_74#_M1013_g 0.00761651f $X=11.71 $Y=0.58
+ $X2=0 $Y2=0
cc_944 N_A_2082_446#_c_1404_n N_A_1824_74#_M1013_g 0.00732912f $X=11.875
+ $Y=0.855 $X2=0 $Y2=0
cc_945 N_A_2082_446#_c_1405_n N_A_1824_74#_M1013_g 0.00376832f $X=12.145 $Y=1.58
+ $X2=0 $Y2=0
cc_946 N_A_2082_446#_c_1401_n N_A_1824_74#_c_1535_n 0.0116511f $X=12.06 $Y=1.665
+ $X2=0 $Y2=0
cc_947 N_A_2082_446#_c_1412_n N_A_1824_74#_c_1537_n 0.00502098f $X=11.41
+ $Y=2.475 $X2=0 $Y2=0
cc_948 N_A_2082_446#_c_1413_n N_A_1824_74#_c_1537_n 0.00496874f $X=11.575
+ $Y=2.75 $X2=0 $Y2=0
cc_949 N_A_2082_446#_c_1401_n N_A_1824_74#_c_1522_n 0.00220284f $X=12.06
+ $Y=1.665 $X2=0 $Y2=0
cc_950 N_A_2082_446#_c_1405_n N_A_1824_74#_c_1522_n 0.022644f $X=12.145 $Y=1.58
+ $X2=0 $Y2=0
cc_951 N_A_2082_446#_c_1401_n N_A_1824_74#_c_1523_n 0.00461365f $X=12.06
+ $Y=1.665 $X2=0 $Y2=0
cc_952 N_A_2082_446#_c_1403_n N_A_1824_74#_c_1523_n 0.0054249f $X=12.06 $Y=0.855
+ $X2=0 $Y2=0
cc_953 N_A_2082_446#_c_1404_n N_A_1824_74#_c_1523_n 0.00561111f $X=11.875
+ $Y=0.855 $X2=0 $Y2=0
cc_954 N_A_2082_446#_c_1401_n N_A_1824_74#_c_1524_n 0.00230014f $X=12.06
+ $Y=1.665 $X2=0 $Y2=0
cc_955 N_A_2082_446#_c_1405_n N_A_1824_74#_c_1524_n 0.0017493f $X=12.145 $Y=1.58
+ $X2=0 $Y2=0
cc_956 N_A_2082_446#_c_1402_n N_A_1824_74#_c_1525_n 0.00350124f $X=11.71 $Y=0.58
+ $X2=0 $Y2=0
cc_957 N_A_2082_446#_c_1403_n N_A_1824_74#_c_1525_n 0.00386679f $X=12.06
+ $Y=0.855 $X2=0 $Y2=0
cc_958 N_A_2082_446#_c_1405_n N_A_1824_74#_c_1525_n 0.00324637f $X=12.145
+ $Y=1.58 $X2=0 $Y2=0
cc_959 N_A_2082_446#_c_1401_n N_A_1824_74#_c_1526_n 0.00573299f $X=12.06
+ $Y=1.665 $X2=0 $Y2=0
cc_960 N_A_2082_446#_c_1405_n N_A_1824_74#_c_1526_n 0.00338011f $X=12.145
+ $Y=1.58 $X2=0 $Y2=0
cc_961 N_A_2082_446#_M1009_g N_A_1824_74#_c_1528_n 0.00114145f $X=10.705 $Y=0.58
+ $X2=0 $Y2=0
cc_962 N_A_2082_446#_c_1408_n N_A_1824_74#_c_1540_n 0.00134164f $X=10.5 $Y=2.465
+ $X2=0 $Y2=0
cc_963 N_A_2082_446#_c_1469_p N_A_1824_74#_c_1540_n 0.00258251f $X=10.85
+ $Y=2.475 $X2=0 $Y2=0
cc_964 N_A_2082_446#_M1009_g N_A_1824_74#_c_1529_n 0.00142814f $X=10.705 $Y=0.58
+ $X2=0 $Y2=0
cc_965 N_A_2082_446#_c_1408_n N_A_1824_74#_c_1530_n 3.62386e-19 $X=10.5 $Y=2.465
+ $X2=0 $Y2=0
cc_966 N_A_2082_446#_M1009_g N_A_1824_74#_c_1530_n 0.00172861f $X=10.705 $Y=0.58
+ $X2=0 $Y2=0
cc_967 N_A_2082_446#_c_1409_n N_A_1824_74#_c_1530_n 0.00168467f $X=10.645
+ $Y=2.23 $X2=0 $Y2=0
cc_968 N_A_2082_446#_c_1469_p N_A_1824_74#_c_1530_n 0.0103077f $X=10.85 $Y=2.475
+ $X2=0 $Y2=0
cc_969 N_A_2082_446#_c_1406_n N_A_1824_74#_c_1530_n 0.074835f $X=10.685 $Y=1.535
+ $X2=0 $Y2=0
cc_970 N_A_2082_446#_c_1407_n N_A_1824_74#_c_1530_n 0.0114396f $X=10.685
+ $Y=1.535 $X2=0 $Y2=0
cc_971 N_A_2082_446#_c_1403_n N_A_1824_74#_c_1531_n 0.00108154f $X=12.06
+ $Y=0.855 $X2=0 $Y2=0
cc_972 N_A_2082_446#_c_1404_n N_A_1824_74#_c_1531_n 0.0272174f $X=11.875
+ $Y=0.855 $X2=0 $Y2=0
cc_973 N_A_2082_446#_c_1405_n N_A_1824_74#_c_1531_n 0.0227002f $X=12.145 $Y=1.58
+ $X2=0 $Y2=0
cc_974 N_A_2082_446#_M1009_g N_A_1824_74#_c_1533_n 0.0143673f $X=10.705 $Y=0.58
+ $X2=0 $Y2=0
cc_975 N_A_2082_446#_c_1401_n N_A_1824_74#_c_1533_n 0.00732151f $X=12.06
+ $Y=1.665 $X2=0 $Y2=0
cc_976 N_A_2082_446#_c_1406_n N_A_1824_74#_c_1533_n 0.0224547f $X=10.685
+ $Y=1.535 $X2=0 $Y2=0
cc_977 N_A_2082_446#_c_1407_n N_A_1824_74#_c_1533_n 0.00598209f $X=10.685
+ $Y=1.535 $X2=0 $Y2=0
cc_978 N_A_2082_446#_M1009_g N_A_1824_74#_c_1534_n 0.0019127f $X=10.705 $Y=0.58
+ $X2=0 $Y2=0
cc_979 N_A_2082_446#_c_1401_n N_A_1824_74#_c_1534_n 0.06452f $X=12.06 $Y=1.665
+ $X2=0 $Y2=0
cc_980 N_A_2082_446#_c_1406_n N_A_1824_74#_c_1534_n 0.00326018f $X=10.685
+ $Y=1.535 $X2=0 $Y2=0
cc_981 N_A_2082_446#_c_1407_n N_A_1824_74#_c_1534_n 2.45278e-19 $X=10.685
+ $Y=1.535 $X2=0 $Y2=0
cc_982 N_A_2082_446#_c_1405_n N_A_2492_392#_c_1667_n 0.0135871f $X=12.145
+ $Y=1.58 $X2=0 $Y2=0
cc_983 N_A_2082_446#_c_1401_n N_A_2492_392#_c_1669_n 0.0058056f $X=12.06
+ $Y=1.665 $X2=0 $Y2=0
cc_984 N_A_2082_446#_c_1401_n N_A_2492_392#_c_1670_n 0.00268745f $X=12.06
+ $Y=1.665 $X2=0 $Y2=0
cc_985 N_A_2082_446#_c_1405_n N_A_2492_392#_c_1670_n 0.0131081f $X=12.145
+ $Y=1.58 $X2=0 $Y2=0
cc_986 N_A_2082_446#_c_1412_n N_VPWR_M1015_d 0.00387797f $X=11.41 $Y=2.475 $X2=0
+ $Y2=0
cc_987 N_A_2082_446#_c_1469_p N_VPWR_M1015_d 0.00236476f $X=10.85 $Y=2.475 $X2=0
+ $Y2=0
cc_988 N_A_2082_446#_c_1401_n N_VPWR_c_1732_n 0.0235807f $X=12.06 $Y=1.665 $X2=0
+ $Y2=0
cc_989 N_A_2082_446#_c_1412_n N_VPWR_c_1732_n 0.012314f $X=11.41 $Y=2.475 $X2=0
+ $Y2=0
cc_990 N_A_2082_446#_c_1413_n N_VPWR_c_1732_n 0.0282274f $X=11.575 $Y=2.75 $X2=0
+ $Y2=0
cc_991 N_A_2082_446#_c_1413_n N_VPWR_c_1740_n 0.0144033f $X=11.575 $Y=2.75 $X2=0
+ $Y2=0
cc_992 N_A_2082_446#_c_1408_n N_VPWR_c_1745_n 0.00415318f $X=10.5 $Y=2.465 $X2=0
+ $Y2=0
cc_993 N_A_2082_446#_c_1408_n N_VPWR_c_1751_n 0.00864935f $X=10.5 $Y=2.465 $X2=0
+ $Y2=0
cc_994 N_A_2082_446#_c_1409_n N_VPWR_c_1751_n 0.00123389f $X=10.645 $Y=2.23
+ $X2=0 $Y2=0
cc_995 N_A_2082_446#_c_1412_n N_VPWR_c_1751_n 0.0288765f $X=11.41 $Y=2.475 $X2=0
+ $Y2=0
cc_996 N_A_2082_446#_c_1469_p N_VPWR_c_1751_n 0.0201549f $X=10.85 $Y=2.475 $X2=0
+ $Y2=0
cc_997 N_A_2082_446#_c_1413_n N_VPWR_c_1751_n 0.0102623f $X=11.575 $Y=2.75 $X2=0
+ $Y2=0
cc_998 N_A_2082_446#_c_1408_n N_VPWR_c_1727_n 0.00817239f $X=10.5 $Y=2.465 $X2=0
+ $Y2=0
cc_999 N_A_2082_446#_c_1409_n N_VPWR_c_1727_n 3.19707e-19 $X=10.645 $Y=2.23
+ $X2=0 $Y2=0
cc_1000 N_A_2082_446#_c_1412_n N_VPWR_c_1727_n 0.00667547f $X=11.41 $Y=2.475
+ $X2=0 $Y2=0
cc_1001 N_A_2082_446#_c_1469_p N_VPWR_c_1727_n 0.00116499f $X=10.85 $Y=2.475
+ $X2=0 $Y2=0
cc_1002 N_A_2082_446#_c_1413_n N_VPWR_c_1727_n 0.0119211f $X=11.575 $Y=2.75
+ $X2=0 $Y2=0
cc_1003 N_A_2082_446#_c_1403_n N_VGND_M1030_s 0.00405314f $X=12.06 $Y=0.855
+ $X2=0 $Y2=0
cc_1004 N_A_2082_446#_c_1405_n N_VGND_M1030_s 8.04296e-19 $X=12.145 $Y=1.58
+ $X2=0 $Y2=0
cc_1005 N_A_2082_446#_M1009_g N_VGND_c_2081_n 0.0119771f $X=10.705 $Y=0.58 $X2=0
+ $Y2=0
cc_1006 N_A_2082_446#_c_1402_n N_VGND_c_2081_n 0.0140354f $X=11.71 $Y=0.58 $X2=0
+ $Y2=0
cc_1007 N_A_2082_446#_c_1404_n N_VGND_c_2081_n 0.00142029f $X=11.875 $Y=0.855
+ $X2=0 $Y2=0
cc_1008 N_A_2082_446#_c_1402_n N_VGND_c_2082_n 0.0168546f $X=11.71 $Y=0.58 $X2=0
+ $Y2=0
cc_1009 N_A_2082_446#_c_1403_n N_VGND_c_2082_n 0.0109002f $X=12.06 $Y=0.855
+ $X2=0 $Y2=0
cc_1010 N_A_2082_446#_M1009_g N_VGND_c_2091_n 0.00383152f $X=10.705 $Y=0.58
+ $X2=0 $Y2=0
cc_1011 N_A_2082_446#_c_1402_n N_VGND_c_2092_n 0.014415f $X=11.71 $Y=0.58 $X2=0
+ $Y2=0
cc_1012 N_A_2082_446#_M1009_g N_VGND_c_2100_n 0.0075725f $X=10.705 $Y=0.58 $X2=0
+ $Y2=0
cc_1013 N_A_2082_446#_c_1402_n N_VGND_c_2100_n 0.0119404f $X=11.71 $Y=0.58 $X2=0
+ $Y2=0
cc_1014 N_A_2082_446#_c_1403_n N_VGND_c_2100_n 0.0092009f $X=12.06 $Y=0.855
+ $X2=0 $Y2=0
cc_1015 N_A_1824_74#_c_1539_n N_A_2492_392#_c_1674_n 0.00352637f $X=12.385
+ $Y=1.885 $X2=0 $Y2=0
cc_1016 N_A_1824_74#_c_1527_n N_A_2492_392#_c_1674_n 0.00239754f $X=12.295
+ $Y=1.095 $X2=0 $Y2=0
cc_1017 N_A_1824_74#_c_1539_n N_A_2492_392#_c_1675_n 0.0089495f $X=12.385
+ $Y=1.885 $X2=0 $Y2=0
cc_1018 N_A_1824_74#_c_1525_n N_A_2492_392#_c_1667_n 0.00769864f $X=12.485
+ $Y=1.095 $X2=0 $Y2=0
cc_1019 N_A_1824_74#_c_1527_n N_A_2492_392#_c_1667_n 0.00167437f $X=12.295
+ $Y=1.095 $X2=0 $Y2=0
cc_1020 N_A_1824_74#_c_1524_n N_A_2492_392#_c_1669_n 0.00768781f $X=12.385
+ $Y=1.795 $X2=0 $Y2=0
cc_1021 N_A_1824_74#_c_1539_n N_A_2492_392#_c_1669_n 0.00189951f $X=12.385
+ $Y=1.885 $X2=0 $Y2=0
cc_1022 N_A_1824_74#_c_1527_n N_A_2492_392#_c_1670_n 0.00471821f $X=12.295
+ $Y=1.095 $X2=0 $Y2=0
cc_1023 N_A_1824_74#_c_1527_n N_A_2492_392#_c_1671_n 0.00503519f $X=12.295
+ $Y=1.095 $X2=0 $Y2=0
cc_1024 N_A_1824_74#_c_1536_n N_VPWR_c_1732_n 0.00975077f $X=11.8 $Y=2.375 $X2=0
+ $Y2=0
cc_1025 N_A_1824_74#_c_1537_n N_VPWR_c_1732_n 0.00807257f $X=11.8 $Y=2.465 $X2=0
+ $Y2=0
cc_1026 N_A_1824_74#_c_1522_n N_VPWR_c_1732_n 7.36409e-19 $X=12.295 $Y=1.26
+ $X2=0 $Y2=0
cc_1027 N_A_1824_74#_c_1539_n N_VPWR_c_1732_n 0.00991624f $X=12.385 $Y=1.885
+ $X2=0 $Y2=0
cc_1028 N_A_1824_74#_c_1539_n N_VPWR_c_1733_n 0.00456767f $X=12.385 $Y=1.885
+ $X2=0 $Y2=0
cc_1029 N_A_1824_74#_c_1537_n N_VPWR_c_1740_n 0.00445602f $X=11.8 $Y=2.465 $X2=0
+ $Y2=0
cc_1030 N_A_1824_74#_c_1540_n N_VPWR_c_1745_n 0.019583f $X=10.22 $Y=2.685 $X2=0
+ $Y2=0
cc_1031 N_A_1824_74#_c_1541_n N_VPWR_c_1745_n 0.00812764f $X=9.6 $Y=2.685 $X2=0
+ $Y2=0
cc_1032 N_A_1824_74#_c_1539_n N_VPWR_c_1746_n 0.00445602f $X=12.385 $Y=1.885
+ $X2=0 $Y2=0
cc_1033 N_A_1824_74#_c_1537_n N_VPWR_c_1727_n 0.00896763f $X=11.8 $Y=2.465 $X2=0
+ $Y2=0
cc_1034 N_A_1824_74#_c_1539_n N_VPWR_c_1727_n 0.00862869f $X=12.385 $Y=1.885
+ $X2=0 $Y2=0
cc_1035 N_A_1824_74#_c_1540_n N_VPWR_c_1727_n 0.025422f $X=10.22 $Y=2.685 $X2=0
+ $Y2=0
cc_1036 N_A_1824_74#_c_1541_n N_VPWR_c_1727_n 0.00936382f $X=9.6 $Y=2.685 $X2=0
+ $Y2=0
cc_1037 N_A_1824_74#_c_1540_n A_2037_508# 0.00191616f $X=10.22 $Y=2.685
+ $X2=-0.19 $Y2=-0.245
cc_1038 N_A_1824_74#_M1013_g N_VGND_c_2081_n 0.00182082f $X=11.495 $Y=0.58 $X2=0
+ $Y2=0
cc_1039 N_A_1824_74#_c_1528_n N_VGND_c_2081_n 0.014224f $X=10.22 $Y=0.645 $X2=0
+ $Y2=0
cc_1040 N_A_1824_74#_c_1533_n N_VGND_c_2081_n 0.0229174f $X=11.02 $Y=1.22 $X2=0
+ $Y2=0
cc_1041 N_A_1824_74#_M1013_g N_VGND_c_2082_n 0.00324482f $X=11.495 $Y=0.58 $X2=0
+ $Y2=0
cc_1042 N_A_1824_74#_c_1522_n N_VGND_c_2082_n 0.00356476f $X=12.295 $Y=1.26
+ $X2=0 $Y2=0
cc_1043 N_A_1824_74#_c_1525_n N_VGND_c_2082_n 0.00936719f $X=12.485 $Y=1.095
+ $X2=0 $Y2=0
cc_1044 N_A_1824_74#_c_1525_n N_VGND_c_2083_n 0.00296233f $X=12.485 $Y=1.095
+ $X2=0 $Y2=0
cc_1045 N_A_1824_74#_c_1528_n N_VGND_c_2091_n 0.0249458f $X=10.22 $Y=0.645 $X2=0
+ $Y2=0
cc_1046 N_A_1824_74#_M1013_g N_VGND_c_2092_n 0.00434272f $X=11.495 $Y=0.58 $X2=0
+ $Y2=0
cc_1047 N_A_1824_74#_c_1525_n N_VGND_c_2093_n 0.00383152f $X=12.485 $Y=1.095
+ $X2=0 $Y2=0
cc_1048 N_A_1824_74#_M1013_g N_VGND_c_2100_n 0.00825669f $X=11.495 $Y=0.58 $X2=0
+ $Y2=0
cc_1049 N_A_1824_74#_c_1525_n N_VGND_c_2100_n 0.00762539f $X=12.485 $Y=1.095
+ $X2=0 $Y2=0
cc_1050 N_A_1824_74#_c_1528_n N_VGND_c_2100_n 0.0310203f $X=10.22 $Y=0.645 $X2=0
+ $Y2=0
cc_1051 N_A_2492_392#_c_1674_n N_VPWR_c_1732_n 0.0405667f $X=12.61 $Y=2.105
+ $X2=0 $Y2=0
cc_1052 N_A_2492_392#_c_1672_n N_VPWR_c_1733_n 0.0180379f $X=13.395 $Y=1.765
+ $X2=0 $Y2=0
cc_1053 N_A_2492_392#_c_1673_n N_VPWR_c_1733_n 7.0907e-19 $X=13.845 $Y=1.765
+ $X2=0 $Y2=0
cc_1054 N_A_2492_392#_c_1668_n N_VPWR_c_1733_n 0.025458f $X=13.19 $Y=1.465 $X2=0
+ $Y2=0
cc_1055 N_A_2492_392#_c_1669_n N_VPWR_c_1733_n 0.0777543f $X=12.61 $Y=1.94 $X2=0
+ $Y2=0
cc_1056 N_A_2492_392#_c_1671_n N_VPWR_c_1733_n 0.00689404f $X=13.845 $Y=1.532
+ $X2=0 $Y2=0
cc_1057 N_A_2492_392#_c_1673_n N_VPWR_c_1735_n 0.0260843f $X=13.845 $Y=1.765
+ $X2=0 $Y2=0
cc_1058 N_A_2492_392#_c_1671_n N_VPWR_c_1735_n 9.39066e-19 $X=13.845 $Y=1.532
+ $X2=0 $Y2=0
cc_1059 N_A_2492_392#_c_1675_n N_VPWR_c_1746_n 0.0145938f $X=12.61 $Y=2.815
+ $X2=0 $Y2=0
cc_1060 N_A_2492_392#_c_1672_n N_VPWR_c_1747_n 0.00413917f $X=13.395 $Y=1.765
+ $X2=0 $Y2=0
cc_1061 N_A_2492_392#_c_1673_n N_VPWR_c_1747_n 0.00445602f $X=13.845 $Y=1.765
+ $X2=0 $Y2=0
cc_1062 N_A_2492_392#_c_1672_n N_VPWR_c_1727_n 0.00817726f $X=13.395 $Y=1.765
+ $X2=0 $Y2=0
cc_1063 N_A_2492_392#_c_1673_n N_VPWR_c_1727_n 0.00860566f $X=13.845 $Y=1.765
+ $X2=0 $Y2=0
cc_1064 N_A_2492_392#_c_1675_n N_VPWR_c_1727_n 0.0120466f $X=12.61 $Y=2.815
+ $X2=0 $Y2=0
cc_1065 N_A_2492_392#_c_1672_n N_Q_c_2057_n 0.00196498f $X=13.395 $Y=1.765 $X2=0
+ $Y2=0
cc_1066 N_A_2492_392#_c_1673_n N_Q_c_2057_n 0.0153501f $X=13.845 $Y=1.765 $X2=0
+ $Y2=0
cc_1067 N_A_2492_392#_c_1671_n N_Q_c_2057_n 0.0338785f $X=13.845 $Y=1.532 $X2=0
+ $Y2=0
cc_1068 N_A_2492_392#_M1001_g Q 0.0138248f $X=13.475 $Y=0.74 $X2=0 $Y2=0
cc_1069 N_A_2492_392#_M1031_g Q 0.0162403f $X=13.905 $Y=0.74 $X2=0 $Y2=0
cc_1070 N_A_2492_392#_c_1667_n Q 0.00465944f $X=12.7 $Y=0.515 $X2=0 $Y2=0
cc_1071 N_A_2492_392#_M1001_g Q 0.0018463f $X=13.475 $Y=0.74 $X2=0 $Y2=0
cc_1072 N_A_2492_392#_M1031_g Q 0.00299044f $X=13.905 $Y=0.74 $X2=0 $Y2=0
cc_1073 N_A_2492_392#_c_1668_n Q 0.02585f $X=13.19 $Y=1.465 $X2=0 $Y2=0
cc_1074 N_A_2492_392#_c_1671_n Q 0.015501f $X=13.845 $Y=1.532 $X2=0 $Y2=0
cc_1075 N_A_2492_392#_c_1667_n N_VGND_c_2082_n 0.0101431f $X=12.7 $Y=0.515 $X2=0
+ $Y2=0
cc_1076 N_A_2492_392#_M1001_g N_VGND_c_2083_n 0.00647412f $X=13.475 $Y=0.74
+ $X2=0 $Y2=0
cc_1077 N_A_2492_392#_c_1667_n N_VGND_c_2083_n 0.0505719f $X=12.7 $Y=0.515 $X2=0
+ $Y2=0
cc_1078 N_A_2492_392#_c_1668_n N_VGND_c_2083_n 0.0209147f $X=13.19 $Y=1.465
+ $X2=0 $Y2=0
cc_1079 N_A_2492_392#_c_1671_n N_VGND_c_2083_n 0.0058967f $X=13.845 $Y=1.532
+ $X2=0 $Y2=0
cc_1080 N_A_2492_392#_M1031_g N_VGND_c_2085_n 0.00647412f $X=13.905 $Y=0.74
+ $X2=0 $Y2=0
cc_1081 N_A_2492_392#_c_1667_n N_VGND_c_2093_n 0.0115122f $X=12.7 $Y=0.515 $X2=0
+ $Y2=0
cc_1082 N_A_2492_392#_M1001_g N_VGND_c_2094_n 0.00434272f $X=13.475 $Y=0.74
+ $X2=0 $Y2=0
cc_1083 N_A_2492_392#_M1031_g N_VGND_c_2094_n 0.00434272f $X=13.905 $Y=0.74
+ $X2=0 $Y2=0
cc_1084 N_A_2492_392#_M1001_g N_VGND_c_2100_n 0.00825283f $X=13.475 $Y=0.74
+ $X2=0 $Y2=0
cc_1085 N_A_2492_392#_M1031_g N_VGND_c_2100_n 0.00823942f $X=13.905 $Y=0.74
+ $X2=0 $Y2=0
cc_1086 N_A_2492_392#_c_1667_n N_VGND_c_2100_n 0.0095288f $X=12.7 $Y=0.515 $X2=0
+ $Y2=0
cc_1087 N_VPWR_M1005_d N_A_390_81#_c_1919_n 0.0110121f $X=3.11 $Y=2.32 $X2=0
+ $Y2=0
cc_1088 N_VPWR_c_1728_n N_A_390_81#_c_1919_n 0.0214041f $X=3.26 $Y=2.79 $X2=0
+ $Y2=0
cc_1089 N_VPWR_c_1727_n N_A_390_81#_c_1919_n 0.0231955f $X=14.16 $Y=3.33 $X2=0
+ $Y2=0
cc_1090 N_VPWR_c_1728_n N_A_390_81#_c_1912_n 0.02127f $X=3.26 $Y=2.79 $X2=0
+ $Y2=0
cc_1091 N_VPWR_c_1736_n N_A_390_81#_c_1912_n 0.0166211f $X=4.705 $Y=3.33 $X2=0
+ $Y2=0
cc_1092 N_VPWR_c_1727_n N_A_390_81#_c_1912_n 0.0136307f $X=14.16 $Y=3.33 $X2=0
+ $Y2=0
cc_1093 N_VPWR_M1018_d N_A_390_81#_c_1913_n 0.00463358f $X=4.72 $Y=1.84 $X2=0
+ $Y2=0
cc_1094 N_VPWR_c_1729_n N_A_390_81#_c_1913_n 0.0166996f $X=4.87 $Y=2.815 $X2=0
+ $Y2=0
cc_1095 N_VPWR_c_1727_n N_A_390_81#_c_1913_n 0.0501229f $X=14.16 $Y=3.33 $X2=0
+ $Y2=0
cc_1096 N_VPWR_M1005_d N_A_390_81#_c_1914_n 8.56696e-19 $X=3.11 $Y=2.32 $X2=0
+ $Y2=0
cc_1097 N_VPWR_c_1727_n N_A_390_81#_c_1914_n 0.00615626f $X=14.16 $Y=3.33 $X2=0
+ $Y2=0
cc_1098 N_VPWR_c_1728_n N_A_390_81#_c_1917_n 0.00713257f $X=3.26 $Y=2.79 $X2=0
+ $Y2=0
cc_1099 N_VPWR_c_1743_n N_A_390_81#_c_1917_n 0.0144799f $X=3.095 $Y=3.33 $X2=0
+ $Y2=0
cc_1100 N_VPWR_c_1748_n N_A_390_81#_c_1917_n 0.0198341f $X=1.4 $Y=2.465 $X2=0
+ $Y2=0
cc_1101 N_VPWR_c_1727_n N_A_390_81#_c_1917_n 0.0119509f $X=14.16 $Y=3.33 $X2=0
+ $Y2=0
cc_1102 N_VPWR_c_1738_n N_A_390_81#_c_1918_n 0.00528674f $X=7.15 $Y=3.33 $X2=0
+ $Y2=0
cc_1103 N_VPWR_c_1727_n N_A_390_81#_c_1918_n 0.00666438f $X=14.16 $Y=3.33 $X2=0
+ $Y2=0
cc_1104 N_VPWR_c_1733_n N_Q_c_2057_n 0.0412253f $X=13.17 $Y=1.985 $X2=0 $Y2=0
cc_1105 N_VPWR_c_1735_n N_Q_c_2057_n 0.0435456f $X=14.12 $Y=1.985 $X2=0 $Y2=0
cc_1106 N_VPWR_c_1747_n N_Q_c_2057_n 0.0114703f $X=13.955 $Y=3.33 $X2=0 $Y2=0
cc_1107 N_VPWR_c_1727_n N_Q_c_2057_n 0.00946127f $X=14.16 $Y=3.33 $X2=0 $Y2=0
cc_1108 N_A_390_81#_c_1919_n A_514_464# 0.013941f $X=3.445 $Y=2.43 $X2=-0.19
+ $Y2=-0.245
cc_1109 N_A_390_81#_M1011_d N_noxref_24_c_2215_n 0.0099946f $X=1.95 $Y=0.405
+ $X2=0 $Y2=0
cc_1110 N_A_390_81#_c_1902_n N_noxref_24_c_2215_n 0.0420252f $X=2.875 $Y=0.72
+ $X2=0 $Y2=0
cc_1111 N_A_390_81#_c_1902_n N_noxref_24_c_2216_n 0.0206309f $X=2.875 $Y=0.72
+ $X2=0 $Y2=0
cc_1112 N_A_390_81#_c_1904_n N_noxref_24_c_2216_n 0.0190079f $X=3.445 $Y=1.225
+ $X2=0 $Y2=0
cc_1113 N_A_390_81#_c_1902_n noxref_26 0.00129814f $X=2.875 $Y=0.72 $X2=-0.19
+ $Y2=-0.245
cc_1114 Q N_VGND_c_2083_n 0.0294122f $X=13.595 $Y=0.47 $X2=0 $Y2=0
cc_1115 Q N_VGND_c_2085_n 0.0294122f $X=13.595 $Y=0.47 $X2=0 $Y2=0
cc_1116 Q N_VGND_c_2094_n 0.0144922f $X=13.595 $Y=0.47 $X2=0 $Y2=0
cc_1117 Q N_VGND_c_2100_n 0.0118826f $X=13.595 $Y=0.47 $X2=0 $Y2=0
cc_1118 N_VGND_c_2079_n N_noxref_24_c_2215_n 0.0134774f $X=3.88 $Y=0.615 $X2=0
+ $Y2=0
cc_1119 N_VGND_c_2086_n N_noxref_24_c_2215_n 0.138041f $X=3.715 $Y=0 $X2=0 $Y2=0
cc_1120 N_VGND_c_2100_n N_noxref_24_c_2215_n 0.0797026f $X=14.16 $Y=0 $X2=0
+ $Y2=0
cc_1121 N_VGND_c_2079_n N_noxref_24_c_2216_n 0.0165124f $X=3.88 $Y=0.615 $X2=0
+ $Y2=0
cc_1122 N_VGND_c_2078_n N_noxref_24_c_2217_n 0.0259561f $X=0.71 $Y=0.555 $X2=0
+ $Y2=0
cc_1123 N_VGND_c_2086_n N_noxref_24_c_2217_n 0.0225398f $X=3.715 $Y=0 $X2=0
+ $Y2=0
cc_1124 N_VGND_c_2100_n N_noxref_24_c_2217_n 0.0125704f $X=14.16 $Y=0 $X2=0
+ $Y2=0
cc_1125 N_noxref_24_c_2215_n noxref_25 0.00198134f $X=3.215 $Y=0.34 $X2=-0.19
+ $Y2=-0.245
cc_1126 N_noxref_24_c_2215_n noxref_26 0.00134156f $X=3.215 $Y=0.34 $X2=-0.19
+ $Y2=-0.245
