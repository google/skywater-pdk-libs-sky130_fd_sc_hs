/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */

`ifndef SKY130_FD_SC_HS__UDP_ISOLATCH_PP_PKG_S_TB_V
`define SKY130_FD_SC_HS__UDP_ISOLATCH_PP_PKG_S_TB_V

/**
 * udp_isolatch_pp$PKG$s: Power isolating latch. Includes VPWR, KAPWR,
 *                        and VGND power pins with active low sleep
 *                        pin (SLEEP_B).
 *
 * Autogenerated test bench.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none

`include "sky130_fd_sc_hs__udp_isolatch_pp_pkg_s.v"

module top();

    // Inputs are registered
    reg D;
    reg SLEEP_B;
    reg KAPWR;
    reg VGND;
    reg VPWR;

    // Outputs are wires
    wire Q;

    initial
    begin
        // Initial state is x for all inputs.
        D       = 1'bX;
        KAPWR   = 1'bX;
        SLEEP_B = 1'bX;
        VGND    = 1'bX;
        VPWR    = 1'bX;

        #20   D       = 1'b0;
        #40   KAPWR   = 1'b0;
        #60   SLEEP_B = 1'b0;
        #80   VGND    = 1'b0;
        #100  VPWR    = 1'b0;
        #120  D       = 1'b1;
        #140  KAPWR   = 1'b1;
        #160  SLEEP_B = 1'b1;
        #180  VGND    = 1'b1;
        #200  VPWR    = 1'b1;
        #220  D       = 1'b0;
        #240  KAPWR   = 1'b0;
        #260  SLEEP_B = 1'b0;
        #280  VGND    = 1'b0;
        #300  VPWR    = 1'b0;
        #320  VPWR    = 1'b1;
        #340  VGND    = 1'b1;
        #360  SLEEP_B = 1'b1;
        #380  KAPWR   = 1'b1;
        #400  D       = 1'b1;
        #420  VPWR    = 1'bx;
        #440  VGND    = 1'bx;
        #460  SLEEP_B = 1'bx;
        #480  KAPWR   = 1'bx;
        #500  D       = 1'bx;
    end

    sky130_fd_sc_hs__udp_isolatch_pp$PKG$s dut (.D(D), .SLEEP_B(SLEEP_B), .KAPWR(KAPWR), .VGND(VGND), .VPWR(VPWR), .Q(Q));

endmodule

`default_nettype wire
`endif  // SKY130_FD_SC_HS__UDP_ISOLATCH_PP_PKG_S_TB_V
