# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_hs__and4bb_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__and4bb_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.800000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A_N
    ANTENNAGATEAREA  0.208500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105000 1.300000 0.400000 1.780000 ;
    END
  END A_N
  PIN B_N
    ANTENNAGATEAREA  0.208500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.400000 1.300000 4.695000 1.780000 ;
    END
  END B_N
  PIN C
    ANTENNAGATEAREA  0.222000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.015000 1.190000 3.345000 1.860000 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  0.222000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.515000 1.190000 3.890000 1.860000 ;
    END
  END D
  PIN X
    ANTENNADIFFAREA  0.692500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.910000 0.960000 1.270000 1.130000 ;
        RECT 0.910000 1.130000 1.080000 1.820000 ;
        RECT 0.910000 1.820000 1.565000 2.150000 ;
        RECT 1.080000 0.350000 1.270000 0.960000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 4.800000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 4.800000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.800000 0.085000 ;
      RECT 0.000000  3.245000 4.800000 3.415000 ;
      RECT 0.115000  0.350000 0.365000 0.960000 ;
      RECT 0.115000  0.960000 0.740000 1.130000 ;
      RECT 0.115000  1.950000 0.740000 2.320000 ;
      RECT 0.115000  2.320000 2.045000 2.490000 ;
      RECT 0.115000  2.490000 0.445000 2.700000 ;
      RECT 0.545000  0.085000 0.875000 0.790000 ;
      RECT 0.570000  1.130000 0.740000 1.950000 ;
      RECT 0.650000  2.660000 0.980000 3.245000 ;
      RECT 1.250000  1.300000 1.610000 1.630000 ;
      RECT 1.440000  0.860000 2.385000 1.030000 ;
      RECT 1.440000  1.030000 1.610000 1.300000 ;
      RECT 1.780000  1.290000 2.045000 2.320000 ;
      RECT 1.795000  2.660000 2.125000 3.245000 ;
      RECT 1.820000  0.350000 2.385000 0.860000 ;
      RECT 2.215000  1.030000 2.385000 2.030000 ;
      RECT 2.215000  2.030000 3.625000 2.200000 ;
      RECT 2.295000  2.200000 2.625000 2.980000 ;
      RECT 2.555000  0.850000 4.685000 1.020000 ;
      RECT 2.555000  1.020000 2.845000 1.790000 ;
      RECT 2.795000  2.370000 3.125000 3.245000 ;
      RECT 3.295000  2.200000 3.625000 2.980000 ;
      RECT 3.720000  0.085000 4.110000 0.680000 ;
      RECT 3.815000  2.290000 4.145000 3.245000 ;
      RECT 4.060000  1.020000 4.685000 1.030000 ;
      RECT 4.060000  1.030000 4.230000 1.950000 ;
      RECT 4.060000  1.950000 4.645000 2.120000 ;
      RECT 4.315000  2.120000 4.645000 2.980000 ;
      RECT 4.355000  0.440000 4.685000 0.850000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
  END
END sky130_fd_sc_hs__and4bb_1
END LIBRARY
