* File: sky130_fd_sc_hs__o2bb2ai_1.spice
* Created: Thu Aug 27 21:01:13 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hs__o2bb2ai_1.pex.spice"
.subckt sky130_fd_sc_hs__o2bb2ai_1  VNB VPB A1_N A2_N B2 B1 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* B1	B1
* B2	B2
* A2_N	A2_N
* A1_N	A1_N
* VPB	VPB
* VNB	VNB
MM1007 A_114_74# N_A1_N_M1007_g N_VGND_M1007_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.0768 AS=0.1824 PD=0.88 PS=1.85 NRD=12.18 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75000.6 A=0.096 P=1.58 MULT=1
MM1003 N_A_131_383#_M1003_d N_A2_N_M1003_g A_114_74# VNB NLOWVT L=0.15 W=0.64
+ AD=0.1824 AS=0.0768 PD=1.85 PS=0.88 NRD=0 NRS=12.18 M=1 R=4.26667 SA=75000.6
+ SB=75000.2 A=0.096 P=1.58 MULT=1
MM1006 N_A_397_74#_M1006_d N_A_131_383#_M1006_g N_Y_M1006_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1295 AS=0.2109 PD=1.09 PS=2.05 NRD=11.34 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75001.1 A=0.111 P=1.78 MULT=1
MM1005 N_VGND_M1005_d N_B2_M1005_g N_A_397_74#_M1006_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1295 PD=1.02 PS=1.09 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.7
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1001 N_A_397_74#_M1001_d N_B1_M1001_g N_VGND_M1005_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.1036 PD=2.05 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.1
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1008 N_A_131_383#_M1008_d N_A1_N_M1008_g N_VPWR_M1008_s VPB PSHORT L=0.15
+ W=0.84 AD=0.126 AS=0.2898 PD=1.14 PS=2.37 NRD=2.3443 NRS=14.0658 M=1 R=5.6
+ SA=75000.3 SB=75002.5 A=0.126 P=1.98 MULT=1
MM1002 N_VPWR_M1002_d N_A2_N_M1002_g N_A_131_383#_M1008_d VPB PSHORT L=0.15
+ W=0.84 AD=0.318011 AS=0.126 PD=1.59857 PS=1.14 NRD=42.5914 NRS=2.3443 M=1
+ R=5.6 SA=75000.7 SB=75002 A=0.126 P=1.98 MULT=1
MM1009 N_Y_M1009_d N_A_131_383#_M1009_g N_VPWR_M1002_d VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.424014 PD=1.42 PS=2.13143 NRD=1.7533 NRS=29.5894 M=1 R=7.46667
+ SA=75001.3 SB=75001.1 A=0.168 P=2.54 MULT=1
MM1000 A_490_368# N_B2_M1000_g N_Y_M1009_d VPB PSHORT L=0.15 W=1.12 AD=0.1848
+ AS=0.168 PD=1.45 PS=1.42 NRD=19.3454 NRS=1.7533 M=1 R=7.46667 SA=75001.7
+ SB=75000.7 A=0.168 P=2.54 MULT=1
MM1004 N_VPWR_M1004_d N_B1_M1004_g A_490_368# VPB PSHORT L=0.15 W=1.12 AD=0.3304
+ AS=0.1848 PD=2.83 PS=1.45 NRD=1.7533 NRS=19.3454 M=1 R=7.46667 SA=75002.2
+ SB=75000.2 A=0.168 P=2.54 MULT=1
DX10_noxref VNB VPB NWDIODE A=6.9564 P=11.2
*
.include "sky130_fd_sc_hs__o2bb2ai_1.pxi.spice"
*
.ends
*
*
