* File: sky130_fd_sc_hs__sdfbbn_1.pex.spice
* Created: Thu Aug 27 21:07:51 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HS__SDFBBN_1%SCD 2 4 5 7 10 12 13 16 17
c34 5 0 8.80698e-20 $X=0.505 $Y=2.245
r35 16 18 45.1558 $w=3.75e-07 $l=1.65e-07 $layer=POLY_cond $X=0.407 $Y=1.37
+ $X2=0.407 $Y2=1.205
r36 16 17 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.385
+ $Y=1.37 $X2=0.385 $Y2=1.37
r37 13 17 2.58853 $w=6.68e-07 $l=1.45e-07 $layer=LI1_cond $X=0.24 $Y=1.54
+ $X2=0.385 $Y2=1.54
r38 10 18 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=0.52 $Y=0.805 $X2=0.52
+ $Y2=1.205
r39 5 7 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=0.505 $Y=2.245
+ $X2=0.505 $Y2=2.64
r40 4 5 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=0.505 $Y=2.155 $X2=0.505
+ $Y2=2.245
r41 4 12 108.839 $w=1.8e-07 $l=2.8e-07 $layer=POLY_cond $X=0.505 $Y=2.155
+ $X2=0.505 $Y2=1.875
r42 2 12 42.8297 $w=3.75e-07 $l=1.87e-07 $layer=POLY_cond $X=0.407 $Y=1.688
+ $X2=0.407 $Y2=1.875
r43 1 16 3.26277 $w=3.75e-07 $l=2.2e-08 $layer=POLY_cond $X=0.407 $Y=1.392
+ $X2=0.407 $Y2=1.37
r44 1 2 43.8991 $w=3.75e-07 $l=2.96e-07 $layer=POLY_cond $X=0.407 $Y=1.392
+ $X2=0.407 $Y2=1.688
.ends

.subckt PM_SKY130_FD_SC_HS__SDFBBN_1%D 3 8 10 11 12 18
c60 12 0 1.09771e-19 $X=1.68 $Y=1.665
r61 16 18 34.9723 $w=3.3e-07 $l=2e-07 $layer=POLY_cond $X=1.45 $Y=1.645 $X2=1.65
+ $Y2=1.645
r62 14 16 5.24584 $w=3.3e-07 $l=3e-08 $layer=POLY_cond $X=1.42 $Y=1.645 $X2=1.45
+ $Y2=1.645
r63 12 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.65
+ $Y=1.645 $X2=1.65 $Y2=1.645
r64 10 11 56.6305 $w=1.65e-07 $l=1.3e-07 $layer=POLY_cond $X=1.412 $Y=2.115
+ $X2=1.412 $Y2=2.245
r65 6 16 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.45 $Y=1.48
+ $X2=1.45 $Y2=1.645
r66 6 8 346.117 $w=1.5e-07 $l=6.75e-07 $layer=POLY_cond $X=1.45 $Y=1.48 $X2=1.45
+ $Y2=0.805
r67 4 14 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.42 $Y=1.81
+ $X2=1.42 $Y2=1.645
r68 4 10 156.394 $w=1.5e-07 $l=3.05e-07 $layer=POLY_cond $X=1.42 $Y=1.81
+ $X2=1.42 $Y2=2.115
r69 3 11 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=1.405 $Y=2.64
+ $X2=1.405 $Y2=2.245
.ends

.subckt PM_SKY130_FD_SC_HS__SDFBBN_1%A_353_93# 1 2 7 9 10 12 14 16 19 21 24 27
+ 35 38 41 42
c90 21 0 5.50415e-20 $X=1.855 $Y=2.147
c91 19 0 1.66897e-19 $X=2.13 $Y=1.165
r92 41 42 8.51103 $w=3.58e-07 $l=1.65e-07 $layer=LI1_cond $X=3.07 $Y=2.465
+ $X2=3.07 $Y2=2.3
r93 37 38 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=2.895 $Y=1.645
+ $X2=2.975 $Y2=1.645
r94 34 37 7.68295 $w=3.28e-07 $l=2.2e-07 $layer=LI1_cond $X=2.675 $Y=1.645
+ $X2=2.895 $Y2=1.645
r95 34 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.675
+ $Y=1.645 $X2=2.675 $Y2=1.645
r96 29 38 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.975 $Y=1.81
+ $X2=2.975 $Y2=1.645
r97 29 42 31.9679 $w=1.68e-07 $l=4.9e-07 $layer=LI1_cond $X=2.975 $Y=1.81
+ $X2=2.975 $Y2=2.3
r98 25 37 0.716491 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=2.895 $Y=1.48
+ $X2=2.895 $Y2=1.645
r99 25 27 23.2235 $w=3.28e-07 $l=6.65e-07 $layer=LI1_cond $X=2.895 $Y=1.48
+ $X2=2.895 $Y2=0.815
r100 23 35 82.1848 $w=3.3e-07 $l=4.7e-07 $layer=POLY_cond $X=2.205 $Y=1.645
+ $X2=2.675 $Y2=1.645
r101 23 24 5.03009 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=2.205 $Y=1.645
+ $X2=2.13 $Y2=1.645
r102 21 22 78.8988 $w=1.68e-07 $l=2.75e-07 $layer=POLY_cond $X=1.855 $Y=2.147
+ $X2=2.13 $Y2=2.147
r103 17 19 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=1.84 $Y=1.165
+ $X2=2.13 $Y2=1.165
r104 16 22 5.52526 $w=1.5e-07 $l=9.7e-08 $layer=POLY_cond $X=2.13 $Y=2.05
+ $X2=2.13 $Y2=2.147
r105 15 24 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.13 $Y=1.81
+ $X2=2.13 $Y2=1.645
r106 15 16 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=2.13 $Y=1.81
+ $X2=2.13 $Y2=2.05
r107 14 24 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.13 $Y=1.48
+ $X2=2.13 $Y2=1.645
r108 13 19 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.13 $Y=1.24
+ $X2=2.13 $Y2=1.165
r109 13 14 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=2.13 $Y=1.24
+ $X2=2.13 $Y2=1.48
r110 10 21 5.52526 $w=1.5e-07 $l=9.8e-08 $layer=POLY_cond $X=1.855 $Y=2.245
+ $X2=1.855 $Y2=2.147
r111 10 12 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=1.855 $Y=2.245
+ $X2=1.855 $Y2=2.64
r112 7 17 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.84 $Y=1.09
+ $X2=1.84 $Y2=1.165
r113 7 9 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=1.84 $Y=1.09 $X2=1.84
+ $Y2=0.805
r114 2 41 300 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=2 $X=2.935
+ $Y=2.32 $X2=3.085 $Y2=2.465
r115 1 27 182 $w=1.7e-07 $l=2.81425e-07 $layer=licon1_NDIFF $count=1 $X=2.755
+ $Y=0.595 $X2=2.895 $Y2=0.815
.ends

.subckt PM_SKY130_FD_SC_HS__SDFBBN_1%SCE 4 6 7 9 10 11 15 16 17 18 20 22 25 26
+ 27 29 32
c105 32 0 8.1544e-20 $X=0.97 $Y=1.37
c106 4 0 2.95072e-20 $X=0.91 $Y=0.805
r107 32 33 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.97
+ $Y=1.37 $X2=0.97 $Y2=1.37
r108 29 33 4.10594 $w=6.68e-07 $l=2.3e-07 $layer=LI1_cond $X=1.2 $Y=1.54
+ $X2=0.97 $Y2=1.54
r109 27 28 85.1437 $w=1.67e-07 $l=2.95e-07 $layer=POLY_cond $X=2.86 $Y=2.147
+ $X2=3.155 $Y2=2.147
r110 25 32 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=0.97 $Y=1.71
+ $X2=0.97 $Y2=1.37
r111 25 26 35.4289 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.97 $Y=1.71
+ $X2=0.97 $Y2=1.875
r112 24 32 41.8716 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.97 $Y=1.205
+ $X2=0.97 $Y2=1.37
r113 22 28 5.38489 $w=1.5e-07 $l=9.7e-08 $layer=POLY_cond $X=3.155 $Y=2.05
+ $X2=3.155 $Y2=2.147
r114 21 22 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=3.155 $Y=1.24
+ $X2=3.155 $Y2=2.05
r115 18 27 5.38489 $w=1.5e-07 $l=9.8e-08 $layer=POLY_cond $X=2.86 $Y=2.245
+ $X2=2.86 $Y2=2.147
r116 18 20 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=2.86 $Y=2.245
+ $X2=2.86 $Y2=2.64
r117 16 21 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.08 $Y=1.165
+ $X2=3.155 $Y2=1.24
r118 16 17 166.649 $w=1.5e-07 $l=3.25e-07 $layer=POLY_cond $X=3.08 $Y=1.165
+ $X2=2.755 $Y2=1.165
r119 13 17 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.68 $Y=1.09
+ $X2=2.755 $Y2=1.165
r120 13 15 146.138 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=2.68 $Y=1.09
+ $X2=2.68 $Y2=0.805
r121 12 15 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=2.68 $Y=0.255
+ $X2=2.68 $Y2=0.805
r122 10 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.605 $Y=0.18
+ $X2=2.68 $Y2=0.255
r123 10 11 830.681 $w=1.5e-07 $l=1.62e-06 $layer=POLY_cond $X=2.605 $Y=0.18
+ $X2=0.985 $Y2=0.18
r124 7 9 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=0.985 $Y=2.245
+ $X2=0.985 $Y2=2.64
r125 6 7 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=0.985 $Y=2.155
+ $X2=0.985 $Y2=2.245
r126 6 26 108.839 $w=1.8e-07 $l=2.8e-07 $layer=POLY_cond $X=0.985 $Y=2.155
+ $X2=0.985 $Y2=1.875
r127 4 24 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=0.91 $Y=0.805 $X2=0.91
+ $Y2=1.205
r128 1 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.91 $Y=0.255
+ $X2=0.985 $Y2=0.18
r129 1 4 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=0.91 $Y=0.255
+ $X2=0.91 $Y2=0.805
.ends

.subckt PM_SKY130_FD_SC_HS__SDFBBN_1%CLK_N 3 5 7 8 12
c39 5 0 1.13441e-19 $X=3.87 $Y=1.765
c40 3 0 1.60531e-19 $X=3.67 $Y=0.78
r41 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.635
+ $Y=1.515 $X2=3.635 $Y2=1.515
r42 8 12 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=3.635 $Y=1.665
+ $X2=3.635 $Y2=1.515
r43 5 11 49.7466 $w=4.26e-07 $l=3.18198e-07 $layer=POLY_cond $X=3.87 $Y=1.765
+ $X2=3.715 $Y2=1.515
r44 5 7 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.87 $Y=1.765
+ $X2=3.87 $Y2=2.4
r45 1 11 40.1292 $w=4.26e-07 $l=1.86145e-07 $layer=POLY_cond $X=3.67 $Y=1.35
+ $X2=3.715 $Y2=1.515
r46 1 3 292.277 $w=1.5e-07 $l=5.7e-07 $layer=POLY_cond $X=3.67 $Y=1.35 $X2=3.67
+ $Y2=0.78
.ends

.subckt PM_SKY130_FD_SC_HS__SDFBBN_1%A_977_243# 1 2 3 12 13 14 16 19 23 25 27 28
+ 29 31 33 36 38 39 42 44 45 49 53 57 58 64 65 67 70 74
c200 57 0 7.19434e-20 $X=5.05 $Y=2.13
c201 53 0 1.7536e-19 $X=9.365 $Y=1.795
c202 42 0 1.77523e-19 $X=7.845 $Y=2.31
c203 31 0 1.02525e-19 $X=5.05 $Y=2.145
c204 29 0 1.49471e-19 $X=5.05 $Y=1.755
c205 25 0 1.74547e-19 $X=9.44 $Y=2.045
c206 19 0 8.96875e-20 $X=5.68 $Y=0.805
r207 72 74 3.904 $w=2.5e-07 $l=8e-08 $layer=LI1_cond $X=8.662 $Y=2.395 $X2=8.662
+ $Y2=2.475
r208 71 72 8.784 $w=2.5e-07 $l=1.8e-07 $layer=LI1_cond $X=8.662 $Y=2.215
+ $X2=8.662 $Y2=2.395
r209 67 69 10.5575 $w=3.28e-07 $l=2.25e-07 $layer=LI1_cond $X=7.925 $Y=0.855
+ $X2=7.925 $Y2=1.08
r210 63 65 8.89604 $w=4.23e-07 $l=1.7e-07 $layer=LI1_cond $X=7.335 $Y=2.862
+ $X2=7.505 $Y2=2.862
r211 63 64 15.404 $w=4.23e-07 $l=4.1e-07 $layer=LI1_cond $X=7.335 $Y=2.862
+ $X2=6.925 $Y2=2.862
r212 57 60 3.47907 $w=2.63e-07 $l=8e-08 $layer=LI1_cond $X=5.082 $Y=2.13
+ $X2=5.082 $Y2=2.21
r213 57 58 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.05
+ $Y=2.13 $X2=5.05 $Y2=2.13
r214 53 54 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.365
+ $Y=1.795 $X2=9.365 $Y2=1.795
r215 51 53 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=9.365 $Y=2.13
+ $X2=9.365 $Y2=1.795
r216 50 71 2.99516 $w=1.7e-07 $l=1.68e-07 $layer=LI1_cond $X=8.83 $Y=2.215
+ $X2=8.662 $Y2=2.215
r217 49 51 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=9.2 $Y=2.215
+ $X2=9.365 $Y2=2.13
r218 49 50 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=9.2 $Y=2.215
+ $X2=8.83 $Y2=2.215
r219 46 70 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.93 $Y=2.395
+ $X2=7.845 $Y2=2.395
r220 45 72 2.99516 $w=1.7e-07 $l=1.67e-07 $layer=LI1_cond $X=8.495 $Y=2.395
+ $X2=8.662 $Y2=2.395
r221 45 46 36.861 $w=1.68e-07 $l=5.65e-07 $layer=LI1_cond $X=8.495 $Y=2.395
+ $X2=7.93 $Y2=2.395
r222 43 70 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.845 $Y=2.48
+ $X2=7.845 $Y2=2.395
r223 43 44 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=7.845 $Y=2.48
+ $X2=7.845 $Y2=2.65
r224 42 70 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.845 $Y=2.31
+ $X2=7.845 $Y2=2.395
r225 42 69 80.246 $w=1.68e-07 $l=1.23e-06 $layer=LI1_cond $X=7.845 $Y=2.31
+ $X2=7.845 $Y2=1.08
r226 39 44 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.76 $Y=2.735
+ $X2=7.845 $Y2=2.65
r227 39 65 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=7.76 $Y=2.735
+ $X2=7.505 $Y2=2.735
r228 38 64 85.7914 $w=1.68e-07 $l=1.315e-06 $layer=LI1_cond $X=5.61 $Y=2.99
+ $X2=6.925 $Y2=2.99
r229 36 38 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.525 $Y=2.905
+ $X2=5.61 $Y2=2.99
r230 35 36 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=5.525 $Y=2.295
+ $X2=5.525 $Y2=2.905
r231 34 60 3.33486 $w=1.7e-07 $l=1.33e-07 $layer=LI1_cond $X=5.215 $Y=2.21
+ $X2=5.082 $Y2=2.21
r232 33 35 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.44 $Y=2.21
+ $X2=5.525 $Y2=2.295
r233 33 34 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=5.44 $Y=2.21
+ $X2=5.215 $Y2=2.21
r234 31 58 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=5.05 $Y=2.145
+ $X2=5.05 $Y2=2.13
r235 31 32 71.7872 $w=1.88e-07 $l=2.8e-07 $layer=POLY_cond $X=5.05 $Y=2.277
+ $X2=5.33 $Y2=2.277
r236 28 58 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=5.05 $Y=1.92
+ $X2=5.05 $Y2=2.13
r237 28 29 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.05 $Y=1.92
+ $X2=5.05 $Y2=1.755
r238 25 54 52.2586 $w=2.99e-07 $l=2.85044e-07 $layer=POLY_cond $X=9.44 $Y=2.045
+ $X2=9.365 $Y2=1.795
r239 25 27 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=9.44 $Y=2.045
+ $X2=9.44 $Y2=2.54
r240 21 54 38.5562 $w=2.99e-07 $l=1.92678e-07 $layer=POLY_cond $X=9.305 $Y=1.63
+ $X2=9.365 $Y2=1.795
r241 21 23 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=9.305 $Y=1.63
+ $X2=9.305 $Y2=0.87
r242 17 19 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=5.68 $Y=1.215
+ $X2=5.68 $Y2=0.805
r243 14 32 8.14712 $w=1.5e-07 $l=1.33e-07 $layer=POLY_cond $X=5.33 $Y=2.41
+ $X2=5.33 $Y2=2.277
r244 14 16 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=5.33 $Y=2.41
+ $X2=5.33 $Y2=2.695
r245 12 17 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.605 $Y=1.29
+ $X2=5.68 $Y2=1.215
r246 12 13 292.277 $w=1.5e-07 $l=5.7e-07 $layer=POLY_cond $X=5.605 $Y=1.29
+ $X2=5.035 $Y2=1.29
r247 10 13 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.96 $Y=1.365
+ $X2=5.035 $Y2=1.29
r248 10 29 199.979 $w=1.5e-07 $l=3.9e-07 $layer=POLY_cond $X=4.96 $Y=1.365
+ $X2=4.96 $Y2=1.755
r249 3 74 300 $w=1.7e-07 $l=4.23409e-07 $layer=licon1_PDIFF $count=2 $X=8.51
+ $Y=2.12 $X2=8.66 $Y2=2.475
r250 2 63 600 $w=1.7e-07 $l=8.00125e-07 $layer=licon1_PDIFF $count=1 $X=7.025
+ $Y=2.12 $X2=7.335 $Y2=2.78
r251 1 67 182 $w=1.7e-07 $l=3.60555e-07 $layer=licon1_NDIFF $count=1 $X=7.685
+ $Y=0.595 $X2=7.925 $Y2=0.855
.ends

.subckt PM_SKY130_FD_SC_HS__SDFBBN_1%A_867_82# 1 2 8 9 11 14 16 18 21 23 26 28
+ 31 36 38 39 45 46 47 50 51 57 58 61 76 77
c221 77 0 1.02525e-19 $X=5.755 $Y=1.727
c222 26 0 1.13441e-19 $X=4.58 $Y=2.04
c223 23 0 1.60531e-19 $X=4.61 $Y=1.045
c224 21 0 3.18534e-20 $X=10.745 $Y=0.805
c225 16 0 1.23448e-20 $X=9.83 $Y=2.045
c226 14 0 2.29882e-20 $X=6.47 $Y=0.805
r227 61 63 20.6118 $w=3.04e-07 $l=1.3e-07 $layer=POLY_cond $X=5.59 $Y=1.74
+ $X2=5.72 $Y2=1.74
r228 58 68 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.905
+ $Y=1.775 $X2=9.905 $Y2=1.775
r229 57 58 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.84 $Y=1.665
+ $X2=9.84 $Y2=1.665
r230 54 77 8.65129 $w=3.53e-07 $l=2.35e-07 $layer=LI1_cond $X=5.52 $Y=1.727
+ $X2=5.755 $Y2=1.727
r231 54 76 6.8759 $w=3.53e-07 $l=1.15e-07 $layer=LI1_cond $X=5.52 $Y=1.727
+ $X2=5.405 $Y2=1.727
r232 54 61 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.59
+ $Y=1.74 $X2=5.59 $Y2=1.74
r233 53 54 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=1.665
+ $X2=5.52 $Y2=1.665
r234 51 53 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.665 $Y=1.665
+ $X2=5.52 $Y2=1.665
r235 50 57 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=9.695 $Y=1.665
+ $X2=9.84 $Y2=1.665
r236 50 51 4.98761 $w=1.4e-07 $l=4.03e-06 $layer=MET1_cond $X=9.695 $Y=1.665
+ $X2=5.665 $Y2=1.665
r237 49 58 3.67446 $w=3.43e-07 $l=1.1e-07 $layer=LI1_cond $X=9.897 $Y=1.555
+ $X2=9.897 $Y2=1.665
r238 47 77 28.8111 $w=2.48e-07 $l=6.25e-07 $layer=LI1_cond $X=6.38 $Y=1.675
+ $X2=5.755 $Y2=1.675
r239 46 65 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.545 $Y=1.635
+ $X2=6.545 $Y2=1.47
r240 45 47 6.46688 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=6.545 $Y=1.635
+ $X2=6.38 $Y2=1.635
r241 45 46 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.545
+ $Y=1.635 $X2=6.545 $Y2=1.635
r242 41 43 16.9064 $w=2.67e-07 $l=3.7e-07 $layer=LI1_cond $X=4.61 $Y=1.635
+ $X2=4.61 $Y2=2.005
r243 39 71 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=10.835 $Y=1.41
+ $X2=10.835 $Y2=1.245
r244 38 39 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.835
+ $Y=1.41 $X2=10.835 $Y2=1.41
r245 36 49 6.87075 $w=2.95e-07 $l=2.35654e-07 $layer=LI1_cond $X=10.07 $Y=1.407
+ $X2=9.897 $Y2=1.555
r246 36 38 29.8854 $w=2.93e-07 $l=7.65e-07 $layer=LI1_cond $X=10.07 $Y=1.407
+ $X2=10.835 $Y2=1.407
r247 33 41 3.37873 $w=1.7e-07 $l=1.8e-07 $layer=LI1_cond $X=4.79 $Y=1.635
+ $X2=4.61 $Y2=1.635
r248 33 76 40.123 $w=1.68e-07 $l=6.15e-07 $layer=LI1_cond $X=4.79 $Y=1.635
+ $X2=5.405 $Y2=1.635
r249 31 41 5.1848 $w=2.67e-07 $l=1.25499e-07 $layer=LI1_cond $X=4.7 $Y=1.55
+ $X2=4.61 $Y2=1.635
r250 30 31 23.4141 $w=1.78e-07 $l=3.8e-07 $layer=LI1_cond $X=4.7 $Y=1.17 $X2=4.7
+ $Y2=1.55
r251 26 43 2.41973 $w=4e-07 $l=4.7697e-08 $layer=LI1_cond $X=4.58 $Y=2.04
+ $X2=4.61 $Y2=2.005
r252 26 28 22.3286 $w=3.98e-07 $l=7.75e-07 $layer=LI1_cond $X=4.58 $Y=2.04
+ $X2=4.58 $Y2=2.815
r253 23 30 7.0541 $w=2.5e-07 $l=1.63936e-07 $layer=LI1_cond $X=4.61 $Y=1.045
+ $X2=4.7 $Y2=1.17
r254 23 25 2.928 $w=2.5e-07 $l=6e-08 $layer=LI1_cond $X=4.61 $Y=1.045 $X2=4.55
+ $Y2=1.045
r255 21 71 225.617 $w=1.5e-07 $l=4.4e-07 $layer=POLY_cond $X=10.745 $Y=0.805
+ $X2=10.745 $Y2=1.245
r256 16 68 55.8646 $w=2.93e-07 $l=3.05205e-07 $layer=POLY_cond $X=9.83 $Y=2.045
+ $X2=9.905 $Y2=1.775
r257 16 18 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=9.83 $Y=2.045
+ $X2=9.83 $Y2=2.54
r258 14 65 340.989 $w=1.5e-07 $l=6.65e-07 $layer=POLY_cond $X=6.47 $Y=0.805
+ $X2=6.47 $Y2=1.47
r259 9 11 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=5.72 $Y=2.41 $X2=5.72
+ $Y2=2.695
r260 8 9 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=5.72 $Y=2.32 $X2=5.72
+ $Y2=2.41
r261 7 63 15.0262 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=5.72 $Y=1.905
+ $X2=5.72 $Y2=1.74
r262 7 8 161.315 $w=1.8e-07 $l=4.15e-07 $layer=POLY_cond $X=5.72 $Y=1.905
+ $X2=5.72 $Y2=2.32
r263 2 43 400 $w=1.7e-07 $l=2.2798e-07 $layer=licon1_PDIFF $count=1 $X=4.395
+ $Y=1.84 $X2=4.545 $Y2=2.005
r264 2 28 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=4.395
+ $Y=1.84 $X2=4.545 $Y2=2.815
r265 1 25 182 $w=1.7e-07 $l=6.94226e-07 $layer=licon1_NDIFF $count=1 $X=4.335
+ $Y=0.41 $X2=4.55 $Y2=1.005
.ends

.subckt PM_SKY130_FD_SC_HS__SDFBBN_1%A_1159_497# 1 2 7 8 10 11 13 14 16 18 21 23
+ 25 26 30 31 32
c97 26 0 8.96875e-20 $X=6.42 $Y=1.215
c98 8 0 2.87426e-20 $X=7.25 $Y=1.33
r99 32 34 19.511 $w=2.72e-07 $l=4.35e-07 $layer=LI1_cond $X=6.03 $Y=2.055
+ $X2=6.03 $Y2=2.49
r100 30 31 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=7.085
+ $Y=1.42 $X2=7.085 $Y2=1.42
r101 28 30 19.2074 $w=3.28e-07 $l=5.5e-07 $layer=LI1_cond $X=7.085 $Y=1.97
+ $X2=7.085 $Y2=1.42
r102 27 30 4.1907 $w=3.28e-07 $l=1.2e-07 $layer=LI1_cond $X=7.085 $Y=1.3
+ $X2=7.085 $Y2=1.42
r103 25 27 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=6.92 $Y=1.215
+ $X2=7.085 $Y2=1.3
r104 25 26 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=6.92 $Y=1.215
+ $X2=6.42 $Y2=1.215
r105 24 32 3.48705 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.195 $Y=2.055
+ $X2=6.03 $Y2=2.055
r106 23 28 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=6.92 $Y=2.055
+ $X2=7.085 $Y2=1.97
r107 23 24 47.2995 $w=1.68e-07 $l=7.25e-07 $layer=LI1_cond $X=6.92 $Y=2.055
+ $X2=6.195 $Y2=2.055
r108 19 26 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=6.295 $Y=1.13
+ $X2=6.42 $Y2=1.215
r109 19 21 14.5208 $w=2.48e-07 $l=3.15e-07 $layer=LI1_cond $X=6.295 $Y=1.13
+ $X2=6.295 $Y2=0.815
r110 17 31 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=7.085 $Y=1.405
+ $X2=7.085 $Y2=1.42
r111 14 18 18.8402 $w=1.65e-07 $l=8.87412e-08 $layer=POLY_cond $X=7.61 $Y=1.255
+ $X2=7.58 $Y2=1.33
r112 14 16 123.713 $w=1.5e-07 $l=3.85e-07 $layer=POLY_cond $X=7.61 $Y=1.255
+ $X2=7.61 $Y2=0.87
r113 11 13 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=7.565 $Y=2.045
+ $X2=7.565 $Y2=2.54
r114 10 11 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=7.565 $Y=1.955
+ $X2=7.565 $Y2=2.045
r115 9 18 18.8402 $w=1.65e-07 $l=8.21584e-08 $layer=POLY_cond $X=7.565 $Y=1.405
+ $X2=7.58 $Y2=1.33
r116 9 10 213.79 $w=1.8e-07 $l=5.5e-07 $layer=POLY_cond $X=7.565 $Y=1.405
+ $X2=7.565 $Y2=1.955
r117 8 17 32.1775 $w=1.5e-07 $l=1.98997e-07 $layer=POLY_cond $X=7.25 $Y=1.33
+ $X2=7.085 $Y2=1.405
r118 7 18 6.66866 $w=1.5e-07 $l=1.05e-07 $layer=POLY_cond $X=7.475 $Y=1.33
+ $X2=7.58 $Y2=1.33
r119 7 8 115.372 $w=1.5e-07 $l=2.25e-07 $layer=POLY_cond $X=7.475 $Y=1.33
+ $X2=7.25 $Y2=1.33
r120 2 34 600 $w=1.7e-07 $l=2.37487e-07 $layer=licon1_PDIFF $count=1 $X=5.795
+ $Y=2.485 $X2=6.03 $Y2=2.49
r121 1 21 182 $w=1.7e-07 $l=2.81425e-07 $layer=licon1_NDIFF $count=1 $X=6.115
+ $Y=0.595 $X2=6.255 $Y2=0.815
.ends

.subckt PM_SKY130_FD_SC_HS__SDFBBN_1%A_1579_258# 1 2 8 9 11 14 16 18 19 20 21 23
+ 24 27 28 29 30 33 34 35 36 39 42 44 46 48 52 54 58 65
c202 58 0 9.562e-20 $X=12.365 $Y=1.215
c203 48 0 1.37535e-19 $X=8.265 $Y=1.375
c204 44 0 7.63376e-20 $X=13.78 $Y=1.915
c205 21 0 3.53982e-19 $X=12.47 $Y=1.885
c206 14 0 4.35224e-20 $X=8.14 $Y=0.87
c207 9 0 1.54972e-19 $X=7.985 $Y=2.045
c208 8 0 1.76028e-19 $X=7.985 $Y=1.955
r209 67 69 27.1035 $w=3.3e-07 $l=1.55e-07 $layer=POLY_cond $X=7.985 $Y=1.455
+ $X2=8.14 $Y2=1.455
r210 64 65 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=13.695 $Y=1.215
+ $X2=13.82 $Y2=1.215
r211 61 62 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=12.365
+ $Y=1.385 $X2=12.365 $Y2=1.385
r212 58 61 5.93683 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=12.365 $Y=1.215
+ $X2=12.365 $Y2=1.385
r213 54 56 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=10.835 $Y=0.45
+ $X2=10.835 $Y2=0.665
r214 52 69 21.8577 $w=3.3e-07 $l=1.25e-07 $layer=POLY_cond $X=8.265 $Y=1.455
+ $X2=8.14 $Y2=1.455
r215 51 52 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.265
+ $Y=1.455 $X2=8.265 $Y2=1.455
r216 48 51 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=8.265 $Y=1.375
+ $X2=8.265 $Y2=1.455
r217 44 46 4.14879 $w=2.48e-07 $l=9e-08 $layer=LI1_cond $X=13.78 $Y=1.915
+ $X2=13.87 $Y2=1.915
r218 40 65 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=13.82 $Y=1.13
+ $X2=13.82 $Y2=1.215
r219 40 42 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=13.82 $Y=1.13
+ $X2=13.82 $Y2=0.9
r220 39 44 7.14316 $w=2.5e-07 $l=1.62019e-07 $layer=LI1_cond $X=13.695 $Y=1.79
+ $X2=13.78 $Y2=1.915
r221 38 64 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=13.695 $Y=1.3
+ $X2=13.695 $Y2=1.215
r222 38 39 31.9679 $w=1.68e-07 $l=4.9e-07 $layer=LI1_cond $X=13.695 $Y=1.3
+ $X2=13.695 $Y2=1.79
r223 37 58 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12.53 $Y=1.215
+ $X2=12.365 $Y2=1.215
r224 36 64 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=13.61 $Y=1.215
+ $X2=13.695 $Y2=1.215
r225 36 37 70.4599 $w=1.68e-07 $l=1.08e-06 $layer=LI1_cond $X=13.61 $Y=1.215
+ $X2=12.53 $Y2=1.215
r226 34 58 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12.2 $Y=1.215
+ $X2=12.365 $Y2=1.215
r227 34 35 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=12.2 $Y=1.215
+ $X2=11.68 $Y2=1.215
r228 33 35 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=11.595 $Y=1.13
+ $X2=11.68 $Y2=1.215
r229 32 33 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=11.595 $Y=0.75
+ $X2=11.595 $Y2=1.13
r230 31 56 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.92 $Y=0.665
+ $X2=10.835 $Y2=0.665
r231 30 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=11.51 $Y=0.665
+ $X2=11.595 $Y2=0.75
r232 30 31 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=11.51 $Y=0.665
+ $X2=10.92 $Y2=0.665
r233 28 54 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.75 $Y=0.45
+ $X2=10.835 $Y2=0.45
r234 28 29 77.9626 $w=1.68e-07 $l=1.195e-06 $layer=LI1_cond $X=10.75 $Y=0.45
+ $X2=9.555 $Y2=0.45
r235 26 29 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.47 $Y=0.535
+ $X2=9.555 $Y2=0.45
r236 26 27 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=9.47 $Y=0.535
+ $X2=9.47 $Y2=1.29
r237 25 48 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.43 $Y=1.375
+ $X2=8.265 $Y2=1.375
r238 24 27 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.385 $Y=1.375
+ $X2=9.47 $Y2=1.29
r239 24 25 62.3048 $w=1.68e-07 $l=9.55e-07 $layer=LI1_cond $X=9.385 $Y=1.375
+ $X2=8.43 $Y2=1.375
r240 21 23 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=12.47 $Y=1.885
+ $X2=12.47 $Y2=2.46
r241 20 21 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=12.47 $Y=1.795
+ $X2=12.47 $Y2=1.885
r242 19 62 34.0194 $w=3.43e-07 $l=2.05122e-07 $layer=POLY_cond $X=12.47 $Y=1.55
+ $X2=12.38 $Y2=1.385
r243 19 20 95.2339 $w=1.8e-07 $l=2.45e-07 $layer=POLY_cond $X=12.47 $Y=1.55
+ $X2=12.47 $Y2=1.795
r244 16 62 38.7084 $w=3.43e-07 $l=1.94808e-07 $layer=POLY_cond $X=12.315 $Y=1.22
+ $X2=12.38 $Y2=1.385
r245 16 18 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=12.315 $Y=1.22
+ $X2=12.315 $Y2=0.74
r246 12 69 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.14 $Y=1.29
+ $X2=8.14 $Y2=1.455
r247 12 14 215.362 $w=1.5e-07 $l=4.2e-07 $layer=POLY_cond $X=8.14 $Y=1.29
+ $X2=8.14 $Y2=0.87
r248 9 11 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=7.985 $Y=2.045
+ $X2=7.985 $Y2=2.54
r249 8 9 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=7.985 $Y=1.955
+ $X2=7.985 $Y2=2.045
r250 7 67 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=7.985 $Y=1.62
+ $X2=7.985 $Y2=1.455
r251 7 8 130.218 $w=1.8e-07 $l=3.35e-07 $layer=POLY_cond $X=7.985 $Y=1.62
+ $X2=7.985 $Y2=1.955
r252 2 46 600 $w=1.7e-07 $l=3.34739e-07 $layer=licon1_PDIFF $count=1 $X=13.6
+ $Y=1.73 $X2=13.87 $Y2=1.875
r253 1 42 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=13.675
+ $Y=0.69 $X2=13.82 $Y2=0.9
.ends

.subckt PM_SKY130_FD_SC_HS__SDFBBN_1%SET_B 1 3 6 8 10 13 15 16 19 21 24 30
c135 24 0 3.15057e-19 $X=8.745 $Y=1.837
c136 21 0 1.48476e-19 $X=11.76 $Y=2.035
c137 6 0 1.76028e-19 $X=8.745 $Y=0.87
r138 30 34 13.969 $w=3.28e-07 $l=4e-07 $layer=LI1_cond $X=11.795 $Y=1.635
+ $X2=11.795 $Y2=2.035
r139 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=11.795
+ $Y=1.635 $X2=11.795 $Y2=1.635
r140 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.825
+ $Y=1.795 $X2=8.825 $Y2=1.795
r141 24 26 13.9206 $w=2.77e-07 $l=8e-08 $layer=POLY_cond $X=8.745 $Y=1.837
+ $X2=8.825 $Y2=1.837
r142 21 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.76 $Y=2.035
+ $X2=11.76 $Y2=2.035
r143 19 27 17.4579 $w=2.97e-07 $l=4.25e-07 $layer=LI1_cond $X=8.4 $Y=1.885
+ $X2=8.825 $Y2=1.885
r144 18 19 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=2.035
+ $X2=8.4 $Y2=2.035
r145 16 18 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=8.545 $Y=2.035
+ $X2=8.4 $Y2=2.035
r146 15 21 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=11.615 $Y=2.035
+ $X2=11.76 $Y2=2.035
r147 15 16 3.7995 $w=1.4e-07 $l=3.07e-06 $layer=MET1_cond $X=11.615 $Y=2.035
+ $X2=8.545 $Y2=2.035
r148 11 29 38.5562 $w=2.99e-07 $l=2.05122e-07 $layer=POLY_cond $X=11.885 $Y=1.47
+ $X2=11.795 $Y2=1.635
r149 11 13 374.319 $w=1.5e-07 $l=7.3e-07 $layer=POLY_cond $X=11.885 $Y=1.47
+ $X2=11.885 $Y2=0.74
r150 8 29 52.2586 $w=2.99e-07 $l=2.76134e-07 $layer=POLY_cond $X=11.85 $Y=1.885
+ $X2=11.795 $Y2=1.635
r151 8 10 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=11.85 $Y=1.885
+ $X2=11.85 $Y2=2.46
r152 4 24 17.1008 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=8.745 $Y=1.63
+ $X2=8.745 $Y2=1.837
r153 4 6 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=8.745 $Y=1.63
+ $X2=8.745 $Y2=0.87
r154 1 24 53.9422 $w=2.77e-07 $l=4.00724e-07 $layer=POLY_cond $X=8.435 $Y=2.045
+ $X2=8.745 $Y2=1.837
r155 1 3 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=8.435 $Y=2.045
+ $X2=8.435 $Y2=2.54
.ends

.subckt PM_SKY130_FD_SC_HS__SDFBBN_1%A_662_82# 1 2 10 11 13 14 15 19 21 22 24 26
+ 30 31 32 35 37 38 40 43 45 46 50 52 54 57 59 65
c184 65 0 1.49471e-19 $X=4.335 $Y=1.505
c185 38 0 4.28297e-20 $X=6.04 $Y=0.18
c186 35 0 3.95129e-20 $X=10.365 $Y=2.465
c187 31 0 1.94296e-19 $X=10.28 $Y=1.295
c188 11 0 7.19434e-20 $X=4.32 $Y=1.765
r189 65 66 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.335
+ $Y=1.505 $X2=4.335 $Y2=1.505
r190 62 65 9.7783 $w=3.28e-07 $l=2.8e-07 $layer=LI1_cond $X=4.055 $Y=1.505
+ $X2=4.335 $Y2=1.505
r191 58 62 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.055 $Y=1.67
+ $X2=4.055 $Y2=1.505
r192 58 59 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=4.055 $Y=1.67
+ $X2=4.055 $Y2=1.95
r193 57 62 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.055 $Y=1.34
+ $X2=4.055 $Y2=1.505
r194 56 57 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=4.055 $Y=1.17
+ $X2=4.055 $Y2=1.34
r195 55 61 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.73 $Y=2.035
+ $X2=3.605 $Y2=2.035
r196 54 59 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.97 $Y=2.035
+ $X2=4.055 $Y2=1.95
r197 54 55 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=3.97 $Y=2.035
+ $X2=3.73 $Y2=2.035
r198 50 61 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.605 $Y=2.12
+ $X2=3.605 $Y2=2.035
r199 50 52 32.0379 $w=2.48e-07 $l=6.95e-07 $layer=LI1_cond $X=3.605 $Y=2.12
+ $X2=3.605 $Y2=2.815
r200 46 56 7.14316 $w=2.5e-07 $l=1.62019e-07 $layer=LI1_cond $X=3.97 $Y=1.045
+ $X2=4.055 $Y2=1.17
r201 46 48 23.7403 $w=2.48e-07 $l=5.15e-07 $layer=LI1_cond $X=3.97 $Y=1.045
+ $X2=3.455 $Y2=1.045
r202 41 43 82.0426 $w=1.5e-07 $l=1.6e-07 $layer=POLY_cond $X=6.095 $Y=2.115
+ $X2=6.255 $Y2=2.115
r203 39 40 48.5235 $w=2.05e-07 $l=1.5e-07 $layer=POLY_cond $X=6.067 $Y=1.09
+ $X2=6.067 $Y2=1.24
r204 35 45 110.782 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=10.365 $Y=2.465
+ $X2=10.365 $Y2=2.18
r205 35 37 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=10.365 $Y=2.465
+ $X2=10.365 $Y2=2.75
r206 33 45 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=10.355 $Y=1.37
+ $X2=10.355 $Y2=2.18
r207 31 33 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=10.28 $Y=1.295
+ $X2=10.355 $Y2=1.37
r208 31 32 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=10.28 $Y=1.295
+ $X2=9.77 $Y2=1.295
r209 28 32 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=9.695 $Y=1.22
+ $X2=9.77 $Y2=1.295
r210 28 30 179.468 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=9.695 $Y=1.22
+ $X2=9.695 $Y2=0.87
r211 27 30 315.351 $w=1.5e-07 $l=6.15e-07 $layer=POLY_cond $X=9.695 $Y=0.255
+ $X2=9.695 $Y2=0.87
r212 24 43 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.255 $Y=2.19
+ $X2=6.255 $Y2=2.115
r213 24 26 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=6.255 $Y=2.19
+ $X2=6.255 $Y2=2.585
r214 23 38 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.115 $Y=0.18
+ $X2=6.04 $Y2=0.18
r215 22 27 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=9.62 $Y=0.18
+ $X2=9.695 $Y2=0.255
r216 22 23 1797.24 $w=1.5e-07 $l=3.505e-06 $layer=POLY_cond $X=9.62 $Y=0.18
+ $X2=6.115 $Y2=0.18
r217 21 41 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.095 $Y=2.04
+ $X2=6.095 $Y2=2.115
r218 21 40 410.213 $w=1.5e-07 $l=8e-07 $layer=POLY_cond $X=6.095 $Y=2.04
+ $X2=6.095 $Y2=1.24
r219 19 39 146.138 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=6.04 $Y=0.805
+ $X2=6.04 $Y2=1.09
r220 16 38 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.04 $Y=0.255
+ $X2=6.04 $Y2=0.18
r221 16 19 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=6.04 $Y=0.255
+ $X2=6.04 $Y2=0.805
r222 14 38 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.965 $Y=0.18
+ $X2=6.04 $Y2=0.18
r223 14 15 835.809 $w=1.5e-07 $l=1.63e-06 $layer=POLY_cond $X=5.965 $Y=0.18
+ $X2=4.335 $Y2=0.18
r224 11 66 54.0414 $w=2.96e-07 $l=2.67395e-07 $layer=POLY_cond $X=4.32 $Y=1.765
+ $X2=4.335 $Y2=1.505
r225 11 13 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=4.32 $Y=1.765
+ $X2=4.32 $Y2=2.4
r226 8 66 38.5718 $w=2.96e-07 $l=1.98997e-07 $layer=POLY_cond $X=4.26 $Y=1.34
+ $X2=4.335 $Y2=1.505
r227 8 10 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=4.26 $Y=1.34
+ $X2=4.26 $Y2=0.78
r228 7 15 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.26 $Y=0.255
+ $X2=4.335 $Y2=0.18
r229 7 10 269.202 $w=1.5e-07 $l=5.25e-07 $layer=POLY_cond $X=4.26 $Y=0.255
+ $X2=4.26 $Y2=0.78
r230 2 61 400 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_PDIFF $count=1 $X=3.5
+ $Y=1.84 $X2=3.645 $Y2=2.115
r231 2 52 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=3.5
+ $Y=1.84 $X2=3.645 $Y2=2.815
r232 1 48 182 $w=1.7e-07 $l=6.63551e-07 $layer=licon1_NDIFF $count=1 $X=3.31
+ $Y=0.41 $X2=3.455 $Y2=1.005
.ends

.subckt PM_SKY130_FD_SC_HS__SDFBBN_1%A_2133_410# 1 2 3 10 12 13 17 19 21 24 26
+ 29 30 32 35 37 40 44 45 47 49 50 51 54 55 56 58 59 60 64 67 68 70 77 79
c234 49 0 1.30488e-19 $X=13.115 $Y=2.38
c235 24 0 1.65234e-19 $X=14.785 $Y=0.74
r236 78 83 5.05594 $w=2.86e-07 $l=3e-08 $layer=POLY_cond $X=14.77 $Y=1.465
+ $X2=14.77 $Y2=1.435
r237 77 80 8.58894 $w=3.83e-07 $l=1.65e-07 $layer=LI1_cond $X=14.742 $Y=1.465
+ $X2=14.742 $Y2=1.63
r238 77 79 8.58894 $w=3.83e-07 $l=1.65e-07 $layer=LI1_cond $X=14.742 $Y=1.465
+ $X2=14.742 $Y2=1.3
r239 77 78 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=14.77
+ $Y=1.465 $X2=14.77 $Y2=1.465
r240 70 72 3.49225 $w=3.28e-07 $l=1e-07 $layer=LI1_cond $X=12.63 $Y=0.775
+ $X2=12.63 $Y2=0.875
r241 66 68 8.48848 $w=3.48e-07 $l=1.65e-07 $layer=LI1_cond $X=11.625 $Y=2.805
+ $X2=11.79 $Y2=2.805
r242 66 67 8.48848 $w=3.48e-07 $l=1.65e-07 $layer=LI1_cond $X=11.625 $Y=2.805
+ $X2=11.46 $Y2=2.805
r243 64 80 37.8396 $w=1.68e-07 $l=5.8e-07 $layer=LI1_cond $X=14.635 $Y=2.21
+ $X2=14.635 $Y2=1.63
r244 61 79 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=14.635 $Y=1.02
+ $X2=14.635 $Y2=1.3
r245 59 61 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=14.55 $Y=0.935
+ $X2=14.635 $Y2=1.02
r246 59 60 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=14.55 $Y=0.935
+ $X2=14.245 $Y2=0.935
r247 58 60 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=14.16 $Y=0.85
+ $X2=14.245 $Y2=0.935
r248 57 58 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=14.16 $Y=0.5
+ $X2=14.16 $Y2=0.85
r249 55 57 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=14.075 $Y=0.415
+ $X2=14.16 $Y2=0.5
r250 55 56 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=14.075 $Y=0.415
+ $X2=13.565 $Y2=0.415
r251 53 56 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=13.48 $Y=0.5
+ $X2=13.565 $Y2=0.415
r252 53 54 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=13.48 $Y=0.5
+ $X2=13.48 $Y2=0.79
r253 52 75 4.65971 $w=1.7e-07 $l=1.98997e-07 $layer=LI1_cond $X=13.28 $Y=2.295
+ $X2=13.115 $Y2=2.22
r254 51 64 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=14.55 $Y=2.295
+ $X2=14.635 $Y2=2.21
r255 51 52 82.8556 $w=1.68e-07 $l=1.27e-06 $layer=LI1_cond $X=14.55 $Y=2.295
+ $X2=13.28 $Y2=2.295
r256 49 75 3.10647 $w=3.3e-07 $l=1.6e-07 $layer=LI1_cond $X=13.115 $Y=2.38
+ $X2=13.115 $Y2=2.22
r257 49 50 8.73063 $w=3.28e-07 $l=2.5e-07 $layer=LI1_cond $X=13.115 $Y=2.38
+ $X2=13.115 $Y2=2.63
r258 48 72 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12.795 $Y=0.875
+ $X2=12.63 $Y2=0.875
r259 47 54 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=13.395 $Y=0.875
+ $X2=13.48 $Y2=0.79
r260 47 48 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=13.395 $Y=0.875
+ $X2=12.795 $Y2=0.875
r261 45 50 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=12.95 $Y=2.715
+ $X2=13.115 $Y2=2.63
r262 45 68 75.6791 $w=1.68e-07 $l=1.16e-06 $layer=LI1_cond $X=12.95 $Y=2.715
+ $X2=11.79 $Y2=2.715
r263 44 67 30.3369 $w=1.68e-07 $l=4.65e-07 $layer=LI1_cond $X=10.995 $Y=2.715
+ $X2=11.46 $Y2=2.715
r264 41 81 14.5084 $w=2.99e-07 $l=9e-08 $layer=POLY_cond $X=10.83 $Y=2.215
+ $X2=10.83 $Y2=2.125
r265 40 41 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.83
+ $Y=2.215 $X2=10.83 $Y2=2.215
r266 38 44 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=10.83 $Y=2.63
+ $X2=10.995 $Y2=2.715
r267 38 40 14.4928 $w=3.28e-07 $l=4.15e-07 $layer=LI1_cond $X=10.83 $Y=2.63
+ $X2=10.83 $Y2=2.215
r268 33 37 30.0832 $w=1.65e-07 $l=1.42302e-07 $layer=POLY_cond $X=15.775 $Y=1.3
+ $X2=15.76 $Y2=1.435
r269 33 35 335.862 $w=1.5e-07 $l=6.55e-07 $layer=POLY_cond $X=15.775 $Y=1.3
+ $X2=15.775 $Y2=0.645
r270 30 32 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=15.76 $Y=1.845
+ $X2=15.76 $Y2=2.34
r271 29 30 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=15.76 $Y=1.755
+ $X2=15.76 $Y2=1.845
r272 28 37 30.0832 $w=1.65e-07 $l=1.35e-07 $layer=POLY_cond $X=15.76 $Y=1.57
+ $X2=15.76 $Y2=1.435
r273 28 29 71.9113 $w=1.8e-07 $l=1.85e-07 $layer=POLY_cond $X=15.76 $Y=1.57
+ $X2=15.76 $Y2=1.755
r274 27 83 4.208 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=14.935 $Y=1.435
+ $X2=14.77 $Y2=1.435
r275 26 37 1.40033 $w=2.7e-07 $l=9e-08 $layer=POLY_cond $X=15.67 $Y=1.435
+ $X2=15.76 $Y2=1.435
r276 26 27 163.298 $w=2.7e-07 $l=7.35e-07 $layer=POLY_cond $X=15.67 $Y=1.435
+ $X2=14.935 $Y2=1.435
r277 22 83 33.5989 $w=2.86e-07 $l=1.42302e-07 $layer=POLY_cond $X=14.785 $Y=1.3
+ $X2=14.77 $Y2=1.435
r278 22 24 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=14.785 $Y=1.3
+ $X2=14.785 $Y2=0.74
r279 19 78 61.4066 $w=2.86e-07 $l=3.09839e-07 $layer=POLY_cond $X=14.75 $Y=1.765
+ $X2=14.77 $Y2=1.465
r280 19 21 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=14.75 $Y=1.765
+ $X2=14.75 $Y2=2.4
r281 15 17 638.394 $w=1.5e-07 $l=1.245e-06 $layer=POLY_cond $X=11.285 $Y=2.05
+ $X2=11.285 $Y2=0.805
r282 14 81 18.89 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=10.995 $Y=2.125
+ $X2=10.83 $Y2=2.125
r283 13 15 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=11.21 $Y=2.125
+ $X2=11.285 $Y2=2.05
r284 13 14 110.245 $w=1.5e-07 $l=2.15e-07 $layer=POLY_cond $X=11.21 $Y=2.125
+ $X2=10.995 $Y2=2.125
r285 10 41 52.2586 $w=2.99e-07 $l=2.85044e-07 $layer=POLY_cond $X=10.755
+ $Y=2.465 $X2=10.83 $Y2=2.215
r286 10 12 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=10.755 $Y=2.465
+ $X2=10.755 $Y2=2.75
r287 3 75 300 $w=1.7e-07 $l=3.31625e-07 $layer=licon1_PDIFF $count=2 $X=12.965
+ $Y=1.96 $X2=13.115 $Y2=2.225
r288 2 66 600 $w=1.7e-07 $l=9.14631e-07 $layer=licon1_PDIFF $count=1 $X=11.48
+ $Y=1.96 $X2=11.625 $Y2=2.805
r289 1 70 182 $w=1.7e-07 $l=5.11102e-07 $layer=licon1_NDIFF $count=1 $X=12.39
+ $Y=0.37 $X2=12.63 $Y2=0.775
.ends

.subckt PM_SKY130_FD_SC_HS__SDFBBN_1%A_1954_119# 1 2 9 11 13 20 23 24 25 26 29
+ 31 32 33 35 36 38 39 44 47 48 49
c145 48 0 1.86341e-19 $X=10.58 $Y=0.897
c146 47 0 1.23448e-20 $X=10.415 $Y=0.87
c147 44 0 1.74547e-19 $X=10.325 $Y=2.195
c148 39 0 7.63376e-20 $X=13.275 $Y=1.635
c149 36 0 7.50187e-20 $X=12.78 $Y=1.68
c150 25 0 1.94296e-19 $X=10.41 $Y=1.81
c151 23 0 3.95129e-20 $X=10.325 $Y=2.11
c152 11 0 9.562e-20 $X=12.89 $Y=1.885
r153 47 48 8.58894 $w=3.83e-07 $l=1.65e-07 $layer=LI1_cond $X=10.415 $Y=0.897
+ $X2=10.58 $Y2=0.897
r154 42 44 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=10.055 $Y=2.195
+ $X2=10.325 $Y2=2.195
r155 38 39 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=13.275
+ $Y=1.635 $X2=13.275 $Y2=1.635
r156 36 38 13.5824 $w=4.18e-07 $l=4.95e-07 $layer=LI1_cond $X=12.78 $Y=1.68
+ $X2=13.275 $Y2=1.68
r157 34 36 7.86469 $w=3.2e-07 $l=2.48898e-07 $layer=LI1_cond $X=12.695 $Y=1.89
+ $X2=12.78 $Y2=1.68
r158 34 35 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=12.695 $Y=1.89
+ $X2=12.695 $Y2=2.29
r159 32 35 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=12.61 $Y=2.375
+ $X2=12.695 $Y2=2.29
r160 32 33 82.8556 $w=1.68e-07 $l=1.27e-06 $layer=LI1_cond $X=12.61 $Y=2.375
+ $X2=11.34 $Y2=2.375
r161 31 33 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=11.255 $Y=2.29
+ $X2=11.34 $Y2=2.375
r162 30 49 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=11.255 $Y=1.895
+ $X2=11.255 $Y2=1.81
r163 30 31 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=11.255 $Y=1.895
+ $X2=11.255 $Y2=2.29
r164 29 49 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=11.255 $Y=1.725
+ $X2=11.255 $Y2=1.81
r165 28 29 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=11.255 $Y=1.09
+ $X2=11.255 $Y2=1.725
r166 26 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=11.17 $Y=1.005
+ $X2=11.255 $Y2=1.09
r167 26 48 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=11.17 $Y=1.005
+ $X2=10.58 $Y2=1.005
r168 24 49 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=11.17 $Y=1.81
+ $X2=11.255 $Y2=1.81
r169 24 25 49.5829 $w=1.68e-07 $l=7.6e-07 $layer=LI1_cond $X=11.17 $Y=1.81
+ $X2=10.41 $Y2=1.81
r170 23 44 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.325 $Y=2.11
+ $X2=10.325 $Y2=2.195
r171 22 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=10.325 $Y=1.895
+ $X2=10.41 $Y2=1.81
r172 22 23 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=10.325 $Y=1.895
+ $X2=10.325 $Y2=2.11
r173 20 42 18.6835 $w=3.28e-07 $l=5.35e-07 $layer=LI1_cond $X=10.055 $Y=2.815
+ $X2=10.055 $Y2=2.28
r174 15 39 51.5841 $w=3.3e-07 $l=2.95e-07 $layer=POLY_cond $X=12.98 $Y=1.635
+ $X2=13.275 $Y2=1.635
r175 11 15 62.743 $w=2.03e-07 $l=2.57391e-07 $layer=POLY_cond $X=12.89 $Y=1.885
+ $X2=12.875 $Y2=1.635
r176 11 13 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=12.89 $Y=1.885
+ $X2=12.89 $Y2=2.46
r177 7 15 42.5607 $w=2.03e-07 $l=1.79374e-07 $layer=POLY_cond $X=12.845 $Y=1.47
+ $X2=12.875 $Y2=1.635
r178 7 9 374.319 $w=1.5e-07 $l=7.3e-07 $layer=POLY_cond $X=12.845 $Y=1.47
+ $X2=12.845 $Y2=0.74
r179 2 42 600 $w=1.7e-07 $l=2.17428e-07 $layer=licon1_PDIFF $count=1 $X=9.905
+ $Y=2.12 $X2=10.055 $Y2=2.275
r180 2 20 600 $w=1.7e-07 $l=7.66339e-07 $layer=licon1_PDIFF $count=1 $X=9.905
+ $Y=2.12 $X2=10.055 $Y2=2.815
r181 1 47 91 $w=1.7e-07 $l=7.70325e-07 $layer=licon1_NDIFF $count=2 $X=9.77
+ $Y=0.595 $X2=10.415 $Y2=0.87
.ends

.subckt PM_SKY130_FD_SC_HS__SDFBBN_1%RESET_B 1 3 4 6 7 8 10 11 18
c53 11 0 1.65234e-19 $X=14.16 $Y=1.295
r54 16 18 5.24584 $w=3.3e-07 $l=3e-08 $layer=POLY_cond $X=14.23 $Y=1.385
+ $X2=14.26 $Y2=1.385
r55 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=14.23
+ $Y=1.385 $X2=14.23 $Y2=1.385
r56 13 16 34.0979 $w=3.3e-07 $l=1.95e-07 $layer=POLY_cond $X=14.035 $Y=1.385
+ $X2=14.23 $Y2=1.385
r57 11 17 3.40065 $w=3.03e-07 $l=9e-08 $layer=LI1_cond $X=14.227 $Y=1.295
+ $X2=14.227 $Y2=1.385
r58 9 18 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=14.26 $Y=1.55
+ $X2=14.26 $Y2=1.385
r59 9 10 279.457 $w=1.5e-07 $l=5.45e-07 $layer=POLY_cond $X=14.26 $Y=1.55
+ $X2=14.26 $Y2=2.095
r60 7 10 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=14.185 $Y=2.17
+ $X2=14.26 $Y2=2.095
r61 7 8 87.1702 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=14.185 $Y=2.17
+ $X2=14.015 $Y2=2.17
r62 4 13 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=14.035 $Y=1.22
+ $X2=14.035 $Y2=1.385
r63 4 6 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=14.035 $Y=1.22
+ $X2=14.035 $Y2=0.9
r64 1 8 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=13.94 $Y=2.245
+ $X2=14.015 $Y2=2.17
r65 1 3 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=13.94 $Y=2.245
+ $X2=13.94 $Y2=2.64
.ends

.subckt PM_SKY130_FD_SC_HS__SDFBBN_1%A_3078_384# 1 2 7 9 10 12 15 19 23 26
r52 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=16.225
+ $Y=1.385 $X2=16.225 $Y2=1.385
r53 21 26 0.533013 $w=3.3e-07 $l=1.38e-07 $layer=LI1_cond $X=15.725 $Y=1.385
+ $X2=15.587 $Y2=1.385
r54 21 23 17.4613 $w=3.28e-07 $l=5e-07 $layer=LI1_cond $X=15.725 $Y=1.385
+ $X2=16.225 $Y2=1.385
r55 17 26 6.22203 $w=2.62e-07 $l=1.70895e-07 $layer=LI1_cond $X=15.575 $Y=1.55
+ $X2=15.587 $Y2=1.385
r56 17 19 23.7403 $w=2.48e-07 $l=5.15e-07 $layer=LI1_cond $X=15.575 $Y=1.55
+ $X2=15.575 $Y2=2.065
r57 13 26 6.22203 $w=2.62e-07 $l=1.65e-07 $layer=LI1_cond $X=15.587 $Y=1.22
+ $X2=15.587 $Y2=1.385
r58 13 15 24.0965 $w=2.73e-07 $l=5.75e-07 $layer=LI1_cond $X=15.587 $Y=1.22
+ $X2=15.587 $Y2=0.645
r59 10 24 77.2841 $w=2.7e-07 $l=4.13521e-07 $layer=POLY_cond $X=16.295 $Y=1.765
+ $X2=16.225 $Y2=1.385
r60 10 12 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=16.295 $Y=1.765
+ $X2=16.295 $Y2=2.4
r61 7 24 38.9026 $w=2.7e-07 $l=1.92678e-07 $layer=POLY_cond $X=16.285 $Y=1.22
+ $X2=16.225 $Y2=1.385
r62 7 9 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=16.285 $Y=1.22
+ $X2=16.285 $Y2=0.74
r63 2 19 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=15.39
+ $Y=1.92 $X2=15.535 $Y2=2.065
r64 1 15 182 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_NDIFF $count=1 $X=15.415
+ $Y=0.37 $X2=15.56 $Y2=0.645
.ends

.subckt PM_SKY130_FD_SC_HS__SDFBBN_1%A_27_464# 1 2 9 11 12 14 15 16 19
c50 16 0 1.00461e-19 $X=1.235 $Y=2.99
c51 14 0 8.80698e-20 $X=1.15 $Y=2.905
r52 17 19 15.3659 $w=3.28e-07 $l=4.4e-07 $layer=LI1_cond $X=2.08 $Y=2.905
+ $X2=2.08 $Y2=2.465
r53 15 17 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.915 $Y=2.99
+ $X2=2.08 $Y2=2.905
r54 15 16 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.915 $Y=2.99
+ $X2=1.235 $Y2=2.99
r55 14 16 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.15 $Y=2.905
+ $X2=1.235 $Y2=2.99
r56 13 14 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.15 $Y=2.215
+ $X2=1.15 $Y2=2.905
r57 11 13 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.065 $Y=2.13
+ $X2=1.15 $Y2=2.215
r58 11 12 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.065 $Y=2.13
+ $X2=0.395 $Y2=2.13
r59 7 12 7.36005 $w=1.7e-07 $l=1.77482e-07 $layer=LI1_cond $X=0.255 $Y=2.215
+ $X2=0.395 $Y2=2.13
r60 7 9 10.2897 $w=2.78e-07 $l=2.5e-07 $layer=LI1_cond $X=0.255 $Y=2.215
+ $X2=0.255 $Y2=2.465
r61 2 19 300 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=2 $X=1.93
+ $Y=2.32 $X2=2.08 $Y2=2.465
r62 1 9 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=2.32 $X2=0.28 $Y2=2.465
.ends

.subckt PM_SKY130_FD_SC_HS__SDFBBN_1%VPWR 1 2 3 4 5 6 7 8 9 10 33 37 41 43 47 51
+ 55 59 63 68 69 71 74 78 79 80 82 87 95 107 115 119 132 133 136 139 142 145 148
+ 151 158
c188 6 0 1.7536e-19 $X=9.07 $Y=2.12
r189 159 161 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=14.64 $Y=3.33
+ $X2=14.16 $Y2=3.33
r190 158 161 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=14.16 $Y=3.33
+ $X2=14.16 $Y2=3.33
r191 158 159 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=14.64 $Y=3.33
+ $X2=14.64 $Y2=3.33
r192 154 155 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.24 $Y=3.33
+ $X2=12.24 $Y2=3.33
r193 151 154 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=12.16 $Y=3.055
+ $X2=12.16 $Y2=3.33
r194 148 149 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.36 $Y=3.33
+ $X2=9.36 $Y2=3.33
r195 145 146 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r196 143 146 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=5.04 $Y2=3.33
r197 142 143 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r198 139 140 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r199 136 137 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r200 132 133 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=16.56 $Y=3.33
+ $X2=16.56 $Y2=3.33
r201 130 133 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=15.6 $Y=3.33
+ $X2=16.56 $Y2=3.33
r202 130 159 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=15.6 $Y=3.33
+ $X2=14.64 $Y2=3.33
r203 129 130 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=15.6 $Y=3.33
+ $X2=15.6 $Y2=3.33
r204 127 158 13.5574 $w=1.7e-07 $l=3.45e-07 $layer=LI1_cond $X=14.69 $Y=3.33
+ $X2=14.345 $Y2=3.33
r205 127 129 59.369 $w=1.68e-07 $l=9.1e-07 $layer=LI1_cond $X=14.69 $Y=3.33
+ $X2=15.6 $Y2=3.33
r206 126 161 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=13.68 $Y=3.33
+ $X2=14.16 $Y2=3.33
r207 125 126 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=13.68 $Y=3.33
+ $X2=13.68 $Y2=3.33
r208 123 126 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=12.72 $Y=3.33
+ $X2=13.68 $Y2=3.33
r209 123 155 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.72 $Y=3.33
+ $X2=12.24 $Y2=3.33
r210 122 125 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=12.72 $Y=3.33
+ $X2=13.68 $Y2=3.33
r211 122 123 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=12.72 $Y=3.33
+ $X2=12.72 $Y2=3.33
r212 120 154 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12.325 $Y=3.33
+ $X2=12.16 $Y2=3.33
r213 120 122 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=12.325 $Y=3.33
+ $X2=12.72 $Y2=3.33
r214 119 158 13.5574 $w=1.7e-07 $l=3.45e-07 $layer=LI1_cond $X=14 $Y=3.33
+ $X2=14.345 $Y2=3.33
r215 119 125 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=14 $Y=3.33
+ $X2=13.68 $Y2=3.33
r216 118 155 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.76 $Y=3.33
+ $X2=12.24 $Y2=3.33
r217 117 118 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=11.76 $Y=3.33
+ $X2=11.76 $Y2=3.33
r218 115 154 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.995 $Y=3.33
+ $X2=12.16 $Y2=3.33
r219 115 117 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=11.995 $Y=3.33
+ $X2=11.76 $Y2=3.33
r220 114 118 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=10.8 $Y=3.33
+ $X2=11.76 $Y2=3.33
r221 114 149 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=10.8 $Y=3.33
+ $X2=9.36 $Y2=3.33
r222 113 114 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.8 $Y=3.33
+ $X2=10.8 $Y2=3.33
r223 111 148 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.38 $Y=3.33
+ $X2=9.215 $Y2=3.33
r224 111 113 92.6417 $w=1.68e-07 $l=1.42e-06 $layer=LI1_cond $X=9.38 $Y=3.33
+ $X2=10.8 $Y2=3.33
r225 110 149 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=3.33
+ $X2=9.36 $Y2=3.33
r226 109 110 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r227 107 148 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.05 $Y=3.33
+ $X2=9.215 $Y2=3.33
r228 107 109 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=9.05 $Y=3.33
+ $X2=8.88 $Y2=3.33
r229 105 106 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r230 103 106 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=7.92 $Y2=3.33
r231 103 146 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=5.04 $Y2=3.33
r232 102 105 156.578 $w=1.68e-07 $l=2.4e-06 $layer=LI1_cond $X=5.52 $Y=3.33
+ $X2=7.92 $Y2=3.33
r233 102 103 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r234 100 145 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.27 $Y=3.33
+ $X2=5.145 $Y2=3.33
r235 100 102 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=5.27 $Y=3.33
+ $X2=5.52 $Y2=3.33
r236 99 143 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.08 $Y2=3.33
r237 99 140 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=2.64 $Y2=3.33
r238 98 99 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r239 96 139 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.72 $Y=3.33
+ $X2=2.595 $Y2=3.33
r240 96 98 57.4118 $w=1.68e-07 $l=8.8e-07 $layer=LI1_cond $X=2.72 $Y=3.33
+ $X2=3.6 $Y2=3.33
r241 95 142 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.93 $Y=3.33
+ $X2=4.055 $Y2=3.33
r242 95 98 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=3.93 $Y=3.33
+ $X2=3.6 $Y2=3.33
r243 94 140 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r244 93 94 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r245 91 94 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.16 $Y2=3.33
r246 91 137 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r247 90 93 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.2 $Y=3.33 $X2=2.16
+ $Y2=3.33
r248 90 91 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r249 88 136 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.895 $Y=3.33
+ $X2=0.73 $Y2=3.33
r250 88 90 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.895 $Y=3.33
+ $X2=1.2 $Y2=3.33
r251 87 139 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.47 $Y=3.33
+ $X2=2.595 $Y2=3.33
r252 87 93 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=2.47 $Y=3.33
+ $X2=2.16 $Y2=3.33
r253 85 137 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r254 84 85 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r255 82 136 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.565 $Y=3.33
+ $X2=0.73 $Y2=3.33
r256 82 84 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.565 $Y=3.33
+ $X2=0.24 $Y2=3.33
r257 80 110 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=3.33
+ $X2=8.88 $Y2=3.33
r258 80 106 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=3.33
+ $X2=7.92 $Y2=3.33
r259 78 129 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=15.905 $Y=3.33
+ $X2=15.6 $Y2=3.33
r260 78 79 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=15.905 $Y=3.33
+ $X2=16.03 $Y2=3.33
r261 77 132 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=16.155 $Y=3.33
+ $X2=16.56 $Y2=3.33
r262 77 79 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=16.155 $Y=3.33
+ $X2=16.03 $Y2=3.33
r263 75 117 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=11.23 $Y=3.33
+ $X2=11.76 $Y2=3.33
r264 74 113 6.52406 $w=1.68e-07 $l=1e-07 $layer=LI1_cond $X=10.9 $Y=3.33
+ $X2=10.8 $Y2=3.33
r265 73 75 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.065 $Y=3.33
+ $X2=11.23 $Y2=3.33
r266 73 74 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.065 $Y=3.33
+ $X2=10.9 $Y2=3.33
r267 71 73 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=11.065 $Y=3.055
+ $X2=11.065 $Y2=3.33
r268 68 105 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=8.125 $Y=3.33
+ $X2=7.92 $Y2=3.33
r269 68 69 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.125 $Y=3.33
+ $X2=8.21 $Y2=3.33
r270 67 109 38.1658 $w=1.68e-07 $l=5.85e-07 $layer=LI1_cond $X=8.295 $Y=3.33
+ $X2=8.88 $Y2=3.33
r271 67 69 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.295 $Y=3.33
+ $X2=8.21 $Y2=3.33
r272 63 66 34.5733 $w=2.48e-07 $l=7.5e-07 $layer=LI1_cond $X=16.03 $Y=2.065
+ $X2=16.03 $Y2=2.815
r273 61 79 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=16.03 $Y=3.245
+ $X2=16.03 $Y2=3.33
r274 61 66 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=16.03 $Y=3.245
+ $X2=16.03 $Y2=2.815
r275 57 158 2.83173 $w=6.9e-07 $l=8.5e-08 $layer=LI1_cond $X=14.345 $Y=3.245
+ $X2=14.345 $Y2=3.33
r276 57 59 9.7073 $w=6.88e-07 $l=5.6e-07 $layer=LI1_cond $X=14.345 $Y=3.245
+ $X2=14.345 $Y2=2.685
r277 53 148 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.215 $Y=3.245
+ $X2=9.215 $Y2=3.33
r278 53 55 21.3027 $w=3.28e-07 $l=6.1e-07 $layer=LI1_cond $X=9.215 $Y=3.245
+ $X2=9.215 $Y2=2.635
r279 49 69 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.21 $Y=3.245
+ $X2=8.21 $Y2=3.33
r280 49 51 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=8.21 $Y=3.245
+ $X2=8.21 $Y2=2.815
r281 45 145 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.145 $Y=3.245
+ $X2=5.145 $Y2=3.33
r282 45 47 25.3537 $w=2.48e-07 $l=5.5e-07 $layer=LI1_cond $X=5.145 $Y=3.245
+ $X2=5.145 $Y2=2.695
r283 44 142 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.18 $Y=3.33
+ $X2=4.055 $Y2=3.33
r284 43 145 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.02 $Y=3.33
+ $X2=5.145 $Y2=3.33
r285 43 44 54.8021 $w=1.68e-07 $l=8.4e-07 $layer=LI1_cond $X=5.02 $Y=3.33
+ $X2=4.18 $Y2=3.33
r286 39 142 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.055 $Y=3.245
+ $X2=4.055 $Y2=3.33
r287 39 41 36.4172 $w=2.48e-07 $l=7.9e-07 $layer=LI1_cond $X=4.055 $Y=3.245
+ $X2=4.055 $Y2=2.455
r288 35 139 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.595 $Y=3.245
+ $X2=2.595 $Y2=3.33
r289 35 37 35.9562 $w=2.48e-07 $l=7.8e-07 $layer=LI1_cond $X=2.595 $Y=3.245
+ $X2=2.595 $Y2=2.465
r290 31 136 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.73 $Y=3.245
+ $X2=0.73 $Y2=3.33
r291 31 33 27.0649 $w=3.28e-07 $l=7.75e-07 $layer=LI1_cond $X=0.73 $Y=3.245
+ $X2=0.73 $Y2=2.47
r292 10 66 600 $w=1.7e-07 $l=1.00566e-06 $layer=licon1_PDIFF $count=1 $X=15.835
+ $Y=1.92 $X2=16.07 $Y2=2.815
r293 10 63 300 $w=1.7e-07 $l=2.98831e-07 $layer=licon1_PDIFF $count=2 $X=15.835
+ $Y=1.92 $X2=16.07 $Y2=2.065
r294 9 59 300 $w=1.7e-07 $l=6.68019e-07 $layer=licon1_PDIFF $count=2 $X=14.015
+ $Y=2.32 $X2=14.525 $Y2=2.685
r295 8 151 600 $w=1.7e-07 $l=1.20679e-06 $layer=licon1_PDIFF $count=1 $X=11.925
+ $Y=1.96 $X2=12.16 $Y2=3.055
r296 7 71 600 $w=1.7e-07 $l=6.2149e-07 $layer=licon1_PDIFF $count=1 $X=10.83
+ $Y=2.54 $X2=11.065 $Y2=3.055
r297 6 55 600 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=1 $X=9.07
+ $Y=2.12 $X2=9.215 $Y2=2.635
r298 5 51 600 $w=1.7e-07 $l=7.66339e-07 $layer=licon1_PDIFF $count=1 $X=8.06
+ $Y=2.12 $X2=8.21 $Y2=2.815
r299 4 47 600 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_PDIFF $count=1 $X=4.96
+ $Y=2.485 $X2=5.105 $Y2=2.695
r300 3 41 300 $w=1.7e-07 $l=6.85912e-07 $layer=licon1_PDIFF $count=2 $X=3.945
+ $Y=1.84 $X2=4.095 $Y2=2.455
r301 2 37 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=2.49
+ $Y=2.32 $X2=2.635 $Y2=2.465
r302 1 33 300 $w=1.7e-07 $l=2.12132e-07 $layer=licon1_PDIFF $count=2 $X=0.58
+ $Y=2.32 $X2=0.73 $Y2=2.47
.ends

.subckt PM_SKY130_FD_SC_HS__SDFBBN_1%A_197_119# 1 2 3 4 13 15 17 21 23 24 26 27
+ 30 31 32 34 35 36 38 39 40 42 43 44 48 49 51 52 54 56 60 61 65 66
c226 61 0 1.93711e-19 $X=1.57 $Y=0.95
c227 54 0 4.35224e-20 $X=7.505 $Y=2.31
c228 52 0 2.87426e-20 $X=6.925 $Y=0.875
c229 49 0 1.54972e-19 $X=7.42 $Y=2.395
c230 44 0 4.28297e-20 $X=5.97 $Y=0.34
c231 39 0 2.29882e-20 $X=5.8 $Y=1.29
c232 13 0 2.95072e-20 $X=1.485 $Y=0.95
r233 66 69 4.36531 $w=3.28e-07 $l=1.25e-07 $layer=LI1_cond $X=6.53 $Y=2.395
+ $X2=6.53 $Y2=2.52
r234 61 63 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=1.57 $Y=0.95
+ $X2=1.57 $Y2=1.225
r235 56 58 5.06376 $w=3.28e-07 $l=1.45e-07 $layer=LI1_cond $X=1.125 $Y=0.805
+ $X2=1.125 $Y2=0.95
r236 53 54 88.0749 $w=1.68e-07 $l=1.35e-06 $layer=LI1_cond $X=7.505 $Y=0.96
+ $X2=7.505 $Y2=2.31
r237 51 53 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.42 $Y=0.875
+ $X2=7.505 $Y2=0.96
r238 51 52 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=7.42 $Y=0.875
+ $X2=6.925 $Y2=0.875
r239 50 66 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.695 $Y=2.395
+ $X2=6.53 $Y2=2.395
r240 49 54 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.42 $Y=2.395
+ $X2=7.505 $Y2=2.31
r241 49 50 47.2995 $w=1.68e-07 $l=7.25e-07 $layer=LI1_cond $X=7.42 $Y=2.395
+ $X2=6.695 $Y2=2.395
r242 46 52 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=6.76 $Y=0.79
+ $X2=6.925 $Y2=0.875
r243 46 48 0.873063 $w=3.28e-07 $l=2.5e-08 $layer=LI1_cond $X=6.76 $Y=0.79
+ $X2=6.76 $Y2=0.765
r244 45 48 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=6.76 $Y=0.425
+ $X2=6.76 $Y2=0.765
r245 43 45 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=6.595 $Y=0.34
+ $X2=6.76 $Y2=0.425
r246 43 44 40.7754 $w=1.68e-07 $l=6.25e-07 $layer=LI1_cond $X=6.595 $Y=0.34
+ $X2=5.97 $Y2=0.34
r247 41 44 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.885 $Y=0.425
+ $X2=5.97 $Y2=0.34
r248 41 42 50.8877 $w=1.68e-07 $l=7.8e-07 $layer=LI1_cond $X=5.885 $Y=0.425
+ $X2=5.885 $Y2=1.205
r249 39 42 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.8 $Y=1.29
+ $X2=5.885 $Y2=1.205
r250 39 40 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.8 $Y=1.29
+ $X2=5.13 $Y2=1.29
r251 38 40 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.045 $Y=1.205
+ $X2=5.13 $Y2=1.29
r252 37 38 29.6845 $w=1.68e-07 $l=4.55e-07 $layer=LI1_cond $X=5.045 $Y=0.75
+ $X2=5.045 $Y2=1.205
r253 35 37 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.96 $Y=0.665
+ $X2=5.045 $Y2=0.75
r254 35 36 101.775 $w=1.68e-07 $l=1.56e-06 $layer=LI1_cond $X=4.96 $Y=0.665
+ $X2=3.4 $Y2=0.665
r255 34 36 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.315 $Y=0.58
+ $X2=3.4 $Y2=0.665
r256 33 34 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=3.315 $Y=0.425
+ $X2=3.315 $Y2=0.58
r257 31 33 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.23 $Y=0.34
+ $X2=3.315 $Y2=0.425
r258 31 32 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.23 $Y=0.34
+ $X2=2.56 $Y2=0.34
r259 29 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.475 $Y=0.425
+ $X2=2.56 $Y2=0.34
r260 29 30 46.6471 $w=1.68e-07 $l=7.15e-07 $layer=LI1_cond $X=2.475 $Y=0.425
+ $X2=2.475 $Y2=1.14
r261 28 65 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.155 $Y=1.225
+ $X2=2.07 $Y2=1.225
r262 27 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.39 $Y=1.225
+ $X2=2.475 $Y2=1.14
r263 27 28 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=2.39 $Y=1.225
+ $X2=2.155 $Y2=1.225
r264 25 65 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.07 $Y=1.31
+ $X2=2.07 $Y2=1.225
r265 25 26 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.07 $Y=1.31
+ $X2=2.07 $Y2=1.98
r266 23 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.985 $Y=2.065
+ $X2=2.07 $Y2=1.98
r267 23 24 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=1.985 $Y=2.065
+ $X2=1.715 $Y2=2.065
r268 22 63 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.655 $Y=1.225
+ $X2=1.57 $Y2=1.225
r269 21 65 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.985 $Y=1.225
+ $X2=2.07 $Y2=1.225
r270 21 22 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=1.985 $Y=1.225
+ $X2=1.655 $Y2=1.225
r271 19 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.63 $Y=2.15
+ $X2=1.715 $Y2=2.065
r272 19 60 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=1.63 $Y=2.15
+ $X2=1.63 $Y2=2.3
r273 15 60 6.94937 $w=2.48e-07 $l=1.25e-07 $layer=LI1_cond $X=1.59 $Y=2.425
+ $X2=1.59 $Y2=2.3
r274 15 17 4.14879 $w=2.48e-07 $l=9e-08 $layer=LI1_cond $X=1.59 $Y=2.425
+ $X2=1.59 $Y2=2.515
r275 14 58 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.29 $Y=0.95
+ $X2=1.125 $Y2=0.95
r276 13 61 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.485 $Y=0.95
+ $X2=1.57 $Y2=0.95
r277 13 14 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=1.485 $Y=0.95
+ $X2=1.29 $Y2=0.95
r278 4 69 600 $w=1.7e-07 $l=3.40624e-07 $layer=licon1_PDIFF $count=1 $X=6.33
+ $Y=2.265 $X2=6.53 $Y2=2.52
r279 3 17 600 $w=1.7e-07 $l=2.59374e-07 $layer=licon1_PDIFF $count=1 $X=1.48
+ $Y=2.32 $X2=1.63 $Y2=2.515
r280 2 48 182 $w=1.7e-07 $l=2.87706e-07 $layer=licon1_NDIFF $count=1 $X=6.545
+ $Y=0.595 $X2=6.76 $Y2=0.765
r281 1 56 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=0.985
+ $Y=0.595 $X2=1.125 $Y2=0.805
.ends

.subckt PM_SKY130_FD_SC_HS__SDFBBN_1%Q_N 1 2 9 13 14 15 16 23 33
r35 21 35 0.808207 $w=3.83e-07 $l=2.7e-08 $layer=LI1_cond $X=15.082 $Y=2.012
+ $X2=15.082 $Y2=1.985
r36 21 23 0.688472 $w=3.83e-07 $l=2.3e-08 $layer=LI1_cond $X=15.082 $Y=2.012
+ $X2=15.082 $Y2=2.035
r37 16 30 1.19734 $w=3.83e-07 $l=4e-08 $layer=LI1_cond $X=15.082 $Y=2.775
+ $X2=15.082 $Y2=2.815
r38 15 16 11.0754 $w=3.83e-07 $l=3.7e-07 $layer=LI1_cond $X=15.082 $Y=2.405
+ $X2=15.082 $Y2=2.775
r39 14 35 0.119734 $w=3.83e-07 $l=4e-09 $layer=LI1_cond $X=15.082 $Y=1.981
+ $X2=15.082 $Y2=1.985
r40 14 33 8.4692 $w=3.83e-07 $l=1.61e-07 $layer=LI1_cond $X=15.082 $Y=1.981
+ $X2=15.082 $Y2=1.82
r41 14 15 10.1475 $w=3.83e-07 $l=3.39e-07 $layer=LI1_cond $X=15.082 $Y=2.066
+ $X2=15.082 $Y2=2.405
r42 14 23 0.927941 $w=3.83e-07 $l=3.1e-08 $layer=LI1_cond $X=15.082 $Y=2.066
+ $X2=15.082 $Y2=2.035
r43 13 33 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=15.19 $Y=1.13
+ $X2=15.19 $Y2=1.82
r44 7 13 8.99121 $w=3.58e-07 $l=1.8e-07 $layer=LI1_cond $X=15.095 $Y=0.95
+ $X2=15.095 $Y2=1.13
r45 7 9 13.9254 $w=3.58e-07 $l=4.35e-07 $layer=LI1_cond $X=15.095 $Y=0.95
+ $X2=15.095 $Y2=0.515
r46 2 35 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=14.825
+ $Y=1.84 $X2=14.975 $Y2=1.985
r47 2 30 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=14.825
+ $Y=1.84 $X2=14.975 $Y2=2.815
r48 1 9 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=14.86
+ $Y=0.37 $X2=15 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__SDFBBN_1%Q 1 2 9 13 14 15 16 23 32
r23 21 23 1.12043 $w=3.58e-07 $l=3.5e-08 $layer=LI1_cond $X=16.535 $Y=2
+ $X2=16.535 $Y2=2.035
r24 15 16 11.8446 $w=3.58e-07 $l=3.7e-07 $layer=LI1_cond $X=16.535 $Y=2.405
+ $X2=16.535 $Y2=2.775
r25 14 21 0.800308 $w=3.58e-07 $l=2.5e-08 $layer=LI1_cond $X=16.535 $Y=1.975
+ $X2=16.535 $Y2=2
r26 14 32 8.1909 $w=3.58e-07 $l=1.55e-07 $layer=LI1_cond $X=16.535 $Y=1.975
+ $X2=16.535 $Y2=1.82
r27 14 15 11.0442 $w=3.58e-07 $l=3.45e-07 $layer=LI1_cond $X=16.535 $Y=2.06
+ $X2=16.535 $Y2=2.405
r28 14 23 0.800308 $w=3.58e-07 $l=2.5e-08 $layer=LI1_cond $X=16.535 $Y=2.06
+ $X2=16.535 $Y2=2.035
r29 13 32 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=16.63 $Y=1.05
+ $X2=16.63 $Y2=1.82
r30 7 13 9.32938 $w=3.78e-07 $l=1.9e-07 $layer=LI1_cond $X=16.525 $Y=0.86
+ $X2=16.525 $Y2=1.05
r31 7 9 10.463 $w=3.78e-07 $l=3.45e-07 $layer=LI1_cond $X=16.525 $Y=0.86
+ $X2=16.525 $Y2=0.515
r32 2 14 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=16.37
+ $Y=1.84 $X2=16.52 $Y2=1.985
r33 2 16 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=16.37
+ $Y=1.84 $X2=16.52 $Y2=2.815
r34 1 9 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=16.36
+ $Y=0.37 $X2=16.5 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__SDFBBN_1%VGND 1 2 3 4 5 6 7 8 25 27 31 35 39 43 47
+ 51 52 59 60 61 63 71 76 81 96 108 109 115 119 125 128 131
c171 109 0 3.18534e-20 $X=16.56 $Y=0
r172 131 132 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=14.64 $Y=0
+ $X2=14.64 $Y2=0
r173 128 129 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=0
+ $X2=8.88 $Y2=0
r174 125 126 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=0
+ $X2=5.52 $Y2=0
r175 119 122 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=3.965 $Y=0
+ $X2=3.965 $Y2=0.325
r176 119 120 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.08 $Y=0
+ $X2=4.08 $Y2=0
r177 115 116 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0
+ $X2=2.16 $Y2=0
r178 112 113 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0
+ $X2=0.24 $Y2=0
r179 108 109 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=16.56 $Y=0
+ $X2=16.56 $Y2=0
r180 106 109 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=15.6 $Y=0
+ $X2=16.56 $Y2=0
r181 106 132 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=15.6 $Y=0
+ $X2=14.64 $Y2=0
r182 105 106 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=15.6 $Y=0
+ $X2=15.6 $Y2=0
r183 103 131 8.42608 $w=1.7e-07 $l=1.6e-07 $layer=LI1_cond $X=14.735 $Y=0
+ $X2=14.575 $Y2=0
r184 103 105 56.4332 $w=1.68e-07 $l=8.65e-07 $layer=LI1_cond $X=14.735 $Y=0
+ $X2=15.6 $Y2=0
r185 102 132 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=14.16 $Y=0
+ $X2=14.64 $Y2=0
r186 101 102 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=14.16 $Y=0
+ $X2=14.16 $Y2=0
r187 99 102 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=11.76 $Y=0
+ $X2=14.16 $Y2=0
r188 98 101 156.578 $w=1.68e-07 $l=2.4e-06 $layer=LI1_cond $X=11.76 $Y=0
+ $X2=14.16 $Y2=0
r189 98 99 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=11.76 $Y=0
+ $X2=11.76 $Y2=0
r190 96 131 8.42608 $w=1.7e-07 $l=1.6e-07 $layer=LI1_cond $X=14.415 $Y=0
+ $X2=14.575 $Y2=0
r191 96 101 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=14.415 $Y=0
+ $X2=14.16 $Y2=0
r192 95 99 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.28 $Y=0
+ $X2=11.76 $Y2=0
r193 94 95 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=11.28 $Y=0
+ $X2=11.28 $Y2=0
r194 92 95 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=9.36 $Y=0
+ $X2=11.28 $Y2=0
r195 92 129 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.36 $Y=0
+ $X2=8.88 $Y2=0
r196 91 94 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=9.36 $Y=0
+ $X2=11.28 $Y2=0
r197 91 92 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=9.36 $Y=0
+ $X2=9.36 $Y2=0
r198 89 128 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.125 $Y=0
+ $X2=8.96 $Y2=0
r199 89 91 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=9.125 $Y=0
+ $X2=9.36 $Y2=0
r200 85 126 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=0 $X2=5.52
+ $Y2=0
r201 84 87 156.578 $w=1.68e-07 $l=2.4e-06 $layer=LI1_cond $X=6 $Y=0 $X2=8.4
+ $Y2=0
r202 84 85 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=6 $Y=0 $X2=6 $Y2=0
r203 82 125 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.63 $Y=0
+ $X2=5.465 $Y2=0
r204 82 84 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=5.63 $Y=0 $X2=6
+ $Y2=0
r205 81 128 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.795 $Y=0
+ $X2=8.96 $Y2=0
r206 81 87 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=8.795 $Y=0 $X2=8.4
+ $Y2=0
r207 80 126 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=0
+ $X2=5.52 $Y2=0
r208 80 120 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.04 $Y=0
+ $X2=4.08 $Y2=0
r209 79 80 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r210 77 119 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.13 $Y=0
+ $X2=3.965 $Y2=0
r211 77 79 59.369 $w=1.68e-07 $l=9.1e-07 $layer=LI1_cond $X=4.13 $Y=0 $X2=5.04
+ $Y2=0
r212 76 125 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.3 $Y=0 $X2=5.465
+ $Y2=0
r213 76 79 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=5.3 $Y=0 $X2=5.04
+ $Y2=0
r214 75 120 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.08
+ $Y2=0
r215 75 116 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=3.6 $Y=0
+ $X2=2.16 $Y2=0
r216 74 75 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r217 72 115 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.22 $Y=0
+ $X2=2.055 $Y2=0
r218 72 74 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=2.22 $Y=0 $X2=3.6
+ $Y2=0
r219 71 119 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.8 $Y=0 $X2=3.965
+ $Y2=0
r220 71 74 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=3.8 $Y=0 $X2=3.6
+ $Y2=0
r221 70 116 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0
+ $X2=2.16 $Y2=0
r222 69 70 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r223 67 70 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r224 67 113 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0
+ $X2=0.24 $Y2=0
r225 66 69 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r226 66 67 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r227 64 112 4.67962 $w=1.7e-07 $l=2.35e-07 $layer=LI1_cond $X=0.47 $Y=0
+ $X2=0.235 $Y2=0
r228 64 66 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=0.47 $Y=0 $X2=0.72
+ $Y2=0
r229 63 115 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.89 $Y=0
+ $X2=2.055 $Y2=0
r230 63 69 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=1.89 $Y=0 $X2=1.68
+ $Y2=0
r231 61 129 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=0 $X2=8.88
+ $Y2=0
r232 61 85 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=8.4 $Y=0 $X2=6
+ $Y2=0
r233 61 87 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r234 59 105 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=15.905 $Y=0
+ $X2=15.6 $Y2=0
r235 59 60 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=15.905 $Y=0
+ $X2=16.03 $Y2=0
r236 58 108 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=16.155 $Y=0
+ $X2=16.56 $Y2=0
r237 58 60 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=16.155 $Y=0
+ $X2=16.03 $Y2=0
r238 54 98 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=11.755 $Y=0
+ $X2=11.76 $Y2=0
r239 52 94 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=11.415 $Y=0
+ $X2=11.28 $Y2=0
r240 51 56 11.016 $w=3.38e-07 $l=3.25e-07 $layer=LI1_cond $X=11.585 $Y=0
+ $X2=11.585 $Y2=0.325
r241 51 54 4.80115 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=11.585 $Y=0
+ $X2=11.755 $Y2=0
r242 51 52 4.80115 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=11.585 $Y=0
+ $X2=11.415 $Y2=0
r243 47 49 17.0562 $w=2.48e-07 $l=3.7e-07 $layer=LI1_cond $X=16.03 $Y=0.515
+ $X2=16.03 $Y2=0.885
r244 45 60 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=16.03 $Y=0.085
+ $X2=16.03 $Y2=0
r245 45 47 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=16.03 $Y=0.085
+ $X2=16.03 $Y2=0.515
r246 41 131 0.800721 $w=3.2e-07 $l=8.5e-08 $layer=LI1_cond $X=14.575 $Y=0.085
+ $X2=14.575 $Y2=0
r247 41 43 15.486 $w=3.18e-07 $l=4.3e-07 $layer=LI1_cond $X=14.575 $Y=0.085
+ $X2=14.575 $Y2=0.515
r248 37 128 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.96 $Y=0.085
+ $X2=8.96 $Y2=0
r249 37 39 26.5411 $w=3.28e-07 $l=7.6e-07 $layer=LI1_cond $X=8.96 $Y=0.085
+ $X2=8.96 $Y2=0.845
r250 33 125 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.465 $Y=0.085
+ $X2=5.465 $Y2=0
r251 33 35 25.1442 $w=3.28e-07 $l=7.2e-07 $layer=LI1_cond $X=5.465 $Y=0.085
+ $X2=5.465 $Y2=0.805
r252 29 115 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.055 $Y=0.085
+ $X2=2.055 $Y2=0
r253 29 31 23.9219 $w=3.28e-07 $l=6.85e-07 $layer=LI1_cond $X=2.055 $Y=0.085
+ $X2=2.055 $Y2=0.77
r254 25 112 3.08656 $w=3.3e-07 $l=1.14782e-07 $layer=LI1_cond $X=0.305 $Y=0.085
+ $X2=0.235 $Y2=0
r255 25 27 25.1442 $w=3.28e-07 $l=7.2e-07 $layer=LI1_cond $X=0.305 $Y=0.085
+ $X2=0.305 $Y2=0.805
r256 8 49 182 $w=1.7e-07 $l=6.15244e-07 $layer=licon1_NDIFF $count=1 $X=15.85
+ $Y=0.37 $X2=16.07 $Y2=0.885
r257 8 47 182 $w=1.7e-07 $l=2.83373e-07 $layer=licon1_NDIFF $count=1 $X=15.85
+ $Y=0.37 $X2=16.07 $Y2=0.515
r258 7 43 182 $w=1.7e-07 $l=5.04975e-07 $layer=licon1_NDIFF $count=1 $X=14.11
+ $Y=0.69 $X2=14.535 $Y2=0.515
r259 6 56 182 $w=1.7e-07 $l=3.65582e-07 $layer=licon1_NDIFF $count=1 $X=11.36
+ $Y=0.595 $X2=11.585 $Y2=0.325
r260 5 39 182 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=1 $X=8.82
+ $Y=0.595 $X2=8.96 $Y2=0.845
r261 4 35 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=5.32
+ $Y=0.595 $X2=5.465 $Y2=0.805
r262 3 122 182 $w=1.7e-07 $l=2.59037e-07 $layer=licon1_NDIFF $count=1 $X=3.745
+ $Y=0.41 $X2=3.965 $Y2=0.325
r263 2 31 182 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_NDIFF $count=1 $X=1.915
+ $Y=0.595 $X2=2.055 $Y2=0.77
r264 1 27 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=0.16
+ $Y=0.595 $X2=0.305 $Y2=0.805
.ends

.subckt PM_SKY130_FD_SC_HS__SDFBBN_1%A_1434_78# 1 2 7 11 13
r29 13 16 6.80989 $w=3.28e-07 $l=1.95e-07 $layer=LI1_cond $X=7.315 $Y=0.34
+ $X2=7.315 $Y2=0.535
r30 9 11 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=8.425 $Y=0.425
+ $X2=8.425 $Y2=0.855
r31 8 13 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.48 $Y=0.34
+ $X2=7.315 $Y2=0.34
r32 7 9 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=8.26 $Y=0.34
+ $X2=8.425 $Y2=0.425
r33 7 8 50.8877 $w=1.68e-07 $l=7.8e-07 $layer=LI1_cond $X=8.26 $Y=0.34 $X2=7.48
+ $Y2=0.34
r34 2 11 182 $w=1.7e-07 $l=3.49571e-07 $layer=licon1_NDIFF $count=1 $X=8.215
+ $Y=0.595 $X2=8.425 $Y2=0.855
r35 1 16 182 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=1 $X=7.17
+ $Y=0.39 $X2=7.315 $Y2=0.535
.ends

.subckt PM_SKY130_FD_SC_HS__SDFBBN_1%A_2392_74# 1 2 9 11 12 13
r31 13 16 5.30124 $w=2.48e-07 $l=1.15e-07 $layer=LI1_cond $X=13.1 $Y=0.34
+ $X2=13.1 $Y2=0.455
r32 11 13 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=12.975 $Y=0.34
+ $X2=13.1 $Y2=0.34
r33 11 12 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=12.975 $Y=0.34
+ $X2=12.265 $Y2=0.34
r34 7 12 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=12.1 $Y=0.425
+ $X2=12.265 $Y2=0.34
r35 7 9 2.44458 $w=3.28e-07 $l=7e-08 $layer=LI1_cond $X=12.1 $Y=0.425 $X2=12.1
+ $Y2=0.495
r36 2 16 182 $w=1.7e-07 $l=2.59037e-07 $layer=licon1_NDIFF $count=1 $X=12.92
+ $Y=0.37 $X2=13.14 $Y2=0.455
r37 1 9 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=11.96
+ $Y=0.37 $X2=12.1 $Y2=0.495
.ends

