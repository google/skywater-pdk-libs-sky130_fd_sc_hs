* File: sky130_fd_sc_hs__sdfsbp_2.spice
* Created: Thu Aug 27 21:09:16 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hs__sdfsbp_2.pex.spice"
.subckt sky130_fd_sc_hs__sdfsbp_2  VNB VPB SCE D SCD CLK SET_B VPWR Q_N Q VGND
* 
* VGND	VGND
* Q	Q
* Q_N	Q_N
* VPWR	VPWR
* SET_B	SET_B
* CLK	CLK
* SCD	SCD
* D	D
* SCE	SCE
* VPB	VPB
* VNB	VNB
MM1046 N_VGND_M1046_d N_SCE_M1046_g N_A_27_74#_M1046_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.08925 AS=0.1197 PD=0.845 PS=1.41 NRD=30 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75002.5 A=0.063 P=1.14 MULT=1
MM1035 A_229_74# N_A_27_74#_M1035_g N_VGND_M1046_d VNB NLOWVT L=0.15 W=0.42
+ AD=0.0504 AS=0.08925 PD=0.66 PS=0.845 NRD=18.564 NRS=11.424 M=1 R=2.8
+ SA=75000.8 SB=75001.9 A=0.063 P=1.14 MULT=1
MM1036 N_A_304_464#_M1036_d N_D_M1036_g A_229_74# VNB NLOWVT L=0.15 W=0.42
+ AD=0.1659 AS=0.0504 PD=1.21 PS=0.66 NRD=137.136 NRS=18.564 M=1 R=2.8
+ SA=75001.2 SB=75001.5 A=0.063 P=1.14 MULT=1
MM1017 A_495_74# N_SCE_M1017_g N_A_304_464#_M1036_d VNB NLOWVT L=0.15 W=0.42
+ AD=0.0504 AS=0.1659 PD=0.66 PS=1.21 NRD=18.564 NRS=8.568 M=1 R=2.8 SA=75002.1
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1014 N_VGND_M1014_d N_SCD_M1014_g A_495_74# VNB NLOWVT L=0.15 W=0.42 AD=0.1197
+ AS=0.0504 PD=1.41 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75002.5 SB=75000.2
+ A=0.063 P=1.14 MULT=1
MM1040 N_VGND_M1040_d N_CLK_M1040_g N_A_619_368#_M1040_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1295 AS=0.2109 PD=1.09 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75000.7 A=0.111 P=1.78 MULT=1
MM1031 N_A_871_74#_M1031_d N_A_619_368#_M1031_g N_VGND_M1040_d VNB NLOWVT L=0.15
+ W=0.74 AD=0.2109 AS=0.1295 PD=2.05 PS=1.09 NRD=0 NRS=11.34 M=1 R=4.93333
+ SA=75000.7 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1020 N_A_1069_81#_M1020_d N_A_619_368#_M1020_g N_A_304_464#_M1020_s VNB NLOWVT
+ L=0.15 W=0.42 AD=0.18375 AS=0.1197 PD=1.295 PS=1.41 NRD=142.848 NRS=0 M=1
+ R=2.8 SA=75000.2 SB=75001.7 A=0.063 P=1.14 MULT=1
MM1028 A_1274_81# N_A_871_74#_M1028_g N_A_1069_81#_M1020_d VNB NLOWVT L=0.15
+ W=0.42 AD=0.0504 AS=0.18375 PD=0.66 PS=1.295 NRD=18.564 NRS=27.132 M=1 R=2.8
+ SA=75001.2 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1025 N_VGND_M1025_d N_A_1252_376#_M1025_g A_1274_81# VNB NLOWVT L=0.15 W=0.42
+ AD=0.1554 AS=0.0504 PD=1.58 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75001.6
+ SB=75000.3 A=0.063 P=1.14 MULT=1
MM1012 A_1567_74# N_A_1069_81#_M1012_g N_A_1252_376#_M1012_s VNB NLOWVT L=0.15
+ W=0.42 AD=0.0504 AS=0.1197 PD=0.66 PS=1.41 NRD=18.564 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75000.8 A=0.063 P=1.14 MULT=1
MM1013 N_VGND_M1013_d N_SET_B_M1013_g A_1567_74# VNB NLOWVT L=0.15 W=0.42
+ AD=0.189 AS=0.0504 PD=1.74 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75000.6
+ SB=75000.4 A=0.063 P=1.14 MULT=1
MM1001 N_VGND_M1001_d N_A_1069_81#_M1001_g N_A_1794_74#_M1001_s VNB NLOWVT
+ L=0.15 W=0.64 AD=0.096 AS=0.2144 PD=0.94 PS=1.95 NRD=3.744 NRS=9.372 M=1
+ R=4.26667 SA=75000.3 SB=75001.7 A=0.096 P=1.58 MULT=1
MM1006 N_VGND_M1001_d N_A_1069_81#_M1006_g N_A_1794_74#_M1006_s VNB NLOWVT
+ L=0.15 W=0.64 AD=0.096 AS=0.0896 PD=0.94 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.7 SB=75001.2 A=0.096 P=1.58 MULT=1
MM1030 N_A_1794_74#_M1006_s N_A_871_74#_M1030_g N_A_2067_74#_M1030_s VNB NLOWVT
+ L=0.15 W=0.64 AD=0.0896 AS=0.112 PD=0.92 PS=0.99 NRD=0 NRS=13.116 M=1
+ R=4.26667 SA=75001.1 SB=75000.8 A=0.096 P=1.58 MULT=1
MM1038 N_A_1794_74#_M1038_d N_A_871_74#_M1038_g N_A_2067_74#_M1030_s VNB NLOWVT
+ L=0.15 W=0.64 AD=0.2272 AS=0.112 PD=1.99 PS=0.99 NRD=13.116 NRS=0 M=1
+ R=4.26667 SA=75001.6 SB=75000.3 A=0.096 P=1.58 MULT=1
MM1003 A_2501_74# N_A_619_368#_M1003_g N_A_2067_74#_M1003_s VNB NLOWVT L=0.15
+ W=0.42 AD=0.0504 AS=0.3759 PD=0.66 PS=2.63 NRD=18.564 NRS=0 M=1 R=2.8
+ SA=75000.8 SB=75001.5 A=0.063 P=1.14 MULT=1
MM1021 A_2579_74# N_A_2513_258#_M1021_g A_2501_74# VNB NLOWVT L=0.15 W=0.42
+ AD=0.0504 AS=0.0504 PD=0.66 PS=0.66 NRD=18.564 NRS=18.564 M=1 R=2.8 SA=75001.2
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1022 N_VGND_M1022_d N_SET_B_M1022_g A_2579_74# VNB NLOWVT L=0.15 W=0.42
+ AD=0.0756 AS=0.0504 PD=0.78 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75001.6
+ SB=75000.7 A=0.063 P=1.14 MULT=1
MM1039 N_A_2513_258#_M1039_d N_A_2067_74#_M1039_g N_VGND_M1022_d VNB NLOWVT
+ L=0.15 W=0.42 AD=0.1197 AS=0.0756 PD=1.41 PS=0.78 NRD=0 NRS=22.848 M=1 R=2.8
+ SA=75002.1 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1024 N_Q_N_M1024_d N_A_2067_74#_M1024_g N_VGND_M1024_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.111 AS=0.2479 PD=1.04 PS=2.15 NRD=3.24 NRS=8.1 M=1 R=4.93333
+ SA=75000.3 SB=75000.7 A=0.111 P=1.78 MULT=1
MM1026 N_Q_N_M1024_d N_A_2067_74#_M1026_g N_VGND_M1026_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.111 AS=0.2442 PD=1.04 PS=2.14 NRD=0 NRS=7.296 M=1 R=4.93333
+ SA=75000.7 SB=75000.3 A=0.111 P=1.78 MULT=1
MM1010 N_VGND_M1010_d N_A_2067_74#_M1010_g N_A_3177_368#_M1010_s VNB NLOWVT
+ L=0.15 W=0.64 AD=0.136394 AS=0.1824 PD=1.0713 PS=1.85 NRD=25.776 NRS=0 M=1
+ R=4.26667 SA=75000.2 SB=75001.2 A=0.096 P=1.58 MULT=1
MM1000 N_VGND_M1010_d N_A_3177_368#_M1000_g N_Q_M1000_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.157706 AS=0.1036 PD=1.2387 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.7
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1023 N_VGND_M1023_d N_A_3177_368#_M1023_g N_Q_M1000_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.1036 PD=2.05 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.1
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1043 N_VPWR_M1043_d N_SCE_M1043_g N_A_27_74#_M1043_s VPB PSHORT L=0.15 W=0.64
+ AD=0.112 AS=0.1888 PD=0.99 PS=1.87 NRD=18.4589 NRS=3.0732 M=1 R=4.26667
+ SA=75000.2 SB=75002.1 A=0.096 P=1.58 MULT=1
MM1037 A_220_464# N_SCE_M1037_g N_VPWR_M1043_d VPB PSHORT L=0.15 W=0.64
+ AD=0.0864 AS=0.112 PD=0.91 PS=0.99 NRD=24.625 NRS=3.0732 M=1 R=4.26667
+ SA=75000.7 SB=75001.6 A=0.096 P=1.58 MULT=1
MM1048 N_A_304_464#_M1048_d N_D_M1048_g A_220_464# VPB PSHORT L=0.15 W=0.64
+ AD=0.1344 AS=0.0864 PD=1.06 PS=0.91 NRD=21.5321 NRS=24.625 M=1 R=4.26667
+ SA=75001.1 SB=75001.2 A=0.096 P=1.58 MULT=1
MM1044 A_418_464# N_A_27_74#_M1044_g N_A_304_464#_M1048_d VPB PSHORT L=0.15
+ W=0.64 AD=0.0864 AS=0.1344 PD=0.91 PS=1.06 NRD=24.625 NRS=21.5321 M=1
+ R=4.26667 SA=75001.7 SB=75000.7 A=0.096 P=1.58 MULT=1
MM1018 N_VPWR_M1018_d N_SCD_M1018_g A_418_464# VPB PSHORT L=0.15 W=0.64
+ AD=0.2016 AS=0.0864 PD=1.91 PS=0.91 NRD=6.1464 NRS=24.625 M=1 R=4.26667
+ SA=75002.1 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1049 N_VPWR_M1049_d N_CLK_M1049_g N_A_619_368#_M1049_s VPB PSHORT L=0.15
+ W=1.12 AD=0.3808 AS=0.3304 PD=1.8 PS=2.83 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75001.1 A=0.168 P=2.54 MULT=1
MM1004 N_A_871_74#_M1004_d N_A_619_368#_M1004_g N_VPWR_M1049_d VPB PSHORT L=0.15
+ W=1.12 AD=0.3696 AS=0.3808 PD=2.9 PS=1.8 NRD=7.8997 NRS=4.3931 M=1 R=7.46667
+ SA=75001 SB=75000.3 A=0.168 P=2.54 MULT=1
MM1033 N_A_1069_81#_M1033_d N_A_871_74#_M1033_g N_A_304_464#_M1033_s VPB PSHORT
+ L=0.15 W=0.42 AD=0.0735 AS=0.1239 PD=0.77 PS=1.43 NRD=28.1316 NRS=4.6886 M=1
+ R=2.8 SA=75000.2 SB=75003.1 A=0.063 P=1.14 MULT=1
MM1034 A_1201_463# N_A_619_368#_M1034_g N_A_1069_81#_M1033_d VPB PSHORT L=0.15
+ W=0.42 AD=0.0567 AS=0.0735 PD=0.69 PS=0.77 NRD=37.5088 NRS=4.6886 M=1 R=2.8
+ SA=75000.7 SB=75002.6 A=0.063 P=1.14 MULT=1
MM1045 N_VPWR_M1045_d N_A_1252_376#_M1045_g A_1201_463# VPB PSHORT L=0.15 W=0.42
+ AD=0.19635 AS=0.0567 PD=1.355 PS=0.69 NRD=60.9715 NRS=37.5088 M=1 R=2.8
+ SA=75001.1 SB=75002.1 A=0.063 P=1.14 MULT=1
MM1019 N_A_1252_376#_M1019_d N_A_1069_81#_M1019_g N_VPWR_M1045_d VPB PSHORT
+ L=0.15 W=0.42 AD=0.084 AS=0.19635 PD=0.82 PS=1.355 NRD=4.6886 NRS=246.25 M=1
+ R=2.8 SA=75002.2 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1007 N_VPWR_M1007_d N_SET_B_M1007_g N_A_1252_376#_M1019_d VPB PSHORT L=0.15
+ W=0.42 AD=0.2457 AS=0.084 PD=2.01 PS=0.82 NRD=140.697 NRS=51.5943 M=1 R=2.8
+ SA=75002.8 SB=75000.5 A=0.063 P=1.14 MULT=1
MM1008 N_VPWR_M1008_d N_A_1069_81#_M1008_g N_A_1789_424#_M1008_s VPB PSHORT
+ L=0.15 W=0.84 AD=0.126 AS=0.2898 PD=1.14 PS=2.37 NRD=2.3443 NRS=14.0658 M=1
+ R=5.6 SA=75000.3 SB=75001.6 A=0.126 P=1.98 MULT=1
MM1015 N_VPWR_M1008_d N_A_1069_81#_M1015_g N_A_1789_424#_M1015_s VPB PSHORT
+ L=0.15 W=0.84 AD=0.126 AS=0.126 PD=1.14 PS=1.14 NRD=2.3443 NRS=2.3443 M=1
+ R=5.6 SA=75000.7 SB=75001.1 A=0.126 P=1.98 MULT=1
MM1041 N_A_2067_74#_M1041_d N_A_619_368#_M1041_g N_A_1789_424#_M1015_s VPB
+ PSHORT L=0.15 W=0.84 AD=0.126 AS=0.126 PD=1.14 PS=1.14 NRD=2.3443 NRS=2.3443
+ M=1 R=5.6 SA=75001.2 SB=75000.7 A=0.126 P=1.98 MULT=1
MM1047 N_A_2067_74#_M1041_d N_A_619_368#_M1047_g N_A_1789_424#_M1047_s VPB
+ PSHORT L=0.15 W=0.84 AD=0.126 AS=0.2478 PD=1.14 PS=2.27 NRD=2.3443 NRS=2.3443
+ M=1 R=5.6 SA=75001.6 SB=75000.2 A=0.126 P=1.98 MULT=1
MM1027 N_A_2067_74#_M1027_d N_A_871_74#_M1027_g N_A_2277_455#_M1027_s VPB PSHORT
+ L=0.15 W=0.42 AD=0.1239 AS=0.126 PD=1.43 PS=1.44 NRD=4.6886 NRS=7.0329 M=1
+ R=2.8 SA=75000.2 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1029 N_VPWR_M1029_d N_A_2513_258#_M1029_g N_A_2277_455#_M1029_s VPB PSHORT
+ L=0.15 W=0.42 AD=0.063 AS=0.1239 PD=0.72 PS=1.43 NRD=4.6886 NRS=4.6886 M=1
+ R=2.8 SA=75000.2 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1032 N_A_2067_74#_M1032_d N_SET_B_M1032_g N_VPWR_M1029_d VPB PSHORT L=0.15
+ W=0.42 AD=0.1239 AS=0.063 PD=1.43 PS=0.72 NRD=4.6886 NRS=4.6886 M=1 R=2.8
+ SA=75000.7 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1002 N_VPWR_M1002_d N_A_2067_74#_M1002_g N_A_2513_258#_M1002_s VPB PSHORT
+ L=0.15 W=0.42 AD=0.100418 AS=0.1239 PD=0.820909 PS=1.43 NRD=119.599 NRS=0 M=1
+ R=2.8 SA=75000.2 SB=75001.2 A=0.063 P=1.14 MULT=1
MM1016 N_Q_N_M1016_d N_A_2067_74#_M1016_g N_VPWR_M1002_d VPB PSHORT L=0.15
+ W=1.12 AD=0.168 AS=0.267782 PD=1.42 PS=2.18909 NRD=1.7533 NRS=1.7533 M=1
+ R=7.46667 SA=75000.4 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1042 N_Q_N_M1016_d N_A_2067_74#_M1042_g N_VPWR_M1042_s VPB PSHORT L=0.15
+ W=1.12 AD=0.168 AS=0.3304 PD=1.42 PS=2.83 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.9 SB=75000.2 A=0.168 P=2.54 MULT=1
MM1011 N_VPWR_M1011_d N_A_2067_74#_M1011_g N_A_3177_368#_M1011_s VPB PSHORT
+ L=0.15 W=1 AD=0.205377 AS=0.295 PD=1.43396 PS=2.59 NRD=21.9852 NRS=1.9503 M=1
+ R=6.66667 SA=75000.2 SB=75001.2 A=0.15 P=2.3 MULT=1
MM1005 N_Q_M1005_d N_A_3177_368#_M1005_g N_VPWR_M1011_d VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.230023 PD=1.42 PS=1.60604 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.7 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1009 N_Q_M1005_d N_A_3177_368#_M1009_g N_VPWR_M1009_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.3304 PD=1.42 PS=2.83 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.2 SB=75000.2 A=0.168 P=2.54 MULT=1
DX50_noxref VNB VPB NWDIODE A=33.7404 P=40
c_372 VPB 0 1.49424e-19 $X=0 $Y=3.085
c_2372 A_1201_463# 0 1.69669e-19 $X=6.005 $Y=2.315
*
.include "sky130_fd_sc_hs__sdfsbp_2.pxi.spice"
*
.ends
*
*
