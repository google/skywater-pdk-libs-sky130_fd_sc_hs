# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_sc_hs__a31o_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__a31o_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.360000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.045000 1.490000 2.405000 1.800000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.535000 1.490000 1.865000 1.800000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.995000 1.490000 1.325000 1.800000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.565000 0.255000 2.815000 0.640000 ;
    END
  END B1
  PIN X
    ANTENNADIFFAREA  0.504100 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.480000 0.450000 1.180000 ;
        RECT 0.085000 1.180000 0.255000 1.850000 ;
        RECT 0.085000 1.850000 0.435000 2.980000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 3.360000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.000000 0.000000 3.360000 0.245000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.660000 3.550000 3.520000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 3.360000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.360000 0.085000 ;
      RECT 0.000000  3.245000 3.360000 3.415000 ;
      RECT 0.425000  1.350000 0.825000 1.680000 ;
      RECT 0.605000  1.970000 1.065000 3.245000 ;
      RECT 0.620000  0.085000 1.200000 0.980000 ;
      RECT 0.620000  1.150000 3.095000 1.320000 ;
      RECT 0.620000  1.320000 0.825000 1.350000 ;
      RECT 1.235000  1.970000 2.645000 2.140000 ;
      RECT 1.235000  2.140000 1.565000 2.980000 ;
      RECT 1.735000  2.310000 2.145000 3.245000 ;
      RECT 2.280000  0.810000 2.610000 1.150000 ;
      RECT 2.315000  2.140000 2.645000 2.980000 ;
      RECT 2.790000  0.810000 3.155000 0.980000 ;
      RECT 2.845000  1.320000 3.095000 2.980000 ;
      RECT 2.985000  0.085000 3.155000 0.810000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
  END
END sky130_fd_sc_hs__a31o_1
END LIBRARY
