* File: sky130_fd_sc_hs__sedfxbp_1.spice
* Created: Tue Sep  1 20:24:20 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hs__sedfxbp_1.pex.spice"
.subckt sky130_fd_sc_hs__sedfxbp_1  VNB VPB D DE SCD SCE CLK VPWR Q Q_N VGND
* 
* VGND	VGND
* Q_N	Q_N
* Q	Q
* VPWR	VPWR
* CLK	CLK
* SCE	SCE
* SCD	SCD
* DE	DE
* D	D
* VPB	VPB
* VNB	VNB
MM1022 A_157_90# N_D_M1022_g N_A_27_90#_M1022_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.0504 AS=0.21 PD=0.66 PS=1.84 NRD=18.564 NRS=0 M=1 R=2.8 SA=75000.4
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1023 N_VGND_M1023_d N_DE_M1023_g A_157_90# VNB NLOWVT L=0.15 W=0.42 AD=0.1197
+ AS=0.0504 PD=1.41 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75000.8 SB=75000.2
+ A=0.063 P=1.14 MULT=1
MM1014 N_VGND_M1014_d N_DE_M1014_g N_A_161_394#_M1014_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.0735 AS=0.1197 PD=0.77 PS=1.41 NRD=19.992 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.6 A=0.063 P=1.14 MULT=1
MM1011 A_533_113# N_A_161_394#_M1011_g N_VGND_M1014_d VNB NLOWVT L=0.15 W=0.42
+ AD=0.0504 AS=0.0735 PD=0.66 PS=0.77 NRD=18.564 NRS=0 M=1 R=2.8 SA=75000.7
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1005 N_A_27_90#_M1005_d N_A_575_305#_M1005_g A_533_113# VNB NLOWVT L=0.15
+ W=0.42 AD=0.0588 AS=0.0504 PD=0.7 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8
+ SA=75001.1 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1036 N_A_697_113#_M1036_d N_A_667_87#_M1036_g N_A_27_90#_M1005_d VNB NLOWVT
+ L=0.15 W=0.42 AD=0.1491 AS=0.0588 PD=1.55 PS=0.7 NRD=19.992 NRS=0 M=1 R=2.8
+ SA=75001.5 SB=75000.3 A=0.063 P=1.14 MULT=1
MM1043 N_VGND_M1043_d N_SCE_M1043_g N_A_667_87#_M1043_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.0756 AS=0.1197 PD=0.78 PS=1.41 NRD=19.992 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1033 A_1075_125# N_SCD_M1033_g N_VGND_M1043_d VNB NLOWVT L=0.15 W=0.42
+ AD=0.0504 AS=0.0756 PD=0.66 PS=0.78 NRD=18.564 NRS=2.856 M=1 R=2.8 SA=75000.7
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1012 N_A_697_113#_M1012_d N_SCE_M1012_g A_1075_125# VNB NLOWVT L=0.15 W=0.42
+ AD=0.1197 AS=0.0504 PD=1.41 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75001.1
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1025 N_A_1348_368#_M1025_d N_CLK_M1025_g N_VGND_M1025_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.2109 AS=0.2109 PD=2.05 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1008 N_A_1549_74#_M1008_d N_A_1348_368#_M1008_g N_VGND_M1008_s VNB NLOWVT
+ L=0.15 W=0.74 AD=0.2109 AS=0.2109 PD=2.05 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1000 N_A_1747_118#_M1000_d N_A_1348_368#_M1000_g N_A_697_113#_M1000_s VNB
+ NLOWVT L=0.15 W=0.42 AD=0.1239 AS=0.1197 PD=1.01 PS=1.41 NRD=79.992 NRS=0 M=1
+ R=2.8 SA=75000.2 SB=75002.3 A=0.063 P=1.14 MULT=1
MM1003 A_1895_118# N_A_1549_74#_M1003_g N_A_1747_118#_M1000_d VNB NLOWVT L=0.15
+ W=0.42 AD=0.08085 AS=0.1239 PD=0.805 PS=1.01 NRD=39.276 NRS=8.568 M=1 R=2.8
+ SA=75000.9 SB=75001.6 A=0.063 P=1.14 MULT=1
MM1031 N_VGND_M1031_d N_A_1972_92#_M1031_g A_1895_118# VNB NLOWVT L=0.15 W=0.42
+ AD=0.163364 AS=0.08085 PD=1.03811 PS=0.805 NRD=34.284 NRS=39.276 M=1 R=2.8
+ SA=75001.5 SB=75001 A=0.063 P=1.14 MULT=1
MM1041 N_A_1972_92#_M1041_d N_A_1747_118#_M1041_g N_VGND_M1031_d VNB NLOWVT
+ L=0.15 W=0.64 AD=0.192 AS=0.248936 PD=1.88 PS=1.58189 NRD=2.808 NRS=51.552 M=1
+ R=4.26667 SA=75001.7 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1026 A_2391_74# N_A_1972_92#_M1026_g N_VGND_M1026_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.0672 AS=0.1824 PD=0.85 PS=1.85 NRD=9.372 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75001.8 A=0.096 P=1.58 MULT=1
MM1028 N_A_2463_74#_M1028_d N_A_1549_74#_M1028_g A_2391_74# VNB NLOWVT L=0.15
+ W=0.64 AD=0.129147 AS=0.0672 PD=1.20755 PS=0.85 NRD=0 NRS=9.372 M=1 R=4.26667
+ SA=75000.6 SB=75001.5 A=0.096 P=1.58 MULT=1
MM1038 A_2565_74# N_A_1348_368#_M1038_g N_A_2463_74#_M1028_d VNB NLOWVT L=0.15
+ W=0.42 AD=0.0504 AS=0.0847528 PD=0.66 PS=0.792453 NRD=18.564 NRS=23.568 M=1
+ R=2.8 SA=75001.1 SB=75001.6 A=0.063 P=1.14 MULT=1
MM1039 N_VGND_M1039_d N_A_575_305#_M1039_g A_2565_74# VNB NLOWVT L=0.15 W=0.42
+ AD=0.165742 AS=0.0504 PD=1.19264 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75001.5
+ SB=75001.2 A=0.063 P=1.14 MULT=1
MM1035 N_A_575_305#_M1035_d N_A_2463_74#_M1035_g N_VGND_M1039_d VNB NLOWVT
+ L=0.15 W=0.64 AD=0.1824 AS=0.252558 PD=1.85 PS=1.81736 NRD=0 NRS=13.116 M=1
+ R=4.26667 SA=75001.7 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1042 N_VGND_M1042_d N_A_2463_74#_M1042_g N_Q_M1042_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1961 AS=0.2109 PD=1.27 PS=2.05 NRD=40.536 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75000.9 A=0.111 P=1.78 MULT=1
MM1004 N_Q_N_M1004_d N_A_575_305#_M1004_g N_VGND_M1042_d VNB NLOWVT L=0.15
+ W=0.74 AD=0.2109 AS=0.1961 PD=2.05 PS=1.27 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.9 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1021 A_116_464# N_D_M1021_g N_A_27_90#_M1021_s VPB PSHORT L=0.15 W=0.64
+ AD=0.0768 AS=0.1888 PD=0.88 PS=1.87 NRD=19.9955 NRS=3.0732 M=1 R=4.26667
+ SA=75000.2 SB=75000.6 A=0.096 P=1.58 MULT=1
MM1001 N_VPWR_M1001_d N_A_161_394#_M1001_g A_116_464# VPB PSHORT L=0.15 W=0.64
+ AD=0.1888 AS=0.0768 PD=1.87 PS=0.88 NRD=3.0732 NRS=19.9955 M=1 R=4.26667
+ SA=75000.6 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1034 N_VPWR_M1034_d N_DE_M1034_g N_A_161_394#_M1034_s VPB PSHORT L=0.15 W=0.64
+ AD=0.1696 AS=0.1888 PD=1.17 PS=1.87 NRD=73.8553 NRS=3.0732 M=1 R=4.26667
+ SA=75000.2 SB=75001.8 A=0.096 P=1.58 MULT=1
MM1037 A_556_464# N_DE_M1037_g N_VPWR_M1034_d VPB PSHORT L=0.15 W=0.64 AD=0.0864
+ AS=0.1696 PD=0.91 PS=1.17 NRD=24.625 NRS=3.0732 M=1 R=4.26667 SA=75000.9
+ SB=75001.1 A=0.096 P=1.58 MULT=1
MM1013 N_A_27_90#_M1013_d N_A_575_305#_M1013_g A_556_464# VPB PSHORT L=0.15
+ W=0.64 AD=0.096 AS=0.0864 PD=0.94 PS=0.91 NRD=3.0732 NRS=24.625 M=1 R=4.26667
+ SA=75001.3 SB=75000.7 A=0.096 P=1.58 MULT=1
MM1017 N_A_697_113#_M1017_d N_SCE_M1017_g N_A_27_90#_M1013_d VPB PSHORT L=0.15
+ W=0.64 AD=0.1888 AS=0.096 PD=1.87 PS=0.94 NRD=3.0732 NRS=3.0732 M=1 R=4.26667
+ SA=75001.8 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1006 N_VPWR_M1006_d N_SCE_M1006_g N_A_667_87#_M1006_s VPB PSHORT L=0.15 W=0.64
+ AD=0.1488 AS=0.2304 PD=1.105 PS=2 NRD=53.8598 NRS=23.0687 M=1 R=4.26667
+ SA=75000.3 SB=75001.2 A=0.096 P=1.58 MULT=1
MM1018 A_1068_462# N_SCD_M1018_g N_VPWR_M1006_d VPB PSHORT L=0.15 W=0.64
+ AD=0.0768 AS=0.1488 PD=0.88 PS=1.105 NRD=19.9955 NRS=3.0732 M=1 R=4.26667
+ SA=75000.9 SB=75000.6 A=0.096 P=1.58 MULT=1
MM1002 N_A_697_113#_M1002_d N_A_667_87#_M1002_g A_1068_462# VPB PSHORT L=0.15
+ W=0.64 AD=0.1888 AS=0.0768 PD=1.87 PS=0.88 NRD=3.0732 NRS=19.9955 M=1
+ R=4.26667 SA=75001.3 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1029 N_A_1348_368#_M1029_d N_CLK_M1029_g N_VPWR_M1029_s VPB PSHORT L=0.15
+ W=1.12 AD=0.3304 AS=0.3304 PD=2.83 PS=2.83 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75000.2 A=0.168 P=2.54 MULT=1
MM1010 N_A_1549_74#_M1010_d N_A_1348_368#_M1010_g N_VPWR_M1010_s VPB PSHORT
+ L=0.15 W=1.12 AD=0.3304 AS=0.3304 PD=2.83 PS=2.83 NRD=1.7533 NRS=1.7533 M=1
+ R=7.46667 SA=75000.2 SB=75000.2 A=0.168 P=2.54 MULT=1
MM1032 N_A_1747_118#_M1032_d N_A_1549_74#_M1032_g N_A_697_113#_M1032_s VPB
+ PSHORT L=0.15 W=0.42 AD=0.0735 AS=0.1302 PD=0.77 PS=1.46 NRD=28.1316
+ NRS=9.3772 M=1 R=2.8 SA=75000.2 SB=75001.5 A=0.063 P=1.14 MULT=1
MM1030 A_1931_508# N_A_1348_368#_M1030_g N_A_1747_118#_M1032_d VPB PSHORT L=0.15
+ W=0.42 AD=0.0588 AS=0.0735 PD=0.7 PS=0.77 NRD=39.8531 NRS=4.6886 M=1 R=2.8
+ SA=75000.7 SB=75001 A=0.063 P=1.14 MULT=1
MM1020 N_VPWR_M1020_d N_A_1972_92#_M1020_g A_1931_508# VPB PSHORT L=0.15 W=0.42
+ AD=0.0999833 AS=0.0588 PD=0.91 PS=0.7 NRD=9.3772 NRS=39.8531 M=1 R=2.8
+ SA=75001.2 SB=75000.6 A=0.063 P=1.14 MULT=1
MM1007 N_A_1972_92#_M1007_d N_A_1747_118#_M1007_g N_VPWR_M1020_d VPB PSHORT
+ L=0.15 W=0.84 AD=0.2478 AS=0.199967 PD=2.27 PS=1.82 NRD=2.3443 NRS=23.443 M=1
+ R=5.6 SA=75000.7 SB=75000.2 A=0.126 P=1.98 MULT=1
MM1009 A_2345_392# N_A_1972_92#_M1009_g N_VPWR_M1009_s VPB PSHORT L=0.15 W=1
+ AD=0.4125 AS=0.4032 PD=1.825 PS=2.92 NRD=70.4078 NRS=19.6803 M=1 R=6.66667
+ SA=75000.3 SB=75001.9 A=0.15 P=2.3 MULT=1
MM1019 N_A_2463_74#_M1019_d N_A_1348_368#_M1019_g A_2345_392# VPB PSHORT L=0.15
+ W=1 AD=0.234366 AS=0.4125 PD=1.9507 PS=1.825 NRD=1.9503 NRS=70.4078 M=1
+ R=6.66667 SA=75001.3 SB=75000.9 A=0.15 P=2.3 MULT=1
MM1015 A_2647_508# N_A_1549_74#_M1015_g N_A_2463_74#_M1019_d VPB PSHORT L=0.15
+ W=0.42 AD=0.0567 AS=0.0984338 PD=0.69 PS=0.819296 NRD=37.5088 NRS=44.5417 M=1
+ R=2.8 SA=75001.8 SB=75001.3 A=0.063 P=1.14 MULT=1
MM1040 N_VPWR_M1040_d N_A_575_305#_M1040_g A_2647_508# VPB PSHORT L=0.15 W=0.42
+ AD=0.115027 AS=0.0567 PD=0.922817 PS=0.69 NRD=65.6601 NRS=37.5088 M=1 R=2.8
+ SA=75002.2 SB=75000.9 A=0.063 P=1.14 MULT=1
MM1016 N_A_575_305#_M1016_d N_A_2463_74#_M1016_g N_VPWR_M1040_d VPB PSHORT
+ L=0.15 W=1 AD=0.295 AS=0.273873 PD=2.59 PS=2.19718 NRD=1.9503 NRS=27.5603 M=1
+ R=6.66667 SA=75001.3 SB=75000.2 A=0.15 P=2.3 MULT=1
MM1027 N_VPWR_M1027_d N_A_2463_74#_M1027_g N_Q_M1027_s VPB PSHORT L=0.15 W=1.12
+ AD=0.196 AS=0.3304 PD=1.47 PS=2.83 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1024 N_Q_N_M1024_d N_A_575_305#_M1024_g N_VPWR_M1027_d VPB PSHORT L=0.15
+ W=1.12 AD=0.3304 AS=0.196 PD=2.83 PS=1.47 NRD=1.7533 NRS=10.5395 M=1 R=7.46667
+ SA=75000.7 SB=75000.2 A=0.168 P=2.54 MULT=1
DX44_noxref VNB VPB NWDIODE A=31.062 P=37.12
c_173 VNB 0 1.45871e-19 $X=0 $Y=0
c_336 VPB 0 1.97671e-19 $X=0 $Y=3.085
*
.include "sky130_fd_sc_hs__sedfxbp_1.pxi.spice"
*
.ends
*
*
