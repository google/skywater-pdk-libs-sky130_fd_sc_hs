* File: sky130_fd_sc_hs__dlxtn_2.pex.spice
* Created: Tue Sep  1 20:03:03 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HS__DLXTN_2%D 3 6 7 9 10 14 17
c32 3 0 1.87332e-19 $X=0.495 $Y=0.875
r33 16 17 27.9778 $w=3.3e-07 $l=1.6e-07 $layer=POLY_cond $X=0.495 $Y=1.465
+ $X2=0.655 $Y2=1.465
r34 13 16 35.8466 $w=3.3e-07 $l=2.05e-07 $layer=POLY_cond $X=0.29 $Y=1.465
+ $X2=0.495 $Y2=1.465
r35 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.29
+ $Y=1.465 $X2=0.29 $Y2=1.465
r36 10 14 6.9845 $w=3.28e-07 $l=2e-07 $layer=LI1_cond $X=0.29 $Y=1.665 $X2=0.29
+ $Y2=1.465
r37 7 9 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=0.655 $Y=2.045
+ $X2=0.655 $Y2=2.54
r38 6 7 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=0.655 $Y=1.955 $X2=0.655
+ $Y2=2.045
r39 5 17 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=0.655 $Y=1.63
+ $X2=0.655 $Y2=1.465
r40 5 6 126.331 $w=1.8e-07 $l=3.25e-07 $layer=POLY_cond $X=0.655 $Y=1.63
+ $X2=0.655 $Y2=1.955
r41 1 16 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.495 $Y=1.3
+ $X2=0.495 $Y2=1.465
r42 1 3 217.926 $w=1.5e-07 $l=4.25e-07 $layer=POLY_cond $X=0.495 $Y=1.3
+ $X2=0.495 $Y2=0.875
.ends

.subckt PM_SKY130_FD_SC_HS__DLXTN_2%GATE_N 3 6 7 9 10 13
c48 13 0 1.38982e-19 $X=1.15 $Y=1.615
r49 13 16 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.15 $Y=1.615
+ $X2=1.15 $Y2=1.78
r50 13 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.15 $Y=1.615
+ $X2=1.15 $Y2=1.45
r51 10 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.15
+ $Y=1.615 $X2=1.15 $Y2=1.615
r52 7 9 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=1.205 $Y=2.045
+ $X2=1.205 $Y2=2.54
r53 6 7 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=1.205 $Y=1.955 $X2=1.205
+ $Y2=2.045
r54 6 16 68.0242 $w=1.8e-07 $l=1.75e-07 $layer=POLY_cond $X=1.205 $Y=1.955
+ $X2=1.205 $Y2=1.78
r55 3 15 343.553 $w=1.5e-07 $l=6.7e-07 $layer=POLY_cond $X=1.085 $Y=0.78
+ $X2=1.085 $Y2=1.45
.ends

.subckt PM_SKY130_FD_SC_HS__DLXTN_2%A_232_82# 1 2 7 10 11 13 14 16 17 19 21 23
+ 24 26 29 31 35 37 41 42 45 48 49 50 52 54 55 60 62 63 66 67
c168 67 0 4.79549e-20 $X=4.185 $Y=1.65
c169 66 0 1.38828e-19 $X=4.185 $Y=1.65
c170 54 0 1.38982e-19 $X=1.43 $Y=2.265
c171 37 0 1.87332e-19 $X=1.485 $Y=1.045
c172 24 0 1.93308e-19 $X=3.88 $Y=2.44
c173 11 0 6.74217e-20 $X=2.215 $Y=1.885
r174 74 76 9.61737 $w=3.3e-07 $l=5.5e-08 $layer=POLY_cond $X=3.825 $Y=1.65
+ $X2=3.88 $Y2=1.65
r175 67 76 53.3327 $w=3.3e-07 $l=3.05e-07 $layer=POLY_cond $X=4.185 $Y=1.65
+ $X2=3.88 $Y2=1.65
r176 66 69 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=4.185 $Y=1.65
+ $X2=4.185 $Y2=1.815
r177 66 67 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.185
+ $Y=1.65 $X2=4.185 $Y2=1.65
r178 62 64 8.64761 $w=3.98e-07 $l=1.65e-07 $layer=LI1_cond $X=1.685 $Y=1.605
+ $X2=1.685 $Y2=1.77
r179 62 63 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.72
+ $Y=1.605 $X2=1.72 $Y2=1.605
r180 59 60 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.72
+ $Y=0.925 $X2=1.72 $Y2=0.925
r181 55 64 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=1.57 $Y=2.1
+ $X2=1.57 $Y2=1.77
r182 54 56 7.68295 $w=3.88e-07 $l=2.6e-07 $layer=LI1_cond $X=1.46 $Y=2.265
+ $X2=1.46 $Y2=2.525
r183 54 55 8.60763 $w=3.88e-07 $l=1.65e-07 $layer=LI1_cond $X=1.46 $Y=2.265
+ $X2=1.46 $Y2=2.1
r184 52 69 71.1123 $w=1.68e-07 $l=1.09e-06 $layer=LI1_cond $X=4.105 $Y=2.905
+ $X2=4.105 $Y2=1.815
r185 49 52 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.02 $Y=2.99
+ $X2=4.105 $Y2=2.905
r186 49 50 63.6096 $w=1.68e-07 $l=9.75e-07 $layer=LI1_cond $X=4.02 $Y=2.99
+ $X2=3.045 $Y2=2.99
r187 48 50 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.96 $Y=2.905
+ $X2=3.045 $Y2=2.99
r188 47 48 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=2.96 $Y=2.61
+ $X2=2.96 $Y2=2.905
r189 46 56 5.6248 $w=1.7e-07 $l=1.95e-07 $layer=LI1_cond $X=1.655 $Y=2.525
+ $X2=1.46 $Y2=2.525
r190 45 47 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.875 $Y=2.525
+ $X2=2.96 $Y2=2.61
r191 45 46 79.5936 $w=1.68e-07 $l=1.22e-06 $layer=LI1_cond $X=2.875 $Y=2.525
+ $X2=1.655 $Y2=2.525
r192 42 62 1.00839 $w=3.98e-07 $l=3.5e-08 $layer=LI1_cond $X=1.685 $Y=1.57
+ $X2=1.685 $Y2=1.605
r193 41 59 3.08538 $w=4e-07 $l=2.05e-07 $layer=LI1_cond $X=1.685 $Y=1.17
+ $X2=1.685 $Y2=0.965
r194 41 42 11.5244 $w=3.98e-07 $l=4e-07 $layer=LI1_cond $X=1.685 $Y=1.17
+ $X2=1.685 $Y2=1.57
r195 37 59 4.21417 $w=2.5e-07 $l=2.36643e-07 $layer=LI1_cond $X=1.485 $Y=1.045
+ $X2=1.685 $Y2=0.965
r196 37 39 8.52808 $w=2.48e-07 $l=1.85e-07 $layer=LI1_cond $X=1.485 $Y=1.045
+ $X2=1.3 $Y2=1.045
r197 33 35 112.809 $w=1.5e-07 $l=2.2e-07 $layer=POLY_cond $X=3.605 $Y=1.185
+ $X2=3.825 $Y2=1.185
r198 28 63 47.2125 $w=3.3e-07 $l=2.7e-07 $layer=POLY_cond $X=1.72 $Y=1.335
+ $X2=1.72 $Y2=1.605
r199 28 29 10.1687 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=1.72 $Y=1.335
+ $X2=1.72 $Y2=1.26
r200 27 60 45.4639 $w=3.3e-07 $l=2.6e-07 $layer=POLY_cond $X=1.72 $Y=1.185
+ $X2=1.72 $Y2=0.925
r201 27 29 10.1687 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=1.72 $Y=1.185
+ $X2=1.72 $Y2=1.26
r202 24 26 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=3.88 $Y=2.44
+ $X2=3.88 $Y2=2.725
r203 23 24 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=3.88 $Y=2.35 $X2=3.88
+ $Y2=2.44
r204 22 76 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=3.88 $Y=1.815
+ $X2=3.88 $Y2=1.65
r205 22 23 207.96 $w=1.8e-07 $l=5.35e-07 $layer=POLY_cond $X=3.88 $Y=1.815
+ $X2=3.88 $Y2=2.35
r206 21 74 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.825 $Y=1.485
+ $X2=3.825 $Y2=1.65
r207 20 35 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.825 $Y=1.26
+ $X2=3.825 $Y2=1.185
r208 20 21 115.372 $w=1.5e-07 $l=2.25e-07 $layer=POLY_cond $X=3.825 $Y=1.26
+ $X2=3.825 $Y2=1.485
r209 17 33 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.605 $Y=1.11
+ $X2=3.605 $Y2=1.185
r210 17 19 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=3.605 $Y=1.11
+ $X2=3.605 $Y2=0.715
r211 14 31 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.355 $Y=1.185
+ $X2=2.355 $Y2=1.26
r212 14 16 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=2.355 $Y=1.185
+ $X2=2.355 $Y2=0.74
r213 11 13 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=2.215 $Y=1.885
+ $X2=2.215 $Y2=2.38
r214 10 11 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=2.215 $Y=1.795
+ $X2=2.215 $Y2=1.885
r215 9 31 71.7872 $w=1.5e-07 $l=1.4e-07 $layer=POLY_cond $X=2.215 $Y=1.26
+ $X2=2.355 $Y2=1.26
r216 9 10 178.806 $w=1.8e-07 $l=4.6e-07 $layer=POLY_cond $X=2.215 $Y=1.335
+ $X2=2.215 $Y2=1.795
r217 8 29 16.9349 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.885 $Y=1.26
+ $X2=1.72 $Y2=1.26
r218 7 9 46.1489 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=2.125 $Y=1.26 $X2=2.215
+ $Y2=1.26
r219 7 8 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=2.125 $Y=1.26
+ $X2=1.885 $Y2=1.26
r220 2 54 300 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=2 $X=1.28
+ $Y=2.12 $X2=1.43 $Y2=2.265
r221 1 39 182 $w=1.7e-07 $l=6.61306e-07 $layer=licon1_NDIFF $count=1 $X=1.16
+ $Y=0.41 $X2=1.3 $Y2=1.005
.ends

.subckt PM_SKY130_FD_SC_HS__DLXTN_2%A_27_120# 1 2 7 8 9 11 12 14 16 19 22 23 26
+ 27 28 30 35 38 43
c120 9 0 1.12757e-19 $X=2.85 $Y=1.885
r121 43 44 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.805
+ $Y=1.465 $X2=2.805 $Y2=1.465
r122 40 43 8.55602 $w=3.28e-07 $l=2.45e-07 $layer=LI1_cond $X=2.56 $Y=1.465
+ $X2=2.805 $Y2=1.465
r123 34 35 8.09223 $w=5.48e-07 $l=8.5e-08 $layer=LI1_cond $X=0.71 $Y=0.855
+ $X2=0.795 $Y2=0.855
r124 32 34 9.35116 $w=5.48e-07 $l=4.3e-07 $layer=LI1_cond $X=0.28 $Y=0.855
+ $X2=0.71 $Y2=0.855
r125 30 40 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.56 $Y=1.3
+ $X2=2.56 $Y2=1.465
r126 29 30 57.0856 $w=1.68e-07 $l=8.75e-07 $layer=LI1_cond $X=2.56 $Y=0.425
+ $X2=2.56 $Y2=1.3
r127 27 29 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.475 $Y=0.34
+ $X2=2.56 $Y2=0.425
r128 27 28 75.6791 $w=1.68e-07 $l=1.16e-06 $layer=LI1_cond $X=2.475 $Y=0.34
+ $X2=1.315 $Y2=0.34
r129 25 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.23 $Y=0.425
+ $X2=1.315 $Y2=0.34
r130 25 26 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=1.23 $Y=0.425
+ $X2=1.23 $Y2=0.58
r131 23 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.145 $Y=0.665
+ $X2=1.23 $Y2=0.58
r132 23 35 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=1.145 $Y=0.665
+ $X2=0.795 $Y2=0.665
r133 22 38 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.71 $Y=1.95
+ $X2=0.71 $Y2=2.035
r134 21 34 7.75927 $w=1.7e-07 $l=2.75e-07 $layer=LI1_cond $X=0.71 $Y=1.13
+ $X2=0.71 $Y2=0.855
r135 21 22 53.4973 $w=1.68e-07 $l=8.2e-07 $layer=LI1_cond $X=0.71 $Y=1.13
+ $X2=0.71 $Y2=1.95
r136 17 38 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=0.43 $Y=2.035
+ $X2=0.71 $Y2=2.035
r137 17 19 5.06376 $w=3.28e-07 $l=1.45e-07 $layer=LI1_cond $X=0.43 $Y=2.12
+ $X2=0.43 $Y2=2.265
r138 14 16 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=3.215 $Y=1.11
+ $X2=3.215 $Y2=0.715
r139 13 44 48.5468 $w=2.78e-07 $l=3.52987e-07 $layer=POLY_cond $X=2.97 $Y=1.185
+ $X2=2.805 $Y2=1.465
r140 12 14 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.14 $Y=1.185
+ $X2=3.215 $Y2=1.11
r141 12 13 87.1702 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=3.14 $Y=1.185
+ $X2=2.97 $Y2=1.185
r142 9 11 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=2.85 $Y=1.885
+ $X2=2.85 $Y2=2.46
r143 8 9 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=2.85 $Y=1.795 $X2=2.85
+ $Y2=1.885
r144 7 44 34.5863 $w=2.78e-07 $l=1.86145e-07 $layer=POLY_cond $X=2.85 $Y=1.63
+ $X2=2.805 $Y2=1.465
r145 7 8 64.1371 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=2.85 $Y=1.63
+ $X2=2.85 $Y2=1.795
r146 2 19 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=0.285
+ $Y=2.12 $X2=0.43 $Y2=2.265
r147 1 32 182 $w=1.7e-07 $l=3.19374e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.6 $X2=0.28 $Y2=0.855
.ends

.subckt PM_SKY130_FD_SC_HS__DLXTN_2%A_369_392# 1 2 7 9 12 15 17 18 21 23 24 30
+ 32 38
c104 38 0 1.38828e-19 $X=4.21 $Y=0.585
c105 30 0 1.60712e-19 $X=3.345 $Y=1.635
c106 23 0 6.89381e-20 $X=4.21 $Y=0.42
c107 21 0 3.15497e-20 $X=3.485 $Y=0.42
c108 15 0 6.74217e-20 $X=2.14 $Y=0.86
r109 30 33 8.73063 $w=3.28e-07 $l=2.5e-07 $layer=LI1_cond $X=3.345 $Y=1.635
+ $X2=3.345 $Y2=1.885
r110 30 32 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=3.345 $Y=1.635
+ $X2=3.345 $Y2=1.47
r111 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.345
+ $Y=1.635 $X2=3.345 $Y2=1.635
r112 27 28 6.58523 $w=3.52e-07 $l=1.9e-07 $layer=LI1_cond $X=1.99 $Y=2.035
+ $X2=2.18 $Y2=2.035
r113 24 38 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.21 $Y=0.42
+ $X2=4.21 $Y2=0.585
r114 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.21
+ $Y=0.42 $X2=4.21 $Y2=0.42
r115 21 23 25.3188 $w=3.28e-07 $l=7.25e-07 $layer=LI1_cond $X=3.485 $Y=0.42
+ $X2=4.21 $Y2=0.42
r116 19 21 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.4 $Y=0.585
+ $X2=3.485 $Y2=0.42
r117 19 32 57.738 $w=1.68e-07 $l=8.85e-07 $layer=LI1_cond $X=3.4 $Y=0.585
+ $X2=3.4 $Y2=1.47
r118 18 28 7.60401 $w=3.52e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.305 $Y=1.885
+ $X2=2.18 $Y2=2.035
r119 17 33 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.18 $Y=1.885
+ $X2=3.345 $Y2=1.885
r120 17 18 57.0856 $w=1.68e-07 $l=8.75e-07 $layer=LI1_cond $X=3.18 $Y=1.885
+ $X2=2.305 $Y2=1.885
r121 13 28 2.74175 $w=2.5e-07 $l=2.35e-07 $layer=LI1_cond $X=2.18 $Y=1.8
+ $X2=2.18 $Y2=2.035
r122 13 15 43.3319 $w=2.48e-07 $l=9.4e-07 $layer=LI1_cond $X=2.18 $Y=1.8
+ $X2=2.18 $Y2=0.86
r123 12 38 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=4.3 $Y=0.905
+ $X2=4.3 $Y2=0.585
r124 7 31 52.2586 $w=2.99e-07 $l=2.85044e-07 $layer=POLY_cond $X=3.27 $Y=1.885
+ $X2=3.345 $Y2=1.635
r125 7 9 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=3.27 $Y=1.885
+ $X2=3.27 $Y2=2.46
r126 2 27 600 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=1.845
+ $Y=1.96 $X2=1.99 $Y2=2.105
r127 1 15 182 $w=1.7e-07 $l=5.57808e-07 $layer=licon1_NDIFF $count=1 $X=1.995
+ $Y=0.37 $X2=2.14 $Y2=0.86
.ends

.subckt PM_SKY130_FD_SC_HS__DLXTN_2%A_842_405# 1 2 7 9 12 16 18 20 23 25 27 28
+ 31 33 36 38 40 44 47 49 52 59 60
c98 49 0 1.98766e-19 $X=5.59 $Y=1.795
c99 12 0 6.89381e-20 $X=4.69 $Y=0.905
r100 58 59 9.02376 $w=2.48e-07 $l=1.7e-07 $layer=LI1_cond $X=5.502 $Y=0.955
+ $X2=5.502 $Y2=1.125
r101 56 57 7.83799 $w=3.58e-07 $l=2.3e-07 $layer=LI1_cond $X=5.462 $Y=1.96
+ $X2=5.462 $Y2=2.19
r102 52 53 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.08
+ $Y=1.46 $X2=6.08 $Y2=1.46
r103 50 60 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.675 $Y=1.46
+ $X2=5.59 $Y2=1.46
r104 50 52 14.1436 $w=3.28e-07 $l=4.05e-07 $layer=LI1_cond $X=5.675 $Y=1.46
+ $X2=6.08 $Y2=1.46
r105 49 56 9.00471 $w=3.58e-07 $l=2.19875e-07 $layer=LI1_cond $X=5.59 $Y=1.795
+ $X2=5.462 $Y2=1.96
r106 48 60 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.59 $Y=1.625
+ $X2=5.59 $Y2=1.46
r107 48 49 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=5.59 $Y=1.625
+ $X2=5.59 $Y2=1.795
r108 47 60 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.59 $Y=1.295
+ $X2=5.59 $Y2=1.46
r109 47 59 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=5.59 $Y=1.295
+ $X2=5.59 $Y2=1.125
r110 44 58 20.0525 $w=2.48e-07 $l=4.35e-07 $layer=LI1_cond $X=5.455 $Y=0.52
+ $X2=5.455 $Y2=0.955
r111 38 57 5.71829 $w=3.58e-07 $l=1.87029e-07 $layer=LI1_cond $X=5.415 $Y=2.355
+ $X2=5.462 $Y2=2.19
r112 38 40 15.1913 $w=3.28e-07 $l=4.35e-07 $layer=LI1_cond $X=5.415 $Y=2.355
+ $X2=5.415 $Y2=2.79
r113 36 65 22.2773 $w=3.57e-07 $l=1.65e-07 $layer=POLY_cond $X=4.525 $Y=2.232
+ $X2=4.69 $Y2=2.232
r114 36 63 30.3782 $w=3.57e-07 $l=2.25e-07 $layer=POLY_cond $X=4.525 $Y=2.232
+ $X2=4.3 $Y2=2.232
r115 35 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.525
+ $Y=2.19 $X2=4.525 $Y2=2.19
r116 33 57 1.20828 $w=3.3e-07 $l=2.12e-07 $layer=LI1_cond $X=5.25 $Y=2.19
+ $X2=5.462 $Y2=2.19
r117 33 35 25.3188 $w=3.28e-07 $l=7.25e-07 $layer=LI1_cond $X=5.25 $Y=2.19
+ $X2=4.525 $Y2=2.19
r118 31 32 1.81658 $w=3.98e-07 $l=1.5e-08 $layer=POLY_cond $X=6.68 $Y=1.53
+ $X2=6.695 $Y2=1.53
r119 30 31 58.1307 $w=3.98e-07 $l=4.8e-07 $layer=POLY_cond $X=6.2 $Y=1.53
+ $X2=6.68 $Y2=1.53
r120 29 30 1.21106 $w=3.98e-07 $l=1e-08 $layer=POLY_cond $X=6.19 $Y=1.53 $X2=6.2
+ $Y2=1.53
r121 28 53 5.24584 $w=3.3e-07 $l=3e-08 $layer=POLY_cond $X=6.11 $Y=1.46 $X2=6.08
+ $Y2=1.46
r122 28 29 11.2379 $w=3.98e-07 $l=1.09545e-07 $layer=POLY_cond $X=6.11 $Y=1.46
+ $X2=6.19 $Y2=1.53
r123 25 32 25.7394 $w=1.5e-07 $l=2.35e-07 $layer=POLY_cond $X=6.695 $Y=1.765
+ $X2=6.695 $Y2=1.53
r124 25 27 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=6.695 $Y=1.765
+ $X2=6.695 $Y2=2.4
r125 21 31 25.7394 $w=1.5e-07 $l=2.35e-07 $layer=POLY_cond $X=6.68 $Y=1.295
+ $X2=6.68 $Y2=1.53
r126 21 23 284.585 $w=1.5e-07 $l=5.55e-07 $layer=POLY_cond $X=6.68 $Y=1.295
+ $X2=6.68 $Y2=0.74
r127 18 30 25.7394 $w=1.5e-07 $l=2.35e-07 $layer=POLY_cond $X=6.2 $Y=1.765
+ $X2=6.2 $Y2=1.53
r128 18 20 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=6.2 $Y=1.765
+ $X2=6.2 $Y2=2.4
r129 14 29 25.7394 $w=1.5e-07 $l=2.35e-07 $layer=POLY_cond $X=6.19 $Y=1.295
+ $X2=6.19 $Y2=1.53
r130 14 16 284.585 $w=1.5e-07 $l=5.55e-07 $layer=POLY_cond $X=6.19 $Y=1.295
+ $X2=6.19 $Y2=0.74
r131 10 65 23.1043 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.69 $Y=2.025
+ $X2=4.69 $Y2=2.232
r132 10 12 574.298 $w=1.5e-07 $l=1.12e-06 $layer=POLY_cond $X=4.69 $Y=2.025
+ $X2=4.69 $Y2=0.905
r133 7 63 23.1043 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=4.3 $Y=2.44 $X2=4.3
+ $Y2=2.232
r134 7 9 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=4.3 $Y=2.44 $X2=4.3
+ $Y2=2.725
r135 2 56 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=5.265
+ $Y=1.815 $X2=5.415 $Y2=1.96
r136 2 40 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=5.265
+ $Y=1.815 $X2=5.415 $Y2=2.79
r137 1 44 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=5.275
+ $Y=0.375 $X2=5.415 $Y2=0.52
.ends

.subckt PM_SKY130_FD_SC_HS__DLXTN_2%A_669_392# 1 2 7 9 12 16 17 19 20
r68 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.17
+ $Y=1.46 $X2=5.17 $Y2=1.46
r69 19 20 7.80118 $w=5.18e-07 $l=8.5e-08 $layer=LI1_cond $X=3.59 $Y=2.225
+ $X2=3.59 $Y2=2.14
r70 17 24 14.0393 $w=3.24e-07 $l=3.77492e-07 $layer=LI1_cond $X=4.25 $Y=1.23
+ $X2=3.95 $Y2=1.055
r71 16 27 9.67586 $w=2.9e-07 $l=3.04072e-07 $layer=LI1_cond $X=4.99 $Y=1.23
+ $X2=5.162 $Y2=1.46
r72 16 17 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=4.99 $Y=1.23
+ $X2=4.25 $Y2=1.23
r73 14 24 6.96605 $w=3.24e-07 $l=1.85e-07 $layer=LI1_cond $X=3.765 $Y=1.055
+ $X2=3.95 $Y2=1.055
r74 14 20 70.7861 $w=1.68e-07 $l=1.085e-06 $layer=LI1_cond $X=3.765 $Y=1.055
+ $X2=3.765 $Y2=2.14
r75 10 28 38.6072 $w=2.91e-07 $l=1.79374e-07 $layer=POLY_cond $X=5.2 $Y=1.295
+ $X2=5.17 $Y2=1.46
r76 10 12 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=5.2 $Y=1.295 $X2=5.2
+ $Y2=0.745
r77 7 28 57.6553 $w=2.91e-07 $l=2.89828e-07 $layer=POLY_cond $X=5.19 $Y=1.74
+ $X2=5.17 $Y2=1.46
r78 7 9 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=5.19 $Y=1.74 $X2=5.19
+ $Y2=2.375
r79 2 19 300 $w=1.7e-07 $l=3.45326e-07 $layer=licon1_PDIFF $count=2 $X=3.345
+ $Y=1.96 $X2=3.53 $Y2=2.225
r80 1 24 182 $w=1.7e-07 $l=6.15366e-07 $layer=licon1_NDIFF $count=1 $X=3.68
+ $Y=0.395 $X2=3.95 $Y2=0.89
.ends

.subckt PM_SKY130_FD_SC_HS__DLXTN_2%VPWR 1 2 3 4 5 18 22 26 30 32 37 38 40 41 42
+ 48 64 69 74 77 80
c82 77 0 1.93308e-19 $X=5.08 $Y=3.02
r83 79 80 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r84 76 77 10.6911 $w=7.88e-07 $l=1.2e-07 $layer=LI1_cond $X=4.96 $Y=3.02
+ $X2=5.08 $Y2=3.02
r85 72 76 6.05609 $w=7.88e-07 $l=4e-07 $layer=LI1_cond $X=4.56 $Y=3.02 $X2=4.96
+ $Y2=3.02
r86 72 74 11.9023 $w=7.88e-07 $l=2e-07 $layer=LI1_cond $X=4.56 $Y=3.02 $X2=4.36
+ $Y2=3.02
r87 72 73 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r88 69 70 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r89 67 80 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=6.96 $Y2=3.33
r90 66 67 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r91 64 79 4.01252 $w=1.7e-07 $l=1.82e-07 $layer=LI1_cond $X=6.835 $Y=3.33
+ $X2=7.017 $Y2=3.33
r92 64 66 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=6.835 $Y=3.33
+ $X2=6.48 $Y2=3.33
r93 63 67 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=6.48 $Y2=3.33
r94 63 73 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=4.56 $Y2=3.33
r95 62 77 28.7059 $w=1.68e-07 $l=4.4e-07 $layer=LI1_cond $X=5.52 $Y=3.33
+ $X2=5.08 $Y2=3.33
r96 62 63 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r97 59 73 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=4.56 $Y2=3.33
r98 58 74 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=4.08 $Y=3.33
+ $X2=4.36 $Y2=3.33
r99 58 59 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r100 56 69 8.88104 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=2.705 $Y=3.33
+ $X2=2.532 $Y2=3.33
r101 56 58 89.7059 $w=1.68e-07 $l=1.375e-06 $layer=LI1_cond $X=2.705 $Y=3.33
+ $X2=4.08 $Y2=3.33
r102 54 70 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r103 53 54 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r104 51 54 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.16 $Y2=3.33
r105 50 53 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.2 $Y=3.33 $X2=2.16
+ $Y2=3.33
r106 50 51 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r107 48 69 8.88104 $w=1.7e-07 $l=1.72e-07 $layer=LI1_cond $X=2.36 $Y=3.33
+ $X2=2.532 $Y2=3.33
r108 48 53 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=2.36 $Y=3.33 $X2=2.16
+ $Y2=3.33
r109 46 51 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r110 45 46 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r111 42 59 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.08 $Y2=3.33
r112 42 70 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=2.64 $Y2=3.33
r113 40 62 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=5.845 $Y=3.33
+ $X2=5.52 $Y2=3.33
r114 40 41 6.25164 $w=1.7e-07 $l=1.07e-07 $layer=LI1_cond $X=5.845 $Y=3.33
+ $X2=5.952 $Y2=3.33
r115 39 66 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=6.06 $Y=3.33
+ $X2=6.48 $Y2=3.33
r116 39 41 6.25164 $w=1.7e-07 $l=1.08e-07 $layer=LI1_cond $X=6.06 $Y=3.33
+ $X2=5.952 $Y2=3.33
r117 37 45 2.93583 $w=1.68e-07 $l=4.5e-08 $layer=LI1_cond $X=0.765 $Y=3.33
+ $X2=0.72 $Y2=3.33
r118 37 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.765 $Y=3.33
+ $X2=0.93 $Y2=3.33
r119 36 50 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=1.095 $Y=3.33
+ $X2=1.2 $Y2=3.33
r120 36 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.095 $Y=3.33
+ $X2=0.93 $Y2=3.33
r121 32 35 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=6.96 $Y=1.985
+ $X2=6.96 $Y2=2.815
r122 30 79 3.13065 $w=2.5e-07 $l=1.09864e-07 $layer=LI1_cond $X=6.96 $Y=3.245
+ $X2=7.017 $Y2=3.33
r123 30 35 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=6.96 $Y=3.245
+ $X2=6.96 $Y2=2.815
r124 26 29 44.4897 $w=2.13e-07 $l=8.3e-07 $layer=LI1_cond $X=5.952 $Y=1.985
+ $X2=5.952 $Y2=2.815
r125 24 41 0.512231 $w=2.15e-07 $l=8.5e-08 $layer=LI1_cond $X=5.952 $Y=3.245
+ $X2=5.952 $Y2=3.33
r126 24 29 23.0489 $w=2.13e-07 $l=4.3e-07 $layer=LI1_cond $X=5.952 $Y=3.245
+ $X2=5.952 $Y2=2.815
r127 20 69 1.03204 $w=3.45e-07 $l=8.5e-08 $layer=LI1_cond $X=2.532 $Y=3.245
+ $X2=2.532 $Y2=3.33
r128 20 22 10.0212 $w=3.43e-07 $l=3e-07 $layer=LI1_cond $X=2.532 $Y=3.245
+ $X2=2.532 $Y2=2.945
r129 16 38 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.93 $Y=3.245
+ $X2=0.93 $Y2=3.33
r130 16 18 29.6841 $w=3.28e-07 $l=8.5e-07 $layer=LI1_cond $X=0.93 $Y=3.245
+ $X2=0.93 $Y2=2.395
r131 5 35 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=6.77
+ $Y=1.84 $X2=6.92 $Y2=2.815
r132 5 32 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=6.77
+ $Y=1.84 $X2=6.92 $Y2=1.985
r133 4 29 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=5.83
+ $Y=1.84 $X2=5.975 $Y2=2.815
r134 4 26 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=5.83
+ $Y=1.84 $X2=5.975 $Y2=1.985
r135 3 76 300 $w=1.7e-07 $l=7.09295e-07 $layer=licon1_PDIFF $count=2 $X=4.375
+ $Y=2.515 $X2=4.96 $Y2=2.79
r136 2 22 600 $w=1.7e-07 $l=1.09846e-06 $layer=licon1_PDIFF $count=1 $X=2.29
+ $Y=1.96 $X2=2.53 $Y2=2.945
r137 1 18 300 $w=1.7e-07 $l=3.61421e-07 $layer=licon1_PDIFF $count=2 $X=0.73
+ $Y=2.12 $X2=0.93 $Y2=2.395
.ends

.subckt PM_SKY130_FD_SC_HS__DLXTN_2%Q 1 2 9 13 14 15 16 29 31
r25 21 31 2.21269 $w=3.73e-07 $l=7.2e-08 $layer=LI1_cond $X=6.447 $Y=2.107
+ $X2=6.447 $Y2=2.035
r26 15 16 11.3708 $w=3.73e-07 $l=3.7e-07 $layer=LI1_cond $X=6.447 $Y=2.405
+ $X2=6.447 $Y2=2.775
r27 14 31 0.215123 $w=3.73e-07 $l=7e-09 $layer=LI1_cond $X=6.447 $Y=2.028
+ $X2=6.447 $Y2=2.035
r28 14 29 6.80275 $w=3.73e-07 $l=1.08e-07 $layer=LI1_cond $X=6.447 $Y=2.028
+ $X2=6.447 $Y2=1.92
r29 14 15 8.97369 $w=3.73e-07 $l=2.92e-07 $layer=LI1_cond $X=6.447 $Y=2.113
+ $X2=6.447 $Y2=2.405
r30 14 21 0.184391 $w=3.73e-07 $l=6e-09 $layer=LI1_cond $X=6.447 $Y=2.113
+ $X2=6.447 $Y2=2.107
r31 13 29 51.8663 $w=1.68e-07 $l=7.95e-07 $layer=LI1_cond $X=6.5 $Y=1.125
+ $X2=6.5 $Y2=1.92
r32 7 13 7.21712 $w=2.63e-07 $l=1.32e-07 $layer=LI1_cond $X=6.452 $Y=0.993
+ $X2=6.452 $Y2=1.125
r33 7 9 20.7875 $w=2.63e-07 $l=4.78e-07 $layer=LI1_cond $X=6.452 $Y=0.993
+ $X2=6.452 $Y2=0.515
r34 2 31 600 $w=1.7e-07 $l=3.18865e-07 $layer=licon1_PDIFF $count=1 $X=6.275
+ $Y=1.84 $X2=6.445 $Y2=2.085
r35 1 9 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=6.265
+ $Y=0.37 $X2=6.41 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__DLXTN_2%VGND 1 2 3 4 5 18 22 28 30 32 34 36 41 49 54
+ 59 66 72 75 78 82
r85 81 82 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=0 $X2=6.96
+ $Y2=0
r86 78 79 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=0 $X2=6 $Y2=0
r87 75 76 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r88 72 73 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r89 66 69 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=0.79 $Y=0 $X2=0.79
+ $Y2=0.325
r90 66 67 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r91 63 82 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=0 $X2=6.96
+ $Y2=0
r92 63 79 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=0 $X2=6
+ $Y2=0
r93 62 63 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=0 $X2=6.48
+ $Y2=0
r94 60 78 7.94884 $w=1.7e-07 $l=1.48e-07 $layer=LI1_cond $X=6.14 $Y=0 $X2=5.992
+ $Y2=0
r95 60 62 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=6.14 $Y=0 $X2=6.48
+ $Y2=0
r96 59 81 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=6.755 $Y=0 $X2=6.977
+ $Y2=0
r97 59 62 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=6.755 $Y=0 $X2=6.48
+ $Y2=0
r98 58 79 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=6
+ $Y2=0
r99 58 76 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=5.04
+ $Y2=0
r100 57 58 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r101 55 75 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.15 $Y=0 $X2=4.985
+ $Y2=0
r102 55 57 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=5.15 $Y=0 $X2=5.52
+ $Y2=0
r103 54 78 7.94884 $w=1.7e-07 $l=1.47e-07 $layer=LI1_cond $X=5.845 $Y=0
+ $X2=5.992 $Y2=0
r104 54 57 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=5.845 $Y=0
+ $X2=5.52 $Y2=0
r105 53 76 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=5.04
+ $Y2=0
r106 52 53 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r107 50 72 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.145 $Y=0 $X2=2.98
+ $Y2=0
r108 50 52 92.3155 $w=1.68e-07 $l=1.415e-06 $layer=LI1_cond $X=3.145 $Y=0
+ $X2=4.56 $Y2=0
r109 49 75 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.82 $Y=0 $X2=4.985
+ $Y2=0
r110 49 52 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=4.82 $Y=0 $X2=4.56
+ $Y2=0
r111 48 73 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r112 47 48 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r113 45 48 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=1.2 $Y=0 $X2=2.64
+ $Y2=0
r114 45 67 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r115 44 47 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.2 $Y=0 $X2=2.64
+ $Y2=0
r116 44 45 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r117 42 66 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.955 $Y=0 $X2=0.79
+ $Y2=0
r118 42 44 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=0.955 $Y=0 $X2=1.2
+ $Y2=0
r119 41 72 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.815 $Y=0 $X2=2.98
+ $Y2=0
r120 41 47 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=2.815 $Y=0
+ $X2=2.64 $Y2=0
r121 39 67 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r122 38 39 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r123 36 66 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.625 $Y=0 $X2=0.79
+ $Y2=0
r124 36 38 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=0.625 $Y=0
+ $X2=0.24 $Y2=0
r125 34 53 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.56
+ $Y2=0
r126 34 73 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=3.12
+ $Y2=0
r127 30 81 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=6.92 $Y=0.085
+ $X2=6.977 $Y2=0
r128 30 32 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=6.92 $Y=0.085
+ $X2=6.92 $Y2=0.515
r129 26 78 0.543863 $w=2.95e-07 $l=8.5e-08 $layer=LI1_cond $X=5.992 $Y=0.085
+ $X2=5.992 $Y2=0
r130 26 28 16.7983 $w=2.93e-07 $l=4.3e-07 $layer=LI1_cond $X=5.992 $Y=0.085
+ $X2=5.992 $Y2=0.515
r131 22 24 13.0959 $w=3.28e-07 $l=3.75e-07 $layer=LI1_cond $X=4.985 $Y=0.515
+ $X2=4.985 $Y2=0.89
r132 20 75 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.985 $Y=0.085
+ $X2=4.985 $Y2=0
r133 20 22 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=4.985 $Y=0.085
+ $X2=4.985 $Y2=0.515
r134 16 72 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.98 $Y=0.085
+ $X2=2.98 $Y2=0
r135 16 18 15.8897 $w=3.28e-07 $l=4.55e-07 $layer=LI1_cond $X=2.98 $Y=0.085
+ $X2=2.98 $Y2=0.54
r136 5 32 91 $w=1.7e-07 $l=2.26164e-07 $layer=licon1_NDIFF $count=2 $X=6.755
+ $Y=0.37 $X2=6.92 $Y2=0.515
r137 4 28 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=5.83
+ $Y=0.37 $X2=5.975 $Y2=0.515
r138 3 24 182 $w=1.7e-07 $l=3.02159e-07 $layer=licon1_NDIFF $count=1 $X=4.765
+ $Y=0.695 $X2=4.985 $Y2=0.89
r139 3 22 182 $w=1.7e-07 $l=2.96648e-07 $layer=licon1_NDIFF $count=1 $X=4.765
+ $Y=0.695 $X2=4.985 $Y2=0.515
r140 2 18 91 $w=1.7e-07 $l=6.29285e-07 $layer=licon1_NDIFF $count=2 $X=2.43
+ $Y=0.37 $X2=2.98 $Y2=0.54
r141 1 69 182 $w=1.7e-07 $l=3.68951e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.6 $X2=0.79 $Y2=0.325
.ends

