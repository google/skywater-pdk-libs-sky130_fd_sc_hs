* File: sky130_fd_sc_hs__o311ai_4.pex.spice
* Created: Thu Aug 27 21:02:19 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HS__O311AI_4%C1 1 3 4 6 7 9 10 12 13 15 16 17 18 20 21
+ 22 33
c66 33 0 7.45181e-20 $X=1.075 $Y=1.465
c67 16 0 4.49374e-20 $X=1.715 $Y=1.26
r68 32 34 11.3986 $w=4.44e-07 $l=1.05e-07 $layer=POLY_cond $X=1.075 $Y=1.475
+ $X2=1.18 $Y2=1.475
r69 32 33 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.075
+ $Y=1.465 $X2=1.075 $Y2=1.465
r70 30 32 15.741 $w=4.44e-07 $l=1.45e-07 $layer=POLY_cond $X=0.93 $Y=1.475
+ $X2=1.075 $Y2=1.475
r71 29 30 46.1374 $w=4.44e-07 $l=4.25e-07 $layer=POLY_cond $X=0.505 $Y=1.475
+ $X2=0.93 $Y2=1.475
r72 28 29 1.08559 $w=4.44e-07 $l=1e-08 $layer=POLY_cond $X=0.495 $Y=1.475
+ $X2=0.505 $Y2=1.475
r73 26 28 10.8559 $w=4.44e-07 $l=1e-07 $layer=POLY_cond $X=0.395 $Y=1.475
+ $X2=0.495 $Y2=1.475
r74 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.395
+ $Y=1.465 $X2=0.395 $Y2=1.465
r75 22 33 8.846 $w=4.78e-07 $l=3.55e-07 $layer=LI1_cond $X=0.72 $Y=1.54
+ $X2=1.075 $Y2=1.54
r76 22 27 8.09845 $w=4.78e-07 $l=3.25e-07 $layer=LI1_cond $X=0.72 $Y=1.54
+ $X2=0.395 $Y2=1.54
r77 21 27 3.86234 $w=4.78e-07 $l=1.55e-07 $layer=LI1_cond $X=0.24 $Y=1.54
+ $X2=0.395 $Y2=1.54
r78 18 20 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=1.79 $Y=1.185
+ $X2=1.79 $Y2=0.74
r79 16 18 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.715 $Y=1.26
+ $X2=1.79 $Y2=1.185
r80 16 17 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=1.715 $Y=1.26
+ $X2=1.435 $Y2=1.26
r81 13 17 30.7687 $w=4.44e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.36 $Y=1.185
+ $X2=1.435 $Y2=1.26
r82 13 34 19.5405 $w=4.44e-07 $l=3.69188e-07 $layer=POLY_cond $X=1.36 $Y=1.185
+ $X2=1.18 $Y2=1.475
r83 13 15 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=1.36 $Y=1.185
+ $X2=1.36 $Y2=0.74
r84 10 34 28.433 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=1.18 $Y=1.765
+ $X2=1.18 $Y2=1.475
r85 10 12 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.18 $Y=1.765
+ $X2=1.18 $Y2=2.4
r86 7 30 28.433 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=0.93 $Y=1.185 $X2=0.93
+ $Y2=1.475
r87 7 9 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=0.93 $Y=1.185
+ $X2=0.93 $Y2=0.74
r88 4 29 28.433 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=0.505 $Y=1.765
+ $X2=0.505 $Y2=1.475
r89 4 6 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.505 $Y=1.765
+ $X2=0.505 $Y2=2.4
r90 1 28 28.433 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=0.495 $Y=1.185
+ $X2=0.495 $Y2=1.475
r91 1 3 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=0.495 $Y=1.185
+ $X2=0.495 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HS__O311AI_4%B1 1 3 4 5 6 8 11 15 19 23 25 26 27 28 41
c66 1 0 7.45181e-20 $X=1.68 $Y=1.765
r67 41 43 11.9176 $w=3.64e-07 $l=9e-08 $layer=POLY_cond $X=3.43 $Y=1.557
+ $X2=3.52 $Y2=1.557
r68 41 42 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.43
+ $Y=1.515 $X2=3.43 $Y2=1.515
r69 39 41 46.3462 $w=3.64e-07 $l=3.5e-07 $layer=POLY_cond $X=3.08 $Y=1.557
+ $X2=3.43 $Y2=1.557
r70 38 39 56.9396 $w=3.64e-07 $l=4.3e-07 $layer=POLY_cond $X=2.65 $Y=1.557
+ $X2=3.08 $Y2=1.557
r71 36 38 31.7802 $w=3.64e-07 $l=2.4e-07 $layer=POLY_cond $X=2.41 $Y=1.557
+ $X2=2.65 $Y2=1.557
r72 36 37 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.41
+ $Y=1.515 $X2=2.41 $Y2=1.515
r73 34 36 25.1593 $w=3.64e-07 $l=1.9e-07 $layer=POLY_cond $X=2.22 $Y=1.557
+ $X2=2.41 $Y2=1.557
r74 27 28 15.8049 $w=3.48e-07 $l=4.8e-07 $layer=LI1_cond $X=3.6 $Y=1.605
+ $X2=4.08 $Y2=1.605
r75 27 42 5.59758 $w=3.48e-07 $l=1.7e-07 $layer=LI1_cond $X=3.6 $Y=1.605
+ $X2=3.43 $Y2=1.605
r76 26 42 10.2074 $w=3.48e-07 $l=3.1e-07 $layer=LI1_cond $X=3.12 $Y=1.605
+ $X2=3.43 $Y2=1.605
r77 25 26 15.8049 $w=3.48e-07 $l=4.8e-07 $layer=LI1_cond $X=2.64 $Y=1.605
+ $X2=3.12 $Y2=1.605
r78 25 37 7.5732 $w=3.48e-07 $l=2.3e-07 $layer=LI1_cond $X=2.64 $Y=1.605
+ $X2=2.41 $Y2=1.605
r79 21 43 23.572 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.52 $Y=1.35
+ $X2=3.52 $Y2=1.557
r80 21 23 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=3.52 $Y=1.35
+ $X2=3.52 $Y2=0.74
r81 17 39 23.572 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.08 $Y=1.35
+ $X2=3.08 $Y2=1.557
r82 17 19 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=3.08 $Y=1.35
+ $X2=3.08 $Y2=0.74
r83 13 38 23.572 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.65 $Y=1.35
+ $X2=2.65 $Y2=1.557
r84 13 15 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.65 $Y=1.35
+ $X2=2.65 $Y2=0.74
r85 9 34 23.572 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.22 $Y=1.35 $X2=2.22
+ $Y2=1.557
r86 9 11 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.22 $Y=1.35 $X2=2.22
+ $Y2=0.74
r87 6 34 11.9176 $w=3.64e-07 $l=2.48966e-07 $layer=POLY_cond $X=2.13 $Y=1.765
+ $X2=2.22 $Y2=1.557
r88 6 8 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.13 $Y=1.765
+ $X2=2.13 $Y2=2.4
r89 4 6 29.035 $w=3.64e-07 $l=1.53542e-07 $layer=POLY_cond $X=2.04 $Y=1.65
+ $X2=2.13 $Y2=1.765
r90 4 5 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=2.04 $Y=1.65 $X2=1.77
+ $Y2=1.65
r91 1 5 26.9307 $w=1.5e-07 $l=1.53542e-07 $layer=POLY_cond $X=1.68 $Y=1.765
+ $X2=1.77 $Y2=1.65
r92 1 3 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.68 $Y=1.765
+ $X2=1.68 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_HS__O311AI_4%A3 1 3 6 8 10 13 15 17 20 22 24 27 34 35 51
+ 52 54 61 64
r98 54 64 0.493904 $w=3.48e-07 $l=1.5e-08 $layer=LI1_cond $X=5.535 $Y=1.605
+ $X2=5.52 $Y2=1.605
r99 52 53 1.99174 $w=3.63e-07 $l=1.5e-08 $layer=POLY_cond $X=6.225 $Y=1.557
+ $X2=6.24 $Y2=1.557
r100 50 52 25.8926 $w=3.63e-07 $l=1.95e-07 $layer=POLY_cond $X=6.03 $Y=1.557
+ $X2=6.225 $Y2=1.557
r101 50 51 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.03
+ $Y=1.515 $X2=6.03 $Y2=1.515
r102 48 50 29.2121 $w=3.63e-07 $l=2.2e-07 $layer=POLY_cond $X=5.81 $Y=1.557
+ $X2=6.03 $Y2=1.557
r103 47 48 28.5482 $w=3.63e-07 $l=2.15e-07 $layer=POLY_cond $X=5.595 $Y=1.557
+ $X2=5.81 $Y2=1.557
r104 46 61 7.26255 $w=3.48e-07 $l=1.65e-07 $layer=LI1_cond $X=5.35 $Y=1.605
+ $X2=5.185 $Y2=1.605
r105 45 47 32.5317 $w=3.63e-07 $l=2.45e-07 $layer=POLY_cond $X=5.35 $Y=1.557
+ $X2=5.595 $Y2=1.557
r106 45 46 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.35
+ $Y=1.515 $X2=5.35 $Y2=1.515
r107 43 45 17.2617 $w=3.63e-07 $l=1.3e-07 $layer=POLY_cond $X=5.22 $Y=1.557
+ $X2=5.35 $Y2=1.557
r108 42 43 19.2534 $w=3.63e-07 $l=1.45e-07 $layer=POLY_cond $X=5.075 $Y=1.557
+ $X2=5.22 $Y2=1.557
r109 39 40 28.5482 $w=3.63e-07 $l=2.15e-07 $layer=POLY_cond $X=4.575 $Y=1.557
+ $X2=4.79 $Y2=1.557
r110 35 51 0.987808 $w=3.48e-07 $l=3e-08 $layer=LI1_cond $X=6 $Y=1.605 $X2=6.03
+ $Y2=1.605
r111 34 64 1.15244 $w=3.48e-07 $l=3.5e-08 $layer=LI1_cond $X=5.485 $Y=1.605
+ $X2=5.52 $Y2=1.605
r112 34 46 4.44514 $w=3.48e-07 $l=1.35e-07 $layer=LI1_cond $X=5.485 $Y=1.605
+ $X2=5.35 $Y2=1.605
r113 34 35 14.1586 $w=3.48e-07 $l=4.3e-07 $layer=LI1_cond $X=5.57 $Y=1.605 $X2=6
+ $Y2=1.605
r114 34 54 1.15244 $w=3.48e-07 $l=3.5e-08 $layer=LI1_cond $X=5.57 $Y=1.605
+ $X2=5.535 $Y2=1.605
r115 32 42 8.63085 $w=3.63e-07 $l=6.5e-08 $layer=POLY_cond $X=5.01 $Y=1.557
+ $X2=5.075 $Y2=1.557
r116 32 40 29.2121 $w=3.63e-07 $l=2.2e-07 $layer=POLY_cond $X=5.01 $Y=1.557
+ $X2=4.79 $Y2=1.557
r117 31 61 9.24242 $w=2.08e-07 $l=1.75e-07 $layer=LI1_cond $X=5.01 $Y=1.535
+ $X2=5.185 $Y2=1.535
r118 31 32 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.01
+ $Y=1.515 $X2=5.01 $Y2=1.515
r119 25 53 23.5056 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=6.24 $Y=1.35
+ $X2=6.24 $Y2=1.557
r120 25 27 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=6.24 $Y=1.35
+ $X2=6.24 $Y2=0.74
r121 22 52 23.5056 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=6.225 $Y=1.765
+ $X2=6.225 $Y2=1.557
r122 22 24 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=6.225 $Y=1.765
+ $X2=6.225 $Y2=2.4
r123 18 48 23.5056 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=5.81 $Y=1.35
+ $X2=5.81 $Y2=1.557
r124 18 20 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=5.81 $Y=1.35
+ $X2=5.81 $Y2=0.74
r125 15 47 23.5056 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=5.595 $Y=1.765
+ $X2=5.595 $Y2=1.557
r126 15 17 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=5.595 $Y=1.765
+ $X2=5.595 $Y2=2.4
r127 11 43 23.5056 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=5.22 $Y=1.35
+ $X2=5.22 $Y2=1.557
r128 11 13 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=5.22 $Y=1.35
+ $X2=5.22 $Y2=0.74
r129 8 42 23.5056 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=5.075 $Y=1.765
+ $X2=5.075 $Y2=1.557
r130 8 10 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=5.075 $Y=1.765
+ $X2=5.075 $Y2=2.4
r131 4 40 23.5056 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.79 $Y=1.35
+ $X2=4.79 $Y2=1.557
r132 4 6 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=4.79 $Y=1.35 $X2=4.79
+ $Y2=0.74
r133 1 39 23.5056 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=4.575 $Y=1.765
+ $X2=4.575 $Y2=1.557
r134 1 3 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=4.575 $Y=1.765
+ $X2=4.575 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_HS__O311AI_4%A2 1 3 6 8 10 13 15 17 18 20 21 23 24 26 27
+ 28 40 43
c89 43 0 1.39068e-19 $X=8.175 $Y=1.482
c90 24 0 5.87245e-20 $X=8.245 $Y=1.2
c91 13 0 1.36796e-19 $X=7.27 $Y=0.74
c92 8 0 9.21518e-20 $X=7.175 $Y=1.765
c93 6 0 5.58611e-20 $X=6.84 $Y=0.74
r94 43 44 8.33086 $w=4.05e-07 $l=7e-08 $layer=POLY_cond $X=8.175 $Y=1.482
+ $X2=8.245 $Y2=1.482
r95 42 43 51.7704 $w=4.05e-07 $l=4.35e-07 $layer=POLY_cond $X=7.74 $Y=1.482
+ $X2=8.175 $Y2=1.482
r96 41 42 1.78519 $w=4.05e-07 $l=1.5e-08 $layer=POLY_cond $X=7.725 $Y=1.482
+ $X2=7.74 $Y2=1.482
r97 39 41 13.6864 $w=4.05e-07 $l=1.15e-07 $layer=POLY_cond $X=7.61 $Y=1.482
+ $X2=7.725 $Y2=1.482
r98 39 40 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=7.61
+ $Y=1.515 $X2=7.61 $Y2=1.515
r99 34 36 29.158 $w=4.05e-07 $l=2.45e-07 $layer=POLY_cond $X=6.93 $Y=1.482
+ $X2=7.175 $Y2=1.482
r100 34 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.93
+ $Y=1.515 $X2=6.93 $Y2=1.515
r101 28 40 4.55617 $w=4.28e-07 $l=1.7e-07 $layer=LI1_cond $X=7.44 $Y=1.565
+ $X2=7.61 $Y2=1.565
r102 27 28 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=6.96 $Y=1.565
+ $X2=7.44 $Y2=1.565
r103 27 35 0.80403 $w=4.28e-07 $l=3e-08 $layer=LI1_cond $X=6.96 $Y=1.565
+ $X2=6.93 $Y2=1.565
r104 24 44 26.1659 $w=1.5e-07 $l=2.82e-07 $layer=POLY_cond $X=8.245 $Y=1.2
+ $X2=8.245 $Y2=1.482
r105 24 26 147.813 $w=1.5e-07 $l=4.6e-07 $layer=POLY_cond $X=8.245 $Y=1.2
+ $X2=8.245 $Y2=0.74
r106 21 43 26.1659 $w=1.5e-07 $l=2.83e-07 $layer=POLY_cond $X=8.175 $Y=1.765
+ $X2=8.175 $Y2=1.482
r107 21 23 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=8.175 $Y=1.765
+ $X2=8.175 $Y2=2.4
r108 18 42 26.1659 $w=1.5e-07 $l=2.82e-07 $layer=POLY_cond $X=7.74 $Y=1.2
+ $X2=7.74 $Y2=1.482
r109 18 20 147.813 $w=1.5e-07 $l=4.6e-07 $layer=POLY_cond $X=7.74 $Y=1.2
+ $X2=7.74 $Y2=0.74
r110 15 41 26.1659 $w=1.5e-07 $l=2.83e-07 $layer=POLY_cond $X=7.725 $Y=1.765
+ $X2=7.725 $Y2=1.482
r111 15 17 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=7.725 $Y=1.765
+ $X2=7.725 $Y2=2.4
r112 11 39 40.4642 $w=4.05e-07 $l=3.4e-07 $layer=POLY_cond $X=7.27 $Y=1.482
+ $X2=7.61 $Y2=1.482
r113 11 36 11.3062 $w=4.05e-07 $l=9.5e-08 $layer=POLY_cond $X=7.27 $Y=1.482
+ $X2=7.175 $Y2=1.482
r114 11 13 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=7.27 $Y=1.35
+ $X2=7.27 $Y2=0.74
r115 8 36 26.1659 $w=1.5e-07 $l=2.83e-07 $layer=POLY_cond $X=7.175 $Y=1.765
+ $X2=7.175 $Y2=1.482
r116 8 10 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=7.175 $Y=1.765
+ $X2=7.175 $Y2=2.4
r117 4 34 10.7111 $w=4.05e-07 $l=9e-08 $layer=POLY_cond $X=6.84 $Y=1.482
+ $X2=6.93 $Y2=1.482
r118 4 31 19.637 $w=4.05e-07 $l=1.65e-07 $layer=POLY_cond $X=6.84 $Y=1.482
+ $X2=6.675 $Y2=1.482
r119 4 6 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=6.84 $Y=1.35 $X2=6.84
+ $Y2=0.74
r120 1 31 26.1659 $w=1.5e-07 $l=2.83e-07 $layer=POLY_cond $X=6.675 $Y=1.765
+ $X2=6.675 $Y2=1.482
r121 1 3 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=6.675 $Y=1.765
+ $X2=6.675 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_HS__O311AI_4%A1 3 5 6 9 11 13 14 16 17 19 20 22 23 25 26
+ 28 29 30 31 45 46
c81 26 0 1.65594e-19 $X=10.545 $Y=1.2
r82 46 47 1.13679 $w=4.24e-07 $l=1e-08 $layer=POLY_cond $X=10.535 $Y=1.482
+ $X2=10.545 $Y2=1.482
r83 44 46 21.0307 $w=4.24e-07 $l=1.85e-07 $layer=POLY_cond $X=10.35 $Y=1.482
+ $X2=10.535 $Y2=1.482
r84 44 45 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=10.35
+ $Y=1.515 $X2=10.35 $Y2=1.515
r85 42 44 28.4198 $w=4.24e-07 $l=2.5e-07 $layer=POLY_cond $X=10.1 $Y=1.482
+ $X2=10.35 $Y2=1.482
r86 41 42 1.70519 $w=4.24e-07 $l=1.5e-08 $layer=POLY_cond $X=10.085 $Y=1.482
+ $X2=10.1 $Y2=1.482
r87 40 41 51.1557 $w=4.24e-07 $l=4.5e-07 $layer=POLY_cond $X=9.635 $Y=1.482
+ $X2=10.085 $Y2=1.482
r88 38 40 34.6722 $w=4.24e-07 $l=3.05e-07 $layer=POLY_cond $X=9.33 $Y=1.482
+ $X2=9.635 $Y2=1.482
r89 38 39 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=9.33
+ $Y=1.515 $X2=9.33 $Y2=1.515
r90 36 38 16.4835 $w=4.24e-07 $l=1.45e-07 $layer=POLY_cond $X=9.185 $Y=1.482
+ $X2=9.33 $Y2=1.482
r91 31 45 0.80403 $w=4.28e-07 $l=3e-08 $layer=LI1_cond $X=10.32 $Y=1.565
+ $X2=10.35 $Y2=1.565
r92 30 31 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=9.84 $Y=1.565
+ $X2=10.32 $Y2=1.565
r93 29 30 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=9.36 $Y=1.565
+ $X2=9.84 $Y2=1.565
r94 29 39 0.80403 $w=4.28e-07 $l=3e-08 $layer=LI1_cond $X=9.36 $Y=1.565 $X2=9.33
+ $Y2=1.565
r95 26 47 27.2926 $w=1.5e-07 $l=2.82e-07 $layer=POLY_cond $X=10.545 $Y=1.2
+ $X2=10.545 $Y2=1.482
r96 26 28 147.813 $w=1.5e-07 $l=4.6e-07 $layer=POLY_cond $X=10.545 $Y=1.2
+ $X2=10.545 $Y2=0.74
r97 23 46 27.2926 $w=1.5e-07 $l=2.83e-07 $layer=POLY_cond $X=10.535 $Y=1.765
+ $X2=10.535 $Y2=1.482
r98 23 25 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=10.535 $Y=1.765
+ $X2=10.535 $Y2=2.4
r99 20 42 27.2926 $w=1.5e-07 $l=2.82e-07 $layer=POLY_cond $X=10.1 $Y=1.2
+ $X2=10.1 $Y2=1.482
r100 20 22 147.813 $w=1.5e-07 $l=4.6e-07 $layer=POLY_cond $X=10.1 $Y=1.2
+ $X2=10.1 $Y2=0.74
r101 17 41 27.2926 $w=1.5e-07 $l=2.83e-07 $layer=POLY_cond $X=10.085 $Y=1.765
+ $X2=10.085 $Y2=1.482
r102 17 19 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=10.085 $Y=1.765
+ $X2=10.085 $Y2=2.4
r103 14 40 27.2926 $w=1.5e-07 $l=2.83e-07 $layer=POLY_cond $X=9.635 $Y=1.765
+ $X2=9.635 $Y2=1.482
r104 14 16 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=9.635 $Y=1.765
+ $X2=9.635 $Y2=2.4
r105 11 36 27.2926 $w=1.5e-07 $l=2.83e-07 $layer=POLY_cond $X=9.185 $Y=1.765
+ $X2=9.185 $Y2=1.482
r106 11 13 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=9.185 $Y=1.765
+ $X2=9.185 $Y2=2.4
r107 7 36 9.09434 $w=4.24e-07 $l=8e-08 $layer=POLY_cond $X=9.105 $Y=1.482
+ $X2=9.185 $Y2=1.482
r108 7 9 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=9.105 $Y=1.35
+ $X2=9.105 $Y2=0.74
r109 5 7 29.854 $w=4.24e-07 $l=1.56058e-07 $layer=POLY_cond $X=9.03 $Y=1.605
+ $X2=9.105 $Y2=1.482
r110 5 6 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=9.03 $Y=1.605
+ $X2=8.75 $Y2=1.605
r111 1 6 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=8.675 $Y=1.53
+ $X2=8.75 $Y2=1.605
r112 1 3 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=8.675 $Y=1.53
+ $X2=8.675 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HS__O311AI_4%VPWR 1 2 3 4 5 6 19 21 27 31 35 37 39 44 45
+ 46 56 64 69 79 88 90 93 97
r113 96 97 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.8 $Y=3.33
+ $X2=10.8 $Y2=3.33
r114 93 94 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.84 $Y=3.33
+ $X2=9.84 $Y2=3.33
r115 90 91 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r116 87 88 13.5255 $w=1.123e-06 $l=1.65e-07 $layer=LI1_cond $X=3.74 $Y=2.852
+ $X2=3.905 $Y2=2.852
r117 84 87 1.51822 $w=1.123e-06 $l=1.4e-07 $layer=LI1_cond $X=3.6 $Y=2.852
+ $X2=3.74 $Y2=2.852
r118 84 85 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r119 82 85 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.6 $Y2=3.33
r120 81 84 10.4107 $w=1.123e-06 $l=9.6e-07 $layer=LI1_cond $X=2.64 $Y=2.852
+ $X2=3.6 $Y2=2.852
r121 81 82 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r122 78 81 3.09067 $w=1.123e-06 $l=2.85e-07 $layer=LI1_cond $X=2.355 $Y=2.852
+ $X2=2.64 $Y2=2.852
r123 78 79 12.9833 $w=1.123e-06 $l=1.15e-07 $layer=LI1_cond $X=2.355 $Y=2.852
+ $X2=2.24 $Y2=2.852
r124 75 76 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r125 73 97 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.32 $Y=3.33
+ $X2=10.8 $Y2=3.33
r126 73 94 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.32 $Y=3.33
+ $X2=9.84 $Y2=3.33
r127 72 73 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.32 $Y=3.33
+ $X2=10.32 $Y2=3.33
r128 70 93 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.025 $Y=3.33
+ $X2=9.86 $Y2=3.33
r129 70 72 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=10.025 $Y=3.33
+ $X2=10.32 $Y2=3.33
r130 69 96 4.01252 $w=1.7e-07 $l=1.82e-07 $layer=LI1_cond $X=10.675 $Y=3.33
+ $X2=10.857 $Y2=3.33
r131 69 72 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=10.675 $Y=3.33
+ $X2=10.32 $Y2=3.33
r132 68 94 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.36 $Y=3.33
+ $X2=9.84 $Y2=3.33
r133 68 91 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.36 $Y=3.33
+ $X2=8.88 $Y2=3.33
r134 67 68 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.36 $Y=3.33
+ $X2=9.36 $Y2=3.33
r135 65 90 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.125 $Y=3.33
+ $X2=8.96 $Y2=3.33
r136 65 67 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=9.125 $Y=3.33
+ $X2=9.36 $Y2=3.33
r137 64 93 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.695 $Y=3.33
+ $X2=9.86 $Y2=3.33
r138 64 67 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=9.695 $Y=3.33
+ $X2=9.36 $Y2=3.33
r139 63 91 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=3.33
+ $X2=8.88 $Y2=3.33
r140 62 63 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=8.4 $Y=3.33
+ $X2=8.4 $Y2=3.33
r141 60 85 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=3.6 $Y2=3.33
r142 59 62 281.84 $w=1.68e-07 $l=4.32e-06 $layer=LI1_cond $X=4.08 $Y=3.33
+ $X2=8.4 $Y2=3.33
r143 59 88 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=4.08 $Y=3.33
+ $X2=3.905 $Y2=3.33
r144 59 60 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r145 56 90 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.795 $Y=3.33
+ $X2=8.96 $Y2=3.33
r146 56 62 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=8.795 $Y=3.33
+ $X2=8.4 $Y2=3.33
r147 55 82 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r148 54 79 5.21925 $w=1.68e-07 $l=8e-08 $layer=LI1_cond $X=2.16 $Y=3.33 $X2=2.24
+ $Y2=3.33
r149 54 55 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r150 51 55 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.16 $Y2=3.33
r151 51 76 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.24 $Y2=3.33
r152 50 51 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r153 48 75 4.73185 $w=1.7e-07 $l=2.23e-07 $layer=LI1_cond $X=0.445 $Y=3.33
+ $X2=0.222 $Y2=3.33
r154 48 50 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=0.445 $Y=3.33
+ $X2=1.2 $Y2=3.33
r155 46 63 0.802756 $w=4.9e-07 $l=2.88e-06 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=8.4 $Y2=3.33
r156 46 60 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=4.08 $Y2=3.33
r157 44 50 2.60963 $w=1.68e-07 $l=4e-08 $layer=LI1_cond $X=1.24 $Y=3.33 $X2=1.2
+ $Y2=3.33
r158 44 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.24 $Y=3.33
+ $X2=1.405 $Y2=3.33
r159 43 54 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=1.57 $Y=3.33
+ $X2=2.16 $Y2=3.33
r160 43 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.57 $Y=3.33
+ $X2=1.405 $Y2=3.33
r161 39 42 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=10.8 $Y=1.985
+ $X2=10.8 $Y2=2.815
r162 37 96 3.13065 $w=2.5e-07 $l=1.09864e-07 $layer=LI1_cond $X=10.8 $Y=3.245
+ $X2=10.857 $Y2=3.33
r163 37 42 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=10.8 $Y=3.245
+ $X2=10.8 $Y2=2.815
r164 33 93 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.86 $Y=3.245
+ $X2=9.86 $Y2=3.33
r165 33 35 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=9.86 $Y=3.245
+ $X2=9.86 $Y2=2.415
r166 29 90 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.96 $Y=3.245
+ $X2=8.96 $Y2=3.33
r167 29 31 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=8.96 $Y=3.245
+ $X2=8.96 $Y2=2.415
r168 25 45 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.405 $Y=3.245
+ $X2=1.405 $Y2=3.33
r169 25 27 27.5888 $w=3.28e-07 $l=7.9e-07 $layer=LI1_cond $X=1.405 $Y=3.245
+ $X2=1.405 $Y2=2.455
r170 21 24 24.4458 $w=3.28e-07 $l=7e-07 $layer=LI1_cond $X=0.28 $Y=2.115
+ $X2=0.28 $Y2=2.815
r171 19 75 3.03433 $w=3.3e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.28 $Y=3.245
+ $X2=0.222 $Y2=3.33
r172 19 24 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=0.28 $Y=3.245
+ $X2=0.28 $Y2=2.815
r173 6 42 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=10.61
+ $Y=1.84 $X2=10.76 $Y2=2.815
r174 6 39 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=10.61
+ $Y=1.84 $X2=10.76 $Y2=1.985
r175 5 35 300 $w=1.7e-07 $l=6.45659e-07 $layer=licon1_PDIFF $count=2 $X=9.71
+ $Y=1.84 $X2=9.86 $Y2=2.415
r176 4 31 300 $w=1.7e-07 $l=6.43428e-07 $layer=licon1_PDIFF $count=2 $X=8.815
+ $Y=1.84 $X2=8.96 $Y2=2.415
r177 3 87 120 $w=1.7e-07 $l=1.81666e-06 $layer=licon1_PDIFF $count=5 $X=2.205
+ $Y=1.84 $X2=3.74 $Y2=2.455
r178 3 78 120 $w=1.7e-07 $l=6.85912e-07 $layer=licon1_PDIFF $count=5 $X=2.205
+ $Y=1.84 $X2=2.355 $Y2=2.455
r179 2 27 300 $w=1.7e-07 $l=6.85912e-07 $layer=licon1_PDIFF $count=2 $X=1.255
+ $Y=1.84 $X2=1.405 $Y2=2.455
r180 1 24 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.815
r181 1 21 400 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.115
.ends

.subckt PM_SKY130_FD_SC_HS__O311AI_4%Y 1 2 3 4 5 6 23 25 27 29 33 35 39 41 45 51
+ 52 54 56 58 60 61 65 67
c137 54 0 4.49374e-20 $X=1.905 $Y=1.985
r138 65 67 1.75372 $w=2.28e-07 $l=3.5e-08 $layer=LI1_cond $X=6.48 $Y=1.26
+ $X2=6.48 $Y2=1.295
r139 60 65 2.9826 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.48 $Y=1.175
+ $X2=6.48 $Y2=1.26
r140 60 61 17.2866 $w=2.28e-07 $l=3.45e-07 $layer=LI1_cond $X=6.48 $Y=1.32
+ $X2=6.48 $Y2=1.665
r141 60 67 1.25266 $w=2.28e-07 $l=2.5e-08 $layer=LI1_cond $X=6.48 $Y=1.32
+ $X2=6.48 $Y2=1.295
r142 59 61 14.2803 $w=2.28e-07 $l=2.85e-07 $layer=LI1_cond $X=6.48 $Y=1.95
+ $X2=6.48 $Y2=1.665
r143 50 52 9.45624 $w=4.88e-07 $l=1.65e-07 $layer=LI1_cond $X=1.575 $Y=1.015
+ $X2=1.74 $Y2=1.015
r144 50 51 5.30815 $w=4.88e-07 $l=1.65e-07 $layer=LI1_cond $X=1.575 $Y=1.015
+ $X2=1.41 $Y2=1.015
r145 46 58 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.015 $Y=2.035
+ $X2=5.85 $Y2=2.035
r146 45 59 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=6.365 $Y=2.035
+ $X2=6.48 $Y2=1.95
r147 45 46 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=6.365 $Y=2.035
+ $X2=6.015 $Y2=2.035
r148 42 56 8.61065 $w=1.7e-07 $l=1.94808e-07 $layer=LI1_cond $X=5.015 $Y=2.035
+ $X2=4.85 $Y2=1.97
r149 41 58 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.685 $Y=2.035
+ $X2=5.85 $Y2=2.035
r150 41 42 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.685 $Y=2.035
+ $X2=5.015 $Y2=2.035
r151 37 56 0.89609 $w=3.3e-07 $l=1.5e-07 $layer=LI1_cond $X=4.85 $Y=2.12
+ $X2=4.85 $Y2=1.97
r152 37 39 6.63528 $w=3.28e-07 $l=1.9e-07 $layer=LI1_cond $X=4.85 $Y=2.12
+ $X2=4.85 $Y2=2.31
r153 36 54 8.61065 $w=1.7e-07 $l=1.94808e-07 $layer=LI1_cond $X=2.07 $Y=2.035
+ $X2=1.905 $Y2=1.97
r154 35 56 8.61065 $w=1.7e-07 $l=1.94808e-07 $layer=LI1_cond $X=4.685 $Y=2.035
+ $X2=4.85 $Y2=1.97
r155 35 36 170.604 $w=1.68e-07 $l=2.615e-06 $layer=LI1_cond $X=4.685 $Y=2.035
+ $X2=2.07 $Y2=2.035
r156 31 54 0.89609 $w=3.3e-07 $l=1.5e-07 $layer=LI1_cond $X=1.905 $Y=2.12
+ $X2=1.905 $Y2=1.97
r157 31 33 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=1.905 $Y=2.12
+ $X2=1.905 $Y2=2.815
r158 29 60 4.03528 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=6.365 $Y=1.175
+ $X2=6.48 $Y2=1.175
r159 29 52 301.738 $w=1.68e-07 $l=4.625e-06 $layer=LI1_cond $X=6.365 $Y=1.175
+ $X2=1.74 $Y2=1.175
r160 28 48 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.07 $Y=2.035
+ $X2=0.905 $Y2=2.035
r161 27 54 8.61065 $w=1.7e-07 $l=1.94808e-07 $layer=LI1_cond $X=1.74 $Y=2.035
+ $X2=1.905 $Y2=1.97
r162 27 28 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.74 $Y=2.035
+ $X2=1.07 $Y2=2.035
r163 23 48 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.905 $Y=2.12
+ $X2=0.905 $Y2=2.035
r164 23 25 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=0.905 $Y=2.12
+ $X2=0.905 $Y2=2.815
r165 21 51 24.4458 $w=3.28e-07 $l=7e-07 $layer=LI1_cond $X=0.71 $Y=0.935
+ $X2=1.41 $Y2=0.935
r166 6 58 300 $w=1.7e-07 $l=3.5373e-07 $layer=licon1_PDIFF $count=2 $X=5.67
+ $Y=1.84 $X2=5.85 $Y2=2.115
r167 5 56 600 $w=1.7e-07 $l=2.56905e-07 $layer=licon1_PDIFF $count=1 $X=4.65
+ $Y=1.84 $X2=4.85 $Y2=1.97
r168 5 39 300 $w=1.7e-07 $l=5.61159e-07 $layer=licon1_PDIFF $count=2 $X=4.65
+ $Y=1.84 $X2=4.85 $Y2=2.31
r169 4 54 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=1.755
+ $Y=1.84 $X2=1.905 $Y2=1.985
r170 4 33 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=1.755
+ $Y=1.84 $X2=1.905 $Y2=2.815
r171 3 48 400 $w=1.7e-07 $l=4.41588e-07 $layer=licon1_PDIFF $count=1 $X=0.58
+ $Y=1.84 $X2=0.905 $Y2=2.115
r172 3 25 400 $w=1.7e-07 $l=1.12583e-06 $layer=licon1_PDIFF $count=1 $X=0.58
+ $Y=1.84 $X2=0.905 $Y2=2.815
r173 2 50 182 $w=1.7e-07 $l=6.4622e-07 $layer=licon1_NDIFF $count=1 $X=1.435
+ $Y=0.37 $X2=1.575 $Y2=0.95
r174 1 21 182 $w=1.7e-07 $l=6.3113e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.37 $X2=0.71 $Y2=0.935
.ends

.subckt PM_SKY130_FD_SC_HS__O311AI_4%A_841_368# 1 2 3 4 5 18 20 21 24 26 30 32
+ 36 38 42 44 45 46
r71 40 42 17.112 $w=3.28e-07 $l=4.9e-07 $layer=LI1_cond $X=8.4 $Y=2.905 $X2=8.4
+ $Y2=2.415
r72 39 46 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.615 $Y=2.99
+ $X2=7.45 $Y2=2.99
r73 38 40 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=8.235 $Y=2.99
+ $X2=8.4 $Y2=2.905
r74 38 39 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=8.235 $Y=2.99
+ $X2=7.615 $Y2=2.99
r75 34 46 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.45 $Y=2.905
+ $X2=7.45 $Y2=2.99
r76 34 36 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=7.45 $Y=2.905
+ $X2=7.45 $Y2=2.455
r77 33 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.615 $Y=2.99
+ $X2=6.45 $Y2=2.99
r78 32 46 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.285 $Y=2.99
+ $X2=7.45 $Y2=2.99
r79 32 33 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=7.285 $Y=2.99
+ $X2=6.615 $Y2=2.99
r80 28 45 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.45 $Y=2.905
+ $X2=6.45 $Y2=2.99
r81 28 30 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=6.45 $Y=2.905
+ $X2=6.45 $Y2=2.455
r82 27 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.515 $Y=2.99
+ $X2=5.35 $Y2=2.99
r83 26 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.285 $Y=2.99
+ $X2=6.45 $Y2=2.99
r84 26 27 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=6.285 $Y=2.99
+ $X2=5.515 $Y2=2.99
r85 22 44 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.35 $Y=2.905
+ $X2=5.35 $Y2=2.99
r86 22 24 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=5.35 $Y=2.905
+ $X2=5.35 $Y2=2.455
r87 20 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.185 $Y=2.99
+ $X2=5.35 $Y2=2.99
r88 20 21 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.185 $Y=2.99
+ $X2=4.515 $Y2=2.99
r89 16 21 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.35 $Y=2.905
+ $X2=4.515 $Y2=2.99
r90 16 18 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=4.35 $Y=2.905
+ $X2=4.35 $Y2=2.455
r91 5 42 300 $w=1.7e-07 $l=6.45659e-07 $layer=licon1_PDIFF $count=2 $X=8.25
+ $Y=1.84 $X2=8.4 $Y2=2.415
r92 4 36 300 $w=1.7e-07 $l=7.07972e-07 $layer=licon1_PDIFF $count=2 $X=7.25
+ $Y=1.84 $X2=7.45 $Y2=2.455
r93 3 30 300 $w=1.7e-07 $l=6.85912e-07 $layer=licon1_PDIFF $count=2 $X=6.3
+ $Y=1.84 $X2=6.45 $Y2=2.455
r94 2 24 300 $w=1.7e-07 $l=7.07972e-07 $layer=licon1_PDIFF $count=2 $X=5.15
+ $Y=1.84 $X2=5.35 $Y2=2.455
r95 1 18 300 $w=1.7e-07 $l=6.83667e-07 $layer=licon1_PDIFF $count=2 $X=4.205
+ $Y=1.84 $X2=4.35 $Y2=2.455
.ends

.subckt PM_SKY130_FD_SC_HS__O311AI_4%A_1350_368# 1 2 3 4 15 19 21 25 27 29 31 34
+ 36 38
c56 36 0 9.21518e-20 $X=7.95 $Y=2.035
c57 21 0 1.39068e-19 $X=9.295 $Y=2.05
r58 29 40 2.94404 $w=2.8e-07 $l=1e-07 $layer=LI1_cond $X=10.335 $Y=2.15
+ $X2=10.335 $Y2=2.05
r59 29 31 12.5534 $w=2.78e-07 $l=3.05e-07 $layer=LI1_cond $X=10.335 $Y=2.15
+ $X2=10.335 $Y2=2.455
r60 28 38 5.79383 $w=2e-07 $l=1.15e-07 $layer=LI1_cond $X=9.525 $Y=2.05 $X2=9.41
+ $Y2=2.05
r61 27 40 4.12165 $w=2e-07 $l=1.4e-07 $layer=LI1_cond $X=10.195 $Y=2.05
+ $X2=10.335 $Y2=2.05
r62 27 28 37.1545 $w=1.98e-07 $l=6.7e-07 $layer=LI1_cond $X=10.195 $Y=2.05
+ $X2=9.525 $Y2=2.05
r63 23 38 0.844453 $w=2.3e-07 $l=1e-07 $layer=LI1_cond $X=9.41 $Y=2.15 $X2=9.41
+ $Y2=2.05
r64 23 25 15.2824 $w=2.28e-07 $l=3.05e-07 $layer=LI1_cond $X=9.41 $Y=2.15
+ $X2=9.41 $Y2=2.455
r65 22 36 7.18321 $w=1.85e-07 $l=1.4e-07 $layer=LI1_cond $X=8.065 $Y=2.05
+ $X2=7.925 $Y2=2.05
r66 21 38 5.79383 $w=2e-07 $l=1.15e-07 $layer=LI1_cond $X=9.295 $Y=2.05 $X2=9.41
+ $Y2=2.05
r67 21 22 68.2091 $w=1.98e-07 $l=1.23e-06 $layer=LI1_cond $X=9.295 $Y=2.05
+ $X2=8.065 $Y2=2.05
r68 17 36 0.097681 $w=2.8e-07 $l=1e-07 $layer=LI1_cond $X=7.925 $Y=2.15
+ $X2=7.925 $Y2=2.05
r69 17 19 17.2866 $w=2.78e-07 $l=4.2e-07 $layer=LI1_cond $X=7.925 $Y=2.15
+ $X2=7.925 $Y2=2.57
r70 16 34 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.115 $Y=2.035
+ $X2=6.95 $Y2=2.035
r71 15 36 7.18321 $w=1.85e-07 $l=1.47309e-07 $layer=LI1_cond $X=7.785 $Y=2.035
+ $X2=7.925 $Y2=2.05
r72 15 16 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=7.785 $Y=2.035
+ $X2=7.115 $Y2=2.035
r73 4 40 600 $w=1.7e-07 $l=2.59374e-07 $layer=licon1_PDIFF $count=1 $X=10.16
+ $Y=1.84 $X2=10.31 $Y2=2.035
r74 4 31 300 $w=1.7e-07 $l=6.85912e-07 $layer=licon1_PDIFF $count=2 $X=10.16
+ $Y=1.84 $X2=10.31 $Y2=2.455
r75 3 38 600 $w=1.7e-07 $l=2.59374e-07 $layer=licon1_PDIFF $count=1 $X=9.26
+ $Y=1.84 $X2=9.41 $Y2=2.035
r76 3 25 300 $w=1.7e-07 $l=6.85912e-07 $layer=licon1_PDIFF $count=2 $X=9.26
+ $Y=1.84 $X2=9.41 $Y2=2.455
r77 2 36 600 $w=1.7e-07 $l=2.59374e-07 $layer=licon1_PDIFF $count=1 $X=7.8
+ $Y=1.84 $X2=7.95 $Y2=2.035
r78 2 19 600 $w=1.7e-07 $l=8.01499e-07 $layer=licon1_PDIFF $count=1 $X=7.8
+ $Y=1.84 $X2=7.95 $Y2=2.57
r79 1 34 300 $w=1.7e-07 $l=3.61421e-07 $layer=licon1_PDIFF $count=2 $X=6.75
+ $Y=1.84 $X2=6.95 $Y2=2.115
.ends

.subckt PM_SKY130_FD_SC_HS__O311AI_4%A_27_74# 1 2 3 4 5 16 18 20 28 32
r40 30 32 56.7594 $w=1.68e-07 $l=8.7e-07 $layer=LI1_cond $X=2.865 $Y=0.835
+ $X2=3.735 $Y2=0.835
r41 28 30 50.5615 $w=1.68e-07 $l=7.75e-07 $layer=LI1_cond $X=2.09 $Y=0.835
+ $X2=2.865 $Y2=0.835
r42 25 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.005 $Y=0.75
+ $X2=2.09 $Y2=0.835
r43 25 27 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=2.005 $Y=0.75
+ $X2=2.005 $Y2=0.635
r44 24 27 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=2.005 $Y=0.6
+ $X2=2.005 $Y2=0.635
r45 21 35 3.40825 $w=2.5e-07 $l=1.25e-07 $layer=LI1_cond $X=0.365 $Y=0.475
+ $X2=0.24 $Y2=0.475
r46 21 23 35.9562 $w=2.48e-07 $l=7.8e-07 $layer=LI1_cond $X=0.365 $Y=0.475
+ $X2=1.145 $Y2=0.475
r47 20 24 7.14316 $w=2.5e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.92 $Y=0.475
+ $X2=2.005 $Y2=0.6
r48 20 23 35.7257 $w=2.48e-07 $l=7.75e-07 $layer=LI1_cond $X=1.92 $Y=0.475
+ $X2=1.145 $Y2=0.475
r49 16 35 3.40825 $w=2.5e-07 $l=1.25e-07 $layer=LI1_cond $X=0.24 $Y=0.6 $X2=0.24
+ $Y2=0.475
r50 16 18 16.8257 $w=2.48e-07 $l=3.65e-07 $layer=LI1_cond $X=0.24 $Y=0.6
+ $X2=0.24 $Y2=0.965
r51 5 32 182 $w=1.7e-07 $l=5.30401e-07 $layer=licon1_NDIFF $count=1 $X=3.595
+ $Y=0.37 $X2=3.735 $Y2=0.835
r52 4 30 182 $w=1.7e-07 $l=5.30401e-07 $layer=licon1_NDIFF $count=1 $X=2.725
+ $Y=0.37 $X2=2.865 $Y2=0.835
r53 3 27 182 $w=1.7e-07 $l=3.27605e-07 $layer=licon1_NDIFF $count=1 $X=1.865
+ $Y=0.37 $X2=2.005 $Y2=0.635
r54 2 23 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=1.005
+ $Y=0.37 $X2=1.145 $Y2=0.515
r55 1 35 182 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.515
r56 1 18 182 $w=1.7e-07 $l=6.63551e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.965
.ends

.subckt PM_SKY130_FD_SC_HS__O311AI_4%A_459_74# 1 2 3 4 5 6 7 8 25 32 33 34 37 39
+ 43 45 49 51 55 57 61 64 65 69 71 72 73 76 79
c149 79 0 5.87245e-20 $X=8.85 $Y=1.045
c150 73 0 1.36796e-19 $X=7.015 $Y=0.835
c151 65 0 1.65594e-19 $X=10.165 $Y=1.045
c152 51 0 5.58611e-20 $X=7.945 $Y=1.095
r153 76 77 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=8.03 $Y=1.095
+ $X2=8.03 $Y2=1.385
r154 73 74 11.9854 $w=2.48e-07 $l=2.6e-07 $layer=LI1_cond $X=7.015 $Y=0.835
+ $X2=7.015 $Y2=1.095
r155 67 69 20.5135 $w=2.48e-07 $l=4.45e-07 $layer=LI1_cond $X=10.29 $Y=0.96
+ $X2=10.29 $Y2=0.515
r156 66 79 2.76166 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.975 $Y=1.045
+ $X2=8.85 $Y2=1.045
r157 65 67 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=10.165 $Y=1.045
+ $X2=10.29 $Y2=0.96
r158 65 66 77.6364 $w=1.68e-07 $l=1.19e-06 $layer=LI1_cond $X=10.165 $Y=1.045
+ $X2=8.975 $Y2=1.045
r159 63 79 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=8.85 $Y=1.13
+ $X2=8.85 $Y2=1.045
r160 63 64 7.83661 $w=2.48e-07 $l=1.7e-07 $layer=LI1_cond $X=8.85 $Y=1.13
+ $X2=8.85 $Y2=1.3
r161 59 79 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=8.85 $Y=0.96
+ $X2=8.85 $Y2=1.045
r162 59 61 20.5135 $w=2.48e-07 $l=4.45e-07 $layer=LI1_cond $X=8.85 $Y=0.96
+ $X2=8.85 $Y2=0.515
r163 58 77 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.115 $Y=1.385
+ $X2=8.03 $Y2=1.385
r164 57 64 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=8.725 $Y=1.385
+ $X2=8.85 $Y2=1.3
r165 57 58 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=8.725 $Y=1.385
+ $X2=8.115 $Y2=1.385
r166 53 76 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=8.03 $Y=1.01
+ $X2=8.03 $Y2=1.095
r167 53 55 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=8.03 $Y=1.01
+ $X2=8.03 $Y2=0.515
r168 52 74 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.14 $Y=1.095
+ $X2=7.015 $Y2=1.095
r169 51 76 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.945 $Y=1.095
+ $X2=8.03 $Y2=1.095
r170 51 52 52.5187 $w=1.68e-07 $l=8.05e-07 $layer=LI1_cond $X=7.945 $Y=1.095
+ $X2=7.14 $Y2=1.095
r171 47 73 3.91831 $w=2.48e-07 $l=8.5e-08 $layer=LI1_cond $X=7.015 $Y=0.75
+ $X2=7.015 $Y2=0.835
r172 47 49 10.833 $w=2.48e-07 $l=2.35e-07 $layer=LI1_cond $X=7.015 $Y=0.75
+ $X2=7.015 $Y2=0.515
r173 46 72 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.19 $Y=0.835
+ $X2=6.025 $Y2=0.835
r174 45 73 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.89 $Y=0.835
+ $X2=7.015 $Y2=0.835
r175 45 46 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=6.89 $Y=0.835
+ $X2=6.19 $Y2=0.835
r176 41 72 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.025 $Y=0.75
+ $X2=6.025 $Y2=0.835
r177 41 43 4.01609 $w=3.28e-07 $l=1.15e-07 $layer=LI1_cond $X=6.025 $Y=0.75
+ $X2=6.025 $Y2=0.635
r178 40 71 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.17 $Y=0.835
+ $X2=5.045 $Y2=0.835
r179 39 72 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.86 $Y=0.835
+ $X2=6.025 $Y2=0.835
r180 39 40 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=5.86 $Y=0.835
+ $X2=5.17 $Y2=0.835
r181 35 71 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.045 $Y=0.75
+ $X2=5.045 $Y2=0.835
r182 35 37 5.30124 $w=2.48e-07 $l=1.15e-07 $layer=LI1_cond $X=5.045 $Y=0.75
+ $X2=5.045 $Y2=0.635
r183 33 71 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.92 $Y=0.835
+ $X2=5.045 $Y2=0.835
r184 33 34 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=4.92 $Y=0.835
+ $X2=4.24 $Y2=0.835
r185 32 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.155 $Y=0.75
+ $X2=4.24 $Y2=0.835
r186 31 32 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=4.155 $Y=0.58
+ $X2=4.155 $Y2=0.75
r187 27 30 39.8745 $w=2.48e-07 $l=8.65e-07 $layer=LI1_cond $X=2.435 $Y=0.455
+ $X2=3.3 $Y2=0.455
r188 25 31 7.14316 $w=2.5e-07 $l=1.62019e-07 $layer=LI1_cond $X=4.07 $Y=0.455
+ $X2=4.155 $Y2=0.58
r189 25 30 35.4952 $w=2.48e-07 $l=7.7e-07 $layer=LI1_cond $X=4.07 $Y=0.455
+ $X2=3.3 $Y2=0.455
r190 8 69 91 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_NDIFF $count=2 $X=10.175
+ $Y=0.37 $X2=10.33 $Y2=0.515
r191 7 61 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=8.75
+ $Y=0.37 $X2=8.89 $Y2=0.515
r192 6 55 91 $w=1.7e-07 $l=2.78209e-07 $layer=licon1_NDIFF $count=2 $X=7.815
+ $Y=0.37 $X2=8.03 $Y2=0.515
r193 5 49 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=6.915
+ $Y=0.37 $X2=7.055 $Y2=0.515
r194 4 43 182 $w=1.7e-07 $l=3.27605e-07 $layer=licon1_NDIFF $count=1 $X=5.885
+ $Y=0.37 $X2=6.025 $Y2=0.635
r195 3 37 182 $w=1.7e-07 $l=3.27605e-07 $layer=licon1_NDIFF $count=1 $X=4.865
+ $Y=0.37 $X2=5.005 $Y2=0.635
r196 2 30 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=3.155
+ $Y=0.37 $X2=3.3 $Y2=0.495
r197 1 27 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=2.295
+ $Y=0.37 $X2=2.435 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_HS__O311AI_4%VGND 1 2 3 4 5 6 7 24 28 32 36 40 42 44 46
+ 48 56 61 66 71 81 87 90 93 96 99 104 110 113
r137 112 113 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.8 $Y=0
+ $X2=10.8 $Y2=0
r138 109 110 11.3568 $w=8.73e-07 $l=1.1e-07 $layer=LI1_cond $X=9.885 $Y=0.352
+ $X2=9.995 $Y2=0.352
r139 106 109 0.627429 $w=8.73e-07 $l=4.5e-08 $layer=LI1_cond $X=9.84 $Y=0.352
+ $X2=9.885 $Y2=0.352
r140 106 107 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.84 $Y=0
+ $X2=9.84 $Y2=0
r141 103 107 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.36 $Y=0
+ $X2=9.84 $Y2=0
r142 102 106 6.69257 $w=8.73e-07 $l=4.8e-07 $layer=LI1_cond $X=9.36 $Y=0.352
+ $X2=9.84 $Y2=0.352
r143 102 104 12.6814 $w=8.73e-07 $l=2.05e-07 $layer=LI1_cond $X=9.36 $Y=0.352
+ $X2=9.155 $Y2=0.352
r144 102 103 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.36 $Y=0
+ $X2=9.36 $Y2=0
r145 99 100 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r146 96 97 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=0 $X2=7.44
+ $Y2=0
r147 93 94 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=0 $X2=6.48
+ $Y2=0
r148 87 88 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r149 85 113 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.32 $Y=0
+ $X2=10.8 $Y2=0
r150 85 107 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.32 $Y=0
+ $X2=9.84 $Y2=0
r151 84 110 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=10.32 $Y=0
+ $X2=9.995 $Y2=0
r152 84 85 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.32 $Y=0
+ $X2=10.32 $Y2=0
r153 81 112 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=10.595 $Y=0
+ $X2=10.817 $Y2=0
r154 81 84 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=10.595 $Y=0
+ $X2=10.32 $Y2=0
r155 80 103 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=0
+ $X2=9.36 $Y2=0
r156 80 100 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=0 $X2=8.4
+ $Y2=0
r157 79 104 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=8.88 $Y=0
+ $X2=9.155 $Y2=0
r158 79 80 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=0 $X2=8.88
+ $Y2=0
r159 77 99 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.545 $Y=0 $X2=8.42
+ $Y2=0
r160 77 79 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=8.545 $Y=0
+ $X2=8.88 $Y2=0
r161 75 100 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=0 $X2=8.4
+ $Y2=0
r162 75 97 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=0 $X2=7.44
+ $Y2=0
r163 74 75 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=0 $X2=7.92
+ $Y2=0
r164 72 96 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.65 $Y=0 $X2=7.485
+ $Y2=0
r165 72 74 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=7.65 $Y=0 $X2=7.92
+ $Y2=0
r166 71 99 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.295 $Y=0 $X2=8.42
+ $Y2=0
r167 71 74 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=8.295 $Y=0
+ $X2=7.92 $Y2=0
r168 70 97 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=0 $X2=7.44
+ $Y2=0
r169 70 94 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=0 $X2=6.48
+ $Y2=0
r170 69 70 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=0 $X2=6.96
+ $Y2=0
r171 67 93 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=6.71 $Y=0 $X2=6.54
+ $Y2=0
r172 67 69 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=6.71 $Y=0 $X2=6.96
+ $Y2=0
r173 66 96 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.32 $Y=0 $X2=7.485
+ $Y2=0
r174 66 69 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=7.32 $Y=0 $X2=6.96
+ $Y2=0
r175 65 94 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=0 $X2=6.48
+ $Y2=0
r176 64 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=0 $X2=6 $Y2=0
r177 62 90 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.68 $Y=0 $X2=5.515
+ $Y2=0
r178 62 64 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=5.68 $Y=0 $X2=6
+ $Y2=0
r179 61 93 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=6.37 $Y=0 $X2=6.54
+ $Y2=0
r180 61 64 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=6.37 $Y=0 $X2=6
+ $Y2=0
r181 60 88 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=4.56
+ $Y2=0
r182 59 60 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r183 57 87 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.74 $Y=0 $X2=4.575
+ $Y2=0
r184 57 59 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=4.74 $Y=0 $X2=5.04
+ $Y2=0
r185 56 90 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.35 $Y=0 $X2=5.515
+ $Y2=0
r186 56 59 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=5.35 $Y=0 $X2=5.04
+ $Y2=0
r187 55 88 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=4.56
+ $Y2=0
r188 54 55 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=4.08 $Y=0
+ $X2=4.08 $Y2=0
r189 51 55 1.07034 $w=4.9e-07 $l=3.84e-06 $layer=MET1_cond $X=0.24 $Y=0 $X2=4.08
+ $Y2=0
r190 50 54 250.524 $w=1.68e-07 $l=3.84e-06 $layer=LI1_cond $X=0.24 $Y=0 $X2=4.08
+ $Y2=0
r191 50 51 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=0.24 $Y=0
+ $X2=0.24 $Y2=0
r192 48 87 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.41 $Y=0 $X2=4.575
+ $Y2=0
r193 48 54 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=4.41 $Y=0 $X2=4.08
+ $Y2=0
r194 46 65 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=6
+ $Y2=0
r195 46 60 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=5.04
+ $Y2=0
r196 46 90 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r197 42 112 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=10.76 $Y=0.085
+ $X2=10.817 $Y2=0
r198 42 44 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=10.76 $Y=0.085
+ $X2=10.76 $Y2=0.515
r199 38 99 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=8.42 $Y=0.085
+ $X2=8.42 $Y2=0
r200 38 40 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=8.42 $Y=0.085
+ $X2=8.42 $Y2=0.515
r201 34 96 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.485 $Y=0.085
+ $X2=7.485 $Y2=0
r202 34 36 20.0804 $w=3.28e-07 $l=5.75e-07 $layer=LI1_cond $X=7.485 $Y=0.085
+ $X2=7.485 $Y2=0.66
r203 30 93 0.987631 $w=3.4e-07 $l=8.5e-08 $layer=LI1_cond $X=6.54 $Y=0.085
+ $X2=6.54 $Y2=0
r204 30 32 11.1855 $w=3.38e-07 $l=3.3e-07 $layer=LI1_cond $X=6.54 $Y=0.085
+ $X2=6.54 $Y2=0.415
r205 26 90 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.515 $Y=0.085
+ $X2=5.515 $Y2=0
r206 26 28 11.5244 $w=3.28e-07 $l=3.3e-07 $layer=LI1_cond $X=5.515 $Y=0.085
+ $X2=5.515 $Y2=0.415
r207 22 87 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.575 $Y=0.085
+ $X2=4.575 $Y2=0
r208 22 24 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=4.575 $Y=0.085
+ $X2=4.575 $Y2=0.495
r209 7 44 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=10.62
+ $Y=0.37 $X2=10.76 $Y2=0.515
r210 6 109 91 $w=1.7e-07 $l=8.22679e-07 $layer=licon1_NDIFF $count=2 $X=9.18
+ $Y=0.37 $X2=9.885 $Y2=0.625
r211 5 40 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=8.32
+ $Y=0.37 $X2=8.46 $Y2=0.515
r212 4 36 182 $w=1.7e-07 $l=3.53129e-07 $layer=licon1_NDIFF $count=1 $X=7.345
+ $Y=0.37 $X2=7.485 $Y2=0.66
r213 3 32 182 $w=1.7e-07 $l=2.46475e-07 $layer=licon1_NDIFF $count=1 $X=6.315
+ $Y=0.37 $X2=6.54 $Y2=0.415
r214 2 28 182 $w=1.7e-07 $l=2.41454e-07 $layer=licon1_NDIFF $count=1 $X=5.295
+ $Y=0.37 $X2=5.515 $Y2=0.415
r215 1 24 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=4.43
+ $Y=0.37 $X2=4.575 $Y2=0.495
.ends

