* NGSPICE file created from sky130_fd_sc_hs__o211ai_1.ext - technology: sky130A

.subckt sky130_fd_sc_hs__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
M1000 Y A2 a_116_368# VPB pshort w=1.12e+06u l=150000u
+  ad=9.688e+11p pd=6.21e+06u as=3.024e+11p ps=2.78e+06u
M1001 a_31_74# A2 VGND VNB nlowvt w=740000u l=150000u
+  ad=4.44e+11p pd=4.16e+06u as=2.59e+11p ps=2.18e+06u
M1002 a_311_74# B1 a_31_74# VNB nlowvt w=740000u l=150000u
+  ad=3.108e+11p pd=2.32e+06u as=0p ps=0u
M1003 Y C1 VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=7.224e+11p ps=5.77e+06u
M1004 VPWR B1 Y VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_116_368# A1 VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VGND A1 a_31_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 Y C1 a_311_74# VNB nlowvt w=740000u l=150000u
+  ad=4.588e+11p pd=2.72e+06u as=0p ps=0u
.ends

