* File: sky130_fd_sc_hs__o2bb2a_1.pxi.spice
* Created: Thu Aug 27 21:00:50 2020
* 
x_PM_SKY130_FD_SC_HS__O2BB2A_1%A_83_260# N_A_83_260#_M1007_s N_A_83_260#_M1001_d
+ N_A_83_260#_M1002_g N_A_83_260#_c_78_n N_A_83_260#_M1006_g N_A_83_260#_c_79_n
+ N_A_83_260#_c_80_n N_A_83_260#_c_81_n N_A_83_260#_c_82_n N_A_83_260#_c_83_n
+ N_A_83_260#_c_84_n N_A_83_260#_c_85_n N_A_83_260#_c_89_n N_A_83_260#_c_90_n
+ N_A_83_260#_c_86_n N_A_83_260#_c_91_n PM_SKY130_FD_SC_HS__O2BB2A_1%A_83_260#
x_PM_SKY130_FD_SC_HS__O2BB2A_1%A1_N N_A1_N_c_176_n N_A1_N_M1003_g N_A1_N_M1004_g
+ A1_N PM_SKY130_FD_SC_HS__O2BB2A_1%A1_N
x_PM_SKY130_FD_SC_HS__O2BB2A_1%A2_N N_A2_N_M1005_g N_A2_N_c_211_n N_A2_N_M1000_g
+ A2_N PM_SKY130_FD_SC_HS__O2BB2A_1%A2_N
x_PM_SKY130_FD_SC_HS__O2BB2A_1%A_233_384# N_A_233_384#_M1005_d
+ N_A_233_384#_M1003_d N_A_233_384#_c_241_n N_A_233_384#_c_242_n
+ N_A_233_384#_c_243_n N_A_233_384#_M1007_g N_A_233_384#_M1001_g
+ N_A_233_384#_c_244_n N_A_233_384#_c_245_n N_A_233_384#_c_249_n
+ N_A_233_384#_c_265_n N_A_233_384#_c_266_n N_A_233_384#_c_250_n
+ N_A_233_384#_c_246_n N_A_233_384#_c_247_n
+ PM_SKY130_FD_SC_HS__O2BB2A_1%A_233_384#
x_PM_SKY130_FD_SC_HS__O2BB2A_1%B2 N_B2_M1010_g N_B2_c_306_n N_B2_c_310_n
+ N_B2_M1008_g B2 B2 N_B2_c_308_n PM_SKY130_FD_SC_HS__O2BB2A_1%B2
x_PM_SKY130_FD_SC_HS__O2BB2A_1%B1 N_B1_M1011_g N_B1_M1009_g N_B1_c_348_n
+ N_B1_c_352_n B1 N_B1_c_350_n PM_SKY130_FD_SC_HS__O2BB2A_1%B1
x_PM_SKY130_FD_SC_HS__O2BB2A_1%X N_X_M1002_s N_X_M1006_s N_X_c_375_n N_X_c_376_n
+ X X X X N_X_c_377_n PM_SKY130_FD_SC_HS__O2BB2A_1%X
x_PM_SKY130_FD_SC_HS__O2BB2A_1%VPWR N_VPWR_M1006_d N_VPWR_M1000_d N_VPWR_M1011_d
+ N_VPWR_c_400_n N_VPWR_c_401_n N_VPWR_c_402_n VPWR N_VPWR_c_403_n
+ N_VPWR_c_404_n N_VPWR_c_405_n N_VPWR_c_406_n N_VPWR_c_407_n N_VPWR_c_399_n
+ PM_SKY130_FD_SC_HS__O2BB2A_1%VPWR
x_PM_SKY130_FD_SC_HS__O2BB2A_1%VGND N_VGND_M1002_d N_VGND_M1010_d N_VGND_c_446_n
+ N_VGND_c_447_n VGND N_VGND_c_448_n N_VGND_c_449_n N_VGND_c_450_n
+ N_VGND_c_451_n N_VGND_c_452_n N_VGND_c_453_n PM_SKY130_FD_SC_HS__O2BB2A_1%VGND
x_PM_SKY130_FD_SC_HS__O2BB2A_1%A_588_74# N_A_588_74#_M1007_d N_A_588_74#_M1009_d
+ N_A_588_74#_c_495_n N_A_588_74#_c_496_n N_A_588_74#_c_497_n
+ N_A_588_74#_c_498_n PM_SKY130_FD_SC_HS__O2BB2A_1%A_588_74#
cc_1 VNB N_A_83_260#_M1002_g 0.0293121f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=0.74
cc_2 VNB N_A_83_260#_c_78_n 0.0353881f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.765
cc_3 VNB N_A_83_260#_c_79_n 0.0138399f $X=-0.19 $Y=-0.245 $X2=1.29 $Y2=1.165
cc_4 VNB N_A_83_260#_c_80_n 0.0094333f $X=-0.19 $Y=-0.245 $X2=0.795 $Y2=1.165
cc_5 VNB N_A_83_260#_c_81_n 6.79008e-19 $X=-0.19 $Y=-0.245 $X2=1.375 $Y2=1.08
cc_6 VNB N_A_83_260#_c_82_n 0.0263861f $X=-0.19 $Y=-0.245 $X2=2.485 $Y2=0.34
cc_7 VNB N_A_83_260#_c_83_n 0.00270027f $X=-0.19 $Y=-0.245 $X2=1.46 $Y2=0.34
cc_8 VNB N_A_83_260#_c_84_n 0.00910354f $X=-0.19 $Y=-0.245 $X2=2.65 $Y2=0.495
cc_9 VNB N_A_83_260#_c_85_n 0.00580571f $X=-0.19 $Y=-0.245 $X2=2.73 $Y2=1.9
cc_10 VNB N_A_83_260#_c_86_n 0.00299619f $X=-0.19 $Y=-0.245 $X2=2.65 $Y2=0.92
cc_11 VNB N_A1_N_c_176_n 0.022695f $X=-0.19 $Y=-0.245 $X2=2.505 $Y2=0.37
cc_12 VNB N_A1_N_M1004_g 0.0235016f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB A1_N 0.0034197f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=0.74
cc_14 VNB N_A2_N_M1005_g 0.0297096f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A2_N_c_211_n 0.0208536f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB A2_N 0.00166191f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=0.74
cc_17 VNB N_A_233_384#_c_241_n 0.0277098f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.3
cc_18 VNB N_A_233_384#_c_242_n 0.0199158f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=0.74
cc_19 VNB N_A_233_384#_c_243_n 0.0185273f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=0.74
cc_20 VNB N_A_233_384#_c_244_n 0.00526231f $X=-0.19 $Y=-0.245 $X2=2.485 $Y2=0.34
cc_21 VNB N_A_233_384#_c_245_n 0.0221028f $X=-0.19 $Y=-0.245 $X2=1.46 $Y2=0.34
cc_22 VNB N_A_233_384#_c_246_n 0.0106619f $X=-0.19 $Y=-0.245 $X2=2.65 $Y2=0.92
cc_23 VNB N_A_233_384#_c_247_n 0.0320751f $X=-0.19 $Y=-0.245 $X2=3.155 $Y2=1.985
cc_24 VNB N_B2_M1010_g 0.0219963f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_B2_c_306_n 0.00895283f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB B2 0.0175784f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.765
cc_27 VNB N_B2_c_308_n 0.0288374f $X=-0.19 $Y=-0.245 $X2=0.795 $Y2=1.165
cc_28 VNB N_B1_M1009_g 0.0297108f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_B1_c_348_n 0.0121866f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB B1 0.00760591f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_31 VNB N_B1_c_350_n 0.0575527f $X=-0.19 $Y=-0.245 $X2=1.375 $Y2=1.08
cc_32 VNB N_X_c_375_n 0.0267746f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=0.74
cc_33 VNB N_X_c_376_n 0.0141322f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_34 VNB N_X_c_377_n 0.0247975f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.465
cc_35 VNB N_VPWR_c_399_n 0.183584f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_446_n 0.0101787f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=0.74
cc_37 VNB N_VGND_c_447_n 0.00963715f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_38 VNB N_VGND_c_448_n 0.0191572f $X=-0.19 $Y=-0.245 $X2=1.375 $Y2=1.08
cc_39 VNB N_VGND_c_449_n 0.0565361f $X=-0.19 $Y=-0.245 $X2=2.65 $Y2=0.495
cc_40 VNB N_VGND_c_450_n 0.018414f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.465
cc_41 VNB N_VGND_c_451_n 0.255724f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.465
cc_42 VNB N_VGND_c_452_n 0.00952121f $X=-0.19 $Y=-0.245 $X2=3.155 $Y2=2.065
cc_43 VNB N_VGND_c_453_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_588_74#_c_495_n 0.00210896f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=0.74
cc_45 VNB N_A_588_74#_c_496_n 0.0085555f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.765
cc_46 VNB N_A_588_74#_c_497_n 0.00180855f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_47 VNB N_A_588_74#_c_498_n 0.0208508f $X=-0.19 $Y=-0.245 $X2=0.795 $Y2=1.165
cc_48 VPB N_A_83_260#_c_78_n 0.0294431f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.765
cc_49 VPB N_A_83_260#_c_85_n 0.00223621f $X=-0.19 $Y=1.66 $X2=2.73 $Y2=1.9
cc_50 VPB N_A_83_260#_c_89_n 0.00116802f $X=-0.19 $Y=1.66 $X2=2.99 $Y2=1.985
cc_51 VPB N_A_83_260#_c_90_n 2.22016e-19 $X=-0.19 $Y=1.66 $X2=2.815 $Y2=1.985
cc_52 VPB N_A_83_260#_c_91_n 0.00500431f $X=-0.19 $Y=1.66 $X2=3.155 $Y2=2.065
cc_53 VPB N_A1_N_c_176_n 0.0338518f $X=-0.19 $Y=1.66 $X2=2.505 $Y2=0.37
cc_54 VPB A1_N 0.00391782f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=0.74
cc_55 VPB N_A2_N_c_211_n 0.0354887f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_56 VPB A2_N 0.0015854f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=0.74
cc_57 VPB N_A_233_384#_c_245_n 0.00497281f $X=-0.19 $Y=1.66 $X2=1.46 $Y2=0.34
cc_58 VPB N_A_233_384#_c_249_n 0.0253878f $X=-0.19 $Y=1.66 $X2=2.65 $Y2=0.425
cc_59 VPB N_A_233_384#_c_250_n 0.00316763f $X=-0.19 $Y=1.66 $X2=0.795 $Y2=1.165
cc_60 VPB N_A_233_384#_c_247_n 0.0167473f $X=-0.19 $Y=1.66 $X2=3.155 $Y2=1.985
cc_61 VPB N_B2_c_306_n 0.00548417f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_62 VPB N_B2_c_310_n 0.0227104f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.3
cc_63 VPB N_B1_c_348_n 0.00727927f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_64 VPB N_B1_c_352_n 0.0269593f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.765
cc_65 VPB X 0.0138461f $X=-0.19 $Y=1.66 $X2=1.29 $Y2=1.165
cc_66 VPB X 0.041687f $X=-0.19 $Y=1.66 $X2=2.65 $Y2=0.495
cc_67 VPB N_X_c_377_n 0.00776054f $X=-0.19 $Y=1.66 $X2=0.59 $Y2=1.465
cc_68 VPB N_VPWR_c_400_n 0.0173145f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.4
cc_69 VPB N_VPWR_c_401_n 0.0123504f $X=-0.19 $Y=1.66 $X2=2.485 $Y2=0.34
cc_70 VPB N_VPWR_c_402_n 0.0549689f $X=-0.19 $Y=1.66 $X2=2.65 $Y2=0.425
cc_71 VPB N_VPWR_c_403_n 0.0189171f $X=-0.19 $Y=1.66 $X2=2.99 $Y2=1.985
cc_72 VPB N_VPWR_c_404_n 0.031591f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=1.465
cc_73 VPB N_VPWR_c_405_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0.585 $Y2=1.465
cc_74 VPB N_VPWR_c_406_n 0.02253f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_75 VPB N_VPWR_c_407_n 0.0547228f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_76 VPB N_VPWR_c_399_n 0.0940406f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_77 N_A_83_260#_c_78_n N_A1_N_c_176_n 0.0446854f $X=0.505 $Y=1.765 $X2=-0.19
+ $Y2=-0.245
cc_78 N_A_83_260#_c_79_n N_A1_N_c_176_n 0.0048691f $X=1.29 $Y=1.165 $X2=-0.19
+ $Y2=-0.245
cc_79 N_A_83_260#_c_80_n N_A1_N_c_176_n 0.00237388f $X=0.795 $Y=1.165 $X2=-0.19
+ $Y2=-0.245
cc_80 N_A_83_260#_M1002_g N_A1_N_M1004_g 0.0102428f $X=0.505 $Y=0.74 $X2=0 $Y2=0
cc_81 N_A_83_260#_c_78_n N_A1_N_M1004_g 0.00148094f $X=0.505 $Y=1.765 $X2=0
+ $Y2=0
cc_82 N_A_83_260#_c_79_n N_A1_N_M1004_g 0.0149897f $X=1.29 $Y=1.165 $X2=0 $Y2=0
cc_83 N_A_83_260#_c_80_n N_A1_N_M1004_g 0.00200333f $X=0.795 $Y=1.165 $X2=0
+ $Y2=0
cc_84 N_A_83_260#_c_81_n N_A1_N_M1004_g 0.0026876f $X=1.375 $Y=1.08 $X2=0 $Y2=0
cc_85 N_A_83_260#_c_83_n N_A1_N_M1004_g 6.82792e-19 $X=1.46 $Y=0.34 $X2=0 $Y2=0
cc_86 N_A_83_260#_c_78_n A1_N 0.00107086f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_87 N_A_83_260#_c_79_n A1_N 0.0261759f $X=1.29 $Y=1.165 $X2=0 $Y2=0
cc_88 N_A_83_260#_c_80_n A1_N 0.0170081f $X=0.795 $Y=1.165 $X2=0 $Y2=0
cc_89 N_A_83_260#_c_79_n N_A2_N_M1005_g 0.00118344f $X=1.29 $Y=1.165 $X2=0 $Y2=0
cc_90 N_A_83_260#_c_81_n N_A2_N_M1005_g 0.00330892f $X=1.375 $Y=1.08 $X2=0 $Y2=0
cc_91 N_A_83_260#_c_82_n N_A2_N_M1005_g 0.0121086f $X=2.485 $Y=0.34 $X2=0 $Y2=0
cc_92 N_A_83_260#_c_85_n N_A_233_384#_c_241_n 0.00944143f $X=2.73 $Y=1.9 $X2=0
+ $Y2=0
cc_93 N_A_83_260#_c_86_n N_A_233_384#_c_241_n 0.00646708f $X=2.65 $Y=0.92 $X2=0
+ $Y2=0
cc_94 N_A_83_260#_c_82_n N_A_233_384#_c_242_n 0.00825806f $X=2.485 $Y=0.34 $X2=0
+ $Y2=0
cc_95 N_A_83_260#_c_82_n N_A_233_384#_c_243_n 0.00534381f $X=2.485 $Y=0.34 $X2=0
+ $Y2=0
cc_96 N_A_83_260#_c_84_n N_A_233_384#_c_243_n 0.00338973f $X=2.65 $Y=0.495 $X2=0
+ $Y2=0
cc_97 N_A_83_260#_c_85_n N_A_233_384#_c_243_n 0.00361776f $X=2.73 $Y=1.9 $X2=0
+ $Y2=0
cc_98 N_A_83_260#_c_86_n N_A_233_384#_c_243_n 0.00170336f $X=2.65 $Y=0.92 $X2=0
+ $Y2=0
cc_99 N_A_83_260#_c_85_n N_A_233_384#_c_244_n 0.00216975f $X=2.73 $Y=1.9 $X2=0
+ $Y2=0
cc_100 N_A_83_260#_c_85_n N_A_233_384#_c_245_n 0.0122328f $X=2.73 $Y=1.9 $X2=0
+ $Y2=0
cc_101 N_A_83_260#_c_85_n N_A_233_384#_c_249_n 0.00542694f $X=2.73 $Y=1.9 $X2=0
+ $Y2=0
cc_102 N_A_83_260#_c_89_n N_A_233_384#_c_249_n 0.0166184f $X=2.99 $Y=1.985 $X2=0
+ $Y2=0
cc_103 N_A_83_260#_c_90_n N_A_233_384#_c_249_n 0.00335121f $X=2.815 $Y=1.985
+ $X2=0 $Y2=0
cc_104 N_A_83_260#_c_91_n N_A_233_384#_c_249_n 0.00393325f $X=3.155 $Y=2.065
+ $X2=0 $Y2=0
cc_105 N_A_83_260#_c_90_n N_A_233_384#_c_265_n 0.00777294f $X=2.815 $Y=1.985
+ $X2=0 $Y2=0
cc_106 N_A_83_260#_c_82_n N_A_233_384#_c_266_n 0.0164516f $X=2.485 $Y=0.34 $X2=0
+ $Y2=0
cc_107 N_A_83_260#_c_84_n N_A_233_384#_c_266_n 0.0104187f $X=2.65 $Y=0.495 $X2=0
+ $Y2=0
cc_108 N_A_83_260#_c_85_n N_A_233_384#_c_250_n 0.035097f $X=2.73 $Y=1.9 $X2=0
+ $Y2=0
cc_109 N_A_83_260#_c_90_n N_A_233_384#_c_250_n 0.00310586f $X=2.815 $Y=1.985
+ $X2=0 $Y2=0
cc_110 N_A_83_260#_c_79_n N_A_233_384#_c_246_n 0.0132372f $X=1.29 $Y=1.165 $X2=0
+ $Y2=0
cc_111 N_A_83_260#_c_82_n N_A_233_384#_c_246_n 0.0132653f $X=2.485 $Y=0.34 $X2=0
+ $Y2=0
cc_112 N_A_83_260#_c_85_n N_A_233_384#_c_246_n 0.00900461f $X=2.73 $Y=1.9 $X2=0
+ $Y2=0
cc_113 N_A_83_260#_c_85_n N_A_233_384#_c_247_n 0.00379203f $X=2.73 $Y=1.9 $X2=0
+ $Y2=0
cc_114 N_A_83_260#_c_82_n N_B2_M1010_g 2.94862e-19 $X=2.485 $Y=0.34 $X2=0 $Y2=0
cc_115 N_A_83_260#_c_85_n N_B2_M1010_g 8.2968e-19 $X=2.73 $Y=1.9 $X2=0 $Y2=0
cc_116 N_A_83_260#_c_85_n N_B2_c_306_n 0.00160643f $X=2.73 $Y=1.9 $X2=0 $Y2=0
cc_117 N_A_83_260#_c_85_n N_B2_c_310_n 2.47254e-19 $X=2.73 $Y=1.9 $X2=0 $Y2=0
cc_118 N_A_83_260#_c_91_n N_B2_c_310_n 0.0173233f $X=3.155 $Y=2.065 $X2=0 $Y2=0
cc_119 N_A_83_260#_c_85_n B2 0.0244039f $X=2.73 $Y=1.9 $X2=0 $Y2=0
cc_120 N_A_83_260#_c_91_n B2 0.0150433f $X=3.155 $Y=2.065 $X2=0 $Y2=0
cc_121 N_A_83_260#_c_85_n N_B2_c_308_n 2.57511e-19 $X=2.73 $Y=1.9 $X2=0 $Y2=0
cc_122 N_A_83_260#_c_91_n N_B2_c_308_n 0.00268889f $X=3.155 $Y=2.065 $X2=0 $Y2=0
cc_123 N_A_83_260#_c_91_n N_B1_c_352_n 0.00249723f $X=3.155 $Y=2.065 $X2=0 $Y2=0
cc_124 N_A_83_260#_M1002_g N_X_c_375_n 0.0084877f $X=0.505 $Y=0.74 $X2=0 $Y2=0
cc_125 N_A_83_260#_M1002_g N_X_c_376_n 0.00427425f $X=0.505 $Y=0.74 $X2=0 $Y2=0
cc_126 N_A_83_260#_c_78_n N_X_c_376_n 5.00255e-19 $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_127 N_A_83_260#_c_80_n N_X_c_376_n 0.00515361f $X=0.795 $Y=1.165 $X2=0 $Y2=0
cc_128 N_A_83_260#_c_78_n X 0.00436092f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_129 N_A_83_260#_c_80_n X 0.001416f $X=0.795 $Y=1.165 $X2=0 $Y2=0
cc_130 N_A_83_260#_c_78_n X 0.0110489f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_131 N_A_83_260#_M1002_g N_X_c_377_n 0.00252147f $X=0.505 $Y=0.74 $X2=0 $Y2=0
cc_132 N_A_83_260#_c_78_n N_X_c_377_n 0.0124517f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_133 N_A_83_260#_c_80_n N_X_c_377_n 0.0307714f $X=0.795 $Y=1.165 $X2=0 $Y2=0
cc_134 N_A_83_260#_c_90_n N_VPWR_M1000_d 0.00371464f $X=2.815 $Y=1.985 $X2=0
+ $Y2=0
cc_135 N_A_83_260#_c_78_n N_VPWR_c_400_n 0.0134468f $X=0.505 $Y=1.765 $X2=0
+ $Y2=0
cc_136 N_A_83_260#_c_80_n N_VPWR_c_400_n 0.0090233f $X=0.795 $Y=1.165 $X2=0
+ $Y2=0
cc_137 N_A_83_260#_c_91_n N_VPWR_c_402_n 0.0254499f $X=3.155 $Y=2.065 $X2=0
+ $Y2=0
cc_138 N_A_83_260#_c_78_n N_VPWR_c_403_n 0.00445602f $X=0.505 $Y=1.765 $X2=0
+ $Y2=0
cc_139 N_A_83_260#_c_91_n N_VPWR_c_404_n 0.00709558f $X=3.155 $Y=2.065 $X2=0
+ $Y2=0
cc_140 N_A_83_260#_c_90_n N_VPWR_c_407_n 0.0055005f $X=2.815 $Y=1.985 $X2=0
+ $Y2=0
cc_141 N_A_83_260#_c_91_n N_VPWR_c_407_n 0.0146526f $X=3.155 $Y=2.065 $X2=0
+ $Y2=0
cc_142 N_A_83_260#_c_78_n N_VPWR_c_399_n 0.00865213f $X=0.505 $Y=1.765 $X2=0
+ $Y2=0
cc_143 N_A_83_260#_c_91_n N_VPWR_c_399_n 0.0105719f $X=3.155 $Y=2.065 $X2=0
+ $Y2=0
cc_144 N_A_83_260#_c_79_n N_VGND_M1002_d 0.00300823f $X=1.29 $Y=1.165 $X2=-0.19
+ $Y2=-0.245
cc_145 N_A_83_260#_c_80_n N_VGND_M1002_d 0.00199955f $X=0.795 $Y=1.165 $X2=-0.19
+ $Y2=-0.245
cc_146 N_A_83_260#_M1002_g N_VGND_c_446_n 0.00660116f $X=0.505 $Y=0.74 $X2=0
+ $Y2=0
cc_147 N_A_83_260#_c_78_n N_VGND_c_446_n 5.97302e-19 $X=0.505 $Y=1.765 $X2=0
+ $Y2=0
cc_148 N_A_83_260#_c_79_n N_VGND_c_446_n 0.0216234f $X=1.29 $Y=1.165 $X2=0 $Y2=0
cc_149 N_A_83_260#_c_80_n N_VGND_c_446_n 0.0140249f $X=0.795 $Y=1.165 $X2=0
+ $Y2=0
cc_150 N_A_83_260#_c_81_n N_VGND_c_446_n 0.0209803f $X=1.375 $Y=1.08 $X2=0 $Y2=0
cc_151 N_A_83_260#_c_83_n N_VGND_c_446_n 0.0151159f $X=1.46 $Y=0.34 $X2=0 $Y2=0
cc_152 N_A_83_260#_c_82_n N_VGND_c_447_n 0.00270678f $X=2.485 $Y=0.34 $X2=0
+ $Y2=0
cc_153 N_A_83_260#_M1002_g N_VGND_c_448_n 0.00434272f $X=0.505 $Y=0.74 $X2=0
+ $Y2=0
cc_154 N_A_83_260#_c_82_n N_VGND_c_449_n 0.08952f $X=2.485 $Y=0.34 $X2=0 $Y2=0
cc_155 N_A_83_260#_c_83_n N_VGND_c_449_n 0.0121867f $X=1.46 $Y=0.34 $X2=0 $Y2=0
cc_156 N_A_83_260#_M1002_g N_VGND_c_451_n 0.00828751f $X=0.505 $Y=0.74 $X2=0
+ $Y2=0
cc_157 N_A_83_260#_c_82_n N_VGND_c_451_n 0.0512413f $X=2.485 $Y=0.34 $X2=0 $Y2=0
cc_158 N_A_83_260#_c_83_n N_VGND_c_451_n 0.00660921f $X=1.46 $Y=0.34 $X2=0 $Y2=0
cc_159 N_A_83_260#_c_81_n A_253_94# 0.00212313f $X=1.375 $Y=1.08 $X2=-0.19
+ $Y2=-0.245
cc_160 N_A_83_260#_c_82_n N_A_588_74#_c_495_n 0.00453469f $X=2.485 $Y=0.34 $X2=0
+ $Y2=0
cc_161 N_A1_N_c_176_n N_A2_N_M1005_g 0.0230306f $X=1.09 $Y=1.845 $X2=0 $Y2=0
cc_162 N_A1_N_M1004_g N_A2_N_M1005_g 0.0466035f $X=1.19 $Y=0.79 $X2=0 $Y2=0
cc_163 A1_N N_A2_N_M1005_g 0.00229645f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_164 N_A1_N_c_176_n N_A2_N_c_211_n 0.0338808f $X=1.09 $Y=1.845 $X2=0 $Y2=0
cc_165 N_A1_N_c_176_n A2_N 4.10857e-19 $X=1.09 $Y=1.845 $X2=0 $Y2=0
cc_166 A1_N A2_N 0.0255486f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_167 N_A1_N_c_176_n N_A_233_384#_c_265_n 0.00490068f $X=1.09 $Y=1.845 $X2=0
+ $Y2=0
cc_168 A1_N N_A_233_384#_c_265_n 0.0111449f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_169 N_A1_N_M1004_g N_X_c_375_n 6.5955e-19 $X=1.19 $Y=0.79 $X2=0 $Y2=0
cc_170 N_A1_N_c_176_n X 7.55204e-19 $X=1.09 $Y=1.845 $X2=0 $Y2=0
cc_171 N_A1_N_c_176_n N_VPWR_c_400_n 0.0205877f $X=1.09 $Y=1.845 $X2=0 $Y2=0
cc_172 N_A1_N_c_176_n N_VPWR_c_406_n 0.00445514f $X=1.09 $Y=1.845 $X2=0 $Y2=0
cc_173 N_A1_N_c_176_n N_VPWR_c_407_n 0.00201773f $X=1.09 $Y=1.845 $X2=0 $Y2=0
cc_174 N_A1_N_c_176_n N_VPWR_c_399_n 0.00484898f $X=1.09 $Y=1.845 $X2=0 $Y2=0
cc_175 N_A1_N_M1004_g N_VGND_c_446_n 0.00998285f $X=1.19 $Y=0.79 $X2=0 $Y2=0
cc_176 N_A1_N_M1004_g N_VGND_c_449_n 0.00489033f $X=1.19 $Y=0.79 $X2=0 $Y2=0
cc_177 N_A1_N_M1004_g N_VGND_c_451_n 0.00500719f $X=1.19 $Y=0.79 $X2=0 $Y2=0
cc_178 N_A2_N_M1005_g N_A_233_384#_c_242_n 0.0105126f $X=1.58 $Y=0.79 $X2=0
+ $Y2=0
cc_179 N_A2_N_c_211_n N_A_233_384#_c_265_n 0.0265025f $X=1.595 $Y=1.845 $X2=0
+ $Y2=0
cc_180 A2_N N_A_233_384#_c_265_n 0.0230711f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_181 N_A2_N_M1005_g N_A_233_384#_c_266_n 0.00735949f $X=1.58 $Y=0.79 $X2=0
+ $Y2=0
cc_182 N_A2_N_M1005_g N_A_233_384#_c_250_n 9.76708e-19 $X=1.58 $Y=0.79 $X2=0
+ $Y2=0
cc_183 N_A2_N_c_211_n N_A_233_384#_c_250_n 0.00635053f $X=1.595 $Y=1.845 $X2=0
+ $Y2=0
cc_184 A2_N N_A_233_384#_c_250_n 0.0219371f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_185 N_A2_N_M1005_g N_A_233_384#_c_246_n 0.00474488f $X=1.58 $Y=0.79 $X2=0
+ $Y2=0
cc_186 N_A2_N_c_211_n N_A_233_384#_c_246_n 0.00126003f $X=1.595 $Y=1.845 $X2=0
+ $Y2=0
cc_187 A2_N N_A_233_384#_c_246_n 0.0153833f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_188 N_A2_N_c_211_n N_A_233_384#_c_247_n 0.0195426f $X=1.595 $Y=1.845 $X2=0
+ $Y2=0
cc_189 A2_N N_A_233_384#_c_247_n 0.00116124f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_190 N_A2_N_c_211_n N_VPWR_c_406_n 0.00399978f $X=1.595 $Y=1.845 $X2=0 $Y2=0
cc_191 N_A2_N_c_211_n N_VPWR_c_407_n 0.0125562f $X=1.595 $Y=1.845 $X2=0 $Y2=0
cc_192 N_A2_N_c_211_n N_VPWR_c_399_n 0.00436409f $X=1.595 $Y=1.845 $X2=0 $Y2=0
cc_193 N_A2_N_M1005_g N_VGND_c_446_n 2.05365e-19 $X=1.58 $Y=0.79 $X2=0 $Y2=0
cc_194 N_A2_N_M1005_g N_VGND_c_449_n 7.64118e-19 $X=1.58 $Y=0.79 $X2=0 $Y2=0
cc_195 N_A_233_384#_c_243_n N_B2_M1010_g 0.0137058f $X=2.865 $Y=1.09 $X2=0 $Y2=0
cc_196 N_A_233_384#_c_245_n N_B2_c_306_n 0.0085276f $X=2.872 $Y=1.75 $X2=0 $Y2=0
cc_197 N_A_233_384#_c_249_n N_B2_c_306_n 0.00356579f $X=2.872 $Y=1.845 $X2=0
+ $Y2=0
cc_198 N_A_233_384#_c_249_n N_B2_c_310_n 0.0195308f $X=2.872 $Y=1.845 $X2=0
+ $Y2=0
cc_199 N_A_233_384#_c_244_n B2 0.0026374f $X=2.865 $Y=1.165 $X2=0 $Y2=0
cc_200 N_A_233_384#_c_244_n N_B2_c_308_n 0.0166018f $X=2.865 $Y=1.165 $X2=0
+ $Y2=0
cc_201 N_A_233_384#_c_265_n N_VPWR_M1000_d 0.0315118f $X=2.05 $Y=2.115 $X2=0
+ $Y2=0
cc_202 N_A_233_384#_c_250_n N_VPWR_M1000_d 9.25727e-19 $X=2.215 $Y=1.95 $X2=0
+ $Y2=0
cc_203 N_A_233_384#_c_265_n N_VPWR_c_400_n 0.0233759f $X=2.05 $Y=2.115 $X2=0
+ $Y2=0
cc_204 N_A_233_384#_c_249_n N_VPWR_c_404_n 0.00399978f $X=2.872 $Y=1.845 $X2=0
+ $Y2=0
cc_205 N_A_233_384#_c_249_n N_VPWR_c_407_n 0.00914735f $X=2.872 $Y=1.845 $X2=0
+ $Y2=0
cc_206 N_A_233_384#_c_265_n N_VPWR_c_407_n 0.0580293f $X=2.05 $Y=2.115 $X2=0
+ $Y2=0
cc_207 N_A_233_384#_c_247_n N_VPWR_c_407_n 9.36276e-19 $X=2.215 $Y=1.255 $X2=0
+ $Y2=0
cc_208 N_A_233_384#_c_249_n N_VPWR_c_399_n 0.00436409f $X=2.872 $Y=1.845 $X2=0
+ $Y2=0
cc_209 N_A_233_384#_c_243_n N_VGND_c_449_n 0.00430908f $X=2.865 $Y=1.09 $X2=0
+ $Y2=0
cc_210 N_A_233_384#_c_243_n N_VGND_c_451_n 0.00821764f $X=2.865 $Y=1.09 $X2=0
+ $Y2=0
cc_211 N_A_233_384#_c_243_n N_A_588_74#_c_495_n 2.18574e-19 $X=2.865 $Y=1.09
+ $X2=0 $Y2=0
cc_212 N_B2_M1010_g N_B1_M1009_g 0.0217086f $X=3.295 $Y=0.69 $X2=0 $Y2=0
cc_213 N_B2_c_306_n N_B1_c_348_n 0.0126967f $X=3.39 $Y=1.755 $X2=0 $Y2=0
cc_214 N_B2_c_306_n N_B1_c_352_n 0.00533542f $X=3.39 $Y=1.755 $X2=0 $Y2=0
cc_215 N_B2_c_310_n N_B1_c_352_n 0.0530345f $X=3.39 $Y=1.845 $X2=0 $Y2=0
cc_216 B2 B1 0.0277564f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_217 N_B2_c_308_n B1 2.37823e-19 $X=3.345 $Y=1.345 $X2=0 $Y2=0
cc_218 B2 N_B1_c_350_n 0.00294527f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_219 N_B2_c_308_n N_B1_c_350_n 0.0175815f $X=3.345 $Y=1.345 $X2=0 $Y2=0
cc_220 N_B2_c_310_n N_VPWR_c_402_n 0.00384728f $X=3.39 $Y=1.845 $X2=0 $Y2=0
cc_221 N_B2_c_310_n N_VPWR_c_404_n 0.00545056f $X=3.39 $Y=1.845 $X2=0 $Y2=0
cc_222 N_B2_c_310_n N_VPWR_c_407_n 0.00511141f $X=3.39 $Y=1.845 $X2=0 $Y2=0
cc_223 N_B2_c_310_n N_VPWR_c_399_n 0.00533081f $X=3.39 $Y=1.845 $X2=0 $Y2=0
cc_224 N_B2_M1010_g N_VGND_c_447_n 0.00363829f $X=3.295 $Y=0.69 $X2=0 $Y2=0
cc_225 N_B2_M1010_g N_VGND_c_449_n 0.00434054f $X=3.295 $Y=0.69 $X2=0 $Y2=0
cc_226 N_B2_M1010_g N_VGND_c_451_n 0.00445726f $X=3.295 $Y=0.69 $X2=0 $Y2=0
cc_227 N_B2_M1010_g N_A_588_74#_c_495_n 0.00711952f $X=3.295 $Y=0.69 $X2=0 $Y2=0
cc_228 N_B2_M1010_g N_A_588_74#_c_496_n 0.0090049f $X=3.295 $Y=0.69 $X2=0 $Y2=0
cc_229 B2 N_A_588_74#_c_496_n 0.0323411f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_230 N_B2_c_308_n N_A_588_74#_c_496_n 0.00344071f $X=3.345 $Y=1.345 $X2=0
+ $Y2=0
cc_231 N_B2_M1010_g N_A_588_74#_c_497_n 7.17385e-19 $X=3.295 $Y=0.69 $X2=0 $Y2=0
cc_232 B2 N_A_588_74#_c_497_n 0.0178517f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_233 N_B1_c_352_n N_VPWR_c_402_n 0.0242829f $X=3.817 $Y=1.845 $X2=0 $Y2=0
cc_234 B1 N_VPWR_c_402_n 0.0142647f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_235 N_B1_c_350_n N_VPWR_c_402_n 0.00211705f $X=4.05 $Y=1.345 $X2=0 $Y2=0
cc_236 N_B1_c_352_n N_VPWR_c_404_n 0.00492531f $X=3.817 $Y=1.845 $X2=0 $Y2=0
cc_237 N_B1_c_352_n N_VPWR_c_399_n 0.00483326f $X=3.817 $Y=1.845 $X2=0 $Y2=0
cc_238 N_B1_M1009_g N_VGND_c_447_n 0.00330983f $X=3.825 $Y=0.69 $X2=0 $Y2=0
cc_239 N_B1_M1009_g N_VGND_c_450_n 0.00461464f $X=3.825 $Y=0.69 $X2=0 $Y2=0
cc_240 N_B1_M1009_g N_VGND_c_451_n 0.00467092f $X=3.825 $Y=0.69 $X2=0 $Y2=0
cc_241 N_B1_M1009_g N_A_588_74#_c_495_n 6.85083e-19 $X=3.825 $Y=0.69 $X2=0 $Y2=0
cc_242 N_B1_M1009_g N_A_588_74#_c_496_n 0.0144732f $X=3.825 $Y=0.69 $X2=0 $Y2=0
cc_243 B1 N_A_588_74#_c_496_n 0.0237154f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_244 N_B1_c_350_n N_A_588_74#_c_496_n 0.00196043f $X=4.05 $Y=1.345 $X2=0 $Y2=0
cc_245 N_B1_M1009_g N_A_588_74#_c_498_n 6.81345e-19 $X=3.825 $Y=0.69 $X2=0 $Y2=0
cc_246 X N_VPWR_c_400_n 0.0399187f $X=0.155 $Y=1.95 $X2=0 $Y2=0
cc_247 X N_VPWR_c_403_n 0.0159324f $X=0.24 $Y=2.035 $X2=0 $Y2=0
cc_248 X N_VPWR_c_399_n 0.0131546f $X=0.24 $Y=2.035 $X2=0 $Y2=0
cc_249 N_X_c_375_n N_VGND_c_446_n 0.0222242f $X=0.29 $Y=0.515 $X2=0 $Y2=0
cc_250 N_X_c_375_n N_VGND_c_448_n 0.0163488f $X=0.29 $Y=0.515 $X2=0 $Y2=0
cc_251 N_X_c_375_n N_VGND_c_451_n 0.0134757f $X=0.29 $Y=0.515 $X2=0 $Y2=0
cc_252 N_VGND_c_447_n N_A_588_74#_c_495_n 0.0130732f $X=3.58 $Y=0.55 $X2=0 $Y2=0
cc_253 N_VGND_c_449_n N_A_588_74#_c_495_n 0.0114427f $X=3.415 $Y=0 $X2=0 $Y2=0
cc_254 N_VGND_c_451_n N_A_588_74#_c_495_n 0.00909435f $X=4.08 $Y=0 $X2=0 $Y2=0
cc_255 N_VGND_M1010_d N_A_588_74#_c_496_n 0.00561113f $X=3.37 $Y=0.37 $X2=0
+ $Y2=0
cc_256 N_VGND_c_447_n N_A_588_74#_c_496_n 0.0211672f $X=3.58 $Y=0.55 $X2=0 $Y2=0
cc_257 N_VGND_c_451_n N_A_588_74#_c_496_n 0.0122262f $X=4.08 $Y=0 $X2=0 $Y2=0
cc_258 N_VGND_c_447_n N_A_588_74#_c_498_n 0.00203724f $X=3.58 $Y=0.55 $X2=0
+ $Y2=0
cc_259 N_VGND_c_450_n N_A_588_74#_c_498_n 0.0115155f $X=4.08 $Y=0 $X2=0 $Y2=0
cc_260 N_VGND_c_451_n N_A_588_74#_c_498_n 0.00920958f $X=4.08 $Y=0 $X2=0 $Y2=0
