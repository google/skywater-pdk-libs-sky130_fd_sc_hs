* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hs__and3b_2 A_N B C VGND VNB VPB VPWR X
X0 a_454_74# C VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X1 a_284_368# C VPWR VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=150000u
X2 X a_284_368# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X3 VPWR a_284_368# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X4 a_284_368# a_27_88# VPWR VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=150000u
X5 X a_284_368# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X6 VPWR B a_284_368# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=150000u
X7 VGND a_284_368# X VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X8 a_376_74# B a_454_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X9 a_27_88# A_N VPWR VPB sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X10 a_27_88# A_N VGND VNB sky130_fd_pr__nfet_01v8_lvt w=550000u l=150000u
X11 a_284_368# a_27_88# a_376_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
.ends
