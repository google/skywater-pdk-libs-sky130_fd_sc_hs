* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hs__or4_2 A B C D VGND VNB VPB VPWR X
X0 a_258_392# B a_342_392# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=150000u
X1 X a_85_392# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X2 a_85_392# C VGND VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X3 VGND a_85_392# X VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X4 a_85_392# D a_174_392# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=150000u
X5 a_174_392# C a_258_392# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=150000u
X6 X a_85_392# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X7 VGND D a_85_392# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X8 VPWR a_85_392# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X9 VGND B a_85_392# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X10 a_342_392# A VPWR VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=150000u
X11 a_85_392# A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
.ends
