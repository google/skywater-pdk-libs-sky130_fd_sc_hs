* File: sky130_fd_sc_hs__o2bb2a_1.pex.spice
* Created: Tue Sep  1 20:16:41 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HS__O2BB2A_1%A_83_260# 1 2 9 11 13 14 15 17 18 19 23 25
+ 26 27 34 36
c99 26 0 1.80776e-19 $X=2.99 $Y=1.985
r100 32 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.59
+ $Y=1.465 $X2=0.59 $Y2=1.465
r101 26 36 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.99 $Y=1.985
+ $X2=3.155 $Y2=1.985
r102 26 27 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=2.99 $Y=1.985
+ $X2=2.815 $Y2=1.985
r103 25 27 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.73 $Y=1.9
+ $X2=2.815 $Y2=1.985
r104 25 34 63.9358 $w=1.68e-07 $l=9.8e-07 $layer=LI1_cond $X=2.73 $Y=1.9
+ $X2=2.73 $Y2=0.92
r105 21 34 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=2.65 $Y=0.755
+ $X2=2.65 $Y2=0.92
r106 21 23 9.07985 $w=3.28e-07 $l=2.6e-07 $layer=LI1_cond $X=2.65 $Y=0.755
+ $X2=2.65 $Y2=0.495
r107 20 23 2.44458 $w=3.28e-07 $l=7e-08 $layer=LI1_cond $X=2.65 $Y=0.425
+ $X2=2.65 $Y2=0.495
r108 18 20 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.485 $Y=0.34
+ $X2=2.65 $Y2=0.425
r109 18 19 66.8717 $w=1.68e-07 $l=1.025e-06 $layer=LI1_cond $X=2.485 $Y=0.34
+ $X2=1.46 $Y2=0.34
r110 16 19 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.375 $Y=0.425
+ $X2=1.46 $Y2=0.34
r111 16 17 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=1.375 $Y=0.425
+ $X2=1.375 $Y2=1.08
r112 15 32 12.6207 $w=2.9e-07 $l=3.81445e-07 $layer=LI1_cond $X=0.795 $Y=1.165
+ $X2=0.61 $Y2=1.465
r113 14 17 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.29 $Y=1.165
+ $X2=1.375 $Y2=1.08
r114 14 15 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=1.29 $Y=1.165
+ $X2=0.795 $Y2=1.165
r115 11 33 60.7998 $w=2.93e-07 $l=3.37639e-07 $layer=POLY_cond $X=0.505 $Y=1.765
+ $X2=0.585 $Y2=1.465
r116 11 13 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.505 $Y=1.765
+ $X2=0.505 $Y2=2.4
r117 7 33 38.5916 $w=2.93e-07 $l=2.0106e-07 $layer=POLY_cond $X=0.505 $Y=1.3
+ $X2=0.585 $Y2=1.465
r118 7 9 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=0.505 $Y=1.3
+ $X2=0.505 $Y2=0.74
r119 2 36 300 $w=1.7e-07 $l=2.62678e-07 $layer=licon1_PDIFF $count=2 $X=2.955
+ $Y=1.92 $X2=3.155 $Y2=2.065
r120 1 23 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=2.505
+ $Y=0.37 $X2=2.65 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_HS__O2BB2A_1%A1_N 1 3 6 8
c34 6 0 3.57487e-19 $X=1.19 $Y=0.79
r35 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.13
+ $Y=1.545 $X2=1.13 $Y2=1.545
r36 8 12 4.4908 $w=3.26e-07 $l=1.2e-07 $layer=LI1_cond $X=1.14 $Y=1.665 $X2=1.14
+ $Y2=1.545
r37 4 11 43.6282 $w=2.89e-07 $l=2.22991e-07 $layer=POLY_cond $X=1.19 $Y=1.35
+ $X2=1.13 $Y2=1.545
r38 4 6 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=1.19 $Y=1.35 $X2=1.19
+ $Y2=0.79
r39 1 11 61.1403 $w=2.89e-07 $l=3.19374e-07 $layer=POLY_cond $X=1.09 $Y=1.845
+ $X2=1.13 $Y2=1.545
r40 1 3 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=1.09 $Y=1.845 $X2=1.09
+ $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_HS__O2BB2A_1%A2_N 3 5 7 8
r31 8 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.67
+ $Y=1.595 $X2=1.67 $Y2=1.595
r32 5 11 52.2586 $w=2.99e-07 $l=2.85044e-07 $layer=POLY_cond $X=1.595 $Y=1.845
+ $X2=1.67 $Y2=1.595
r33 5 7 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=1.595 $Y=1.845
+ $X2=1.595 $Y2=2.34
r34 1 11 38.5562 $w=2.99e-07 $l=2.05122e-07 $layer=POLY_cond $X=1.58 $Y=1.43
+ $X2=1.67 $Y2=1.595
r35 1 3 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=1.58 $Y=1.43 $X2=1.58
+ $Y2=0.79
.ends

.subckt PM_SKY130_FD_SC_HS__O2BB2A_1%A_233_384# 1 2 7 8 9 11 16 18 19 20 21 27
+ 30 34 35
c64 34 0 1.64798e-19 $X=2.215 $Y=1.255
c65 27 0 1.63523e-19 $X=1.795 $Y=0.86
r66 34 35 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.215
+ $Y=1.255 $X2=2.215 $Y2=1.255
r67 30 34 24.0965 $w=3.28e-07 $l=6.9e-07 $layer=LI1_cond $X=2.215 $Y=1.95
+ $X2=2.215 $Y2=1.26
r68 25 34 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=1.755 $Y=1.175
+ $X2=2.215 $Y2=1.175
r69 25 27 10.6025 $w=2.48e-07 $l=2.3e-07 $layer=LI1_cond $X=1.755 $Y=1.09
+ $X2=1.755 $Y2=0.86
r70 21 30 6.81649 $w=3.3e-07 $l=2.33345e-07 $layer=LI1_cond $X=2.05 $Y=2.115
+ $X2=2.215 $Y2=1.95
r71 21 23 25.668 $w=3.28e-07 $l=7.35e-07 $layer=LI1_cond $X=2.05 $Y=2.115
+ $X2=1.315 $Y2=2.115
r72 19 20 41.3838 $w=1.65e-07 $l=9.5e-08 $layer=POLY_cond $X=2.872 $Y=1.75
+ $X2=2.872 $Y2=1.845
r73 17 35 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=2.215 $Y=1.24
+ $X2=2.215 $Y2=1.255
r74 16 20 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=2.88 $Y=2.34
+ $X2=2.88 $Y2=1.845
r75 12 18 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.865 $Y=1.24
+ $X2=2.865 $Y2=1.165
r76 12 19 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=2.865 $Y=1.24
+ $X2=2.865 $Y2=1.75
r77 9 18 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.865 $Y=1.09
+ $X2=2.865 $Y2=1.165
r78 9 11 128.533 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=2.865 $Y=1.09 $X2=2.865
+ $Y2=0.69
r79 8 17 32.1775 $w=1.5e-07 $l=1.98997e-07 $layer=POLY_cond $X=2.38 $Y=1.165
+ $X2=2.215 $Y2=1.24
r80 7 18 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.79 $Y=1.165
+ $X2=2.865 $Y2=1.165
r81 7 8 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=2.79 $Y=1.165 $X2=2.38
+ $Y2=1.165
r82 2 23 600 $w=1.7e-07 $l=2.59374e-07 $layer=licon1_PDIFF $count=1 $X=1.165
+ $Y=1.92 $X2=1.315 $Y2=2.115
r83 1 27 182 $w=1.7e-07 $l=4.54643e-07 $layer=licon1_NDIFF $count=1 $X=1.655
+ $Y=0.47 $X2=1.795 $Y2=0.86
.ends

.subckt PM_SKY130_FD_SC_HS__O2BB2A_1%B2 3 6 7 9 10 11 15
r42 15 18 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.345 $Y=1.345
+ $X2=3.345 $Y2=1.51
r43 15 17 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.345 $Y=1.345
+ $X2=3.345 $Y2=1.18
r44 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.345
+ $Y=1.345 $X2=3.345 $Y2=1.345
r45 11 16 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=3.6 $Y=1.345
+ $X2=3.345 $Y2=1.345
r46 10 16 7.85757 $w=3.28e-07 $l=2.25e-07 $layer=LI1_cond $X=3.12 $Y=1.345
+ $X2=3.345 $Y2=1.345
r47 7 9 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=3.39 $Y=1.845
+ $X2=3.39 $Y2=2.42
r48 6 7 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=3.39 $Y=1.755 $X2=3.39
+ $Y2=1.845
r49 6 18 95.2339 $w=1.8e-07 $l=2.45e-07 $layer=POLY_cond $X=3.39 $Y=1.755
+ $X2=3.39 $Y2=1.51
r50 3 17 251.255 $w=1.5e-07 $l=4.9e-07 $layer=POLY_cond $X=3.295 $Y=0.69
+ $X2=3.295 $Y2=1.18
.ends

.subckt PM_SKY130_FD_SC_HS__O2BB2A_1%B1 3 6 10 11 12 17
r28 14 17 39.3438 $w=3.3e-07 $l=2.25e-07 $layer=POLY_cond $X=3.825 $Y=1.345
+ $X2=4.05 $Y2=1.345
r29 12 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.05
+ $Y=1.345 $X2=4.05 $Y2=1.345
r30 10 11 41.3838 $w=1.65e-07 $l=9.5e-08 $layer=POLY_cond $X=3.817 $Y=1.75
+ $X2=3.817 $Y2=1.845
r31 8 14 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.825 $Y=1.51
+ $X2=3.825 $Y2=1.345
r32 8 10 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=3.825 $Y=1.51
+ $X2=3.825 $Y2=1.75
r33 4 14 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.825 $Y=1.18
+ $X2=3.825 $Y2=1.345
r34 4 6 251.255 $w=1.5e-07 $l=4.9e-07 $layer=POLY_cond $X=3.825 $Y=1.18
+ $X2=3.825 $Y2=0.69
r35 3 11 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=3.81 $Y=2.42
+ $X2=3.81 $Y2=1.845
.ends

.subckt PM_SKY130_FD_SC_HS__O2BB2A_1%X 1 2 9 13 14 15 16 23 32
c24 13 0 2.91662e-20 $X=0.27 $Y=1.13
r25 21 23 1.12043 $w=3.58e-07 $l=3.5e-08 $layer=LI1_cond $X=0.265 $Y=2 $X2=0.265
+ $Y2=2.035
r26 15 16 11.8446 $w=3.58e-07 $l=3.7e-07 $layer=LI1_cond $X=0.265 $Y=2.405
+ $X2=0.265 $Y2=2.775
r27 14 21 0.800308 $w=3.58e-07 $l=2.5e-08 $layer=LI1_cond $X=0.265 $Y=1.975
+ $X2=0.265 $Y2=2
r28 14 32 8.1909 $w=3.58e-07 $l=1.55e-07 $layer=LI1_cond $X=0.265 $Y=1.975
+ $X2=0.265 $Y2=1.82
r29 14 15 11.0442 $w=3.58e-07 $l=3.45e-07 $layer=LI1_cond $X=0.265 $Y=2.06
+ $X2=0.265 $Y2=2.405
r30 14 23 0.800308 $w=3.58e-07 $l=2.5e-08 $layer=LI1_cond $X=0.265 $Y=2.06
+ $X2=0.265 $Y2=2.035
r31 13 32 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=0.17 $Y=1.13 $X2=0.17
+ $Y2=1.82
r32 7 13 9.16175 $w=3.68e-07 $l=1.85e-07 $layer=LI1_cond $X=0.27 $Y=0.945
+ $X2=0.27 $Y2=1.13
r33 7 9 13.3933 $w=3.68e-07 $l=4.3e-07 $layer=LI1_cond $X=0.27 $Y=0.945 $X2=0.27
+ $Y2=0.515
r34 2 14 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=1.985
r35 2 16 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.815
r36 1 9 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.145
+ $Y=0.37 $X2=0.29 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__O2BB2A_1%VPWR 1 2 3 12 18 20 24 26 31 37 42 50 53
c47 50 0 1.80776e-19 $X=2.82 $Y=2.932
r48 52 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r49 49 50 12.652 $w=9.63e-07 $l=1.65e-07 $layer=LI1_cond $X=2.655 $Y=2.932
+ $X2=2.82 $Y2=2.932
r50 46 49 0.189637 $w=9.63e-07 $l=1.5e-08 $layer=LI1_cond $X=2.64 $Y=2.932
+ $X2=2.655 $Y2=2.932
r51 46 47 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r52 44 46 10.3668 $w=9.63e-07 $l=8.2e-07 $layer=LI1_cond $X=1.82 $Y=2.932
+ $X2=2.64 $Y2=2.932
r53 40 44 1.76995 $w=9.63e-07 $l=1.4e-07 $layer=LI1_cond $X=1.68 $Y=2.932
+ $X2=1.82 $Y2=2.932
r54 40 42 10.8821 $w=9.63e-07 $l=2.5e-08 $layer=LI1_cond $X=1.68 $Y=2.932
+ $X2=1.655 $Y2=2.932
r55 40 41 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r56 38 41 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.68 $Y2=3.33
r57 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r58 35 53 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.08 $Y2=3.33
r59 35 47 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=2.64 $Y2=3.33
r60 34 50 50.8877 $w=1.68e-07 $l=7.8e-07 $layer=LI1_cond $X=3.6 $Y=3.33 $X2=2.82
+ $Y2=3.33
r61 34 35 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r62 31 52 4.72267 $w=1.7e-07 $l=2.25e-07 $layer=LI1_cond $X=3.87 $Y=3.33
+ $X2=4.095 $Y2=3.33
r63 31 34 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=3.87 $Y=3.33 $X2=3.6
+ $Y2=3.33
r64 29 38 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r65 28 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r66 26 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.615 $Y=3.33
+ $X2=0.78 $Y2=3.33
r67 26 28 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=0.615 $Y=3.33
+ $X2=0.24 $Y2=3.33
r68 24 47 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r69 24 41 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.68 $Y2=3.33
r70 20 23 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=4.035 $Y=2.065
+ $X2=4.035 $Y2=2.775
r71 18 52 3.0435 $w=3.3e-07 $l=1.11018e-07 $layer=LI1_cond $X=4.035 $Y=3.245
+ $X2=4.095 $Y2=3.33
r72 18 23 16.4136 $w=3.28e-07 $l=4.7e-07 $layer=LI1_cond $X=4.035 $Y=3.245
+ $X2=4.035 $Y2=2.775
r73 17 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.945 $Y=3.33
+ $X2=0.78 $Y2=3.33
r74 17 42 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=0.945 $Y=3.33
+ $X2=1.655 $Y2=3.33
r75 12 15 26.8903 $w=3.28e-07 $l=7.7e-07 $layer=LI1_cond $X=0.78 $Y=2.045
+ $X2=0.78 $Y2=2.815
r76 10 37 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.78 $Y=3.245
+ $X2=0.78 $Y2=3.33
r77 10 15 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=0.78 $Y=3.245
+ $X2=0.78 $Y2=2.815
r78 3 23 400 $w=1.7e-07 $l=9.26971e-07 $layer=licon1_PDIFF $count=1 $X=3.885
+ $Y=1.92 $X2=4.035 $Y2=2.775
r79 3 20 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=3.885
+ $Y=1.92 $X2=4.035 $Y2=2.065
r80 2 49 400 $w=1.7e-07 $l=1.27292e-06 $layer=licon1_PDIFF $count=1 $X=1.67
+ $Y=1.92 $X2=2.655 $Y2=2.58
r81 2 44 400 $w=1.7e-07 $l=7.31163e-07 $layer=licon1_PDIFF $count=1 $X=1.67
+ $Y=1.92 $X2=1.82 $Y2=2.58
r82 1 15 600 $w=1.7e-07 $l=1.07034e-06 $layer=licon1_PDIFF $count=1 $X=0.58
+ $Y=1.84 $X2=0.78 $Y2=2.815
r83 1 12 300 $w=1.7e-07 $l=2.88141e-07 $layer=licon1_PDIFF $count=2 $X=0.58
+ $Y=1.84 $X2=0.78 $Y2=2.045
.ends

.subckt PM_SKY130_FD_SC_HS__O2BB2A_1%VGND 1 2 9 13 15 17 22 32 33 36 39
r48 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r49 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r50 33 40 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=3.6
+ $Y2=0
r51 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r52 30 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.745 $Y=0 $X2=3.58
+ $Y2=0
r53 30 32 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=3.745 $Y=0 $X2=4.08
+ $Y2=0
r54 29 40 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=3.6
+ $Y2=0
r55 28 29 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r56 26 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r57 25 28 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=1.2 $Y=0 $X2=3.12
+ $Y2=0
r58 25 26 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r59 23 36 11.2236 $w=1.7e-07 $l=2.48e-07 $layer=LI1_cond $X=1.12 $Y=0 $X2=0.872
+ $Y2=0
r60 23 25 5.21925 $w=1.68e-07 $l=8e-08 $layer=LI1_cond $X=1.12 $Y=0 $X2=1.2
+ $Y2=0
r61 22 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.415 $Y=0 $X2=3.58
+ $Y2=0
r62 22 28 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=3.415 $Y=0 $X2=3.12
+ $Y2=0
r63 20 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r64 19 20 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r65 17 36 11.2236 $w=1.7e-07 $l=2.47e-07 $layer=LI1_cond $X=0.625 $Y=0 $X2=0.872
+ $Y2=0
r66 17 19 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=0.625 $Y=0 $X2=0.24
+ $Y2=0
r67 15 29 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=3.12
+ $Y2=0
r68 15 26 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.2
+ $Y2=0
r69 11 39 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.58 $Y=0.085
+ $X2=3.58 $Y2=0
r70 11 13 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=3.58 $Y=0.085
+ $X2=3.58 $Y2=0.55
r71 7 36 2.04857 $w=4.95e-07 $l=8.5e-08 $layer=LI1_cond $X=0.872 $Y=0.085
+ $X2=0.872 $Y2=0
r72 7 9 9.90691 $w=4.93e-07 $l=4.1e-07 $layer=LI1_cond $X=0.872 $Y=0.085
+ $X2=0.872 $Y2=0.495
r73 2 13 182 $w=1.7e-07 $l=2.86182e-07 $layer=licon1_NDIFF $count=1 $X=3.37
+ $Y=0.37 $X2=3.58 $Y2=0.55
r74 1 9 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=0.58
+ $Y=0.37 $X2=0.72 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_HS__O2BB2A_1%A_588_74# 1 2 9 11 12 15
r26 13 15 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=4.08 $Y=0.84
+ $X2=4.08 $Y2=0.505
r27 11 13 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=3.955 $Y=0.925
+ $X2=4.08 $Y2=0.84
r28 11 12 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=3.955 $Y=0.925
+ $X2=3.245 $Y2=0.925
r29 7 12 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=3.12 $Y=0.84
+ $X2=3.245 $Y2=0.925
r30 7 9 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=3.12 $Y=0.84 $X2=3.12
+ $Y2=0.505
r31 2 15 91 $w=1.7e-07 $l=1.96214e-07 $layer=licon1_NDIFF $count=2 $X=3.9
+ $Y=0.37 $X2=4.04 $Y2=0.505
r32 1 9 91 $w=1.7e-07 $l=1.96214e-07 $layer=licon1_NDIFF $count=2 $X=2.94
+ $Y=0.37 $X2=3.08 $Y2=0.505
.ends

