* File: sky130_fd_sc_hs__dfrtn_1.spice
* Created: Thu Aug 27 20:38:30 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hs__dfrtn_1.pex.spice"
.subckt sky130_fd_sc_hs__dfrtn_1  VNB VPB D RESET_B CLK_N VPWR Q VGND
* 
* VGND	VGND
* Q	Q
* VPWR	VPWR
* CLK_N	CLK_N
* RESET_B	RESET_B
* D	D
* VPB	VPB
* VNB	VNB
MM1029 A_120_74# N_D_M1029_g N_A_33_74#_M1029_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.0504 AS=0.1197 PD=0.66 PS=1.41 NRD=18.564 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1024 N_VGND_M1024_d N_RESET_B_M1024_g A_120_74# VNB NLOWVT L=0.15 W=0.42
+ AD=0.0877655 AS=0.0504 PD=0.796552 PS=0.66 NRD=22.848 NRS=18.564 M=1 R=2.8
+ SA=75000.6 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1027 N_A_300_74#_M1027_d N_CLK_N_M1027_g N_VGND_M1024_d VNB NLOWVT L=0.15
+ W=0.74 AD=0.2035 AS=0.154634 PD=2.03 PS=1.40345 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.7 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1010 N_A_507_368#_M1010_d N_A_300_74#_M1010_g N_VGND_M1010_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.2596 AS=0.3593 PD=2.24 PS=2.88 NRD=11.34 NRS=69.816 M=1 R=4.93333
+ SA=75000.3 SB=75000.3 A=0.111 P=1.78 MULT=1
MM1013 N_A_714_127#_M1013_d N_A_507_368#_M1013_g N_A_33_74#_M1013_s VNB NLOWVT
+ L=0.15 W=0.42 AD=0.1113 AS=0.1113 PD=0.95 PS=1.37 NRD=71.424 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75005.4 A=0.063 P=1.14 MULT=1
MM1030 A_850_127# N_A_300_74#_M1030_g N_A_714_127#_M1013_d VNB NLOWVT L=0.15
+ W=0.42 AD=0.0441 AS=0.1113 PD=0.63 PS=0.95 NRD=14.28 NRS=0 M=1 R=2.8
+ SA=75000.9 SB=75004.8 A=0.063 P=1.14 MULT=1
MM1026 A_922_127# N_A_856_304#_M1026_g A_850_127# VNB NLOWVT L=0.15 W=0.42
+ AD=0.0441 AS=0.0441 PD=0.63 PS=0.63 NRD=14.28 NRS=14.28 M=1 R=2.8 SA=75001.2
+ SB=75004.4 A=0.063 P=1.14 MULT=1
MM1015 N_VGND_M1015_d N_RESET_B_M1015_g A_922_127# VNB NLOWVT L=0.15 W=0.42
+ AD=0.174028 AS=0.0441 PD=1.2419 PS=0.63 NRD=102.672 NRS=14.28 M=1 R=2.8
+ SA=75001.6 SB=75004 A=0.063 P=1.14 MULT=1
MM1019 N_A_856_304#_M1019_d N_A_714_127#_M1019_g N_VGND_M1015_d VNB NLOWVT
+ L=0.15 W=0.74 AD=0.1073 AS=0.306622 PD=1.03 PS=2.1881 NRD=0 NRS=58.272 M=1
+ R=4.93333 SA=75001.5 SB=75002.2 A=0.111 P=1.78 MULT=1
MM1005 N_A_1266_119#_M1005_d N_A_300_74#_M1005_g N_A_856_304#_M1019_d VNB NLOWVT
+ L=0.15 W=0.74 AD=0.391307 AS=0.1073 PD=2.56448 PS=1.03 NRD=51.888 NRS=1.62 M=1
+ R=4.93333 SA=75002 SB=75001.7 A=0.111 P=1.78 MULT=1
MM1021 A_1550_119# N_A_507_368#_M1021_g N_A_1266_119#_M1005_d VNB NLOWVT L=0.15
+ W=0.42 AD=0.0504 AS=0.222093 PD=0.66 PS=1.45552 NRD=18.564 NRS=0 M=1 R=2.8
+ SA=75004.2 SB=75001.5 A=0.063 P=1.14 MULT=1
MM1000 N_VGND_M1000_d N_A_1598_93#_M1000_g A_1550_119# VNB NLOWVT L=0.15 W=0.42
+ AD=0.0819 AS=0.0504 PD=0.81 PS=0.66 NRD=15.708 NRS=18.564 M=1 R=2.8 SA=75004.6
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1012 A_1736_119# N_RESET_B_M1012_g N_VGND_M1000_d VNB NLOWVT L=0.15 W=0.42
+ AD=0.0504 AS=0.0819 PD=0.66 PS=0.81 NRD=18.564 NRS=15.708 M=1 R=2.8 SA=75005.1
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1002 N_A_1598_93#_M1002_d N_A_1266_119#_M1002_g A_1736_119# VNB NLOWVT L=0.15
+ W=0.42 AD=0.1197 AS=0.0504 PD=1.41 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8
+ SA=75005.5 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1020 N_VGND_M1020_d N_A_1266_119#_M1020_g N_A_1934_94#_M1020_s VNB NLOWVT
+ L=0.15 W=0.55 AD=0.107506 AS=0.15675 PD=0.937984 PS=1.67 NRD=18 NRS=0 M=1
+ R=3.66667 SA=75000.2 SB=75000.7 A=0.0825 P=1.4 MULT=1
MM1028 N_Q_M1028_d N_A_1934_94#_M1028_g N_VGND_M1020_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.2146 AS=0.144644 PD=2.06 PS=1.26202 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.6
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1008 N_A_33_74#_M1008_d N_D_M1008_g N_VPWR_M1008_s VPB PSHORT L=0.15 W=0.42
+ AD=0.063 AS=0.1218 PD=0.72 PS=1.42 NRD=4.6886 NRS=4.6886 M=1 R=2.8 SA=75000.2
+ SB=75001.2 A=0.063 P=1.14 MULT=1
MM1007 N_VPWR_M1007_d N_RESET_B_M1007_g N_A_33_74#_M1008_d VPB PSHORT L=0.15
+ W=0.42 AD=0.0912545 AS=0.063 PD=0.804545 PS=0.72 NRD=28.1316 NRS=4.6886 M=1
+ R=2.8 SA=75000.7 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1017 N_A_300_74#_M1017_d N_CLK_N_M1017_g N_VPWR_M1007_d VPB PSHORT L=0.15
+ W=1.12 AD=0.3248 AS=0.243345 PD=2.82 PS=2.14545 NRD=1.7533 NRS=2.6201 M=1
+ R=7.46667 SA=75000.6 SB=75000.2 A=0.168 P=2.54 MULT=1
MM1009 N_A_507_368#_M1009_d N_A_300_74#_M1009_g N_VPWR_M1009_s VPB PSHORT L=0.15
+ W=1.12 AD=0.4312 AS=0.3304 PD=3.01 PS=2.83 NRD=15.8191 NRS=1.7533 M=1
+ R=7.46667 SA=75000.2 SB=75000.3 A=0.168 P=2.54 MULT=1
MM1014 N_A_714_127#_M1014_d N_A_300_74#_M1014_g N_A_33_74#_M1014_s VPB PSHORT
+ L=0.15 W=0.42 AD=0.063 AS=0.1239 PD=0.72 PS=1.43 NRD=4.6886 NRS=4.6886 M=1
+ R=2.8 SA=75000.2 SB=75001.6 A=0.063 P=1.14 MULT=1
MM1016 A_817_508# N_A_507_368#_M1016_g N_A_714_127#_M1014_d VPB PSHORT L=0.15
+ W=0.42 AD=0.0504 AS=0.063 PD=0.66 PS=0.72 NRD=30.4759 NRS=4.6886 M=1 R=2.8
+ SA=75000.7 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1004 N_VPWR_M1004_d N_A_856_304#_M1004_g A_817_508# VPB PSHORT L=0.15 W=0.42
+ AD=0.0756 AS=0.0504 PD=0.78 PS=0.66 NRD=4.6886 NRS=30.4759 M=1 R=2.8
+ SA=75001.1 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1022 N_A_714_127#_M1022_d N_RESET_B_M1022_g N_VPWR_M1004_d VPB PSHORT L=0.15
+ W=0.42 AD=0.1155 AS=0.0756 PD=1.39 PS=0.78 NRD=4.6886 NRS=32.8202 M=1 R=2.8
+ SA=75001.6 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1018 N_A_856_304#_M1018_d N_A_714_127#_M1018_g N_VPWR_M1018_s VPB PSHORT
+ L=0.15 W=1 AD=0.39 AS=0.275 PD=1.78 PS=2.55 NRD=2.9353 NRS=1.9503 M=1
+ R=6.66667 SA=75000.2 SB=75002.1 A=0.15 P=2.3 MULT=1
MM1011 N_A_1266_119#_M1011_d N_A_507_368#_M1011_g N_A_856_304#_M1018_d VPB
+ PSHORT L=0.15 W=1 AD=0.315282 AS=0.39 PD=2.39437 PS=1.78 NRD=1.9503 NRS=2.9353
+ M=1 R=6.66667 SA=75001.1 SB=75001.1 A=0.15 P=2.3 MULT=1
MM1006 A_1547_508# N_A_300_74#_M1006_g N_A_1266_119#_M1011_d VPB PSHORT L=0.15
+ W=0.42 AD=0.0567 AS=0.132418 PD=0.69 PS=1.00563 NRD=37.5088 NRS=4.6886 M=1
+ R=2.8 SA=75002 SB=75001.6 A=0.063 P=1.14 MULT=1
MM1023 N_VPWR_M1023_d N_A_1598_93#_M1023_g A_1547_508# VPB PSHORT L=0.15 W=0.42
+ AD=0.0819 AS=0.0567 PD=0.81 PS=0.69 NRD=4.6886 NRS=37.5088 M=1 R=2.8
+ SA=75002.4 SB=75001.2 A=0.063 P=1.14 MULT=1
MM1025 N_A_1598_93#_M1025_d N_RESET_B_M1025_g N_VPWR_M1023_d VPB PSHORT L=0.15
+ W=0.42 AD=0.063 AS=0.0819 PD=0.72 PS=0.81 NRD=4.6886 NRS=46.886 M=1 R=2.8
+ SA=75002.9 SB=75000.6 A=0.063 P=1.14 MULT=1
MM1031 N_VPWR_M1031_d N_A_1266_119#_M1031_g N_A_1598_93#_M1025_d VPB PSHORT
+ L=0.15 W=0.42 AD=0.1155 AS=0.063 PD=1.39 PS=0.72 NRD=4.6886 NRS=4.6886 M=1
+ R=2.8 SA=75003.4 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1003 N_VPWR_M1003_d N_A_1266_119#_M1003_g N_A_1934_94#_M1003_s VPB PSHORT
+ L=0.15 W=0.84 AD=0.1596 AS=0.231 PD=1.26429 PS=2.23 NRD=14.0658 NRS=2.3443 M=1
+ R=5.6 SA=75000.2 SB=75000.7 A=0.126 P=1.98 MULT=1
MM1001 N_Q_M1001_d N_A_1934_94#_M1001_g N_VPWR_M1003_d VPB PSHORT L=0.15 W=1.12
+ AD=0.3192 AS=0.2128 PD=2.81 PS=1.68571 NRD=1.7533 NRS=2.6201 M=1 R=7.46667
+ SA=75000.6 SB=75000.2 A=0.168 P=2.54 MULT=1
DX32_noxref VNB VPB NWDIODE A=21.1858 P=26.59
c_121 VNB 0 2.87859e-19 $X=0 $Y=0
c_1702 A_120_74# 0 1.52323e-19 $X=0.6 $Y=0.37
*
.include "sky130_fd_sc_hs__dfrtn_1.pxi.spice"
*
.ends
*
*
