* File: sky130_fd_sc_hs__inv_2.pex.spice
* Created: Thu Aug 27 20:47:56 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HS__INV_2%A 1 3 6 8 11 14 16 18 19 20 25
r39 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.27
+ $Y=1.465 $X2=0.27 $Y2=1.465
r40 22 24 11.0663 $w=3.92e-07 $l=9e-08 $layer=POLY_cond $X=0.345 $Y=1.375
+ $X2=0.345 $Y2=1.465
r41 20 25 6.9845 $w=3.28e-07 $l=2e-07 $layer=LI1_cond $X=0.27 $Y=1.665 $X2=0.27
+ $Y2=1.465
r42 16 18 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.945 $Y=1.765
+ $X2=0.945 $Y2=2.4
r43 12 19 18.8402 $w=1.65e-07 $l=7.74597e-08 $layer=POLY_cond $X=0.94 $Y=1.3
+ $X2=0.945 $Y2=1.375
r44 12 14 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=0.94 $Y=1.3 $X2=0.94
+ $Y2=0.74
r45 11 16 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=0.945 $Y=1.675
+ $X2=0.945 $Y2=1.765
r46 10 19 18.8402 $w=1.65e-07 $l=7.5e-08 $layer=POLY_cond $X=0.945 $Y=1.45
+ $X2=0.945 $Y2=1.375
r47 10 11 87.4597 $w=1.8e-07 $l=2.25e-07 $layer=POLY_cond $X=0.945 $Y=1.45
+ $X2=0.945 $Y2=1.675
r48 9 22 25.3688 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=0.585 $Y=1.375
+ $X2=0.345 $Y2=1.375
r49 8 19 6.66866 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=0.855 $Y=1.375
+ $X2=0.945 $Y2=1.375
r50 8 9 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=0.855 $Y=1.375
+ $X2=0.585 $Y2=1.375
r51 4 22 28.3659 $w=3.92e-07 $l=1.98997e-07 $layer=POLY_cond $X=0.51 $Y=1.3
+ $X2=0.345 $Y2=1.375
r52 4 6 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=0.51 $Y=1.3 $X2=0.51
+ $Y2=0.74
r53 1 24 56.0318 $w=3.92e-07 $l=3.67423e-07 $layer=POLY_cond $X=0.495 $Y=1.765
+ $X2=0.345 $Y2=1.465
r54 1 3 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.495 $Y=1.765
+ $X2=0.495 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_HS__INV_2%VPWR 1 2 7 9 13 15 19 21 31
r19 30 31 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r20 27 28 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r21 22 27 4.75569 $w=1.7e-07 $l=2.18e-07 $layer=LI1_cond $X=0.435 $Y=3.33
+ $X2=0.217 $Y2=3.33
r22 22 24 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.435 $Y=3.33
+ $X2=0.72 $Y2=3.33
r23 21 30 4.02656 $w=1.7e-07 $l=1.77e-07 $layer=LI1_cond $X=1.085 $Y=3.33
+ $X2=1.262 $Y2=3.33
r24 21 24 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=1.085 $Y=3.33
+ $X2=0.72 $Y2=3.33
r25 19 31 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r26 19 28 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r27 19 24 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r28 15 18 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=1.21 $Y=1.985
+ $X2=1.21 $Y2=2.815
r29 13 30 3.1166 $w=2.5e-07 $l=1.07912e-07 $layer=LI1_cond $X=1.21 $Y=3.245
+ $X2=1.262 $Y2=3.33
r30 13 18 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=1.21 $Y=3.245
+ $X2=1.21 $Y2=2.815
r31 9 12 24.4458 $w=3.28e-07 $l=7e-07 $layer=LI1_cond $X=0.27 $Y=2.115 $X2=0.27
+ $Y2=2.815
r32 7 27 3.01048 $w=3.3e-07 $l=1.08305e-07 $layer=LI1_cond $X=0.27 $Y=3.245
+ $X2=0.217 $Y2=3.33
r33 7 12 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=0.27 $Y=3.245
+ $X2=0.27 $Y2=2.815
r34 2 18 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=1.02
+ $Y=1.84 $X2=1.17 $Y2=2.815
r35 2 15 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=1.02
+ $Y=1.84 $X2=1.17 $Y2=1.985
r36 1 12 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.27 $Y2=2.815
r37 1 9 400 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.27 $Y2=2.115
.ends

.subckt PM_SKY130_FD_SC_HS__INV_2%Y 1 2 7 8 9 10 11 12 13 29
r24 22 29 1.3969 $w=3.28e-07 $l=4e-08 $layer=LI1_cond $X=0.725 $Y=0.965
+ $X2=0.725 $Y2=0.925
r25 12 13 14.9615 $w=2.83e-07 $l=3.7e-07 $layer=LI1_cond $X=0.747 $Y=2.405
+ $X2=0.747 $Y2=2.775
r26 11 12 16.9834 $w=2.83e-07 $l=4.2e-07 $layer=LI1_cond $X=0.747 $Y=1.985
+ $X2=0.747 $Y2=2.405
r27 10 11 12.9397 $w=2.83e-07 $l=3.2e-07 $layer=LI1_cond $X=0.747 $Y=1.665
+ $X2=0.747 $Y2=1.985
r28 9 10 14.9615 $w=2.83e-07 $l=3.7e-07 $layer=LI1_cond $X=0.747 $Y=1.295
+ $X2=0.747 $Y2=1.665
r29 9 45 6.67204 $w=2.83e-07 $l=1.65e-07 $layer=LI1_cond $X=0.747 $Y=1.295
+ $X2=0.747 $Y2=1.13
r30 8 45 5.23984 $w=3.28e-07 $l=1.43e-07 $layer=LI1_cond $X=0.725 $Y=0.987
+ $X2=0.725 $Y2=1.13
r31 8 22 0.768295 $w=3.28e-07 $l=2.2e-08 $layer=LI1_cond $X=0.725 $Y=0.987
+ $X2=0.725 $Y2=0.965
r32 8 29 0.803218 $w=3.28e-07 $l=2.3e-08 $layer=LI1_cond $X=0.725 $Y=0.902
+ $X2=0.725 $Y2=0.925
r33 7 8 13.515 $w=3.28e-07 $l=3.87e-07 $layer=LI1_cond $X=0.725 $Y=0.515
+ $X2=0.725 $Y2=0.902
r34 2 13 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=0.57
+ $Y=1.84 $X2=0.72 $Y2=2.815
r35 2 11 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=0.57
+ $Y=1.84 $X2=0.72 $Y2=1.985
r36 1 7 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=0.585
+ $Y=0.37 $X2=0.725 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__INV_2%VGND 1 2 7 9 11 13 15 17 27
r18 26 27 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r19 23 24 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r20 18 23 3.99177 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.38 $Y=0 $X2=0.19
+ $Y2=0
r21 18 20 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=0.38 $Y=0 $X2=0.72
+ $Y2=0
r22 17 26 4.0045 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=1.07 $Y=0 $X2=1.255
+ $Y2=0
r23 17 20 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=1.07 $Y=0 $X2=0.72
+ $Y2=0
r24 15 27 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r25 15 24 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r26 15 20 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r27 11 26 3.13866 $w=2.5e-07 $l=1.11018e-07 $layer=LI1_cond $X=1.195 $Y=0.085
+ $X2=1.255 $Y2=0
r28 11 13 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=1.195 $Y=0.085
+ $X2=1.195 $Y2=0.515
r29 7 23 3.1514 $w=2.5e-07 $l=1.12916e-07 $layer=LI1_cond $X=0.255 $Y=0.085
+ $X2=0.19 $Y2=0
r30 7 9 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=0.255 $Y=0.085
+ $X2=0.255 $Y2=0.515
r31 2 13 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.015
+ $Y=0.37 $X2=1.155 $Y2=0.515
r32 1 9 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.15
+ $Y=0.37 $X2=0.295 $Y2=0.515
.ends

