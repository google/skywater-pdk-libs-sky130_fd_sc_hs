* File: sky130_fd_sc_hs__clkbuf_1.pex.spice
* Created: Thu Aug 27 20:35:29 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HS__CLKBUF_1%A 3 5 7 8 9 14
c34 5 0 1.38478e-19 $X=0.735 $Y=1.765
r35 14 16 9.87705 $w=3.66e-07 $l=7.5e-08 $layer=POLY_cond $X=0.66 $Y=1.532
+ $X2=0.735 $Y2=1.532
r36 14 15 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.66
+ $Y=1.465 $X2=0.66 $Y2=1.465
r37 12 14 21.7295 $w=3.66e-07 $l=1.65e-07 $layer=POLY_cond $X=0.495 $Y=1.532
+ $X2=0.66 $Y2=1.532
r38 9 15 1.4951 $w=4.78e-07 $l=6e-08 $layer=LI1_cond $X=0.72 $Y=1.54 $X2=0.66
+ $Y2=1.54
r39 8 15 10.4657 $w=4.78e-07 $l=4.2e-07 $layer=LI1_cond $X=0.24 $Y=1.54 $X2=0.66
+ $Y2=1.54
r40 5 16 23.7042 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=0.735 $Y=1.765
+ $X2=0.735 $Y2=1.532
r41 5 7 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.735 $Y=1.765
+ $X2=0.735 $Y2=2.4
r42 1 12 23.7042 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=0.495 $Y=1.3
+ $X2=0.495 $Y2=1.532
r43 1 3 369.191 $w=1.5e-07 $l=7.2e-07 $layer=POLY_cond $X=0.495 $Y=1.3 $X2=0.495
+ $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_HS__CLKBUF_1%A_27_74# 1 2 8 9 11 14 18 20 22 24 25 26 28
+ 29 31 36 37
r68 36 39 46.536 $w=4.35e-07 $l=1.65e-07 $layer=POLY_cond $X=1.282 $Y=1.125
+ $X2=1.282 $Y2=0.96
r69 35 36 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.23
+ $Y=1.125 $X2=1.23 $Y2=1.125
r70 31 37 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=1.09 $Y=1.95 $X2=1.09
+ $Y2=1.63
r71 29 37 9.49412 $w=3.88e-07 $l=1.95e-07 $layer=LI1_cond $X=1.2 $Y=1.435
+ $X2=1.2 $Y2=1.63
r72 28 35 2.51472 $w=3.9e-07 $l=8.5e-08 $layer=LI1_cond $X=1.2 $Y=1.13 $X2=1.2
+ $Y2=1.045
r73 28 29 9.0127 $w=3.88e-07 $l=3.05e-07 $layer=LI1_cond $X=1.2 $Y=1.13 $X2=1.2
+ $Y2=1.435
r74 27 33 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.675 $Y=2.035
+ $X2=0.51 $Y2=2.035
r75 26 31 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.005 $Y=2.035
+ $X2=1.09 $Y2=1.95
r76 26 27 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=1.005 $Y=2.035
+ $X2=0.675 $Y2=2.035
r77 24 35 5.76906 $w=1.7e-07 $l=1.95e-07 $layer=LI1_cond $X=1.005 $Y=1.045
+ $X2=1.2 $Y2=1.045
r78 24 25 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=1.005 $Y=1.045
+ $X2=0.445 $Y2=1.045
r79 20 33 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.51 $Y=2.12 $X2=0.51
+ $Y2=2.035
r80 20 22 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=0.51 $Y=2.12
+ $X2=0.51 $Y2=2.815
r81 16 25 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.28 $Y=0.96
+ $X2=0.445 $Y2=1.045
r82 16 18 13.2706 $w=3.28e-07 $l=3.8e-07 $layer=LI1_cond $X=0.28 $Y=0.96
+ $X2=0.28 $Y2=0.58
r83 14 39 194.851 $w=1.5e-07 $l=3.8e-07 $layer=POLY_cond $X=1.425 $Y=0.58
+ $X2=1.425 $Y2=0.96
r84 9 11 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.285 $Y=1.765
+ $X2=1.285 $Y2=2.4
r85 8 9 50.3454 $w=3.37e-07 $l=3.53497e-07 $layer=POLY_cond $X=1.282 $Y=1.413
+ $X2=1.285 $Y2=1.765
r86 7 36 6.64828 $w=4.35e-07 $l=5.2e-08 $layer=POLY_cond $X=1.282 $Y=1.177
+ $X2=1.282 $Y2=1.125
r87 7 8 30.1729 $w=4.35e-07 $l=2.36e-07 $layer=POLY_cond $X=1.282 $Y=1.177
+ $X2=1.282 $Y2=1.413
r88 2 33 400 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_PDIFF $count=1 $X=0.365
+ $Y=1.84 $X2=0.51 $Y2=2.115
r89 2 22 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=0.365
+ $Y=1.84 $X2=0.51 $Y2=2.815
r90 1 18 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_HS__CLKBUF_1%VPWR 1 6 9 10 11 18 19
r22 18 19 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r23 14 15 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r24 11 19 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=0.96 $Y=3.33
+ $X2=1.68 $Y2=3.33
r25 11 15 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=0.96 $Y=3.33
+ $X2=0.72 $Y2=3.33
r26 9 14 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=0.845 $Y=3.33
+ $X2=0.72 $Y2=3.33
r27 9 10 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.845 $Y=3.33
+ $X2=1.01 $Y2=3.33
r28 8 18 32.9465 $w=1.68e-07 $l=5.05e-07 $layer=LI1_cond $X=1.175 $Y=3.33
+ $X2=1.68 $Y2=3.33
r29 8 10 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.175 $Y=3.33
+ $X2=1.01 $Y2=3.33
r30 4 10 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.01 $Y=3.245 $X2=1.01
+ $Y2=3.33
r31 4 6 27.5888 $w=3.28e-07 $l=7.9e-07 $layer=LI1_cond $X=1.01 $Y=3.245 $X2=1.01
+ $Y2=2.455
r32 1 6 300 $w=1.7e-07 $l=7.07972e-07 $layer=licon1_PDIFF $count=2 $X=0.81
+ $Y=1.84 $X2=1.01 $Y2=2.455
.ends

.subckt PM_SKY130_FD_SC_HS__CLKBUF_1%X 1 2 7 8 9 10 11 12 13 45 49
c25 45 0 1.38478e-19 $X=1.51 $Y=1.985
r26 45 46 7.01411 $w=4.58e-07 $l=1.65e-07 $layer=LI1_cond $X=1.575 $Y=1.985
+ $X2=1.575 $Y2=1.82
r27 30 49 0.390026 $w=4.58e-07 $l=1.5e-08 $layer=LI1_cond $X=1.575 $Y=2.05
+ $X2=1.575 $Y2=2.035
r28 13 37 1.04007 $w=4.58e-07 $l=4e-08 $layer=LI1_cond $X=1.575 $Y=2.775
+ $X2=1.575 $Y2=2.815
r29 12 13 9.62063 $w=4.58e-07 $l=3.7e-07 $layer=LI1_cond $X=1.575 $Y=2.405
+ $X2=1.575 $Y2=2.775
r30 11 49 0.91006 $w=4.58e-07 $l=3.5e-08 $layer=LI1_cond $X=1.575 $Y=2 $X2=1.575
+ $Y2=2.035
r31 11 45 0.390026 $w=4.58e-07 $l=1.5e-08 $layer=LI1_cond $X=1.575 $Y=2
+ $X2=1.575 $Y2=1.985
r32 11 12 8.32055 $w=4.58e-07 $l=3.2e-07 $layer=LI1_cond $X=1.575 $Y=2.085
+ $X2=1.575 $Y2=2.405
r33 11 30 0.91006 $w=4.58e-07 $l=3.5e-08 $layer=LI1_cond $X=1.575 $Y=2.085
+ $X2=1.575 $Y2=2.05
r34 10 46 7.44286 $w=2.38e-07 $l=1.55e-07 $layer=LI1_cond $X=1.685 $Y=1.665
+ $X2=1.685 $Y2=1.82
r35 9 10 17.7668 $w=2.38e-07 $l=3.7e-07 $layer=LI1_cond $X=1.685 $Y=1.295
+ $X2=1.685 $Y2=1.665
r36 8 9 17.7668 $w=2.38e-07 $l=3.7e-07 $layer=LI1_cond $X=1.685 $Y=0.925
+ $X2=1.685 $Y2=1.295
r37 8 43 6.48249 $w=2.38e-07 $l=1.35e-07 $layer=LI1_cond $X=1.685 $Y=0.925
+ $X2=1.685 $Y2=0.79
r38 7 43 9.08452 $w=3.28e-07 $l=2.35e-07 $layer=LI1_cond $X=1.64 $Y=0.555
+ $X2=1.64 $Y2=0.79
r39 2 45 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=1.36
+ $Y=1.84 $X2=1.51 $Y2=1.985
r40 2 37 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=1.36
+ $Y=1.84 $X2=1.51 $Y2=2.815
r41 1 7 182 $w=1.7e-07 $l=2.60768e-07 $layer=licon1_NDIFF $count=1 $X=1.5
+ $Y=0.37 $X2=1.64 $Y2=0.57
.ends

.subckt PM_SKY130_FD_SC_HS__CLKBUF_1%VGND 1 4 13 14 19 25
r19 23 25 10.279 $w=7.63e-07 $l=1.05e-07 $layer=LI1_cond $X=1.2 $Y=0.297
+ $X2=1.305 $Y2=0.297
r20 23 24 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r21 21 23 0.938101 $w=7.63e-07 $l=6e-08 $layer=LI1_cond $X=1.14 $Y=0.297 $X2=1.2
+ $Y2=0.297
r22 17 21 6.5667 $w=7.63e-07 $l=4.2e-07 $layer=LI1_cond $X=0.72 $Y=0.297
+ $X2=1.14 $Y2=0.297
r23 17 19 10.279 $w=7.63e-07 $l=1.05e-07 $layer=LI1_cond $X=0.72 $Y=0.297
+ $X2=0.615 $Y2=0.297
r24 17 18 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r25 14 24 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r26 13 25 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=1.68 $Y=0 $X2=1.305
+ $Y2=0
r27 13 14 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r28 9 18 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r29 8 19 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=0.24 $Y=0 $X2=0.615
+ $Y2=0
r30 8 9 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r31 4 24 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=0.96 $Y=0 $X2=1.2
+ $Y2=0
r32 4 18 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=0.96 $Y=0 $X2=0.72
+ $Y2=0
r33 1 21 91 $w=1.7e-07 $l=6.38396e-07 $layer=licon1_NDIFF $count=2 $X=0.57
+ $Y=0.37 $X2=1.14 $Y2=0.515
.ends

