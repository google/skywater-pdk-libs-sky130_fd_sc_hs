* File: sky130_fd_sc_hs__fahcon_1.spice
* Created: Thu Aug 27 20:46:43 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hs__fahcon_1.pex.spice"
.subckt sky130_fd_sc_hs__fahcon_1  VNB VPB A B CI VPWR COUT_N SUM VGND
* 
* VGND	VGND
* SUM	SUM
* COUT_N	COUT_N
* VPWR	VPWR
* CI	CI
* B	B
* A	A
* VPB	VPB
* VNB	VNB
MM1013 N_VGND_M1013_d N_A_M1013_g N_A_27_100#_M1013_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.263987 AS=0.2109 PD=1.5658 PS=2.05 NRD=2.424 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75002.6 A=0.111 P=1.78 MULT=1
MM1000 N_A_241_368#_M1000_d N_A_27_100#_M1000_g N_VGND_M1013_d VNB NLOWVT L=0.15
+ W=0.64 AD=0.0896 AS=0.228313 PD=0.92 PS=1.3542 NRD=0 NRS=80.616 M=1 R=4.26667
+ SA=75001.1 SB=75002.1 A=0.096 P=1.58 MULT=1
MM1001 N_A_374_120#_M1001_d N_A_336_263#_M1001_g N_A_241_368#_M1000_d VNB NLOWVT
+ L=0.15 W=0.64 AD=0.150225 AS=0.0896 PD=1.145 PS=0.92 NRD=14.988 NRS=0 M=1
+ R=4.26667 SA=75001.5 SB=75001.7 A=0.096 P=1.58 MULT=1
MM1010 N_A_27_100#_M1010_d N_B_M1010_g N_A_374_120#_M1001_d VNB NLOWVT L=0.15
+ W=0.64 AD=0.0928 AS=0.150225 PD=0.93 PS=1.145 NRD=1.872 NRS=14.988 M=1
+ R=4.26667 SA=75001.9 SB=75001.3 A=0.096 P=1.58 MULT=1
MM1029 N_A_369_365#_M1029_d N_A_336_263#_M1029_g N_A_27_100#_M1010_d VNB NLOWVT
+ L=0.15 W=0.64 AD=0.1456 AS=0.0928 PD=1.095 PS=0.93 NRD=13.116 NRS=0 M=1
+ R=4.26667 SA=75002.4 SB=75000.8 A=0.096 P=1.58 MULT=1
MM1016 N_A_241_368#_M1016_d N_B_M1016_g N_A_369_365#_M1029_d VNB NLOWVT L=0.15
+ W=0.64 AD=0.1824 AS=0.1456 PD=1.85 PS=1.095 NRD=0 NRS=19.68 M=1 R=4.26667
+ SA=75003 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1024 N_VGND_M1024_d N_B_M1024_g N_A_336_263#_M1024_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.124942 AS=0.4662 PD=1.14217 PS=2.74 NRD=7.296 NRS=2.016 M=1 R=4.93333
+ SA=75000.6 SB=75005.2 A=0.111 P=1.78 MULT=1
MM1031 N_A_1023_389#_M1031_d N_B_M1031_g N_VGND_M1024_d VNB NLOWVT L=0.15 W=0.64
+ AD=0.2496 AS=0.108058 PD=1.42 PS=0.987826 NRD=0 NRS=0 M=1 R=4.26667 SA=75001
+ SB=75005.5 A=0.096 P=1.58 MULT=1
MM1017 N_COUT_N_M1017_d N_A_369_365#_M1017_g N_A_1023_389#_M1031_d VNB NLOWVT
+ L=0.15 W=0.64 AD=0.1792 AS=0.2496 PD=1.2 PS=1.42 NRD=10.308 NRS=2.808 M=1
+ R=4.26667 SA=75002 SB=75004.6 A=0.096 P=1.58 MULT=1
MM1022 N_A_1261_421#_M1022_d N_A_374_120#_M1022_g N_COUT_N_M1017_d VNB NLOWVT
+ L=0.15 W=0.64 AD=0.176 AS=0.1792 PD=1.19 PS=1.2 NRD=50.616 NRS=42.18 M=1
+ R=4.26667 SA=75002.7 SB=75003.9 A=0.096 P=1.58 MULT=1
MM1025 N_VGND_M1025_d N_CI_M1025_g N_A_1261_421#_M1022_d VNB NLOWVT L=0.15
+ W=0.64 AD=0.118446 AS=0.176 PD=1.02029 PS=1.19 NRD=13.116 NRS=0 M=1 R=4.26667
+ SA=75003.4 SB=75003.2 A=0.096 P=1.58 MULT=1
MM1003 N_A_1606_368#_M1003_d N_CI_M1003_g N_VGND_M1025_d VNB NLOWVT L=0.15
+ W=0.74 AD=0.13883 AS=0.136954 PD=1.17971 PS=1.17971 NRD=0 NRS=1.62 M=1
+ R=4.93333 SA=75003.4 SB=75002.7 A=0.111 P=1.78 MULT=1
MM1026 N_A_1744_94#_M1026_d N_A_369_365#_M1026_g N_A_1606_368#_M1003_d VNB
+ NLOWVT L=0.15 W=0.64 AD=0.2112 AS=0.12007 PD=1.3 PS=1.02029 NRD=14.988
+ NRS=15.468 M=1 R=4.26667 SA=75003.8 SB=75002.6 A=0.096 P=1.58 MULT=1
MM1023 N_A_1719_368#_M1023_d N_A_374_120#_M1023_g N_A_1744_94#_M1026_d VNB
+ NLOWVT L=0.15 W=0.64 AD=0.1632 AS=0.2112 PD=1.15 PS=1.3 NRD=43.116 NRS=56.244
+ M=1 R=4.26667 SA=75004.6 SB=75001.8 A=0.096 P=1.58 MULT=1
MM1018 N_VGND_M1018_d N_A_1606_368#_M1018_g N_A_1719_368#_M1023_d VNB NLOWVT
+ L=0.15 W=0.64 AD=0.277472 AS=0.1632 PD=1.56754 PS=1.15 NRD=70.968 NRS=0 M=1
+ R=4.26667 SA=75005.3 SB=75001.1 A=0.096 P=1.58 MULT=1
MM1006 N_SUM_M1006_d N_A_1744_94#_M1006_g N_VGND_M1018_d VNB NLOWVT L=0.15
+ W=0.74 AD=0.2109 AS=0.320828 PD=2.05 PS=1.81246 NRD=0 NRS=61.38 M=1 R=4.93333
+ SA=75005.4 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1030 N_VPWR_M1030_d N_A_M1030_g N_A_27_100#_M1030_s VPB PSHORT L=0.15 W=1.12
+ AD=0.251683 AS=0.3304 PD=1.64302 PS=2.83 NRD=10.5395 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75002.4 A=0.168 P=2.54 MULT=1
MM1008 N_A_241_368#_M1008_d N_A_27_100#_M1008_g N_VPWR_M1030_d VPB PSHORT L=0.15
+ W=1 AD=0.249918 AS=0.224717 PD=1.63587 PS=1.46698 NRD=1.9503 NRS=19.0302 M=1
+ R=6.66667 SA=75000.8 SB=75002.1 A=0.15 P=2.3 MULT=1
MM1007 N_A_369_365#_M1007_d N_A_336_263#_M1007_g N_A_241_368#_M1008_d VPB PSHORT
+ L=0.15 W=0.84 AD=0.1764 AS=0.209932 PD=1.26 PS=1.37413 NRD=30.4759 NRS=47.28
+ M=1 R=5.6 SA=75001.4 SB=75001.8 A=0.126 P=1.98 MULT=1
MM1019 N_A_27_100#_M1019_d N_B_M1019_g N_A_369_365#_M1007_d VPB PSHORT L=0.15
+ W=0.84 AD=0.126 AS=0.1764 PD=1.14 PS=1.26 NRD=2.3443 NRS=2.3443 M=1 R=5.6
+ SA=75002 SB=75001.3 A=0.126 P=1.98 MULT=1
MM1021 N_A_374_120#_M1021_d N_A_336_263#_M1021_g N_A_27_100#_M1019_d VPB PSHORT
+ L=0.15 W=0.84 AD=0.2114 AS=0.126 PD=1.43 PS=1.14 NRD=22.261 NRS=2.3443 M=1
+ R=5.6 SA=75002.4 SB=75000.8 A=0.126 P=1.98 MULT=1
MM1027 N_A_241_368#_M1027_d N_B_M1027_g N_A_374_120#_M1021_d VPB PSHORT L=0.15
+ W=0.84 AD=0.2436 AS=0.2114 PD=2.26 PS=1.43 NRD=2.3443 NRS=22.261 M=1 R=5.6
+ SA=75003.1 SB=75000.2 A=0.126 P=1.98 MULT=1
MM1015 N_VPWR_M1015_d N_B_M1015_g N_A_336_263#_M1015_s VPB PSHORT L=0.15 W=1.12
+ AD=0.262249 AS=0.3304 PD=1.66415 PS=2.83 NRD=10.5395 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75003 A=0.168 P=2.54 MULT=1
MM1005 N_A_1023_389#_M1005_d N_B_M1005_g N_VPWR_M1015_d VPB PSHORT L=0.15 W=1
+ AD=0.201413 AS=0.234151 PD=1.50543 PS=1.48585 NRD=1.9503 NRS=22.9702 M=1
+ R=6.66667 SA=75000.8 SB=75002.7 A=0.15 P=2.3 MULT=1
MM1028 N_COUT_N_M1028_d N_A_374_120#_M1028_g N_A_1023_389#_M1005_d VPB PSHORT
+ L=0.15 W=0.84 AD=0.2121 AS=0.169187 PD=1.345 PS=1.26457 NRD=38.6908 NRS=22.655
+ M=1 R=5.6 SA=75001.4 SB=75002.6 A=0.126 P=1.98 MULT=1
MM1009 N_A_1261_421#_M1009_d N_A_369_365#_M1009_g N_COUT_N_M1028_d VPB PSHORT
+ L=0.15 W=0.84 AD=0.429678 AS=0.2121 PD=1.89 PS=1.345 NRD=2.3443 NRS=14.0658
+ M=1 R=5.6 SA=75002 SB=75001.9 A=0.126 P=1.98 MULT=1
MM1012 N_VPWR_M1012_d N_CI_M1012_g N_A_1261_421#_M1009_d VPB PSHORT L=0.15 W=1
+ AD=0.182453 AS=0.511522 PD=1.39151 PS=2.25 NRD=12.7853 NRS=1.9503 M=1
+ R=6.66667 SA=75002.7 SB=75000.7 A=0.15 P=2.3 MULT=1
MM1011 N_A_1606_368#_M1011_d N_CI_M1011_g N_VPWR_M1012_d VPB PSHORT L=0.15
+ W=1.12 AD=0.3304 AS=0.204347 PD=2.83 PS=1.55849 NRD=1.7533 NRS=1.7533 M=1
+ R=7.46667 SA=75002.9 SB=75000.2 A=0.168 P=2.54 MULT=1
MM1014 N_A_1744_94#_M1014_d N_A_369_365#_M1014_g N_A_1719_368#_M1014_s VPB
+ PSHORT L=0.15 W=0.84 AD=0.126 AS=0.4033 PD=1.14 PS=3.02 NRD=2.3443 NRS=99.682
+ M=1 R=5.6 SA=75000.3 SB=75000.7 A=0.126 P=1.98 MULT=1
MM1020 N_A_1606_368#_M1020_d N_A_374_120#_M1020_g N_A_1744_94#_M1014_d VPB
+ PSHORT L=0.15 W=0.84 AD=0.2478 AS=0.126 PD=2.27 PS=1.14 NRD=2.3443 NRS=2.3443
+ M=1 R=5.6 SA=75000.8 SB=75000.2 A=0.126 P=1.98 MULT=1
MM1004 N_VPWR_M1004_d N_A_1606_368#_M1004_g N_A_1719_368#_M1004_s VPB PSHORT
+ L=0.15 W=1 AD=0.182453 AS=0.295 PD=1.39151 PS=2.59 NRD=1.9503 NRS=1.9503 M=1
+ R=6.66667 SA=75000.2 SB=75000.7 A=0.15 P=2.3 MULT=1
MM1002 N_SUM_M1002_d N_A_1744_94#_M1002_g N_VPWR_M1004_d VPB PSHORT L=0.15
+ W=1.12 AD=0.3304 AS=0.204347 PD=2.83 PS=1.55849 NRD=1.7533 NRS=11.426 M=1
+ R=7.46667 SA=75000.7 SB=75000.2 A=0.168 P=2.54 MULT=1
DX32_noxref VNB VPB NWDIODE A=22.1908 P=27.55
c_226 VPB 0 1.25754e-19 $X=0 $Y=3.085
*
.include "sky130_fd_sc_hs__fahcon_1.pxi.spice"
*
.ends
*
*
