* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hs__dlrtn_1 D GATE_N RESET_B VGND VNB VPB VPWR Q
M1000 VPWR D a_27_136# VPB pshort w=840000u l=150000u
+  ad=1.81275e+12p pd=1.271e+07u as=2.478e+11p ps=2.27e+06u
M1001 a_232_98# GATE_N VPWR VPB pshort w=840000u l=150000u
+  ad=2.478e+11p pd=2.27e+06u as=0p ps=0u
M1002 a_232_98# GATE_N VGND VNB nlowvt w=740000u l=150000u
+  ad=1.961e+11p pd=2.01e+06u as=1.64835e+12p ps=1.063e+07u
M1003 VGND a_897_406# a_854_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.155e+11p ps=1.39e+06u
M1004 a_654_392# a_357_392# a_570_392# VPB pshort w=1e+06u l=150000u
+  ad=4.029e+11p pd=3.09e+06u as=2.7e+11p ps=2.54e+06u
M1005 a_897_406# a_654_392# VPWR VPB pshort w=1e+06u l=150000u
+  ad=4.7e+11p pd=2.94e+06u as=0p ps=0u
M1006 a_854_74# a_357_392# a_654_392# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.915e+11p ps=1.93e+06u
M1007 Q a_897_406# VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=3.304e+11p pd=2.83e+06u as=0p ps=0u
M1008 VGND RESET_B a_1139_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=1.776e+11p ps=1.96e+06u
M1009 a_681_74# a_27_136# VGND VNB nlowvt w=640000u l=150000u
+  ad=1.536e+11p pd=1.76e+06u as=0p ps=0u
M1010 a_793_508# a_232_98# a_654_392# VPB pshort w=420000u l=150000u
+  ad=2.247e+11p pd=1.91e+06u as=0p ps=0u
M1011 VGND D a_27_136# VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=1.5675e+11p ps=1.67e+06u
M1012 a_1139_74# a_654_392# a_897_406# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1013 Q a_897_406# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.701e+11p pd=2.21e+06u as=0p ps=0u
M1014 VPWR a_232_98# a_357_392# VPB pshort w=840000u l=150000u
+  ad=0p pd=0u as=2.478e+11p ps=2.27e+06u
M1015 VGND a_232_98# a_357_392# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1016 a_654_392# a_232_98# a_681_74# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 VPWR a_897_406# a_793_508# VPB pshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 VPWR RESET_B a_897_406# VPB pshort w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_570_392# a_27_136# VPWR VPB pshort w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
