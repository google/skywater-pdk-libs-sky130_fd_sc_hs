* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hs__sdlclkp_1 CLK GATE SCE VGND VNB VPB VPWR GCLK
X0 VGND a_288_48# a_318_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X1 VGND a_1238_94# GCLK VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X2 a_722_492# a_709_54# VPWR VPB sky130_fd_pr__pfet_01v8 w=420000u l=150000u
X3 VPWR CLK a_1238_94# VPB sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X4 a_1166_94# a_709_54# a_1238_94# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X5 a_116_424# GATE a_114_112# VPB sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X6 VPWR a_288_48# a_318_74# VPB sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X7 a_288_48# CLK VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X8 a_114_112# a_288_48# a_566_74# VNB sky130_fd_pr__nfet_01v8_lvt w=550000u l=150000u
X9 VPWR a_566_74# a_709_54# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X10 a_566_74# a_318_74# a_667_80# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X11 a_288_48# CLK VPWR VPB sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X12 a_114_112# a_318_74# a_566_74# VPB sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X13 VGND SCE a_114_112# VNB sky130_fd_pr__nfet_01v8_lvt w=550000u l=150000u
X14 a_1238_94# a_709_54# VPWR VPB sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X15 a_114_112# GATE VGND VNB sky130_fd_pr__nfet_01v8_lvt w=550000u l=150000u
X16 VGND CLK a_1166_94# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X17 VPWR a_1238_94# GCLK VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X18 a_667_80# a_709_54# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X19 VPWR SCE a_116_424# VPB sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X20 a_566_74# a_288_48# a_722_492# VPB sky130_fd_pr__pfet_01v8 w=420000u l=150000u
X21 VGND a_566_74# a_709_54# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
.ends
