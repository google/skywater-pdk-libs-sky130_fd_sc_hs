* File: sky130_fd_sc_hs__maj3_4.pex.spice
* Created: Thu Aug 27 20:48:38 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HS__MAJ3_4%B 1 3 4 6 7 9 10 12 13 15 16 18 19 21 22 24
+ 27 31 32 33 39 46 49
c114 16 0 1.44963e-19 $X=2.935 $Y=1.375
c115 1 0 1.94433e-19 $X=1.02 $Y=1.885
r116 46 47 1.72967 $w=4.18e-07 $l=1.5e-08 $layer=POLY_cond $X=3.365 $Y=1.63
+ $X2=3.38 $Y2=1.63
r117 44 46 47.2775 $w=4.18e-07 $l=4.1e-07 $layer=POLY_cond $X=2.955 $Y=1.63
+ $X2=3.365 $Y2=1.63
r118 44 45 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.955
+ $Y=1.54 $X2=2.955 $Y2=1.54
r119 42 44 2.30622 $w=4.18e-07 $l=2e-08 $layer=POLY_cond $X=2.935 $Y=1.63
+ $X2=2.955 $Y2=1.63
r120 41 42 6.34211 $w=4.18e-07 $l=5.5e-08 $layer=POLY_cond $X=2.88 $Y=1.63
+ $X2=2.935 $Y2=1.63
r121 39 40 5.25182 $w=4.13e-07 $l=4.5e-08 $layer=POLY_cond $X=1.47 $Y=1.63
+ $X2=1.515 $Y2=1.63
r122 36 37 7.58596 $w=4.13e-07 $l=6.5e-08 $layer=POLY_cond $X=1.02 $Y=1.63
+ $X2=1.085 $Y2=1.63
r123 33 45 3.43222 $w=5.73e-07 $l=1.65e-07 $layer=LI1_cond $X=3.12 $Y=1.417
+ $X2=2.955 $Y2=1.417
r124 32 45 6.55243 $w=5.73e-07 $l=3.15e-07 $layer=LI1_cond $X=2.64 $Y=1.417
+ $X2=2.955 $Y2=1.417
r125 32 49 8.95336 $w=5.73e-07 $l=1.15e-07 $layer=LI1_cond $X=2.64 $Y=1.417
+ $X2=2.525 $Y2=1.417
r126 31 49 69.1551 $w=1.68e-07 $l=1.06e-06 $layer=LI1_cond $X=1.465 $Y=1.215
+ $X2=2.525 $Y2=1.215
r127 28 39 19.8402 $w=4.13e-07 $l=1.7e-07 $layer=POLY_cond $X=1.3 $Y=1.63
+ $X2=1.47 $Y2=1.63
r128 28 37 25.092 $w=4.13e-07 $l=2.15e-07 $layer=POLY_cond $X=1.3 $Y=1.63
+ $X2=1.085 $Y2=1.63
r129 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.3
+ $Y=1.54 $X2=1.3 $Y2=1.54
r130 25 31 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.3 $Y=1.3
+ $X2=1.465 $Y2=1.215
r131 25 27 8.3814 $w=3.28e-07 $l=2.4e-07 $layer=LI1_cond $X=1.3 $Y=1.3 $X2=1.3
+ $Y2=1.54
r132 22 47 26.9416 $w=1.5e-07 $l=2.55e-07 $layer=POLY_cond $X=3.38 $Y=1.885
+ $X2=3.38 $Y2=1.63
r133 22 24 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=3.38 $Y=1.885
+ $X2=3.38 $Y2=2.46
r134 19 46 26.9416 $w=1.5e-07 $l=2.55e-07 $layer=POLY_cond $X=3.365 $Y=1.375
+ $X2=3.365 $Y2=1.63
r135 19 21 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=3.365 $Y=1.375
+ $X2=3.365 $Y2=0.945
r136 16 42 26.9416 $w=1.5e-07 $l=2.55e-07 $layer=POLY_cond $X=2.935 $Y=1.375
+ $X2=2.935 $Y2=1.63
r137 16 18 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=2.935 $Y=1.375
+ $X2=2.935 $Y2=0.945
r138 13 41 26.9416 $w=1.5e-07 $l=2.55e-07 $layer=POLY_cond $X=2.88 $Y=1.885
+ $X2=2.88 $Y2=1.63
r139 13 15 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=2.88 $Y=1.885
+ $X2=2.88 $Y2=2.46
r140 10 40 26.6457 $w=1.5e-07 $l=2.55e-07 $layer=POLY_cond $X=1.515 $Y=1.375
+ $X2=1.515 $Y2=1.63
r141 10 12 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=1.515 $Y=1.375
+ $X2=1.515 $Y2=0.945
r142 7 39 26.6457 $w=1.5e-07 $l=2.55e-07 $layer=POLY_cond $X=1.47 $Y=1.885
+ $X2=1.47 $Y2=1.63
r143 7 9 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=1.47 $Y=1.885
+ $X2=1.47 $Y2=2.46
r144 4 37 26.6457 $w=1.5e-07 $l=2.55e-07 $layer=POLY_cond $X=1.085 $Y=1.375
+ $X2=1.085 $Y2=1.63
r145 4 6 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=1.085 $Y=1.375
+ $X2=1.085 $Y2=0.945
r146 1 36 26.6457 $w=1.5e-07 $l=2.55e-07 $layer=POLY_cond $X=1.02 $Y=1.885
+ $X2=1.02 $Y2=1.63
r147 1 3 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=1.02 $Y=1.885
+ $X2=1.02 $Y2=2.46
.ends

.subckt PM_SKY130_FD_SC_HS__MAJ3_4%A 4 6 7 9 10 11 12 14 18 19 21 25 26 27 29 30
+ 32 36 38 40 41 45 48
c159 29 0 1.41402e-19 $X=5.8 $Y=1.795
c160 18 0 9.20449e-20 $X=2.015 $Y=0.945
r161 51 52 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.965
+ $Y=1.635 $X2=1.965 $Y2=1.635
r162 48 52 1.06087 $w=3.45e-07 $l=3e-08 $layer=LI1_cond $X=2.037 $Y=1.665
+ $X2=2.037 $Y2=1.635
r163 45 46 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.405
+ $Y=1.635 $X2=4.405 $Y2=1.635
r164 43 45 8.3814 $w=3.28e-07 $l=2.4e-07 $layer=LI1_cond $X=4.405 $Y=1.875
+ $X2=4.405 $Y2=1.635
r165 42 48 10.4319 $w=3.45e-07 $l=3.96529e-07 $layer=LI1_cond $X=2.275 $Y=1.96
+ $X2=2.037 $Y2=1.665
r166 41 43 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.24 $Y=1.96
+ $X2=4.405 $Y2=1.875
r167 41 42 128.198 $w=1.68e-07 $l=1.965e-06 $layer=LI1_cond $X=4.24 $Y=1.96
+ $X2=2.275 $Y2=1.96
r168 39 40 60.4563 $w=1.8e-07 $l=1.5e-07 $layer=POLY_cond $X=5.805 $Y=1.31
+ $X2=5.805 $Y2=1.46
r169 37 38 60.4563 $w=1.8e-07 $l=1.5e-07 $layer=POLY_cond $X=0.515 $Y=1.34
+ $X2=0.515 $Y2=1.49
r170 36 39 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=5.825 $Y=0.915
+ $X2=5.825 $Y2=1.31
r171 33 36 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=5.825 $Y=0.255
+ $X2=5.825 $Y2=0.915
r172 30 32 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=5.8 $Y=1.885
+ $X2=5.8 $Y2=2.46
r173 29 30 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=5.8 $Y=1.795 $X2=5.8
+ $Y2=1.885
r174 29 40 130.218 $w=1.8e-07 $l=3.35e-07 $layer=POLY_cond $X=5.8 $Y=1.795
+ $X2=5.8 $Y2=1.46
r175 26 33 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.75 $Y=0.18
+ $X2=5.825 $Y2=0.255
r176 26 27 625.574 $w=1.5e-07 $l=1.22e-06 $layer=POLY_cond $X=5.75 $Y=0.18
+ $X2=4.53 $Y2=0.18
r177 23 46 38.5562 $w=2.99e-07 $l=1.88348e-07 $layer=POLY_cond $X=4.455 $Y=1.47
+ $X2=4.405 $Y2=1.635
r178 23 25 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=4.455 $Y=1.47
+ $X2=4.455 $Y2=0.71
r179 22 27 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.455 $Y=0.255
+ $X2=4.53 $Y2=0.18
r180 22 25 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=4.455 $Y=0.255
+ $X2=4.455 $Y2=0.71
r181 19 46 52.2586 $w=2.99e-07 $l=2.7157e-07 $layer=POLY_cond $X=4.45 $Y=1.885
+ $X2=4.405 $Y2=1.635
r182 19 21 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=4.45 $Y=1.885
+ $X2=4.45 $Y2=2.46
r183 16 51 38.5562 $w=2.99e-07 $l=1.88348e-07 $layer=POLY_cond $X=2.015 $Y=1.47
+ $X2=1.965 $Y2=1.635
r184 16 18 269.202 $w=1.5e-07 $l=5.25e-07 $layer=POLY_cond $X=2.015 $Y=1.47
+ $X2=2.015 $Y2=0.945
r185 15 18 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=2.015 $Y=0.255
+ $X2=2.015 $Y2=0.945
r186 12 51 52.2586 $w=2.99e-07 $l=2.7157e-07 $layer=POLY_cond $X=1.92 $Y=1.885
+ $X2=1.965 $Y2=1.635
r187 12 14 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=1.92 $Y=1.885
+ $X2=1.92 $Y2=2.46
r188 10 15 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.94 $Y=0.18
+ $X2=2.015 $Y2=0.255
r189 10 11 702.489 $w=1.5e-07 $l=1.37e-06 $layer=POLY_cond $X=1.94 $Y=0.18
+ $X2=0.57 $Y2=0.18
r190 7 9 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=0.52 $Y=1.885
+ $X2=0.52 $Y2=2.46
r191 6 7 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=0.52 $Y=1.795 $X2=0.52
+ $Y2=1.885
r192 6 38 118.556 $w=1.8e-07 $l=3.05e-07 $layer=POLY_cond $X=0.52 $Y=1.795
+ $X2=0.52 $Y2=1.49
r193 4 37 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=0.495 $Y=0.945
+ $X2=0.495 $Y2=1.34
r194 1 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.495 $Y=0.255
+ $X2=0.57 $Y2=0.18
r195 1 4 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=0.495 $Y=0.255
+ $X2=0.495 $Y2=0.945
.ends

.subckt PM_SKY130_FD_SC_HS__MAJ3_4%C 1 2 3 5 9 10 11 12 14 18 19 21 24 26 28 31
+ 34 37 41 44 52 54
c139 41 0 1.41402e-19 $X=5.055 $Y=1.635
c140 18 0 1.46446e-19 $X=3.955 $Y=0.71
r141 52 53 5.89402 $w=3.68e-07 $l=4.5e-08 $layer=POLY_cond $X=5.35 $Y=1.677
+ $X2=5.395 $Y2=1.677
r142 49 50 8.51359 $w=3.68e-07 $l=6.5e-08 $layer=POLY_cond $X=4.9 $Y=1.677
+ $X2=4.965 $Y2=1.677
r143 47 48 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.845
+ $Y=1.54 $X2=3.845 $Y2=1.54
r144 44 48 5.5817 $w=5.23e-07 $l=2.45e-07 $layer=LI1_cond $X=3.747 $Y=1.295
+ $X2=3.747 $Y2=1.54
r145 44 54 1.8226 $w=5.23e-07 $l=8e-08 $layer=LI1_cond $X=3.747 $Y=1.295
+ $X2=3.747 $Y2=1.215
r146 42 52 38.6386 $w=3.68e-07 $l=2.95e-07 $layer=POLY_cond $X=5.055 $Y=1.677
+ $X2=5.35 $Y2=1.677
r147 42 50 11.788 $w=3.68e-07 $l=9e-08 $layer=POLY_cond $X=5.055 $Y=1.677
+ $X2=4.965 $Y2=1.677
r148 41 42 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.055
+ $Y=1.635 $X2=5.055 $Y2=1.635
r149 38 41 7.50834 $w=3.28e-07 $l=2.15e-07 $layer=LI1_cond $X=4.84 $Y=1.635
+ $X2=5.055 $Y2=1.635
r150 37 38 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.84 $Y=1.47
+ $X2=4.84 $Y2=1.635
r151 36 37 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=4.84 $Y=1.3
+ $X2=4.84 $Y2=1.47
r152 35 54 7.46409 $w=1.7e-07 $l=2.63e-07 $layer=LI1_cond $X=4.01 $Y=1.215
+ $X2=3.747 $Y2=1.215
r153 34 36 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.755 $Y=1.215
+ $X2=4.84 $Y2=1.3
r154 34 35 48.6043 $w=1.68e-07 $l=7.45e-07 $layer=LI1_cond $X=4.755 $Y=1.215
+ $X2=4.01 $Y2=1.215
r155 29 53 23.8357 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=5.395 $Y=1.47
+ $X2=5.395 $Y2=1.677
r156 29 31 284.585 $w=1.5e-07 $l=5.55e-07 $layer=POLY_cond $X=5.395 $Y=1.47
+ $X2=5.395 $Y2=0.915
r157 26 52 23.8357 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=5.35 $Y=1.885
+ $X2=5.35 $Y2=1.677
r158 26 28 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=5.35 $Y=1.885
+ $X2=5.35 $Y2=2.46
r159 22 50 23.8357 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.965 $Y=1.47
+ $X2=4.965 $Y2=1.677
r160 22 24 284.585 $w=1.5e-07 $l=5.55e-07 $layer=POLY_cond $X=4.965 $Y=1.47
+ $X2=4.965 $Y2=0.915
r161 19 49 23.8357 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=4.9 $Y=1.885
+ $X2=4.9 $Y2=1.677
r162 19 21 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=4.9 $Y=1.885
+ $X2=4.9 $Y2=2.46
r163 16 47 38.6157 $w=2.9e-07 $l=2.09105e-07 $layer=POLY_cond $X=3.955 $Y=1.375
+ $X2=3.855 $Y2=1.54
r164 16 18 340.989 $w=1.5e-07 $l=6.65e-07 $layer=POLY_cond $X=3.955 $Y=1.375
+ $X2=3.955 $Y2=0.71
r165 15 18 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=3.955 $Y=0.255
+ $X2=3.955 $Y2=0.71
r166 12 47 68.5329 $w=2.9e-07 $l=3.57281e-07 $layer=POLY_cond $X=3.88 $Y=1.885
+ $X2=3.855 $Y2=1.54
r167 12 14 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=3.88 $Y=1.885
+ $X2=3.88 $Y2=2.46
r168 10 15 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.88 $Y=0.18
+ $X2=3.955 $Y2=0.255
r169 10 11 697.362 $w=1.5e-07 $l=1.36e-06 $layer=POLY_cond $X=3.88 $Y=0.18
+ $X2=2.52 $Y2=0.18
r170 9 33 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=2.445 $Y=0.945
+ $X2=2.445 $Y2=1.34
r171 6 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.445 $Y=0.255
+ $X2=2.52 $Y2=0.18
r172 6 9 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=2.445 $Y=0.255
+ $X2=2.445 $Y2=0.945
r173 3 5 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=2.43 $Y=1.885
+ $X2=2.43 $Y2=2.46
r174 2 3 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=2.43 $Y=1.795 $X2=2.43
+ $Y2=1.885
r175 1 33 37.1337 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=2.43 $Y=1.43 $X2=2.43
+ $Y2=1.34
r176 1 2 141.879 $w=1.8e-07 $l=3.65e-07 $layer=POLY_cond $X=2.43 $Y=1.43
+ $X2=2.43 $Y2=1.795
.ends

.subckt PM_SKY130_FD_SC_HS__MAJ3_4%A_219_392# 1 2 3 4 5 6 19 21 22 24 25 27 28
+ 30 31 33 34 36 37 39 40 42 43 44 45 48 51 53 57 59 61 67 68 74 84 86 88 93 96
+ 107
c220 88 0 1.44963e-19 $X=3.15 $Y=0.78
c221 84 0 1.94433e-19 $X=1.252 $Y=2.3
c222 68 0 1.04924e-19 $X=5.475 $Y=1.97
c223 43 0 9.20449e-20 $X=0.88 $Y=0.96
c224 28 0 1.55372e-19 $X=6.805 $Y=1.345
c225 22 0 1.82103e-19 $X=6.335 $Y=1.345
r226 107 108 1.30623 $w=3.69e-07 $l=1e-08 $layer=POLY_cond $X=7.655 $Y=1.555
+ $X2=7.665 $Y2=1.555
r227 106 107 54.8618 $w=3.69e-07 $l=4.2e-07 $layer=POLY_cond $X=7.235 $Y=1.555
+ $X2=7.655 $Y2=1.555
r228 105 106 3.9187 $w=3.69e-07 $l=3e-08 $layer=POLY_cond $X=7.205 $Y=1.555
+ $X2=7.235 $Y2=1.555
r229 102 103 6.53117 $w=3.69e-07 $l=5e-08 $layer=POLY_cond $X=6.755 $Y=1.555
+ $X2=6.805 $Y2=1.555
r230 101 102 54.8618 $w=3.69e-07 $l=4.2e-07 $layer=POLY_cond $X=6.335 $Y=1.555
+ $X2=6.755 $Y2=1.555
r231 96 98 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=5.18 $Y=0.76
+ $X2=5.18 $Y2=0.875
r232 88 90 4.37928 $w=2.48e-07 $l=9.5e-08 $layer=LI1_cond $X=3.19 $Y=0.78
+ $X2=3.19 $Y2=0.875
r233 75 105 28.7371 $w=3.69e-07 $l=2.2e-07 $layer=POLY_cond $X=6.985 $Y=1.555
+ $X2=7.205 $Y2=1.555
r234 75 103 23.5122 $w=3.69e-07 $l=1.8e-07 $layer=POLY_cond $X=6.985 $Y=1.555
+ $X2=6.805 $Y2=1.555
r235 74 75 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=6.985
+ $Y=1.51 $X2=6.985 $Y2=1.51
r236 72 101 3.9187 $w=3.69e-07 $l=3e-08 $layer=POLY_cond $X=6.305 $Y=1.555
+ $X2=6.335 $Y2=1.555
r237 71 74 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=6.305 $Y=1.51
+ $X2=6.985 $Y2=1.51
r238 71 72 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=6.305
+ $Y=1.51 $X2=6.305 $Y2=1.51
r239 69 71 26.0173 $w=3.28e-07 $l=7.45e-07 $layer=LI1_cond $X=5.56 $Y=1.51
+ $X2=6.305 $Y2=1.51
r240 68 93 14.0461 $w=3.04e-07 $l=4.41531e-07 $layer=LI1_cond $X=5.475 $Y=1.97
+ $X2=5.125 $Y2=2.177
r241 67 69 9.18505 $w=2.62e-07 $l=2.03101e-07 $layer=LI1_cond $X=5.475 $Y=1.675
+ $X2=5.39 $Y2=1.51
r242 67 68 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=5.475 $Y=1.675
+ $X2=5.475 $Y2=1.97
r243 64 69 19.1965 $w=2.62e-07 $l=4.73498e-07 $layer=LI1_cond $X=5.18 $Y=1.13
+ $X2=5.39 $Y2=1.51
r244 64 66 1.95722 $w=1.68e-07 $l=3e-08 $layer=LI1_cond $X=5.18 $Y=1.13 $X2=5.18
+ $Y2=1.1
r245 63 98 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=5.18 $Y=0.96
+ $X2=5.18 $Y2=0.875
r246 63 66 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=5.18 $Y=0.96
+ $X2=5.18 $Y2=1.1
r247 62 86 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.32 $Y=2.3
+ $X2=3.155 $Y2=2.3
r248 61 93 8.97325 $w=3.04e-07 $l=2.17991e-07 $layer=LI1_cond $X=4.96 $Y=2.3
+ $X2=5.125 $Y2=2.177
r249 61 62 106.995 $w=1.68e-07 $l=1.64e-06 $layer=LI1_cond $X=4.96 $Y=2.3
+ $X2=3.32 $Y2=2.3
r250 60 90 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.315 $Y=0.875
+ $X2=3.19 $Y2=0.875
r251 59 98 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.095 $Y=0.875
+ $X2=5.18 $Y2=0.875
r252 59 60 116.128 $w=1.68e-07 $l=1.78e-06 $layer=LI1_cond $X=5.095 $Y=0.875
+ $X2=3.315 $Y2=0.875
r253 55 86 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.155 $Y=2.385
+ $X2=3.155 $Y2=2.3
r254 55 57 9.25447 $w=3.28e-07 $l=2.65e-07 $layer=LI1_cond $X=3.155 $Y=2.385
+ $X2=3.155 $Y2=2.65
r255 54 84 3.25423 $w=1.7e-07 $l=1.58e-07 $layer=LI1_cond $X=1.41 $Y=2.3
+ $X2=1.252 $Y2=2.3
r256 53 86 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.99 $Y=2.3
+ $X2=3.155 $Y2=2.3
r257 53 54 103.08 $w=1.68e-07 $l=1.58e-06 $layer=LI1_cond $X=2.99 $Y=2.3
+ $X2=1.41 $Y2=2.3
r258 49 84 3.29812 $w=2.85e-07 $l=9.88686e-08 $layer=LI1_cond $X=1.222 $Y=2.385
+ $X2=1.252 $Y2=2.3
r259 49 51 8.36086 $w=2.53e-07 $l=1.85e-07 $layer=LI1_cond $X=1.222 $Y=2.385
+ $X2=1.222 $Y2=2.57
r260 46 84 3.29812 $w=2.85e-07 $l=8.5e-08 $layer=LI1_cond $X=1.252 $Y=2.215
+ $X2=1.252 $Y2=2.3
r261 46 48 2.0122 $w=3.13e-07 $l=5.5e-08 $layer=LI1_cond $X=1.252 $Y=2.215
+ $X2=1.252 $Y2=2.16
r262 45 80 24.2695 $w=1.68e-07 $l=3.72e-07 $layer=LI1_cond $X=1.252 $Y=1.96
+ $X2=0.88 $Y2=1.96
r263 45 48 4.20733 $w=3.13e-07 $l=1.15e-07 $layer=LI1_cond $X=1.252 $Y=2.045
+ $X2=1.252 $Y2=2.16
r264 44 80 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.88 $Y=1.875
+ $X2=0.88 $Y2=1.96
r265 43 79 19.6322 $w=2.61e-07 $l=5.35593e-07 $layer=LI1_cond $X=0.88 $Y=0.96
+ $X2=1.3 $Y2=0.697
r266 43 44 59.6952 $w=1.68e-07 $l=9.15e-07 $layer=LI1_cond $X=0.88 $Y=0.96
+ $X2=0.88 $Y2=1.875
r267 40 108 23.9013 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=7.665 $Y=1.345
+ $X2=7.665 $Y2=1.555
r268 40 42 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=7.665 $Y=1.345
+ $X2=7.665 $Y2=0.865
r269 37 107 23.9013 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=7.655 $Y=1.765
+ $X2=7.655 $Y2=1.555
r270 37 39 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=7.655 $Y=1.765
+ $X2=7.655 $Y2=2.4
r271 34 106 23.9013 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=7.235 $Y=1.345
+ $X2=7.235 $Y2=1.555
r272 34 36 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=7.235 $Y=1.345
+ $X2=7.235 $Y2=0.865
r273 31 105 23.9013 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=7.205 $Y=1.765
+ $X2=7.205 $Y2=1.555
r274 31 33 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=7.205 $Y=1.765
+ $X2=7.205 $Y2=2.4
r275 28 103 23.9013 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=6.805 $Y=1.345
+ $X2=6.805 $Y2=1.555
r276 28 30 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=6.805 $Y=1.345
+ $X2=6.805 $Y2=0.865
r277 25 102 23.9013 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=6.755 $Y=1.765
+ $X2=6.755 $Y2=1.555
r278 25 27 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=6.755 $Y=1.765
+ $X2=6.755 $Y2=2.4
r279 22 101 23.9013 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=6.335 $Y=1.345
+ $X2=6.335 $Y2=1.555
r280 22 24 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=6.335 $Y=1.345
+ $X2=6.335 $Y2=0.865
r281 19 72 23.9013 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=6.305 $Y=1.765
+ $X2=6.305 $Y2=1.555
r282 19 21 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=6.305 $Y=1.765
+ $X2=6.305 $Y2=2.4
r283 6 93 600 $w=1.7e-07 $l=3.21364e-07 $layer=licon1_PDIFF $count=1 $X=4.975
+ $Y=1.96 $X2=5.125 $Y2=2.215
r284 5 86 600 $w=1.7e-07 $l=4.28486e-07 $layer=licon1_PDIFF $count=1 $X=2.955
+ $Y=1.96 $X2=3.155 $Y2=2.3
r285 5 57 600 $w=1.7e-07 $l=7.83645e-07 $layer=licon1_PDIFF $count=1 $X=2.955
+ $Y=1.96 $X2=3.155 $Y2=2.65
r286 4 51 600 $w=1.7e-07 $l=6.80882e-07 $layer=licon1_PDIFF $count=1 $X=1.095
+ $Y=1.96 $X2=1.245 $Y2=2.57
r287 4 48 600 $w=1.7e-07 $l=2.64575e-07 $layer=licon1_PDIFF $count=1 $X=1.095
+ $Y=1.96 $X2=1.245 $Y2=2.16
r288 3 96 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=5.04
+ $Y=0.595 $X2=5.18 $Y2=0.76
r289 3 66 182 $w=1.7e-07 $l=5.70723e-07 $layer=licon1_NDIFF $count=1 $X=5.04
+ $Y=0.595 $X2=5.18 $Y2=1.1
r290 2 88 182 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_NDIFF $count=1 $X=3.01
+ $Y=0.625 $X2=3.15 $Y2=0.78
r291 1 79 182 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_NDIFF $count=1 $X=1.16
+ $Y=0.625 $X2=1.3 $Y2=0.78
.ends

.subckt PM_SKY130_FD_SC_HS__MAJ3_4%VPWR 1 2 3 4 5 6 19 21 27 31 35 39 43 45 47
+ 51 53 61 69 74 83 86 89 92 96
r112 95 96 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r113 92 93 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r114 90 93 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6 $Y=3.33 $X2=6.96
+ $Y2=3.33
r115 89 90 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r116 83 84 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r117 80 81 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r118 78 96 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=7.92 $Y2=3.33
r119 78 93 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=6.96 $Y2=3.33
r120 77 78 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r121 75 92 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.145 $Y=3.33
+ $X2=7.02 $Y2=3.33
r122 75 77 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=7.145 $Y=3.33
+ $X2=7.44 $Y2=3.33
r123 74 95 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=7.715 $Y=3.33
+ $X2=7.937 $Y2=3.33
r124 74 77 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=7.715 $Y=3.33
+ $X2=7.44 $Y2=3.33
r125 73 90 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=6 $Y2=3.33
r126 72 73 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r127 70 86 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.32 $Y=3.33
+ $X2=4.155 $Y2=3.33
r128 70 72 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=4.32 $Y=3.33
+ $X2=4.56 $Y2=3.33
r129 69 89 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.94 $Y=3.33
+ $X2=6.065 $Y2=3.33
r130 69 72 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=5.94 $Y=3.33
+ $X2=4.56 $Y2=3.33
r131 67 68 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r132 65 68 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.6 $Y2=3.33
r133 65 84 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=2.16 $Y2=3.33
r134 64 67 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=2.64 $Y=3.33 $X2=3.6
+ $Y2=3.33
r135 64 65 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r136 62 83 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.32 $Y=3.33
+ $X2=2.19 $Y2=3.33
r137 62 64 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=2.32 $Y=3.33
+ $X2=2.64 $Y2=3.33
r138 61 86 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.99 $Y=3.33
+ $X2=4.155 $Y2=3.33
r139 61 67 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=3.99 $Y=3.33
+ $X2=3.6 $Y2=3.33
r140 60 84 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r141 59 60 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r142 57 60 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.68 $Y2=3.33
r143 57 81 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r144 56 59 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.72 $Y=3.33
+ $X2=1.68 $Y2=3.33
r145 56 57 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r146 54 80 3.99177 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.38 $Y=3.33
+ $X2=0.19 $Y2=3.33
r147 54 56 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=0.38 $Y=3.33
+ $X2=0.72 $Y2=3.33
r148 53 83 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.06 $Y=3.33
+ $X2=2.19 $Y2=3.33
r149 53 59 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=2.06 $Y=3.33
+ $X2=1.68 $Y2=3.33
r150 51 73 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=4.56 $Y2=3.33
r151 51 68 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=3.6 $Y2=3.33
r152 51 86 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r153 47 50 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=7.88 $Y=1.985
+ $X2=7.88 $Y2=2.815
r154 45 95 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=7.88 $Y=3.245
+ $X2=7.937 $Y2=3.33
r155 45 50 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=7.88 $Y=3.245
+ $X2=7.88 $Y2=2.815
r156 41 92 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=7.02 $Y=3.245
+ $X2=7.02 $Y2=3.33
r157 41 43 41.2575 $w=2.48e-07 $l=8.95e-07 $layer=LI1_cond $X=7.02 $Y=3.245
+ $X2=7.02 $Y2=2.35
r158 40 89 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.19 $Y=3.33
+ $X2=6.065 $Y2=3.33
r159 39 92 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.895 $Y=3.33
+ $X2=7.02 $Y2=3.33
r160 39 40 45.9947 $w=1.68e-07 $l=7.05e-07 $layer=LI1_cond $X=6.895 $Y=3.33
+ $X2=6.19 $Y2=3.33
r161 35 38 32.7294 $w=2.48e-07 $l=7.1e-07 $layer=LI1_cond $X=6.065 $Y=2.105
+ $X2=6.065 $Y2=2.815
r162 33 89 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.065 $Y=3.245
+ $X2=6.065 $Y2=3.33
r163 33 38 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=6.065 $Y=3.245
+ $X2=6.065 $Y2=2.815
r164 29 86 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.155 $Y=3.245
+ $X2=4.155 $Y2=3.33
r165 29 31 18.3343 $w=3.28e-07 $l=5.25e-07 $layer=LI1_cond $X=4.155 $Y=3.245
+ $X2=4.155 $Y2=2.72
r166 25 83 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=2.19 $Y=3.245
+ $X2=2.19 $Y2=3.33
r167 25 27 23.2705 $w=2.58e-07 $l=5.25e-07 $layer=LI1_cond $X=2.19 $Y=3.245
+ $X2=2.19 $Y2=2.72
r168 21 24 32.7294 $w=2.48e-07 $l=7.1e-07 $layer=LI1_cond $X=0.255 $Y=2.105
+ $X2=0.255 $Y2=2.815
r169 19 80 3.1514 $w=2.5e-07 $l=1.12916e-07 $layer=LI1_cond $X=0.255 $Y=3.245
+ $X2=0.19 $Y2=3.33
r170 19 24 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=0.255 $Y=3.245
+ $X2=0.255 $Y2=2.815
r171 6 50 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=7.73
+ $Y=1.84 $X2=7.88 $Y2=2.815
r172 6 47 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=7.73
+ $Y=1.84 $X2=7.88 $Y2=1.985
r173 5 43 300 $w=1.7e-07 $l=5.80172e-07 $layer=licon1_PDIFF $count=2 $X=6.83
+ $Y=1.84 $X2=6.98 $Y2=2.35
r174 4 38 400 $w=1.7e-07 $l=9.26971e-07 $layer=licon1_PDIFF $count=1 $X=5.875
+ $Y=1.96 $X2=6.025 $Y2=2.815
r175 4 35 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=5.875
+ $Y=1.96 $X2=6.025 $Y2=2.105
r176 3 31 600 $w=1.7e-07 $l=8.54166e-07 $layer=licon1_PDIFF $count=1 $X=3.955
+ $Y=1.96 $X2=4.155 $Y2=2.72
r177 2 27 600 $w=1.7e-07 $l=8.33906e-07 $layer=licon1_PDIFF $count=1 $X=1.995
+ $Y=1.96 $X2=2.15 $Y2=2.72
r178 1 24 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=0.15
+ $Y=1.96 $X2=0.295 $Y2=2.815
r179 1 21 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.15
+ $Y=1.96 $X2=0.295 $Y2=2.105
.ends

.subckt PM_SKY130_FD_SC_HS__MAJ3_4%A_119_392# 1 2 9 11 12 15
r26 13 15 4.88915 $w=3.28e-07 $l=1.4e-07 $layer=LI1_cond $X=1.695 $Y=2.905
+ $X2=1.695 $Y2=2.765
r27 11 13 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.53 $Y=2.99
+ $X2=1.695 $Y2=2.905
r28 11 12 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=1.53 $Y=2.99
+ $X2=0.91 $Y2=2.99
r29 7 12 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.745 $Y=2.905
+ $X2=0.91 $Y2=2.99
r30 7 9 18.3343 $w=3.28e-07 $l=5.25e-07 $layer=LI1_cond $X=0.745 $Y=2.905
+ $X2=0.745 $Y2=2.38
r31 2 15 600 $w=1.7e-07 $l=8.76798e-07 $layer=licon1_PDIFF $count=1 $X=1.545
+ $Y=1.96 $X2=1.695 $Y2=2.765
r32 1 9 300 $w=1.7e-07 $l=4.89285e-07 $layer=licon1_PDIFF $count=2 $X=0.595
+ $Y=1.96 $X2=0.745 $Y2=2.38
.ends

.subckt PM_SKY130_FD_SC_HS__MAJ3_4%A_501_392# 1 2 9 11 12 15
r27 13 15 6.46067 $w=3.28e-07 $l=1.85e-07 $layer=LI1_cond $X=3.655 $Y=2.905
+ $X2=3.655 $Y2=2.72
r28 11 13 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.49 $Y=2.99
+ $X2=3.655 $Y2=2.905
r29 11 12 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.49 $Y=2.99
+ $X2=2.82 $Y2=2.99
r30 7 12 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.655 $Y=2.905
+ $X2=2.82 $Y2=2.99
r31 7 9 6.46067 $w=3.28e-07 $l=1.85e-07 $layer=LI1_cond $X=2.655 $Y=2.905
+ $X2=2.655 $Y2=2.72
r32 2 15 600 $w=1.7e-07 $l=8.54166e-07 $layer=licon1_PDIFF $count=1 $X=3.455
+ $Y=1.96 $X2=3.655 $Y2=2.72
r33 1 9 600 $w=1.7e-07 $l=8.31625e-07 $layer=licon1_PDIFF $count=1 $X=2.505
+ $Y=1.96 $X2=2.655 $Y2=2.72
.ends

.subckt PM_SKY130_FD_SC_HS__MAJ3_4%A_905_392# 1 2 7 9 14
c25 2 0 1.04924e-19 $X=5.425 $Y=1.96
r26 14 17 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=5.575 $Y=2.64 $X2=5.575
+ $Y2=2.72
r27 9 12 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=4.675 $Y=2.64 $X2=4.675
+ $Y2=2.72
r28 8 9 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.84 $Y=2.64 $X2=4.675
+ $Y2=2.64
r29 7 14 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.41 $Y=2.64
+ $X2=5.575 $Y2=2.64
r30 7 8 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=5.41 $Y=2.64 $X2=4.84
+ $Y2=2.64
r31 2 17 600 $w=1.7e-07 $l=8.31625e-07 $layer=licon1_PDIFF $count=1 $X=5.425
+ $Y=1.96 $X2=5.575 $Y2=2.72
r32 1 12 600 $w=1.7e-07 $l=8.31625e-07 $layer=licon1_PDIFF $count=1 $X=4.525
+ $Y=1.96 $X2=4.675 $Y2=2.72
.ends

.subckt PM_SKY130_FD_SC_HS__MAJ3_4%X 1 2 3 4 13 15 19 21 22 25 28 31 33 34 38 41
c59 19 0 3.37475e-19 $X=6.59 $Y=0.64
r60 40 41 9.26965 $w=2.28e-07 $l=1.85e-07 $layer=LI1_cond $X=7.92 $Y=1.48
+ $X2=7.92 $Y2=1.295
r61 39 41 6.01275 $w=2.28e-07 $l=1.2e-07 $layer=LI1_cond $X=7.92 $Y=1.175
+ $X2=7.92 $Y2=1.295
r62 33 40 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=7.805 $Y=1.565
+ $X2=7.92 $Y2=1.48
r63 33 34 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=7.805 $Y=1.565
+ $X2=7.515 $Y2=1.565
r64 29 38 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.43 $Y=2.015
+ $X2=7.43 $Y2=1.93
r65 29 31 52.1925 $w=1.68e-07 $l=8e-07 $layer=LI1_cond $X=7.43 $Y=2.015 $X2=7.43
+ $Y2=2.815
r66 28 38 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.43 $Y=1.845
+ $X2=7.43 $Y2=1.93
r67 27 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.43 $Y=1.65
+ $X2=7.515 $Y2=1.565
r68 27 28 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=7.43 $Y=1.65
+ $X2=7.43 $Y2=1.845
r69 26 36 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.695 $Y=1.93
+ $X2=6.53 $Y2=1.93
r70 25 38 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.345 $Y=1.93
+ $X2=7.43 $Y2=1.93
r71 25 26 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=7.345 $Y=1.93
+ $X2=6.695 $Y2=1.93
r72 22 24 50.5615 $w=1.68e-07 $l=7.75e-07 $layer=LI1_cond $X=6.675 $Y=1.09
+ $X2=7.45 $Y2=1.09
r73 21 39 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=7.805 $Y=1.09
+ $X2=7.92 $Y2=1.175
r74 21 24 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=7.805 $Y=1.09
+ $X2=7.45 $Y2=1.09
r75 17 22 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=6.55 $Y=1.005
+ $X2=6.675 $Y2=1.09
r76 17 19 16.8257 $w=2.48e-07 $l=3.65e-07 $layer=LI1_cond $X=6.55 $Y=1.005
+ $X2=6.55 $Y2=0.64
r77 13 36 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.53 $Y=2.015 $X2=6.53
+ $Y2=1.93
r78 13 15 27.938 $w=3.28e-07 $l=8e-07 $layer=LI1_cond $X=6.53 $Y=2.015 $X2=6.53
+ $Y2=2.815
r79 4 38 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=7.28
+ $Y=1.84 $X2=7.43 $Y2=1.985
r80 4 31 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=7.28
+ $Y=1.84 $X2=7.43 $Y2=2.815
r81 3 36 400 $w=1.7e-07 $l=2.33238e-07 $layer=licon1_PDIFF $count=1 $X=6.38
+ $Y=1.84 $X2=6.53 $Y2=2.01
r82 3 15 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=6.38
+ $Y=1.84 $X2=6.53 $Y2=2.815
r83 2 24 182 $w=1.7e-07 $l=6.61306e-07 $layer=licon1_NDIFF $count=1 $X=7.31
+ $Y=0.495 $X2=7.45 $Y2=1.09
r84 1 19 91 $w=1.7e-07 $l=2.41868e-07 $layer=licon1_NDIFF $count=2 $X=6.41
+ $Y=0.495 $X2=6.59 $Y2=0.64
.ends

.subckt PM_SKY130_FD_SC_HS__MAJ3_4%VGND 1 2 3 4 5 6 19 21 25 29 33 37 39 41 43
+ 45 50 55 60 65 74 77 80 83 87
r94 86 87 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=0 $X2=7.92
+ $Y2=0
r95 83 84 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=0 $X2=6.96
+ $Y2=0
r96 80 81 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6 $Y=0 $X2=6 $Y2=0
r97 74 75 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r98 71 72 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r99 69 87 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=0 $X2=7.92
+ $Y2=0
r100 69 84 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=0 $X2=6.96
+ $Y2=0
r101 68 69 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=0 $X2=7.44
+ $Y2=0
r102 66 83 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.185 $Y=0 $X2=7.02
+ $Y2=0
r103 66 68 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=7.185 $Y=0
+ $X2=7.44 $Y2=0
r104 65 86 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=7.715 $Y=0
+ $X2=7.937 $Y2=0
r105 65 68 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=7.715 $Y=0
+ $X2=7.44 $Y2=0
r106 64 84 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=0 $X2=6.96
+ $Y2=0
r107 64 81 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=0 $X2=6
+ $Y2=0
r108 63 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=0 $X2=6.48
+ $Y2=0
r109 61 80 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.205 $Y=0 $X2=6.08
+ $Y2=0
r110 61 63 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=6.205 $Y=0
+ $X2=6.48 $Y2=0
r111 60 83 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.855 $Y=0 $X2=7.02
+ $Y2=0
r112 60 63 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=6.855 $Y=0
+ $X2=6.48 $Y2=0
r113 59 81 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=4.56 $Y=0 $X2=6
+ $Y2=0
r114 58 59 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r115 56 77 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.335 $Y=0 $X2=4.17
+ $Y2=0
r116 56 58 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=4.335 $Y=0
+ $X2=4.56 $Y2=0
r117 55 80 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.955 $Y=0 $X2=6.08
+ $Y2=0
r118 55 58 91.0107 $w=1.68e-07 $l=1.395e-06 $layer=LI1_cond $X=5.955 $Y=0
+ $X2=4.56 $Y2=0
r119 54 75 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=2.16
+ $Y2=0
r120 53 54 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r121 51 74 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.315 $Y=0 $X2=2.23
+ $Y2=0
r122 51 53 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=2.315 $Y=0
+ $X2=2.64 $Y2=0
r123 50 77 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.005 $Y=0 $X2=4.17
+ $Y2=0
r124 50 53 89.0535 $w=1.68e-07 $l=1.365e-06 $layer=LI1_cond $X=4.005 $Y=0
+ $X2=2.64 $Y2=0
r125 49 75 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=0.72 $Y=0
+ $X2=2.16 $Y2=0
r126 49 72 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r127 48 49 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r128 46 71 4.73185 $w=1.7e-07 $l=2.23e-07 $layer=LI1_cond $X=0.445 $Y=0
+ $X2=0.222 $Y2=0
r129 46 48 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=0.445 $Y=0
+ $X2=0.72 $Y2=0
r130 45 74 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.145 $Y=0 $X2=2.23
+ $Y2=0
r131 45 48 92.9679 $w=1.68e-07 $l=1.425e-06 $layer=LI1_cond $X=2.145 $Y=0
+ $X2=0.72 $Y2=0
r132 43 59 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=4.56
+ $Y2=0
r133 43 54 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=4.08 $Y=0
+ $X2=2.64 $Y2=0
r134 43 77 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r135 39 86 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=7.88 $Y=0.085
+ $X2=7.937 $Y2=0
r136 39 41 20.4297 $w=3.28e-07 $l=5.85e-07 $layer=LI1_cond $X=7.88 $Y=0.085
+ $X2=7.88 $Y2=0.67
r137 35 83 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.02 $Y=0.085
+ $X2=7.02 $Y2=0
r138 35 37 20.4297 $w=3.28e-07 $l=5.85e-07 $layer=LI1_cond $X=7.02 $Y=0.085
+ $X2=7.02 $Y2=0.67
r139 31 80 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.08 $Y=0.085
+ $X2=6.08 $Y2=0
r140 31 33 25.5842 $w=2.48e-07 $l=5.55e-07 $layer=LI1_cond $X=6.08 $Y=0.085
+ $X2=6.08 $Y2=0.64
r141 27 77 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.17 $Y=0.085
+ $X2=4.17 $Y2=0
r142 27 29 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=4.17 $Y=0.085
+ $X2=4.17 $Y2=0.535
r143 23 74 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.23 $Y=0.085
+ $X2=2.23 $Y2=0
r144 23 25 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=2.23 $Y=0.085
+ $X2=2.23 $Y2=0.78
r145 19 71 3.03433 $w=3.3e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.28 $Y=0.085
+ $X2=0.222 $Y2=0
r146 19 21 23.9219 $w=3.28e-07 $l=6.85e-07 $layer=LI1_cond $X=0.28 $Y=0.085
+ $X2=0.28 $Y2=0.77
r147 6 41 182 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_NDIFF $count=1 $X=7.74
+ $Y=0.495 $X2=7.88 $Y2=0.67
r148 5 37 182 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_NDIFF $count=1 $X=6.88
+ $Y=0.495 $X2=7.02 $Y2=0.67
r149 4 33 91 $w=1.7e-07 $l=2.41454e-07 $layer=licon1_NDIFF $count=2 $X=5.9
+ $Y=0.595 $X2=6.12 $Y2=0.64
r150 3 29 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=4.03
+ $Y=0.39 $X2=4.17 $Y2=0.535
r151 2 25 182 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_NDIFF $count=1 $X=2.09
+ $Y=0.625 $X2=2.23 $Y2=0.78
r152 1 21 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.625 $X2=0.28 $Y2=0.77
.ends

.subckt PM_SKY130_FD_SC_HS__MAJ3_4%A_114_125# 1 2 7 11 13
r26 13 16 6.46067 $w=3.28e-07 $l=1.85e-07 $layer=LI1_cond $X=0.79 $Y=0.35
+ $X2=0.79 $Y2=0.535
r27 9 11 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=1.8 $Y=0.435 $X2=1.8
+ $Y2=0.78
r28 8 13 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.955 $Y=0.35
+ $X2=0.79 $Y2=0.35
r29 7 9 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.635 $Y=0.35
+ $X2=1.8 $Y2=0.435
r30 7 8 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.635 $Y=0.35
+ $X2=0.955 $Y2=0.35
r31 2 11 182 $w=1.7e-07 $l=2.76857e-07 $layer=licon1_NDIFF $count=1 $X=1.59
+ $Y=0.625 $X2=1.8 $Y2=0.78
r32 1 16 182 $w=1.7e-07 $l=2.61151e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.625 $X2=0.79 $Y2=0.535
.ends

.subckt PM_SKY130_FD_SC_HS__MAJ3_4%A_504_125# 1 2 9 11 12 13
r34 13 16 6.28605 $w=3.28e-07 $l=1.8e-07 $layer=LI1_cond $X=3.66 $Y=0.35
+ $X2=3.66 $Y2=0.53
r35 11 13 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.495 $Y=0.35
+ $X2=3.66 $Y2=0.35
r36 11 12 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=3.495 $Y=0.35
+ $X2=2.885 $Y2=0.35
r37 7 12 8.28377 $w=1.7e-07 $l=2.33666e-07 $layer=LI1_cond $X=2.69 $Y=0.435
+ $X2=2.885 $Y2=0.35
r38 7 9 9.89919 $w=3.88e-07 $l=3.35e-07 $layer=LI1_cond $X=2.69 $Y=0.435
+ $X2=2.69 $Y2=0.77
r39 2 16 182 $w=1.7e-07 $l=2.63249e-07 $layer=licon1_NDIFF $count=1 $X=3.44
+ $Y=0.625 $X2=3.66 $Y2=0.53
r40 1 9 182 $w=1.7e-07 $l=2.31409e-07 $layer=licon1_NDIFF $count=1 $X=2.52
+ $Y=0.625 $X2=2.69 $Y2=0.77
.ends

.subckt PM_SKY130_FD_SC_HS__MAJ3_4%A_906_78# 1 2 7 11 13
c30 13 0 1.46446e-19 $X=4.67 $Y=0.34
r31 13 16 6.80989 $w=3.28e-07 $l=1.95e-07 $layer=LI1_cond $X=4.67 $Y=0.34
+ $X2=4.67 $Y2=0.535
r32 9 11 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=5.61 $Y=0.425
+ $X2=5.61 $Y2=0.795
r33 8 13 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.835 $Y=0.34
+ $X2=4.67 $Y2=0.34
r34 7 9 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=5.445 $Y=0.34
+ $X2=5.61 $Y2=0.425
r35 7 8 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=5.445 $Y=0.34
+ $X2=4.835 $Y2=0.34
r36 2 11 182 $w=1.7e-07 $l=2.60768e-07 $layer=licon1_NDIFF $count=1 $X=5.47
+ $Y=0.595 $X2=5.61 $Y2=0.795
r37 1 16 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=4.53
+ $Y=0.39 $X2=4.67 $Y2=0.535
.ends

