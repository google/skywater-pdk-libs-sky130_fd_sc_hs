* File: sky130_fd_sc_hs__dfrbp_1.pxi.spice
* Created: Thu Aug 27 20:38:15 2020
* 
x_PM_SKY130_FD_SC_HS__DFRBP_1%D N_D_c_241_n N_D_M1000_g N_D_M1011_g N_D_c_242_n
+ D D D N_D_c_238_n N_D_c_239_n N_D_c_240_n PM_SKY130_FD_SC_HS__DFRBP_1%D
x_PM_SKY130_FD_SC_HS__DFRBP_1%RESET_B N_RESET_B_M1033_g N_RESET_B_c_269_n
+ N_RESET_B_c_277_n N_RESET_B_c_278_n N_RESET_B_M1001_g N_RESET_B_M1022_g
+ N_RESET_B_c_270_n N_RESET_B_c_280_n N_RESET_B_M1027_g N_RESET_B_M1030_g
+ N_RESET_B_c_282_n N_RESET_B_M1016_g N_RESET_B_c_272_n N_RESET_B_c_273_n
+ N_RESET_B_c_283_n N_RESET_B_c_284_n N_RESET_B_c_285_n N_RESET_B_c_286_n
+ N_RESET_B_c_287_n N_RESET_B_c_288_n RESET_B N_RESET_B_c_289_n
+ N_RESET_B_c_290_n N_RESET_B_c_274_n N_RESET_B_c_275_n N_RESET_B_c_292_n
+ N_RESET_B_c_293_n PM_SKY130_FD_SC_HS__DFRBP_1%RESET_B
x_PM_SKY130_FD_SC_HS__DFRBP_1%CLK N_CLK_c_459_n N_CLK_M1017_g N_CLK_M1002_g CLK
+ PM_SKY130_FD_SC_HS__DFRBP_1%CLK
x_PM_SKY130_FD_SC_HS__DFRBP_1%A_498_360# N_A_498_360#_M1013_d
+ N_A_498_360#_M1023_d N_A_498_360#_c_519_n N_A_498_360#_c_520_n
+ N_A_498_360#_M1021_g N_A_498_360#_c_502_n N_A_498_360#_c_503_n
+ N_A_498_360#_c_504_n N_A_498_360#_M1018_g N_A_498_360#_c_505_n
+ N_A_498_360#_M1007_g N_A_498_360#_c_506_n N_A_498_360#_c_507_n
+ N_A_498_360#_c_522_n N_A_498_360#_M1015_g N_A_498_360#_c_508_n
+ N_A_498_360#_c_509_n N_A_498_360#_c_510_n N_A_498_360#_c_523_n
+ N_A_498_360#_c_511_n N_A_498_360#_c_512_n N_A_498_360#_c_513_n
+ N_A_498_360#_c_546_p N_A_498_360#_c_572_p N_A_498_360#_c_514_n
+ N_A_498_360#_c_558_p N_A_498_360#_c_515_n N_A_498_360#_c_516_n
+ N_A_498_360#_c_535_n N_A_498_360#_c_526_n N_A_498_360#_c_517_n
+ N_A_498_360#_c_518_n PM_SKY130_FD_SC_HS__DFRBP_1%A_498_360#
x_PM_SKY130_FD_SC_HS__DFRBP_1%A_841_401# N_A_841_401#_M1004_d
+ N_A_841_401#_M1028_d N_A_841_401#_c_709_n N_A_841_401#_M1005_g
+ N_A_841_401#_M1006_g N_A_841_401#_c_710_n N_A_841_401#_c_701_n
+ N_A_841_401#_c_702_n N_A_841_401#_c_703_n N_A_841_401#_c_704_n
+ N_A_841_401#_c_705_n N_A_841_401#_c_706_n N_A_841_401#_c_707_n
+ N_A_841_401#_c_708_n N_A_841_401#_c_714_n
+ PM_SKY130_FD_SC_HS__DFRBP_1%A_841_401#
x_PM_SKY130_FD_SC_HS__DFRBP_1%A_706_463# N_A_706_463#_M1020_d
+ N_A_706_463#_M1021_d N_A_706_463#_M1027_d N_A_706_463#_M1004_g
+ N_A_706_463#_c_814_n N_A_706_463#_c_820_n N_A_706_463#_M1028_g
+ N_A_706_463#_c_815_n N_A_706_463#_c_833_n N_A_706_463#_c_822_n
+ N_A_706_463#_c_823_n N_A_706_463#_c_816_n N_A_706_463#_c_817_n
+ N_A_706_463#_c_818_n N_A_706_463#_c_825_n
+ PM_SKY130_FD_SC_HS__DFRBP_1%A_706_463#
x_PM_SKY130_FD_SC_HS__DFRBP_1%A_319_360# N_A_319_360#_M1002_s
+ N_A_319_360#_M1017_s N_A_319_360#_c_955_n N_A_319_360#_M1023_g
+ N_A_319_360#_c_942_n N_A_319_360#_M1013_g N_A_319_360#_c_943_n
+ N_A_319_360#_c_944_n N_A_319_360#_c_945_n N_A_319_360#_c_958_n
+ N_A_319_360#_c_959_n N_A_319_360#_M1020_g N_A_319_360#_c_960_n
+ N_A_319_360#_c_961_n N_A_319_360#_c_962_n N_A_319_360#_M1025_g
+ N_A_319_360#_c_963_n N_A_319_360#_c_964_n N_A_319_360#_c_965_n
+ N_A_319_360#_M1032_g N_A_319_360#_c_947_n N_A_319_360#_c_948_n
+ N_A_319_360#_M1003_g N_A_319_360#_c_969_n N_A_319_360#_c_950_n
+ N_A_319_360#_c_951_n N_A_319_360#_c_952_n N_A_319_360#_c_953_n
+ N_A_319_360#_c_954_n N_A_319_360#_c_971_n
+ PM_SKY130_FD_SC_HS__DFRBP_1%A_319_360#
x_PM_SKY130_FD_SC_HS__DFRBP_1%A_1482_48# N_A_1482_48#_M1031_d
+ N_A_1482_48#_M1016_d N_A_1482_48#_c_1132_n N_A_1482_48#_M1029_g
+ N_A_1482_48#_c_1133_n N_A_1482_48#_c_1141_n N_A_1482_48#_M1026_g
+ N_A_1482_48#_c_1134_n N_A_1482_48#_c_1142_n N_A_1482_48#_c_1135_n
+ N_A_1482_48#_c_1136_n N_A_1482_48#_c_1137_n N_A_1482_48#_c_1144_n
+ N_A_1482_48#_c_1138_n N_A_1482_48#_c_1139_n
+ PM_SKY130_FD_SC_HS__DFRBP_1%A_1482_48#
x_PM_SKY130_FD_SC_HS__DFRBP_1%A_1224_74# N_A_1224_74#_M1007_d
+ N_A_1224_74#_M1032_d N_A_1224_74#_M1031_g N_A_1224_74#_c_1228_n
+ N_A_1224_74#_c_1245_n N_A_1224_74#_M1019_g N_A_1224_74#_c_1229_n
+ N_A_1224_74#_c_1230_n N_A_1224_74#_c_1231_n N_A_1224_74#_M1024_g
+ N_A_1224_74#_M1014_g N_A_1224_74#_c_1233_n N_A_1224_74#_c_1234_n
+ N_A_1224_74#_c_1248_n N_A_1224_74#_M1008_g N_A_1224_74#_M1012_g
+ N_A_1224_74#_c_1236_n N_A_1224_74#_c_1277_n N_A_1224_74#_c_1257_n
+ N_A_1224_74#_c_1237_n N_A_1224_74#_c_1238_n N_A_1224_74#_c_1239_n
+ N_A_1224_74#_c_1240_n N_A_1224_74#_c_1241_n N_A_1224_74#_c_1242_n
+ N_A_1224_74#_c_1243_n PM_SKY130_FD_SC_HS__DFRBP_1%A_1224_74#
x_PM_SKY130_FD_SC_HS__DFRBP_1%A_2026_424# N_A_2026_424#_M1012_s
+ N_A_2026_424#_M1008_s N_A_2026_424#_M1009_g N_A_2026_424#_c_1392_n
+ N_A_2026_424#_M1010_g N_A_2026_424#_c_1393_n N_A_2026_424#_c_1394_n
+ N_A_2026_424#_c_1395_n N_A_2026_424#_c_1396_n
+ PM_SKY130_FD_SC_HS__DFRBP_1%A_2026_424#
x_PM_SKY130_FD_SC_HS__DFRBP_1%VPWR N_VPWR_M1000_s N_VPWR_M1001_d N_VPWR_M1017_d
+ N_VPWR_M1005_d N_VPWR_M1028_s N_VPWR_M1026_d N_VPWR_M1019_d N_VPWR_M1008_d
+ N_VPWR_c_1442_n N_VPWR_c_1443_n N_VPWR_c_1444_n N_VPWR_c_1445_n
+ N_VPWR_c_1446_n N_VPWR_c_1447_n N_VPWR_c_1448_n N_VPWR_c_1449_n
+ N_VPWR_c_1450_n N_VPWR_c_1451_n VPWR N_VPWR_c_1452_n N_VPWR_c_1453_n
+ N_VPWR_c_1454_n N_VPWR_c_1455_n N_VPWR_c_1456_n N_VPWR_c_1457_n
+ N_VPWR_c_1458_n N_VPWR_c_1441_n N_VPWR_c_1460_n N_VPWR_c_1461_n
+ N_VPWR_c_1462_n N_VPWR_c_1463_n N_VPWR_c_1464_n N_VPWR_c_1465_n
+ N_VPWR_c_1466_n PM_SKY130_FD_SC_HS__DFRBP_1%VPWR
x_PM_SKY130_FD_SC_HS__DFRBP_1%A_38_78# N_A_38_78#_M1011_s N_A_38_78#_M1020_s
+ N_A_38_78#_M1000_d N_A_38_78#_M1021_s N_A_38_78#_c_1581_n N_A_38_78#_c_1582_n
+ N_A_38_78#_c_1588_n N_A_38_78#_c_1583_n N_A_38_78#_c_1589_n
+ N_A_38_78#_c_1584_n N_A_38_78#_c_1585_n N_A_38_78#_c_1591_n
+ N_A_38_78#_c_1592_n N_A_38_78#_c_1586_n PM_SKY130_FD_SC_HS__DFRBP_1%A_38_78#
x_PM_SKY130_FD_SC_HS__DFRBP_1%Q_N N_Q_N_M1014_d N_Q_N_M1024_d N_Q_N_c_1691_n Q_N
+ Q_N Q_N N_Q_N_c_1694_n PM_SKY130_FD_SC_HS__DFRBP_1%Q_N
x_PM_SKY130_FD_SC_HS__DFRBP_1%Q N_Q_M1009_d N_Q_M1010_d Q Q Q Q Q N_Q_c_1717_n
+ PM_SKY130_FD_SC_HS__DFRBP_1%Q
x_PM_SKY130_FD_SC_HS__DFRBP_1%VGND N_VGND_M1033_d N_VGND_M1002_d N_VGND_M1022_d
+ N_VGND_M1029_d N_VGND_M1014_s N_VGND_M1012_d N_VGND_c_1738_n N_VGND_c_1739_n
+ N_VGND_c_1740_n N_VGND_c_1741_n N_VGND_c_1742_n N_VGND_c_1743_n VGND
+ N_VGND_c_1744_n N_VGND_c_1745_n N_VGND_c_1746_n N_VGND_c_1747_n
+ N_VGND_c_1748_n N_VGND_c_1749_n N_VGND_c_1750_n N_VGND_c_1751_n
+ N_VGND_c_1752_n N_VGND_c_1753_n N_VGND_c_1754_n N_VGND_c_1755_n
+ N_VGND_c_1756_n PM_SKY130_FD_SC_HS__DFRBP_1%VGND
cc_1 VNB N_D_M1011_g 0.0286427f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=0.6
cc_2 VNB N_D_c_238_n 0.0408539f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.845
cc_3 VNB N_D_c_239_n 0.0253354f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.165
cc_4 VNB N_D_c_240_n 0.0298264f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.165
cc_5 VNB N_RESET_B_M1033_g 0.0302438f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.75
cc_6 VNB N_RESET_B_c_269_n 0.0275049f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=0.6
cc_7 VNB N_RESET_B_c_270_n 0.0190115f $X=-0.19 $Y=-0.245 $X2=0.422 $Y2=1.845
cc_8 VNB N_RESET_B_M1030_g 0.0515393f $X=-0.19 $Y=-0.245 $X2=0.422 $Y2=1
cc_9 VNB N_RESET_B_c_272_n 0.0152827f $X=-0.19 $Y=-0.245 $X2=0.322 $Y2=1.665
cc_10 VNB N_RESET_B_c_273_n 0.0133173f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_RESET_B_c_274_n 0.0321958f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_RESET_B_c_275_n 0.00371377f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_CLK_c_459_n 0.026783f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.465
cc_14 VNB N_CLK_M1002_g 0.0265726f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=0.6
cc_15 VNB CLK 0.00502284f $X=-0.19 $Y=-0.245 $X2=0.422 $Y2=2.148
cc_16 VNB N_A_498_360#_c_502_n 0.0116282f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_498_360#_c_503_n 0.0167298f $X=-0.19 $Y=-0.245 $X2=0.422 $Y2=1.202
cc_18 VNB N_A_498_360#_c_504_n 0.0148131f $X=-0.19 $Y=-0.245 $X2=0.422 $Y2=1.845
cc_19 VNB N_A_498_360#_c_505_n 0.0205313f $X=-0.19 $Y=-0.245 $X2=0.422 $Y2=1.165
cc_20 VNB N_A_498_360#_c_506_n 0.0187502f $X=-0.19 $Y=-0.245 $X2=0.422 $Y2=1
cc_21 VNB N_A_498_360#_c_507_n 0.00880336f $X=-0.19 $Y=-0.245 $X2=0.322
+ $Y2=1.165
cc_22 VNB N_A_498_360#_c_508_n 0.0143796f $X=-0.19 $Y=-0.245 $X2=0.322 $Y2=1.845
cc_23 VNB N_A_498_360#_c_509_n 0.010555f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_498_360#_c_510_n 0.0403927f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_498_360#_c_511_n 0.00114194f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_498_360#_c_512_n 0.00349432f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_498_360#_c_513_n 0.00368177f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_498_360#_c_514_n 0.00621215f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_498_360#_c_515_n 0.0316981f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_498_360#_c_516_n 0.00782104f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_498_360#_c_517_n 0.0140979f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_498_360#_c_518_n 0.00789534f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_841_401#_M1006_g 0.0301498f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_841_401#_c_701_n 0.00632861f $X=-0.19 $Y=-0.245 $X2=0.422
+ $Y2=1.165
cc_35 VNB N_A_841_401#_c_702_n 0.015896f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.165
cc_36 VNB N_A_841_401#_c_703_n 0.0101533f $X=-0.19 $Y=-0.245 $X2=0.422 $Y2=1
cc_37 VNB N_A_841_401#_c_704_n 4.83161e-19 $X=-0.19 $Y=-0.245 $X2=0.322
+ $Y2=1.165
cc_38 VNB N_A_841_401#_c_705_n 4.96212e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_841_401#_c_706_n 0.00934369f $X=-0.19 $Y=-0.245 $X2=0.322
+ $Y2=1.295
cc_40 VNB N_A_841_401#_c_707_n 0.00496873f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_841_401#_c_708_n 4.11682e-19 $X=-0.19 $Y=-0.245 $X2=0.322
+ $Y2=1.665
cc_42 VNB N_A_706_463#_M1004_g 0.0294971f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_706_463#_c_814_n 0.0206988f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_706_463#_c_815_n 0.00364311f $X=-0.19 $Y=-0.245 $X2=0.385
+ $Y2=1.165
cc_45 VNB N_A_706_463#_c_816_n 0.00333952f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_A_706_463#_c_817_n 0.0104779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_706_463#_c_818_n 0.0286964f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_319_360#_c_942_n 0.018582f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_49 VNB N_A_319_360#_c_943_n 0.0036222f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_A_319_360#_c_944_n 0.0379132f $X=-0.19 $Y=-0.245 $X2=0.422 $Y2=1.202
cc_51 VNB N_A_319_360#_c_945_n 0.0627021f $X=-0.19 $Y=-0.245 $X2=0.422 $Y2=1.845
cc_52 VNB N_A_319_360#_M1020_g 0.0231068f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.165
cc_53 VNB N_A_319_360#_c_947_n 0.021569f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_A_319_360#_c_948_n 0.00563426f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_A_319_360#_M1003_g 0.0529012f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_A_319_360#_c_950_n 0.012043f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_A_319_360#_c_951_n 0.00908852f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_A_319_360#_c_952_n 0.00499474f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_A_319_360#_c_953_n 0.00330536f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_A_319_360#_c_954_n 0.00578626f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_A_1482_48#_c_1132_n 0.0177983f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_A_1482_48#_c_1133_n 0.0233363f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.95
cc_63 VNB N_A_1482_48#_c_1134_n 0.0157083f $X=-0.19 $Y=-0.245 $X2=0.422
+ $Y2=1.202
cc_64 VNB N_A_1482_48#_c_1135_n 0.0117659f $X=-0.19 $Y=-0.245 $X2=0.385
+ $Y2=1.165
cc_65 VNB N_A_1482_48#_c_1136_n 0.00518085f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_A_1482_48#_c_1137_n 0.00346875f $X=-0.19 $Y=-0.245 $X2=0.322
+ $Y2=1.295
cc_67 VNB N_A_1482_48#_c_1138_n 0.00600532f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_A_1482_48#_c_1139_n 0.0330587f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_A_1224_74#_M1031_g 0.0408739f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_70 VNB N_A_1224_74#_c_1228_n 0.00400132f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_A_1224_74#_c_1229_n 0.0327014f $X=-0.19 $Y=-0.245 $X2=0.422
+ $Y2=1.845
cc_72 VNB N_A_1224_74#_c_1230_n 0.0281282f $X=-0.19 $Y=-0.245 $X2=0.385
+ $Y2=1.845
cc_73 VNB N_A_1224_74#_c_1231_n 0.0364438f $X=-0.19 $Y=-0.245 $X2=0.385
+ $Y2=1.845
cc_74 VNB N_A_1224_74#_M1014_g 0.0260029f $X=-0.19 $Y=-0.245 $X2=0.322 $Y2=1.165
cc_75 VNB N_A_1224_74#_c_1233_n 0.0888375f $X=-0.19 $Y=-0.245 $X2=0.322
+ $Y2=1.295
cc_76 VNB N_A_1224_74#_c_1234_n 0.00400127f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_A_1224_74#_M1012_g 0.0355065f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_A_1224_74#_c_1236_n 0.0100839f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VNB N_A_1224_74#_c_1237_n 0.00749917f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_A_1224_74#_c_1238_n 0.0120508f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_81 VNB N_A_1224_74#_c_1239_n 4.69525e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_82 VNB N_A_1224_74#_c_1240_n 9.056e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_83 VNB N_A_1224_74#_c_1241_n 0.00965329f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_84 VNB N_A_1224_74#_c_1242_n 5.50055e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_85 VNB N_A_1224_74#_c_1243_n 0.00638783f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_86 VNB N_A_2026_424#_M1009_g 0.0282052f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_87 VNB N_A_2026_424#_c_1392_n 0.0344608f $X=-0.19 $Y=-0.245 $X2=0.155
+ $Y2=1.95
cc_88 VNB N_A_2026_424#_c_1393_n 0.00968545f $X=-0.19 $Y=-0.245 $X2=0.422
+ $Y2=1.845
cc_89 VNB N_A_2026_424#_c_1394_n 3.04122e-19 $X=-0.19 $Y=-0.245 $X2=0.385
+ $Y2=1.165
cc_90 VNB N_A_2026_424#_c_1395_n 0.00611923f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_91 VNB N_A_2026_424#_c_1396_n 3.73161e-19 $X=-0.19 $Y=-0.245 $X2=0.322
+ $Y2=1.665
cc_92 VNB N_VPWR_c_1441_n 0.48212f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_93 VNB N_A_38_78#_c_1581_n 0.00234225f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_94 VNB N_A_38_78#_c_1582_n 0.0151449f $X=-0.19 $Y=-0.245 $X2=0.422 $Y2=1.845
cc_95 VNB N_A_38_78#_c_1583_n 0.00135826f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.165
cc_96 VNB N_A_38_78#_c_1584_n 0.00432348f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_97 VNB N_A_38_78#_c_1585_n 0.0222631f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_98 VNB N_A_38_78#_c_1586_n 0.0065782f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_99 VNB N_Q_N_c_1691_n 0.0157896f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_100 VNB Q 0.0267746f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_101 VNB Q 0.0133985f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_102 VNB N_Q_c_1717_n 0.0249767f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_103 VNB N_VGND_c_1738_n 0.0129144f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.165
cc_104 VNB N_VGND_c_1739_n 0.0222124f $X=-0.19 $Y=-0.245 $X2=0.322 $Y2=1.165
cc_105 VNB N_VGND_c_1740_n 0.0093032f $X=-0.19 $Y=-0.245 $X2=0.322 $Y2=1.665
cc_106 VNB N_VGND_c_1741_n 0.00450041f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_107 VNB N_VGND_c_1742_n 0.00944343f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_108 VNB N_VGND_c_1743_n 0.0125104f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_109 VNB N_VGND_c_1744_n 0.0309201f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_110 VNB N_VGND_c_1745_n 0.0613f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_111 VNB N_VGND_c_1746_n 0.0603291f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_112 VNB N_VGND_c_1747_n 0.0324414f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_113 VNB N_VGND_c_1748_n 0.0347338f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_114 VNB N_VGND_c_1749_n 0.0191572f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_115 VNB N_VGND_c_1750_n 0.64872f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_116 VNB N_VGND_c_1751_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_117 VNB N_VGND_c_1752_n 0.00634414f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_118 VNB N_VGND_c_1753_n 0.0158757f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_119 VNB N_VGND_c_1754_n 0.00846888f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_120 VNB N_VGND_c_1755_n 0.00461913f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_121 VNB N_VGND_c_1756_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_122 VPB N_D_c_241_n 0.0179054f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.465
cc_123 VPB N_D_c_242_n 0.0399063f $X=-0.19 $Y=1.66 $X2=0.422 $Y2=2.148
cc_124 VPB N_D_c_238_n 0.0435358f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.845
cc_125 VPB N_D_c_240_n 0.0215212f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.165
cc_126 VPB N_RESET_B_c_269_n 0.0234437f $X=-0.19 $Y=1.66 $X2=0.55 $Y2=0.6
cc_127 VPB N_RESET_B_c_277_n 0.0179996f $X=-0.19 $Y=1.66 $X2=0.422 $Y2=2.148
cc_128 VPB N_RESET_B_c_278_n 0.0242054f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.21
cc_129 VPB N_RESET_B_c_270_n 0.0124021f $X=-0.19 $Y=1.66 $X2=0.422 $Y2=1.845
cc_130 VPB N_RESET_B_c_280_n 0.0192017f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.845
cc_131 VPB N_RESET_B_M1030_g 0.00974243f $X=-0.19 $Y=1.66 $X2=0.422 $Y2=1
cc_132 VPB N_RESET_B_c_282_n 0.052471f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_133 VPB N_RESET_B_c_283_n 0.0189222f $X=-0.19 $Y=1.66 $X2=0.322 $Y2=2.035
cc_134 VPB N_RESET_B_c_284_n 0.0277677f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_135 VPB N_RESET_B_c_285_n 0.00343269f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_136 VPB N_RESET_B_c_286_n 0.00537181f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_137 VPB N_RESET_B_c_287_n 0.00350644f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_138 VPB N_RESET_B_c_288_n 0.00338092f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_139 VPB N_RESET_B_c_289_n 0.0554752f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_140 VPB N_RESET_B_c_290_n 0.00383188f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_141 VPB N_RESET_B_c_275_n 9.2757e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_142 VPB N_RESET_B_c_292_n 0.0291504f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_143 VPB N_RESET_B_c_293_n 0.00608672f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_144 VPB N_CLK_c_459_n 0.0278698f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.465
cc_145 VPB CLK 0.00526029f $X=-0.19 $Y=1.66 $X2=0.422 $Y2=2.148
cc_146 VPB N_A_498_360#_c_519_n 0.0150349f $X=-0.19 $Y=1.66 $X2=0.422 $Y2=2.148
cc_147 VPB N_A_498_360#_c_520_n 0.0192995f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.21
cc_148 VPB N_A_498_360#_c_502_n 0.0203903f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_149 VPB N_A_498_360#_c_522_n 0.0569971f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_150 VPB N_A_498_360#_c_523_n 0.00670952f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_151 VPB N_A_498_360#_c_511_n 7.52671e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_152 VPB N_A_498_360#_c_516_n 0.0024834f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_153 VPB N_A_498_360#_c_526_n 0.00306084f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_154 VPB N_A_498_360#_c_518_n 0.0207328f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_155 VPB N_A_841_401#_c_709_n 0.0144605f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_156 VPB N_A_841_401#_c_710_n 0.0554176f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_157 VPB N_A_841_401#_c_701_n 0.0026876f $X=-0.19 $Y=1.66 $X2=0.422 $Y2=1.165
cc_158 VPB N_A_841_401#_c_702_n 0.00209419f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.165
cc_159 VPB N_A_841_401#_c_707_n 6.92353e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_160 VPB N_A_841_401#_c_714_n 0.00398554f $X=-0.19 $Y=1.66 $X2=0.322 $Y2=2.035
cc_161 VPB N_A_706_463#_c_814_n 0.0214001f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_162 VPB N_A_706_463#_c_820_n 0.0168657f $X=-0.19 $Y=1.66 $X2=0.422 $Y2=1.845
cc_163 VPB N_A_706_463#_c_815_n 0.00977738f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.165
cc_164 VPB N_A_706_463#_c_822_n 0.00239542f $X=-0.19 $Y=1.66 $X2=0.422 $Y2=1
cc_165 VPB N_A_706_463#_c_823_n 0.0104778f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_166 VPB N_A_706_463#_c_818_n 3.30851e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_167 VPB N_A_706_463#_c_825_n 0.00486691f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_168 VPB N_A_319_360#_c_955_n 0.0144896f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_169 VPB N_A_319_360#_c_943_n 0.0795561f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_170 VPB N_A_319_360#_c_945_n 0.00692409f $X=-0.19 $Y=1.66 $X2=0.422 $Y2=1.845
cc_171 VPB N_A_319_360#_c_958_n 0.0555942f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.845
cc_172 VPB N_A_319_360#_c_959_n 0.0125859f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.845
cc_173 VPB N_A_319_360#_c_960_n 0.00711139f $X=-0.19 $Y=1.66 $X2=0.322 $Y2=1.165
cc_174 VPB N_A_319_360#_c_961_n 0.0163876f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_175 VPB N_A_319_360#_c_962_n 0.0142197f $X=-0.19 $Y=1.66 $X2=0.322 $Y2=1.295
cc_176 VPB N_A_319_360#_c_963_n 0.200784f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_177 VPB N_A_319_360#_c_964_n 0.00738389f $X=-0.19 $Y=1.66 $X2=0.322 $Y2=2.035
cc_178 VPB N_A_319_360#_c_965_n 0.0161081f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_179 VPB N_A_319_360#_M1032_g 0.00837835f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_180 VPB N_A_319_360#_c_947_n 0.0142262f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_181 VPB N_A_319_360#_c_948_n 0.00505238f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_182 VPB N_A_319_360#_c_969_n 0.0089864f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_183 VPB N_A_319_360#_c_951_n 0.00397652f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_184 VPB N_A_319_360#_c_971_n 0.00442119f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_185 VPB N_A_1482_48#_c_1133_n 0.0272407f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.95
cc_186 VPB N_A_1482_48#_c_1141_n 0.0213103f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_187 VPB N_A_1482_48#_c_1142_n 0.0103983f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.845
cc_188 VPB N_A_1482_48#_c_1136_n 0.00239847f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_189 VPB N_A_1482_48#_c_1144_n 0.00655902f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_190 VPB N_A_1224_74#_c_1228_n 0.0278194f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_191 VPB N_A_1224_74#_c_1245_n 0.021316f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_192 VPB N_A_1224_74#_c_1231_n 0.0280594f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.845
cc_193 VPB N_A_1224_74#_c_1234_n 0.0203227f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_194 VPB N_A_1224_74#_c_1248_n 0.0278562f $X=-0.19 $Y=1.66 $X2=0.322 $Y2=1.845
cc_195 VPB N_A_1224_74#_c_1240_n 0.00656652f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_196 VPB N_A_2026_424#_c_1392_n 0.0290451f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.95
cc_197 VPB N_A_2026_424#_c_1394_n 0.00753336f $X=-0.19 $Y=1.66 $X2=0.385
+ $Y2=1.165
cc_198 VPB N_VPWR_c_1442_n 0.0106521f $X=-0.19 $Y=1.66 $X2=0.322 $Y2=1.295
cc_199 VPB N_VPWR_c_1443_n 0.0314176f $X=-0.19 $Y=1.66 $X2=0.322 $Y2=1.665
cc_200 VPB N_VPWR_c_1444_n 0.0150499f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_201 VPB N_VPWR_c_1445_n 0.00605696f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_202 VPB N_VPWR_c_1446_n 0.013849f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_203 VPB N_VPWR_c_1447_n 0.0156795f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_204 VPB N_VPWR_c_1448_n 0.0249508f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_205 VPB N_VPWR_c_1449_n 0.021993f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_206 VPB N_VPWR_c_1450_n 0.0118234f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_207 VPB N_VPWR_c_1451_n 0.0143642f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_208 VPB N_VPWR_c_1452_n 0.0205885f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_209 VPB N_VPWR_c_1453_n 0.0215753f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_210 VPB N_VPWR_c_1454_n 0.0602093f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_211 VPB N_VPWR_c_1455_n 0.0273297f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_212 VPB N_VPWR_c_1456_n 0.0507873f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_213 VPB N_VPWR_c_1457_n 0.0430282f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_214 VPB N_VPWR_c_1458_n 0.0189171f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_215 VPB N_VPWR_c_1441_n 0.127213f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_216 VPB N_VPWR_c_1460_n 0.0047828f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_217 VPB N_VPWR_c_1461_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_218 VPB N_VPWR_c_1462_n 0.00456739f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_219 VPB N_VPWR_c_1463_n 0.00330333f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_220 VPB N_VPWR_c_1464_n 0.00430193f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_221 VPB N_VPWR_c_1465_n 0.00410958f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_222 VPB N_VPWR_c_1466_n 0.00564836f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_223 VPB N_A_38_78#_c_1582_n 0.0107742f $X=-0.19 $Y=1.66 $X2=0.422 $Y2=1.845
cc_224 VPB N_A_38_78#_c_1588_n 0.0176488f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.845
cc_225 VPB N_A_38_78#_c_1589_n 0.00661138f $X=-0.19 $Y=1.66 $X2=0.322 $Y2=1.165
cc_226 VPB N_A_38_78#_c_1584_n 0.00548757f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_227 VPB N_A_38_78#_c_1591_n 0.00798703f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_228 VPB N_A_38_78#_c_1592_n 0.00917021f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_229 VPB N_Q_N_c_1691_n 0.00323856f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.21
cc_230 VPB Q_N 0.0168178f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_231 VPB N_Q_N_c_1694_n 0.00844312f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_232 VPB Q 0.0131162f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.95
cc_233 VPB Q 0.041687f $X=-0.19 $Y=1.66 $X2=0.322 $Y2=1.665
cc_234 VPB N_Q_c_1717_n 0.00776073f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_235 N_D_M1011_g N_RESET_B_M1033_g 0.0258218f $X=0.55 $Y=0.6 $X2=0 $Y2=0
cc_236 N_D_c_238_n N_RESET_B_c_269_n 0.0258218f $X=0.385 $Y=1.845 $X2=0 $Y2=0
cc_237 N_D_c_242_n N_RESET_B_c_277_n 0.00488452f $X=0.422 $Y=2.148 $X2=0 $Y2=0
cc_238 N_D_c_241_n N_RESET_B_c_278_n 0.00917787f $X=0.505 $Y=2.465 $X2=0 $Y2=0
cc_239 N_D_c_239_n N_RESET_B_c_274_n 0.0258218f $X=0.385 $Y=1.165 $X2=0 $Y2=0
cc_240 N_D_c_242_n N_RESET_B_c_292_n 0.0258218f $X=0.422 $Y=2.148 $X2=0 $Y2=0
cc_241 N_D_c_241_n N_VPWR_c_1443_n 0.00729224f $X=0.505 $Y=2.465 $X2=0 $Y2=0
cc_242 N_D_c_242_n N_VPWR_c_1443_n 0.0042702f $X=0.422 $Y=2.148 $X2=0 $Y2=0
cc_243 N_D_c_240_n N_VPWR_c_1443_n 0.013492f $X=0.385 $Y=1.165 $X2=0 $Y2=0
cc_244 N_D_c_241_n N_VPWR_c_1452_n 0.00444469f $X=0.505 $Y=2.465 $X2=0 $Y2=0
cc_245 N_D_c_241_n N_VPWR_c_1441_n 0.00857499f $X=0.505 $Y=2.465 $X2=0 $Y2=0
cc_246 N_D_c_242_n N_VPWR_c_1441_n 3.7828e-19 $X=0.422 $Y=2.148 $X2=0 $Y2=0
cc_247 N_D_M1011_g N_A_38_78#_c_1581_n 0.0116103f $X=0.55 $Y=0.6 $X2=0 $Y2=0
cc_248 N_D_c_240_n N_A_38_78#_c_1581_n 0.00144733f $X=0.385 $Y=1.165 $X2=0 $Y2=0
cc_249 N_D_M1011_g N_A_38_78#_c_1582_n 0.0152564f $X=0.55 $Y=0.6 $X2=0 $Y2=0
cc_250 N_D_c_240_n N_A_38_78#_c_1582_n 0.0904243f $X=0.385 $Y=1.165 $X2=0 $Y2=0
cc_251 N_D_M1011_g N_A_38_78#_c_1585_n 0.0078958f $X=0.55 $Y=0.6 $X2=0 $Y2=0
cc_252 N_D_c_239_n N_A_38_78#_c_1585_n 0.00191909f $X=0.385 $Y=1.165 $X2=0 $Y2=0
cc_253 N_D_c_240_n N_A_38_78#_c_1585_n 0.028486f $X=0.385 $Y=1.165 $X2=0 $Y2=0
cc_254 N_D_c_241_n N_A_38_78#_c_1591_n 0.00810441f $X=0.505 $Y=2.465 $X2=0 $Y2=0
cc_255 N_D_c_242_n N_A_38_78#_c_1591_n 0.00689915f $X=0.422 $Y=2.148 $X2=0 $Y2=0
cc_256 N_D_M1011_g N_VGND_c_1744_n 0.00429844f $X=0.55 $Y=0.6 $X2=0 $Y2=0
cc_257 N_D_M1011_g N_VGND_c_1750_n 0.00539454f $X=0.55 $Y=0.6 $X2=0 $Y2=0
cc_258 N_RESET_B_c_269_n N_CLK_c_459_n 0.00558152f $X=1.097 $Y=1.908 $X2=-0.19
+ $Y2=-0.245
cc_259 N_RESET_B_c_284_n N_CLK_c_459_n 0.00512823f $X=5.375 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_260 N_RESET_B_c_274_n N_CLK_c_459_n 0.00656816f $X=1.165 $Y=1.295 $X2=-0.19
+ $Y2=-0.245
cc_261 N_RESET_B_c_274_n N_CLK_M1002_g 0.00246398f $X=1.165 $Y=1.295 $X2=0 $Y2=0
cc_262 N_RESET_B_c_284_n CLK 0.0124675f $X=5.375 $Y=2.035 $X2=0 $Y2=0
cc_263 N_RESET_B_c_284_n N_A_498_360#_c_519_n 0.00396118f $X=5.375 $Y=2.035
+ $X2=0 $Y2=0
cc_264 N_RESET_B_c_284_n N_A_498_360#_c_502_n 0.00522086f $X=5.375 $Y=2.035
+ $X2=0 $Y2=0
cc_265 N_RESET_B_c_286_n N_A_498_360#_c_522_n 0.00152844f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_266 N_RESET_B_c_284_n N_A_498_360#_c_523_n 0.0311928f $X=5.375 $Y=2.035 $X2=0
+ $Y2=0
cc_267 N_RESET_B_c_284_n N_A_498_360#_c_511_n 0.0105554f $X=5.375 $Y=2.035 $X2=0
+ $Y2=0
cc_268 N_RESET_B_c_272_n N_A_498_360#_c_512_n 7.29156e-19 $X=4.89 $Y=1.085 $X2=0
+ $Y2=0
cc_269 N_RESET_B_c_272_n N_A_498_360#_c_513_n 0.0112129f $X=4.89 $Y=1.085 $X2=0
+ $Y2=0
cc_270 N_RESET_B_c_286_n N_A_498_360#_c_535_n 0.0123453f $X=7.775 $Y=2.035 $X2=0
+ $Y2=0
cc_271 N_RESET_B_c_286_n N_A_498_360#_c_526_n 0.0237639f $X=7.775 $Y=2.035 $X2=0
+ $Y2=0
cc_272 N_RESET_B_c_284_n N_A_498_360#_c_518_n 0.0038641f $X=5.375 $Y=2.035 $X2=0
+ $Y2=0
cc_273 N_RESET_B_c_286_n N_A_841_401#_M1028_d 0.00313731f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_274 N_RESET_B_c_280_n N_A_841_401#_c_709_n 0.013563f $X=4.93 $Y=2.24 $X2=0
+ $Y2=0
cc_275 N_RESET_B_c_270_n N_A_841_401#_M1006_g 0.00971829f $X=4.915 $Y=1.825
+ $X2=0 $Y2=0
cc_276 N_RESET_B_c_272_n N_A_841_401#_M1006_g 0.0416068f $X=4.89 $Y=1.085 $X2=0
+ $Y2=0
cc_277 N_RESET_B_c_283_n N_A_841_401#_c_710_n 0.0230883f $X=4.93 $Y=2.032 $X2=0
+ $Y2=0
cc_278 N_RESET_B_c_284_n N_A_841_401#_c_710_n 0.00672549f $X=5.375 $Y=2.035
+ $X2=0 $Y2=0
cc_279 N_RESET_B_c_270_n N_A_841_401#_c_701_n 0.00534914f $X=4.915 $Y=1.825
+ $X2=0 $Y2=0
cc_280 N_RESET_B_c_273_n N_A_841_401#_c_701_n 0.00329036f $X=4.89 $Y=1.235 $X2=0
+ $Y2=0
cc_281 N_RESET_B_c_284_n N_A_841_401#_c_701_n 0.0258991f $X=5.375 $Y=2.035 $X2=0
+ $Y2=0
cc_282 N_RESET_B_c_270_n N_A_841_401#_c_702_n 0.0210965f $X=4.915 $Y=1.825 $X2=0
+ $Y2=0
cc_283 N_RESET_B_c_272_n N_A_841_401#_c_703_n 0.00865825f $X=4.89 $Y=1.085 $X2=0
+ $Y2=0
cc_284 N_RESET_B_c_273_n N_A_841_401#_c_703_n 0.00713061f $X=4.89 $Y=1.235 $X2=0
+ $Y2=0
cc_285 N_RESET_B_c_286_n N_A_841_401#_c_707_n 0.0067544f $X=7.775 $Y=2.035 $X2=0
+ $Y2=0
cc_286 N_RESET_B_c_286_n N_A_841_401#_c_708_n 0.00201833f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_287 N_RESET_B_c_286_n N_A_841_401#_c_714_n 0.0328549f $X=7.775 $Y=2.035 $X2=0
+ $Y2=0
cc_288 N_RESET_B_c_272_n N_A_706_463#_M1004_g 0.0177824f $X=4.89 $Y=1.085 $X2=0
+ $Y2=0
cc_289 N_RESET_B_c_273_n N_A_706_463#_M1004_g 0.0075767f $X=4.89 $Y=1.235 $X2=0
+ $Y2=0
cc_290 N_RESET_B_c_286_n N_A_706_463#_c_814_n 0.00249739f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_291 N_RESET_B_c_287_n N_A_706_463#_c_814_n 0.00116431f $X=5.665 $Y=2.035
+ $X2=0 $Y2=0
cc_292 N_RESET_B_c_290_n N_A_706_463#_c_814_n 0.0017604f $X=5.395 $Y=1.99 $X2=0
+ $Y2=0
cc_293 N_RESET_B_c_286_n N_A_706_463#_c_820_n 0.0069988f $X=7.775 $Y=2.035 $X2=0
+ $Y2=0
cc_294 N_RESET_B_c_284_n N_A_706_463#_c_815_n 0.0215965f $X=5.375 $Y=2.035 $X2=0
+ $Y2=0
cc_295 N_RESET_B_c_280_n N_A_706_463#_c_833_n 0.00472575f $X=4.93 $Y=2.24 $X2=0
+ $Y2=0
cc_296 N_RESET_B_c_284_n N_A_706_463#_c_833_n 0.0175481f $X=5.375 $Y=2.035 $X2=0
+ $Y2=0
cc_297 N_RESET_B_c_284_n N_A_706_463#_c_822_n 0.00764153f $X=5.375 $Y=2.035
+ $X2=0 $Y2=0
cc_298 N_RESET_B_c_270_n N_A_706_463#_c_823_n 0.00710021f $X=4.915 $Y=1.825
+ $X2=0 $Y2=0
cc_299 N_RESET_B_c_280_n N_A_706_463#_c_823_n 0.0043958f $X=4.93 $Y=2.24 $X2=0
+ $Y2=0
cc_300 N_RESET_B_c_283_n N_A_706_463#_c_823_n 0.0106103f $X=4.93 $Y=2.032 $X2=0
+ $Y2=0
cc_301 N_RESET_B_c_284_n N_A_706_463#_c_823_n 0.0226098f $X=5.375 $Y=2.035 $X2=0
+ $Y2=0
cc_302 N_RESET_B_c_287_n N_A_706_463#_c_823_n 4.39853e-19 $X=5.665 $Y=2.035
+ $X2=0 $Y2=0
cc_303 N_RESET_B_c_289_n N_A_706_463#_c_823_n 0.00639141f $X=5.395 $Y=1.99 $X2=0
+ $Y2=0
cc_304 N_RESET_B_c_290_n N_A_706_463#_c_823_n 0.0224281f $X=5.395 $Y=1.99 $X2=0
+ $Y2=0
cc_305 N_RESET_B_c_270_n N_A_706_463#_c_817_n 0.0074551f $X=4.915 $Y=1.825 $X2=0
+ $Y2=0
cc_306 N_RESET_B_c_284_n N_A_706_463#_c_817_n 0.00666358f $X=5.375 $Y=2.035
+ $X2=0 $Y2=0
cc_307 N_RESET_B_c_287_n N_A_706_463#_c_817_n 0.00107679f $X=5.665 $Y=2.035
+ $X2=0 $Y2=0
cc_308 N_RESET_B_c_289_n N_A_706_463#_c_817_n 0.00728227f $X=5.395 $Y=1.99 $X2=0
+ $Y2=0
cc_309 N_RESET_B_c_290_n N_A_706_463#_c_817_n 0.0190365f $X=5.395 $Y=1.99 $X2=0
+ $Y2=0
cc_310 N_RESET_B_c_270_n N_A_706_463#_c_818_n 0.0174208f $X=4.915 $Y=1.825 $X2=0
+ $Y2=0
cc_311 N_RESET_B_c_289_n N_A_706_463#_c_818_n 0.0207972f $X=5.395 $Y=1.99 $X2=0
+ $Y2=0
cc_312 N_RESET_B_c_290_n N_A_706_463#_c_818_n 4.14991e-19 $X=5.395 $Y=1.99 $X2=0
+ $Y2=0
cc_313 N_RESET_B_c_280_n N_A_706_463#_c_825_n 0.00782859f $X=4.93 $Y=2.24 $X2=0
+ $Y2=0
cc_314 N_RESET_B_c_284_n N_A_706_463#_c_825_n 0.00769568f $X=5.375 $Y=2.035
+ $X2=0 $Y2=0
cc_315 N_RESET_B_c_289_n N_A_706_463#_c_825_n 0.00879621f $X=5.395 $Y=1.99 $X2=0
+ $Y2=0
cc_316 N_RESET_B_c_290_n N_A_706_463#_c_825_n 0.00602228f $X=5.395 $Y=1.99 $X2=0
+ $Y2=0
cc_317 N_RESET_B_c_284_n N_A_319_360#_M1017_s 0.00113357f $X=5.375 $Y=2.035
+ $X2=0 $Y2=0
cc_318 N_RESET_B_c_284_n N_A_319_360#_c_955_n 0.00711303f $X=5.375 $Y=2.035
+ $X2=0 $Y2=0
cc_319 N_RESET_B_c_284_n N_A_319_360#_c_943_n 0.00517522f $X=5.375 $Y=2.035
+ $X2=0 $Y2=0
cc_320 N_RESET_B_c_284_n N_A_319_360#_c_945_n 3.7969e-19 $X=5.375 $Y=2.035 $X2=0
+ $Y2=0
cc_321 N_RESET_B_c_284_n N_A_319_360#_c_962_n 0.00238834f $X=5.375 $Y=2.035
+ $X2=0 $Y2=0
cc_322 N_RESET_B_c_280_n N_A_319_360#_c_963_n 0.00992461f $X=4.93 $Y=2.24 $X2=0
+ $Y2=0
cc_323 N_RESET_B_c_286_n N_A_319_360#_M1032_g 0.0118743f $X=7.775 $Y=2.035 $X2=0
+ $Y2=0
cc_324 N_RESET_B_c_286_n N_A_319_360#_c_947_n 3.83564e-19 $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_325 N_RESET_B_c_286_n N_A_319_360#_c_948_n 3.03408e-19 $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_326 N_RESET_B_M1033_g N_A_319_360#_c_950_n 0.00331172f $X=0.94 $Y=0.6 $X2=0
+ $Y2=0
cc_327 N_RESET_B_c_284_n N_A_319_360#_c_951_n 8.85602e-19 $X=5.375 $Y=2.035
+ $X2=0 $Y2=0
cc_328 N_RESET_B_c_274_n N_A_319_360#_c_951_n 0.00664799f $X=1.165 $Y=1.295
+ $X2=0 $Y2=0
cc_329 N_RESET_B_c_275_n N_A_319_360#_c_951_n 0.0495178f $X=1.165 $Y=1.295 $X2=0
+ $Y2=0
cc_330 N_RESET_B_c_284_n N_A_319_360#_c_953_n 0.00239237f $X=5.375 $Y=2.035
+ $X2=0 $Y2=0
cc_331 N_RESET_B_M1033_g N_A_319_360#_c_954_n 0.00289085f $X=0.94 $Y=0.6 $X2=0
+ $Y2=0
cc_332 N_RESET_B_c_275_n N_A_319_360#_c_954_n 8.31882e-19 $X=1.165 $Y=1.295
+ $X2=0 $Y2=0
cc_333 N_RESET_B_c_269_n N_A_319_360#_c_971_n 0.0030016f $X=1.097 $Y=1.908 $X2=0
+ $Y2=0
cc_334 N_RESET_B_c_284_n N_A_319_360#_c_971_n 0.0235177f $X=5.375 $Y=2.035 $X2=0
+ $Y2=0
cc_335 N_RESET_B_c_285_n N_A_319_360#_c_971_n 0.00241767f $X=1.345 $Y=2.035
+ $X2=0 $Y2=0
cc_336 N_RESET_B_c_275_n N_A_319_360#_c_971_n 0.0234848f $X=1.165 $Y=1.295 $X2=0
+ $Y2=0
cc_337 N_RESET_B_M1030_g N_A_1482_48#_c_1132_n 0.0196155f $X=8.045 $Y=0.58 $X2=0
+ $Y2=0
cc_338 N_RESET_B_c_282_n N_A_1482_48#_c_1133_n 0.044692f $X=8.18 $Y=2.28 $X2=0
+ $Y2=0
cc_339 N_RESET_B_c_286_n N_A_1482_48#_c_1133_n 0.00564012f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_340 N_RESET_B_c_288_n N_A_1482_48#_c_1133_n 0.00149248f $X=7.92 $Y=2.035
+ $X2=0 $Y2=0
cc_341 N_RESET_B_c_293_n N_A_1482_48#_c_1133_n 0.00190186f $X=8.135 $Y=2 $X2=0
+ $Y2=0
cc_342 N_RESET_B_c_282_n N_A_1482_48#_c_1141_n 0.00623945f $X=8.18 $Y=2.28 $X2=0
+ $Y2=0
cc_343 N_RESET_B_M1030_g N_A_1482_48#_c_1134_n 0.0144302f $X=8.045 $Y=0.58 $X2=0
+ $Y2=0
cc_344 N_RESET_B_c_282_n N_A_1482_48#_c_1142_n 0.00528461f $X=8.18 $Y=2.28 $X2=0
+ $Y2=0
cc_345 N_RESET_B_c_288_n N_A_1482_48#_c_1142_n 9.35982e-19 $X=7.92 $Y=2.035
+ $X2=0 $Y2=0
cc_346 N_RESET_B_c_293_n N_A_1482_48#_c_1142_n 0.0201792f $X=8.135 $Y=2 $X2=0
+ $Y2=0
cc_347 N_RESET_B_M1030_g N_A_1482_48#_c_1135_n 0.00201284f $X=8.045 $Y=0.58
+ $X2=0 $Y2=0
cc_348 N_RESET_B_M1030_g N_A_1482_48#_c_1137_n 0.00118187f $X=8.045 $Y=0.58
+ $X2=0 $Y2=0
cc_349 N_RESET_B_M1030_g N_A_1482_48#_c_1144_n 0.00150115f $X=8.045 $Y=0.58
+ $X2=0 $Y2=0
cc_350 N_RESET_B_c_282_n N_A_1482_48#_c_1144_n 3.55688e-19 $X=8.18 $Y=2.28 $X2=0
+ $Y2=0
cc_351 N_RESET_B_c_293_n N_A_1482_48#_c_1144_n 0.00823641f $X=8.135 $Y=2 $X2=0
+ $Y2=0
cc_352 N_RESET_B_M1030_g N_A_1482_48#_c_1139_n 0.0401889f $X=8.045 $Y=0.58 $X2=0
+ $Y2=0
cc_353 N_RESET_B_c_286_n N_A_1224_74#_M1032_d 0.00185339f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_354 N_RESET_B_M1030_g N_A_1224_74#_M1031_g 0.0533792f $X=8.045 $Y=0.58 $X2=0
+ $Y2=0
cc_355 N_RESET_B_M1030_g N_A_1224_74#_c_1228_n 0.00701487f $X=8.045 $Y=0.58
+ $X2=0 $Y2=0
cc_356 N_RESET_B_c_282_n N_A_1224_74#_c_1228_n 0.0230744f $X=8.18 $Y=2.28 $X2=0
+ $Y2=0
cc_357 N_RESET_B_c_293_n N_A_1224_74#_c_1228_n 3.64033e-19 $X=8.135 $Y=2 $X2=0
+ $Y2=0
cc_358 N_RESET_B_c_282_n N_A_1224_74#_c_1245_n 0.00895543f $X=8.18 $Y=2.28 $X2=0
+ $Y2=0
cc_359 N_RESET_B_M1030_g N_A_1224_74#_c_1230_n 0.0220605f $X=8.045 $Y=0.58 $X2=0
+ $Y2=0
cc_360 N_RESET_B_c_286_n N_A_1224_74#_c_1257_n 0.0113671f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_361 N_RESET_B_c_286_n N_A_1224_74#_c_1238_n 0.00715094f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_362 N_RESET_B_c_286_n N_A_1224_74#_c_1239_n 0.00106639f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_363 N_RESET_B_M1030_g N_A_1224_74#_c_1240_n 0.00129569f $X=8.045 $Y=0.58
+ $X2=0 $Y2=0
cc_364 N_RESET_B_c_282_n N_A_1224_74#_c_1240_n 0.00121033f $X=8.18 $Y=2.28 $X2=0
+ $Y2=0
cc_365 N_RESET_B_c_286_n N_A_1224_74#_c_1240_n 0.0226223f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_366 N_RESET_B_c_288_n N_A_1224_74#_c_1240_n 0.00270727f $X=7.92 $Y=2.035
+ $X2=0 $Y2=0
cc_367 N_RESET_B_c_293_n N_A_1224_74#_c_1240_n 0.0230781f $X=8.135 $Y=2 $X2=0
+ $Y2=0
cc_368 N_RESET_B_M1030_g N_A_1224_74#_c_1241_n 0.0108822f $X=8.045 $Y=0.58 $X2=0
+ $Y2=0
cc_369 N_RESET_B_c_282_n N_A_1224_74#_c_1241_n 0.00436274f $X=8.18 $Y=2.28 $X2=0
+ $Y2=0
cc_370 N_RESET_B_c_286_n N_A_1224_74#_c_1241_n 0.00339956f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_371 N_RESET_B_c_288_n N_A_1224_74#_c_1241_n 0.00379913f $X=7.92 $Y=2.035
+ $X2=0 $Y2=0
cc_372 N_RESET_B_c_293_n N_A_1224_74#_c_1241_n 0.0255102f $X=8.135 $Y=2 $X2=0
+ $Y2=0
cc_373 N_RESET_B_M1030_g N_A_1224_74#_c_1243_n 0.00118353f $X=8.045 $Y=0.58
+ $X2=0 $Y2=0
cc_374 N_RESET_B_c_284_n N_VPWR_M1017_d 0.00649671f $X=5.375 $Y=2.035 $X2=0
+ $Y2=0
cc_375 N_RESET_B_c_286_n N_VPWR_M1028_s 0.00310864f $X=7.775 $Y=2.035 $X2=0
+ $Y2=0
cc_376 N_RESET_B_c_278_n N_VPWR_c_1444_n 0.00589882f $X=0.955 $Y=2.465 $X2=0
+ $Y2=0
cc_377 N_RESET_B_c_280_n N_VPWR_c_1446_n 0.00321752f $X=4.93 $Y=2.24 $X2=0 $Y2=0
cc_378 N_RESET_B_c_286_n N_VPWR_c_1447_n 0.0237051f $X=7.775 $Y=2.035 $X2=0
+ $Y2=0
cc_379 N_RESET_B_c_287_n N_VPWR_c_1447_n 0.00275995f $X=5.665 $Y=2.035 $X2=0
+ $Y2=0
cc_380 N_RESET_B_c_289_n N_VPWR_c_1447_n 0.00101439f $X=5.395 $Y=1.99 $X2=0
+ $Y2=0
cc_381 N_RESET_B_c_290_n N_VPWR_c_1447_n 0.0239958f $X=5.395 $Y=1.99 $X2=0 $Y2=0
cc_382 N_RESET_B_c_282_n N_VPWR_c_1448_n 0.0062044f $X=8.18 $Y=2.28 $X2=0 $Y2=0
cc_383 N_RESET_B_c_288_n N_VPWR_c_1448_n 0.00183431f $X=7.92 $Y=2.035 $X2=0
+ $Y2=0
cc_384 N_RESET_B_c_293_n N_VPWR_c_1448_n 0.0174647f $X=8.135 $Y=2 $X2=0 $Y2=0
cc_385 N_RESET_B_c_282_n N_VPWR_c_1449_n 0.00454183f $X=8.18 $Y=2.28 $X2=0 $Y2=0
cc_386 N_RESET_B_c_278_n N_VPWR_c_1452_n 0.00444469f $X=0.955 $Y=2.465 $X2=0
+ $Y2=0
cc_387 N_RESET_B_c_278_n N_VPWR_c_1441_n 0.0046079f $X=0.955 $Y=2.465 $X2=0
+ $Y2=0
cc_388 N_RESET_B_c_280_n N_VPWR_c_1441_n 9.39239e-19 $X=4.93 $Y=2.24 $X2=0 $Y2=0
cc_389 N_RESET_B_c_282_n N_VPWR_c_1441_n 0.00489211f $X=8.18 $Y=2.28 $X2=0 $Y2=0
cc_390 N_RESET_B_M1033_g N_A_38_78#_c_1581_n 7.65322e-19 $X=0.94 $Y=0.6 $X2=0
+ $Y2=0
cc_391 N_RESET_B_M1033_g N_A_38_78#_c_1582_n 0.016607f $X=0.94 $Y=0.6 $X2=0
+ $Y2=0
cc_392 N_RESET_B_c_285_n N_A_38_78#_c_1582_n 0.00199354f $X=1.345 $Y=2.035 $X2=0
+ $Y2=0
cc_393 N_RESET_B_c_275_n N_A_38_78#_c_1582_n 0.0731888f $X=1.165 $Y=1.295 $X2=0
+ $Y2=0
cc_394 N_RESET_B_c_277_n N_A_38_78#_c_1588_n 0.00857116f $X=0.955 $Y=2.375 $X2=0
+ $Y2=0
cc_395 N_RESET_B_c_278_n N_A_38_78#_c_1588_n 0.00725597f $X=0.955 $Y=2.465 $X2=0
+ $Y2=0
cc_396 N_RESET_B_c_284_n N_A_38_78#_c_1588_n 0.0370624f $X=5.375 $Y=2.035 $X2=0
+ $Y2=0
cc_397 N_RESET_B_c_285_n N_A_38_78#_c_1588_n 0.00899314f $X=1.345 $Y=2.035 $X2=0
+ $Y2=0
cc_398 N_RESET_B_c_275_n N_A_38_78#_c_1588_n 0.0173863f $X=1.165 $Y=1.295 $X2=0
+ $Y2=0
cc_399 N_RESET_B_c_292_n N_A_38_78#_c_1588_n 0.00281001f $X=1.165 $Y=1.975 $X2=0
+ $Y2=0
cc_400 N_RESET_B_c_284_n N_A_38_78#_c_1589_n 0.0181085f $X=5.375 $Y=2.035 $X2=0
+ $Y2=0
cc_401 N_RESET_B_c_284_n N_A_38_78#_c_1584_n 0.0105056f $X=5.375 $Y=2.035 $X2=0
+ $Y2=0
cc_402 N_RESET_B_M1033_g N_A_38_78#_c_1585_n 8.39005e-19 $X=0.94 $Y=0.6 $X2=0
+ $Y2=0
cc_403 N_RESET_B_c_277_n N_A_38_78#_c_1591_n 0.00220362f $X=0.955 $Y=2.375 $X2=0
+ $Y2=0
cc_404 N_RESET_B_c_278_n N_A_38_78#_c_1591_n 0.0135313f $X=0.955 $Y=2.465 $X2=0
+ $Y2=0
cc_405 N_RESET_B_c_284_n N_A_38_78#_c_1592_n 0.0207866f $X=5.375 $Y=2.035 $X2=0
+ $Y2=0
cc_406 N_RESET_B_c_284_n N_A_38_78#_c_1586_n 0.00574905f $X=5.375 $Y=2.035 $X2=0
+ $Y2=0
cc_407 N_RESET_B_M1033_g N_VGND_c_1738_n 0.00630196f $X=0.94 $Y=0.6 $X2=0 $Y2=0
cc_408 N_RESET_B_c_274_n N_VGND_c_1738_n 0.00181416f $X=1.165 $Y=1.295 $X2=0
+ $Y2=0
cc_409 N_RESET_B_c_275_n N_VGND_c_1738_n 0.0144384f $X=1.165 $Y=1.295 $X2=0
+ $Y2=0
cc_410 N_RESET_B_M1030_g N_VGND_c_1741_n 0.0152783f $X=8.045 $Y=0.58 $X2=0 $Y2=0
cc_411 N_RESET_B_M1033_g N_VGND_c_1744_n 0.00563421f $X=0.94 $Y=0.6 $X2=0 $Y2=0
cc_412 N_RESET_B_c_272_n N_VGND_c_1745_n 0.0033127f $X=4.89 $Y=1.085 $X2=0 $Y2=0
cc_413 N_RESET_B_M1030_g N_VGND_c_1747_n 0.00383152f $X=8.045 $Y=0.58 $X2=0
+ $Y2=0
cc_414 N_RESET_B_M1033_g N_VGND_c_1750_n 0.00539454f $X=0.94 $Y=0.6 $X2=0 $Y2=0
cc_415 N_RESET_B_M1030_g N_VGND_c_1750_n 0.0075725f $X=8.045 $Y=0.58 $X2=0 $Y2=0
cc_416 N_RESET_B_c_272_n N_VGND_c_1750_n 0.00479212f $X=4.89 $Y=1.085 $X2=0
+ $Y2=0
cc_417 CLK N_A_498_360#_c_509_n 6.59991e-19 $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_418 N_CLK_c_459_n N_A_498_360#_c_523_n 0.00121483f $X=1.965 $Y=1.725 $X2=0
+ $Y2=0
cc_419 CLK N_A_498_360#_c_523_n 0.00781881f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_420 N_CLK_c_459_n N_A_319_360#_c_955_n 0.0410783f $X=1.965 $Y=1.725 $X2=0
+ $Y2=0
cc_421 CLK N_A_319_360#_c_955_n 4.81376e-19 $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_422 N_CLK_M1002_g N_A_319_360#_c_942_n 0.0212584f $X=1.97 $Y=0.74 $X2=0 $Y2=0
cc_423 N_CLK_c_459_n N_A_319_360#_c_945_n 0.0245971f $X=1.965 $Y=1.725 $X2=0
+ $Y2=0
cc_424 N_CLK_M1002_g N_A_319_360#_c_945_n 0.0060685f $X=1.97 $Y=0.74 $X2=0 $Y2=0
cc_425 CLK N_A_319_360#_c_945_n 0.0044697f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_426 N_CLK_M1002_g N_A_319_360#_c_950_n 0.0101587f $X=1.97 $Y=0.74 $X2=0 $Y2=0
cc_427 N_CLK_c_459_n N_A_319_360#_c_951_n 0.00476904f $X=1.965 $Y=1.725 $X2=0
+ $Y2=0
cc_428 N_CLK_M1002_g N_A_319_360#_c_951_n 0.00355229f $X=1.97 $Y=0.74 $X2=0
+ $Y2=0
cc_429 CLK N_A_319_360#_c_951_n 0.031171f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_430 N_CLK_c_459_n N_A_319_360#_c_952_n 4.93185e-19 $X=1.965 $Y=1.725 $X2=0
+ $Y2=0
cc_431 N_CLK_M1002_g N_A_319_360#_c_952_n 0.0117933f $X=1.97 $Y=0.74 $X2=0 $Y2=0
cc_432 CLK N_A_319_360#_c_952_n 0.0274826f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_433 N_CLK_M1002_g N_A_319_360#_c_953_n 0.00145065f $X=1.97 $Y=0.74 $X2=0
+ $Y2=0
cc_434 CLK N_A_319_360#_c_953_n 0.0196155f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_435 N_CLK_c_459_n N_A_319_360#_c_954_n 0.00142627f $X=1.965 $Y=1.725 $X2=0
+ $Y2=0
cc_436 N_CLK_M1002_g N_A_319_360#_c_954_n 0.00133296f $X=1.97 $Y=0.74 $X2=0
+ $Y2=0
cc_437 CLK N_A_319_360#_c_954_n 0.00920934f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_438 N_CLK_c_459_n N_A_319_360#_c_971_n 8.2387e-19 $X=1.965 $Y=1.725 $X2=0
+ $Y2=0
cc_439 CLK N_A_319_360#_c_971_n 0.00109875f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_440 N_CLK_c_459_n N_VPWR_c_1444_n 0.00969432f $X=1.965 $Y=1.725 $X2=0 $Y2=0
cc_441 N_CLK_c_459_n N_VPWR_c_1445_n 0.0190995f $X=1.965 $Y=1.725 $X2=0 $Y2=0
cc_442 N_CLK_c_459_n N_VPWR_c_1453_n 0.00492531f $X=1.965 $Y=1.725 $X2=0 $Y2=0
cc_443 N_CLK_c_459_n N_VPWR_c_1441_n 0.00483326f $X=1.965 $Y=1.725 $X2=0 $Y2=0
cc_444 N_CLK_c_459_n N_A_38_78#_c_1588_n 0.0159566f $X=1.965 $Y=1.725 $X2=0
+ $Y2=0
cc_445 CLK N_A_38_78#_c_1588_n 0.00483858f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_446 N_CLK_M1002_g N_VGND_c_1738_n 0.00316318f $X=1.97 $Y=0.74 $X2=0 $Y2=0
cc_447 N_CLK_M1002_g N_VGND_c_1739_n 0.00434272f $X=1.97 $Y=0.74 $X2=0 $Y2=0
cc_448 N_CLK_M1002_g N_VGND_c_1740_n 0.00598308f $X=1.97 $Y=0.74 $X2=0 $Y2=0
cc_449 N_CLK_M1002_g N_VGND_c_1750_n 0.00826311f $X=1.97 $Y=0.74 $X2=0 $Y2=0
cc_450 N_A_498_360#_c_513_n N_A_841_401#_M1004_d 0.0095109f $X=6.085 $Y=0.665
+ $X2=-0.19 $Y2=-0.245
cc_451 N_A_498_360#_c_503_n N_A_841_401#_M1006_g 0.00801556f $X=3.975 $Y=1.575
+ $X2=0 $Y2=0
cc_452 N_A_498_360#_c_504_n N_A_841_401#_M1006_g 0.0414117f $X=4.085 $Y=1.095
+ $X2=0 $Y2=0
cc_453 N_A_498_360#_c_512_n N_A_841_401#_M1006_g 0.00547982f $X=4.435 $Y=0.58
+ $X2=0 $Y2=0
cc_454 N_A_498_360#_c_513_n N_A_841_401#_M1006_g 0.00301737f $X=6.085 $Y=0.665
+ $X2=0 $Y2=0
cc_455 N_A_498_360#_c_546_p N_A_841_401#_M1006_g 0.00422982f $X=4.52 $Y=0.665
+ $X2=0 $Y2=0
cc_456 N_A_498_360#_c_519_n N_A_841_401#_c_710_n 0.00243638f $X=3.455 $Y=2.15
+ $X2=0 $Y2=0
cc_457 N_A_498_360#_c_502_n N_A_841_401#_c_710_n 0.00593179f $X=3.9 $Y=1.65
+ $X2=0 $Y2=0
cc_458 N_A_498_360#_c_503_n N_A_841_401#_c_701_n 8.60057e-19 $X=3.975 $Y=1.575
+ $X2=0 $Y2=0
cc_459 N_A_498_360#_c_504_n N_A_841_401#_c_701_n 4.83625e-19 $X=4.085 $Y=1.095
+ $X2=0 $Y2=0
cc_460 N_A_498_360#_c_503_n N_A_841_401#_c_702_n 0.00593179f $X=3.975 $Y=1.575
+ $X2=0 $Y2=0
cc_461 N_A_498_360#_c_513_n N_A_841_401#_c_703_n 0.0628972f $X=6.085 $Y=0.665
+ $X2=0 $Y2=0
cc_462 N_A_498_360#_c_504_n N_A_841_401#_c_704_n 3.61442e-19 $X=4.085 $Y=1.095
+ $X2=0 $Y2=0
cc_463 N_A_498_360#_c_513_n N_A_841_401#_c_704_n 0.00412245f $X=6.085 $Y=0.665
+ $X2=0 $Y2=0
cc_464 N_A_498_360#_c_546_p N_A_841_401#_c_704_n 0.00987819f $X=4.52 $Y=0.665
+ $X2=0 $Y2=0
cc_465 N_A_498_360#_c_505_n N_A_841_401#_c_705_n 0.00136384f $X=6.045 $Y=1.085
+ $X2=0 $Y2=0
cc_466 N_A_498_360#_c_513_n N_A_841_401#_c_705_n 0.0136179f $X=6.085 $Y=0.665
+ $X2=0 $Y2=0
cc_467 N_A_498_360#_c_558_p N_A_841_401#_c_705_n 0.0108515f $X=6.255 $Y=1.065
+ $X2=0 $Y2=0
cc_468 N_A_498_360#_c_507_n N_A_841_401#_c_706_n 0.00176493f $X=6.12 $Y=1.16
+ $X2=0 $Y2=0
cc_469 N_A_498_360#_c_558_p N_A_841_401#_c_706_n 0.011149f $X=6.255 $Y=1.065
+ $X2=0 $Y2=0
cc_470 N_A_498_360#_c_506_n N_A_841_401#_c_707_n 0.00507154f $X=6.48 $Y=1.16
+ $X2=0 $Y2=0
cc_471 N_A_498_360#_c_507_n N_A_841_401#_c_707_n 0.00303743f $X=6.12 $Y=1.16
+ $X2=0 $Y2=0
cc_472 N_A_498_360#_c_513_n N_A_841_401#_c_707_n 0.00373373f $X=6.085 $Y=0.665
+ $X2=0 $Y2=0
cc_473 N_A_498_360#_c_514_n N_A_841_401#_c_707_n 0.0188995f $X=6.65 $Y=1.065
+ $X2=0 $Y2=0
cc_474 N_A_498_360#_c_558_p N_A_841_401#_c_707_n 0.0136879f $X=6.255 $Y=1.065
+ $X2=0 $Y2=0
cc_475 N_A_498_360#_c_516_n N_A_841_401#_c_707_n 0.0135711f $X=6.735 $Y=1.865
+ $X2=0 $Y2=0
cc_476 N_A_498_360#_c_522_n N_A_841_401#_c_714_n 0.00141721f $X=7.25 $Y=2.28
+ $X2=0 $Y2=0
cc_477 N_A_498_360#_c_516_n N_A_841_401#_c_714_n 0.016501f $X=6.735 $Y=1.865
+ $X2=0 $Y2=0
cc_478 N_A_498_360#_c_535_n N_A_841_401#_c_714_n 0.0140459f $X=6.82 $Y=2.03
+ $X2=0 $Y2=0
cc_479 N_A_498_360#_c_505_n N_A_706_463#_M1004_g 0.0261676f $X=6.045 $Y=1.085
+ $X2=0 $Y2=0
cc_480 N_A_498_360#_c_513_n N_A_706_463#_M1004_g 0.0128398f $X=6.085 $Y=0.665
+ $X2=0 $Y2=0
cc_481 N_A_498_360#_c_572_p N_A_706_463#_M1004_g 6.89487e-19 $X=6.17 $Y=0.9
+ $X2=0 $Y2=0
cc_482 N_A_498_360#_c_558_p N_A_706_463#_M1004_g 2.33891e-19 $X=6.255 $Y=1.065
+ $X2=0 $Y2=0
cc_483 N_A_498_360#_c_507_n N_A_706_463#_c_814_n 0.0123428f $X=6.12 $Y=1.16
+ $X2=0 $Y2=0
cc_484 N_A_498_360#_c_519_n N_A_706_463#_c_815_n 4.02488e-19 $X=3.455 $Y=2.15
+ $X2=0 $Y2=0
cc_485 N_A_498_360#_c_502_n N_A_706_463#_c_815_n 0.00449587f $X=3.9 $Y=1.65
+ $X2=0 $Y2=0
cc_486 N_A_498_360#_c_503_n N_A_706_463#_c_815_n 0.00635368f $X=3.975 $Y=1.575
+ $X2=0 $Y2=0
cc_487 N_A_498_360#_c_504_n N_A_706_463#_c_815_n 0.00267225f $X=4.085 $Y=1.095
+ $X2=0 $Y2=0
cc_488 N_A_498_360#_c_508_n N_A_706_463#_c_815_n 0.00702274f $X=4.085 $Y=1.17
+ $X2=0 $Y2=0
cc_489 N_A_498_360#_c_520_n N_A_706_463#_c_822_n 0.00141905f $X=3.455 $Y=2.24
+ $X2=0 $Y2=0
cc_490 N_A_498_360#_c_502_n N_A_706_463#_c_822_n 0.00106793f $X=3.9 $Y=1.65
+ $X2=0 $Y2=0
cc_491 N_A_498_360#_c_502_n N_A_706_463#_c_816_n 0.00155973f $X=3.9 $Y=1.65
+ $X2=0 $Y2=0
cc_492 N_A_498_360#_c_504_n N_A_706_463#_c_816_n 0.00947091f $X=4.085 $Y=1.095
+ $X2=0 $Y2=0
cc_493 N_A_498_360#_c_508_n N_A_706_463#_c_816_n 0.00554532f $X=4.085 $Y=1.17
+ $X2=0 $Y2=0
cc_494 N_A_498_360#_c_510_n N_A_706_463#_c_816_n 0.0317578f $X=4.35 $Y=0.34
+ $X2=0 $Y2=0
cc_495 N_A_498_360#_c_523_n N_A_319_360#_c_955_n 0.0079624f $X=3.115 $Y=1.74
+ $X2=0 $Y2=0
cc_496 N_A_498_360#_c_509_n N_A_319_360#_c_942_n 0.0059419f $X=3.03 $Y=1.575
+ $X2=0 $Y2=0
cc_497 N_A_498_360#_c_510_n N_A_319_360#_c_942_n 2.90433e-19 $X=4.35 $Y=0.34
+ $X2=0 $Y2=0
cc_498 N_A_498_360#_c_517_n N_A_319_360#_c_942_n 0.00956439f $X=2.852 $Y=0.34
+ $X2=0 $Y2=0
cc_499 N_A_498_360#_c_519_n N_A_319_360#_c_943_n 0.0111591f $X=3.455 $Y=2.15
+ $X2=0 $Y2=0
cc_500 N_A_498_360#_c_520_n N_A_319_360#_c_943_n 0.0128837f $X=3.455 $Y=2.24
+ $X2=0 $Y2=0
cc_501 N_A_498_360#_c_509_n N_A_319_360#_c_943_n 8.99067e-19 $X=3.03 $Y=1.575
+ $X2=0 $Y2=0
cc_502 N_A_498_360#_c_523_n N_A_319_360#_c_943_n 0.0229657f $X=3.115 $Y=1.74
+ $X2=0 $Y2=0
cc_503 N_A_498_360#_c_518_n N_A_319_360#_c_943_n 0.021379f $X=3.385 $Y=1.65
+ $X2=0 $Y2=0
cc_504 N_A_498_360#_c_503_n N_A_319_360#_c_944_n 0.00605671f $X=3.975 $Y=1.575
+ $X2=0 $Y2=0
cc_505 N_A_498_360#_c_509_n N_A_319_360#_c_944_n 0.00834646f $X=3.03 $Y=1.575
+ $X2=0 $Y2=0
cc_506 N_A_498_360#_c_511_n N_A_319_360#_c_944_n 0.00427309f $X=3.385 $Y=1.74
+ $X2=0 $Y2=0
cc_507 N_A_498_360#_c_518_n N_A_319_360#_c_944_n 0.0237371f $X=3.385 $Y=1.65
+ $X2=0 $Y2=0
cc_508 N_A_498_360#_c_509_n N_A_319_360#_c_945_n 0.0109326f $X=3.03 $Y=1.575
+ $X2=0 $Y2=0
cc_509 N_A_498_360#_c_523_n N_A_319_360#_c_945_n 0.00633977f $X=3.115 $Y=1.74
+ $X2=0 $Y2=0
cc_510 N_A_498_360#_c_517_n N_A_319_360#_c_945_n 0.0064559f $X=2.852 $Y=0.34
+ $X2=0 $Y2=0
cc_511 N_A_498_360#_c_520_n N_A_319_360#_c_958_n 0.0103487f $X=3.455 $Y=2.24
+ $X2=0 $Y2=0
cc_512 N_A_498_360#_c_504_n N_A_319_360#_M1020_g 0.0132831f $X=4.085 $Y=1.095
+ $X2=0 $Y2=0
cc_513 N_A_498_360#_c_508_n N_A_319_360#_M1020_g 0.00605671f $X=4.085 $Y=1.17
+ $X2=0 $Y2=0
cc_514 N_A_498_360#_c_510_n N_A_319_360#_M1020_g 0.00680216f $X=4.35 $Y=0.34
+ $X2=0 $Y2=0
cc_515 N_A_498_360#_c_517_n N_A_319_360#_M1020_g 0.005681f $X=2.852 $Y=0.34
+ $X2=0 $Y2=0
cc_516 N_A_498_360#_c_520_n N_A_319_360#_c_960_n 0.00278823f $X=3.455 $Y=2.24
+ $X2=0 $Y2=0
cc_517 N_A_498_360#_c_520_n N_A_319_360#_c_962_n 0.0114271f $X=3.455 $Y=2.24
+ $X2=0 $Y2=0
cc_518 N_A_498_360#_c_502_n N_A_319_360#_c_962_n 0.00429214f $X=3.9 $Y=1.65
+ $X2=0 $Y2=0
cc_519 N_A_498_360#_c_522_n N_A_319_360#_c_964_n 0.002647f $X=7.25 $Y=2.28 $X2=0
+ $Y2=0
cc_520 N_A_498_360#_c_522_n N_A_319_360#_M1032_g 0.0194051f $X=7.25 $Y=2.28
+ $X2=0 $Y2=0
cc_521 N_A_498_360#_c_516_n N_A_319_360#_M1032_g 0.0042093f $X=6.735 $Y=1.865
+ $X2=0 $Y2=0
cc_522 N_A_498_360#_c_535_n N_A_319_360#_M1032_g 0.00216411f $X=6.82 $Y=2.03
+ $X2=0 $Y2=0
cc_523 N_A_498_360#_c_522_n N_A_319_360#_c_947_n 0.00720172f $X=7.25 $Y=2.28
+ $X2=0 $Y2=0
cc_524 N_A_498_360#_c_515_n N_A_319_360#_c_947_n 0.0103797f $X=6.645 $Y=1.065
+ $X2=0 $Y2=0
cc_525 N_A_498_360#_c_516_n N_A_319_360#_c_947_n 0.0123591f $X=6.735 $Y=1.865
+ $X2=0 $Y2=0
cc_526 N_A_498_360#_c_526_n N_A_319_360#_c_947_n 0.00746766f $X=7.205 $Y=2.03
+ $X2=0 $Y2=0
cc_527 N_A_498_360#_c_506_n N_A_319_360#_c_948_n 0.0103797f $X=6.48 $Y=1.16
+ $X2=0 $Y2=0
cc_528 N_A_498_360#_c_514_n N_A_319_360#_c_948_n 0.00126209f $X=6.65 $Y=1.065
+ $X2=0 $Y2=0
cc_529 N_A_498_360#_c_516_n N_A_319_360#_c_948_n 8.31237e-19 $X=6.735 $Y=1.865
+ $X2=0 $Y2=0
cc_530 N_A_498_360#_c_514_n N_A_319_360#_M1003_g 0.00116888f $X=6.65 $Y=1.065
+ $X2=0 $Y2=0
cc_531 N_A_498_360#_c_515_n N_A_319_360#_M1003_g 0.0216896f $X=6.645 $Y=1.065
+ $X2=0 $Y2=0
cc_532 N_A_498_360#_c_516_n N_A_319_360#_M1003_g 0.00159607f $X=6.735 $Y=1.865
+ $X2=0 $Y2=0
cc_533 N_A_498_360#_M1013_d N_A_319_360#_c_952_n 0.00267638f $X=2.615 $Y=0.37
+ $X2=0 $Y2=0
cc_534 N_A_498_360#_c_509_n N_A_319_360#_c_952_n 0.0141097f $X=3.03 $Y=1.575
+ $X2=0 $Y2=0
cc_535 N_A_498_360#_c_517_n N_A_319_360#_c_952_n 0.0110032f $X=2.852 $Y=0.34
+ $X2=0 $Y2=0
cc_536 N_A_498_360#_c_509_n N_A_319_360#_c_953_n 0.0295916f $X=3.03 $Y=1.575
+ $X2=0 $Y2=0
cc_537 N_A_498_360#_c_523_n N_A_319_360#_c_953_n 0.0223623f $X=3.115 $Y=1.74
+ $X2=0 $Y2=0
cc_538 N_A_498_360#_c_523_n N_A_319_360#_c_971_n 0.00673278f $X=3.115 $Y=1.74
+ $X2=0 $Y2=0
cc_539 N_A_498_360#_c_522_n N_A_1482_48#_c_1133_n 0.0212122f $X=7.25 $Y=2.28
+ $X2=0 $Y2=0
cc_540 N_A_498_360#_c_526_n N_A_1482_48#_c_1133_n 4.05192e-19 $X=7.205 $Y=2.03
+ $X2=0 $Y2=0
cc_541 N_A_498_360#_c_522_n N_A_1482_48#_c_1141_n 0.0335632f $X=7.25 $Y=2.28
+ $X2=0 $Y2=0
cc_542 N_A_498_360#_c_513_n N_A_1224_74#_M1007_d 0.00392413f $X=6.085 $Y=0.665
+ $X2=-0.19 $Y2=-0.245
cc_543 N_A_498_360#_c_572_p N_A_1224_74#_M1007_d 0.00564702f $X=6.17 $Y=0.9
+ $X2=-0.19 $Y2=-0.245
cc_544 N_A_498_360#_c_514_n N_A_1224_74#_M1007_d 0.00471261f $X=6.65 $Y=1.065
+ $X2=-0.19 $Y2=-0.245
cc_545 N_A_498_360#_c_516_n N_A_1224_74#_M1032_d 0.00321319f $X=6.735 $Y=1.865
+ $X2=0 $Y2=0
cc_546 N_A_498_360#_c_535_n N_A_1224_74#_M1032_d 0.00528653f $X=6.82 $Y=2.03
+ $X2=0 $Y2=0
cc_547 N_A_498_360#_c_526_n N_A_1224_74#_M1032_d 0.00213077f $X=7.205 $Y=2.03
+ $X2=0 $Y2=0
cc_548 N_A_498_360#_c_505_n N_A_1224_74#_c_1277_n 0.00722906f $X=6.045 $Y=1.085
+ $X2=0 $Y2=0
cc_549 N_A_498_360#_c_513_n N_A_1224_74#_c_1277_n 0.013434f $X=6.085 $Y=0.665
+ $X2=0 $Y2=0
cc_550 N_A_498_360#_c_514_n N_A_1224_74#_c_1277_n 0.0317086f $X=6.65 $Y=1.065
+ $X2=0 $Y2=0
cc_551 N_A_498_360#_c_515_n N_A_1224_74#_c_1277_n 0.00506999f $X=6.645 $Y=1.065
+ $X2=0 $Y2=0
cc_552 N_A_498_360#_c_522_n N_A_1224_74#_c_1257_n 0.0215946f $X=7.25 $Y=2.28
+ $X2=0 $Y2=0
cc_553 N_A_498_360#_c_535_n N_A_1224_74#_c_1257_n 0.00944134f $X=6.82 $Y=2.03
+ $X2=0 $Y2=0
cc_554 N_A_498_360#_c_526_n N_A_1224_74#_c_1257_n 0.0346045f $X=7.205 $Y=2.03
+ $X2=0 $Y2=0
cc_555 N_A_498_360#_c_514_n N_A_1224_74#_c_1237_n 0.0278616f $X=6.65 $Y=1.065
+ $X2=0 $Y2=0
cc_556 N_A_498_360#_c_515_n N_A_1224_74#_c_1237_n 9.55385e-19 $X=6.645 $Y=1.065
+ $X2=0 $Y2=0
cc_557 N_A_498_360#_c_516_n N_A_1224_74#_c_1237_n 0.0146057f $X=6.735 $Y=1.865
+ $X2=0 $Y2=0
cc_558 N_A_498_360#_c_522_n N_A_1224_74#_c_1238_n 0.00534955f $X=7.25 $Y=2.28
+ $X2=0 $Y2=0
cc_559 N_A_498_360#_c_526_n N_A_1224_74#_c_1238_n 0.00761315f $X=7.205 $Y=2.03
+ $X2=0 $Y2=0
cc_560 N_A_498_360#_c_522_n N_A_1224_74#_c_1239_n 4.21127e-19 $X=7.25 $Y=2.28
+ $X2=0 $Y2=0
cc_561 N_A_498_360#_c_516_n N_A_1224_74#_c_1239_n 0.0133634f $X=6.735 $Y=1.865
+ $X2=0 $Y2=0
cc_562 N_A_498_360#_c_526_n N_A_1224_74#_c_1239_n 0.00832552f $X=7.205 $Y=2.03
+ $X2=0 $Y2=0
cc_563 N_A_498_360#_c_522_n N_A_1224_74#_c_1240_n 0.005245f $X=7.25 $Y=2.28
+ $X2=0 $Y2=0
cc_564 N_A_498_360#_c_516_n N_A_1224_74#_c_1240_n 0.00741853f $X=6.735 $Y=1.865
+ $X2=0 $Y2=0
cc_565 N_A_498_360#_c_526_n N_A_1224_74#_c_1240_n 0.0242903f $X=7.205 $Y=2.03
+ $X2=0 $Y2=0
cc_566 N_A_498_360#_c_522_n N_VPWR_c_1456_n 0.00349642f $X=7.25 $Y=2.28 $X2=0
+ $Y2=0
cc_567 N_A_498_360#_c_520_n N_VPWR_c_1441_n 9.39239e-19 $X=3.455 $Y=2.24 $X2=0
+ $Y2=0
cc_568 N_A_498_360#_c_522_n N_VPWR_c_1441_n 0.00489211f $X=7.25 $Y=2.28 $X2=0
+ $Y2=0
cc_569 N_A_498_360#_M1023_d N_A_38_78#_c_1588_n 0.00723917f $X=2.49 $Y=1.8 $X2=0
+ $Y2=0
cc_570 N_A_498_360#_c_523_n N_A_38_78#_c_1588_n 0.0245465f $X=3.115 $Y=1.74
+ $X2=0 $Y2=0
cc_571 N_A_498_360#_c_504_n N_A_38_78#_c_1583_n 3.16057e-19 $X=4.085 $Y=1.095
+ $X2=0 $Y2=0
cc_572 N_A_498_360#_c_508_n N_A_38_78#_c_1583_n 3.23037e-19 $X=4.085 $Y=1.17
+ $X2=0 $Y2=0
cc_573 N_A_498_360#_c_510_n N_A_38_78#_c_1583_n 0.0167583f $X=4.35 $Y=0.34 $X2=0
+ $Y2=0
cc_574 N_A_498_360#_c_517_n N_A_38_78#_c_1583_n 0.0476134f $X=2.852 $Y=0.34
+ $X2=0 $Y2=0
cc_575 N_A_498_360#_c_519_n N_A_38_78#_c_1589_n 0.00418749f $X=3.455 $Y=2.15
+ $X2=0 $Y2=0
cc_576 N_A_498_360#_c_520_n N_A_38_78#_c_1589_n 0.00876534f $X=3.455 $Y=2.24
+ $X2=0 $Y2=0
cc_577 N_A_498_360#_c_502_n N_A_38_78#_c_1589_n 0.00284282f $X=3.9 $Y=1.65 $X2=0
+ $Y2=0
cc_578 N_A_498_360#_c_511_n N_A_38_78#_c_1589_n 0.0064771f $X=3.385 $Y=1.74
+ $X2=0 $Y2=0
cc_579 N_A_498_360#_c_519_n N_A_38_78#_c_1584_n 0.00482637f $X=3.455 $Y=2.15
+ $X2=0 $Y2=0
cc_580 N_A_498_360#_c_502_n N_A_38_78#_c_1584_n 0.0131596f $X=3.9 $Y=1.65 $X2=0
+ $Y2=0
cc_581 N_A_498_360#_c_503_n N_A_38_78#_c_1584_n 0.00444981f $X=3.975 $Y=1.575
+ $X2=0 $Y2=0
cc_582 N_A_498_360#_c_509_n N_A_38_78#_c_1584_n 0.00677786f $X=3.03 $Y=1.575
+ $X2=0 $Y2=0
cc_583 N_A_498_360#_c_511_n N_A_38_78#_c_1584_n 0.0254503f $X=3.385 $Y=1.74
+ $X2=0 $Y2=0
cc_584 N_A_498_360#_c_518_n N_A_38_78#_c_1584_n 0.00429414f $X=3.385 $Y=1.65
+ $X2=0 $Y2=0
cc_585 N_A_498_360#_c_519_n N_A_38_78#_c_1592_n 0.00144717f $X=3.455 $Y=2.15
+ $X2=0 $Y2=0
cc_586 N_A_498_360#_c_520_n N_A_38_78#_c_1592_n 0.0102027f $X=3.455 $Y=2.24
+ $X2=0 $Y2=0
cc_587 N_A_498_360#_c_523_n N_A_38_78#_c_1592_n 0.00722647f $X=3.115 $Y=1.74
+ $X2=0 $Y2=0
cc_588 N_A_498_360#_c_511_n N_A_38_78#_c_1592_n 0.0187455f $X=3.385 $Y=1.74
+ $X2=0 $Y2=0
cc_589 N_A_498_360#_c_518_n N_A_38_78#_c_1592_n 0.00323248f $X=3.385 $Y=1.65
+ $X2=0 $Y2=0
cc_590 N_A_498_360#_c_502_n N_A_38_78#_c_1586_n 7.4782e-19 $X=3.9 $Y=1.65 $X2=0
+ $Y2=0
cc_591 N_A_498_360#_c_508_n N_A_38_78#_c_1586_n 0.00175844f $X=4.085 $Y=1.17
+ $X2=0 $Y2=0
cc_592 N_A_498_360#_c_509_n N_A_38_78#_c_1586_n 0.0128596f $X=3.03 $Y=1.575
+ $X2=0 $Y2=0
cc_593 N_A_498_360#_c_511_n N_A_38_78#_c_1586_n 0.0134538f $X=3.385 $Y=1.74
+ $X2=0 $Y2=0
cc_594 N_A_498_360#_c_518_n N_A_38_78#_c_1586_n 0.00482607f $X=3.385 $Y=1.65
+ $X2=0 $Y2=0
cc_595 N_A_498_360#_c_513_n N_VGND_M1022_d 0.00722747f $X=6.085 $Y=0.665 $X2=0
+ $Y2=0
cc_596 N_A_498_360#_c_517_n N_VGND_c_1740_n 0.0266974f $X=2.852 $Y=0.34 $X2=0
+ $Y2=0
cc_597 N_A_498_360#_c_510_n N_VGND_c_1745_n 0.0914273f $X=4.35 $Y=0.34 $X2=0
+ $Y2=0
cc_598 N_A_498_360#_c_513_n N_VGND_c_1745_n 0.00941901f $X=6.085 $Y=0.665 $X2=0
+ $Y2=0
cc_599 N_A_498_360#_c_517_n N_VGND_c_1745_n 0.0369908f $X=2.852 $Y=0.34 $X2=0
+ $Y2=0
cc_600 N_A_498_360#_c_505_n N_VGND_c_1746_n 0.00320103f $X=6.045 $Y=1.085 $X2=0
+ $Y2=0
cc_601 N_A_498_360#_c_513_n N_VGND_c_1746_n 0.0163564f $X=6.085 $Y=0.665 $X2=0
+ $Y2=0
cc_602 N_A_498_360#_c_505_n N_VGND_c_1750_n 0.00407044f $X=6.045 $Y=1.085 $X2=0
+ $Y2=0
cc_603 N_A_498_360#_c_510_n N_VGND_c_1750_n 0.0529847f $X=4.35 $Y=0.34 $X2=0
+ $Y2=0
cc_604 N_A_498_360#_c_513_n N_VGND_c_1750_n 0.0422032f $X=6.085 $Y=0.665 $X2=0
+ $Y2=0
cc_605 N_A_498_360#_c_517_n N_VGND_c_1750_n 0.0201445f $X=2.852 $Y=0.34 $X2=0
+ $Y2=0
cc_606 N_A_498_360#_c_510_n N_VGND_c_1753_n 0.00672073f $X=4.35 $Y=0.34 $X2=0
+ $Y2=0
cc_607 N_A_498_360#_c_513_n N_VGND_c_1753_n 0.0245264f $X=6.085 $Y=0.665 $X2=0
+ $Y2=0
cc_608 N_A_498_360#_c_513_n A_910_118# 0.00134207f $X=6.085 $Y=0.665 $X2=-0.19
+ $Y2=-0.245
cc_609 N_A_841_401#_c_703_n N_A_706_463#_M1004_g 0.0117829f $X=5.745 $Y=1.005
+ $X2=0 $Y2=0
cc_610 N_A_841_401#_c_706_n N_A_706_463#_M1004_g 0.0046522f $X=5.83 $Y=1.4 $X2=0
+ $Y2=0
cc_611 N_A_841_401#_c_703_n N_A_706_463#_c_814_n 0.00506798f $X=5.745 $Y=1.005
+ $X2=0 $Y2=0
cc_612 N_A_841_401#_c_707_n N_A_706_463#_c_814_n 0.00925955f $X=6.23 $Y=1.485
+ $X2=0 $Y2=0
cc_613 N_A_841_401#_c_708_n N_A_706_463#_c_814_n 0.00867517f $X=5.915 $Y=1.485
+ $X2=0 $Y2=0
cc_614 N_A_841_401#_c_714_n N_A_706_463#_c_814_n 0.00185802f $X=6.315 $Y=1.88
+ $X2=0 $Y2=0
cc_615 N_A_841_401#_c_714_n N_A_706_463#_c_820_n 0.00551932f $X=6.315 $Y=1.88
+ $X2=0 $Y2=0
cc_616 N_A_841_401#_c_709_n N_A_706_463#_c_815_n 0.00213772f $X=4.295 $Y=2.24
+ $X2=0 $Y2=0
cc_617 N_A_841_401#_M1006_g N_A_706_463#_c_815_n 0.00129073f $X=4.475 $Y=0.8
+ $X2=0 $Y2=0
cc_618 N_A_841_401#_c_710_n N_A_706_463#_c_815_n 0.0040903f $X=4.465 $Y=2.005
+ $X2=0 $Y2=0
cc_619 N_A_841_401#_c_701_n N_A_706_463#_c_815_n 0.0796667f $X=4.465 $Y=1.65
+ $X2=0 $Y2=0
cc_620 N_A_841_401#_c_702_n N_A_706_463#_c_815_n 0.00795351f $X=4.465 $Y=1.65
+ $X2=0 $Y2=0
cc_621 N_A_841_401#_c_704_n N_A_706_463#_c_815_n 0.0050659f $X=4.63 $Y=1.005
+ $X2=0 $Y2=0
cc_622 N_A_841_401#_c_709_n N_A_706_463#_c_833_n 0.0125311f $X=4.295 $Y=2.24
+ $X2=0 $Y2=0
cc_623 N_A_841_401#_c_710_n N_A_706_463#_c_833_n 0.00144235f $X=4.465 $Y=2.005
+ $X2=0 $Y2=0
cc_624 N_A_841_401#_c_701_n N_A_706_463#_c_833_n 0.0126181f $X=4.465 $Y=1.65
+ $X2=0 $Y2=0
cc_625 N_A_841_401#_c_709_n N_A_706_463#_c_822_n 8.31361e-19 $X=4.295 $Y=2.24
+ $X2=0 $Y2=0
cc_626 N_A_841_401#_c_709_n N_A_706_463#_c_823_n 5.53787e-19 $X=4.295 $Y=2.24
+ $X2=0 $Y2=0
cc_627 N_A_841_401#_c_710_n N_A_706_463#_c_823_n 4.44352e-19 $X=4.465 $Y=2.005
+ $X2=0 $Y2=0
cc_628 N_A_841_401#_c_701_n N_A_706_463#_c_823_n 0.0259264f $X=4.465 $Y=1.65
+ $X2=0 $Y2=0
cc_629 N_A_841_401#_c_702_n N_A_706_463#_c_823_n 0.00173976f $X=4.465 $Y=1.65
+ $X2=0 $Y2=0
cc_630 N_A_841_401#_c_704_n N_A_706_463#_c_816_n 0.00164172f $X=4.63 $Y=1.005
+ $X2=0 $Y2=0
cc_631 N_A_841_401#_c_701_n N_A_706_463#_c_817_n 0.0144822f $X=4.465 $Y=1.65
+ $X2=0 $Y2=0
cc_632 N_A_841_401#_c_702_n N_A_706_463#_c_817_n 4.19328e-19 $X=4.465 $Y=1.65
+ $X2=0 $Y2=0
cc_633 N_A_841_401#_c_703_n N_A_706_463#_c_817_n 0.0373672f $X=5.745 $Y=1.005
+ $X2=0 $Y2=0
cc_634 N_A_841_401#_c_706_n N_A_706_463#_c_817_n 0.00811118f $X=5.83 $Y=1.4
+ $X2=0 $Y2=0
cc_635 N_A_841_401#_c_708_n N_A_706_463#_c_817_n 0.0135374f $X=5.915 $Y=1.485
+ $X2=0 $Y2=0
cc_636 N_A_841_401#_c_714_n N_A_706_463#_c_817_n 0.0012591f $X=6.315 $Y=1.88
+ $X2=0 $Y2=0
cc_637 N_A_841_401#_c_703_n N_A_706_463#_c_818_n 0.00123201f $X=5.745 $Y=1.005
+ $X2=0 $Y2=0
cc_638 N_A_841_401#_c_706_n N_A_706_463#_c_818_n 7.93674e-19 $X=5.83 $Y=1.4
+ $X2=0 $Y2=0
cc_639 N_A_841_401#_c_708_n N_A_706_463#_c_818_n 5.0886e-19 $X=5.915 $Y=1.485
+ $X2=0 $Y2=0
cc_640 N_A_841_401#_c_709_n N_A_706_463#_c_825_n 7.43442e-19 $X=4.295 $Y=2.24
+ $X2=0 $Y2=0
cc_641 N_A_841_401#_c_709_n N_A_319_360#_c_960_n 0.00323347f $X=4.295 $Y=2.24
+ $X2=0 $Y2=0
cc_642 N_A_841_401#_c_709_n N_A_319_360#_c_962_n 0.0288994f $X=4.295 $Y=2.24
+ $X2=0 $Y2=0
cc_643 N_A_841_401#_c_710_n N_A_319_360#_c_962_n 0.0026362f $X=4.465 $Y=2.005
+ $X2=0 $Y2=0
cc_644 N_A_841_401#_c_709_n N_A_319_360#_c_963_n 0.00993882f $X=4.295 $Y=2.24
+ $X2=0 $Y2=0
cc_645 N_A_841_401#_c_714_n N_A_319_360#_c_963_n 0.00262042f $X=6.315 $Y=1.88
+ $X2=0 $Y2=0
cc_646 N_A_841_401#_c_714_n N_A_319_360#_c_964_n 5.08057e-19 $X=6.315 $Y=1.88
+ $X2=0 $Y2=0
cc_647 N_A_841_401#_c_714_n N_A_319_360#_M1032_g 0.0143858f $X=6.315 $Y=1.88
+ $X2=0 $Y2=0
cc_648 N_A_841_401#_c_707_n N_A_319_360#_c_948_n 0.00287849f $X=6.23 $Y=1.485
+ $X2=0 $Y2=0
cc_649 N_A_841_401#_c_714_n N_A_319_360#_c_948_n 0.00245265f $X=6.315 $Y=1.88
+ $X2=0 $Y2=0
cc_650 N_A_841_401#_c_714_n N_A_1224_74#_c_1257_n 0.0217845f $X=6.315 $Y=1.88
+ $X2=0 $Y2=0
cc_651 N_A_841_401#_c_709_n N_VPWR_c_1446_n 0.00321752f $X=4.295 $Y=2.24 $X2=0
+ $Y2=0
cc_652 N_A_841_401#_c_707_n N_VPWR_c_1447_n 0.00590731f $X=6.23 $Y=1.485 $X2=0
+ $Y2=0
cc_653 N_A_841_401#_c_708_n N_VPWR_c_1447_n 0.0111121f $X=5.915 $Y=1.485 $X2=0
+ $Y2=0
cc_654 N_A_841_401#_c_714_n N_VPWR_c_1447_n 0.0651453f $X=6.315 $Y=1.88 $X2=0
+ $Y2=0
cc_655 N_A_841_401#_c_714_n N_VPWR_c_1456_n 0.00567879f $X=6.315 $Y=1.88 $X2=0
+ $Y2=0
cc_656 N_A_841_401#_c_709_n N_VPWR_c_1441_n 9.39239e-19 $X=4.295 $Y=2.24 $X2=0
+ $Y2=0
cc_657 N_A_841_401#_c_714_n N_VPWR_c_1441_n 0.00684413f $X=6.315 $Y=1.88 $X2=0
+ $Y2=0
cc_658 N_A_841_401#_c_703_n N_VGND_M1022_d 0.00362168f $X=5.745 $Y=1.005 $X2=0
+ $Y2=0
cc_659 N_A_841_401#_M1006_g N_VGND_c_1745_n 0.00113933f $X=4.475 $Y=0.8 $X2=0
+ $Y2=0
cc_660 N_A_841_401#_M1006_g N_VGND_c_1750_n 9.75345e-19 $X=4.475 $Y=0.8 $X2=0
+ $Y2=0
cc_661 N_A_841_401#_c_703_n A_910_118# 0.00108692f $X=5.745 $Y=1.005 $X2=-0.19
+ $Y2=-0.245
cc_662 N_A_841_401#_c_704_n A_910_118# 2.5515e-19 $X=4.63 $Y=1.005 $X2=-0.19
+ $Y2=-0.245
cc_663 N_A_706_463#_c_822_n N_A_319_360#_c_958_n 0.0025201f $X=4.18 $Y=2.5 $X2=0
+ $Y2=0
cc_664 N_A_706_463#_c_815_n N_A_319_360#_M1020_g 5.66449e-19 $X=4.095 $Y=2.415
+ $X2=0 $Y2=0
cc_665 N_A_706_463#_c_816_n N_A_319_360#_M1020_g 0.00232642f $X=4.095 $Y=0.812
+ $X2=0 $Y2=0
cc_666 N_A_706_463#_c_822_n N_A_319_360#_c_960_n 4.85207e-19 $X=4.18 $Y=2.5
+ $X2=0 $Y2=0
cc_667 N_A_706_463#_c_815_n N_A_319_360#_c_962_n 0.00165201f $X=4.095 $Y=2.415
+ $X2=0 $Y2=0
cc_668 N_A_706_463#_c_822_n N_A_319_360#_c_962_n 0.012138f $X=4.18 $Y=2.5 $X2=0
+ $Y2=0
cc_669 N_A_706_463#_c_820_n N_A_319_360#_c_963_n 0.0103562f $X=6.09 $Y=1.66
+ $X2=0 $Y2=0
cc_670 N_A_706_463#_c_833_n N_A_319_360#_c_963_n 0.00347672f $X=4.89 $Y=2.5
+ $X2=0 $Y2=0
cc_671 N_A_706_463#_c_822_n N_A_319_360#_c_963_n 0.00158973f $X=4.18 $Y=2.5
+ $X2=0 $Y2=0
cc_672 N_A_706_463#_c_825_n N_A_319_360#_c_963_n 0.00580249f $X=4.975 $Y=2.515
+ $X2=0 $Y2=0
cc_673 N_A_706_463#_c_820_n N_A_319_360#_c_964_n 0.00249951f $X=6.09 $Y=1.66
+ $X2=0 $Y2=0
cc_674 N_A_706_463#_c_820_n N_A_319_360#_M1032_g 0.00575058f $X=6.09 $Y=1.66
+ $X2=0 $Y2=0
cc_675 N_A_706_463#_c_814_n N_A_319_360#_c_948_n 0.00860655f $X=6 $Y=1.54 $X2=0
+ $Y2=0
cc_676 N_A_706_463#_c_833_n N_VPWR_M1005_d 0.00921529f $X=4.89 $Y=2.5 $X2=0
+ $Y2=0
cc_677 N_A_706_463#_c_833_n N_VPWR_c_1446_n 0.0270329f $X=4.89 $Y=2.5 $X2=0
+ $Y2=0
cc_678 N_A_706_463#_c_814_n N_VPWR_c_1447_n 0.00446017f $X=6 $Y=1.54 $X2=0 $Y2=0
cc_679 N_A_706_463#_c_820_n N_VPWR_c_1447_n 0.0144868f $X=6.09 $Y=1.66 $X2=0
+ $Y2=0
cc_680 N_A_706_463#_c_825_n N_VPWR_c_1447_n 0.0135993f $X=4.975 $Y=2.515 $X2=0
+ $Y2=0
cc_681 N_A_706_463#_c_833_n N_VPWR_c_1454_n 0.00280825f $X=4.89 $Y=2.5 $X2=0
+ $Y2=0
cc_682 N_A_706_463#_c_822_n N_VPWR_c_1454_n 0.00966244f $X=4.18 $Y=2.5 $X2=0
+ $Y2=0
cc_683 N_A_706_463#_c_833_n N_VPWR_c_1455_n 0.00103577f $X=4.89 $Y=2.5 $X2=0
+ $Y2=0
cc_684 N_A_706_463#_c_825_n N_VPWR_c_1455_n 0.00688776f $X=4.975 $Y=2.515 $X2=0
+ $Y2=0
cc_685 N_A_706_463#_c_820_n N_VPWR_c_1441_n 8.51577e-19 $X=6.09 $Y=1.66 $X2=0
+ $Y2=0
cc_686 N_A_706_463#_c_833_n N_VPWR_c_1441_n 0.00928815f $X=4.89 $Y=2.5 $X2=0
+ $Y2=0
cc_687 N_A_706_463#_c_822_n N_VPWR_c_1441_n 0.0142735f $X=4.18 $Y=2.5 $X2=0
+ $Y2=0
cc_688 N_A_706_463#_c_825_n N_VPWR_c_1441_n 0.010728f $X=4.975 $Y=2.515 $X2=0
+ $Y2=0
cc_689 N_A_706_463#_c_815_n N_A_38_78#_c_1583_n 0.00511985f $X=4.095 $Y=2.415
+ $X2=0 $Y2=0
cc_690 N_A_706_463#_c_816_n N_A_38_78#_c_1583_n 0.0164395f $X=4.095 $Y=0.812
+ $X2=0 $Y2=0
cc_691 N_A_706_463#_c_815_n N_A_38_78#_c_1589_n 0.0133272f $X=4.095 $Y=2.415
+ $X2=0 $Y2=0
cc_692 N_A_706_463#_c_822_n N_A_38_78#_c_1589_n 0.0172937f $X=4.18 $Y=2.5 $X2=0
+ $Y2=0
cc_693 N_A_706_463#_c_815_n N_A_38_78#_c_1584_n 0.0505899f $X=4.095 $Y=2.415
+ $X2=0 $Y2=0
cc_694 N_A_706_463#_c_815_n N_A_38_78#_c_1592_n 0.00325632f $X=4.095 $Y=2.415
+ $X2=0 $Y2=0
cc_695 N_A_706_463#_c_822_n N_A_38_78#_c_1592_n 0.0238608f $X=4.18 $Y=2.5 $X2=0
+ $Y2=0
cc_696 N_A_706_463#_c_815_n N_A_38_78#_c_1586_n 0.0132832f $X=4.095 $Y=2.415
+ $X2=0 $Y2=0
cc_697 N_A_706_463#_c_816_n N_A_38_78#_c_1586_n 0.0109432f $X=4.095 $Y=0.812
+ $X2=0 $Y2=0
cc_698 N_A_706_463#_c_822_n A_796_463# 0.0022949f $X=4.18 $Y=2.5 $X2=-0.19
+ $Y2=-0.245
cc_699 N_A_706_463#_M1004_g N_VGND_c_1746_n 0.00320129f $X=5.455 $Y=0.69 $X2=0
+ $Y2=0
cc_700 N_A_706_463#_M1004_g N_VGND_c_1750_n 0.00406112f $X=5.455 $Y=0.69 $X2=0
+ $Y2=0
cc_701 N_A_706_463#_M1004_g N_VGND_c_1753_n 0.00617301f $X=5.455 $Y=0.69 $X2=0
+ $Y2=0
cc_702 N_A_319_360#_M1003_g N_A_1482_48#_c_1132_n 0.0495982f $X=7.095 $Y=0.58
+ $X2=0 $Y2=0
cc_703 N_A_319_360#_M1003_g N_A_1482_48#_c_1133_n 0.0112982f $X=7.095 $Y=0.58
+ $X2=0 $Y2=0
cc_704 N_A_319_360#_M1003_g N_A_1482_48#_c_1137_n 0.00102678f $X=7.095 $Y=0.58
+ $X2=0 $Y2=0
cc_705 N_A_319_360#_M1003_g N_A_1224_74#_c_1277_n 0.0169263f $X=7.095 $Y=0.58
+ $X2=0 $Y2=0
cc_706 N_A_319_360#_M1032_g N_A_1224_74#_c_1257_n 0.00382767f $X=6.54 $Y=2.235
+ $X2=0 $Y2=0
cc_707 N_A_319_360#_M1003_g N_A_1224_74#_c_1237_n 0.0221333f $X=7.095 $Y=0.58
+ $X2=0 $Y2=0
cc_708 N_A_319_360#_c_947_n N_A_1224_74#_c_1238_n 0.00206465f $X=7.02 $Y=1.55
+ $X2=0 $Y2=0
cc_709 N_A_319_360#_M1003_g N_A_1224_74#_c_1238_n 0.0011854f $X=7.095 $Y=0.58
+ $X2=0 $Y2=0
cc_710 N_A_319_360#_c_947_n N_A_1224_74#_c_1239_n 0.00561544f $X=7.02 $Y=1.55
+ $X2=0 $Y2=0
cc_711 N_A_319_360#_M1003_g N_A_1224_74#_c_1239_n 0.00135722f $X=7.095 $Y=0.58
+ $X2=0 $Y2=0
cc_712 N_A_319_360#_c_947_n N_A_1224_74#_c_1240_n 3.07924e-19 $X=7.02 $Y=1.55
+ $X2=0 $Y2=0
cc_713 N_A_319_360#_c_955_n N_VPWR_c_1445_n 0.00963453f $X=2.415 $Y=1.725 $X2=0
+ $Y2=0
cc_714 N_A_319_360#_c_943_n N_VPWR_c_1445_n 0.00539724f $X=2.935 $Y=3.075 $X2=0
+ $Y2=0
cc_715 N_A_319_360#_c_960_n N_VPWR_c_1446_n 0.00604299f $X=3.905 $Y=2.9 $X2=0
+ $Y2=0
cc_716 N_A_319_360#_c_963_n N_VPWR_c_1446_n 0.0257522f $X=6.45 $Y=3.15 $X2=0
+ $Y2=0
cc_717 N_A_319_360#_c_963_n N_VPWR_c_1447_n 0.0213056f $X=6.45 $Y=3.15 $X2=0
+ $Y2=0
cc_718 N_A_319_360#_c_964_n N_VPWR_c_1447_n 0.00613773f $X=6.54 $Y=2.9 $X2=0
+ $Y2=0
cc_719 N_A_319_360#_M1032_g N_VPWR_c_1447_n 6.32588e-19 $X=6.54 $Y=2.235 $X2=0
+ $Y2=0
cc_720 N_A_319_360#_c_955_n N_VPWR_c_1454_n 0.00492531f $X=2.415 $Y=1.725 $X2=0
+ $Y2=0
cc_721 N_A_319_360#_c_959_n N_VPWR_c_1454_n 0.0456126f $X=3.01 $Y=3.15 $X2=0
+ $Y2=0
cc_722 N_A_319_360#_c_963_n N_VPWR_c_1455_n 0.0295821f $X=6.45 $Y=3.15 $X2=0
+ $Y2=0
cc_723 N_A_319_360#_c_963_n N_VPWR_c_1456_n 0.0193014f $X=6.45 $Y=3.15 $X2=0
+ $Y2=0
cc_724 N_A_319_360#_c_955_n N_VPWR_c_1441_n 0.00483326f $X=2.415 $Y=1.725 $X2=0
+ $Y2=0
cc_725 N_A_319_360#_c_958_n N_VPWR_c_1441_n 0.0241512f $X=3.815 $Y=3.15 $X2=0
+ $Y2=0
cc_726 N_A_319_360#_c_959_n N_VPWR_c_1441_n 0.00718166f $X=3.01 $Y=3.15 $X2=0
+ $Y2=0
cc_727 N_A_319_360#_c_963_n N_VPWR_c_1441_n 0.077543f $X=6.45 $Y=3.15 $X2=0
+ $Y2=0
cc_728 N_A_319_360#_c_969_n N_VPWR_c_1441_n 0.00536159f $X=3.905 $Y=3.15 $X2=0
+ $Y2=0
cc_729 N_A_319_360#_c_950_n N_A_38_78#_c_1582_n 0.0046003f $X=1.755 $Y=0.515
+ $X2=0 $Y2=0
cc_730 N_A_319_360#_c_954_n N_A_38_78#_c_1582_n 0.00548739f $X=1.695 $Y=1.055
+ $X2=0 $Y2=0
cc_731 N_A_319_360#_M1017_s N_A_38_78#_c_1588_n 0.0082374f $X=1.595 $Y=1.8 $X2=0
+ $Y2=0
cc_732 N_A_319_360#_c_955_n N_A_38_78#_c_1588_n 0.0126077f $X=2.415 $Y=1.725
+ $X2=0 $Y2=0
cc_733 N_A_319_360#_c_943_n N_A_38_78#_c_1588_n 0.0127092f $X=2.935 $Y=3.075
+ $X2=0 $Y2=0
cc_734 N_A_319_360#_c_971_n N_A_38_78#_c_1588_n 0.025151f $X=1.74 $Y=1.975 $X2=0
+ $Y2=0
cc_735 N_A_319_360#_c_942_n N_A_38_78#_c_1583_n 2.54456e-19 $X=2.54 $Y=1.185
+ $X2=0 $Y2=0
cc_736 N_A_319_360#_c_944_n N_A_38_78#_c_1583_n 0.00462134f $X=3.51 $Y=1.26
+ $X2=0 $Y2=0
cc_737 N_A_319_360#_M1020_g N_A_38_78#_c_1583_n 0.0109364f $X=3.585 $Y=0.8 $X2=0
+ $Y2=0
cc_738 N_A_319_360#_c_962_n N_A_38_78#_c_1589_n 0.00153498f $X=3.905 $Y=2.81
+ $X2=0 $Y2=0
cc_739 N_A_319_360#_c_945_n N_A_38_78#_c_1584_n 6.6894e-19 $X=3.01 $Y=1.26 $X2=0
+ $Y2=0
cc_740 N_A_319_360#_c_943_n N_A_38_78#_c_1592_n 0.0136255f $X=2.935 $Y=3.075
+ $X2=0 $Y2=0
cc_741 N_A_319_360#_c_958_n N_A_38_78#_c_1592_n 0.00570622f $X=3.815 $Y=3.15
+ $X2=0 $Y2=0
cc_742 N_A_319_360#_c_962_n N_A_38_78#_c_1592_n 5.94401e-19 $X=3.905 $Y=2.81
+ $X2=0 $Y2=0
cc_743 N_A_319_360#_c_944_n N_A_38_78#_c_1586_n 0.0151003f $X=3.51 $Y=1.26 $X2=0
+ $Y2=0
cc_744 N_A_319_360#_c_952_n N_VGND_M1002_d 0.00360404f $X=2.445 $Y=1.055 $X2=0
+ $Y2=0
cc_745 N_A_319_360#_c_950_n N_VGND_c_1738_n 0.0364619f $X=1.755 $Y=0.515 $X2=0
+ $Y2=0
cc_746 N_A_319_360#_c_950_n N_VGND_c_1739_n 0.0199184f $X=1.755 $Y=0.515 $X2=0
+ $Y2=0
cc_747 N_A_319_360#_c_942_n N_VGND_c_1740_n 0.0040978f $X=2.54 $Y=1.185 $X2=0
+ $Y2=0
cc_748 N_A_319_360#_c_950_n N_VGND_c_1740_n 0.018496f $X=1.755 $Y=0.515 $X2=0
+ $Y2=0
cc_749 N_A_319_360#_c_952_n N_VGND_c_1740_n 0.0248957f $X=2.445 $Y=1.055 $X2=0
+ $Y2=0
cc_750 N_A_319_360#_M1003_g N_VGND_c_1741_n 0.00154981f $X=7.095 $Y=0.58 $X2=0
+ $Y2=0
cc_751 N_A_319_360#_c_942_n N_VGND_c_1745_n 0.0043213f $X=2.54 $Y=1.185 $X2=0
+ $Y2=0
cc_752 N_A_319_360#_M1003_g N_VGND_c_1746_n 0.00309049f $X=7.095 $Y=0.58 $X2=0
+ $Y2=0
cc_753 N_A_319_360#_c_942_n N_VGND_c_1750_n 0.00825415f $X=2.54 $Y=1.185 $X2=0
+ $Y2=0
cc_754 N_A_319_360#_M1003_g N_VGND_c_1750_n 0.0040628f $X=7.095 $Y=0.58 $X2=0
+ $Y2=0
cc_755 N_A_319_360#_c_950_n N_VGND_c_1750_n 0.0164304f $X=1.755 $Y=0.515 $X2=0
+ $Y2=0
cc_756 N_A_1482_48#_c_1134_n N_A_1224_74#_M1031_g 0.0108008f $X=8.485 $Y=0.985
+ $X2=0 $Y2=0
cc_757 N_A_1482_48#_c_1135_n N_A_1224_74#_M1031_g 0.0132755f $X=8.65 $Y=0.58
+ $X2=0 $Y2=0
cc_758 N_A_1482_48#_c_1136_n N_A_1224_74#_M1031_g 0.00584201f $X=8.885 $Y=1.765
+ $X2=0 $Y2=0
cc_759 N_A_1482_48#_c_1138_n N_A_1224_74#_M1031_g 0.0045388f $X=8.727 $Y=0.985
+ $X2=0 $Y2=0
cc_760 N_A_1482_48#_c_1142_n N_A_1224_74#_c_1228_n 0.00705834f $X=8.555 $Y=2.335
+ $X2=0 $Y2=0
cc_761 N_A_1482_48#_c_1136_n N_A_1224_74#_c_1228_n 0.00407488f $X=8.885 $Y=1.765
+ $X2=0 $Y2=0
cc_762 N_A_1482_48#_c_1144_n N_A_1224_74#_c_1228_n 0.0144908f $X=8.885 $Y=1.85
+ $X2=0 $Y2=0
cc_763 N_A_1482_48#_c_1142_n N_A_1224_74#_c_1245_n 0.0115505f $X=8.555 $Y=2.335
+ $X2=0 $Y2=0
cc_764 N_A_1482_48#_c_1136_n N_A_1224_74#_c_1229_n 0.0256662f $X=8.885 $Y=1.765
+ $X2=0 $Y2=0
cc_765 N_A_1482_48#_c_1144_n N_A_1224_74#_c_1229_n 0.00384268f $X=8.885 $Y=1.85
+ $X2=0 $Y2=0
cc_766 N_A_1482_48#_c_1144_n N_A_1224_74#_c_1230_n 4.86873e-19 $X=8.885 $Y=1.85
+ $X2=0 $Y2=0
cc_767 N_A_1482_48#_c_1138_n N_A_1224_74#_c_1230_n 0.00795f $X=8.727 $Y=0.985
+ $X2=0 $Y2=0
cc_768 N_A_1482_48#_c_1142_n N_A_1224_74#_c_1231_n 5.60188e-19 $X=8.555 $Y=2.335
+ $X2=0 $Y2=0
cc_769 N_A_1482_48#_c_1136_n N_A_1224_74#_c_1231_n 0.00210772f $X=8.885 $Y=1.765
+ $X2=0 $Y2=0
cc_770 N_A_1482_48#_c_1144_n N_A_1224_74#_c_1231_n 0.00185013f $X=8.885 $Y=1.85
+ $X2=0 $Y2=0
cc_771 N_A_1482_48#_c_1135_n N_A_1224_74#_M1014_g 0.00122775f $X=8.65 $Y=0.58
+ $X2=0 $Y2=0
cc_772 N_A_1482_48#_c_1136_n N_A_1224_74#_M1014_g 0.00251042f $X=8.885 $Y=1.765
+ $X2=0 $Y2=0
cc_773 N_A_1482_48#_c_1132_n N_A_1224_74#_c_1277_n 0.0012657f $X=7.485 $Y=0.9
+ $X2=0 $Y2=0
cc_774 N_A_1482_48#_c_1141_n N_A_1224_74#_c_1257_n 0.00944193f $X=7.67 $Y=2.28
+ $X2=0 $Y2=0
cc_775 N_A_1482_48#_c_1132_n N_A_1224_74#_c_1237_n 0.00230939f $X=7.485 $Y=0.9
+ $X2=0 $Y2=0
cc_776 N_A_1482_48#_c_1133_n N_A_1224_74#_c_1237_n 0.00111943f $X=7.67 $Y=2.19
+ $X2=0 $Y2=0
cc_777 N_A_1482_48#_c_1137_n N_A_1224_74#_c_1237_n 0.0162835f $X=7.595 $Y=0.985
+ $X2=0 $Y2=0
cc_778 N_A_1482_48#_c_1137_n N_A_1224_74#_c_1238_n 0.00432309f $X=7.595 $Y=0.985
+ $X2=0 $Y2=0
cc_779 N_A_1482_48#_c_1139_n N_A_1224_74#_c_1238_n 0.00127859f $X=7.67 $Y=1.065
+ $X2=0 $Y2=0
cc_780 N_A_1482_48#_c_1133_n N_A_1224_74#_c_1240_n 0.0153989f $X=7.67 $Y=2.19
+ $X2=0 $Y2=0
cc_781 N_A_1482_48#_c_1141_n N_A_1224_74#_c_1240_n 0.00481867f $X=7.67 $Y=2.28
+ $X2=0 $Y2=0
cc_782 N_A_1482_48#_c_1133_n N_A_1224_74#_c_1241_n 0.00617973f $X=7.67 $Y=2.19
+ $X2=0 $Y2=0
cc_783 N_A_1482_48#_c_1134_n N_A_1224_74#_c_1241_n 0.0246405f $X=8.485 $Y=0.985
+ $X2=0 $Y2=0
cc_784 N_A_1482_48#_c_1137_n N_A_1224_74#_c_1241_n 0.00601156f $X=7.595 $Y=0.985
+ $X2=0 $Y2=0
cc_785 N_A_1482_48#_c_1133_n N_A_1224_74#_c_1242_n 0.0053332f $X=7.67 $Y=2.19
+ $X2=0 $Y2=0
cc_786 N_A_1482_48#_c_1137_n N_A_1224_74#_c_1242_n 0.0125972f $X=7.595 $Y=0.985
+ $X2=0 $Y2=0
cc_787 N_A_1482_48#_c_1139_n N_A_1224_74#_c_1242_n 6.55449e-19 $X=7.67 $Y=1.065
+ $X2=0 $Y2=0
cc_788 N_A_1482_48#_c_1134_n N_A_1224_74#_c_1243_n 0.00997859f $X=8.485 $Y=0.985
+ $X2=0 $Y2=0
cc_789 N_A_1482_48#_c_1136_n N_A_1224_74#_c_1243_n 0.0233867f $X=8.885 $Y=1.765
+ $X2=0 $Y2=0
cc_790 N_A_1482_48#_c_1144_n N_A_1224_74#_c_1243_n 0.0116759f $X=8.885 $Y=1.85
+ $X2=0 $Y2=0
cc_791 N_A_1482_48#_c_1138_n N_A_1224_74#_c_1243_n 0.0109402f $X=8.727 $Y=0.985
+ $X2=0 $Y2=0
cc_792 N_A_1482_48#_c_1144_n N_VPWR_M1019_d 0.00365297f $X=8.885 $Y=1.85 $X2=0
+ $Y2=0
cc_793 N_A_1482_48#_c_1141_n N_VPWR_c_1448_n 0.00610146f $X=7.67 $Y=2.28 $X2=0
+ $Y2=0
cc_794 N_A_1482_48#_c_1142_n N_VPWR_c_1448_n 0.00131777f $X=8.555 $Y=2.335 $X2=0
+ $Y2=0
cc_795 N_A_1482_48#_c_1142_n N_VPWR_c_1449_n 0.00646407f $X=8.555 $Y=2.335 $X2=0
+ $Y2=0
cc_796 N_A_1482_48#_c_1142_n N_VPWR_c_1450_n 0.0463782f $X=8.555 $Y=2.335 $X2=0
+ $Y2=0
cc_797 N_A_1482_48#_c_1144_n N_VPWR_c_1450_n 0.012936f $X=8.885 $Y=1.85 $X2=0
+ $Y2=0
cc_798 N_A_1482_48#_c_1141_n N_VPWR_c_1456_n 0.00405364f $X=7.67 $Y=2.28 $X2=0
+ $Y2=0
cc_799 N_A_1482_48#_c_1141_n N_VPWR_c_1441_n 0.00489211f $X=7.67 $Y=2.28 $X2=0
+ $Y2=0
cc_800 N_A_1482_48#_c_1142_n N_VPWR_c_1441_n 0.011426f $X=8.555 $Y=2.335 $X2=0
+ $Y2=0
cc_801 N_A_1482_48#_c_1136_n N_Q_N_c_1691_n 0.018767f $X=8.885 $Y=1.765 $X2=0
+ $Y2=0
cc_802 N_A_1482_48#_c_1144_n N_Q_N_c_1691_n 0.00158159f $X=8.885 $Y=1.85 $X2=0
+ $Y2=0
cc_803 N_A_1482_48#_c_1144_n N_Q_N_c_1694_n 0.00456533f $X=8.885 $Y=1.85 $X2=0
+ $Y2=0
cc_804 N_A_1482_48#_c_1132_n N_VGND_c_1741_n 0.0147674f $X=7.485 $Y=0.9 $X2=0
+ $Y2=0
cc_805 N_A_1482_48#_c_1134_n N_VGND_c_1741_n 0.0137782f $X=8.485 $Y=0.985 $X2=0
+ $Y2=0
cc_806 N_A_1482_48#_c_1135_n N_VGND_c_1741_n 0.0110441f $X=8.65 $Y=0.58 $X2=0
+ $Y2=0
cc_807 N_A_1482_48#_c_1137_n N_VGND_c_1741_n 0.0129689f $X=7.595 $Y=0.985 $X2=0
+ $Y2=0
cc_808 N_A_1482_48#_c_1139_n N_VGND_c_1741_n 0.00131228f $X=7.67 $Y=1.065 $X2=0
+ $Y2=0
cc_809 N_A_1482_48#_c_1135_n N_VGND_c_1742_n 0.0454165f $X=8.65 $Y=0.58 $X2=0
+ $Y2=0
cc_810 N_A_1482_48#_c_1136_n N_VGND_c_1742_n 0.00455872f $X=8.885 $Y=1.765 $X2=0
+ $Y2=0
cc_811 N_A_1482_48#_c_1138_n N_VGND_c_1742_n 0.0145003f $X=8.727 $Y=0.985 $X2=0
+ $Y2=0
cc_812 N_A_1482_48#_c_1132_n N_VGND_c_1746_n 0.00383152f $X=7.485 $Y=0.9 $X2=0
+ $Y2=0
cc_813 N_A_1482_48#_c_1135_n N_VGND_c_1747_n 0.0215384f $X=8.65 $Y=0.58 $X2=0
+ $Y2=0
cc_814 N_A_1482_48#_c_1132_n N_VGND_c_1750_n 0.0075725f $X=7.485 $Y=0.9 $X2=0
+ $Y2=0
cc_815 N_A_1482_48#_c_1135_n N_VGND_c_1750_n 0.0177458f $X=8.65 $Y=0.58 $X2=0
+ $Y2=0
cc_816 N_A_1224_74#_M1012_g N_A_2026_424#_M1009_g 0.0197956f $X=10.515 $Y=0.645
+ $X2=0 $Y2=0
cc_817 N_A_1224_74#_c_1234_n N_A_2026_424#_c_1392_n 0.00994164f $X=10.5 $Y=1.955
+ $X2=0 $Y2=0
cc_818 N_A_1224_74#_c_1248_n N_A_2026_424#_c_1392_n 0.00588428f $X=10.5 $Y=2.045
+ $X2=0 $Y2=0
cc_819 N_A_1224_74#_c_1236_n N_A_2026_424#_c_1392_n 0.0214662f $X=10.5 $Y=1.43
+ $X2=0 $Y2=0
cc_820 N_A_1224_74#_c_1233_n N_A_2026_424#_c_1393_n 0.00517977f $X=10.41 $Y=1.43
+ $X2=0 $Y2=0
cc_821 N_A_1224_74#_M1012_g N_A_2026_424#_c_1393_n 0.0146713f $X=10.515 $Y=0.645
+ $X2=0 $Y2=0
cc_822 N_A_1224_74#_c_1236_n N_A_2026_424#_c_1393_n 6.73726e-19 $X=10.5 $Y=1.43
+ $X2=0 $Y2=0
cc_823 N_A_1224_74#_c_1234_n N_A_2026_424#_c_1394_n 0.0112992f $X=10.5 $Y=1.955
+ $X2=0 $Y2=0
cc_824 N_A_1224_74#_c_1248_n N_A_2026_424#_c_1394_n 0.0166377f $X=10.5 $Y=2.045
+ $X2=0 $Y2=0
cc_825 N_A_1224_74#_c_1234_n N_A_2026_424#_c_1395_n 0.00782285f $X=10.5 $Y=1.955
+ $X2=0 $Y2=0
cc_826 N_A_1224_74#_c_1236_n N_A_2026_424#_c_1395_n 0.0139388f $X=10.5 $Y=1.43
+ $X2=0 $Y2=0
cc_827 N_A_1224_74#_c_1233_n N_A_2026_424#_c_1396_n 0.0166486f $X=10.41 $Y=1.43
+ $X2=0 $Y2=0
cc_828 N_A_1224_74#_c_1234_n N_A_2026_424#_c_1396_n 7.34008e-19 $X=10.5 $Y=1.955
+ $X2=0 $Y2=0
cc_829 N_A_1224_74#_c_1236_n N_A_2026_424#_c_1396_n 8.33355e-19 $X=10.5 $Y=1.43
+ $X2=0 $Y2=0
cc_830 N_A_1224_74#_c_1257_n N_VPWR_c_1448_n 0.0264538f $X=7.495 $Y=2.53 $X2=0
+ $Y2=0
cc_831 N_A_1224_74#_c_1240_n N_VPWR_c_1448_n 0.0021468f $X=7.58 $Y=2.365 $X2=0
+ $Y2=0
cc_832 N_A_1224_74#_c_1245_n N_VPWR_c_1449_n 0.00393528f $X=8.63 $Y=2.28 $X2=0
+ $Y2=0
cc_833 N_A_1224_74#_c_1228_n N_VPWR_c_1450_n 0.0013401f $X=8.63 $Y=2.19 $X2=0
+ $Y2=0
cc_834 N_A_1224_74#_c_1245_n N_VPWR_c_1450_n 0.00764221f $X=8.63 $Y=2.28 $X2=0
+ $Y2=0
cc_835 N_A_1224_74#_c_1229_n N_VPWR_c_1450_n 0.00151008f $X=9.055 $Y=1.43 $X2=0
+ $Y2=0
cc_836 N_A_1224_74#_c_1231_n N_VPWR_c_1450_n 0.00556331f $X=9.145 $Y=1.765 $X2=0
+ $Y2=0
cc_837 N_A_1224_74#_c_1234_n N_VPWR_c_1451_n 0.00204674f $X=10.5 $Y=1.955 $X2=0
+ $Y2=0
cc_838 N_A_1224_74#_c_1248_n N_VPWR_c_1451_n 0.00449437f $X=10.5 $Y=2.045 $X2=0
+ $Y2=0
cc_839 N_A_1224_74#_c_1257_n N_VPWR_c_1456_n 0.0159863f $X=7.495 $Y=2.53 $X2=0
+ $Y2=0
cc_840 N_A_1224_74#_c_1231_n N_VPWR_c_1457_n 0.00461464f $X=9.145 $Y=1.765 $X2=0
+ $Y2=0
cc_841 N_A_1224_74#_c_1248_n N_VPWR_c_1457_n 0.00445665f $X=10.5 $Y=2.045 $X2=0
+ $Y2=0
cc_842 N_A_1224_74#_c_1245_n N_VPWR_c_1441_n 0.00489211f $X=8.63 $Y=2.28 $X2=0
+ $Y2=0
cc_843 N_A_1224_74#_c_1231_n N_VPWR_c_1441_n 0.00918106f $X=9.145 $Y=1.765 $X2=0
+ $Y2=0
cc_844 N_A_1224_74#_c_1248_n N_VPWR_c_1441_n 0.00862405f $X=10.5 $Y=2.045 $X2=0
+ $Y2=0
cc_845 N_A_1224_74#_c_1257_n N_VPWR_c_1441_n 0.0282176f $X=7.495 $Y=2.53 $X2=0
+ $Y2=0
cc_846 N_A_1224_74#_c_1257_n A_1465_471# 0.00449141f $X=7.495 $Y=2.53 $X2=-0.19
+ $Y2=-0.245
cc_847 N_A_1224_74#_c_1231_n N_Q_N_c_1691_n 0.0044298f $X=9.145 $Y=1.765 $X2=0
+ $Y2=0
cc_848 N_A_1224_74#_M1014_g N_Q_N_c_1691_n 0.0191689f $X=9.44 $Y=0.74 $X2=0
+ $Y2=0
cc_849 N_A_1224_74#_c_1233_n N_Q_N_c_1691_n 0.0449729f $X=10.41 $Y=1.43 $X2=0
+ $Y2=0
cc_850 N_A_1224_74#_c_1234_n N_Q_N_c_1691_n 0.0010753f $X=10.5 $Y=1.955 $X2=0
+ $Y2=0
cc_851 N_A_1224_74#_c_1231_n N_Q_N_c_1694_n 0.014297f $X=9.145 $Y=1.765 $X2=0
+ $Y2=0
cc_852 N_A_1224_74#_c_1248_n N_Q_N_c_1694_n 0.00385512f $X=10.5 $Y=2.045 $X2=0
+ $Y2=0
cc_853 N_A_1224_74#_M1031_g N_VGND_c_1741_n 0.0014914f $X=8.435 $Y=0.58 $X2=0
+ $Y2=0
cc_854 N_A_1224_74#_c_1277_n N_VGND_c_1741_n 0.0120929f $X=6.99 $Y=0.565 $X2=0
+ $Y2=0
cc_855 N_A_1224_74#_M1031_g N_VGND_c_1742_n 0.00378178f $X=8.435 $Y=0.58 $X2=0
+ $Y2=0
cc_856 N_A_1224_74#_c_1231_n N_VGND_c_1742_n 0.00633828f $X=9.145 $Y=1.765 $X2=0
+ $Y2=0
cc_857 N_A_1224_74#_M1014_g N_VGND_c_1742_n 0.017876f $X=9.44 $Y=0.74 $X2=0
+ $Y2=0
cc_858 N_A_1224_74#_M1012_g N_VGND_c_1743_n 0.00770628f $X=10.515 $Y=0.645 $X2=0
+ $Y2=0
cc_859 N_A_1224_74#_c_1277_n N_VGND_c_1746_n 0.0242914f $X=6.99 $Y=0.565 $X2=0
+ $Y2=0
cc_860 N_A_1224_74#_M1031_g N_VGND_c_1747_n 0.00434272f $X=8.435 $Y=0.58 $X2=0
+ $Y2=0
cc_861 N_A_1224_74#_M1014_g N_VGND_c_1748_n 0.00383152f $X=9.44 $Y=0.74 $X2=0
+ $Y2=0
cc_862 N_A_1224_74#_M1012_g N_VGND_c_1748_n 0.00461464f $X=10.515 $Y=0.645 $X2=0
+ $Y2=0
cc_863 N_A_1224_74#_M1031_g N_VGND_c_1750_n 0.00825979f $X=8.435 $Y=0.58 $X2=0
+ $Y2=0
cc_864 N_A_1224_74#_M1014_g N_VGND_c_1750_n 0.00762539f $X=9.44 $Y=0.74 $X2=0
+ $Y2=0
cc_865 N_A_1224_74#_M1012_g N_VGND_c_1750_n 0.00914043f $X=10.515 $Y=0.645 $X2=0
+ $Y2=0
cc_866 N_A_1224_74#_c_1277_n N_VGND_c_1750_n 0.02509f $X=6.99 $Y=0.565 $X2=0
+ $Y2=0
cc_867 N_A_2026_424#_c_1392_n N_VPWR_c_1451_n 0.00610705f $X=11.015 $Y=1.765
+ $X2=0 $Y2=0
cc_868 N_A_2026_424#_c_1394_n N_VPWR_c_1451_n 0.0542643f $X=10.275 $Y=2.27 $X2=0
+ $Y2=0
cc_869 N_A_2026_424#_c_1395_n N_VPWR_c_1451_n 0.0235211f $X=10.965 $Y=1.465
+ $X2=0 $Y2=0
cc_870 N_A_2026_424#_c_1394_n N_VPWR_c_1457_n 0.0108068f $X=10.275 $Y=2.27 $X2=0
+ $Y2=0
cc_871 N_A_2026_424#_c_1392_n N_VPWR_c_1458_n 0.00445602f $X=11.015 $Y=1.765
+ $X2=0 $Y2=0
cc_872 N_A_2026_424#_c_1392_n N_VPWR_c_1441_n 0.00861048f $X=11.015 $Y=1.765
+ $X2=0 $Y2=0
cc_873 N_A_2026_424#_c_1394_n N_VPWR_c_1441_n 0.00906421f $X=10.275 $Y=2.27
+ $X2=0 $Y2=0
cc_874 N_A_2026_424#_c_1393_n N_Q_N_c_1691_n 0.0605318f $X=10.3 $Y=0.64 $X2=0
+ $Y2=0
cc_875 N_A_2026_424#_c_1394_n N_Q_N_c_1691_n 0.0894769f $X=10.275 $Y=2.27 $X2=0
+ $Y2=0
cc_876 N_A_2026_424#_c_1396_n N_Q_N_c_1691_n 0.0205307f $X=10.315 $Y=1.465 $X2=0
+ $Y2=0
cc_877 N_A_2026_424#_M1009_g Q 0.00795463f $X=11.015 $Y=0.74 $X2=0 $Y2=0
cc_878 N_A_2026_424#_M1009_g Q 0.00263483f $X=11.015 $Y=0.74 $X2=0 $Y2=0
cc_879 N_A_2026_424#_c_1392_n Q 0.00169664f $X=11.015 $Y=1.765 $X2=0 $Y2=0
cc_880 N_A_2026_424#_c_1395_n Q 0.00233746f $X=10.965 $Y=1.465 $X2=0 $Y2=0
cc_881 N_A_2026_424#_c_1392_n Q 0.00408255f $X=11.015 $Y=1.765 $X2=0 $Y2=0
cc_882 N_A_2026_424#_c_1395_n Q 0.00140951f $X=10.965 $Y=1.465 $X2=0 $Y2=0
cc_883 N_A_2026_424#_c_1392_n Q 0.0109295f $X=11.015 $Y=1.765 $X2=0 $Y2=0
cc_884 N_A_2026_424#_M1009_g N_Q_c_1717_n 0.00406947f $X=11.015 $Y=0.74 $X2=0
+ $Y2=0
cc_885 N_A_2026_424#_c_1392_n N_Q_c_1717_n 0.0126603f $X=11.015 $Y=1.765 $X2=0
+ $Y2=0
cc_886 N_A_2026_424#_c_1395_n N_Q_c_1717_n 0.0262113f $X=10.965 $Y=1.465 $X2=0
+ $Y2=0
cc_887 N_A_2026_424#_M1009_g N_VGND_c_1743_n 0.00357902f $X=11.015 $Y=0.74 $X2=0
+ $Y2=0
cc_888 N_A_2026_424#_c_1392_n N_VGND_c_1743_n 0.00218979f $X=11.015 $Y=1.765
+ $X2=0 $Y2=0
cc_889 N_A_2026_424#_c_1393_n N_VGND_c_1743_n 0.0295846f $X=10.3 $Y=0.64 $X2=0
+ $Y2=0
cc_890 N_A_2026_424#_c_1395_n N_VGND_c_1743_n 0.0215504f $X=10.965 $Y=1.465
+ $X2=0 $Y2=0
cc_891 N_A_2026_424#_c_1393_n N_VGND_c_1748_n 0.011066f $X=10.3 $Y=0.64 $X2=0
+ $Y2=0
cc_892 N_A_2026_424#_M1009_g N_VGND_c_1749_n 0.00434272f $X=11.015 $Y=0.74 $X2=0
+ $Y2=0
cc_893 N_A_2026_424#_M1009_g N_VGND_c_1750_n 0.00824463f $X=11.015 $Y=0.74 $X2=0
+ $Y2=0
cc_894 N_A_2026_424#_c_1393_n N_VGND_c_1750_n 0.00915947f $X=10.3 $Y=0.64 $X2=0
+ $Y2=0
cc_895 N_VPWR_M1017_d N_A_38_78#_c_1588_n 0.00485884f $X=2.04 $Y=1.8 $X2=0 $Y2=0
cc_896 N_VPWR_c_1444_n N_A_38_78#_c_1588_n 0.0193188f $X=1.18 $Y=2.815 $X2=0
+ $Y2=0
cc_897 N_VPWR_c_1445_n N_A_38_78#_c_1588_n 0.0162579f $X=2.19 $Y=2.755 $X2=0
+ $Y2=0
cc_898 N_VPWR_c_1441_n N_A_38_78#_c_1588_n 0.0532271f $X=11.28 $Y=3.33 $X2=0
+ $Y2=0
cc_899 N_VPWR_c_1443_n N_A_38_78#_c_1591_n 0.0310355f $X=0.28 $Y=2.75 $X2=0
+ $Y2=0
cc_900 N_VPWR_c_1444_n N_A_38_78#_c_1591_n 0.0222518f $X=1.18 $Y=2.815 $X2=0
+ $Y2=0
cc_901 N_VPWR_c_1452_n N_A_38_78#_c_1591_n 0.0144812f $X=1.095 $Y=3.33 $X2=0
+ $Y2=0
cc_902 N_VPWR_c_1441_n N_A_38_78#_c_1591_n 0.0119834f $X=11.28 $Y=3.33 $X2=0
+ $Y2=0
cc_903 N_VPWR_c_1454_n N_A_38_78#_c_1592_n 0.00751951f $X=4.44 $Y=3.33 $X2=0
+ $Y2=0
cc_904 N_VPWR_c_1441_n N_A_38_78#_c_1592_n 0.00908407f $X=11.28 $Y=3.33 $X2=0
+ $Y2=0
cc_905 N_VPWR_c_1450_n Q_N 0.00163554f $X=8.92 $Y=2.27 $X2=0 $Y2=0
cc_906 N_VPWR_c_1451_n Q_N 3.35434e-19 $X=10.79 $Y=1.985 $X2=0 $Y2=0
cc_907 N_VPWR_c_1457_n Q_N 0.0313273f $X=10.61 $Y=3.33 $X2=0 $Y2=0
cc_908 N_VPWR_c_1441_n Q_N 0.0254862f $X=11.28 $Y=3.33 $X2=0 $Y2=0
cc_909 N_VPWR_c_1451_n Q 0.0456259f $X=10.79 $Y=1.985 $X2=0 $Y2=0
cc_910 N_VPWR_c_1458_n Q 0.0159324f $X=11.28 $Y=3.33 $X2=0 $Y2=0
cc_911 N_VPWR_c_1441_n Q 0.0131546f $X=11.28 $Y=3.33 $X2=0 $Y2=0
cc_912 N_A_38_78#_c_1581_n A_125_78# 0.00236678f $X=0.69 $Y=0.745 $X2=-0.19
+ $Y2=-0.245
cc_913 N_A_38_78#_c_1581_n N_VGND_c_1738_n 0.00157034f $X=0.69 $Y=0.745 $X2=0
+ $Y2=0
cc_914 N_A_38_78#_c_1585_n N_VGND_c_1738_n 0.00465719f $X=0.335 $Y=0.6 $X2=0
+ $Y2=0
cc_915 N_A_38_78#_c_1581_n N_VGND_c_1744_n 0.00520932f $X=0.69 $Y=0.745 $X2=0
+ $Y2=0
cc_916 N_A_38_78#_c_1585_n N_VGND_c_1744_n 0.0131067f $X=0.335 $Y=0.6 $X2=0
+ $Y2=0
cc_917 N_A_38_78#_c_1581_n N_VGND_c_1750_n 0.0102476f $X=0.69 $Y=0.745 $X2=0
+ $Y2=0
cc_918 N_A_38_78#_c_1585_n N_VGND_c_1750_n 0.0117869f $X=0.335 $Y=0.6 $X2=0
+ $Y2=0
cc_919 N_Q_N_c_1691_n N_VGND_c_1742_n 0.0296698f $X=9.725 $Y=0.515 $X2=0 $Y2=0
cc_920 N_Q_N_c_1694_n N_VGND_c_1742_n 0.00437693f $X=9.37 $Y=1.985 $X2=0 $Y2=0
cc_921 N_Q_N_c_1691_n N_VGND_c_1748_n 0.0173129f $X=9.725 $Y=0.515 $X2=0 $Y2=0
cc_922 N_Q_N_c_1691_n N_VGND_c_1750_n 0.0143301f $X=9.725 $Y=0.515 $X2=0 $Y2=0
cc_923 Q N_VGND_c_1743_n 0.0312622f $X=11.195 $Y=0.47 $X2=0 $Y2=0
cc_924 Q N_VGND_c_1749_n 0.0163488f $X=11.195 $Y=0.47 $X2=0 $Y2=0
cc_925 Q N_VGND_c_1750_n 0.0134757f $X=11.195 $Y=0.47 $X2=0 $Y2=0
