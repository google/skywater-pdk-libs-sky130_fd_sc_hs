* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hs__nand2b_1 A_N B VGND VNB VPB VPWR Y
M1000 Y a_27_112# a_269_74# VNB nlowvt w=740000u l=150000u
+  ad=3.182e+11p pd=2.34e+06u as=1.776e+11p ps=1.96e+06u
M1001 a_269_74# B VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=4.4825e+11p ps=2.73e+06u
M1002 VPWR a_27_112# Y VPB pshort w=1.12e+06u l=150000u
+  ad=8.932e+11p pd=6.12e+06u as=3.92e+11p ps=2.94e+06u
M1003 Y B VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 VGND A_N a_27_112# VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=1.5675e+11p ps=1.67e+06u
M1005 VPWR A_N a_27_112# VPB pshort w=840000u l=150000u
+  ad=0p pd=0u as=2.478e+11p ps=2.27e+06u
.ends
