* File: sky130_fd_sc_hs__a311o_4.pex.spice
* Created: Thu Aug 27 20:28:39 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HS__A311O_4%C1 1 3 6 8 10 13 15 22
r60 22 23 7.49223 $w=3.86e-07 $l=6e-08 $layer=POLY_cond $X=1.145 $Y=1.662
+ $X2=1.205 $Y2=1.662
r61 21 22 46.2021 $w=3.86e-07 $l=3.7e-07 $layer=POLY_cond $X=0.775 $Y=1.662
+ $X2=1.145 $Y2=1.662
r62 20 21 9.98964 $w=3.86e-07 $l=8e-08 $layer=POLY_cond $X=0.695 $Y=1.662
+ $X2=0.775 $Y2=1.662
r63 18 20 4.37047 $w=3.86e-07 $l=3.5e-08 $layer=POLY_cond $X=0.66 $Y=1.662
+ $X2=0.695 $Y2=1.662
r64 15 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.66
+ $Y=1.635 $X2=0.66 $Y2=1.635
r65 11 23 24.9932 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=1.205 $Y=1.44
+ $X2=1.205 $Y2=1.662
r66 11 13 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=1.205 $Y=1.44
+ $X2=1.205 $Y2=0.73
r67 8 22 24.9932 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=1.145 $Y=1.885
+ $X2=1.145 $Y2=1.662
r68 8 10 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=1.145 $Y=1.885
+ $X2=1.145 $Y2=2.46
r69 4 21 24.9932 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=0.775 $Y=1.44
+ $X2=0.775 $Y2=1.662
r70 4 6 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=0.775 $Y=1.44
+ $X2=0.775 $Y2=0.73
r71 1 20 24.9932 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=0.695 $Y=1.885
+ $X2=0.695 $Y2=1.662
r72 1 3 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=0.695 $Y=1.885
+ $X2=0.695 $Y2=2.46
.ends

.subckt PM_SKY130_FD_SC_HS__A311O_4%B1 1 3 6 8 10 13 15 22
c62 1 0 1.22191e-19 $X=1.595 $Y=1.885
r63 22 23 2.56383 $w=3.76e-07 $l=2e-08 $layer=POLY_cond $X=2.045 $Y=1.677
+ $X2=2.065 $Y2=1.677
r64 20 22 44.2261 $w=3.76e-07 $l=3.45e-07 $layer=POLY_cond $X=1.7 $Y=1.677
+ $X2=2.045 $Y2=1.677
r65 18 20 8.33245 $w=3.76e-07 $l=6.5e-08 $layer=POLY_cond $X=1.635 $Y=1.677
+ $X2=1.7 $Y2=1.677
r66 17 18 5.12766 $w=3.76e-07 $l=4e-08 $layer=POLY_cond $X=1.595 $Y=1.677
+ $X2=1.635 $Y2=1.677
r67 15 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.7
+ $Y=1.635 $X2=1.7 $Y2=1.635
r68 11 23 24.356 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.065 $Y=1.47
+ $X2=2.065 $Y2=1.677
r69 11 13 379.447 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=2.065 $Y=1.47
+ $X2=2.065 $Y2=0.73
r70 8 22 24.356 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=2.045 $Y=1.885
+ $X2=2.045 $Y2=1.677
r71 8 10 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=2.045 $Y=1.885
+ $X2=2.045 $Y2=2.46
r72 4 18 24.356 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.635 $Y=1.47
+ $X2=1.635 $Y2=1.677
r73 4 6 379.447 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=1.635 $Y=1.47
+ $X2=1.635 $Y2=0.73
r74 1 17 24.356 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=1.595 $Y=1.885
+ $X2=1.595 $Y2=1.677
r75 1 3 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=1.595 $Y=1.885
+ $X2=1.595 $Y2=2.46
.ends

.subckt PM_SKY130_FD_SC_HS__A311O_4%A_154_392# 1 2 3 4 15 19 21 23 26 28 30 33
+ 35 37 38 39 40 42 45 48 49 53 56 60 63 64 65 67 71 73 76 78 82
c213 71 0 1.22191e-19 $X=1.08 $Y=2.105
c214 64 0 5.4224e-20 $X=5.545 $Y=2.035
c215 63 0 1.44209e-19 $X=4.56 $Y=1.95
c216 53 0 1.88456e-19 $X=1.85 $Y=0.555
c217 40 0 1.37258e-19 $X=4.365 $Y=1.765
c218 38 0 1.4091e-19 $X=4.275 $Y=1.675
r219 91 92 4.43218 $w=4.35e-07 $l=4e-08 $layer=POLY_cond $X=3.875 $Y=1.542
+ $X2=3.915 $Y2=1.542
r220 88 89 2.21609 $w=4.35e-07 $l=2e-08 $layer=POLY_cond $X=3.445 $Y=1.542
+ $X2=3.465 $Y2=1.542
r221 87 88 47.646 $w=4.35e-07 $l=4.3e-07 $layer=POLY_cond $X=3.015 $Y=1.542
+ $X2=3.445 $Y2=1.542
r222 86 87 4.98621 $w=4.35e-07 $l=4.5e-08 $layer=POLY_cond $X=2.97 $Y=1.542
+ $X2=3.015 $Y2=1.542
r223 79 82 13.6198 $w=3.28e-07 $l=3.9e-07 $layer=LI1_cond $X=5.63 $Y=1.1
+ $X2=6.02 $Y2=1.1
r224 77 91 14.9586 $w=4.35e-07 $l=1.35e-07 $layer=POLY_cond $X=3.74 $Y=1.542
+ $X2=3.875 $Y2=1.542
r225 77 89 30.4713 $w=4.35e-07 $l=2.75e-07 $layer=POLY_cond $X=3.74 $Y=1.542
+ $X2=3.465 $Y2=1.542
r226 76 78 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=3.74 $Y=1.485
+ $X2=3.905 $Y2=1.485
r227 76 77 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.74
+ $Y=1.485 $X2=3.74 $Y2=1.485
r228 69 71 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=0.92 $Y=2.105
+ $X2=1.08 $Y2=2.105
r229 66 79 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.63 $Y=1.265
+ $X2=5.63 $Y2=1.1
r230 66 67 44.6898 $w=1.68e-07 $l=6.85e-07 $layer=LI1_cond $X=5.63 $Y=1.265
+ $X2=5.63 $Y2=1.95
r231 64 67 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.545 $Y=2.035
+ $X2=5.63 $Y2=1.95
r232 64 65 58.7166 $w=1.68e-07 $l=9e-07 $layer=LI1_cond $X=5.545 $Y=2.035
+ $X2=4.645 $Y2=2.035
r233 63 65 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.56 $Y=1.95
+ $X2=4.645 $Y2=2.035
r234 62 63 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=4.56 $Y=1.65 $X2=4.56
+ $Y2=1.95
r235 60 62 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.475 $Y=1.565
+ $X2=4.56 $Y2=1.65
r236 60 78 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=4.475 $Y=1.565
+ $X2=3.905 $Y2=1.565
r237 59 86 27.7011 $w=4.35e-07 $l=2.5e-07 $layer=POLY_cond $X=2.72 $Y=1.542
+ $X2=2.97 $Y2=1.542
r238 59 84 19.9448 $w=4.35e-07 $l=1.8e-07 $layer=POLY_cond $X=2.72 $Y=1.542
+ $X2=2.54 $Y2=1.542
r239 58 76 35.621 $w=3.28e-07 $l=1.02e-06 $layer=LI1_cond $X=2.72 $Y=1.485
+ $X2=3.74 $Y2=1.485
r240 58 59 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.72
+ $Y=1.485 $X2=2.72 $Y2=1.485
r241 56 58 13.7944 $w=3.28e-07 $l=3.95e-07 $layer=LI1_cond $X=2.325 $Y=1.485
+ $X2=2.72 $Y2=1.485
r242 51 56 17.4806 $w=3.35e-07 $l=6.33088e-07 $layer=LI1_cond $X=1.845 $Y=1.13
+ $X2=2.325 $Y2=1.485
r243 51 53 35.4293 $w=1.78e-07 $l=5.75e-07 $layer=LI1_cond $X=1.845 $Y=1.13
+ $X2=1.845 $Y2=0.555
r244 50 73 1.44715 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.165 $Y=1.215
+ $X2=1.035 $Y2=1.215
r245 49 51 6.23108 $w=3.35e-07 $l=1.25499e-07 $layer=LI1_cond $X=1.755 $Y=1.215
+ $X2=1.845 $Y2=1.13
r246 49 50 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=1.755 $Y=1.215
+ $X2=1.165 $Y2=1.215
r247 48 71 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.08 $Y=2.02
+ $X2=1.08 $Y2=2.105
r248 47 73 5.04255 $w=1.75e-07 $l=1.05119e-07 $layer=LI1_cond $X=1.08 $Y=1.3
+ $X2=1.035 $Y2=1.215
r249 47 48 46.9733 $w=1.68e-07 $l=7.2e-07 $layer=LI1_cond $X=1.08 $Y=1.3
+ $X2=1.08 $Y2=2.02
r250 43 73 5.04255 $w=1.75e-07 $l=1.03078e-07 $layer=LI1_cond $X=0.995 $Y=1.13
+ $X2=1.035 $Y2=1.215
r251 43 45 35.4293 $w=1.78e-07 $l=5.75e-07 $layer=LI1_cond $X=0.995 $Y=1.13
+ $X2=0.995 $Y2=0.555
r252 40 42 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=4.365 $Y=1.765
+ $X2=4.365 $Y2=2.4
r253 39 92 32.0209 $w=4.35e-07 $l=1.72218e-07 $layer=POLY_cond $X=4.005 $Y=1.675
+ $X2=3.915 $Y2=1.542
r254 38 40 26.9307 $w=1.5e-07 $l=1.27279e-07 $layer=POLY_cond $X=4.275 $Y=1.675
+ $X2=4.365 $Y2=1.765
r255 38 39 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=4.275 $Y=1.675
+ $X2=4.005 $Y2=1.675
r256 35 92 27.9254 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=3.915 $Y=1.765
+ $X2=3.915 $Y2=1.542
r257 35 37 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.915 $Y=1.765
+ $X2=3.915 $Y2=2.4
r258 31 91 27.9254 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=3.875 $Y=1.32
+ $X2=3.875 $Y2=1.542
r259 31 33 269.202 $w=1.5e-07 $l=5.25e-07 $layer=POLY_cond $X=3.875 $Y=1.32
+ $X2=3.875 $Y2=0.795
r260 28 89 27.9254 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=3.465 $Y=1.765
+ $X2=3.465 $Y2=1.542
r261 28 30 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.465 $Y=1.765
+ $X2=3.465 $Y2=2.4
r262 24 88 27.9254 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=3.445 $Y=1.32
+ $X2=3.445 $Y2=1.542
r263 24 26 269.202 $w=1.5e-07 $l=5.25e-07 $layer=POLY_cond $X=3.445 $Y=1.32
+ $X2=3.445 $Y2=0.795
r264 21 87 27.9254 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=3.015 $Y=1.765
+ $X2=3.015 $Y2=1.542
r265 21 23 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.015 $Y=1.765
+ $X2=3.015 $Y2=2.4
r266 17 86 27.9254 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=2.97 $Y=1.32
+ $X2=2.97 $Y2=1.542
r267 17 19 276.894 $w=1.5e-07 $l=5.4e-07 $layer=POLY_cond $X=2.97 $Y=1.32
+ $X2=2.97 $Y2=0.78
r268 13 84 27.9254 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=2.54 $Y=1.32
+ $X2=2.54 $Y2=1.542
r269 13 15 276.894 $w=1.5e-07 $l=5.4e-07 $layer=POLY_cond $X=2.54 $Y=1.32
+ $X2=2.54 $Y2=0.78
r270 4 69 600 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=0.77
+ $Y=1.96 $X2=0.92 $Y2=2.105
r271 3 82 182 $w=1.7e-07 $l=5.80797e-07 $layer=licon1_NDIFF $count=1 $X=5.88
+ $Y=0.585 $X2=6.02 $Y2=1.1
r272 2 53 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.71
+ $Y=0.41 $X2=1.85 $Y2=0.555
r273 1 45 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=0.85
+ $Y=0.41 $X2=0.99 $Y2=0.555
.ends

.subckt PM_SKY130_FD_SC_HS__A311O_4%A3 1 3 4 5 6 8 9 11 12 14 15 20 21
c65 21 0 8.68168e-20 $X=5.13 $Y=1.585
r66 20 22 22.9524 $w=4.2e-07 $l=2e-07 $layer=POLY_cond $X=5.13 $Y=1.562 $X2=5.33
+ $Y2=1.562
r67 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.13
+ $Y=1.585 $X2=5.13 $Y2=1.585
r68 18 20 28.6905 $w=4.2e-07 $l=2.5e-07 $layer=POLY_cond $X=4.88 $Y=1.562
+ $X2=5.13 $Y2=1.562
r69 17 18 9.75476 $w=4.2e-07 $l=8.5e-08 $layer=POLY_cond $X=4.795 $Y=1.562
+ $X2=4.88 $Y2=1.562
r70 15 21 2.88111 $w=3.58e-07 $l=9e-08 $layer=LI1_cond $X=5.04 $Y=1.6 $X2=5.13
+ $Y2=1.6
r71 12 22 27.059 $w=1.5e-07 $l=3.23e-07 $layer=POLY_cond $X=5.33 $Y=1.885
+ $X2=5.33 $Y2=1.562
r72 12 14 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=5.33 $Y=1.885
+ $X2=5.33 $Y2=2.46
r73 9 18 27.059 $w=1.5e-07 $l=3.23e-07 $layer=POLY_cond $X=4.88 $Y=1.885
+ $X2=4.88 $Y2=1.562
r74 9 11 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=4.88 $Y=1.885
+ $X2=4.88 $Y2=2.46
r75 6 17 27.059 $w=1.5e-07 $l=3.22e-07 $layer=POLY_cond $X=4.795 $Y=1.24
+ $X2=4.795 $Y2=1.562
r76 6 8 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=4.795 $Y=1.24
+ $X2=4.795 $Y2=0.845
r77 4 17 29.6695 $w=4.2e-07 $l=2.82018e-07 $layer=POLY_cond $X=4.72 $Y=1.315
+ $X2=4.795 $Y2=1.562
r78 4 5 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=4.72 $Y=1.315 $X2=4.44
+ $Y2=1.315
r79 1 5 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.365 $Y=1.24
+ $X2=4.44 $Y2=1.315
r80 1 3 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=4.365 $Y=1.24
+ $X2=4.365 $Y2=0.845
.ends

.subckt PM_SKY130_FD_SC_HS__A311O_4%A1 1 3 6 8 10 13 15 16 17 24
c57 8 0 5.4224e-20 $X=6.23 $Y=1.885
c58 6 0 8.35615e-20 $X=5.805 $Y=0.905
c59 1 0 9.08767e-20 $X=5.78 $Y=1.885
r60 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.245
+ $Y=1.615 $X2=6.245 $Y2=1.615
r61 24 26 1.26178 $w=3.82e-07 $l=1e-08 $layer=POLY_cond $X=6.235 $Y=1.667
+ $X2=6.245 $Y2=1.667
r62 23 24 0.63089 $w=3.82e-07 $l=5e-09 $layer=POLY_cond $X=6.23 $Y=1.667
+ $X2=6.235 $Y2=1.667
r63 22 23 53.6257 $w=3.82e-07 $l=4.25e-07 $layer=POLY_cond $X=5.805 $Y=1.667
+ $X2=6.23 $Y2=1.667
r64 21 22 3.15445 $w=3.82e-07 $l=2.5e-08 $layer=POLY_cond $X=5.78 $Y=1.667
+ $X2=5.805 $Y2=1.667
r65 16 17 16.7628 $w=3.28e-07 $l=4.8e-07 $layer=LI1_cond $X=6.48 $Y=1.615
+ $X2=6.96 $Y2=1.615
r66 16 27 8.20679 $w=3.28e-07 $l=2.35e-07 $layer=LI1_cond $X=6.48 $Y=1.615
+ $X2=6.245 $Y2=1.615
r67 15 27 8.55602 $w=3.28e-07 $l=2.45e-07 $layer=LI1_cond $X=6 $Y=1.615
+ $X2=6.245 $Y2=1.615
r68 11 24 24.74 $w=1.5e-07 $l=2.17e-07 $layer=POLY_cond $X=6.235 $Y=1.45
+ $X2=6.235 $Y2=1.667
r69 11 13 279.457 $w=1.5e-07 $l=5.45e-07 $layer=POLY_cond $X=6.235 $Y=1.45
+ $X2=6.235 $Y2=0.905
r70 8 23 24.74 $w=1.5e-07 $l=2.18e-07 $layer=POLY_cond $X=6.23 $Y=1.885 $X2=6.23
+ $Y2=1.667
r71 8 10 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=6.23 $Y=1.885
+ $X2=6.23 $Y2=2.46
r72 4 22 24.74 $w=1.5e-07 $l=2.17e-07 $layer=POLY_cond $X=5.805 $Y=1.45
+ $X2=5.805 $Y2=1.667
r73 4 6 279.457 $w=1.5e-07 $l=5.45e-07 $layer=POLY_cond $X=5.805 $Y=1.45
+ $X2=5.805 $Y2=0.905
r74 1 21 24.74 $w=1.5e-07 $l=2.18e-07 $layer=POLY_cond $X=5.78 $Y=1.885 $X2=5.78
+ $Y2=1.667
r75 1 3 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=5.78 $Y=1.885
+ $X2=5.78 $Y2=2.46
.ends

.subckt PM_SKY130_FD_SC_HS__A311O_4%A2 1 3 6 10 12 14 15 20
r41 20 22 33.1044 $w=3.64e-07 $l=2.5e-07 $layer=POLY_cond $X=7.16 $Y=1.667
+ $X2=7.41 $Y2=1.667
r42 19 20 0.662088 $w=3.64e-07 $l=5e-09 $layer=POLY_cond $X=7.155 $Y=1.667
+ $X2=7.16 $Y2=1.667
r43 18 19 56.9396 $w=3.64e-07 $l=4.3e-07 $layer=POLY_cond $X=6.725 $Y=1.667
+ $X2=7.155 $Y2=1.667
r44 17 18 1.98626 $w=3.64e-07 $l=1.5e-08 $layer=POLY_cond $X=6.71 $Y=1.667
+ $X2=6.725 $Y2=1.667
r45 15 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.41
+ $Y=1.615 $X2=7.41 $Y2=1.615
r46 12 20 23.572 $w=1.5e-07 $l=2.18e-07 $layer=POLY_cond $X=7.16 $Y=1.885
+ $X2=7.16 $Y2=1.667
r47 12 14 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=7.16 $Y=1.885
+ $X2=7.16 $Y2=2.46
r48 8 19 23.572 $w=1.5e-07 $l=2.17e-07 $layer=POLY_cond $X=7.155 $Y=1.45
+ $X2=7.155 $Y2=1.667
r49 8 10 279.457 $w=1.5e-07 $l=5.45e-07 $layer=POLY_cond $X=7.155 $Y=1.45
+ $X2=7.155 $Y2=0.905
r50 4 18 23.572 $w=1.5e-07 $l=2.17e-07 $layer=POLY_cond $X=6.725 $Y=1.45
+ $X2=6.725 $Y2=1.667
r51 4 6 279.457 $w=1.5e-07 $l=5.45e-07 $layer=POLY_cond $X=6.725 $Y=1.45
+ $X2=6.725 $Y2=0.905
r52 1 17 23.572 $w=1.5e-07 $l=2.18e-07 $layer=POLY_cond $X=6.71 $Y=1.885
+ $X2=6.71 $Y2=1.667
r53 1 3 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=6.71 $Y=1.885
+ $X2=6.71 $Y2=2.46
.ends

.subckt PM_SKY130_FD_SC_HS__A311O_4%A_69_392# 1 2 3 14 18 19 21
r38 21 23 7.33373 $w=3.28e-07 $l=2.1e-07 $layer=LI1_cond $X=2.27 $Y=2.78
+ $X2=2.27 $Y2=2.99
r39 17 19 8.55446 $w=3.73e-07 $l=1.65e-07 $layer=LI1_cond $X=1.37 $Y=2.887
+ $X2=1.535 $Y2=2.887
r40 17 18 5.8355 $w=3.73e-07 $l=1.65e-07 $layer=LI1_cond $X=1.37 $Y=2.887
+ $X2=1.205 $Y2=2.887
r41 14 23 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.105 $Y=2.99
+ $X2=2.27 $Y2=2.99
r42 14 19 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=2.105 $Y=2.99
+ $X2=1.535 $Y2=2.99
r43 12 18 30.2516 $w=2.78e-07 $l=7.35e-07 $layer=LI1_cond $X=0.47 $Y=2.84
+ $X2=1.205 $Y2=2.84
r44 3 21 600 $w=1.7e-07 $l=8.91852e-07 $layer=licon1_PDIFF $count=1 $X=2.12
+ $Y=1.96 $X2=2.27 $Y2=2.78
r45 2 17 600 $w=1.7e-07 $l=9.11921e-07 $layer=licon1_PDIFF $count=1 $X=1.22
+ $Y=1.96 $X2=1.37 $Y2=2.8
r46 1 12 600 $w=1.7e-07 $l=9.00333e-07 $layer=licon1_PDIFF $count=1 $X=0.345
+ $Y=1.96 $X2=0.47 $Y2=2.8
.ends

.subckt PM_SKY130_FD_SC_HS__A311O_4%A_334_392# 1 2 3 4 13 17 19 23 25 27 29 31
+ 37 40
c83 37 0 2.28135e-19 $X=5.105 $Y=2.455
r84 31 34 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=1.82 $Y=2.405
+ $X2=1.82 $Y2=2.52
r85 27 42 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.935 $Y=2.12
+ $X2=6.935 $Y2=2.035
r86 27 29 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=6.935 $Y=2.12
+ $X2=6.935 $Y2=2.815
r87 26 39 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.09 $Y=2.035
+ $X2=6.005 $Y2=2.035
r88 25 42 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.85 $Y=2.035
+ $X2=6.935 $Y2=2.035
r89 25 26 49.5829 $w=1.68e-07 $l=7.6e-07 $layer=LI1_cond $X=6.85 $Y=2.035
+ $X2=6.09 $Y2=2.035
r90 21 40 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.005 $Y=2.46
+ $X2=6.005 $Y2=2.375
r91 21 23 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=6.005 $Y=2.46
+ $X2=6.005 $Y2=2.465
r92 20 40 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.005 $Y=2.29
+ $X2=6.005 $Y2=2.375
r93 19 39 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.005 $Y=2.12
+ $X2=6.005 $Y2=2.035
r94 19 20 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=6.005 $Y=2.12
+ $X2=6.005 $Y2=2.29
r95 18 37 8.61065 $w=1.7e-07 $l=1.72337e-07 $layer=LI1_cond $X=5.27 $Y=2.375
+ $X2=5.105 $Y2=2.39
r96 17 40 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.92 $Y=2.375
+ $X2=6.005 $Y2=2.375
r97 17 18 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=5.92 $Y=2.375
+ $X2=5.27 $Y2=2.375
r98 14 31 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.905 $Y=2.405
+ $X2=1.82 $Y2=2.405
r99 13 37 8.61065 $w=1.7e-07 $l=1.72337e-07 $layer=LI1_cond $X=4.94 $Y=2.405
+ $X2=5.105 $Y2=2.39
r100 13 14 198.005 $w=1.68e-07 $l=3.035e-06 $layer=LI1_cond $X=4.94 $Y=2.405
+ $X2=1.905 $Y2=2.405
r101 4 42 400 $w=1.7e-07 $l=2.17428e-07 $layer=licon1_PDIFF $count=1 $X=6.785
+ $Y=1.96 $X2=6.935 $Y2=2.115
r102 4 29 400 $w=1.7e-07 $l=9.26971e-07 $layer=licon1_PDIFF $count=1 $X=6.785
+ $Y=1.96 $X2=6.935 $Y2=2.815
r103 3 39 600 $w=1.7e-07 $l=2.17428e-07 $layer=licon1_PDIFF $count=1 $X=5.855
+ $Y=1.96 $X2=6.005 $Y2=2.115
r104 3 23 300 $w=1.7e-07 $l=5.7513e-07 $layer=licon1_PDIFF $count=2 $X=5.855
+ $Y=1.96 $X2=6.005 $Y2=2.465
r105 2 37 300 $w=1.7e-07 $l=5.65044e-07 $layer=licon1_PDIFF $count=2 $X=4.955
+ $Y=1.96 $X2=5.105 $Y2=2.455
r106 1 34 600 $w=1.7e-07 $l=6.30555e-07 $layer=licon1_PDIFF $count=1 $X=1.67
+ $Y=1.96 $X2=1.82 $Y2=2.52
.ends

.subckt PM_SKY130_FD_SC_HS__A311O_4%VPWR 1 2 3 4 5 6 21 23 27 31 33 37 41 43 45
+ 49 51 56 61 66 72 75 78 81 84 88
r110 87 88 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r111 84 85 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r112 81 82 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r113 79 82 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=5.52 $Y2=3.33
r114 78 79 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r115 75 76 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r116 73 76 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.6 $Y2=3.33
r117 72 73 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r118 70 88 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=7.44 $Y2=3.33
r119 70 85 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=6.48 $Y2=3.33
r120 69 70 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r121 67 84 9.14399 $w=1.7e-07 $l=1.8e-07 $layer=LI1_cond $X=6.65 $Y=3.33
+ $X2=6.47 $Y2=3.33
r122 67 69 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=6.65 $Y=3.33
+ $X2=6.96 $Y2=3.33
r123 66 87 4.70058 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=7.22 $Y=3.33
+ $X2=7.45 $Y2=3.33
r124 66 69 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=7.22 $Y=3.33
+ $X2=6.96 $Y2=3.33
r125 65 85 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=3.33 $X2=6.48
+ $Y2=3.33
r126 65 82 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=3.33 $X2=5.52
+ $Y2=3.33
r127 64 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r128 62 81 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.72 $Y=3.33
+ $X2=5.595 $Y2=3.33
r129 62 64 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=5.72 $Y=3.33 $X2=6
+ $Y2=3.33
r130 61 84 9.14399 $w=1.7e-07 $l=1.8e-07 $layer=LI1_cond $X=6.29 $Y=3.33
+ $X2=6.47 $Y2=3.33
r131 61 64 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=6.29 $Y=3.33 $X2=6
+ $Y2=3.33
r132 60 79 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=4.56 $Y2=3.33
r133 59 60 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r134 57 75 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.855 $Y=3.33
+ $X2=3.69 $Y2=3.33
r135 57 59 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=3.855 $Y=3.33
+ $X2=4.08 $Y2=3.33
r136 56 78 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.425 $Y=3.33
+ $X2=4.59 $Y2=3.33
r137 56 59 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=4.425 $Y=3.33
+ $X2=4.08 $Y2=3.33
r138 54 73 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=2.64 $Y2=3.33
r139 53 54 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r140 51 72 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.625 $Y=3.33
+ $X2=2.79 $Y2=3.33
r141 51 53 155.599 $w=1.68e-07 $l=2.385e-06 $layer=LI1_cond $X=2.625 $Y=3.33
+ $X2=0.24 $Y2=3.33
r142 49 60 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=3.84 $Y=3.33
+ $X2=4.08 $Y2=3.33
r143 49 76 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=3.84 $Y=3.33
+ $X2=3.6 $Y2=3.33
r144 45 48 24.4458 $w=3.28e-07 $l=7e-07 $layer=LI1_cond $X=7.385 $Y=2.115
+ $X2=7.385 $Y2=2.815
r145 43 87 3.0656 $w=3.3e-07 $l=1.12916e-07 $layer=LI1_cond $X=7.385 $Y=3.245
+ $X2=7.45 $Y2=3.33
r146 43 48 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=7.385 $Y=3.245
+ $X2=7.385 $Y2=2.815
r147 39 84 1.16013 $w=3.6e-07 $l=8.5e-08 $layer=LI1_cond $X=6.47 $Y=3.245
+ $X2=6.47 $Y2=3.33
r148 39 41 25.2897 $w=3.58e-07 $l=7.9e-07 $layer=LI1_cond $X=6.47 $Y=3.245
+ $X2=6.47 $Y2=2.455
r149 35 81 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.595 $Y=3.245
+ $X2=5.595 $Y2=3.33
r150 35 37 20.283 $w=2.48e-07 $l=4.4e-07 $layer=LI1_cond $X=5.595 $Y=3.245
+ $X2=5.595 $Y2=2.805
r151 34 78 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.755 $Y=3.33
+ $X2=4.59 $Y2=3.33
r152 33 81 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.47 $Y=3.33
+ $X2=5.595 $Y2=3.33
r153 33 34 46.6471 $w=1.68e-07 $l=7.15e-07 $layer=LI1_cond $X=5.47 $Y=3.33
+ $X2=4.755 $Y2=3.33
r154 29 78 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.59 $Y=3.245
+ $X2=4.59 $Y2=3.33
r155 29 31 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=4.59 $Y=3.245
+ $X2=4.59 $Y2=2.78
r156 25 75 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.69 $Y=3.245
+ $X2=3.69 $Y2=3.33
r157 25 27 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=3.69 $Y=3.245
+ $X2=3.69 $Y2=2.78
r158 24 72 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.955 $Y=3.33
+ $X2=2.79 $Y2=3.33
r159 23 75 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.525 $Y=3.33
+ $X2=3.69 $Y2=3.33
r160 23 24 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=3.525 $Y=3.33
+ $X2=2.955 $Y2=3.33
r161 19 72 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.79 $Y=3.245
+ $X2=2.79 $Y2=3.33
r162 19 21 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=2.79 $Y=3.245
+ $X2=2.79 $Y2=2.78
r163 6 48 400 $w=1.7e-07 $l=9.26971e-07 $layer=licon1_PDIFF $count=1 $X=7.235
+ $Y=1.96 $X2=7.385 $Y2=2.815
r164 6 45 400 $w=1.7e-07 $l=2.17428e-07 $layer=licon1_PDIFF $count=1 $X=7.235
+ $Y=1.96 $X2=7.385 $Y2=2.115
r165 5 41 300 $w=1.7e-07 $l=5.71577e-07 $layer=licon1_PDIFF $count=2 $X=6.305
+ $Y=1.96 $X2=6.47 $Y2=2.455
r166 4 37 600 $w=1.7e-07 $l=9.16938e-07 $layer=licon1_PDIFF $count=1 $X=5.405
+ $Y=1.96 $X2=5.555 $Y2=2.805
r167 3 31 600 $w=1.7e-07 $l=1.01223e-06 $layer=licon1_PDIFF $count=1 $X=4.44
+ $Y=1.84 $X2=4.59 $Y2=2.78
r168 2 27 600 $w=1.7e-07 $l=1.01223e-06 $layer=licon1_PDIFF $count=1 $X=3.54
+ $Y=1.84 $X2=3.69 $Y2=2.78
r169 1 21 600 $w=1.7e-07 $l=1.00055e-06 $layer=licon1_PDIFF $count=1 $X=2.665
+ $Y=1.84 $X2=2.79 $Y2=2.78
.ends

.subckt PM_SKY130_FD_SC_HS__A311O_4%X 1 2 3 4 14 15 16 18 20 21 25 27 28 31 33
+ 35 36 38 41 44 48
c132 44 0 1.88456e-19 $X=2.755 $Y=0.555
r133 48 51 6.56993 $w=2.28e-07 $l=1.15e-07 $layer=LI1_cond $X=0.24 $Y=0.925
+ $X2=0.24 $Y2=1.04
r134 41 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0.925
+ $X2=0.24 $Y2=0.925
r135 39 44 11.0754 $w=3.83e-07 $l=3.7e-07 $layer=LI1_cond $X=2.727 $Y=0.925
+ $X2=2.727 $Y2=0.555
r136 38 39 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0.925
+ $X2=2.64 $Y2=0.925
r137 36 41 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=0.385 $Y=0.925
+ $X2=0.24 $Y2=0.925
r138 35 38 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.495 $Y=0.925
+ $X2=2.64 $Y2=0.925
r139 35 36 2.61138 $w=1.4e-07 $l=2.11e-06 $layer=MET1_cond $X=2.495 $Y=0.925
+ $X2=0.385 $Y2=0.925
r140 34 39 1.64635 $w=3.83e-07 $l=5.5e-08 $layer=LI1_cond $X=2.727 $Y=0.98
+ $X2=2.727 $Y2=0.925
r141 29 31 18.9001 $w=2.48e-07 $l=4.1e-07 $layer=LI1_cond $X=3.62 $Y=0.98
+ $X2=3.62 $Y2=0.57
r142 28 34 8.24022 $w=1.7e-07 $l=2.31633e-07 $layer=LI1_cond $X=2.92 $Y=1.065
+ $X2=2.727 $Y2=0.98
r143 27 29 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=3.495 $Y=1.065
+ $X2=3.62 $Y2=0.98
r144 27 28 37.5134 $w=1.68e-07 $l=5.75e-07 $layer=LI1_cond $X=3.495 $Y=1.065
+ $X2=2.92 $Y2=1.065
r145 23 25 31.4303 $w=3.28e-07 $l=9e-07 $layer=LI1_cond $X=3.24 $Y=1.985
+ $X2=4.14 $Y2=1.985
r146 21 33 8.16218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=2.69 $Y=1.985
+ $X2=2.525 $Y2=1.985
r147 21 23 19.2074 $w=3.28e-07 $l=5.5e-07 $layer=LI1_cond $X=2.69 $Y=1.985
+ $X2=3.24 $Y2=1.985
r148 20 33 66.5455 $w=1.68e-07 $l=1.02e-06 $layer=LI1_cond $X=1.505 $Y=2.055
+ $X2=2.525 $Y2=2.055
r149 17 20 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.42 $Y=2.14
+ $X2=1.505 $Y2=2.055
r150 17 18 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=1.42 $Y=2.14
+ $X2=1.42 $Y2=2.36
r151 15 18 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.335 $Y=2.445
+ $X2=1.42 $Y2=2.36
r152 15 16 67.8503 $w=1.68e-07 $l=1.04e-06 $layer=LI1_cond $X=1.335 $Y=2.445
+ $X2=0.295 $Y2=2.445
r153 14 16 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.21 $Y=2.36
+ $X2=0.295 $Y2=2.445
r154 14 51 86.1176 $w=1.68e-07 $l=1.32e-06 $layer=LI1_cond $X=0.21 $Y=2.36
+ $X2=0.21 $Y2=1.04
r155 4 25 600 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=3.99
+ $Y=1.84 $X2=4.14 $Y2=1.985
r156 3 23 600 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=3.09
+ $Y=1.84 $X2=3.24 $Y2=1.985
r157 2 31 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.52
+ $Y=0.425 $X2=3.66 $Y2=0.57
r158 1 44 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.615
+ $Y=0.41 $X2=2.755 $Y2=0.555
.ends

.subckt PM_SKY130_FD_SC_HS__A311O_4%VGND 1 2 3 4 5 6 21 25 27 31 33 37 42 43 45
+ 48 49 50 51 53 62 72 73 76 79 82
c107 45 0 5.40935e-20 $X=5.01 $Y=1.02
r108 82 83 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r109 79 80 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r110 77 80 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=3.12
+ $Y2=0
r111 76 77 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r112 72 73 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=7.44 $Y=0
+ $X2=7.44 $Y2=0
r113 70 73 0.802756 $w=4.9e-07 $l=2.88e-06 $layer=MET1_cond $X=4.56 $Y=0
+ $X2=7.44 $Y2=0
r114 70 83 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=4.08
+ $Y2=0
r115 69 72 187.893 $w=1.68e-07 $l=2.88e-06 $layer=LI1_cond $X=4.56 $Y=0 $X2=7.44
+ $Y2=0
r116 69 70 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=4.56 $Y=0
+ $X2=4.56 $Y2=0
r117 67 82 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.175 $Y=0 $X2=4.05
+ $Y2=0
r118 67 69 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=4.175 $Y=0
+ $X2=4.56 $Y2=0
r119 66 80 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=3.12
+ $Y2=0
r120 65 66 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r121 63 79 6.25164 $w=1.7e-07 $l=1.08e-07 $layer=LI1_cond $X=3.315 $Y=0
+ $X2=3.207 $Y2=0
r122 63 65 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=3.315 $Y=0 $X2=3.6
+ $Y2=0
r123 62 82 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.925 $Y=0 $X2=4.05
+ $Y2=0
r124 62 65 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=3.925 $Y=0 $X2=3.6
+ $Y2=0
r125 61 77 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r126 60 61 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r127 57 61 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=1.2
+ $Y2=0
r128 56 57 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r129 53 83 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=3.84 $Y=0
+ $X2=4.08 $Y2=0
r130 53 66 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=3.84 $Y=0 $X2=3.6
+ $Y2=0
r131 50 60 3.58824 $w=1.68e-07 $l=5.5e-08 $layer=LI1_cond $X=1.255 $Y=0 $X2=1.2
+ $Y2=0
r132 50 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.255 $Y=0 $X2=1.42
+ $Y2=0
r133 48 56 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=0.395 $Y=0
+ $X2=0.24 $Y2=0
r134 48 49 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.395 $Y=0 $X2=0.56
+ $Y2=0
r135 47 60 30.9893 $w=1.68e-07 $l=4.75e-07 $layer=LI1_cond $X=0.725 $Y=0 $X2=1.2
+ $Y2=0
r136 47 49 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.725 $Y=0 $X2=0.56
+ $Y2=0
r137 43 52 18.3822 $w=2.5e-07 $l=3.75e-07 $layer=LI1_cond $X=4.425 $Y=1.06
+ $X2=4.05 $Y2=1.06
r138 43 45 26.9672 $w=2.48e-07 $l=5.85e-07 $layer=LI1_cond $X=4.425 $Y=1.06
+ $X2=5.01 $Y2=1.06
r139 40 52 0.255588 $w=2.5e-07 $l=1.25e-07 $layer=LI1_cond $X=4.05 $Y=0.935
+ $X2=4.05 $Y2=1.06
r140 40 42 16.8257 $w=2.48e-07 $l=3.65e-07 $layer=LI1_cond $X=4.05 $Y=0.935
+ $X2=4.05 $Y2=0.57
r141 39 82 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.05 $Y=0.085
+ $X2=4.05 $Y2=0
r142 39 42 22.3574 $w=2.48e-07 $l=4.85e-07 $layer=LI1_cond $X=4.05 $Y=0.085
+ $X2=4.05 $Y2=0.57
r143 35 79 0.512231 $w=2.15e-07 $l=8.5e-08 $layer=LI1_cond $X=3.207 $Y=0.085
+ $X2=3.207 $Y2=0
r144 35 37 27.873 $w=2.13e-07 $l=5.2e-07 $layer=LI1_cond $X=3.207 $Y=0.085
+ $X2=3.207 $Y2=0.605
r145 34 76 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.365 $Y=0 $X2=2.24
+ $Y2=0
r146 33 79 6.25164 $w=1.7e-07 $l=1.07e-07 $layer=LI1_cond $X=3.1 $Y=0 $X2=3.207
+ $Y2=0
r147 33 34 47.9519 $w=1.68e-07 $l=7.35e-07 $layer=LI1_cond $X=3.1 $Y=0 $X2=2.365
+ $Y2=0
r148 29 76 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.24 $Y=0.085
+ $X2=2.24 $Y2=0
r149 29 31 32.7294 $w=2.48e-07 $l=7.1e-07 $layer=LI1_cond $X=2.24 $Y=0.085
+ $X2=2.24 $Y2=0.795
r150 28 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.585 $Y=0 $X2=1.42
+ $Y2=0
r151 27 76 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.115 $Y=0 $X2=2.24
+ $Y2=0
r152 27 28 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=2.115 $Y=0
+ $X2=1.585 $Y2=0
r153 23 51 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.42 $Y=0.085
+ $X2=1.42 $Y2=0
r154 23 25 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=1.42 $Y=0.085
+ $X2=1.42 $Y2=0.535
r155 19 49 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.56 $Y=0.085
+ $X2=0.56 $Y2=0
r156 19 21 16.4136 $w=3.28e-07 $l=4.7e-07 $layer=LI1_cond $X=0.56 $Y=0.085
+ $X2=0.56 $Y2=0.555
r157 6 45 182 $w=1.7e-07 $l=5.60647e-07 $layer=licon1_NDIFF $count=1 $X=4.87
+ $Y=0.525 $X2=5.01 $Y2=1.02
r158 5 42 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.95
+ $Y=0.425 $X2=4.09 $Y2=0.57
r159 4 37 182 $w=1.7e-07 $l=2.63106e-07 $layer=licon1_NDIFF $count=1 $X=3.045
+ $Y=0.41 $X2=3.205 $Y2=0.605
r160 3 31 182 $w=1.7e-07 $l=4.49583e-07 $layer=licon1_NDIFF $count=1 $X=2.14
+ $Y=0.41 $X2=2.28 $Y2=0.795
r161 2 25 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=1.28
+ $Y=0.41 $X2=1.42 $Y2=0.535
r162 1 21 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=0.435
+ $Y=0.41 $X2=0.56 $Y2=0.555
.ends

.subckt PM_SKY130_FD_SC_HS__A311O_4%A_888_105# 1 2 12 14 15
r30 14 15 9.26861 $w=2.18e-07 $l=1.65e-07 $layer=LI1_cond $X=6.94 $Y=0.705
+ $X2=6.775 $Y2=0.705
r31 12 15 132.439 $w=1.68e-07 $l=2.03e-06 $layer=LI1_cond $X=4.745 $Y=0.68
+ $X2=6.775 $Y2=0.68
r32 10 12 8.69362 $w=2.58e-07 $l=1.65e-07 $layer=LI1_cond $X=4.58 $Y=0.635
+ $X2=4.745 $Y2=0.635
r33 2 14 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=6.8
+ $Y=0.585 $X2=6.94 $Y2=0.73
r34 1 10 182 $w=1.7e-07 $l=2.08567e-07 $layer=licon1_NDIFF $count=1 $X=4.44
+ $Y=0.525 $X2=4.58 $Y2=0.675
.ends

.subckt PM_SKY130_FD_SC_HS__A311O_4%A_1081_39# 1 2 3 10 14 19 21
c30 14 0 8.35615e-20 $X=7.285 $Y=1.115
r31 19 23 3.47681 $w=2.5e-07 $l=1.3e-07 $layer=LI1_cond $X=7.41 $Y=0.985
+ $X2=7.41 $Y2=1.115
r32 19 21 11.7549 $w=2.48e-07 $l=2.55e-07 $layer=LI1_cond $X=7.41 $Y=0.985
+ $X2=7.41 $Y2=0.73
r33 18 21 14.0598 $w=2.48e-07 $l=3.05e-07 $layer=LI1_cond $X=7.41 $Y=0.425
+ $X2=7.41 $Y2=0.73
r34 14 23 3.34309 $w=2.6e-07 $l=1.25e-07 $layer=LI1_cond $X=7.285 $Y=1.115
+ $X2=7.41 $Y2=1.115
r35 14 16 37.0112 $w=2.58e-07 $l=8.35e-07 $layer=LI1_cond $X=7.285 $Y=1.115
+ $X2=6.45 $Y2=1.115
r36 10 18 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=7.285 $Y=0.34
+ $X2=7.41 $Y2=0.425
r37 10 12 114.497 $w=1.68e-07 $l=1.755e-06 $layer=LI1_cond $X=7.285 $Y=0.34
+ $X2=5.53 $Y2=0.34
r38 3 23 182 $w=1.7e-07 $l=5.60647e-07 $layer=licon1_NDIFF $count=1 $X=7.23
+ $Y=0.585 $X2=7.37 $Y2=1.08
r39 3 21 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=7.23
+ $Y=0.585 $X2=7.37 $Y2=0.73
r40 2 16 182 $w=1.7e-07 $l=5.55608e-07 $layer=licon1_NDIFF $count=1 $X=6.31
+ $Y=0.585 $X2=6.45 $Y2=1.075
r41 1 12 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=5.405
+ $Y=0.195 $X2=5.53 $Y2=0.34
.ends

