# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_hs__fah_4
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_hs__fah_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  15.36000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425000 1.510000 1.095000 1.800000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.723000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.675000 1.220000 4.925000 2.290000 ;
        RECT 4.675000 2.290000 5.155000 2.910000 ;
    END
  END B
  PIN CI
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 12.635000 1.350000 12.980000 1.780000 ;
    END
  END CI
  PIN COUT
    ANTENNADIFFAREA  1.086400 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT  9.890000 1.850000 11.395000 2.100000 ;
        RECT 10.475000 1.010000 11.785000 1.180000 ;
        RECT 10.960000 1.180000 11.785000 1.260000 ;
        RECT 10.960000 1.260000 11.395000 1.850000 ;
    END
  END COUT
  PIN SUM
    ANTENNADIFFAREA  1.097600 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 13.420000 1.850000 14.755000 2.020000 ;
        RECT 13.420000 2.020000 13.750000 2.980000 ;
        RECT 13.555000 0.480000 13.805000 1.010000 ;
        RECT 13.555000 1.010000 14.745000 1.180000 ;
        RECT 14.420000 2.020000 14.755000 2.980000 ;
        RECT 14.495000 0.480000 14.745000 1.010000 ;
        RECT 14.495000 1.180000 14.745000 1.850000 ;
    END
  END SUM
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT  0.000000 -0.085000 15.360000 0.085000 ;
        RECT  0.545000  0.085000  0.795000 1.000000 ;
        RECT  1.535000  0.085000  1.795000 0.620000 ;
        RECT  4.585000  0.085000  4.915000 0.535000 ;
        RECT 10.065000  0.085000 10.315000 0.500000 ;
        RECT 10.965000  0.085000 11.295000 0.500000 ;
        RECT 11.965000  0.085000 12.295000 0.500000 ;
        RECT 13.035000  0.085000 13.375000 0.500000 ;
        RECT 13.985000  0.085000 14.315000 0.840000 ;
        RECT 14.915000  0.085000 15.245000 1.260000 ;
      LAYER mcon ;
        RECT  0.155000 -0.085000  0.325000 0.085000 ;
        RECT  0.635000 -0.085000  0.805000 0.085000 ;
        RECT  1.115000 -0.085000  1.285000 0.085000 ;
        RECT  1.595000 -0.085000  1.765000 0.085000 ;
        RECT  2.075000 -0.085000  2.245000 0.085000 ;
        RECT  2.555000 -0.085000  2.725000 0.085000 ;
        RECT  3.035000 -0.085000  3.205000 0.085000 ;
        RECT  3.515000 -0.085000  3.685000 0.085000 ;
        RECT  3.995000 -0.085000  4.165000 0.085000 ;
        RECT  4.475000 -0.085000  4.645000 0.085000 ;
        RECT  4.955000 -0.085000  5.125000 0.085000 ;
        RECT  5.435000 -0.085000  5.605000 0.085000 ;
        RECT  5.915000 -0.085000  6.085000 0.085000 ;
        RECT  6.395000 -0.085000  6.565000 0.085000 ;
        RECT  6.875000 -0.085000  7.045000 0.085000 ;
        RECT  7.355000 -0.085000  7.525000 0.085000 ;
        RECT  7.835000 -0.085000  8.005000 0.085000 ;
        RECT  8.315000 -0.085000  8.485000 0.085000 ;
        RECT  8.795000 -0.085000  8.965000 0.085000 ;
        RECT  9.275000 -0.085000  9.445000 0.085000 ;
        RECT  9.755000 -0.085000  9.925000 0.085000 ;
        RECT 10.235000 -0.085000 10.405000 0.085000 ;
        RECT 10.715000 -0.085000 10.885000 0.085000 ;
        RECT 11.195000 -0.085000 11.365000 0.085000 ;
        RECT 11.675000 -0.085000 11.845000 0.085000 ;
        RECT 12.155000 -0.085000 12.325000 0.085000 ;
        RECT 12.635000 -0.085000 12.805000 0.085000 ;
        RECT 13.115000 -0.085000 13.285000 0.085000 ;
        RECT 13.595000 -0.085000 13.765000 0.085000 ;
        RECT 14.075000 -0.085000 14.245000 0.085000 ;
        RECT 14.555000 -0.085000 14.725000 0.085000 ;
        RECT 15.035000 -0.085000 15.205000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.245000 15.360000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT  0.000000 3.245000 15.360000 3.415000 ;
        RECT  0.565000 1.970000  0.815000 3.245000 ;
        RECT  1.575000 2.970000  1.915000 3.245000 ;
        RECT  5.325000 2.290000  5.655000 3.245000 ;
        RECT  9.115000 2.950000  9.685000 3.245000 ;
        RECT 10.425000 2.950000 10.755000 3.245000 ;
        RECT 11.495000 2.950000 12.125000 3.245000 ;
        RECT 12.920000 1.950000 13.250000 3.245000 ;
        RECT 13.920000 2.190000 14.250000 3.245000 ;
        RECT 14.950000 1.820000 15.200000 3.245000 ;
      LAYER mcon ;
        RECT  0.155000 3.245000  0.325000 3.415000 ;
        RECT  0.635000 3.245000  0.805000 3.415000 ;
        RECT  1.115000 3.245000  1.285000 3.415000 ;
        RECT  1.595000 3.245000  1.765000 3.415000 ;
        RECT  2.075000 3.245000  2.245000 3.415000 ;
        RECT  2.555000 3.245000  2.725000 3.415000 ;
        RECT  3.035000 3.245000  3.205000 3.415000 ;
        RECT  3.515000 3.245000  3.685000 3.415000 ;
        RECT  3.995000 3.245000  4.165000 3.415000 ;
        RECT  4.475000 3.245000  4.645000 3.415000 ;
        RECT  4.955000 3.245000  5.125000 3.415000 ;
        RECT  5.435000 3.245000  5.605000 3.415000 ;
        RECT  5.915000 3.245000  6.085000 3.415000 ;
        RECT  6.395000 3.245000  6.565000 3.415000 ;
        RECT  6.875000 3.245000  7.045000 3.415000 ;
        RECT  7.355000 3.245000  7.525000 3.415000 ;
        RECT  7.835000 3.245000  8.005000 3.415000 ;
        RECT  8.315000 3.245000  8.485000 3.415000 ;
        RECT  8.795000 3.245000  8.965000 3.415000 ;
        RECT  9.275000 3.245000  9.445000 3.415000 ;
        RECT  9.755000 3.245000  9.925000 3.415000 ;
        RECT 10.235000 3.245000 10.405000 3.415000 ;
        RECT 10.715000 3.245000 10.885000 3.415000 ;
        RECT 11.195000 3.245000 11.365000 3.415000 ;
        RECT 11.675000 3.245000 11.845000 3.415000 ;
        RECT 12.155000 3.245000 12.325000 3.415000 ;
        RECT 12.635000 3.245000 12.805000 3.415000 ;
        RECT 13.115000 3.245000 13.285000 3.415000 ;
        RECT 13.595000 3.245000 13.765000 3.415000 ;
        RECT 14.075000 3.245000 14.245000 3.415000 ;
        RECT 14.555000 3.245000 14.725000 3.415000 ;
        RECT 15.035000 3.245000 15.205000 3.415000 ;
      LAYER met1 ;
        RECT 0.000000 3.085000 15.360000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.085000 0.350000  0.365000 1.170000 ;
      RECT  0.085000 1.170000  1.665000 1.340000 ;
      RECT  0.085000 1.340000  0.255000 1.970000 ;
      RECT  0.085000 1.970000  0.365000 2.980000 ;
      RECT  0.975000 0.350000  1.305000 0.790000 ;
      RECT  0.975000 0.790000  2.135000 0.960000 ;
      RECT  0.975000 0.960000  2.005000 1.000000 ;
      RECT  1.015000 1.970000  1.345000 2.630000 ;
      RECT  1.015000 2.630000  3.495000 2.800000 ;
      RECT  1.015000 2.800000  1.345000 2.980000 ;
      RECT  1.335000 1.340000  1.665000 1.650000 ;
      RECT  1.835000 1.000000  2.005000 2.630000 ;
      RECT  1.965000 0.255000  3.415000 0.425000 ;
      RECT  1.965000 0.425000  2.135000 0.790000 ;
      RECT  2.175000 1.790000  2.505000 2.290000 ;
      RECT  2.175000 2.290000  4.505000 2.460000 ;
      RECT  2.305000 0.625000  2.475000 1.790000 ;
      RECT  2.655000 0.625000  2.985000 1.210000 ;
      RECT  2.655000 1.210000  3.545000 1.380000 ;
      RECT  2.705000 1.550000  3.205000 1.780000 ;
      RECT  2.705000 1.780000  2.960000 2.120000 ;
      RECT  3.155000 0.425000  3.415000 1.040000 ;
      RECT  3.165000 2.800000  3.495000 2.960000 ;
      RECT  3.375000 1.380000  3.545000 1.935000 ;
      RECT  3.375000 1.935000  4.030000 2.120000 ;
      RECT  3.715000 0.630000  3.885000 1.550000 ;
      RECT  3.715000 1.550000  4.165000 1.765000 ;
      RECT  4.055000 0.255000  4.385000 0.705000 ;
      RECT  4.055000 0.705000  5.405000 0.875000 ;
      RECT  4.065000 1.045000  4.505000 1.310000 ;
      RECT  4.230000 1.935000  4.505000 2.290000 ;
      RECT  4.230000 2.460000  4.505000 2.670000 ;
      RECT  4.335000 1.310000  4.505000 1.935000 ;
      RECT  5.095000 0.255000  8.195000 0.425000 ;
      RECT  5.095000 0.425000  5.405000 0.705000 ;
      RECT  5.095000 0.875000  5.405000 0.920000 ;
      RECT  5.095000 0.920000  5.265000 1.950000 ;
      RECT  5.095000 1.950000  6.025000 2.120000 ;
      RECT  5.435000 1.090000  5.805000 1.375000 ;
      RECT  5.435000 1.375000  5.635000 1.780000 ;
      RECT  5.855000 2.120000  6.025000 2.980000 ;
      RECT  5.875000 0.595000  6.205000 0.875000 ;
      RECT  5.885000 1.550000  6.145000 1.780000 ;
      RECT  5.975000 0.875000  6.145000 1.550000 ;
      RECT  6.195000 1.980000  6.485000 2.150000 ;
      RECT  6.195000 2.150000  6.365000 2.905000 ;
      RECT  6.195000 2.905000  8.715000 3.075000 ;
      RECT  6.315000 1.045000  7.195000 1.215000 ;
      RECT  6.315000 1.215000  6.485000 1.980000 ;
      RECT  6.375000 0.595000  8.535000 0.765000 ;
      RECT  6.375000 0.765000  6.705000 0.845000 ;
      RECT  6.535000 2.320000  7.535000 2.490000 ;
      RECT  6.535000 2.490000  6.785000 2.735000 ;
      RECT  6.655000 1.405000  7.075000 2.150000 ;
      RECT  6.865000 1.015000  7.195000 1.045000 ;
      RECT  6.990000 2.725000  7.875000 2.905000 ;
      RECT  7.365000 0.935000  8.875000 1.105000 ;
      RECT  7.365000 1.105000  7.685000 1.285000 ;
      RECT  7.365000 1.285000  7.535000 2.320000 ;
      RECT  7.705000 1.480000  8.875000 1.650000 ;
      RECT  7.705000 1.650000  7.875000 2.725000 ;
      RECT  8.045000 2.095000  8.375000 2.270000 ;
      RECT  8.045000 2.270000 12.125000 2.440000 ;
      RECT  8.045000 2.440000  8.375000 2.735000 ;
      RECT  8.205000 1.320000  8.875000 1.480000 ;
      RECT  8.365000 0.255000  9.895000 0.425000 ;
      RECT  8.365000 0.425000  8.535000 0.595000 ;
      RECT  8.545000 2.610000 12.715000 2.780000 ;
      RECT  8.545000 2.780000  8.715000 2.905000 ;
      RECT  8.580000 1.900000  9.215000 2.100000 ;
      RECT  8.705000 0.595000  9.555000 0.765000 ;
      RECT  8.705000 0.765000  8.875000 0.935000 ;
      RECT  9.045000 0.935000  9.215000 1.550000 ;
      RECT  9.045000 1.550000  9.475000 1.775000 ;
      RECT  9.045000 1.775000  9.215000 1.900000 ;
      RECT  9.385000 0.765000  9.555000 1.010000 ;
      RECT  9.385000 1.010000  9.950000 1.180000 ;
      RECT  9.725000 0.425000  9.895000 0.670000 ;
      RECT  9.725000 0.670000 13.385000 0.840000 ;
      RECT  9.780000 1.180000  9.950000 1.350000 ;
      RECT  9.780000 1.350000 10.710000 1.680000 ;
      RECT 11.955000 0.840000 12.125000 2.270000 ;
      RECT 12.295000 1.010000 12.855000 1.180000 ;
      RECT 12.295000 1.180000 12.465000 1.950000 ;
      RECT 12.295000 1.950000 12.715000 2.610000 ;
      RECT 12.295000 2.780000 12.715000 2.860000 ;
      RECT 13.215000 0.840000 13.385000 1.350000 ;
      RECT 13.215000 1.350000 14.325000 1.680000 ;
    LAYER mcon ;
      RECT 3.035000 1.580000 3.205000 1.750000 ;
      RECT 3.515000 1.950000 3.685000 2.120000 ;
      RECT 3.995000 1.580000 4.165000 1.750000 ;
      RECT 5.435000 1.580000 5.605000 1.750000 ;
      RECT 5.915000 1.580000 6.085000 1.750000 ;
      RECT 6.875000 1.950000 7.045000 2.120000 ;
      RECT 9.275000 1.580000 9.445000 1.750000 ;
    LAYER met1 ;
      RECT 2.975000 1.550000 3.265000 1.595000 ;
      RECT 2.975000 1.595000 5.665000 1.735000 ;
      RECT 2.975000 1.735000 3.265000 1.780000 ;
      RECT 3.455000 1.920000 3.745000 1.965000 ;
      RECT 3.455000 1.965000 7.105000 2.105000 ;
      RECT 3.455000 2.105000 3.745000 2.150000 ;
      RECT 3.935000 1.550000 4.225000 1.595000 ;
      RECT 3.935000 1.735000 4.225000 1.780000 ;
      RECT 5.375000 1.550000 5.665000 1.595000 ;
      RECT 5.375000 1.735000 5.665000 1.780000 ;
      RECT 5.855000 1.550000 6.145000 1.595000 ;
      RECT 5.855000 1.595000 9.505000 1.735000 ;
      RECT 5.855000 1.735000 6.145000 1.780000 ;
      RECT 6.815000 1.920000 7.105000 1.965000 ;
      RECT 6.815000 2.105000 7.105000 2.150000 ;
      RECT 9.215000 1.550000 9.505000 1.595000 ;
      RECT 9.215000 1.735000 9.505000 1.780000 ;
  END
END sky130_fd_sc_hs__fah_4
