* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hs__o22a_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
X0 VPWR a_82_48# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X1 X a_82_48# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X2 X a_82_48# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X3 a_82_48# A2 a_575_384# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=150000u
X4 VGND a_82_48# X VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X5 a_383_384# B2 a_82_48# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=150000u
X6 a_575_384# A1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=150000u
X7 a_307_74# B1 a_82_48# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X8 VGND A1 a_307_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X9 a_307_74# A2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X10 VPWR B1 a_383_384# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=150000u
X11 a_82_48# B2 a_307_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
.ends
