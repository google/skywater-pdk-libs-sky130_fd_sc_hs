* File: sky130_fd_sc_hs__dfbbn_2.pex.spice
* Created: Tue Sep  1 19:59:27 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HS__DFBBN_2%CLK_N 3 5 7 8 12
c31 5 0 1.54296e-19 $X=0.495 $Y=1.765
r32 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.33
+ $Y=1.465 $X2=0.33 $Y2=1.465
r33 8 12 6.22942 $w=3.68e-07 $l=2e-07 $layer=LI1_cond $X=0.31 $Y=1.665 $X2=0.31
+ $Y2=1.465
r34 5 11 57.3754 $w=3.5e-07 $l=3.54965e-07 $layer=POLY_cond $X=0.495 $Y=1.765
+ $X2=0.375 $Y2=1.465
r35 5 7 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.495 $Y=1.765
+ $X2=0.495 $Y2=2.4
r36 1 11 38.7839 $w=3.5e-07 $l=2.16852e-07 $layer=POLY_cond $X=0.495 $Y=1.3
+ $X2=0.375 $Y2=1.465
r37 1 3 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=0.495 $Y=1.3 $X2=0.495
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HS__DFBBN_2%D 3 6 7 9 10 11 18
r43 16 18 19.2347 $w=3.3e-07 $l=1.1e-07 $layer=POLY_cond $X=2.01 $Y=1.345
+ $X2=2.12 $Y2=1.345
r44 14 16 16.6118 $w=3.3e-07 $l=9.5e-08 $layer=POLY_cond $X=1.915 $Y=1.345
+ $X2=2.01 $Y2=1.345
r45 10 11 18.1597 $w=3.28e-07 $l=5.2e-07 $layer=LI1_cond $X=2.12 $Y=1.345
+ $X2=2.64 $Y2=1.345
r46 10 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.12
+ $Y=1.345 $X2=2.12 $Y2=1.345
r47 7 9 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=2.01 $Y=2.44 $X2=2.01
+ $Y2=2.725
r48 6 7 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=2.01 $Y=2.35 $X2=2.01
+ $Y2=2.44
r49 5 16 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=2.01 $Y=1.51
+ $X2=2.01 $Y2=1.345
r50 5 6 326.516 $w=1.8e-07 $l=8.4e-07 $layer=POLY_cond $X=2.01 $Y=1.51 $X2=2.01
+ $Y2=2.35
r51 1 14 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.915 $Y=1.18
+ $X2=1.915 $Y2=1.345
r52 1 3 192.287 $w=1.5e-07 $l=3.75e-07 $layer=POLY_cond $X=1.915 $Y=1.18
+ $X2=1.915 $Y2=0.805
.ends

.subckt PM_SKY130_FD_SC_HS__DFBBN_2%A_473_405# 1 2 3 12 14 16 19 21 23 25 26 27
+ 29 31 32 34 36 40 42 43 49 52 54
c177 34 0 1.08905e-19 $X=4.91 $Y=0.86
c178 19 0 1.32682e-19 $X=6.125 $Y=0.9
c179 14 0 1.48509e-19 $X=2.605 $Y=2.44
c180 12 0 4.5553e-21 $X=2.57 $Y=0.805
r181 46 49 6.63528 $w=3.28e-07 $l=1.9e-07 $layer=LI1_cond $X=2.53 $Y=2.19
+ $X2=2.72 $Y2=2.19
r182 46 47 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.53
+ $Y=2.19 $X2=2.53 $Y2=2.19
r183 43 60 36.2507 $w=3.59e-07 $l=2.7e-07 $layer=POLY_cond $X=6.215 $Y=1.837
+ $X2=6.485 $Y2=1.837
r184 43 58 12.0836 $w=3.59e-07 $l=9e-08 $layer=POLY_cond $X=6.215 $Y=1.837
+ $X2=6.125 $Y2=1.837
r185 42 43 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.215
+ $Y=1.795 $X2=6.215 $Y2=1.795
r186 40 54 31.6417 $w=1.68e-07 $l=4.85e-07 $layer=LI1_cond $X=6.215 $Y=2.405
+ $X2=5.73 $Y2=2.405
r187 40 42 18.3343 $w=3.28e-07 $l=5.25e-07 $layer=LI1_cond $X=6.215 $Y=2.32
+ $X2=6.215 $Y2=1.795
r188 37 52 3.3845 $w=1.7e-07 $l=2.98973e-07 $layer=LI1_cond $X=4.775 $Y=2.405
+ $X2=4.48 $Y2=2.397
r189 36 54 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=5.565 $Y=2.405
+ $X2=5.73 $Y2=2.405
r190 36 37 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=5.565 $Y=2.405
+ $X2=4.775 $Y2=2.405
r191 32 34 3.05058 $w=3.38e-07 $l=9e-08 $layer=LI1_cond $X=4.905 $Y=0.95
+ $X2=4.905 $Y2=0.86
r192 31 52 3.19717 $w=2.95e-07 $l=2.51833e-07 $layer=LI1_cond $X=4.69 $Y=2.305
+ $X2=4.48 $Y2=2.397
r193 30 32 13.2776 $w=3.17e-07 $l=4.39545e-07 $layer=LI1_cond $X=4.69 $Y=1.295
+ $X2=4.905 $Y2=0.95
r194 30 31 65.8931 $w=1.68e-07 $l=1.01e-06 $layer=LI1_cond $X=4.69 $Y=1.295
+ $X2=4.69 $Y2=2.305
r195 28 52 3.19717 $w=2.95e-07 $l=1.28662e-07 $layer=LI1_cond $X=4.395 $Y=2.49
+ $X2=4.48 $Y2=2.397
r196 28 29 11.3872 $w=4.18e-07 $l=4.15e-07 $layer=LI1_cond $X=4.395 $Y=2.49
+ $X2=4.395 $Y2=2.905
r197 26 29 8.54503 $w=1.7e-07 $l=2.48898e-07 $layer=LI1_cond $X=4.185 $Y=2.99
+ $X2=4.395 $Y2=2.905
r198 26 27 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=4.185 $Y=2.99
+ $X2=2.805 $Y2=2.99
r199 25 27 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.72 $Y=2.905
+ $X2=2.805 $Y2=2.99
r200 24 49 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.72 $Y=2.355
+ $X2=2.72 $Y2=2.19
r201 24 25 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=2.72 $Y=2.355
+ $X2=2.72 $Y2=2.905
r202 21 60 23.2387 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=6.485 $Y=2.045
+ $X2=6.485 $Y2=1.837
r203 21 23 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=6.485 $Y=2.045
+ $X2=6.485 $Y2=2.54
r204 17 58 23.2387 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=6.125 $Y=1.63
+ $X2=6.125 $Y2=1.837
r205 17 19 374.319 $w=1.5e-07 $l=7.3e-07 $layer=POLY_cond $X=6.125 $Y=1.63
+ $X2=6.125 $Y2=0.9
r206 14 47 52.2586 $w=2.99e-07 $l=2.85044e-07 $layer=POLY_cond $X=2.605 $Y=2.44
+ $X2=2.53 $Y2=2.19
r207 14 16 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=2.605 $Y=2.44
+ $X2=2.605 $Y2=2.725
r208 10 47 38.5562 $w=2.99e-07 $l=1.83916e-07 $layer=POLY_cond $X=2.57 $Y=2.025
+ $X2=2.53 $Y2=2.19
r209 10 12 625.574 $w=1.5e-07 $l=1.22e-06 $layer=POLY_cond $X=2.57 $Y=2.025
+ $X2=2.57 $Y2=0.805
r210 3 54 300 $w=1.7e-07 $l=3.52101e-07 $layer=licon1_PDIFF $count=2 $X=5.58
+ $Y=2.12 $X2=5.73 $Y2=2.405
r211 2 52 300 $w=1.7e-07 $l=3.28634e-07 $layer=licon1_PDIFF $count=2 $X=4.22
+ $Y=2.12 $X2=4.35 $Y2=2.39
r212 1 34 182 $w=1.7e-07 $l=2.96859e-07 $layer=licon1_NDIFF $count=1 $X=4.77
+ $Y=0.625 $X2=4.91 $Y2=0.86
.ends

.subckt PM_SKY130_FD_SC_HS__DFBBN_2%A_200_74# 1 2 7 9 12 13 15 16 18 22 25 29 30
+ 32 33 34 37 41 42 44 47 50 51 52 53 54 58 60 61 67 72 73 74
c228 61 0 4.5553e-21 $X=3.265 $Y=1.295
c229 58 0 1.03189e-19 $X=7.85 $Y=1.385
c230 54 0 1.71006e-19 $X=7.81 $Y=1.295
c231 53 0 4.11442e-20 $X=3.102 $Y=1.77
c232 50 0 1.54296e-19 $X=1.17 $Y=1.985
c233 42 0 1.06658e-19 $X=6.95 $Y=1.41
c234 41 0 9.60143e-20 $X=3.117 $Y=1.685
c235 34 0 1.55193e-19 $X=2.125 $Y=1.77
c236 16 0 1.87607e-19 $X=8.125 $Y=1.22
r237 72 74 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.38 $Y=1.29
+ $X2=3.38 $Y2=1.125
r238 72 73 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.38
+ $Y=1.29 $X2=3.38 $Y2=1.29
r239 67 68 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=1.295
+ $X2=6.96 $Y2=1.295
r240 64 73 9.07985 $w=3.28e-07 $l=2.6e-07 $layer=LI1_cond $X=3.12 $Y=1.29
+ $X2=3.38 $Y2=1.29
r241 64 79 0.104768 $w=3.28e-07 $l=3e-09 $layer=LI1_cond $X=3.12 $Y=1.29
+ $X2=3.117 $Y2=1.29
r242 63 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=1.295
+ $X2=3.12 $Y2=1.295
r243 61 63 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.265 $Y=1.295
+ $X2=3.12 $Y2=1.295
r244 60 67 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.815 $Y=1.295
+ $X2=6.96 $Y2=1.295
r245 60 61 4.39356 $w=1.4e-07 $l=3.55e-06 $layer=MET1_cond $X=6.815 $Y=1.295
+ $X2=3.265 $Y2=1.295
r246 57 58 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.85
+ $Y=1.385 $X2=7.85 $Y2=1.385
r247 54 57 4.14879 $w=2.48e-07 $l=9e-08 $layer=LI1_cond $X=7.81 $Y=1.295
+ $X2=7.81 $Y2=1.385
r248 51 52 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.36 $Y=1.82
+ $X2=1.36 $Y2=1.13
r249 50 51 8.83531 $w=4.38e-07 $l=1.65e-07 $layer=LI1_cond $X=1.225 $Y=1.985
+ $X2=1.225 $Y2=1.82
r250 48 68 4.18573 $w=2.3e-07 $l=1.65e-07 $layer=LI1_cond $X=7.115 $Y=1.295
+ $X2=6.95 $Y2=1.295
r251 47 54 1.2199 $w=2.3e-07 $l=1.25e-07 $layer=LI1_cond $X=7.685 $Y=1.295
+ $X2=7.81 $Y2=1.295
r252 47 48 28.5605 $w=2.28e-07 $l=5.7e-07 $layer=LI1_cond $X=7.685 $Y=1.295
+ $X2=7.115 $Y2=1.295
r253 44 45 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.95
+ $Y=1.745 $X2=6.95 $Y2=1.745
r254 42 68 2.91733 $w=3.3e-07 $l=1.15e-07 $layer=LI1_cond $X=6.95 $Y=1.41
+ $X2=6.95 $Y2=1.295
r255 42 44 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=6.95 $Y=1.41
+ $X2=6.95 $Y2=1.745
r256 41 53 3.84343 $w=2.4e-07 $l=9.21954e-08 $layer=LI1_cond $X=3.117 $Y=1.685
+ $X2=3.102 $Y2=1.77
r257 40 79 2.99809 $w=2.25e-07 $l=1.65e-07 $layer=LI1_cond $X=3.117 $Y=1.455
+ $X2=3.117 $Y2=1.29
r258 40 41 11.7805 $w=2.23e-07 $l=2.3e-07 $layer=LI1_cond $X=3.117 $Y=1.455
+ $X2=3.117 $Y2=1.685
r259 37 38 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.07
+ $Y=2.19 $X2=3.07 $Y2=2.19
r260 35 53 3.84343 $w=2.4e-07 $l=8.5e-08 $layer=LI1_cond $X=3.102 $Y=1.855
+ $X2=3.102 $Y2=1.77
r261 35 37 15.1399 $w=2.53e-07 $l=3.35e-07 $layer=LI1_cond $X=3.102 $Y=1.855
+ $X2=3.102 $Y2=2.19
r262 33 53 2.60907 $w=1.7e-07 $l=1.27e-07 $layer=LI1_cond $X=2.975 $Y=1.77
+ $X2=3.102 $Y2=1.77
r263 33 34 55.4545 $w=1.68e-07 $l=8.5e-07 $layer=LI1_cond $X=2.975 $Y=1.77
+ $X2=2.125 $Y2=1.77
r264 31 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.04 $Y=1.855
+ $X2=2.125 $Y2=1.77
r265 31 32 68.5027 $w=1.68e-07 $l=1.05e-06 $layer=LI1_cond $X=2.04 $Y=1.855
+ $X2=2.04 $Y2=2.905
r266 29 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.955 $Y=2.99
+ $X2=2.04 $Y2=2.905
r267 29 30 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=1.955 $Y=2.99
+ $X2=1.445 $Y2=2.99
r268 23 52 9.49412 $w=3.88e-07 $l=1.95e-07 $layer=LI1_cond $X=1.25 $Y=0.935
+ $X2=1.25 $Y2=1.13
r269 23 25 12.4109 $w=3.88e-07 $l=4.2e-07 $layer=LI1_cond $X=1.25 $Y=0.935
+ $X2=1.25 $Y2=0.515
r270 20 30 8.71846 $w=1.7e-07 $l=2.59037e-07 $layer=LI1_cond $X=1.225 $Y=2.905
+ $X2=1.445 $Y2=2.99
r271 20 22 2.35727 $w=4.38e-07 $l=9e-08 $layer=LI1_cond $X=1.225 $Y=2.905
+ $X2=1.225 $Y2=2.815
r272 19 50 1.44055 $w=4.38e-07 $l=5.5e-08 $layer=LI1_cond $X=1.225 $Y=2.04
+ $X2=1.225 $Y2=1.985
r273 19 22 20.2987 $w=4.38e-07 $l=7.75e-07 $layer=LI1_cond $X=1.225 $Y=2.04
+ $X2=1.225 $Y2=2.815
r274 16 58 50.0189 $w=2.65e-07 $l=3.47851e-07 $layer=POLY_cond $X=8.125 $Y=1.22
+ $X2=7.85 $Y2=1.385
r275 16 18 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=8.125 $Y=1.22
+ $X2=8.125 $Y2=0.9
r276 13 45 61.4066 $w=2.86e-07 $l=3.21714e-07 $layer=POLY_cond $X=6.905 $Y=2.045
+ $X2=6.95 $Y2=1.745
r277 13 15 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=6.905 $Y=2.045
+ $X2=6.905 $Y2=2.54
r278 12 74 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=3.36 $Y=0.805
+ $X2=3.36 $Y2=1.125
r279 7 38 52.2586 $w=2.99e-07 $l=2.7157e-07 $layer=POLY_cond $X=3.025 $Y=2.44
+ $X2=3.07 $Y2=2.19
r280 7 9 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=3.025 $Y=2.44
+ $X2=3.025 $Y2=2.725
r281 2 50 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=1.02
+ $Y=1.84 $X2=1.17 $Y2=1.985
r282 2 22 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=1.02
+ $Y=1.84 $X2=1.17 $Y2=2.815
r283 1 25 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1 $Y=0.37
+ $X2=1.14 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__DFBBN_2%A_601_119# 1 2 7 8 9 11 12 14 16 17 21 24 26
+ 28 33
c107 17 0 1.48509e-19 $X=3.4 $Y=2.65
c108 16 0 4.11442e-20 $X=4.485 $Y=1.63
c109 7 0 1.56987e-19 $X=4.575 $Y=1.795
r110 35 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4 $Y=1.63
+ $X2=4 $Y2=1.63
r111 33 35 9.49416 $w=2.57e-07 $l=2e-07 $layer=LI1_cond $X=3.8 $Y=1.63 $X2=4
+ $Y2=1.63
r112 32 33 14.9533 $w=2.57e-07 $l=3.15e-07 $layer=LI1_cond $X=3.485 $Y=1.63
+ $X2=3.8 $Y2=1.63
r113 28 30 3.31764 $w=3.28e-07 $l=9.5e-08 $layer=LI1_cond $X=3.145 $Y=0.775
+ $X2=3.145 $Y2=0.87
r114 26 33 3.1561 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.8 $Y=1.465 $X2=3.8
+ $Y2=1.63
r115 25 26 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=3.8 $Y=0.955
+ $X2=3.8 $Y2=1.465
r116 23 32 3.1561 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.485 $Y=1.795
+ $X2=3.485 $Y2=1.63
r117 23 24 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=3.485 $Y=1.795
+ $X2=3.485 $Y2=2.565
r118 22 30 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.31 $Y=0.87
+ $X2=3.145 $Y2=0.87
r119 21 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.715 $Y=0.87
+ $X2=3.8 $Y2=0.955
r120 21 22 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=3.715 $Y=0.87
+ $X2=3.31 $Y2=0.87
r121 17 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.4 $Y=2.65
+ $X2=3.485 $Y2=2.565
r122 17 19 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=3.4 $Y=2.65
+ $X2=3.28 $Y2=2.65
r123 16 36 84.8077 $w=3.3e-07 $l=4.85e-07 $layer=POLY_cond $X=4.485 $Y=1.63
+ $X2=4 $Y2=1.63
r124 12 16 95.8357 $w=1.97e-07 $l=4.12602e-07 $layer=POLY_cond $X=4.695 $Y=1.25
+ $X2=4.627 $Y2=1.63
r125 12 14 112.467 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=4.695 $Y=1.25
+ $X2=4.695 $Y2=0.9
r126 9 11 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=4.575 $Y=2.045
+ $X2=4.575 $Y2=2.54
r127 8 9 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=4.575 $Y=1.955
+ $X2=4.575 $Y2=2.045
r128 7 16 40.8205 $w=1.97e-07 $l=1.89222e-07 $layer=POLY_cond $X=4.575 $Y=1.795
+ $X2=4.627 $Y2=1.63
r129 7 8 62.1936 $w=1.8e-07 $l=1.6e-07 $layer=POLY_cond $X=4.575 $Y=1.795
+ $X2=4.575 $Y2=1.955
r130 2 19 600 $w=1.7e-07 $l=2.38118e-07 $layer=licon1_PDIFF $count=1 $X=3.1
+ $Y=2.515 $X2=3.28 $Y2=2.65
r131 1 28 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=3.005
+ $Y=0.595 $X2=3.145 $Y2=0.775
.ends

.subckt PM_SKY130_FD_SC_HS__DFBBN_2%A_975_322# 1 2 7 9 12 16 18 19 21 23 24 25
+ 27 28 29 31 32 33 36 37 39 42 45 47 49 55 57 58 61
c185 57 0 1.31864e-19 $X=9.535 $Y=1.095
c186 49 0 1.49644e-19 $X=10.755 $Y=2.035
c187 37 0 6.04573e-20 $X=9.535 $Y=1.385
c188 36 0 2.26093e-19 $X=9.535 $Y=1.385
c189 33 0 1.87607e-19 $X=8.615 $Y=1.095
c190 29 0 1.32682e-19 $X=6.415 $Y=0.425
c191 23 0 1.56987e-19 $X=5.16 $Y=1.61
c192 19 0 2.60146e-19 $X=9.58 $Y=1.885
r193 52 55 4.1907 $w=3.28e-07 $l=1.2e-07 $layer=LI1_cond $X=5.04 $Y=1.775
+ $X2=5.16 $Y2=1.775
r194 52 53 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.04
+ $Y=1.775 $X2=5.04 $Y2=1.775
r195 47 49 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=10.545 $Y=2.035
+ $X2=10.755 $Y2=2.035
r196 43 58 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.545 $Y=1.095
+ $X2=10.46 $Y2=1.095
r197 43 45 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=10.545 $Y=1.095
+ $X2=10.825 $Y2=1.095
r198 42 47 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=10.46 $Y=1.95
+ $X2=10.545 $Y2=2.035
r199 41 58 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.46 $Y=1.18
+ $X2=10.46 $Y2=1.095
r200 41 42 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=10.46 $Y=1.18
+ $X2=10.46 $Y2=1.95
r201 40 57 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.7 $Y=1.095
+ $X2=9.535 $Y2=1.095
r202 39 58 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.375 $Y=1.095
+ $X2=10.46 $Y2=1.095
r203 39 40 44.0374 $w=1.68e-07 $l=6.75e-07 $layer=LI1_cond $X=10.375 $Y=1.095
+ $X2=9.7 $Y2=1.095
r204 37 62 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=9.535 $Y=1.385
+ $X2=9.535 $Y2=1.55
r205 37 61 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=9.535 $Y=1.385
+ $X2=9.535 $Y2=1.22
r206 36 37 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.535
+ $Y=1.385 $X2=9.535 $Y2=1.385
r207 34 57 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.535 $Y=1.18
+ $X2=9.535 $Y2=1.095
r208 34 36 7.15912 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=9.535 $Y=1.18
+ $X2=9.535 $Y2=1.385
r209 32 57 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.37 $Y=1.095
+ $X2=9.535 $Y2=1.095
r210 32 33 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=9.37 $Y=1.095
+ $X2=8.615 $Y2=1.095
r211 31 33 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.53 $Y=1.01
+ $X2=8.615 $Y2=1.095
r212 30 31 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=8.53 $Y=0.51 $X2=8.53
+ $Y2=1.01
r213 28 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.445 $Y=0.425
+ $X2=8.53 $Y2=0.51
r214 28 29 132.439 $w=1.68e-07 $l=2.03e-06 $layer=LI1_cond $X=8.445 $Y=0.425
+ $X2=6.415 $Y2=0.425
r215 26 29 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.33 $Y=0.51
+ $X2=6.415 $Y2=0.425
r216 26 27 50.8877 $w=1.68e-07 $l=7.8e-07 $layer=LI1_cond $X=6.33 $Y=0.51
+ $X2=6.33 $Y2=1.29
r217 24 27 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.245 $Y=1.375
+ $X2=6.33 $Y2=1.29
r218 24 25 65.2406 $w=1.68e-07 $l=1e-06 $layer=LI1_cond $X=6.245 $Y=1.375
+ $X2=5.245 $Y2=1.375
r219 23 55 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.16 $Y=1.61
+ $X2=5.16 $Y2=1.775
r220 22 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.16 $Y=1.46
+ $X2=5.245 $Y2=1.375
r221 22 23 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=5.16 $Y=1.46
+ $X2=5.16 $Y2=1.61
r222 19 21 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=9.58 $Y=1.885
+ $X2=9.58 $Y2=2.46
r223 18 19 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=9.58 $Y=1.795
+ $X2=9.58 $Y2=1.885
r224 18 62 95.2339 $w=1.8e-07 $l=2.45e-07 $layer=POLY_cond $X=9.58 $Y=1.795
+ $X2=9.58 $Y2=1.55
r225 16 61 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=9.515 $Y=0.74
+ $X2=9.515 $Y2=1.22
r226 10 53 38.5916 $w=2.93e-07 $l=2.03101e-07 $layer=POLY_cond $X=5.125 $Y=1.61
+ $X2=5.04 $Y2=1.775
r227 10 12 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=5.125 $Y=1.61
+ $X2=5.125 $Y2=0.9
r228 7 53 55.8646 $w=2.93e-07 $l=2.91633e-07 $layer=POLY_cond $X=4.995 $Y=2.045
+ $X2=5.04 $Y2=1.775
r229 7 9 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=4.995 $Y=2.045
+ $X2=4.995 $Y2=2.54
r230 2 49 600 $w=1.7e-07 $l=2.51744e-07 $layer=licon1_PDIFF $count=1 $X=10.625
+ $Y=1.84 $X2=10.755 $Y2=2.035
r231 1 45 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=10.685
+ $Y=0.82 $X2=10.825 $Y2=1.095
.ends

.subckt PM_SKY130_FD_SC_HS__DFBBN_2%SET_B 1 3 6 8 10 13 19 22 23 28 32 39
c128 8 0 1.25046e-19 $X=8.96 $Y=1.885
c129 6 0 1.08905e-19 $X=5.625 $Y=0.9
r130 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.58
+ $Y=1.795 $X2=5.58 $Y2=1.795
r131 28 39 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=2.035
+ $X2=8.88 $Y2=2.035
r132 26 32 8.3814 $w=3.28e-07 $l=2.4e-07 $layer=LI1_cond $X=5.58 $Y=2.035
+ $X2=5.58 $Y2=1.795
r133 25 26 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=2.035
+ $X2=5.52 $Y2=2.035
r134 23 25 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.665 $Y=2.035
+ $X2=5.52 $Y2=2.035
r135 22 28 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=8.735 $Y=2.035
+ $X2=8.88 $Y2=2.035
r136 22 23 3.7995 $w=1.4e-07 $l=3.07e-06 $layer=MET1_cond $X=8.735 $Y=2.035
+ $X2=5.665 $Y2=2.035
r137 19 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.995
+ $Y=1.615 $X2=8.995 $Y2=1.615
r138 16 39 12.7771 $w=2.28e-07 $l=2.55e-07 $layer=LI1_cond $X=8.88 $Y=1.78
+ $X2=8.88 $Y2=2.035
r139 15 19 4.01609 $w=3.28e-07 $l=1.15e-07 $layer=LI1_cond $X=8.88 $Y=1.615
+ $X2=8.995 $Y2=1.615
r140 15 16 2.85155 $w=2.3e-07 $l=1.65e-07 $layer=LI1_cond $X=8.88 $Y=1.615
+ $X2=8.88 $Y2=1.78
r141 11 20 38.5916 $w=2.93e-07 $l=2.05122e-07 $layer=POLY_cond $X=9.085 $Y=1.45
+ $X2=8.995 $Y2=1.615
r142 11 13 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=9.085 $Y=1.45
+ $X2=9.085 $Y2=0.74
r143 8 20 55.8646 $w=2.93e-07 $l=2.86967e-07 $layer=POLY_cond $X=8.96 $Y=1.885
+ $X2=8.995 $Y2=1.615
r144 8 10 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=8.96 $Y=1.885
+ $X2=8.96 $Y2=2.46
r145 4 31 38.5562 $w=2.99e-07 $l=1.86145e-07 $layer=POLY_cond $X=5.625 $Y=1.63
+ $X2=5.58 $Y2=1.795
r146 4 6 374.319 $w=1.5e-07 $l=7.3e-07 $layer=POLY_cond $X=5.625 $Y=1.63
+ $X2=5.625 $Y2=0.9
r147 1 31 52.2586 $w=2.99e-07 $l=2.85044e-07 $layer=POLY_cond $X=5.505 $Y=2.045
+ $X2=5.58 $Y2=1.795
r148 1 3 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=5.505 $Y=2.045
+ $X2=5.505 $Y2=2.54
.ends

.subckt PM_SKY130_FD_SC_HS__DFBBN_2%A_27_74# 1 2 10 11 13 14 15 19 20 22 23 25
+ 26 28 32 33 34 38 39 41 42 43 44 45 47 51 53 54 55 58 60 66
c191 33 0 1.71006e-19 $X=7.325 $Y=1.26
c192 32 0 1.06658e-19 $X=6.6 $Y=0.835
c193 19 0 6.36774e-20 $X=2.93 $Y=0.805
r194 66 67 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.96
+ $Y=1.465 $X2=0.96 $Y2=1.465
r195 63 66 7.33373 $w=3.28e-07 $l=2.1e-07 $layer=LI1_cond $X=0.75 $Y=1.465
+ $X2=0.96 $Y2=1.465
r196 59 63 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.75 $Y=1.63
+ $X2=0.75 $Y2=1.465
r197 59 60 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=0.75 $Y=1.63
+ $X2=0.75 $Y2=1.95
r198 58 63 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.75 $Y=1.3
+ $X2=0.75 $Y2=1.465
r199 57 58 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=0.75 $Y=1.13
+ $X2=0.75 $Y2=1.3
r200 56 62 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.435 $Y=2.035
+ $X2=0.27 $Y2=2.035
r201 55 60 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.665 $Y=2.035
+ $X2=0.75 $Y2=1.95
r202 55 56 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=0.665 $Y=2.035
+ $X2=0.435 $Y2=2.035
r203 53 57 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.665 $Y=1.045
+ $X2=0.75 $Y2=1.13
r204 53 54 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=0.665 $Y=1.045
+ $X2=0.365 $Y2=1.045
r205 49 54 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.24 $Y=0.96
+ $X2=0.365 $Y2=1.045
r206 49 51 20.5135 $w=2.48e-07 $l=4.45e-07 $layer=LI1_cond $X=0.24 $Y=0.96
+ $X2=0.24 $Y2=0.515
r207 45 62 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.27 $Y=2.12 $X2=0.27
+ $Y2=2.035
r208 45 47 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=0.27 $Y=2.12
+ $X2=0.27 $Y2=2.815
r209 43 44 60.4563 $w=1.8e-07 $l=1.5e-07 $layer=POLY_cond $X=7.43 $Y=1.79
+ $X2=7.43 $Y2=1.94
r210 39 41 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=7.445 $Y=2.465
+ $X2=7.445 $Y2=2.75
r211 38 39 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=7.445 $Y=2.375
+ $X2=7.445 $Y2=2.465
r212 38 44 169.089 $w=1.8e-07 $l=4.35e-07 $layer=POLY_cond $X=7.445 $Y=2.375
+ $X2=7.445 $Y2=1.94
r213 35 43 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=7.4 $Y=1.335
+ $X2=7.4 $Y2=1.79
r214 33 35 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=7.325 $Y=1.26
+ $X2=7.4 $Y2=1.335
r215 33 34 333.298 $w=1.5e-07 $l=6.5e-07 $layer=POLY_cond $X=7.325 $Y=1.26
+ $X2=6.675 $Y2=1.26
r216 30 34 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=6.6 $Y=1.185
+ $X2=6.675 $Y2=1.26
r217 30 32 179.468 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=6.6 $Y=1.185
+ $X2=6.6 $Y2=0.835
r218 29 32 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=6.6 $Y=0.255
+ $X2=6.6 $Y2=0.835
r219 26 28 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=3.535 $Y=2.44
+ $X2=3.535 $Y2=2.725
r220 25 26 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=3.535 $Y=2.35
+ $X2=3.535 $Y2=2.44
r221 24 25 207.96 $w=1.8e-07 $l=5.35e-07 $layer=POLY_cond $X=3.535 $Y=1.815
+ $X2=3.535 $Y2=2.35
r222 22 24 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=3.445 $Y=1.74
+ $X2=3.535 $Y2=1.815
r223 22 23 225.617 $w=1.5e-07 $l=4.4e-07 $layer=POLY_cond $X=3.445 $Y=1.74
+ $X2=3.005 $Y2=1.74
r224 21 42 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.005 $Y=0.18
+ $X2=2.93 $Y2=0.18
r225 20 29 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=6.525 $Y=0.18
+ $X2=6.6 $Y2=0.255
r226 20 21 1804.94 $w=1.5e-07 $l=3.52e-06 $layer=POLY_cond $X=6.525 $Y=0.18
+ $X2=3.005 $Y2=0.18
r227 17 23 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.93 $Y=1.665
+ $X2=3.005 $Y2=1.74
r228 17 19 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=2.93 $Y=1.665
+ $X2=2.93 $Y2=0.805
r229 16 42 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.93 $Y=0.255
+ $X2=2.93 $Y2=0.18
r230 16 19 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=2.93 $Y=0.255
+ $X2=2.93 $Y2=0.805
r231 14 42 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.855 $Y=0.18
+ $X2=2.93 $Y2=0.18
r232 14 15 951.181 $w=1.5e-07 $l=1.855e-06 $layer=POLY_cond $X=2.855 $Y=0.18
+ $X2=1 $Y2=0.18
r233 11 67 61.4066 $w=2.86e-07 $l=3.07409e-07 $layer=POLY_cond $X=0.945 $Y=1.765
+ $X2=0.96 $Y2=1.465
r234 11 13 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.945 $Y=1.765
+ $X2=0.945 $Y2=2.4
r235 8 67 38.6549 $w=2.86e-07 $l=1.81659e-07 $layer=POLY_cond $X=0.925 $Y=1.3
+ $X2=0.96 $Y2=1.465
r236 8 10 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=0.925 $Y=1.3
+ $X2=0.925 $Y2=0.74
r237 7 15 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.925 $Y=0.255
+ $X2=1 $Y2=0.18
r238 7 10 248.691 $w=1.5e-07 $l=4.85e-07 $layer=POLY_cond $X=0.925 $Y=0.255
+ $X2=0.925 $Y2=0.74
r239 2 62 400 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.27 $Y2=2.115
r240 2 47 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.27 $Y2=2.815
r241 1 51 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__DFBBN_2%A_1555_410# 1 2 3 10 12 14 17 19 21 22 24 25
+ 27 28 30 31 32 33 35 38 42 47 48 51 52 54 56 57 58 63 66 67 71 75 77
c223 56 0 1.20203e-19 $X=10.225 $Y=2.46
c224 33 0 1.79505e-19 $X=12.935 $Y=1.765
c225 19 0 1.91438e-19 $X=11.505 $Y=1.765
c226 2 0 4.70478e-20 $X=8.59 $Y=1.96
r227 85 86 7.16487 $w=3.7e-07 $l=5.5e-08 $layer=POLY_cond $X=11.955 $Y=1.557
+ $X2=12.01 $Y2=1.557
r228 84 85 48.8514 $w=3.7e-07 $l=3.75e-07 $layer=POLY_cond $X=11.58 $Y=1.557
+ $X2=11.955 $Y2=1.557
r229 83 84 9.77027 $w=3.7e-07 $l=7.5e-08 $layer=POLY_cond $X=11.505 $Y=1.557
+ $X2=11.58 $Y2=1.557
r230 76 83 1.95405 $w=3.7e-07 $l=1.5e-08 $layer=POLY_cond $X=11.49 $Y=1.557
+ $X2=11.505 $Y2=1.557
r231 75 78 8.49906 $w=3.53e-07 $l=1.65e-07 $layer=LI1_cond $X=11.467 $Y=1.515
+ $X2=11.467 $Y2=1.68
r232 75 77 8.49906 $w=3.53e-07 $l=1.65e-07 $layer=LI1_cond $X=11.467 $Y=1.515
+ $X2=11.467 $Y2=1.35
r233 75 76 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=11.49
+ $Y=1.515 $X2=11.49 $Y2=1.515
r234 69 71 8.85254 $w=2.43e-07 $l=1.65e-07 $layer=LI1_cond $X=9.77 $Y=0.717
+ $X2=9.935 $Y2=0.717
r235 65 67 8.48848 $w=3.48e-07 $l=1.65e-07 $layer=LI1_cond $X=8.735 $Y=2.805
+ $X2=8.9 $Y2=2.805
r236 65 66 8.48848 $w=3.48e-07 $l=1.65e-07 $layer=LI1_cond $X=8.735 $Y=2.805
+ $X2=8.57 $Y2=2.805
r237 63 78 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=11.375 $Y=2.29
+ $X2=11.375 $Y2=1.68
r238 60 77 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=11.375 $Y=0.84
+ $X2=11.375 $Y2=1.35
r239 59 73 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.39 $Y=2.375
+ $X2=10.225 $Y2=2.375
r240 58 63 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=11.29 $Y=2.375
+ $X2=11.375 $Y2=2.29
r241 58 59 58.7166 $w=1.68e-07 $l=9e-07 $layer=LI1_cond $X=11.29 $Y=2.375
+ $X2=10.39 $Y2=2.375
r242 56 73 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=10.225 $Y=2.46
+ $X2=10.225 $Y2=2.375
r243 56 57 5.93683 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=10.225 $Y=2.46
+ $X2=10.225 $Y2=2.63
r244 54 60 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=11.29 $Y=0.755
+ $X2=11.375 $Y2=0.84
r245 54 71 88.4011 $w=1.68e-07 $l=1.355e-06 $layer=LI1_cond $X=11.29 $Y=0.755
+ $X2=9.935 $Y2=0.755
r246 52 57 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=10.06 $Y=2.715
+ $X2=10.225 $Y2=2.63
r247 52 67 75.6791 $w=1.68e-07 $l=1.16e-06 $layer=LI1_cond $X=10.06 $Y=2.715
+ $X2=8.9 $Y2=2.715
r248 51 66 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=8.255 $Y=2.715
+ $X2=8.57 $Y2=2.715
r249 48 81 32.678 $w=3.54e-07 $l=2.4e-07 $layer=POLY_cond $X=8.09 $Y=2.257
+ $X2=8.33 $Y2=2.257
r250 48 79 30.6356 $w=3.54e-07 $l=2.25e-07 $layer=POLY_cond $X=8.09 $Y=2.257
+ $X2=7.865 $Y2=2.257
r251 47 48 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.09
+ $Y=2.215 $X2=8.09 $Y2=2.215
r252 45 51 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=8.09 $Y=2.63
+ $X2=8.255 $Y2=2.715
r253 45 47 14.4928 $w=3.28e-07 $l=4.15e-07 $layer=LI1_cond $X=8.09 $Y=2.63
+ $X2=8.09 $Y2=2.215
r254 40 42 94.8617 $w=1.5e-07 $l=1.85e-07 $layer=POLY_cond $X=8.33 $Y=1.81
+ $X2=8.515 $Y2=1.81
r255 36 38 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=13.015 $Y=1.35
+ $X2=13.015 $Y2=0.69
r256 33 35 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=12.935 $Y=1.765
+ $X2=12.935 $Y2=2.34
r257 32 86 10.4461 $w=3.7e-07 $l=9.3675e-08 $layer=POLY_cond $X=12.085 $Y=1.515
+ $X2=12.01 $Y2=1.557
r258 31 33 62.743 $w=2.03e-07 $l=2.65518e-07 $layer=POLY_cond $X=12.967 $Y=1.515
+ $X2=12.935 $Y2=1.765
r259 31 36 42.5607 $w=2.03e-07 $l=1.8747e-07 $layer=POLY_cond $X=12.967 $Y=1.515
+ $X2=13.015 $Y2=1.35
r260 31 32 132.895 $w=3.3e-07 $l=7.6e-07 $layer=POLY_cond $X=12.845 $Y=1.515
+ $X2=12.085 $Y2=1.515
r261 28 86 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=12.01 $Y=1.35
+ $X2=12.01 $Y2=1.557
r262 28 30 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=12.01 $Y=1.35
+ $X2=12.01 $Y2=0.87
r263 25 85 23.9667 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=11.955 $Y=1.765
+ $X2=11.955 $Y2=1.557
r264 25 27 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=11.955 $Y=1.765
+ $X2=11.955 $Y2=2.4
r265 22 84 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=11.58 $Y=1.35
+ $X2=11.58 $Y2=1.557
r266 22 24 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=11.58 $Y=1.35
+ $X2=11.58 $Y2=0.87
r267 19 83 23.9667 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=11.505 $Y=1.765
+ $X2=11.505 $Y2=1.557
r268 19 21 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=11.505 $Y=1.765
+ $X2=11.505 $Y2=2.4
r269 15 42 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=8.515 $Y=1.735
+ $X2=8.515 $Y2=1.81
r270 15 17 428.16 $w=1.5e-07 $l=8.35e-07 $layer=POLY_cond $X=8.515 $Y=1.735
+ $X2=8.515 $Y2=0.9
r271 14 81 22.9014 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=8.33 $Y=2.05
+ $X2=8.33 $Y2=2.257
r272 13 40 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=8.33 $Y=1.885
+ $X2=8.33 $Y2=1.81
r273 13 14 84.6064 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.33 $Y=1.885
+ $X2=8.33 $Y2=2.05
r274 10 79 22.9014 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=7.865 $Y=2.465
+ $X2=7.865 $Y2=2.257
r275 10 12 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=7.865 $Y=2.465
+ $X2=7.865 $Y2=2.75
r276 3 73 300 $w=1.7e-07 $l=5.65044e-07 $layer=licon1_PDIFF $count=2 $X=10.075
+ $Y=1.96 $X2=10.225 $Y2=2.455
r277 2 65 600 $w=1.7e-07 $l=9.14631e-07 $layer=licon1_PDIFF $count=1 $X=8.59
+ $Y=1.96 $X2=8.735 $Y2=2.805
r278 1 69 182 $w=1.7e-07 $l=4.25588e-07 $layer=licon1_NDIFF $count=1 $X=9.59
+ $Y=0.37 $X2=9.77 $Y2=0.715
.ends

.subckt PM_SKY130_FD_SC_HS__DFBBN_2%A_1335_112# 1 2 9 11 13 14 24 28 29 31 33 34
+ 35 36 37 39 40 42
c139 42 0 1.03189e-19 $X=8.51 $Y=1.805
c140 36 0 1.39943e-19 $X=9.805 $Y=1.89
c141 35 0 4.70478e-20 $X=8.595 $Y=2.375
c142 11 0 1.01047e-19 $X=10 $Y=1.885
r143 46 47 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.075
+ $Y=1.635 $X2=10.075 $Y2=1.635
r144 41 42 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=8.19 $Y=1.805
+ $X2=8.51 $Y2=1.805
r145 39 40 9.45624 $w=4.88e-07 $l=1.65e-07 $layer=LI1_cond $X=7.21 $Y=2.265
+ $X2=7.21 $Y2=2.1
r146 36 46 10.2298 $w=3.22e-07 $l=3.6e-07 $layer=LI1_cond $X=9.805 $Y=1.89
+ $X2=10.075 $Y2=1.68
r147 36 37 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=9.805 $Y=1.89
+ $X2=9.805 $Y2=2.29
r148 34 37 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.72 $Y=2.375
+ $X2=9.805 $Y2=2.29
r149 34 35 73.3957 $w=1.68e-07 $l=1.125e-06 $layer=LI1_cond $X=9.72 $Y=2.375
+ $X2=8.595 $Y2=2.375
r150 33 35 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.51 $Y=2.29
+ $X2=8.595 $Y2=2.375
r151 32 42 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.51 $Y=1.89
+ $X2=8.51 $Y2=1.805
r152 32 33 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=8.51 $Y=1.89 $X2=8.51
+ $Y2=2.29
r153 31 41 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.19 $Y=1.72
+ $X2=8.19 $Y2=1.805
r154 30 31 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=8.19 $Y=1.01
+ $X2=8.19 $Y2=1.72
r155 28 41 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=8.105 $Y=1.805
+ $X2=8.19 $Y2=1.805
r156 28 29 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=8.105 $Y=1.805
+ $X2=7.455 $Y2=1.805
r157 26 29 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.37 $Y=1.89
+ $X2=7.455 $Y2=1.805
r158 26 40 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=7.37 $Y=1.89
+ $X2=7.37 $Y2=2.1
r159 22 39 1.95278 $w=4.88e-07 $l=8e-08 $layer=LI1_cond $X=7.21 $Y=2.345
+ $X2=7.21 $Y2=2.265
r160 22 24 11.4726 $w=4.88e-07 $l=4.7e-07 $layer=LI1_cond $X=7.21 $Y=2.345
+ $X2=7.21 $Y2=2.815
r161 19 21 25.4934 $w=3.28e-07 $l=7.3e-07 $layer=LI1_cond $X=7.18 $Y=0.845
+ $X2=7.91 $Y2=0.845
r162 16 19 12.7467 $w=3.28e-07 $l=3.65e-07 $layer=LI1_cond $X=6.815 $Y=0.845
+ $X2=7.18 $Y2=0.845
r163 14 30 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=8.105 $Y=0.845
+ $X2=8.19 $Y2=1.01
r164 14 21 6.80989 $w=3.28e-07 $l=1.95e-07 $layer=LI1_cond $X=8.105 $Y=0.845
+ $X2=7.91 $Y2=0.845
r165 11 47 52.2586 $w=2.99e-07 $l=2.85044e-07 $layer=POLY_cond $X=10 $Y=1.885
+ $X2=10.075 $Y2=1.635
r166 11 13 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=10 $Y=1.885 $X2=10
+ $Y2=2.46
r167 7 47 38.5562 $w=2.99e-07 $l=2.05122e-07 $layer=POLY_cond $X=9.985 $Y=1.47
+ $X2=10.075 $Y2=1.635
r168 7 9 374.319 $w=1.5e-07 $l=7.3e-07 $layer=POLY_cond $X=9.985 $Y=1.47
+ $X2=9.985 $Y2=0.74
r169 2 39 600 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=6.98
+ $Y=2.12 $X2=7.13 $Y2=2.265
r170 2 24 600 $w=1.7e-07 $l=7.66339e-07 $layer=licon1_PDIFF $count=1 $X=6.98
+ $Y=2.12 $X2=7.13 $Y2=2.815
r171 1 21 121.333 $w=1.7e-07 $l=1.37011e-06 $layer=licon1_NDIFF $count=1
+ $X=6.675 $Y=0.56 $X2=7.91 $Y2=0.845
r172 1 19 121.333 $w=1.7e-07 $l=6.31625e-07 $layer=licon1_NDIFF $count=1
+ $X=6.675 $Y=0.56 $X2=7.18 $Y2=0.845
r173 1 16 182 $w=1.7e-07 $l=3.4803e-07 $layer=licon1_NDIFF $count=1 $X=6.675
+ $Y=0.56 $X2=6.815 $Y2=0.845
.ends

.subckt PM_SKY130_FD_SC_HS__DFBBN_2%RESET_B 1 3 4 6 7 11
c30 11 0 4.17943e-20 $X=10.95 $Y=1.515
c31 4 0 1.75691e-19 $X=11.04 $Y=1.35
r32 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.95
+ $Y=1.515 $X2=10.95 $Y2=1.515
r33 7 11 4.32166 $w=3.98e-07 $l=1.5e-07 $layer=LI1_cond $X=10.915 $Y=1.665
+ $X2=10.915 $Y2=1.515
r34 4 10 38.5562 $w=2.99e-07 $l=2.05122e-07 $layer=POLY_cond $X=11.04 $Y=1.35
+ $X2=10.95 $Y2=1.515
r35 4 6 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=11.04 $Y=1.35
+ $X2=11.04 $Y2=1.03
r36 1 10 52.2586 $w=2.99e-07 $l=2.64575e-07 $layer=POLY_cond $X=10.98 $Y=1.765
+ $X2=10.95 $Y2=1.515
r37 1 3 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=10.98 $Y=1.765
+ $X2=10.98 $Y2=2.16
.ends

.subckt PM_SKY130_FD_SC_HS__DFBBN_2%A_2516_368# 1 2 7 9 12 14 16 19 23 25 29 35
+ 38 39 43
c79 7 0 2.31826e-20 $X=13.455 $Y=1.765
r80 43 44 1.70519 $w=4.24e-07 $l=1.5e-08 $layer=POLY_cond $X=13.905 $Y=1.517
+ $X2=13.92 $Y2=1.517
r81 40 41 3.97877 $w=4.24e-07 $l=3.5e-08 $layer=POLY_cond $X=13.455 $Y=1.517
+ $X2=13.49 $Y2=1.517
r82 36 43 42.6297 $w=4.24e-07 $l=3.75e-07 $layer=POLY_cond $X=13.53 $Y=1.517
+ $X2=13.905 $Y2=1.517
r83 36 41 4.54717 $w=4.24e-07 $l=4e-08 $layer=POLY_cond $X=13.53 $Y=1.517
+ $X2=13.49 $Y2=1.517
r84 35 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=13.53
+ $Y=1.435 $X2=13.53 $Y2=1.435
r85 33 39 0.295496 $w=3.3e-07 $l=1.25e-07 $layer=LI1_cond $X=12.885 $Y=1.435
+ $X2=12.76 $Y2=1.435
r86 33 35 22.525 $w=3.28e-07 $l=6.45e-07 $layer=LI1_cond $X=12.885 $Y=1.435
+ $X2=13.53 $Y2=1.435
r87 31 39 6.56857 $w=2.45e-07 $l=1.67481e-07 $layer=LI1_cond $X=12.755 $Y=1.6
+ $X2=12.76 $Y2=1.435
r88 31 38 10.5641 $w=2.38e-07 $l=2.2e-07 $layer=LI1_cond $X=12.755 $Y=1.6
+ $X2=12.755 $Y2=1.82
r89 27 39 6.56857 $w=2.45e-07 $l=1.65e-07 $layer=LI1_cond $X=12.76 $Y=1.27
+ $X2=12.76 $Y2=1.435
r90 27 29 34.8038 $w=2.48e-07 $l=7.55e-07 $layer=LI1_cond $X=12.76 $Y=1.27
+ $X2=12.76 $Y2=0.515
r91 23 38 6.63994 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=12.71 $Y=1.985
+ $X2=12.71 $Y2=1.82
r92 23 25 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=12.71 $Y=1.985
+ $X2=12.71 $Y2=2.695
r93 17 44 27.2926 $w=1.5e-07 $l=2.47e-07 $layer=POLY_cond $X=13.92 $Y=1.27
+ $X2=13.92 $Y2=1.517
r94 17 19 271.766 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=13.92 $Y=1.27
+ $X2=13.92 $Y2=0.74
r95 14 43 27.2926 $w=1.5e-07 $l=2.48e-07 $layer=POLY_cond $X=13.905 $Y=1.765
+ $X2=13.905 $Y2=1.517
r96 14 16 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=13.905 $Y=1.765
+ $X2=13.905 $Y2=2.4
r97 10 41 27.2926 $w=1.5e-07 $l=2.47e-07 $layer=POLY_cond $X=13.49 $Y=1.27
+ $X2=13.49 $Y2=1.517
r98 10 12 271.766 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=13.49 $Y=1.27
+ $X2=13.49 $Y2=0.74
r99 7 40 27.2926 $w=1.5e-07 $l=2.48e-07 $layer=POLY_cond $X=13.455 $Y=1.765
+ $X2=13.455 $Y2=1.517
r100 7 9 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=13.455 $Y=1.765
+ $X2=13.455 $Y2=2.4
r101 2 25 400 $w=1.7e-07 $l=9.17701e-07 $layer=licon1_PDIFF $count=1 $X=12.58
+ $Y=1.84 $X2=12.71 $Y2=2.695
r102 2 23 400 $w=1.7e-07 $l=1.99687e-07 $layer=licon1_PDIFF $count=1 $X=12.58
+ $Y=1.84 $X2=12.71 $Y2=1.985
r103 1 29 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=12.655
+ $Y=0.37 $X2=12.8 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__DFBBN_2%VPWR 1 2 3 4 5 6 7 8 9 10 33 37 41 45 49 53
+ 57 61 63 66 67 69 70 72 73 75 78 81 83 110 114 119 124 129 135 138 145 148 151
+ 155
r173 154 155 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=14.16 $Y=3.33
+ $X2=14.16 $Y2=3.33
r174 151 152 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.2 $Y=3.33
+ $X2=13.2 $Y2=3.33
r175 148 149 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.24 $Y=3.33
+ $X2=12.24 $Y2=3.33
r176 145 146 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.28 $Y=3.33
+ $X2=11.28 $Y2=3.33
r177 141 142 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.36 $Y=3.33
+ $X2=9.36 $Y2=3.33
r178 138 141 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=9.27 $Y=3.055
+ $X2=9.27 $Y2=3.33
r179 135 136 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r180 133 155 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=13.68 $Y=3.33
+ $X2=14.16 $Y2=3.33
r181 133 152 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=13.68 $Y=3.33
+ $X2=13.2 $Y2=3.33
r182 132 133 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.68 $Y=3.33
+ $X2=13.68 $Y2=3.33
r183 130 151 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=13.315 $Y=3.33
+ $X2=13.19 $Y2=3.33
r184 130 132 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=13.315 $Y=3.33
+ $X2=13.68 $Y2=3.33
r185 129 154 4.02656 $w=1.7e-07 $l=1.77e-07 $layer=LI1_cond $X=14.045 $Y=3.33
+ $X2=14.222 $Y2=3.33
r186 129 132 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=14.045 $Y=3.33
+ $X2=13.68 $Y2=3.33
r187 128 152 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.72 $Y=3.33
+ $X2=13.2 $Y2=3.33
r188 128 149 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.72 $Y=3.33
+ $X2=12.24 $Y2=3.33
r189 127 128 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.72 $Y=3.33
+ $X2=12.72 $Y2=3.33
r190 125 148 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12.345 $Y=3.33
+ $X2=12.18 $Y2=3.33
r191 125 127 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=12.345 $Y=3.33
+ $X2=12.72 $Y2=3.33
r192 124 151 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=13.065 $Y=3.33
+ $X2=13.19 $Y2=3.33
r193 124 127 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=13.065 $Y=3.33
+ $X2=12.72 $Y2=3.33
r194 123 149 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.76 $Y=3.33
+ $X2=12.24 $Y2=3.33
r195 123 146 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.76 $Y=3.33
+ $X2=11.28 $Y2=3.33
r196 122 123 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.76 $Y=3.33
+ $X2=11.76 $Y2=3.33
r197 120 145 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.445 $Y=3.33
+ $X2=11.28 $Y2=3.33
r198 120 122 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=11.445 $Y=3.33
+ $X2=11.76 $Y2=3.33
r199 119 148 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12.015 $Y=3.33
+ $X2=12.18 $Y2=3.33
r200 119 122 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=12.015 $Y=3.33
+ $X2=11.76 $Y2=3.33
r201 118 146 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.8 $Y=3.33
+ $X2=11.28 $Y2=3.33
r202 118 142 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=10.8 $Y=3.33
+ $X2=9.36 $Y2=3.33
r203 117 118 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.8 $Y=3.33
+ $X2=10.8 $Y2=3.33
r204 115 141 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.435 $Y=3.33
+ $X2=9.27 $Y2=3.33
r205 115 117 89.0535 $w=1.68e-07 $l=1.365e-06 $layer=LI1_cond $X=9.435 $Y=3.33
+ $X2=10.8 $Y2=3.33
r206 114 145 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.115 $Y=3.33
+ $X2=11.28 $Y2=3.33
r207 114 117 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=11.115 $Y=3.33
+ $X2=10.8 $Y2=3.33
r208 113 142 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=3.33
+ $X2=9.36 $Y2=3.33
r209 112 113 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r210 110 141 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.105 $Y=3.33
+ $X2=9.27 $Y2=3.33
r211 110 112 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=9.105 $Y=3.33
+ $X2=8.88 $Y2=3.33
r212 109 113 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=7.92 $Y=3.33
+ $X2=8.88 $Y2=3.33
r213 108 109 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r214 105 108 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=6.48 $Y=3.33
+ $X2=7.92 $Y2=3.33
r215 105 106 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r216 103 106 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=3.33
+ $X2=6.48 $Y2=3.33
r217 102 103 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r218 100 103 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=6 $Y2=3.33
r219 99 100 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r220 97 100 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=5.04 $Y2=3.33
r221 96 99 156.578 $w=1.68e-07 $l=2.4e-06 $layer=LI1_cond $X=2.64 $Y=3.33
+ $X2=5.04 $Y2=3.33
r222 96 97 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r223 94 97 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r224 93 94 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r225 91 94 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.16 $Y2=3.33
r226 91 136 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r227 90 93 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.2 $Y=3.33 $X2=2.16
+ $Y2=3.33
r228 90 91 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r229 88 135 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.805 $Y=3.33
+ $X2=0.72 $Y2=3.33
r230 88 90 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=0.805 $Y=3.33
+ $X2=1.2 $Y2=3.33
r231 86 136 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r232 85 86 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r233 83 135 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.635 $Y=3.33
+ $X2=0.72 $Y2=3.33
r234 83 85 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=0.635 $Y=3.33
+ $X2=0.24 $Y2=3.33
r235 81 109 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=7.2 $Y=3.33
+ $X2=7.92 $Y2=3.33
r236 81 106 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=7.2 $Y=3.33
+ $X2=6.48 $Y2=3.33
r237 79 112 35.2299 $w=1.68e-07 $l=5.4e-07 $layer=LI1_cond $X=8.34 $Y=3.33
+ $X2=8.88 $Y2=3.33
r238 78 108 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=8.01 $Y=3.33
+ $X2=7.92 $Y2=3.33
r239 77 79 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.175 $Y=3.33
+ $X2=8.34 $Y2=3.33
r240 77 78 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.175 $Y=3.33
+ $X2=8.01 $Y2=3.33
r241 75 77 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=8.175 $Y=3.055
+ $X2=8.175 $Y2=3.33
r242 72 102 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=6.095 $Y=3.33
+ $X2=6 $Y2=3.33
r243 72 73 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.095 $Y=3.33
+ $X2=6.26 $Y2=3.33
r244 71 105 3.58824 $w=1.68e-07 $l=5.5e-08 $layer=LI1_cond $X=6.425 $Y=3.33
+ $X2=6.48 $Y2=3.33
r245 71 73 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.425 $Y=3.33
+ $X2=6.26 $Y2=3.33
r246 69 99 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=5.055 $Y=3.33
+ $X2=5.04 $Y2=3.33
r247 69 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.055 $Y=3.33
+ $X2=5.22 $Y2=3.33
r248 68 102 40.123 $w=1.68e-07 $l=6.15e-07 $layer=LI1_cond $X=5.385 $Y=3.33
+ $X2=6 $Y2=3.33
r249 68 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.385 $Y=3.33
+ $X2=5.22 $Y2=3.33
r250 66 93 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=2.295 $Y=3.33
+ $X2=2.16 $Y2=3.33
r251 66 67 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.295 $Y=3.33
+ $X2=2.38 $Y2=3.33
r252 65 96 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=2.465 $Y=3.33
+ $X2=2.64 $Y2=3.33
r253 65 67 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.465 $Y=3.33
+ $X2=2.38 $Y2=3.33
r254 61 154 3.1166 $w=2.5e-07 $l=1.07912e-07 $layer=LI1_cond $X=14.17 $Y=3.245
+ $X2=14.222 $Y2=3.33
r255 61 63 44.7148 $w=2.48e-07 $l=9.7e-07 $layer=LI1_cond $X=14.17 $Y=3.245
+ $X2=14.17 $Y2=2.275
r256 57 60 32.7294 $w=2.48e-07 $l=7.1e-07 $layer=LI1_cond $X=13.19 $Y=1.985
+ $X2=13.19 $Y2=2.695
r257 55 151 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=13.19 $Y=3.245
+ $X2=13.19 $Y2=3.33
r258 55 60 25.3537 $w=2.48e-07 $l=5.5e-07 $layer=LI1_cond $X=13.19 $Y=3.245
+ $X2=13.19 $Y2=2.695
r259 51 148 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=12.18 $Y=3.245
+ $X2=12.18 $Y2=3.33
r260 51 53 31.081 $w=3.28e-07 $l=8.9e-07 $layer=LI1_cond $X=12.18 $Y=3.245
+ $X2=12.18 $Y2=2.355
r261 47 145 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=11.28 $Y=3.245
+ $X2=11.28 $Y2=3.33
r262 47 49 15.3659 $w=3.28e-07 $l=4.4e-07 $layer=LI1_cond $X=11.28 $Y=3.245
+ $X2=11.28 $Y2=2.805
r263 43 73 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.26 $Y=3.245
+ $X2=6.26 $Y2=3.33
r264 43 45 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=6.26 $Y=3.245
+ $X2=6.26 $Y2=2.78
r265 39 70 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.22 $Y=3.245
+ $X2=5.22 $Y2=3.33
r266 39 41 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=5.22 $Y=3.245
+ $X2=5.22 $Y2=2.78
r267 35 67 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.38 $Y=3.245
+ $X2=2.38 $Y2=3.33
r268 35 37 32.9465 $w=1.68e-07 $l=5.05e-07 $layer=LI1_cond $X=2.38 $Y=3.245
+ $X2=2.38 $Y2=2.74
r269 31 135 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.72 $Y=3.245
+ $X2=0.72 $Y2=3.33
r270 31 33 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=0.72 $Y=3.245
+ $X2=0.72 $Y2=2.455
r271 10 63 300 $w=1.7e-07 $l=5.04455e-07 $layer=licon1_PDIFF $count=2 $X=13.98
+ $Y=1.84 $X2=14.13 $Y2=2.275
r272 9 60 400 $w=1.7e-07 $l=9.5871e-07 $layer=licon1_PDIFF $count=1 $X=13.01
+ $Y=1.84 $X2=13.23 $Y2=2.695
r273 9 57 400 $w=1.7e-07 $l=2.83373e-07 $layer=licon1_PDIFF $count=1 $X=13.01
+ $Y=1.84 $X2=13.23 $Y2=1.985
r274 8 53 300 $w=1.7e-07 $l=5.85214e-07 $layer=licon1_PDIFF $count=2 $X=12.03
+ $Y=1.84 $X2=12.18 $Y2=2.355
r275 7 49 600 $w=1.7e-07 $l=1.07161e-06 $layer=licon1_PDIFF $count=1 $X=11.055
+ $Y=1.84 $X2=11.28 $Y2=2.805
r276 6 138 600 $w=1.7e-07 $l=1.20679e-06 $layer=licon1_PDIFF $count=1 $X=9.035
+ $Y=1.96 $X2=9.27 $Y2=3.055
r277 5 75 600 $w=1.7e-07 $l=6.2149e-07 $layer=licon1_PDIFF $count=1 $X=7.94
+ $Y=2.54 $X2=8.175 $Y2=3.055
r278 4 45 600 $w=1.7e-07 $l=7.2208e-07 $layer=licon1_PDIFF $count=1 $X=6.13
+ $Y=2.12 $X2=6.26 $Y2=2.78
r279 3 41 600 $w=1.7e-07 $l=7.31163e-07 $layer=licon1_PDIFF $count=1 $X=5.07
+ $Y=2.12 $X2=5.22 $Y2=2.78
r280 2 37 600 $w=1.7e-07 $l=3.91663e-07 $layer=licon1_PDIFF $count=1 $X=2.085
+ $Y=2.515 $X2=2.38 $Y2=2.74
r281 1 33 300 $w=1.7e-07 $l=6.85912e-07 $layer=licon1_PDIFF $count=2 $X=0.57
+ $Y=1.84 $X2=0.72 $Y2=2.455
.ends

.subckt PM_SKY130_FD_SC_HS__DFBBN_2%A_311_119# 1 2 3 4 15 17 20 22 23 24 29 31
+ 32 34 36 38 42 45
r121 43 45 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=4.14 $Y=1.21
+ $X2=4.35 $Y2=1.21
r122 40 41 5.10546 $w=2.48e-07 $l=8.5e-08 $layer=LI1_cond $X=1.74 $Y=0.925
+ $X2=1.74 $Y2=1.01
r123 38 40 6.22319 $w=2.48e-07 $l=1.35e-07 $layer=LI1_cond $X=1.74 $Y=0.79
+ $X2=1.74 $Y2=0.925
r124 35 45 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.35 $Y=1.295
+ $X2=4.35 $Y2=1.21
r125 35 36 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.35 $Y=1.295
+ $X2=4.35 $Y2=1.965
r126 34 43 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.14 $Y=1.125
+ $X2=4.14 $Y2=1.21
r127 33 34 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=4.14 $Y=0.615
+ $X2=4.14 $Y2=1.125
r128 31 36 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.265 $Y=2.05
+ $X2=4.35 $Y2=1.965
r129 31 32 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=4.265 $Y=2.05
+ $X2=3.99 $Y2=2.05
r130 27 32 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=3.865 $Y=2.135
+ $X2=3.99 $Y2=2.05
r131 27 29 20.0525 $w=2.48e-07 $l=4.35e-07 $layer=LI1_cond $X=3.865 $Y=2.135
+ $X2=3.865 $Y2=2.57
r132 24 42 8.99121 $w=3.58e-07 $l=1.8e-07 $layer=LI1_cond $X=3.67 $Y=0.435
+ $X2=3.49 $Y2=0.435
r133 24 26 3.68142 $w=3.58e-07 $l=1.15e-07 $layer=LI1_cond $X=3.67 $Y=0.435
+ $X2=3.785 $Y2=0.435
r134 23 33 8.02311 $w=3.6e-07 $l=2.18403e-07 $layer=LI1_cond $X=4.055 $Y=0.435
+ $X2=4.14 $Y2=0.615
r135 23 26 8.64332 $w=3.58e-07 $l=2.7e-07 $layer=LI1_cond $X=4.055 $Y=0.435
+ $X2=3.785 $Y2=0.435
r136 22 42 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=2.78 $Y=0.34
+ $X2=3.49 $Y2=0.34
r137 19 22 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.695 $Y=0.425
+ $X2=2.78 $Y2=0.34
r138 19 20 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=2.695 $Y=0.425
+ $X2=2.695 $Y2=0.84
r139 18 40 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.865 $Y=0.925
+ $X2=1.74 $Y2=0.925
r140 17 20 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.61 $Y=0.925
+ $X2=2.695 $Y2=0.84
r141 17 18 48.6043 $w=1.68e-07 $l=7.45e-07 $layer=LI1_cond $X=2.61 $Y=0.925
+ $X2=1.865 $Y2=0.925
r142 15 41 101.775 $w=1.68e-07 $l=1.56e-06 $layer=LI1_cond $X=1.7 $Y=2.57
+ $X2=1.7 $Y2=1.01
r143 4 29 600 $w=1.7e-07 $l=2.40936e-07 $layer=licon1_PDIFF $count=1 $X=3.61
+ $Y=2.515 $X2=3.825 $Y2=2.57
r144 3 15 600 $w=1.7e-07 $l=1.99687e-07 $layer=licon1_PDIFF $count=1 $X=1.57
+ $Y=2.425 $X2=1.7 $Y2=2.57
r145 2 26 182 $w=1.7e-07 $l=3.81117e-07 $layer=licon1_NDIFF $count=1 $X=3.435
+ $Y=0.595 $X2=3.785 $Y2=0.53
r146 1 38 182 $w=1.7e-07 $l=2.57488e-07 $layer=licon1_NDIFF $count=1 $X=1.555
+ $Y=0.595 $X2=1.7 $Y2=0.79
.ends

.subckt PM_SKY130_FD_SC_HS__DFBBN_2%Q_N 1 2 9 12 16 18 19 31
c38 18 0 1.75691e-19 $X=11.76 $Y=0.555
r39 23 31 2.53213 $w=3.53e-07 $l=7.8e-08 $layer=LI1_cond $X=11.807 $Y=1.003
+ $X2=11.807 $Y2=0.925
r40 19 33 8.79122 $w=3.53e-07 $l=1.74e-07 $layer=LI1_cond $X=11.807 $Y=1.006
+ $X2=11.807 $Y2=1.18
r41 19 23 0.0973895 $w=3.53e-07 $l=3e-09 $layer=LI1_cond $X=11.807 $Y=1.006
+ $X2=11.807 $Y2=1.003
r42 19 31 0.129853 $w=3.53e-07 $l=4e-09 $layer=LI1_cond $X=11.807 $Y=0.921
+ $X2=11.807 $Y2=0.925
r43 19 28 8.95984 $w=3.53e-07 $l=2.76e-07 $layer=LI1_cond $X=11.807 $Y=0.921
+ $X2=11.807 $Y2=0.645
r44 18 28 2.92169 $w=3.53e-07 $l=9e-08 $layer=LI1_cond $X=11.807 $Y=0.555
+ $X2=11.807 $Y2=0.645
r45 14 16 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=11.73 $Y=1.935
+ $X2=11.9 $Y2=1.935
r46 12 16 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=11.9 $Y=1.85
+ $X2=11.9 $Y2=1.935
r47 12 33 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=11.9 $Y=1.85
+ $X2=11.9 $Y2=1.18
r48 7 14 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=11.73 $Y=2.02
+ $X2=11.73 $Y2=1.935
r49 7 9 51.8663 $w=1.68e-07 $l=7.95e-07 $layer=LI1_cond $X=11.73 $Y=2.02
+ $X2=11.73 $Y2=2.815
r50 2 14 400 $w=1.7e-07 $l=2.38485e-07 $layer=licon1_PDIFF $count=1 $X=11.58
+ $Y=1.84 $X2=11.73 $Y2=2.015
r51 2 9 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=11.58
+ $Y=1.84 $X2=11.73 $Y2=2.815
r52 1 28 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=11.655
+ $Y=0.5 $X2=11.795 $Y2=0.645
.ends

.subckt PM_SKY130_FD_SC_HS__DFBBN_2%Q 1 2 9 12 16 21 23 24 25
c36 16 0 1.79505e-19 $X=13.95 $Y=1.855
c37 12 0 2.31826e-20 $X=13.95 $Y=1.77
r38 24 25 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=13.68 $Y=2.405
+ $X2=13.68 $Y2=2.775
r39 23 24 14.6675 $w=3.28e-07 $l=4.2e-07 $layer=LI1_cond $X=13.68 $Y=1.985
+ $X2=13.68 $Y2=2.405
r40 20 21 12.9074 $w=2.48e-07 $l=2.8e-07 $layer=LI1_cond $X=13.67 $Y=0.975
+ $X2=13.95 $Y2=0.975
r41 14 23 1.57151 $w=3.28e-07 $l=4.5e-08 $layer=LI1_cond $X=13.68 $Y=1.94
+ $X2=13.68 $Y2=1.985
r42 14 16 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=13.68 $Y=1.855
+ $X2=13.95 $Y2=1.855
r43 12 16 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=13.95 $Y=1.77
+ $X2=13.95 $Y2=1.855
r44 11 21 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=13.95 $Y=1.1
+ $X2=13.95 $Y2=0.975
r45 11 12 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=13.95 $Y=1.1
+ $X2=13.95 $Y2=1.77
r46 7 20 0.475901 $w=2.6e-07 $l=1.25e-07 $layer=LI1_cond $X=13.67 $Y=0.85
+ $X2=13.67 $Y2=0.975
r47 7 9 14.8488 $w=2.58e-07 $l=3.35e-07 $layer=LI1_cond $X=13.67 $Y=0.85
+ $X2=13.67 $Y2=0.515
r48 2 25 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=13.53
+ $Y=1.84 $X2=13.68 $Y2=2.815
r49 2 23 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=13.53
+ $Y=1.84 $X2=13.68 $Y2=1.985
r50 1 20 182 $w=1.7e-07 $l=6.3113e-07 $layer=licon1_NDIFF $count=1 $X=13.565
+ $Y=0.37 $X2=13.705 $Y2=0.935
r51 1 9 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=13.565
+ $Y=0.37 $X2=13.705 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__DFBBN_2%VGND 1 2 3 4 5 6 7 8 27 31 35 39 43 47 49 51
+ 53 55 60 65 73 83 88 93 99 102 105 108 113 119 121 124 128
r145 127 128 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=14.16 $Y=0
+ $X2=14.16 $Y2=0
r146 124 125 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.2 $Y=0
+ $X2=13.2 $Y2=0
r147 121 122 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.24 $Y=0
+ $X2=12.24 $Y2=0
r148 118 119 10.0584 $w=5.83e-07 $l=1.65e-07 $layer=LI1_cond $X=11.285 $Y=0.207
+ $X2=11.45 $Y2=0.207
r149 115 118 0.102229 $w=5.83e-07 $l=5e-09 $layer=LI1_cond $X=11.28 $Y=0.207
+ $X2=11.285 $Y2=0.207
r150 115 116 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.28 $Y=0
+ $X2=11.28 $Y2=0
r151 112 116 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.8 $Y=0
+ $X2=11.28 $Y2=0
r152 111 115 9.81398 $w=5.83e-07 $l=4.8e-07 $layer=LI1_cond $X=10.8 $Y=0.207
+ $X2=11.28 $Y2=0.207
r153 111 113 9.44502 $w=5.83e-07 $l=1.35e-07 $layer=LI1_cond $X=10.8 $Y=0.207
+ $X2=10.665 $Y2=0.207
r154 111 112 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.8 $Y=0
+ $X2=10.8 $Y2=0
r155 108 109 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.88 $Y=0
+ $X2=8.88 $Y2=0
r156 105 106 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=6 $Y=0 $X2=6
+ $Y2=0
r157 102 103 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0
+ $X2=2.16 $Y2=0
r158 99 100 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r159 97 128 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=13.68 $Y=0
+ $X2=14.16 $Y2=0
r160 97 125 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=13.68 $Y=0
+ $X2=13.2 $Y2=0
r161 96 97 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.68 $Y=0
+ $X2=13.68 $Y2=0
r162 94 124 7.54988 $w=1.7e-07 $l=1.38e-07 $layer=LI1_cond $X=13.37 $Y=0
+ $X2=13.232 $Y2=0
r163 94 96 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=13.37 $Y=0
+ $X2=13.68 $Y2=0
r164 93 127 4.77065 $w=1.7e-07 $l=2.15e-07 $layer=LI1_cond $X=13.97 $Y=0
+ $X2=14.185 $Y2=0
r165 93 96 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=13.97 $Y=0
+ $X2=13.68 $Y2=0
r166 92 125 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.72 $Y=0
+ $X2=13.2 $Y2=0
r167 92 122 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.72 $Y=0
+ $X2=12.24 $Y2=0
r168 91 92 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.72 $Y=0
+ $X2=12.72 $Y2=0
r169 89 121 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=12.405 $Y=0
+ $X2=12.28 $Y2=0
r170 89 91 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=12.405 $Y=0
+ $X2=12.72 $Y2=0
r171 88 124 7.54988 $w=1.7e-07 $l=1.37e-07 $layer=LI1_cond $X=13.095 $Y=0
+ $X2=13.232 $Y2=0
r172 88 91 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=13.095 $Y=0
+ $X2=12.72 $Y2=0
r173 87 122 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.76 $Y=0
+ $X2=12.24 $Y2=0
r174 87 116 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.76 $Y=0
+ $X2=11.28 $Y2=0
r175 86 119 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=11.76 $Y=0
+ $X2=11.45 $Y2=0
r176 86 87 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.76 $Y=0
+ $X2=11.76 $Y2=0
r177 83 121 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=12.155 $Y=0
+ $X2=12.28 $Y2=0
r178 83 86 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=12.155 $Y=0
+ $X2=11.76 $Y2=0
r179 82 112 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.32 $Y=0
+ $X2=10.8 $Y2=0
r180 82 109 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=10.32 $Y=0
+ $X2=8.88 $Y2=0
r181 81 113 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=10.32 $Y=0
+ $X2=10.665 $Y2=0
r182 81 82 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.32 $Y=0
+ $X2=10.32 $Y2=0
r183 79 108 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.955 $Y=0 $X2=8.87
+ $Y2=0
r184 79 81 89.0535 $w=1.68e-07 $l=1.365e-06 $layer=LI1_cond $X=8.955 $Y=0
+ $X2=10.32 $Y2=0
r185 77 109 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=0 $X2=8.88
+ $Y2=0
r186 76 77 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r187 74 105 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.075 $Y=0
+ $X2=5.91 $Y2=0
r188 74 76 151.684 $w=1.68e-07 $l=2.325e-06 $layer=LI1_cond $X=6.075 $Y=0
+ $X2=8.4 $Y2=0
r189 73 108 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.785 $Y=0 $X2=8.87
+ $Y2=0
r190 73 76 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=8.785 $Y=0 $X2=8.4
+ $Y2=0
r191 72 106 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=6
+ $Y2=0
r192 71 72 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=5.52 $Y=0
+ $X2=5.52 $Y2=0
r193 69 72 0.802756 $w=4.9e-07 $l=2.88e-06 $layer=MET1_cond $X=2.64 $Y=0
+ $X2=5.52 $Y2=0
r194 69 103 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0
+ $X2=2.16 $Y2=0
r195 68 71 187.893 $w=1.68e-07 $l=2.88e-06 $layer=LI1_cond $X=2.64 $Y=0 $X2=5.52
+ $Y2=0
r196 68 69 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=2.64 $Y=0
+ $X2=2.64 $Y2=0
r197 66 102 9.73034 $w=1.7e-07 $l=1.98e-07 $layer=LI1_cond $X=2.44 $Y=0
+ $X2=2.242 $Y2=0
r198 66 68 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=2.44 $Y=0 $X2=2.64
+ $Y2=0
r199 65 105 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.745 $Y=0
+ $X2=5.91 $Y2=0
r200 65 71 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=5.745 $Y=0
+ $X2=5.52 $Y2=0
r201 64 103 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0
+ $X2=2.16 $Y2=0
r202 64 100 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0
+ $X2=0.72 $Y2=0
r203 63 64 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r204 61 99 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.875 $Y=0 $X2=0.71
+ $Y2=0
r205 61 63 52.5187 $w=1.68e-07 $l=8.05e-07 $layer=LI1_cond $X=0.875 $Y=0
+ $X2=1.68 $Y2=0
r206 60 102 9.73034 $w=1.7e-07 $l=1.97e-07 $layer=LI1_cond $X=2.045 $Y=0
+ $X2=2.242 $Y2=0
r207 60 63 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=2.045 $Y=0
+ $X2=1.68 $Y2=0
r208 58 100 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0
+ $X2=0.72 $Y2=0
r209 57 58 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r210 55 99 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.545 $Y=0 $X2=0.71
+ $Y2=0
r211 55 57 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.545 $Y=0
+ $X2=0.24 $Y2=0
r212 53 77 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=7.2 $Y=0 $X2=8.4
+ $Y2=0
r213 53 106 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=7.2 $Y=0 $X2=6
+ $Y2=0
r214 49 127 2.99552 $w=3.3e-07 $l=1.07121e-07 $layer=LI1_cond $X=14.135 $Y=0.085
+ $X2=14.185 $Y2=0
r215 49 51 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=14.135 $Y=0.085
+ $X2=14.135 $Y2=0.515
r216 45 124 0.316938 $w=2.75e-07 $l=8.5e-08 $layer=LI1_cond $X=13.232 $Y=0.085
+ $X2=13.232 $Y2=0
r217 45 47 17.1819 $w=2.73e-07 $l=4.1e-07 $layer=LI1_cond $X=13.232 $Y=0.085
+ $X2=13.232 $Y2=0.495
r218 41 121 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=12.28 $Y=0.085
+ $X2=12.28 $Y2=0
r219 41 43 25.8147 $w=2.48e-07 $l=5.6e-07 $layer=LI1_cond $X=12.28 $Y=0.085
+ $X2=12.28 $Y2=0.645
r220 37 108 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.87 $Y=0.085
+ $X2=8.87 $Y2=0
r221 37 39 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=8.87 $Y=0.085
+ $X2=8.87 $Y2=0.595
r222 33 105 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.91 $Y=0.085
+ $X2=5.91 $Y2=0
r223 33 35 27.0649 $w=3.28e-07 $l=7.75e-07 $layer=LI1_cond $X=5.91 $Y=0.085
+ $X2=5.91 $Y2=0.86
r224 29 102 1.43204 $w=3.95e-07 $l=8.5e-08 $layer=LI1_cond $X=2.242 $Y=0.085
+ $X2=2.242 $Y2=0
r225 29 31 14.5879 $w=3.93e-07 $l=5e-07 $layer=LI1_cond $X=2.242 $Y=0.085
+ $X2=2.242 $Y2=0.585
r226 25 99 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.71 $Y=0.085
+ $X2=0.71 $Y2=0
r227 25 27 18.8582 $w=3.28e-07 $l=5.4e-07 $layer=LI1_cond $X=0.71 $Y=0.085
+ $X2=0.71 $Y2=0.625
r228 8 51 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=13.995
+ $Y=0.37 $X2=14.135 $Y2=0.515
r229 7 47 91 $w=1.7e-07 $l=2.23942e-07 $layer=licon1_NDIFF $count=2 $X=13.09
+ $Y=0.37 $X2=13.26 $Y2=0.495
r230 6 43 91 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_NDIFF $count=2 $X=12.085
+ $Y=0.5 $X2=12.24 $Y2=0.645
r231 5 118 91 $w=1.7e-07 $l=6.68581e-07 $layer=licon1_NDIFF $count=2 $X=10.685
+ $Y=0.19 $X2=11.285 $Y2=0.335
r232 4 39 182 $w=1.7e-07 $l=3.24037e-07 $layer=licon1_NDIFF $count=1 $X=8.59
+ $Y=0.69 $X2=8.87 $Y2=0.595
r233 3 35 182 $w=1.7e-07 $l=3.23381e-07 $layer=licon1_NDIFF $count=1 $X=5.7
+ $Y=0.625 $X2=5.91 $Y2=0.86
r234 2 31 182 $w=1.7e-07 $l=2.54951e-07 $layer=licon1_NDIFF $count=1 $X=1.99
+ $Y=0.595 $X2=2.24 $Y2=0.585
r235 1 27 182 $w=1.7e-07 $l=3.17372e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.37 $X2=0.71 $Y2=0.625
.ends

.subckt PM_SKY130_FD_SC_HS__DFBBN_2%A_867_125# 1 2 9 11 12 15
r31 13 15 14.8421 $w=3.28e-07 $l=4.25e-07 $layer=LI1_cond $X=5.41 $Y=0.435
+ $X2=5.41 $Y2=0.86
r32 11 13 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=5.245 $Y=0.35
+ $X2=5.41 $Y2=0.435
r33 11 12 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=5.245 $Y=0.35
+ $X2=4.565 $Y2=0.35
r34 7 12 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.48 $Y=0.435
+ $X2=4.565 $Y2=0.35
r35 7 9 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=4.48 $Y=0.435 $X2=4.48
+ $Y2=0.78
r36 2 15 182 $w=1.7e-07 $l=3.23381e-07 $layer=licon1_NDIFF $count=1 $X=5.2
+ $Y=0.625 $X2=5.41 $Y2=0.86
r37 1 9 182 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_NDIFF $count=1 $X=4.335
+ $Y=0.625 $X2=4.48 $Y2=0.78
.ends

.subckt PM_SKY130_FD_SC_HS__DFBBN_2%A_1832_74# 1 2 9 12 14 15
c24 9 0 6.04573e-20 $X=9.3 $Y=0.595
c25 1 0 1.31864e-19 $X=9.16 $Y=0.37
r26 14 15 8.85254 $w=2.43e-07 $l=1.65e-07 $layer=LI1_cond $X=10.275 $Y=0.377
+ $X2=10.11 $Y2=0.377
r27 12 15 47.2995 $w=1.68e-07 $l=7.25e-07 $layer=LI1_cond $X=9.385 $Y=0.34
+ $X2=10.11 $Y2=0.34
r28 7 12 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=9.26 $Y=0.425
+ $X2=9.385 $Y2=0.34
r29 7 9 7.83661 $w=2.48e-07 $l=1.7e-07 $layer=LI1_cond $X=9.26 $Y=0.425 $X2=9.26
+ $Y2=0.595
r30 2 14 182 $w=1.7e-07 $l=2.36432e-07 $layer=licon1_NDIFF $count=1 $X=10.06
+ $Y=0.37 $X2=10.275 $Y2=0.415
r31 1 9 182 $w=1.7e-07 $l=2.86575e-07 $layer=licon1_NDIFF $count=1 $X=9.16
+ $Y=0.37 $X2=9.3 $Y2=0.595
.ends

