* File: sky130_fd_sc_hs__dlygate4sd3_1.pxi.spice
* Created: Thu Aug 27 20:43:24 2020
* 
x_PM_SKY130_FD_SC_HS__DLYGATE4SD3_1%A N_A_M1004_g N_A_c_64_n N_A_c_68_n
+ N_A_M1007_g A A N_A_c_66_n PM_SKY130_FD_SC_HS__DLYGATE4SD3_1%A
x_PM_SKY130_FD_SC_HS__DLYGATE4SD3_1%A_28_74# N_A_28_74#_M1004_s
+ N_A_28_74#_M1007_s N_A_28_74#_M1003_g N_A_28_74#_M1000_g N_A_28_74#_c_101_n
+ N_A_28_74#_c_107_n N_A_28_74#_c_108_n N_A_28_74#_c_109_n N_A_28_74#_c_102_n
+ N_A_28_74#_c_103_n N_A_28_74#_c_104_n N_A_28_74#_c_105_n
+ PM_SKY130_FD_SC_HS__DLYGATE4SD3_1%A_28_74#
x_PM_SKY130_FD_SC_HS__DLYGATE4SD3_1%A_289_74# N_A_289_74#_M1000_d
+ N_A_289_74#_M1003_d N_A_289_74#_M1001_g N_A_289_74#_M1005_g
+ N_A_289_74#_c_160_n N_A_289_74#_c_161_n N_A_289_74#_c_162_n
+ N_A_289_74#_c_163_n N_A_289_74#_c_167_n N_A_289_74#_c_164_n
+ N_A_289_74#_c_165_n PM_SKY130_FD_SC_HS__DLYGATE4SD3_1%A_289_74#
x_PM_SKY130_FD_SC_HS__DLYGATE4SD3_1%A_405_138# N_A_405_138#_M1005_s
+ N_A_405_138#_M1001_s N_A_405_138#_M1006_g N_A_405_138#_c_213_n
+ N_A_405_138#_M1002_g N_A_405_138#_c_214_n N_A_405_138#_c_219_n
+ N_A_405_138#_c_215_n N_A_405_138#_c_216_n N_A_405_138#_c_217_n
+ N_A_405_138#_c_221_n PM_SKY130_FD_SC_HS__DLYGATE4SD3_1%A_405_138#
x_PM_SKY130_FD_SC_HS__DLYGATE4SD3_1%VPWR N_VPWR_M1007_d N_VPWR_M1001_d
+ N_VPWR_c_269_n N_VPWR_c_270_n N_VPWR_c_271_n N_VPWR_c_272_n VPWR
+ N_VPWR_c_273_n N_VPWR_c_274_n N_VPWR_c_268_n N_VPWR_c_276_n
+ PM_SKY130_FD_SC_HS__DLYGATE4SD3_1%VPWR
x_PM_SKY130_FD_SC_HS__DLYGATE4SD3_1%X N_X_M1006_d N_X_M1002_d X X X X X X X
+ N_X_c_301_n X X N_X_c_305_n PM_SKY130_FD_SC_HS__DLYGATE4SD3_1%X
x_PM_SKY130_FD_SC_HS__DLYGATE4SD3_1%VGND N_VGND_M1004_d N_VGND_M1005_d
+ N_VGND_c_321_n N_VGND_c_322_n N_VGND_c_323_n N_VGND_c_324_n VGND
+ N_VGND_c_325_n N_VGND_c_326_n N_VGND_c_327_n N_VGND_c_328_n
+ PM_SKY130_FD_SC_HS__DLYGATE4SD3_1%VGND
cc_1 VNB N_A_M1004_g 0.0471271f $X=-0.19 $Y=-0.245 $X2=0.48 $Y2=0.58
cc_2 VNB N_A_c_64_n 0.00890285f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.17
cc_3 VNB A 0.0265853f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_4 VNB N_A_c_66_n 0.0358668f $X=-0.19 $Y=-0.245 $X2=0.57 $Y2=1.355
cc_5 VNB N_A_28_74#_M1003_g 0.0282514f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.545
cc_6 VNB N_A_28_74#_M1000_g 0.0395872f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_7 VNB N_A_28_74#_c_101_n 0.0226356f $X=-0.19 $Y=-0.245 $X2=0.57 $Y2=1.19
cc_8 VNB N_A_28_74#_c_102_n 0.0207876f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A_28_74#_c_103_n 0.0121635f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_28_74#_c_104_n 0.00140945f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_28_74#_c_105_n 0.0333044f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_289_74#_M1001_g 0.00313542f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.545
cc_13 VNB N_A_289_74#_M1005_g 0.0313942f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_289_74#_c_160_n 0.0147468f $X=-0.19 $Y=-0.245 $X2=0.57 $Y2=1.355
cc_15 VNB N_A_289_74#_c_161_n 0.020833f $X=-0.19 $Y=-0.245 $X2=0.57 $Y2=1.355
cc_16 VNB N_A_289_74#_c_162_n 0.0219379f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_289_74#_c_163_n 0.0575836f $X=-0.19 $Y=-0.245 $X2=0.415 $Y2=1.355
cc_18 VNB N_A_289_74#_c_164_n 0.00135856f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_289_74#_c_165_n 0.00336402f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_405_138#_M1006_g 0.0275176f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.545
cc_21 VNB N_A_405_138#_c_213_n 0.0358021f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_22 VNB N_A_405_138#_c_214_n 0.00382325f $X=-0.19 $Y=-0.245 $X2=0.57 $Y2=1.355
cc_23 VNB N_A_405_138#_c_215_n 0.00323188f $X=-0.19 $Y=-0.245 $X2=0.57 $Y2=1.52
cc_24 VNB N_A_405_138#_c_216_n 2.9305e-19 $X=-0.19 $Y=-0.245 $X2=0.415 $Y2=1.295
cc_25 VNB N_A_405_138#_c_217_n 0.00925722f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_VPWR_c_268_n 0.163682f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB X 0.0286532f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.545
cc_28 VNB N_X_c_301_n 0.029118f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB X 0.0145768f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_321_n 0.00984874f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.545
cc_31 VNB N_VGND_c_322_n 0.0187989f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_323_n 0.0567418f $X=-0.19 $Y=-0.245 $X2=0.57 $Y2=1.355
cc_33 VNB N_VGND_c_324_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0.57 $Y2=1.19
cc_34 VNB N_VGND_c_325_n 0.0180717f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_326_n 0.0205885f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_327_n 0.253699f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_328_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VPB N_A_c_64_n 0.0368635f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=2.17
cc_39 VPB N_A_c_68_n 0.0270096f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=2.26
cc_40 VPB A 0.0145994f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.21
cc_41 VPB N_A_28_74#_M1003_g 0.0637558f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=2.545
cc_42 VPB N_A_28_74#_c_107_n 0.0222081f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_43 VPB N_A_28_74#_c_108_n 0.00180999f $X=-0.19 $Y=1.66 $X2=0.415 $Y2=1.665
cc_44 VPB N_A_28_74#_c_109_n 0.0109668f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_45 VPB N_A_289_74#_M1001_g 0.0499439f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=2.545
cc_46 VPB N_A_289_74#_c_167_n 0.00516643f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_47 VPB N_A_289_74#_c_164_n 0.0129551f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_48 VPB N_A_405_138#_c_213_n 0.0265074f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_49 VPB N_A_405_138#_c_219_n 0.00175644f $X=-0.19 $Y=1.66 $X2=0.57 $Y2=1.355
cc_50 VPB N_A_405_138#_c_216_n 0.00160201f $X=-0.19 $Y=1.66 $X2=0.415 $Y2=1.295
cc_51 VPB N_A_405_138#_c_221_n 0.00745707f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_52 VPB N_VPWR_c_269_n 0.0183719f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=2.545
cc_53 VPB N_VPWR_c_270_n 0.0111617f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_54 VPB N_VPWR_c_271_n 0.0596029f $X=-0.19 $Y=1.66 $X2=0.57 $Y2=1.52
cc_55 VPB N_VPWR_c_272_n 0.00614127f $X=-0.19 $Y=1.66 $X2=0.415 $Y2=1.295
cc_56 VPB N_VPWR_c_273_n 0.018958f $X=-0.19 $Y=1.66 $X2=0.415 $Y2=1.355
cc_57 VPB N_VPWR_c_274_n 0.0200102f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_58 VPB N_VPWR_c_268_n 0.0940165f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_59 VPB N_VPWR_c_276_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_60 VPB X 0.00819691f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=2.545
cc_61 VPB X 0.0507685f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_62 VPB N_X_c_305_n 0.0146297f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_63 N_A_c_64_n N_A_28_74#_M1003_g 0.0251826f $X=0.495 $Y=2.17 $X2=0 $Y2=0
cc_64 N_A_c_68_n N_A_28_74#_M1003_g 0.012328f $X=0.495 $Y=2.26 $X2=0 $Y2=0
cc_65 A N_A_28_74#_M1003_g 0.00299941f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_66 N_A_M1004_g N_A_28_74#_M1000_g 0.00799939f $X=0.48 $Y=0.58 $X2=0 $Y2=0
cc_67 N_A_M1004_g N_A_28_74#_c_101_n 0.0127782f $X=0.48 $Y=0.58 $X2=0 $Y2=0
cc_68 N_A_c_68_n N_A_28_74#_c_107_n 0.00624408f $X=0.495 $Y=2.26 $X2=0 $Y2=0
cc_69 N_A_c_64_n N_A_28_74#_c_108_n 0.00956435f $X=0.495 $Y=2.17 $X2=0 $Y2=0
cc_70 N_A_c_68_n N_A_28_74#_c_108_n 0.00925083f $X=0.495 $Y=2.26 $X2=0 $Y2=0
cc_71 A N_A_28_74#_c_108_n 0.0262324f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_72 N_A_c_66_n N_A_28_74#_c_108_n 6.49888e-19 $X=0.57 $Y=1.355 $X2=0 $Y2=0
cc_73 A N_A_28_74#_c_109_n 0.0280303f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_74 N_A_M1004_g N_A_28_74#_c_102_n 0.012097f $X=0.48 $Y=0.58 $X2=0 $Y2=0
cc_75 A N_A_28_74#_c_102_n 0.0251751f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_76 N_A_c_66_n N_A_28_74#_c_102_n 0.00146766f $X=0.57 $Y=1.355 $X2=0 $Y2=0
cc_77 N_A_M1004_g N_A_28_74#_c_103_n 0.00415005f $X=0.48 $Y=0.58 $X2=0 $Y2=0
cc_78 A N_A_28_74#_c_103_n 0.0289843f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_79 N_A_M1004_g N_A_28_74#_c_104_n 0.00253208f $X=0.48 $Y=0.58 $X2=0 $Y2=0
cc_80 N_A_c_64_n N_A_28_74#_c_104_n 0.0013064f $X=0.495 $Y=2.17 $X2=0 $Y2=0
cc_81 A N_A_28_74#_c_104_n 0.0410413f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_82 N_A_c_66_n N_A_28_74#_c_104_n 0.00110237f $X=0.57 $Y=1.355 $X2=0 $Y2=0
cc_83 N_A_M1004_g N_A_28_74#_c_105_n 0.0021171f $X=0.48 $Y=0.58 $X2=0 $Y2=0
cc_84 A N_A_28_74#_c_105_n 0.00125289f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_85 N_A_c_66_n N_A_28_74#_c_105_n 0.0208561f $X=0.57 $Y=1.355 $X2=0 $Y2=0
cc_86 N_A_c_68_n N_VPWR_c_269_n 0.00399172f $X=0.495 $Y=2.26 $X2=0 $Y2=0
cc_87 N_A_c_68_n N_VPWR_c_273_n 0.00442668f $X=0.495 $Y=2.26 $X2=0 $Y2=0
cc_88 N_A_c_68_n N_VPWR_c_268_n 0.0048347f $X=0.495 $Y=2.26 $X2=0 $Y2=0
cc_89 N_A_M1004_g N_VGND_c_321_n 0.00294484f $X=0.48 $Y=0.58 $X2=0 $Y2=0
cc_90 N_A_M1004_g N_VGND_c_325_n 0.00456766f $X=0.48 $Y=0.58 $X2=0 $Y2=0
cc_91 N_A_M1004_g N_VGND_c_327_n 0.00456459f $X=0.48 $Y=0.58 $X2=0 $Y2=0
cc_92 N_A_28_74#_M1000_g N_A_289_74#_c_160_n 0.00977792f $X=1.355 $Y=0.58 $X2=0
+ $Y2=0
cc_93 N_A_28_74#_M1000_g N_A_289_74#_c_161_n 0.0149882f $X=1.355 $Y=0.58 $X2=0
+ $Y2=0
cc_94 N_A_28_74#_c_102_n N_A_289_74#_c_161_n 0.0164121f $X=0.975 $Y=0.92 $X2=0
+ $Y2=0
cc_95 N_A_28_74#_c_104_n N_A_289_74#_c_161_n 0.0277104f $X=1.14 $Y=1.295 $X2=0
+ $Y2=0
cc_96 N_A_28_74#_c_105_n N_A_289_74#_c_163_n 0.00415635f $X=1.14 $Y=1.295 $X2=0
+ $Y2=0
cc_97 N_A_28_74#_M1003_g N_A_289_74#_c_167_n 0.0102218f $X=1.195 $Y=2.46 $X2=0
+ $Y2=0
cc_98 N_A_28_74#_M1003_g N_A_289_74#_c_164_n 0.0203813f $X=1.195 $Y=2.46 $X2=0
+ $Y2=0
cc_99 N_A_28_74#_c_104_n N_A_289_74#_c_164_n 0.0295618f $X=1.14 $Y=1.295 $X2=0
+ $Y2=0
cc_100 N_A_28_74#_M1003_g N_A_289_74#_c_165_n 0.00351799f $X=1.195 $Y=2.46 $X2=0
+ $Y2=0
cc_101 N_A_28_74#_c_104_n N_A_289_74#_c_165_n 0.0193558f $X=1.14 $Y=1.295 $X2=0
+ $Y2=0
cc_102 N_A_28_74#_c_108_n N_VPWR_M1007_d 0.00835292f $X=0.975 $Y=2.117 $X2=-0.19
+ $Y2=-0.245
cc_103 N_A_28_74#_M1003_g N_VPWR_c_269_n 0.0119144f $X=1.195 $Y=2.46 $X2=0 $Y2=0
cc_104 N_A_28_74#_c_108_n N_VPWR_c_269_n 0.0227744f $X=0.975 $Y=2.117 $X2=0
+ $Y2=0
cc_105 N_A_28_74#_M1003_g N_VPWR_c_271_n 0.0151141f $X=1.195 $Y=2.46 $X2=0 $Y2=0
cc_106 N_A_28_74#_c_107_n N_VPWR_c_273_n 0.00593336f $X=0.265 $Y=2.56 $X2=0
+ $Y2=0
cc_107 N_A_28_74#_M1003_g N_VPWR_c_268_n 0.0292865f $X=1.195 $Y=2.46 $X2=0 $Y2=0
cc_108 N_A_28_74#_c_107_n N_VPWR_c_268_n 0.00940928f $X=0.265 $Y=2.56 $X2=0
+ $Y2=0
cc_109 N_A_28_74#_M1000_g N_VGND_c_321_n 0.00494615f $X=1.355 $Y=0.58 $X2=0
+ $Y2=0
cc_110 N_A_28_74#_c_101_n N_VGND_c_321_n 0.0151665f $X=0.265 $Y=0.58 $X2=0 $Y2=0
cc_111 N_A_28_74#_c_102_n N_VGND_c_321_n 0.0255952f $X=0.975 $Y=0.92 $X2=0 $Y2=0
cc_112 N_A_28_74#_M1000_g N_VGND_c_323_n 0.00518524f $X=1.355 $Y=0.58 $X2=0
+ $Y2=0
cc_113 N_A_28_74#_c_101_n N_VGND_c_325_n 0.0170785f $X=0.265 $Y=0.58 $X2=0 $Y2=0
cc_114 N_A_28_74#_M1000_g N_VGND_c_327_n 0.00867081f $X=1.355 $Y=0.58 $X2=0
+ $Y2=0
cc_115 N_A_28_74#_c_101_n N_VGND_c_327_n 0.0118627f $X=0.265 $Y=0.58 $X2=0 $Y2=0
cc_116 N_A_28_74#_c_102_n N_VGND_c_327_n 0.0214056f $X=0.975 $Y=0.92 $X2=0 $Y2=0
cc_117 N_A_289_74#_M1005_g N_A_405_138#_M1006_g 0.0198704f $X=2.695 $Y=0.9 $X2=0
+ $Y2=0
cc_118 N_A_289_74#_M1001_g N_A_405_138#_c_213_n 0.0313737f $X=2.535 $Y=2.34
+ $X2=0 $Y2=0
cc_119 N_A_289_74#_M1005_g N_A_405_138#_c_213_n 2.62551e-19 $X=2.695 $Y=0.9
+ $X2=0 $Y2=0
cc_120 N_A_289_74#_c_162_n N_A_405_138#_c_213_n 2.17534e-19 $X=2.575 $Y=1.465
+ $X2=0 $Y2=0
cc_121 N_A_289_74#_c_163_n N_A_405_138#_c_213_n 0.0215648f $X=2.575 $Y=1.465
+ $X2=0 $Y2=0
cc_122 N_A_289_74#_M1005_g N_A_405_138#_c_214_n 0.0189992f $X=2.695 $Y=0.9 $X2=0
+ $Y2=0
cc_123 N_A_289_74#_c_162_n N_A_405_138#_c_214_n 0.0283815f $X=2.575 $Y=1.465
+ $X2=0 $Y2=0
cc_124 N_A_289_74#_c_163_n N_A_405_138#_c_214_n 0.00767481f $X=2.575 $Y=1.465
+ $X2=0 $Y2=0
cc_125 N_A_289_74#_M1001_g N_A_405_138#_c_219_n 0.0366973f $X=2.535 $Y=2.34
+ $X2=0 $Y2=0
cc_126 N_A_289_74#_c_162_n N_A_405_138#_c_219_n 0.0227169f $X=2.575 $Y=1.465
+ $X2=0 $Y2=0
cc_127 N_A_289_74#_M1005_g N_A_405_138#_c_215_n 0.00219888f $X=2.695 $Y=0.9
+ $X2=0 $Y2=0
cc_128 N_A_289_74#_c_162_n N_A_405_138#_c_215_n 0.0193923f $X=2.575 $Y=1.465
+ $X2=0 $Y2=0
cc_129 N_A_289_74#_c_163_n N_A_405_138#_c_215_n 0.00410963f $X=2.575 $Y=1.465
+ $X2=0 $Y2=0
cc_130 N_A_289_74#_M1001_g N_A_405_138#_c_216_n 0.00496065f $X=2.535 $Y=2.34
+ $X2=0 $Y2=0
cc_131 N_A_289_74#_M1005_g N_A_405_138#_c_217_n 0.0100145f $X=2.695 $Y=0.9 $X2=0
+ $Y2=0
cc_132 N_A_289_74#_c_161_n N_A_405_138#_c_217_n 0.0301033f $X=1.597 $Y=1.38
+ $X2=0 $Y2=0
cc_133 N_A_289_74#_c_162_n N_A_405_138#_c_217_n 0.0290383f $X=2.575 $Y=1.465
+ $X2=0 $Y2=0
cc_134 N_A_289_74#_c_163_n N_A_405_138#_c_217_n 0.00721063f $X=2.575 $Y=1.465
+ $X2=0 $Y2=0
cc_135 N_A_289_74#_M1001_g N_A_405_138#_c_221_n 0.0147779f $X=2.535 $Y=2.34
+ $X2=0 $Y2=0
cc_136 N_A_289_74#_c_162_n N_A_405_138#_c_221_n 0.0235446f $X=2.575 $Y=1.465
+ $X2=0 $Y2=0
cc_137 N_A_289_74#_c_163_n N_A_405_138#_c_221_n 0.00490082f $X=2.575 $Y=1.465
+ $X2=0 $Y2=0
cc_138 N_A_289_74#_c_164_n N_A_405_138#_c_221_n 0.021975f $X=1.567 $Y=2.395
+ $X2=0 $Y2=0
cc_139 N_A_289_74#_M1001_g N_VPWR_c_270_n 0.00865052f $X=2.535 $Y=2.34 $X2=0
+ $Y2=0
cc_140 N_A_289_74#_M1001_g N_VPWR_c_271_n 0.0164683f $X=2.535 $Y=2.34 $X2=0
+ $Y2=0
cc_141 N_A_289_74#_c_167_n N_VPWR_c_271_n 0.00561205f $X=1.58 $Y=2.56 $X2=0
+ $Y2=0
cc_142 N_A_289_74#_M1001_g N_VPWR_c_268_n 0.016946f $X=2.535 $Y=2.34 $X2=0 $Y2=0
cc_143 N_A_289_74#_c_167_n N_VPWR_c_268_n 0.00918412f $X=1.58 $Y=2.56 $X2=0
+ $Y2=0
cc_144 N_A_289_74#_c_160_n N_VGND_c_321_n 0.0111541f $X=1.597 $Y=0.635 $X2=0
+ $Y2=0
cc_145 N_A_289_74#_M1005_g N_VGND_c_322_n 0.00468436f $X=2.695 $Y=0.9 $X2=0
+ $Y2=0
cc_146 N_A_289_74#_M1005_g N_VGND_c_323_n 0.00459186f $X=2.695 $Y=0.9 $X2=0
+ $Y2=0
cc_147 N_A_289_74#_c_160_n N_VGND_c_323_n 0.0163385f $X=1.597 $Y=0.635 $X2=0
+ $Y2=0
cc_148 N_A_289_74#_M1005_g N_VGND_c_327_n 0.00542201f $X=2.695 $Y=0.9 $X2=0
+ $Y2=0
cc_149 N_A_289_74#_c_160_n N_VGND_c_327_n 0.0113715f $X=1.597 $Y=0.635 $X2=0
+ $Y2=0
cc_150 N_A_405_138#_c_219_n N_VPWR_M1001_d 0.00262668f $X=2.91 $Y=1.91 $X2=0
+ $Y2=0
cc_151 N_A_405_138#_c_213_n N_VPWR_c_270_n 0.0153694f $X=3.215 $Y=1.765 $X2=0
+ $Y2=0
cc_152 N_A_405_138#_c_219_n N_VPWR_c_270_n 0.0222367f $X=2.91 $Y=1.91 $X2=0
+ $Y2=0
cc_153 N_A_405_138#_c_213_n N_VPWR_c_274_n 0.00413917f $X=3.215 $Y=1.765 $X2=0
+ $Y2=0
cc_154 N_A_405_138#_c_213_n N_VPWR_c_268_n 0.00821556f $X=3.215 $Y=1.765 $X2=0
+ $Y2=0
cc_155 N_A_405_138#_M1006_g X 0.00260428f $X=3.205 $Y=0.74 $X2=0 $Y2=0
cc_156 N_A_405_138#_c_213_n X 0.0110819f $X=3.215 $Y=1.765 $X2=0 $Y2=0
cc_157 N_A_405_138#_c_215_n X 0.0327059f $X=3.032 $Y=1.625 $X2=0 $Y2=0
cc_158 N_A_405_138#_c_216_n X 0.00709928f $X=3.032 $Y=1.825 $X2=0 $Y2=0
cc_159 N_A_405_138#_M1006_g N_X_c_301_n 0.00143568f $X=3.205 $Y=0.74 $X2=0 $Y2=0
cc_160 N_A_405_138#_c_215_n X 0.0037592f $X=3.032 $Y=1.625 $X2=0 $Y2=0
cc_161 N_A_405_138#_c_213_n N_X_c_305_n 0.00396238f $X=3.215 $Y=1.765 $X2=0
+ $Y2=0
cc_162 N_A_405_138#_c_219_n N_X_c_305_n 0.00776663f $X=2.91 $Y=1.91 $X2=0 $Y2=0
cc_163 N_A_405_138#_c_216_n N_X_c_305_n 7.53348e-19 $X=3.032 $Y=1.825 $X2=0
+ $Y2=0
cc_164 N_A_405_138#_c_214_n N_VGND_M1005_d 7.12223e-19 $X=2.91 $Y=1.125 $X2=0
+ $Y2=0
cc_165 N_A_405_138#_c_215_n N_VGND_M1005_d 0.0018038f $X=3.032 $Y=1.625 $X2=0
+ $Y2=0
cc_166 N_A_405_138#_M1006_g N_VGND_c_322_n 0.0156117f $X=3.205 $Y=0.74 $X2=0
+ $Y2=0
cc_167 N_A_405_138#_c_213_n N_VGND_c_322_n 4.77198e-19 $X=3.215 $Y=1.765 $X2=0
+ $Y2=0
cc_168 N_A_405_138#_c_214_n N_VGND_c_322_n 0.00549591f $X=2.91 $Y=1.125 $X2=0
+ $Y2=0
cc_169 N_A_405_138#_c_215_n N_VGND_c_322_n 0.016728f $X=3.032 $Y=1.625 $X2=0
+ $Y2=0
cc_170 N_A_405_138#_c_217_n N_VGND_c_323_n 0.00580898f $X=2.15 $Y=0.875 $X2=0
+ $Y2=0
cc_171 N_A_405_138#_M1006_g N_VGND_c_326_n 0.00383152f $X=3.205 $Y=0.74 $X2=0
+ $Y2=0
cc_172 N_A_405_138#_M1006_g N_VGND_c_327_n 0.00761589f $X=3.205 $Y=0.74 $X2=0
+ $Y2=0
cc_173 N_A_405_138#_c_217_n N_VGND_c_327_n 0.0101265f $X=2.15 $Y=0.875 $X2=0
+ $Y2=0
cc_174 N_VPWR_c_270_n X 0.0378466f $X=2.99 $Y=2.27 $X2=0 $Y2=0
cc_175 N_VPWR_c_274_n X 0.0270407f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_176 N_VPWR_c_268_n X 0.0159412f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_177 N_X_c_301_n N_VGND_c_322_n 0.019927f $X=3.42 $Y=0.52 $X2=0 $Y2=0
cc_178 N_X_c_301_n N_VGND_c_326_n 0.0180659f $X=3.42 $Y=0.52 $X2=0 $Y2=0
cc_179 N_X_c_301_n N_VGND_c_327_n 0.0152075f $X=3.42 $Y=0.52 $X2=0 $Y2=0
