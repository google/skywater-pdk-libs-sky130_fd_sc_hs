# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_sc_hs__dfxtp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__dfxtp_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  8.160000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.870000 2.025000 2.250000 2.355000 ;
        RECT 1.970000 1.125000 2.250000 2.025000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.541300 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.715000 0.350000 8.075000 1.130000 ;
        RECT 7.715000 2.030000 8.075000 2.980000 ;
        RECT 7.905000 1.130000 8.075000 2.030000 ;
    END
  END Q
  PIN CLK
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.300000 0.505000 1.780000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 8.160000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.000000 0.000000 8.160000 0.245000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.660000 8.350000 3.520000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 8.160000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 8.160000 0.085000 ;
      RECT 0.000000  3.245000 8.160000 3.415000 ;
      RECT 0.115000  0.350000 0.365000 0.960000 ;
      RECT 0.115000  0.960000 1.135000 1.130000 ;
      RECT 0.115000  1.950000 0.845000 2.120000 ;
      RECT 0.115000  2.120000 0.445000 2.980000 ;
      RECT 0.545000  0.085000 0.795000 0.790000 ;
      RECT 0.645000  2.290000 0.815000 3.245000 ;
      RECT 0.675000  1.130000 1.135000 1.550000 ;
      RECT 0.675000  1.550000 0.845000 1.950000 ;
      RECT 0.965000  0.255000 1.815000 0.425000 ;
      RECT 0.965000  0.425000 1.135000 0.960000 ;
      RECT 1.015000  1.820000 1.475000 2.625000 ;
      RECT 1.015000  2.625000 2.250000 2.795000 ;
      RECT 1.015000  2.795000 1.345000 2.980000 ;
      RECT 1.305000  0.595000 1.475000 1.350000 ;
      RECT 1.305000  1.350000 1.760000 1.680000 ;
      RECT 1.305000  1.680000 1.475000 1.820000 ;
      RECT 1.575000  2.965000 1.910000 3.245000 ;
      RECT 1.645000  0.425000 1.815000 0.730000 ;
      RECT 1.645000  0.730000 2.655000 0.900000 ;
      RECT 1.985000  0.085000 2.315000 0.560000 ;
      RECT 2.080000  2.795000 3.460000 2.965000 ;
      RECT 2.420000  1.070000 2.975000 1.240000 ;
      RECT 2.420000  1.240000 2.590000 2.625000 ;
      RECT 2.485000  0.275000 3.760000 0.445000 ;
      RECT 2.485000  0.445000 2.655000 0.730000 ;
      RECT 2.760000  1.410000 3.420000 1.580000 ;
      RECT 2.760000  1.580000 2.930000 2.285000 ;
      RECT 2.760000  2.285000 4.140000 2.455000 ;
      RECT 2.760000  2.455000 3.120000 2.625000 ;
      RECT 3.100000  1.750000 3.760000 2.080000 ;
      RECT 3.155000  0.615000 3.420000 1.410000 ;
      RECT 3.290000  2.625000 4.950000 2.795000 ;
      RECT 3.590000  0.445000 3.760000 0.690000 ;
      RECT 3.590000  0.690000 4.660000 0.860000 ;
      RECT 3.590000  0.860000 3.760000 1.750000 ;
      RECT 3.800000  2.965000 4.130000 3.245000 ;
      RECT 3.930000  1.030000 5.000000 1.200000 ;
      RECT 3.930000  1.200000 4.260000 1.415000 ;
      RECT 3.970000  1.625000 4.270000 1.955000 ;
      RECT 3.970000  1.955000 4.140000 2.285000 ;
      RECT 4.070000  0.085000 4.320000 0.520000 ;
      RECT 4.335000  2.125000 4.610000 2.455000 ;
      RECT 4.440000  1.200000 4.610000 2.125000 ;
      RECT 4.490000  0.255000 5.895000 0.425000 ;
      RECT 4.490000  0.425000 4.660000 0.690000 ;
      RECT 4.780000  1.370000 5.480000 1.540000 ;
      RECT 4.780000  1.540000 4.950000 2.625000 ;
      RECT 4.780000  2.795000 4.950000 2.905000 ;
      RECT 4.780000  2.905000 5.840000 3.075000 ;
      RECT 4.830000  0.595000 5.000000 1.030000 ;
      RECT 5.120000  1.710000 5.820000 1.880000 ;
      RECT 5.120000  1.880000 5.290000 2.735000 ;
      RECT 5.170000  1.150000 5.480000 1.370000 ;
      RECT 5.220000  0.730000 5.820000 0.980000 ;
      RECT 5.510000  2.050000 5.840000 2.905000 ;
      RECT 5.565000  0.425000 5.895000 0.510000 ;
      RECT 5.650000  0.980000 5.820000 1.230000 ;
      RECT 5.650000  1.230000 7.205000 1.400000 ;
      RECT 5.650000  1.400000 5.820000 1.710000 ;
      RECT 6.050000  1.570000 6.380000 1.690000 ;
      RECT 6.050000  1.690000 7.735000 1.860000 ;
      RECT 6.050000  1.860000 6.380000 2.240000 ;
      RECT 6.200000  2.520000 6.530000 3.245000 ;
      RECT 6.230000  0.085000 6.560000 1.060000 ;
      RECT 6.760000  1.860000 7.010000 2.700000 ;
      RECT 6.790000  0.350000 7.040000 0.850000 ;
      RECT 6.790000  0.850000 7.545000 1.020000 ;
      RECT 6.875000  1.190000 7.205000 1.230000 ;
      RECT 6.875000  1.400000 7.205000 1.520000 ;
      RECT 7.210000  2.030000 7.540000 3.245000 ;
      RECT 7.220000  0.085000 7.535000 0.680000 ;
      RECT 7.375000  1.020000 7.545000 1.350000 ;
      RECT 7.375000  1.350000 7.735000 1.690000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
      RECT 7.835000 -0.085000 8.005000 0.085000 ;
      RECT 7.835000  3.245000 8.005000 3.415000 ;
  END
END sky130_fd_sc_hs__dfxtp_1
END LIBRARY
