* File: sky130_fd_sc_hs__a221oi_1.pex.spice
* Created: Tue Sep  1 19:50:25 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HS__A221OI_1%C1 1 3 6 8 12 13
c27 13 0 1.63146e-19 $X=0.71 $Y=1.515
c28 1 0 5.89647e-20 $X=0.515 $Y=1.765
r29 12 14 60.9588 $w=3.4e-07 $l=4.3e-07 $layer=POLY_cond $X=0.71 $Y=1.557
+ $X2=1.14 $Y2=1.557
r30 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.71
+ $Y=1.515 $X2=0.71 $Y2=1.515
r31 10 12 27.6441 $w=3.4e-07 $l=1.95e-07 $layer=POLY_cond $X=0.515 $Y=1.557
+ $X2=0.71 $Y2=1.557
r32 8 13 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=0.71 $Y=1.665
+ $X2=0.71 $Y2=1.515
r33 4 14 21.9347 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.14 $Y=1.35
+ $X2=1.14 $Y2=1.557
r34 4 6 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.14 $Y=1.35 $X2=1.14
+ $Y2=0.74
r35 1 10 21.9347 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=0.515 $Y=1.765
+ $X2=0.515 $Y2=1.557
r36 1 3 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.515 $Y=1.765
+ $X2=0.515 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_HS__A221OI_1%B2 1 3 6 8 9
c30 9 0 5.89647e-20 $X=1.68 $Y=1.665
c31 1 0 1.63146e-19 $X=1.665 $Y=1.765
r32 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.59
+ $Y=1.515 $X2=1.59 $Y2=1.515
r33 9 14 2.41209 $w=4.28e-07 $l=9e-08 $layer=LI1_cond $X=1.68 $Y=1.565 $X2=1.59
+ $Y2=1.565
r34 8 14 10.4524 $w=4.28e-07 $l=3.9e-07 $layer=LI1_cond $X=1.2 $Y=1.565 $X2=1.59
+ $Y2=1.565
r35 4 13 38.5562 $w=2.99e-07 $l=2.05122e-07 $layer=POLY_cond $X=1.68 $Y=1.35
+ $X2=1.59 $Y2=1.515
r36 4 6 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.68 $Y=1.35 $X2=1.68
+ $Y2=0.74
r37 1 13 52.2586 $w=2.99e-07 $l=2.85044e-07 $layer=POLY_cond $X=1.665 $Y=1.765
+ $X2=1.59 $Y2=1.515
r38 1 3 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.665 $Y=1.765
+ $X2=1.665 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_HS__A221OI_1%B1 3 5 7 8 12
r31 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.13
+ $Y=1.515 $X2=2.13 $Y2=1.515
r32 8 12 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=2.13 $Y=1.665
+ $X2=2.13 $Y2=1.515
r33 5 11 52.2586 $w=2.99e-07 $l=2.57391e-07 $layer=POLY_cond $X=2.115 $Y=1.765
+ $X2=2.13 $Y2=1.515
r34 5 7 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.115 $Y=1.765
+ $X2=2.115 $Y2=2.4
r35 1 11 38.5562 $w=2.99e-07 $l=2.05122e-07 $layer=POLY_cond $X=2.04 $Y=1.35
+ $X2=2.13 $Y2=1.515
r36 1 3 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.04 $Y=1.35 $X2=2.04
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HS__A221OI_1%A1 1 3 6 8 12
r31 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.67
+ $Y=1.515 $X2=2.67 $Y2=1.515
r32 8 12 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=2.67 $Y=1.665
+ $X2=2.67 $Y2=1.515
r33 4 11 38.5562 $w=2.99e-07 $l=2.05122e-07 $layer=POLY_cond $X=2.76 $Y=1.35
+ $X2=2.67 $Y2=1.515
r34 4 6 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.76 $Y=1.35 $X2=2.76
+ $Y2=0.74
r35 1 11 52.2586 $w=2.99e-07 $l=2.85044e-07 $layer=POLY_cond $X=2.595 $Y=1.765
+ $X2=2.67 $Y2=1.515
r36 1 3 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.595 $Y=1.765
+ $X2=2.595 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_HS__A221OI_1%A2 1 3 4 6 7 8
r22 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.21
+ $Y=1.385 $X2=3.21 $Y2=1.385
r23 8 13 12.1474 $w=3.68e-07 $l=3.9e-07 $layer=LI1_cond $X=3.6 $Y=1.365 $X2=3.21
+ $Y2=1.365
r24 7 13 2.80324 $w=3.68e-07 $l=9e-08 $layer=LI1_cond $X=3.12 $Y=1.365 $X2=3.21
+ $Y2=1.365
r25 4 12 77.2841 $w=2.7e-07 $l=4.15812e-07 $layer=POLY_cond $X=3.135 $Y=1.765
+ $X2=3.21 $Y2=1.385
r26 4 6 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.135 $Y=1.765
+ $X2=3.135 $Y2=2.4
r27 1 12 38.9026 $w=2.7e-07 $l=2.05122e-07 $layer=POLY_cond $X=3.12 $Y=1.22
+ $X2=3.21 $Y2=1.385
r28 1 3 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=3.12 $Y=1.22 $X2=3.12
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HS__A221OI_1%Y 1 2 3 10 14 16 18 19 20 21 22 51
r39 50 51 11.617 $w=8.28e-07 $l=1.65e-07 $layer=LI1_cond $X=0.925 $Y=0.765
+ $X2=1.09 $Y2=0.765
r40 48 50 9.72714 $w=8.28e-07 $l=6.75e-07 $layer=LI1_cond $X=0.25 $Y=0.765
+ $X2=0.925 $Y2=0.765
r41 30 48 7.92413 $w=2.5e-07 $l=4.15e-07 $layer=LI1_cond $X=0.25 $Y=1.18
+ $X2=0.25 $Y2=0.765
r42 21 22 17.0562 $w=2.48e-07 $l=3.7e-07 $layer=LI1_cond $X=0.25 $Y=2.405
+ $X2=0.25 $Y2=2.775
r43 20 21 19.361 $w=2.48e-07 $l=4.2e-07 $layer=LI1_cond $X=0.25 $Y=1.985
+ $X2=0.25 $Y2=2.405
r44 19 20 14.7513 $w=2.48e-07 $l=3.2e-07 $layer=LI1_cond $X=0.25 $Y=1.665
+ $X2=0.25 $Y2=1.985
r45 18 19 17.0562 $w=2.48e-07 $l=3.7e-07 $layer=LI1_cond $X=0.25 $Y=1.295
+ $X2=0.25 $Y2=1.665
r46 18 30 5.30124 $w=2.48e-07 $l=1.15e-07 $layer=LI1_cond $X=0.25 $Y=1.295
+ $X2=0.25 $Y2=1.18
r47 16 48 0.144106 $w=8.28e-07 $l=1e-08 $layer=LI1_cond $X=0.24 $Y=0.765
+ $X2=0.25 $Y2=0.765
r48 12 14 14.3014 $w=4.13e-07 $l=5.15e-07 $layer=LI1_cond $X=2.367 $Y=1.01
+ $X2=2.367 $Y2=0.495
r49 10 12 8.50155 $w=1.7e-07 $l=2.45854e-07 $layer=LI1_cond $X=2.16 $Y=1.095
+ $X2=2.367 $Y2=1.01
r50 10 51 69.8075 $w=1.68e-07 $l=1.07e-06 $layer=LI1_cond $X=2.16 $Y=1.095
+ $X2=1.09 $Y2=1.095
r51 3 22 400 $w=1.7e-07 $l=1.03562e-06 $layer=licon1_PDIFF $count=1 $X=0.165
+ $Y=1.84 $X2=0.29 $Y2=2.815
r52 3 20 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.165
+ $Y=1.84 $X2=0.29 $Y2=1.985
r53 2 14 91 $w=1.7e-07 $l=3.16386e-07 $layer=licon1_NDIFF $count=2 $X=2.115
+ $Y=0.37 $X2=2.375 $Y2=0.495
r54 1 50 45.5 $w=1.7e-07 $l=5.32588e-07 $layer=licon1_NDIFF $count=4 $X=0.46
+ $Y=0.37 $X2=0.925 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__A221OI_1%A_118_368# 1 2 9 13 14 17
r28 15 17 17.6359 $w=3.28e-07 $l=5.05e-07 $layer=LI1_cond $X=1.89 $Y=2.905
+ $X2=1.89 $Y2=2.4
r29 13 15 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.725 $Y=2.99
+ $X2=1.89 $Y2=2.905
r30 13 14 53.4973 $w=1.68e-07 $l=8.2e-07 $layer=LI1_cond $X=1.725 $Y=2.99
+ $X2=0.905 $Y2=2.99
r31 9 12 24.4458 $w=3.28e-07 $l=7e-07 $layer=LI1_cond $X=0.74 $Y=2.115 $X2=0.74
+ $Y2=2.815
r32 7 14 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.74 $Y=2.905
+ $X2=0.905 $Y2=2.99
r33 7 12 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=0.74 $Y=2.905 $X2=0.74
+ $Y2=2.815
r34 2 17 300 $w=1.7e-07 $l=6.30555e-07 $layer=licon1_PDIFF $count=2 $X=1.74
+ $Y=1.84 $X2=1.89 $Y2=2.4
r35 1 12 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=0.59
+ $Y=1.84 $X2=0.74 $Y2=2.815
r36 1 9 400 $w=1.7e-07 $l=3.4187e-07 $layer=licon1_PDIFF $count=1 $X=0.59
+ $Y=1.84 $X2=0.74 $Y2=2.115
.ends

.subckt PM_SKY130_FD_SC_HS__A221OI_1%A_263_368# 1 2 3 10 12 14 18 20 22 24 29
r40 22 31 3.0656 $w=3.3e-07 $l=1.5e-07 $layer=LI1_cond $X=3.36 $Y=2.12 $X2=3.36
+ $Y2=1.97
r41 22 24 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=3.36 $Y=2.12
+ $X2=3.36 $Y2=2.815
r42 21 29 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.505 $Y=2.035
+ $X2=2.38 $Y2=2.035
r43 20 31 4.70058 $w=1.7e-07 $l=1.94808e-07 $layer=LI1_cond $X=3.195 $Y=2.035
+ $X2=3.36 $Y2=1.97
r44 20 21 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=3.195 $Y=2.035
+ $X2=2.505 $Y2=2.035
r45 16 29 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.38 $Y=2.12
+ $X2=2.38 $Y2=2.035
r46 16 18 14.7513 $w=2.48e-07 $l=3.2e-07 $layer=LI1_cond $X=2.38 $Y=2.12
+ $X2=2.38 $Y2=2.44
r47 15 27 4.47015 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=1.545 $Y=2.035
+ $X2=1.41 $Y2=2.035
r48 14 29 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.255 $Y=2.035
+ $X2=2.38 $Y2=2.035
r49 14 15 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=2.255 $Y=2.035
+ $X2=1.545 $Y2=2.035
r50 10 27 2.81454 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.41 $Y=2.12 $X2=1.41
+ $Y2=2.035
r51 10 12 19.2074 $w=2.68e-07 $l=4.5e-07 $layer=LI1_cond $X=1.41 $Y=2.12
+ $X2=1.41 $Y2=2.57
r52 3 31 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=3.21
+ $Y=1.84 $X2=3.36 $Y2=1.985
r53 3 24 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=3.21
+ $Y=1.84 $X2=3.36 $Y2=2.815
r54 2 29 600 $w=1.7e-07 $l=2.59374e-07 $layer=licon1_PDIFF $count=1 $X=2.19
+ $Y=1.84 $X2=2.34 $Y2=2.035
r55 2 18 300 $w=1.7e-07 $l=6.7082e-07 $layer=licon1_PDIFF $count=2 $X=2.19
+ $Y=1.84 $X2=2.34 $Y2=2.44
r56 1 27 600 $w=1.7e-07 $l=2.498e-07 $layer=licon1_PDIFF $count=1 $X=1.315
+ $Y=1.84 $X2=1.44 $Y2=2.035
r57 1 12 600 $w=1.7e-07 $l=7.90032e-07 $layer=licon1_PDIFF $count=1 $X=1.315
+ $Y=1.84 $X2=1.44 $Y2=2.57
.ends

.subckt PM_SKY130_FD_SC_HS__A221OI_1%VPWR 1 6 9 10 11 21 22
r33 21 22 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r34 19 22 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.6 $Y2=3.33
r35 18 19 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r36 14 18 156.578 $w=1.68e-07 $l=2.4e-06 $layer=LI1_cond $X=0.24 $Y=3.33
+ $X2=2.64 $Y2=3.33
r37 14 15 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r38 11 19 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=2.64 $Y2=3.33
r39 11 15 0.468274 $w=4.9e-07 $l=1.68e-06 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=0.24 $Y2=3.33
r40 9 18 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=2.675 $Y=3.33
+ $X2=2.64 $Y2=3.33
r41 9 10 8.9695 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=2.675 $Y=3.33 $X2=2.85
+ $Y2=3.33
r42 8 21 37.5134 $w=1.68e-07 $l=5.75e-07 $layer=LI1_cond $X=3.025 $Y=3.33
+ $X2=3.6 $Y2=3.33
r43 8 10 8.9695 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=3.025 $Y=3.33 $X2=2.85
+ $Y2=3.33
r44 4 10 1.07557 $w=3.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.85 $Y=3.245 $X2=2.85
+ $Y2=3.33
r45 4 6 27.8233 $w=3.48e-07 $l=8.45e-07 $layer=LI1_cond $X=2.85 $Y=3.245
+ $X2=2.85 $Y2=2.4
r46 1 6 300 $w=1.7e-07 $l=6.43739e-07 $layer=licon1_PDIFF $count=2 $X=2.67
+ $Y=1.84 $X2=2.85 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_HS__A221OI_1%VGND 1 2 9 13 16 17 19 20 21 37 38
r34 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r35 35 38 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=3.6
+ $Y2=0
r36 34 35 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r37 31 34 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.68 $Y=0 $X2=3.12
+ $Y2=0
r38 31 32 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r39 29 32 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=1.68
+ $Y2=0
r40 28 29 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r41 25 29 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=1.2
+ $Y2=0
r42 24 28 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.24 $Y=0 $X2=1.2
+ $Y2=0
r43 24 25 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r44 21 35 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=1.92 $Y=0 $X2=3.12
+ $Y2=0
r45 21 32 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=1.68
+ $Y2=0
r46 19 34 3.26203 $w=1.68e-07 $l=5e-08 $layer=LI1_cond $X=3.17 $Y=0 $X2=3.12
+ $Y2=0
r47 19 20 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.17 $Y=0 $X2=3.335
+ $Y2=0
r48 18 37 6.52406 $w=1.68e-07 $l=1e-07 $layer=LI1_cond $X=3.5 $Y=0 $X2=3.6 $Y2=0
r49 18 20 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.5 $Y=0 $X2=3.335
+ $Y2=0
r50 16 28 3.91444 $w=1.68e-07 $l=6e-08 $layer=LI1_cond $X=1.26 $Y=0 $X2=1.2
+ $Y2=0
r51 16 17 9.31531 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=1.26 $Y=0 $X2=1.445
+ $Y2=0
r52 15 31 3.26203 $w=1.68e-07 $l=5e-08 $layer=LI1_cond $X=1.63 $Y=0 $X2=1.68
+ $Y2=0
r53 15 17 9.31531 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=1.63 $Y=0 $X2=1.445
+ $Y2=0
r54 11 20 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.335 $Y=0.085
+ $X2=3.335 $Y2=0
r55 11 13 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=3.335 $Y=0.085
+ $X2=3.335 $Y2=0.515
r56 7 17 1.24149 $w=3.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.445 $Y=0.085
+ $X2=1.445 $Y2=0
r57 7 9 18.3768 $w=3.68e-07 $l=5.9e-07 $layer=LI1_cond $X=1.445 $Y=0.085
+ $X2=1.445 $Y2=0.675
r58 2 13 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.195
+ $Y=0.37 $X2=3.335 $Y2=0.515
r59 1 9 182 $w=1.7e-07 $l=4.03949e-07 $layer=licon1_NDIFF $count=1 $X=1.215
+ $Y=0.37 $X2=1.445 $Y2=0.675
.ends

