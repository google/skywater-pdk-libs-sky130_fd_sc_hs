* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hs__nand3b_4 A_N B C VGND VNB VPB VPWR Y
M1000 VGND A_N a_89_172# VNB nlowvt w=740000u l=150000u
+  ad=1.1492e+12p pd=8.02e+06u as=1.9515e+11p ps=2.05e+06u
M1001 a_744_74# B a_297_82# VNB nlowvt w=740000u l=150000u
+  ad=1.0672e+12p pd=1.036e+07u as=8.806e+11p ps=8.3e+06u
M1002 a_744_74# a_89_172# Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=4.329e+11p ps=4.13e+06u
M1003 a_89_172# A_N VPWR VPB pshort w=840000u l=150000u
+  ad=2.52e+11p pd=2.28e+06u as=4.9686e+12p ps=1.99e+07u
M1004 a_297_82# C VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_744_74# B a_297_82# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VPWR A_N a_89_172# VPB pshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 Y B VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=1.4336e+12p pd=9.28e+06u as=0p ps=0u
M1008 VPWR B Y VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VGND C a_297_82# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 Y C VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VGND C a_297_82# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VPWR C Y VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_297_82# C VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 VPWR a_89_172# Y VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 Y a_89_172# VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 Y a_89_172# a_744_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 Y a_89_172# a_744_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_297_82# B a_744_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_297_82# B a_744_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_744_74# a_89_172# Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
