* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hs__and2b_4 A_N B VGND VNB VPB VPWR X
M1000 VGND a_218_424# X VNB nlowvt w=740000u l=150000u
+  ad=9.074e+11p pd=8.29e+06u as=4.218e+11p ps=4.1e+06u
M1001 a_218_424# a_27_392# VPWR VPB pshort w=840000u l=150000u
+  ad=5.04e+11p pd=4.56e+06u as=1.7066e+12p ps=1.379e+07u
M1002 VPWR a_27_392# a_218_424# VPB pshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1003 VGND a_218_424# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 X a_218_424# VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=6.72e+11p pd=5.68e+06u as=0p ps=0u
M1005 a_218_424# a_27_392# a_233_74# VNB nlowvt w=640000u l=150000u
+  ad=1.792e+11p pd=1.84e+06u as=4.16e+11p ps=3.86e+06u
M1006 VPWR a_218_424# X VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_233_74# B VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_218_424# B VPWR VPB pshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 X a_218_424# VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VPWR B a_218_424# VPB pshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VGND A_N a_27_392# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=1.824e+11p ps=1.85e+06u
M1012 VPWR a_218_424# X VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 X a_218_424# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 X a_218_424# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_233_74# a_27_392# a_218_424# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VPWR A_N a_27_392# VPB pshort w=1e+06u l=150000u
+  ad=0p pd=0u as=2.85e+11p ps=2.57e+06u
M1017 VGND B a_233_74# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
