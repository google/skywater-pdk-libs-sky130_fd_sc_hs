* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hs__nor2b_4 A B_N VGND VNB VPB VPWR Y
X0 VPWR A a_116_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X1 a_353_323# B_N VPWR VPB sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X2 Y a_353_323# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X3 VPWR A a_116_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X4 Y a_353_323# a_116_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X5 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X6 Y a_353_323# a_116_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X7 VGND B_N a_353_323# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X8 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X9 VPWR B_N a_353_323# VPB sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X10 a_116_368# A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X11 a_116_368# A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X12 a_116_368# a_353_323# Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X13 a_116_368# a_353_323# Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X14 VGND a_353_323# Y VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
.ends
