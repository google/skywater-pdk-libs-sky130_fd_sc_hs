* File: sky130_fd_sc_hs__a21boi_2.spice
* Created: Tue Sep  1 19:49:22 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hs__a21boi_2.pex.spice"
.subckt sky130_fd_sc_hs__a21boi_2  VNB VPB B1_N A1 A2 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A2	A2
* A1	A1
* B1_N	B1_N
* VPB	VPB
* VNB	VNB
MM1002 N_VGND_M1002_d N_B1_N_M1002_g N_A_62_94#_M1002_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.113206 AS=0.1696 PD=1.00174 PS=1.81 NRD=11.712 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75001.1 A=0.096 P=1.58 MULT=1
MM1003 N_Y_M1003_d N_A_62_94#_M1003_g N_VGND_M1002_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.130894 PD=1.02 PS=1.15826 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.6
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1009 N_Y_M1003_d N_A_62_94#_M1009_g N_VGND_M1009_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1961 PD=1.02 PS=2.01 NRD=0 NRS=0 M=1 R=4.93333 SA=75001
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1000 N_A_436_74#_M1000_d N_A1_M1000_g N_Y_M1000_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1961 AS=0.1036 PD=2.01 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75001.5 A=0.111 P=1.78 MULT=1
MM1011 N_A_436_74#_M1011_d N_A1_M1011_g N_Y_M1000_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.6
+ SB=75001.1 A=0.111 P=1.78 MULT=1
MM1004 N_VGND_M1004_d N_A2_M1004_g N_A_436_74#_M1011_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.1
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1013 N_VGND_M1004_d N_A2_M1013_g N_A_436_74#_M1013_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1961 PD=1.02 PS=2.01 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.5
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1012 N_A_62_94#_M1012_d N_B1_N_M1012_g N_VPWR_M1012_s VPB PSHORT L=0.15 W=1
+ AD=0.275 AS=0.275 PD=2.55 PS=2.55 NRD=1.9503 NRS=1.9503 M=1 R=6.66667
+ SA=75000.2 SB=75000.2 A=0.15 P=2.3 MULT=1
MM1005 N_Y_M1005_d N_A_62_94#_M1005_g N_A_241_368#_M1005_s VPB PSHORT L=0.15
+ W=1.12 AD=0.168 AS=0.308 PD=1.42 PS=2.79 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75002.5 A=0.168 P=2.54 MULT=1
MM1006 N_Y_M1005_d N_A_62_94#_M1006_g N_A_241_368#_M1006_s VPB PSHORT L=0.15
+ W=1.12 AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.6 SB=75002 A=0.168 P=2.54 MULT=1
MM1007 N_VPWR_M1007_d N_A1_M1007_g N_A_241_368#_M1006_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.1 SB=75001.6 A=0.168 P=2.54 MULT=1
MM1008 N_VPWR_M1007_d N_A1_M1008_g N_A_241_368#_M1008_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.5 SB=75001.1 A=0.168 P=2.54 MULT=1
MM1001 N_A_241_368#_M1008_s N_A2_M1001_g N_VPWR_M1001_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.1792 PD=1.42 PS=1.44 NRD=1.7533 NRS=3.5066 M=1 R=7.46667
+ SA=75002 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1010 N_A_241_368#_M1010_d N_A2_M1010_g N_VPWR_M1001_s VPB PSHORT L=0.15 W=1.12
+ AD=0.308 AS=0.1792 PD=2.79 PS=1.44 NRD=1.7533 NRS=3.5066 M=1 R=7.46667
+ SA=75002.5 SB=75000.2 A=0.168 P=2.54 MULT=1
DX14_noxref VNB VPB NWDIODE A=8.742 P=13.12
c_44 VNB 0 1.97879e-19 $X=0 $Y=0
*
.include "sky130_fd_sc_hs__a21boi_2.pxi.spice"
*
.ends
*
*
