* File: sky130_fd_sc_hs__a211o_2.pxi.spice
* Created: Tue Sep  1 19:48:30 2020
* 
x_PM_SKY130_FD_SC_HS__A211O_2%A_85_270# N_A_85_270#_M1000_d N_A_85_270#_M1010_d
+ N_A_85_270#_M1011_d N_A_85_270#_c_75_n N_A_85_270#_c_84_n N_A_85_270#_M1001_g
+ N_A_85_270#_M1005_g N_A_85_270#_c_85_n N_A_85_270#_M1002_g N_A_85_270#_M1009_g
+ N_A_85_270#_c_86_n N_A_85_270#_c_94_p N_A_85_270#_c_177_p N_A_85_270#_c_87_n
+ N_A_85_270#_c_88_n N_A_85_270#_c_78_n N_A_85_270#_c_79_n N_A_85_270#_c_89_n
+ N_A_85_270#_c_90_n N_A_85_270#_c_80_n N_A_85_270#_c_91_n N_A_85_270#_c_81_n
+ N_A_85_270#_c_113_p N_A_85_270#_c_82_n PM_SKY130_FD_SC_HS__A211O_2%A_85_270#
x_PM_SKY130_FD_SC_HS__A211O_2%A2 N_A2_M1003_g N_A2_c_207_n N_A2_M1004_g
+ N_A2_c_204_n A2 N_A2_c_205_n N_A2_c_206_n PM_SKY130_FD_SC_HS__A211O_2%A2
x_PM_SKY130_FD_SC_HS__A211O_2%A1 N_A1_M1000_g N_A1_c_251_n N_A1_M1007_g
+ N_A1_c_248_n A1 N_A1_c_249_n N_A1_c_250_n PM_SKY130_FD_SC_HS__A211O_2%A1
x_PM_SKY130_FD_SC_HS__A211O_2%B1 N_B1_M1006_g N_B1_c_294_n N_B1_c_298_n
+ N_B1_M1008_g B1 N_B1_c_295_n N_B1_c_296_n PM_SKY130_FD_SC_HS__A211O_2%B1
x_PM_SKY130_FD_SC_HS__A211O_2%C1 N_C1_c_333_n N_C1_M1011_g N_C1_M1010_g C1
+ PM_SKY130_FD_SC_HS__A211O_2%C1
x_PM_SKY130_FD_SC_HS__A211O_2%VPWR N_VPWR_M1001_s N_VPWR_M1002_s N_VPWR_M1004_d
+ N_VPWR_c_361_n N_VPWR_c_362_n N_VPWR_c_363_n N_VPWR_c_364_n VPWR
+ N_VPWR_c_365_n N_VPWR_c_366_n N_VPWR_c_367_n N_VPWR_c_360_n N_VPWR_c_369_n
+ N_VPWR_c_370_n PM_SKY130_FD_SC_HS__A211O_2%VPWR
x_PM_SKY130_FD_SC_HS__A211O_2%X N_X_M1005_s N_X_M1001_d N_X_c_411_n N_X_c_412_n
+ X X X X X PM_SKY130_FD_SC_HS__A211O_2%X
x_PM_SKY130_FD_SC_HS__A211O_2%A_317_392# N_A_317_392#_M1004_s
+ N_A_317_392#_M1007_d N_A_317_392#_c_443_n N_A_317_392#_c_439_n
+ N_A_317_392#_c_440_n PM_SKY130_FD_SC_HS__A211O_2%A_317_392#
x_PM_SKY130_FD_SC_HS__A211O_2%VGND N_VGND_M1005_d N_VGND_M1009_d N_VGND_M1006_d
+ N_VGND_c_466_n N_VGND_c_467_n N_VGND_c_468_n N_VGND_c_490_n N_VGND_c_469_n
+ N_VGND_c_470_n N_VGND_c_471_n N_VGND_c_472_n N_VGND_c_473_n N_VGND_c_474_n
+ N_VGND_c_475_n VGND N_VGND_c_476_n N_VGND_c_477_n N_VGND_c_478_n
+ PM_SKY130_FD_SC_HS__A211O_2%VGND
cc_1 VNB N_A_85_270#_c_75_n 0.01271f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=1.675
cc_2 VNB N_A_85_270#_M1005_g 0.0266606f $X=-0.19 $Y=-0.245 $X2=0.68 $Y2=0.74
cc_3 VNB N_A_85_270#_M1009_g 0.0250288f $X=-0.19 $Y=-0.245 $X2=1.11 $Y2=0.74
cc_4 VNB N_A_85_270#_c_78_n 0.00317075f $X=-0.19 $Y=-0.245 $X2=2.515 $Y2=0.515
cc_5 VNB N_A_85_270#_c_79_n 0.0111838f $X=-0.19 $Y=-0.245 $X2=3.49 $Y2=1.005
cc_6 VNB N_A_85_270#_c_80_n 0.0237055f $X=-0.19 $Y=-0.245 $X2=3.575 $Y2=0.515
cc_7 VNB N_A_85_270#_c_81_n 0.00252387f $X=-0.19 $Y=-0.245 $X2=1.17 $Y2=1.35
cc_8 VNB N_A_85_270#_c_82_n 0.0543481f $X=-0.19 $Y=-0.245 $X2=1.11 $Y2=1.557
cc_9 VNB N_A2_M1003_g 0.0222885f $X=-0.19 $Y=-0.245 $X2=3.42 $Y2=1.96
cc_10 VNB N_A2_c_204_n 0.00405643f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=1.5
cc_11 VNB N_A2_c_205_n 0.0032582f $X=-0.19 $Y=-0.245 $X2=0.68 $Y2=1.35
cc_12 VNB N_A2_c_206_n 0.0443914f $X=-0.19 $Y=-0.245 $X2=0.68 $Y2=0.74
cc_13 VNB N_A1_M1000_g 0.0203333f $X=-0.19 $Y=-0.245 $X2=3.42 $Y2=1.96
cc_14 VNB N_A1_c_248_n 0.00364784f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=1.5
cc_15 VNB N_A1_c_249_n 0.0306419f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=2.4
cc_16 VNB N_A1_c_250_n 0.00551212f $X=-0.19 $Y=-0.245 $X2=0.68 $Y2=1.35
cc_17 VNB N_B1_M1006_g 0.0214297f $X=-0.19 $Y=-0.245 $X2=3.42 $Y2=1.96
cc_18 VNB N_B1_c_294_n 0.00318739f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_B1_c_295_n 0.0297888f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=2.4
cc_20 VNB N_B1_c_296_n 0.00683457f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=2.4
cc_21 VNB N_C1_c_333_n 0.0333068f $X=-0.19 $Y=-0.245 $X2=2.355 $Y2=0.37
cc_22 VNB N_C1_M1010_g 0.0428504f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB C1 0.0035847f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_VPWR_c_360_n 0.163682f $X=-0.19 $Y=-0.245 $X2=3.57 $Y2=2.815
cc_25 VNB N_X_c_411_n 0.0017881f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_X_c_412_n 0.00593091f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=2.4
cc_27 VNB X 0.00870155f $X=-0.19 $Y=-0.245 $X2=0.68 $Y2=0.74
cc_28 VNB N_VGND_c_466_n 0.0290431f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=1.765
cc_29 VNB N_VGND_c_467_n 0.0151736f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=2.4
cc_30 VNB N_VGND_c_468_n 0.00464087f $X=-0.19 $Y=-0.245 $X2=0.68 $Y2=0.74
cc_31 VNB N_VGND_c_469_n 0.00356735f $X=-0.19 $Y=-0.245 $X2=0.965 $Y2=2.4
cc_32 VNB N_VGND_c_470_n 0.00548601f $X=-0.19 $Y=-0.245 $X2=1.11 $Y2=0.74
cc_33 VNB N_VGND_c_471_n 0.0116899f $X=-0.19 $Y=-0.245 $X2=1.11 $Y2=0.74
cc_34 VNB N_VGND_c_472_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_473_n 0.0415749f $X=-0.19 $Y=-0.245 $X2=1.25 $Y2=1.35
cc_36 VNB N_VGND_c_474_n 0.00307912f $X=-0.19 $Y=-0.245 $X2=1.25 $Y2=1.68
cc_37 VNB N_VGND_c_475_n 0.00195927f $X=-0.19 $Y=-0.245 $X2=3.405 $Y2=2.035
cc_38 VNB N_VGND_c_476_n 0.0234852f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_477_n 0.244793f $X=-0.19 $Y=-0.245 $X2=1.17 $Y2=1.515
cc_40 VNB N_VGND_c_478_n 0.00311272f $X=-0.19 $Y=-0.245 $X2=1.17 $Y2=1.35
cc_41 VPB N_A_85_270#_c_75_n 0.00111912f $X=-0.19 $Y=1.66 $X2=0.515 $Y2=1.675
cc_42 VPB N_A_85_270#_c_84_n 0.0258384f $X=-0.19 $Y=1.66 $X2=0.515 $Y2=1.765
cc_43 VPB N_A_85_270#_c_85_n 0.0172159f $X=-0.19 $Y=1.66 $X2=0.965 $Y2=1.765
cc_44 VPB N_A_85_270#_c_86_n 0.00419525f $X=-0.19 $Y=1.66 $X2=1.25 $Y2=1.95
cc_45 VPB N_A_85_270#_c_87_n 0.0313759f $X=-0.19 $Y=1.66 $X2=3.405 $Y2=2.035
cc_46 VPB N_A_85_270#_c_88_n 3.13193e-19 $X=-0.19 $Y=1.66 $X2=1.335 $Y2=2.035
cc_47 VPB N_A_85_270#_c_89_n 0.00908171f $X=-0.19 $Y=1.66 $X2=3.57 $Y2=2.12
cc_48 VPB N_A_85_270#_c_90_n 0.0360166f $X=-0.19 $Y=1.66 $X2=3.57 $Y2=2.815
cc_49 VPB N_A_85_270#_c_91_n 0.00178597f $X=-0.19 $Y=1.66 $X2=1.17 $Y2=1.515
cc_50 VPB N_A_85_270#_c_82_n 0.0160011f $X=-0.19 $Y=1.66 $X2=1.11 $Y2=1.557
cc_51 VPB N_A2_c_207_n 0.0311719f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_52 VPB N_A2_c_204_n 0.00445766f $X=-0.19 $Y=1.66 $X2=0.515 $Y2=1.5
cc_53 VPB N_A2_c_205_n 0.00374417f $X=-0.19 $Y=1.66 $X2=0.68 $Y2=1.35
cc_54 VPB N_A1_c_251_n 0.0274273f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_55 VPB N_A1_c_248_n 0.00364784f $X=-0.19 $Y=1.66 $X2=0.515 $Y2=1.5
cc_56 VPB N_A1_c_250_n 0.00388517f $X=-0.19 $Y=1.66 $X2=0.68 $Y2=1.35
cc_57 VPB N_B1_c_294_n 0.00619599f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_58 VPB N_B1_c_298_n 0.0216637f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_59 VPB N_B1_c_296_n 0.00437976f $X=-0.19 $Y=1.66 $X2=0.515 $Y2=2.4
cc_60 VPB N_C1_c_333_n 0.0546125f $X=-0.19 $Y=1.66 $X2=2.355 $Y2=0.37
cc_61 VPB C1 0.00276779f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_62 VPB N_VPWR_c_361_n 0.0109711f $X=-0.19 $Y=1.66 $X2=0.515 $Y2=1.5
cc_63 VPB N_VPWR_c_362_n 0.0647053f $X=-0.19 $Y=1.66 $X2=0.515 $Y2=1.765
cc_64 VPB N_VPWR_c_363_n 0.0128119f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_65 VPB N_VPWR_c_364_n 0.0093235f $X=-0.19 $Y=1.66 $X2=1.11 $Y2=1.35
cc_66 VPB N_VPWR_c_365_n 0.0184472f $X=-0.19 $Y=1.66 $X2=1.25 $Y2=1.09
cc_67 VPB N_VPWR_c_366_n 0.0202859f $X=-0.19 $Y=1.66 $X2=1.335 $Y2=1.005
cc_68 VPB N_VPWR_c_367_n 0.0439561f $X=-0.19 $Y=1.66 $X2=3.57 $Y2=2.815
cc_69 VPB N_VPWR_c_360_n 0.0819269f $X=-0.19 $Y=1.66 $X2=3.57 $Y2=2.815
cc_70 VPB N_VPWR_c_369_n 0.00614127f $X=-0.19 $Y=1.66 $X2=1.17 $Y2=1.515
cc_71 VPB N_VPWR_c_370_n 0.00555219f $X=-0.19 $Y=1.66 $X2=1.17 $Y2=1.35
cc_72 VPB X 0.0037735f $X=-0.19 $Y=1.66 $X2=0.68 $Y2=0.74
cc_73 VPB N_A_317_392#_c_439_n 0.00927352f $X=-0.19 $Y=1.66 $X2=0.515 $Y2=2.4
cc_74 VPB N_A_317_392#_c_440_n 0.00257417f $X=-0.19 $Y=1.66 $X2=0.68 $Y2=0.74
cc_75 N_A_85_270#_M1009_g N_A2_M1003_g 0.00936275f $X=1.11 $Y=0.74 $X2=0 $Y2=0
cc_76 N_A_85_270#_c_94_p N_A2_M1003_g 0.0188837f $X=2.33 $Y=1.005 $X2=0 $Y2=0
cc_77 N_A_85_270#_c_78_n N_A2_M1003_g 0.00193971f $X=2.515 $Y=0.515 $X2=0 $Y2=0
cc_78 N_A_85_270#_c_81_n N_A2_M1003_g 0.0026977f $X=1.17 $Y=1.35 $X2=0 $Y2=0
cc_79 N_A_85_270#_c_86_n N_A2_c_207_n 0.00408199f $X=1.25 $Y=1.95 $X2=0 $Y2=0
cc_80 N_A_85_270#_c_87_n N_A2_c_207_n 0.0181021f $X=3.405 $Y=2.035 $X2=0 $Y2=0
cc_81 N_A_85_270#_c_86_n N_A2_c_204_n 3.67047e-19 $X=1.25 $Y=1.95 $X2=0 $Y2=0
cc_82 N_A_85_270#_c_82_n N_A2_c_204_n 0.00161944f $X=1.11 $Y=1.557 $X2=0 $Y2=0
cc_83 N_A_85_270#_c_94_p N_A2_c_205_n 0.0230785f $X=2.33 $Y=1.005 $X2=0 $Y2=0
cc_84 N_A_85_270#_c_87_n N_A2_c_205_n 0.0269175f $X=3.405 $Y=2.035 $X2=0 $Y2=0
cc_85 N_A_85_270#_c_81_n N_A2_c_205_n 0.0338358f $X=1.17 $Y=1.35 $X2=0 $Y2=0
cc_86 N_A_85_270#_c_82_n N_A2_c_205_n 0.00179973f $X=1.11 $Y=1.557 $X2=0 $Y2=0
cc_87 N_A_85_270#_M1009_g N_A2_c_206_n 0.00279477f $X=1.11 $Y=0.74 $X2=0 $Y2=0
cc_88 N_A_85_270#_c_94_p N_A2_c_206_n 0.00198342f $X=2.33 $Y=1.005 $X2=0 $Y2=0
cc_89 N_A_85_270#_c_87_n N_A2_c_206_n 0.00134333f $X=3.405 $Y=2.035 $X2=0 $Y2=0
cc_90 N_A_85_270#_c_91_n N_A2_c_206_n 8.85995e-19 $X=1.17 $Y=1.515 $X2=0 $Y2=0
cc_91 N_A_85_270#_c_81_n N_A2_c_206_n 6.65509e-19 $X=1.17 $Y=1.35 $X2=0 $Y2=0
cc_92 N_A_85_270#_c_82_n N_A2_c_206_n 0.0156904f $X=1.11 $Y=1.557 $X2=0 $Y2=0
cc_93 N_A_85_270#_c_94_p N_A1_M1000_g 0.0106432f $X=2.33 $Y=1.005 $X2=0 $Y2=0
cc_94 N_A_85_270#_c_78_n N_A1_M1000_g 0.0100536f $X=2.515 $Y=0.515 $X2=0 $Y2=0
cc_95 N_A_85_270#_c_113_p N_A1_M1000_g 7.3104e-19 $X=2.515 $Y=1.005 $X2=0 $Y2=0
cc_96 N_A_85_270#_c_87_n N_A1_c_251_n 0.0124566f $X=3.405 $Y=2.035 $X2=0 $Y2=0
cc_97 N_A_85_270#_c_113_p N_A1_c_251_n 8.26903e-19 $X=2.515 $Y=1.005 $X2=0 $Y2=0
cc_98 N_A_85_270#_c_87_n N_A1_c_249_n 8.00066e-19 $X=3.405 $Y=2.035 $X2=0 $Y2=0
cc_99 N_A_85_270#_c_113_p N_A1_c_249_n 0.00123018f $X=2.515 $Y=1.005 $X2=0 $Y2=0
cc_100 N_A_85_270#_c_94_p N_A1_c_250_n 0.0199035f $X=2.33 $Y=1.005 $X2=0 $Y2=0
cc_101 N_A_85_270#_c_87_n N_A1_c_250_n 0.0391613f $X=3.405 $Y=2.035 $X2=0 $Y2=0
cc_102 N_A_85_270#_c_113_p N_A1_c_250_n 0.0148045f $X=2.515 $Y=1.005 $X2=0 $Y2=0
cc_103 N_A_85_270#_c_78_n N_B1_M1006_g 0.00333996f $X=2.515 $Y=0.515 $X2=0 $Y2=0
cc_104 N_A_85_270#_c_79_n N_B1_M1006_g 0.0153168f $X=3.49 $Y=1.005 $X2=0 $Y2=0
cc_105 N_A_85_270#_c_87_n N_B1_c_298_n 0.0154523f $X=3.405 $Y=2.035 $X2=0 $Y2=0
cc_106 N_A_85_270#_c_90_n N_B1_c_298_n 0.00280499f $X=3.57 $Y=2.815 $X2=0 $Y2=0
cc_107 N_A_85_270#_c_87_n N_B1_c_295_n 6.643e-19 $X=3.405 $Y=2.035 $X2=0 $Y2=0
cc_108 N_A_85_270#_c_79_n N_B1_c_295_n 0.00113349f $X=3.49 $Y=1.005 $X2=0 $Y2=0
cc_109 N_A_85_270#_c_87_n N_B1_c_296_n 0.0389655f $X=3.405 $Y=2.035 $X2=0 $Y2=0
cc_110 N_A_85_270#_c_79_n N_B1_c_296_n 0.03557f $X=3.49 $Y=1.005 $X2=0 $Y2=0
cc_111 N_A_85_270#_c_87_n N_C1_c_333_n 0.016376f $X=3.405 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_112 N_A_85_270#_c_79_n N_C1_c_333_n 0.00178482f $X=3.49 $Y=1.005 $X2=-0.19
+ $Y2=-0.245
cc_113 N_A_85_270#_c_89_n N_C1_c_333_n 0.00344035f $X=3.57 $Y=2.12 $X2=-0.19
+ $Y2=-0.245
cc_114 N_A_85_270#_c_90_n N_C1_c_333_n 0.0151081f $X=3.57 $Y=2.815 $X2=-0.19
+ $Y2=-0.245
cc_115 N_A_85_270#_c_79_n N_C1_M1010_g 0.0174318f $X=3.49 $Y=1.005 $X2=0 $Y2=0
cc_116 N_A_85_270#_c_80_n N_C1_M1010_g 0.00161119f $X=3.575 $Y=0.515 $X2=0 $Y2=0
cc_117 N_A_85_270#_c_79_n C1 0.0151444f $X=3.49 $Y=1.005 $X2=0 $Y2=0
cc_118 N_A_85_270#_c_89_n C1 0.0277331f $X=3.57 $Y=2.12 $X2=0 $Y2=0
cc_119 N_A_85_270#_c_86_n N_VPWR_M1002_s 0.00191369f $X=1.25 $Y=1.95 $X2=0 $Y2=0
cc_120 N_A_85_270#_c_88_n N_VPWR_M1002_s 0.00495189f $X=1.335 $Y=2.035 $X2=0
+ $Y2=0
cc_121 N_A_85_270#_c_87_n N_VPWR_M1004_d 0.00320511f $X=3.405 $Y=2.035 $X2=0
+ $Y2=0
cc_122 N_A_85_270#_c_84_n N_VPWR_c_362_n 0.008783f $X=0.515 $Y=1.765 $X2=0 $Y2=0
cc_123 N_A_85_270#_c_84_n N_VPWR_c_363_n 5.56513e-19 $X=0.515 $Y=1.765 $X2=0
+ $Y2=0
cc_124 N_A_85_270#_c_85_n N_VPWR_c_363_n 0.0121809f $X=0.965 $Y=1.765 $X2=0
+ $Y2=0
cc_125 N_A_85_270#_c_87_n N_VPWR_c_363_n 0.00156694f $X=3.405 $Y=2.035 $X2=0
+ $Y2=0
cc_126 N_A_85_270#_c_88_n N_VPWR_c_363_n 0.0153531f $X=1.335 $Y=2.035 $X2=0
+ $Y2=0
cc_127 N_A_85_270#_c_91_n N_VPWR_c_363_n 0.00317781f $X=1.17 $Y=1.515 $X2=0
+ $Y2=0
cc_128 N_A_85_270#_c_82_n N_VPWR_c_363_n 0.00105405f $X=1.11 $Y=1.557 $X2=0
+ $Y2=0
cc_129 N_A_85_270#_c_84_n N_VPWR_c_365_n 0.00445602f $X=0.515 $Y=1.765 $X2=0
+ $Y2=0
cc_130 N_A_85_270#_c_85_n N_VPWR_c_365_n 0.00413917f $X=0.965 $Y=1.765 $X2=0
+ $Y2=0
cc_131 N_A_85_270#_c_90_n N_VPWR_c_367_n 0.0145938f $X=3.57 $Y=2.815 $X2=0 $Y2=0
cc_132 N_A_85_270#_c_84_n N_VPWR_c_360_n 0.00861117f $X=0.515 $Y=1.765 $X2=0
+ $Y2=0
cc_133 N_A_85_270#_c_85_n N_VPWR_c_360_n 0.00817726f $X=0.965 $Y=1.765 $X2=0
+ $Y2=0
cc_134 N_A_85_270#_c_90_n N_VPWR_c_360_n 0.0120466f $X=3.57 $Y=2.815 $X2=0 $Y2=0
cc_135 N_A_85_270#_M1005_g N_X_c_411_n 3.92313e-19 $X=0.68 $Y=0.74 $X2=0 $Y2=0
cc_136 N_A_85_270#_M1009_g N_X_c_411_n 3.92031e-19 $X=1.11 $Y=0.74 $X2=0 $Y2=0
cc_137 N_A_85_270#_M1005_g N_X_c_412_n 0.0117483f $X=0.68 $Y=0.74 $X2=0 $Y2=0
cc_138 N_A_85_270#_M1009_g N_X_c_412_n 5.39763e-19 $X=1.11 $Y=0.74 $X2=0 $Y2=0
cc_139 N_A_85_270#_c_81_n N_X_c_412_n 0.00556069f $X=1.17 $Y=1.35 $X2=0 $Y2=0
cc_140 N_A_85_270#_c_82_n N_X_c_412_n 0.00424762f $X=1.11 $Y=1.557 $X2=0 $Y2=0
cc_141 N_A_85_270#_c_75_n X 0.00899625f $X=0.515 $Y=1.675 $X2=0 $Y2=0
cc_142 N_A_85_270#_c_84_n X 0.0213056f $X=0.515 $Y=1.765 $X2=0 $Y2=0
cc_143 N_A_85_270#_M1005_g X 0.0062358f $X=0.68 $Y=0.74 $X2=0 $Y2=0
cc_144 N_A_85_270#_c_85_n X 0.0011171f $X=0.965 $Y=1.765 $X2=0 $Y2=0
cc_145 N_A_85_270#_M1009_g X 0.00123769f $X=1.11 $Y=0.74 $X2=0 $Y2=0
cc_146 N_A_85_270#_c_86_n X 0.0102211f $X=1.25 $Y=1.95 $X2=0 $Y2=0
cc_147 N_A_85_270#_c_91_n X 0.0250323f $X=1.17 $Y=1.515 $X2=0 $Y2=0
cc_148 N_A_85_270#_c_81_n X 0.00767189f $X=1.17 $Y=1.35 $X2=0 $Y2=0
cc_149 N_A_85_270#_c_82_n X 0.0169711f $X=1.11 $Y=1.557 $X2=0 $Y2=0
cc_150 N_A_85_270#_c_87_n N_A_317_392#_M1004_s 0.00315345f $X=3.405 $Y=2.035
+ $X2=-0.19 $Y2=-0.245
cc_151 N_A_85_270#_c_87_n N_A_317_392#_M1007_d 0.00197722f $X=3.405 $Y=2.035
+ $X2=0 $Y2=0
cc_152 N_A_85_270#_c_87_n N_A_317_392#_c_443_n 0.0382797f $X=3.405 $Y=2.035
+ $X2=0 $Y2=0
cc_153 N_A_85_270#_c_85_n N_A_317_392#_c_439_n 8.39569e-19 $X=0.965 $Y=1.765
+ $X2=0 $Y2=0
cc_154 N_A_85_270#_c_87_n N_A_317_392#_c_439_n 0.0221949f $X=3.405 $Y=2.035
+ $X2=0 $Y2=0
cc_155 N_A_85_270#_c_87_n N_A_317_392#_c_440_n 0.0173542f $X=3.405 $Y=2.035
+ $X2=0 $Y2=0
cc_156 N_A_85_270#_c_90_n N_A_317_392#_c_440_n 0.0203497f $X=3.57 $Y=2.815 $X2=0
+ $Y2=0
cc_157 N_A_85_270#_c_87_n A_600_392# 0.00595227f $X=3.405 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_158 N_A_85_270#_c_94_p N_VGND_M1009_d 0.0174908f $X=2.33 $Y=1.005 $X2=0 $Y2=0
cc_159 N_A_85_270#_c_177_p N_VGND_M1009_d 0.0010293f $X=1.335 $Y=1.005 $X2=0
+ $Y2=0
cc_160 N_A_85_270#_c_81_n N_VGND_M1009_d 2.95258e-19 $X=1.17 $Y=1.35 $X2=0 $Y2=0
cc_161 N_A_85_270#_c_79_n N_VGND_M1006_d 0.00585867f $X=3.49 $Y=1.005 $X2=0
+ $Y2=0
cc_162 N_A_85_270#_M1005_g N_VGND_c_466_n 0.0120602f $X=0.68 $Y=0.74 $X2=0 $Y2=0
cc_163 N_A_85_270#_M1009_g N_VGND_c_466_n 4.71636e-19 $X=1.11 $Y=0.74 $X2=0
+ $Y2=0
cc_164 N_A_85_270#_c_82_n N_VGND_c_466_n 0.00461225f $X=1.11 $Y=1.557 $X2=0
+ $Y2=0
cc_165 N_A_85_270#_M1005_g N_VGND_c_467_n 0.00383152f $X=0.68 $Y=0.74 $X2=0
+ $Y2=0
cc_166 N_A_85_270#_M1009_g N_VGND_c_467_n 0.00383152f $X=1.11 $Y=0.74 $X2=0
+ $Y2=0
cc_167 N_A_85_270#_M1005_g N_VGND_c_468_n 3.2548e-19 $X=0.68 $Y=0.74 $X2=0 $Y2=0
cc_168 N_A_85_270#_M1009_g N_VGND_c_468_n 0.00384973f $X=1.11 $Y=0.74 $X2=0
+ $Y2=0
cc_169 N_A_85_270#_M1009_g N_VGND_c_490_n 0.00491108f $X=1.11 $Y=0.74 $X2=0
+ $Y2=0
cc_170 N_A_85_270#_c_177_p N_VGND_c_490_n 0.00962725f $X=1.335 $Y=1.005 $X2=0
+ $Y2=0
cc_171 N_A_85_270#_c_82_n N_VGND_c_490_n 4.02474e-19 $X=1.11 $Y=1.557 $X2=0
+ $Y2=0
cc_172 N_A_85_270#_c_94_p N_VGND_c_469_n 0.0369249f $X=2.33 $Y=1.005 $X2=0 $Y2=0
cc_173 N_A_85_270#_c_177_p N_VGND_c_469_n 3.90227e-19 $X=1.335 $Y=1.005 $X2=0
+ $Y2=0
cc_174 N_A_85_270#_c_78_n N_VGND_c_469_n 0.0142905f $X=2.515 $Y=0.515 $X2=0
+ $Y2=0
cc_175 N_A_85_270#_c_78_n N_VGND_c_473_n 0.0163488f $X=2.515 $Y=0.515 $X2=0
+ $Y2=0
cc_176 N_A_85_270#_c_78_n N_VGND_c_475_n 0.0164559f $X=2.515 $Y=0.515 $X2=0
+ $Y2=0
cc_177 N_A_85_270#_c_79_n N_VGND_c_475_n 0.0250026f $X=3.49 $Y=1.005 $X2=0 $Y2=0
cc_178 N_A_85_270#_c_80_n N_VGND_c_475_n 0.0156761f $X=3.575 $Y=0.515 $X2=0
+ $Y2=0
cc_179 N_A_85_270#_c_80_n N_VGND_c_476_n 0.011066f $X=3.575 $Y=0.515 $X2=0 $Y2=0
cc_180 N_A_85_270#_M1005_g N_VGND_c_477_n 0.0075754f $X=0.68 $Y=0.74 $X2=0 $Y2=0
cc_181 N_A_85_270#_M1009_g N_VGND_c_477_n 0.0075754f $X=1.11 $Y=0.74 $X2=0 $Y2=0
cc_182 N_A_85_270#_c_78_n N_VGND_c_477_n 0.0134757f $X=2.515 $Y=0.515 $X2=0
+ $Y2=0
cc_183 N_A_85_270#_c_80_n N_VGND_c_477_n 0.00915947f $X=3.575 $Y=0.515 $X2=0
+ $Y2=0
cc_184 N_A_85_270#_c_94_p A_399_74# 0.00468343f $X=2.33 $Y=1.005 $X2=-0.19
+ $Y2=-0.245
cc_185 N_A2_M1003_g N_A1_M1000_g 0.0416311f $X=1.92 $Y=0.74 $X2=0 $Y2=0
cc_186 N_A2_c_207_n N_A1_c_251_n 0.0351454f $X=1.935 $Y=1.885 $X2=0 $Y2=0
cc_187 N_A2_c_204_n N_A1_c_248_n 0.0034522f $X=1.935 $Y=1.73 $X2=0 $Y2=0
cc_188 N_A2_c_205_n N_A1_c_249_n 2.5478e-19 $X=1.71 $Y=1.425 $X2=0 $Y2=0
cc_189 N_A2_c_206_n N_A1_c_249_n 0.0416311f $X=1.92 $Y=1.425 $X2=0 $Y2=0
cc_190 N_A2_c_207_n N_A1_c_250_n 4.83978e-19 $X=1.935 $Y=1.885 $X2=0 $Y2=0
cc_191 N_A2_c_205_n N_A1_c_250_n 0.0424031f $X=1.71 $Y=1.425 $X2=0 $Y2=0
cc_192 N_A2_c_206_n N_A1_c_250_n 0.00385707f $X=1.92 $Y=1.425 $X2=0 $Y2=0
cc_193 N_A2_c_207_n N_VPWR_c_363_n 0.00391987f $X=1.935 $Y=1.885 $X2=0 $Y2=0
cc_194 N_A2_c_207_n N_VPWR_c_364_n 0.0043537f $X=1.935 $Y=1.885 $X2=0 $Y2=0
cc_195 N_A2_c_207_n N_VPWR_c_366_n 0.00445602f $X=1.935 $Y=1.885 $X2=0 $Y2=0
cc_196 N_A2_c_207_n N_VPWR_c_360_n 0.00863223f $X=1.935 $Y=1.885 $X2=0 $Y2=0
cc_197 N_A2_c_207_n N_A_317_392#_c_443_n 0.0121961f $X=1.935 $Y=1.885 $X2=0
+ $Y2=0
cc_198 N_A2_c_207_n N_A_317_392#_c_439_n 0.00781981f $X=1.935 $Y=1.885 $X2=0
+ $Y2=0
cc_199 N_A2_c_207_n N_A_317_392#_c_440_n 5.47349e-19 $X=1.935 $Y=1.885 $X2=0
+ $Y2=0
cc_200 N_A2_M1003_g N_VGND_c_468_n 0.00170329f $X=1.92 $Y=0.74 $X2=0 $Y2=0
cc_201 N_A2_M1003_g N_VGND_c_469_n 0.00732382f $X=1.92 $Y=0.74 $X2=0 $Y2=0
cc_202 N_A2_M1003_g N_VGND_c_473_n 0.00433162f $X=1.92 $Y=0.74 $X2=0 $Y2=0
cc_203 N_A2_M1003_g N_VGND_c_477_n 0.00819679f $X=1.92 $Y=0.74 $X2=0 $Y2=0
cc_204 N_A1_M1000_g N_B1_M1006_g 0.018661f $X=2.28 $Y=0.74 $X2=0 $Y2=0
cc_205 N_A1_c_251_n N_B1_c_294_n 0.00780146f $X=2.475 $Y=1.885 $X2=0 $Y2=0
cc_206 N_A1_c_248_n N_B1_c_294_n 0.00517221f $X=2.475 $Y=1.73 $X2=0 $Y2=0
cc_207 N_A1_c_250_n N_B1_c_294_n 2.06886e-19 $X=2.37 $Y=1.425 $X2=0 $Y2=0
cc_208 N_A1_c_251_n N_B1_c_298_n 0.0223339f $X=2.475 $Y=1.885 $X2=0 $Y2=0
cc_209 N_A1_c_249_n N_B1_c_295_n 0.0201104f $X=2.37 $Y=1.425 $X2=0 $Y2=0
cc_210 N_A1_c_250_n N_B1_c_295_n 0.00114728f $X=2.37 $Y=1.425 $X2=0 $Y2=0
cc_211 N_A1_c_251_n N_B1_c_296_n 3.31736e-19 $X=2.475 $Y=1.885 $X2=0 $Y2=0
cc_212 N_A1_c_248_n N_B1_c_296_n 8.93334e-19 $X=2.475 $Y=1.73 $X2=0 $Y2=0
cc_213 N_A1_c_249_n N_B1_c_296_n 0.00114728f $X=2.37 $Y=1.425 $X2=0 $Y2=0
cc_214 N_A1_c_250_n N_B1_c_296_n 0.0357827f $X=2.37 $Y=1.425 $X2=0 $Y2=0
cc_215 N_A1_c_251_n N_VPWR_c_364_n 0.0052183f $X=2.475 $Y=1.885 $X2=0 $Y2=0
cc_216 N_A1_c_251_n N_VPWR_c_367_n 0.00445602f $X=2.475 $Y=1.885 $X2=0 $Y2=0
cc_217 N_A1_c_251_n N_VPWR_c_360_n 0.00857833f $X=2.475 $Y=1.885 $X2=0 $Y2=0
cc_218 N_A1_c_251_n N_A_317_392#_c_443_n 0.0121961f $X=2.475 $Y=1.885 $X2=0
+ $Y2=0
cc_219 N_A1_c_251_n N_A_317_392#_c_439_n 6.06825e-19 $X=2.475 $Y=1.885 $X2=0
+ $Y2=0
cc_220 N_A1_c_251_n N_A_317_392#_c_440_n 0.00741768f $X=2.475 $Y=1.885 $X2=0
+ $Y2=0
cc_221 N_A1_M1000_g N_VGND_c_469_n 0.00107858f $X=2.28 $Y=0.74 $X2=0 $Y2=0
cc_222 N_A1_M1000_g N_VGND_c_470_n 5.22255e-19 $X=2.28 $Y=0.74 $X2=0 $Y2=0
cc_223 N_A1_M1000_g N_VGND_c_473_n 0.00434272f $X=2.28 $Y=0.74 $X2=0 $Y2=0
cc_224 N_A1_M1000_g N_VGND_c_477_n 0.00821699f $X=2.28 $Y=0.74 $X2=0 $Y2=0
cc_225 N_B1_c_294_n N_C1_c_333_n 0.0152523f $X=2.925 $Y=1.795 $X2=-0.19
+ $Y2=-0.245
cc_226 N_B1_c_298_n N_C1_c_333_n 0.0544725f $X=2.925 $Y=1.885 $X2=-0.19
+ $Y2=-0.245
cc_227 N_B1_c_296_n N_C1_c_333_n 4.48526e-19 $X=2.91 $Y=1.425 $X2=-0.19
+ $Y2=-0.245
cc_228 N_B1_M1006_g N_C1_M1010_g 0.0195423f $X=2.82 $Y=0.74 $X2=0 $Y2=0
cc_229 N_B1_c_295_n N_C1_M1010_g 0.0199123f $X=2.91 $Y=1.425 $X2=0 $Y2=0
cc_230 N_B1_c_296_n N_C1_M1010_g 0.00774557f $X=2.91 $Y=1.425 $X2=0 $Y2=0
cc_231 N_B1_c_296_n C1 0.0269573f $X=2.91 $Y=1.425 $X2=0 $Y2=0
cc_232 N_B1_c_298_n N_VPWR_c_367_n 0.00445602f $X=2.925 $Y=1.885 $X2=0 $Y2=0
cc_233 N_B1_c_298_n N_VPWR_c_360_n 0.00858241f $X=2.925 $Y=1.885 $X2=0 $Y2=0
cc_234 N_B1_c_298_n N_A_317_392#_c_440_n 0.0122028f $X=2.925 $Y=1.885 $X2=0
+ $Y2=0
cc_235 N_B1_M1006_g N_VGND_c_470_n 0.00368901f $X=2.82 $Y=0.74 $X2=0 $Y2=0
cc_236 N_B1_M1006_g N_VGND_c_473_n 0.00383152f $X=2.82 $Y=0.74 $X2=0 $Y2=0
cc_237 N_B1_M1006_g N_VGND_c_475_n 0.00479502f $X=2.82 $Y=0.74 $X2=0 $Y2=0
cc_238 N_B1_M1006_g N_VGND_c_477_n 0.00758569f $X=2.82 $Y=0.74 $X2=0 $Y2=0
cc_239 N_C1_c_333_n N_VPWR_c_367_n 0.00445602f $X=3.345 $Y=1.885 $X2=0 $Y2=0
cc_240 N_C1_c_333_n N_VPWR_c_360_n 0.00861618f $X=3.345 $Y=1.885 $X2=0 $Y2=0
cc_241 N_C1_c_333_n N_A_317_392#_c_440_n 0.00198831f $X=3.345 $Y=1.885 $X2=0
+ $Y2=0
cc_242 N_C1_M1010_g N_VGND_c_470_n 0.00216113f $X=3.36 $Y=0.74 $X2=0 $Y2=0
cc_243 N_C1_M1010_g N_VGND_c_475_n 0.00523524f $X=3.36 $Y=0.74 $X2=0 $Y2=0
cc_244 N_C1_M1010_g N_VGND_c_476_n 0.00433162f $X=3.36 $Y=0.74 $X2=0 $Y2=0
cc_245 N_C1_M1010_g N_VGND_c_477_n 0.00822253f $X=3.36 $Y=0.74 $X2=0 $Y2=0
cc_246 N_VPWR_c_362_n X 0.0764675f $X=0.29 $Y=1.985 $X2=0 $Y2=0
cc_247 N_VPWR_c_363_n X 0.0243883f $X=1.19 $Y=2.455 $X2=0 $Y2=0
cc_248 N_VPWR_c_365_n X 0.0114703f $X=1.025 $Y=3.33 $X2=0 $Y2=0
cc_249 N_VPWR_c_360_n X 0.00946127f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_250 N_VPWR_M1004_d N_A_317_392#_c_443_n 0.00640171f $X=2.01 $Y=1.96 $X2=0
+ $Y2=0
cc_251 N_VPWR_c_364_n N_A_317_392#_c_443_n 0.0217227f $X=2.18 $Y=2.805 $X2=0
+ $Y2=0
cc_252 N_VPWR_c_363_n N_A_317_392#_c_439_n 0.0539029f $X=1.19 $Y=2.455 $X2=0
+ $Y2=0
cc_253 N_VPWR_c_364_n N_A_317_392#_c_439_n 0.023766f $X=2.18 $Y=2.805 $X2=0
+ $Y2=0
cc_254 N_VPWR_c_366_n N_A_317_392#_c_439_n 0.0146094f $X=2.075 $Y=3.33 $X2=0
+ $Y2=0
cc_255 N_VPWR_c_360_n N_A_317_392#_c_439_n 0.0120527f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_256 N_VPWR_c_364_n N_A_317_392#_c_440_n 0.013908f $X=2.18 $Y=2.805 $X2=0
+ $Y2=0
cc_257 N_VPWR_c_367_n N_A_317_392#_c_440_n 0.0145674f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_258 N_VPWR_c_360_n N_A_317_392#_c_440_n 0.0119851f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_259 N_X_c_411_n N_VGND_c_466_n 0.0182488f $X=0.895 $Y=0.515 $X2=0 $Y2=0
cc_260 N_X_c_412_n N_VGND_c_466_n 0.00182821f $X=0.895 $Y=1.095 $X2=0 $Y2=0
cc_261 N_X_c_411_n N_VGND_c_467_n 0.00747999f $X=0.895 $Y=0.515 $X2=0 $Y2=0
cc_262 N_X_c_411_n N_VGND_c_490_n 0.0168852f $X=0.895 $Y=0.515 $X2=0 $Y2=0
cc_263 N_X_c_411_n N_VGND_c_477_n 0.00619848f $X=0.895 $Y=0.515 $X2=0 $Y2=0
