* File: sky130_fd_sc_hs__o311ai_2.pxi.spice
* Created: Tue Sep  1 20:17:43 2020
* 
x_PM_SKY130_FD_SC_HS__O311AI_2%A1 N_A1_M1000_g N_A1_c_103_n N_A1_M1009_g
+ N_A1_c_104_n N_A1_M1018_g N_A1_M1019_g A1 A1 N_A1_c_102_n
+ PM_SKY130_FD_SC_HS__O311AI_2%A1
x_PM_SKY130_FD_SC_HS__O311AI_2%A2 N_A2_c_145_n N_A2_M1007_g N_A2_M1012_g
+ N_A2_M1013_g N_A2_c_146_n N_A2_M1015_g A2 A2 A2 N_A2_c_144_n
+ PM_SKY130_FD_SC_HS__O311AI_2%A2
x_PM_SKY130_FD_SC_HS__O311AI_2%A3 N_A3_M1005_g N_A3_M1017_g N_A3_c_200_n
+ N_A3_M1002_g N_A3_c_197_n N_A3_c_198_n N_A3_c_203_n N_A3_M1004_g A3 A3
+ PM_SKY130_FD_SC_HS__O311AI_2%A3
x_PM_SKY130_FD_SC_HS__O311AI_2%B1 N_B1_c_257_n N_B1_M1003_g N_B1_c_258_n
+ N_B1_c_259_n N_B1_c_260_n N_B1_M1014_g N_B1_c_265_n N_B1_M1006_g N_B1_c_266_n
+ N_B1_M1008_g N_B1_c_261_n N_B1_c_262_n B1 B1 N_B1_c_264_n
+ PM_SKY130_FD_SC_HS__O311AI_2%B1
x_PM_SKY130_FD_SC_HS__O311AI_2%C1 N_C1_c_331_n N_C1_M1010_g N_C1_M1001_g
+ N_C1_c_332_n N_C1_M1016_g N_C1_M1011_g C1 C1 N_C1_c_330_n
+ PM_SKY130_FD_SC_HS__O311AI_2%C1
x_PM_SKY130_FD_SC_HS__O311AI_2%A_28_368# N_A_28_368#_M1009_s N_A_28_368#_M1018_s
+ N_A_28_368#_M1015_s N_A_28_368#_c_377_n N_A_28_368#_c_378_n
+ N_A_28_368#_c_385_n N_A_28_368#_c_379_n N_A_28_368#_c_391_n
+ N_A_28_368#_c_395_n N_A_28_368#_c_380_n PM_SKY130_FD_SC_HS__O311AI_2%A_28_368#
x_PM_SKY130_FD_SC_HS__O311AI_2%VPWR N_VPWR_M1009_d N_VPWR_M1006_d N_VPWR_M1010_d
+ N_VPWR_c_417_n N_VPWR_c_418_n N_VPWR_c_419_n N_VPWR_c_420_n N_VPWR_c_421_n
+ VPWR N_VPWR_c_422_n N_VPWR_c_423_n N_VPWR_c_416_n N_VPWR_c_425_n
+ N_VPWR_c_426_n PM_SKY130_FD_SC_HS__O311AI_2%VPWR
x_PM_SKY130_FD_SC_HS__O311AI_2%A_307_368# N_A_307_368#_M1007_d
+ N_A_307_368#_M1002_d N_A_307_368#_c_486_n N_A_307_368#_c_484_n
+ N_A_307_368#_c_485_n N_A_307_368#_c_505_p
+ PM_SKY130_FD_SC_HS__O311AI_2%A_307_368#
x_PM_SKY130_FD_SC_HS__O311AI_2%Y N_Y_M1001_s N_Y_M1011_s N_Y_M1002_s N_Y_M1004_s
+ N_Y_M1008_s N_Y_M1016_s N_Y_c_519_n N_Y_c_514_n N_Y_c_533_n N_Y_c_515_n
+ N_Y_c_510_n N_Y_c_553_n N_Y_c_516_n N_Y_c_517_n N_Y_c_511_n N_Y_c_518_n
+ N_Y_c_529_n N_Y_c_539_n Y Y Y Y PM_SKY130_FD_SC_HS__O311AI_2%Y
x_PM_SKY130_FD_SC_HS__O311AI_2%A_27_74# N_A_27_74#_M1000_d N_A_27_74#_M1019_d
+ N_A_27_74#_M1013_s N_A_27_74#_M1017_s N_A_27_74#_M1014_s N_A_27_74#_c_602_n
+ N_A_27_74#_c_603_n N_A_27_74#_c_604_n N_A_27_74#_c_605_n N_A_27_74#_c_606_n
+ N_A_27_74#_c_607_n N_A_27_74#_c_608_n N_A_27_74#_c_609_n N_A_27_74#_c_610_n
+ N_A_27_74#_c_611_n N_A_27_74#_c_612_n N_A_27_74#_c_613_n N_A_27_74#_c_614_n
+ PM_SKY130_FD_SC_HS__O311AI_2%A_27_74#
x_PM_SKY130_FD_SC_HS__O311AI_2%VGND N_VGND_M1000_s N_VGND_M1012_d N_VGND_M1005_d
+ N_VGND_c_683_n N_VGND_c_684_n N_VGND_c_685_n VGND N_VGND_c_686_n
+ N_VGND_c_687_n N_VGND_c_688_n N_VGND_c_689_n N_VGND_c_690_n N_VGND_c_691_n
+ N_VGND_c_692_n N_VGND_c_693_n PM_SKY130_FD_SC_HS__O311AI_2%VGND
x_PM_SKY130_FD_SC_HS__O311AI_2%A_670_74# N_A_670_74#_M1003_d N_A_670_74#_M1001_d
+ N_A_670_74#_c_765_n N_A_670_74#_c_750_n N_A_670_74#_c_751_n
+ N_A_670_74#_c_756_n PM_SKY130_FD_SC_HS__O311AI_2%A_670_74#
cc_1 VNB N_A1_M1000_g 0.0327337f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_2 VNB N_A1_M1019_g 0.0253298f $X=-0.19 $Y=-0.245 $X2=0.985 $Y2=0.74
cc_3 VNB A1 0.0167148f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_4 VNB N_A1_c_102_n 0.0404672f $X=-0.19 $Y=-0.245 $X2=0.97 $Y2=1.557
cc_5 VNB N_A2_M1012_g 0.0240209f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=2.4
cc_6 VNB N_A2_M1013_g 0.0237011f $X=-0.19 $Y=-0.245 $X2=0.97 $Y2=2.4
cc_7 VNB A2 0.0106647f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_A2_c_144_n 0.0351644f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.565
cc_9 VNB N_A3_M1005_g 0.0246497f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_10 VNB N_A3_M1017_g 0.0238365f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=2.4
cc_11 VNB N_A3_c_197_n 0.0138261f $X=-0.19 $Y=-0.245 $X2=0.985 $Y2=0.74
cc_12 VNB N_A3_c_198_n 0.0412386f $X=-0.19 $Y=-0.245 $X2=0.985 $Y2=0.74
cc_13 VNB A3 0.00488881f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_B1_c_257_n 0.0157815f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.35
cc_15 VNB N_B1_c_258_n 0.0203202f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_B1_c_259_n 0.00814437f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=1.765
cc_17 VNB N_B1_c_260_n 0.0179631f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=2.4
cc_18 VNB N_B1_c_261_n 0.0142118f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_19 VNB N_B1_c_262_n 0.0267906f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.557
cc_20 VNB B1 0.006035f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.515
cc_21 VNB N_B1_c_264_n 0.0170025f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.565
cc_22 VNB N_C1_M1001_g 0.0239843f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=2.4
cc_23 VNB N_C1_M1011_g 0.0291604f $X=-0.19 $Y=-0.245 $X2=0.985 $Y2=0.74
cc_24 VNB C1 0.0152566f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_25 VNB N_C1_c_330_n 0.0758738f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.515
cc_26 VNB N_VPWR_c_416_n 0.243291f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_Y_c_510_n 0.012331f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_Y_c_511_n 0.0247743f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB Y 0.0060107f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB Y 0.00619631f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_27_74#_c_602_n 0.0266107f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_27_74#_c_603_n 0.00612368f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=1.557
cc_33 VNB N_A_27_74#_c_604_n 0.00998227f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.557
cc_34 VNB N_A_27_74#_c_605_n 0.00253842f $X=-0.19 $Y=-0.245 $X2=0.97 $Y2=1.557
cc_35 VNB N_A_27_74#_c_606_n 0.0029209f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.565
cc_36 VNB N_A_27_74#_c_607_n 0.00253214f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.565
cc_37 VNB N_A_27_74#_c_608_n 0.00491768f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_27_74#_c_609_n 0.00206666f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_27_74#_c_610_n 0.00725544f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_27_74#_c_611_n 0.00351892f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_27_74#_c_612_n 0.00234762f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_27_74#_c_613_n 0.0028931f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_27_74#_c_614_n 0.00155944f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_683_n 0.00576795f $X=-0.19 $Y=-0.245 $X2=0.985 $Y2=0.74
cc_45 VNB N_VGND_c_684_n 0.00276855f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_46 VNB N_VGND_c_685_n 0.00563529f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=1.557
cc_47 VNB N_VGND_c_686_n 0.0173909f $X=-0.19 $Y=-0.245 $X2=0.97 $Y2=1.557
cc_48 VNB N_VGND_c_687_n 0.0188435f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.565
cc_49 VNB N_VGND_c_688_n 0.016883f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_VGND_c_689_n 0.0749446f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_VGND_c_690_n 0.326435f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_VGND_c_691_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_VGND_c_692_n 0.00604233f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_VGND_c_693_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_A_670_74#_c_750_n 0.0178206f $X=-0.19 $Y=-0.245 $X2=0.985 $Y2=1.35
cc_56 VNB N_A_670_74#_c_751_n 0.00417668f $X=-0.19 $Y=-0.245 $X2=0.985 $Y2=0.74
cc_57 VPB N_A1_c_103_n 0.0209395f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=1.765
cc_58 VPB N_A1_c_104_n 0.0157395f $X=-0.19 $Y=1.66 $X2=0.97 $Y2=1.765
cc_59 VPB A1 0.011263f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_60 VPB N_A1_c_102_n 0.0219936f $X=-0.19 $Y=1.66 $X2=0.97 $Y2=1.557
cc_61 VPB N_A2_c_145_n 0.0166076f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.35
cc_62 VPB N_A2_c_146_n 0.0191885f $X=-0.19 $Y=1.66 $X2=0.985 $Y2=0.74
cc_63 VPB A2 0.0106081f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_64 VPB N_A2_c_144_n 0.0221042f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=1.565
cc_65 VPB N_A3_c_200_n 0.0186669f $X=-0.19 $Y=1.66 $X2=0.97 $Y2=2.4
cc_66 VPB N_A3_c_197_n 0.013671f $X=-0.19 $Y=1.66 $X2=0.985 $Y2=0.74
cc_67 VPB N_A3_c_198_n 0.0306696f $X=-0.19 $Y=1.66 $X2=0.985 $Y2=0.74
cc_68 VPB N_A3_c_203_n 0.0158385f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_69 VPB A3 0.00821766f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_70 VPB N_B1_c_265_n 0.0153024f $X=-0.19 $Y=1.66 $X2=0.97 $Y2=2.4
cc_71 VPB N_B1_c_266_n 0.0149853f $X=-0.19 $Y=1.66 $X2=0.985 $Y2=0.74
cc_72 VPB N_B1_c_262_n 0.0198076f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.557
cc_73 VPB B1 0.00556484f $X=-0.19 $Y=1.66 $X2=0.585 $Y2=1.515
cc_74 VPB N_C1_c_331_n 0.0149852f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.35
cc_75 VPB N_C1_c_332_n 0.0208567f $X=-0.19 $Y=1.66 $X2=0.97 $Y2=1.765
cc_76 VPB C1 0.0109861f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_77 VPB N_C1_c_330_n 0.0131664f $X=-0.19 $Y=1.66 $X2=0.585 $Y2=1.515
cc_78 VPB N_A_28_368#_c_377_n 0.00739392f $X=-0.19 $Y=1.66 $X2=0.97 $Y2=2.4
cc_79 VPB N_A_28_368#_c_378_n 0.0353617f $X=-0.19 $Y=1.66 $X2=0.985 $Y2=0.74
cc_80 VPB N_A_28_368#_c_379_n 0.00289674f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_81 VPB N_A_28_368#_c_380_n 0.00735526f $X=-0.19 $Y=1.66 $X2=0.585 $Y2=1.565
cc_82 VPB N_VPWR_c_417_n 0.00581775f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_83 VPB N_VPWR_c_418_n 0.00329129f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_84 VPB N_VPWR_c_419_n 0.00504372f $X=-0.19 $Y=1.66 $X2=0.585 $Y2=1.515
cc_85 VPB N_VPWR_c_420_n 0.0164465f $X=-0.19 $Y=1.66 $X2=0.985 $Y2=1.557
cc_86 VPB N_VPWR_c_421_n 0.00460249f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=1.565
cc_87 VPB N_VPWR_c_422_n 0.0757972f $X=-0.19 $Y=1.66 $X2=0.585 $Y2=1.565
cc_88 VPB N_VPWR_c_423_n 0.0205835f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_89 VPB N_VPWR_c_416_n 0.0865852f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_90 VPB N_VPWR_c_425_n 0.024857f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_91 VPB N_VPWR_c_426_n 0.00601644f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_92 VPB N_A_307_368#_c_484_n 0.0200646f $X=-0.19 $Y=1.66 $X2=0.985 $Y2=1.35
cc_93 VPB N_A_307_368#_c_485_n 0.00400615f $X=-0.19 $Y=1.66 $X2=0.985 $Y2=0.74
cc_94 VPB N_Y_c_514_n 0.00216998f $X=-0.19 $Y=1.66 $X2=0.985 $Y2=1.557
cc_95 VPB N_Y_c_515_n 0.00180921f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_96 VPB N_Y_c_516_n 0.00723723f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_97 VPB N_Y_c_517_n 0.035396f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_98 VPB N_Y_c_518_n 0.00725308f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_99 N_A1_c_104_n N_A2_c_145_n 0.0107286f $X=0.97 $Y=1.765 $X2=-0.19 $Y2=-0.245
cc_100 N_A1_M1019_g N_A2_M1012_g 0.0179972f $X=0.985 $Y=0.74 $X2=0 $Y2=0
cc_101 A1 A2 0.0290771f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_102 N_A1_c_102_n A2 0.00529096f $X=0.97 $Y=1.557 $X2=0 $Y2=0
cc_103 A1 N_A2_c_144_n 2.03322e-19 $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_104 N_A1_c_102_n N_A2_c_144_n 0.0207993f $X=0.97 $Y=1.557 $X2=0 $Y2=0
cc_105 N_A1_c_103_n N_A_28_368#_c_377_n 4.27055e-19 $X=0.51 $Y=1.765 $X2=0 $Y2=0
cc_106 A1 N_A_28_368#_c_377_n 0.0260502f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_107 N_A1_c_103_n N_A_28_368#_c_378_n 0.0106409f $X=0.51 $Y=1.765 $X2=0 $Y2=0
cc_108 N_A1_c_104_n N_A_28_368#_c_378_n 6.58912e-19 $X=0.97 $Y=1.765 $X2=0 $Y2=0
cc_109 N_A1_c_103_n N_A_28_368#_c_385_n 0.012065f $X=0.51 $Y=1.765 $X2=0 $Y2=0
cc_110 N_A1_c_104_n N_A_28_368#_c_385_n 0.0175448f $X=0.97 $Y=1.765 $X2=0 $Y2=0
cc_111 A1 N_A_28_368#_c_385_n 0.0276588f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_112 N_A1_c_102_n N_A_28_368#_c_385_n 0.00222405f $X=0.97 $Y=1.557 $X2=0 $Y2=0
cc_113 N_A1_c_103_n N_VPWR_c_417_n 0.00527858f $X=0.51 $Y=1.765 $X2=0 $Y2=0
cc_114 N_A1_c_104_n N_VPWR_c_417_n 0.00930375f $X=0.97 $Y=1.765 $X2=0 $Y2=0
cc_115 N_A1_c_104_n N_VPWR_c_422_n 0.00444681f $X=0.97 $Y=1.765 $X2=0 $Y2=0
cc_116 N_A1_c_103_n N_VPWR_c_416_n 0.00861196f $X=0.51 $Y=1.765 $X2=0 $Y2=0
cc_117 N_A1_c_104_n N_VPWR_c_416_n 0.00878147f $X=0.97 $Y=1.765 $X2=0 $Y2=0
cc_118 N_A1_c_103_n N_VPWR_c_425_n 0.00445602f $X=0.51 $Y=1.765 $X2=0 $Y2=0
cc_119 N_A1_M1000_g N_A_27_74#_c_602_n 0.00159319f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_120 N_A1_M1000_g N_A_27_74#_c_603_n 0.013995f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_121 N_A1_M1019_g N_A_27_74#_c_603_n 0.018835f $X=0.985 $Y=0.74 $X2=0 $Y2=0
cc_122 A1 N_A_27_74#_c_603_n 0.0356901f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_123 N_A1_c_102_n N_A_27_74#_c_603_n 0.00358729f $X=0.97 $Y=1.557 $X2=0 $Y2=0
cc_124 A1 N_A_27_74#_c_604_n 0.0216404f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_125 N_A1_M1019_g N_A_27_74#_c_605_n 4.77375e-19 $X=0.985 $Y=0.74 $X2=0 $Y2=0
cc_126 N_A1_M1000_g N_VGND_c_683_n 0.0133418f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_127 N_A1_M1019_g N_VGND_c_683_n 0.00435015f $X=0.985 $Y=0.74 $X2=0 $Y2=0
cc_128 N_A1_M1019_g N_VGND_c_684_n 4.54333e-19 $X=0.985 $Y=0.74 $X2=0 $Y2=0
cc_129 N_A1_M1000_g N_VGND_c_686_n 0.00383152f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_130 N_A1_M1019_g N_VGND_c_687_n 0.00461464f $X=0.985 $Y=0.74 $X2=0 $Y2=0
cc_131 N_A1_M1000_g N_VGND_c_690_n 0.00761198f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_132 N_A1_M1019_g N_VGND_c_690_n 0.00909082f $X=0.985 $Y=0.74 $X2=0 $Y2=0
cc_133 N_A2_M1013_g N_A3_M1005_g 0.0164357f $X=1.915 $Y=0.74 $X2=0 $Y2=0
cc_134 A2 N_A3_c_198_n 0.00428545f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_135 N_A2_c_144_n N_A3_c_198_n 0.0205288f $X=1.915 $Y=1.557 $X2=0 $Y2=0
cc_136 A2 A3 0.0288737f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_137 N_A2_c_144_n A3 4.57332e-19 $X=1.915 $Y=1.557 $X2=0 $Y2=0
cc_138 N_A2_c_145_n N_A_28_368#_c_379_n 0.0104685f $X=1.46 $Y=1.765 $X2=0 $Y2=0
cc_139 N_A2_c_146_n N_A_28_368#_c_379_n 8.86279e-19 $X=1.98 $Y=1.765 $X2=0 $Y2=0
cc_140 N_A2_c_145_n N_A_28_368#_c_391_n 0.0123801f $X=1.46 $Y=1.765 $X2=0 $Y2=0
cc_141 N_A2_c_146_n N_A_28_368#_c_391_n 0.013058f $X=1.98 $Y=1.765 $X2=0 $Y2=0
cc_142 A2 N_A_28_368#_c_391_n 0.0491284f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_143 N_A2_c_144_n N_A_28_368#_c_391_n 0.00168607f $X=1.915 $Y=1.557 $X2=0
+ $Y2=0
cc_144 N_A2_c_145_n N_A_28_368#_c_395_n 4.27055e-19 $X=1.46 $Y=1.765 $X2=0 $Y2=0
cc_145 A2 N_A_28_368#_c_395_n 0.0243766f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_146 N_A2_c_146_n N_A_28_368#_c_380_n 0.0063565f $X=1.98 $Y=1.765 $X2=0 $Y2=0
cc_147 A2 N_A_28_368#_c_380_n 0.0137016f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_148 N_A2_c_145_n N_VPWR_c_417_n 6.85334e-19 $X=1.46 $Y=1.765 $X2=0 $Y2=0
cc_149 N_A2_c_145_n N_VPWR_c_422_n 0.00445602f $X=1.46 $Y=1.765 $X2=0 $Y2=0
cc_150 N_A2_c_146_n N_VPWR_c_422_n 0.00278257f $X=1.98 $Y=1.765 $X2=0 $Y2=0
cc_151 N_A2_c_145_n N_VPWR_c_416_n 0.00859416f $X=1.46 $Y=1.765 $X2=0 $Y2=0
cc_152 N_A2_c_146_n N_VPWR_c_416_n 0.00359257f $X=1.98 $Y=1.765 $X2=0 $Y2=0
cc_153 N_A2_c_146_n N_A_307_368#_c_486_n 0.0121561f $X=1.98 $Y=1.765 $X2=0 $Y2=0
cc_154 N_A2_c_146_n N_A_307_368#_c_484_n 0.012762f $X=1.98 $Y=1.765 $X2=0 $Y2=0
cc_155 N_A2_c_145_n N_A_307_368#_c_485_n 0.00359877f $X=1.46 $Y=1.765 $X2=0
+ $Y2=0
cc_156 N_A2_c_146_n N_A_307_368#_c_485_n 0.0017422f $X=1.98 $Y=1.765 $X2=0 $Y2=0
cc_157 A2 N_A_27_74#_c_603_n 0.0023919f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_158 N_A2_M1012_g N_A_27_74#_c_605_n 0.00348659f $X=1.475 $Y=0.74 $X2=0 $Y2=0
cc_159 N_A2_M1012_g N_A_27_74#_c_606_n 0.014989f $X=1.475 $Y=0.74 $X2=0 $Y2=0
cc_160 N_A2_M1013_g N_A_27_74#_c_606_n 0.0132249f $X=1.915 $Y=0.74 $X2=0 $Y2=0
cc_161 A2 N_A_27_74#_c_606_n 0.0511151f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_162 N_A2_c_144_n N_A_27_74#_c_606_n 0.00396531f $X=1.915 $Y=1.557 $X2=0 $Y2=0
cc_163 N_A2_M1013_g N_A_27_74#_c_607_n 4.39117e-19 $X=1.915 $Y=0.74 $X2=0 $Y2=0
cc_164 A2 N_A_27_74#_c_612_n 0.0225421f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_165 A2 N_A_27_74#_c_613_n 0.0206318f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_166 N_A2_c_144_n N_A_27_74#_c_613_n 6.38135e-19 $X=1.915 $Y=1.557 $X2=0 $Y2=0
cc_167 N_A2_M1012_g N_VGND_c_684_n 0.00983261f $X=1.475 $Y=0.74 $X2=0 $Y2=0
cc_168 N_A2_M1013_g N_VGND_c_684_n 0.0105836f $X=1.915 $Y=0.74 $X2=0 $Y2=0
cc_169 N_A2_M1012_g N_VGND_c_687_n 0.00413917f $X=1.475 $Y=0.74 $X2=0 $Y2=0
cc_170 N_A2_M1013_g N_VGND_c_688_n 0.00383152f $X=1.915 $Y=0.74 $X2=0 $Y2=0
cc_171 N_A2_M1012_g N_VGND_c_690_n 0.00818158f $X=1.475 $Y=0.74 $X2=0 $Y2=0
cc_172 N_A2_M1013_g N_VGND_c_690_n 0.00757998f $X=1.915 $Y=0.74 $X2=0 $Y2=0
cc_173 N_A3_M1017_g N_B1_c_257_n 0.0198315f $X=2.845 $Y=0.74 $X2=-0.19
+ $Y2=-0.245
cc_174 N_A3_c_197_n N_B1_c_259_n 0.0190635f $X=3.35 $Y=1.65 $X2=0 $Y2=0
cc_175 A3 N_B1_c_259_n 3.30527e-19 $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_176 N_A3_c_203_n N_B1_c_265_n 0.0122788f $X=3.44 $Y=1.765 $X2=0 $Y2=0
cc_177 N_A3_c_197_n N_B1_c_262_n 0.00984806f $X=3.35 $Y=1.65 $X2=0 $Y2=0
cc_178 N_A3_c_197_n B1 0.00652232f $X=3.35 $Y=1.65 $X2=0 $Y2=0
cc_179 N_A3_c_198_n B1 9.57942e-19 $X=3.08 $Y=1.65 $X2=0 $Y2=0
cc_180 N_A3_c_203_n B1 7.49256e-19 $X=3.44 $Y=1.765 $X2=0 $Y2=0
cc_181 A3 B1 0.0290571f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_182 A3 N_B1_c_264_n 9.7564e-19 $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_183 N_A3_c_200_n N_A_28_368#_c_380_n 0.00112319f $X=2.99 $Y=1.765 $X2=0 $Y2=0
cc_184 N_A3_c_198_n N_A_28_368#_c_380_n 0.00273636f $X=3.08 $Y=1.65 $X2=0 $Y2=0
cc_185 N_A3_c_203_n N_VPWR_c_418_n 5.91791e-19 $X=3.44 $Y=1.765 $X2=0 $Y2=0
cc_186 N_A3_c_200_n N_VPWR_c_422_n 0.00278271f $X=2.99 $Y=1.765 $X2=0 $Y2=0
cc_187 N_A3_c_203_n N_VPWR_c_422_n 0.00445602f $X=3.44 $Y=1.765 $X2=0 $Y2=0
cc_188 N_A3_c_200_n N_VPWR_c_416_n 0.00358624f $X=2.99 $Y=1.765 $X2=0 $Y2=0
cc_189 N_A3_c_203_n N_VPWR_c_416_n 0.00858435f $X=3.44 $Y=1.765 $X2=0 $Y2=0
cc_190 N_A3_c_200_n N_A_307_368#_c_484_n 0.0144245f $X=2.99 $Y=1.765 $X2=0 $Y2=0
cc_191 N_A3_c_203_n N_A_307_368#_c_484_n 0.001955f $X=3.44 $Y=1.765 $X2=0 $Y2=0
cc_192 N_A3_c_200_n N_Y_c_519_n 0.0120074f $X=2.99 $Y=1.765 $X2=0 $Y2=0
cc_193 N_A3_c_197_n N_Y_c_519_n 0.00387625f $X=3.35 $Y=1.65 $X2=0 $Y2=0
cc_194 N_A3_c_203_n N_Y_c_519_n 0.0126452f $X=3.44 $Y=1.765 $X2=0 $Y2=0
cc_195 A3 N_Y_c_519_n 0.0212867f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_196 N_A3_c_200_n N_Y_c_514_n 6.56812e-19 $X=2.99 $Y=1.765 $X2=0 $Y2=0
cc_197 N_A3_c_203_n N_Y_c_514_n 0.0102765f $X=3.44 $Y=1.765 $X2=0 $Y2=0
cc_198 N_A3_c_200_n N_Y_c_518_n 0.00941736f $X=2.99 $Y=1.765 $X2=0 $Y2=0
cc_199 N_A3_c_198_n N_Y_c_518_n 0.00192242f $X=3.08 $Y=1.65 $X2=0 $Y2=0
cc_200 N_A3_c_203_n N_Y_c_518_n 5.7112e-19 $X=3.44 $Y=1.765 $X2=0 $Y2=0
cc_201 A3 N_Y_c_518_n 0.0265005f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_202 N_A3_c_203_n N_Y_c_529_n 4.20803e-19 $X=3.44 $Y=1.765 $X2=0 $Y2=0
cc_203 N_A3_M1005_g N_A_27_74#_c_607_n 4.73925e-19 $X=2.385 $Y=0.74 $X2=0 $Y2=0
cc_204 N_A3_M1005_g N_A_27_74#_c_608_n 0.018337f $X=2.385 $Y=0.74 $X2=0 $Y2=0
cc_205 N_A3_M1017_g N_A_27_74#_c_608_n 0.0132506f $X=2.845 $Y=0.74 $X2=0 $Y2=0
cc_206 N_A3_c_198_n N_A_27_74#_c_608_n 0.00321928f $X=3.08 $Y=1.65 $X2=0 $Y2=0
cc_207 A3 N_A_27_74#_c_608_n 0.034156f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_208 N_A3_M1017_g N_A_27_74#_c_609_n 3.97481e-19 $X=2.845 $Y=0.74 $X2=0 $Y2=0
cc_209 N_A3_c_197_n N_A_27_74#_c_610_n 0.00213563f $X=3.35 $Y=1.65 $X2=0 $Y2=0
cc_210 A3 N_A_27_74#_c_610_n 7.38037e-19 $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_211 N_A3_c_198_n N_A_27_74#_c_614_n 0.00107191f $X=3.08 $Y=1.65 $X2=0 $Y2=0
cc_212 A3 N_A_27_74#_c_614_n 0.0224275f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_213 N_A3_M1005_g N_VGND_c_684_n 4.69274e-19 $X=2.385 $Y=0.74 $X2=0 $Y2=0
cc_214 N_A3_M1005_g N_VGND_c_685_n 0.00227662f $X=2.385 $Y=0.74 $X2=0 $Y2=0
cc_215 N_A3_M1017_g N_VGND_c_685_n 0.0103163f $X=2.845 $Y=0.74 $X2=0 $Y2=0
cc_216 N_A3_M1005_g N_VGND_c_688_n 0.00461464f $X=2.385 $Y=0.74 $X2=0 $Y2=0
cc_217 N_A3_M1017_g N_VGND_c_689_n 0.00383152f $X=2.845 $Y=0.74 $X2=0 $Y2=0
cc_218 N_A3_M1005_g N_VGND_c_690_n 0.00907963f $X=2.385 $Y=0.74 $X2=0 $Y2=0
cc_219 N_A3_M1017_g N_VGND_c_690_n 0.00757637f $X=2.845 $Y=0.74 $X2=0 $Y2=0
cc_220 N_B1_c_266_n N_C1_c_331_n 0.00943412f $X=4.34 $Y=1.765 $X2=-0.19
+ $Y2=-0.245
cc_221 N_B1_c_261_n N_C1_M1001_g 0.00126295f $X=3.935 $Y=1.26 $X2=0 $Y2=0
cc_222 N_B1_c_261_n N_C1_c_330_n 0.00317238f $X=3.935 $Y=1.26 $X2=0 $Y2=0
cc_223 N_B1_c_262_n N_C1_c_330_n 0.0111776f $X=3.935 $Y=1.53 $X2=0 $Y2=0
cc_224 B1 N_C1_c_330_n 5.56398e-19 $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_225 N_B1_c_265_n N_VPWR_c_418_n 0.0111808f $X=3.89 $Y=1.765 $X2=0 $Y2=0
cc_226 N_B1_c_266_n N_VPWR_c_418_n 0.0110266f $X=4.34 $Y=1.765 $X2=0 $Y2=0
cc_227 N_B1_c_266_n N_VPWR_c_419_n 5.37805e-19 $X=4.34 $Y=1.765 $X2=0 $Y2=0
cc_228 N_B1_c_266_n N_VPWR_c_420_n 0.00413917f $X=4.34 $Y=1.765 $X2=0 $Y2=0
cc_229 N_B1_c_265_n N_VPWR_c_422_n 0.00413917f $X=3.89 $Y=1.765 $X2=0 $Y2=0
cc_230 N_B1_c_265_n N_VPWR_c_416_n 0.0081781f $X=3.89 $Y=1.765 $X2=0 $Y2=0
cc_231 N_B1_c_266_n N_VPWR_c_416_n 0.0081781f $X=4.34 $Y=1.765 $X2=0 $Y2=0
cc_232 N_B1_c_258_n N_Y_c_519_n 4.321e-19 $X=3.77 $Y=1.26 $X2=0 $Y2=0
cc_233 B1 N_Y_c_519_n 0.00106056f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_234 N_B1_c_265_n N_Y_c_514_n 0.00605728f $X=3.89 $Y=1.765 $X2=0 $Y2=0
cc_235 N_B1_c_265_n N_Y_c_533_n 0.0126853f $X=3.89 $Y=1.765 $X2=0 $Y2=0
cc_236 N_B1_c_266_n N_Y_c_533_n 0.0152577f $X=4.34 $Y=1.765 $X2=0 $Y2=0
cc_237 N_B1_c_262_n N_Y_c_533_n 0.00213646f $X=3.935 $Y=1.53 $X2=0 $Y2=0
cc_238 B1 N_Y_c_533_n 0.0302312f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_239 N_B1_c_266_n N_Y_c_515_n 0.00576879f $X=4.34 $Y=1.765 $X2=0 $Y2=0
cc_240 B1 N_Y_c_529_n 0.0193938f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_241 N_B1_c_266_n N_Y_c_539_n 8.9901e-19 $X=4.34 $Y=1.765 $X2=0 $Y2=0
cc_242 N_B1_c_260_n Y 0.00117611f $X=3.845 $Y=1.185 $X2=0 $Y2=0
cc_243 N_B1_c_260_n Y 3.14144e-19 $X=3.845 $Y=1.185 $X2=0 $Y2=0
cc_244 N_B1_c_265_n Y 8.1906e-19 $X=3.89 $Y=1.765 $X2=0 $Y2=0
cc_245 N_B1_c_266_n Y 0.00407086f $X=4.34 $Y=1.765 $X2=0 $Y2=0
cc_246 N_B1_c_261_n Y 0.00415302f $X=3.935 $Y=1.26 $X2=0 $Y2=0
cc_247 N_B1_c_262_n Y 0.00755495f $X=3.935 $Y=1.53 $X2=0 $Y2=0
cc_248 B1 Y 0.031504f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_249 N_B1_c_264_n Y 6.27941e-19 $X=3.935 $Y=1.515 $X2=0 $Y2=0
cc_250 N_B1_c_257_n N_A_27_74#_c_609_n 0.00944442f $X=3.275 $Y=1.185 $X2=0 $Y2=0
cc_251 N_B1_c_260_n N_A_27_74#_c_609_n 6.66923e-19 $X=3.845 $Y=1.185 $X2=0 $Y2=0
cc_252 N_B1_c_257_n N_A_27_74#_c_610_n 0.011964f $X=3.275 $Y=1.185 $X2=0 $Y2=0
cc_253 N_B1_c_258_n N_A_27_74#_c_610_n 0.0063964f $X=3.77 $Y=1.26 $X2=0 $Y2=0
cc_254 N_B1_c_260_n N_A_27_74#_c_610_n 0.0129915f $X=3.845 $Y=1.185 $X2=0 $Y2=0
cc_255 N_B1_c_261_n N_A_27_74#_c_610_n 0.00564918f $X=3.935 $Y=1.26 $X2=0 $Y2=0
cc_256 N_B1_c_262_n N_A_27_74#_c_610_n 0.00148214f $X=3.935 $Y=1.53 $X2=0 $Y2=0
cc_257 B1 N_A_27_74#_c_610_n 0.0579009f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_258 N_B1_c_257_n N_A_27_74#_c_611_n 5.80141e-19 $X=3.275 $Y=1.185 $X2=0 $Y2=0
cc_259 N_B1_c_260_n N_A_27_74#_c_611_n 0.0077283f $X=3.845 $Y=1.185 $X2=0 $Y2=0
cc_260 N_B1_c_257_n N_A_27_74#_c_614_n 0.0014099f $X=3.275 $Y=1.185 $X2=0 $Y2=0
cc_261 N_B1_c_257_n N_VGND_c_685_n 5.57463e-19 $X=3.275 $Y=1.185 $X2=0 $Y2=0
cc_262 N_B1_c_257_n N_VGND_c_689_n 0.00434272f $X=3.275 $Y=1.185 $X2=0 $Y2=0
cc_263 N_B1_c_260_n N_VGND_c_689_n 0.00278271f $X=3.845 $Y=1.185 $X2=0 $Y2=0
cc_264 N_B1_c_257_n N_VGND_c_690_n 0.00822601f $X=3.275 $Y=1.185 $X2=0 $Y2=0
cc_265 N_B1_c_260_n N_VGND_c_690_n 0.00359661f $X=3.845 $Y=1.185 $X2=0 $Y2=0
cc_266 N_B1_c_260_n N_A_670_74#_c_750_n 0.0132715f $X=3.845 $Y=1.185 $X2=0 $Y2=0
cc_267 N_B1_c_257_n N_A_670_74#_c_751_n 0.00220721f $X=3.275 $Y=1.185 $X2=0
+ $Y2=0
cc_268 N_C1_c_331_n N_VPWR_c_418_n 5.35985e-19 $X=4.79 $Y=1.765 $X2=0 $Y2=0
cc_269 N_C1_c_331_n N_VPWR_c_419_n 0.0106464f $X=4.79 $Y=1.765 $X2=0 $Y2=0
cc_270 N_C1_c_332_n N_VPWR_c_419_n 0.00526215f $X=5.24 $Y=1.765 $X2=0 $Y2=0
cc_271 N_C1_c_331_n N_VPWR_c_420_n 0.00413917f $X=4.79 $Y=1.765 $X2=0 $Y2=0
cc_272 N_C1_c_332_n N_VPWR_c_423_n 0.00445602f $X=5.24 $Y=1.765 $X2=0 $Y2=0
cc_273 N_C1_c_331_n N_VPWR_c_416_n 0.0081781f $X=4.79 $Y=1.765 $X2=0 $Y2=0
cc_274 N_C1_c_332_n N_VPWR_c_416_n 0.00861133f $X=5.24 $Y=1.765 $X2=0 $Y2=0
cc_275 N_C1_c_331_n N_Y_c_515_n 0.0039133f $X=4.79 $Y=1.765 $X2=0 $Y2=0
cc_276 N_C1_M1001_g N_Y_c_510_n 0.015974f $X=4.835 $Y=0.74 $X2=0 $Y2=0
cc_277 N_C1_M1011_g N_Y_c_510_n 0.0126386f $X=5.265 $Y=0.74 $X2=0 $Y2=0
cc_278 C1 N_Y_c_510_n 0.0567145f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_279 N_C1_c_330_n N_Y_c_510_n 0.00935997f $X=5.265 $Y=1.532 $X2=0 $Y2=0
cc_280 N_C1_c_331_n N_Y_c_553_n 0.0156295f $X=4.79 $Y=1.765 $X2=0 $Y2=0
cc_281 N_C1_c_332_n N_Y_c_553_n 0.0120074f $X=5.24 $Y=1.765 $X2=0 $Y2=0
cc_282 C1 N_Y_c_553_n 0.027126f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_283 N_C1_c_330_n N_Y_c_553_n 0.00199349f $X=5.265 $Y=1.532 $X2=0 $Y2=0
cc_284 N_C1_c_332_n N_Y_c_516_n 4.27055e-19 $X=5.24 $Y=1.765 $X2=0 $Y2=0
cc_285 C1 N_Y_c_516_n 0.0267405f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_286 N_C1_c_330_n N_Y_c_516_n 0.00136954f $X=5.265 $Y=1.532 $X2=0 $Y2=0
cc_287 N_C1_c_331_n N_Y_c_517_n 6.69308e-19 $X=4.79 $Y=1.765 $X2=0 $Y2=0
cc_288 N_C1_c_332_n N_Y_c_517_n 0.0106911f $X=5.24 $Y=1.765 $X2=0 $Y2=0
cc_289 N_C1_M1011_g N_Y_c_511_n 0.00159289f $X=5.265 $Y=0.74 $X2=0 $Y2=0
cc_290 N_C1_c_331_n N_Y_c_539_n 8.9901e-19 $X=4.79 $Y=1.765 $X2=0 $Y2=0
cc_291 N_C1_c_331_n Y 0.00406785f $X=4.79 $Y=1.765 $X2=0 $Y2=0
cc_292 N_C1_M1001_g Y 0.0060753f $X=4.835 $Y=0.74 $X2=0 $Y2=0
cc_293 N_C1_c_332_n Y 8.18876e-19 $X=5.24 $Y=1.765 $X2=0 $Y2=0
cc_294 C1 Y 0.0349366f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_295 N_C1_c_330_n Y 0.0148268f $X=5.265 $Y=1.532 $X2=0 $Y2=0
cc_296 N_C1_M1001_g N_A_27_74#_c_610_n 4.45329e-19 $X=4.835 $Y=0.74 $X2=0 $Y2=0
cc_297 N_C1_M1001_g N_VGND_c_689_n 0.00278247f $X=4.835 $Y=0.74 $X2=0 $Y2=0
cc_298 N_C1_M1011_g N_VGND_c_689_n 0.00430908f $X=5.265 $Y=0.74 $X2=0 $Y2=0
cc_299 N_C1_M1001_g N_VGND_c_690_n 0.00358425f $X=4.835 $Y=0.74 $X2=0 $Y2=0
cc_300 N_C1_M1011_g N_VGND_c_690_n 0.00820326f $X=5.265 $Y=0.74 $X2=0 $Y2=0
cc_301 N_C1_M1001_g N_A_670_74#_c_750_n 0.0117594f $X=4.835 $Y=0.74 $X2=0 $Y2=0
cc_302 N_C1_M1011_g N_A_670_74#_c_750_n 0.00685665f $X=5.265 $Y=0.74 $X2=0 $Y2=0
cc_303 N_C1_M1001_g N_A_670_74#_c_756_n 0.0100975f $X=4.835 $Y=0.74 $X2=0 $Y2=0
cc_304 N_C1_M1011_g N_A_670_74#_c_756_n 0.00461693f $X=5.265 $Y=0.74 $X2=0 $Y2=0
cc_305 N_A_28_368#_c_385_n N_VPWR_M1009_d 0.00400851f $X=1.07 $Y=2.035 $X2=-0.19
+ $Y2=1.66
cc_306 N_A_28_368#_c_378_n N_VPWR_c_417_n 0.0462948f $X=0.285 $Y=2.815 $X2=0
+ $Y2=0
cc_307 N_A_28_368#_c_385_n N_VPWR_c_417_n 0.0154766f $X=1.07 $Y=2.035 $X2=0
+ $Y2=0
cc_308 N_A_28_368#_c_379_n N_VPWR_c_417_n 0.0256025f $X=1.235 $Y=2.815 $X2=0
+ $Y2=0
cc_309 N_A_28_368#_c_379_n N_VPWR_c_422_n 0.0145938f $X=1.235 $Y=2.815 $X2=0
+ $Y2=0
cc_310 N_A_28_368#_c_378_n N_VPWR_c_416_n 0.0120466f $X=0.285 $Y=2.815 $X2=0
+ $Y2=0
cc_311 N_A_28_368#_c_379_n N_VPWR_c_416_n 0.0120466f $X=1.235 $Y=2.815 $X2=0
+ $Y2=0
cc_312 N_A_28_368#_c_378_n N_VPWR_c_425_n 0.0145938f $X=0.285 $Y=2.815 $X2=0
+ $Y2=0
cc_313 N_A_28_368#_c_391_n N_A_307_368#_M1007_d 0.00503909f $X=2.12 $Y=2.035
+ $X2=-0.19 $Y2=1.66
cc_314 N_A_28_368#_c_391_n N_A_307_368#_c_486_n 0.0218521f $X=2.12 $Y=2.035
+ $X2=0 $Y2=0
cc_315 N_A_28_368#_c_380_n N_A_307_368#_c_486_n 0.0298377f $X=2.205 $Y=2.115
+ $X2=0 $Y2=0
cc_316 N_A_28_368#_M1015_s N_A_307_368#_c_484_n 0.00312144f $X=2.055 $Y=1.84
+ $X2=0 $Y2=0
cc_317 N_A_28_368#_c_380_n N_A_307_368#_c_484_n 0.018931f $X=2.205 $Y=2.115
+ $X2=0 $Y2=0
cc_318 N_A_28_368#_c_379_n N_A_307_368#_c_485_n 0.00340374f $X=1.235 $Y=2.815
+ $X2=0 $Y2=0
cc_319 N_A_28_368#_c_380_n N_Y_c_518_n 0.0534095f $X=2.205 $Y=2.115 $X2=0 $Y2=0
cc_320 N_VPWR_c_418_n N_A_307_368#_c_484_n 0.00286602f $X=4.115 $Y=2.455 $X2=0
+ $Y2=0
cc_321 N_VPWR_c_422_n N_A_307_368#_c_484_n 0.0892479f $X=3.95 $Y=3.33 $X2=0
+ $Y2=0
cc_322 N_VPWR_c_416_n N_A_307_368#_c_484_n 0.0507982f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_323 N_VPWR_c_422_n N_A_307_368#_c_485_n 0.0236039f $X=3.95 $Y=3.33 $X2=0
+ $Y2=0
cc_324 N_VPWR_c_416_n N_A_307_368#_c_485_n 0.012761f $X=5.52 $Y=3.33 $X2=0 $Y2=0
cc_325 N_VPWR_c_418_n N_Y_c_514_n 0.0462948f $X=4.115 $Y=2.455 $X2=0 $Y2=0
cc_326 N_VPWR_c_422_n N_Y_c_514_n 0.0110241f $X=3.95 $Y=3.33 $X2=0 $Y2=0
cc_327 N_VPWR_c_416_n N_Y_c_514_n 0.00909194f $X=5.52 $Y=3.33 $X2=0 $Y2=0
cc_328 N_VPWR_M1006_d N_Y_c_533_n 0.00364355f $X=3.965 $Y=1.84 $X2=0 $Y2=0
cc_329 N_VPWR_c_418_n N_Y_c_533_n 0.0171813f $X=4.115 $Y=2.455 $X2=0 $Y2=0
cc_330 N_VPWR_c_418_n N_Y_c_515_n 0.0449718f $X=4.115 $Y=2.455 $X2=0 $Y2=0
cc_331 N_VPWR_c_419_n N_Y_c_515_n 0.0440249f $X=5.015 $Y=2.455 $X2=0 $Y2=0
cc_332 N_VPWR_c_420_n N_Y_c_515_n 0.00749631f $X=4.85 $Y=3.33 $X2=0 $Y2=0
cc_333 N_VPWR_c_416_n N_Y_c_515_n 0.0062048f $X=5.52 $Y=3.33 $X2=0 $Y2=0
cc_334 N_VPWR_M1010_d N_Y_c_553_n 0.00384766f $X=4.865 $Y=1.84 $X2=0 $Y2=0
cc_335 N_VPWR_c_419_n N_Y_c_553_n 0.0154248f $X=5.015 $Y=2.455 $X2=0 $Y2=0
cc_336 N_VPWR_c_419_n N_Y_c_517_n 0.0462948f $X=5.015 $Y=2.455 $X2=0 $Y2=0
cc_337 N_VPWR_c_423_n N_Y_c_517_n 0.0145938f $X=5.52 $Y=3.33 $X2=0 $Y2=0
cc_338 N_VPWR_c_416_n N_Y_c_517_n 0.0120466f $X=5.52 $Y=3.33 $X2=0 $Y2=0
cc_339 N_A_307_368#_c_484_n N_Y_M1002_s 0.00287371f $X=3.13 $Y=2.99 $X2=0 $Y2=0
cc_340 N_A_307_368#_M1002_d N_Y_c_519_n 0.00431876f $X=3.065 $Y=1.84 $X2=0 $Y2=0
cc_341 N_A_307_368#_c_505_p N_Y_c_519_n 0.0136682f $X=3.215 $Y=2.455 $X2=0 $Y2=0
cc_342 N_A_307_368#_c_484_n N_Y_c_514_n 0.00539515f $X=3.13 $Y=2.99 $X2=0 $Y2=0
cc_343 N_A_307_368#_c_505_p N_Y_c_514_n 0.039183f $X=3.215 $Y=2.455 $X2=0 $Y2=0
cc_344 N_A_307_368#_c_484_n N_Y_c_518_n 0.0205764f $X=3.13 $Y=2.99 $X2=0 $Y2=0
cc_345 N_A_307_368#_c_505_p N_Y_c_518_n 0.0289859f $X=3.215 $Y=2.455 $X2=0 $Y2=0
cc_346 Y N_A_27_74#_c_610_n 0.011013f $X=4.475 $Y=0.84 $X2=0 $Y2=0
cc_347 Y N_A_27_74#_c_610_n 0.00429194f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_348 Y N_A_27_74#_c_611_n 0.0338529f $X=4.475 $Y=0.84 $X2=0 $Y2=0
cc_349 N_Y_c_511_n N_VGND_c_689_n 0.011066f $X=5.48 $Y=0.515 $X2=0 $Y2=0
cc_350 N_Y_c_511_n N_VGND_c_690_n 0.00915947f $X=5.48 $Y=0.515 $X2=0 $Y2=0
cc_351 N_Y_c_510_n N_A_670_74#_M1001_d 0.00176461f $X=5.395 $Y=1.045 $X2=0 $Y2=0
cc_352 N_Y_M1001_s N_A_670_74#_c_750_n 0.00273752f $X=4.475 $Y=0.37 $X2=0 $Y2=0
cc_353 N_Y_c_510_n N_A_670_74#_c_750_n 0.0032855f $X=5.395 $Y=1.045 $X2=0 $Y2=0
cc_354 N_Y_c_511_n N_A_670_74#_c_750_n 0.00374778f $X=5.48 $Y=0.515 $X2=0 $Y2=0
cc_355 Y N_A_670_74#_c_750_n 0.0232003f $X=4.475 $Y=0.84 $X2=0 $Y2=0
cc_356 N_Y_c_510_n N_A_670_74#_c_756_n 0.0168291f $X=5.395 $Y=1.045 $X2=0 $Y2=0
cc_357 N_A_27_74#_c_603_n N_VGND_M1000_s 0.00240242f $X=1.115 $Y=1.095 $X2=-0.19
+ $Y2=-0.245
cc_358 N_A_27_74#_c_606_n N_VGND_M1012_d 0.00187091f $X=2.045 $Y=1.095 $X2=0
+ $Y2=0
cc_359 N_A_27_74#_c_608_n N_VGND_M1005_d 0.00208352f $X=2.975 $Y=1.095 $X2=0
+ $Y2=0
cc_360 N_A_27_74#_c_602_n N_VGND_c_683_n 0.0182902f $X=0.28 $Y=0.515 $X2=0 $Y2=0
cc_361 N_A_27_74#_c_603_n N_VGND_c_683_n 0.0202152f $X=1.115 $Y=1.095 $X2=0
+ $Y2=0
cc_362 N_A_27_74#_c_605_n N_VGND_c_683_n 0.00121634f $X=1.2 $Y=0.515 $X2=0 $Y2=0
cc_363 N_A_27_74#_c_605_n N_VGND_c_684_n 0.0191439f $X=1.2 $Y=0.515 $X2=0 $Y2=0
cc_364 N_A_27_74#_c_606_n N_VGND_c_684_n 0.0172138f $X=2.045 $Y=1.095 $X2=0
+ $Y2=0
cc_365 N_A_27_74#_c_607_n N_VGND_c_684_n 0.0182902f $X=2.13 $Y=0.515 $X2=0 $Y2=0
cc_366 N_A_27_74#_c_607_n N_VGND_c_685_n 0.00154841f $X=2.13 $Y=0.515 $X2=0
+ $Y2=0
cc_367 N_A_27_74#_c_608_n N_VGND_c_685_n 0.0177745f $X=2.975 $Y=1.095 $X2=0
+ $Y2=0
cc_368 N_A_27_74#_c_609_n N_VGND_c_685_n 0.0182902f $X=3.06 $Y=0.515 $X2=0 $Y2=0
cc_369 N_A_27_74#_c_602_n N_VGND_c_686_n 0.011066f $X=0.28 $Y=0.515 $X2=0 $Y2=0
cc_370 N_A_27_74#_c_605_n N_VGND_c_687_n 0.011066f $X=1.2 $Y=0.515 $X2=0 $Y2=0
cc_371 N_A_27_74#_c_607_n N_VGND_c_688_n 0.011066f $X=2.13 $Y=0.515 $X2=0 $Y2=0
cc_372 N_A_27_74#_c_609_n N_VGND_c_689_n 0.0109942f $X=3.06 $Y=0.515 $X2=0 $Y2=0
cc_373 N_A_27_74#_c_602_n N_VGND_c_690_n 0.00915947f $X=0.28 $Y=0.515 $X2=0
+ $Y2=0
cc_374 N_A_27_74#_c_605_n N_VGND_c_690_n 0.00915947f $X=1.2 $Y=0.515 $X2=0 $Y2=0
cc_375 N_A_27_74#_c_607_n N_VGND_c_690_n 0.00915947f $X=2.13 $Y=0.515 $X2=0
+ $Y2=0
cc_376 N_A_27_74#_c_609_n N_VGND_c_690_n 0.00904371f $X=3.06 $Y=0.515 $X2=0
+ $Y2=0
cc_377 N_A_27_74#_c_610_n N_A_670_74#_M1003_d 0.00358162f $X=3.895 $Y=1.095
+ $X2=-0.19 $Y2=-0.245
cc_378 N_A_27_74#_c_610_n N_A_670_74#_c_765_n 0.0245925f $X=3.895 $Y=1.095 $X2=0
+ $Y2=0
cc_379 N_A_27_74#_M1014_s N_A_670_74#_c_750_n 0.00273752f $X=3.92 $Y=0.37 $X2=0
+ $Y2=0
cc_380 N_A_27_74#_c_610_n N_A_670_74#_c_750_n 0.00304353f $X=3.895 $Y=1.095
+ $X2=0 $Y2=0
cc_381 N_A_27_74#_c_611_n N_A_670_74#_c_750_n 0.0203278f $X=4.06 $Y=0.86 $X2=0
+ $Y2=0
cc_382 N_A_27_74#_c_609_n N_A_670_74#_c_751_n 0.00359554f $X=3.06 $Y=0.515 $X2=0
+ $Y2=0
cc_383 N_VGND_c_689_n N_A_670_74#_c_750_n 0.096935f $X=5.52 $Y=0 $X2=0 $Y2=0
cc_384 N_VGND_c_690_n N_A_670_74#_c_750_n 0.0548766f $X=5.52 $Y=0 $X2=0 $Y2=0
cc_385 N_VGND_c_685_n N_A_670_74#_c_751_n 0.00306547f $X=2.63 $Y=0.595 $X2=0
+ $Y2=0
cc_386 N_VGND_c_689_n N_A_670_74#_c_751_n 0.023391f $X=5.52 $Y=0 $X2=0 $Y2=0
cc_387 N_VGND_c_690_n N_A_670_74#_c_751_n 0.0127797f $X=5.52 $Y=0 $X2=0 $Y2=0
