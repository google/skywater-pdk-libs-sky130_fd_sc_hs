* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hs__a31o_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
M1000 a_529_392# B1 a_83_274# VPB pshort w=1e+06u l=150000u
+  ad=1.69e+12p pd=1.338e+07u as=3.7e+11p ps=2.74e+06u
M1001 a_529_392# A3 VPWR VPB pshort w=1e+06u l=150000u
+  ad=0p pd=0u as=2.3248e+12p ps=1.712e+07u
M1002 a_83_274# B1 VGND VNB nlowvt w=640000u l=150000u
+  ad=5.888e+11p pd=5.68e+06u as=1.0507e+12p ps=1.001e+07u
M1003 VGND A3 a_1000_74# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=5.44e+11p ps=5.54e+06u
M1004 a_529_392# A2 VPWR VPB pshort w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VPWR A3 a_529_392# VPB pshort w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_775_74# A2 a_1000_74# VNB nlowvt w=640000u l=150000u
+  ad=4.032e+11p pd=3.82e+06u as=0p ps=0u
M1007 VGND B1 a_83_274# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 X a_83_274# VGND VNB nlowvt w=740000u l=150000u
+  ad=4.662e+11p pd=4.22e+06u as=0p ps=0u
M1009 VGND a_83_274# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 X a_83_274# VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=6.72e+11p pd=5.68e+06u as=0p ps=0u
M1011 a_83_274# A1 a_775_74# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VPWR a_83_274# X VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_775_74# A1 a_83_274# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_1000_74# A3 VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VPWR a_83_274# X VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_529_392# A1 VPWR VPB pshort w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 X a_83_274# VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_1000_74# A2 a_775_74# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VGND a_83_274# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_83_274# B1 a_529_392# VPB pshort w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 VPWR A1 a_529_392# VPB pshort w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 X a_83_274# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 VPWR A2 a_529_392# VPB pshort w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
