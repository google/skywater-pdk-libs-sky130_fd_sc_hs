* File: sky130_fd_sc_hs__and4b_4.pex.spice
* Created: Thu Aug 27 20:33:40 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HS__AND4B_4%A_N 1 3 4 6 7
r32 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.59
+ $Y=1.385 $X2=0.59 $Y2=1.385
r33 7 11 4.1616 $w=3.58e-07 $l=1.3e-07 $layer=LI1_cond $X=0.72 $Y=1.37 $X2=0.59
+ $Y2=1.37
r34 4 10 38.7914 $w=2.76e-07 $l=1.88348e-07 $layer=POLY_cond $X=0.535 $Y=1.22
+ $X2=0.585 $Y2=1.385
r35 4 6 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=0.535 $Y=1.22
+ $X2=0.535 $Y2=0.79
r36 1 10 76.3385 $w=2.76e-07 $l=4.18091e-07 $layer=POLY_cond $X=0.505 $Y=1.765
+ $X2=0.585 $Y2=1.385
r37 1 3 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=0.505 $Y=1.765
+ $X2=0.505 $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_HS__AND4B_4%A_199_294# 1 2 3 4 5 16 18 21 23 27 29 31 32
+ 34 37 39 41 44 47 56 57 58 65 66 69 71 74 76 86
c154 76 0 4.33893e-19 $X=6.08 $Y=2.08
c155 74 0 1.24153e-19 $X=5.65 $Y=2.08
c156 71 0 8.61189e-20 $X=3.515 $Y=2.085
c157 56 0 5.40706e-20 $X=2.66 $Y=1.95
c158 39 0 4.4621e-20 $X=2.575 $Y=1.765
r159 86 87 1.90263 $w=3.8e-07 $l=1.5e-08 $layer=POLY_cond $X=2.575 $Y=1.542
+ $X2=2.59 $Y2=1.542
r160 83 84 18.3921 $w=3.8e-07 $l=1.45e-07 $layer=POLY_cond $X=2.015 $Y=1.542
+ $X2=2.16 $Y2=1.542
r161 80 81 1.90263 $w=3.8e-07 $l=1.5e-08 $layer=POLY_cond $X=1.52 $Y=1.542
+ $X2=1.535 $Y2=1.542
r162 75 76 3.65747 $w=2.78e-07 $l=8.5e-08 $layer=LI1_cond $X=5.995 $Y=2.08
+ $X2=6.08 $Y2=2.08
r163 73 75 7.40856 $w=2.78e-07 $l=1.8e-07 $layer=LI1_cond $X=5.815 $Y=2.08
+ $X2=5.995 $Y2=2.08
r164 73 74 6.95017 $w=2.78e-07 $l=1.65e-07 $layer=LI1_cond $X=5.815 $Y=2.08
+ $X2=5.65 $Y2=2.08
r165 69 76 29.2721 $w=2.48e-07 $l=6.35e-07 $layer=LI1_cond $X=6.715 $Y=2.095
+ $X2=6.08 $Y2=2.095
r166 66 75 3.65648 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=5.995 $Y=1.94
+ $X2=5.995 $Y2=2.08
r167 65 79 10.8397 $w=2.87e-07 $l=3.34201e-07 $layer=LI1_cond $X=5.995 $Y=1.3
+ $X2=6.25 $Y2=1.117
r168 65 66 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=5.995 $Y=1.3
+ $X2=5.995 $Y2=1.94
r169 64 74 34.8038 $w=2.48e-07 $l=7.55e-07 $layer=LI1_cond $X=4.895 $Y=2.095
+ $X2=5.65 $Y2=2.095
r170 64 71 63.6149 $w=2.48e-07 $l=1.38e-06 $layer=LI1_cond $X=4.895 $Y=2.095
+ $X2=3.515 $Y2=2.095
r171 58 60 25.8233 $w=2.68e-07 $l=6.05e-07 $layer=LI1_cond $X=2.745 $Y=2.085
+ $X2=3.35 $Y2=2.085
r172 57 71 5.8439 $w=2.68e-07 $l=1.35e-07 $layer=LI1_cond $X=3.38 $Y=2.085
+ $X2=3.515 $Y2=2.085
r173 57 60 1.28049 $w=2.68e-07 $l=3e-08 $layer=LI1_cond $X=3.38 $Y=2.085
+ $X2=3.35 $Y2=2.085
r174 56 58 7.28469 $w=2.7e-07 $l=1.72337e-07 $layer=LI1_cond $X=2.66 $Y=1.95
+ $X2=2.745 $Y2=2.085
r175 55 56 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=2.66 $Y=1.65 $X2=2.66
+ $Y2=1.95
r176 54 86 31.0763 $w=3.8e-07 $l=2.45e-07 $layer=POLY_cond $X=2.33 $Y=1.542
+ $X2=2.575 $Y2=1.542
r177 54 84 21.5632 $w=3.8e-07 $l=1.7e-07 $layer=POLY_cond $X=2.33 $Y=1.542
+ $X2=2.16 $Y2=1.542
r178 53 54 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=2.33
+ $Y=1.485 $X2=2.33 $Y2=1.485
r179 50 83 46.2974 $w=3.8e-07 $l=3.65e-07 $layer=POLY_cond $X=1.65 $Y=1.542
+ $X2=2.015 $Y2=1.542
r180 50 81 14.5868 $w=3.8e-07 $l=1.15e-07 $layer=POLY_cond $X=1.65 $Y=1.542
+ $X2=1.535 $Y2=1.542
r181 49 53 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=1.65 $Y=1.485
+ $X2=2.33 $Y2=1.485
r182 49 50 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.65
+ $Y=1.485 $X2=1.65 $Y2=1.485
r183 47 55 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.575 $Y=1.485
+ $X2=2.66 $Y2=1.65
r184 47 53 8.55602 $w=3.28e-07 $l=2.45e-07 $layer=LI1_cond $X=2.575 $Y=1.485
+ $X2=2.33 $Y2=1.485
r185 42 87 24.6126 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=2.59 $Y=1.32
+ $X2=2.59 $Y2=1.542
r186 42 44 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=2.59 $Y=1.32
+ $X2=2.59 $Y2=0.74
r187 39 86 24.6126 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=2.575 $Y=1.765
+ $X2=2.575 $Y2=1.542
r188 39 41 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.575 $Y=1.765
+ $X2=2.575 $Y2=2.4
r189 35 84 24.6126 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=2.16 $Y=1.32
+ $X2=2.16 $Y2=1.542
r190 35 37 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=2.16 $Y=1.32
+ $X2=2.16 $Y2=0.74
r191 32 83 24.6126 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=2.015 $Y=1.765
+ $X2=2.015 $Y2=1.542
r192 32 34 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.015 $Y=1.765
+ $X2=2.015 $Y2=2.4
r193 29 81 24.6126 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=1.535 $Y=1.765
+ $X2=1.535 $Y2=1.542
r194 29 31 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.535 $Y=1.765
+ $X2=1.535 $Y2=2.4
r195 25 80 24.6126 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=1.52 $Y=1.32
+ $X2=1.52 $Y2=1.542
r196 25 27 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=1.52 $Y=1.32
+ $X2=1.52 $Y2=0.74
r197 24 46 6.21277 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=1.175 $Y=1.395
+ $X2=1.085 $Y2=1.395
r198 23 80 27.8023 $w=3.8e-07 $l=1.80649e-07 $layer=POLY_cond $X=1.445 $Y=1.395
+ $X2=1.52 $Y2=1.542
r199 23 24 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=1.445 $Y=1.395
+ $X2=1.175 $Y2=1.395
r200 19 46 21.8783 $w=1.73e-07 $l=7.74597e-08 $layer=POLY_cond $X=1.09 $Y=1.32
+ $X2=1.085 $Y2=1.395
r201 19 21 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=1.09 $Y=1.32
+ $X2=1.09 $Y2=0.74
r202 16 46 104.069 $w=1.73e-07 $l=3.7e-07 $layer=POLY_cond $X=1.085 $Y=1.765
+ $X2=1.085 $Y2=1.395
r203 16 18 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.085 $Y=1.765
+ $X2=1.085 $Y2=2.4
r204 5 69 600 $w=1.7e-07 $l=2.38485e-07 $layer=licon1_PDIFF $count=1 $X=6.565
+ $Y=1.96 $X2=6.715 $Y2=2.135
r205 4 73 600 $w=1.7e-07 $l=2.22711e-07 $layer=licon1_PDIFF $count=1 $X=5.665
+ $Y=1.96 $X2=5.815 $Y2=2.12
r206 3 64 300 $w=1.7e-07 $l=7.92685e-07 $layer=licon1_PDIFF $count=2 $X=4.185
+ $Y=1.96 $X2=4.895 $Y2=2.135
r207 2 60 600 $w=1.7e-07 $l=2.2798e-07 $layer=licon1_PDIFF $count=1 $X=3.2
+ $Y=1.96 $X2=3.35 $Y2=2.125
r208 1 79 182 $w=1.7e-07 $l=5.50568e-07 $layer=licon1_NDIFF $count=1 $X=6.11
+ $Y=0.625 $X2=6.25 $Y2=1.11
.ends

.subckt PM_SKY130_FD_SC_HS__AND4B_4%D 1 3 4 6 8 9 11 12 14 15 17 18 19 26
c60 6 0 8.61189e-20 $X=4.11 $Y=1.885
r61 26 28 18.1887 $w=4.24e-07 $l=1.6e-07 $layer=POLY_cond $X=4.585 $Y=1.615
+ $X2=4.745 $Y2=1.615
r62 24 26 48.8821 $w=4.24e-07 $l=4.3e-07 $layer=POLY_cond $X=4.155 $Y=1.615
+ $X2=4.585 $Y2=1.615
r63 23 24 5.11557 $w=4.24e-07 $l=4.5e-08 $layer=POLY_cond $X=4.11 $Y=1.615
+ $X2=4.155 $Y2=1.615
r64 18 19 16.7628 $w=3.28e-07 $l=4.8e-07 $layer=LI1_cond $X=4.56 $Y=1.635
+ $X2=5.04 $Y2=1.635
r65 18 26 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.585
+ $Y=1.635 $X2=4.585 $Y2=1.635
r66 17 18 16.7628 $w=3.28e-07 $l=4.8e-07 $layer=LI1_cond $X=4.08 $Y=1.635
+ $X2=4.56 $Y2=1.635
r67 12 28 27.2926 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=4.745 $Y=1.345
+ $X2=4.745 $Y2=1.615
r68 12 14 128.533 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=4.745 $Y=1.345
+ $X2=4.745 $Y2=0.945
r69 9 24 27.2926 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=4.155 $Y=1.345
+ $X2=4.155 $Y2=1.615
r70 9 11 128.533 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=4.155 $Y=1.345
+ $X2=4.155 $Y2=0.945
r71 6 23 27.2926 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=4.11 $Y=1.885
+ $X2=4.11 $Y2=1.615
r72 6 8 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=4.11 $Y=1.885
+ $X2=4.11 $Y2=2.46
r73 5 15 7.1379 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=3.665 $Y=1.725 $X2=3.575
+ $Y2=1.725
r74 4 23 31.5592 $w=4.24e-07 $l=1.48324e-07 $layer=POLY_cond $X=4.02 $Y=1.725
+ $X2=4.11 $Y2=1.615
r75 4 5 182.032 $w=1.5e-07 $l=3.55e-07 $layer=POLY_cond $X=4.02 $Y=1.725
+ $X2=3.665 $Y2=1.725
r76 1 15 64.3434 $w=1.8e-07 $l=1.6e-07 $layer=POLY_cond $X=3.575 $Y=1.885
+ $X2=3.575 $Y2=1.725
r77 1 3 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=3.575 $Y=1.885
+ $X2=3.575 $Y2=2.46
.ends

.subckt PM_SKY130_FD_SC_HS__AND4B_4%C 1 3 5 6 7 10 12 14 16 22 23 24 26 27 31
c81 31 0 4.4621e-20 $X=3.08 $Y=1.515
c82 14 0 2.5326e-19 $X=5.12 $Y=1.885
c83 10 0 1.24153e-19 $X=3.68 $Y=0.945
c84 5 0 1.18606e-19 $X=3.17 $Y=1.35
r85 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.08
+ $Y=1.515 $X2=3.08 $Y2=1.515
r86 27 31 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=3.08 $Y=1.665
+ $X2=3.08 $Y2=1.515
r87 25 26 53.9552 $w=1.9e-07 $l=1.5e-07 $layer=POLY_cond $X=5.155 $Y=1.34
+ $X2=5.155 $Y2=1.49
r88 24 26 125.628 $w=1.5e-07 $l=2.45e-07 $layer=POLY_cond $X=5.135 $Y=1.735
+ $X2=5.135 $Y2=1.49
r89 22 25 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=5.175 $Y=0.945
+ $X2=5.175 $Y2=1.34
r90 19 22 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=5.175 $Y=0.255
+ $X2=5.175 $Y2=0.945
r91 14 24 58.3064 $w=1.8e-07 $l=1.5e-07 $layer=POLY_cond $X=5.12 $Y=1.885
+ $X2=5.12 $Y2=1.735
r92 14 16 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=5.12 $Y=1.885
+ $X2=5.12 $Y2=2.46
r93 13 23 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.755 $Y=0.18
+ $X2=3.68 $Y2=0.18
r94 12 19 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.1 $Y=0.18
+ $X2=5.175 $Y2=0.255
r95 12 13 689.67 $w=1.5e-07 $l=1.345e-06 $layer=POLY_cond $X=5.1 $Y=0.18
+ $X2=3.755 $Y2=0.18
r96 8 23 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.68 $Y=0.255
+ $X2=3.68 $Y2=0.18
r97 8 10 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=3.68 $Y=0.255
+ $X2=3.68 $Y2=0.945
r98 6 23 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.605 $Y=0.18
+ $X2=3.68 $Y2=0.18
r99 6 7 184.596 $w=1.5e-07 $l=3.6e-07 $layer=POLY_cond $X=3.605 $Y=0.18
+ $X2=3.245 $Y2=0.18
r100 5 30 38.8629 $w=2.72e-07 $l=2.05122e-07 $layer=POLY_cond $X=3.17 $Y=1.35
+ $X2=3.08 $Y2=1.515
r101 4 7 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.17 $Y=0.255
+ $X2=3.245 $Y2=0.18
r102 4 5 561.479 $w=1.5e-07 $l=1.095e-06 $layer=POLY_cond $X=3.17 $Y=0.255
+ $X2=3.17 $Y2=1.35
r103 1 30 75.1901 $w=2.72e-07 $l=3.91855e-07 $layer=POLY_cond $X=3.125 $Y=1.885
+ $X2=3.08 $Y2=1.515
r104 1 3 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=3.125 $Y=1.885
+ $X2=3.125 $Y2=2.46
.ends

.subckt PM_SKY130_FD_SC_HS__AND4B_4%A_27_368# 1 2 9 11 13 16 18 20 21 27 28 31
+ 32 33 35 36 38 39 40 48 53
c133 53 0 1.31377e-19 $X=6.465 $Y=1.677
c134 18 0 1.66257e-19 $X=6.49 $Y=1.885
c135 9 0 5.7483e-20 $X=6.035 $Y=0.945
r136 53 54 3.20479 $w=3.76e-07 $l=2.5e-08 $layer=POLY_cond $X=6.465 $Y=1.677
+ $X2=6.49 $Y2=1.677
r137 50 51 0.640957 $w=3.76e-07 $l=5e-09 $layer=POLY_cond $X=6.035 $Y=1.677
+ $X2=6.04 $Y2=1.677
r138 46 53 6.40957 $w=3.76e-07 $l=5e-08 $layer=POLY_cond $X=6.415 $Y=1.677
+ $X2=6.465 $Y2=1.677
r139 46 51 48.0718 $w=3.76e-07 $l=3.75e-07 $layer=POLY_cond $X=6.415 $Y=1.677
+ $X2=6.04 $Y2=1.677
r140 45 48 6.11144 $w=3.28e-07 $l=1.75e-07 $layer=LI1_cond $X=6.415 $Y=1.635
+ $X2=6.59 $Y2=1.635
r141 45 46 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.415
+ $Y=1.635 $X2=6.415 $Y2=1.635
r142 40 42 7.04271 $w=3.58e-07 $l=2.2e-07 $layer=LI1_cond $X=0.265 $Y=2.475
+ $X2=0.265 $Y2=2.695
r143 38 39 8.51103 $w=3.58e-07 $l=1.65e-07 $layer=LI1_cond $X=0.265 $Y=1.985
+ $X2=0.265 $Y2=1.82
r144 36 39 52.1925 $w=1.68e-07 $l=8e-07 $layer=LI1_cond $X=0.17 $Y=1.02 $X2=0.17
+ $Y2=1.82
r145 34 35 71.1123 $w=1.68e-07 $l=1.09e-06 $layer=LI1_cond $X=7.435 $Y=1.3
+ $X2=7.435 $Y2=2.39
r146 32 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.35 $Y=1.215
+ $X2=7.435 $Y2=1.3
r147 32 33 44.0374 $w=1.68e-07 $l=6.75e-07 $layer=LI1_cond $X=7.35 $Y=1.215
+ $X2=6.675 $Y2=1.215
r148 31 48 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.59 $Y=1.47
+ $X2=6.59 $Y2=1.635
r149 30 33 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.59 $Y=1.3
+ $X2=6.675 $Y2=1.215
r150 30 31 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=6.59 $Y=1.3
+ $X2=6.59 $Y2=1.47
r151 29 40 5.14255 $w=1.7e-07 $l=1.8e-07 $layer=LI1_cond $X=0.445 $Y=2.475
+ $X2=0.265 $Y2=2.475
r152 28 35 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.35 $Y=2.475
+ $X2=7.435 $Y2=2.39
r153 28 29 450.487 $w=1.68e-07 $l=6.905e-06 $layer=LI1_cond $X=7.35 $Y=2.475
+ $X2=0.445 $Y2=2.475
r154 27 40 2.72105 $w=3.58e-07 $l=8.5e-08 $layer=LI1_cond $X=0.265 $Y=2.39
+ $X2=0.265 $Y2=2.475
r155 26 38 0.480185 $w=3.58e-07 $l=1.5e-08 $layer=LI1_cond $X=0.265 $Y=2
+ $X2=0.265 $Y2=1.985
r156 26 27 12.4848 $w=3.58e-07 $l=3.9e-07 $layer=LI1_cond $X=0.265 $Y=2
+ $X2=0.265 $Y2=2.39
r157 21 36 8.28018 $w=3.18e-07 $l=1.6e-07 $layer=LI1_cond $X=0.245 $Y=0.86
+ $X2=0.245 $Y2=1.02
r158 21 23 4.38438 $w=3.2e-07 $l=1.15e-07 $layer=LI1_cond $X=0.245 $Y=0.86
+ $X2=0.245 $Y2=0.745
r159 18 54 24.356 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=6.49 $Y=1.885
+ $X2=6.49 $Y2=1.677
r160 18 20 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=6.49 $Y=1.885
+ $X2=6.49 $Y2=2.46
r161 14 53 24.356 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=6.465 $Y=1.47
+ $X2=6.465 $Y2=1.677
r162 14 16 269.202 $w=1.5e-07 $l=5.25e-07 $layer=POLY_cond $X=6.465 $Y=1.47
+ $X2=6.465 $Y2=0.945
r163 11 51 24.356 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=6.04 $Y=1.885
+ $X2=6.04 $Y2=1.677
r164 11 13 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=6.04 $Y=1.885
+ $X2=6.04 $Y2=2.46
r165 7 50 24.356 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=6.035 $Y=1.47
+ $X2=6.035 $Y2=1.677
r166 7 9 269.202 $w=1.5e-07 $l=5.25e-07 $layer=POLY_cond $X=6.035 $Y=1.47
+ $X2=6.035 $Y2=0.945
r167 2 42 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.695
r168 2 38 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=1.985
r169 1 23 182 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_NDIFF $count=1 $X=0.175
+ $Y=0.47 $X2=0.32 $Y2=0.745
.ends

.subckt PM_SKY130_FD_SC_HS__AND4B_4%B 1 2 3 5 9 10 11 12 14 18 20
c66 9 0 2.3468e-20 $X=5.605 $Y=0.945
r67 20 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.015
+ $Y=1.635 $X2=7.015 $Y2=1.635
r68 16 23 38.5336 $w=3.07e-07 $l=2.07123e-07 $layer=POLY_cond $X=7.115 $Y=1.47
+ $X2=7.02 $Y2=1.635
r69 16 18 269.202 $w=1.5e-07 $l=5.25e-07 $layer=POLY_cond $X=7.115 $Y=1.47
+ $X2=7.115 $Y2=0.945
r70 15 18 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=7.115 $Y=0.255
+ $X2=7.115 $Y2=0.945
r71 12 23 51.8789 $w=3.07e-07 $l=2.87228e-07 $layer=POLY_cond $X=6.94 $Y=1.885
+ $X2=7.02 $Y2=1.635
r72 12 14 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=6.94 $Y=1.885
+ $X2=6.94 $Y2=2.46
r73 10 15 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=7.04 $Y=0.18
+ $X2=7.115 $Y2=0.255
r74 10 11 697.362 $w=1.5e-07 $l=1.36e-06 $layer=POLY_cond $X=7.04 $Y=0.18
+ $X2=5.68 $Y2=0.18
r75 9 19 230.745 $w=1.5e-07 $l=4.5e-07 $layer=POLY_cond $X=5.605 $Y=0.945
+ $X2=5.605 $Y2=1.395
r76 6 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.605 $Y=0.255
+ $X2=5.68 $Y2=0.18
r77 6 9 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=5.605 $Y=0.255
+ $X2=5.605 $Y2=0.945
r78 3 5 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=5.59 $Y=1.885
+ $X2=5.59 $Y2=2.46
r79 2 3 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=5.59 $Y=1.795 $X2=5.59
+ $Y2=1.885
r80 1 19 37.1337 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=5.59 $Y=1.485 $X2=5.59
+ $Y2=1.395
r81 1 2 120.5 $w=1.8e-07 $l=3.1e-07 $layer=POLY_cond $X=5.59 $Y=1.485 $X2=5.59
+ $Y2=1.795
.ends

.subckt PM_SKY130_FD_SC_HS__AND4B_4%VPWR 1 2 3 4 5 6 7 26 30 32 36 40 44 48 51
+ 52 54 55 57 58 59 61 79 84 87 90 95 96
r94 95 96 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r95 93 95 10.5953 $w=5.93e-07 $l=5.15e-07 $layer=LI1_cond $X=7.34 $Y=2.815
+ $X2=7.34 $Y2=3.33
r96 90 91 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r97 88 91 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.64 $Y2=3.33
r98 87 88 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r99 84 85 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r100 82 96 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=7.44 $Y2=3.33
r101 81 82 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r102 79 95 8.24118 $w=1.7e-07 $l=3.4e-07 $layer=LI1_cond $X=7 $Y=3.33 $X2=7.34
+ $Y2=3.33
r103 79 81 2.60963 $w=1.68e-07 $l=4e-08 $layer=LI1_cond $X=7 $Y=3.33 $X2=6.96
+ $Y2=3.33
r104 78 82 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6 $Y=3.33 $X2=6.96
+ $Y2=3.33
r105 77 78 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r106 75 78 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.04 $Y=3.33 $X2=6
+ $Y2=3.33
r107 74 75 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r108 72 75 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=5.04 $Y2=3.33
r109 71 74 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=4.08 $Y=3.33
+ $X2=5.04 $Y2=3.33
r110 71 72 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r111 69 91 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=2.64 $Y2=3.33
r112 68 69 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r113 66 90 8.88104 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=2.98 $Y=3.33
+ $X2=2.807 $Y2=3.33
r114 66 68 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=2.98 $Y=3.33
+ $X2=3.6 $Y2=3.33
r115 65 88 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=1.68 $Y2=3.33
r116 65 85 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r117 64 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r118 62 84 9.39981 $w=1.7e-07 $l=1.88e-07 $layer=LI1_cond $X=1.025 $Y=3.33
+ $X2=0.837 $Y2=3.33
r119 62 64 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=1.025 $Y=3.33
+ $X2=1.2 $Y2=3.33
r120 61 87 9.14399 $w=1.7e-07 $l=1.8e-07 $layer=LI1_cond $X=1.595 $Y=3.33
+ $X2=1.775 $Y2=3.33
r121 61 64 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=1.595 $Y=3.33
+ $X2=1.2 $Y2=3.33
r122 59 72 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=3.84 $Y=3.33
+ $X2=4.08 $Y2=3.33
r123 59 69 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=3.84 $Y=3.33
+ $X2=3.6 $Y2=3.33
r124 57 77 6.52406 $w=1.68e-07 $l=1e-07 $layer=LI1_cond $X=6.1 $Y=3.33 $X2=6
+ $Y2=3.33
r125 57 58 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.1 $Y=3.33
+ $X2=6.265 $Y2=3.33
r126 56 81 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=6.43 $Y=3.33
+ $X2=6.96 $Y2=3.33
r127 56 58 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.43 $Y=3.33
+ $X2=6.265 $Y2=3.33
r128 54 74 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=5.18 $Y=3.33
+ $X2=5.04 $Y2=3.33
r129 54 55 8.9695 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=5.18 $Y=3.33
+ $X2=5.355 $Y2=3.33
r130 53 77 30.6631 $w=1.68e-07 $l=4.7e-07 $layer=LI1_cond $X=5.53 $Y=3.33 $X2=6
+ $Y2=3.33
r131 53 55 8.9695 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=5.53 $Y=3.33
+ $X2=5.355 $Y2=3.33
r132 51 68 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=3.72 $Y=3.33
+ $X2=3.6 $Y2=3.33
r133 51 52 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.72 $Y=3.33
+ $X2=3.885 $Y2=3.33
r134 50 71 1.95722 $w=1.68e-07 $l=3e-08 $layer=LI1_cond $X=4.05 $Y=3.33 $X2=4.08
+ $Y2=3.33
r135 50 52 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.05 $Y=3.33
+ $X2=3.885 $Y2=3.33
r136 46 58 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.265 $Y=3.245
+ $X2=6.265 $Y2=3.33
r137 46 48 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=6.265 $Y=3.245
+ $X2=6.265 $Y2=2.815
r138 42 55 1.07557 $w=3.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.355 $Y=3.245
+ $X2=5.355 $Y2=3.33
r139 42 44 14.1586 $w=3.48e-07 $l=4.3e-07 $layer=LI1_cond $X=5.355 $Y=3.245
+ $X2=5.355 $Y2=2.815
r140 38 52 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.885 $Y=3.245
+ $X2=3.885 $Y2=3.33
r141 38 40 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=3.885 $Y=3.245
+ $X2=3.885 $Y2=2.815
r142 34 90 1.03204 $w=3.45e-07 $l=8.5e-08 $layer=LI1_cond $X=2.807 $Y=3.245
+ $X2=2.807 $Y2=3.33
r143 34 36 14.3638 $w=3.43e-07 $l=4.3e-07 $layer=LI1_cond $X=2.807 $Y=3.245
+ $X2=2.807 $Y2=2.815
r144 33 87 9.14399 $w=1.7e-07 $l=1.8e-07 $layer=LI1_cond $X=1.955 $Y=3.33
+ $X2=1.775 $Y2=3.33
r145 32 90 8.88104 $w=1.7e-07 $l=1.72e-07 $layer=LI1_cond $X=2.635 $Y=3.33
+ $X2=2.807 $Y2=3.33
r146 32 33 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=2.635 $Y=3.33
+ $X2=1.955 $Y2=3.33
r147 28 87 1.16013 $w=3.6e-07 $l=8.5e-08 $layer=LI1_cond $X=1.775 $Y=3.245
+ $X2=1.775 $Y2=3.33
r148 28 30 13.7653 $w=3.58e-07 $l=4.3e-07 $layer=LI1_cond $X=1.775 $Y=3.245
+ $X2=1.775 $Y2=2.815
r149 24 84 1.28102 $w=3.75e-07 $l=8.5e-08 $layer=LI1_cond $X=0.837 $Y=3.245
+ $X2=0.837 $Y2=3.33
r150 24 26 13.2147 $w=3.73e-07 $l=4.3e-07 $layer=LI1_cond $X=0.837 $Y=3.245
+ $X2=0.837 $Y2=2.815
r151 7 93 600 $w=1.7e-07 $l=9.7857e-07 $layer=licon1_PDIFF $count=1 $X=7.015
+ $Y=1.96 $X2=7.28 $Y2=2.815
r152 6 48 600 $w=1.7e-07 $l=9.26971e-07 $layer=licon1_PDIFF $count=1 $X=6.115
+ $Y=1.96 $X2=6.265 $Y2=2.815
r153 5 44 600 $w=1.7e-07 $l=9.31571e-07 $layer=licon1_PDIFF $count=1 $X=5.195
+ $Y=1.96 $X2=5.355 $Y2=2.815
r154 4 40 600 $w=1.7e-07 $l=9.65376e-07 $layer=licon1_PDIFF $count=1 $X=3.65
+ $Y=1.96 $X2=3.885 $Y2=2.815
r155 3 36 600 $w=1.7e-07 $l=1.04964e-06 $layer=licon1_PDIFF $count=1 $X=2.65
+ $Y=1.84 $X2=2.805 $Y2=2.815
r156 2 30 600 $w=1.7e-07 $l=1.05428e-06 $layer=licon1_PDIFF $count=1 $X=1.61
+ $Y=1.84 $X2=1.775 $Y2=2.815
r157 1 26 600 $w=1.7e-07 $l=1.0951e-06 $layer=licon1_PDIFF $count=1 $X=0.58
+ $Y=1.84 $X2=0.835 $Y2=2.815
.ends

.subckt PM_SKY130_FD_SC_HS__AND4B_4%X 1 2 3 4 15 17 21 23 24 25 26 27 36 42 44
c61 17 0 1.18606e-19 $X=2.21 $Y=1.065
r62 34 42 1.64635 $w=3.83e-07 $l=5.5e-08 $layer=LI1_cond $X=1.277 $Y=0.98
+ $X2=1.277 $Y2=0.925
r63 27 44 4.75094 $w=2.3e-07 $l=2e-07 $layer=LI1_cond $X=1.2 $Y=2.02 $X2=1.2
+ $Y2=1.82
r64 26 44 7.76646 $w=2.28e-07 $l=1.55e-07 $layer=LI1_cond $X=1.2 $Y=1.665
+ $X2=1.2 $Y2=1.82
r65 25 26 18.5393 $w=2.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.2 $Y=1.295 $X2=1.2
+ $Y2=1.665
r66 25 43 7.2654 $w=2.28e-07 $l=1.45e-07 $layer=LI1_cond $X=1.2 $Y=1.295 $X2=1.2
+ $Y2=1.15
r67 24 34 3.0793 $w=3.07e-07 $l=8.5e-08 $layer=LI1_cond $X=1.277 $Y=1.065
+ $X2=1.277 $Y2=0.98
r68 24 43 3.0793 $w=3.07e-07 $l=1.17346e-07 $layer=LI1_cond $X=1.277 $Y=1.065
+ $X2=1.2 $Y2=1.15
r69 24 42 0.449004 $w=3.83e-07 $l=1.5e-08 $layer=LI1_cond $X=1.277 $Y=0.91
+ $X2=1.277 $Y2=0.925
r70 23 24 10.6264 $w=3.83e-07 $l=3.55e-07 $layer=LI1_cond $X=1.277 $Y=0.555
+ $X2=1.277 $Y2=0.91
r71 23 36 1.19734 $w=3.83e-07 $l=4e-08 $layer=LI1_cond $X=1.277 $Y=0.555
+ $X2=1.277 $Y2=0.515
r72 19 21 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=2.375 $Y=0.98
+ $X2=2.375 $Y2=0.515
r73 18 24 3.54158 $w=1.7e-07 $l=1.93e-07 $layer=LI1_cond $X=1.47 $Y=1.065
+ $X2=1.277 $Y2=1.065
r74 17 19 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.21 $Y=1.065
+ $X2=2.375 $Y2=0.98
r75 17 18 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=2.21 $Y=1.065
+ $X2=1.47 $Y2=1.065
r76 13 27 2.73179 $w=4e-07 $l=1.15e-07 $layer=LI1_cond $X=1.315 $Y=2.02 $X2=1.2
+ $Y2=2.02
r77 13 15 26.6502 $w=3.98e-07 $l=9.25e-07 $layer=LI1_cond $X=1.315 $Y=2.02
+ $X2=2.24 $Y2=2.02
r78 4 15 600 $w=1.7e-07 $l=2.43721e-07 $layer=licon1_PDIFF $count=1 $X=2.09
+ $Y=1.84 $X2=2.24 $Y2=2.02
r79 3 27 600 $w=1.7e-07 $l=2.43721e-07 $layer=licon1_PDIFF $count=1 $X=1.16
+ $Y=1.84 $X2=1.31 $Y2=2.02
r80 2 21 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.235
+ $Y=0.37 $X2=2.375 $Y2=0.515
r81 1 36 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.165
+ $Y=0.37 $X2=1.305 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__AND4B_4%VGND 1 2 3 4 15 17 21 25 29 32 33 34 36 45
+ 54 55 58 61 64
r83 64 65 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=4.56 $Y=0
+ $X2=4.56 $Y2=0
r84 61 62 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r85 59 62 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r86 58 59 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r87 55 65 0.802756 $w=4.9e-07 $l=2.88e-06 $layer=MET1_cond $X=7.44 $Y=0 $X2=4.56
+ $Y2=0
r88 54 55 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=7.44 $Y=0
+ $X2=7.44 $Y2=0
r89 52 64 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.615 $Y=0 $X2=4.45
+ $Y2=0
r90 52 54 184.305 $w=1.68e-07 $l=2.825e-06 $layer=LI1_cond $X=4.615 $Y=0
+ $X2=7.44 $Y2=0
r91 51 65 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=4.56
+ $Y2=0
r92 50 51 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r93 47 50 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=3.12 $Y=0 $X2=4.08
+ $Y2=0
r94 47 48 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r95 45 64 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.285 $Y=0 $X2=4.45
+ $Y2=0
r96 45 50 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=4.285 $Y=0 $X2=4.08
+ $Y2=0
r97 44 48 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r98 44 62 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=1.68
+ $Y2=0
r99 43 44 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r100 41 61 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2 $Y=0 $X2=1.835
+ $Y2=0
r101 41 43 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=2 $Y=0 $X2=2.64
+ $Y2=0
r102 39 59 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r103 38 39 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r104 36 58 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.585 $Y=0 $X2=0.75
+ $Y2=0
r105 36 38 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.585 $Y=0 $X2=0.24
+ $Y2=0
r106 34 51 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=3.84 $Y=0
+ $X2=4.08 $Y2=0
r107 34 48 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=3.84 $Y=0 $X2=3.12
+ $Y2=0
r108 32 43 4.56684 $w=1.68e-07 $l=7e-08 $layer=LI1_cond $X=2.71 $Y=0 $X2=2.64
+ $Y2=0
r109 32 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.71 $Y=0 $X2=2.875
+ $Y2=0
r110 31 47 5.21925 $w=1.68e-07 $l=8e-08 $layer=LI1_cond $X=3.04 $Y=0 $X2=3.12
+ $Y2=0
r111 31 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.04 $Y=0 $X2=2.875
+ $Y2=0
r112 27 64 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.45 $Y=0.085
+ $X2=4.45 $Y2=0
r113 27 29 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=4.45 $Y=0.085
+ $X2=4.45 $Y2=0.535
r114 23 33 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.875 $Y=0.085
+ $X2=2.875 $Y2=0
r115 23 25 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=2.875 $Y=0.085
+ $X2=2.875 $Y2=0.515
r116 19 61 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.835 $Y=0.085
+ $X2=1.835 $Y2=0
r117 19 21 19.5566 $w=3.28e-07 $l=5.6e-07 $layer=LI1_cond $X=1.835 $Y=0.085
+ $X2=1.835 $Y2=0.645
r118 18 58 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.915 $Y=0 $X2=0.75
+ $Y2=0
r119 17 61 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.67 $Y=0 $X2=1.835
+ $Y2=0
r120 17 18 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=1.67 $Y=0
+ $X2=0.915 $Y2=0
r121 13 58 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.75 $Y=0.085
+ $X2=0.75 $Y2=0
r122 13 15 17.8105 $w=3.28e-07 $l=5.1e-07 $layer=LI1_cond $X=0.75 $Y=0.085
+ $X2=0.75 $Y2=0.595
r123 4 29 182 $w=1.7e-07 $l=2.61151e-07 $layer=licon1_NDIFF $count=1 $X=4.23
+ $Y=0.625 $X2=4.45 $Y2=0.535
r124 3 25 91 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=2 $X=2.665
+ $Y=0.37 $X2=2.875 $Y2=0.515
r125 2 21 182 $w=1.7e-07 $l=3.76331e-07 $layer=licon1_NDIFF $count=1 $X=1.595
+ $Y=0.37 $X2=1.835 $Y2=0.645
r126 1 15 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=0.61
+ $Y=0.47 $X2=0.75 $Y2=0.595
.ends

.subckt PM_SKY130_FD_SC_HS__AND4B_4%A_664_125# 1 2 3 12 14 15 19 20 21 24
c59 14 0 1.17001e-19 $X=5.305 $Y=1.215
r60 22 24 12.3975 $w=3.28e-07 $l=3.55e-07 $layer=LI1_cond $X=7.33 $Y=0.425
+ $X2=7.33 $Y2=0.78
r61 20 22 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=7.165 $Y=0.34
+ $X2=7.33 $Y2=0.425
r62 20 21 110.257 $w=1.68e-07 $l=1.69e-06 $layer=LI1_cond $X=7.165 $Y=0.34
+ $X2=5.475 $Y2=0.34
r63 17 19 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=5.39 $Y=1.13
+ $X2=5.39 $Y2=0.77
r64 16 21 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.39 $Y=0.425
+ $X2=5.475 $Y2=0.34
r65 16 19 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=5.39 $Y=0.425
+ $X2=5.39 $Y2=0.77
r66 14 17 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.305 $Y=1.215
+ $X2=5.39 $Y2=1.13
r67 14 15 109.278 $w=1.68e-07 $l=1.675e-06 $layer=LI1_cond $X=5.305 $Y=1.215
+ $X2=3.63 $Y2=1.215
r68 10 15 22.9197 $w=8.4e-08 $l=2.03101e-07 $layer=LI1_cond $X=3.465 $Y=1.13
+ $X2=3.63 $Y2=1.215
r69 10 12 8.3814 $w=3.28e-07 $l=2.4e-07 $layer=LI1_cond $X=3.465 $Y=1.13
+ $X2=3.465 $Y2=0.89
r70 3 24 182 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_NDIFF $count=1 $X=7.19
+ $Y=0.625 $X2=7.33 $Y2=0.78
r71 2 19 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=5.25
+ $Y=0.625 $X2=5.39 $Y2=0.77
r72 1 12 182 $w=1.7e-07 $l=3.29621e-07 $layer=licon1_NDIFF $count=1 $X=3.32
+ $Y=0.625 $X2=3.465 $Y2=0.89
.ends

.subckt PM_SKY130_FD_SC_HS__AND4B_4%A_751_125# 1 2 7 12 14
r24 14 16 3.31764 $w=3.28e-07 $l=9.5e-08 $layer=LI1_cond $X=4.96 $Y=0.78
+ $X2=4.96 $Y2=0.875
r25 10 12 9.33524 $w=3.28e-07 $l=1.9e-07 $layer=LI1_cond $X=3.915 $Y=0.795
+ $X2=4.105 $Y2=0.795
r26 7 16 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.795 $Y=0.875
+ $X2=4.96 $Y2=0.875
r27 7 12 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=4.795 $Y=0.875
+ $X2=4.105 $Y2=0.875
r28 2 14 182 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_NDIFF $count=1 $X=4.82
+ $Y=0.625 $X2=4.96 $Y2=0.78
r29 1 10 182 $w=1.7e-07 $l=2.36854e-07 $layer=licon1_NDIFF $count=1 $X=3.755
+ $Y=0.625 $X2=3.915 $Y2=0.795
.ends

.subckt PM_SKY130_FD_SC_HS__AND4B_4%A_1136_125# 1 2 7 9 14
c20 9 0 5.7483e-20 $X=5.78 $Y=0.68
c21 7 0 2.3468e-20 $X=6.625 $Y=0.68
r22 14 17 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=6.79 $Y=0.68 $X2=6.79
+ $Y2=0.77
r23 9 12 4.60977 $w=2.48e-07 $l=1e-07 $layer=LI1_cond $X=5.78 $Y=0.68 $X2=5.78
+ $Y2=0.78
r24 8 9 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.905 $Y=0.68 $X2=5.78
+ $Y2=0.68
r25 7 14 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.625 $Y=0.68
+ $X2=6.79 $Y2=0.68
r26 7 8 46.9733 $w=1.68e-07 $l=7.2e-07 $layer=LI1_cond $X=6.625 $Y=0.68
+ $X2=5.905 $Y2=0.68
r27 2 17 182 $w=1.7e-07 $l=3.14245e-07 $layer=licon1_NDIFF $count=1 $X=6.54
+ $Y=0.625 $X2=6.79 $Y2=0.77
r28 1 12 182 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_NDIFF $count=1 $X=5.68
+ $Y=0.625 $X2=5.82 $Y2=0.78
.ends

