* File: sky130_fd_sc_hs__fah_4.spice
* Created: Thu Aug 27 20:46:28 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hs__fah_4.pex.spice"
.subckt sky130_fd_sc_hs__fah_4  VNB VPB A B CI VPWR COUT SUM VGND
* 
* VGND	VGND
* SUM	SUM
* COUT	COUT
* VPWR	VPWR
* CI	CI
* B	B
* A	A
* VPB	VPB
* VNB	VNB
MM1038 N_VGND_M1038_d N_A_M1038_g N_A_27_74#_M1038_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.0896 AS=0.1824 PD=0.92 PS=1.85 NRD=0 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75000.6 A=0.096 P=1.58 MULT=1
MM1039 N_A_200_74#_M1039_d N_A_M1039_g N_VGND_M1038_d VNB NLOWVT L=0.15 W=0.64
+ AD=0.1824 AS=0.0896 PD=1.85 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667 SA=75000.6
+ SB=75000.2 A=0.096 P=1.58 MULT=1
MM1004 N_A_427_362#_M1004_d N_A_27_74#_M1004_g N_VGND_M1004_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.124942 AS=0.418 PD=1.14217 PS=2.8 NRD=7.296 NRS=34.86 M=1
+ R=4.93333 SA=75000.4 SB=75001.7 A=0.111 P=1.78 MULT=1
MM1020 N_A_536_114#_M1020_d N_B_M1020_g N_A_427_362#_M1004_d VNB NLOWVT L=0.15
+ W=0.64 AD=0.0896 AS=0.108058 PD=0.92 PS=0.987826 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.9 SB=75001.5 A=0.096 P=1.58 MULT=1
MM1033 N_A_200_74#_M1033_d N_A_586_257#_M1033_g N_A_536_114#_M1020_d VNB NLOWVT
+ L=0.15 W=0.64 AD=0.1222 AS=0.0896 PD=1.08 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75001.3 SB=75001 A=0.096 P=1.58 MULT=1
MM1030 N_A_528_362#_M1030_d N_B_M1030_g N_A_200_74#_M1033_d VNB NLOWVT L=0.15
+ W=0.64 AD=0.1024 AS=0.1222 PD=0.96 PS=1.08 NRD=7.488 NRS=14.988 M=1 R=4.26667
+ SA=75001.6 SB=75000.7 A=0.096 P=1.58 MULT=1
MM1036 N_A_427_362#_M1036_d N_A_586_257#_M1036_g N_A_528_362#_M1030_d VNB NLOWVT
+ L=0.15 W=0.64 AD=0.1696 AS=0.1024 PD=1.81 PS=0.96 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75002.1 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1028 N_A_586_257#_M1028_d N_B_M1028_g N_VGND_M1028_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.2035 AS=0.27675 PD=2.05 PS=2.42 NRD=0 NRS=10.536 M=1 R=4.93333 SA=75000.2
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1025 N_A_1278_102#_M1025_d N_A_528_362#_M1025_g N_A_1183_102#_M1025_s VNB
+ NLOWVT L=0.15 W=0.64 AD=0.122062 AS=0.208 PD=1.105 PS=1.93 NRD=1.872 NRS=9.372
+ M=1 R=4.26667 SA=75000.2 SB=75001.3 A=0.096 P=1.58 MULT=1
MM1040 N_A_1378_125#_M1040_d N_A_536_114#_M1040_g N_A_1278_102#_M1025_d VNB
+ NLOWVT L=0.15 W=0.64 AD=0.0896 AS=0.122062 PD=0.92 PS=1.105 NRD=0 NRS=12.18
+ M=1 R=4.26667 SA=75000.6 SB=75001.1 A=0.096 P=1.58 MULT=1
MM1041 N_A_1265_379#_M1041_d N_A_528_362#_M1041_g N_A_1378_125#_M1040_d VNB
+ NLOWVT L=0.15 W=0.64 AD=0.118425 AS=0.0896 PD=1.09 PS=0.92 NRD=11.244 NRS=0
+ M=1 R=4.26667 SA=75001.1 SB=75000.7 A=0.096 P=1.58 MULT=1
MM1029 N_A_586_257#_M1029_d N_A_536_114#_M1029_g N_A_1265_379#_M1041_d VNB
+ NLOWVT L=0.15 W=0.64 AD=0.356425 AS=0.118425 PD=3.14 PS=1.09 NRD=94.104 NRS=0
+ M=1 R=4.26667 SA=75001.3 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1023 N_VGND_M1023_d N_A_1378_125#_M1023_g N_A_1183_102#_M1023_s VNB NLOWVT
+ L=0.15 W=0.64 AD=0.307107 AS=0.23505 PD=1.76232 PS=2.02 NRD=79.656 NRS=14.988
+ M=1 R=4.26667 SA=75000.3 SB=75002.7 A=0.096 P=1.58 MULT=1
MM1007 N_COUT_M1007_d N_A_1265_379#_M1007_g N_VGND_M1023_d VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.355093 PD=1.02 PS=2.03768 NRD=0 NRS=68.892 M=1 R=4.93333
+ SA=75001.2 SB=75001.7 A=0.111 P=1.78 MULT=1
MM1009 N_COUT_M1007_d N_A_1265_379#_M1009_g N_VGND_M1009_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.18675 PD=1.02 PS=1.45 NRD=0 NRS=32.004 M=1 R=4.93333
+ SA=75001.6 SB=75001.3 A=0.111 P=1.78 MULT=1
MM1015 N_COUT_M1015_d N_A_1265_379#_M1015_g N_VGND_M1009_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.18675 PD=1.02 PS=1.45 NRD=0 NRS=32.004 M=1 R=4.93333
+ SA=75002.1 SB=75000.7 A=0.111 P=1.78 MULT=1
MM1026 N_COUT_M1015_d N_A_1265_379#_M1026_g N_VGND_M1026_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.36 PD=1.02 PS=2.83 NRD=0 NRS=69.96 M=1 R=4.93333
+ SA=75002.6 SB=75000.3 A=0.111 P=1.78 MULT=1
MM1018 N_VGND_M1018_d N_CI_M1018_g N_A_1378_125#_M1018_s VNB NLOWVT L=0.15
+ W=0.64 AD=0.194087 AS=0.1824 PD=1.3913 PS=1.85 NRD=46.548 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75002.2 A=0.096 P=1.58 MULT=1
MM1002 N_VGND_M1018_d N_A_1278_102#_M1002_g N_SUM_M1002_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.224413 AS=0.1036 PD=1.6087 PS=1.02 NRD=40.248 NRS=0 M=1 R=4.93333
+ SA=75000.7 SB=75001.6 A=0.111 P=1.78 MULT=1
MM1032 N_VGND_M1032_d N_A_1278_102#_M1032_g N_SUM_M1002_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75001.2 SB=75001.1 A=0.111 P=1.78 MULT=1
MM1034 N_VGND_M1032_d N_A_1278_102#_M1034_g N_SUM_M1034_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75001.6 SB=75000.7 A=0.111 P=1.78 MULT=1
MM1043 N_VGND_M1043_d N_A_1278_102#_M1043_g N_SUM_M1034_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.2627 AS=0.1036 PD=2.19 PS=1.02 NRD=11.34 NRS=0 M=1 R=4.93333
+ SA=75002 SB=75000.3 A=0.111 P=1.78 MULT=1
MM1011 N_VPWR_M1011_d N_A_M1011_g N_A_27_74#_M1011_s VPB PSHORT L=0.15 W=1
+ AD=0.15 AS=0.295 PD=1.3 PS=2.59 NRD=1.9503 NRS=1.9503 M=1 R=6.66667 SA=75000.2
+ SB=75000.7 A=0.15 P=2.3 MULT=1
MM1012 N_A_200_74#_M1012_d N_A_M1012_g N_VPWR_M1011_d VPB PSHORT L=0.15 W=1
+ AD=0.295 AS=0.15 PD=2.59 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=6.66667 SA=75000.7
+ SB=75000.2 A=0.15 P=2.3 MULT=1
MM1013 N_A_427_362#_M1013_d N_A_27_74#_M1013_g N_VPWR_M1013_s VPB PSHORT L=0.15
+ W=1.12 AD=0.2128 AS=0.5163 PD=1.68571 PS=3.55 NRD=11.426 NRS=71.3928 M=1
+ R=7.46667 SA=75000.3 SB=75001.7 A=0.168 P=2.54 MULT=1
MM1003 N_A_528_362#_M1003_d N_B_M1003_g N_A_427_362#_M1013_d VPB PSHORT L=0.15
+ W=0.84 AD=0.1281 AS=0.1596 PD=1.145 PS=1.26429 NRD=2.3443 NRS=2.3443 M=1 R=5.6
+ SA=75000.8 SB=75001.7 A=0.126 P=1.98 MULT=1
MM1037 N_A_200_74#_M1037_d N_A_586_257#_M1037_g N_A_528_362#_M1003_d VPB PSHORT
+ L=0.15 W=0.84 AD=0.23945 AS=0.1281 PD=1.6 PS=1.145 NRD=53.9386 NRS=3.5066 M=1
+ R=5.6 SA=75001.3 SB=75001.3 A=0.126 P=1.98 MULT=1
MM1042 N_A_536_114#_M1042_d N_B_M1042_g N_A_200_74#_M1037_d VPB PSHORT L=0.15
+ W=0.84 AD=0.126 AS=0.23945 PD=1.14 PS=1.6 NRD=2.3443 NRS=53.9386 M=1 R=5.6
+ SA=75001.9 SB=75000.7 A=0.126 P=1.98 MULT=1
MM1000 N_A_427_362#_M1000_d N_A_586_257#_M1000_g N_A_536_114#_M1042_d VPB PSHORT
+ L=0.15 W=0.84 AD=0.2478 AS=0.126 PD=2.27 PS=1.14 NRD=2.3443 NRS=2.3443 M=1
+ R=5.6 SA=75002.3 SB=75000.2 A=0.126 P=1.98 MULT=1
MM1017 N_A_586_257#_M1017_d N_B_M1017_g N_VPWR_M1017_s VPB PSHORT L=0.15 W=1.12
+ AD=0.231057 AS=0.3304 PD=1.72 PS=2.83 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75003.8 A=0.168 P=2.54 MULT=1
MM1010 N_A_1265_379#_M1010_d N_A_528_362#_M1010_g N_A_586_257#_M1017_d VPB
+ PSHORT L=0.15 W=0.84 AD=0.1869 AS=0.173293 PD=1.285 PS=1.29 NRD=36.3465
+ NRS=22.261 M=1 R=5.6 SA=75000.8 SB=75004.4 A=0.126 P=1.98 MULT=1
MM1014 N_A_1378_125#_M1014_d N_A_536_114#_M1014_g N_A_1265_379#_M1010_d VPB
+ PSHORT L=0.15 W=0.84 AD=0.22505 AS=0.1869 PD=1.55 PS=1.285 NRD=49.9198 NRS=0
+ M=1 R=5.6 SA=75001.3 SB=75003.8 A=0.126 P=1.98 MULT=1
MM1019 N_A_1278_102#_M1019_d N_A_528_362#_M1019_g N_A_1378_125#_M1014_d VPB
+ PSHORT L=0.15 W=0.84 AD=0.336 AS=0.22505 PD=1.64 PS=1.55 NRD=119.599
+ NRS=15.2281 M=1 R=5.6 SA=75001.6 SB=75004 A=0.126 P=1.98 MULT=1
MM1024 N_A_1183_102#_M1024_d N_A_536_114#_M1024_g N_A_1278_102#_M1019_d VPB
+ PSHORT L=0.15 W=0.84 AD=0.178374 AS=0.336 PD=1.36957 PS=1.64 NRD=36.8981
+ NRS=2.3443 M=1 R=5.6 SA=75002.5 SB=75003.1 A=0.126 P=1.98 MULT=1
MM1031 N_VPWR_M1031_d N_A_1378_125#_M1031_g N_A_1183_102#_M1024_d VPB PSHORT
+ L=0.15 W=1 AD=0.425 AS=0.212351 PD=1.93396 PS=1.63043 NRD=72.8703 NRS=1.9503
+ M=1 R=6.66667 SA=75002.4 SB=75003 A=0.15 P=2.3 MULT=1
MM1005 N_COUT_M1005_d N_A_1265_379#_M1005_g N_VPWR_M1031_d VPB PSHORT L=0.15
+ W=1.12 AD=0.168 AS=0.476 PD=1.42 PS=2.16604 NRD=0 NRS=65.0691 M=1 R=7.46667
+ SA=75003 SB=75002.1 A=0.168 P=2.54 MULT=1
MM1006 N_COUT_M1005_d N_A_1265_379#_M1006_g N_VPWR_M1006_s VPB PSHORT L=0.15
+ W=1.12 AD=0.168 AS=0.297275 PD=1.42 PS=1.825 NRD=1.7533 NRS=36.9966 M=1
+ R=7.46667 SA=75003.4 SB=75001.7 A=0.168 P=2.54 MULT=1
MM1008 N_COUT_M1008_d N_A_1265_379#_M1008_g N_VPWR_M1006_s VPB PSHORT L=0.15
+ W=1.12 AD=0.168 AS=0.297275 PD=1.42 PS=1.825 NRD=1.7533 NRS=36.9966 M=1
+ R=7.46667 SA=75004 SB=75001.1 A=0.168 P=2.54 MULT=1
MM1035 N_COUT_M1008_d N_A_1265_379#_M1035_g N_VPWR_M1035_s VPB PSHORT L=0.15
+ W=1.12 AD=0.168 AS=0.8914 PD=1.42 PS=4.04 NRD=0 NRS=130.315 M=1 R=7.46667
+ SA=75004.5 SB=75000.6 A=0.168 P=2.54 MULT=1
MM1016 N_VPWR_M1016_d N_CI_M1016_g N_A_1378_125#_M1016_s VPB PSHORT L=0.15 W=1
+ AD=0.224717 AS=0.295 PD=1.46698 PS=2.59 NRD=19.0302 NRS=1.9503 M=1 R=6.66667
+ SA=75000.2 SB=75002.3 A=0.15 P=2.3 MULT=1
MM1001 N_SUM_M1001_d N_A_1278_102#_M1001_g N_VPWR_M1016_d VPB PSHORT L=0.15
+ W=1.12 AD=0.168 AS=0.251683 PD=1.42 PS=1.64302 NRD=1.7533 NRS=10.5395 M=1
+ R=7.46667 SA=75000.7 SB=75001.7 A=0.168 P=2.54 MULT=1
MM1021 N_SUM_M1001_d N_A_1278_102#_M1021_g N_VPWR_M1021_s VPB PSHORT L=0.15
+ W=1.12 AD=0.168 AS=0.2184 PD=1.42 PS=1.51 NRD=1.7533 NRS=10.5395 M=1 R=7.46667
+ SA=75001.2 SB=75001.2 A=0.168 P=2.54 MULT=1
MM1022 N_SUM_M1022_d N_A_1278_102#_M1022_g N_VPWR_M1021_s VPB PSHORT L=0.15
+ W=1.12 AD=0.1736 AS=0.2184 PD=1.43 PS=1.51 NRD=3.5066 NRS=8.7862 M=1 R=7.46667
+ SA=75001.7 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1027 N_SUM_M1022_d N_A_1278_102#_M1027_g N_VPWR_M1027_s VPB PSHORT L=0.15
+ W=1.12 AD=0.1736 AS=0.3304 PD=1.43 PS=2.83 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75002.2 SB=75000.2 A=0.168 P=2.54 MULT=1
DX44_noxref VNB VPB NWDIODE A=29.3716 P=35.37
c_161 VNB 0 3.55461e-19 $X=0 $Y=0
*
.include "sky130_fd_sc_hs__fah_4.pxi.spice"
*
.ends
*
*
