* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hs__dlxtp_1 D GATE VGND VNB VPB VPWR Q
M1000 VGND a_116_424# a_239_85# VNB nlowvt w=740000u l=150000u
+  ad=1.47895e+12p pd=1.06e+07u as=4.458e+11p ps=4.22e+06u
M1001 VPWR GATE a_562_123# VPB pshort w=840000u l=150000u
+  ad=1.69967e+12p pd=1.266e+07u as=2.478e+11p ps=2.27e+06u
M1002 a_419_392# a_685_59# a_592_149# VPB pshort w=420000u l=150000u
+  ad=3.1685e+11p pd=3.26e+06u as=3.328e+11p ps=2.77e+06u
M1003 a_592_149# a_562_123# a_229_392# VPB pshort w=1e+06u l=150000u
+  ad=0p pd=0u as=5.9e+11p ps=5.18e+06u
M1004 Q a_386_326# VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=3.304e+11p pd=2.83e+06u as=0p ps=0u
M1005 a_685_59# a_562_123# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1006 a_592_149# a_562_123# a_514_149# VNB nlowvt w=420000u l=150000u
+  ad=2.753e+11p pd=2.41e+06u as=1.008e+11p ps=1.32e+06u
M1007 Q a_386_326# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1008 a_116_424# D VGND VNB nlowvt w=550000u l=150000u
+  ad=1.815e+11p pd=1.76e+06u as=0p ps=0u
M1009 a_419_392# a_386_326# VPWR VPB pshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VGND a_592_149# a_386_326# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1011 a_514_149# a_386_326# VGND VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VPWR a_116_424# a_229_392# VPB pshort w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_116_424# D VPWR VPB pshort w=840000u l=150000u
+  ad=2.478e+11p pd=2.27e+06u as=0p ps=0u
M1014 a_239_85# a_685_59# a_592_149# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VGND GATE a_562_123# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.22e+11p ps=2.08e+06u
M1016 VPWR a_592_149# a_386_326# VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=3.696e+11p ps=2.9e+06u
M1017 a_685_59# a_562_123# VPWR VPB pshort w=840000u l=150000u
+  ad=2.478e+11p pd=2.27e+06u as=0p ps=0u
.ends
