* File: sky130_fd_sc_hs__bufinv_8.spice
* Created: Thu Aug 27 20:35:14 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hs__bufinv_8.pex.spice"
.subckt sky130_fd_sc_hs__bufinv_8  VNB VPB A VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A	A
* VPB	VPB
* VNB	VNB
MM1023 N_VGND_M1023_d N_A_M1023_g N_A_27_368#_M1023_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1221 AS=0.2109 PD=1.07 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75005.4 A=0.111 P=1.78 MULT=1
MM1000 N_Y_M1000_d N_A_183_48#_M1000_g N_VGND_M1023_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.111 AS=0.1221 PD=1.04 PS=1.07 NRD=3.24 NRS=8.1 M=1 R=4.93333 SA=75000.7
+ SB=75005 A=0.111 P=1.78 MULT=1
MM1001 N_Y_M1000_d N_A_183_48#_M1001_g N_VGND_M1001_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.111 AS=0.1295 PD=1.04 PS=1.09 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75001.1
+ SB=75004.5 A=0.111 P=1.78 MULT=1
MM1004 N_Y_M1004_d N_A_183_48#_M1004_g N_VGND_M1001_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1295 PD=1.02 PS=1.09 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.6
+ SB=75004 A=0.111 P=1.78 MULT=1
MM1005 N_Y_M1004_d N_A_183_48#_M1005_g N_VGND_M1005_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1295 PD=1.02 PS=1.09 NRD=0 NRS=0 M=1 R=4.93333 SA=75002.1
+ SB=75003.6 A=0.111 P=1.78 MULT=1
MM1011 N_Y_M1011_d N_A_183_48#_M1011_g N_VGND_M1005_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1295 PD=1.02 PS=1.09 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75002.6
+ SB=75003.1 A=0.111 P=1.78 MULT=1
MM1015 N_Y_M1011_d N_A_183_48#_M1015_g N_VGND_M1015_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1295 PD=1.02 PS=1.09 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75003
+ SB=75002.7 A=0.111 P=1.78 MULT=1
MM1017 N_Y_M1017_d N_A_183_48#_M1017_g N_VGND_M1015_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1295 AS=0.1295 PD=1.09 PS=1.09 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75003.5
+ SB=75002.2 A=0.111 P=1.78 MULT=1
MM1020 N_Y_M1017_d N_A_183_48#_M1020_g N_VGND_M1020_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1295 AS=0.1295 PD=1.09 PS=1.09 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75004
+ SB=75001.7 A=0.111 P=1.78 MULT=1
MM1002 N_A_183_48#_M1002_d N_A_27_368#_M1002_g N_VGND_M1020_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.10915 AS=0.1295 PD=1.035 PS=1.09 NRD=0.804 NRS=0 M=1 R=4.93333
+ SA=75004.5 SB=75001.2 A=0.111 P=1.78 MULT=1
MM1006 N_A_183_48#_M1002_d N_A_27_368#_M1006_g N_VGND_M1006_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.10915 AS=0.1295 PD=1.035 PS=1.09 NRD=1.62 NRS=0 M=1 R=4.93333
+ SA=75004.9 SB=75000.7 A=0.111 P=1.78 MULT=1
MM1012 N_A_183_48#_M1012_d N_A_27_368#_M1012_g N_VGND_M1006_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.2109 AS=0.1295 PD=2.05 PS=1.09 NRD=0 NRS=11.34 M=1 R=4.93333
+ SA=75005.4 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1008 N_VPWR_M1008_d N_A_M1008_g N_A_27_368#_M1008_s VPB PSHORT L=0.15 W=1.12
+ AD=0.196 AS=0.3304 PD=1.47 PS=2.83 NRD=10.5395 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75005.4 A=0.168 P=2.54 MULT=1
MM1003 N_Y_M1003_d N_A_183_48#_M1003_g N_VPWR_M1008_d VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.196 PD=1.42 PS=1.47 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.7 SB=75004.9 A=0.168 P=2.54 MULT=1
MM1007 N_Y_M1003_d N_A_183_48#_M1007_g N_VPWR_M1007_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.2 SB=75004.5 A=0.168 P=2.54 MULT=1
MM1009 N_Y_M1009_d N_A_183_48#_M1009_g N_VPWR_M1007_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.6 SB=75004 A=0.168 P=2.54 MULT=1
MM1013 N_Y_M1009_d N_A_183_48#_M1013_g N_VPWR_M1013_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75002.1 SB=75003.6 A=0.168 P=2.54 MULT=1
MM1014 N_Y_M1014_d N_A_183_48#_M1014_g N_VPWR_M1013_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75002.5 SB=75003.1 A=0.168 P=2.54 MULT=1
MM1016 N_Y_M1014_d N_A_183_48#_M1016_g N_VPWR_M1016_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667 SA=75003
+ SB=75002.7 A=0.168 P=2.54 MULT=1
MM1018 N_Y_M1018_d N_A_183_48#_M1018_g N_VPWR_M1016_s VPB PSHORT L=0.15 W=1.12
+ AD=0.2408 AS=0.168 PD=1.55 PS=1.42 NRD=13.1793 NRS=1.7533 M=1 R=7.46667
+ SA=75003.4 SB=75002.2 A=0.168 P=2.54 MULT=1
MM1021 N_Y_M1018_d N_A_183_48#_M1021_g N_VPWR_M1021_s VPB PSHORT L=0.15 W=1.12
+ AD=0.2408 AS=0.196 PD=1.55 PS=1.47 NRD=13.1793 NRS=1.7533 M=1 R=7.46667
+ SA=75004 SB=75001.7 A=0.168 P=2.54 MULT=1
MM1010 N_A_183_48#_M1010_d N_A_27_368#_M1010_g N_VPWR_M1021_s VPB PSHORT L=0.15
+ W=1.12 AD=0.168 AS=0.196 PD=1.42 PS=1.47 NRD=1.7533 NRS=10.5395 M=1 R=7.46667
+ SA=75004.5 SB=75001.2 A=0.168 P=2.54 MULT=1
MM1019 N_A_183_48#_M1010_d N_A_27_368#_M1019_g N_VPWR_M1019_s VPB PSHORT L=0.15
+ W=1.12 AD=0.168 AS=0.196 PD=1.42 PS=1.47 NRD=1.7533 NRS=10.5395 M=1 R=7.46667
+ SA=75004.9 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1022 N_A_183_48#_M1022_d N_A_27_368#_M1022_g N_VPWR_M1019_s VPB PSHORT L=0.15
+ W=1.12 AD=0.3304 AS=0.196 PD=2.83 PS=1.47 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75005.4 SB=75000.2 A=0.168 P=2.54 MULT=1
DX24_noxref VNB VPB NWDIODE A=12.3132 P=16.96
*
.include "sky130_fd_sc_hs__bufinv_8.pxi.spice"
*
.ends
*
*
