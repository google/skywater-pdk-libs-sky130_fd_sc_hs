* File: sky130_fd_sc_hs__dlrtn_2.spice
* Created: Thu Aug 27 20:41:32 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hs__dlrtn_2.pex.spice"
.subckt sky130_fd_sc_hs__dlrtn_2  VNB VPB D GATE_N RESET_B VPWR Q VGND
* 
* VGND	VGND
* Q	Q
* VPWR	VPWR
* RESET_B	RESET_B
* GATE_N	GATE_N
* D	D
* VPB	VPB
* VNB	VNB
MM1018 N_VGND_M1018_d N_D_M1018_g N_A_27_136#_M1018_s VNB NLOWVT L=0.15 W=0.55
+ AD=0.171076 AS=0.15675 PD=1.27054 PS=1.67 NRD=55.86 NRS=0 M=1 R=3.66667
+ SA=75000.2 SB=75000.8 A=0.0825 P=1.4 MULT=1
MM1002 N_A_232_98#_M1002_d N_GATE_N_M1002_g N_VGND_M1018_d VNB NLOWVT L=0.15
+ W=0.74 AD=0.2257 AS=0.230174 PD=2.09 PS=1.70946 NRD=0 NRS=41.52 M=1 R=4.93333
+ SA=75000.7 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1007 N_VGND_M1007_d N_A_232_98#_M1007_g N_A_373_82#_M1007_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.4514 AS=0.2294 PD=2.12348 PS=2.1 NRD=89.988 NRS=2.424 M=1
+ R=4.93333 SA=75000.2 SB=75001.9 A=0.111 P=1.78 MULT=1
MM1015 A_697_74# N_A_27_136#_M1015_g N_VGND_M1007_d VNB NLOWVT L=0.15 W=0.64
+ AD=0.0768 AS=0.3904 PD=0.88 PS=1.83652 NRD=12.18 NRS=15.936 M=1 R=4.26667
+ SA=75001.4 SB=75001.2 A=0.096 P=1.58 MULT=1
MM1012 N_A_670_392#_M1012_d N_A_232_98#_M1012_g A_697_74# VNB NLOWVT L=0.15
+ W=0.64 AD=0.115623 AS=0.0768 PD=1.16528 PS=0.88 NRD=8.436 NRS=12.18 M=1
+ R=4.26667 SA=75001.8 SB=75000.8 A=0.096 P=1.58 MULT=1
MM1021 A_870_74# N_A_373_82#_M1021_g N_A_670_392#_M1012_d VNB NLOWVT L=0.15
+ W=0.42 AD=0.05775 AS=0.0758774 PD=0.695 PS=0.764717 NRD=23.568 NRS=0 M=1 R=2.8
+ SA=75002.2 SB=75000.6 A=0.063 P=1.14 MULT=1
MM1019 N_VGND_M1019_d N_A_913_406#_M1019_g A_870_74# VNB NLOWVT L=0.15 W=0.42
+ AD=0.1197 AS=0.05775 PD=1.41 PS=0.695 NRD=0 NRS=23.568 M=1 R=2.8 SA=75002.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1003 A_1153_74# N_A_670_392#_M1003_g N_A_913_406#_M1003_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.0888 AS=0.2109 PD=0.98 PS=2.05 NRD=10.536 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75002.2 A=0.111 P=1.78 MULT=1
MM1001 N_VGND_M1001_d N_RESET_B_M1001_g A_1153_74# VNB NLOWVT L=0.15 W=0.74
+ AD=0.34225 AS=0.0888 PD=1.665 PS=0.98 NRD=0 NRS=10.536 M=1 R=4.93333
+ SA=75000.6 SB=75001.8 A=0.111 P=1.78 MULT=1
MM1006 N_Q_M1006_d N_A_913_406#_M1006_g N_VGND_M1001_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.34225 PD=1.02 PS=1.665 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75001.7
+ SB=75000.7 A=0.111 P=1.78 MULT=1
MM1011 N_Q_M1006_d N_A_913_406#_M1011_g N_VGND_M1011_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.2627 PD=1.02 PS=2.19 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75002.1
+ SB=75000.3 A=0.111 P=1.78 MULT=1
MM1004 N_VPWR_M1004_d N_D_M1004_g N_A_27_136#_M1004_s VPB PSHORT L=0.15 W=0.84
+ AD=0.168 AS=0.2478 PD=1.24 PS=2.27 NRD=14.0658 NRS=2.3443 M=1 R=5.6 SA=75000.2
+ SB=75000.8 A=0.126 P=1.98 MULT=1
MM1000 N_A_232_98#_M1000_d N_GATE_N_M1000_g N_VPWR_M1004_d VPB PSHORT L=0.15
+ W=0.84 AD=0.2478 AS=0.168 PD=2.27 PS=1.24 NRD=2.3443 NRS=14.0658 M=1 R=5.6
+ SA=75000.8 SB=75000.2 A=0.126 P=1.98 MULT=1
MM1016 N_VPWR_M1016_d N_A_232_98#_M1016_g N_A_373_82#_M1016_s VPB PSHORT L=0.15
+ W=0.84 AD=0.235793 AS=0.2478 PD=1.53391 PS=2.27 NRD=52.9142 NRS=2.3443 M=1
+ R=5.6 SA=75000.2 SB=75002.7 A=0.126 P=1.98 MULT=1
MM1008 A_586_392# N_A_27_136#_M1008_g N_VPWR_M1016_d VPB PSHORT L=0.15 W=1
+ AD=0.135 AS=0.280707 PD=1.27 PS=1.82609 NRD=15.7403 NRS=19.6803 M=1 R=6.66667
+ SA=75000.8 SB=75002.5 A=0.15 P=2.3 MULT=1
MM1020 N_A_670_392#_M1020_d N_A_373_82#_M1020_g A_586_392# VPB PSHORT L=0.15 W=1
+ AD=0.237394 AS=0.135 PD=1.95775 PS=1.27 NRD=1.9503 NRS=15.7403 M=1 R=6.66667
+ SA=75001.2 SB=75002.1 A=0.15 P=2.3 MULT=1
MM1017 A_778_504# N_A_232_98#_M1017_g N_A_670_392#_M1020_d VPB PSHORT L=0.15
+ W=0.42 AD=0.1449 AS=0.0997056 PD=1.11 PS=0.822254 NRD=136.009 NRS=85.5374 M=1
+ R=2.8 SA=75001.6 SB=75004.1 A=0.063 P=1.14 MULT=1
MM1009 N_VPWR_M1009_d N_A_913_406#_M1009_g A_778_504# VPB PSHORT L=0.15 W=0.42
+ AD=0.146809 AS=0.1449 PD=1.06909 PS=1.11 NRD=4.6886 NRS=136.009 M=1 R=2.8
+ SA=75002.5 SB=75003.2 A=0.063 P=1.14 MULT=1
MM1013 N_A_913_406#_M1013_d N_A_670_392#_M1013_g N_VPWR_M1009_d VPB PSHORT
+ L=0.15 W=1.12 AD=0.1736 AS=0.391491 PD=1.43 PS=2.85091 NRD=3.5066 NRS=8.7862
+ M=1 R=7.46667 SA=75001.4 SB=75002.2 A=0.168 P=2.54 MULT=1
MM1005 N_VPWR_M1005_d N_RESET_B_M1005_g N_A_913_406#_M1013_d VPB PSHORT L=0.15
+ W=1.12 AD=0.4984 AS=0.1736 PD=2.01 PS=1.43 NRD=29.0181 NRS=1.7533 M=1
+ R=7.46667 SA=75001.9 SB=75001.8 A=0.168 P=2.54 MULT=1
MM1010 N_Q_M1010_d N_A_913_406#_M1010_g N_VPWR_M1005_d VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.4984 PD=1.42 PS=2.01 NRD=1.7533 NRS=78.2681 M=1 R=7.46667
+ SA=75002.9 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1014 N_Q_M1010_d N_A_913_406#_M1014_g N_VPWR_M1014_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.3976 PD=1.42 PS=2.95 NRD=1.7533 NRS=11.426 M=1 R=7.46667
+ SA=75003.4 SB=75000.3 A=0.168 P=2.54 MULT=1
DX22_noxref VNB VPB NWDIODE A=15.8844 P=20.8
*
.include "sky130_fd_sc_hs__dlrtn_2.pxi.spice"
*
.ends
*
*
