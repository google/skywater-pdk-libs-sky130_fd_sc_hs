* File: sky130_fd_sc_hs__a211o_2.spice
* Created: Tue Sep  1 19:48:30 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hs__a211o_2.pex.spice"
.subckt sky130_fd_sc_hs__a211o_2  VNB VPB A2 A1 B1 C1 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* C1	C1
* B1	B1
* A1	A1
* A2	A2
* VPB	VPB
* VNB	VNB
MM1005 N_VGND_M1005_d N_A_85_270#_M1005_g N_X_M1005_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1961 AS=0.1036 PD=2.01 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75002.9 A=0.111 P=1.78 MULT=1
MM1009 N_VGND_M1009_d N_A_85_270#_M1009_g N_X_M1005_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.2442 AS=0.1036 PD=1.4 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.6
+ SB=75002.4 A=0.111 P=1.78 MULT=1
MM1003 A_399_74# N_A2_M1003_g N_VGND_M1009_d VNB NLOWVT L=0.15 W=0.74 AD=0.0777
+ AS=0.2442 PD=0.95 PS=1.4 NRD=8.1 NRS=0 M=1 R=4.93333 SA=75001.4 SB=75001.6
+ A=0.111 P=1.78 MULT=1
MM1000 N_A_85_270#_M1000_d N_A1_M1000_g A_399_74# VNB NLOWVT L=0.15 W=0.74
+ AD=0.1443 AS=0.0777 PD=1.13 PS=0.95 NRD=3.24 NRS=8.1 M=1 R=4.93333 SA=75001.8
+ SB=75001.3 A=0.111 P=1.78 MULT=1
MM1006 N_VGND_M1006_d N_B1_M1006_g N_A_85_270#_M1000_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.1443 AS=0.1443 PD=1.13 PS=1.13 NRD=8.916 NRS=14.592 M=1 R=4.93333
+ SA=75002.3 SB=75000.7 A=0.111 P=1.78 MULT=1
MM1010 N_A_85_270#_M1010_d N_C1_M1010_g N_VGND_M1006_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.1961 AS=0.1443 PD=2.01 PS=1.13 NRD=0 NRS=8.916 M=1 R=4.93333 SA=75002.9
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1001 N_X_M1001_d N_A_85_270#_M1001_g N_VPWR_M1001_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.308 PD=1.42 PS=2.79 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75000.6 A=0.168 P=2.54 MULT=1
MM1002 N_X_M1001_d N_A_85_270#_M1002_g N_VPWR_M1002_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.308 PD=1.42 PS=2.79 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.6 SB=75000.2 A=0.168 P=2.54 MULT=1
MM1004 N_VPWR_M1004_d N_A2_M1004_g N_A_317_392#_M1004_s VPB PSHORT L=0.15 W=1
+ AD=0.195 AS=0.275 PD=1.39 PS=2.55 NRD=5.8903 NRS=1.9503 M=1 R=6.66667
+ SA=75000.2 SB=75001.6 A=0.15 P=2.3 MULT=1
MM1007 N_A_317_392#_M1007_d N_A1_M1007_g N_VPWR_M1004_d VPB PSHORT L=0.15 W=1
+ AD=0.15 AS=0.195 PD=1.3 PS=1.39 NRD=1.9503 NRS=15.7403 M=1 R=6.66667
+ SA=75000.7 SB=75001.1 A=0.15 P=2.3 MULT=1
MM1008 A_600_392# N_B1_M1008_g N_A_317_392#_M1007_d VPB PSHORT L=0.15 W=1
+ AD=0.135 AS=0.15 PD=1.27 PS=1.3 NRD=15.7403 NRS=1.9503 M=1 R=6.66667
+ SA=75001.2 SB=75000.6 A=0.15 P=2.3 MULT=1
MM1011 N_A_85_270#_M1011_d N_C1_M1011_g A_600_392# VPB PSHORT L=0.15 W=1
+ AD=0.275 AS=0.135 PD=2.55 PS=1.27 NRD=1.9503 NRS=15.7403 M=1 R=6.66667
+ SA=75001.6 SB=75000.2 A=0.15 P=2.3 MULT=1
DX12_noxref VNB VPB NWDIODE A=7.8492 P=12.16
*
.include "sky130_fd_sc_hs__a211o_2.pxi.spice"
*
.ends
*
*
