* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hs__edfxtp_1 CLK D DE VGND VNB VPB VPWR Q
M1000 a_1156_90# a_958_74# a_27_508# VPB pshort w=420000u l=150000u
+  ad=1.26e+11p pd=1.44e+06u as=3.528e+11p ps=4.2e+06u
M1001 VGND a_1409_64# a_1349_90# VNB nlowvt w=420000u l=150000u
+  ad=1.8056e+12p pd=1.622e+07u as=1.26e+11p ps=1.44e+06u
M1002 a_763_74# CLK VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=3.08e+11p pd=2.79e+06u as=2.22792e+12p ps=1.982e+07u
M1003 VPWR a_159_446# a_114_508# VPB pshort w=420000u l=150000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1004 a_1382_508# a_763_74# a_1156_90# VPB pshort w=420000u l=150000u
+  ad=1.491e+11p pd=1.55e+06u as=0p ps=0u
M1005 VGND a_533_61# a_1997_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1006 a_2088_502# a_958_74# a_1895_74# VPB pshort w=420000u l=150000u
+  ad=1.134e+11p pd=1.38e+06u as=3.328e+11p ps=2.77e+06u
M1007 a_533_61# a_1895_74# VGND VNB nlowvt w=420000u l=150000u
+  ad=1.197e+11p pd=1.41e+06u as=0p ps=0u
M1008 a_1409_64# a_1156_90# VGND VNB nlowvt w=640000u l=150000u
+  ad=1.824e+11p pd=1.85e+06u as=0p ps=0u
M1009 VGND DE a_131_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1010 VPWR a_1895_74# Q VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=3.08e+11p ps=2.79e+06u
M1011 a_1997_74# a_763_74# a_1895_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=2.424e+11p ps=2.2e+06u
M1012 VPWR DE a_159_446# VPB pshort w=640000u l=150000u
+  ad=0p pd=0u as=1.888e+11p ps=1.87e+06u
M1013 a_131_74# D a_27_508# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=3.591e+11p ps=4.23e+06u
M1014 VGND DE a_159_446# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.176e+11p ps=1.4e+06u
M1015 a_1409_64# a_1156_90# VPWR VPB pshort w=840000u l=150000u
+  ad=2.478e+11p pd=2.27e+06u as=0p ps=0u
M1016 a_27_508# a_533_61# a_554_436# VPB pshort w=420000u l=150000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1017 a_763_74# CLK VGND VNB nlowvt w=740000u l=150000u
+  ad=2.035e+11p pd=2.03e+06u as=0p ps=0u
M1018 a_1797_74# a_1409_64# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.516e+11p pd=2.16e+06u as=0p ps=0u
M1019 a_958_74# a_763_74# VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=3.08e+11p pd=2.79e+06u as=0p ps=0u
M1020 a_114_508# D a_27_508# VPB pshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_1895_74# a_763_74# a_1794_392# VPB pshort w=1e+06u l=150000u
+  ad=0p pd=0u as=7.85e+11p ps=3.57e+06u
M1022 VGND a_1895_74# Q VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1023 a_491_87# a_159_446# VGND VNB nlowvt w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1024 VPWR a_533_61# a_2088_502# VPB pshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 a_27_508# a_533_61# a_491_87# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 a_554_436# DE VPWR VPB pshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 a_533_61# a_1895_74# VPWR VPB pshort w=640000u l=150000u
+  ad=1.76e+11p pd=1.83e+06u as=0p ps=0u
M1028 a_1156_90# a_763_74# a_27_508# VNB nlowvt w=420000u l=150000u
+  ad=3.423e+11p pd=2.47e+06u as=0p ps=0u
M1029 a_1794_392# a_1409_64# VPWR VPB pshort w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1030 VPWR a_1409_64# a_1382_508# VPB pshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1031 a_1349_90# a_958_74# a_1156_90# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1032 a_1895_74# a_958_74# a_1797_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1033 a_958_74# a_763_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
.ends
