* File: sky130_fd_sc_hs__nor3_4.pxi.spice
* Created: Tue Sep  1 20:11:38 2020
* 
x_PM_SKY130_FD_SC_HS__NOR3_4%A N_A_M1004_g N_A_c_115_n N_A_M1005_g N_A_M1016_g
+ N_A_c_116_n N_A_M1006_g N_A_c_117_n N_A_M1012_g N_A_c_118_n N_A_M1013_g
+ N_A_c_169_p N_A_c_110_n N_A_c_145_p N_A_c_130_p N_A_c_111_n N_A_c_112_n
+ N_A_c_113_n N_A_c_131_p A A A N_A_c_114_n N_A_c_128_p
+ PM_SKY130_FD_SC_HS__NOR3_4%A
x_PM_SKY130_FD_SC_HS__NOR3_4%B N_B_c_246_n N_B_c_247_n N_B_M1003_g N_B_c_248_n
+ N_B_M1007_g N_B_c_249_n N_B_c_250_n N_B_M1011_g N_B_c_251_n N_B_c_263_n
+ N_B_M1014_g N_B_c_252_n N_B_c_265_n N_B_M1015_g N_B_c_253_n N_B_c_267_n
+ N_B_M1017_g N_B_c_254_n N_B_c_255_n N_B_c_268_n B B N_B_c_256_n N_B_c_257_n
+ N_B_c_258_n N_B_c_259_n B B N_B_c_260_n PM_SKY130_FD_SC_HS__NOR3_4%B
x_PM_SKY130_FD_SC_HS__NOR3_4%C N_C_c_385_n N_C_M1000_g N_C_c_372_n N_C_c_373_n
+ N_C_M1001_g N_C_c_388_n N_C_M1002_g N_C_c_375_n N_C_c_376_n N_C_M1010_g
+ N_C_c_391_n N_C_M1008_g N_C_c_378_n N_C_c_379_n N_C_c_394_n N_C_M1009_g
+ N_C_c_380_n N_C_c_381_n N_C_c_382_n C C C C N_C_c_384_n
+ PM_SKY130_FD_SC_HS__NOR3_4%C
x_PM_SKY130_FD_SC_HS__NOR3_4%A_27_368# N_A_27_368#_M1005_s N_A_27_368#_M1006_s
+ N_A_27_368#_M1014_d N_A_27_368#_M1017_d N_A_27_368#_M1013_s
+ N_A_27_368#_c_485_n N_A_27_368#_c_486_n N_A_27_368#_c_499_n
+ N_A_27_368#_c_487_n N_A_27_368#_c_504_n N_A_27_368#_c_509_n
+ N_A_27_368#_c_488_n N_A_27_368#_c_511_n N_A_27_368#_c_489_n
+ N_A_27_368#_c_490_n N_A_27_368#_c_491_n N_A_27_368#_c_518_n
+ N_A_27_368#_c_520_n N_A_27_368#_c_521_n N_A_27_368#_c_492_n
+ PM_SKY130_FD_SC_HS__NOR3_4%A_27_368#
x_PM_SKY130_FD_SC_HS__NOR3_4%VPWR N_VPWR_M1005_d N_VPWR_M1012_d N_VPWR_c_574_n
+ N_VPWR_c_575_n VPWR N_VPWR_c_576_n N_VPWR_c_577_n N_VPWR_c_578_n
+ N_VPWR_c_573_n N_VPWR_c_580_n N_VPWR_c_581_n PM_SKY130_FD_SC_HS__NOR3_4%VPWR
x_PM_SKY130_FD_SC_HS__NOR3_4%A_295_368# N_A_295_368#_M1003_s
+ N_A_295_368#_M1002_d N_A_295_368#_M1009_d N_A_295_368#_M1015_s
+ N_A_295_368#_c_642_n N_A_295_368#_c_643_n N_A_295_368#_c_656_n
+ N_A_295_368#_c_644_n PM_SKY130_FD_SC_HS__NOR3_4%A_295_368#
x_PM_SKY130_FD_SC_HS__NOR3_4%Y N_Y_M1004_s N_Y_M1007_d N_Y_M1001_d N_Y_M1000_s
+ N_Y_M1008_s N_Y_c_688_n N_Y_c_689_n N_Y_c_690_n N_Y_c_727_n N_Y_c_691_n
+ N_Y_c_692_n N_Y_c_696_n N_Y_c_693_n N_Y_c_694_n N_Y_c_746_n N_Y_c_697_n
+ N_Y_c_698_n Y PM_SKY130_FD_SC_HS__NOR3_4%Y
x_PM_SKY130_FD_SC_HS__NOR3_4%VGND N_VGND_M1004_d N_VGND_M1016_d N_VGND_M1011_s
+ N_VGND_M1010_s N_VGND_c_806_n N_VGND_c_807_n N_VGND_c_808_n N_VGND_c_809_n
+ N_VGND_c_810_n N_VGND_c_811_n VGND N_VGND_c_812_n N_VGND_c_813_n
+ N_VGND_c_814_n N_VGND_c_815_n N_VGND_c_816_n N_VGND_c_817_n N_VGND_c_818_n
+ PM_SKY130_FD_SC_HS__NOR3_4%VGND
cc_1 VNB N_A_M1004_g 0.0307057f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_2 VNB N_A_M1016_g 0.024721f $X=-0.19 $Y=-0.245 $X2=0.935 $Y2=0.74
cc_3 VNB N_A_c_110_n 0.00103091f $X=-0.19 $Y=-0.245 $X2=0.77 $Y2=1.515
cc_4 VNB N_A_c_111_n 0.0027193f $X=-0.19 $Y=-0.245 $X2=5.97 $Y2=0.495
cc_5 VNB N_A_c_112_n 0.16813f $X=-0.19 $Y=-0.245 $X2=5.97 $Y2=0.495
cc_6 VNB N_A_c_113_n 0.0357942f $X=-0.19 $Y=-0.245 $X2=5.97 $Y2=1.515
cc_7 VNB N_A_c_114_n 0.0478585f $X=-0.19 $Y=-0.245 $X2=0.935 $Y2=1.557
cc_8 VNB N_B_c_246_n 0.0147148f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_9 VNB N_B_c_247_n 0.0114101f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_10 VNB N_B_c_248_n 0.0156992f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=2.4
cc_11 VNB N_B_c_249_n 0.0193149f $X=-0.19 $Y=-0.245 $X2=0.935 $Y2=0.74
cc_12 VNB N_B_c_250_n 0.0161096f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_B_c_251_n 0.00903762f $X=-0.19 $Y=-0.245 $X2=5.775 $Y2=1.765
cc_14 VNB N_B_c_252_n 0.00789458f $X=-0.19 $Y=-0.245 $X2=6.225 $Y2=2.4
cc_15 VNB N_B_c_253_n 0.00773158f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_B_c_254_n 0.0110988f $X=-0.19 $Y=-0.245 $X2=4.02 $Y2=2.105
cc_17 VNB N_B_c_255_n 0.0256494f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_B_c_256_n 0.0861866f $X=-0.19 $Y=-0.245 $X2=0.77 $Y2=1.557
cc_19 VNB N_B_c_257_n 0.0037819f $X=-0.19 $Y=-0.245 $X2=0.95 $Y2=1.557
cc_20 VNB N_B_c_258_n 0.00684755f $X=-0.19 $Y=-0.245 $X2=6 $Y2=1.515
cc_21 VNB N_B_c_259_n 0.00930406f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_B_c_260_n 0.00306353f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_C_c_372_n 0.00838125f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_C_c_373_n 0.00549055f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=1.765
cc_25 VNB N_C_M1001_g 0.0363229f $X=-0.19 $Y=-0.245 $X2=0.935 $Y2=1.35
cc_26 VNB N_C_c_375_n 0.00208586f $X=-0.19 $Y=-0.245 $X2=0.95 $Y2=2.4
cc_27 VNB N_C_c_376_n 0.00214066f $X=-0.19 $Y=-0.245 $X2=0.95 $Y2=2.4
cc_28 VNB N_C_M1010_g 0.0396304f $X=-0.19 $Y=-0.245 $X2=5.775 $Y2=2.4
cc_29 VNB N_C_c_378_n 0.00960643f $X=-0.19 $Y=-0.245 $X2=0.77 $Y2=1.515
cc_30 VNB N_C_c_379_n 0.00730873f $X=-0.19 $Y=-0.245 $X2=0.77 $Y2=1.515
cc_31 VNB N_C_c_380_n 0.00435531f $X=-0.19 $Y=-0.245 $X2=5.97 $Y2=0.495
cc_32 VNB N_C_c_381_n 0.0732211f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_C_c_382_n 0.0194928f $X=-0.19 $Y=-0.245 $X2=5.97 $Y2=1.515
cc_34 VNB C 0.00924763f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_C_c_384_n 0.14102f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_VPWR_c_573_n 0.283096f $X=-0.19 $Y=-0.245 $X2=5.97 $Y2=0.495
cc_37 VNB N_Y_c_688_n 0.0103011f $X=-0.19 $Y=-0.245 $X2=5.775 $Y2=2.4
cc_38 VNB N_Y_c_689_n 0.00348993f $X=-0.19 $Y=-0.245 $X2=5.775 $Y2=2.4
cc_39 VNB N_Y_c_690_n 0.00240191f $X=-0.19 $Y=-0.245 $X2=6.225 $Y2=2.4
cc_40 VNB N_Y_c_691_n 0.0024006f $X=-0.19 $Y=-0.245 $X2=5.97 $Y2=2.02
cc_41 VNB N_Y_c_692_n 0.0314239f $X=-0.19 $Y=-0.245 $X2=5.97 $Y2=0.495
cc_42 VNB N_Y_c_693_n 0.00896499f $X=-0.19 $Y=-0.245 $X2=5.97 $Y2=1.515
cc_43 VNB N_Y_c_694_n 0.00226854f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB Y 0.00248769f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_VGND_c_806_n 0.010678f $X=-0.19 $Y=-0.245 $X2=0.95 $Y2=2.4
cc_46 VNB N_VGND_c_807_n 0.0505972f $X=-0.19 $Y=-0.245 $X2=5.775 $Y2=1.765
cc_47 VNB N_VGND_c_808_n 0.00900483f $X=-0.19 $Y=-0.245 $X2=6.225 $Y2=2.4
cc_48 VNB N_VGND_c_809_n 0.00900728f $X=-0.19 $Y=-0.245 $X2=0.77 $Y2=1.515
cc_49 VNB N_VGND_c_810_n 0.019013f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_VGND_c_811_n 0.0120529f $X=-0.19 $Y=-0.245 $X2=4.02 $Y2=2.105
cc_51 VNB N_VGND_c_812_n 0.019013f $X=-0.19 $Y=-0.245 $X2=5.97 $Y2=0.495
cc_52 VNB N_VGND_c_813_n 0.0186948f $X=-0.19 $Y=-0.245 $X2=3.935 $Y2=2.105
cc_53 VNB N_VGND_c_814_n 0.0915322f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_VGND_c_815_n 0.388363f $X=-0.19 $Y=-0.245 $X2=6 $Y2=1.395
cc_55 VNB N_VGND_c_816_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0.935 $Y2=1.557
cc_56 VNB N_VGND_c_817_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=1.625 $Y2=2.045
cc_57 VNB N_VGND_c_818_n 0.00596278f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VPB N_A_c_115_n 0.0198916f $X=-0.19 $Y=1.66 $X2=0.5 $Y2=1.765
cc_59 VPB N_A_c_116_n 0.0151062f $X=-0.19 $Y=1.66 $X2=0.95 $Y2=1.765
cc_60 VPB N_A_c_117_n 0.0150909f $X=-0.19 $Y=1.66 $X2=5.775 $Y2=1.765
cc_61 VPB N_A_c_118_n 0.0198913f $X=-0.19 $Y=1.66 $X2=6.225 $Y2=1.765
cc_62 VPB N_A_c_110_n 0.00149582f $X=-0.19 $Y=1.66 $X2=0.77 $Y2=1.515
cc_63 VPB N_A_c_111_n 0.00149165f $X=-0.19 $Y=1.66 $X2=5.97 $Y2=0.495
cc_64 VPB N_A_c_113_n 0.0241722f $X=-0.19 $Y=1.66 $X2=5.97 $Y2=1.515
cc_65 VPB N_A_c_114_n 0.0239136f $X=-0.19 $Y=1.66 $X2=0.935 $Y2=1.557
cc_66 VPB N_B_c_247_n 0.0289938f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.74
cc_67 VPB N_B_c_251_n 8.49173e-19 $X=-0.19 $Y=1.66 $X2=5.775 $Y2=1.765
cc_68 VPB N_B_c_263_n 0.0206111f $X=-0.19 $Y=1.66 $X2=5.775 $Y2=2.4
cc_69 VPB N_B_c_252_n 7.41773e-19 $X=-0.19 $Y=1.66 $X2=6.225 $Y2=2.4
cc_70 VPB N_B_c_265_n 0.0190288f $X=-0.19 $Y=1.66 $X2=0.77 $Y2=1.92
cc_71 VPB N_B_c_253_n 7.26457e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_72 VPB N_B_c_267_n 0.0206215f $X=-0.19 $Y=1.66 $X2=3.85 $Y2=2.255
cc_73 VPB N_B_c_268_n 0.00155728f $X=-0.19 $Y=1.66 $X2=5.97 $Y2=1.515
cc_74 VPB N_C_c_385_n 0.0169332f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.35
cc_75 VPB N_C_c_372_n 0.0107554f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_76 VPB N_C_c_373_n 0.00960415f $X=-0.19 $Y=1.66 $X2=0.5 $Y2=1.765
cc_77 VPB N_C_c_388_n 0.0161554f $X=-0.19 $Y=1.66 $X2=0.935 $Y2=0.74
cc_78 VPB N_C_c_375_n 0.00528909f $X=-0.19 $Y=1.66 $X2=0.95 $Y2=2.4
cc_79 VPB N_C_c_376_n 0.0106858f $X=-0.19 $Y=1.66 $X2=0.95 $Y2=2.4
cc_80 VPB N_C_c_391_n 0.0161554f $X=-0.19 $Y=1.66 $X2=6.225 $Y2=2.4
cc_81 VPB N_C_c_378_n 0.0162707f $X=-0.19 $Y=1.66 $X2=0.77 $Y2=1.515
cc_82 VPB N_C_c_379_n 0.0170207f $X=-0.19 $Y=1.66 $X2=0.77 $Y2=1.515
cc_83 VPB N_C_c_394_n 0.0161691f $X=-0.19 $Y=1.66 $X2=0.77 $Y2=1.515
cc_84 VPB N_C_c_380_n 0.00699923f $X=-0.19 $Y=1.66 $X2=5.97 $Y2=0.495
cc_85 VPB N_A_27_368#_c_485_n 0.0295533f $X=-0.19 $Y=1.66 $X2=6.225 $Y2=1.765
cc_86 VPB N_A_27_368#_c_486_n 0.0197262f $X=-0.19 $Y=1.66 $X2=0.77 $Y2=1.515
cc_87 VPB N_A_27_368#_c_487_n 0.00216775f $X=-0.19 $Y=1.66 $X2=5.805 $Y2=2.105
cc_88 VPB N_A_27_368#_c_488_n 0.00212741f $X=-0.19 $Y=1.66 $X2=5.97 $Y2=1.515
cc_89 VPB N_A_27_368#_c_489_n 0.0303846f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.95
cc_90 VPB N_A_27_368#_c_490_n 0.0190674f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_91 VPB N_A_27_368#_c_491_n 0.00708086f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_92 VPB N_A_27_368#_c_492_n 0.0071123f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_93 VPB N_VPWR_c_574_n 0.00396467f $X=-0.19 $Y=1.66 $X2=0.935 $Y2=0.74
cc_94 VPB N_VPWR_c_575_n 0.00396467f $X=-0.19 $Y=1.66 $X2=0.95 $Y2=2.4
cc_95 VPB N_VPWR_c_576_n 0.0178682f $X=-0.19 $Y=1.66 $X2=5.775 $Y2=2.4
cc_96 VPB N_VPWR_c_577_n 0.116818f $X=-0.19 $Y=1.66 $X2=0.77 $Y2=1.515
cc_97 VPB N_VPWR_c_578_n 0.0177091f $X=-0.19 $Y=1.66 $X2=5.97 $Y2=0.495
cc_98 VPB N_VPWR_c_573_n 0.0774077f $X=-0.19 $Y=1.66 $X2=5.97 $Y2=0.495
cc_99 VPB N_VPWR_c_580_n 0.00601644f $X=-0.19 $Y=1.66 $X2=5.97 $Y2=1.515
cc_100 VPB N_VPWR_c_581_n 0.00601813f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_101 VPB N_A_295_368#_c_642_n 0.0110966f $X=-0.19 $Y=1.66 $X2=0.95 $Y2=2.4
cc_102 VPB N_A_295_368#_c_643_n 0.00259172f $X=-0.19 $Y=1.66 $X2=0.77 $Y2=1.92
cc_103 VPB N_A_295_368#_c_644_n 0.00216178f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_104 VPB N_Y_c_696_n 0.00849352f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_105 VPB N_Y_c_697_n 0.00688612f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_106 VPB N_Y_c_698_n 5.90677e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_107 N_A_c_110_n N_B_c_246_n 0.00151667f $X=0.77 $Y=1.515 $X2=0 $Y2=0
cc_108 N_A_c_114_n N_B_c_246_n 0.0200095f $X=0.935 $Y=1.557 $X2=0 $Y2=0
cc_109 N_A_c_116_n N_B_c_247_n 0.0244645f $X=0.95 $Y=1.765 $X2=0 $Y2=0
cc_110 N_A_c_110_n N_B_c_247_n 7.91761e-19 $X=0.77 $Y=1.515 $X2=0 $Y2=0
cc_111 A N_B_c_247_n 0.00443308f $X=1.595 $Y=1.95 $X2=0 $Y2=0
cc_112 N_A_c_128_p N_B_c_247_n 0.0154871f $X=1.625 $Y=2.045 $X2=0 $Y2=0
cc_113 N_A_M1016_g N_B_c_248_n 0.0209692f $X=0.935 $Y=0.74 $X2=0 $Y2=0
cc_114 N_A_c_130_p N_B_c_263_n 0.011766f $X=5.805 $Y=2.105 $X2=0 $Y2=0
cc_115 N_A_c_131_p N_B_c_263_n 0.0029335f $X=3.935 $Y=2.105 $X2=0 $Y2=0
cc_116 N_A_c_130_p N_B_c_265_n 0.0107326f $X=5.805 $Y=2.105 $X2=0 $Y2=0
cc_117 N_A_c_113_n N_B_c_253_n 0.011057f $X=5.97 $Y=1.515 $X2=0 $Y2=0
cc_118 N_A_c_117_n N_B_c_267_n 0.0249034f $X=5.775 $Y=1.765 $X2=0 $Y2=0
cc_119 N_A_c_130_p N_B_c_267_n 0.0135807f $X=5.805 $Y=2.105 $X2=0 $Y2=0
cc_120 N_A_c_111_n N_B_c_267_n 0.00110585f $X=5.97 $Y=0.495 $X2=0 $Y2=0
cc_121 N_A_c_113_n N_B_c_267_n 0.00340713f $X=5.97 $Y=1.515 $X2=0 $Y2=0
cc_122 N_A_M1016_g N_B_c_254_n 0.00879955f $X=0.935 $Y=0.74 $X2=0 $Y2=0
cc_123 N_A_c_110_n N_B_c_268_n 0.0130906f $X=0.77 $Y=1.515 $X2=0 $Y2=0
cc_124 A N_B_c_268_n 7.95053e-19 $X=1.595 $Y=1.95 $X2=0 $Y2=0
cc_125 N_A_c_114_n N_B_c_268_n 0.00150439f $X=0.935 $Y=1.557 $X2=0 $Y2=0
cc_126 N_A_c_128_p N_B_c_268_n 0.0158741f $X=1.625 $Y=2.045 $X2=0 $Y2=0
cc_127 N_A_c_111_n N_B_c_256_n 0.00218149f $X=5.97 $Y=0.495 $X2=0 $Y2=0
cc_128 N_A_c_112_n N_B_c_256_n 0.011057f $X=5.97 $Y=0.495 $X2=0 $Y2=0
cc_129 N_A_c_145_p N_B_c_259_n 0.00790273f $X=3.85 $Y=2.255 $X2=0 $Y2=0
cc_130 A N_B_c_259_n 0.00663543f $X=1.595 $Y=1.95 $X2=0 $Y2=0
cc_131 N_A_c_145_p N_C_c_385_n 0.0130085f $X=3.85 $Y=2.255 $X2=-0.19 $Y2=-0.245
cc_132 A N_C_c_385_n 0.00510773f $X=1.595 $Y=1.95 $X2=-0.19 $Y2=-0.245
cc_133 N_A_c_145_p N_C_c_372_n 9.66579e-19 $X=3.85 $Y=2.255 $X2=0 $Y2=0
cc_134 N_A_c_145_p N_C_c_388_n 0.0122132f $X=3.85 $Y=2.255 $X2=0 $Y2=0
cc_135 N_A_c_145_p N_C_c_391_n 0.0122132f $X=3.85 $Y=2.255 $X2=0 $Y2=0
cc_136 N_A_c_131_p N_C_c_391_n 7.80042e-19 $X=3.935 $Y=2.105 $X2=0 $Y2=0
cc_137 N_A_c_145_p N_C_c_378_n 0.00133602f $X=3.85 $Y=2.255 $X2=0 $Y2=0
cc_138 N_A_c_145_p N_C_c_394_n 0.00873106f $X=3.85 $Y=2.255 $X2=0 $Y2=0
cc_139 N_A_c_130_p N_C_c_394_n 3.09461e-19 $X=5.805 $Y=2.105 $X2=0 $Y2=0
cc_140 N_A_c_131_p N_C_c_394_n 0.00866814f $X=3.935 $Y=2.105 $X2=0 $Y2=0
cc_141 N_A_c_111_n C 0.0276579f $X=5.97 $Y=0.495 $X2=0 $Y2=0
cc_142 N_A_c_112_n C 0.00275385f $X=5.97 $Y=0.495 $X2=0 $Y2=0
cc_143 N_A_c_111_n N_C_c_384_n 2.67785e-19 $X=5.97 $Y=0.495 $X2=0 $Y2=0
cc_144 N_A_c_112_n N_C_c_384_n 0.0179842f $X=5.97 $Y=0.495 $X2=0 $Y2=0
cc_145 N_A_c_128_p N_A_27_368#_M1006_s 0.0094261f $X=1.625 $Y=2.045 $X2=0 $Y2=0
cc_146 N_A_c_130_p N_A_27_368#_M1014_d 0.00384479f $X=5.805 $Y=2.105 $X2=0 $Y2=0
cc_147 N_A_c_130_p N_A_27_368#_M1017_d 0.00907456f $X=5.805 $Y=2.105 $X2=0 $Y2=0
cc_148 N_A_c_115_n N_A_27_368#_c_485_n 0.00588726f $X=0.5 $Y=1.765 $X2=0 $Y2=0
cc_149 N_A_c_110_n N_A_27_368#_c_485_n 0.00358027f $X=0.77 $Y=1.515 $X2=0 $Y2=0
cc_150 N_A_c_115_n N_A_27_368#_c_486_n 0.00547771f $X=0.5 $Y=1.765 $X2=0 $Y2=0
cc_151 N_A_c_115_n N_A_27_368#_c_499_n 0.01427f $X=0.5 $Y=1.765 $X2=0 $Y2=0
cc_152 N_A_c_116_n N_A_27_368#_c_499_n 0.00975433f $X=0.95 $Y=1.765 $X2=0 $Y2=0
cc_153 N_A_c_169_p N_A_27_368#_c_499_n 0.0196611f $X=0.77 $Y=1.92 $X2=0 $Y2=0
cc_154 N_A_c_114_n N_A_27_368#_c_499_n 6.0988e-19 $X=0.935 $Y=1.557 $X2=0 $Y2=0
cc_155 N_A_c_128_p N_A_27_368#_c_499_n 0.00681496f $X=1.625 $Y=2.045 $X2=0 $Y2=0
cc_156 N_A_c_145_p N_A_27_368#_c_504_n 0.117563f $X=3.85 $Y=2.255 $X2=0 $Y2=0
cc_157 N_A_c_130_p N_A_27_368#_c_504_n 0.0179717f $X=5.805 $Y=2.105 $X2=0 $Y2=0
cc_158 N_A_c_131_p N_A_27_368#_c_504_n 0.00830881f $X=3.935 $Y=2.105 $X2=0 $Y2=0
cc_159 A N_A_27_368#_c_504_n 0.0131482f $X=1.595 $Y=1.95 $X2=0 $Y2=0
cc_160 N_A_c_128_p N_A_27_368#_c_504_n 0.00958959f $X=1.625 $Y=2.045 $X2=0 $Y2=0
cc_161 N_A_c_130_p N_A_27_368#_c_509_n 0.0349019f $X=5.805 $Y=2.105 $X2=0 $Y2=0
cc_162 N_A_c_117_n N_A_27_368#_c_488_n 0.00440717f $X=5.775 $Y=1.765 $X2=0 $Y2=0
cc_163 N_A_c_117_n N_A_27_368#_c_511_n 0.00969265f $X=5.775 $Y=1.765 $X2=0 $Y2=0
cc_164 N_A_c_118_n N_A_27_368#_c_511_n 0.0142588f $X=6.225 $Y=1.765 $X2=0 $Y2=0
cc_165 N_A_c_130_p N_A_27_368#_c_511_n 0.0261124f $X=5.805 $Y=2.105 $X2=0 $Y2=0
cc_166 N_A_c_113_n N_A_27_368#_c_511_n 6.12681e-19 $X=5.97 $Y=1.515 $X2=0 $Y2=0
cc_167 N_A_c_118_n N_A_27_368#_c_489_n 0.00588736f $X=6.225 $Y=1.765 $X2=0 $Y2=0
cc_168 N_A_c_111_n N_A_27_368#_c_489_n 0.00682412f $X=5.97 $Y=0.495 $X2=0 $Y2=0
cc_169 N_A_c_118_n N_A_27_368#_c_490_n 0.00540876f $X=6.225 $Y=1.765 $X2=0 $Y2=0
cc_170 N_A_c_116_n N_A_27_368#_c_518_n 0.00475181f $X=0.95 $Y=1.765 $X2=0 $Y2=0
cc_171 N_A_c_128_p N_A_27_368#_c_518_n 0.0157617f $X=1.625 $Y=2.045 $X2=0 $Y2=0
cc_172 N_A_c_130_p N_A_27_368#_c_520_n 0.0147062f $X=5.805 $Y=2.105 $X2=0 $Y2=0
cc_173 N_A_c_130_p N_A_27_368#_c_521_n 0.0137635f $X=5.805 $Y=2.105 $X2=0 $Y2=0
cc_174 N_A_c_169_p N_VPWR_M1005_d 0.00288301f $X=0.77 $Y=1.92 $X2=-0.19
+ $Y2=-0.245
cc_175 N_A_c_130_p N_VPWR_M1012_d 0.0026248f $X=5.805 $Y=2.105 $X2=0 $Y2=0
cc_176 N_A_c_111_n N_VPWR_M1012_d 4.83872e-19 $X=5.97 $Y=0.495 $X2=0 $Y2=0
cc_177 N_A_c_115_n N_VPWR_c_574_n 0.00991225f $X=0.5 $Y=1.765 $X2=0 $Y2=0
cc_178 N_A_c_116_n N_VPWR_c_574_n 0.00722226f $X=0.95 $Y=1.765 $X2=0 $Y2=0
cc_179 N_A_c_117_n N_VPWR_c_575_n 0.00676092f $X=5.775 $Y=1.765 $X2=0 $Y2=0
cc_180 N_A_c_118_n N_VPWR_c_575_n 0.00969781f $X=6.225 $Y=1.765 $X2=0 $Y2=0
cc_181 N_A_c_115_n N_VPWR_c_576_n 0.00413917f $X=0.5 $Y=1.765 $X2=0 $Y2=0
cc_182 N_A_c_116_n N_VPWR_c_577_n 0.00413917f $X=0.95 $Y=1.765 $X2=0 $Y2=0
cc_183 N_A_c_117_n N_VPWR_c_577_n 0.00413917f $X=5.775 $Y=1.765 $X2=0 $Y2=0
cc_184 N_A_c_118_n N_VPWR_c_578_n 0.00413917f $X=6.225 $Y=1.765 $X2=0 $Y2=0
cc_185 N_A_c_115_n N_VPWR_c_573_n 0.00413459f $X=0.5 $Y=1.765 $X2=0 $Y2=0
cc_186 N_A_c_116_n N_VPWR_c_573_n 0.00410066f $X=0.95 $Y=1.765 $X2=0 $Y2=0
cc_187 N_A_c_117_n N_VPWR_c_573_n 0.00405533f $X=5.775 $Y=1.765 $X2=0 $Y2=0
cc_188 N_A_c_118_n N_VPWR_c_573_n 0.0040891f $X=6.225 $Y=1.765 $X2=0 $Y2=0
cc_189 N_A_c_145_p N_A_295_368#_M1003_s 0.00287876f $X=3.85 $Y=2.255 $X2=-0.19
+ $Y2=-0.245
cc_190 A N_A_295_368#_M1003_s 0.0123756f $X=1.595 $Y=1.95 $X2=-0.19 $Y2=-0.245
cc_191 N_A_c_128_p N_A_295_368#_M1003_s 0.00294192f $X=1.625 $Y=2.045 $X2=-0.19
+ $Y2=-0.245
cc_192 N_A_c_145_p N_A_295_368#_M1002_d 0.00786725f $X=3.85 $Y=2.255 $X2=0 $Y2=0
cc_193 N_A_c_130_p N_A_295_368#_M1009_d 0.00814261f $X=5.805 $Y=2.105 $X2=0
+ $Y2=0
cc_194 N_A_c_131_p N_A_295_368#_M1009_d 0.00398493f $X=3.935 $Y=2.105 $X2=0
+ $Y2=0
cc_195 N_A_c_130_p N_A_295_368#_M1015_s 0.00384909f $X=5.805 $Y=2.105 $X2=0
+ $Y2=0
cc_196 N_A_c_117_n N_A_295_368#_c_644_n 3.12716e-19 $X=5.775 $Y=1.765 $X2=0
+ $Y2=0
cc_197 N_A_c_145_p N_Y_M1000_s 0.00751361f $X=3.85 $Y=2.255 $X2=0 $Y2=0
cc_198 N_A_c_145_p N_Y_M1008_s 0.0075174f $X=3.85 $Y=2.255 $X2=0 $Y2=0
cc_199 N_A_M1016_g N_Y_c_688_n 0.0148128f $X=0.935 $Y=0.74 $X2=0 $Y2=0
cc_200 N_A_c_110_n N_Y_c_688_n 0.00446029f $X=0.77 $Y=1.515 $X2=0 $Y2=0
cc_201 N_A_c_114_n N_Y_c_688_n 0.00120237f $X=0.935 $Y=1.557 $X2=0 $Y2=0
cc_202 N_A_M1004_g N_Y_c_689_n 0.00582181f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_203 N_A_M1016_g N_Y_c_689_n 0.00129659f $X=0.935 $Y=0.74 $X2=0 $Y2=0
cc_204 N_A_c_110_n N_Y_c_689_n 0.0239178f $X=0.77 $Y=1.515 $X2=0 $Y2=0
cc_205 N_A_c_114_n N_Y_c_689_n 8.70621e-19 $X=0.935 $Y=1.557 $X2=0 $Y2=0
cc_206 N_A_M1016_g N_Y_c_690_n 6.36864e-19 $X=0.935 $Y=0.74 $X2=0 $Y2=0
cc_207 N_A_c_111_n N_Y_c_692_n 0.00639395f $X=5.97 $Y=0.495 $X2=0 $Y2=0
cc_208 N_A_c_112_n N_Y_c_692_n 0.00389741f $X=5.97 $Y=0.495 $X2=0 $Y2=0
cc_209 N_A_c_145_p N_Y_c_696_n 0.00456214f $X=3.85 $Y=2.255 $X2=0 $Y2=0
cc_210 N_A_c_130_p N_Y_c_696_n 0.071842f $X=5.805 $Y=2.105 $X2=0 $Y2=0
cc_211 N_A_c_111_n N_Y_c_696_n 0.00557926f $X=5.97 $Y=0.495 $X2=0 $Y2=0
cc_212 N_A_c_113_n N_Y_c_696_n 5.18523e-19 $X=5.97 $Y=1.515 $X2=0 $Y2=0
cc_213 N_A_c_131_p N_Y_c_696_n 0.00830881f $X=3.935 $Y=2.105 $X2=0 $Y2=0
cc_214 N_A_c_111_n N_Y_c_693_n 0.0204114f $X=5.97 $Y=0.495 $X2=0 $Y2=0
cc_215 N_A_c_112_n N_Y_c_693_n 0.00555926f $X=5.97 $Y=0.495 $X2=0 $Y2=0
cc_216 N_A_c_145_p N_Y_c_697_n 0.0970067f $X=3.85 $Y=2.255 $X2=0 $Y2=0
cc_217 A N_Y_c_697_n 0.00380783f $X=1.595 $Y=1.95 $X2=0 $Y2=0
cc_218 N_A_M1004_g Y 0.00840664f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_219 N_A_M1016_g Y 0.00914611f $X=0.935 $Y=0.74 $X2=0 $Y2=0
cc_220 N_A_M1004_g N_VGND_c_807_n 0.00647381f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_221 N_A_M1016_g N_VGND_c_808_n 0.00625757f $X=0.935 $Y=0.74 $X2=0 $Y2=0
cc_222 N_A_M1004_g N_VGND_c_812_n 0.00434272f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_223 N_A_M1016_g N_VGND_c_812_n 0.00445602f $X=0.935 $Y=0.74 $X2=0 $Y2=0
cc_224 N_A_c_111_n N_VGND_c_814_n 0.0148959f $X=5.97 $Y=0.495 $X2=0 $Y2=0
cc_225 N_A_c_112_n N_VGND_c_814_n 0.0101867f $X=5.97 $Y=0.495 $X2=0 $Y2=0
cc_226 N_A_M1004_g N_VGND_c_815_n 0.00824041f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_227 N_A_M1016_g N_VGND_c_815_n 0.00857802f $X=0.935 $Y=0.74 $X2=0 $Y2=0
cc_228 N_A_c_111_n N_VGND_c_815_n 0.0120047f $X=5.97 $Y=0.495 $X2=0 $Y2=0
cc_229 N_A_c_112_n N_VGND_c_815_n 0.00834893f $X=5.97 $Y=0.495 $X2=0 $Y2=0
cc_230 N_B_c_247_n N_C_c_385_n 0.0309323f $X=1.4 $Y=1.765 $X2=-0.19 $Y2=-0.245
cc_231 N_B_c_258_n N_C_c_372_n 0.00642948f $X=2.215 $Y=1.35 $X2=0 $Y2=0
cc_232 N_B_c_247_n N_C_c_373_n 0.0102931f $X=1.4 $Y=1.765 $X2=0 $Y2=0
cc_233 N_B_c_249_n N_C_c_373_n 0.00550534f $X=1.85 $Y=1.26 $X2=0 $Y2=0
cc_234 N_B_c_268_n N_C_c_373_n 0.00100564f $X=1.475 $Y=1.435 $X2=0 $Y2=0
cc_235 N_B_c_259_n N_C_c_373_n 0.00642948f $X=2.045 $Y=1.35 $X2=0 $Y2=0
cc_236 N_B_c_250_n N_C_M1001_g 0.0257968f $X=1.925 $Y=1.185 $X2=0 $Y2=0
cc_237 N_B_c_257_n N_C_M1001_g 0.0194702f $X=2.585 $Y=1.35 $X2=0 $Y2=0
cc_238 N_B_c_260_n N_C_c_376_n 0.0024922f $X=2.755 $Y=1.35 $X2=0 $Y2=0
cc_239 N_B_c_255_n N_C_M1010_g 0.0203249f $X=4.8 $Y=1.345 $X2=0 $Y2=0
cc_240 N_B_c_260_n N_C_M1010_g 2.71203e-19 $X=2.755 $Y=1.35 $X2=0 $Y2=0
cc_241 N_B_c_255_n N_C_c_379_n 0.0148196f $X=4.8 $Y=1.345 $X2=0 $Y2=0
cc_242 N_B_c_263_n N_C_c_394_n 0.0326923f $X=4.425 $Y=1.765 $X2=0 $Y2=0
cc_243 N_B_c_263_n N_C_c_380_n 0.00431398f $X=4.425 $Y=1.765 $X2=0 $Y2=0
cc_244 N_B_c_251_n N_C_c_381_n 0.00431398f $X=4.425 $Y=1.675 $X2=0 $Y2=0
cc_245 N_B_c_255_n N_C_c_381_n 0.0216801f $X=4.8 $Y=1.345 $X2=0 $Y2=0
cc_246 N_B_c_256_n N_C_c_381_n 0.00958311f $X=5.325 $Y=1.345 $X2=0 $Y2=0
cc_247 N_B_c_256_n C 0.00104974f $X=5.325 $Y=1.345 $X2=0 $Y2=0
cc_248 N_B_c_256_n N_C_c_384_n 0.0204898f $X=5.325 $Y=1.345 $X2=0 $Y2=0
cc_249 N_B_c_247_n N_A_27_368#_c_487_n 0.004986f $X=1.4 $Y=1.765 $X2=0 $Y2=0
cc_250 N_B_c_247_n N_A_27_368#_c_504_n 0.0110965f $X=1.4 $Y=1.765 $X2=0 $Y2=0
cc_251 N_B_c_263_n N_A_27_368#_c_504_n 0.0105921f $X=4.425 $Y=1.765 $X2=0 $Y2=0
cc_252 N_B_c_265_n N_A_27_368#_c_509_n 0.00951207f $X=4.875 $Y=1.765 $X2=0 $Y2=0
cc_253 N_B_c_267_n N_A_27_368#_c_509_n 0.00965708f $X=5.325 $Y=1.765 $X2=0 $Y2=0
cc_254 N_B_c_267_n N_A_27_368#_c_488_n 0.00440717f $X=5.325 $Y=1.765 $X2=0 $Y2=0
cc_255 N_B_c_247_n N_A_27_368#_c_518_n 0.00425721f $X=1.4 $Y=1.765 $X2=0 $Y2=0
cc_256 N_B_c_263_n N_A_27_368#_c_520_n 0.00515187f $X=4.425 $Y=1.765 $X2=0 $Y2=0
cc_257 N_B_c_247_n N_VPWR_c_574_n 4.74948e-19 $X=1.4 $Y=1.765 $X2=0 $Y2=0
cc_258 N_B_c_267_n N_VPWR_c_575_n 3.97026e-19 $X=5.325 $Y=1.765 $X2=0 $Y2=0
cc_259 N_B_c_247_n N_VPWR_c_577_n 0.00325313f $X=1.4 $Y=1.765 $X2=0 $Y2=0
cc_260 N_B_c_263_n N_VPWR_c_577_n 0.00278271f $X=4.425 $Y=1.765 $X2=0 $Y2=0
cc_261 N_B_c_265_n N_VPWR_c_577_n 0.00279479f $X=4.875 $Y=1.765 $X2=0 $Y2=0
cc_262 N_B_c_267_n N_VPWR_c_577_n 0.00444353f $X=5.325 $Y=1.765 $X2=0 $Y2=0
cc_263 N_B_c_247_n N_VPWR_c_573_n 0.00412334f $X=1.4 $Y=1.765 $X2=0 $Y2=0
cc_264 N_B_c_263_n N_VPWR_c_573_n 0.00354248f $X=4.425 $Y=1.765 $X2=0 $Y2=0
cc_265 N_B_c_265_n N_VPWR_c_573_n 0.00352913f $X=4.875 $Y=1.765 $X2=0 $Y2=0
cc_266 N_B_c_267_n N_VPWR_c_573_n 0.00445635f $X=5.325 $Y=1.765 $X2=0 $Y2=0
cc_267 N_B_c_247_n N_A_295_368#_c_642_n 0.00306738f $X=1.4 $Y=1.765 $X2=0 $Y2=0
cc_268 N_B_c_263_n N_A_295_368#_c_643_n 0.0103927f $X=4.425 $Y=1.765 $X2=0 $Y2=0
cc_269 N_B_c_265_n N_A_295_368#_c_643_n 0.00876256f $X=4.875 $Y=1.765 $X2=0
+ $Y2=0
cc_270 N_B_c_263_n N_A_295_368#_c_656_n 9.77496e-19 $X=4.425 $Y=1.765 $X2=0
+ $Y2=0
cc_271 N_B_c_263_n N_A_295_368#_c_644_n 7.8402e-19 $X=4.425 $Y=1.765 $X2=0 $Y2=0
cc_272 N_B_c_265_n N_A_295_368#_c_644_n 0.00585602f $X=4.875 $Y=1.765 $X2=0
+ $Y2=0
cc_273 N_B_c_267_n N_A_295_368#_c_644_n 0.00605224f $X=5.325 $Y=1.765 $X2=0
+ $Y2=0
cc_274 N_B_c_248_n N_Y_c_688_n 0.0128008f $X=1.495 $Y=1.185 $X2=0 $Y2=0
cc_275 N_B_c_254_n N_Y_c_688_n 0.00352001f $X=1.475 $Y=1.26 $X2=0 $Y2=0
cc_276 N_B_c_268_n N_Y_c_688_n 0.0172045f $X=1.475 $Y=1.435 $X2=0 $Y2=0
cc_277 N_B_c_248_n N_Y_c_690_n 0.00622488f $X=1.495 $Y=1.185 $X2=0 $Y2=0
cc_278 N_B_c_250_n N_Y_c_690_n 0.0079293f $X=1.925 $Y=1.185 $X2=0 $Y2=0
cc_279 N_B_c_250_n N_Y_c_727_n 0.0105176f $X=1.925 $Y=1.185 $X2=0 $Y2=0
cc_280 N_B_c_258_n N_Y_c_727_n 0.035669f $X=2.215 $Y=1.35 $X2=0 $Y2=0
cc_281 N_B_c_259_n N_Y_c_727_n 0.00635832f $X=2.045 $Y=1.35 $X2=0 $Y2=0
cc_282 N_B_c_250_n N_Y_c_691_n 5.95058e-19 $X=1.925 $Y=1.185 $X2=0 $Y2=0
cc_283 N_B_c_255_n N_Y_c_692_n 0.157951f $X=4.8 $Y=1.345 $X2=0 $Y2=0
cc_284 N_B_c_256_n N_Y_c_692_n 0.00908482f $X=5.325 $Y=1.345 $X2=0 $Y2=0
cc_285 N_B_c_263_n N_Y_c_696_n 0.0123387f $X=4.425 $Y=1.765 $X2=0 $Y2=0
cc_286 N_B_c_265_n N_Y_c_696_n 0.0116345f $X=4.875 $Y=1.765 $X2=0 $Y2=0
cc_287 N_B_c_267_n N_Y_c_696_n 0.00647517f $X=5.325 $Y=1.765 $X2=0 $Y2=0
cc_288 N_B_c_256_n N_Y_c_696_n 0.00509515f $X=5.325 $Y=1.345 $X2=0 $Y2=0
cc_289 N_B_c_252_n N_Y_c_693_n 0.00349655f $X=4.875 $Y=1.675 $X2=0 $Y2=0
cc_290 N_B_c_253_n N_Y_c_693_n 0.00436904f $X=5.325 $Y=1.675 $X2=0 $Y2=0
cc_291 N_B_c_255_n N_Y_c_693_n 0.0249855f $X=4.8 $Y=1.345 $X2=0 $Y2=0
cc_292 N_B_c_256_n N_Y_c_693_n 0.0172245f $X=5.325 $Y=1.345 $X2=0 $Y2=0
cc_293 N_B_c_248_n N_Y_c_694_n 0.00551466f $X=1.495 $Y=1.185 $X2=0 $Y2=0
cc_294 N_B_c_249_n N_Y_c_694_n 0.00245638f $X=1.85 $Y=1.26 $X2=0 $Y2=0
cc_295 N_B_c_250_n N_Y_c_694_n 0.00540275f $X=1.925 $Y=1.185 $X2=0 $Y2=0
cc_296 N_B_c_268_n N_Y_c_694_n 0.00777454f $X=1.475 $Y=1.435 $X2=0 $Y2=0
cc_297 N_B_c_259_n N_Y_c_694_n 0.0196452f $X=2.045 $Y=1.35 $X2=0 $Y2=0
cc_298 N_B_c_257_n N_Y_c_746_n 0.0229777f $X=2.585 $Y=1.35 $X2=0 $Y2=0
cc_299 N_B_c_255_n N_Y_c_697_n 0.0366801f $X=4.8 $Y=1.345 $X2=0 $Y2=0
cc_300 N_B_c_258_n N_Y_c_697_n 0.0392244f $X=2.215 $Y=1.35 $X2=0 $Y2=0
cc_301 N_B_c_255_n N_Y_c_698_n 0.122294f $X=4.8 $Y=1.345 $X2=0 $Y2=0
cc_302 N_B_c_248_n Y 6.20067e-19 $X=1.495 $Y=1.185 $X2=0 $Y2=0
cc_303 N_B_c_248_n N_VGND_c_808_n 0.00477239f $X=1.495 $Y=1.185 $X2=0 $Y2=0
cc_304 N_B_c_250_n N_VGND_c_809_n 0.00381161f $X=1.925 $Y=1.185 $X2=0 $Y2=0
cc_305 N_B_c_248_n N_VGND_c_813_n 0.00434272f $X=1.495 $Y=1.185 $X2=0 $Y2=0
cc_306 N_B_c_250_n N_VGND_c_813_n 0.00434272f $X=1.925 $Y=1.185 $X2=0 $Y2=0
cc_307 N_B_c_248_n N_VGND_c_815_n 0.00821239f $X=1.495 $Y=1.185 $X2=0 $Y2=0
cc_308 N_B_c_250_n N_VGND_c_815_n 0.0044609f $X=1.925 $Y=1.185 $X2=0 $Y2=0
cc_309 N_C_c_385_n N_A_27_368#_c_504_n 0.0120974f $X=2.005 $Y=1.765 $X2=0 $Y2=0
cc_310 N_C_c_388_n N_A_27_368#_c_504_n 0.0121912f $X=2.605 $Y=1.765 $X2=0 $Y2=0
cc_311 N_C_c_391_n N_A_27_368#_c_504_n 0.0121912f $X=3.215 $Y=1.765 $X2=0 $Y2=0
cc_312 N_C_c_394_n N_A_27_368#_c_504_n 0.0121008f $X=3.815 $Y=1.765 $X2=0 $Y2=0
cc_313 N_C_c_385_n N_A_27_368#_c_518_n 0.0015897f $X=2.005 $Y=1.765 $X2=0 $Y2=0
cc_314 N_C_c_394_n N_A_27_368#_c_520_n 9.87881e-19 $X=3.815 $Y=1.765 $X2=0 $Y2=0
cc_315 N_C_c_385_n N_VPWR_c_577_n 0.00278271f $X=2.005 $Y=1.765 $X2=0 $Y2=0
cc_316 N_C_c_388_n N_VPWR_c_577_n 0.00278271f $X=2.605 $Y=1.765 $X2=0 $Y2=0
cc_317 N_C_c_391_n N_VPWR_c_577_n 0.00278271f $X=3.215 $Y=1.765 $X2=0 $Y2=0
cc_318 N_C_c_394_n N_VPWR_c_577_n 0.00278271f $X=3.815 $Y=1.765 $X2=0 $Y2=0
cc_319 N_C_c_385_n N_VPWR_c_573_n 0.00356384f $X=2.005 $Y=1.765 $X2=0 $Y2=0
cc_320 N_C_c_388_n N_VPWR_c_573_n 0.00356415f $X=2.605 $Y=1.765 $X2=0 $Y2=0
cc_321 N_C_c_391_n N_VPWR_c_573_n 0.00356415f $X=3.215 $Y=1.765 $X2=0 $Y2=0
cc_322 N_C_c_394_n N_VPWR_c_573_n 0.00356417f $X=3.815 $Y=1.765 $X2=0 $Y2=0
cc_323 N_C_c_385_n N_A_295_368#_c_642_n 0.013127f $X=2.005 $Y=1.765 $X2=0 $Y2=0
cc_324 N_C_c_388_n N_A_295_368#_c_642_n 0.0135873f $X=2.605 $Y=1.765 $X2=0 $Y2=0
cc_325 N_C_c_391_n N_A_295_368#_c_642_n 0.0135873f $X=3.215 $Y=1.765 $X2=0 $Y2=0
cc_326 N_C_c_394_n N_A_295_368#_c_642_n 0.0133941f $X=3.815 $Y=1.765 $X2=0 $Y2=0
cc_327 N_C_M1001_g N_Y_c_690_n 5.99621e-19 $X=2.495 $Y=0.74 $X2=0 $Y2=0
cc_328 N_C_M1001_g N_Y_c_727_n 0.00917824f $X=2.495 $Y=0.74 $X2=0 $Y2=0
cc_329 N_C_M1001_g N_Y_c_691_n 0.00744777f $X=2.495 $Y=0.74 $X2=0 $Y2=0
cc_330 N_C_M1010_g N_Y_c_691_n 0.0115222f $X=2.925 $Y=0.74 $X2=0 $Y2=0
cc_331 N_C_M1010_g N_Y_c_692_n 0.0105704f $X=2.925 $Y=0.74 $X2=0 $Y2=0
cc_332 N_C_c_381_n N_Y_c_692_n 0.0148401f $X=3.815 $Y=1.545 $X2=0 $Y2=0
cc_333 C N_Y_c_692_n 0.112382f $X=5.435 $Y=0.47 $X2=0 $Y2=0
cc_334 N_C_c_384_n N_Y_c_692_n 0.0178347f $X=5.31 $Y=0.505 $X2=0 $Y2=0
cc_335 N_C_c_378_n N_Y_c_696_n 0.00139555f $X=3.725 $Y=1.62 $X2=0 $Y2=0
cc_336 N_C_c_394_n N_Y_c_696_n 0.0066238f $X=3.815 $Y=1.765 $X2=0 $Y2=0
cc_337 N_C_c_380_n N_Y_c_696_n 0.00675241f $X=3.815 $Y=1.62 $X2=0 $Y2=0
cc_338 N_C_M1001_g N_Y_c_694_n 8.58155e-19 $X=2.495 $Y=0.74 $X2=0 $Y2=0
cc_339 N_C_M1001_g N_Y_c_746_n 7.17169e-19 $X=2.495 $Y=0.74 $X2=0 $Y2=0
cc_340 N_C_M1010_g N_Y_c_746_n 7.17169e-19 $X=2.925 $Y=0.74 $X2=0 $Y2=0
cc_341 N_C_c_385_n N_Y_c_697_n 0.00625046f $X=2.005 $Y=1.765 $X2=0 $Y2=0
cc_342 N_C_c_372_n N_Y_c_697_n 0.00944381f $X=2.42 $Y=1.62 $X2=0 $Y2=0
cc_343 N_C_c_373_n N_Y_c_697_n 4.77037e-19 $X=2.095 $Y=1.62 $X2=0 $Y2=0
cc_344 N_C_c_388_n N_Y_c_697_n 0.012885f $X=2.605 $Y=1.765 $X2=0 $Y2=0
cc_345 N_C_c_375_n N_Y_c_697_n 0.0126832f $X=2.85 $Y=1.62 $X2=0 $Y2=0
cc_346 N_C_c_376_n N_Y_c_697_n 0.00402531f $X=2.695 $Y=1.62 $X2=0 $Y2=0
cc_347 N_C_c_391_n N_Y_c_697_n 0.0130459f $X=3.215 $Y=1.765 $X2=0 $Y2=0
cc_348 N_C_c_378_n N_Y_c_697_n 0.00102525f $X=3.725 $Y=1.62 $X2=0 $Y2=0
cc_349 N_C_c_379_n N_Y_c_697_n 0.00345577f $X=3.305 $Y=1.62 $X2=0 $Y2=0
cc_350 N_C_c_378_n N_Y_c_698_n 0.0107878f $X=3.725 $Y=1.62 $X2=0 $Y2=0
cc_351 N_C_c_379_n N_Y_c_698_n 0.00187408f $X=3.305 $Y=1.62 $X2=0 $Y2=0
cc_352 N_C_c_394_n N_Y_c_698_n 0.00499512f $X=3.815 $Y=1.765 $X2=0 $Y2=0
cc_353 N_C_M1001_g N_VGND_c_809_n 0.00519354f $X=2.495 $Y=0.74 $X2=0 $Y2=0
cc_354 N_C_M1001_g N_VGND_c_810_n 0.00434272f $X=2.495 $Y=0.74 $X2=0 $Y2=0
cc_355 N_C_M1010_g N_VGND_c_810_n 0.00434272f $X=2.925 $Y=0.74 $X2=0 $Y2=0
cc_356 N_C_M1010_g N_VGND_c_811_n 0.00500066f $X=2.925 $Y=0.74 $X2=0 $Y2=0
cc_357 N_C_c_382_n N_VGND_c_811_n 0.00758204f $X=3.905 $Y=0.505 $X2=0 $Y2=0
cc_358 C N_VGND_c_811_n 0.0133731f $X=5.435 $Y=0.47 $X2=0 $Y2=0
cc_359 N_C_c_382_n N_VGND_c_814_n 0.0360112f $X=3.905 $Y=0.505 $X2=0 $Y2=0
cc_360 C N_VGND_c_814_n 0.0766498f $X=5.435 $Y=0.47 $X2=0 $Y2=0
cc_361 N_C_M1001_g N_VGND_c_815_n 0.0044609f $X=2.495 $Y=0.74 $X2=0 $Y2=0
cc_362 N_C_M1010_g N_VGND_c_815_n 0.0045006f $X=2.925 $Y=0.74 $X2=0 $Y2=0
cc_363 N_C_c_382_n N_VGND_c_815_n 0.0528683f $X=3.905 $Y=0.505 $X2=0 $Y2=0
cc_364 C N_VGND_c_815_n 0.0658172f $X=5.435 $Y=0.47 $X2=0 $Y2=0
cc_365 N_A_27_368#_c_499_n N_VPWR_M1005_d 0.00378122f $X=1.09 $Y=2.425 $X2=-0.19
+ $Y2=1.66
cc_366 N_A_27_368#_c_511_n N_VPWR_M1012_d 0.00378564f $X=6.365 $Y=2.445 $X2=0
+ $Y2=0
cc_367 N_A_27_368#_c_486_n N_VPWR_c_574_n 0.0201449f $X=0.275 $Y=2.815 $X2=0
+ $Y2=0
cc_368 N_A_27_368#_c_499_n N_VPWR_c_574_n 0.0167733f $X=1.09 $Y=2.425 $X2=0
+ $Y2=0
cc_369 N_A_27_368#_c_487_n N_VPWR_c_574_n 0.0201107f $X=1.175 $Y=2.815 $X2=0
+ $Y2=0
cc_370 N_A_27_368#_c_488_n N_VPWR_c_575_n 0.0195957f $X=5.55 $Y=2.835 $X2=0
+ $Y2=0
cc_371 N_A_27_368#_c_511_n N_VPWR_c_575_n 0.0168121f $X=6.365 $Y=2.445 $X2=0
+ $Y2=0
cc_372 N_A_27_368#_c_490_n N_VPWR_c_575_n 0.0188038f $X=6.45 $Y=2.815 $X2=0
+ $Y2=0
cc_373 N_A_27_368#_c_486_n N_VPWR_c_576_n 0.011066f $X=0.275 $Y=2.815 $X2=0
+ $Y2=0
cc_374 N_A_27_368#_c_487_n N_VPWR_c_577_n 0.0109757f $X=1.175 $Y=2.815 $X2=0
+ $Y2=0
cc_375 N_A_27_368#_c_504_n N_VPWR_c_577_n 0.0028011f $X=4.485 $Y=2.595 $X2=0
+ $Y2=0
cc_376 N_A_27_368#_c_488_n N_VPWR_c_577_n 0.00811275f $X=5.55 $Y=2.835 $X2=0
+ $Y2=0
cc_377 N_A_27_368#_c_490_n N_VPWR_c_578_n 0.011066f $X=6.45 $Y=2.815 $X2=0 $Y2=0
cc_378 N_A_27_368#_c_486_n N_VPWR_c_573_n 0.00915947f $X=0.275 $Y=2.815 $X2=0
+ $Y2=0
cc_379 N_A_27_368#_c_499_n N_VPWR_c_573_n 0.0131813f $X=1.09 $Y=2.425 $X2=0
+ $Y2=0
cc_380 N_A_27_368#_c_487_n N_VPWR_c_573_n 0.00907307f $X=1.175 $Y=2.815 $X2=0
+ $Y2=0
cc_381 N_A_27_368#_c_504_n N_VPWR_c_573_n 0.010442f $X=4.485 $Y=2.595 $X2=0
+ $Y2=0
cc_382 N_A_27_368#_c_509_n N_VPWR_c_573_n 0.00720248f $X=5.465 $Y=2.445 $X2=0
+ $Y2=0
cc_383 N_A_27_368#_c_488_n N_VPWR_c_573_n 0.006266f $X=5.55 $Y=2.835 $X2=0 $Y2=0
cc_384 N_A_27_368#_c_511_n N_VPWR_c_573_n 0.0134397f $X=6.365 $Y=2.445 $X2=0
+ $Y2=0
cc_385 N_A_27_368#_c_490_n N_VPWR_c_573_n 0.00915947f $X=6.45 $Y=2.815 $X2=0
+ $Y2=0
cc_386 N_A_27_368#_c_504_n N_A_295_368#_M1003_s 0.00843301f $X=4.485 $Y=2.595
+ $X2=-0.19 $Y2=1.66
cc_387 N_A_27_368#_c_504_n N_A_295_368#_M1002_d 0.00817018f $X=4.485 $Y=2.595
+ $X2=0 $Y2=0
cc_388 N_A_27_368#_c_504_n N_A_295_368#_M1009_d 0.00916087f $X=4.485 $Y=2.595
+ $X2=0 $Y2=0
cc_389 N_A_27_368#_c_509_n N_A_295_368#_M1015_s 0.00392599f $X=5.465 $Y=2.445
+ $X2=0 $Y2=0
cc_390 N_A_27_368#_c_487_n N_A_295_368#_c_642_n 0.00925377f $X=1.175 $Y=2.815
+ $X2=0 $Y2=0
cc_391 N_A_27_368#_c_504_n N_A_295_368#_c_642_n 0.158778f $X=4.485 $Y=2.595
+ $X2=0 $Y2=0
cc_392 N_A_27_368#_M1014_d N_A_295_368#_c_643_n 0.00200562f $X=4.5 $Y=1.84 $X2=0
+ $Y2=0
cc_393 N_A_27_368#_c_504_n N_A_295_368#_c_643_n 0.00708332f $X=4.485 $Y=2.595
+ $X2=0 $Y2=0
cc_394 N_A_27_368#_c_509_n N_A_295_368#_c_643_n 0.0044524f $X=5.465 $Y=2.445
+ $X2=0 $Y2=0
cc_395 N_A_27_368#_c_520_n N_A_295_368#_c_643_n 0.0137977f $X=4.61 $Y=2.445
+ $X2=0 $Y2=0
cc_396 N_A_27_368#_c_509_n N_A_295_368#_c_644_n 0.0159412f $X=5.465 $Y=2.445
+ $X2=0 $Y2=0
cc_397 N_A_27_368#_c_488_n N_A_295_368#_c_644_n 0.0195957f $X=5.55 $Y=2.835
+ $X2=0 $Y2=0
cc_398 N_A_27_368#_c_520_n N_A_295_368#_c_644_n 0.00234679f $X=4.61 $Y=2.445
+ $X2=0 $Y2=0
cc_399 N_A_27_368#_c_504_n N_Y_M1000_s 0.00780516f $X=4.485 $Y=2.595 $X2=0 $Y2=0
cc_400 N_A_27_368#_c_504_n N_Y_M1008_s 0.00783597f $X=4.485 $Y=2.595 $X2=0 $Y2=0
cc_401 N_A_27_368#_M1014_d N_Y_c_696_n 0.00197138f $X=4.5 $Y=1.84 $X2=0 $Y2=0
cc_402 N_VPWR_c_574_n N_A_295_368#_c_642_n 0.00283585f $X=0.725 $Y=2.79 $X2=0
+ $Y2=0
cc_403 N_VPWR_c_577_n N_A_295_368#_c_642_n 0.218565f $X=5.835 $Y=3.33 $X2=0
+ $Y2=0
cc_404 N_VPWR_c_573_n N_A_295_368#_c_642_n 0.124232f $X=6.48 $Y=3.33 $X2=0 $Y2=0
cc_405 N_VPWR_c_575_n N_A_295_368#_c_644_n 0.00207751f $X=6 $Y=2.8 $X2=0 $Y2=0
cc_406 N_VPWR_c_577_n N_A_295_368#_c_644_n 0.0224058f $X=5.835 $Y=3.33 $X2=0
+ $Y2=0
cc_407 N_VPWR_c_573_n N_A_295_368#_c_644_n 0.0124346f $X=6.48 $Y=3.33 $X2=0
+ $Y2=0
cc_408 N_A_295_368#_c_642_n N_Y_M1000_s 0.00412228f $X=4.173 $Y=2.962 $X2=0
+ $Y2=0
cc_409 N_A_295_368#_c_642_n N_Y_M1008_s 0.00415452f $X=4.173 $Y=2.962 $X2=0
+ $Y2=0
cc_410 N_A_295_368#_M1009_d N_Y_c_696_n 0.00370936f $X=3.89 $Y=1.84 $X2=0 $Y2=0
cc_411 N_A_295_368#_M1015_s N_Y_c_696_n 0.00199675f $X=4.95 $Y=1.84 $X2=0 $Y2=0
cc_412 N_A_295_368#_M1002_d N_Y_c_697_n 0.00443682f $X=2.68 $Y=1.84 $X2=0 $Y2=0
cc_413 N_Y_c_688_n N_VGND_M1016_d 0.00342052f $X=1.545 $Y=1.095 $X2=0 $Y2=0
cc_414 N_Y_c_727_n N_VGND_M1011_s 0.00669573f $X=2.545 $Y=0.925 $X2=0 $Y2=0
cc_415 N_Y_c_692_n N_VGND_M1010_s 0.0147644f $X=5.135 $Y=0.925 $X2=0 $Y2=0
cc_416 N_Y_c_689_n N_VGND_c_807_n 0.00555794f $X=0.875 $Y=1.095 $X2=0 $Y2=0
cc_417 Y N_VGND_c_807_n 0.0243474f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_418 N_Y_c_688_n N_VGND_c_808_n 0.0240821f $X=1.545 $Y=1.095 $X2=0 $Y2=0
cc_419 N_Y_c_690_n N_VGND_c_808_n 0.0191389f $X=1.71 $Y=0.515 $X2=0 $Y2=0
cc_420 Y N_VGND_c_808_n 0.0191765f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_421 N_Y_c_690_n N_VGND_c_809_n 0.0127977f $X=1.71 $Y=0.515 $X2=0 $Y2=0
cc_422 N_Y_c_727_n N_VGND_c_809_n 0.0243503f $X=2.545 $Y=0.925 $X2=0 $Y2=0
cc_423 N_Y_c_691_n N_VGND_c_809_n 0.0127977f $X=2.71 $Y=0.515 $X2=0 $Y2=0
cc_424 N_Y_c_691_n N_VGND_c_810_n 0.0144609f $X=2.71 $Y=0.515 $X2=0 $Y2=0
cc_425 N_Y_c_691_n N_VGND_c_811_n 0.0122213f $X=2.71 $Y=0.515 $X2=0 $Y2=0
cc_426 N_Y_c_692_n N_VGND_c_811_n 0.0244298f $X=5.135 $Y=0.925 $X2=0 $Y2=0
cc_427 Y N_VGND_c_812_n 0.0145221f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_428 N_Y_c_690_n N_VGND_c_813_n 0.0144922f $X=1.71 $Y=0.515 $X2=0 $Y2=0
cc_429 N_Y_c_690_n N_VGND_c_815_n 0.0118826f $X=1.71 $Y=0.515 $X2=0 $Y2=0
cc_430 N_Y_c_727_n N_VGND_c_815_n 0.0110662f $X=2.545 $Y=0.925 $X2=0 $Y2=0
cc_431 N_Y_c_691_n N_VGND_c_815_n 0.0118703f $X=2.71 $Y=0.515 $X2=0 $Y2=0
cc_432 N_Y_c_692_n N_VGND_c_815_n 0.0226485f $X=5.135 $Y=0.925 $X2=0 $Y2=0
cc_433 Y N_VGND_c_815_n 0.0119308f $X=0.635 $Y=0.47 $X2=0 $Y2=0
