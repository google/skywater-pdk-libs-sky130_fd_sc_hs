* File: sky130_fd_sc_hs__fah_2.spice
* Created: Tue Sep  1 20:05:45 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hs__fah_2.pex.spice"
.subckt sky130_fd_sc_hs__fah_2  VNB VPB A B CI VPWR COUT SUM VGND
* 
* VGND	VGND
* SUM	SUM
* COUT	COUT
* VPWR	VPWR
* CI	CI
* B	B
* A	A
* VPB	VPB
* VNB	VNB
MM1034 N_A_114_368#_M1034_d N_A_81_260#_M1034_g N_VGND_M1034_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1961 AS=0.222 PD=2.01 PS=2.08 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1017 N_VGND_M1017_d N_A_M1017_g N_A_81_260#_M1017_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.0896 AS=0.2272 PD=0.92 PS=1.99 NRD=0 NRS=13.116 M=1 R=4.26667 SA=75000.3
+ SB=75003.8 A=0.096 P=1.58 MULT=1
MM1005 N_A_413_392#_M1005_d N_A_M1005_g N_VGND_M1017_d VNB NLOWVT L=0.15 W=0.64
+ AD=0.0896 AS=0.0896 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667 SA=75000.7
+ SB=75003.3 A=0.096 P=1.58 MULT=1
MM1006 N_A_514_424#_M1006_d N_B_M1006_g N_A_413_392#_M1005_d VNB NLOWVT L=0.15
+ W=0.64 AD=0.1952 AS=0.0896 PD=1.25 PS=0.92 NRD=61.872 NRS=0 M=1 R=4.26667
+ SA=75001.1 SB=75002.9 A=0.096 P=1.58 MULT=1
MM1008 N_A_114_368#_M1008_d N_A_481_379#_M1008_g N_A_514_424#_M1006_d VNB NLOWVT
+ L=0.15 W=0.64 AD=0.272 AS=0.1952 PD=1.49 PS=1.25 NRD=76.872 NRS=0 M=1
+ R=4.26667 SA=75001.9 SB=75002.2 A=0.096 P=1.58 MULT=1
MM1007 N_A_849_424#_M1007_d N_B_M1007_g N_A_114_368#_M1008_d VNB NLOWVT L=0.15
+ W=0.64 AD=0.2224 AS=0.272 PD=1.335 PS=1.49 NRD=50.616 NRS=29.988 M=1 R=4.26667
+ SA=75002.9 SB=75001.2 A=0.096 P=1.58 MULT=1
MM1025 N_A_413_392#_M1025_d N_A_481_379#_M1025_g N_A_849_424#_M1007_d VNB NLOWVT
+ L=0.15 W=0.64 AD=0.2455 AS=0.2224 PD=2.38 PS=1.335 NRD=49.68 NRS=27.18 M=1
+ R=4.26667 SA=75003.7 SB=75000.3 A=0.096 P=1.58 MULT=1
MM1033 N_A_481_379#_M1033_d N_B_M1033_g N_VGND_M1033_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.124942 AS=0.31405 PD=1.14217 PS=2.87 NRD=0 NRS=66.48 M=1 R=4.93333
+ SA=75000.3 SB=75004 A=0.111 P=1.78 MULT=1
MM1019 N_A_1451_424#_M1019_d N_A_849_424#_M1019_g N_A_481_379#_M1033_d VNB
+ NLOWVT L=0.15 W=0.64 AD=0.28 AS=0.108058 PD=1.515 PS=0.987826 NRD=88.116
+ NRS=8.436 M=1 R=4.26667 SA=75000.8 SB=75004.1 A=0.096 P=1.58 MULT=1
MM1020 N_A_1689_424#_M1020_d N_A_514_424#_M1020_g N_A_1451_424#_M1019_d VNB
+ NLOWVT L=0.15 W=0.64 AD=0.2176 AS=0.28 PD=1.32 PS=1.515 NRD=13.116 NRS=23.436
+ M=1 R=4.26667 SA=75001.9 SB=75003.1 A=0.096 P=1.58 MULT=1
MM1009 N_A_1895_424#_M1009_d N_A_849_424#_M1009_g N_A_1689_424#_M1020_d VNB
+ NLOWVT L=0.15 W=0.64 AD=0.23645 AS=0.2176 PD=1.45 PS=1.32 NRD=15.936
+ NRS=61.872 M=1 R=4.26667 SA=75002.7 SB=75002.2 A=0.096 P=1.58 MULT=1
MM1027 N_A_2052_424#_M1027_d N_A_514_424#_M1027_g N_A_1895_424#_M1009_d VNB
+ NLOWVT L=0.15 W=0.64 AD=0.1344 AS=0.23645 PD=1.06 PS=1.45 NRD=1.872 NRS=60.936
+ M=1 R=4.26667 SA=75003.5 SB=75001.4 A=0.096 P=1.58 MULT=1
MM1011 N_VGND_M1011_d N_A_1689_424#_M1011_g N_A_2052_424#_M1027_d VNB NLOWVT
+ L=0.15 W=0.64 AD=0.1826 AS=0.1344 PD=1.32 PS=1.06 NRD=43.176 NRS=7.02 M=1
+ R=4.26667 SA=75004.1 SB=75000.8 A=0.096 P=1.58 MULT=1
MM1021 N_A_1689_424#_M1021_d N_CI_M1021_g N_VGND_M1011_d VNB NLOWVT L=0.15
+ W=0.64 AD=0.176 AS=0.1826 PD=1.83 PS=1.32 NRD=0 NRS=43.176 M=1 R=4.26667
+ SA=75004.7 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1014 N_COUT_M1014_d N_A_1451_424#_M1014_g N_VGND_M1014_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.2739 PD=1.02 PS=2.27 NRD=0 NRS=12.972 M=1 R=4.93333
+ SA=75000.3 SB=75001.6 A=0.111 P=1.78 MULT=1
MM1035 N_COUT_M1014_d N_A_1451_424#_M1035_g N_VGND_M1035_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.1295 PD=1.02 PS=1.09 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.7 SB=75001.1 A=0.111 P=1.78 MULT=1
MM1022 N_VGND_M1035_s N_A_1895_424#_M1022_g N_SUM_M1022_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1295 AS=0.1073 PD=1.09 PS=1.03 NRD=11.34 NRS=0.804 M=1 R=4.93333
+ SA=75001.2 SB=75000.6 A=0.111 P=1.78 MULT=1
MM1029 N_VGND_M1029_d N_A_1895_424#_M1029_g N_SUM_M1022_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.2109 AS=0.1073 PD=2.05 PS=1.03 NRD=0 NRS=0.804 M=1 R=4.93333
+ SA=75001.6 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1002 N_A_114_368#_M1002_d N_A_81_260#_M1002_g N_VPWR_M1002_s VPB PSHORT L=0.15
+ W=1.12 AD=0.3136 AS=0.3192 PD=2.8 PS=2.81 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75000.2 A=0.168 P=2.54 MULT=1
MM1015 N_VPWR_M1015_d N_A_M1015_g N_A_81_260#_M1015_s VPB PSHORT L=0.15 W=1
+ AD=0.18 AS=0.285 PD=1.36 PS=2.57 NRD=1.9503 NRS=1.9503 M=1 R=6.66667
+ SA=75000.2 SB=75003.8 A=0.15 P=2.3 MULT=1
MM1030 N_A_413_392#_M1030_d N_A_M1030_g N_VPWR_M1015_d VPB PSHORT L=0.15 W=1
+ AD=0.185109 AS=0.18 PD=1.47283 PS=1.36 NRD=2.9353 NRS=13.7703 M=1 R=6.66667
+ SA=75000.7 SB=75003.3 A=0.15 P=2.3 MULT=1
MM1003 N_A_514_424#_M1003_d N_A_481_379#_M1003_g N_A_413_392#_M1030_d VPB PSHORT
+ L=0.15 W=0.84 AD=0.3843 AS=0.155491 PD=1.755 PS=1.23717 NRD=2.3443 NRS=14.0658
+ M=1 R=5.6 SA=75001.2 SB=75003.4 A=0.126 P=1.98 MULT=1
MM1010 N_A_114_368#_M1010_d N_B_M1010_g N_A_514_424#_M1003_d VPB PSHORT L=0.15
+ W=0.84 AD=0.1932 AS=0.3843 PD=1.3 PS=1.755 NRD=21.0987 NRS=14.0658 M=1 R=5.6
+ SA=75002.3 SB=75002.3 A=0.126 P=1.98 MULT=1
MM1016 N_A_849_424#_M1016_d N_A_481_379#_M1016_g N_A_114_368#_M1010_d VPB PSHORT
+ L=0.15 W=0.84 AD=0.5649 AS=0.1932 PD=2.185 PS=1.3 NRD=14.0658 NRS=21.0987 M=1
+ R=5.6 SA=75002.9 SB=75001.7 A=0.126 P=1.98 MULT=1
MM1024 N_A_413_392#_M1024_d N_B_M1024_g N_A_849_424#_M1016_d VPB PSHORT L=0.15
+ W=0.84 AD=0.2394 AS=0.5649 PD=2.25 PS=2.185 NRD=2.3443 NRS=93.7917 M=1 R=5.6
+ SA=75004.4 SB=75000.2 A=0.126 P=1.98 MULT=1
MM1000 N_A_481_379#_M1000_d N_B_M1000_g N_VPWR_M1000_s VPB PSHORT L=0.15 W=1.12
+ AD=0.2256 AS=0.3192 PD=1.70857 PS=2.81 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75003.9 A=0.168 P=2.54 MULT=1
MM1012 N_A_1451_424#_M1012_d N_A_514_424#_M1012_g N_A_481_379#_M1000_d VPB
+ PSHORT L=0.15 W=0.84 AD=0.4368 AS=0.1692 PD=1.88 PS=1.28143 NRD=76.2193
+ NRS=34.3371 M=1 R=5.6 SA=75000.7 SB=75004.6 A=0.126 P=1.98 MULT=1
MM1004 N_A_1689_424#_M1004_d N_A_849_424#_M1004_g N_A_1451_424#_M1012_d VPB
+ PSHORT L=0.15 W=0.84 AD=0.3696 AS=0.4368 PD=1.72 PS=1.88 NRD=113.728
+ NRS=2.3443 M=1 R=5.6 SA=75001.9 SB=75003.4 A=0.126 P=1.98 MULT=1
MM1031 N_A_1895_424#_M1031_d N_A_514_424#_M1031_g N_A_1689_424#_M1004_d VPB
+ PSHORT L=0.15 W=0.84 AD=0.2667 AS=0.3696 PD=1.475 PS=1.72 NRD=69.1667
+ NRS=26.9693 M=1 R=5.6 SA=75003 SB=75002.3 A=0.126 P=1.98 MULT=1
MM1013 N_A_2052_424#_M1013_d N_A_849_424#_M1013_g N_A_1895_424#_M1031_d VPB
+ PSHORT L=0.15 W=0.84 AD=0.224517 AS=0.2667 PD=1.40152 PS=1.475 NRD=22.261
+ NRS=14.0658 M=1 R=5.6 SA=75003.7 SB=75001.6 A=0.126 P=1.98 MULT=1
MM1032 N_VPWR_M1032_d N_A_1689_424#_M1032_g N_A_2052_424#_M1013_d VPB PSHORT
+ L=0.15 W=1 AD=0.2957 AS=0.267283 PD=1.73 PS=1.66848 NRD=47.3982 NRS=10.3228
+ M=1 R=6.66667 SA=75003.7 SB=75000.9 A=0.15 P=2.3 MULT=1
MM1001 N_A_1689_424#_M1001_d N_CI_M1001_g N_VPWR_M1032_d VPB PSHORT L=0.15 W=1
+ AD=0.285 AS=0.2957 PD=2.57 PS=1.73 NRD=0 NRS=47.3982 M=1 R=6.66667 SA=75004.4
+ SB=75000.2 A=0.15 P=2.3 MULT=1
MM1023 N_COUT_M1023_d N_A_1451_424#_M1023_g N_VPWR_M1023_s VPB PSHORT L=0.15
+ W=1.12 AD=0.168 AS=0.303 PD=1.42 PS=2.81 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75001.6 A=0.168 P=2.54 MULT=1
MM1026 N_COUT_M1023_d N_A_1451_424#_M1026_g N_VPWR_M1026_s VPB PSHORT L=0.15
+ W=1.12 AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.6 SB=75001.1 A=0.168 P=2.54 MULT=1
MM1018 N_VPWR_M1026_s N_A_1895_424#_M1018_g N_SUM_M1018_s VPB PSHORT L=0.15
+ W=1.12 AD=0.168 AS=0.1736 PD=1.42 PS=1.43 NRD=1.7533 NRS=2.6201 M=1 R=7.46667
+ SA=75001.1 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1028 N_VPWR_M1028_d N_A_1895_424#_M1028_g N_SUM_M1018_s VPB PSHORT L=0.15
+ W=1.12 AD=0.336 AS=0.1736 PD=2.84 PS=1.43 NRD=4.3931 NRS=2.6201 M=1 R=7.46667
+ SA=75001.6 SB=75000.2 A=0.168 P=2.54 MULT=1
DX36_noxref VNB VPB NWDIODE A=27.4908 P=33.28
c_147 VNB 0 7.1893e-20 $X=0 $Y=0
c_257 VPB 0 5.31033e-20 $X=0 $Y=3.085
*
.include "sky130_fd_sc_hs__fah_2.pxi.spice"
*
.ends
*
*
