* File: sky130_fd_sc_hs__dfrtp_2.pex.spice
* Created: Thu Aug 27 20:38:45 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HS__DFRTP_2%D 2 4 5 7 10 12 13 14 19 20 23
r34 23 25 40.9207 $w=3.65e-07 $l=1.65e-07 $layer=POLY_cond $X=0.402 $Y=1.845
+ $X2=0.402 $Y2=2.01
r35 23 24 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=0.385
+ $Y=1.845 $X2=0.385 $Y2=1.845
r36 19 21 46.6671 $w=3.65e-07 $l=1.65e-07 $layer=POLY_cond $X=0.402 $Y=1.165
+ $X2=0.402 $Y2=1
r37 19 20 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=0.385
+ $Y=1.165 $X2=0.385 $Y2=1.165
r38 14 24 5.91795 $w=3.68e-07 $l=1.9e-07 $layer=LI1_cond $X=0.31 $Y=2.035
+ $X2=0.31 $Y2=1.845
r39 13 24 5.60648 $w=3.68e-07 $l=1.8e-07 $layer=LI1_cond $X=0.31 $Y=1.665
+ $X2=0.31 $Y2=1.845
r40 12 13 11.5244 $w=3.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.31 $Y=1.295
+ $X2=0.31 $Y2=1.665
r41 12 20 4.04912 $w=3.68e-07 $l=1.3e-07 $layer=LI1_cond $X=0.31 $Y=1.295
+ $X2=0.31 $Y2=1.165
r42 10 21 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=0.51 $Y=0.6 $X2=0.51
+ $Y2=1
r43 5 7 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=0.495 $Y=2.465
+ $X2=0.495 $Y2=2.75
r44 4 5 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=0.495 $Y=2.375 $X2=0.495
+ $Y2=2.465
r45 4 25 141.879 $w=1.8e-07 $l=3.65e-07 $layer=POLY_cond $X=0.495 $Y=2.375
+ $X2=0.495 $Y2=2.01
r46 2 23 2.68759 $w=3.65e-07 $l=1.7e-08 $layer=POLY_cond $X=0.402 $Y=1.828
+ $X2=0.402 $Y2=1.845
r47 1 19 2.68759 $w=3.65e-07 $l=1.7e-08 $layer=POLY_cond $X=0.402 $Y=1.182
+ $X2=0.402 $Y2=1.165
r48 1 2 102.129 $w=3.65e-07 $l=6.46e-07 $layer=POLY_cond $X=0.402 $Y=1.182
+ $X2=0.402 $Y2=1.828
.ends

.subckt PM_SKY130_FD_SC_HS__DFRTP_2%RESET_B 3 6 8 9 11 12 14 16 17 19 20 22 25
+ 29 31 32 33 34 37 39 42 45 46 49 57
c190 46 0 7.91465e-21 $X=1.12 $Y=1.305
c191 45 0 1.04983e-19 $X=1.12 $Y=1.305
c192 39 0 3.83476e-20 $X=7.92 $Y=2.035
c193 33 0 4.38853e-20 $X=7.775 $Y=2.035
c194 29 0 4.03239e-20 $X=4.88 $Y=1.26
r195 56 57 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.23
+ $Y=2.11 $X2=8.23 $Y2=2.11
r196 49 51 41.3282 $w=4.6e-07 $l=1.65e-07 $layer=POLY_cond $X=1.055 $Y=1.985
+ $X2=1.055 $Y2=2.15
r197 49 50 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.12
+ $Y=1.985 $X2=1.12 $Y2=1.985
r198 46 50 27.9879 $w=2.78e-07 $l=6.8e-07 $layer=LI1_cond $X=1.145 $Y=1.305
+ $X2=1.145 $Y2=1.985
r199 45 47 47.2161 $w=4.6e-07 $l=1.65e-07 $layer=POLY_cond $X=1.055 $Y=1.305
+ $X2=1.055 $Y2=1.14
r200 45 46 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.12
+ $Y=1.305 $X2=1.12 $Y2=1.305
r201 42 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=2.035
+ $X2=1.2 $Y2=2.035
r202 40 57 10.0636 $w=3.53e-07 $l=3.1e-07 $layer=LI1_cond $X=7.92 $Y=2.097
+ $X2=8.23 $Y2=2.097
r203 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=2.035
+ $X2=7.92 $Y2=2.035
r204 37 53 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.12
+ $Y=1.96 $X2=5.12 $Y2=1.96
r205 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=2.035
+ $X2=5.04 $Y2=2.035
r206 34 36 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.185 $Y=2.035
+ $X2=5.04 $Y2=2.035
r207 33 39 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=7.775 $Y=2.035
+ $X2=7.92 $Y2=2.035
r208 33 34 3.20544 $w=1.4e-07 $l=2.59e-06 $layer=MET1_cond $X=7.775 $Y=2.035
+ $X2=5.185 $Y2=2.035
r209 32 42 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.345 $Y=2.035
+ $X2=1.2 $Y2=2.035
r210 31 36 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.895 $Y=2.035
+ $X2=5.04 $Y2=2.035
r211 31 32 4.39356 $w=1.4e-07 $l=3.55e-06 $layer=MET1_cond $X=4.895 $Y=2.035
+ $X2=1.345 $Y2=2.035
r212 27 29 46.1489 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=4.79 $Y=1.26 $X2=4.88
+ $Y2=1.26
r213 23 56 38.6072 $w=2.91e-07 $l=1.69926e-07 $layer=POLY_cond $X=8.24 $Y=1.945
+ $X2=8.23 $Y2=2.11
r214 23 25 681.979 $w=1.5e-07 $l=1.33e-06 $layer=POLY_cond $X=8.24 $Y=1.945
+ $X2=8.24 $Y2=0.615
r215 20 56 57.6553 $w=2.91e-07 $l=2.82489e-07 $layer=POLY_cond $X=8.235 $Y=2.39
+ $X2=8.23 $Y2=2.11
r216 20 22 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=8.235 $Y=2.39
+ $X2=8.235 $Y2=2.675
r217 17 53 49.7565 $w=4.18e-07 $l=3.16228e-07 $layer=POLY_cond $X=4.895 $Y=2.21
+ $X2=5.045 $Y2=1.96
r218 17 19 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=4.895 $Y=2.21
+ $X2=4.895 $Y2=2.495
r219 16 53 39.9551 $w=4.18e-07 $l=2.33345e-07 $layer=POLY_cond $X=4.88 $Y=1.795
+ $X2=5.045 $Y2=1.96
r220 15 29 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.88 $Y=1.335
+ $X2=4.88 $Y2=1.26
r221 15 16 235.872 $w=1.5e-07 $l=4.6e-07 $layer=POLY_cond $X=4.88 $Y=1.335
+ $X2=4.88 $Y2=1.795
r222 12 27 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.79 $Y=1.185
+ $X2=4.79 $Y2=1.26
r223 12 14 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=4.79 $Y=1.185
+ $X2=4.79 $Y2=0.9
r224 9 11 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=0.945 $Y=2.465
+ $X2=0.945 $Y2=2.75
r225 8 9 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=0.945 $Y=2.375
+ $X2=0.945 $Y2=2.465
r226 8 51 87.4597 $w=1.8e-07 $l=2.25e-07 $layer=POLY_cond $X=0.945 $Y=2.375
+ $X2=0.945 $Y2=2.15
r227 6 49 7.8587 $w=4.6e-07 $l=6.5e-08 $layer=POLY_cond $X=1.055 $Y=1.92
+ $X2=1.055 $Y2=1.985
r228 5 45 7.8587 $w=4.6e-07 $l=6.5e-08 $layer=POLY_cond $X=1.055 $Y=1.37
+ $X2=1.055 $Y2=1.305
r229 5 6 66.4967 $w=4.6e-07 $l=5.5e-07 $layer=POLY_cond $X=1.055 $Y=1.37
+ $X2=1.055 $Y2=1.92
r230 3 47 276.894 $w=1.5e-07 $l=5.4e-07 $layer=POLY_cond $X=0.9 $Y=0.6 $X2=0.9
+ $Y2=1.14
.ends

.subckt PM_SKY130_FD_SC_HS__DFRTP_2%CLK 3 5 7 8
c43 5 0 1.57874e-19 $X=1.925 $Y=1.735
c44 3 0 7.91465e-21 $X=1.89 $Y=0.74
r45 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.91
+ $Y=1.485 $X2=1.91 $Y2=1.485
r46 8 12 7.78061 $w=3.92e-07 $l=2.5e-07 $layer=LI1_cond $X=2.16 $Y=1.55 $X2=1.91
+ $Y2=1.55
r47 5 11 52.2586 $w=2.99e-07 $l=2.57391e-07 $layer=POLY_cond $X=1.925 $Y=1.735
+ $X2=1.91 $Y2=1.485
r48 5 7 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.925 $Y=1.735
+ $X2=1.925 $Y2=2.37
r49 1 11 38.5562 $w=2.99e-07 $l=1.74714e-07 $layer=POLY_cond $X=1.89 $Y=1.32
+ $X2=1.91 $Y2=1.485
r50 1 3 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=1.89 $Y=1.32 $X2=1.89
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HS__DFRTP_2%A_490_362# 1 2 8 9 11 12 14 16 18 20 21 22
+ 23 25 28 29 31 33 36 39 40 41 44 45 48 49 57 63 66 68
c193 44 0 1.33493e-19 $X=7.12 $Y=2.14
c194 22 0 4.38853e-20 $X=6.355 $Y=1.27
c195 16 0 8.97095e-20 $X=4.01 $Y=0.9
r196 65 66 8.73063 $w=3.28e-07 $l=2.5e-07 $layer=LI1_cond $X=7.12 $Y=1.18
+ $X2=7.37 $Y2=1.18
r197 63 74 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=6.88 $Y=1.18 $X2=6.88
+ $Y2=1.27
r198 62 65 8.3814 $w=3.28e-07 $l=2.4e-07 $layer=LI1_cond $X=6.88 $Y=1.18
+ $X2=7.12 $Y2=1.18
r199 62 63 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.88
+ $Y=1.18 $X2=6.88 $Y2=1.18
r200 57 59 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=4.355 $Y=0.415
+ $X2=4.355 $Y2=0.7
r201 55 56 11.8011 $w=3.67e-07 $l=3.55e-07 $layer=LI1_cond $X=2.6 $Y=1.847
+ $X2=2.955 $Y2=1.847
r202 52 53 10.2686 $w=5.28e-07 $l=1.9e-07 $layer=LI1_cond $X=2.775 $Y=0.62
+ $X2=2.775 $Y2=0.81
r203 49 52 4.62634 $w=5.28e-07 $l=2.05e-07 $layer=LI1_cond $X=2.775 $Y=0.415
+ $X2=2.775 $Y2=0.62
r204 48 66 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.37 $Y=1.015
+ $X2=7.37 $Y2=1.18
r205 47 48 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=7.37 $Y=0.425
+ $X2=7.37 $Y2=1.015
r206 45 77 25.8214 $w=3.64e-07 $l=1.95e-07 $layer=POLY_cond $X=7.12 $Y=2.182
+ $X2=7.315 $Y2=2.182
r207 44 45 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.12
+ $Y=2.14 $X2=7.12 $Y2=2.14
r208 42 65 0.716491 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=7.12 $Y=1.345
+ $X2=7.12 $Y2=1.18
r209 42 44 27.7634 $w=3.28e-07 $l=7.95e-07 $layer=LI1_cond $X=7.12 $Y=1.345
+ $X2=7.12 $Y2=2.14
r210 40 47 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.285 $Y=0.34
+ $X2=7.37 $Y2=0.425
r211 40 41 104.385 $w=1.68e-07 $l=1.6e-06 $layer=LI1_cond $X=7.285 $Y=0.34
+ $X2=5.685 $Y2=0.34
r212 38 41 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.6 $Y=0.425
+ $X2=5.685 $Y2=0.34
r213 38 39 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=5.6 $Y=0.425
+ $X2=5.6 $Y2=0.615
r214 37 59 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.44 $Y=0.7
+ $X2=4.355 $Y2=0.7
r215 36 39 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.515 $Y=0.7
+ $X2=5.6 $Y2=0.615
r216 36 37 70.1337 $w=1.68e-07 $l=1.075e-06 $layer=LI1_cond $X=5.515 $Y=0.7
+ $X2=4.44 $Y2=0.7
r217 34 71 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.33 $Y=1.74
+ $X2=3.33 $Y2=1.905
r218 34 68 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=3.33 $Y=1.74 $X2=3.33
+ $Y2=1.65
r219 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.33
+ $Y=1.74 $X2=3.33 $Y2=1.74
r220 31 56 2.97641 $w=3.67e-07 $l=1.43332e-07 $layer=LI1_cond $X=3.04 $Y=1.74
+ $X2=2.955 $Y2=1.847
r221 31 33 10.1275 $w=3.28e-07 $l=2.9e-07 $layer=LI1_cond $X=3.04 $Y=1.74
+ $X2=3.33 $Y2=1.74
r222 30 49 7.52407 $w=1.7e-07 $l=2.65e-07 $layer=LI1_cond $X=3.04 $Y=0.415
+ $X2=2.775 $Y2=0.415
r223 29 57 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.27 $Y=0.415
+ $X2=4.355 $Y2=0.415
r224 29 30 80.246 $w=1.68e-07 $l=1.23e-06 $layer=LI1_cond $X=4.27 $Y=0.415
+ $X2=3.04 $Y2=0.415
r225 28 56 5.25812 $w=1.7e-07 $l=2.72e-07 $layer=LI1_cond $X=2.955 $Y=1.575
+ $X2=2.955 $Y2=1.847
r226 28 53 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=2.955 $Y=1.575
+ $X2=2.955 $Y2=0.81
r227 23 77 23.572 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=7.315 $Y=2.39
+ $X2=7.315 $Y2=2.182
r228 23 25 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=7.315 $Y=2.39
+ $X2=7.315 $Y2=2.675
r229 21 74 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.715 $Y=1.27
+ $X2=6.88 $Y2=1.27
r230 21 22 184.596 $w=1.5e-07 $l=3.6e-07 $layer=POLY_cond $X=6.715 $Y=1.27
+ $X2=6.355 $Y2=1.27
r231 18 22 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=6.28 $Y=1.195
+ $X2=6.355 $Y2=1.27
r232 18 20 146.207 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=6.28 $Y=1.195
+ $X2=6.28 $Y2=0.74
r233 14 26 61.9591 $w=2.01e-07 $l=2.71109e-07 $layer=POLY_cond $X=4.01 $Y=1.405
+ $X2=3.955 $Y2=1.65
r234 14 16 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=4.01 $Y=1.405
+ $X2=4.01 $Y2=0.9
r235 13 68 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.495 $Y=1.65
+ $X2=3.33 $Y2=1.65
r236 12 26 9.69179 $w=1.5e-07 $l=1.3e-07 $layer=POLY_cond $X=3.825 $Y=1.65
+ $X2=3.955 $Y2=1.65
r237 12 13 169.213 $w=1.5e-07 $l=3.3e-07 $layer=POLY_cond $X=3.825 $Y=1.65
+ $X2=3.495 $Y2=1.65
r238 9 11 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=3.405 $Y=2.21
+ $X2=3.405 $Y2=2.495
r239 8 9 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=3.405 $Y=2.12 $X2=3.405
+ $Y2=2.21
r240 8 71 83.5726 $w=1.8e-07 $l=2.15e-07 $layer=POLY_cond $X=3.405 $Y=2.12
+ $X2=3.405 $Y2=1.905
r241 2 55 600 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=2.45
+ $Y=1.81 $X2=2.6 $Y2=1.955
r242 1 52 182 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=1 $X=2.535
+ $Y=0.37 $X2=2.675 $Y2=0.62
.ends

.subckt PM_SKY130_FD_SC_HS__DFRTP_2%A_837_359# 1 2 7 9 12 16 19 20 23 29 31 32
c82 20 0 1.7626e-19 $X=4.445 $Y=1.04
c83 16 0 4.03239e-20 $X=4.36 $Y=1.96
c84 12 0 1.23255e-19 $X=4.4 $Y=0.9
r85 29 32 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=6.18 $Y=2.02
+ $X2=6.18 $Y2=1.855
r86 25 31 3.70735 $w=2.5e-07 $l=1.21589e-07 $layer=LI1_cond $X=6.1 $Y=1.13
+ $X2=6.02 $Y2=1.042
r87 25 32 47.2995 $w=1.68e-07 $l=7.25e-07 $layer=LI1_cond $X=6.1 $Y=1.13 $X2=6.1
+ $Y2=1.855
r88 21 31 3.70735 $w=2.5e-07 $l=8.7e-08 $layer=LI1_cond $X=6.02 $Y=0.955
+ $X2=6.02 $Y2=1.042
r89 21 23 3.31764 $w=3.28e-07 $l=9.5e-08 $layer=LI1_cond $X=6.02 $Y=0.955
+ $X2=6.02 $Y2=0.86
r90 19 31 2.76166 $w=1.7e-07 $l=1.65997e-07 $layer=LI1_cond $X=5.855 $Y=1.04
+ $X2=6.02 $Y2=1.042
r91 19 20 91.9893 $w=1.68e-07 $l=1.41e-06 $layer=LI1_cond $X=5.855 $Y=1.04
+ $X2=4.445 $Y2=1.04
r92 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.36
+ $Y=1.96 $X2=4.36 $Y2=1.96
r93 14 20 6.81835 $w=1.7e-07 $l=1.23386e-07 $layer=LI1_cond $X=4.357 $Y=1.125
+ $X2=4.445 $Y2=1.04
r94 14 16 52.9195 $w=1.73e-07 $l=8.35e-07 $layer=LI1_cond $X=4.357 $Y=1.125
+ $X2=4.357 $Y2=1.96
r95 10 17 38.5336 $w=3.07e-07 $l=1.86145e-07 $layer=POLY_cond $X=4.4 $Y=1.795
+ $X2=4.355 $Y2=1.96
r96 10 12 458.926 $w=1.5e-07 $l=8.95e-07 $layer=POLY_cond $X=4.4 $Y=1.795
+ $X2=4.4 $Y2=0.9
r97 7 17 51.8789 $w=3.07e-07 $l=2.87228e-07 $layer=POLY_cond $X=4.275 $Y=2.21
+ $X2=4.355 $Y2=1.96
r98 7 9 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=4.275 $Y=2.21 $X2=4.275
+ $Y2=2.495
r99 2 29 300 $w=1.7e-07 $l=3.71786e-07 $layer=licon1_PDIFF $count=2 $X=5.98
+ $Y=1.735 $X2=6.18 $Y2=2.02
r100 1 23 182 $w=1.7e-07 $l=5.55608e-07 $layer=licon1_NDIFF $count=1 $X=5.88
+ $Y=0.37 $X2=6.02 $Y2=0.86
.ends

.subckt PM_SKY130_FD_SC_HS__DFRTP_2%A_696_457# 1 2 3 12 14 16 18 20 21 22 24 25
+ 27 32 40 42
c121 40 0 1.23255e-19 $X=4.015 $Y=0.867
c122 25 0 1.21261e-19 $X=4.785 $Y=1.435
c123 22 0 1.12683e-19 $X=4.1 $Y=2.5
r124 38 40 6.41867 $w=3.93e-07 $l=2.2e-07 $layer=LI1_cond $X=3.795 $Y=0.867
+ $X2=4.015 $Y2=0.867
r125 35 36 19.4091 $w=2.42e-07 $l=3.85e-07 $layer=LI1_cond $X=3.63 $Y=2.57
+ $X2=4.015 $Y2=2.57
r126 30 42 4.18896 $w=2.17e-07 $l=8.5e-08 $layer=LI1_cond $X=4.785 $Y=2.452
+ $X2=4.7 $Y2=2.452
r127 30 32 14.5686 $w=2.63e-07 $l=3.35e-07 $layer=LI1_cond $X=4.785 $Y=2.452
+ $X2=5.12 $Y2=2.452
r128 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.52
+ $Y=1.41 $X2=5.52 $Y2=1.41
r129 25 27 30.2516 $w=2.78e-07 $l=7.35e-07 $layer=LI1_cond $X=4.785 $Y=1.435
+ $X2=5.52 $Y2=1.435
r130 24 42 2.24312 $w=1.7e-07 $l=1.32e-07 $layer=LI1_cond $X=4.7 $Y=2.32 $X2=4.7
+ $Y2=2.452
r131 23 25 7.36005 $w=2.8e-07 $l=1.77482e-07 $layer=LI1_cond $X=4.7 $Y=1.575
+ $X2=4.785 $Y2=1.435
r132 23 24 48.6043 $w=1.68e-07 $l=7.45e-07 $layer=LI1_cond $X=4.7 $Y=1.575
+ $X2=4.7 $Y2=2.32
r133 22 36 5.3796 $w=2.42e-07 $l=1.14782e-07 $layer=LI1_cond $X=4.1 $Y=2.5
+ $X2=4.015 $Y2=2.57
r134 21 42 4.18896 $w=2.17e-07 $l=1.06325e-07 $layer=LI1_cond $X=4.615 $Y=2.5
+ $X2=4.7 $Y2=2.452
r135 21 22 33.5989 $w=1.68e-07 $l=5.15e-07 $layer=LI1_cond $X=4.615 $Y=2.5
+ $X2=4.1 $Y2=2.5
r136 20 36 2.80567 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=4.015 $Y=2.415
+ $X2=4.015 $Y2=2.57
r137 19 40 5.70203 $w=1.7e-07 $l=1.98e-07 $layer=LI1_cond $X=4.015 $Y=1.065
+ $X2=4.015 $Y2=0.867
r138 19 20 88.0749 $w=1.68e-07 $l=1.35e-06 $layer=LI1_cond $X=4.015 $Y=1.065
+ $X2=4.015 $Y2=2.415
r139 18 28 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=5.73 $Y=1.41
+ $X2=5.52 $Y2=1.41
r140 14 18 64.0286 $w=1.97e-07 $l=2.70647e-07 $layer=POLY_cond $X=5.905 $Y=1.66
+ $X2=5.862 $Y2=1.41
r141 14 16 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=5.905 $Y=1.66
+ $X2=5.905 $Y2=2.235
r142 10 18 43.2316 $w=1.97e-07 $l=1.9139e-07 $layer=POLY_cond $X=5.805 $Y=1.245
+ $X2=5.862 $Y2=1.41
r143 10 12 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=5.805 $Y=1.245
+ $X2=5.805 $Y2=0.74
r144 3 32 600 $w=1.7e-07 $l=2.69768e-07 $layer=licon1_PDIFF $count=1 $X=4.97
+ $Y=2.285 $X2=5.12 $Y2=2.49
r145 2 35 600 $w=1.7e-07 $l=3.11087e-07 $layer=licon1_PDIFF $count=1 $X=3.48
+ $Y=2.285 $X2=3.63 $Y2=2.53
r146 1 38 182 $w=1.7e-07 $l=2.84341e-07 $layer=licon1_NDIFF $count=1 $X=3.585
+ $Y=0.69 $X2=3.795 $Y2=0.865
.ends

.subckt PM_SKY130_FD_SC_HS__DFRTP_2%A_306_74# 1 2 7 9 10 12 13 16 17 18 19 21 22
+ 23 24 26 27 32 33 34 37 40 41 42 43 47 50 51 55 56 58 62
c182 58 0 1.04983e-19 $X=1.647 $Y=1.065
c183 55 0 1.57874e-19 $X=2.57 $Y=1.385
c184 41 0 5.51194e-20 $X=2.51 $Y=1.575
c185 33 0 3.77492e-20 $X=7.255 $Y=1.66
c186 16 0 1.12683e-19 $X=2.88 $Y=3.075
r187 59 62 5.5876 $w=3.28e-07 $l=1.6e-07 $layer=LI1_cond $X=1.54 $Y=1.985
+ $X2=1.7 $Y2=1.985
r188 55 56 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.57
+ $Y=1.385 $X2=2.57 $Y2=1.385
r189 53 55 10.6206 $w=2.53e-07 $l=2.35e-07 $layer=LI1_cond $X=2.572 $Y=1.15
+ $X2=2.572 $Y2=1.385
r190 52 58 3.15366 $w=1.7e-07 $l=1.93e-07 $layer=LI1_cond $X=1.84 $Y=1.065
+ $X2=1.647 $Y2=1.065
r191 51 53 7.17723 $w=1.7e-07 $l=1.64085e-07 $layer=LI1_cond $X=2.445 $Y=1.065
+ $X2=2.572 $Y2=1.15
r192 51 52 39.4706 $w=1.68e-07 $l=6.05e-07 $layer=LI1_cond $X=2.445 $Y=1.065
+ $X2=1.84 $Y2=1.065
r193 50 59 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.54 $Y=1.82
+ $X2=1.54 $Y2=1.985
r194 49 58 3.37808 $w=2.77e-07 $l=1.43332e-07 $layer=LI1_cond $X=1.54 $Y=1.15
+ $X2=1.647 $Y2=1.065
r195 49 50 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.54 $Y=1.15
+ $X2=1.54 $Y2=1.82
r196 45 58 3.37808 $w=2.77e-07 $l=8.5e-08 $layer=LI1_cond $X=1.647 $Y=0.98
+ $X2=1.647 $Y2=1.065
r197 45 47 13.9191 $w=3.83e-07 $l=4.65e-07 $layer=LI1_cond $X=1.647 $Y=0.98
+ $X2=1.647 $Y2=0.515
r198 41 56 23.4821 $w=4.5e-07 $l=1.9e-07 $layer=POLY_cond $X=2.51 $Y=1.575
+ $X2=2.51 $Y2=1.385
r199 39 56 6.17949 $w=4.5e-07 $l=5e-08 $layer=POLY_cond $X=2.51 $Y=1.335
+ $X2=2.51 $Y2=1.385
r200 39 40 11.1008 $w=3e-07 $l=7.5e-08 $layer=POLY_cond $X=2.51 $Y=1.335
+ $X2=2.51 $Y2=1.26
r201 35 37 497.383 $w=1.5e-07 $l=9.7e-07 $layer=POLY_cond $X=7.33 $Y=1.585
+ $X2=7.33 $Y2=0.615
r202 33 35 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=7.255 $Y=1.66
+ $X2=7.33 $Y2=1.585
r203 33 34 394.83 $w=1.5e-07 $l=7.7e-07 $layer=POLY_cond $X=7.255 $Y=1.66
+ $X2=6.485 $Y2=1.66
r204 30 43 105.158 $w=1.8e-07 $l=2.65e-07 $layer=POLY_cond $X=6.41 $Y=2.885
+ $X2=6.41 $Y2=3.15
r205 30 32 294.84 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=6.41 $Y=2.885
+ $X2=6.41 $Y2=2.31
r206 29 34 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=6.41 $Y=1.735
+ $X2=6.485 $Y2=1.66
r207 29 32 294.84 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=6.41 $Y=1.735
+ $X2=6.41 $Y2=2.31
r208 28 42 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=3.945 $Y=3.15
+ $X2=3.855 $Y2=3.15
r209 27 43 7.1379 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=6.32 $Y=3.15 $X2=6.41
+ $Y2=3.15
r210 27 28 1217.82 $w=1.5e-07 $l=2.375e-06 $layer=POLY_cond $X=6.32 $Y=3.15
+ $X2=3.945 $Y2=3.15
r211 24 26 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=3.855 $Y=2.78
+ $X2=3.855 $Y2=2.495
r212 23 42 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=3.855 $Y=3.075
+ $X2=3.855 $Y2=3.15
r213 22 24 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=3.855 $Y=2.87
+ $X2=3.855 $Y2=2.78
r214 22 23 79.6855 $w=1.8e-07 $l=2.05e-07 $layer=POLY_cond $X=3.855 $Y=2.87
+ $X2=3.855 $Y2=3.075
r215 19 21 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=3.51 $Y=1.185
+ $X2=3.51 $Y2=0.9
r216 17 42 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=3.765 $Y=3.15
+ $X2=3.855 $Y2=3.15
r217 17 18 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=3.765 $Y=3.15
+ $X2=2.955 $Y2=3.15
r218 16 18 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.88 $Y=3.075
+ $X2=2.955 $Y2=3.15
r219 14 40 15.4994 $w=1.5e-07 $l=2.25e-07 $layer=POLY_cond $X=2.735 $Y=1.26
+ $X2=2.51 $Y2=1.26
r220 13 19 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.435 $Y=1.26
+ $X2=3.51 $Y2=1.185
r221 13 14 358.936 $w=1.5e-07 $l=7e-07 $layer=POLY_cond $X=3.435 $Y=1.26
+ $X2=2.735 $Y2=1.26
r222 10 40 11.1008 $w=3e-07 $l=9.68246e-08 $layer=POLY_cond $X=2.46 $Y=1.185
+ $X2=2.51 $Y2=1.26
r223 10 12 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=2.46 $Y=1.185
+ $X2=2.46 $Y2=0.74
r224 7 41 11.3146 $w=6.39e-07 $l=4.38634e-07 $layer=POLY_cond $X=2.88 $Y=1.725
+ $X2=2.51 $Y2=1.575
r225 7 16 692.234 $w=1.5e-07 $l=1.35e-06 $layer=POLY_cond $X=2.88 $Y=1.725
+ $X2=2.88 $Y2=3.075
r226 7 9 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.375 $Y=1.735
+ $X2=2.375 $Y2=2.37
r227 2 62 600 $w=1.7e-07 $l=2.3103e-07 $layer=licon1_PDIFF $count=1 $X=1.57
+ $Y=1.81 $X2=1.7 $Y2=1.985
r228 1 47 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=1.53
+ $Y=0.37 $X2=1.675 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__DFRTP_2%A_1525_212# 1 2 9 13 14 15 17 18 19 21 27 30
+ 31 32 33 36 38 39 43
c118 39 0 1.33493e-19 $X=7.79 $Y=1.225
c119 36 0 4.37308e-20 $X=9.29 $Y=2.105
c120 21 0 4.77539e-20 $X=8.715 $Y=2.61
c121 13 0 3.83476e-20 $X=7.735 $Y=2.065
r122 39 46 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=7.79 $Y=1.225
+ $X2=7.79 $Y2=1.39
r123 39 45 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=7.79 $Y=1.225
+ $X2=7.79 $Y2=1.06
r124 38 41 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=7.79 $Y=1.225 $X2=7.79
+ $Y2=1.305
r125 38 39 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.79
+ $Y=1.225 $X2=7.79 $Y2=1.225
r126 35 36 46.6471 $w=1.68e-07 $l=7.15e-07 $layer=LI1_cond $X=9.29 $Y=1.39
+ $X2=9.29 $Y2=2.105
r127 34 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.01 $Y=1.305
+ $X2=8.845 $Y2=1.305
r128 33 35 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.205 $Y=1.305
+ $X2=9.29 $Y2=1.39
r129 33 34 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=9.205 $Y=1.305
+ $X2=9.01 $Y2=1.305
r130 31 36 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.205 $Y=2.19
+ $X2=9.29 $Y2=2.105
r131 31 32 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=9.205 $Y=2.19
+ $X2=8.885 $Y2=2.19
r132 29 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.8 $Y=2.275
+ $X2=8.885 $Y2=2.19
r133 29 30 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=8.8 $Y=2.275
+ $X2=8.8 $Y2=2.445
r134 25 43 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.845 $Y=1.22
+ $X2=8.845 $Y2=1.305
r135 25 27 21.1281 $w=3.28e-07 $l=6.05e-07 $layer=LI1_cond $X=8.845 $Y=1.22
+ $X2=8.845 $Y2=0.615
r136 21 30 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=8.715 $Y=2.61
+ $X2=8.8 $Y2=2.445
r137 21 23 4.36531 $w=3.28e-07 $l=1.25e-07 $layer=LI1_cond $X=8.715 $Y=2.61
+ $X2=8.59 $Y2=2.61
r138 20 41 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.955 $Y=1.305
+ $X2=7.79 $Y2=1.305
r139 19 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.68 $Y=1.305
+ $X2=8.845 $Y2=1.305
r140 19 20 47.2995 $w=1.68e-07 $l=7.25e-07 $layer=LI1_cond $X=8.68 $Y=1.305
+ $X2=7.955 $Y2=1.305
r141 18 46 299.968 $w=1.5e-07 $l=5.85e-07 $layer=POLY_cond $X=7.72 $Y=1.975
+ $X2=7.72 $Y2=1.39
r142 15 17 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=7.735 $Y=2.39
+ $X2=7.735 $Y2=2.675
r143 14 15 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=7.735 $Y=2.3
+ $X2=7.735 $Y2=2.39
r144 13 18 37.1337 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=7.735 $Y=2.065
+ $X2=7.735 $Y2=1.975
r145 13 14 91.3468 $w=1.8e-07 $l=2.35e-07 $layer=POLY_cond $X=7.735 $Y=2.065
+ $X2=7.735 $Y2=2.3
r146 9 45 228.181 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=7.72 $Y=0.615
+ $X2=7.72 $Y2=1.06
r147 2 23 600 $w=1.7e-07 $l=3.44964e-07 $layer=licon1_PDIFF $count=1 $X=8.31
+ $Y=2.465 $X2=8.59 $Y2=2.61
r148 1 27 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=8.705
+ $Y=0.405 $X2=8.845 $Y2=0.615
.ends

.subckt PM_SKY130_FD_SC_HS__DFRTP_2%A_1271_74# 1 2 9 12 13 15 16 17 19 20 22 25
+ 27 28 29 31 34 36 37 41 42 43 48 50
c148 41 0 1.53326e-19 $X=7.54 $Y=2.475
c149 17 0 4.77539e-20 $X=9.035 $Y=1.63
c150 12 0 1.36674e-19 $X=8.945 $Y=2.3
r151 54 58 13.0505 $w=2.77e-07 $l=7.5e-08 $layer=POLY_cond $X=8.87 $Y=1.722
+ $X2=8.945 $Y2=1.722
r152 53 54 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.87
+ $Y=1.725 $X2=8.87 $Y2=1.725
r153 50 53 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=8.87 $Y=1.645 $X2=8.87
+ $Y2=1.725
r154 46 48 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=6.44 $Y=1.6 $X2=6.6
+ $Y2=1.6
r155 42 50 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.705 $Y=1.645
+ $X2=8.87 $Y2=1.645
r156 42 43 70.4599 $w=1.68e-07 $l=1.08e-06 $layer=LI1_cond $X=8.705 $Y=1.645
+ $X2=7.625 $Y2=1.645
r157 40 43 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.54 $Y=1.73
+ $X2=7.625 $Y2=1.645
r158 40 41 48.6043 $w=1.68e-07 $l=7.45e-07 $layer=LI1_cond $X=7.54 $Y=1.73
+ $X2=7.54 $Y2=2.475
r159 37 39 14.1436 $w=3.28e-07 $l=4.05e-07 $layer=LI1_cond $X=6.685 $Y=2.64
+ $X2=7.09 $Y2=2.64
r160 36 41 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=7.455 $Y=2.64
+ $X2=7.54 $Y2=2.475
r161 36 39 12.7467 $w=3.28e-07 $l=3.65e-07 $layer=LI1_cond $X=7.455 $Y=2.64
+ $X2=7.09 $Y2=2.64
r162 32 45 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.525 $Y=0.72
+ $X2=6.44 $Y2=0.72
r163 32 34 19.5915 $w=2.48e-07 $l=4.25e-07 $layer=LI1_cond $X=6.525 $Y=0.72
+ $X2=6.95 $Y2=0.72
r164 31 37 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=6.6 $Y=2.475
+ $X2=6.685 $Y2=2.64
r165 30 48 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.6 $Y=1.685
+ $X2=6.6 $Y2=1.6
r166 30 31 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=6.6 $Y=1.685
+ $X2=6.6 $Y2=2.475
r167 29 46 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.44 $Y=1.515
+ $X2=6.44 $Y2=1.6
r168 28 45 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.44 $Y=0.845
+ $X2=6.44 $Y2=0.72
r169 28 29 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=6.44 $Y=0.845
+ $X2=6.44 $Y2=1.515
r170 23 27 18.8402 $w=1.65e-07 $l=9.60469e-08 $layer=POLY_cond $X=9.61 $Y=1.555
+ $X2=9.562 $Y2=1.63
r171 23 25 417.904 $w=1.5e-07 $l=8.15e-07 $layer=POLY_cond $X=9.61 $Y=1.555
+ $X2=9.61 $Y2=0.74
r172 20 22 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=9.53 $Y=1.97
+ $X2=9.53 $Y2=2.465
r173 19 20 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=9.53 $Y=1.88 $X2=9.53
+ $Y2=1.97
r174 18 27 18.8402 $w=1.65e-07 $l=8.95824e-08 $layer=POLY_cond $X=9.53 $Y=1.705
+ $X2=9.562 $Y2=1.63
r175 18 19 68.0242 $w=1.8e-07 $l=1.75e-07 $layer=POLY_cond $X=9.53 $Y=1.705
+ $X2=9.53 $Y2=1.88
r176 17 58 25.7246 $w=2.77e-07 $l=1.29399e-07 $layer=POLY_cond $X=9.035 $Y=1.63
+ $X2=8.945 $Y2=1.722
r177 16 27 6.66866 $w=1.5e-07 $l=1.22e-07 $layer=POLY_cond $X=9.44 $Y=1.63
+ $X2=9.562 $Y2=1.63
r178 16 17 207.67 $w=1.5e-07 $l=4.05e-07 $layer=POLY_cond $X=9.44 $Y=1.63
+ $X2=9.035 $Y2=1.63
r179 13 15 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=8.945 $Y=2.39
+ $X2=8.945 $Y2=2.675
r180 12 13 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=8.945 $Y=2.3
+ $X2=8.945 $Y2=2.39
r181 11 58 12.8788 $w=1.8e-07 $l=1.68e-07 $layer=POLY_cond $X=8.945 $Y=1.89
+ $X2=8.945 $Y2=1.722
r182 11 12 159.371 $w=1.8e-07 $l=4.1e-07 $layer=POLY_cond $X=8.945 $Y=1.89
+ $X2=8.945 $Y2=2.3
r183 7 54 41.7617 $w=2.77e-07 $l=3.12538e-07 $layer=POLY_cond $X=8.63 $Y=1.555
+ $X2=8.87 $Y2=1.722
r184 7 9 482 $w=1.5e-07 $l=9.4e-07 $layer=POLY_cond $X=8.63 $Y=1.555 $X2=8.63
+ $Y2=0.615
r185 2 39 300 $w=1.7e-07 $l=1.09135e-06 $layer=licon1_PDIFF $count=2 $X=6.485
+ $Y=1.81 $X2=7.09 $Y2=2.64
r186 1 45 182 $w=1.7e-07 $l=3.83732e-07 $layer=licon1_NDIFF $count=1 $X=6.355
+ $Y=0.37 $X2=6.52 $Y2=0.68
r187 1 34 182 $w=1.7e-07 $l=7.33809e-07 $layer=licon1_NDIFF $count=1 $X=6.355
+ $Y=0.37 $X2=6.95 $Y2=0.68
.ends

.subckt PM_SKY130_FD_SC_HS__DFRTP_2%A_1921_409# 1 2 7 10 11 13 16 18 21 22 24 27
+ 29 30 33 37 41 46 49
c72 49 0 4.37308e-20 $X=10.09 $Y=1.375
c73 33 0 1.36674e-19 $X=9.755 $Y=2.195
r74 47 49 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=10.09 $Y=1.465
+ $X2=10.09 $Y2=1.375
r75 46 47 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.09
+ $Y=1.465 $X2=10.09 $Y2=1.465
r76 44 46 9.25447 $w=3.28e-07 $l=2.65e-07 $layer=LI1_cond $X=9.825 $Y=1.465
+ $X2=10.09 $Y2=1.465
r77 42 44 1.22229 $w=3.28e-07 $l=3.5e-08 $layer=LI1_cond $X=9.79 $Y=1.465
+ $X2=9.825 $Y2=1.465
r78 39 42 2.13598 $w=2.6e-07 $l=1.65e-07 $layer=LI1_cond $X=9.79 $Y=1.63
+ $X2=9.79 $Y2=1.465
r79 39 41 17.7299 $w=2.58e-07 $l=4e-07 $layer=LI1_cond $X=9.79 $Y=1.63 $X2=9.79
+ $Y2=2.03
r80 35 44 0.716491 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=9.825 $Y=1.3
+ $X2=9.825 $Y2=1.465
r81 35 37 27.4142 $w=3.28e-07 $l=7.85e-07 $layer=LI1_cond $X=9.825 $Y=1.3
+ $X2=9.825 $Y2=0.515
r82 33 41 6.31279 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=9.755 $Y=2.195
+ $X2=9.755 $Y2=2.03
r83 25 30 18.8402 $w=1.65e-07 $l=8.21584e-08 $layer=POLY_cond $X=11.03 $Y=1.3
+ $X2=11.015 $Y2=1.375
r84 25 27 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=11.03 $Y=1.3
+ $X2=11.03 $Y2=0.74
r85 22 24 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=11.015 $Y=1.765
+ $X2=11.015 $Y2=2.4
r86 21 22 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=11.015 $Y=1.675
+ $X2=11.015 $Y2=1.765
r87 20 30 18.8402 $w=1.65e-07 $l=7.5e-08 $layer=POLY_cond $X=11.015 $Y=1.45
+ $X2=11.015 $Y2=1.375
r88 20 21 87.4597 $w=1.8e-07 $l=2.25e-07 $layer=POLY_cond $X=11.015 $Y=1.45
+ $X2=11.015 $Y2=1.675
r89 19 29 13.2179 $w=1.5e-07 $l=1e-07 $layer=POLY_cond $X=10.675 $Y=1.375
+ $X2=10.575 $Y2=1.375
r90 18 30 6.66866 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=10.925 $Y=1.375
+ $X2=11.015 $Y2=1.375
r91 18 19 128.191 $w=1.5e-07 $l=2.5e-07 $layer=POLY_cond $X=10.925 $Y=1.375
+ $X2=10.675 $Y2=1.375
r92 14 29 10.9219 $w=1.5e-07 $l=8.66025e-08 $layer=POLY_cond $X=10.6 $Y=1.3
+ $X2=10.575 $Y2=1.375
r93 14 16 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=10.6 $Y=1.3 $X2=10.6
+ $Y2=0.74
r94 11 13 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=10.565 $Y=1.765
+ $X2=10.565 $Y2=2.4
r95 10 11 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=10.565 $Y=1.675
+ $X2=10.565 $Y2=1.765
r96 9 29 10.9219 $w=1.8e-07 $l=7.98436e-08 $layer=POLY_cond $X=10.565 $Y=1.45
+ $X2=10.575 $Y2=1.375
r97 9 10 87.4597 $w=1.8e-07 $l=2.25e-07 $layer=POLY_cond $X=10.565 $Y=1.45
+ $X2=10.565 $Y2=1.675
r98 8 49 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=10.255 $Y=1.375
+ $X2=10.09 $Y2=1.375
r99 7 29 13.2179 $w=1.5e-07 $l=1e-07 $layer=POLY_cond $X=10.475 $Y=1.375
+ $X2=10.575 $Y2=1.375
r100 7 8 112.809 $w=1.5e-07 $l=2.2e-07 $layer=POLY_cond $X=10.475 $Y=1.375
+ $X2=10.255 $Y2=1.375
r101 2 33 300 $w=1.7e-07 $l=2.12132e-07 $layer=licon1_PDIFF $count=2 $X=9.605
+ $Y=2.045 $X2=9.755 $Y2=2.195
r102 1 37 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=9.685
+ $Y=0.37 $X2=9.825 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__DFRTP_2%VPWR 1 2 3 4 5 6 7 8 9 28 30 34 38 42 44 48
+ 54 58 62 66 68 73 74 75 77 82 87 95 107 111 120 123 126 129 132 135 139
r150 138 139 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.28 $Y=3.33
+ $X2=11.28 $Y2=3.33
r151 135 136 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.32 $Y=3.33
+ $X2=10.32 $Y2=3.33
r152 132 133 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r153 129 130 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r154 127 130 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=5.52 $Y2=3.33
r155 126 127 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r156 123 124 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r157 120 121 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r158 117 118 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r159 115 139 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.8 $Y=3.33
+ $X2=11.28 $Y2=3.33
r160 115 136 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.8 $Y=3.33
+ $X2=10.32 $Y2=3.33
r161 114 115 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.8 $Y=3.33
+ $X2=10.8 $Y2=3.33
r162 112 135 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.48 $Y=3.33
+ $X2=10.315 $Y2=3.33
r163 112 114 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=10.48 $Y=3.33
+ $X2=10.8 $Y2=3.33
r164 111 138 4.01252 $w=1.7e-07 $l=1.82e-07 $layer=LI1_cond $X=11.155 $Y=3.33
+ $X2=11.337 $Y2=3.33
r165 111 114 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=11.155 $Y=3.33
+ $X2=10.8 $Y2=3.33
r166 110 136 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.84 $Y=3.33
+ $X2=10.32 $Y2=3.33
r167 109 110 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.84 $Y=3.33
+ $X2=9.84 $Y2=3.33
r168 107 135 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.15 $Y=3.33
+ $X2=10.315 $Y2=3.33
r169 107 109 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=10.15 $Y=3.33
+ $X2=9.84 $Y2=3.33
r170 106 110 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=8.88 $Y=3.33
+ $X2=9.84 $Y2=3.33
r171 106 133 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=8.88 $Y=3.33
+ $X2=7.92 $Y2=3.33
r172 105 106 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r173 103 132 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.125 $Y=3.33
+ $X2=7.96 $Y2=3.33
r174 103 105 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=8.125 $Y=3.33
+ $X2=8.88 $Y2=3.33
r175 102 133 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=7.92 $Y2=3.33
r176 101 102 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r177 99 102 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=6 $Y=3.33
+ $X2=7.44 $Y2=3.33
r178 98 101 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=6 $Y=3.33
+ $X2=7.44 $Y2=3.33
r179 98 99 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r180 96 129 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.845 $Y=3.33
+ $X2=5.68 $Y2=3.33
r181 96 98 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=5.845 $Y=3.33
+ $X2=6 $Y2=3.33
r182 95 132 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.795 $Y=3.33
+ $X2=7.96 $Y2=3.33
r183 95 101 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=7.795 $Y=3.33
+ $X2=7.44 $Y2=3.33
r184 94 127 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=4.56 $Y2=3.33
r185 93 94 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r186 91 94 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=4.08 $Y2=3.33
r187 91 124 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=2.16 $Y2=3.33
r188 90 93 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=2.64 $Y=3.33
+ $X2=4.08 $Y2=3.33
r189 90 91 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r190 88 123 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.315 $Y=3.33
+ $X2=2.15 $Y2=3.33
r191 88 90 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=2.315 $Y=3.33
+ $X2=2.64 $Y2=3.33
r192 87 126 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.42 $Y=3.33
+ $X2=4.585 $Y2=3.33
r193 87 93 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=4.42 $Y=3.33
+ $X2=4.08 $Y2=3.33
r194 86 124 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r195 86 121 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r196 85 86 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r197 83 120 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.335 $Y=3.33
+ $X2=1.17 $Y2=3.33
r198 83 85 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.335 $Y=3.33
+ $X2=1.68 $Y2=3.33
r199 82 123 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.985 $Y=3.33
+ $X2=2.15 $Y2=3.33
r200 82 85 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.985 $Y=3.33
+ $X2=1.68 $Y2=3.33
r201 81 121 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r202 81 118 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r203 80 81 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r204 78 117 4.75569 $w=1.7e-07 $l=2.18e-07 $layer=LI1_cond $X=0.435 $Y=3.33
+ $X2=0.217 $Y2=3.33
r205 78 80 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.435 $Y=3.33
+ $X2=0.72 $Y2=3.33
r206 77 120 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.005 $Y=3.33
+ $X2=1.17 $Y2=3.33
r207 77 80 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=1.005 $Y=3.33
+ $X2=0.72 $Y2=3.33
r208 75 99 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=5.76 $Y=3.33
+ $X2=6 $Y2=3.33
r209 75 130 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=5.76 $Y=3.33
+ $X2=5.52 $Y2=3.33
r210 73 105 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=9.09 $Y=3.33
+ $X2=8.88 $Y2=3.33
r211 73 74 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.09 $Y=3.33
+ $X2=9.255 $Y2=3.33
r212 72 109 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=9.42 $Y=3.33
+ $X2=9.84 $Y2=3.33
r213 72 74 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.42 $Y=3.33
+ $X2=9.255 $Y2=3.33
r214 68 71 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=11.28 $Y=1.985
+ $X2=11.28 $Y2=2.815
r215 66 138 3.13065 $w=2.5e-07 $l=1.09864e-07 $layer=LI1_cond $X=11.28 $Y=3.245
+ $X2=11.337 $Y2=3.33
r216 66 71 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=11.28 $Y=3.245
+ $X2=11.28 $Y2=2.815
r217 62 65 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=10.315 $Y=1.985
+ $X2=10.315 $Y2=2.815
r218 60 135 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=10.315 $Y=3.245
+ $X2=10.315 $Y2=3.33
r219 60 65 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=10.315 $Y=3.245
+ $X2=10.315 $Y2=2.815
r220 56 74 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.255 $Y=3.245
+ $X2=9.255 $Y2=3.33
r221 56 58 19.9058 $w=3.28e-07 $l=5.7e-07 $layer=LI1_cond $X=9.255 $Y=3.245
+ $X2=9.255 $Y2=2.675
r222 52 132 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.96 $Y=3.245
+ $X2=7.96 $Y2=3.33
r223 52 54 19.9058 $w=3.28e-07 $l=5.7e-07 $layer=LI1_cond $X=7.96 $Y=3.245
+ $X2=7.96 $Y2=2.675
r224 48 51 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=5.68 $Y=1.91
+ $X2=5.68 $Y2=2.59
r225 46 129 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.68 $Y=3.245
+ $X2=5.68 $Y2=3.33
r226 46 51 22.8742 $w=3.28e-07 $l=6.55e-07 $layer=LI1_cond $X=5.68 $Y=3.245
+ $X2=5.68 $Y2=2.59
r227 45 126 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.75 $Y=3.33
+ $X2=4.585 $Y2=3.33
r228 44 129 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.515 $Y=3.33
+ $X2=5.68 $Y2=3.33
r229 44 45 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=5.515 $Y=3.33
+ $X2=4.75 $Y2=3.33
r230 40 126 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.585 $Y=3.245
+ $X2=4.585 $Y2=3.33
r231 40 42 14.1436 $w=3.28e-07 $l=4.05e-07 $layer=LI1_cond $X=4.585 $Y=3.245
+ $X2=4.585 $Y2=2.84
r232 36 123 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.15 $Y=3.245
+ $X2=2.15 $Y2=3.33
r233 36 38 16.7628 $w=3.28e-07 $l=4.8e-07 $layer=LI1_cond $X=2.15 $Y=3.245
+ $X2=2.15 $Y2=2.765
r234 32 120 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.17 $Y=3.245
+ $X2=1.17 $Y2=3.33
r235 32 34 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=1.17 $Y=3.245
+ $X2=1.17 $Y2=2.78
r236 28 117 3.01048 $w=3.3e-07 $l=1.08305e-07 $layer=LI1_cond $X=0.27 $Y=3.245
+ $X2=0.217 $Y2=3.33
r237 28 30 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=0.27 $Y=3.245
+ $X2=0.27 $Y2=2.75
r238 9 71 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=11.09
+ $Y=1.84 $X2=11.24 $Y2=2.815
r239 9 68 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=11.09
+ $Y=1.84 $X2=11.24 $Y2=1.985
r240 8 65 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=10.17
+ $Y=1.84 $X2=10.315 $Y2=2.815
r241 8 62 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=10.17
+ $Y=1.84 $X2=10.315 $Y2=1.985
r242 7 58 600 $w=1.7e-07 $l=3.23381e-07 $layer=licon1_PDIFF $count=1 $X=9.02
+ $Y=2.465 $X2=9.255 $Y2=2.675
r243 6 54 600 $w=1.7e-07 $l=2.74955e-07 $layer=licon1_PDIFF $count=1 $X=7.81
+ $Y=2.465 $X2=7.96 $Y2=2.675
r244 5 51 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=5.535
+ $Y=1.735 $X2=5.68 $Y2=2.59
r245 5 48 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=5.535
+ $Y=1.735 $X2=5.68 $Y2=1.91
r246 4 42 600 $w=1.7e-07 $l=6.62156e-07 $layer=licon1_PDIFF $count=1 $X=4.35
+ $Y=2.285 $X2=4.585 $Y2=2.84
r247 3 38 600 $w=1.7e-07 $l=1.02727e-06 $layer=licon1_PDIFF $count=1 $X=2
+ $Y=1.81 $X2=2.15 $Y2=2.765
r248 2 34 600 $w=1.7e-07 $l=3.05941e-07 $layer=licon1_PDIFF $count=1 $X=1.02
+ $Y=2.54 $X2=1.17 $Y2=2.78
r249 1 30 600 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.54 $X2=0.27 $Y2=2.75
.ends

.subckt PM_SKY130_FD_SC_HS__DFRTP_2%A_30_78# 1 2 3 4 13 15 17 20 21 25 27 30 32
+ 38 43
c110 30 0 5.51194e-20 $X=3.675 $Y=2.075
r111 38 40 5.47085 $w=2.23e-07 $l=1e-07 $layer=LI1_cond $X=3.14 $Y=2.405
+ $X2=3.14 $Y2=2.505
r112 37 38 13.4036 $w=2.23e-07 $l=2.45e-07 $layer=LI1_cond $X=3.14 $Y=2.16
+ $X2=3.14 $Y2=2.405
r113 32 34 5.06376 $w=3.28e-07 $l=1.45e-07 $layer=LI1_cond $X=0.295 $Y=0.6
+ $X2=0.295 $Y2=0.745
r114 29 43 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.675 $Y=1.405
+ $X2=3.675 $Y2=1.32
r115 29 30 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.675 $Y=1.405
+ $X2=3.675 $Y2=2.075
r116 28 37 2.32876 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.265 $Y=2.16
+ $X2=3.14 $Y2=2.16
r117 27 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.59 $Y=2.16
+ $X2=3.675 $Y2=2.075
r118 27 28 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=3.59 $Y=2.16
+ $X2=3.265 $Y2=2.16
r119 23 43 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=3.335 $Y=1.32
+ $X2=3.675 $Y2=1.32
r120 23 25 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=3.335 $Y=1.235
+ $X2=3.335 $Y2=0.9
r121 22 36 1.06262 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=0.835 $Y=2.405
+ $X2=0.735 $Y2=2.405
r122 21 38 2.32876 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.015 $Y=2.405
+ $X2=3.14 $Y2=2.405
r123 21 22 142.225 $w=1.68e-07 $l=2.18e-06 $layer=LI1_cond $X=3.015 $Y=2.405
+ $X2=0.835 $Y2=2.405
r124 20 36 5.81257 $w=1.8e-07 $l=9.21954e-08 $layer=LI1_cond $X=0.75 $Y=2.32
+ $X2=0.735 $Y2=2.405
r125 19 20 97.2086 $w=1.68e-07 $l=1.49e-06 $layer=LI1_cond $X=0.75 $Y=0.83
+ $X2=0.75 $Y2=2.32
r126 15 36 13.2636 $w=2e-07 $l=2.15e-07 $layer=LI1_cond $X=0.735 $Y=2.62
+ $X2=0.735 $Y2=2.405
r127 15 17 7.20909 $w=1.98e-07 $l=1.3e-07 $layer=LI1_cond $X=0.735 $Y=2.62
+ $X2=0.735 $Y2=2.75
r128 14 34 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.46 $Y=0.745
+ $X2=0.295 $Y2=0.745
r129 13 19 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.665 $Y=0.745
+ $X2=0.75 $Y2=0.83
r130 13 14 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=0.665 $Y=0.745
+ $X2=0.46 $Y2=0.745
r131 4 40 600 $w=1.7e-07 $l=2.81425e-07 $layer=licon1_PDIFF $count=1 $X=3.04
+ $Y=2.285 $X2=3.18 $Y2=2.505
r132 3 17 600 $w=1.7e-07 $l=2.74955e-07 $layer=licon1_PDIFF $count=1 $X=0.57
+ $Y=2.54 $X2=0.72 $Y2=2.75
r133 2 25 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=3.15
+ $Y=0.69 $X2=3.295 $Y2=0.9
r134 1 32 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=0.15
+ $Y=0.39 $X2=0.295 $Y2=0.6
.ends

.subckt PM_SKY130_FD_SC_HS__DFRTP_2%Q 1 2 7 8 9 10 11 12 13
r22 12 13 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=10.815 $Y=2.405
+ $X2=10.815 $Y2=2.775
r23 11 12 14.6675 $w=3.28e-07 $l=4.2e-07 $layer=LI1_cond $X=10.815 $Y=1.985
+ $X2=10.815 $Y2=2.405
r24 10 11 11.1752 $w=3.28e-07 $l=3.2e-07 $layer=LI1_cond $X=10.815 $Y=1.665
+ $X2=10.815 $Y2=1.985
r25 9 10 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=10.815 $Y=1.295
+ $X2=10.815 $Y2=1.665
r26 8 9 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=10.815 $Y=0.925
+ $X2=10.815 $Y2=1.295
r27 7 8 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=10.815 $Y=0.515
+ $X2=10.815 $Y2=0.925
r28 2 13 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=10.64
+ $Y=1.84 $X2=10.79 $Y2=2.815
r29 2 11 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=10.64
+ $Y=1.84 $X2=10.79 $Y2=1.985
r30 1 7 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=10.675
+ $Y=0.37 $X2=10.815 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__DFRTP_2%VGND 1 2 3 4 5 6 7 24 28 32 36 40 42 44 47
+ 48 49 55 59 67 75 80 85 91 101 104 107 111
r116 110 111 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.28 $Y=0
+ $X2=11.28 $Y2=0
r117 107 108 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.32 $Y=0
+ $X2=10.32 $Y2=0
r118 104 105 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.36 $Y=0
+ $X2=9.36 $Y2=0
r119 101 102 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=0
+ $X2=7.92 $Y2=0
r120 91 92 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r121 89 111 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.8 $Y=0
+ $X2=11.28 $Y2=0
r122 89 108 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.8 $Y=0
+ $X2=10.32 $Y2=0
r123 88 89 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.8 $Y=0 $X2=10.8
+ $Y2=0
r124 86 107 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=10.47 $Y=0
+ $X2=10.345 $Y2=0
r125 86 88 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=10.47 $Y=0 $X2=10.8
+ $Y2=0
r126 85 110 4.01803 $w=1.7e-07 $l=1.8e-07 $layer=LI1_cond $X=11.16 $Y=0
+ $X2=11.34 $Y2=0
r127 85 88 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=11.16 $Y=0 $X2=10.8
+ $Y2=0
r128 84 108 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.84 $Y=0
+ $X2=10.32 $Y2=0
r129 84 105 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.84 $Y=0
+ $X2=9.36 $Y2=0
r130 83 84 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.84 $Y=0 $X2=9.84
+ $Y2=0
r131 81 104 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=9.48 $Y=0
+ $X2=9.355 $Y2=0
r132 81 83 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=9.48 $Y=0 $X2=9.84
+ $Y2=0
r133 80 107 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=10.22 $Y=0
+ $X2=10.345 $Y2=0
r134 80 83 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=10.22 $Y=0 $X2=9.84
+ $Y2=0
r135 79 105 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=0
+ $X2=9.36 $Y2=0
r136 79 102 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=8.88 $Y=0
+ $X2=7.92 $Y2=0
r137 78 79 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.88 $Y=0 $X2=8.88
+ $Y2=0
r138 76 101 10.1275 $w=1.7e-07 $l=2.1e-07 $layer=LI1_cond $X=8.19 $Y=0 $X2=7.98
+ $Y2=0
r139 76 78 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=8.19 $Y=0 $X2=8.88
+ $Y2=0
r140 75 104 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=9.23 $Y=0
+ $X2=9.355 $Y2=0
r141 75 78 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=9.23 $Y=0 $X2=8.88
+ $Y2=0
r142 74 102 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=0
+ $X2=7.92 $Y2=0
r143 73 74 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=7.44 $Y=0
+ $X2=7.44 $Y2=0
r144 71 96 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=5.04
+ $Y2=0
r145 70 73 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=5.52 $Y=0 $X2=7.44
+ $Y2=0
r146 70 71 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=5.52 $Y=0
+ $X2=5.52 $Y2=0
r147 68 70 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=5.345 $Y=0
+ $X2=5.52 $Y2=0
r148 67 101 10.1275 $w=1.7e-07 $l=2.1e-07 $layer=LI1_cond $X=7.77 $Y=0 $X2=7.98
+ $Y2=0
r149 67 73 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=7.77 $Y=0 $X2=7.44
+ $Y2=0
r150 66 96 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=5.04
+ $Y2=0
r151 65 66 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.56 $Y=0
+ $X2=4.56 $Y2=0
r152 63 66 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=2.64 $Y=0
+ $X2=4.56 $Y2=0
r153 63 92 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=2.16
+ $Y2=0
r154 62 65 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=2.64 $Y=0 $X2=4.56
+ $Y2=0
r155 62 63 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.64 $Y=0
+ $X2=2.64 $Y2=0
r156 60 91 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.34 $Y=0 $X2=2.175
+ $Y2=0
r157 60 62 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=2.34 $Y=0 $X2=2.64
+ $Y2=0
r158 59 98 7.59257 $w=4.23e-07 $l=2.8e-07 $layer=LI1_cond $X=5.132 $Y=0
+ $X2=5.132 $Y2=0.28
r159 59 68 6.14847 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=5.132 $Y=0
+ $X2=5.345 $Y2=0
r160 59 96 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r161 59 65 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=4.92 $Y=0 $X2=4.56
+ $Y2=0
r162 58 92 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r163 57 58 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r164 55 91 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.01 $Y=0 $X2=2.175
+ $Y2=0
r165 55 57 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=2.01 $Y=0 $X2=1.68
+ $Y2=0
r166 53 58 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r167 52 53 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r168 49 74 0.468274 $w=4.9e-07 $l=1.68e-06 $layer=MET1_cond $X=5.76 $Y=0
+ $X2=7.44 $Y2=0
r169 49 71 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=5.76 $Y=0
+ $X2=5.52 $Y2=0
r170 47 52 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=1.03 $Y=0 $X2=0.72
+ $Y2=0
r171 47 48 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.03 $Y=0 $X2=1.155
+ $Y2=0
r172 46 57 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=1.28 $Y=0 $X2=1.68
+ $Y2=0
r173 46 48 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.28 $Y=0 $X2=1.155
+ $Y2=0
r174 42 110 3.12513 $w=2.5e-07 $l=1.09087e-07 $layer=LI1_cond $X=11.285 $Y=0.085
+ $X2=11.34 $Y2=0
r175 42 44 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=11.285 $Y=0.085
+ $X2=11.285 $Y2=0.515
r176 38 107 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=10.345 $Y=0.085
+ $X2=10.345 $Y2=0
r177 38 40 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=10.345 $Y=0.085
+ $X2=10.345 $Y2=0.515
r178 34 104 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=9.355 $Y=0.085
+ $X2=9.355 $Y2=0
r179 34 36 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=9.355 $Y=0.085
+ $X2=9.355 $Y2=0.515
r180 30 101 1.60615 $w=4.2e-07 $l=8.5e-08 $layer=LI1_cond $X=7.98 $Y=0.085
+ $X2=7.98 $Y2=0
r181 30 32 12.7592 $w=4.18e-07 $l=4.65e-07 $layer=LI1_cond $X=7.98 $Y=0.085
+ $X2=7.98 $Y2=0.55
r182 26 91 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.175 $Y=0.085
+ $X2=2.175 $Y2=0
r183 26 28 18.6835 $w=3.28e-07 $l=5.35e-07 $layer=LI1_cond $X=2.175 $Y=0.085
+ $X2=2.175 $Y2=0.62
r184 22 48 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.155 $Y=0.085
+ $X2=1.155 $Y2=0
r185 22 24 23.5098 $w=2.48e-07 $l=5.1e-07 $layer=LI1_cond $X=1.155 $Y=0.085
+ $X2=1.155 $Y2=0.595
r186 7 44 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=11.105
+ $Y=0.37 $X2=11.245 $Y2=0.515
r187 6 40 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=10.24
+ $Y=0.37 $X2=10.385 $Y2=0.515
r188 5 36 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=9.255
+ $Y=0.37 $X2=9.395 $Y2=0.515
r189 4 32 182 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=1 $X=7.795
+ $Y=0.405 $X2=7.98 $Y2=0.55
r190 3 98 182 $w=1.7e-07 $l=5.2607e-07 $layer=licon1_NDIFF $count=1 $X=4.865
+ $Y=0.69 $X2=5.13 $Y2=0.28
r191 2 28 182 $w=1.7e-07 $l=3.39116e-07 $layer=licon1_NDIFF $count=1 $X=1.965
+ $Y=0.37 $X2=2.175 $Y2=0.62
r192 1 24 182 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_NDIFF $count=1 $X=0.975
+ $Y=0.39 $X2=1.115 $Y2=0.595
.ends

