# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_hs__or4b_4
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_hs__or4b_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  7.200000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.411000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.005000 1.450000 1.335000 1.780000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.411000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.110000 2.035000 1.280000 ;
        RECT 0.125000 1.280000 0.835000 1.550000 ;
        RECT 1.705000 1.280000 2.035000 1.550000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.411000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2.495000 1.180000 2.785000 1.225000 ;
        RECT 2.495000 1.225000 4.225000 1.365000 ;
        RECT 2.495000 1.365000 2.785000 1.410000 ;
        RECT 3.935000 1.180000 4.225000 1.225000 ;
        RECT 3.935000 1.365000 4.225000 1.410000 ;
    END
  END C
  PIN D_N
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.445000 1.180000 4.815000 1.550000 ;
    END
  END D_N
  PIN X
    ANTENNADIFFAREA  1.178900 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.325000 0.350000 5.655000 0.980000 ;
        RECT 5.325000 0.980000 6.575000 1.150000 ;
        RECT 5.410000 1.820000 7.075000 2.150000 ;
        RECT 5.410000 2.150000 5.690000 2.980000 ;
        RECT 6.325000 0.350000 6.575000 0.980000 ;
        RECT 6.325000 1.150000 6.575000 1.300000 ;
        RECT 6.325000 1.300000 6.655000 1.470000 ;
        RECT 6.360000 2.150000 6.590000 2.980000 ;
        RECT 6.365000 1.470000 6.655000 1.820000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 7.200000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 7.200000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 7.200000 0.085000 ;
      RECT 0.000000  3.245000 7.200000 3.415000 ;
      RECT 0.115000  0.350000 0.445000 0.770000 ;
      RECT 0.115000  0.770000 3.270000 0.840000 ;
      RECT 0.115000  0.840000 5.155000 0.940000 ;
      RECT 0.115000  1.940000 0.445000 1.950000 ;
      RECT 0.115000  1.950000 2.345000 2.120000 ;
      RECT 0.115000  2.120000 0.445000 2.980000 ;
      RECT 0.615000  0.085000 0.945000 0.600000 ;
      RECT 0.645000  2.290000 1.845000 2.460000 ;
      RECT 0.645000  2.460000 0.815000 2.980000 ;
      RECT 1.015000  2.630000 1.345000 3.245000 ;
      RECT 1.115000  0.350000 2.200000 0.770000 ;
      RECT 1.515000  2.460000 1.845000 2.980000 ;
      RECT 2.015000  2.120000 2.345000 2.360000 ;
      RECT 2.015000  2.360000 4.195000 2.530000 ;
      RECT 2.015000  2.530000 2.345000 2.980000 ;
      RECT 2.245000  1.180000 2.725000 1.780000 ;
      RECT 2.370000  0.085000 2.725000 0.600000 ;
      RECT 2.515000  2.700000 3.745000 2.980000 ;
      RECT 2.895000  0.350000 3.270000 0.770000 ;
      RECT 2.895000  0.940000 5.155000 1.010000 ;
      RECT 2.895000  1.010000 3.270000 1.130000 ;
      RECT 2.895000  1.130000 3.065000 2.020000 ;
      RECT 2.895000  2.020000 3.295000 2.190000 ;
      RECT 3.235000  1.470000 3.635000 1.720000 ;
      RECT 3.235000  1.720000 4.755000 1.800000 ;
      RECT 3.440000  0.340000 4.565000 0.670000 ;
      RECT 3.465000  1.800000 4.755000 1.890000 ;
      RECT 3.865000  1.180000 4.195000 1.510000 ;
      RECT 3.945000  2.060000 4.195000 2.360000 ;
      RECT 3.945000  2.530000 4.195000 2.980000 ;
      RECT 4.425000  1.890000 4.755000 2.860000 ;
      RECT 4.825000  0.085000 5.155000 0.670000 ;
      RECT 4.960000  1.820000 5.210000 3.245000 ;
      RECT 4.985000  1.010000 5.155000 1.320000 ;
      RECT 4.985000  1.320000 6.155000 1.650000 ;
      RECT 5.825000  0.085000 6.155000 0.810000 ;
      RECT 5.860000  2.320000 6.190000 3.245000 ;
      RECT 6.755000  0.085000 7.085000 1.130000 ;
      RECT 6.760000  2.320000 7.090000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  1.210000 2.725000 1.380000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  1.210000 4.165000 1.380000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
  END
END sky130_fd_sc_hs__or4b_4
END LIBRARY
