# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_hs__o21ba_1
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_hs__o21ba_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.840000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.130000 0.550000 1.800000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.835000 1.130000 1.315000 1.800000 ;
    END
  END A2
  PIN B1_N
    ANTENNAGATEAREA  0.208500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.515000 1.180000 2.845000 1.550000 ;
    END
  END B1_N
  PIN X
    ANTENNADIFFAREA  0.541300 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.390000 0.350000 3.755000 1.130000 ;
        RECT 3.395000 1.820000 3.755000 2.980000 ;
        RECT 3.585000 1.130000 3.755000 1.820000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 3.840000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 3.840000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.840000 0.085000 ;
      RECT 0.000000  3.245000 3.840000 3.415000 ;
      RECT 0.115000  0.350000 0.445000 0.790000 ;
      RECT 0.115000  0.790000 1.445000 0.960000 ;
      RECT 0.115000  1.970000 0.445000 3.245000 ;
      RECT 0.615000  0.085000 0.945000 0.620000 ;
      RECT 1.055000  1.970000 1.785000 2.320000 ;
      RECT 1.055000  2.320000 3.225000 2.490000 ;
      RECT 1.055000  2.490000 1.385000 2.980000 ;
      RECT 1.115000  0.350000 1.445000 0.790000 ;
      RECT 1.555000  2.660000 1.885000 3.245000 ;
      RECT 1.615000  0.350000 1.945000 1.030000 ;
      RECT 1.615000  1.030000 1.785000 1.970000 ;
      RECT 1.975000  1.220000 2.305000 1.820000 ;
      RECT 1.975000  1.820000 2.690000 2.150000 ;
      RECT 2.135000  0.680000 2.720000 1.010000 ;
      RECT 2.135000  1.010000 2.305000 1.220000 ;
      RECT 2.890000  0.085000 3.220000 1.010000 ;
      RECT 2.895000  2.660000 3.225000 3.245000 ;
      RECT 3.055000  1.320000 3.415000 1.650000 ;
      RECT 3.055000  1.650000 3.225000 2.320000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
  END
END sky130_fd_sc_hs__o21ba_1
