* NGSPICE file created from sky130_fd_sc_hs__o32a_2.ext - technology: sky130A

.subckt sky130_fd_sc_hs__o32a_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
M1000 a_346_368# A1 VPWR VPB pshort w=1e+06u l=150000u
+  ad=2.7e+11p pd=2.54e+06u as=1.2072e+12p ps=8.76e+06u
M1001 a_83_264# B2 a_349_74# VNB nlowvt w=740000u l=150000u
+  ad=6.771e+11p pd=3.31e+06u as=7.289e+11p ps=6.41e+06u
M1002 a_349_74# A3 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=9.62e+11p ps=7.04e+06u
M1003 a_349_74# A1 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 VPWR a_83_264# X VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=3.36e+11p ps=2.84e+06u
M1005 X a_83_264# VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_430_368# A2 a_346_368# VPB pshort w=1e+06u l=150000u
+  ad=3.9e+11p pd=2.78e+06u as=0p ps=0u
M1007 a_349_74# B1 a_83_264# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_83_264# A3 a_430_368# VPB pshort w=1e+06u l=150000u
+  ad=4.2e+11p pd=2.84e+06u as=0p ps=0u
M1009 X a_83_264# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.072e+11p pd=2.04e+06u as=0p ps=0u
M1010 VGND A2 a_349_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VPWR B1 a_652_368# VPB pshort w=1e+06u l=150000u
+  ad=0p pd=0u as=4.2e+11p ps=2.84e+06u
M1012 a_652_368# B2 a_83_264# VPB pshort w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VGND a_83_264# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

