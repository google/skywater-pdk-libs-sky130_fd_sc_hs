* File: sky130_fd_sc_hs__a2bb2oi_1.pex.spice
* Created: Thu Aug 27 20:27:59 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HS__A2BB2OI_1%A1_N 2 3 5 8 10 14 15
r28 15 16 6.79937 $w=3.19e-07 $l=4.5e-08 $layer=POLY_cond $X=0.51 $Y=1.425
+ $X2=0.555 $Y2=1.425
r29 13 15 36.2633 $w=3.19e-07 $l=2.4e-07 $layer=POLY_cond $X=0.27 $Y=1.425
+ $X2=0.51 $Y2=1.425
r30 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.27
+ $Y=1.425 $X2=0.27 $Y2=1.425
r31 10 14 8.3814 $w=3.28e-07 $l=2.4e-07 $layer=LI1_cond $X=0.27 $Y=1.665
+ $X2=0.27 $Y2=1.425
r32 6 16 20.418 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.555 $Y=1.26
+ $X2=0.555 $Y2=1.425
r33 6 8 217.926 $w=1.5e-07 $l=4.25e-07 $layer=POLY_cond $X=0.555 $Y=1.26
+ $X2=0.555 $Y2=0.835
r34 3 5 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=0.51 $Y=1.885
+ $X2=0.51 $Y2=2.46
r35 2 3 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=0.51 $Y=1.795 $X2=0.51
+ $Y2=1.885
r36 1 15 16.143 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=0.51 $Y=1.59 $X2=0.51
+ $Y2=1.425
r37 1 2 79.6855 $w=1.8e-07 $l=2.05e-07 $layer=POLY_cond $X=0.51 $Y=1.59 $X2=0.51
+ $Y2=1.795
.ends

.subckt PM_SKY130_FD_SC_HS__A2BB2OI_1%A2_N 1 3 6 8 12
c39 12 0 8.79615e-20 $X=1.005 $Y=1.615
r40 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.005
+ $Y=1.615 $X2=1.005 $Y2=1.615
r41 8 12 9.95292 $w=3.28e-07 $l=2.85e-07 $layer=LI1_cond $X=0.72 $Y=1.615
+ $X2=1.005 $Y2=1.615
r42 4 11 38.6139 $w=3.32e-07 $l=1.67481e-07 $layer=POLY_cond $X=0.985 $Y=1.45
+ $X2=0.99 $Y2=1.615
r43 4 6 315.351 $w=1.5e-07 $l=6.15e-07 $layer=POLY_cond $X=0.985 $Y=1.45
+ $X2=0.985 $Y2=0.835
r44 1 11 53.8579 $w=3.32e-07 $l=3.11769e-07 $layer=POLY_cond $X=0.9 $Y=1.885
+ $X2=0.99 $Y2=1.615
r45 1 3 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=0.9 $Y=1.885 $X2=0.9
+ $Y2=2.46
.ends

.subckt PM_SKY130_FD_SC_HS__A2BB2OI_1%A_126_112# 1 2 7 9 12 14 15 18 20 21 24 26
+ 29 30
c70 15 0 1.45091e-19 $X=1.92 $Y=1.22
c71 14 0 9.59822e-20 $X=1.83 $Y=1.385
c72 7 0 1.19409e-19 $X=1.92 $Y=1.765
r73 34 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.545
+ $Y=1.385 $X2=1.545 $Y2=1.385
r74 29 31 1.30231 $w=4.78e-07 $l=5e-09 $layer=LI1_cond $X=1.2 $Y=2.115 $X2=1.2
+ $Y2=2.12
r75 29 30 9.39634 $w=4.78e-07 $l=1.65e-07 $layer=LI1_cond $X=1.2 $Y=2.115
+ $X2=1.2 $Y2=1.95
r76 26 34 8.95599 $w=3.21e-07 $l=2.22486e-07 $layer=LI1_cond $X=1.355 $Y=1.55
+ $X2=1.49 $Y2=1.385
r77 26 30 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=1.355 $Y=1.55
+ $X2=1.355 $Y2=1.95
r78 24 31 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=1.125 $Y=2.815
+ $X2=1.125 $Y2=2.12
r79 20 34 12.9221 $w=3.21e-07 $l=4.36348e-07 $layer=LI1_cond $X=1.27 $Y=1.045
+ $X2=1.49 $Y2=1.385
r80 20 21 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=1.27 $Y=1.045
+ $X2=0.935 $Y2=1.045
r81 16 21 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.77 $Y=0.96
+ $X2=0.935 $Y2=1.045
r82 16 18 4.36531 $w=3.28e-07 $l=1.25e-07 $layer=LI1_cond $X=0.77 $Y=0.96
+ $X2=0.77 $Y2=0.835
r83 14 35 49.8355 $w=3.3e-07 $l=2.85e-07 $layer=POLY_cond $X=1.83 $Y=1.385
+ $X2=1.545 $Y2=1.385
r84 14 15 66.2869 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.92 $Y=1.385
+ $X2=1.92 $Y2=1.22
r85 12 15 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.935 $Y=0.74
+ $X2=1.935 $Y2=1.22
r86 7 14 149.859 $w=1.8e-07 $l=3.8e-07 $layer=POLY_cond $X=1.92 $Y=1.765
+ $X2=1.92 $Y2=1.385
r87 7 9 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.92 $Y=1.765
+ $X2=1.92 $Y2=2.4
r88 2 29 400 $w=1.7e-07 $l=2.17428e-07 $layer=licon1_PDIFF $count=1 $X=0.975
+ $Y=1.96 $X2=1.125 $Y2=2.115
r89 2 24 400 $w=1.7e-07 $l=9.26971e-07 $layer=licon1_PDIFF $count=1 $X=0.975
+ $Y=1.96 $X2=1.125 $Y2=2.815
r90 1 18 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=0.63
+ $Y=0.56 $X2=0.77 $Y2=0.835
.ends

.subckt PM_SKY130_FD_SC_HS__A2BB2OI_1%B2 1 3 4 6 11 14 15
c41 14 0 8.02067e-21 $X=2.64 $Y=1.665
r42 14 15 18.5393 $w=2.28e-07 $l=3.7e-07 $layer=LI1_cond $X=2.64 $Y=1.665
+ $X2=2.64 $Y2=2.035
r43 12 14 6.26328 $w=2.28e-07 $l=1.25e-07 $layer=LI1_cond $X=2.64 $Y=1.54
+ $X2=2.64 $Y2=1.665
r44 11 12 2.67223 $w=2.3e-07 $l=1.6e-07 $layer=LI1_cond $X=2.64 $Y=1.38 $X2=2.64
+ $Y2=1.54
r45 8 11 9.18353 $w=3.18e-07 $l=2.55e-07 $layer=LI1_cond $X=2.385 $Y=1.38
+ $X2=2.64 $Y2=1.38
r46 8 9 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.385
+ $Y=1.385 $X2=2.385 $Y2=1.385
r47 4 9 77.2841 $w=2.7e-07 $l=3.87427e-07 $layer=POLY_cond $X=2.37 $Y=1.765
+ $X2=2.385 $Y2=1.385
r48 4 6 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.37 $Y=1.765
+ $X2=2.37 $Y2=2.4
r49 1 9 38.9026 $w=2.7e-07 $l=1.74714e-07 $layer=POLY_cond $X=2.365 $Y=1.22
+ $X2=2.385 $Y2=1.385
r50 1 3 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=2.365 $Y=1.22 $X2=2.365
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HS__A2BB2OI_1%B1 1 3 4 6 7
r26 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.09
+ $Y=1.385 $X2=3.09 $Y2=1.385
r27 7 11 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=3.09 $Y=1.295 $X2=3.09
+ $Y2=1.385
r28 4 10 67.0639 $w=3.7e-07 $l=4.5173e-07 $layer=POLY_cond $X=2.85 $Y=1.765
+ $X2=3.007 $Y2=1.385
r29 4 6 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.85 $Y=1.765
+ $X2=2.85 $Y2=2.4
r30 1 10 39.0558 $w=3.7e-07 $l=2.40757e-07 $layer=POLY_cond $X=2.835 $Y=1.22
+ $X2=3.007 $Y2=1.385
r31 1 3 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=2.835 $Y=1.22 $X2=2.835
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HS__A2BB2OI_1%VPWR 1 2 7 9 14 18 21 22 23 33 34
c43 18 0 1.19409e-19 $X=2.61 $Y=2.815
r44 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r45 33 34 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r46 31 34 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=3.12 $Y2=3.33
r47 30 31 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r48 28 38 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r49 27 30 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=0.72 $Y=3.33
+ $X2=2.16 $Y2=3.33
r50 27 28 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r51 25 37 4.72267 $w=1.7e-07 $l=2.25e-07 $layer=LI1_cond $X=0.45 $Y=3.33
+ $X2=0.225 $Y2=3.33
r52 25 27 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=0.45 $Y=3.33 $X2=0.72
+ $Y2=3.33
r53 23 31 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r54 23 28 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=0.72 $Y2=3.33
r55 21 30 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=2.43 $Y=3.33 $X2=2.16
+ $Y2=3.33
r56 21 22 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.43 $Y=3.33
+ $X2=2.515 $Y2=3.33
r57 20 33 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=2.6 $Y=3.33 $X2=3.12
+ $Y2=3.33
r58 20 22 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.6 $Y=3.33 $X2=2.515
+ $Y2=3.33
r59 15 18 4.37928 $w=2.48e-07 $l=9.5e-08 $layer=LI1_cond $X=2.515 $Y=2.855
+ $X2=2.61 $Y2=2.855
r60 14 22 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.515 $Y=3.245
+ $X2=2.515 $Y2=3.33
r61 13 15 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.515 $Y=2.98
+ $X2=2.515 $Y2=2.855
r62 13 14 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=2.515 $Y=2.98
+ $X2=2.515 $Y2=3.245
r63 9 12 24.4458 $w=3.28e-07 $l=7e-07 $layer=LI1_cond $X=0.285 $Y=2.115
+ $X2=0.285 $Y2=2.815
r64 7 37 3.0435 $w=3.3e-07 $l=1.11018e-07 $layer=LI1_cond $X=0.285 $Y=3.245
+ $X2=0.225 $Y2=3.33
r65 7 12 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=0.285 $Y=3.245
+ $X2=0.285 $Y2=2.815
r66 2 18 600 $w=1.7e-07 $l=1.05428e-06 $layer=licon1_PDIFF $count=1 $X=2.445
+ $Y=1.84 $X2=2.61 $Y2=2.815
r67 1 12 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=0.16
+ $Y=1.96 $X2=0.285 $Y2=2.815
r68 1 9 400 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_PDIFF $count=1 $X=0.16
+ $Y=1.96 $X2=0.285 $Y2=2.115
.ends

.subckt PM_SKY130_FD_SC_HS__A2BB2OI_1%Y 1 2 10 11 13 19 23
c46 13 0 1.45091e-19 $X=2.15 $Y=0.515
r47 23 25 7.73239 $w=4.26e-07 $l=2.7e-07 $layer=LI1_cond $X=1.695 $Y=2.082
+ $X2=1.965 $Y2=2.082
r48 19 25 5.58451 $w=4.26e-07 $l=1.95e-07 $layer=LI1_cond $X=2.16 $Y=2.082
+ $X2=1.965 $Y2=2.082
r49 11 15 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=2.185 $Y=0.965
+ $X2=1.965 $Y2=0.965
r50 11 13 16.1785 $w=2.58e-07 $l=3.65e-07 $layer=LI1_cond $X=2.185 $Y=0.88
+ $X2=2.185 $Y2=0.515
r51 10 25 6.16288 $w=1.7e-07 $l=3.32e-07 $layer=LI1_cond $X=1.965 $Y=1.75
+ $X2=1.965 $Y2=2.082
r52 9 15 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.965 $Y=1.05
+ $X2=1.965 $Y2=0.965
r53 9 10 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=1.965 $Y=1.05 $X2=1.965
+ $Y2=1.75
r54 2 23 300 $w=1.7e-07 $l=6.19354e-07 $layer=licon1_PDIFF $count=2 $X=1.57
+ $Y=1.84 $X2=1.695 $Y2=2.4
r55 2 23 600 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=1.57
+ $Y=1.84 $X2=1.695 $Y2=1.985
r56 1 13 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.01
+ $Y=0.37 $X2=2.15 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__A2BB2OI_1%A_399_368# 1 2 9 11 12 15 19 21
r28 17 21 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.115 $Y=2.56
+ $X2=3.115 $Y2=2.475
r29 17 19 11.7549 $w=2.48e-07 $l=2.55e-07 $layer=LI1_cond $X=3.115 $Y=2.56
+ $X2=3.115 $Y2=2.815
r30 13 21 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.115 $Y=2.39
+ $X2=3.115 $Y2=2.475
r31 13 15 18.6696 $w=2.48e-07 $l=4.05e-07 $layer=LI1_cond $X=3.115 $Y=2.39
+ $X2=3.115 $Y2=1.985
r32 11 21 2.76166 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.99 $Y=2.475
+ $X2=3.115 $Y2=2.475
r33 11 12 49.5829 $w=1.68e-07 $l=7.6e-07 $layer=LI1_cond $X=2.99 $Y=2.475
+ $X2=2.23 $Y2=2.475
r34 7 12 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=2.105 $Y=2.56
+ $X2=2.23 $Y2=2.475
r35 7 9 5.76222 $w=2.48e-07 $l=1.25e-07 $layer=LI1_cond $X=2.105 $Y=2.56
+ $X2=2.105 $Y2=2.685
r36 2 19 600 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=2.925
+ $Y=1.84 $X2=3.075 $Y2=2.815
r37 2 15 300 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=2 $X=2.925
+ $Y=1.84 $X2=3.075 $Y2=1.985
r38 1 9 600 $w=1.7e-07 $l=9.16938e-07 $layer=licon1_PDIFF $count=1 $X=1.995
+ $Y=1.84 $X2=2.145 $Y2=2.685
.ends

.subckt PM_SKY130_FD_SC_HS__A2BB2OI_1%VGND 1 2 3 10 12 14 16 18 20 25 39 44
r43 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r44 39 41 1.27749 $w=7.64e-07 $l=8e-08 $layer=LI1_cond $X=1.495 $Y=0.625
+ $X2=1.495 $Y2=0.705
r45 34 39 9.98037 $w=7.64e-07 $l=6.25e-07 $layer=LI1_cond $X=1.495 $Y=0
+ $X2=1.495 $Y2=0.625
r46 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r47 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r48 29 44 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r49 28 29 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r50 26 34 9.90117 $w=1.7e-07 $l=3.9e-07 $layer=LI1_cond $X=1.885 $Y=0 $X2=1.495
+ $Y2=0
r51 26 28 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=1.885 $Y=0 $X2=2.64
+ $Y2=0
r52 25 43 4.67153 $w=1.7e-07 $l=2.37e-07 $layer=LI1_cond $X=2.885 $Y=0 $X2=3.122
+ $Y2=0
r53 25 28 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=2.885 $Y=0 $X2=2.64
+ $Y2=0
r54 24 35 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r55 24 32 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r56 23 24 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r57 21 31 3.94169 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=0.425 $Y=0 $X2=0.212
+ $Y2=0
r58 21 23 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.425 $Y=0 $X2=0.72
+ $Y2=0
r59 20 34 9.90117 $w=1.7e-07 $l=3.9e-07 $layer=LI1_cond $X=1.105 $Y=0 $X2=1.495
+ $Y2=0
r60 20 23 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=1.105 $Y=0 $X2=0.72
+ $Y2=0
r61 18 29 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.64
+ $Y2=0
r62 18 35 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r63 18 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r64 14 43 3.09464 $w=3.3e-07 $l=1.15521e-07 $layer=LI1_cond $X=3.05 $Y=0.085
+ $X2=3.122 $Y2=0
r65 14 16 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=3.05 $Y=0.085
+ $X2=3.05 $Y2=0.515
r66 10 31 3.20147 $w=2.5e-07 $l=1.23386e-07 $layer=LI1_cond $X=0.3 $Y=0.085
+ $X2=0.212 $Y2=0
r67 10 12 33.6513 $w=2.48e-07 $l=7.3e-07 $layer=LI1_cond $X=0.3 $Y=0.085 $X2=0.3
+ $Y2=0.815
r68 3 16 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.91
+ $Y=0.37 $X2=3.05 $Y2=0.515
r69 2 41 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=1.06
+ $Y=0.56 $X2=1.27 $Y2=0.705
r70 2 39 182 $w=1.7e-07 $l=6.91737e-07 $layer=licon1_NDIFF $count=1 $X=1.06
+ $Y=0.56 $X2=1.72 $Y2=0.625
r71 1 12 182 $w=1.7e-07 $l=3.11288e-07 $layer=licon1_NDIFF $count=1 $X=0.215
+ $Y=0.56 $X2=0.34 $Y2=0.815
.ends

