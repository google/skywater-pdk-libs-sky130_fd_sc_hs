* File: sky130_fd_sc_hs__clkinv_4.spice
* Created: Tue Sep  1 19:58:52 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hs__clkinv_4.pex.spice"
.subckt sky130_fd_sc_hs__clkinv_4  VNB VPB A VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A	A
* VPB	VPB
* VNB	VNB
MM1000 N_Y_M1000_d N_A_M1000_g N_VGND_M1000_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.14805 AS=0.3066 PD=1.125 PS=2.3 NRD=0 NRS=19.992 M=1 R=2.8 SA=75000.7
+ SB=75002.1 A=0.063 P=1.14 MULT=1
MM1001 N_Y_M1000_d N_A_M1001_g N_VGND_M1001_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.14805 AS=0.0882 PD=1.125 PS=0.84 NRD=0 NRS=19.992 M=1 R=2.8 SA=75001.5
+ SB=75001.3 A=0.063 P=1.14 MULT=1
MM1002 N_Y_M1002_d N_A_M1002_g N_VGND_M1001_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.06405 AS=0.0882 PD=0.725 PS=0.84 NRD=0 NRS=19.992 M=1 R=2.8 SA=75002.1
+ SB=75000.7 A=0.063 P=1.14 MULT=1
MM1009 N_Y_M1002_d N_A_M1009_g N_VGND_M1009_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.06405 AS=0.1386 PD=0.725 PS=1.5 NRD=7.14 NRS=12.852 M=1 R=2.8 SA=75002.5
+ SB=75000.3 A=0.063 P=1.14 MULT=1
MM1003 N_VPWR_M1003_d N_A_M1003_g N_Y_M1003_s VPB PSHORT L=0.15 W=1.12 AD=0.3304
+ AS=0.168 PD=2.83 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667 SA=75000.2
+ SB=75002.6 A=0.168 P=2.54 MULT=1
MM1004 N_VPWR_M1004_d N_A_M1004_g N_Y_M1003_s VPB PSHORT L=0.15 W=1.12 AD=0.168
+ AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667 SA=75000.7
+ SB=75002.1 A=0.168 P=2.54 MULT=1
MM1005 N_VPWR_M1004_d N_A_M1005_g N_Y_M1005_s VPB PSHORT L=0.15 W=1.12 AD=0.168
+ AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667 SA=75001.1
+ SB=75001.7 A=0.168 P=2.54 MULT=1
MM1006 N_VPWR_M1006_d N_A_M1006_g N_Y_M1005_s VPB PSHORT L=0.15 W=1.12 AD=0.196
+ AS=0.168 PD=1.47 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667 SA=75001.6
+ SB=75001.2 A=0.168 P=2.54 MULT=1
MM1007 N_VPWR_M1006_d N_A_M1007_g N_Y_M1007_s VPB PSHORT L=0.15 W=1.12 AD=0.196
+ AS=0.168 PD=1.47 PS=1.42 NRD=10.5395 NRS=1.7533 M=1 R=7.46667 SA=75002.1
+ SB=75000.7 A=0.168 P=2.54 MULT=1
MM1008 N_VPWR_M1008_d N_A_M1008_g N_Y_M1007_s VPB PSHORT L=0.15 W=1.12 AD=0.3864
+ AS=0.168 PD=2.93 PS=1.42 NRD=10.5395 NRS=1.7533 M=1 R=7.46667 SA=75002.5
+ SB=75000.3 A=0.168 P=2.54 MULT=1
DX10_noxref VNB VPB NWDIODE A=6.9564 P=11.2
*
.include "sky130_fd_sc_hs__clkinv_4.pxi.spice"
*
.ends
*
*
