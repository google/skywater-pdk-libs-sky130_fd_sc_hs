* NGSPICE file created from sky130_fd_sc_hs__o221a_4.ext - technology: sky130A

.subckt sky130_fd_sc_hs__o221a_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
M1000 a_114_125# B2 a_297_387# VPB pshort w=1e+06u l=150000u
+  ad=9.25e+11p pd=7.85e+06u as=6.45e+11p ps=5.29e+06u
M1001 a_297_387# B2 a_114_125# VPB pshort w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1002 a_27_125# B1 a_300_125# VNB nlowvt w=640000u l=150000u
+  ad=7.904e+11p pd=7.59e+06u as=7.456e+11p ps=7.45e+06u
M1003 VPWR B1 a_297_387# VPB pshort w=1e+06u l=150000u
+  ad=2.4382e+12p pd=1.739e+07u as=0p ps=0u
M1004 VPWR A1 a_763_387# VPB pshort w=1e+06u l=150000u
+  ad=0p pd=0u as=6.75e+11p ps=5.35e+06u
M1005 VGND a_114_125# X VNB nlowvt w=740000u l=150000u
+  ad=1.2421e+12p pd=1.053e+07u as=4.181e+11p ps=4.09e+06u
M1006 VPWR a_114_125# X VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=8.176e+11p ps=5.94e+06u
M1007 a_300_125# B2 a_27_125# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 X a_114_125# VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VPWR a_114_125# X VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 X a_114_125# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 X a_114_125# VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VGND A1 a_300_125# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VGND A2 a_300_125# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_300_125# A2 VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_300_125# B1 a_27_125# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_27_125# C1 a_114_125# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=1.792e+11p ps=1.84e+06u
M1017 a_114_125# C1 a_27_125# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_300_125# A1 VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_297_387# B1 VPWR VPB pshort w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_114_125# A2 a_763_387# VPB pshort w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 X a_114_125# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_763_387# A1 VPWR VPB pshort w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_27_125# B2 a_300_125# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 a_114_125# C1 VPWR VPB pshort w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 VPWR C1 a_114_125# VPB pshort w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 a_763_387# A2 a_114_125# VPB pshort w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 VGND a_114_125# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

