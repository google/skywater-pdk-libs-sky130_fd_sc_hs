* File: sky130_fd_sc_hs__edfxtp_1.pxi.spice
* Created: Tue Sep  1 20:04:27 2020
* 
x_PM_SKY130_FD_SC_HS__EDFXTP_1%D N_D_c_269_n N_D_c_270_n N_D_M1020_g N_D_M1013_g
+ D D N_D_c_266_n N_D_c_267_n N_D_c_268_n N_D_c_273_n
+ PM_SKY130_FD_SC_HS__EDFXTP_1%D
x_PM_SKY130_FD_SC_HS__EDFXTP_1%A_159_446# N_A_159_446#_M1014_s
+ N_A_159_446#_M1012_s N_A_159_446#_c_322_n N_A_159_446#_M1003_g
+ N_A_159_446#_c_323_n N_A_159_446#_M1023_g N_A_159_446#_c_324_n
+ N_A_159_446#_c_325_n N_A_159_446#_c_312_n N_A_159_446#_c_313_n
+ N_A_159_446#_c_314_n N_A_159_446#_c_343_n N_A_159_446#_c_315_n
+ N_A_159_446#_c_316_n N_A_159_446#_c_317_n N_A_159_446#_c_329_n
+ N_A_159_446#_c_318_n N_A_159_446#_c_319_n N_A_159_446#_c_320_n
+ N_A_159_446#_c_321_n PM_SKY130_FD_SC_HS__EDFXTP_1%A_159_446#
x_PM_SKY130_FD_SC_HS__EDFXTP_1%DE N_DE_M1009_g N_DE_c_439_n N_DE_c_440_n
+ N_DE_c_441_n N_DE_c_442_n N_DE_M1014_g N_DE_c_448_n N_DE_M1012_g N_DE_c_449_n
+ N_DE_c_450_n N_DE_c_451_n N_DE_M1026_g N_DE_c_443_n DE N_DE_c_445_n
+ N_DE_c_446_n PM_SKY130_FD_SC_HS__EDFXTP_1%DE
x_PM_SKY130_FD_SC_HS__EDFXTP_1%A_533_61# N_A_533_61#_M1007_d N_A_533_61#_M1027_d
+ N_A_533_61#_M1025_g N_A_533_61#_c_540_n N_A_533_61#_c_541_n
+ N_A_533_61#_M1016_g N_A_533_61#_c_528_n N_A_533_61#_M1005_g
+ N_A_533_61#_c_529_n N_A_533_61#_c_530_n N_A_533_61#_c_542_n
+ N_A_533_61#_M1024_g N_A_533_61#_c_531_n N_A_533_61#_c_544_n
+ N_A_533_61#_c_545_n N_A_533_61#_c_546_n N_A_533_61#_c_532_n
+ N_A_533_61#_c_547_n N_A_533_61#_c_533_n N_A_533_61#_c_534_n
+ N_A_533_61#_c_535_n N_A_533_61#_c_536_n N_A_533_61#_c_537_n
+ N_A_533_61#_c_538_n N_A_533_61#_c_539_n PM_SKY130_FD_SC_HS__EDFXTP_1%A_533_61#
x_PM_SKY130_FD_SC_HS__EDFXTP_1%CLK N_CLK_M1017_g N_CLK_c_728_n N_CLK_c_733_n
+ N_CLK_M1002_g N_CLK_c_729_n CLK N_CLK_c_731_n N_CLK_c_732_n
+ PM_SKY130_FD_SC_HS__EDFXTP_1%CLK
x_PM_SKY130_FD_SC_HS__EDFXTP_1%A_958_74# N_A_958_74#_M1033_d N_A_958_74#_M1019_d
+ N_A_958_74#_c_794_n N_A_958_74#_M1000_g N_A_958_74#_c_771_n
+ N_A_958_74#_M1031_g N_A_958_74#_M1032_g N_A_958_74#_c_772_n
+ N_A_958_74#_c_796_n N_A_958_74#_M1006_g N_A_958_74#_c_773_n
+ N_A_958_74#_c_774_n N_A_958_74#_c_775_n N_A_958_74#_c_797_n
+ N_A_958_74#_c_776_n N_A_958_74#_c_777_n N_A_958_74#_c_778_n
+ N_A_958_74#_c_779_n N_A_958_74#_c_868_p N_A_958_74#_c_780_n
+ N_A_958_74#_c_781_n N_A_958_74#_c_782_n N_A_958_74#_c_783_n
+ N_A_958_74#_c_784_n N_A_958_74#_c_785_n N_A_958_74#_c_786_n
+ N_A_958_74#_c_799_n N_A_958_74#_c_800_n N_A_958_74#_c_787_n
+ N_A_958_74#_c_788_n N_A_958_74#_c_789_n N_A_958_74#_c_790_n
+ N_A_958_74#_c_791_n N_A_958_74#_c_792_n N_A_958_74#_c_793_n
+ PM_SKY130_FD_SC_HS__EDFXTP_1%A_958_74#
x_PM_SKY130_FD_SC_HS__EDFXTP_1%A_763_74# N_A_763_74#_M1017_d N_A_763_74#_M1002_d
+ N_A_763_74#_M1033_g N_A_763_74#_c_995_n N_A_763_74#_c_1009_n
+ N_A_763_74#_M1019_g N_A_763_74#_M1028_g N_A_763_74#_c_997_n
+ N_A_763_74#_c_998_n N_A_763_74#_c_1012_n N_A_763_74#_c_1013_n
+ N_A_763_74#_M1004_g N_A_763_74#_c_999_n N_A_763_74#_M1021_g
+ N_A_763_74#_M1011_g N_A_763_74#_c_1001_n N_A_763_74#_c_1002_n
+ N_A_763_74#_c_1003_n N_A_763_74#_c_1004_n N_A_763_74#_c_1005_n
+ N_A_763_74#_c_1018_n N_A_763_74#_c_1019_n N_A_763_74#_c_1006_n
+ N_A_763_74#_c_1020_n N_A_763_74#_c_1007_n N_A_763_74#_c_1022_n
+ PM_SKY130_FD_SC_HS__EDFXTP_1%A_763_74#
x_PM_SKY130_FD_SC_HS__EDFXTP_1%A_1409_64# N_A_1409_64#_M1008_d
+ N_A_1409_64#_M1015_d N_A_1409_64#_M1001_g N_A_1409_64#_c_1181_n
+ N_A_1409_64#_c_1192_n N_A_1409_64#_M1030_g N_A_1409_64#_c_1182_n
+ N_A_1409_64#_c_1194_n N_A_1409_64#_M1029_g N_A_1409_64#_M1018_g
+ N_A_1409_64#_c_1184_n N_A_1409_64#_c_1185_n N_A_1409_64#_c_1186_n
+ N_A_1409_64#_c_1187_n N_A_1409_64#_c_1195_n N_A_1409_64#_c_1188_n
+ N_A_1409_64#_c_1189_n N_A_1409_64#_c_1205_n N_A_1409_64#_c_1206_n
+ N_A_1409_64#_c_1190_n PM_SKY130_FD_SC_HS__EDFXTP_1%A_1409_64#
x_PM_SKY130_FD_SC_HS__EDFXTP_1%A_1156_90# N_A_1156_90#_M1028_d
+ N_A_1156_90#_M1000_d N_A_1156_90#_M1008_g N_A_1156_90#_c_1285_n
+ N_A_1156_90#_M1015_g N_A_1156_90#_c_1286_n N_A_1156_90#_c_1312_n
+ N_A_1156_90#_c_1290_n N_A_1156_90#_c_1291_n N_A_1156_90#_c_1292_n
+ N_A_1156_90#_c_1287_n N_A_1156_90#_c_1288_n
+ PM_SKY130_FD_SC_HS__EDFXTP_1%A_1156_90#
x_PM_SKY130_FD_SC_HS__EDFXTP_1%A_1895_74# N_A_1895_74#_M1032_d
+ N_A_1895_74#_M1021_d N_A_1895_74#_M1007_g N_A_1895_74#_c_1378_n
+ N_A_1895_74#_c_1390_n N_A_1895_74#_M1027_g N_A_1895_74#_c_1379_n
+ N_A_1895_74#_c_1380_n N_A_1895_74#_M1022_g N_A_1895_74#_c_1381_n
+ N_A_1895_74#_c_1392_n N_A_1895_74#_M1010_g N_A_1895_74#_c_1382_n
+ N_A_1895_74#_c_1383_n N_A_1895_74#_c_1384_n N_A_1895_74#_c_1451_n
+ N_A_1895_74#_c_1393_n N_A_1895_74#_c_1394_n N_A_1895_74#_c_1395_n
+ N_A_1895_74#_c_1385_n N_A_1895_74#_c_1386_n N_A_1895_74#_c_1387_n
+ N_A_1895_74#_c_1388_n PM_SKY130_FD_SC_HS__EDFXTP_1%A_1895_74#
x_PM_SKY130_FD_SC_HS__EDFXTP_1%A_27_508# N_A_27_508#_M1013_s N_A_27_508#_M1025_d
+ N_A_27_508#_M1028_s N_A_27_508#_M1020_s N_A_27_508#_M1016_d
+ N_A_27_508#_M1000_s N_A_27_508#_c_1514_n N_A_27_508#_c_1521_n
+ N_A_27_508#_c_1522_n N_A_27_508#_c_1523_n N_A_27_508#_c_1524_n
+ N_A_27_508#_c_1525_n N_A_27_508#_c_1526_n N_A_27_508#_c_1527_n
+ N_A_27_508#_c_1528_n N_A_27_508#_c_1515_n N_A_27_508#_c_1530_n
+ N_A_27_508#_c_1531_n N_A_27_508#_c_1516_n N_A_27_508#_c_1517_n
+ N_A_27_508#_c_1532_n N_A_27_508#_c_1600_n N_A_27_508#_c_1533_n
+ N_A_27_508#_c_1518_n N_A_27_508#_c_1534_n N_A_27_508#_c_1519_n
+ N_A_27_508#_c_1535_n PM_SKY130_FD_SC_HS__EDFXTP_1%A_27_508#
x_PM_SKY130_FD_SC_HS__EDFXTP_1%VPWR N_VPWR_M1003_d N_VPWR_M1012_d N_VPWR_M1002_s
+ N_VPWR_M1019_s N_VPWR_M1030_d N_VPWR_M1029_s N_VPWR_M1024_d N_VPWR_M1010_d
+ N_VPWR_c_1693_n N_VPWR_c_1694_n N_VPWR_c_1695_n N_VPWR_c_1696_n
+ N_VPWR_c_1697_n N_VPWR_c_1698_n N_VPWR_c_1699_n N_VPWR_c_1700_n
+ N_VPWR_c_1701_n N_VPWR_c_1702_n N_VPWR_c_1703_n N_VPWR_c_1704_n
+ N_VPWR_c_1705_n N_VPWR_c_1706_n N_VPWR_c_1707_n N_VPWR_c_1708_n
+ N_VPWR_c_1709_n VPWR N_VPWR_c_1710_n N_VPWR_c_1711_n N_VPWR_c_1712_n
+ N_VPWR_c_1713_n N_VPWR_c_1714_n N_VPWR_c_1715_n N_VPWR_c_1716_n
+ N_VPWR_c_1692_n PM_SKY130_FD_SC_HS__EDFXTP_1%VPWR
x_PM_SKY130_FD_SC_HS__EDFXTP_1%Q N_Q_M1022_s N_Q_M1010_s N_Q_c_1831_n
+ N_Q_c_1832_n Q Q Q Q N_Q_c_1834_n Q PM_SKY130_FD_SC_HS__EDFXTP_1%Q
x_PM_SKY130_FD_SC_HS__EDFXTP_1%VGND N_VGND_M1009_d N_VGND_M1014_d N_VGND_M1017_s
+ N_VGND_M1033_s N_VGND_M1001_d N_VGND_M1018_s N_VGND_M1005_d N_VGND_M1022_d
+ N_VGND_c_1861_n N_VGND_c_1862_n N_VGND_c_1863_n N_VGND_c_1864_n
+ N_VGND_c_1865_n N_VGND_c_1866_n N_VGND_c_1867_n N_VGND_c_1868_n
+ N_VGND_c_1869_n N_VGND_c_1870_n N_VGND_c_1871_n N_VGND_c_1872_n
+ N_VGND_c_1873_n N_VGND_c_1874_n VGND N_VGND_c_1875_n N_VGND_c_1876_n
+ N_VGND_c_1877_n N_VGND_c_1878_n N_VGND_c_1879_n N_VGND_c_1880_n
+ N_VGND_c_1881_n N_VGND_c_1882_n N_VGND_c_1883_n N_VGND_c_1884_n
+ PM_SKY130_FD_SC_HS__EDFXTP_1%VGND
cc_1 VNB N_D_M1013_g 0.025709f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=0.58
cc_2 VNB N_D_c_266_n 0.0171113f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=1.145
cc_3 VNB N_D_c_267_n 0.0117045f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=1.145
cc_4 VNB N_D_c_268_n 0.0399559f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=1.825
cc_5 VNB N_A_159_446#_M1023_g 0.0386628f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_6 VNB N_A_159_446#_c_312_n 0.00331491f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=1.99
cc_7 VNB N_A_159_446#_c_313_n 0.0273265f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=1.145
cc_8 VNB N_A_159_446#_c_314_n 0.00951957f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A_159_446#_c_315_n 0.00319209f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_159_446#_c_316_n 3.2668e-19 $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=1.665
cc_11 VNB N_A_159_446#_c_317_n 0.00674726f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_159_446#_c_318_n 0.0029594f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_159_446#_c_319_n 6.37728e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_159_446#_c_320_n 0.0037051f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_159_446#_c_321_n 0.0279463f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_DE_M1009_g 0.0227548f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.465
cc_17 VNB N_DE_c_439_n 0.0256476f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.75
cc_18 VNB N_DE_c_440_n 0.0101882f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=0.98
cc_19 VNB N_DE_c_441_n 0.0115035f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=1.145
cc_20 VNB N_DE_c_442_n 0.0166758f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=0.98
cc_21 VNB N_DE_c_443_n 0.0236907f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=1.825
cc_22 VNB DE 0.00159289f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=1.295
cc_23 VNB N_DE_c_445_n 0.0148266f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_DE_c_446_n 0.0176647f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_533_61#_M1025_g 0.0228356f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_533_61#_c_528_n 0.0182482f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=1.825
cc_27 VNB N_A_533_61#_c_529_n 0.0406862f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=1.145
cc_28 VNB N_A_533_61#_c_530_n 0.00732576f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=1.825
cc_29 VNB N_A_533_61#_c_531_n 0.0325649f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_533_61#_c_532_n 0.0108941f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_533_61#_c_533_n 0.028351f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_533_61#_c_534_n 0.00306562f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_533_61#_c_535_n 0.00462585f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_533_61#_c_536_n 0.0036769f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_533_61#_c_537_n 0.0603477f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_533_61#_c_538_n 0.010322f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_533_61#_c_539_n 0.010666f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_CLK_c_728_n 0.0114076f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.75
cc_39 VNB N_CLK_c_729_n 0.0140862f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB CLK 0.00749125f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=0.98
cc_41 VNB N_CLK_c_731_n 0.0403775f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_CLK_c_732_n 0.0204272f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=1.825
cc_43 VNB N_A_958_74#_c_771_n 0.0184494f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=1.145
cc_44 VNB N_A_958_74#_c_772_n 0.00355316f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=1.145
cc_45 VNB N_A_958_74#_c_773_n 0.00945287f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=1.99
cc_46 VNB N_A_958_74#_c_774_n 0.0195832f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_958_74#_c_775_n 0.00279267f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=1.295
cc_48 VNB N_A_958_74#_c_776_n 0.0134814f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A_958_74#_c_777_n 0.0210336f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_A_958_74#_c_778_n 0.00189334f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_A_958_74#_c_779_n 0.012232f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_A_958_74#_c_780_n 0.0177357f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_A_958_74#_c_781_n 0.00257567f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_A_958_74#_c_782_n 0.011221f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_A_958_74#_c_783_n 0.0049927f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_A_958_74#_c_784_n 0.00315025f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_A_958_74#_c_785_n 0.0115318f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_A_958_74#_c_786_n 0.00145761f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_A_958_74#_c_787_n 0.0357913f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_A_958_74#_c_788_n 0.00837626f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_A_958_74#_c_789_n 0.00984652f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_A_958_74#_c_790_n 0.0355682f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_A_958_74#_c_791_n 0.00360052f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_A_958_74#_c_792_n 0.0305607f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_A_958_74#_c_793_n 0.0188906f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_A_763_74#_M1033_g 0.039916f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=0.98
cc_67 VNB N_A_763_74#_c_995_n 0.0159104f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_68 VNB N_A_763_74#_M1028_g 0.060147f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=1.825
cc_69 VNB N_A_763_74#_c_997_n 0.044652f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=1.825
cc_70 VNB N_A_763_74#_c_998_n 0.0127683f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=1.99
cc_71 VNB N_A_763_74#_c_999_n 0.0178472f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_A_763_74#_M1011_g 0.0523977f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_A_763_74#_c_1001_n 0.00710918f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_A_763_74#_c_1002_n 0.00706889f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_A_763_74#_c_1003_n 0.00122182f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_A_763_74#_c_1004_n 0.0118574f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_A_763_74#_c_1005_n 0.0182436f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_A_763_74#_c_1006_n 0.00148024f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VNB N_A_763_74#_c_1007_n 0.00381083f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_A_1409_64#_M1001_g 0.0291657f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_81 VNB N_A_1409_64#_c_1181_n 0.00834433f $X=-0.19 $Y=-0.245 $X2=0.635
+ $Y2=1.21
cc_82 VNB N_A_1409_64#_c_1182_n 0.00468362f $X=-0.19 $Y=-0.245 $X2=0.52
+ $Y2=1.145
cc_83 VNB N_A_1409_64#_M1018_g 0.0269585f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=1.99
cc_84 VNB N_A_1409_64#_c_1184_n 0.0548296f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_85 VNB N_A_1409_64#_c_1185_n 0.013644f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=1.295
cc_86 VNB N_A_1409_64#_c_1186_n 0.00646005f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_87 VNB N_A_1409_64#_c_1187_n 0.00782438f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_88 VNB N_A_1409_64#_c_1188_n 0.00102187f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_89 VNB N_A_1409_64#_c_1189_n 0.0127351f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_90 VNB N_A_1409_64#_c_1190_n 0.0452693f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_91 VNB N_A_1156_90#_M1008_g 0.0366237f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_92 VNB N_A_1156_90#_c_1285_n 0.013567f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=0.98
cc_93 VNB N_A_1156_90#_c_1286_n 0.02004f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_94 VNB N_A_1156_90#_c_1287_n 3.83683e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_95 VNB N_A_1156_90#_c_1288_n 0.00354447f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_96 VNB N_A_1895_74#_M1007_g 0.0293184f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_97 VNB N_A_1895_74#_c_1378_n 0.0216858f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_98 VNB N_A_1895_74#_c_1379_n 0.0559245f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=1.825
cc_99 VNB N_A_1895_74#_c_1380_n 0.0215641f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=1.145
cc_100 VNB N_A_1895_74#_c_1381_n 0.0295f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=1.825
cc_101 VNB N_A_1895_74#_c_1382_n 0.0155398f $X=-0.19 $Y=-0.245 $X2=0.615
+ $Y2=1.295
cc_102 VNB N_A_1895_74#_c_1383_n 0.00329363f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_103 VNB N_A_1895_74#_c_1384_n 0.0109396f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_104 VNB N_A_1895_74#_c_1385_n 0.00243682f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_105 VNB N_A_1895_74#_c_1386_n 0.00510635f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_106 VNB N_A_1895_74#_c_1387_n 0.0384052f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_107 VNB N_A_1895_74#_c_1388_n 0.0106154f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_108 VNB N_A_27_508#_c_1514_n 0.0404044f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=1.825
cc_109 VNB N_A_27_508#_c_1515_n 0.00984382f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_110 VNB N_A_27_508#_c_1516_n 0.00828722f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_111 VNB N_A_27_508#_c_1517_n 0.0125822f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_112 VNB N_A_27_508#_c_1518_n 0.0297869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_113 VNB N_A_27_508#_c_1519_n 0.013391f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_114 VNB N_VPWR_c_1692_n 0.541827f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_115 VNB N_Q_c_1831_n 0.00764267f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_116 VNB N_Q_c_1832_n 0.0018251f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_117 VNB Q 0.00236984f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_118 VNB N_Q_c_1834_n 0.00432377f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_119 VNB N_VGND_c_1861_n 0.00867737f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_120 VNB N_VGND_c_1862_n 0.0111489f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_121 VNB N_VGND_c_1863_n 0.00989189f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_122 VNB N_VGND_c_1864_n 0.018697f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_123 VNB N_VGND_c_1865_n 0.00789365f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_124 VNB N_VGND_c_1866_n 0.00590394f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_125 VNB N_VGND_c_1867_n 0.0122168f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_126 VNB N_VGND_c_1868_n 0.0546602f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_127 VNB N_VGND_c_1869_n 0.0319647f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_128 VNB N_VGND_c_1870_n 0.00326991f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_129 VNB N_VGND_c_1871_n 0.0614466f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_130 VNB N_VGND_c_1872_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_131 VNB N_VGND_c_1873_n 0.0298174f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_132 VNB N_VGND_c_1874_n 0.00461913f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_133 VNB N_VGND_c_1875_n 0.0309056f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_134 VNB N_VGND_c_1876_n 0.0189154f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_135 VNB N_VGND_c_1877_n 0.020445f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_136 VNB N_VGND_c_1878_n 0.0328797f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_137 VNB N_VGND_c_1879_n 0.00613227f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_138 VNB N_VGND_c_1880_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_139 VNB N_VGND_c_1881_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_140 VNB N_VGND_c_1882_n 0.0444719f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_141 VNB N_VGND_c_1883_n 0.0314426f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_142 VNB N_VGND_c_1884_n 0.729984f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_143 VPB N_D_c_269_n 0.023966f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=2.375
cc_144 VPB N_D_c_270_n 0.0264927f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=2.465
cc_145 VPB N_D_c_267_n 0.00411548f $X=-0.19 $Y=1.66 $X2=0.52 $Y2=1.145
cc_146 VPB N_D_c_268_n 0.0118292f $X=-0.19 $Y=1.66 $X2=0.52 $Y2=1.825
cc_147 VPB N_D_c_273_n 0.0160786f $X=-0.19 $Y=1.66 $X2=0.52 $Y2=1.99
cc_148 VPB N_A_159_446#_c_322_n 0.017454f $X=-0.19 $Y=1.66 $X2=0.58 $Y2=0.58
cc_149 VPB N_A_159_446#_c_323_n 0.0144439f $X=-0.19 $Y=1.66 $X2=0.52 $Y2=0.98
cc_150 VPB N_A_159_446#_c_324_n 0.0263038f $X=-0.19 $Y=1.66 $X2=0.52 $Y2=1.825
cc_151 VPB N_A_159_446#_c_325_n 0.0159417f $X=-0.19 $Y=1.66 $X2=0.52 $Y2=1.145
cc_152 VPB N_A_159_446#_c_313_n 0.0119695f $X=-0.19 $Y=1.66 $X2=0.615 $Y2=1.145
cc_153 VPB N_A_159_446#_c_315_n 0.00744243f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_154 VPB N_A_159_446#_c_316_n 0.00580517f $X=-0.19 $Y=1.66 $X2=0.615 $Y2=1.665
cc_155 VPB N_A_159_446#_c_329_n 0.00731855f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_156 VPB N_A_159_446#_c_318_n 0.00185815f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_157 VPB N_A_159_446#_c_320_n 0.00251827f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_158 VPB N_A_159_446#_c_321_n 0.00894816f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_159 VPB N_DE_c_441_n 0.0177427f $X=-0.19 $Y=1.66 $X2=0.52 $Y2=1.145
cc_160 VPB N_DE_c_448_n 0.0177379f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_161 VPB N_DE_c_449_n 0.0345564f $X=-0.19 $Y=1.66 $X2=0.52 $Y2=1.145
cc_162 VPB N_DE_c_450_n 0.0272677f $X=-0.19 $Y=1.66 $X2=0.52 $Y2=1.145
cc_163 VPB N_DE_c_451_n 0.016174f $X=-0.19 $Y=1.66 $X2=0.52 $Y2=1.145
cc_164 VPB N_A_533_61#_c_540_n 0.0246199f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.21
cc_165 VPB N_A_533_61#_c_541_n 0.0241533f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_166 VPB N_A_533_61#_c_542_n 0.0540732f $X=-0.19 $Y=1.66 $X2=0.52 $Y2=1.825
cc_167 VPB N_A_533_61#_c_531_n 0.0205345f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_168 VPB N_A_533_61#_c_544_n 0.00967562f $X=-0.19 $Y=1.66 $X2=0.615 $Y2=1.295
cc_169 VPB N_A_533_61#_c_545_n 0.00854453f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_170 VPB N_A_533_61#_c_546_n 0.0100761f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_171 VPB N_A_533_61#_c_547_n 0.00356208f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_172 VPB N_A_533_61#_c_533_n 0.0654153f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_173 VPB N_A_533_61#_c_534_n 0.00294976f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_174 VPB N_A_533_61#_c_535_n 0.00262327f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_175 VPB N_A_533_61#_c_536_n 2.54227e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_176 VPB N_A_533_61#_c_537_n 0.01285f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_177 VPB N_A_533_61#_c_538_n 0.00287546f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_178 VPB N_CLK_c_733_n 0.0205746f $X=-0.19 $Y=1.66 $X2=0.58 $Y2=0.98
cc_179 VPB N_CLK_c_729_n 0.00777712f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_180 VPB N_A_958_74#_c_794_n 0.0194889f $X=-0.19 $Y=1.66 $X2=0.58 $Y2=0.58
cc_181 VPB N_A_958_74#_c_772_n 0.0368565f $X=-0.19 $Y=1.66 $X2=0.52 $Y2=1.145
cc_182 VPB N_A_958_74#_c_796_n 0.0225521f $X=-0.19 $Y=1.66 $X2=0.52 $Y2=1.145
cc_183 VPB N_A_958_74#_c_797_n 0.00210791f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_184 VPB N_A_958_74#_c_776_n 0.00159321f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_185 VPB N_A_958_74#_c_799_n 0.00862439f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_186 VPB N_A_958_74#_c_800_n 0.0595516f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_187 VPB N_A_763_74#_c_995_n 0.0162963f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_188 VPB N_A_763_74#_c_1009_n 0.020397f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_189 VPB N_A_763_74#_c_997_n 0.0271937f $X=-0.19 $Y=1.66 $X2=0.52 $Y2=1.825
cc_190 VPB N_A_763_74#_c_998_n 0.016033f $X=-0.19 $Y=1.66 $X2=0.52 $Y2=1.99
cc_191 VPB N_A_763_74#_c_1012_n 0.0165753f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_192 VPB N_A_763_74#_c_1013_n 0.0585063f $X=-0.19 $Y=1.66 $X2=0.615 $Y2=1.295
cc_193 VPB N_A_763_74#_c_999_n 0.0448045f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_194 VPB N_A_763_74#_c_1003_n 0.00340096f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_195 VPB N_A_763_74#_c_1004_n 0.00506357f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_196 VPB N_A_763_74#_c_1005_n 0.00535596f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_197 VPB N_A_763_74#_c_1018_n 0.0140888f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_198 VPB N_A_763_74#_c_1019_n 0.00340905f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_199 VPB N_A_763_74#_c_1020_n 0.00877063f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_200 VPB N_A_763_74#_c_1007_n 0.00165135f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_201 VPB N_A_763_74#_c_1022_n 0.0379962f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_202 VPB N_A_1409_64#_c_1181_n 0.041826f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.21
cc_203 VPB N_A_1409_64#_c_1192_n 0.022599f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_204 VPB N_A_1409_64#_c_1182_n 0.0110002f $X=-0.19 $Y=1.66 $X2=0.52 $Y2=1.145
cc_205 VPB N_A_1409_64#_c_1194_n 0.0301291f $X=-0.19 $Y=1.66 $X2=0.52 $Y2=1.145
cc_206 VPB N_A_1409_64#_c_1195_n 0.00522514f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_207 VPB N_A_1409_64#_c_1188_n 0.0100806f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_208 VPB N_A_1156_90#_c_1285_n 0.0444055f $X=-0.19 $Y=1.66 $X2=0.52 $Y2=0.98
cc_209 VPB N_A_1156_90#_c_1290_n 0.00333956f $X=-0.19 $Y=1.66 $X2=0.52 $Y2=1.825
cc_210 VPB N_A_1156_90#_c_1291_n 0.00723895f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_211 VPB N_A_1156_90#_c_1292_n 0.00900971f $X=-0.19 $Y=1.66 $X2=0.615
+ $Y2=1.665
cc_212 VPB N_A_1156_90#_c_1287_n 0.00167199f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_213 VPB N_A_1156_90#_c_1288_n 0.0121922f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_214 VPB N_A_1895_74#_c_1378_n 0.0308459f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.21
cc_215 VPB N_A_1895_74#_c_1390_n 0.0260142f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_216 VPB N_A_1895_74#_c_1381_n 0.00133984f $X=-0.19 $Y=1.66 $X2=0.52 $Y2=1.825
cc_217 VPB N_A_1895_74#_c_1392_n 0.0317221f $X=-0.19 $Y=1.66 $X2=0.52 $Y2=1.99
cc_218 VPB N_A_1895_74#_c_1393_n 0.00729312f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_219 VPB N_A_1895_74#_c_1394_n 0.0104845f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_220 VPB N_A_1895_74#_c_1395_n 0.00680098f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_221 VPB N_A_1895_74#_c_1385_n 0.00116664f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_222 VPB N_A_27_508#_c_1514_n 0.0244832f $X=-0.19 $Y=1.66 $X2=0.52 $Y2=1.825
cc_223 VPB N_A_27_508#_c_1521_n 0.0283234f $X=-0.19 $Y=1.66 $X2=0.52 $Y2=1.99
cc_224 VPB N_A_27_508#_c_1522_n 0.0279615f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_225 VPB N_A_27_508#_c_1523_n 0.0121061f $X=-0.19 $Y=1.66 $X2=0.615 $Y2=1.665
cc_226 VPB N_A_27_508#_c_1524_n 0.0174906f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_227 VPB N_A_27_508#_c_1525_n 0.00349119f $X=-0.19 $Y=1.66 $X2=0.615 $Y2=1.825
cc_228 VPB N_A_27_508#_c_1526_n 0.00146513f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_229 VPB N_A_27_508#_c_1527_n 0.0224096f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_230 VPB N_A_27_508#_c_1528_n 0.00113173f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_231 VPB N_A_27_508#_c_1515_n 0.00831197f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_232 VPB N_A_27_508#_c_1530_n 0.0281515f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_233 VPB N_A_27_508#_c_1531_n 0.00161431f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_234 VPB N_A_27_508#_c_1532_n 0.00892442f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_235 VPB N_A_27_508#_c_1533_n 0.00666749f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_236 VPB N_A_27_508#_c_1534_n 0.0124532f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_237 VPB N_A_27_508#_c_1535_n 0.0162464f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_238 VPB N_VPWR_c_1693_n 0.00772185f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_239 VPB N_VPWR_c_1694_n 0.0243274f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_240 VPB N_VPWR_c_1695_n 0.0240424f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_241 VPB N_VPWR_c_1696_n 0.0243657f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_242 VPB N_VPWR_c_1697_n 0.0102489f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_243 VPB N_VPWR_c_1698_n 0.0126657f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_244 VPB N_VPWR_c_1699_n 0.0113109f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_245 VPB N_VPWR_c_1700_n 0.0103331f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_246 VPB N_VPWR_c_1701_n 0.0649899f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_247 VPB N_VPWR_c_1702_n 0.0293385f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_248 VPB N_VPWR_c_1703_n 0.00460249f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_249 VPB N_VPWR_c_1704_n 0.0298174f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_250 VPB N_VPWR_c_1705_n 0.0047828f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_251 VPB N_VPWR_c_1706_n 0.0314345f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_252 VPB N_VPWR_c_1707_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_253 VPB N_VPWR_c_1708_n 0.0215854f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_254 VPB N_VPWR_c_1709_n 0.00614052f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_255 VPB N_VPWR_c_1710_n 0.0323948f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_256 VPB N_VPWR_c_1711_n 0.0590477f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_257 VPB N_VPWR_c_1712_n 0.0583199f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_258 VPB N_VPWR_c_1713_n 0.033781f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_259 VPB N_VPWR_c_1714_n 0.0047828f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_260 VPB N_VPWR_c_1715_n 0.00614976f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_261 VPB N_VPWR_c_1716_n 0.0103609f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_262 VPB N_VPWR_c_1692_n 0.194712f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_263 VPB Q 0.0151107f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_264 N_D_c_270_n N_A_159_446#_c_322_n 0.031194f $X=0.495 $Y=2.465 $X2=0 $Y2=0
cc_265 N_D_c_269_n N_A_159_446#_c_324_n 0.0150942f $X=0.495 $Y=2.375 $X2=0 $Y2=0
cc_266 N_D_c_269_n N_A_159_446#_c_325_n 0.00843883f $X=0.495 $Y=2.375 $X2=0
+ $Y2=0
cc_267 N_D_c_273_n N_A_159_446#_c_325_n 0.0137702f $X=0.52 $Y=1.99 $X2=0 $Y2=0
cc_268 N_D_M1013_g N_A_159_446#_c_312_n 2.08437e-19 $X=0.58 $Y=0.58 $X2=0 $Y2=0
cc_269 N_D_c_266_n N_A_159_446#_c_312_n 0.00142126f $X=0.52 $Y=1.145 $X2=0 $Y2=0
cc_270 N_D_c_267_n N_A_159_446#_c_312_n 0.0513743f $X=0.52 $Y=1.145 $X2=0 $Y2=0
cc_271 N_D_c_268_n N_A_159_446#_c_312_n 2.79757e-19 $X=0.52 $Y=1.825 $X2=0 $Y2=0
cc_272 N_D_c_267_n N_A_159_446#_c_313_n 0.00320031f $X=0.52 $Y=1.145 $X2=0 $Y2=0
cc_273 N_D_c_268_n N_A_159_446#_c_313_n 0.0137702f $X=0.52 $Y=1.825 $X2=0 $Y2=0
cc_274 N_D_M1013_g N_A_159_446#_c_343_n 8.2231e-19 $X=0.58 $Y=0.58 $X2=0 $Y2=0
cc_275 N_D_c_267_n N_A_159_446#_c_316_n 0.0312709f $X=0.52 $Y=1.145 $X2=0 $Y2=0
cc_276 N_D_c_268_n N_A_159_446#_c_316_n 3.92359e-19 $X=0.52 $Y=1.825 $X2=0 $Y2=0
cc_277 N_D_M1013_g N_DE_M1009_g 0.0377085f $X=0.58 $Y=0.58 $X2=0 $Y2=0
cc_278 N_D_c_266_n N_DE_c_440_n 0.00787042f $X=0.52 $Y=1.145 $X2=0 $Y2=0
cc_279 N_D_c_267_n N_DE_c_440_n 8.91711e-19 $X=0.52 $Y=1.145 $X2=0 $Y2=0
cc_280 N_D_c_269_n N_A_27_508#_c_1514_n 0.00675092f $X=0.495 $Y=2.375 $X2=0
+ $Y2=0
cc_281 N_D_M1013_g N_A_27_508#_c_1514_n 0.0053259f $X=0.58 $Y=0.58 $X2=0 $Y2=0
cc_282 N_D_c_266_n N_A_27_508#_c_1514_n 0.0245541f $X=0.52 $Y=1.145 $X2=0 $Y2=0
cc_283 N_D_c_267_n N_A_27_508#_c_1514_n 0.0766518f $X=0.52 $Y=1.145 $X2=0 $Y2=0
cc_284 N_D_c_269_n N_A_27_508#_c_1521_n 8.93269e-19 $X=0.495 $Y=2.375 $X2=0
+ $Y2=0
cc_285 N_D_c_270_n N_A_27_508#_c_1521_n 0.0149319f $X=0.495 $Y=2.465 $X2=0 $Y2=0
cc_286 N_D_c_269_n N_A_27_508#_c_1522_n 0.0128162f $X=0.495 $Y=2.375 $X2=0 $Y2=0
cc_287 N_D_c_267_n N_A_27_508#_c_1522_n 0.0270499f $X=0.52 $Y=1.145 $X2=0 $Y2=0
cc_288 N_D_c_273_n N_A_27_508#_c_1522_n 6.79407e-19 $X=0.52 $Y=1.99 $X2=0 $Y2=0
cc_289 N_D_M1013_g N_A_27_508#_c_1518_n 0.0103351f $X=0.58 $Y=0.58 $X2=0 $Y2=0
cc_290 N_D_c_266_n N_A_27_508#_c_1518_n 0.00386592f $X=0.52 $Y=1.145 $X2=0 $Y2=0
cc_291 N_D_c_267_n N_A_27_508#_c_1518_n 0.00885856f $X=0.52 $Y=1.145 $X2=0 $Y2=0
cc_292 N_D_c_269_n N_A_27_508#_c_1534_n 0.00518121f $X=0.495 $Y=2.375 $X2=0
+ $Y2=0
cc_293 N_D_c_267_n N_A_27_508#_c_1534_n 6.96185e-19 $X=0.52 $Y=1.145 $X2=0 $Y2=0
cc_294 N_D_c_273_n N_A_27_508#_c_1534_n 0.00236763f $X=0.52 $Y=1.99 $X2=0 $Y2=0
cc_295 N_D_c_270_n N_VPWR_c_1693_n 0.0018421f $X=0.495 $Y=2.465 $X2=0 $Y2=0
cc_296 N_D_c_270_n N_VPWR_c_1702_n 0.00445602f $X=0.495 $Y=2.465 $X2=0 $Y2=0
cc_297 N_D_c_270_n N_VPWR_c_1692_n 0.00899152f $X=0.495 $Y=2.465 $X2=0 $Y2=0
cc_298 N_D_M1013_g N_VGND_c_1861_n 0.00124923f $X=0.58 $Y=0.58 $X2=0 $Y2=0
cc_299 N_D_M1013_g N_VGND_c_1875_n 0.00432935f $X=0.58 $Y=0.58 $X2=0 $Y2=0
cc_300 N_D_M1013_g N_VGND_c_1884_n 0.00821075f $X=0.58 $Y=0.58 $X2=0 $Y2=0
cc_301 N_A_159_446#_c_312_n N_DE_M1009_g 3.25298e-19 $X=1.14 $Y=1.505 $X2=0
+ $Y2=0
cc_302 N_A_159_446#_c_343_n N_DE_M1009_g 0.0092911f $X=1.305 $Y=0.855 $X2=0
+ $Y2=0
cc_303 N_A_159_446#_c_317_n N_DE_M1009_g 0.00290865f $X=1.735 $Y=0.645 $X2=0
+ $Y2=0
cc_304 N_A_159_446#_c_312_n N_DE_c_439_n 0.0164959f $X=1.14 $Y=1.505 $X2=0 $Y2=0
cc_305 N_A_159_446#_c_314_n N_DE_c_439_n 0.0078387f $X=1.57 $Y=0.855 $X2=0 $Y2=0
cc_306 N_A_159_446#_c_315_n N_DE_c_439_n 0.00330448f $X=1.705 $Y=1.695 $X2=0
+ $Y2=0
cc_307 N_A_159_446#_c_312_n N_DE_c_440_n 0.00292959f $X=1.14 $Y=1.505 $X2=0
+ $Y2=0
cc_308 N_A_159_446#_c_313_n N_DE_c_440_n 0.0182201f $X=1.14 $Y=1.505 $X2=0 $Y2=0
cc_309 N_A_159_446#_c_312_n N_DE_c_441_n 9.98266e-19 $X=1.14 $Y=1.505 $X2=0
+ $Y2=0
cc_310 N_A_159_446#_c_313_n N_DE_c_441_n 0.0094379f $X=1.14 $Y=1.505 $X2=0 $Y2=0
cc_311 N_A_159_446#_c_315_n N_DE_c_441_n 0.00510837f $X=1.705 $Y=1.695 $X2=0
+ $Y2=0
cc_312 N_A_159_446#_c_316_n N_DE_c_441_n 9.01876e-19 $X=1.305 $Y=1.695 $X2=0
+ $Y2=0
cc_313 N_A_159_446#_c_329_n N_DE_c_441_n 0.00622022f $X=1.79 $Y=2.495 $X2=0
+ $Y2=0
cc_314 N_A_159_446#_c_319_n N_DE_c_441_n 0.00563344f $X=1.79 $Y=1.695 $X2=0
+ $Y2=0
cc_315 N_A_159_446#_c_320_n N_DE_c_441_n 0.00145247f $X=2.22 $Y=1.55 $X2=0 $Y2=0
cc_316 N_A_159_446#_c_321_n N_DE_c_441_n 0.0154054f $X=2.38 $Y=1.55 $X2=0 $Y2=0
cc_317 N_A_159_446#_M1023_g N_DE_c_442_n 0.0199563f $X=2.38 $Y=0.645 $X2=0 $Y2=0
cc_318 N_A_159_446#_c_312_n N_DE_c_442_n 2.20134e-19 $X=1.14 $Y=1.505 $X2=0
+ $Y2=0
cc_319 N_A_159_446#_c_314_n N_DE_c_442_n 0.00377761f $X=1.57 $Y=0.855 $X2=0
+ $Y2=0
cc_320 N_A_159_446#_c_317_n N_DE_c_442_n 7.31217e-19 $X=1.735 $Y=0.645 $X2=0
+ $Y2=0
cc_321 N_A_159_446#_c_329_n N_DE_c_448_n 0.00624167f $X=1.79 $Y=2.495 $X2=0
+ $Y2=0
cc_322 N_A_159_446#_c_323_n N_DE_c_450_n 0.00250929f $X=1.05 $Y=2.23 $X2=0 $Y2=0
cc_323 N_A_159_446#_c_325_n N_DE_c_450_n 0.0094379f $X=1.14 $Y=2.01 $X2=0 $Y2=0
cc_324 N_A_159_446#_c_329_n N_DE_c_450_n 0.0116006f $X=1.79 $Y=2.495 $X2=0 $Y2=0
cc_325 N_A_159_446#_c_318_n N_DE_c_450_n 0.00659937f $X=2.055 $Y=1.695 $X2=0
+ $Y2=0
cc_326 N_A_159_446#_c_320_n N_DE_c_450_n 0.00113317f $X=2.22 $Y=1.55 $X2=0 $Y2=0
cc_327 N_A_159_446#_c_321_n N_DE_c_450_n 0.0220693f $X=2.38 $Y=1.55 $X2=0 $Y2=0
cc_328 N_A_159_446#_c_314_n N_DE_c_443_n 0.00681326f $X=1.57 $Y=0.855 $X2=0
+ $Y2=0
cc_329 N_A_159_446#_c_318_n N_DE_c_443_n 0.00434828f $X=2.055 $Y=1.695 $X2=0
+ $Y2=0
cc_330 N_A_159_446#_c_319_n N_DE_c_443_n 0.00101655f $X=1.79 $Y=1.695 $X2=0
+ $Y2=0
cc_331 N_A_159_446#_M1023_g DE 0.00150886f $X=2.38 $Y=0.645 $X2=0 $Y2=0
cc_332 N_A_159_446#_c_312_n DE 0.0218472f $X=1.14 $Y=1.505 $X2=0 $Y2=0
cc_333 N_A_159_446#_c_313_n DE 3.48291e-19 $X=1.14 $Y=1.505 $X2=0 $Y2=0
cc_334 N_A_159_446#_c_314_n DE 0.0247809f $X=1.57 $Y=0.855 $X2=0 $Y2=0
cc_335 N_A_159_446#_c_315_n DE 0.014091f $X=1.705 $Y=1.695 $X2=0 $Y2=0
cc_336 N_A_159_446#_c_319_n DE 0.0112841f $X=1.79 $Y=1.695 $X2=0 $Y2=0
cc_337 N_A_159_446#_c_320_n DE 0.00348554f $X=2.22 $Y=1.55 $X2=0 $Y2=0
cc_338 N_A_159_446#_M1023_g N_DE_c_445_n 0.00817197f $X=2.38 $Y=0.645 $X2=0
+ $Y2=0
cc_339 N_A_159_446#_c_312_n N_DE_c_445_n 0.00546415f $X=1.14 $Y=1.505 $X2=0
+ $Y2=0
cc_340 N_A_159_446#_c_312_n N_DE_c_446_n 3.48291e-19 $X=1.14 $Y=1.505 $X2=0
+ $Y2=0
cc_341 N_A_159_446#_c_313_n N_DE_c_446_n 0.00609406f $X=1.14 $Y=1.505 $X2=0
+ $Y2=0
cc_342 N_A_159_446#_c_315_n N_DE_c_446_n 0.00104323f $X=1.705 $Y=1.695 $X2=0
+ $Y2=0
cc_343 N_A_159_446#_c_321_n N_DE_c_446_n 0.0034012f $X=2.38 $Y=1.55 $X2=0 $Y2=0
cc_344 N_A_159_446#_M1023_g N_A_533_61#_M1025_g 0.0421816f $X=2.38 $Y=0.645
+ $X2=0 $Y2=0
cc_345 N_A_159_446#_c_320_n N_A_533_61#_c_534_n 0.00774583f $X=2.22 $Y=1.55
+ $X2=0 $Y2=0
cc_346 N_A_159_446#_c_321_n N_A_533_61#_c_534_n 0.00333561f $X=2.38 $Y=1.55
+ $X2=0 $Y2=0
cc_347 N_A_159_446#_c_320_n N_A_533_61#_c_537_n 2.95947e-19 $X=2.22 $Y=1.55
+ $X2=0 $Y2=0
cc_348 N_A_159_446#_c_321_n N_A_533_61#_c_537_n 0.0421816f $X=2.38 $Y=1.55 $X2=0
+ $Y2=0
cc_349 N_A_159_446#_M1023_g N_A_533_61#_c_538_n 0.0107379f $X=2.38 $Y=0.645
+ $X2=0 $Y2=0
cc_350 N_A_159_446#_c_320_n N_A_533_61#_c_538_n 0.0285435f $X=2.22 $Y=1.55 $X2=0
+ $Y2=0
cc_351 N_A_159_446#_c_322_n N_A_27_508#_c_1521_n 0.00154959f $X=0.885 $Y=2.465
+ $X2=0 $Y2=0
cc_352 N_A_159_446#_c_324_n N_A_27_508#_c_1521_n 5.59111e-19 $X=0.885 $Y=2.347
+ $X2=0 $Y2=0
cc_353 N_A_159_446#_c_323_n N_A_27_508#_c_1522_n 0.00448415f $X=1.05 $Y=2.23
+ $X2=0 $Y2=0
cc_354 N_A_159_446#_c_324_n N_A_27_508#_c_1522_n 0.0178082f $X=0.885 $Y=2.347
+ $X2=0 $Y2=0
cc_355 N_A_159_446#_c_325_n N_A_27_508#_c_1522_n 0.00125351f $X=1.14 $Y=2.01
+ $X2=0 $Y2=0
cc_356 N_A_159_446#_c_315_n N_A_27_508#_c_1522_n 0.0103913f $X=1.705 $Y=1.695
+ $X2=0 $Y2=0
cc_357 N_A_159_446#_c_316_n N_A_27_508#_c_1522_n 0.0258112f $X=1.305 $Y=1.695
+ $X2=0 $Y2=0
cc_358 N_A_159_446#_c_329_n N_A_27_508#_c_1522_n 0.0141316f $X=1.79 $Y=2.495
+ $X2=0 $Y2=0
cc_359 N_A_159_446#_c_322_n N_A_27_508#_c_1523_n 0.00209312f $X=0.885 $Y=2.465
+ $X2=0 $Y2=0
cc_360 N_A_159_446#_c_324_n N_A_27_508#_c_1523_n 0.00338256f $X=0.885 $Y=2.347
+ $X2=0 $Y2=0
cc_361 N_A_159_446#_c_329_n N_A_27_508#_c_1523_n 0.028439f $X=1.79 $Y=2.495
+ $X2=0 $Y2=0
cc_362 N_A_159_446#_c_329_n N_A_27_508#_c_1524_n 0.0130106f $X=1.79 $Y=2.495
+ $X2=0 $Y2=0
cc_363 N_A_159_446#_c_322_n N_A_27_508#_c_1525_n 6.93242e-19 $X=0.885 $Y=2.465
+ $X2=0 $Y2=0
cc_364 N_A_159_446#_c_329_n N_A_27_508#_c_1526_n 0.0432202f $X=1.79 $Y=2.495
+ $X2=0 $Y2=0
cc_365 N_A_159_446#_c_320_n N_A_27_508#_c_1527_n 0.013613f $X=2.22 $Y=1.55 $X2=0
+ $Y2=0
cc_366 N_A_159_446#_c_321_n N_A_27_508#_c_1527_n 0.00183975f $X=2.38 $Y=1.55
+ $X2=0 $Y2=0
cc_367 N_A_159_446#_c_329_n N_A_27_508#_c_1528_n 0.013005f $X=1.79 $Y=2.495
+ $X2=0 $Y2=0
cc_368 N_A_159_446#_c_318_n N_A_27_508#_c_1528_n 8.44449e-19 $X=2.055 $Y=1.695
+ $X2=0 $Y2=0
cc_369 N_A_159_446#_c_320_n N_A_27_508#_c_1528_n 0.0143089f $X=2.22 $Y=1.55
+ $X2=0 $Y2=0
cc_370 N_A_159_446#_c_321_n N_A_27_508#_c_1528_n 5.27783e-19 $X=2.38 $Y=1.55
+ $X2=0 $Y2=0
cc_371 N_A_159_446#_c_343_n N_A_27_508#_c_1518_n 0.00145863f $X=1.305 $Y=0.855
+ $X2=0 $Y2=0
cc_372 N_A_159_446#_M1023_g N_A_27_508#_c_1519_n 0.00124492f $X=2.38 $Y=0.645
+ $X2=0 $Y2=0
cc_373 N_A_159_446#_c_322_n N_VPWR_c_1693_n 0.0132287f $X=0.885 $Y=2.465 $X2=0
+ $Y2=0
cc_374 N_A_159_446#_c_324_n N_VPWR_c_1693_n 0.00461083f $X=0.885 $Y=2.347 $X2=0
+ $Y2=0
cc_375 N_A_159_446#_c_322_n N_VPWR_c_1702_n 0.00413917f $X=0.885 $Y=2.465 $X2=0
+ $Y2=0
cc_376 N_A_159_446#_c_322_n N_VPWR_c_1692_n 0.00817239f $X=0.885 $Y=2.465 $X2=0
+ $Y2=0
cc_377 N_A_159_446#_c_324_n N_VPWR_c_1692_n 3.19707e-19 $X=0.885 $Y=2.347 $X2=0
+ $Y2=0
cc_378 N_A_159_446#_c_343_n N_VGND_M1009_d 0.00220205f $X=1.305 $Y=0.855
+ $X2=-0.19 $Y2=-0.245
cc_379 N_A_159_446#_c_314_n N_VGND_c_1861_n 0.00351808f $X=1.57 $Y=0.855 $X2=0
+ $Y2=0
cc_380 N_A_159_446#_c_343_n N_VGND_c_1861_n 0.0196647f $X=1.305 $Y=0.855 $X2=0
+ $Y2=0
cc_381 N_A_159_446#_c_317_n N_VGND_c_1861_n 0.0125975f $X=1.735 $Y=0.645 $X2=0
+ $Y2=0
cc_382 N_A_159_446#_M1023_g N_VGND_c_1862_n 0.012473f $X=2.38 $Y=0.645 $X2=0
+ $Y2=0
cc_383 N_A_159_446#_c_314_n N_VGND_c_1862_n 0.00463069f $X=1.57 $Y=0.855 $X2=0
+ $Y2=0
cc_384 N_A_159_446#_c_317_n N_VGND_c_1862_n 0.0134516f $X=1.735 $Y=0.645 $X2=0
+ $Y2=0
cc_385 N_A_159_446#_c_320_n N_VGND_c_1862_n 0.0101419f $X=2.22 $Y=1.55 $X2=0
+ $Y2=0
cc_386 N_A_159_446#_c_321_n N_VGND_c_1862_n 0.00165606f $X=2.38 $Y=1.55 $X2=0
+ $Y2=0
cc_387 N_A_159_446#_M1023_g N_VGND_c_1869_n 0.00441186f $X=2.38 $Y=0.645 $X2=0
+ $Y2=0
cc_388 N_A_159_446#_c_317_n N_VGND_c_1876_n 0.00860429f $X=1.735 $Y=0.645 $X2=0
+ $Y2=0
cc_389 N_A_159_446#_M1023_g N_VGND_c_1884_n 0.0044119f $X=2.38 $Y=0.645 $X2=0
+ $Y2=0
cc_390 N_A_159_446#_c_314_n N_VGND_c_1884_n 0.00826433f $X=1.57 $Y=0.855 $X2=0
+ $Y2=0
cc_391 N_A_159_446#_c_343_n N_VGND_c_1884_n 0.00271168f $X=1.305 $Y=0.855 $X2=0
+ $Y2=0
cc_392 N_A_159_446#_c_317_n N_VGND_c_1884_n 0.00870705f $X=1.735 $Y=0.645 $X2=0
+ $Y2=0
cc_393 N_DE_c_449_n N_A_533_61#_c_540_n 0.00970968f $X=2.62 $Y=2.03 $X2=0 $Y2=0
cc_394 N_DE_c_451_n N_A_533_61#_c_541_n 0.031582f $X=2.695 $Y=2.105 $X2=0 $Y2=0
cc_395 N_DE_c_449_n N_A_533_61#_c_537_n 0.00664698f $X=2.62 $Y=2.03 $X2=0 $Y2=0
cc_396 N_DE_c_449_n N_A_533_61#_c_538_n 0.0010711f $X=2.62 $Y=2.03 $X2=0 $Y2=0
cc_397 N_DE_c_448_n N_A_27_508#_c_1523_n 0.00341917f $X=2.015 $Y=2.105 $X2=0
+ $Y2=0
cc_398 N_DE_c_448_n N_A_27_508#_c_1524_n 0.00949792f $X=2.015 $Y=2.105 $X2=0
+ $Y2=0
cc_399 N_DE_c_448_n N_A_27_508#_c_1526_n 0.0207293f $X=2.015 $Y=2.105 $X2=0
+ $Y2=0
cc_400 N_DE_c_451_n N_A_27_508#_c_1526_n 0.00353893f $X=2.695 $Y=2.105 $X2=0
+ $Y2=0
cc_401 N_DE_c_449_n N_A_27_508#_c_1527_n 0.0176401f $X=2.62 $Y=2.03 $X2=0 $Y2=0
cc_402 N_DE_c_451_n N_A_27_508#_c_1527_n 0.00653291f $X=2.695 $Y=2.105 $X2=0
+ $Y2=0
cc_403 N_DE_c_448_n N_A_27_508#_c_1528_n 4.308e-19 $X=2.015 $Y=2.105 $X2=0 $Y2=0
cc_404 N_DE_c_449_n N_A_27_508#_c_1528_n 0.00284546f $X=2.62 $Y=2.03 $X2=0 $Y2=0
cc_405 N_DE_c_450_n N_A_27_508#_c_1528_n 0.00301735f $X=2.09 $Y=2.03 $X2=0 $Y2=0
cc_406 N_DE_M1009_g N_A_27_508#_c_1518_n 0.00168095f $X=0.97 $Y=0.58 $X2=0 $Y2=0
cc_407 N_DE_c_451_n N_A_27_508#_c_1535_n 0.00189511f $X=2.695 $Y=2.105 $X2=0
+ $Y2=0
cc_408 N_DE_c_448_n N_VPWR_c_1694_n 0.00250187f $X=2.015 $Y=2.105 $X2=0 $Y2=0
cc_409 N_DE_c_449_n N_VPWR_c_1694_n 0.00110823f $X=2.62 $Y=2.03 $X2=0 $Y2=0
cc_410 N_DE_c_451_n N_VPWR_c_1694_n 0.00921909f $X=2.695 $Y=2.105 $X2=0 $Y2=0
cc_411 N_DE_c_448_n N_VPWR_c_1704_n 7.0893e-19 $X=2.015 $Y=2.105 $X2=0 $Y2=0
cc_412 N_DE_c_451_n N_VPWR_c_1706_n 0.00326897f $X=2.695 $Y=2.105 $X2=0 $Y2=0
cc_413 N_DE_c_451_n N_VPWR_c_1692_n 0.00400166f $X=2.695 $Y=2.105 $X2=0 $Y2=0
cc_414 N_DE_M1009_g N_VGND_c_1861_n 0.00953711f $X=0.97 $Y=0.58 $X2=0 $Y2=0
cc_415 N_DE_c_439_n N_VGND_c_1861_n 9.9363e-19 $X=1.515 $Y=1.025 $X2=0 $Y2=0
cc_416 N_DE_c_442_n N_VGND_c_1861_n 0.00208085f $X=1.95 $Y=0.95 $X2=0 $Y2=0
cc_417 N_DE_c_442_n N_VGND_c_1862_n 0.0111681f $X=1.95 $Y=0.95 $X2=0 $Y2=0
cc_418 N_DE_M1009_g N_VGND_c_1875_n 0.00383152f $X=0.97 $Y=0.58 $X2=0 $Y2=0
cc_419 N_DE_c_442_n N_VGND_c_1876_n 0.00441186f $X=1.95 $Y=0.95 $X2=0 $Y2=0
cc_420 N_DE_M1009_g N_VGND_c_1884_n 0.00615424f $X=0.97 $Y=0.58 $X2=0 $Y2=0
cc_421 N_DE_c_442_n N_VGND_c_1884_n 0.0044119f $X=1.95 $Y=0.95 $X2=0 $Y2=0
cc_422 N_A_533_61#_c_533_n CLK 0.0167f $X=11.615 $Y=1.665 $X2=0 $Y2=0
cc_423 N_A_533_61#_c_537_n CLK 4.84099e-19 $X=2.83 $Y=1.21 $X2=0 $Y2=0
cc_424 N_A_533_61#_c_533_n N_CLK_c_731_n 0.00417411f $X=11.615 $Y=1.665 $X2=0
+ $Y2=0
cc_425 N_A_533_61#_c_537_n N_CLK_c_731_n 0.0150512f $X=2.83 $Y=1.21 $X2=0 $Y2=0
cc_426 N_A_533_61#_c_537_n N_CLK_c_732_n 0.00337304f $X=2.83 $Y=1.21 $X2=0 $Y2=0
cc_427 N_A_533_61#_c_542_n N_A_958_74#_c_772_n 0.0204153f $X=10.785 $Y=2.435
+ $X2=0 $Y2=0
cc_428 N_A_533_61#_c_531_n N_A_958_74#_c_772_n 0.0146467f $X=10.89 $Y=2.02 $X2=0
+ $Y2=0
cc_429 N_A_533_61#_c_544_n N_A_958_74#_c_772_n 8.23648e-19 $X=11.555 $Y=2.207
+ $X2=0 $Y2=0
cc_430 N_A_533_61#_c_533_n N_A_958_74#_c_772_n 0.00564714f $X=11.615 $Y=1.665
+ $X2=0 $Y2=0
cc_431 N_A_533_61#_c_542_n N_A_958_74#_c_796_n 0.0324155f $X=10.785 $Y=2.435
+ $X2=0 $Y2=0
cc_432 N_A_533_61#_c_533_n N_A_958_74#_c_773_n 0.00789556f $X=11.615 $Y=1.665
+ $X2=0 $Y2=0
cc_433 N_A_533_61#_c_533_n N_A_958_74#_c_797_n 0.0140605f $X=11.615 $Y=1.665
+ $X2=0 $Y2=0
cc_434 N_A_533_61#_c_533_n N_A_958_74#_c_776_n 0.0221532f $X=11.615 $Y=1.665
+ $X2=0 $Y2=0
cc_435 N_A_533_61#_c_533_n N_A_958_74#_c_779_n 0.00423047f $X=11.615 $Y=1.665
+ $X2=0 $Y2=0
cc_436 N_A_533_61#_c_533_n N_A_958_74#_c_783_n 0.00730168f $X=11.615 $Y=1.665
+ $X2=0 $Y2=0
cc_437 N_A_533_61#_c_533_n N_A_958_74#_c_784_n 7.61262e-19 $X=11.615 $Y=1.665
+ $X2=0 $Y2=0
cc_438 N_A_533_61#_c_530_n N_A_958_74#_c_785_n 0.00130497f $X=10.375 $Y=0.94
+ $X2=0 $Y2=0
cc_439 N_A_533_61#_c_533_n N_A_958_74#_c_785_n 0.015916f $X=11.615 $Y=1.665
+ $X2=0 $Y2=0
cc_440 N_A_533_61#_c_533_n N_A_958_74#_c_799_n 0.00761408f $X=11.615 $Y=1.665
+ $X2=0 $Y2=0
cc_441 N_A_533_61#_c_533_n N_A_958_74#_c_787_n 0.00190225f $X=11.615 $Y=1.665
+ $X2=0 $Y2=0
cc_442 N_A_533_61#_c_533_n N_A_958_74#_c_788_n 0.0098216f $X=11.615 $Y=1.665
+ $X2=0 $Y2=0
cc_443 N_A_533_61#_c_533_n N_A_958_74#_c_789_n 0.01903f $X=11.615 $Y=1.665 $X2=0
+ $Y2=0
cc_444 N_A_533_61#_c_533_n N_A_958_74#_c_790_n 0.00174952f $X=11.615 $Y=1.665
+ $X2=0 $Y2=0
cc_445 N_A_533_61#_c_530_n N_A_958_74#_c_791_n 0.0019999f $X=10.375 $Y=0.94
+ $X2=0 $Y2=0
cc_446 N_A_533_61#_c_531_n N_A_958_74#_c_791_n 7.22432e-19 $X=10.89 $Y=2.02
+ $X2=0 $Y2=0
cc_447 N_A_533_61#_c_533_n N_A_958_74#_c_791_n 0.00931256f $X=11.615 $Y=1.665
+ $X2=0 $Y2=0
cc_448 N_A_533_61#_c_530_n N_A_958_74#_c_792_n 0.017152f $X=10.375 $Y=0.94 $X2=0
+ $Y2=0
cc_449 N_A_533_61#_c_531_n N_A_958_74#_c_792_n 0.0205371f $X=10.89 $Y=2.02 $X2=0
+ $Y2=0
cc_450 N_A_533_61#_c_533_n N_A_763_74#_c_995_n 0.00550162f $X=11.615 $Y=1.665
+ $X2=0 $Y2=0
cc_451 N_A_533_61#_c_533_n N_A_763_74#_c_997_n 0.0172604f $X=11.615 $Y=1.665
+ $X2=0 $Y2=0
cc_452 N_A_533_61#_c_533_n N_A_763_74#_c_998_n 0.00980106f $X=11.615 $Y=1.665
+ $X2=0 $Y2=0
cc_453 N_A_533_61#_c_533_n N_A_763_74#_c_999_n 0.00811584f $X=11.615 $Y=1.665
+ $X2=0 $Y2=0
cc_454 N_A_533_61#_c_528_n N_A_763_74#_M1011_g 0.0406264f $X=10.3 $Y=0.865 $X2=0
+ $Y2=0
cc_455 N_A_533_61#_c_533_n N_A_763_74#_c_1003_n 0.0193665f $X=11.615 $Y=1.665
+ $X2=0 $Y2=0
cc_456 N_A_533_61#_c_533_n N_A_763_74#_c_1004_n 0.0523905f $X=11.615 $Y=1.665
+ $X2=0 $Y2=0
cc_457 N_A_533_61#_c_533_n N_A_763_74#_c_1019_n 0.00977116f $X=11.615 $Y=1.665
+ $X2=0 $Y2=0
cc_458 N_A_533_61#_c_533_n N_A_763_74#_c_1006_n 0.00551289f $X=11.615 $Y=1.665
+ $X2=0 $Y2=0
cc_459 N_A_533_61#_c_533_n N_A_763_74#_c_1020_n 0.00239393f $X=11.615 $Y=1.665
+ $X2=0 $Y2=0
cc_460 N_A_533_61#_c_533_n N_A_763_74#_c_1007_n 0.0217703f $X=11.615 $Y=1.665
+ $X2=0 $Y2=0
cc_461 N_A_533_61#_c_533_n N_A_1409_64#_c_1181_n 0.00192057f $X=11.615 $Y=1.665
+ $X2=0 $Y2=0
cc_462 N_A_533_61#_c_533_n N_A_1409_64#_c_1182_n 0.0116494f $X=11.615 $Y=1.665
+ $X2=0 $Y2=0
cc_463 N_A_533_61#_c_533_n N_A_1409_64#_c_1184_n 0.00379165f $X=11.615 $Y=1.665
+ $X2=0 $Y2=0
cc_464 N_A_533_61#_c_533_n N_A_1409_64#_c_1185_n 7.57862e-19 $X=11.615 $Y=1.665
+ $X2=0 $Y2=0
cc_465 N_A_533_61#_c_533_n N_A_1409_64#_c_1186_n 0.0112543f $X=11.615 $Y=1.665
+ $X2=0 $Y2=0
cc_466 N_A_533_61#_c_533_n N_A_1409_64#_c_1195_n 0.00667603f $X=11.615 $Y=1.665
+ $X2=0 $Y2=0
cc_467 N_A_533_61#_c_533_n N_A_1409_64#_c_1188_n 0.0170068f $X=11.615 $Y=1.665
+ $X2=0 $Y2=0
cc_468 N_A_533_61#_c_533_n N_A_1409_64#_c_1189_n 0.0135625f $X=11.615 $Y=1.665
+ $X2=0 $Y2=0
cc_469 N_A_533_61#_c_533_n N_A_1409_64#_c_1205_n 0.0170777f $X=11.615 $Y=1.665
+ $X2=0 $Y2=0
cc_470 N_A_533_61#_c_533_n N_A_1409_64#_c_1206_n 0.00784482f $X=11.615 $Y=1.665
+ $X2=0 $Y2=0
cc_471 N_A_533_61#_c_533_n N_A_1409_64#_c_1190_n 0.0066297f $X=11.615 $Y=1.665
+ $X2=0 $Y2=0
cc_472 N_A_533_61#_c_533_n N_A_1156_90#_c_1285_n 0.00508221f $X=11.615 $Y=1.665
+ $X2=0 $Y2=0
cc_473 N_A_533_61#_c_533_n N_A_1156_90#_c_1286_n 0.010891f $X=11.615 $Y=1.665
+ $X2=0 $Y2=0
cc_474 N_A_533_61#_c_533_n N_A_1156_90#_c_1290_n 0.0151876f $X=11.615 $Y=1.665
+ $X2=0 $Y2=0
cc_475 N_A_533_61#_c_533_n N_A_1156_90#_c_1292_n 0.00152612f $X=11.615 $Y=1.665
+ $X2=0 $Y2=0
cc_476 N_A_533_61#_c_533_n N_A_1156_90#_c_1287_n 0.0186899f $X=11.615 $Y=1.665
+ $X2=0 $Y2=0
cc_477 N_A_533_61#_c_533_n N_A_1156_90#_c_1288_n 0.0554077f $X=11.615 $Y=1.665
+ $X2=0 $Y2=0
cc_478 N_A_533_61#_c_529_n N_A_1895_74#_M1007_g 0.0054796f $X=10.815 $Y=0.94
+ $X2=0 $Y2=0
cc_479 N_A_533_61#_c_532_n N_A_1895_74#_M1007_g 0.00230527f $X=11.62 $Y=0.57
+ $X2=0 $Y2=0
cc_480 N_A_533_61#_c_539_n N_A_1895_74#_M1007_g 0.00646527f $X=11.765 $Y=1.55
+ $X2=0 $Y2=0
cc_481 N_A_533_61#_c_542_n N_A_1895_74#_c_1378_n 0.00575402f $X=10.785 $Y=2.435
+ $X2=0 $Y2=0
cc_482 N_A_533_61#_c_531_n N_A_1895_74#_c_1378_n 0.0187228f $X=10.89 $Y=2.02
+ $X2=0 $Y2=0
cc_483 N_A_533_61#_c_544_n N_A_1895_74#_c_1378_n 0.00377771f $X=11.555 $Y=2.207
+ $X2=0 $Y2=0
cc_484 N_A_533_61#_c_547_n N_A_1895_74#_c_1378_n 0.00133931f $X=11.72 $Y=2.207
+ $X2=0 $Y2=0
cc_485 N_A_533_61#_c_533_n N_A_1895_74#_c_1378_n 0.0101744f $X=11.615 $Y=1.665
+ $X2=0 $Y2=0
cc_486 N_A_533_61#_c_535_n N_A_1895_74#_c_1378_n 0.00239059f $X=11.76 $Y=1.665
+ $X2=0 $Y2=0
cc_487 N_A_533_61#_c_536_n N_A_1895_74#_c_1378_n 0.0209862f $X=11.76 $Y=1.665
+ $X2=0 $Y2=0
cc_488 N_A_533_61#_c_539_n N_A_1895_74#_c_1378_n 0.00816022f $X=11.765 $Y=1.55
+ $X2=0 $Y2=0
cc_489 N_A_533_61#_c_542_n N_A_1895_74#_c_1390_n 0.014924f $X=10.785 $Y=2.435
+ $X2=0 $Y2=0
cc_490 N_A_533_61#_c_544_n N_A_1895_74#_c_1390_n 0.011974f $X=11.555 $Y=2.207
+ $X2=0 $Y2=0
cc_491 N_A_533_61#_c_545_n N_A_1895_74#_c_1390_n 0.00904298f $X=11.72 $Y=2.435
+ $X2=0 $Y2=0
cc_492 N_A_533_61#_c_547_n N_A_1895_74#_c_1390_n 0.00407264f $X=11.72 $Y=2.207
+ $X2=0 $Y2=0
cc_493 N_A_533_61#_c_532_n N_A_1895_74#_c_1379_n 0.00332519f $X=11.62 $Y=0.57
+ $X2=0 $Y2=0
cc_494 N_A_533_61#_c_535_n N_A_1895_74#_c_1379_n 4.89582e-19 $X=11.76 $Y=1.665
+ $X2=0 $Y2=0
cc_495 N_A_533_61#_c_536_n N_A_1895_74#_c_1379_n 0.0012174f $X=11.76 $Y=1.665
+ $X2=0 $Y2=0
cc_496 N_A_533_61#_c_539_n N_A_1895_74#_c_1379_n 0.0149104f $X=11.765 $Y=1.55
+ $X2=0 $Y2=0
cc_497 N_A_533_61#_c_532_n N_A_1895_74#_c_1380_n 0.00180935f $X=11.62 $Y=0.57
+ $X2=0 $Y2=0
cc_498 N_A_533_61#_c_536_n N_A_1895_74#_c_1381_n 3.51301e-19 $X=11.76 $Y=1.665
+ $X2=0 $Y2=0
cc_499 N_A_533_61#_c_545_n N_A_1895_74#_c_1392_n 0.00101927f $X=11.72 $Y=2.435
+ $X2=0 $Y2=0
cc_500 N_A_533_61#_c_546_n N_A_1895_74#_c_1392_n 9.80733e-19 $X=11.765 $Y=2.095
+ $X2=0 $Y2=0
cc_501 N_A_533_61#_c_547_n N_A_1895_74#_c_1392_n 4.67954e-19 $X=11.72 $Y=2.207
+ $X2=0 $Y2=0
cc_502 N_A_533_61#_c_528_n N_A_1895_74#_c_1384_n 0.00454092f $X=10.3 $Y=0.865
+ $X2=0 $Y2=0
cc_503 N_A_533_61#_c_529_n N_A_1895_74#_c_1384_n 0.0155364f $X=10.815 $Y=0.94
+ $X2=0 $Y2=0
cc_504 N_A_533_61#_c_530_n N_A_1895_74#_c_1384_n 0.00422433f $X=10.375 $Y=0.94
+ $X2=0 $Y2=0
cc_505 N_A_533_61#_c_533_n N_A_1895_74#_c_1384_n 0.00541203f $X=11.615 $Y=1.665
+ $X2=0 $Y2=0
cc_506 N_A_533_61#_c_544_n N_A_1895_74#_c_1393_n 0.00884557f $X=11.555 $Y=2.207
+ $X2=0 $Y2=0
cc_507 N_A_533_61#_c_542_n N_A_1895_74#_c_1394_n 0.00417634f $X=10.785 $Y=2.435
+ $X2=0 $Y2=0
cc_508 N_A_533_61#_c_531_n N_A_1895_74#_c_1394_n 0.00941512f $X=10.89 $Y=2.02
+ $X2=0 $Y2=0
cc_509 N_A_533_61#_c_544_n N_A_1895_74#_c_1394_n 0.0202046f $X=11.555 $Y=2.207
+ $X2=0 $Y2=0
cc_510 N_A_533_61#_c_533_n N_A_1895_74#_c_1394_n 0.0147772f $X=11.615 $Y=1.665
+ $X2=0 $Y2=0
cc_511 N_A_533_61#_c_542_n N_A_1895_74#_c_1395_n 4.73647e-19 $X=10.785 $Y=2.435
+ $X2=0 $Y2=0
cc_512 N_A_533_61#_c_531_n N_A_1895_74#_c_1395_n 5.07165e-19 $X=10.89 $Y=2.02
+ $X2=0 $Y2=0
cc_513 N_A_533_61#_c_533_n N_A_1895_74#_c_1395_n 0.0124112f $X=11.615 $Y=1.665
+ $X2=0 $Y2=0
cc_514 N_A_533_61#_c_531_n N_A_1895_74#_c_1385_n 0.0132717f $X=10.89 $Y=2.02
+ $X2=0 $Y2=0
cc_515 N_A_533_61#_c_533_n N_A_1895_74#_c_1385_n 0.0215477f $X=11.615 $Y=1.665
+ $X2=0 $Y2=0
cc_516 N_A_533_61#_c_529_n N_A_1895_74#_c_1386_n 3.34269e-19 $X=10.815 $Y=0.94
+ $X2=0 $Y2=0
cc_517 N_A_533_61#_c_542_n N_A_1895_74#_c_1386_n 7.13955e-19 $X=10.785 $Y=2.435
+ $X2=0 $Y2=0
cc_518 N_A_533_61#_c_531_n N_A_1895_74#_c_1386_n 0.00376914f $X=10.89 $Y=2.02
+ $X2=0 $Y2=0
cc_519 N_A_533_61#_c_532_n N_A_1895_74#_c_1386_n 0.00103395f $X=11.62 $Y=0.57
+ $X2=0 $Y2=0
cc_520 N_A_533_61#_c_533_n N_A_1895_74#_c_1386_n 0.0230881f $X=11.615 $Y=1.665
+ $X2=0 $Y2=0
cc_521 N_A_533_61#_c_539_n N_A_1895_74#_c_1386_n 0.0256537f $X=11.765 $Y=1.55
+ $X2=0 $Y2=0
cc_522 N_A_533_61#_c_529_n N_A_1895_74#_c_1387_n 0.0213762f $X=10.815 $Y=0.94
+ $X2=0 $Y2=0
cc_523 N_A_533_61#_c_532_n N_A_1895_74#_c_1387_n 0.00396895f $X=11.62 $Y=0.57
+ $X2=0 $Y2=0
cc_524 N_A_533_61#_c_533_n N_A_1895_74#_c_1387_n 0.00552909f $X=11.615 $Y=1.665
+ $X2=0 $Y2=0
cc_525 N_A_533_61#_c_539_n N_A_1895_74#_c_1387_n 0.00465196f $X=11.765 $Y=1.55
+ $X2=0 $Y2=0
cc_526 N_A_533_61#_c_529_n N_A_1895_74#_c_1388_n 0.00859599f $X=10.815 $Y=0.94
+ $X2=0 $Y2=0
cc_527 N_A_533_61#_c_531_n N_A_1895_74#_c_1388_n 0.00762021f $X=10.89 $Y=2.02
+ $X2=0 $Y2=0
cc_528 N_A_533_61#_c_540_n N_A_27_508#_c_1527_n 0.00284577f $X=3.085 $Y=2.015
+ $X2=0 $Y2=0
cc_529 N_A_533_61#_c_541_n N_A_27_508#_c_1527_n 0.00592753f $X=3.085 $Y=2.105
+ $X2=0 $Y2=0
cc_530 N_A_533_61#_c_533_n N_A_27_508#_c_1527_n 0.00761887f $X=11.615 $Y=1.665
+ $X2=0 $Y2=0
cc_531 N_A_533_61#_c_534_n N_A_27_508#_c_1527_n 0.00466191f $X=2.785 $Y=1.665
+ $X2=0 $Y2=0
cc_532 N_A_533_61#_c_537_n N_A_27_508#_c_1527_n 0.00316757f $X=2.83 $Y=1.21
+ $X2=0 $Y2=0
cc_533 N_A_533_61#_c_538_n N_A_27_508#_c_1527_n 0.0267574f $X=2.83 $Y=1.21 $X2=0
+ $Y2=0
cc_534 N_A_533_61#_M1025_g N_A_27_508#_c_1515_n 0.00513151f $X=2.74 $Y=0.645
+ $X2=0 $Y2=0
cc_535 N_A_533_61#_c_540_n N_A_27_508#_c_1515_n 0.0122012f $X=3.085 $Y=2.015
+ $X2=0 $Y2=0
cc_536 N_A_533_61#_c_533_n N_A_27_508#_c_1515_n 0.0266392f $X=11.615 $Y=1.665
+ $X2=0 $Y2=0
cc_537 N_A_533_61#_c_534_n N_A_27_508#_c_1515_n 4.40756e-19 $X=2.785 $Y=1.665
+ $X2=0 $Y2=0
cc_538 N_A_533_61#_c_537_n N_A_27_508#_c_1515_n 0.0205144f $X=2.83 $Y=1.21 $X2=0
+ $Y2=0
cc_539 N_A_533_61#_c_538_n N_A_27_508#_c_1515_n 0.0519058f $X=2.83 $Y=1.21 $X2=0
+ $Y2=0
cc_540 N_A_533_61#_c_533_n N_A_27_508#_c_1530_n 0.0250611f $X=11.615 $Y=1.665
+ $X2=0 $Y2=0
cc_541 N_A_533_61#_c_533_n N_A_27_508#_c_1531_n 0.0133932f $X=11.615 $Y=1.665
+ $X2=0 $Y2=0
cc_542 N_A_533_61#_c_533_n N_A_27_508#_c_1516_n 0.0194929f $X=11.615 $Y=1.665
+ $X2=0 $Y2=0
cc_543 N_A_533_61#_c_533_n N_A_27_508#_c_1517_n 0.0020928f $X=11.615 $Y=1.665
+ $X2=0 $Y2=0
cc_544 N_A_533_61#_c_533_n N_A_27_508#_c_1600_n 0.00303214f $X=11.615 $Y=1.665
+ $X2=0 $Y2=0
cc_545 N_A_533_61#_M1025_g N_A_27_508#_c_1519_n 0.00946606f $X=2.74 $Y=0.645
+ $X2=0 $Y2=0
cc_546 N_A_533_61#_c_537_n N_A_27_508#_c_1519_n 0.0090921f $X=2.83 $Y=1.21 $X2=0
+ $Y2=0
cc_547 N_A_533_61#_c_538_n N_A_27_508#_c_1519_n 0.0118563f $X=2.83 $Y=1.21 $X2=0
+ $Y2=0
cc_548 N_A_533_61#_c_540_n N_A_27_508#_c_1535_n 0.00148404f $X=3.085 $Y=2.015
+ $X2=0 $Y2=0
cc_549 N_A_533_61#_c_541_n N_A_27_508#_c_1535_n 0.0157086f $X=3.085 $Y=2.105
+ $X2=0 $Y2=0
cc_550 N_A_533_61#_c_533_n N_A_27_508#_c_1535_n 0.00808113f $X=11.615 $Y=1.665
+ $X2=0 $Y2=0
cc_551 N_A_533_61#_c_544_n N_VPWR_M1024_d 0.00249823f $X=11.555 $Y=2.207 $X2=0
+ $Y2=0
cc_552 N_A_533_61#_c_541_n N_VPWR_c_1694_n 0.00144182f $X=3.085 $Y=2.105 $X2=0
+ $Y2=0
cc_553 N_A_533_61#_c_541_n N_VPWR_c_1695_n 0.00207844f $X=3.085 $Y=2.105 $X2=0
+ $Y2=0
cc_554 N_A_533_61#_c_542_n N_VPWR_c_1699_n 0.0229807f $X=10.785 $Y=2.435 $X2=0
+ $Y2=0
cc_555 N_A_533_61#_c_544_n N_VPWR_c_1699_n 0.03489f $X=11.555 $Y=2.207 $X2=0
+ $Y2=0
cc_556 N_A_533_61#_c_545_n N_VPWR_c_1699_n 0.0167986f $X=11.72 $Y=2.435 $X2=0
+ $Y2=0
cc_557 N_A_533_61#_c_541_n N_VPWR_c_1706_n 0.00333198f $X=3.085 $Y=2.105 $X2=0
+ $Y2=0
cc_558 N_A_533_61#_c_542_n N_VPWR_c_1712_n 0.0049908f $X=10.785 $Y=2.435 $X2=0
+ $Y2=0
cc_559 N_A_533_61#_c_545_n N_VPWR_c_1713_n 0.0130196f $X=11.72 $Y=2.435 $X2=0
+ $Y2=0
cc_560 N_A_533_61#_c_541_n N_VPWR_c_1692_n 0.00441359f $X=3.085 $Y=2.105 $X2=0
+ $Y2=0
cc_561 N_A_533_61#_c_542_n N_VPWR_c_1692_n 0.00486206f $X=10.785 $Y=2.435 $X2=0
+ $Y2=0
cc_562 N_A_533_61#_c_545_n N_VPWR_c_1692_n 0.0118804f $X=11.72 $Y=2.435 $X2=0
+ $Y2=0
cc_563 N_A_533_61#_c_532_n N_Q_c_1831_n 0.0319039f $X=11.62 $Y=0.57 $X2=0 $Y2=0
cc_564 N_A_533_61#_c_539_n N_Q_c_1832_n 0.0319039f $X=11.765 $Y=1.55 $X2=0 $Y2=0
cc_565 N_A_533_61#_c_545_n Q 0.0484731f $X=11.72 $Y=2.435 $X2=0 $Y2=0
cc_566 N_A_533_61#_c_546_n Q 0.0188963f $X=11.765 $Y=2.095 $X2=0 $Y2=0
cc_567 N_A_533_61#_c_547_n Q 0.0183971f $X=11.72 $Y=2.207 $X2=0 $Y2=0
cc_568 N_A_533_61#_c_535_n Q 0.00740378f $X=11.76 $Y=1.665 $X2=0 $Y2=0
cc_569 N_A_533_61#_c_536_n Q 0.0188963f $X=11.76 $Y=1.665 $X2=0 $Y2=0
cc_570 N_A_533_61#_c_539_n N_Q_c_1834_n 0.0252426f $X=11.765 $Y=1.55 $X2=0 $Y2=0
cc_571 N_A_533_61#_M1025_g N_VGND_c_1862_n 0.00180764f $X=2.74 $Y=0.645 $X2=0
+ $Y2=0
cc_572 N_A_533_61#_M1025_g N_VGND_c_1863_n 0.00309386f $X=2.74 $Y=0.645 $X2=0
+ $Y2=0
cc_573 N_A_533_61#_c_533_n N_VGND_c_1863_n 6.4869e-19 $X=11.615 $Y=1.665 $X2=0
+ $Y2=0
cc_574 N_A_533_61#_c_533_n N_VGND_c_1864_n 0.00166402f $X=11.615 $Y=1.665 $X2=0
+ $Y2=0
cc_575 N_A_533_61#_c_532_n N_VGND_c_1868_n 4.75821e-19 $X=11.62 $Y=0.57 $X2=0
+ $Y2=0
cc_576 N_A_533_61#_M1025_g N_VGND_c_1869_n 0.00506571f $X=2.74 $Y=0.645 $X2=0
+ $Y2=0
cc_577 N_A_533_61#_c_532_n N_VGND_c_1878_n 0.0165341f $X=11.62 $Y=0.57 $X2=0
+ $Y2=0
cc_578 N_A_533_61#_c_528_n N_VGND_c_1882_n 0.00383152f $X=10.3 $Y=0.865 $X2=0
+ $Y2=0
cc_579 N_A_533_61#_c_528_n N_VGND_c_1883_n 0.011715f $X=10.3 $Y=0.865 $X2=0
+ $Y2=0
cc_580 N_A_533_61#_c_529_n N_VGND_c_1883_n 0.00459991f $X=10.815 $Y=0.94 $X2=0
+ $Y2=0
cc_581 N_A_533_61#_c_532_n N_VGND_c_1883_n 0.00290096f $X=11.62 $Y=0.57 $X2=0
+ $Y2=0
cc_582 N_A_533_61#_M1025_g N_VGND_c_1884_n 0.00525227f $X=2.74 $Y=0.645 $X2=0
+ $Y2=0
cc_583 N_A_533_61#_c_528_n N_VGND_c_1884_n 0.00380989f $X=10.3 $Y=0.865 $X2=0
+ $Y2=0
cc_584 N_A_533_61#_c_532_n N_VGND_c_1884_n 0.013075f $X=11.62 $Y=0.57 $X2=0
+ $Y2=0
cc_585 N_CLK_c_729_n N_A_763_74#_M1033_g 0.00202801f $X=4.06 $Y=1.475 $X2=0
+ $Y2=0
cc_586 N_CLK_c_732_n N_A_763_74#_c_1001_n 0.0064177f $X=3.632 $Y=1.22 $X2=0
+ $Y2=0
cc_587 N_CLK_c_728_n N_A_763_74#_c_1002_n 0.00149505f $X=3.97 $Y=1.475 $X2=0
+ $Y2=0
cc_588 N_CLK_c_729_n N_A_763_74#_c_1002_n 0.0058044f $X=4.06 $Y=1.475 $X2=0
+ $Y2=0
cc_589 CLK N_A_763_74#_c_1002_n 0.0214612f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_590 N_CLK_c_732_n N_A_763_74#_c_1002_n 0.00934401f $X=3.632 $Y=1.22 $X2=0
+ $Y2=0
cc_591 N_CLK_c_728_n N_A_763_74#_c_1003_n 0.00174372f $X=3.97 $Y=1.475 $X2=0
+ $Y2=0
cc_592 N_CLK_c_733_n N_A_763_74#_c_1003_n 0.014377f $X=4.06 $Y=1.685 $X2=0 $Y2=0
cc_593 N_CLK_c_729_n N_A_763_74#_c_1003_n 0.00529254f $X=4.06 $Y=1.475 $X2=0
+ $Y2=0
cc_594 CLK N_A_763_74#_c_1003_n 0.00638598f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_595 N_CLK_c_733_n N_A_763_74#_c_1004_n 0.00194519f $X=4.06 $Y=1.685 $X2=0
+ $Y2=0
cc_596 N_CLK_c_729_n N_A_763_74#_c_1004_n 0.00560965f $X=4.06 $Y=1.475 $X2=0
+ $Y2=0
cc_597 N_CLK_c_733_n N_A_763_74#_c_1005_n 0.00653404f $X=4.06 $Y=1.685 $X2=0
+ $Y2=0
cc_598 N_CLK_c_729_n N_A_763_74#_c_1005_n 0.0055879f $X=4.06 $Y=1.475 $X2=0
+ $Y2=0
cc_599 N_CLK_c_728_n N_A_763_74#_c_1006_n 0.00326043f $X=3.97 $Y=1.475 $X2=0
+ $Y2=0
cc_600 N_CLK_c_732_n N_A_763_74#_c_1006_n 0.00239841f $X=3.632 $Y=1.22 $X2=0
+ $Y2=0
cc_601 CLK N_A_27_508#_c_1515_n 0.0268019f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_602 N_CLK_c_731_n N_A_27_508#_c_1515_n 0.00214569f $X=3.615 $Y=1.385 $X2=0
+ $Y2=0
cc_603 N_CLK_c_732_n N_A_27_508#_c_1515_n 0.00316008f $X=3.632 $Y=1.22 $X2=0
+ $Y2=0
cc_604 N_CLK_c_733_n N_A_27_508#_c_1530_n 0.0158311f $X=4.06 $Y=1.685 $X2=0
+ $Y2=0
cc_605 N_CLK_c_733_n N_A_27_508#_c_1535_n 0.00736782f $X=4.06 $Y=1.685 $X2=0
+ $Y2=0
cc_606 CLK N_A_27_508#_c_1535_n 3.50421e-19 $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_607 N_CLK_c_733_n N_VPWR_c_1695_n 0.0184362f $X=4.06 $Y=1.685 $X2=0 $Y2=0
cc_608 N_CLK_c_733_n N_VPWR_c_1710_n 0.00467292f $X=4.06 $Y=1.685 $X2=0 $Y2=0
cc_609 N_CLK_c_733_n N_VPWR_c_1692_n 0.00471987f $X=4.06 $Y=1.685 $X2=0 $Y2=0
cc_610 CLK N_VGND_c_1863_n 0.0134779f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_611 N_CLK_c_731_n N_VGND_c_1863_n 0.0011191f $X=3.615 $Y=1.385 $X2=0 $Y2=0
cc_612 N_CLK_c_732_n N_VGND_c_1863_n 0.00467989f $X=3.632 $Y=1.22 $X2=0 $Y2=0
cc_613 N_CLK_c_732_n N_VGND_c_1864_n 0.00380993f $X=3.632 $Y=1.22 $X2=0 $Y2=0
cc_614 N_CLK_c_732_n N_VGND_c_1877_n 0.00434272f $X=3.632 $Y=1.22 $X2=0 $Y2=0
cc_615 N_CLK_c_732_n N_VGND_c_1884_n 0.00830282f $X=3.632 $Y=1.22 $X2=0 $Y2=0
cc_616 N_A_958_74#_c_773_n N_A_763_74#_M1033_g 0.00978502f $X=4.93 $Y=0.515
+ $X2=0 $Y2=0
cc_617 N_A_958_74#_c_775_n N_A_763_74#_M1033_g 0.00474255f $X=5.095 $Y=0.34
+ $X2=0 $Y2=0
cc_618 N_A_958_74#_c_773_n N_A_763_74#_c_995_n 0.00592455f $X=4.93 $Y=0.515
+ $X2=0 $Y2=0
cc_619 N_A_958_74#_c_797_n N_A_763_74#_c_1009_n 0.00388708f $X=5.825 $Y=1.98
+ $X2=0 $Y2=0
cc_620 N_A_958_74#_c_776_n N_A_763_74#_c_1009_n 9.95108e-19 $X=5.91 $Y=1.82
+ $X2=0 $Y2=0
cc_621 N_A_958_74#_c_799_n N_A_763_74#_c_1009_n 0.00115889f $X=5.91 $Y=2.06
+ $X2=0 $Y2=0
cc_622 N_A_958_74#_c_800_n N_A_763_74#_c_1009_n 0.00493673f $X=6.085 $Y=2.135
+ $X2=0 $Y2=0
cc_623 N_A_958_74#_c_773_n N_A_763_74#_M1028_g 0.00475197f $X=4.93 $Y=0.515
+ $X2=0 $Y2=0
cc_624 N_A_958_74#_c_774_n N_A_763_74#_M1028_g 0.0146867f $X=5.825 $Y=0.34 $X2=0
+ $Y2=0
cc_625 N_A_958_74#_c_776_n N_A_763_74#_M1028_g 0.0248347f $X=5.91 $Y=1.82 $X2=0
+ $Y2=0
cc_626 N_A_958_74#_c_776_n N_A_763_74#_c_997_n 0.0126149f $X=5.91 $Y=1.82 $X2=0
+ $Y2=0
cc_627 N_A_958_74#_c_799_n N_A_763_74#_c_997_n 0.00108974f $X=5.91 $Y=2.06 $X2=0
+ $Y2=0
cc_628 N_A_958_74#_c_800_n N_A_763_74#_c_997_n 0.0243286f $X=6.085 $Y=2.135
+ $X2=0 $Y2=0
cc_629 N_A_958_74#_c_787_n N_A_763_74#_c_997_n 0.01534f $X=6.67 $Y=1.145 $X2=0
+ $Y2=0
cc_630 N_A_958_74#_c_788_n N_A_763_74#_c_997_n 0.00129792f $X=6.96 $Y=1.122
+ $X2=0 $Y2=0
cc_631 N_A_958_74#_c_797_n N_A_763_74#_c_998_n 0.010024f $X=5.825 $Y=1.98 $X2=0
+ $Y2=0
cc_632 N_A_958_74#_c_776_n N_A_763_74#_c_998_n 6.4931e-19 $X=5.91 $Y=1.82 $X2=0
+ $Y2=0
cc_633 N_A_958_74#_c_776_n N_A_763_74#_c_1012_n 2.32223e-19 $X=5.91 $Y=1.82
+ $X2=0 $Y2=0
cc_634 N_A_958_74#_c_800_n N_A_763_74#_c_1012_n 0.0037154f $X=6.085 $Y=2.135
+ $X2=0 $Y2=0
cc_635 N_A_958_74#_c_794_n N_A_763_74#_c_1013_n 0.0101282f $X=6.385 $Y=2.465
+ $X2=0 $Y2=0
cc_636 N_A_958_74#_c_800_n N_A_763_74#_c_1013_n 0.0170478f $X=6.085 $Y=2.135
+ $X2=0 $Y2=0
cc_637 N_A_958_74#_c_772_n N_A_763_74#_c_999_n 0.010824f $X=10.365 $Y=2.345
+ $X2=0 $Y2=0
cc_638 N_A_958_74#_c_796_n N_A_763_74#_c_999_n 0.00887659f $X=10.365 $Y=2.435
+ $X2=0 $Y2=0
cc_639 N_A_958_74#_c_785_n N_A_763_74#_c_999_n 0.00476967f $X=10.275 $Y=1.29
+ $X2=0 $Y2=0
cc_640 N_A_958_74#_c_789_n N_A_763_74#_c_999_n 4.65488e-19 $X=9.285 $Y=1.29
+ $X2=0 $Y2=0
cc_641 N_A_958_74#_c_790_n N_A_763_74#_c_999_n 0.00547187f $X=9.36 $Y=1.385
+ $X2=0 $Y2=0
cc_642 N_A_958_74#_c_791_n N_A_763_74#_c_999_n 5.91559e-19 $X=10.44 $Y=1.29
+ $X2=0 $Y2=0
cc_643 N_A_958_74#_c_792_n N_A_763_74#_c_999_n 0.0217713f $X=10.44 $Y=1.42 $X2=0
+ $Y2=0
cc_644 N_A_958_74#_c_785_n N_A_763_74#_M1011_g 0.011158f $X=10.275 $Y=1.29 $X2=0
+ $Y2=0
cc_645 N_A_958_74#_c_789_n N_A_763_74#_M1011_g 5.09316e-19 $X=9.285 $Y=1.29
+ $X2=0 $Y2=0
cc_646 N_A_958_74#_c_790_n N_A_763_74#_M1011_g 0.0102681f $X=9.36 $Y=1.385 $X2=0
+ $Y2=0
cc_647 N_A_958_74#_c_791_n N_A_763_74#_M1011_g 8.46596e-19 $X=10.44 $Y=1.29
+ $X2=0 $Y2=0
cc_648 N_A_958_74#_c_792_n N_A_763_74#_M1011_g 0.00953531f $X=10.44 $Y=1.42
+ $X2=0 $Y2=0
cc_649 N_A_958_74#_c_793_n N_A_763_74#_M1011_g 0.0190284f $X=9.36 $Y=1.22 $X2=0
+ $Y2=0
cc_650 N_A_958_74#_c_773_n N_A_763_74#_c_1004_n 0.00591734f $X=4.93 $Y=0.515
+ $X2=0 $Y2=0
cc_651 N_A_958_74#_c_773_n N_A_763_74#_c_1005_n 0.00264098f $X=4.93 $Y=0.515
+ $X2=0 $Y2=0
cc_652 N_A_958_74#_c_772_n N_A_763_74#_c_1019_n 4.30958e-19 $X=10.365 $Y=2.345
+ $X2=0 $Y2=0
cc_653 N_A_958_74#_c_785_n N_A_763_74#_c_1007_n 0.0283969f $X=10.275 $Y=1.29
+ $X2=0 $Y2=0
cc_654 N_A_958_74#_c_791_n N_A_763_74#_c_1007_n 0.00253545f $X=10.44 $Y=1.29
+ $X2=0 $Y2=0
cc_655 N_A_958_74#_c_792_n N_A_763_74#_c_1007_n 0.00164371f $X=10.44 $Y=1.42
+ $X2=0 $Y2=0
cc_656 N_A_958_74#_c_771_n N_A_1409_64#_M1001_g 0.0218463f $X=6.67 $Y=0.98 $X2=0
+ $Y2=0
cc_657 N_A_958_74#_c_777_n N_A_1409_64#_M1001_g 9.04159e-19 $X=6.79 $Y=0.34
+ $X2=0 $Y2=0
cc_658 N_A_958_74#_c_778_n N_A_1409_64#_M1001_g 0.00456962f $X=6.875 $Y=0.935
+ $X2=0 $Y2=0
cc_659 N_A_958_74#_c_779_n N_A_1409_64#_M1001_g 0.0155025f $X=7.59 $Y=1.02 $X2=0
+ $Y2=0
cc_660 N_A_958_74#_c_868_p N_A_1409_64#_M1001_g 0.00183812f $X=7.675 $Y=0.935
+ $X2=0 $Y2=0
cc_661 N_A_958_74#_c_781_n N_A_1409_64#_M1001_g 2.95155e-19 $X=7.76 $Y=0.34
+ $X2=0 $Y2=0
cc_662 N_A_958_74#_c_787_n N_A_1409_64#_M1001_g 0.0205478f $X=6.67 $Y=1.145
+ $X2=0 $Y2=0
cc_663 N_A_958_74#_c_788_n N_A_1409_64#_M1001_g 0.00490258f $X=6.96 $Y=1.122
+ $X2=0 $Y2=0
cc_664 N_A_958_74#_c_780_n N_A_1409_64#_M1018_g 6.63977e-19 $X=8.27 $Y=0.34
+ $X2=0 $Y2=0
cc_665 N_A_958_74#_c_782_n N_A_1409_64#_M1018_g 0.00510095f $X=8.355 $Y=0.935
+ $X2=0 $Y2=0
cc_666 N_A_958_74#_c_783_n N_A_1409_64#_M1018_g 0.0165155f $X=9.11 $Y=1.02 $X2=0
+ $Y2=0
cc_667 N_A_958_74#_c_789_n N_A_1409_64#_M1018_g 0.00621114f $X=9.285 $Y=1.29
+ $X2=0 $Y2=0
cc_668 N_A_958_74#_c_790_n N_A_1409_64#_M1018_g 0.0213033f $X=9.36 $Y=1.385
+ $X2=0 $Y2=0
cc_669 N_A_958_74#_c_793_n N_A_1409_64#_M1018_g 0.0321202f $X=9.36 $Y=1.22 $X2=0
+ $Y2=0
cc_670 N_A_958_74#_c_783_n N_A_1409_64#_c_1184_n 0.00881339f $X=9.11 $Y=1.02
+ $X2=0 $Y2=0
cc_671 N_A_958_74#_c_784_n N_A_1409_64#_c_1184_n 0.00134551f $X=8.44 $Y=1.02
+ $X2=0 $Y2=0
cc_672 N_A_958_74#_c_779_n N_A_1409_64#_c_1186_n 0.0135045f $X=7.59 $Y=1.02
+ $X2=0 $Y2=0
cc_673 N_A_958_74#_c_779_n N_A_1409_64#_c_1187_n 0.00769005f $X=7.59 $Y=1.02
+ $X2=0 $Y2=0
cc_674 N_A_958_74#_c_780_n N_A_1409_64#_c_1187_n 0.012971f $X=8.27 $Y=0.34 $X2=0
+ $Y2=0
cc_675 N_A_958_74#_c_782_n N_A_1409_64#_c_1187_n 0.0251105f $X=8.355 $Y=0.935
+ $X2=0 $Y2=0
cc_676 N_A_958_74#_c_784_n N_A_1409_64#_c_1187_n 0.0141515f $X=8.44 $Y=1.02
+ $X2=0 $Y2=0
cc_677 N_A_958_74#_c_784_n N_A_1409_64#_c_1189_n 0.0145877f $X=8.44 $Y=1.02
+ $X2=0 $Y2=0
cc_678 N_A_958_74#_c_783_n N_A_1409_64#_c_1205_n 0.0334569f $X=9.11 $Y=1.02
+ $X2=0 $Y2=0
cc_679 N_A_958_74#_c_789_n N_A_1409_64#_c_1205_n 0.0236381f $X=9.285 $Y=1.29
+ $X2=0 $Y2=0
cc_680 N_A_958_74#_c_790_n N_A_1409_64#_c_1205_n 2.66003e-19 $X=9.36 $Y=1.385
+ $X2=0 $Y2=0
cc_681 N_A_958_74#_c_779_n N_A_1409_64#_c_1206_n 0.0319684f $X=7.59 $Y=1.02
+ $X2=0 $Y2=0
cc_682 N_A_958_74#_c_788_n N_A_1409_64#_c_1206_n 0.0028512f $X=6.96 $Y=1.122
+ $X2=0 $Y2=0
cc_683 N_A_958_74#_c_779_n N_A_1409_64#_c_1190_n 0.00726198f $X=7.59 $Y=1.02
+ $X2=0 $Y2=0
cc_684 N_A_958_74#_c_776_n N_A_1156_90#_M1028_d 0.00768863f $X=5.91 $Y=1.82
+ $X2=-0.19 $Y2=-0.245
cc_685 N_A_958_74#_c_779_n N_A_1156_90#_M1008_g 0.00553873f $X=7.59 $Y=1.02
+ $X2=0 $Y2=0
cc_686 N_A_958_74#_c_868_p N_A_1156_90#_M1008_g 0.0131174f $X=7.675 $Y=0.935
+ $X2=0 $Y2=0
cc_687 N_A_958_74#_c_780_n N_A_1156_90#_M1008_g 0.0103073f $X=8.27 $Y=0.34 $X2=0
+ $Y2=0
cc_688 N_A_958_74#_c_781_n N_A_1156_90#_M1008_g 0.00210537f $X=7.76 $Y=0.34
+ $X2=0 $Y2=0
cc_689 N_A_958_74#_c_782_n N_A_1156_90#_M1008_g 0.00339873f $X=8.355 $Y=0.935
+ $X2=0 $Y2=0
cc_690 N_A_958_74#_c_771_n N_A_1156_90#_c_1286_n 0.00363252f $X=6.67 $Y=0.98
+ $X2=0 $Y2=0
cc_691 N_A_958_74#_c_776_n N_A_1156_90#_c_1286_n 0.06434f $X=5.91 $Y=1.82 $X2=0
+ $Y2=0
cc_692 N_A_958_74#_c_778_n N_A_1156_90#_c_1286_n 0.00426874f $X=6.875 $Y=0.935
+ $X2=0 $Y2=0
cc_693 N_A_958_74#_c_787_n N_A_1156_90#_c_1286_n 0.00231928f $X=6.67 $Y=1.145
+ $X2=0 $Y2=0
cc_694 N_A_958_74#_c_788_n N_A_1156_90#_c_1286_n 0.0294985f $X=6.96 $Y=1.122
+ $X2=0 $Y2=0
cc_695 N_A_958_74#_c_771_n N_A_1156_90#_c_1312_n 0.00607399f $X=6.67 $Y=0.98
+ $X2=0 $Y2=0
cc_696 N_A_958_74#_c_776_n N_A_1156_90#_c_1312_n 0.0133947f $X=5.91 $Y=1.82
+ $X2=0 $Y2=0
cc_697 N_A_958_74#_c_777_n N_A_1156_90#_c_1312_n 0.0310197f $X=6.79 $Y=0.34
+ $X2=0 $Y2=0
cc_698 N_A_958_74#_c_787_n N_A_1156_90#_c_1312_n 4.46549e-19 $X=6.67 $Y=1.145
+ $X2=0 $Y2=0
cc_699 N_A_958_74#_c_788_n N_A_1156_90#_c_1312_n 0.00682255f $X=6.96 $Y=1.122
+ $X2=0 $Y2=0
cc_700 N_A_958_74#_c_776_n N_A_1156_90#_c_1290_n 0.0122725f $X=5.91 $Y=1.82
+ $X2=0 $Y2=0
cc_701 N_A_958_74#_c_799_n N_A_1156_90#_c_1290_n 0.00555219f $X=5.91 $Y=2.06
+ $X2=0 $Y2=0
cc_702 N_A_958_74#_c_800_n N_A_1156_90#_c_1290_n 0.00349883f $X=6.085 $Y=2.135
+ $X2=0 $Y2=0
cc_703 N_A_958_74#_c_787_n N_A_1156_90#_c_1290_n 0.00149648f $X=6.67 $Y=1.145
+ $X2=0 $Y2=0
cc_704 N_A_958_74#_c_788_n N_A_1156_90#_c_1290_n 0.0145923f $X=6.96 $Y=1.122
+ $X2=0 $Y2=0
cc_705 N_A_958_74#_c_794_n N_A_1156_90#_c_1291_n 0.00682633f $X=6.385 $Y=2.465
+ $X2=0 $Y2=0
cc_706 N_A_958_74#_c_794_n N_A_1156_90#_c_1292_n 0.00260822f $X=6.385 $Y=2.465
+ $X2=0 $Y2=0
cc_707 N_A_958_74#_c_776_n N_A_1156_90#_c_1292_n 7.8612e-19 $X=5.91 $Y=1.82
+ $X2=0 $Y2=0
cc_708 N_A_958_74#_c_799_n N_A_1156_90#_c_1292_n 0.0319585f $X=5.91 $Y=2.06
+ $X2=0 $Y2=0
cc_709 N_A_958_74#_c_800_n N_A_1156_90#_c_1292_n 0.0143546f $X=6.085 $Y=2.135
+ $X2=0 $Y2=0
cc_710 N_A_958_74#_c_779_n N_A_1156_90#_c_1288_n 0.00326485f $X=7.59 $Y=1.02
+ $X2=0 $Y2=0
cc_711 N_A_958_74#_c_793_n N_A_1895_74#_c_1383_n 0.00968523f $X=9.36 $Y=1.22
+ $X2=0 $Y2=0
cc_712 N_A_958_74#_c_785_n N_A_1895_74#_c_1384_n 0.0306291f $X=10.275 $Y=1.29
+ $X2=0 $Y2=0
cc_713 N_A_958_74#_c_791_n N_A_1895_74#_c_1384_n 0.021501f $X=10.44 $Y=1.29
+ $X2=0 $Y2=0
cc_714 N_A_958_74#_c_792_n N_A_1895_74#_c_1384_n 3.74086e-19 $X=10.44 $Y=1.42
+ $X2=0 $Y2=0
cc_715 N_A_958_74#_c_785_n N_A_1895_74#_c_1451_n 0.020247f $X=10.275 $Y=1.29
+ $X2=0 $Y2=0
cc_716 N_A_958_74#_c_789_n N_A_1895_74#_c_1451_n 6.75349e-19 $X=9.285 $Y=1.29
+ $X2=0 $Y2=0
cc_717 N_A_958_74#_c_793_n N_A_1895_74#_c_1451_n 0.00314181f $X=9.36 $Y=1.22
+ $X2=0 $Y2=0
cc_718 N_A_958_74#_c_772_n N_A_1895_74#_c_1393_n 0.00594809f $X=10.365 $Y=2.345
+ $X2=0 $Y2=0
cc_719 N_A_958_74#_c_796_n N_A_1895_74#_c_1393_n 0.00915762f $X=10.365 $Y=2.435
+ $X2=0 $Y2=0
cc_720 N_A_958_74#_c_772_n N_A_1895_74#_c_1394_n 0.00593412f $X=10.365 $Y=2.345
+ $X2=0 $Y2=0
cc_721 N_A_958_74#_c_791_n N_A_1895_74#_c_1394_n 0.0116227f $X=10.44 $Y=1.29
+ $X2=0 $Y2=0
cc_722 N_A_958_74#_c_792_n N_A_1895_74#_c_1394_n 0.00105037f $X=10.44 $Y=1.42
+ $X2=0 $Y2=0
cc_723 N_A_958_74#_c_772_n N_A_1895_74#_c_1395_n 0.0176301f $X=10.365 $Y=2.345
+ $X2=0 $Y2=0
cc_724 N_A_958_74#_c_785_n N_A_1895_74#_c_1395_n 0.00357633f $X=10.275 $Y=1.29
+ $X2=0 $Y2=0
cc_725 N_A_958_74#_c_791_n N_A_1895_74#_c_1395_n 0.00771291f $X=10.44 $Y=1.29
+ $X2=0 $Y2=0
cc_726 N_A_958_74#_c_772_n N_A_1895_74#_c_1385_n 0.00231398f $X=10.365 $Y=2.345
+ $X2=0 $Y2=0
cc_727 N_A_958_74#_c_791_n N_A_1895_74#_c_1385_n 0.0187515f $X=10.44 $Y=1.29
+ $X2=0 $Y2=0
cc_728 N_A_958_74#_c_792_n N_A_1895_74#_c_1385_n 0.00131611f $X=10.44 $Y=1.42
+ $X2=0 $Y2=0
cc_729 N_A_958_74#_c_791_n N_A_1895_74#_c_1388_n 0.0111691f $X=10.44 $Y=1.29
+ $X2=0 $Y2=0
cc_730 N_A_958_74#_c_792_n N_A_1895_74#_c_1388_n 4.90605e-19 $X=10.44 $Y=1.42
+ $X2=0 $Y2=0
cc_731 N_A_958_74#_c_797_n N_A_27_508#_c_1531_n 0.0138333f $X=5.825 $Y=1.98
+ $X2=0 $Y2=0
cc_732 N_A_958_74#_c_776_n N_A_27_508#_c_1531_n 0.00412304f $X=5.91 $Y=1.82
+ $X2=0 $Y2=0
cc_733 N_A_958_74#_c_797_n N_A_27_508#_c_1516_n 0.0119639f $X=5.825 $Y=1.98
+ $X2=0 $Y2=0
cc_734 N_A_958_74#_c_776_n N_A_27_508#_c_1516_n 0.0123714f $X=5.91 $Y=1.82 $X2=0
+ $Y2=0
cc_735 N_A_958_74#_c_773_n N_A_27_508#_c_1517_n 0.0360689f $X=4.93 $Y=0.515
+ $X2=0 $Y2=0
cc_736 N_A_958_74#_c_774_n N_A_27_508#_c_1517_n 0.0229863f $X=5.825 $Y=0.34
+ $X2=0 $Y2=0
cc_737 N_A_958_74#_c_776_n N_A_27_508#_c_1517_n 0.0561201f $X=5.91 $Y=1.82 $X2=0
+ $Y2=0
cc_738 N_A_958_74#_M1019_d N_A_27_508#_c_1532_n 0.00581991f $X=5.485 $Y=1.84
+ $X2=0 $Y2=0
cc_739 N_A_958_74#_c_794_n N_A_27_508#_c_1532_n 0.00130627f $X=6.385 $Y=2.465
+ $X2=0 $Y2=0
cc_740 N_A_958_74#_c_797_n N_A_27_508#_c_1532_n 0.00923409f $X=5.825 $Y=1.98
+ $X2=0 $Y2=0
cc_741 N_A_958_74#_c_799_n N_A_27_508#_c_1532_n 0.0284908f $X=5.91 $Y=2.06 $X2=0
+ $Y2=0
cc_742 N_A_958_74#_c_800_n N_A_27_508#_c_1532_n 0.00233063f $X=6.085 $Y=2.135
+ $X2=0 $Y2=0
cc_743 N_A_958_74#_M1019_d N_A_27_508#_c_1600_n 0.00621451f $X=5.485 $Y=1.84
+ $X2=0 $Y2=0
cc_744 N_A_958_74#_c_794_n N_A_27_508#_c_1600_n 0.00114433f $X=6.385 $Y=2.465
+ $X2=0 $Y2=0
cc_745 N_A_958_74#_c_797_n N_A_27_508#_c_1600_n 0.00645106f $X=5.825 $Y=1.98
+ $X2=0 $Y2=0
cc_746 N_A_958_74#_c_800_n N_A_27_508#_c_1600_n 0.0038162f $X=6.085 $Y=2.135
+ $X2=0 $Y2=0
cc_747 N_A_958_74#_c_794_n N_A_27_508#_c_1533_n 0.00152236f $X=6.385 $Y=2.465
+ $X2=0 $Y2=0
cc_748 N_A_958_74#_c_796_n N_VPWR_c_1699_n 0.00169994f $X=10.365 $Y=2.435 $X2=0
+ $Y2=0
cc_749 N_A_958_74#_c_794_n N_VPWR_c_1711_n 0.00411612f $X=6.385 $Y=2.465 $X2=0
+ $Y2=0
cc_750 N_A_958_74#_c_796_n N_VPWR_c_1712_n 0.0055601f $X=10.365 $Y=2.435 $X2=0
+ $Y2=0
cc_751 N_A_958_74#_c_794_n N_VPWR_c_1692_n 0.00753176f $X=6.385 $Y=2.465 $X2=0
+ $Y2=0
cc_752 N_A_958_74#_c_796_n N_VPWR_c_1692_n 0.00536257f $X=10.365 $Y=2.435 $X2=0
+ $Y2=0
cc_753 N_A_958_74#_c_800_n N_VPWR_c_1692_n 3.33135e-19 $X=6.085 $Y=2.135 $X2=0
+ $Y2=0
cc_754 N_A_958_74#_c_779_n N_VGND_M1001_d 0.00494641f $X=7.59 $Y=1.02 $X2=0
+ $Y2=0
cc_755 N_A_958_74#_c_868_p N_VGND_M1001_d 0.00544252f $X=7.675 $Y=0.935 $X2=0
+ $Y2=0
cc_756 N_A_958_74#_c_783_n N_VGND_M1018_s 0.0068916f $X=9.11 $Y=1.02 $X2=0 $Y2=0
cc_757 N_A_958_74#_c_773_n N_VGND_c_1864_n 0.0259603f $X=4.93 $Y=0.515 $X2=0
+ $Y2=0
cc_758 N_A_958_74#_c_775_n N_VGND_c_1864_n 0.0112234f $X=5.095 $Y=0.34 $X2=0
+ $Y2=0
cc_759 N_A_958_74#_c_777_n N_VGND_c_1865_n 0.0122752f $X=6.79 $Y=0.34 $X2=0
+ $Y2=0
cc_760 N_A_958_74#_c_778_n N_VGND_c_1865_n 0.0208855f $X=6.875 $Y=0.935 $X2=0
+ $Y2=0
cc_761 N_A_958_74#_c_779_n N_VGND_c_1865_n 0.0177503f $X=7.59 $Y=1.02 $X2=0
+ $Y2=0
cc_762 N_A_958_74#_c_868_p N_VGND_c_1865_n 0.025461f $X=7.675 $Y=0.935 $X2=0
+ $Y2=0
cc_763 N_A_958_74#_c_781_n N_VGND_c_1865_n 0.014745f $X=7.76 $Y=0.34 $X2=0 $Y2=0
cc_764 N_A_958_74#_c_780_n N_VGND_c_1866_n 0.0146661f $X=8.27 $Y=0.34 $X2=0
+ $Y2=0
cc_765 N_A_958_74#_c_782_n N_VGND_c_1866_n 0.0258447f $X=8.355 $Y=0.935 $X2=0
+ $Y2=0
cc_766 N_A_958_74#_c_783_n N_VGND_c_1866_n 0.0154151f $X=9.11 $Y=1.02 $X2=0
+ $Y2=0
cc_767 N_A_958_74#_c_793_n N_VGND_c_1866_n 0.00180636f $X=9.36 $Y=1.22 $X2=0
+ $Y2=0
cc_768 N_A_958_74#_c_771_n N_VGND_c_1871_n 8.05596e-19 $X=6.67 $Y=0.98 $X2=0
+ $Y2=0
cc_769 N_A_958_74#_c_774_n N_VGND_c_1871_n 0.0469671f $X=5.825 $Y=0.34 $X2=0
+ $Y2=0
cc_770 N_A_958_74#_c_775_n N_VGND_c_1871_n 0.0235688f $X=5.095 $Y=0.34 $X2=0
+ $Y2=0
cc_771 N_A_958_74#_c_777_n N_VGND_c_1871_n 0.063341f $X=6.79 $Y=0.34 $X2=0 $Y2=0
cc_772 N_A_958_74#_c_786_n N_VGND_c_1871_n 0.0121867f $X=5.91 $Y=0.34 $X2=0
+ $Y2=0
cc_773 N_A_958_74#_c_780_n N_VGND_c_1873_n 0.0449818f $X=8.27 $Y=0.34 $X2=0
+ $Y2=0
cc_774 N_A_958_74#_c_781_n N_VGND_c_1873_n 0.0121867f $X=7.76 $Y=0.34 $X2=0
+ $Y2=0
cc_775 N_A_958_74#_c_793_n N_VGND_c_1882_n 0.00434272f $X=9.36 $Y=1.22 $X2=0
+ $Y2=0
cc_776 N_A_958_74#_c_774_n N_VGND_c_1884_n 0.0274384f $X=5.825 $Y=0.34 $X2=0
+ $Y2=0
cc_777 N_A_958_74#_c_775_n N_VGND_c_1884_n 0.0127152f $X=5.095 $Y=0.34 $X2=0
+ $Y2=0
cc_778 N_A_958_74#_c_777_n N_VGND_c_1884_n 0.0364914f $X=6.79 $Y=0.34 $X2=0
+ $Y2=0
cc_779 N_A_958_74#_c_780_n N_VGND_c_1884_n 0.025776f $X=8.27 $Y=0.34 $X2=0 $Y2=0
cc_780 N_A_958_74#_c_781_n N_VGND_c_1884_n 0.00660921f $X=7.76 $Y=0.34 $X2=0
+ $Y2=0
cc_781 N_A_958_74#_c_786_n N_VGND_c_1884_n 0.00660921f $X=5.91 $Y=0.34 $X2=0
+ $Y2=0
cc_782 N_A_958_74#_c_793_n N_VGND_c_1884_n 0.00822691f $X=9.36 $Y=1.22 $X2=0
+ $Y2=0
cc_783 N_A_958_74#_c_778_n A_1349_90# 0.00579581f $X=6.875 $Y=0.935 $X2=-0.19
+ $Y2=-0.245
cc_784 N_A_958_74#_c_783_n A_1797_74# 0.00378025f $X=9.11 $Y=1.02 $X2=-0.19
+ $Y2=-0.245
cc_785 N_A_958_74#_c_789_n A_1797_74# 0.00761182f $X=9.285 $Y=1.29 $X2=-0.19
+ $Y2=-0.245
cc_786 N_A_763_74#_c_1018_n N_A_1409_64#_M1015_d 0.00826597f $X=9.63 $Y=2.495
+ $X2=0 $Y2=0
cc_787 N_A_763_74#_c_997_n N_A_1409_64#_c_1181_n 0.0125636f $X=6.685 $Y=1.655
+ $X2=0 $Y2=0
cc_788 N_A_763_74#_c_1013_n N_A_1409_64#_c_1181_n 0.0238077f $X=6.835 $Y=2.465
+ $X2=0 $Y2=0
cc_789 N_A_763_74#_c_1020_n N_A_1409_64#_c_1181_n 0.00981344f $X=6.875 $Y=2.165
+ $X2=0 $Y2=0
cc_790 N_A_763_74#_c_1013_n N_A_1409_64#_c_1192_n 0.0204155f $X=6.835 $Y=2.465
+ $X2=0 $Y2=0
cc_791 N_A_763_74#_c_1018_n N_A_1409_64#_c_1192_n 0.0161215f $X=9.63 $Y=2.495
+ $X2=0 $Y2=0
cc_792 N_A_763_74#_c_1019_n N_A_1409_64#_c_1182_n 0.00331754f $X=9.715 $Y=2.41
+ $X2=0 $Y2=0
cc_793 N_A_763_74#_c_1018_n N_A_1409_64#_c_1194_n 0.0206687f $X=9.63 $Y=2.495
+ $X2=0 $Y2=0
cc_794 N_A_763_74#_c_1019_n N_A_1409_64#_c_1194_n 0.0108219f $X=9.715 $Y=2.41
+ $X2=0 $Y2=0
cc_795 N_A_763_74#_c_1007_n N_A_1409_64#_c_1185_n 0.00294553f $X=9.9 $Y=1.635
+ $X2=0 $Y2=0
cc_796 N_A_763_74#_c_1018_n N_A_1409_64#_c_1195_n 0.0336264f $X=9.63 $Y=2.495
+ $X2=0 $Y2=0
cc_797 N_A_763_74#_c_1018_n N_A_1156_90#_c_1285_n 0.0180488f $X=9.63 $Y=2.495
+ $X2=0 $Y2=0
cc_798 N_A_763_74#_c_997_n N_A_1156_90#_c_1286_n 0.00673678f $X=6.685 $Y=1.655
+ $X2=0 $Y2=0
cc_799 N_A_763_74#_c_997_n N_A_1156_90#_c_1290_n 0.0119426f $X=6.685 $Y=1.655
+ $X2=0 $Y2=0
cc_800 N_A_763_74#_c_1013_n N_A_1156_90#_c_1291_n 0.0126906f $X=6.835 $Y=2.465
+ $X2=0 $Y2=0
cc_801 N_A_763_74#_c_1020_n N_A_1156_90#_c_1291_n 0.00455051f $X=6.875 $Y=2.165
+ $X2=0 $Y2=0
cc_802 N_A_763_74#_c_997_n N_A_1156_90#_c_1292_n 0.00102203f $X=6.685 $Y=1.655
+ $X2=0 $Y2=0
cc_803 N_A_763_74#_c_1012_n N_A_1156_90#_c_1292_n 0.00950617f $X=6.76 $Y=2 $X2=0
+ $Y2=0
cc_804 N_A_763_74#_c_1013_n N_A_1156_90#_c_1292_n 0.00147297f $X=6.835 $Y=2.465
+ $X2=0 $Y2=0
cc_805 N_A_763_74#_c_1020_n N_A_1156_90#_c_1292_n 0.0341447f $X=6.875 $Y=2.165
+ $X2=0 $Y2=0
cc_806 N_A_763_74#_c_1018_n N_A_1156_90#_c_1287_n 0.00556244f $X=9.63 $Y=2.495
+ $X2=0 $Y2=0
cc_807 N_A_763_74#_c_997_n N_A_1156_90#_c_1288_n 0.00664733f $X=6.685 $Y=1.655
+ $X2=0 $Y2=0
cc_808 N_A_763_74#_c_1012_n N_A_1156_90#_c_1288_n 0.00770657f $X=6.76 $Y=2 $X2=0
+ $Y2=0
cc_809 N_A_763_74#_c_1013_n N_A_1156_90#_c_1288_n 0.0013887f $X=6.835 $Y=2.465
+ $X2=0 $Y2=0
cc_810 N_A_763_74#_c_1018_n N_A_1156_90#_c_1288_n 0.0165064f $X=9.63 $Y=2.495
+ $X2=0 $Y2=0
cc_811 N_A_763_74#_c_1020_n N_A_1156_90#_c_1288_n 0.0220457f $X=6.875 $Y=2.165
+ $X2=0 $Y2=0
cc_812 N_A_763_74#_M1011_g N_A_1895_74#_c_1383_n 0.00369459f $X=9.91 $Y=0.58
+ $X2=0 $Y2=0
cc_813 N_A_763_74#_M1011_g N_A_1895_74#_c_1384_n 0.0121459f $X=9.91 $Y=0.58
+ $X2=0 $Y2=0
cc_814 N_A_763_74#_c_999_n N_A_1895_74#_c_1393_n 0.0105775f $X=9.83 $Y=1.885
+ $X2=0 $Y2=0
cc_815 N_A_763_74#_c_1018_n N_A_1895_74#_c_1393_n 0.0137304f $X=9.63 $Y=2.495
+ $X2=0 $Y2=0
cc_816 N_A_763_74#_c_1019_n N_A_1895_74#_c_1393_n 0.0227221f $X=9.715 $Y=2.41
+ $X2=0 $Y2=0
cc_817 N_A_763_74#_c_999_n N_A_1895_74#_c_1395_n 0.00472833f $X=9.83 $Y=1.885
+ $X2=0 $Y2=0
cc_818 N_A_763_74#_c_1019_n N_A_1895_74#_c_1395_n 0.0198165f $X=9.715 $Y=2.41
+ $X2=0 $Y2=0
cc_819 N_A_763_74#_c_1007_n N_A_1895_74#_c_1395_n 0.0056188f $X=9.9 $Y=1.635
+ $X2=0 $Y2=0
cc_820 N_A_763_74#_M1002_d N_A_27_508#_c_1530_n 0.0075824f $X=4.135 $Y=1.76
+ $X2=0 $Y2=0
cc_821 N_A_763_74#_c_995_n N_A_27_508#_c_1530_n 0.00408844f $X=5.32 $Y=1.655
+ $X2=0 $Y2=0
cc_822 N_A_763_74#_c_1003_n N_A_27_508#_c_1530_n 0.0100413f $X=4.12 $Y=1.805
+ $X2=0 $Y2=0
cc_823 N_A_763_74#_c_1004_n N_A_27_508#_c_1530_n 0.0569398f $X=4.735 $Y=1.635
+ $X2=0 $Y2=0
cc_824 N_A_763_74#_c_1022_n N_A_27_508#_c_1530_n 0.00862812f $X=4.735 $Y=1.655
+ $X2=0 $Y2=0
cc_825 N_A_763_74#_c_995_n N_A_27_508#_c_1531_n 0.00757173f $X=5.32 $Y=1.655
+ $X2=0 $Y2=0
cc_826 N_A_763_74#_c_1009_n N_A_27_508#_c_1531_n 0.00620601f $X=5.41 $Y=1.765
+ $X2=0 $Y2=0
cc_827 N_A_763_74#_c_998_n N_A_27_508#_c_1531_n 4.98583e-19 $X=5.78 $Y=1.655
+ $X2=0 $Y2=0
cc_828 N_A_763_74#_c_1004_n N_A_27_508#_c_1531_n 0.0292713f $X=4.735 $Y=1.635
+ $X2=0 $Y2=0
cc_829 N_A_763_74#_c_1022_n N_A_27_508#_c_1531_n 0.00150053f $X=4.735 $Y=1.655
+ $X2=0 $Y2=0
cc_830 N_A_763_74#_c_995_n N_A_27_508#_c_1516_n 0.00531088f $X=5.32 $Y=1.655
+ $X2=0 $Y2=0
cc_831 N_A_763_74#_M1028_g N_A_27_508#_c_1516_n 0.00334012f $X=5.705 $Y=0.66
+ $X2=0 $Y2=0
cc_832 N_A_763_74#_c_998_n N_A_27_508#_c_1516_n 0.0113819f $X=5.78 $Y=1.655
+ $X2=0 $Y2=0
cc_833 N_A_763_74#_c_1004_n N_A_27_508#_c_1516_n 0.0104131f $X=4.735 $Y=1.635
+ $X2=0 $Y2=0
cc_834 N_A_763_74#_c_1005_n N_A_27_508#_c_1516_n 7.30496e-19 $X=4.735 $Y=1.635
+ $X2=0 $Y2=0
cc_835 N_A_763_74#_M1033_g N_A_27_508#_c_1517_n 0.00970544f $X=4.715 $Y=0.74
+ $X2=0 $Y2=0
cc_836 N_A_763_74#_M1028_g N_A_27_508#_c_1517_n 0.0222528f $X=5.705 $Y=0.66
+ $X2=0 $Y2=0
cc_837 N_A_763_74#_c_998_n N_A_27_508#_c_1517_n 0.00199723f $X=5.78 $Y=1.655
+ $X2=0 $Y2=0
cc_838 N_A_763_74#_c_1004_n N_A_27_508#_c_1517_n 3.79465e-19 $X=4.735 $Y=1.635
+ $X2=0 $Y2=0
cc_839 N_A_763_74#_c_1009_n N_A_27_508#_c_1600_n 0.02998f $X=5.41 $Y=1.765 $X2=0
+ $Y2=0
cc_840 N_A_763_74#_c_1009_n N_A_27_508#_c_1533_n 0.0072676f $X=5.41 $Y=1.765
+ $X2=0 $Y2=0
cc_841 N_A_763_74#_c_1018_n N_VPWR_M1030_d 0.00720873f $X=9.63 $Y=2.495 $X2=0
+ $Y2=0
cc_842 N_A_763_74#_c_1018_n N_VPWR_M1029_s 0.012625f $X=9.63 $Y=2.495 $X2=0
+ $Y2=0
cc_843 N_A_763_74#_c_1009_n N_VPWR_c_1696_n 0.0110465f $X=5.41 $Y=1.765 $X2=0
+ $Y2=0
cc_844 N_A_763_74#_c_1013_n N_VPWR_c_1697_n 0.00120039f $X=6.835 $Y=2.465 $X2=0
+ $Y2=0
cc_845 N_A_763_74#_c_1018_n N_VPWR_c_1697_n 0.0212695f $X=9.63 $Y=2.495 $X2=0
+ $Y2=0
cc_846 N_A_763_74#_c_1018_n N_VPWR_c_1698_n 0.0212764f $X=9.63 $Y=2.495 $X2=0
+ $Y2=0
cc_847 N_A_763_74#_c_1018_n N_VPWR_c_1708_n 0.00979113f $X=9.63 $Y=2.495 $X2=0
+ $Y2=0
cc_848 N_A_763_74#_c_1009_n N_VPWR_c_1711_n 0.00421014f $X=5.41 $Y=1.765 $X2=0
+ $Y2=0
cc_849 N_A_763_74#_c_1013_n N_VPWR_c_1711_n 0.00445602f $X=6.835 $Y=2.465 $X2=0
+ $Y2=0
cc_850 N_A_763_74#_c_1018_n N_VPWR_c_1711_n 0.00351679f $X=9.63 $Y=2.495 $X2=0
+ $Y2=0
cc_851 N_A_763_74#_c_1020_n N_VPWR_c_1711_n 0.00239222f $X=6.875 $Y=2.165 $X2=0
+ $Y2=0
cc_852 N_A_763_74#_c_999_n N_VPWR_c_1712_n 0.00424414f $X=9.83 $Y=1.885 $X2=0
+ $Y2=0
cc_853 N_A_763_74#_c_1018_n N_VPWR_c_1712_n 0.0124686f $X=9.63 $Y=2.495 $X2=0
+ $Y2=0
cc_854 N_A_763_74#_c_1009_n N_VPWR_c_1692_n 0.00460416f $X=5.41 $Y=1.765 $X2=0
+ $Y2=0
cc_855 N_A_763_74#_c_1013_n N_VPWR_c_1692_n 0.00894287f $X=6.835 $Y=2.465 $X2=0
+ $Y2=0
cc_856 N_A_763_74#_c_999_n N_VPWR_c_1692_n 0.00779072f $X=9.83 $Y=1.885 $X2=0
+ $Y2=0
cc_857 N_A_763_74#_c_1018_n N_VPWR_c_1692_n 0.0539395f $X=9.63 $Y=2.495 $X2=0
+ $Y2=0
cc_858 N_A_763_74#_c_1020_n N_VPWR_c_1692_n 0.00470026f $X=6.875 $Y=2.165 $X2=0
+ $Y2=0
cc_859 N_A_763_74#_c_1018_n A_1382_508# 0.00180683f $X=9.63 $Y=2.495 $X2=-0.19
+ $Y2=-0.245
cc_860 N_A_763_74#_c_1020_n A_1382_508# 0.00326318f $X=6.875 $Y=2.165 $X2=-0.19
+ $Y2=-0.245
cc_861 N_A_763_74#_c_1018_n A_1794_392# 0.0401264f $X=9.63 $Y=2.495 $X2=-0.19
+ $Y2=-0.245
cc_862 N_A_763_74#_c_1019_n A_1794_392# 0.00789352f $X=9.715 $Y=2.41 $X2=-0.19
+ $Y2=-0.245
cc_863 N_A_763_74#_c_1001_n N_VGND_c_1863_n 0.024306f $X=3.955 $Y=0.515 $X2=0
+ $Y2=0
cc_864 N_A_763_74#_M1033_g N_VGND_c_1864_n 0.00473533f $X=4.715 $Y=0.74 $X2=0
+ $Y2=0
cc_865 N_A_763_74#_c_1001_n N_VGND_c_1864_n 0.0534949f $X=3.955 $Y=0.515 $X2=0
+ $Y2=0
cc_866 N_A_763_74#_c_1004_n N_VGND_c_1864_n 0.0122043f $X=4.735 $Y=1.635 $X2=0
+ $Y2=0
cc_867 N_A_763_74#_c_1005_n N_VGND_c_1864_n 3.36125e-19 $X=4.735 $Y=1.635 $X2=0
+ $Y2=0
cc_868 N_A_763_74#_M1033_g N_VGND_c_1871_n 0.00430908f $X=4.715 $Y=0.74 $X2=0
+ $Y2=0
cc_869 N_A_763_74#_M1028_g N_VGND_c_1871_n 8.05596e-19 $X=5.705 $Y=0.66 $X2=0
+ $Y2=0
cc_870 N_A_763_74#_c_1001_n N_VGND_c_1877_n 0.0145488f $X=3.955 $Y=0.515 $X2=0
+ $Y2=0
cc_871 N_A_763_74#_M1011_g N_VGND_c_1882_n 0.00461464f $X=9.91 $Y=0.58 $X2=0
+ $Y2=0
cc_872 N_A_763_74#_M1011_g N_VGND_c_1883_n 0.00147769f $X=9.91 $Y=0.58 $X2=0
+ $Y2=0
cc_873 N_A_763_74#_M1033_g N_VGND_c_1884_n 0.0082568f $X=4.715 $Y=0.74 $X2=0
+ $Y2=0
cc_874 N_A_763_74#_M1011_g N_VGND_c_1884_n 0.00463846f $X=9.91 $Y=0.58 $X2=0
+ $Y2=0
cc_875 N_A_763_74#_c_1001_n N_VGND_c_1884_n 0.0119924f $X=3.955 $Y=0.515 $X2=0
+ $Y2=0
cc_876 N_A_1409_64#_M1001_g N_A_1156_90#_M1008_g 0.0132329f $X=7.12 $Y=0.66
+ $X2=0 $Y2=0
cc_877 N_A_1409_64#_c_1184_n N_A_1156_90#_M1008_g 0.00723897f $X=8.805 $Y=1.44
+ $X2=0 $Y2=0
cc_878 N_A_1409_64#_c_1186_n N_A_1156_90#_M1008_g 0.0143234f $X=7.93 $Y=1.36
+ $X2=0 $Y2=0
cc_879 N_A_1409_64#_c_1187_n N_A_1156_90#_M1008_g 0.00891563f $X=8.015 $Y=0.85
+ $X2=0 $Y2=0
cc_880 N_A_1409_64#_c_1189_n N_A_1156_90#_M1008_g 5.12204e-19 $X=8.44 $Y=1.44
+ $X2=0 $Y2=0
cc_881 N_A_1409_64#_c_1190_n N_A_1156_90#_M1008_g 0.0169447f $X=7.34 $Y=1.365
+ $X2=0 $Y2=0
cc_882 N_A_1409_64#_c_1181_n N_A_1156_90#_c_1285_n 0.0372188f $X=7.34 $Y=2.375
+ $X2=0 $Y2=0
cc_883 N_A_1409_64#_c_1192_n N_A_1156_90#_c_1285_n 0.0105777f $X=7.34 $Y=2.465
+ $X2=0 $Y2=0
cc_884 N_A_1409_64#_c_1184_n N_A_1156_90#_c_1285_n 0.0037983f $X=8.805 $Y=1.44
+ $X2=0 $Y2=0
cc_885 N_A_1409_64#_c_1186_n N_A_1156_90#_c_1285_n 0.00220559f $X=7.93 $Y=1.36
+ $X2=0 $Y2=0
cc_886 N_A_1409_64#_c_1195_n N_A_1156_90#_c_1285_n 0.00487808f $X=8.27 $Y=2.155
+ $X2=0 $Y2=0
cc_887 N_A_1409_64#_c_1188_n N_A_1156_90#_c_1285_n 0.008291f $X=8.355 $Y=2.07
+ $X2=0 $Y2=0
cc_888 N_A_1409_64#_c_1189_n N_A_1156_90#_c_1285_n 0.00324239f $X=8.44 $Y=1.44
+ $X2=0 $Y2=0
cc_889 N_A_1409_64#_c_1192_n N_A_1156_90#_c_1291_n 0.00153047f $X=7.34 $Y=2.465
+ $X2=0 $Y2=0
cc_890 N_A_1409_64#_c_1181_n N_A_1156_90#_c_1287_n 3.28132e-19 $X=7.34 $Y=2.375
+ $X2=0 $Y2=0
cc_891 N_A_1409_64#_c_1186_n N_A_1156_90#_c_1287_n 0.0139504f $X=7.93 $Y=1.36
+ $X2=0 $Y2=0
cc_892 N_A_1409_64#_c_1195_n N_A_1156_90#_c_1287_n 0.00282923f $X=8.27 $Y=2.155
+ $X2=0 $Y2=0
cc_893 N_A_1409_64#_c_1188_n N_A_1156_90#_c_1287_n 0.0113679f $X=8.355 $Y=2.07
+ $X2=0 $Y2=0
cc_894 N_A_1409_64#_c_1189_n N_A_1156_90#_c_1287_n 0.00702578f $X=8.44 $Y=1.44
+ $X2=0 $Y2=0
cc_895 N_A_1409_64#_c_1181_n N_A_1156_90#_c_1288_n 0.0137102f $X=7.34 $Y=2.375
+ $X2=0 $Y2=0
cc_896 N_A_1409_64#_c_1186_n N_A_1156_90#_c_1288_n 0.0143302f $X=7.93 $Y=1.36
+ $X2=0 $Y2=0
cc_897 N_A_1409_64#_c_1206_n N_A_1156_90#_c_1288_n 0.0201775f $X=7.46 $Y=1.367
+ $X2=0 $Y2=0
cc_898 N_A_1409_64#_c_1190_n N_A_1156_90#_c_1288_n 0.00655078f $X=7.34 $Y=1.365
+ $X2=0 $Y2=0
cc_899 N_A_1409_64#_M1018_g N_A_1895_74#_c_1383_n 0.00159894f $X=8.91 $Y=0.74
+ $X2=0 $Y2=0
cc_900 N_A_1409_64#_M1018_g N_A_1895_74#_c_1451_n 5.21752e-19 $X=8.91 $Y=0.74
+ $X2=0 $Y2=0
cc_901 N_A_1409_64#_c_1192_n N_VPWR_c_1697_n 0.0085563f $X=7.34 $Y=2.465 $X2=0
+ $Y2=0
cc_902 N_A_1409_64#_c_1194_n N_VPWR_c_1698_n 0.0174616f $X=8.895 $Y=1.885 $X2=0
+ $Y2=0
cc_903 N_A_1409_64#_c_1192_n N_VPWR_c_1711_n 0.00326216f $X=7.34 $Y=2.465 $X2=0
+ $Y2=0
cc_904 N_A_1409_64#_c_1194_n N_VPWR_c_1712_n 0.00303678f $X=8.895 $Y=1.885 $X2=0
+ $Y2=0
cc_905 N_A_1409_64#_c_1192_n N_VPWR_c_1692_n 0.004235f $X=7.34 $Y=2.465 $X2=0
+ $Y2=0
cc_906 N_A_1409_64#_c_1194_n N_VPWR_c_1692_n 0.00398906f $X=8.895 $Y=1.885 $X2=0
+ $Y2=0
cc_907 N_A_1409_64#_M1001_g N_VGND_c_1865_n 0.00752223f $X=7.12 $Y=0.66 $X2=0
+ $Y2=0
cc_908 N_A_1409_64#_M1018_g N_VGND_c_1866_n 0.0133979f $X=8.91 $Y=0.74 $X2=0
+ $Y2=0
cc_909 N_A_1409_64#_M1001_g N_VGND_c_1871_n 0.00432588f $X=7.12 $Y=0.66 $X2=0
+ $Y2=0
cc_910 N_A_1409_64#_M1018_g N_VGND_c_1882_n 0.00383152f $X=8.91 $Y=0.74 $X2=0
+ $Y2=0
cc_911 N_A_1409_64#_M1001_g N_VGND_c_1884_n 0.00437282f $X=7.12 $Y=0.66 $X2=0
+ $Y2=0
cc_912 N_A_1409_64#_M1018_g N_VGND_c_1884_n 0.00758168f $X=8.91 $Y=0.74 $X2=0
+ $Y2=0
cc_913 N_A_1156_90#_c_1291_n N_A_27_508#_c_1532_n 0.0141592f $X=6.61 $Y=2.75
+ $X2=0 $Y2=0
cc_914 N_A_1156_90#_c_1291_n N_A_27_508#_c_1533_n 0.0221746f $X=6.61 $Y=2.75
+ $X2=0 $Y2=0
cc_915 N_A_1156_90#_c_1285_n N_VPWR_c_1697_n 0.00686287f $X=7.885 $Y=1.95 $X2=0
+ $Y2=0
cc_916 N_A_1156_90#_c_1291_n N_VPWR_c_1697_n 0.00580593f $X=6.61 $Y=2.75 $X2=0
+ $Y2=0
cc_917 N_A_1156_90#_c_1285_n N_VPWR_c_1698_n 0.00614449f $X=7.885 $Y=1.95 $X2=0
+ $Y2=0
cc_918 N_A_1156_90#_c_1285_n N_VPWR_c_1708_n 0.00401159f $X=7.885 $Y=1.95 $X2=0
+ $Y2=0
cc_919 N_A_1156_90#_c_1291_n N_VPWR_c_1711_n 0.015569f $X=6.61 $Y=2.75 $X2=0
+ $Y2=0
cc_920 N_A_1156_90#_c_1285_n N_VPWR_c_1692_n 0.00515964f $X=7.885 $Y=1.95 $X2=0
+ $Y2=0
cc_921 N_A_1156_90#_c_1291_n N_VPWR_c_1692_n 0.0128526f $X=6.61 $Y=2.75 $X2=0
+ $Y2=0
cc_922 N_A_1156_90#_M1008_g N_VGND_c_1865_n 0.00129371f $X=7.8 $Y=0.77 $X2=0
+ $Y2=0
cc_923 N_A_1156_90#_M1008_g N_VGND_c_1873_n 8.23937e-19 $X=7.8 $Y=0.77 $X2=0
+ $Y2=0
cc_924 N_A_1895_74#_c_1390_n N_VPWR_c_1699_n 0.00712319f $X=11.495 $Y=2.215
+ $X2=0 $Y2=0
cc_925 N_A_1895_74#_c_1393_n N_VPWR_c_1699_n 0.0134376f $X=10.055 $Y=2.105 $X2=0
+ $Y2=0
cc_926 N_A_1895_74#_c_1392_n N_VPWR_c_1701_n 0.0100916f $X=12.465 $Y=1.765 $X2=0
+ $Y2=0
cc_927 N_A_1895_74#_c_1393_n N_VPWR_c_1712_n 0.0120294f $X=10.055 $Y=2.105 $X2=0
+ $Y2=0
cc_928 N_A_1895_74#_c_1390_n N_VPWR_c_1713_n 0.00541219f $X=11.495 $Y=2.215
+ $X2=0 $Y2=0
cc_929 N_A_1895_74#_c_1392_n N_VPWR_c_1713_n 0.00445602f $X=12.465 $Y=1.765
+ $X2=0 $Y2=0
cc_930 N_A_1895_74#_c_1390_n N_VPWR_c_1692_n 0.00536257f $X=11.495 $Y=2.215
+ $X2=0 $Y2=0
cc_931 N_A_1895_74#_c_1392_n N_VPWR_c_1692_n 0.00865852f $X=12.465 $Y=1.765
+ $X2=0 $Y2=0
cc_932 N_A_1895_74#_c_1393_n N_VPWR_c_1692_n 0.00926813f $X=10.055 $Y=2.105
+ $X2=0 $Y2=0
cc_933 N_A_1895_74#_c_1380_n N_Q_c_1831_n 0.00837961f $X=12.395 $Y=1.185 $X2=0
+ $Y2=0
cc_934 N_A_1895_74#_c_1379_n N_Q_c_1832_n 0.00274954f $X=12.32 $Y=1.26 $X2=0
+ $Y2=0
cc_935 N_A_1895_74#_c_1380_n N_Q_c_1832_n 0.00214314f $X=12.395 $Y=1.185 $X2=0
+ $Y2=0
cc_936 N_A_1895_74#_c_1378_n Q 4.67537e-19 $X=11.495 $Y=2.125 $X2=0 $Y2=0
cc_937 N_A_1895_74#_c_1390_n Q 0.0021229f $X=11.495 $Y=2.215 $X2=0 $Y2=0
cc_938 N_A_1895_74#_c_1381_n Q 0.00948321f $X=12.465 $Y=1.675 $X2=0 $Y2=0
cc_939 N_A_1895_74#_c_1392_n Q 0.0239007f $X=12.465 $Y=1.765 $X2=0 $Y2=0
cc_940 N_A_1895_74#_c_1379_n N_Q_c_1834_n 0.0167995f $X=12.32 $Y=1.26 $X2=0
+ $Y2=0
cc_941 N_A_1895_74#_c_1380_n N_Q_c_1834_n 0.00326896f $X=12.395 $Y=1.185 $X2=0
+ $Y2=0
cc_942 N_A_1895_74#_c_1381_n N_Q_c_1834_n 0.00920291f $X=12.465 $Y=1.675 $X2=0
+ $Y2=0
cc_943 N_A_1895_74#_c_1382_n N_Q_c_1834_n 0.00652656f $X=12.437 $Y=1.26 $X2=0
+ $Y2=0
cc_944 N_A_1895_74#_c_1383_n N_VGND_c_1866_n 0.0109084f $X=9.615 $Y=0.515 $X2=0
+ $Y2=0
cc_945 N_A_1895_74#_c_1380_n N_VGND_c_1868_n 0.0196825f $X=12.395 $Y=1.185 $X2=0
+ $Y2=0
cc_946 N_A_1895_74#_c_1382_n N_VGND_c_1868_n 0.00211944f $X=12.437 $Y=1.26 $X2=0
+ $Y2=0
cc_947 N_A_1895_74#_M1007_g N_VGND_c_1878_n 0.00461464f $X=11.405 $Y=0.58 $X2=0
+ $Y2=0
cc_948 N_A_1895_74#_c_1380_n N_VGND_c_1878_n 0.00434272f $X=12.395 $Y=1.185
+ $X2=0 $Y2=0
cc_949 N_A_1895_74#_c_1383_n N_VGND_c_1882_n 0.0145243f $X=9.615 $Y=0.515 $X2=0
+ $Y2=0
cc_950 N_A_1895_74#_M1007_g N_VGND_c_1883_n 0.00540028f $X=11.405 $Y=0.58 $X2=0
+ $Y2=0
cc_951 N_A_1895_74#_c_1383_n N_VGND_c_1883_n 0.00520222f $X=9.615 $Y=0.515 $X2=0
+ $Y2=0
cc_952 N_A_1895_74#_c_1384_n N_VGND_c_1883_n 0.0313981f $X=10.775 $Y=0.92 $X2=0
+ $Y2=0
cc_953 N_A_1895_74#_c_1386_n N_VGND_c_1883_n 0.0175339f $X=11.34 $Y=1.17 $X2=0
+ $Y2=0
cc_954 N_A_1895_74#_c_1387_n N_VGND_c_1883_n 0.00268565f $X=11.34 $Y=1.17 $X2=0
+ $Y2=0
cc_955 N_A_1895_74#_c_1388_n N_VGND_c_1883_n 0.0151641f $X=10.86 $Y=1.085 $X2=0
+ $Y2=0
cc_956 N_A_1895_74#_M1007_g N_VGND_c_1884_n 0.00917524f $X=11.405 $Y=0.58 $X2=0
+ $Y2=0
cc_957 N_A_1895_74#_c_1380_n N_VGND_c_1884_n 0.00828933f $X=12.395 $Y=1.185
+ $X2=0 $Y2=0
cc_958 N_A_1895_74#_c_1383_n N_VGND_c_1884_n 0.0119829f $X=9.615 $Y=0.515 $X2=0
+ $Y2=0
cc_959 N_A_1895_74#_c_1384_n N_VGND_c_1884_n 0.0191617f $X=10.775 $Y=0.92 $X2=0
+ $Y2=0
cc_960 N_A_1895_74#_c_1388_n N_VGND_c_1884_n 6.25089e-19 $X=10.86 $Y=1.085 $X2=0
+ $Y2=0
cc_961 N_A_27_508#_c_1526_n N_VPWR_M1012_d 0.00654762f $X=2.13 $Y=2.905 $X2=0
+ $Y2=0
cc_962 N_A_27_508#_c_1530_n N_VPWR_M1002_s 0.00767671f $X=5.13 $Y=2.395 $X2=0
+ $Y2=0
cc_963 N_A_27_508#_c_1530_n N_VPWR_M1019_s 0.00194622f $X=5.13 $Y=2.395 $X2=0
+ $Y2=0
cc_964 N_A_27_508#_c_1531_n N_VPWR_M1019_s 0.0113914f $X=5.215 $Y=2.31 $X2=0
+ $Y2=0
cc_965 N_A_27_508#_c_1600_n N_VPWR_M1019_s 0.0019583f $X=5.61 $Y=2.605 $X2=0
+ $Y2=0
cc_966 N_A_27_508#_c_1521_n N_VPWR_c_1693_n 0.0138422f $X=0.27 $Y=2.75 $X2=0
+ $Y2=0
cc_967 N_A_27_508#_c_1522_n N_VPWR_c_1693_n 0.0202063f $X=1.365 $Y=2.265 $X2=0
+ $Y2=0
cc_968 N_A_27_508#_c_1523_n N_VPWR_c_1693_n 0.0292993f $X=1.45 $Y=2.905 $X2=0
+ $Y2=0
cc_969 N_A_27_508#_c_1525_n N_VPWR_c_1693_n 0.0146662f $X=1.535 $Y=2.99 $X2=0
+ $Y2=0
cc_970 N_A_27_508#_c_1524_n N_VPWR_c_1694_n 0.0147456f $X=2.045 $Y=2.99 $X2=0
+ $Y2=0
cc_971 N_A_27_508#_c_1526_n N_VPWR_c_1694_n 0.0465119f $X=2.13 $Y=2.905 $X2=0
+ $Y2=0
cc_972 N_A_27_508#_c_1527_n N_VPWR_c_1694_n 0.0175725f $X=3.1 $Y=2.035 $X2=0
+ $Y2=0
cc_973 N_A_27_508#_c_1535_n N_VPWR_c_1694_n 0.0111172f $X=3.31 $Y=2.39 $X2=0
+ $Y2=0
cc_974 N_A_27_508#_c_1530_n N_VPWR_c_1695_n 0.0215735f $X=5.13 $Y=2.395 $X2=0
+ $Y2=0
cc_975 N_A_27_508#_c_1530_n N_VPWR_c_1696_n 0.00876485f $X=5.13 $Y=2.395 $X2=0
+ $Y2=0
cc_976 N_A_27_508#_c_1600_n N_VPWR_c_1696_n 0.0154296f $X=5.61 $Y=2.605 $X2=0
+ $Y2=0
cc_977 N_A_27_508#_c_1521_n N_VPWR_c_1702_n 0.0154862f $X=0.27 $Y=2.75 $X2=0
+ $Y2=0
cc_978 N_A_27_508#_c_1524_n N_VPWR_c_1704_n 0.0449818f $X=2.045 $Y=2.99 $X2=0
+ $Y2=0
cc_979 N_A_27_508#_c_1525_n N_VPWR_c_1704_n 0.0121867f $X=1.535 $Y=2.99 $X2=0
+ $Y2=0
cc_980 N_A_27_508#_c_1535_n N_VPWR_c_1706_n 0.00632564f $X=3.31 $Y=2.39 $X2=0
+ $Y2=0
cc_981 N_A_27_508#_c_1532_n N_VPWR_c_1711_n 0.00681477f $X=5.995 $Y=2.605 $X2=0
+ $Y2=0
cc_982 N_A_27_508#_c_1600_n N_VPWR_c_1711_n 0.00256262f $X=5.61 $Y=2.605 $X2=0
+ $Y2=0
cc_983 N_A_27_508#_c_1533_n N_VPWR_c_1711_n 0.0107588f $X=6.16 $Y=2.75 $X2=0
+ $Y2=0
cc_984 N_A_27_508#_c_1521_n N_VPWR_c_1692_n 0.0127853f $X=0.27 $Y=2.75 $X2=0
+ $Y2=0
cc_985 N_A_27_508#_c_1524_n N_VPWR_c_1692_n 0.025776f $X=2.045 $Y=2.99 $X2=0
+ $Y2=0
cc_986 N_A_27_508#_c_1525_n N_VPWR_c_1692_n 0.00660921f $X=1.535 $Y=2.99 $X2=0
+ $Y2=0
cc_987 N_A_27_508#_c_1530_n N_VPWR_c_1692_n 0.0426254f $X=5.13 $Y=2.395 $X2=0
+ $Y2=0
cc_988 N_A_27_508#_c_1532_n N_VPWR_c_1692_n 0.0109468f $X=5.995 $Y=2.605 $X2=0
+ $Y2=0
cc_989 N_A_27_508#_c_1600_n N_VPWR_c_1692_n 0.0105038f $X=5.61 $Y=2.605 $X2=0
+ $Y2=0
cc_990 N_A_27_508#_c_1533_n N_VPWR_c_1692_n 0.00904147f $X=6.16 $Y=2.75 $X2=0
+ $Y2=0
cc_991 N_A_27_508#_c_1535_n N_VPWR_c_1692_n 0.0106028f $X=3.31 $Y=2.39 $X2=0
+ $Y2=0
cc_992 N_A_27_508#_c_1518_n N_VGND_c_1861_n 0.00841519f $X=0.365 $Y=0.575 $X2=0
+ $Y2=0
cc_993 N_A_27_508#_c_1519_n N_VGND_c_1862_n 0.01581f $X=3.185 $Y=0.645 $X2=0
+ $Y2=0
cc_994 N_A_27_508#_c_1515_n N_VGND_c_1863_n 0.00998528f $X=3.185 $Y=1.95 $X2=0
+ $Y2=0
cc_995 N_A_27_508#_c_1519_n N_VGND_c_1863_n 0.0369819f $X=3.185 $Y=0.645 $X2=0
+ $Y2=0
cc_996 N_A_27_508#_c_1519_n N_VGND_c_1869_n 0.0163765f $X=3.185 $Y=0.645 $X2=0
+ $Y2=0
cc_997 N_A_27_508#_c_1518_n N_VGND_c_1875_n 0.0199786f $X=0.365 $Y=0.575 $X2=0
+ $Y2=0
cc_998 N_A_27_508#_c_1518_n N_VGND_c_1884_n 0.0162038f $X=0.365 $Y=0.575 $X2=0
+ $Y2=0
cc_999 N_A_27_508#_c_1519_n N_VGND_c_1884_n 0.0167347f $X=3.185 $Y=0.645 $X2=0
+ $Y2=0
cc_1000 N_VPWR_c_1701_n Q 0.0778383f $X=12.69 $Y=1.985 $X2=0 $Y2=0
cc_1001 N_VPWR_c_1713_n Q 0.0145938f $X=12.605 $Y=3.33 $X2=0 $Y2=0
cc_1002 N_VPWR_c_1692_n Q 0.0120466f $X=12.72 $Y=3.33 $X2=0 $Y2=0
cc_1003 N_Q_c_1831_n N_VGND_c_1868_n 0.0308109f $X=12.18 $Y=0.515 $X2=0 $Y2=0
cc_1004 N_Q_c_1831_n N_VGND_c_1878_n 0.0145639f $X=12.18 $Y=0.515 $X2=0 $Y2=0
cc_1005 N_Q_c_1831_n N_VGND_c_1884_n 0.0119984f $X=12.18 $Y=0.515 $X2=0 $Y2=0
