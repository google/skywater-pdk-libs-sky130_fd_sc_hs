# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_hs__a2111o_4
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_hs__a2111o_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  8.160000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.285000 1.450000 7.075000 1.780000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.245000 1.260000 8.035000 1.780000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.405000 1.450000 6.115000 1.780000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.965000 1.450000 5.155000 1.780000 ;
    END
  END C1
  PIN D1
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.385000 1.260000 3.715000 1.780000 ;
    END
  END D1
  PIN X
    ANTENNADIFFAREA  1.086400 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 0.960000 2.445000 1.130000 ;
        RECT 0.125000 1.130000 0.650000 1.800000 ;
        RECT 0.125000 1.800000 2.065000 1.970000 ;
        RECT 0.835000 1.970000 1.165000 2.980000 ;
        RECT 1.415000 0.350000 1.665000 0.960000 ;
        RECT 1.735000 1.970000 2.065000 2.980000 ;
        RECT 2.195000 0.350000 2.445000 0.960000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 8.160000 0.085000 ;
        RECT 0.905000  0.085000 1.235000 0.790000 ;
        RECT 1.845000  0.085000 2.015000 0.790000 ;
        RECT 2.625000  0.085000 2.875000 1.030000 ;
        RECT 3.530000  0.085000 3.870000 0.750000 ;
        RECT 4.400000  0.085000 4.740000 0.940000 ;
        RECT 5.270000  0.085000 5.600000 0.940000 ;
        RECT 7.300000  0.085000 7.630000 0.750000 ;
      LAYER mcon ;
        RECT 0.155000 -0.085000 0.325000 0.085000 ;
        RECT 0.635000 -0.085000 0.805000 0.085000 ;
        RECT 1.115000 -0.085000 1.285000 0.085000 ;
        RECT 1.595000 -0.085000 1.765000 0.085000 ;
        RECT 2.075000 -0.085000 2.245000 0.085000 ;
        RECT 2.555000 -0.085000 2.725000 0.085000 ;
        RECT 3.035000 -0.085000 3.205000 0.085000 ;
        RECT 3.515000 -0.085000 3.685000 0.085000 ;
        RECT 3.995000 -0.085000 4.165000 0.085000 ;
        RECT 4.475000 -0.085000 4.645000 0.085000 ;
        RECT 4.955000 -0.085000 5.125000 0.085000 ;
        RECT 5.435000 -0.085000 5.605000 0.085000 ;
        RECT 5.915000 -0.085000 6.085000 0.085000 ;
        RECT 6.395000 -0.085000 6.565000 0.085000 ;
        RECT 6.875000 -0.085000 7.045000 0.085000 ;
        RECT 7.355000 -0.085000 7.525000 0.085000 ;
        RECT 7.835000 -0.085000 8.005000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.245000 8.160000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 3.245000 8.160000 3.415000 ;
        RECT 0.385000 2.140000 0.635000 3.245000 ;
        RECT 1.365000 2.140000 1.535000 3.245000 ;
        RECT 2.265000 1.820000 2.515000 3.245000 ;
        RECT 6.375000 2.290000 6.705000 3.245000 ;
        RECT 7.275000 2.290000 7.525000 3.245000 ;
      LAYER mcon ;
        RECT 0.155000 3.245000 0.325000 3.415000 ;
        RECT 0.635000 3.245000 0.805000 3.415000 ;
        RECT 1.115000 3.245000 1.285000 3.415000 ;
        RECT 1.595000 3.245000 1.765000 3.415000 ;
        RECT 2.075000 3.245000 2.245000 3.415000 ;
        RECT 2.555000 3.245000 2.725000 3.415000 ;
        RECT 3.035000 3.245000 3.205000 3.415000 ;
        RECT 3.515000 3.245000 3.685000 3.415000 ;
        RECT 3.995000 3.245000 4.165000 3.415000 ;
        RECT 4.475000 3.245000 4.645000 3.415000 ;
        RECT 4.955000 3.245000 5.125000 3.415000 ;
        RECT 5.435000 3.245000 5.605000 3.415000 ;
        RECT 5.915000 3.245000 6.085000 3.415000 ;
        RECT 6.395000 3.245000 6.565000 3.415000 ;
        RECT 6.875000 3.245000 7.045000 3.415000 ;
        RECT 7.355000 3.245000 7.525000 3.415000 ;
        RECT 7.835000 3.245000 8.005000 3.415000 ;
      LAYER met1 ;
        RECT 0.000000 3.085000 8.160000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.870000 1.300000 3.215000 1.630000 ;
      RECT 2.705000 2.290000 3.035000 2.905000 ;
      RECT 2.705000 2.905000 4.835000 3.075000 ;
      RECT 3.045000 0.350000 3.350000 0.920000 ;
      RECT 3.045000 0.920000 4.220000 1.090000 ;
      RECT 3.045000 1.090000 3.215000 1.300000 ;
      RECT 3.045000 1.630000 3.215000 1.950000 ;
      RECT 3.045000 1.950000 3.405000 2.120000 ;
      RECT 3.235000 2.120000 3.405000 2.735000 ;
      RECT 3.605000 1.950000 3.935000 2.905000 ;
      RECT 4.050000 0.350000 4.220000 0.920000 ;
      RECT 4.050000 1.090000 4.220000 1.110000 ;
      RECT 4.050000 1.110000 6.770000 1.280000 ;
      RECT 4.135000 1.950000 5.805000 2.120000 ;
      RECT 4.135000 2.120000 4.305000 2.735000 ;
      RECT 4.505000 2.290000 4.835000 2.905000 ;
      RECT 4.920000 0.350000 5.090000 1.110000 ;
      RECT 5.025000 2.290000 5.305000 2.905000 ;
      RECT 5.025000 2.905000 6.175000 3.075000 ;
      RECT 5.475000 2.120000 5.805000 2.735000 ;
      RECT 6.005000 1.950000 8.055000 2.120000 ;
      RECT 6.005000 2.120000 6.175000 2.905000 ;
      RECT 6.010000 0.285000 7.120000 0.455000 ;
      RECT 6.010000 0.455000 6.340000 0.940000 ;
      RECT 6.510000 0.625000 6.770000 1.110000 ;
      RECT 6.905000 2.120000 7.075000 2.980000 ;
      RECT 6.950000 0.455000 7.120000 0.920000 ;
      RECT 6.950000 0.920000 8.060000 1.090000 ;
      RECT 7.725000 2.120000 8.055000 2.980000 ;
      RECT 7.810000 0.350000 8.060000 0.920000 ;
  END
END sky130_fd_sc_hs__a2111o_4
