* File: sky130_fd_sc_hs__o2bb2ai_4.pxi.spice
* Created: Tue Sep  1 20:17:12 2020
* 
x_PM_SKY130_FD_SC_HS__O2BB2AI_4%A1_N N_A1_N_M1009_g N_A1_N_c_173_n
+ N_A1_N_M1001_g N_A1_N_M1032_g N_A1_N_c_174_n N_A1_N_M1002_g N_A1_N_M1033_g
+ N_A1_N_c_175_n N_A1_N_M1004_g N_A1_N_M1034_g N_A1_N_c_176_n N_A1_N_M1008_g
+ A1_N A1_N A1_N A1_N N_A1_N_c_171_n N_A1_N_c_172_n
+ PM_SKY130_FD_SC_HS__O2BB2AI_4%A1_N
x_PM_SKY130_FD_SC_HS__O2BB2AI_4%A2_N N_A2_N_M1006_g N_A2_N_c_257_n
+ N_A2_N_M1011_g N_A2_N_M1013_g N_A2_N_c_258_n N_A2_N_M1014_g N_A2_N_M1021_g
+ N_A2_N_c_259_n N_A2_N_M1015_g N_A2_N_c_253_n N_A2_N_c_254_n N_A2_N_c_255_n
+ N_A2_N_M1017_g N_A2_N_M1039_g A2_N A2_N PM_SKY130_FD_SC_HS__O2BB2AI_4%A2_N
x_PM_SKY130_FD_SC_HS__O2BB2AI_4%A_114_368# N_A_114_368#_M1006_s
+ N_A_114_368#_M1021_s N_A_114_368#_M1001_d N_A_114_368#_M1004_d
+ N_A_114_368#_M1011_d N_A_114_368#_M1015_d N_A_114_368#_c_355_n
+ N_A_114_368#_M1003_g N_A_114_368#_c_356_n N_A_114_368#_M1019_g
+ N_A_114_368#_M1007_g N_A_114_368#_c_357_n N_A_114_368#_M1026_g
+ N_A_114_368#_M1016_g N_A_114_368#_c_358_n N_A_114_368#_M1028_g
+ N_A_114_368#_M1022_g N_A_114_368#_c_348_n N_A_114_368#_c_349_n
+ N_A_114_368#_M1030_g N_A_114_368#_c_365_n N_A_114_368#_c_360_n
+ N_A_114_368#_c_372_n N_A_114_368#_c_361_n N_A_114_368#_c_379_n
+ N_A_114_368#_c_393_n N_A_114_368#_c_362_n N_A_114_368#_c_351_n
+ N_A_114_368#_c_352_n N_A_114_368#_c_407_n N_A_114_368#_c_363_n
+ N_A_114_368#_c_414_n N_A_114_368#_c_353_n N_A_114_368#_c_364_n
+ N_A_114_368#_c_354_n N_A_114_368#_c_382_n N_A_114_368#_c_427_n
+ N_A_114_368#_c_431_n PM_SKY130_FD_SC_HS__O2BB2AI_4%A_114_368#
x_PM_SKY130_FD_SC_HS__O2BB2AI_4%B2 N_B2_M1000_g N_B2_c_558_n N_B2_M1018_g
+ N_B2_M1024_g N_B2_c_559_n N_B2_M1020_g N_B2_M1027_g N_B2_c_560_n N_B2_M1023_g
+ N_B2_c_561_n N_B2_M1025_g N_B2_M1037_g B2 B2 B2 B2 N_B2_c_556_n N_B2_c_557_n
+ PM_SKY130_FD_SC_HS__O2BB2AI_4%B2
x_PM_SKY130_FD_SC_HS__O2BB2AI_4%B1 N_B1_M1005_g N_B1_c_649_n N_B1_M1029_g
+ N_B1_M1010_g N_B1_c_650_n N_B1_M1031_g N_B1_M1012_g N_B1_c_651_n N_B1_M1036_g
+ N_B1_M1035_g N_B1_c_652_n N_B1_M1038_g B1 B1 B1 B1 N_B1_c_648_n
+ PM_SKY130_FD_SC_HS__O2BB2AI_4%B1
x_PM_SKY130_FD_SC_HS__O2BB2AI_4%VPWR N_VPWR_M1001_s N_VPWR_M1002_s
+ N_VPWR_M1008_s N_VPWR_M1014_s N_VPWR_M1017_s N_VPWR_M1019_d N_VPWR_M1028_d
+ N_VPWR_M1029_d N_VPWR_M1036_d N_VPWR_c_725_n N_VPWR_c_726_n N_VPWR_c_727_n
+ N_VPWR_c_728_n N_VPWR_c_729_n N_VPWR_c_730_n N_VPWR_c_731_n N_VPWR_c_732_n
+ N_VPWR_c_733_n N_VPWR_c_734_n N_VPWR_c_735_n N_VPWR_c_736_n N_VPWR_c_737_n
+ N_VPWR_c_738_n N_VPWR_c_739_n N_VPWR_c_740_n N_VPWR_c_741_n N_VPWR_c_742_n
+ N_VPWR_c_743_n N_VPWR_c_744_n N_VPWR_c_745_n VPWR N_VPWR_c_746_n
+ N_VPWR_c_747_n N_VPWR_c_748_n N_VPWR_c_724_n N_VPWR_c_750_n N_VPWR_c_751_n
+ N_VPWR_c_752_n PM_SKY130_FD_SC_HS__O2BB2AI_4%VPWR
x_PM_SKY130_FD_SC_HS__O2BB2AI_4%Y N_Y_M1007_s N_Y_M1022_s N_Y_M1003_s
+ N_Y_M1026_s N_Y_M1018_d N_Y_M1023_d N_Y_c_881_n N_Y_c_882_n N_Y_c_883_n
+ N_Y_c_900_n N_Y_c_877_n N_Y_c_878_n N_Y_c_884_n N_Y_c_913_n N_Y_c_879_n
+ N_Y_c_886_n N_Y_c_887_n N_Y_c_939_n N_Y_c_880_n N_Y_c_943_n N_Y_c_948_n Y
+ PM_SKY130_FD_SC_HS__O2BB2AI_4%Y
x_PM_SKY130_FD_SC_HS__O2BB2AI_4%A_1215_368# N_A_1215_368#_M1018_s
+ N_A_1215_368#_M1020_s N_A_1215_368#_M1025_s N_A_1215_368#_M1031_s
+ N_A_1215_368#_M1038_s N_A_1215_368#_c_988_n N_A_1215_368#_c_989_n
+ N_A_1215_368#_c_990_n N_A_1215_368#_c_1051_n N_A_1215_368#_c_991_n
+ N_A_1215_368#_c_1003_n N_A_1215_368#_c_992_n N_A_1215_368#_c_1011_n
+ N_A_1215_368#_c_993_n N_A_1215_368#_c_994_n N_A_1215_368#_c_995_n
+ N_A_1215_368#_c_1020_n PM_SKY130_FD_SC_HS__O2BB2AI_4%A_1215_368#
x_PM_SKY130_FD_SC_HS__O2BB2AI_4%A_27_74# N_A_27_74#_M1009_d N_A_27_74#_M1032_d
+ N_A_27_74#_M1034_d N_A_27_74#_M1013_d N_A_27_74#_M1039_d N_A_27_74#_c_1054_n
+ N_A_27_74#_c_1055_n N_A_27_74#_c_1056_n N_A_27_74#_c_1057_n
+ N_A_27_74#_c_1058_n N_A_27_74#_c_1059_n N_A_27_74#_c_1060_n
+ N_A_27_74#_c_1093_n N_A_27_74#_c_1061_n N_A_27_74#_c_1062_n
+ N_A_27_74#_c_1063_n N_A_27_74#_c_1064_n PM_SKY130_FD_SC_HS__O2BB2AI_4%A_27_74#
x_PM_SKY130_FD_SC_HS__O2BB2AI_4%VGND N_VGND_M1009_s N_VGND_M1033_s
+ N_VGND_M1000_d N_VGND_M1027_d N_VGND_M1005_s N_VGND_M1012_s N_VGND_c_1122_n
+ N_VGND_c_1123_n N_VGND_c_1124_n N_VGND_c_1125_n N_VGND_c_1126_n
+ N_VGND_c_1127_n N_VGND_c_1128_n VGND N_VGND_c_1129_n N_VGND_c_1130_n
+ N_VGND_c_1131_n N_VGND_c_1132_n N_VGND_c_1133_n N_VGND_c_1134_n
+ N_VGND_c_1135_n N_VGND_c_1136_n N_VGND_c_1137_n N_VGND_c_1138_n
+ N_VGND_c_1139_n N_VGND_c_1140_n N_VGND_c_1141_n
+ PM_SKY130_FD_SC_HS__O2BB2AI_4%VGND
x_PM_SKY130_FD_SC_HS__O2BB2AI_4%A_857_74# N_A_857_74#_M1007_d
+ N_A_857_74#_M1016_d N_A_857_74#_M1030_d N_A_857_74#_M1024_s
+ N_A_857_74#_M1037_s N_A_857_74#_M1010_d N_A_857_74#_M1035_d
+ N_A_857_74#_c_1251_n N_A_857_74#_c_1252_n N_A_857_74#_c_1253_n
+ N_A_857_74#_c_1318_n N_A_857_74#_c_1254_n N_A_857_74#_c_1255_n
+ N_A_857_74#_c_1256_n N_A_857_74#_c_1257_n N_A_857_74#_c_1258_n
+ N_A_857_74#_c_1259_n N_A_857_74#_c_1260_n N_A_857_74#_c_1261_n
+ N_A_857_74#_c_1262_n N_A_857_74#_c_1263_n N_A_857_74#_c_1264_n
+ N_A_857_74#_c_1265_n N_A_857_74#_c_1266_n N_A_857_74#_c_1267_n
+ PM_SKY130_FD_SC_HS__O2BB2AI_4%A_857_74#
cc_1 VNB N_A1_N_M1009_g 0.0318708f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_2 VNB N_A1_N_M1032_g 0.0226407f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=0.74
cc_3 VNB N_A1_N_M1033_g 0.0226407f $X=-0.19 $Y=-0.245 $X2=1.365 $Y2=0.74
cc_4 VNB N_A1_N_M1034_g 0.0229726f $X=-0.19 $Y=-0.245 $X2=1.795 $Y2=0.74
cc_5 VNB N_A1_N_c_171_n 0.0160224f $X=-0.19 $Y=-0.245 $X2=1.77 $Y2=1.515
cc_6 VNB N_A1_N_c_172_n 0.0810377f $X=-0.19 $Y=-0.245 $X2=1.795 $Y2=1.557
cc_7 VNB N_A2_N_M1006_g 0.0213573f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_8 VNB N_A2_N_M1013_g 0.0218695f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=0.74
cc_9 VNB N_A2_N_M1021_g 0.0224304f $X=-0.19 $Y=-0.245 $X2=1.365 $Y2=0.74
cc_10 VNB N_A2_N_c_253_n 0.0106061f $X=-0.19 $Y=-0.245 $X2=1.795 $Y2=1.35
cc_11 VNB N_A2_N_c_254_n 0.0571439f $X=-0.19 $Y=-0.245 $X2=1.795 $Y2=0.74
cc_12 VNB N_A2_N_c_255_n 0.0140026f $X=-0.19 $Y=-0.245 $X2=1.795 $Y2=0.74
cc_13 VNB N_A2_N_M1039_g 0.0282424f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_14 VNB N_A_114_368#_M1007_g 0.027434f $X=-0.19 $Y=-0.245 $X2=1.845 $Y2=2.4
cc_15 VNB N_A_114_368#_M1016_g 0.0200535f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_114_368#_M1022_g 0.0193643f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=1.557
cc_17 VNB N_A_114_368#_c_348_n 0.0243374f $X=-0.19 $Y=-0.245 $X2=1.365 $Y2=1.557
cc_18 VNB N_A_114_368#_c_349_n 0.117009f $X=-0.19 $Y=-0.245 $X2=1.395 $Y2=1.557
cc_19 VNB N_A_114_368#_M1030_g 0.020471f $X=-0.19 $Y=-0.245 $X2=1.77 $Y2=1.515
cc_20 VNB N_A_114_368#_c_351_n 0.00349695f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_114_368#_c_352_n 0.00229069f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_114_368#_c_353_n 0.00589432f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_114_368#_c_354_n 0.0113354f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_B2_M1000_g 0.0239651f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_25 VNB N_B2_M1024_g 0.0240453f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=0.74
cc_26 VNB N_B2_M1027_g 0.0234895f $X=-0.19 $Y=-0.245 $X2=1.365 $Y2=0.74
cc_27 VNB N_B2_M1037_g 0.0245189f $X=-0.19 $Y=-0.245 $X2=1.845 $Y2=2.4
cc_28 VNB N_B2_c_556_n 0.00585801f $X=-0.19 $Y=-0.245 $X2=1.795 $Y2=1.557
cc_29 VNB N_B2_c_557_n 0.0755667f $X=-0.19 $Y=-0.245 $X2=1.845 $Y2=1.557
cc_30 VNB N_B1_M1005_g 0.0230003f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_31 VNB N_B1_M1010_g 0.0224928f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=0.74
cc_32 VNB N_B1_M1012_g 0.0240453f $X=-0.19 $Y=-0.245 $X2=1.365 $Y2=0.74
cc_33 VNB N_B1_M1035_g 0.0328675f $X=-0.19 $Y=-0.245 $X2=1.795 $Y2=0.74
cc_34 VNB B1 0.0153948f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=1.58
cc_35 VNB N_B1_c_648_n 0.082811f $X=-0.19 $Y=-0.245 $X2=1.77 $Y2=1.515
cc_36 VNB N_VPWR_c_724_n 0.422413f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_Y_c_877_n 0.00258452f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.58
cc_38 VNB N_Y_c_878_n 0.00229484f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=1.58
cc_39 VNB N_Y_c_879_n 0.00349117f $X=-0.19 $Y=-0.245 $X2=0.945 $Y2=1.557
cc_40 VNB N_Y_c_880_n 0.00416741f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_27_74#_c_1054_n 0.0266107f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_27_74#_c_1055_n 0.00307486f $X=-0.19 $Y=-0.245 $X2=1.395 $Y2=2.4
cc_43 VNB N_A_27_74#_c_1056_n 0.00955057f $X=-0.19 $Y=-0.245 $X2=1.395 $Y2=2.4
cc_44 VNB N_A_27_74#_c_1057_n 0.00188248f $X=-0.19 $Y=-0.245 $X2=1.795 $Y2=0.74
cc_45 VNB N_A_27_74#_c_1058_n 0.0101688f $X=-0.19 $Y=-0.245 $X2=1.845 $Y2=1.765
cc_46 VNB N_A_27_74#_c_1059_n 0.0026914f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=1.58
cc_47 VNB N_A_27_74#_c_1060_n 0.00211517f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_27_74#_c_1061_n 0.00647211f $X=-0.19 $Y=-0.245 $X2=0.41 $Y2=1.515
cc_49 VNB N_A_27_74#_c_1062_n 0.00865153f $X=-0.19 $Y=-0.245 $X2=0.945 $Y2=1.557
cc_50 VNB N_A_27_74#_c_1063_n 0.00133271f $X=-0.19 $Y=-0.245 $X2=1.395 $Y2=1.557
cc_51 VNB N_A_27_74#_c_1064_n 0.00244965f $X=-0.19 $Y=-0.245 $X2=1.77 $Y2=1.557
cc_52 VNB N_VGND_c_1122_n 0.00324953f $X=-0.19 $Y=-0.245 $X2=1.395 $Y2=2.4
cc_53 VNB N_VGND_c_1123_n 0.00324953f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_VGND_c_1124_n 0.108794f $X=-0.19 $Y=-0.245 $X2=1.845 $Y2=2.4
cc_55 VNB N_VGND_c_1125_n 0.00558127f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.58
cc_56 VNB N_VGND_c_1126_n 0.00494723f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_VGND_c_1127_n 0.00269659f $X=-0.19 $Y=-0.245 $X2=0.41 $Y2=1.515
cc_58 VNB N_VGND_c_1128_n 0.00558127f $X=-0.19 $Y=-0.245 $X2=1.365 $Y2=1.557
cc_59 VNB N_VGND_c_1129_n 0.0173909f $X=-0.19 $Y=-0.245 $X2=1.77 $Y2=1.515
cc_60 VNB N_VGND_c_1130_n 0.0154137f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_VGND_c_1131_n 0.0169342f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_VGND_c_1132_n 0.0169342f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_VGND_c_1133_n 0.0169342f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_VGND_c_1134_n 0.0173909f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_VGND_c_1135_n 0.534813f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_VGND_c_1136_n 0.00604233f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_VGND_c_1137_n 0.00604233f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_VGND_c_1138_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_VGND_c_1139_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_VGND_c_1140_n 0.00604233f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_VGND_c_1141_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_A_857_74#_c_1251_n 0.00792168f $X=-0.19 $Y=-0.245 $X2=1.795 $Y2=0.74
cc_73 VNB N_A_857_74#_c_1252_n 0.0027626f $X=-0.19 $Y=-0.245 $X2=1.845 $Y2=1.765
cc_74 VNB N_A_857_74#_c_1253_n 0.00377359f $X=-0.19 $Y=-0.245 $X2=1.845 $Y2=2.4
cc_75 VNB N_A_857_74#_c_1254_n 0.00487777f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=1.58
cc_76 VNB N_A_857_74#_c_1255_n 0.00317099f $X=-0.19 $Y=-0.245 $X2=0.41 $Y2=1.515
cc_77 VNB N_A_857_74#_c_1256_n 0.00219196f $X=-0.19 $Y=-0.245 $X2=0.41 $Y2=1.515
cc_78 VNB N_A_857_74#_c_1257_n 0.00206666f $X=-0.19 $Y=-0.245 $X2=0.945
+ $Y2=1.557
cc_79 VNB N_A_857_74#_c_1258_n 0.00518435f $X=-0.19 $Y=-0.245 $X2=1.395
+ $Y2=1.557
cc_80 VNB N_A_857_74#_c_1259_n 0.00206666f $X=-0.19 $Y=-0.245 $X2=1.795
+ $Y2=1.557
cc_81 VNB N_A_857_74#_c_1260_n 0.00448959f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.565
cc_82 VNB N_A_857_74#_c_1261_n 0.00206666f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.565
cc_83 VNB N_A_857_74#_c_1262_n 0.0125337f $X=-0.19 $Y=-0.245 $X2=1.2 $Y2=1.565
cc_84 VNB N_A_857_74#_c_1263_n 0.0266107f $X=-0.19 $Y=-0.245 $X2=1.77 $Y2=1.565
cc_85 VNB N_A_857_74#_c_1264_n 0.00121798f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_86 VNB N_A_857_74#_c_1265_n 0.00178779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_87 VNB N_A_857_74#_c_1266_n 0.0090169f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_88 VNB N_A_857_74#_c_1267_n 0.00178779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_89 VPB N_A1_N_c_173_n 0.0179811f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.765
cc_90 VPB N_A1_N_c_174_n 0.0155127f $X=-0.19 $Y=1.66 $X2=0.945 $Y2=1.765
cc_91 VPB N_A1_N_c_175_n 0.0155127f $X=-0.19 $Y=1.66 $X2=1.395 $Y2=1.765
cc_92 VPB N_A1_N_c_176_n 0.0158162f $X=-0.19 $Y=1.66 $X2=1.845 $Y2=1.765
cc_93 VPB N_A1_N_c_171_n 0.0189682f $X=-0.19 $Y=1.66 $X2=1.77 $Y2=1.515
cc_94 VPB N_A1_N_c_172_n 0.0519715f $X=-0.19 $Y=1.66 $X2=1.795 $Y2=1.557
cc_95 VPB N_A2_N_c_257_n 0.0158886f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.765
cc_96 VPB N_A2_N_c_258_n 0.0155113f $X=-0.19 $Y=1.66 $X2=0.945 $Y2=1.765
cc_97 VPB N_A2_N_c_259_n 0.0155447f $X=-0.19 $Y=1.66 $X2=1.395 $Y2=1.765
cc_98 VPB N_A2_N_c_254_n 0.0348179f $X=-0.19 $Y=1.66 $X2=1.795 $Y2=0.74
cc_99 VPB N_A2_N_c_255_n 0.0221829f $X=-0.19 $Y=1.66 $X2=1.795 $Y2=0.74
cc_100 VPB A2_N 0.00559536f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_101 VPB N_A_114_368#_c_355_n 0.0157503f $X=-0.19 $Y=1.66 $X2=1.395 $Y2=1.765
cc_102 VPB N_A_114_368#_c_356_n 0.015247f $X=-0.19 $Y=1.66 $X2=1.795 $Y2=1.35
cc_103 VPB N_A_114_368#_c_357_n 0.015242f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_104 VPB N_A_114_368#_c_358_n 0.0172702f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_105 VPB N_A_114_368#_c_349_n 0.0263278f $X=-0.19 $Y=1.66 $X2=1.395 $Y2=1.557
cc_106 VPB N_A_114_368#_c_360_n 0.00257348f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_107 VPB N_A_114_368#_c_361_n 0.00257348f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_108 VPB N_A_114_368#_c_362_n 0.00257348f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_109 VPB N_A_114_368#_c_363_n 0.00257348f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_110 VPB N_A_114_368#_c_364_n 0.00129086f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_111 VPB N_B2_c_558_n 0.0174849f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.765
cc_112 VPB N_B2_c_559_n 0.014664f $X=-0.19 $Y=1.66 $X2=0.945 $Y2=1.765
cc_113 VPB N_B2_c_560_n 0.014664f $X=-0.19 $Y=1.66 $X2=1.395 $Y2=1.765
cc_114 VPB N_B2_c_561_n 0.0149125f $X=-0.19 $Y=1.66 $X2=1.795 $Y2=1.35
cc_115 VPB N_B2_c_556_n 0.0148402f $X=-0.19 $Y=1.66 $X2=1.795 $Y2=1.557
cc_116 VPB N_B2_c_557_n 0.0501886f $X=-0.19 $Y=1.66 $X2=1.845 $Y2=1.557
cc_117 VPB N_B1_c_649_n 0.0152732f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.765
cc_118 VPB N_B1_c_650_n 0.0155114f $X=-0.19 $Y=1.66 $X2=0.945 $Y2=1.765
cc_119 VPB N_B1_c_651_n 0.0155114f $X=-0.19 $Y=1.66 $X2=1.395 $Y2=1.765
cc_120 VPB N_B1_c_652_n 0.02086f $X=-0.19 $Y=1.66 $X2=1.845 $Y2=1.765
cc_121 VPB B1 0.0162213f $X=-0.19 $Y=1.66 $X2=1.595 $Y2=1.58
cc_122 VPB N_B1_c_648_n 0.0529031f $X=-0.19 $Y=1.66 $X2=1.77 $Y2=1.515
cc_123 VPB N_VPWR_c_725_n 0.0103331f $X=-0.19 $Y=1.66 $X2=1.845 $Y2=2.4
cc_124 VPB N_VPWR_c_726_n 0.0506502f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_125 VPB N_VPWR_c_727_n 0.00799266f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_126 VPB N_VPWR_c_728_n 0.00799266f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.557
cc_127 VPB N_VPWR_c_729_n 0.00799266f $X=-0.19 $Y=1.66 $X2=1.395 $Y2=1.557
cc_128 VPB N_VPWR_c_730_n 0.0100001f $X=-0.19 $Y=1.66 $X2=1.795 $Y2=1.557
cc_129 VPB N_VPWR_c_731_n 0.00734662f $X=-0.19 $Y=1.66 $X2=0.72 $Y2=1.565
cc_130 VPB N_VPWR_c_732_n 0.0185253f $X=-0.19 $Y=1.66 $X2=1.2 $Y2=1.565
cc_131 VPB N_VPWR_c_733_n 0.0118925f $X=-0.19 $Y=1.66 $X2=1.77 $Y2=1.565
cc_132 VPB N_VPWR_c_734_n 0.00586597f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_133 VPB N_VPWR_c_735_n 0.00838286f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_134 VPB N_VPWR_c_736_n 0.0206041f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_135 VPB N_VPWR_c_737_n 0.00324402f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_136 VPB N_VPWR_c_738_n 0.0206041f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_137 VPB N_VPWR_c_739_n 0.00324402f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_138 VPB N_VPWR_c_740_n 0.0206041f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_139 VPB N_VPWR_c_741_n 0.00324402f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_140 VPB N_VPWR_c_742_n 0.0206041f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_141 VPB N_VPWR_c_743_n 0.00324402f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_142 VPB N_VPWR_c_744_n 0.0206041f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_143 VPB N_VPWR_c_745_n 0.00324402f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_144 VPB N_VPWR_c_746_n 0.058109f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_145 VPB N_VPWR_c_747_n 0.0196495f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_146 VPB N_VPWR_c_748_n 0.0191515f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_147 VPB N_VPWR_c_724_n 0.121483f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_148 VPB N_VPWR_c_750_n 0.00614127f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_149 VPB N_VPWR_c_751_n 0.00489101f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_150 VPB N_VPWR_c_752_n 0.00391723f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_151 VPB N_Y_c_881_n 0.00257348f $X=-0.19 $Y=1.66 $X2=1.395 $Y2=2.4
cc_152 VPB N_Y_c_882_n 0.00179527f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_153 VPB N_Y_c_883_n 0.00183475f $X=-0.19 $Y=1.66 $X2=1.845 $Y2=1.765
cc_154 VPB N_Y_c_884_n 0.00216998f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_155 VPB N_Y_c_879_n 0.00245343f $X=-0.19 $Y=1.66 $X2=0.945 $Y2=1.557
cc_156 VPB N_Y_c_886_n 0.0120271f $X=-0.19 $Y=1.66 $X2=1.365 $Y2=1.557
cc_157 VPB N_Y_c_887_n 0.0027601f $X=-0.19 $Y=1.66 $X2=1.395 $Y2=1.557
cc_158 VPB N_A_1215_368#_c_988_n 0.00591568f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_159 VPB N_A_1215_368#_c_989_n 0.0028338f $X=-0.19 $Y=1.66 $X2=1.395 $Y2=2.4
cc_160 VPB N_A_1215_368#_c_990_n 0.00391405f $X=-0.19 $Y=1.66 $X2=1.395 $Y2=2.4
cc_161 VPB N_A_1215_368#_c_991_n 0.00527877f $X=-0.19 $Y=1.66 $X2=1.845
+ $Y2=1.765
cc_162 VPB N_A_1215_368#_c_992_n 0.00257348f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_163 VPB N_A_1215_368#_c_993_n 0.00802076f $X=-0.19 $Y=1.66 $X2=0.495
+ $Y2=1.557
cc_164 VPB N_A_1215_368#_c_994_n 0.0357063f $X=-0.19 $Y=1.66 $X2=0.945 $Y2=1.557
cc_165 VPB N_A_1215_368#_c_995_n 0.00145593f $X=-0.19 $Y=1.66 $X2=1.395
+ $Y2=1.557
cc_166 N_A1_N_M1034_g N_A2_N_M1006_g 0.0189918f $X=1.795 $Y=0.74 $X2=0 $Y2=0
cc_167 N_A1_N_c_176_n N_A2_N_c_257_n 0.025113f $X=1.845 $Y=1.765 $X2=0 $Y2=0
cc_168 N_A1_N_c_171_n N_A2_N_c_254_n 0.0016977f $X=1.77 $Y=1.515 $X2=0 $Y2=0
cc_169 N_A1_N_c_172_n N_A2_N_c_254_n 0.025232f $X=1.795 $Y=1.557 $X2=0 $Y2=0
cc_170 N_A1_N_c_171_n A2_N 0.0235847f $X=1.77 $Y=1.515 $X2=0 $Y2=0
cc_171 N_A1_N_c_172_n A2_N 4.71205e-19 $X=1.795 $Y=1.557 $X2=0 $Y2=0
cc_172 N_A1_N_c_173_n N_A_114_368#_c_365_n 0.00203651f $X=0.495 $Y=1.765 $X2=0
+ $Y2=0
cc_173 N_A1_N_c_174_n N_A_114_368#_c_365_n 4.27055e-19 $X=0.945 $Y=1.765 $X2=0
+ $Y2=0
cc_174 N_A1_N_c_171_n N_A_114_368#_c_365_n 0.0237598f $X=1.77 $Y=1.515 $X2=0
+ $Y2=0
cc_175 N_A1_N_c_172_n N_A_114_368#_c_365_n 0.00144162f $X=1.795 $Y=1.557 $X2=0
+ $Y2=0
cc_176 N_A1_N_c_173_n N_A_114_368#_c_360_n 0.00979955f $X=0.495 $Y=1.765 $X2=0
+ $Y2=0
cc_177 N_A1_N_c_174_n N_A_114_368#_c_360_n 0.0105344f $X=0.945 $Y=1.765 $X2=0
+ $Y2=0
cc_178 N_A1_N_c_175_n N_A_114_368#_c_360_n 6.45594e-19 $X=1.395 $Y=1.765 $X2=0
+ $Y2=0
cc_179 N_A1_N_c_174_n N_A_114_368#_c_372_n 0.0120074f $X=0.945 $Y=1.765 $X2=0
+ $Y2=0
cc_180 N_A1_N_c_175_n N_A_114_368#_c_372_n 0.0120074f $X=1.395 $Y=1.765 $X2=0
+ $Y2=0
cc_181 N_A1_N_c_171_n N_A_114_368#_c_372_n 0.0393875f $X=1.77 $Y=1.515 $X2=0
+ $Y2=0
cc_182 N_A1_N_c_172_n N_A_114_368#_c_372_n 0.0013093f $X=1.795 $Y=1.557 $X2=0
+ $Y2=0
cc_183 N_A1_N_c_174_n N_A_114_368#_c_361_n 6.45594e-19 $X=0.945 $Y=1.765 $X2=0
+ $Y2=0
cc_184 N_A1_N_c_175_n N_A_114_368#_c_361_n 0.0105344f $X=1.395 $Y=1.765 $X2=0
+ $Y2=0
cc_185 N_A1_N_c_176_n N_A_114_368#_c_361_n 0.0105344f $X=1.845 $Y=1.765 $X2=0
+ $Y2=0
cc_186 N_A1_N_c_176_n N_A_114_368#_c_379_n 0.0119563f $X=1.845 $Y=1.765 $X2=0
+ $Y2=0
cc_187 N_A1_N_c_171_n N_A_114_368#_c_379_n 0.0104662f $X=1.77 $Y=1.515 $X2=0
+ $Y2=0
cc_188 N_A1_N_c_176_n N_A_114_368#_c_362_n 6.45594e-19 $X=1.845 $Y=1.765 $X2=0
+ $Y2=0
cc_189 N_A1_N_c_175_n N_A_114_368#_c_382_n 4.27055e-19 $X=1.395 $Y=1.765 $X2=0
+ $Y2=0
cc_190 N_A1_N_c_176_n N_A_114_368#_c_382_n 4.27055e-19 $X=1.845 $Y=1.765 $X2=0
+ $Y2=0
cc_191 N_A1_N_c_171_n N_A_114_368#_c_382_n 0.0237598f $X=1.77 $Y=1.515 $X2=0
+ $Y2=0
cc_192 N_A1_N_c_172_n N_A_114_368#_c_382_n 0.00144162f $X=1.795 $Y=1.557 $X2=0
+ $Y2=0
cc_193 N_A1_N_c_173_n N_VPWR_c_726_n 0.00831454f $X=0.495 $Y=1.765 $X2=0 $Y2=0
cc_194 N_A1_N_c_171_n N_VPWR_c_726_n 0.0202607f $X=1.77 $Y=1.515 $X2=0 $Y2=0
cc_195 N_A1_N_c_172_n N_VPWR_c_726_n 6.71896e-19 $X=1.795 $Y=1.557 $X2=0 $Y2=0
cc_196 N_A1_N_c_174_n N_VPWR_c_727_n 0.00486623f $X=0.945 $Y=1.765 $X2=0 $Y2=0
cc_197 N_A1_N_c_175_n N_VPWR_c_727_n 0.00486623f $X=1.395 $Y=1.765 $X2=0 $Y2=0
cc_198 N_A1_N_c_176_n N_VPWR_c_728_n 0.00486623f $X=1.845 $Y=1.765 $X2=0 $Y2=0
cc_199 N_A1_N_c_173_n N_VPWR_c_736_n 0.00445602f $X=0.495 $Y=1.765 $X2=0 $Y2=0
cc_200 N_A1_N_c_174_n N_VPWR_c_736_n 0.00445602f $X=0.945 $Y=1.765 $X2=0 $Y2=0
cc_201 N_A1_N_c_175_n N_VPWR_c_738_n 0.00445602f $X=1.395 $Y=1.765 $X2=0 $Y2=0
cc_202 N_A1_N_c_176_n N_VPWR_c_738_n 0.00445602f $X=1.845 $Y=1.765 $X2=0 $Y2=0
cc_203 N_A1_N_c_173_n N_VPWR_c_724_n 0.0086105f $X=0.495 $Y=1.765 $X2=0 $Y2=0
cc_204 N_A1_N_c_174_n N_VPWR_c_724_n 0.00857589f $X=0.945 $Y=1.765 $X2=0 $Y2=0
cc_205 N_A1_N_c_175_n N_VPWR_c_724_n 0.00857589f $X=1.395 $Y=1.765 $X2=0 $Y2=0
cc_206 N_A1_N_c_176_n N_VPWR_c_724_n 0.00857673f $X=1.845 $Y=1.765 $X2=0 $Y2=0
cc_207 N_A1_N_M1009_g N_A_27_74#_c_1054_n 0.00159319f $X=0.495 $Y=0.74 $X2=0
+ $Y2=0
cc_208 N_A1_N_M1009_g N_A_27_74#_c_1055_n 0.0136535f $X=0.495 $Y=0.74 $X2=0
+ $Y2=0
cc_209 N_A1_N_M1032_g N_A_27_74#_c_1055_n 0.0131164f $X=0.925 $Y=0.74 $X2=0
+ $Y2=0
cc_210 N_A1_N_c_171_n N_A_27_74#_c_1055_n 0.0517333f $X=1.77 $Y=1.515 $X2=0
+ $Y2=0
cc_211 N_A1_N_c_172_n N_A_27_74#_c_1055_n 0.00348928f $X=1.795 $Y=1.557 $X2=0
+ $Y2=0
cc_212 N_A1_N_c_171_n N_A_27_74#_c_1056_n 0.0211272f $X=1.77 $Y=1.515 $X2=0
+ $Y2=0
cc_213 N_A1_N_c_172_n N_A_27_74#_c_1056_n 0.00279548f $X=1.795 $Y=1.557 $X2=0
+ $Y2=0
cc_214 N_A1_N_M1032_g N_A_27_74#_c_1057_n 4.03599e-19 $X=0.925 $Y=0.74 $X2=0
+ $Y2=0
cc_215 N_A1_N_M1033_g N_A_27_74#_c_1057_n 4.03599e-19 $X=1.365 $Y=0.74 $X2=0
+ $Y2=0
cc_216 N_A1_N_M1033_g N_A_27_74#_c_1058_n 0.0130699f $X=1.365 $Y=0.74 $X2=0
+ $Y2=0
cc_217 N_A1_N_M1034_g N_A_27_74#_c_1058_n 0.0128967f $X=1.795 $Y=0.74 $X2=0
+ $Y2=0
cc_218 N_A1_N_c_171_n N_A_27_74#_c_1058_n 0.0525922f $X=1.77 $Y=1.515 $X2=0
+ $Y2=0
cc_219 N_A1_N_c_172_n N_A_27_74#_c_1058_n 0.00391924f $X=1.795 $Y=1.557 $X2=0
+ $Y2=0
cc_220 N_A1_N_M1034_g N_A_27_74#_c_1060_n 9.48753e-19 $X=1.795 $Y=0.74 $X2=0
+ $Y2=0
cc_221 N_A1_N_c_171_n N_A_27_74#_c_1063_n 0.0154618f $X=1.77 $Y=1.515 $X2=0
+ $Y2=0
cc_222 N_A1_N_c_172_n N_A_27_74#_c_1063_n 0.00256252f $X=1.795 $Y=1.557 $X2=0
+ $Y2=0
cc_223 N_A1_N_M1009_g N_VGND_c_1122_n 0.0133724f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_224 N_A1_N_M1032_g N_VGND_c_1122_n 0.0103611f $X=0.925 $Y=0.74 $X2=0 $Y2=0
cc_225 N_A1_N_M1033_g N_VGND_c_1122_n 4.7018e-19 $X=1.365 $Y=0.74 $X2=0 $Y2=0
cc_226 N_A1_N_M1032_g N_VGND_c_1123_n 4.7018e-19 $X=0.925 $Y=0.74 $X2=0 $Y2=0
cc_227 N_A1_N_M1033_g N_VGND_c_1123_n 0.0103611f $X=1.365 $Y=0.74 $X2=0 $Y2=0
cc_228 N_A1_N_M1034_g N_VGND_c_1123_n 0.00968343f $X=1.795 $Y=0.74 $X2=0 $Y2=0
cc_229 N_A1_N_M1034_g N_VGND_c_1124_n 0.00383152f $X=1.795 $Y=0.74 $X2=0 $Y2=0
cc_230 N_A1_N_M1009_g N_VGND_c_1129_n 0.00383152f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_231 N_A1_N_M1032_g N_VGND_c_1130_n 0.00383152f $X=0.925 $Y=0.74 $X2=0 $Y2=0
cc_232 N_A1_N_M1033_g N_VGND_c_1130_n 0.00383152f $X=1.365 $Y=0.74 $X2=0 $Y2=0
cc_233 N_A1_N_M1009_g N_VGND_c_1135_n 0.00761198f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_234 N_A1_N_M1032_g N_VGND_c_1135_n 0.0075764f $X=0.925 $Y=0.74 $X2=0 $Y2=0
cc_235 N_A1_N_M1033_g N_VGND_c_1135_n 0.0075764f $X=1.365 $Y=0.74 $X2=0 $Y2=0
cc_236 N_A1_N_M1034_g N_VGND_c_1135_n 0.00757637f $X=1.795 $Y=0.74 $X2=0 $Y2=0
cc_237 N_A2_N_c_255_n N_A_114_368#_c_355_n 0.00861049f $X=3.645 $Y=1.765 $X2=0
+ $Y2=0
cc_238 N_A2_N_c_255_n N_A_114_368#_c_349_n 0.0141027f $X=3.645 $Y=1.765 $X2=0
+ $Y2=0
cc_239 N_A2_N_M1039_g N_A_114_368#_c_349_n 0.00590113f $X=3.655 $Y=0.74 $X2=0
+ $Y2=0
cc_240 N_A2_N_c_257_n N_A_114_368#_c_361_n 6.45594e-19 $X=2.295 $Y=1.765 $X2=0
+ $Y2=0
cc_241 N_A2_N_c_257_n N_A_114_368#_c_379_n 0.012109f $X=2.295 $Y=1.765 $X2=0
+ $Y2=0
cc_242 N_A2_N_c_254_n N_A_114_368#_c_379_n 0.00139665f $X=3.285 $Y=1.395 $X2=0
+ $Y2=0
cc_243 A2_N N_A_114_368#_c_379_n 0.00945133f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_244 N_A2_N_M1006_g N_A_114_368#_c_393_n 0.00498003f $X=2.225 $Y=0.74 $X2=0
+ $Y2=0
cc_245 N_A2_N_M1013_g N_A_114_368#_c_393_n 0.00661392f $X=2.655 $Y=0.74 $X2=0
+ $Y2=0
cc_246 N_A2_N_M1021_g N_A_114_368#_c_393_n 5.87434e-19 $X=3.18 $Y=0.74 $X2=0
+ $Y2=0
cc_247 N_A2_N_c_257_n N_A_114_368#_c_362_n 0.0105344f $X=2.295 $Y=1.765 $X2=0
+ $Y2=0
cc_248 N_A2_N_c_258_n N_A_114_368#_c_362_n 0.0105344f $X=2.745 $Y=1.765 $X2=0
+ $Y2=0
cc_249 N_A2_N_c_259_n N_A_114_368#_c_362_n 6.45594e-19 $X=3.195 $Y=1.765 $X2=0
+ $Y2=0
cc_250 N_A2_N_M1013_g N_A_114_368#_c_351_n 0.00952207f $X=2.655 $Y=0.74 $X2=0
+ $Y2=0
cc_251 N_A2_N_M1021_g N_A_114_368#_c_351_n 0.0132432f $X=3.18 $Y=0.74 $X2=0
+ $Y2=0
cc_252 N_A2_N_c_254_n N_A_114_368#_c_351_n 0.00462638f $X=3.285 $Y=1.395 $X2=0
+ $Y2=0
cc_253 A2_N N_A_114_368#_c_351_n 0.0473393f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_254 N_A2_N_M1006_g N_A_114_368#_c_352_n 0.00407645f $X=2.225 $Y=0.74 $X2=0
+ $Y2=0
cc_255 N_A2_N_M1013_g N_A_114_368#_c_352_n 0.00271614f $X=2.655 $Y=0.74 $X2=0
+ $Y2=0
cc_256 N_A2_N_c_254_n N_A_114_368#_c_352_n 0.00244236f $X=3.285 $Y=1.395 $X2=0
+ $Y2=0
cc_257 A2_N N_A_114_368#_c_352_n 0.027784f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_258 N_A2_N_c_258_n N_A_114_368#_c_407_n 0.0120074f $X=2.745 $Y=1.765 $X2=0
+ $Y2=0
cc_259 N_A2_N_c_259_n N_A_114_368#_c_407_n 0.0125877f $X=3.195 $Y=1.765 $X2=0
+ $Y2=0
cc_260 N_A2_N_c_254_n N_A_114_368#_c_407_n 0.00131281f $X=3.285 $Y=1.395 $X2=0
+ $Y2=0
cc_261 A2_N N_A_114_368#_c_407_n 0.0379621f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_262 N_A2_N_c_258_n N_A_114_368#_c_363_n 6.45594e-19 $X=2.745 $Y=1.765 $X2=0
+ $Y2=0
cc_263 N_A2_N_c_259_n N_A_114_368#_c_363_n 0.0105344f $X=3.195 $Y=1.765 $X2=0
+ $Y2=0
cc_264 N_A2_N_c_255_n N_A_114_368#_c_363_n 0.0092887f $X=3.645 $Y=1.765 $X2=0
+ $Y2=0
cc_265 N_A2_N_M1039_g N_A_114_368#_c_414_n 0.00567006f $X=3.655 $Y=0.74 $X2=0
+ $Y2=0
cc_266 N_A2_N_M1021_g N_A_114_368#_c_353_n 0.00319592f $X=3.18 $Y=0.74 $X2=0
+ $Y2=0
cc_267 N_A2_N_c_253_n N_A_114_368#_c_353_n 0.0114992f $X=3.555 $Y=1.395 $X2=0
+ $Y2=0
cc_268 N_A2_N_c_254_n N_A_114_368#_c_353_n 0.00135651f $X=3.285 $Y=1.395 $X2=0
+ $Y2=0
cc_269 N_A2_N_c_255_n N_A_114_368#_c_353_n 0.00360771f $X=3.645 $Y=1.765 $X2=0
+ $Y2=0
cc_270 N_A2_N_M1039_g N_A_114_368#_c_353_n 0.0115523f $X=3.655 $Y=0.74 $X2=0
+ $Y2=0
cc_271 A2_N N_A_114_368#_c_353_n 0.0232738f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_272 N_A2_N_c_259_n N_A_114_368#_c_364_n 0.00333846f $X=3.195 $Y=1.765 $X2=0
+ $Y2=0
cc_273 N_A2_N_c_254_n N_A_114_368#_c_364_n 8.94325e-19 $X=3.285 $Y=1.395 $X2=0
+ $Y2=0
cc_274 N_A2_N_c_255_n N_A_114_368#_c_364_n 0.0065214f $X=3.645 $Y=1.765 $X2=0
+ $Y2=0
cc_275 A2_N N_A_114_368#_c_364_n 0.0113235f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_276 N_A2_N_c_255_n N_A_114_368#_c_354_n 0.0137803f $X=3.645 $Y=1.765 $X2=0
+ $Y2=0
cc_277 N_A2_N_M1039_g N_A_114_368#_c_354_n 0.00637964f $X=3.655 $Y=0.74 $X2=0
+ $Y2=0
cc_278 N_A2_N_c_257_n N_A_114_368#_c_427_n 4.27055e-19 $X=2.295 $Y=1.765 $X2=0
+ $Y2=0
cc_279 N_A2_N_c_258_n N_A_114_368#_c_427_n 4.27055e-19 $X=2.745 $Y=1.765 $X2=0
+ $Y2=0
cc_280 N_A2_N_c_254_n N_A_114_368#_c_427_n 0.00144082f $X=3.285 $Y=1.395 $X2=0
+ $Y2=0
cc_281 A2_N N_A_114_368#_c_427_n 0.0237598f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_282 N_A2_N_c_259_n N_A_114_368#_c_431_n 9.50925e-19 $X=3.195 $Y=1.765 $X2=0
+ $Y2=0
cc_283 N_A2_N_c_253_n N_A_114_368#_c_431_n 0.00118718f $X=3.555 $Y=1.395 $X2=0
+ $Y2=0
cc_284 N_A2_N_c_255_n N_A_114_368#_c_431_n 0.0017329f $X=3.645 $Y=1.765 $X2=0
+ $Y2=0
cc_285 N_A2_N_c_257_n N_VPWR_c_728_n 0.00486623f $X=2.295 $Y=1.765 $X2=0 $Y2=0
cc_286 N_A2_N_c_258_n N_VPWR_c_729_n 0.00486623f $X=2.745 $Y=1.765 $X2=0 $Y2=0
cc_287 N_A2_N_c_259_n N_VPWR_c_729_n 0.00486623f $X=3.195 $Y=1.765 $X2=0 $Y2=0
cc_288 N_A2_N_c_255_n N_VPWR_c_730_n 0.00665298f $X=3.645 $Y=1.765 $X2=0 $Y2=0
cc_289 N_A2_N_c_257_n N_VPWR_c_740_n 0.00445602f $X=2.295 $Y=1.765 $X2=0 $Y2=0
cc_290 N_A2_N_c_258_n N_VPWR_c_740_n 0.00445602f $X=2.745 $Y=1.765 $X2=0 $Y2=0
cc_291 N_A2_N_c_259_n N_VPWR_c_742_n 0.00445602f $X=3.195 $Y=1.765 $X2=0 $Y2=0
cc_292 N_A2_N_c_255_n N_VPWR_c_742_n 0.00445602f $X=3.645 $Y=1.765 $X2=0 $Y2=0
cc_293 N_A2_N_c_257_n N_VPWR_c_724_n 0.00857673f $X=2.295 $Y=1.765 $X2=0 $Y2=0
cc_294 N_A2_N_c_258_n N_VPWR_c_724_n 0.00857589f $X=2.745 $Y=1.765 $X2=0 $Y2=0
cc_295 N_A2_N_c_259_n N_VPWR_c_724_n 0.00857589f $X=3.195 $Y=1.765 $X2=0 $Y2=0
cc_296 N_A2_N_c_255_n N_VPWR_c_724_n 0.00857673f $X=3.645 $Y=1.765 $X2=0 $Y2=0
cc_297 N_A2_N_M1006_g N_A_27_74#_c_1058_n 5.7448e-19 $X=2.225 $Y=0.74 $X2=0
+ $Y2=0
cc_298 N_A2_N_M1006_g N_A_27_74#_c_1059_n 0.0120041f $X=2.225 $Y=0.74 $X2=0
+ $Y2=0
cc_299 N_A2_N_M1013_g N_A_27_74#_c_1059_n 0.0112986f $X=2.655 $Y=0.74 $X2=0
+ $Y2=0
cc_300 N_A2_N_M1021_g N_A_27_74#_c_1061_n 0.00938114f $X=3.18 $Y=0.74 $X2=0
+ $Y2=0
cc_301 N_A2_N_M1039_g N_A_27_74#_c_1061_n 0.0135229f $X=3.655 $Y=0.74 $X2=0
+ $Y2=0
cc_302 N_A2_N_M1039_g N_A_27_74#_c_1062_n 0.00159289f $X=3.655 $Y=0.74 $X2=0
+ $Y2=0
cc_303 N_A2_N_M1021_g N_A_27_74#_c_1064_n 0.00217786f $X=3.18 $Y=0.74 $X2=0
+ $Y2=0
cc_304 N_A2_N_M1006_g N_VGND_c_1124_n 0.00278271f $X=2.225 $Y=0.74 $X2=0 $Y2=0
cc_305 N_A2_N_M1013_g N_VGND_c_1124_n 0.00278271f $X=2.655 $Y=0.74 $X2=0 $Y2=0
cc_306 N_A2_N_M1021_g N_VGND_c_1124_n 0.00278271f $X=3.18 $Y=0.74 $X2=0 $Y2=0
cc_307 N_A2_N_M1039_g N_VGND_c_1124_n 0.00278271f $X=3.655 $Y=0.74 $X2=0 $Y2=0
cc_308 N_A2_N_M1006_g N_VGND_c_1135_n 0.00353526f $X=2.225 $Y=0.74 $X2=0 $Y2=0
cc_309 N_A2_N_M1013_g N_VGND_c_1135_n 0.00354301f $X=2.655 $Y=0.74 $X2=0 $Y2=0
cc_310 N_A2_N_M1021_g N_VGND_c_1135_n 0.00354734f $X=3.18 $Y=0.74 $X2=0 $Y2=0
cc_311 N_A2_N_M1039_g N_VGND_c_1135_n 0.0035886f $X=3.655 $Y=0.74 $X2=0 $Y2=0
cc_312 N_A2_N_M1039_g N_A_857_74#_c_1253_n 5.96586e-19 $X=3.655 $Y=0.74 $X2=0
+ $Y2=0
cc_313 N_A_114_368#_M1030_g N_B2_M1000_g 0.0115453f $X=5.935 $Y=0.74 $X2=0 $Y2=0
cc_314 N_A_114_368#_c_348_n N_B2_c_556_n 0.0125083f $X=5.86 $Y=1.375 $X2=0 $Y2=0
cc_315 N_A_114_368#_c_349_n N_B2_c_556_n 5.44913e-19 $X=5.58 $Y=1.375 $X2=0
+ $Y2=0
cc_316 N_A_114_368#_c_348_n N_B2_c_557_n 0.0115453f $X=5.86 $Y=1.375 $X2=0 $Y2=0
cc_317 N_A_114_368#_c_349_n N_B2_c_557_n 0.00141988f $X=5.58 $Y=1.375 $X2=0
+ $Y2=0
cc_318 N_A_114_368#_c_372_n N_VPWR_M1002_s 0.00408911f $X=1.455 $Y=2.035 $X2=0
+ $Y2=0
cc_319 N_A_114_368#_c_379_n N_VPWR_M1008_s 0.00923646f $X=2.355 $Y=2.035 $X2=0
+ $Y2=0
cc_320 N_A_114_368#_c_407_n N_VPWR_M1014_s 0.00408911f $X=3.255 $Y=2.035 $X2=0
+ $Y2=0
cc_321 N_A_114_368#_c_365_n N_VPWR_c_726_n 0.0121024f $X=0.72 $Y=2.12 $X2=0
+ $Y2=0
cc_322 N_A_114_368#_c_360_n N_VPWR_c_726_n 0.0576605f $X=0.72 $Y=2.815 $X2=0
+ $Y2=0
cc_323 N_A_114_368#_c_360_n N_VPWR_c_727_n 0.0449718f $X=0.72 $Y=2.815 $X2=0
+ $Y2=0
cc_324 N_A_114_368#_c_372_n N_VPWR_c_727_n 0.0136682f $X=1.455 $Y=2.035 $X2=0
+ $Y2=0
cc_325 N_A_114_368#_c_361_n N_VPWR_c_727_n 0.0449718f $X=1.62 $Y=2.815 $X2=0
+ $Y2=0
cc_326 N_A_114_368#_c_361_n N_VPWR_c_728_n 0.0449718f $X=1.62 $Y=2.815 $X2=0
+ $Y2=0
cc_327 N_A_114_368#_c_379_n N_VPWR_c_728_n 0.0136682f $X=2.355 $Y=2.035 $X2=0
+ $Y2=0
cc_328 N_A_114_368#_c_362_n N_VPWR_c_728_n 0.0449718f $X=2.52 $Y=2.815 $X2=0
+ $Y2=0
cc_329 N_A_114_368#_c_362_n N_VPWR_c_729_n 0.0449718f $X=2.52 $Y=2.815 $X2=0
+ $Y2=0
cc_330 N_A_114_368#_c_407_n N_VPWR_c_729_n 0.0136682f $X=3.255 $Y=2.035 $X2=0
+ $Y2=0
cc_331 N_A_114_368#_c_363_n N_VPWR_c_729_n 0.0449718f $X=3.42 $Y=2.815 $X2=0
+ $Y2=0
cc_332 N_A_114_368#_c_355_n N_VPWR_c_730_n 0.00665327f $X=4.095 $Y=1.765 $X2=0
+ $Y2=0
cc_333 N_A_114_368#_c_363_n N_VPWR_c_730_n 0.0560121f $X=3.42 $Y=2.815 $X2=0
+ $Y2=0
cc_334 N_A_114_368#_c_364_n N_VPWR_c_730_n 0.00805078f $X=3.5 $Y=1.95 $X2=0
+ $Y2=0
cc_335 N_A_114_368#_c_354_n N_VPWR_c_730_n 0.0137368f $X=5.26 $Y=1.465 $X2=0
+ $Y2=0
cc_336 N_A_114_368#_c_431_n N_VPWR_c_730_n 0.0117758f $X=3.42 $Y=2.035 $X2=0
+ $Y2=0
cc_337 N_A_114_368#_c_356_n N_VPWR_c_731_n 0.00586501f $X=4.545 $Y=1.765 $X2=0
+ $Y2=0
cc_338 N_A_114_368#_c_357_n N_VPWR_c_731_n 0.00466569f $X=4.995 $Y=1.765 $X2=0
+ $Y2=0
cc_339 N_A_114_368#_c_357_n N_VPWR_c_732_n 0.00445602f $X=4.995 $Y=1.765 $X2=0
+ $Y2=0
cc_340 N_A_114_368#_c_358_n N_VPWR_c_732_n 0.00413917f $X=5.445 $Y=1.765 $X2=0
+ $Y2=0
cc_341 N_A_114_368#_c_357_n N_VPWR_c_733_n 5.57166e-19 $X=4.995 $Y=1.765 $X2=0
+ $Y2=0
cc_342 N_A_114_368#_c_358_n N_VPWR_c_733_n 0.0122524f $X=5.445 $Y=1.765 $X2=0
+ $Y2=0
cc_343 N_A_114_368#_c_360_n N_VPWR_c_736_n 0.014552f $X=0.72 $Y=2.815 $X2=0
+ $Y2=0
cc_344 N_A_114_368#_c_361_n N_VPWR_c_738_n 0.014552f $X=1.62 $Y=2.815 $X2=0
+ $Y2=0
cc_345 N_A_114_368#_c_362_n N_VPWR_c_740_n 0.014552f $X=2.52 $Y=2.815 $X2=0
+ $Y2=0
cc_346 N_A_114_368#_c_363_n N_VPWR_c_742_n 0.014552f $X=3.42 $Y=2.815 $X2=0
+ $Y2=0
cc_347 N_A_114_368#_c_355_n N_VPWR_c_744_n 0.00445602f $X=4.095 $Y=1.765 $X2=0
+ $Y2=0
cc_348 N_A_114_368#_c_356_n N_VPWR_c_744_n 0.00445602f $X=4.545 $Y=1.765 $X2=0
+ $Y2=0
cc_349 N_A_114_368#_c_355_n N_VPWR_c_724_n 0.00857673f $X=4.095 $Y=1.765 $X2=0
+ $Y2=0
cc_350 N_A_114_368#_c_356_n N_VPWR_c_724_n 0.00857589f $X=4.545 $Y=1.765 $X2=0
+ $Y2=0
cc_351 N_A_114_368#_c_357_n N_VPWR_c_724_n 0.00857589f $X=4.995 $Y=1.765 $X2=0
+ $Y2=0
cc_352 N_A_114_368#_c_358_n N_VPWR_c_724_n 0.00817726f $X=5.445 $Y=1.765 $X2=0
+ $Y2=0
cc_353 N_A_114_368#_c_360_n N_VPWR_c_724_n 0.0119791f $X=0.72 $Y=2.815 $X2=0
+ $Y2=0
cc_354 N_A_114_368#_c_361_n N_VPWR_c_724_n 0.0119791f $X=1.62 $Y=2.815 $X2=0
+ $Y2=0
cc_355 N_A_114_368#_c_362_n N_VPWR_c_724_n 0.0119791f $X=2.52 $Y=2.815 $X2=0
+ $Y2=0
cc_356 N_A_114_368#_c_363_n N_VPWR_c_724_n 0.0119791f $X=3.42 $Y=2.815 $X2=0
+ $Y2=0
cc_357 N_A_114_368#_c_355_n N_Y_c_881_n 0.0112572f $X=4.095 $Y=1.765 $X2=0 $Y2=0
cc_358 N_A_114_368#_c_356_n N_Y_c_881_n 0.0125003f $X=4.545 $Y=1.765 $X2=0 $Y2=0
cc_359 N_A_114_368#_c_357_n N_Y_c_881_n 6.91e-19 $X=4.995 $Y=1.765 $X2=0 $Y2=0
cc_360 N_A_114_368#_c_356_n N_Y_c_882_n 0.0120074f $X=4.545 $Y=1.765 $X2=0 $Y2=0
cc_361 N_A_114_368#_c_357_n N_Y_c_882_n 0.0120074f $X=4.995 $Y=1.765 $X2=0 $Y2=0
cc_362 N_A_114_368#_c_349_n N_Y_c_882_n 0.00765693f $X=5.58 $Y=1.375 $X2=0 $Y2=0
cc_363 N_A_114_368#_c_354_n N_Y_c_882_n 0.0417603f $X=5.26 $Y=1.465 $X2=0 $Y2=0
cc_364 N_A_114_368#_c_355_n N_Y_c_883_n 0.00259534f $X=4.095 $Y=1.765 $X2=0
+ $Y2=0
cc_365 N_A_114_368#_c_356_n N_Y_c_883_n 9.3899e-19 $X=4.545 $Y=1.765 $X2=0 $Y2=0
cc_366 N_A_114_368#_c_349_n N_Y_c_883_n 0.00717196f $X=5.58 $Y=1.375 $X2=0 $Y2=0
cc_367 N_A_114_368#_c_364_n N_Y_c_883_n 5.60583e-19 $X=3.5 $Y=1.95 $X2=0 $Y2=0
cc_368 N_A_114_368#_c_354_n N_Y_c_883_n 0.0276943f $X=5.26 $Y=1.465 $X2=0 $Y2=0
cc_369 N_A_114_368#_M1007_g N_Y_c_900_n 0.00515339f $X=4.645 $Y=0.74 $X2=0 $Y2=0
cc_370 N_A_114_368#_M1016_g N_Y_c_900_n 0.00611761f $X=5.075 $Y=0.74 $X2=0 $Y2=0
cc_371 N_A_114_368#_M1022_g N_Y_c_900_n 5.55764e-19 $X=5.505 $Y=0.74 $X2=0 $Y2=0
cc_372 N_A_114_368#_M1016_g N_Y_c_877_n 0.00885064f $X=5.075 $Y=0.74 $X2=0 $Y2=0
cc_373 N_A_114_368#_M1022_g N_Y_c_877_n 0.00992864f $X=5.505 $Y=0.74 $X2=0 $Y2=0
cc_374 N_A_114_368#_c_349_n N_Y_c_877_n 0.00224206f $X=5.58 $Y=1.375 $X2=0 $Y2=0
cc_375 N_A_114_368#_c_354_n N_Y_c_877_n 0.0258049f $X=5.26 $Y=1.465 $X2=0 $Y2=0
cc_376 N_A_114_368#_M1007_g N_Y_c_878_n 0.00310933f $X=4.645 $Y=0.74 $X2=0 $Y2=0
cc_377 N_A_114_368#_M1016_g N_Y_c_878_n 0.00163137f $X=5.075 $Y=0.74 $X2=0 $Y2=0
cc_378 N_A_114_368#_c_349_n N_Y_c_878_n 0.00231784f $X=5.58 $Y=1.375 $X2=0 $Y2=0
cc_379 N_A_114_368#_c_354_n N_Y_c_878_n 0.0270731f $X=5.26 $Y=1.465 $X2=0 $Y2=0
cc_380 N_A_114_368#_c_357_n N_Y_c_884_n 0.0092272f $X=4.995 $Y=1.765 $X2=0 $Y2=0
cc_381 N_A_114_368#_c_358_n N_Y_c_884_n 0.00617286f $X=5.445 $Y=1.765 $X2=0
+ $Y2=0
cc_382 N_A_114_368#_M1016_g N_Y_c_913_n 5.64138e-19 $X=5.075 $Y=0.74 $X2=0 $Y2=0
cc_383 N_A_114_368#_M1022_g N_Y_c_913_n 0.00646632f $X=5.505 $Y=0.74 $X2=0 $Y2=0
cc_384 N_A_114_368#_M1030_g N_Y_c_913_n 0.00494352f $X=5.935 $Y=0.74 $X2=0 $Y2=0
cc_385 N_A_114_368#_M1016_g N_Y_c_879_n 8.44792e-19 $X=5.075 $Y=0.74 $X2=0 $Y2=0
cc_386 N_A_114_368#_c_358_n N_Y_c_879_n 0.001364f $X=5.445 $Y=1.765 $X2=0 $Y2=0
cc_387 N_A_114_368#_M1022_g N_Y_c_879_n 0.00419028f $X=5.505 $Y=0.74 $X2=0 $Y2=0
cc_388 N_A_114_368#_c_348_n N_Y_c_879_n 0.00830694f $X=5.86 $Y=1.375 $X2=0 $Y2=0
cc_389 N_A_114_368#_c_349_n N_Y_c_879_n 0.0144772f $X=5.58 $Y=1.375 $X2=0 $Y2=0
cc_390 N_A_114_368#_M1030_g N_Y_c_879_n 0.00294584f $X=5.935 $Y=0.74 $X2=0 $Y2=0
cc_391 N_A_114_368#_c_354_n N_Y_c_879_n 0.0250936f $X=5.26 $Y=1.465 $X2=0 $Y2=0
cc_392 N_A_114_368#_c_348_n N_Y_c_886_n 0.00510836f $X=5.86 $Y=1.375 $X2=0 $Y2=0
cc_393 N_A_114_368#_c_356_n N_Y_c_887_n 4.37811e-19 $X=4.545 $Y=1.765 $X2=0
+ $Y2=0
cc_394 N_A_114_368#_c_357_n N_Y_c_887_n 0.00401618f $X=4.995 $Y=1.765 $X2=0
+ $Y2=0
cc_395 N_A_114_368#_c_358_n N_Y_c_887_n 0.0236248f $X=5.445 $Y=1.765 $X2=0 $Y2=0
cc_396 N_A_114_368#_c_349_n N_Y_c_887_n 0.00878722f $X=5.58 $Y=1.375 $X2=0 $Y2=0
cc_397 N_A_114_368#_c_354_n N_Y_c_887_n 0.0265878f $X=5.26 $Y=1.465 $X2=0 $Y2=0
cc_398 N_A_114_368#_M1022_g N_Y_c_880_n 0.00144713f $X=5.505 $Y=0.74 $X2=0 $Y2=0
cc_399 N_A_114_368#_c_348_n N_Y_c_880_n 0.00217378f $X=5.86 $Y=1.375 $X2=0 $Y2=0
cc_400 N_A_114_368#_M1030_g N_Y_c_880_n 0.00375789f $X=5.935 $Y=0.74 $X2=0 $Y2=0
cc_401 N_A_114_368#_c_358_n N_A_1215_368#_c_988_n 9.45414e-19 $X=5.445 $Y=1.765
+ $X2=0 $Y2=0
cc_402 N_A_114_368#_c_358_n N_A_1215_368#_c_990_n 5.85502e-19 $X=5.445 $Y=1.765
+ $X2=0 $Y2=0
cc_403 N_A_114_368#_c_351_n N_A_27_74#_M1013_d 0.00285668f $X=3.275 $Y=1.095
+ $X2=0 $Y2=0
cc_404 N_A_114_368#_c_352_n N_A_27_74#_c_1058_n 0.00997012f $X=2.605 $Y=1.095
+ $X2=0 $Y2=0
cc_405 N_A_114_368#_M1006_s N_A_27_74#_c_1059_n 0.00176461f $X=2.3 $Y=0.37 $X2=0
+ $Y2=0
cc_406 N_A_114_368#_c_393_n N_A_27_74#_c_1059_n 0.0158692f $X=2.44 $Y=0.82 $X2=0
+ $Y2=0
cc_407 N_A_114_368#_c_351_n N_A_27_74#_c_1059_n 0.00304353f $X=3.275 $Y=1.095
+ $X2=0 $Y2=0
cc_408 N_A_114_368#_c_351_n N_A_27_74#_c_1093_n 0.020976f $X=3.275 $Y=1.095
+ $X2=0 $Y2=0
cc_409 N_A_114_368#_M1021_s N_A_27_74#_c_1061_n 0.00224297f $X=3.255 $Y=0.37
+ $X2=0 $Y2=0
cc_410 N_A_114_368#_M1007_g N_A_27_74#_c_1061_n 5.96586e-19 $X=4.645 $Y=0.74
+ $X2=0 $Y2=0
cc_411 N_A_114_368#_c_351_n N_A_27_74#_c_1061_n 0.00364245f $X=3.275 $Y=1.095
+ $X2=0 $Y2=0
cc_412 N_A_114_368#_c_414_n N_A_27_74#_c_1061_n 0.0176798f $X=3.44 $Y=0.86 $X2=0
+ $Y2=0
cc_413 N_A_114_368#_c_353_n N_A_27_74#_c_1062_n 0.00555794f $X=3.5 $Y=1.63 $X2=0
+ $Y2=0
cc_414 N_A_114_368#_c_354_n N_A_27_74#_c_1062_n 0.0219383f $X=5.26 $Y=1.465
+ $X2=0 $Y2=0
cc_415 N_A_114_368#_M1007_g N_VGND_c_1124_n 0.00278271f $X=4.645 $Y=0.74 $X2=0
+ $Y2=0
cc_416 N_A_114_368#_M1016_g N_VGND_c_1124_n 0.00278271f $X=5.075 $Y=0.74 $X2=0
+ $Y2=0
cc_417 N_A_114_368#_M1022_g N_VGND_c_1124_n 0.00278271f $X=5.505 $Y=0.74 $X2=0
+ $Y2=0
cc_418 N_A_114_368#_M1030_g N_VGND_c_1124_n 0.00278271f $X=5.935 $Y=0.74 $X2=0
+ $Y2=0
cc_419 N_A_114_368#_M1007_g N_VGND_c_1135_n 0.00358427f $X=4.645 $Y=0.74 $X2=0
+ $Y2=0
cc_420 N_A_114_368#_M1016_g N_VGND_c_1135_n 0.00353428f $X=5.075 $Y=0.74 $X2=0
+ $Y2=0
cc_421 N_A_114_368#_M1022_g N_VGND_c_1135_n 0.00353428f $X=5.505 $Y=0.74 $X2=0
+ $Y2=0
cc_422 N_A_114_368#_M1030_g N_VGND_c_1135_n 0.00353526f $X=5.935 $Y=0.74 $X2=0
+ $Y2=0
cc_423 N_A_114_368#_M1007_g N_A_857_74#_c_1251_n 0.00159289f $X=4.645 $Y=0.74
+ $X2=0 $Y2=0
cc_424 N_A_114_368#_c_349_n N_A_857_74#_c_1251_n 0.00597558f $X=5.58 $Y=1.375
+ $X2=0 $Y2=0
cc_425 N_A_114_368#_c_354_n N_A_857_74#_c_1251_n 0.0209147f $X=5.26 $Y=1.465
+ $X2=0 $Y2=0
cc_426 N_A_114_368#_M1007_g N_A_857_74#_c_1252_n 0.0132617f $X=4.645 $Y=0.74
+ $X2=0 $Y2=0
cc_427 N_A_114_368#_M1016_g N_A_857_74#_c_1252_n 0.0100569f $X=5.075 $Y=0.74
+ $X2=0 $Y2=0
cc_428 N_A_114_368#_M1022_g N_A_857_74#_c_1254_n 0.00988997f $X=5.505 $Y=0.74
+ $X2=0 $Y2=0
cc_429 N_A_114_368#_M1030_g N_A_857_74#_c_1254_n 0.0120041f $X=5.935 $Y=0.74
+ $X2=0 $Y2=0
cc_430 N_A_114_368#_M1030_g N_A_857_74#_c_1256_n 7.38995e-19 $X=5.935 $Y=0.74
+ $X2=0 $Y2=0
cc_431 N_B2_M1037_g N_B1_M1005_g 0.0195038f $X=7.795 $Y=0.74 $X2=0 $Y2=0
cc_432 N_B2_c_561_n N_B1_c_649_n 0.0120684f $X=7.785 $Y=1.765 $X2=0 $Y2=0
cc_433 N_B2_c_556_n B1 0.0151763f $X=7.475 $Y=1.515 $X2=0 $Y2=0
cc_434 N_B2_c_557_n B1 0.0019406f $X=7.785 $Y=1.557 $X2=0 $Y2=0
cc_435 N_B2_c_556_n N_B1_c_648_n 6.26242e-19 $X=7.475 $Y=1.515 $X2=0 $Y2=0
cc_436 N_B2_c_557_n N_B1_c_648_n 0.0203273f $X=7.785 $Y=1.557 $X2=0 $Y2=0
cc_437 N_B2_c_558_n N_VPWR_c_733_n 8.69902e-19 $X=6.435 $Y=1.765 $X2=0 $Y2=0
cc_438 N_B2_c_558_n N_VPWR_c_746_n 0.00278271f $X=6.435 $Y=1.765 $X2=0 $Y2=0
cc_439 N_B2_c_559_n N_VPWR_c_746_n 0.00278271f $X=6.885 $Y=1.765 $X2=0 $Y2=0
cc_440 N_B2_c_560_n N_VPWR_c_746_n 0.00278271f $X=7.335 $Y=1.765 $X2=0 $Y2=0
cc_441 N_B2_c_561_n N_VPWR_c_746_n 0.00278271f $X=7.785 $Y=1.765 $X2=0 $Y2=0
cc_442 N_B2_c_558_n N_VPWR_c_724_n 0.00358624f $X=6.435 $Y=1.765 $X2=0 $Y2=0
cc_443 N_B2_c_559_n N_VPWR_c_724_n 0.00353823f $X=6.885 $Y=1.765 $X2=0 $Y2=0
cc_444 N_B2_c_560_n N_VPWR_c_724_n 0.00353823f $X=7.335 $Y=1.765 $X2=0 $Y2=0
cc_445 N_B2_c_561_n N_VPWR_c_724_n 0.00353907f $X=7.785 $Y=1.765 $X2=0 $Y2=0
cc_446 N_B2_c_558_n N_Y_c_879_n 4.66361e-19 $X=6.435 $Y=1.765 $X2=0 $Y2=0
cc_447 N_B2_c_556_n N_Y_c_879_n 0.035327f $X=7.475 $Y=1.515 $X2=0 $Y2=0
cc_448 N_B2_c_557_n N_Y_c_879_n 7.82002e-19 $X=7.785 $Y=1.557 $X2=0 $Y2=0
cc_449 N_B2_c_558_n N_Y_c_886_n 0.0139279f $X=6.435 $Y=1.765 $X2=0 $Y2=0
cc_450 N_B2_c_556_n N_Y_c_886_n 0.0458338f $X=7.475 $Y=1.515 $X2=0 $Y2=0
cc_451 N_B2_c_557_n N_Y_c_886_n 2.20176e-19 $X=7.785 $Y=1.557 $X2=0 $Y2=0
cc_452 N_B2_c_558_n N_Y_c_887_n 0.00377434f $X=6.435 $Y=1.765 $X2=0 $Y2=0
cc_453 N_B2_c_559_n N_Y_c_939_n 0.0120074f $X=6.885 $Y=1.765 $X2=0 $Y2=0
cc_454 N_B2_c_560_n N_Y_c_939_n 0.0120074f $X=7.335 $Y=1.765 $X2=0 $Y2=0
cc_455 N_B2_c_556_n N_Y_c_939_n 0.0393875f $X=7.475 $Y=1.515 $X2=0 $Y2=0
cc_456 N_B2_c_557_n N_Y_c_939_n 0.00130859f $X=7.785 $Y=1.557 $X2=0 $Y2=0
cc_457 N_B2_c_558_n N_Y_c_943_n 0.014383f $X=6.435 $Y=1.765 $X2=0 $Y2=0
cc_458 N_B2_c_559_n N_Y_c_943_n 0.00991071f $X=6.885 $Y=1.765 $X2=0 $Y2=0
cc_459 N_B2_c_560_n N_Y_c_943_n 5.61652e-19 $X=7.335 $Y=1.765 $X2=0 $Y2=0
cc_460 N_B2_c_556_n N_Y_c_943_n 0.0237598f $X=7.475 $Y=1.515 $X2=0 $Y2=0
cc_461 N_B2_c_557_n N_Y_c_943_n 0.00144657f $X=7.785 $Y=1.557 $X2=0 $Y2=0
cc_462 N_B2_c_559_n N_Y_c_948_n 5.61652e-19 $X=6.885 $Y=1.765 $X2=0 $Y2=0
cc_463 N_B2_c_560_n N_Y_c_948_n 0.00991071f $X=7.335 $Y=1.765 $X2=0 $Y2=0
cc_464 N_B2_c_561_n N_Y_c_948_n 0.0105586f $X=7.785 $Y=1.765 $X2=0 $Y2=0
cc_465 N_B2_c_556_n N_Y_c_948_n 0.0189517f $X=7.475 $Y=1.515 $X2=0 $Y2=0
cc_466 N_B2_c_557_n N_Y_c_948_n 0.00269473f $X=7.785 $Y=1.557 $X2=0 $Y2=0
cc_467 N_B2_c_558_n N_A_1215_368#_c_989_n 0.0137046f $X=6.435 $Y=1.765 $X2=0
+ $Y2=0
cc_468 N_B2_c_559_n N_A_1215_368#_c_989_n 0.0128349f $X=6.885 $Y=1.765 $X2=0
+ $Y2=0
cc_469 N_B2_c_560_n N_A_1215_368#_c_991_n 0.0127839f $X=7.335 $Y=1.765 $X2=0
+ $Y2=0
cc_470 N_B2_c_561_n N_A_1215_368#_c_991_n 0.0125358f $X=7.785 $Y=1.765 $X2=0
+ $Y2=0
cc_471 N_B2_M1000_g N_VGND_c_1124_n 0.00383152f $X=6.365 $Y=0.74 $X2=0 $Y2=0
cc_472 N_B2_M1000_g N_VGND_c_1125_n 0.00964869f $X=6.365 $Y=0.74 $X2=0 $Y2=0
cc_473 N_B2_M1024_g N_VGND_c_1125_n 0.00418685f $X=6.865 $Y=0.74 $X2=0 $Y2=0
cc_474 N_B2_M1024_g N_VGND_c_1126_n 5.14838e-19 $X=6.865 $Y=0.74 $X2=0 $Y2=0
cc_475 N_B2_M1027_g N_VGND_c_1126_n 0.010415f $X=7.295 $Y=0.74 $X2=0 $Y2=0
cc_476 N_B2_M1037_g N_VGND_c_1126_n 0.00418685f $X=7.795 $Y=0.74 $X2=0 $Y2=0
cc_477 N_B2_M1037_g N_VGND_c_1127_n 5.14838e-19 $X=7.795 $Y=0.74 $X2=0 $Y2=0
cc_478 N_B2_M1024_g N_VGND_c_1131_n 0.00434272f $X=6.865 $Y=0.74 $X2=0 $Y2=0
cc_479 N_B2_M1027_g N_VGND_c_1131_n 0.00383152f $X=7.295 $Y=0.74 $X2=0 $Y2=0
cc_480 N_B2_M1037_g N_VGND_c_1132_n 0.00434272f $X=7.795 $Y=0.74 $X2=0 $Y2=0
cc_481 N_B2_M1000_g N_VGND_c_1135_n 0.00757637f $X=6.365 $Y=0.74 $X2=0 $Y2=0
cc_482 N_B2_M1024_g N_VGND_c_1135_n 0.00820718f $X=6.865 $Y=0.74 $X2=0 $Y2=0
cc_483 N_B2_M1027_g N_VGND_c_1135_n 0.0075754f $X=7.295 $Y=0.74 $X2=0 $Y2=0
cc_484 N_B2_M1037_g N_VGND_c_1135_n 0.00820816f $X=7.795 $Y=0.74 $X2=0 $Y2=0
cc_485 N_B2_M1000_g N_A_857_74#_c_1254_n 9.48753e-19 $X=6.365 $Y=0.74 $X2=0
+ $Y2=0
cc_486 N_B2_M1000_g N_A_857_74#_c_1255_n 0.0132997f $X=6.365 $Y=0.74 $X2=0 $Y2=0
cc_487 N_B2_M1024_g N_A_857_74#_c_1255_n 0.0115433f $X=6.865 $Y=0.74 $X2=0 $Y2=0
cc_488 N_B2_c_556_n N_A_857_74#_c_1255_n 0.051298f $X=7.475 $Y=1.515 $X2=0 $Y2=0
cc_489 N_B2_c_557_n N_A_857_74#_c_1255_n 0.00381149f $X=7.785 $Y=1.557 $X2=0
+ $Y2=0
cc_490 N_B2_c_556_n N_A_857_74#_c_1256_n 0.0153286f $X=7.475 $Y=1.515 $X2=0
+ $Y2=0
cc_491 N_B2_M1000_g N_A_857_74#_c_1257_n 9.78807e-19 $X=6.365 $Y=0.74 $X2=0
+ $Y2=0
cc_492 N_B2_M1024_g N_A_857_74#_c_1257_n 0.00922099f $X=6.865 $Y=0.74 $X2=0
+ $Y2=0
cc_493 N_B2_M1027_g N_A_857_74#_c_1257_n 3.97481e-19 $X=7.295 $Y=0.74 $X2=0
+ $Y2=0
cc_494 N_B2_M1027_g N_A_857_74#_c_1258_n 0.0134949f $X=7.295 $Y=0.74 $X2=0 $Y2=0
cc_495 N_B2_M1037_g N_A_857_74#_c_1258_n 0.0153304f $X=7.795 $Y=0.74 $X2=0 $Y2=0
cc_496 N_B2_c_556_n N_A_857_74#_c_1258_n 0.0358392f $X=7.475 $Y=1.515 $X2=0
+ $Y2=0
cc_497 N_B2_c_557_n N_A_857_74#_c_1258_n 0.00381149f $X=7.785 $Y=1.557 $X2=0
+ $Y2=0
cc_498 N_B2_M1027_g N_A_857_74#_c_1259_n 9.78807e-19 $X=7.295 $Y=0.74 $X2=0
+ $Y2=0
cc_499 N_B2_M1037_g N_A_857_74#_c_1259_n 0.00922099f $X=7.795 $Y=0.74 $X2=0
+ $Y2=0
cc_500 N_B2_M1024_g N_A_857_74#_c_1265_n 0.00157732f $X=6.865 $Y=0.74 $X2=0
+ $Y2=0
cc_501 N_B2_c_556_n N_A_857_74#_c_1265_n 0.0213626f $X=7.475 $Y=1.515 $X2=0
+ $Y2=0
cc_502 N_B2_c_557_n N_A_857_74#_c_1265_n 0.00232957f $X=7.785 $Y=1.557 $X2=0
+ $Y2=0
cc_503 N_B2_M1037_g N_A_857_74#_c_1266_n 0.0024689f $X=7.795 $Y=0.74 $X2=0 $Y2=0
cc_504 N_B2_c_557_n N_A_857_74#_c_1266_n 2.2764e-19 $X=7.785 $Y=1.557 $X2=0
+ $Y2=0
cc_505 N_B1_c_649_n N_VPWR_c_734_n 0.00972561f $X=8.235 $Y=1.765 $X2=0 $Y2=0
cc_506 N_B1_c_650_n N_VPWR_c_734_n 0.00303585f $X=8.685 $Y=1.765 $X2=0 $Y2=0
cc_507 N_B1_c_651_n N_VPWR_c_735_n 0.00289754f $X=9.135 $Y=1.765 $X2=0 $Y2=0
cc_508 N_B1_c_652_n N_VPWR_c_735_n 0.00291556f $X=9.585 $Y=1.765 $X2=0 $Y2=0
cc_509 N_B1_c_649_n N_VPWR_c_746_n 0.00413917f $X=8.235 $Y=1.765 $X2=0 $Y2=0
cc_510 N_B1_c_650_n N_VPWR_c_747_n 0.00445602f $X=8.685 $Y=1.765 $X2=0 $Y2=0
cc_511 N_B1_c_651_n N_VPWR_c_747_n 0.00445602f $X=9.135 $Y=1.765 $X2=0 $Y2=0
cc_512 N_B1_c_652_n N_VPWR_c_748_n 0.00445602f $X=9.585 $Y=1.765 $X2=0 $Y2=0
cc_513 N_B1_c_649_n N_VPWR_c_724_n 0.0081781f $X=8.235 $Y=1.765 $X2=0 $Y2=0
cc_514 N_B1_c_650_n N_VPWR_c_724_n 0.00857253f $X=8.685 $Y=1.765 $X2=0 $Y2=0
cc_515 N_B1_c_651_n N_VPWR_c_724_n 0.00857253f $X=9.135 $Y=1.765 $X2=0 $Y2=0
cc_516 N_B1_c_652_n N_VPWR_c_724_n 0.00860602f $X=9.585 $Y=1.765 $X2=0 $Y2=0
cc_517 N_B1_c_649_n N_A_1215_368#_c_991_n 0.0010012f $X=8.235 $Y=1.765 $X2=0
+ $Y2=0
cc_518 N_B1_c_649_n N_A_1215_368#_c_1003_n 0.0126853f $X=8.235 $Y=1.765 $X2=0
+ $Y2=0
cc_519 N_B1_c_650_n N_A_1215_368#_c_1003_n 0.0119563f $X=8.685 $Y=1.765 $X2=0
+ $Y2=0
cc_520 B1 N_A_1215_368#_c_1003_n 0.0409153f $X=9.755 $Y=1.58 $X2=0 $Y2=0
cc_521 N_B1_c_648_n N_A_1215_368#_c_1003_n 0.00130859f $X=9.585 $Y=1.557 $X2=0
+ $Y2=0
cc_522 N_B1_c_649_n N_A_1215_368#_c_992_n 6.51912e-19 $X=8.235 $Y=1.765 $X2=0
+ $Y2=0
cc_523 N_B1_c_650_n N_A_1215_368#_c_992_n 0.0103961f $X=8.685 $Y=1.765 $X2=0
+ $Y2=0
cc_524 N_B1_c_651_n N_A_1215_368#_c_992_n 0.0102302f $X=9.135 $Y=1.765 $X2=0
+ $Y2=0
cc_525 N_B1_c_652_n N_A_1215_368#_c_992_n 6.30912e-19 $X=9.585 $Y=1.765 $X2=0
+ $Y2=0
cc_526 N_B1_c_651_n N_A_1215_368#_c_1011_n 0.0120074f $X=9.135 $Y=1.765 $X2=0
+ $Y2=0
cc_527 N_B1_c_652_n N_A_1215_368#_c_1011_n 0.0120074f $X=9.585 $Y=1.765 $X2=0
+ $Y2=0
cc_528 B1 N_A_1215_368#_c_1011_n 0.0393875f $X=9.755 $Y=1.58 $X2=0 $Y2=0
cc_529 N_B1_c_648_n N_A_1215_368#_c_1011_n 0.00131353f $X=9.585 $Y=1.557 $X2=0
+ $Y2=0
cc_530 N_B1_c_652_n N_A_1215_368#_c_993_n 4.27055e-19 $X=9.585 $Y=1.765 $X2=0
+ $Y2=0
cc_531 B1 N_A_1215_368#_c_993_n 0.0247152f $X=9.755 $Y=1.58 $X2=0 $Y2=0
cc_532 N_B1_c_648_n N_A_1215_368#_c_993_n 9.11744e-19 $X=9.585 $Y=1.557 $X2=0
+ $Y2=0
cc_533 N_B1_c_651_n N_A_1215_368#_c_994_n 6.25988e-19 $X=9.135 $Y=1.765 $X2=0
+ $Y2=0
cc_534 N_B1_c_652_n N_A_1215_368#_c_994_n 0.0103728f $X=9.585 $Y=1.765 $X2=0
+ $Y2=0
cc_535 N_B1_c_650_n N_A_1215_368#_c_1020_n 4.27055e-19 $X=8.685 $Y=1.765 $X2=0
+ $Y2=0
cc_536 N_B1_c_651_n N_A_1215_368#_c_1020_n 4.27055e-19 $X=9.135 $Y=1.765 $X2=0
+ $Y2=0
cc_537 B1 N_A_1215_368#_c_1020_n 0.0237598f $X=9.755 $Y=1.58 $X2=0 $Y2=0
cc_538 N_B1_c_648_n N_A_1215_368#_c_1020_n 0.00144162f $X=9.585 $Y=1.557 $X2=0
+ $Y2=0
cc_539 N_B1_M1005_g N_VGND_c_1127_n 0.0104021f $X=8.225 $Y=0.74 $X2=0 $Y2=0
cc_540 N_B1_M1010_g N_VGND_c_1127_n 0.0104021f $X=8.655 $Y=0.74 $X2=0 $Y2=0
cc_541 N_B1_M1012_g N_VGND_c_1127_n 5.14838e-19 $X=9.085 $Y=0.74 $X2=0 $Y2=0
cc_542 N_B1_M1012_g N_VGND_c_1128_n 0.00418685f $X=9.085 $Y=0.74 $X2=0 $Y2=0
cc_543 N_B1_M1035_g N_VGND_c_1128_n 0.0133319f $X=9.585 $Y=0.74 $X2=0 $Y2=0
cc_544 N_B1_M1005_g N_VGND_c_1132_n 0.00383152f $X=8.225 $Y=0.74 $X2=0 $Y2=0
cc_545 N_B1_M1010_g N_VGND_c_1133_n 0.00383152f $X=8.655 $Y=0.74 $X2=0 $Y2=0
cc_546 N_B1_M1012_g N_VGND_c_1133_n 0.00434272f $X=9.085 $Y=0.74 $X2=0 $Y2=0
cc_547 N_B1_M1035_g N_VGND_c_1134_n 0.00383152f $X=9.585 $Y=0.74 $X2=0 $Y2=0
cc_548 N_B1_M1005_g N_VGND_c_1135_n 0.00757637f $X=8.225 $Y=0.74 $X2=0 $Y2=0
cc_549 N_B1_M1010_g N_VGND_c_1135_n 0.0075754f $X=8.655 $Y=0.74 $X2=0 $Y2=0
cc_550 N_B1_M1012_g N_VGND_c_1135_n 0.00820718f $X=9.085 $Y=0.74 $X2=0 $Y2=0
cc_551 N_B1_M1035_g N_VGND_c_1135_n 0.00761198f $X=9.585 $Y=0.74 $X2=0 $Y2=0
cc_552 N_B1_M1005_g N_A_857_74#_c_1259_n 3.97481e-19 $X=8.225 $Y=0.74 $X2=0
+ $Y2=0
cc_553 N_B1_M1005_g N_A_857_74#_c_1260_n 0.0130828f $X=8.225 $Y=0.74 $X2=0 $Y2=0
cc_554 N_B1_M1010_g N_A_857_74#_c_1260_n 0.0131017f $X=8.655 $Y=0.74 $X2=0 $Y2=0
cc_555 B1 N_A_857_74#_c_1260_n 0.0475521f $X=9.755 $Y=1.58 $X2=0 $Y2=0
cc_556 N_B1_c_648_n N_A_857_74#_c_1260_n 0.00239094f $X=9.585 $Y=1.557 $X2=0
+ $Y2=0
cc_557 N_B1_M1010_g N_A_857_74#_c_1261_n 3.97481e-19 $X=8.655 $Y=0.74 $X2=0
+ $Y2=0
cc_558 N_B1_M1012_g N_A_857_74#_c_1261_n 0.00922099f $X=9.085 $Y=0.74 $X2=0
+ $Y2=0
cc_559 N_B1_M1035_g N_A_857_74#_c_1261_n 9.78807e-19 $X=9.585 $Y=0.74 $X2=0
+ $Y2=0
cc_560 N_B1_M1012_g N_A_857_74#_c_1262_n 0.0115433f $X=9.085 $Y=0.74 $X2=0 $Y2=0
cc_561 N_B1_M1035_g N_A_857_74#_c_1262_n 0.0140566f $X=9.585 $Y=0.74 $X2=0 $Y2=0
cc_562 B1 N_A_857_74#_c_1262_n 0.0721685f $X=9.755 $Y=1.58 $X2=0 $Y2=0
cc_563 N_B1_c_648_n N_A_857_74#_c_1262_n 0.00797067f $X=9.585 $Y=1.557 $X2=0
+ $Y2=0
cc_564 N_B1_M1035_g N_A_857_74#_c_1263_n 0.00159319f $X=9.585 $Y=0.74 $X2=0
+ $Y2=0
cc_565 N_B1_M1012_g N_A_857_74#_c_1267_n 0.00157732f $X=9.085 $Y=0.74 $X2=0
+ $Y2=0
cc_566 B1 N_A_857_74#_c_1267_n 0.0213626f $X=9.755 $Y=1.58 $X2=0 $Y2=0
cc_567 N_B1_c_648_n N_A_857_74#_c_1267_n 0.00232957f $X=9.585 $Y=1.557 $X2=0
+ $Y2=0
cc_568 N_VPWR_c_730_n N_Y_c_881_n 0.0657826f $X=3.87 $Y=1.985 $X2=0 $Y2=0
cc_569 N_VPWR_c_731_n N_Y_c_881_n 0.0547423f $X=4.77 $Y=2.305 $X2=0 $Y2=0
cc_570 N_VPWR_c_744_n N_Y_c_881_n 0.014552f $X=4.685 $Y=3.33 $X2=0 $Y2=0
cc_571 N_VPWR_c_724_n N_Y_c_881_n 0.0119791f $X=9.84 $Y=3.33 $X2=0 $Y2=0
cc_572 N_VPWR_M1019_d N_Y_c_882_n 0.00247267f $X=4.62 $Y=1.84 $X2=0 $Y2=0
cc_573 N_VPWR_c_731_n N_Y_c_882_n 0.0136682f $X=4.77 $Y=2.305 $X2=0 $Y2=0
cc_574 N_VPWR_c_730_n N_Y_c_883_n 0.0104177f $X=3.87 $Y=1.985 $X2=0 $Y2=0
cc_575 N_VPWR_c_731_n N_Y_c_884_n 0.0529204f $X=4.77 $Y=2.305 $X2=0 $Y2=0
cc_576 N_VPWR_c_732_n N_Y_c_884_n 0.0110241f $X=5.505 $Y=3.33 $X2=0 $Y2=0
cc_577 N_VPWR_c_733_n N_Y_c_884_n 0.0442833f $X=5.67 $Y=2.405 $X2=0 $Y2=0
cc_578 N_VPWR_c_724_n N_Y_c_884_n 0.00909194f $X=9.84 $Y=3.33 $X2=0 $Y2=0
cc_579 N_VPWR_M1028_d N_Y_c_886_n 0.00321299f $X=5.52 $Y=1.84 $X2=0 $Y2=0
cc_580 N_VPWR_c_733_n N_Y_c_886_n 0.00863845f $X=5.67 $Y=2.405 $X2=0 $Y2=0
cc_581 N_VPWR_M1028_d N_Y_c_887_n 0.0054101f $X=5.52 $Y=1.84 $X2=0 $Y2=0
cc_582 N_VPWR_c_731_n N_Y_c_887_n 6.83856e-19 $X=4.77 $Y=2.305 $X2=0 $Y2=0
cc_583 N_VPWR_c_733_n N_Y_c_887_n 0.0127008f $X=5.67 $Y=2.405 $X2=0 $Y2=0
cc_584 N_VPWR_c_733_n N_A_1215_368#_c_988_n 0.0412871f $X=5.67 $Y=2.405 $X2=0
+ $Y2=0
cc_585 N_VPWR_c_746_n N_A_1215_368#_c_989_n 0.0441612f $X=8.295 $Y=3.33 $X2=0
+ $Y2=0
cc_586 N_VPWR_c_724_n N_A_1215_368#_c_989_n 0.0249452f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_587 N_VPWR_c_733_n N_A_1215_368#_c_990_n 0.0129575f $X=5.67 $Y=2.405 $X2=0
+ $Y2=0
cc_588 N_VPWR_c_746_n N_A_1215_368#_c_990_n 0.018997f $X=8.295 $Y=3.33 $X2=0
+ $Y2=0
cc_589 N_VPWR_c_724_n N_A_1215_368#_c_990_n 0.0103026f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_590 N_VPWR_c_734_n N_A_1215_368#_c_991_n 0.0107938f $X=8.46 $Y=2.455 $X2=0
+ $Y2=0
cc_591 N_VPWR_c_746_n N_A_1215_368#_c_991_n 0.0584986f $X=8.295 $Y=3.33 $X2=0
+ $Y2=0
cc_592 N_VPWR_c_724_n N_A_1215_368#_c_991_n 0.0327208f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_593 N_VPWR_M1029_d N_A_1215_368#_c_1003_n 0.00359365f $X=8.31 $Y=1.84 $X2=0
+ $Y2=0
cc_594 N_VPWR_c_734_n N_A_1215_368#_c_1003_n 0.016157f $X=8.46 $Y=2.455 $X2=0
+ $Y2=0
cc_595 N_VPWR_c_734_n N_A_1215_368#_c_992_n 0.0249143f $X=8.46 $Y=2.455 $X2=0
+ $Y2=0
cc_596 N_VPWR_c_735_n N_A_1215_368#_c_992_n 0.0248868f $X=9.36 $Y=2.455 $X2=0
+ $Y2=0
cc_597 N_VPWR_c_747_n N_A_1215_368#_c_992_n 0.014552f $X=9.26 $Y=3.33 $X2=0
+ $Y2=0
cc_598 N_VPWR_c_724_n N_A_1215_368#_c_992_n 0.0119791f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_599 N_VPWR_M1036_d N_A_1215_368#_c_1011_n 0.00359365f $X=9.21 $Y=1.84 $X2=0
+ $Y2=0
cc_600 N_VPWR_c_735_n N_A_1215_368#_c_1011_n 0.0151327f $X=9.36 $Y=2.455 $X2=0
+ $Y2=0
cc_601 N_VPWR_c_735_n N_A_1215_368#_c_994_n 0.0254369f $X=9.36 $Y=2.455 $X2=0
+ $Y2=0
cc_602 N_VPWR_c_748_n N_A_1215_368#_c_994_n 0.0145938f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_603 N_VPWR_c_724_n N_A_1215_368#_c_994_n 0.0120466f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_604 N_VPWR_c_746_n N_A_1215_368#_c_995_n 0.0143373f $X=8.295 $Y=3.33 $X2=0
+ $Y2=0
cc_605 N_VPWR_c_724_n N_A_1215_368#_c_995_n 0.00777554f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_606 N_Y_c_886_n N_A_1215_368#_M1018_s 0.0058041f $X=6.495 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_607 N_Y_c_939_n N_A_1215_368#_M1020_s 0.00359365f $X=7.395 $Y=2.035 $X2=0
+ $Y2=0
cc_608 N_Y_c_886_n N_A_1215_368#_c_988_n 0.0209991f $X=6.495 $Y=2.035 $X2=0
+ $Y2=0
cc_609 N_Y_M1018_d N_A_1215_368#_c_989_n 0.00197722f $X=6.51 $Y=1.84 $X2=0 $Y2=0
cc_610 N_Y_c_943_n N_A_1215_368#_c_989_n 0.0160777f $X=6.66 $Y=2.055 $X2=0 $Y2=0
cc_611 N_Y_c_939_n N_A_1215_368#_c_1051_n 0.0151327f $X=7.395 $Y=2.035 $X2=0
+ $Y2=0
cc_612 N_Y_M1023_d N_A_1215_368#_c_991_n 0.00197722f $X=7.41 $Y=1.84 $X2=0 $Y2=0
cc_613 N_Y_c_948_n N_A_1215_368#_c_991_n 0.0160777f $X=7.56 $Y=2.055 $X2=0 $Y2=0
cc_614 N_Y_c_877_n N_A_857_74#_M1016_d 0.00176461f $X=5.545 $Y=1.045 $X2=0 $Y2=0
cc_615 N_Y_c_878_n N_A_857_74#_c_1251_n 0.00756924f $X=5.025 $Y=1.045 $X2=0
+ $Y2=0
cc_616 N_Y_M1007_s N_A_857_74#_c_1252_n 0.00176461f $X=4.72 $Y=0.37 $X2=0 $Y2=0
cc_617 N_Y_c_900_n N_A_857_74#_c_1252_n 0.0157609f $X=4.86 $Y=0.86 $X2=0 $Y2=0
cc_618 N_Y_c_877_n N_A_857_74#_c_1252_n 0.0032855f $X=5.545 $Y=1.045 $X2=0 $Y2=0
cc_619 N_Y_c_877_n N_A_857_74#_c_1318_n 0.0132452f $X=5.545 $Y=1.045 $X2=0 $Y2=0
cc_620 N_Y_M1022_s N_A_857_74#_c_1254_n 0.00176461f $X=5.58 $Y=0.37 $X2=0 $Y2=0
cc_621 N_Y_c_877_n N_A_857_74#_c_1254_n 0.00302054f $X=5.545 $Y=1.045 $X2=0
+ $Y2=0
cc_622 N_Y_c_913_n N_A_857_74#_c_1254_n 0.0166135f $X=5.72 $Y=0.86 $X2=0 $Y2=0
cc_623 N_Y_c_879_n N_A_857_74#_c_1256_n 0.00252526f $X=5.63 $Y=1.8 $X2=0 $Y2=0
cc_624 N_Y_c_880_n N_A_857_74#_c_1256_n 0.00570271f $X=5.715 $Y=1.045 $X2=0
+ $Y2=0
cc_625 N_A_27_74#_c_1055_n N_VGND_M1009_s 0.00176461f $X=1.055 $Y=1.095
+ $X2=-0.19 $Y2=-0.245
cc_626 N_A_27_74#_c_1058_n N_VGND_M1033_s 0.00176461f $X=1.925 $Y=1.095 $X2=0
+ $Y2=0
cc_627 N_A_27_74#_c_1054_n N_VGND_c_1122_n 0.0182902f $X=0.28 $Y=0.515 $X2=0
+ $Y2=0
cc_628 N_A_27_74#_c_1055_n N_VGND_c_1122_n 0.0171619f $X=1.055 $Y=1.095 $X2=0
+ $Y2=0
cc_629 N_A_27_74#_c_1057_n N_VGND_c_1122_n 0.0182548f $X=1.145 $Y=0.515 $X2=0
+ $Y2=0
cc_630 N_A_27_74#_c_1057_n N_VGND_c_1123_n 0.0182548f $X=1.145 $Y=0.515 $X2=0
+ $Y2=0
cc_631 N_A_27_74#_c_1058_n N_VGND_c_1123_n 0.0171619f $X=1.925 $Y=1.095 $X2=0
+ $Y2=0
cc_632 N_A_27_74#_c_1060_n N_VGND_c_1123_n 0.0112234f $X=2.095 $Y=0.34 $X2=0
+ $Y2=0
cc_633 N_A_27_74#_c_1059_n N_VGND_c_1124_n 0.0428729f $X=2.775 $Y=0.34 $X2=0
+ $Y2=0
cc_634 N_A_27_74#_c_1060_n N_VGND_c_1124_n 0.0121867f $X=2.095 $Y=0.34 $X2=0
+ $Y2=0
cc_635 N_A_27_74#_c_1061_n N_VGND_c_1124_n 0.0607975f $X=3.785 $Y=0.34 $X2=0
+ $Y2=0
cc_636 N_A_27_74#_c_1064_n N_VGND_c_1124_n 0.023391f $X=2.94 $Y=0.34 $X2=0 $Y2=0
cc_637 N_A_27_74#_c_1054_n N_VGND_c_1129_n 0.011066f $X=0.28 $Y=0.515 $X2=0
+ $Y2=0
cc_638 N_A_27_74#_c_1057_n N_VGND_c_1130_n 0.00794252f $X=1.145 $Y=0.515 $X2=0
+ $Y2=0
cc_639 N_A_27_74#_c_1054_n N_VGND_c_1135_n 0.00915947f $X=0.28 $Y=0.515 $X2=0
+ $Y2=0
cc_640 N_A_27_74#_c_1057_n N_VGND_c_1135_n 0.00657413f $X=1.145 $Y=0.515 $X2=0
+ $Y2=0
cc_641 N_A_27_74#_c_1059_n N_VGND_c_1135_n 0.0241933f $X=2.775 $Y=0.34 $X2=0
+ $Y2=0
cc_642 N_A_27_74#_c_1060_n N_VGND_c_1135_n 0.00660921f $X=2.095 $Y=0.34 $X2=0
+ $Y2=0
cc_643 N_A_27_74#_c_1061_n N_VGND_c_1135_n 0.0339133f $X=3.785 $Y=0.34 $X2=0
+ $Y2=0
cc_644 N_A_27_74#_c_1064_n N_VGND_c_1135_n 0.0127797f $X=2.94 $Y=0.34 $X2=0
+ $Y2=0
cc_645 N_A_27_74#_c_1062_n N_A_857_74#_c_1251_n 0.0455088f $X=3.87 $Y=0.515
+ $X2=0 $Y2=0
cc_646 N_A_27_74#_c_1061_n N_A_857_74#_c_1253_n 0.0128665f $X=3.785 $Y=0.34
+ $X2=0 $Y2=0
cc_647 N_VGND_c_1124_n N_A_857_74#_c_1252_n 0.043517f $X=6.415 $Y=0 $X2=0 $Y2=0
cc_648 N_VGND_c_1135_n N_A_857_74#_c_1252_n 0.0245693f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_649 N_VGND_c_1124_n N_A_857_74#_c_1253_n 0.0179217f $X=6.415 $Y=0 $X2=0 $Y2=0
cc_650 N_VGND_c_1135_n N_A_857_74#_c_1253_n 0.00971942f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_651 N_VGND_c_1124_n N_A_857_74#_c_1254_n 0.0557038f $X=6.415 $Y=0 $X2=0 $Y2=0
cc_652 N_VGND_c_1125_n N_A_857_74#_c_1254_n 0.0112234f $X=6.58 $Y=0.65 $X2=0
+ $Y2=0
cc_653 N_VGND_c_1135_n N_A_857_74#_c_1254_n 0.0311785f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_654 N_VGND_M1000_d N_A_857_74#_c_1255_n 0.00256964f $X=6.44 $Y=0.37 $X2=0
+ $Y2=0
cc_655 N_VGND_c_1125_n N_A_857_74#_c_1255_n 0.0201026f $X=6.58 $Y=0.65 $X2=0
+ $Y2=0
cc_656 N_VGND_c_1125_n N_A_857_74#_c_1257_n 0.018051f $X=6.58 $Y=0.65 $X2=0
+ $Y2=0
cc_657 N_VGND_c_1126_n N_A_857_74#_c_1257_n 0.0179318f $X=7.51 $Y=0.65 $X2=0
+ $Y2=0
cc_658 N_VGND_c_1131_n N_A_857_74#_c_1257_n 0.0109942f $X=7.345 $Y=0 $X2=0 $Y2=0
cc_659 N_VGND_c_1135_n N_A_857_74#_c_1257_n 0.00904371f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_660 N_VGND_M1027_d N_A_857_74#_c_1258_n 0.00256964f $X=7.37 $Y=0.37 $X2=0
+ $Y2=0
cc_661 N_VGND_c_1126_n N_A_857_74#_c_1258_n 0.0201026f $X=7.51 $Y=0.65 $X2=0
+ $Y2=0
cc_662 N_VGND_c_1126_n N_A_857_74#_c_1259_n 0.018051f $X=7.51 $Y=0.65 $X2=0
+ $Y2=0
cc_663 N_VGND_c_1127_n N_A_857_74#_c_1259_n 0.0179318f $X=8.44 $Y=0.65 $X2=0
+ $Y2=0
cc_664 N_VGND_c_1132_n N_A_857_74#_c_1259_n 0.0109942f $X=8.275 $Y=0 $X2=0 $Y2=0
cc_665 N_VGND_c_1135_n N_A_857_74#_c_1259_n 0.00904371f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_666 N_VGND_M1005_s N_A_857_74#_c_1260_n 0.00180746f $X=8.3 $Y=0.37 $X2=0
+ $Y2=0
cc_667 N_VGND_c_1127_n N_A_857_74#_c_1260_n 0.0163515f $X=8.44 $Y=0.65 $X2=0
+ $Y2=0
cc_668 N_VGND_c_1127_n N_A_857_74#_c_1261_n 0.0179318f $X=8.44 $Y=0.65 $X2=0
+ $Y2=0
cc_669 N_VGND_c_1128_n N_A_857_74#_c_1261_n 0.018051f $X=9.37 $Y=0.65 $X2=0
+ $Y2=0
cc_670 N_VGND_c_1133_n N_A_857_74#_c_1261_n 0.0109942f $X=9.205 $Y=0 $X2=0 $Y2=0
cc_671 N_VGND_c_1135_n N_A_857_74#_c_1261_n 0.00904371f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_672 N_VGND_M1012_s N_A_857_74#_c_1262_n 0.00256964f $X=9.16 $Y=0.37 $X2=0
+ $Y2=0
cc_673 N_VGND_c_1128_n N_A_857_74#_c_1262_n 0.0201026f $X=9.37 $Y=0.65 $X2=0
+ $Y2=0
cc_674 N_VGND_c_1128_n N_A_857_74#_c_1263_n 0.0179318f $X=9.37 $Y=0.65 $X2=0
+ $Y2=0
cc_675 N_VGND_c_1134_n N_A_857_74#_c_1263_n 0.011066f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_676 N_VGND_c_1135_n N_A_857_74#_c_1263_n 0.00915947f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_677 N_VGND_c_1124_n N_A_857_74#_c_1264_n 0.0119713f $X=6.415 $Y=0 $X2=0 $Y2=0
cc_678 N_VGND_c_1135_n N_A_857_74#_c_1264_n 0.00656877f $X=9.84 $Y=0 $X2=0 $Y2=0
