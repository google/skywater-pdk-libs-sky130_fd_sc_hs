* File: sky130_fd_sc_hs__a41o_4.spice
* Created: Tue Sep  1 19:54:11 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hs__a41o_4.pex.spice"
.subckt sky130_fd_sc_hs__a41o_4  VNB VPB B1 A1 A2 A3 A4 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A4	A4
* A3	A3
* A2	A2
* A1	A1
* B1	B1
* VPB	VPB
* VNB	VNB
MM1012 N_A_113_98#_M1012_d N_B1_M1012_g N_VGND_M1012_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.2072 PD=1.02 PS=2.04 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75002.7 A=0.111 P=1.78 MULT=1
MM1017 N_A_113_98#_M1012_d N_B1_M1017_g N_VGND_M1017_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1955 PD=1.02 PS=1.43 NRD=0 NRS=33.912 M=1 R=4.93333 SA=75000.6
+ SB=75002.3 A=0.111 P=1.78 MULT=1
MM1002 N_VGND_M1017_s N_A_113_98#_M1002_g N_X_M1002_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1955 AS=0.1036 PD=1.43 PS=1.02 NRD=33.912 NRS=0 M=1 R=4.93333 SA=75001.2
+ SB=75001.7 A=0.111 P=1.78 MULT=1
MM1009 N_VGND_M1009_d N_A_113_98#_M1009_g N_X_M1002_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.193 AS=0.1036 PD=1.425 PS=1.02 NRD=33.372 NRS=0 M=1 R=4.93333 SA=75001.6
+ SB=75001.3 A=0.111 P=1.78 MULT=1
MM1016 N_VGND_M1009_d N_A_113_98#_M1016_g N_X_M1016_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.193 AS=0.1036 PD=1.425 PS=1.02 NRD=33.372 NRS=0 M=1 R=4.93333 SA=75002.2
+ SB=75000.7 A=0.111 P=1.78 MULT=1
MM1023 N_VGND_M1023_d N_A_113_98#_M1023_g N_X_M1016_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.3495 AS=0.1036 PD=2.81 PS=1.02 NRD=67.668 NRS=0 M=1 R=4.93333 SA=75002.6
+ SB=75000.3 A=0.111 P=1.78 MULT=1
MM1013 N_A_113_98#_M1013_d N_A1_M1013_g N_A_751_74#_M1013_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.2109 PD=1.02 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75001.5 A=0.111 P=1.78 MULT=1
MM1014 N_A_113_98#_M1013_d N_A1_M1014_g N_A_751_74#_M1014_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.6 SB=75001.1 A=0.111 P=1.78 MULT=1
MM1011 N_A_751_74#_M1014_s N_A2_M1011_g N_A_1010_74#_M1011_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75001.1 SB=75000.6 A=0.111 P=1.78 MULT=1
MM1026 N_A_751_74#_M1026_d N_A2_M1026_g N_A_1010_74#_M1011_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.2035 AS=0.1036 PD=2.03 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75001.5 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1007 N_A_1205_74#_M1007_d N_A3_M1007_g N_A_1010_74#_M1007_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.2072 AS=0.1036 PD=2.04 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75001.5 A=0.111 P=1.78 MULT=1
MM1018 N_A_1205_74#_M1018_d N_A3_M1018_g N_A_1010_74#_M1007_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.6 SB=75001.1 A=0.111 P=1.78 MULT=1
MM1004 N_A_1205_74#_M1018_d N_A4_M1004_g N_VGND_M1004_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.1
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1015 N_A_1205_74#_M1015_d N_A4_M1015_g N_VGND_M1004_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.2072 AS=0.1036 PD=2.04 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.5
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1006 N_A_27_392#_M1006_d N_B1_M1006_g N_A_113_98#_M1006_s VPB PSHORT L=0.15
+ W=1 AD=0.295 AS=0.175 PD=2.59 PS=1.35 NRD=1.9503 NRS=11.8003 M=1 R=6.66667
+ SA=75000.2 SB=75000.7 A=0.15 P=2.3 MULT=1
MM1010 N_A_27_392#_M1010_d N_B1_M1010_g N_A_113_98#_M1006_s VPB PSHORT L=0.15
+ W=1 AD=0.295 AS=0.175 PD=2.59 PS=1.35 NRD=1.9503 NRS=1.9503 M=1 R=6.66667
+ SA=75000.7 SB=75000.2 A=0.15 P=2.3 MULT=1
MM1000 N_VPWR_M1000_d N_A_113_98#_M1000_g N_X_M1000_s VPB PSHORT L=0.15 W=1.12
+ AD=0.3304 AS=0.168 PD=2.83 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75005.4 A=0.168 P=2.54 MULT=1
MM1001 N_VPWR_M1001_d N_A_113_98#_M1001_g N_X_M1000_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.7 SB=75004.9 A=0.168 P=2.54 MULT=1
MM1003 N_VPWR_M1001_d N_A_113_98#_M1003_g N_X_M1003_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.1 SB=75004.5 A=0.168 P=2.54 MULT=1
MM1027 N_VPWR_M1027_d N_A_113_98#_M1027_g N_X_M1003_s VPB PSHORT L=0.15 W=1.12
+ AD=0.212272 AS=0.168 PD=1.57434 PS=1.42 NRD=3.5066 NRS=1.7533 M=1 R=7.46667
+ SA=75001.6 SB=75004 A=0.168 P=2.54 MULT=1
MM1005 N_VPWR_M1027_d N_A1_M1005_g N_A_27_392#_M1005_s VPB PSHORT L=0.15 W=1
+ AD=0.189528 AS=0.2475 PD=1.40566 PS=1.495 NRD=13.7703 NRS=21.67 M=1 R=6.66667
+ SA=75002.1 SB=75004 A=0.15 P=2.3 MULT=1
MM1008 N_VPWR_M1008_d N_A1_M1008_g N_A_27_392#_M1005_s VPB PSHORT L=0.15 W=1
+ AD=0.2625 AS=0.2475 PD=1.525 PS=1.495 NRD=23.6203 NRS=20.685 M=1 R=6.66667
+ SA=75002.7 SB=75003.3 A=0.15 P=2.3 MULT=1
MM1024 N_A_27_392#_M1024_d N_A2_M1024_g N_VPWR_M1008_d VPB PSHORT L=0.15 W=1
+ AD=0.15 AS=0.2625 PD=1.3 PS=1.525 NRD=1.9503 NRS=24.6053 M=1 R=6.66667
+ SA=75003.4 SB=75002.7 A=0.15 P=2.3 MULT=1
MM1025 N_A_27_392#_M1024_d N_A2_M1025_g N_VPWR_M1025_s VPB PSHORT L=0.15 W=1
+ AD=0.15 AS=0.2 PD=1.3 PS=1.4 NRD=1.9503 NRS=11.8003 M=1 R=6.66667 SA=75003.9
+ SB=75002.2 A=0.15 P=2.3 MULT=1
MM1019 N_VPWR_M1025_s N_A3_M1019_g N_A_27_392#_M1019_s VPB PSHORT L=0.15 W=1
+ AD=0.2 AS=0.175 PD=1.4 PS=1.35 NRD=11.8003 NRS=1.9503 M=1 R=6.66667 SA=75004.4
+ SB=75001.7 A=0.15 P=2.3 MULT=1
MM1021 N_VPWR_M1021_d N_A3_M1021_g N_A_27_392#_M1019_s VPB PSHORT L=0.15 W=1
+ AD=0.175 AS=0.175 PD=1.35 PS=1.35 NRD=1.9503 NRS=11.8003 M=1 R=6.66667
+ SA=75004.9 SB=75001.2 A=0.15 P=2.3 MULT=1
MM1020 N_A_27_392#_M1020_d N_A4_M1020_g N_VPWR_M1021_d VPB PSHORT L=0.15 W=1
+ AD=0.15 AS=0.175 PD=1.3 PS=1.35 NRD=1.9503 NRS=11.8003 M=1 R=6.66667
+ SA=75005.4 SB=75000.7 A=0.15 P=2.3 MULT=1
MM1022 N_A_27_392#_M1020_d N_A4_M1022_g N_VPWR_M1022_s VPB PSHORT L=0.15 W=1
+ AD=0.15 AS=0.295 PD=1.3 PS=2.59 NRD=1.9503 NRS=1.9503 M=1 R=6.66667 SA=75005.9
+ SB=75000.2 A=0.15 P=2.3 MULT=1
DX28_noxref VNB VPB NWDIODE A=15.8844 P=20.8
c_134 VPB 0 1.25754e-19 $X=0 $Y=3.085
*
.include "sky130_fd_sc_hs__a41o_4.pxi.spice"
*
.ends
*
*
