* File: sky130_fd_sc_hs__dfxbp_2.spice
* Created: Thu Aug 27 20:39:49 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hs__dfxbp_2.pex.spice"
.subckt sky130_fd_sc_hs__dfxbp_2  VNB VPB CLK D VPWR Q Q_N VGND
* 
* VGND	VGND
* Q_N	Q_N
* Q	Q
* VPWR	VPWR
* D	D
* CLK	CLK
* VPB	VPB
* VNB	VNB
MM1025 N_VGND_M1025_d N_CLK_M1025_g N_A_27_74#_M1025_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.20385 AS=0.2109 PD=1.355 PS=2.05 NRD=17.832 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75000.9 A=0.111 P=1.78 MULT=1
MM1011 N_A_206_368#_M1011_d N_A_27_74#_M1011_g N_VGND_M1025_d VNB NLOWVT L=0.15
+ W=0.74 AD=0.3252 AS=0.20385 PD=2.59 PS=1.355 NRD=62.34 NRS=4.86 M=1 R=4.93333
+ SA=75000.9 SB=75000.3 A=0.111 P=1.78 MULT=1
MM1024 N_A_451_503#_M1024_d N_D_M1024_g N_VGND_M1024_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.0588 AS=0.35635 PD=0.7 PS=2.6 NRD=0 NRS=226.692 M=1 R=2.8 SA=75000.5
+ SB=75003.3 A=0.063 P=1.14 MULT=1
MM1026 N_A_558_445#_M1026_d N_A_27_74#_M1026_g N_A_451_503#_M1024_d VNB NLOWVT
+ L=0.15 W=0.42 AD=0.0830375 AS=0.0588 PD=0.865 PS=0.7 NRD=0 NRS=0 M=1 R=2.8
+ SA=75001 SB=75002.9 A=0.063 P=1.14 MULT=1
MM1014 A_717_102# N_A_206_368#_M1014_g N_A_558_445#_M1026_d VNB NLOWVT L=0.15
+ W=0.42 AD=0.0504 AS=0.0830375 PD=0.66 PS=0.865 NRD=18.564 NRS=22.848 M=1 R=2.8
+ SA=75001.2 SB=75002.8 A=0.063 P=1.14 MULT=1
MM1004 N_VGND_M1004_d N_A_753_284#_M1004_g A_717_102# VNB NLOWVT L=0.15 W=0.42
+ AD=0.0850825 AS=0.0504 PD=0.801031 PS=0.66 NRD=25.704 NRS=18.564 M=1 R=2.8
+ SA=75001.6 SB=75002.4 A=0.063 P=1.14 MULT=1
MM1007 N_A_753_284#_M1007_d N_A_558_445#_M1007_g N_VGND_M1004_d VNB NLOWVT
+ L=0.15 W=0.55 AD=0.1935 AS=0.111418 PD=1.49 PS=1.04897 NRD=64.752 NRS=2.172
+ M=1 R=3.66667 SA=75001.7 SB=75001.6 A=0.0825 P=1.4 MULT=1
MM1012 N_A_1000_424#_M1012_d N_A_206_368#_M1012_g N_A_753_284#_M1007_d VNB
+ NLOWVT L=0.15 W=0.55 AD=0.222296 AS=0.1935 PD=1.90515 PS=1.49 NRD=157.08
+ NRS=64.752 M=1 R=3.66667 SA=75002.3 SB=75001 A=0.0825 P=1.4 MULT=1
MM1002 A_1248_128# N_A_27_74#_M1002_g N_A_1000_424#_M1012_d VNB NLOWVT L=0.15
+ W=0.42 AD=0.0441 AS=0.169754 PD=0.63 PS=1.45485 NRD=14.28 NRS=0 M=1 R=2.8
+ SA=75002.9 SB=75000.6 A=0.063 P=1.14 MULT=1
MM1010 N_VGND_M1010_d N_A_1290_102#_M1010_g A_1248_128# VNB NLOWVT L=0.15 W=0.42
+ AD=0.1533 AS=0.0441 PD=1.57 PS=0.63 NRD=22.848 NRS=14.28 M=1 R=2.8 SA=75003.3
+ SB=75000.3 A=0.063 P=1.14 MULT=1
MM1021 N_VGND_M1021_d N_A_1000_424#_M1021_g N_A_1290_102#_M1021_s VNB NLOWVT
+ L=0.15 W=0.74 AD=0.12025 AS=0.2109 PD=1.065 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75001.2 A=0.111 P=1.78 MULT=1
MM1003 N_Q_M1003_d N_A_1290_102#_M1003_g N_VGND_M1021_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.12025 PD=1.02 PS=1.065 NRD=0 NRS=7.296 M=1 R=4.93333 SA=75000.7
+ SB=75000.7 A=0.111 P=1.78 MULT=1
MM1013 N_Q_M1003_d N_A_1290_102#_M1013_g N_VGND_M1013_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.2627 PD=1.02 PS=2.19 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75001.1
+ SB=75000.3 A=0.111 P=1.78 MULT=1
MM1027 N_VGND_M1027_d N_A_1290_102#_M1027_g N_A_1835_368#_M1027_s VNB NLOWVT
+ L=0.15 W=0.64 AD=0.133426 AS=0.1824 PD=1.06203 PS=1.85 NRD=23.904 NRS=0 M=1
+ R=4.26667 SA=75000.2 SB=75001.2 A=0.096 P=1.58 MULT=1
MM1006 N_Q_N_M1006_d N_A_1835_368#_M1006_g N_VGND_M1027_d VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.154274 PD=1.02 PS=1.22797 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.7 SB=75000.6 A=0.111 P=1.78 MULT=1
MM1008 N_Q_N_M1006_d N_A_1835_368#_M1008_g N_VGND_M1008_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.2109 PD=1.02 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75001.1 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1017 N_VPWR_M1017_d N_CLK_M1017_g N_A_27_74#_M1017_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.3304 PD=1.42 PS=2.83 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1016 N_A_206_368#_M1016_d N_A_27_74#_M1016_g N_VPWR_M1017_d VPB PSHORT L=0.15
+ W=1.12 AD=0.3304 AS=0.168 PD=2.83 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.7 SB=75000.2 A=0.168 P=2.54 MULT=1
MM1022 N_A_451_503#_M1022_d N_D_M1022_g N_VPWR_M1022_s VPB PSHORT L=0.15 W=0.42
+ AD=0.106225 AS=0.3234 PD=1.095 PS=2.38 NRD=92.8264 NRS=335.353 M=1 R=2.8
+ SA=75000.4 SB=75002.2 A=0.063 P=1.14 MULT=1
MM1028 N_A_558_445#_M1028_d N_A_206_368#_M1028_g N_A_451_503#_M1022_d VPB PSHORT
+ L=0.15 W=0.42 AD=0.1197 AS=0.106225 PD=0.99 PS=1.095 NRD=72.693 NRS=4.6886 M=1
+ R=2.8 SA=75000.5 SB=75004.6 A=0.063 P=1.14 MULT=1
MM1029 A_702_445# N_A_27_74#_M1029_g N_A_558_445#_M1028_d VPB PSHORT L=0.15
+ W=0.42 AD=0.0567 AS=0.1197 PD=0.69 PS=0.99 NRD=37.5088 NRS=63.3158 M=1 R=2.8
+ SA=75001.2 SB=75003.8 A=0.063 P=1.14 MULT=1
MM1005 N_VPWR_M1005_d N_A_753_284#_M1005_g A_702_445# VPB PSHORT L=0.15 W=0.42
+ AD=0.137692 AS=0.0567 PD=1.03 PS=0.69 NRD=127.971 NRS=37.5088 M=1 R=2.8
+ SA=75001.6 SB=75003.4 A=0.063 P=1.14 MULT=1
MM1031 N_A_753_284#_M1031_d N_A_558_445#_M1031_g N_VPWR_M1005_d VPB PSHORT
+ L=0.15 W=0.84 AD=0.126 AS=0.275383 PD=1.14 PS=2.06 NRD=2.3443 NRS=63.9856 M=1
+ R=5.6 SA=75001.2 SB=75002.5 A=0.126 P=1.98 MULT=1
MM1000 N_A_1000_424#_M1000_d N_A_27_74#_M1000_g N_A_753_284#_M1031_d VPB PSHORT
+ L=0.15 W=0.84 AD=0.3234 AS=0.126 PD=2.30667 PS=1.14 NRD=93.7917 NRS=2.3443 M=1
+ R=5.6 SA=75001.7 SB=75002 A=0.126 P=1.98 MULT=1
MM1030 A_1208_479# N_A_206_368#_M1030_g N_A_1000_424#_M1000_d VPB PSHORT L=0.15
+ W=0.42 AD=0.08925 AS=0.1617 PD=0.845 PS=1.15333 NRD=73.875 NRS=98.4803 M=1
+ R=2.8 SA=75003 SB=75002.8 A=0.063 P=1.14 MULT=1
MM1032 N_VPWR_M1032_d N_A_1290_102#_M1032_g A_1208_479# VPB PSHORT L=0.15 W=0.42
+ AD=0.0945 AS=0.08925 PD=0.833333 PS=0.845 NRD=4.6886 NRS=73.875 M=1 R=2.8
+ SA=75003.6 SB=75002.2 A=0.063 P=1.14 MULT=1
MM1015 N_A_1290_102#_M1015_d N_A_1000_424#_M1015_g N_VPWR_M1032_d VPB PSHORT
+ L=0.15 W=0.84 AD=0.126 AS=0.189 PD=1.14 PS=1.66667 NRD=2.3443 NRS=28.1316 M=1
+ R=5.6 SA=75002.2 SB=75001.7 A=0.126 P=1.98 MULT=1
MM1020 N_A_1290_102#_M1015_d N_A_1000_424#_M1020_g N_VPWR_M1020_s VPB PSHORT
+ L=0.15 W=0.84 AD=0.126 AS=0.1704 PD=1.14 PS=1.29 NRD=2.3443 NRS=22.261 M=1
+ R=5.6 SA=75002.6 SB=75001.2 A=0.126 P=1.98 MULT=1
MM1001 N_Q_M1001_d N_A_1290_102#_M1001_g N_VPWR_M1020_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.2272 PD=1.42 PS=1.72 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75002.4 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1009 N_Q_M1001_d N_A_1290_102#_M1009_g N_VPWR_M1009_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.3304 PD=1.42 PS=2.83 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75002.9 SB=75000.2 A=0.168 P=2.54 MULT=1
MM1019 N_VPWR_M1019_d N_A_1290_102#_M1019_g N_A_1835_368#_M1019_s VPB PSHORT
+ L=0.15 W=1 AD=0.198302 AS=0.295 PD=1.41981 PS=2.59 NRD=19.0302 NRS=1.9503 M=1
+ R=6.66667 SA=75000.2 SB=75001.2 A=0.15 P=2.3 MULT=1
MM1018 N_Q_N_M1018_d N_A_1835_368#_M1018_g N_VPWR_M1019_d VPB PSHORT L=0.15
+ W=1.12 AD=0.168 AS=0.222098 PD=1.42 PS=1.59019 NRD=1.7533 NRS=1.7533 M=1
+ R=7.46667 SA=75000.7 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1023 N_Q_N_M1018_d N_A_1835_368#_M1023_g N_VPWR_M1023_s VPB PSHORT L=0.15
+ W=1.12 AD=0.168 AS=0.336 PD=1.42 PS=2.84 NRD=1.7533 NRS=2.6201 M=1 R=7.46667
+ SA=75001.1 SB=75000.2 A=0.168 P=2.54 MULT=1
DX33_noxref VNB VPB NWDIODE A=20.8198 P=27.12
c_128 VNB 0 8.25183e-20 $X=0 $Y=0
c_220 VPB 0 6.95252e-20 $X=0 $Y=3.085
*
.include "sky130_fd_sc_hs__dfxbp_2.pxi.spice"
*
.ends
*
*
