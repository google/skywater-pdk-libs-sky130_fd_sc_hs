* File: sky130_fd_sc_hs__dlygate4sd1_1.spice
* Created: Tue Sep  1 20:03:21 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hs__dlygate4sd1_1.pex.spice"
.subckt sky130_fd_sc_hs__dlygate4sd1_1  VNB VPB A VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A	A
* VPB	VPB
* VNB	VNB
MM1004 N_VGND_M1004_d N_A_M1004_g N_A_28_74#_M1004_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.15435 AS=0.1113 PD=1.155 PS=1.37 NRD=15.708 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1007 N_A_288_74#_M1007_d N_A_28_74#_M1007_g N_VGND_M1004_d VNB NLOWVT L=0.15
+ W=0.42 AD=0.1113 AS=0.15435 PD=1.37 PS=1.155 NRD=0 NRS=114.276 M=1 R=2.8
+ SA=75001.1 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1002 N_VGND_M1002_d N_A_288_74#_M1002_g N_A_405_138#_M1002_s VNB NLOWVT L=0.15
+ W=0.42 AD=0.0831672 AS=0.2562 PD=0.78569 PS=2.06 NRD=40.86 NRS=41.424 M=1
+ R=2.8 SA=75000.5 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1005 N_X_M1005_d N_A_405_138#_M1005_g N_VGND_M1002_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.1961 AS=0.146533 PD=2.01 PS=1.38431 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.7
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1006 N_VPWR_M1006_d N_A_M1006_g N_A_28_74#_M1006_s VPB PSHORT L=0.15 W=0.42
+ AD=0.18412 AS=0.1176 PD=1.00268 PS=1.4 NRD=14.0658 NRS=7.0329 M=1 R=2.8
+ SA=75000.2 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1001 N_A_288_74#_M1001_d N_A_28_74#_M1001_g N_VPWR_M1006_d VPB PSHORT L=0.18
+ W=1 AD=0.26 AS=0.43838 PD=2.52 PS=2.38732 NRD=0 NRS=75.8253 M=1 R=5.55556
+ SA=90000.7 SB=90000.2 A=0.18 P=2.36 MULT=1
MM1000 N_VPWR_M1000_d N_A_288_74#_M1000_g N_A_405_138#_M1000_s VPB PSHORT L=0.18
+ W=1 AD=0.183019 AS=0.58 PD=1.39151 PS=3.16 NRD=13.2778 NRS=62.0353 M=1
+ R=5.55556 SA=90000.5 SB=90000.7 A=0.18 P=2.36 MULT=1
MM1003 N_X_M1003_d N_A_405_138#_M1003_g N_VPWR_M1000_d VPB PSHORT L=0.15 W=1.12
+ AD=0.3136 AS=0.204981 PD=2.8 PS=1.55849 NRD=2.6201 NRS=1.7533 M=1 R=7.46667
+ SA=75000.9 SB=75000.2 A=0.168 P=2.54 MULT=1
DX8_noxref VNB VPB NWDIODE A=7.8492 P=12.16
*
.include "sky130_fd_sc_hs__dlygate4sd1_1.pxi.spice"
*
.ends
*
*
