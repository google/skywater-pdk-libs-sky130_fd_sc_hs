* File: sky130_fd_sc_hs__nand3b_4.pex.spice
* Created: Tue Sep  1 20:09:43 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HS__NAND3B_4%A_N 3 5 7 8 10 12 13 20 21
c51 20 0 5.29186e-20 $X=0.93 $Y=1.515
c52 10 0 9.68625e-20 $X=1.345 $Y=1.765
r53 19 21 46.0284 $w=4.15e-07 $l=1.65e-07 $layer=POLY_cond $X=0.93 $Y=1.557
+ $X2=1.095 $Y2=1.557
r54 19 20 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.93
+ $Y=1.515 $X2=0.93 $Y2=1.515
r55 17 19 4.69045 $w=4.15e-07 $l=3.5e-08 $layer=POLY_cond $X=0.895 $Y=1.557
+ $X2=0.93 $Y2=1.557
r56 13 20 2.67779 $w=6.68e-07 $l=1.5e-07 $layer=LI1_cond $X=0.76 $Y=1.665
+ $X2=0.76 $Y2=1.515
r57 10 12 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=1.345 $Y=1.765
+ $X2=1.345 $Y2=2.26
r58 8 10 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.27 $Y=1.69
+ $X2=1.345 $Y2=1.765
r59 8 21 89.734 $w=1.5e-07 $l=1.75e-07 $layer=POLY_cond $X=1.27 $Y=1.69
+ $X2=1.095 $Y2=1.69
r60 5 17 26.7644 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=0.895 $Y=1.765
+ $X2=0.895 $Y2=1.557
r61 5 7 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=0.895 $Y=1.765
+ $X2=0.895 $Y2=2.26
r62 1 17 12.0612 $w=4.15e-07 $l=9e-08 $layer=POLY_cond $X=0.805 $Y=1.557
+ $X2=0.895 $Y2=1.557
r63 1 3 292.277 $w=1.5e-07 $l=5.7e-07 $layer=POLY_cond $X=0.805 $Y=1.35
+ $X2=0.805 $Y2=0.78
.ends

.subckt PM_SKY130_FD_SC_HS__NAND3B_4%C 1 3 4 5 6 8 9 11 12 14 15 17 18 20 22 23
+ 24 25 29 41
c82 25 0 9.68625e-20 $X=3.12 $Y=1.665
c83 5 0 2.71579e-20 $X=1.485 $Y=1.3
r84 41 42 1.44024 $w=5.02e-07 $l=1.5e-08 $layer=POLY_cond $X=3.075 $Y=1.495
+ $X2=3.09 $Y2=1.495
r85 39 41 12.002 $w=5.02e-07 $l=1.25e-07 $layer=POLY_cond $X=2.95 $Y=1.495
+ $X2=3.075 $Y2=1.495
r86 39 40 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.95
+ $Y=1.515 $X2=2.95 $Y2=1.515
r87 37 39 31.2052 $w=5.02e-07 $l=3.25e-07 $layer=POLY_cond $X=2.625 $Y=1.495
+ $X2=2.95 $Y2=1.495
r88 35 37 1.44024 $w=5.02e-07 $l=1.5e-08 $layer=POLY_cond $X=2.61 $Y=1.495
+ $X2=2.625 $Y2=1.495
r89 35 36 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=2.61
+ $Y=1.515 $X2=2.61 $Y2=1.515
r90 33 35 1.92032 $w=5.02e-07 $l=2e-08 $layer=POLY_cond $X=2.59 $Y=1.495
+ $X2=2.61 $Y2=1.495
r91 31 32 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.93
+ $Y=1.515 $X2=1.93 $Y2=1.515
r92 29 33 7.72247 $w=5.02e-07 $l=9.40744e-08 $layer=POLY_cond $X=2.515 $Y=1.452
+ $X2=2.59 $Y2=1.495
r93 29 31 71.5055 $w=4.55e-07 $l=5.85e-07 $layer=POLY_cond $X=2.515 $Y=1.452
+ $X2=1.93 $Y2=1.452
r94 25 40 4.55617 $w=4.28e-07 $l=1.7e-07 $layer=LI1_cond $X=3.12 $Y=1.565
+ $X2=2.95 $Y2=1.565
r95 24 40 8.30831 $w=4.28e-07 $l=3.1e-07 $layer=LI1_cond $X=2.64 $Y=1.565
+ $X2=2.95 $Y2=1.565
r96 24 36 0.80403 $w=4.28e-07 $l=3e-08 $layer=LI1_cond $X=2.64 $Y=1.565 $X2=2.61
+ $Y2=1.565
r97 23 36 12.0604 $w=4.28e-07 $l=4.5e-07 $layer=LI1_cond $X=2.16 $Y=1.565
+ $X2=2.61 $Y2=1.565
r98 23 32 6.16423 $w=4.28e-07 $l=2.3e-07 $layer=LI1_cond $X=2.16 $Y=1.565
+ $X2=1.93 $Y2=1.565
r99 21 31 1.83347 $w=4.55e-07 $l=1.5e-08 $layer=POLY_cond $X=1.915 $Y=1.452
+ $X2=1.93 $Y2=1.452
r100 21 22 11.0167 $w=3.02e-07 $l=7.5e-08 $layer=POLY_cond $X=1.915 $Y=1.452
+ $X2=1.84 $Y2=1.452
r101 18 42 31.5089 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=3.09 $Y=1.225
+ $X2=3.09 $Y2=1.495
r102 18 20 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=3.09 $Y=1.225
+ $X2=3.09 $Y2=0.78
r103 15 41 31.5089 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=3.075 $Y=1.765
+ $X2=3.075 $Y2=1.495
r104 15 17 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.075 $Y=1.765
+ $X2=3.075 $Y2=2.4
r105 12 37 31.5089 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=2.625 $Y=1.765
+ $X2=2.625 $Y2=1.495
r106 12 14 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.625 $Y=1.765
+ $X2=2.625 $Y2=2.4
r107 9 33 31.5089 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=2.59 $Y=1.225
+ $X2=2.59 $Y2=1.495
r108 9 11 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=2.59 $Y=1.225
+ $X2=2.59 $Y2=0.78
r109 6 22 15.6242 $w=1.5e-07 $l=2.27e-07 $layer=POLY_cond $X=1.84 $Y=1.225
+ $X2=1.84 $Y2=1.452
r110 6 8 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=1.84 $Y=1.225
+ $X2=1.84 $Y2=0.78
r111 4 22 11.0167 $w=3.02e-07 $l=1.85753e-07 $layer=POLY_cond $X=1.765 $Y=1.3
+ $X2=1.84 $Y2=1.452
r112 4 5 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=1.765 $Y=1.3
+ $X2=1.485 $Y2=1.3
r113 1 5 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.41 $Y=1.225
+ $X2=1.485 $Y2=1.3
r114 1 3 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=1.41 $Y=1.225
+ $X2=1.41 $Y2=0.78
.ends

.subckt PM_SKY130_FD_SC_HS__NAND3B_4%A_89_172# 1 2 7 9 10 12 13 15 16 18 19 20
+ 21 23 24 26 28 29 30 32 37 38 42 46 50 51
c132 50 0 1.74867e-19 $X=1.35 $Y=1.095
c133 24 0 2.37294e-19 $X=5.32 $Y=1.26
c134 16 0 3.1443e-19 $X=4.535 $Y=1.185
r135 61 62 1.46653 $w=4.93e-07 $l=1.5e-08 $layer=POLY_cond $X=4.52 $Y=1.475
+ $X2=4.535 $Y2=1.475
r136 55 59 30.7972 $w=4.93e-07 $l=3.15e-07 $layer=POLY_cond $X=3.765 $Y=1.475
+ $X2=4.08 $Y2=1.475
r137 55 57 7.33266 $w=4.93e-07 $l=7.5e-08 $layer=POLY_cond $X=3.765 $Y=1.475
+ $X2=3.69 $Y2=1.475
r138 54 55 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=3.765
+ $Y=1.465 $X2=3.765 $Y2=1.465
r139 51 54 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=3.685 $Y=1.095
+ $X2=3.685 $Y2=1.465
r140 46 48 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=0.59 $Y=1.005
+ $X2=0.59 $Y2=1.095
r141 43 61 7.33266 $w=4.93e-07 $l=7.5e-08 $layer=POLY_cond $X=4.445 $Y=1.475
+ $X2=4.52 $Y2=1.475
r142 43 59 35.6856 $w=4.93e-07 $l=3.65e-07 $layer=POLY_cond $X=4.445 $Y=1.475
+ $X2=4.08 $Y2=1.475
r143 42 54 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=4.445 $Y=1.465
+ $X2=3.77 $Y2=1.465
r144 42 43 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=4.445
+ $Y=1.465 $X2=4.445 $Y2=1.465
r145 39 50 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.435 $Y=1.095
+ $X2=1.35 $Y2=1.095
r146 38 51 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.6 $Y=1.095
+ $X2=3.685 $Y2=1.095
r147 38 39 141.246 $w=1.68e-07 $l=2.165e-06 $layer=LI1_cond $X=3.6 $Y=1.095
+ $X2=1.435 $Y2=1.095
r148 36 50 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.35 $Y=1.18
+ $X2=1.35 $Y2=1.095
r149 36 37 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=1.35 $Y=1.18
+ $X2=1.35 $Y2=1.95
r150 32 37 6.84389 $w=1.9e-07 $l=1.30767e-07 $layer=LI1_cond $X=1.265 $Y=2.045
+ $X2=1.35 $Y2=1.95
r151 32 34 8.46412 $w=1.88e-07 $l=1.45e-07 $layer=LI1_cond $X=1.265 $Y=2.045
+ $X2=1.12 $Y2=2.045
r152 31 48 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.755 $Y=1.095
+ $X2=0.59 $Y2=1.095
r153 30 50 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.265 $Y=1.095
+ $X2=1.35 $Y2=1.095
r154 30 31 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=1.265 $Y=1.095
+ $X2=0.755 $Y2=1.095
r155 26 28 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=5.395 $Y=1.185
+ $X2=5.395 $Y2=0.74
r156 25 29 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.04 $Y=1.26
+ $X2=4.965 $Y2=1.26
r157 24 26 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.32 $Y=1.26
+ $X2=5.395 $Y2=1.185
r158 24 25 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=5.32 $Y=1.26
+ $X2=5.04 $Y2=1.26
r159 21 29 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.965 $Y=1.185
+ $X2=4.965 $Y2=1.26
r160 21 23 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=4.965 $Y=1.185
+ $X2=4.965 $Y2=0.74
r161 20 62 32.9464 $w=4.93e-07 $l=2.497e-07 $layer=POLY_cond $X=4.61 $Y=1.26
+ $X2=4.535 $Y2=1.475
r162 19 29 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.89 $Y=1.26
+ $X2=4.965 $Y2=1.26
r163 19 20 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=4.89 $Y=1.26
+ $X2=4.61 $Y2=1.26
r164 16 62 31.0522 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=4.535 $Y=1.185
+ $X2=4.535 $Y2=1.475
r165 16 18 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=4.535 $Y=1.185
+ $X2=4.535 $Y2=0.74
r166 13 61 31.0522 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=4.52 $Y=1.765
+ $X2=4.52 $Y2=1.475
r167 13 15 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=4.52 $Y=1.765
+ $X2=4.52 $Y2=2.4
r168 10 59 31.0522 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=4.08 $Y=1.185
+ $X2=4.08 $Y2=1.475
r169 10 12 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=4.08 $Y=1.185
+ $X2=4.08 $Y2=0.74
r170 7 57 31.0522 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=3.69 $Y=1.765
+ $X2=3.69 $Y2=1.475
r171 7 9 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.69 $Y=1.765
+ $X2=3.69 $Y2=2.4
r172 2 34 600 $w=1.7e-07 $l=2.69768e-07 $layer=licon1_PDIFF $count=1 $X=0.97
+ $Y=1.84 $X2=1.12 $Y2=2.045
r173 1 46 182 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=1 $X=0.445
+ $Y=0.86 $X2=0.59 $Y2=1.005
.ends

.subckt PM_SKY130_FD_SC_HS__NAND3B_4%B 1 3 4 5 8 10 12 15 19 23 25 26 27 39 40
c71 40 0 6.5646e-20 $X=6.965 $Y=1.485
c72 39 0 1.64144e-19 $X=6.965 $Y=1.485
c73 8 0 1.10856e-19 $X=5.895 $Y=0.74
r74 39 40 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.965
+ $Y=1.485 $X2=6.965 $Y2=1.485
r75 37 39 25.8214 $w=3.92e-07 $l=2.1e-07 $layer=POLY_cond $X=6.755 $Y=1.542
+ $X2=6.965 $Y2=1.542
r76 36 37 52.8724 $w=3.92e-07 $l=4.3e-07 $layer=POLY_cond $X=6.325 $Y=1.542
+ $X2=6.755 $Y2=1.542
r77 34 36 46.7245 $w=3.92e-07 $l=3.8e-07 $layer=POLY_cond $X=5.945 $Y=1.542
+ $X2=6.325 $Y2=1.542
r78 34 35 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.945
+ $Y=1.485 $X2=5.945 $Y2=1.485
r79 32 34 4.30357 $w=3.92e-07 $l=3.5e-08 $layer=POLY_cond $X=5.91 $Y=1.542
+ $X2=5.945 $Y2=1.542
r80 31 32 1.84439 $w=3.92e-07 $l=1.5e-08 $layer=POLY_cond $X=5.895 $Y=1.542
+ $X2=5.91 $Y2=1.542
r81 27 40 0.127242 $w=4.68e-07 $l=5e-09 $layer=LI1_cond $X=6.96 $Y=1.415
+ $X2=6.965 $Y2=1.415
r82 26 27 12.2153 $w=4.68e-07 $l=4.8e-07 $layer=LI1_cond $X=6.48 $Y=1.415
+ $X2=6.96 $Y2=1.415
r83 25 26 12.2153 $w=4.68e-07 $l=4.8e-07 $layer=LI1_cond $X=6 $Y=1.415 $X2=6.48
+ $Y2=1.415
r84 25 35 1.39967 $w=4.68e-07 $l=5.5e-08 $layer=LI1_cond $X=6 $Y=1.415 $X2=5.945
+ $Y2=1.415
r85 21 39 27.051 $w=3.92e-07 $l=3.13247e-07 $layer=POLY_cond $X=7.185 $Y=1.32
+ $X2=6.965 $Y2=1.542
r86 21 23 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=7.185 $Y=1.32
+ $X2=7.185 $Y2=0.74
r87 17 37 25.3688 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=6.755 $Y=1.32
+ $X2=6.755 $Y2=1.542
r88 17 19 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=6.755 $Y=1.32
+ $X2=6.755 $Y2=0.74
r89 13 36 25.3688 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=6.325 $Y=1.32
+ $X2=6.325 $Y2=1.542
r90 13 15 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=6.325 $Y=1.32
+ $X2=6.325 $Y2=0.74
r91 10 32 25.3688 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=5.91 $Y=1.765
+ $X2=5.91 $Y2=1.542
r92 10 12 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=5.91 $Y=1.765
+ $X2=5.91 $Y2=2.4
r93 6 31 25.3688 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=5.895 $Y=1.32
+ $X2=5.895 $Y2=1.542
r94 6 8 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=5.895 $Y=1.32
+ $X2=5.895 $Y2=0.74
r95 4 31 38.2027 $w=3.92e-07 $l=2.01903e-07 $layer=POLY_cond $X=5.74 $Y=1.65
+ $X2=5.895 $Y2=1.542
r96 4 5 97.4255 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=5.74 $Y=1.65 $X2=5.55
+ $Y2=1.65
r97 1 5 26.9307 $w=1.5e-07 $l=1.53542e-07 $layer=POLY_cond $X=5.46 $Y=1.765
+ $X2=5.55 $Y2=1.65
r98 1 3 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=5.46 $Y=1.765
+ $X2=5.46 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_HS__NAND3B_4%VPWR 1 2 3 4 5 16 18 22 24 26 33 48 54 56
+ 61 64 76 79
c69 76 0 1.64144e-19 $X=7.4 $Y=2.325
r70 78 79 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r71 76 78 0.461248 $w=1.058e-06 $l=4e-08 $layer=LI1_cond $X=7.4 $Y=2.787
+ $X2=7.44 $Y2=2.787
r72 74 76 9.74386 $w=1.058e-06 $l=8.45e-07 $layer=LI1_cond $X=6.555 $Y=2.787
+ $X2=7.4 $Y2=2.787
r73 72 79 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=7.44 $Y2=3.33
r74 71 74 0.864839 $w=1.058e-06 $l=7.5e-08 $layer=LI1_cond $X=6.48 $Y=2.787
+ $X2=6.555 $Y2=2.787
r75 71 72 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r76 69 71 3.97826 $w=1.058e-06 $l=3.45e-07 $layer=LI1_cond $X=6.135 $Y=2.787
+ $X2=6.48 $Y2=2.787
r77 67 72 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=3.33 $X2=6.48
+ $Y2=3.33
r78 66 69 1.55671 $w=1.058e-06 $l=1.35e-07 $layer=LI1_cond $X=6 $Y=2.787
+ $X2=6.135 $Y2=2.787
r79 66 67 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r80 63 64 11.2171 $w=7.63e-07 $l=1.65e-07 $layer=LI1_cond $X=5.235 $Y=3.032
+ $X2=5.4 $Y2=3.032
r81 60 67 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.04 $Y=3.33 $X2=6
+ $Y2=3.33
r82 59 63 3.04883 $w=7.63e-07 $l=1.95e-07 $layer=LI1_cond $X=5.04 $Y=3.032
+ $X2=5.235 $Y2=3.032
r83 59 61 15.8294 $w=7.63e-07 $l=4.6e-07 $layer=LI1_cond $X=5.04 $Y=3.032
+ $X2=4.58 $Y2=3.032
r84 59 60 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r85 56 57 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r86 53 54 11.2171 $w=7.63e-07 $l=1.65e-07 $layer=LI1_cond $X=2.4 $Y=3.032
+ $X2=2.565 $Y2=3.032
r87 50 53 3.7524 $w=7.63e-07 $l=2.4e-07 $layer=LI1_cond $X=2.16 $Y=3.032 $X2=2.4
+ $Y2=3.032
r88 50 51 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r89 47 50 7.89568 $w=7.63e-07 $l=5.05e-07 $layer=LI1_cond $X=1.655 $Y=3.032
+ $X2=2.16 $Y2=3.032
r90 47 48 11.2171 $w=7.63e-07 $l=1.65e-07 $layer=LI1_cond $X=1.655 $Y=3.032
+ $X2=1.49 $Y2=3.032
r91 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r92 42 60 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=5.04 $Y2=3.33
r93 41 61 1.30481 $w=1.68e-07 $l=2e-08 $layer=LI1_cond $X=4.56 $Y=3.33 $X2=4.58
+ $Y2=3.33
r94 41 42 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r95 39 56 11.2236 $w=1.7e-07 $l=2.48e-07 $layer=LI1_cond $X=3.63 $Y=3.33
+ $X2=3.382 $Y2=3.33
r96 39 41 60.6738 $w=1.68e-07 $l=9.3e-07 $layer=LI1_cond $X=3.63 $Y=3.33
+ $X2=4.56 $Y2=3.33
r97 37 57 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=3.6 $Y2=3.33
r98 37 51 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=2.16 $Y2=3.33
r99 36 54 36.2086 $w=1.68e-07 $l=5.55e-07 $layer=LI1_cond $X=3.12 $Y=3.33
+ $X2=2.565 $Y2=3.33
r100 36 37 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r101 33 56 11.2236 $w=1.7e-07 $l=2.47e-07 $layer=LI1_cond $X=3.135 $Y=3.33
+ $X2=3.382 $Y2=3.33
r102 33 36 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=3.135 $Y=3.33
+ $X2=3.12 $Y2=3.33
r103 32 51 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.16 $Y2=3.33
r104 32 45 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.24 $Y2=3.33
r105 31 48 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=1.2 $Y=3.33
+ $X2=1.49 $Y2=3.33
r106 31 32 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r107 29 44 4.73185 $w=1.7e-07 $l=2.23e-07 $layer=LI1_cond $X=0.445 $Y=3.33
+ $X2=0.222 $Y2=3.33
r108 29 31 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=0.445 $Y=3.33
+ $X2=1.2 $Y2=3.33
r109 26 42 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=3.84 $Y=3.33
+ $X2=4.56 $Y2=3.33
r110 26 57 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=3.84 $Y=3.33
+ $X2=3.6 $Y2=3.33
r111 24 66 11.613 $w=1.058e-06 $l=5.57798e-07 $layer=LI1_cond $X=5.97 $Y=3.33
+ $X2=6 $Y2=2.787
r112 24 64 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=5.97 $Y=3.33
+ $X2=5.4 $Y2=3.33
r113 20 56 2.04857 $w=4.95e-07 $l=8.5e-08 $layer=LI1_cond $X=3.382 $Y=3.245
+ $X2=3.382 $Y2=3.33
r114 20 22 10.3902 $w=4.93e-07 $l=4.3e-07 $layer=LI1_cond $X=3.382 $Y=3.245
+ $X2=3.382 $Y2=2.815
r115 16 44 3.03433 $w=3.3e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.28 $Y=3.245
+ $X2=0.222 $Y2=3.33
r116 16 18 26.1919 $w=3.28e-07 $l=7.5e-07 $layer=LI1_cond $X=0.28 $Y=3.245
+ $X2=0.28 $Y2=2.495
r117 5 76 200 $w=1.7e-07 $l=1.63966e-06 $layer=licon1_PDIFF $count=3 $X=5.985
+ $Y=1.84 $X2=7.4 $Y2=2.325
r118 5 74 200 $w=1.7e-07 $l=7.75468e-07 $layer=licon1_PDIFF $count=3 $X=5.985
+ $Y=1.84 $X2=6.555 $Y2=2.325
r119 5 69 600 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=5.985
+ $Y=1.84 $X2=6.135 $Y2=2.815
r120 4 63 300 $w=1.7e-07 $l=1.25484e-06 $layer=licon1_PDIFF $count=2 $X=4.595
+ $Y=1.84 $X2=5.235 $Y2=2.815
r121 3 22 600 $w=1.7e-07 $l=1.08392e-06 $layer=licon1_PDIFF $count=1 $X=3.15
+ $Y=1.84 $X2=3.38 $Y2=2.815
r122 2 53 300 $w=1.7e-07 $l=1.38416e-06 $layer=licon1_PDIFF $count=2 $X=1.42
+ $Y=1.84 $X2=2.4 $Y2=2.815
r123 2 47 600 $w=1.7e-07 $l=1.08616e-06 $layer=licon1_PDIFF $count=1 $X=1.42
+ $Y=1.84 $X2=1.655 $Y2=2.815
r124 1 18 600 $w=1.7e-07 $l=7.23878e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.495
.ends

.subckt PM_SKY130_FD_SC_HS__NAND3B_4%Y 1 2 3 4 5 20 21 24 30 32 34 35 36 37 41
c70 41 0 1.74292e-19 $X=5.04 $Y=1.13
c71 36 0 1.10856e-19 $X=5.04 $Y=1.295
c72 34 0 1.70138e-19 $X=5.04 $Y=1.98
r73 36 37 18.5393 $w=2.28e-07 $l=3.7e-07 $layer=LI1_cond $X=5.04 $Y=1.295
+ $X2=5.04 $Y2=1.665
r74 36 41 8.26753 $w=2.28e-07 $l=1.65e-07 $layer=LI1_cond $X=5.04 $Y=1.295
+ $X2=5.04 $Y2=1.13
r75 35 41 3.90668 $w=2.3e-07 $l=2.22486e-07 $layer=LI1_cond $X=5.135 $Y=0.95
+ $X2=5.04 $Y2=1.13
r76 33 37 7.76646 $w=2.28e-07 $l=1.55e-07 $layer=LI1_cond $X=5.04 $Y=1.82
+ $X2=5.04 $Y2=1.665
r77 33 34 2.55462 $w=2.3e-07 $l=1.6e-07 $layer=LI1_cond $X=5.04 $Y=1.82 $X2=5.04
+ $Y2=1.98
r78 28 34 3.89311 $w=3.2e-07 $l=1.15e-07 $layer=LI1_cond $X=5.155 $Y=1.98
+ $X2=5.04 $Y2=1.98
r79 28 30 19.0873 $w=3.18e-07 $l=5.3e-07 $layer=LI1_cond $X=5.155 $Y=1.98
+ $X2=5.685 $Y2=1.98
r80 24 35 3.19638 $w=3.3e-07 $l=2.17371e-07 $layer=LI1_cond $X=4.925 $Y=0.965
+ $X2=5.135 $Y2=0.95
r81 24 26 21.652 $w=3.28e-07 $l=6.2e-07 $layer=LI1_cond $X=4.925 $Y=0.965
+ $X2=4.305 $Y2=0.965
r82 21 32 7.64885 $w=3.18e-07 $l=1.6e-07 $layer=LI1_cond $X=3.91 $Y=1.98
+ $X2=3.75 $Y2=1.98
r83 21 23 13.8653 $w=3.18e-07 $l=3.85e-07 $layer=LI1_cond $X=3.91 $Y=1.98
+ $X2=4.295 $Y2=1.98
r84 20 34 3.89311 $w=3.2e-07 $l=1.15e-07 $layer=LI1_cond $X=4.925 $Y=1.98
+ $X2=5.04 $Y2=1.98
r85 20 23 22.6887 $w=3.18e-07 $l=6.3e-07 $layer=LI1_cond $X=4.925 $Y=1.98
+ $X2=4.295 $Y2=1.98
r86 18 32 52.5359 $w=1.88e-07 $l=9e-07 $layer=LI1_cond $X=2.85 $Y=2.045 $X2=3.75
+ $Y2=2.045
r87 5 30 600 $w=1.7e-07 $l=2.43721e-07 $layer=licon1_PDIFF $count=1 $X=5.535
+ $Y=1.84 $X2=5.685 $Y2=2.02
r88 4 23 300 $w=1.7e-07 $l=5.98122e-07 $layer=licon1_PDIFF $count=2 $X=3.765
+ $Y=1.84 $X2=4.295 $Y2=1.985
r89 3 18 600 $w=1.7e-07 $l=2.69768e-07 $layer=licon1_PDIFF $count=1 $X=2.7
+ $Y=1.84 $X2=2.85 $Y2=2.045
r90 2 35 182 $w=1.7e-07 $l=6.0597e-07 $layer=licon1_NDIFF $count=1 $X=5.04
+ $Y=0.37 $X2=5.18 $Y2=0.91
r91 1 26 182 $w=1.7e-07 $l=6.65789e-07 $layer=licon1_NDIFF $count=1 $X=4.155
+ $Y=0.37 $X2=4.305 $Y2=0.965
.ends

.subckt PM_SKY130_FD_SC_HS__NAND3B_4%VGND 1 2 3 12 15 22 23 24 30 42 43 47
c67 1 0 1.74867e-19 $X=0.88 $Y=0.41
r68 47 50 8.17727 $w=4.88e-07 $l=3.35e-07 $layer=LI1_cond $X=2.215 $Y=0
+ $X2=2.215 $Y2=0.335
r69 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r70 42 43 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=7.44 $Y=0
+ $X2=7.44 $Y2=0
r71 39 42 250.524 $w=1.68e-07 $l=3.84e-06 $layer=LI1_cond $X=3.6 $Y=0 $X2=7.44
+ $Y2=0
r72 39 40 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=3.6 $Y=0
+ $X2=3.6 $Y2=0
r73 37 40 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=3.6
+ $Y2=0
r74 37 48 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=2.16
+ $Y2=0
r75 36 37 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r76 34 47 7.03003 $w=1.7e-07 $l=2.45e-07 $layer=LI1_cond $X=2.46 $Y=0 $X2=2.215
+ $Y2=0
r77 34 36 43.0588 $w=1.68e-07 $l=6.6e-07 $layer=LI1_cond $X=2.46 $Y=0 $X2=3.12
+ $Y2=0
r78 33 48 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r79 32 33 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r80 30 47 7.03003 $w=1.7e-07 $l=2.45e-07 $layer=LI1_cond $X=1.97 $Y=0 $X2=2.215
+ $Y2=0
r81 30 32 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=1.97 $Y=0 $X2=1.68
+ $Y2=0
r82 28 33 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r83 27 28 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r84 24 43 1.00344 $w=4.9e-07 $l=3.6e-06 $layer=MET1_cond $X=3.84 $Y=0 $X2=7.44
+ $Y2=0
r85 24 40 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=3.84 $Y=0 $X2=3.6
+ $Y2=0
r86 22 36 1.30481 $w=1.68e-07 $l=2e-08 $layer=LI1_cond $X=3.14 $Y=0 $X2=3.12
+ $Y2=0
r87 22 23 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.14 $Y=0 $X2=3.305
+ $Y2=0
r88 21 39 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=3.47 $Y=0 $X2=3.6
+ $Y2=0
r89 21 23 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.47 $Y=0 $X2=3.305
+ $Y2=0
r90 17 32 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=1.28 $Y=0 $X2=1.68
+ $Y2=0
r91 15 27 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=0.935 $Y=0 $X2=0.72
+ $Y2=0
r92 15 19 10.8563 $w=3.43e-07 $l=3.25e-07 $layer=LI1_cond $X=1.107 $Y=0
+ $X2=1.107 $Y2=0.325
r93 15 17 4.88813 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=1.107 $Y=0 $X2=1.28
+ $Y2=0
r94 10 23 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.305 $Y=0.085
+ $X2=3.305 $Y2=0
r95 10 12 18.5089 $w=3.28e-07 $l=5.3e-07 $layer=LI1_cond $X=3.305 $Y=0.085
+ $X2=3.305 $Y2=0.615
r96 3 12 182 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_NDIFF $count=1 $X=3.165
+ $Y=0.41 $X2=3.305 $Y2=0.615
r97 2 50 182 $w=1.7e-07 $l=3.3541e-07 $layer=licon1_NDIFF $count=1 $X=1.915
+ $Y=0.41 $X2=2.215 $Y2=0.335
r98 1 19 182 $w=1.7e-07 $l=2.64102e-07 $layer=licon1_NDIFF $count=1 $X=0.88
+ $Y=0.41 $X2=1.105 $Y2=0.325
.ends

.subckt PM_SKY130_FD_SC_HS__NAND3B_4%A_297_82# 1 2 3 4 14 16 17 18 20 21 22 23
+ 25 32 33 34 36 39 40 42
c126 39 0 2.57607e-20 $X=1.46 $Y=0.615
r127 42 44 4.88915 $w=3.28e-07 $l=1.4e-07 $layer=LI1_cond $X=2.805 $Y=0.615
+ $X2=2.805 $Y2=0.755
r128 38 40 9.22412 $w=4.48e-07 $l=1.65e-07 $layer=LI1_cond $X=1.625 $Y=0.615
+ $X2=1.79 $Y2=0.615
r129 38 39 9.22412 $w=4.48e-07 $l=1.65e-07 $layer=LI1_cond $X=1.625 $Y=0.615
+ $X2=1.46 $Y2=0.615
r130 35 36 52.8449 $w=1.68e-07 $l=8.1e-07 $layer=LI1_cond $X=7.33 $Y=1.01
+ $X2=7.33 $Y2=1.82
r131 33 36 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.245 $Y=1.905
+ $X2=7.33 $Y2=1.82
r132 33 34 66.2193 $w=1.68e-07 $l=1.015e-06 $layer=LI1_cond $X=7.245 $Y=1.905
+ $X2=6.23 $Y2=1.905
r133 31 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.145 $Y=1.99
+ $X2=6.23 $Y2=1.905
r134 31 32 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=6.145 $Y=1.99
+ $X2=6.145 $Y2=2.31
r135 27 30 56.107 $w=1.68e-07 $l=8.6e-07 $layer=LI1_cond $X=6.11 $Y=0.925
+ $X2=6.97 $Y2=0.925
r136 25 35 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.245 $Y=0.925
+ $X2=7.33 $Y2=1.01
r137 25 30 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=7.245 $Y=0.925
+ $X2=6.97 $Y2=0.925
r138 23 44 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.64 $Y=0.755
+ $X2=2.805 $Y2=0.755
r139 23 40 55.4545 $w=1.68e-07 $l=8.5e-07 $layer=LI1_cond $X=2.64 $Y=0.755
+ $X2=1.79 $Y2=0.755
r140 21 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.06 $Y=2.395
+ $X2=6.145 $Y2=2.31
r141 21 22 344.144 $w=1.68e-07 $l=5.275e-06 $layer=LI1_cond $X=6.06 $Y=2.395
+ $X2=0.785 $Y2=2.395
r142 20 22 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.7 $Y=2.31
+ $X2=0.785 $Y2=2.395
r143 19 20 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=0.7 $Y=2.12 $X2=0.7
+ $Y2=2.31
r144 17 19 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.615 $Y=2.035
+ $X2=0.7 $Y2=2.12
r145 17 18 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=0.615 $Y=2.035
+ $X2=0.255 $Y2=2.035
r146 16 39 78.615 $w=1.68e-07 $l=1.205e-06 $layer=LI1_cond $X=0.255 $Y=0.665
+ $X2=1.46 $Y2=0.665
r147 14 18 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.17 $Y=1.95
+ $X2=0.255 $Y2=2.035
r148 13 16 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.17 $Y=0.75
+ $X2=0.255 $Y2=0.665
r149 13 14 78.2888 $w=1.68e-07 $l=1.2e-06 $layer=LI1_cond $X=0.17 $Y=0.75
+ $X2=0.17 $Y2=1.95
r150 4 30 182 $w=1.7e-07 $l=6.21068e-07 $layer=licon1_NDIFF $count=1 $X=6.83
+ $Y=0.37 $X2=6.97 $Y2=0.925
r151 3 27 182 $w=1.7e-07 $l=6.21068e-07 $layer=licon1_NDIFF $count=1 $X=5.97
+ $Y=0.37 $X2=6.11 $Y2=0.925
r152 2 42 182 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_NDIFF $count=1 $X=2.665
+ $Y=0.41 $X2=2.805 $Y2=0.615
r153 1 38 182 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_NDIFF $count=1 $X=1.485
+ $Y=0.41 $X2=1.625 $Y2=0.615
.ends

.subckt PM_SKY130_FD_SC_HS__NAND3B_4%A_744_74# 1 2 3 4 5 20 24 29 32
c35 32 0 1.71648e-19 $X=5.515 $Y=0.51
c36 29 0 1.40137e-19 $X=4.03 $Y=0.49
r37 31 32 6.52497 $w=3.18e-07 $l=1.65e-07 $layer=LI1_cond $X=5.68 $Y=0.51
+ $X2=5.515 $Y2=0.51
r38 27 29 6.95017 $w=2.78e-07 $l=1.65e-07 $layer=LI1_cond $X=3.865 $Y=0.49
+ $X2=4.03 $Y2=0.49
r39 22 24 30.9719 $w=3.18e-07 $l=8.6e-07 $layer=LI1_cond $X=6.54 $Y=0.51 $X2=7.4
+ $Y2=0.51
r40 20 31 5.58215 $w=3.18e-07 $l=1.55e-07 $layer=LI1_cond $X=5.835 $Y=0.51
+ $X2=5.68 $Y2=0.51
r41 20 22 25.3898 $w=3.18e-07 $l=7.05e-07 $layer=LI1_cond $X=5.835 $Y=0.51
+ $X2=6.54 $Y2=0.51
r42 19 32 35.2648 $w=2.48e-07 $l=7.65e-07 $layer=LI1_cond $X=4.75 $Y=0.475
+ $X2=5.515 $Y2=0.475
r43 19 29 33.1904 $w=2.48e-07 $l=7.2e-07 $layer=LI1_cond $X=4.75 $Y=0.475
+ $X2=4.03 $Y2=0.475
r44 5 24 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=7.26 $Y=0.37
+ $X2=7.4 $Y2=0.55
r45 4 22 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=6.4 $Y=0.37
+ $X2=6.54 $Y2=0.55
r46 3 31 182 $w=1.7e-07 $l=2.86182e-07 $layer=licon1_NDIFF $count=1 $X=5.47
+ $Y=0.37 $X2=5.68 $Y2=0.55
r47 2 19 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=4.61
+ $Y=0.37 $X2=4.75 $Y2=0.515
r48 1 27 182 $w=1.7e-07 $l=2.20907e-07 $layer=licon1_NDIFF $count=1 $X=3.72
+ $Y=0.37 $X2=3.865 $Y2=0.53
.ends

