* File: sky130_fd_sc_hs__nand4bb_4.spice
* Created: Thu Aug 27 20:52:46 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hs__nand4bb_4.pex.spice"
.subckt sky130_fd_sc_hs__nand4bb_4  VNB VPB A_N B_N C D VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* D	D
* C	C
* B_N	B_N
* A_N	A_N
* VPB	VPB
* VNB	VNB
MM1019 N_VGND_M1019_d N_A_N_M1019_g N_A_27_114#_M1019_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.21935 AS=0.2109 PD=1.57 PS=2.05 NRD=39.144 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75000.8 A=0.111 P=1.78 MULT=1
MM1022 N_A_232_114#_M1022_d N_B_N_M1022_g N_VGND_M1019_d VNB NLOWVT L=0.15
+ W=0.74 AD=0.2368 AS=0.21935 PD=2.12 PS=1.57 NRD=2.424 NRS=39.144 M=1 R=4.93333
+ SA=75000.8 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1000 N_A_374_74#_M1000_d N_A_27_114#_M1000_g N_Y_M1000_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.2109 AS=0.14245 PD=2.05 PS=1.125 NRD=0 NRS=6.48 M=1 R=4.93333
+ SA=75000.2 SB=75003.5 A=0.111 P=1.78 MULT=1
MM1005 N_A_374_74#_M1005_d N_A_27_114#_M1005_g N_Y_M1000_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1073 AS=0.14245 PD=1.03 PS=1.125 NRD=0.804 NRS=10.536 M=1
+ R=4.93333 SA=75000.7 SB=75003 A=0.111 P=1.78 MULT=1
MM1011 N_A_374_74#_M1005_d N_A_27_114#_M1011_g N_Y_M1011_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1073 AS=0.1036 PD=1.03 PS=1.02 NRD=0.804 NRS=0 M=1 R=4.93333
+ SA=75001.2 SB=75002.5 A=0.111 P=1.78 MULT=1
MM1031 N_A_374_74#_M1031_d N_A_27_114#_M1031_g N_Y_M1011_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75001.6 SB=75002.1 A=0.111 P=1.78 MULT=1
MM1002 N_A_828_74#_M1002_d N_A_232_114#_M1002_g N_A_374_74#_M1031_d VNB NLOWVT
+ L=0.15 W=0.74 AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75002 SB=75001.7 A=0.111 P=1.78 MULT=1
MM1007 N_A_828_74#_M1002_d N_A_232_114#_M1007_g N_A_374_74#_M1007_s VNB NLOWVT
+ L=0.15 W=0.74 AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75002.5 SB=75001.2 A=0.111 P=1.78 MULT=1
MM1017 N_A_828_74#_M1017_d N_A_232_114#_M1017_g N_A_374_74#_M1007_s VNB NLOWVT
+ L=0.15 W=0.74 AD=0.1657 AS=0.1036 PD=1.2 PS=1.02 NRD=12.972 NRS=0 M=1
+ R=4.93333 SA=75002.9 SB=75000.8 A=0.111 P=1.78 MULT=1
MM1028 N_A_828_74#_M1017_d N_A_232_114#_M1028_g N_A_374_74#_M1028_s VNB NLOWVT
+ L=0.15 W=0.74 AD=0.1657 AS=0.2109 PD=1.2 PS=2.05 NRD=12.972 NRS=0 M=1
+ R=4.93333 SA=75003.5 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1023 N_A_828_74#_M1023_d N_C_M1023_g N_A_1229_74#_M1023_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.2109 PD=1.02 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75003.3 A=0.111 P=1.78 MULT=1
MM1024 N_A_828_74#_M1023_d N_C_M1024_g N_A_1229_74#_M1024_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.6 SB=75002.9 A=0.111 P=1.78 MULT=1
MM1036 N_A_828_74#_M1036_d N_C_M1036_g N_A_1229_74#_M1024_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75001.1 SB=75002.4 A=0.111 P=1.78 MULT=1
MM1037 N_A_828_74#_M1036_d N_C_M1037_g N_A_1229_74#_M1037_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75001.5 SB=75002 A=0.111 P=1.78 MULT=1
MM1003 N_A_1229_74#_M1037_s N_D_M1003_g N_VGND_M1003_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.9
+ SB=75001.6 A=0.111 P=1.78 MULT=1
MM1008 N_A_1229_74#_M1008_d N_D_M1008_g N_VGND_M1003_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75002.4
+ SB=75001.1 A=0.111 P=1.78 MULT=1
MM1013 N_A_1229_74#_M1008_d N_D_M1013_g N_VGND_M1013_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1295 PD=1.02 PS=1.09 NRD=0 NRS=0 M=1 R=4.93333 SA=75002.8
+ SB=75000.7 A=0.111 P=1.78 MULT=1
MM1034 N_A_1229_74#_M1034_d N_D_M1034_g N_VGND_M1013_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.1295 PD=2.05 PS=1.09 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75003.3
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1025 N_A_27_114#_M1025_d N_A_N_M1025_g N_VPWR_M1025_s VPB PSHORT L=0.15 W=0.84
+ AD=0.126 AS=0.2478 PD=1.14 PS=2.27 NRD=2.3443 NRS=2.3443 M=1 R=5.6 SA=75000.2
+ SB=75009.3 A=0.126 P=1.98 MULT=1
MM1026 N_A_27_114#_M1025_d N_A_N_M1026_g N_VPWR_M1026_s VPB PSHORT L=0.15 W=0.84
+ AD=0.126 AS=0.126 PD=1.14 PS=1.14 NRD=2.3443 NRS=2.3443 M=1 R=5.6 SA=75000.7
+ SB=75008.8 A=0.126 P=1.98 MULT=1
MM1029 N_A_232_114#_M1029_d N_B_N_M1029_g N_VPWR_M1026_s VPB PSHORT L=0.15
+ W=0.84 AD=0.126 AS=0.126 PD=1.14 PS=1.14 NRD=2.3443 NRS=2.3443 M=1 R=5.6
+ SA=75001.1 SB=75008.4 A=0.126 P=1.98 MULT=1
MM1032 N_A_232_114#_M1029_d N_B_N_M1032_g N_VPWR_M1032_s VPB PSHORT L=0.15
+ W=0.84 AD=0.126 AS=0.237 PD=1.14 PS=1.44857 NRD=2.3443 NRS=23.443 M=1 R=5.6
+ SA=75001.6 SB=75007.9 A=0.126 P=1.98 MULT=1
MM1020 N_Y_M1020_d N_A_27_114#_M1020_g N_VPWR_M1032_s VPB PSHORT L=0.15 W=1.12
+ AD=0.196 AS=0.316 PD=1.47 PS=1.93143 NRD=1.7533 NRS=33.4112 M=1 R=7.46667
+ SA=75001.8 SB=75007.2 A=0.168 P=2.54 MULT=1
MM1021 N_Y_M1020_d N_A_27_114#_M1021_g N_VPWR_M1021_s VPB PSHORT L=0.15 W=1.12
+ AD=0.196 AS=0.168 PD=1.47 PS=1.42 NRD=10.5395 NRS=1.7533 M=1 R=7.46667
+ SA=75002.3 SB=75006.7 A=0.168 P=2.54 MULT=1
MM1027 N_Y_M1027_d N_A_27_114#_M1027_g N_VPWR_M1021_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75002.7 SB=75006.3 A=0.168 P=2.54 MULT=1
MM1030 N_Y_M1027_d N_A_27_114#_M1030_g N_VPWR_M1030_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75003.2 SB=75005.8 A=0.168 P=2.54 MULT=1
MM1001 N_Y_M1001_d N_A_232_114#_M1001_g N_VPWR_M1030_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75003.6 SB=75005.4 A=0.168 P=2.54 MULT=1
MM1004 N_Y_M1001_d N_A_232_114#_M1004_g N_VPWR_M1004_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.196 PD=1.42 PS=1.47 NRD=1.7533 NRS=10.5395 M=1 R=7.46667
+ SA=75004.1 SB=75004.9 A=0.168 P=2.54 MULT=1
MM1033 N_Y_M1033_d N_A_232_114#_M1033_g N_VPWR_M1004_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.196 PD=1.42 PS=1.47 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75004.6 SB=75004.4 A=0.168 P=2.54 MULT=1
MM1035 N_Y_M1033_d N_A_232_114#_M1035_g N_VPWR_M1035_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667 SA=75005
+ SB=75004 A=0.168 P=2.54 MULT=1
MM1006 N_Y_M1006_d N_C_M1006_g N_VPWR_M1035_s VPB PSHORT L=0.15 W=1.12 AD=0.168
+ AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667 SA=75005.5
+ SB=75003.5 A=0.168 P=2.54 MULT=1
MM1009 N_Y_M1006_d N_C_M1009_g N_VPWR_M1009_s VPB PSHORT L=0.15 W=1.12 AD=0.168
+ AS=0.224 PD=1.42 PS=1.52 NRD=1.7533 NRS=10.5395 M=1 R=7.46667 SA=75005.9
+ SB=75003.1 A=0.168 P=2.54 MULT=1
MM1012 N_Y_M1012_d N_C_M1012_g N_VPWR_M1009_s VPB PSHORT L=0.15 W=1.12 AD=0.168
+ AS=0.224 PD=1.42 PS=1.52 NRD=1.7533 NRS=10.5395 M=1 R=7.46667 SA=75006.5
+ SB=75002.5 A=0.168 P=2.54 MULT=1
MM1014 N_Y_M1012_d N_C_M1014_g N_VPWR_M1014_s VPB PSHORT L=0.15 W=1.12 AD=0.168
+ AS=0.196 PD=1.42 PS=1.47 NRD=1.7533 NRS=1.7533 M=1 R=7.46667 SA=75006.9
+ SB=75002.1 A=0.168 P=2.54 MULT=1
MM1010 N_Y_M1010_d N_D_M1010_g N_VPWR_M1014_s VPB PSHORT L=0.15 W=1.12 AD=0.168
+ AS=0.196 PD=1.42 PS=1.47 NRD=1.7533 NRS=10.5395 M=1 R=7.46667 SA=75007.4
+ SB=75001.6 A=0.168 P=2.54 MULT=1
MM1015 N_Y_M1010_d N_D_M1015_g N_VPWR_M1015_s VPB PSHORT L=0.15 W=1.12 AD=0.168
+ AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667 SA=75007.9
+ SB=75001.1 A=0.168 P=2.54 MULT=1
MM1016 N_Y_M1016_d N_D_M1016_g N_VPWR_M1015_s VPB PSHORT L=0.15 W=1.12 AD=0.168
+ AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667 SA=75008.3
+ SB=75000.7 A=0.168 P=2.54 MULT=1
MM1018 N_Y_M1016_d N_D_M1018_g N_VPWR_M1018_s VPB PSHORT L=0.15 W=1.12 AD=0.168
+ AS=0.3304 PD=1.42 PS=2.83 NRD=1.7533 NRS=1.7533 M=1 R=7.46667 SA=75008.8
+ SB=75000.2 A=0.168 P=2.54 MULT=1
DX38_noxref VNB VPB NWDIODE A=19.4556 P=24.64
c_85 VNB 0 1.90128e-19 $X=0 $Y=0
*
.include "sky130_fd_sc_hs__nand4bb_4.pxi.spice"
*
.ends
*
*
