* File: sky130_fd_sc_hs__dlrbp_1.spice
* Created: Tue Sep  1 20:01:51 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hs__dlrbp_1.pex.spice"
.subckt sky130_fd_sc_hs__dlrbp_1  VNB VPB D GATE RESET_B VPWR Q Q_N VGND
* 
* VGND	VGND
* Q_N	Q_N
* Q	Q
* VPWR	VPWR
* RESET_B	RESET_B
* GATE	GATE
* D	D
* VPB	VPB
* VNB	VNB
MM1006 N_VGND_M1006_d N_D_M1006_g N_A_27_142#_M1006_s VNB NLOWVT L=0.15 W=0.55
+ AD=0.123281 AS=0.15675 PD=0.98062 PS=1.67 NRD=18 NRS=0 M=1 R=3.66667
+ SA=75000.2 SB=75000.8 A=0.0825 P=1.4 MULT=1
MM1016 N_A_226_104#_M1016_d N_GATE_M1016_g N_VGND_M1006_d VNB NLOWVT L=0.15
+ W=0.74 AD=0.2701 AS=0.165869 PD=2.21 PS=1.31938 NRD=12.972 NRS=8.1 M=1
+ R=4.93333 SA=75000.6 SB=75000.3 A=0.111 P=1.78 MULT=1
MM1007 N_VGND_M1007_d N_A_226_104#_M1007_g N_A_353_98#_M1007_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.207066 AS=0.259 PD=1.59797 PS=2.18 NRD=36.456 NRS=5.664 M=1
+ R=4.93333 SA=75000.3 SB=75001.5 A=0.111 P=1.78 MULT=1
MM1009 A_571_80# N_A_27_142#_M1009_g N_VGND_M1007_d VNB NLOWVT L=0.15 W=0.64
+ AD=0.0672 AS=0.179084 PD=0.85 PS=1.38203 NRD=9.372 NRS=15.936 M=1 R=4.26667
+ SA=75000.8 SB=75001.2 A=0.096 P=1.58 MULT=1
MM1010 N_A_642_392#_M1010_d N_A_353_98#_M1010_g A_571_80# VNB NLOWVT L=0.15
+ W=0.64 AD=0.162536 AS=0.0672 PD=1.38868 PS=0.85 NRD=21.552 NRS=9.372 M=1
+ R=4.26667 SA=75001.1 SB=75000.9 A=0.096 P=1.58 MULT=1
MM1014 A_775_124# N_A_226_104#_M1014_g N_A_642_392#_M1010_d VNB NLOWVT L=0.15
+ W=0.42 AD=0.0504 AS=0.106664 PD=0.66 PS=0.911321 NRD=18.564 NRS=32.856 M=1
+ R=2.8 SA=75001.9 SB=75000.6 A=0.063 P=1.14 MULT=1
MM1008 N_VGND_M1008_d N_A_823_98#_M1008_g A_775_124# VNB NLOWVT L=0.15 W=0.42
+ AD=0.1197 AS=0.0504 PD=1.41 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75002.3
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1021 A_1051_74# N_A_642_392#_M1021_g N_A_823_98#_M1021_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.0888 AS=0.2109 PD=0.98 PS=2.05 NRD=10.536 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75001.1 A=0.111 P=1.78 MULT=1
MM1017 N_VGND_M1017_d N_RESET_B_M1017_g A_1051_74# VNB NLOWVT L=0.15 W=0.74
+ AD=0.1332 AS=0.0888 PD=1.1 PS=0.98 NRD=0 NRS=10.536 M=1 R=4.93333 SA=75000.6
+ SB=75000.7 A=0.111 P=1.78 MULT=1
MM1002 N_Q_M1002_d N_A_823_98#_M1002_g N_VGND_M1017_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.1332 PD=2.05 PS=1.1 NRD=0 NRS=12.972 M=1 R=4.93333 SA=75001.1
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1011 N_VGND_M1011_d N_A_823_98#_M1011_g N_A_1342_74#_M1011_s VNB NLOWVT L=0.15
+ W=0.55 AD=0.105886 AS=0.15675 PD=0.937984 PS=1.67 NRD=18 NRS=0 M=1 R=3.66667
+ SA=75000.2 SB=75000.8 A=0.0825 P=1.4 MULT=1
MM1023 N_Q_N_M1023_d N_A_1342_74#_M1023_g N_VGND_M1011_d VNB NLOWVT L=0.15
+ W=0.74 AD=0.2738 AS=0.142464 PD=2.22 PS=1.26202 NRD=12.972 NRS=0 M=1 R=4.93333
+ SA=75000.6 SB=75000.3 A=0.111 P=1.78 MULT=1
MM1005 N_VPWR_M1005_d N_D_M1005_g N_A_27_142#_M1005_s VPB PSHORT L=0.15 W=0.84
+ AD=0.22785 AS=0.2478 PD=1.52 PS=2.27 NRD=50.7078 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75000.9 A=0.126 P=1.98 MULT=1
MM1003 N_A_226_104#_M1003_d N_GATE_M1003_g N_VPWR_M1005_d VPB PSHORT L=0.15
+ W=0.84 AD=0.3066 AS=0.22785 PD=2.41 PS=1.52 NRD=0 NRS=50.7078 M=1 R=5.6
+ SA=75000.8 SB=75000.3 A=0.126 P=1.98 MULT=1
MM1018 N_VPWR_M1018_d N_A_226_104#_M1018_g N_A_353_98#_M1018_s VPB PSHORT L=0.15
+ W=0.84 AD=0.17147 AS=0.2478 PD=1.26913 PS=2.27 NRD=23.443 NRS=2.3443 M=1 R=5.6
+ SA=75000.2 SB=75002.1 A=0.126 P=1.98 MULT=1
MM1004 A_564_392# N_A_27_142#_M1004_g N_VPWR_M1018_d VPB PSHORT L=0.15 W=1
+ AD=0.12 AS=0.20413 PD=1.24 PS=1.51087 NRD=12.7853 NRS=2.9353 M=1 R=6.66667
+ SA=75000.7 SB=75001.9 A=0.15 P=2.3 MULT=1
MM1019 N_A_642_392#_M1019_d N_A_226_104#_M1019_g A_564_392# VPB PSHORT L=0.15
+ W=1 AD=0.248451 AS=0.12 PD=1.97887 PS=1.24 NRD=3.9203 NRS=12.7853 M=1
+ R=6.66667 SA=75001.1 SB=75001.5 A=0.15 P=2.3 MULT=1
MM1001 A_753_508# N_A_353_98#_M1001_g N_A_642_392#_M1019_d VPB PSHORT L=0.15
+ W=0.42 AD=0.10605 AS=0.104349 PD=0.925 PS=0.831127 NRD=92.6294 NRS=51.5943 M=1
+ R=2.8 SA=75001.5 SB=75002.7 A=0.063 P=1.14 MULT=1
MM1013 N_VPWR_M1013_d N_A_823_98#_M1013_g A_753_508# VPB PSHORT L=0.15 W=0.42
+ AD=0.127336 AS=0.10605 PD=0.976364 PS=0.925 NRD=4.6886 NRS=92.6294 M=1 R=2.8
+ SA=75002.2 SB=75002 A=0.063 P=1.14 MULT=1
MM1015 N_A_823_98#_M1015_d N_A_642_392#_M1015_g N_VPWR_M1013_d VPB PSHORT L=0.15
+ W=1.12 AD=0.182 AS=0.339564 PD=1.445 PS=2.60364 NRD=6.1464 NRS=6.1464 M=1
+ R=7.46667 SA=75001.2 SB=75001.2 A=0.168 P=2.54 MULT=1
MM1022 N_VPWR_M1022_d N_RESET_B_M1022_g N_A_823_98#_M1015_d VPB PSHORT L=0.15
+ W=1.12 AD=0.196 AS=0.182 PD=1.47 PS=1.445 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75001.7 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1020 N_Q_M1020_d N_A_823_98#_M1020_g N_VPWR_M1022_d VPB PSHORT L=0.15 W=1.12
+ AD=0.3304 AS=0.196 PD=2.83 PS=1.47 NRD=1.7533 NRS=10.5395 M=1 R=7.46667
+ SA=75002.2 SB=75000.2 A=0.168 P=2.54 MULT=1
MM1012 N_VPWR_M1012_d N_A_823_98#_M1012_g N_A_1342_74#_M1012_s VPB PSHORT L=0.15
+ W=0.84 AD=0.1596 AS=0.2478 PD=1.26429 PS=2.27 NRD=2.3443 NRS=2.3443 M=1 R=5.6
+ SA=75000.2 SB=75000.7 A=0.126 P=1.98 MULT=1
MM1000 N_Q_N_M1000_d N_A_1342_74#_M1000_g N_VPWR_M1012_d VPB PSHORT L=0.15
+ W=1.12 AD=0.3304 AS=0.2128 PD=2.83 PS=1.68571 NRD=1.7533 NRS=11.426 M=1
+ R=7.46667 SA=75000.6 SB=75000.2 A=0.168 P=2.54 MULT=1
DX24_noxref VNB VPB NWDIODE A=15.8844 P=20.8
c_88 VNB 0 6.46507e-20 $X=0 $Y=0
*
.include "sky130_fd_sc_hs__dlrbp_1.pxi.spice"
*
.ends
*
*
