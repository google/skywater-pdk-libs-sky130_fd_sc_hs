* File: sky130_fd_sc_hs__dlrtp_4.pxi.spice
* Created: Thu Aug 27 20:42:03 2020
* 
x_PM_SKY130_FD_SC_HS__DLRTP_4%D N_D_M1019_g N_D_c_179_n N_D_M1009_g D
+ N_D_c_180_n PM_SKY130_FD_SC_HS__DLRTP_4%D
x_PM_SKY130_FD_SC_HS__DLRTP_4%GATE N_GATE_c_204_n N_GATE_M1007_g N_GATE_M1004_g
+ GATE PM_SKY130_FD_SC_HS__DLRTP_4%GATE
x_PM_SKY130_FD_SC_HS__DLRTP_4%A_240_394# N_A_240_394#_M1004_d
+ N_A_240_394#_M1007_d N_A_240_394#_c_251_n N_A_240_394#_M1016_g
+ N_A_240_394#_c_237_n N_A_240_394#_M1024_g N_A_240_394#_c_252_n
+ N_A_240_394#_M1008_g N_A_240_394#_c_253_n N_A_240_394#_c_254_n
+ N_A_240_394#_M1002_g N_A_240_394#_c_239_n N_A_240_394#_c_240_n
+ N_A_240_394#_c_257_n N_A_240_394#_c_241_n N_A_240_394#_c_242_n
+ N_A_240_394#_c_243_n N_A_240_394#_c_382_p N_A_240_394#_c_244_n
+ N_A_240_394#_c_245_n N_A_240_394#_c_246_n N_A_240_394#_c_247_n
+ N_A_240_394#_c_248_n N_A_240_394#_c_249_n N_A_240_394#_c_250_n
+ PM_SKY130_FD_SC_HS__DLRTP_4%A_240_394#
x_PM_SKY130_FD_SC_HS__DLRTP_4%A_27_126# N_A_27_126#_M1019_s N_A_27_126#_M1009_s
+ N_A_27_126#_M1001_g N_A_27_126#_c_387_n N_A_27_126#_M1018_g
+ N_A_27_126#_c_388_n N_A_27_126#_c_389_n N_A_27_126#_c_390_n
+ N_A_27_126#_c_391_n N_A_27_126#_c_395_n N_A_27_126#_c_396_n
+ N_A_27_126#_c_397_n N_A_27_126#_c_392_n PM_SKY130_FD_SC_HS__DLRTP_4%A_27_126#
x_PM_SKY130_FD_SC_HS__DLRTP_4%A_364_120# N_A_364_120#_M1024_s
+ N_A_364_120#_M1016_s N_A_364_120#_M1027_g N_A_364_120#_c_481_n
+ N_A_364_120#_M1005_g N_A_364_120#_c_475_n N_A_364_120#_c_476_n
+ N_A_364_120#_c_477_n N_A_364_120#_c_572_p N_A_364_120#_c_478_n
+ N_A_364_120#_c_484_n N_A_364_120#_c_485_n N_A_364_120#_c_486_n
+ N_A_364_120#_c_487_n N_A_364_120#_c_518_n N_A_364_120#_c_479_n
+ N_A_364_120#_c_480_n PM_SKY130_FD_SC_HS__DLRTP_4%A_364_120#
x_PM_SKY130_FD_SC_HS__DLRTP_4%A_797_48# N_A_797_48#_M1000_s N_A_797_48#_M1017_d
+ N_A_797_48#_M1021_d N_A_797_48#_c_581_n N_A_797_48#_M1026_g
+ N_A_797_48#_c_582_n N_A_797_48#_c_583_n N_A_797_48#_c_597_n
+ N_A_797_48#_M1003_g N_A_797_48#_c_584_n N_A_797_48#_c_599_n
+ N_A_797_48#_M1010_g N_A_797_48#_M1011_g N_A_797_48#_c_600_n
+ N_A_797_48#_M1012_g N_A_797_48#_M1015_g N_A_797_48#_c_601_n
+ N_A_797_48#_M1013_g N_A_797_48#_M1023_g N_A_797_48#_c_602_n
+ N_A_797_48#_M1014_g N_A_797_48#_M1029_g N_A_797_48#_c_603_n
+ N_A_797_48#_c_589_n N_A_797_48#_c_604_n N_A_797_48#_c_590_n
+ N_A_797_48#_c_606_n N_A_797_48#_c_591_n N_A_797_48#_c_769_p
+ N_A_797_48#_c_592_n N_A_797_48#_c_593_n N_A_797_48#_c_594_n
+ N_A_797_48#_c_595_n N_A_797_48#_c_596_n PM_SKY130_FD_SC_HS__DLRTP_4%A_797_48#
x_PM_SKY130_FD_SC_HS__DLRTP_4%A_640_74# N_A_640_74#_M1027_d N_A_640_74#_M1008_d
+ N_A_640_74#_M1000_g N_A_640_74#_c_774_n N_A_640_74#_M1017_g
+ N_A_640_74#_c_775_n N_A_640_74#_M1006_g N_A_640_74#_c_777_n
+ N_A_640_74#_c_783_n N_A_640_74#_M1025_g N_A_640_74#_c_778_n
+ N_A_640_74#_c_790_n N_A_640_74#_c_779_n N_A_640_74#_c_785_n
+ N_A_640_74#_c_786_n N_A_640_74#_c_780_n N_A_640_74#_c_803_n
+ N_A_640_74#_c_788_n PM_SKY130_FD_SC_HS__DLRTP_4%A_640_74#
x_PM_SKY130_FD_SC_HS__DLRTP_4%RESET_B N_RESET_B_c_883_n N_RESET_B_M1020_g
+ N_RESET_B_c_884_n N_RESET_B_c_890_n N_RESET_B_M1021_g N_RESET_B_c_885_n
+ N_RESET_B_M1028_g N_RESET_B_c_886_n N_RESET_B_c_892_n N_RESET_B_M1022_g
+ RESET_B RESET_B N_RESET_B_c_888_n PM_SKY130_FD_SC_HS__DLRTP_4%RESET_B
x_PM_SKY130_FD_SC_HS__DLRTP_4%VPWR N_VPWR_M1009_d N_VPWR_M1016_d N_VPWR_M1003_d
+ N_VPWR_M1025_s N_VPWR_M1022_s N_VPWR_M1012_s N_VPWR_M1014_s N_VPWR_c_948_n
+ N_VPWR_c_949_n N_VPWR_c_950_n N_VPWR_c_951_n N_VPWR_c_952_n N_VPWR_c_953_n
+ N_VPWR_c_954_n N_VPWR_c_955_n N_VPWR_c_956_n N_VPWR_c_957_n N_VPWR_c_958_n
+ N_VPWR_c_959_n N_VPWR_c_960_n N_VPWR_c_961_n VPWR N_VPWR_c_962_n
+ N_VPWR_c_963_n N_VPWR_c_964_n N_VPWR_c_965_n N_VPWR_c_966_n N_VPWR_c_967_n
+ N_VPWR_c_947_n PM_SKY130_FD_SC_HS__DLRTP_4%VPWR
x_PM_SKY130_FD_SC_HS__DLRTP_4%Q N_Q_M1011_d N_Q_M1023_d N_Q_M1010_d N_Q_M1013_d
+ N_Q_c_1072_n N_Q_c_1065_n N_Q_c_1066_n N_Q_c_1073_n N_Q_c_1074_n N_Q_c_1067_n
+ N_Q_c_1075_n N_Q_c_1068_n N_Q_c_1076_n N_Q_c_1069_n N_Q_c_1077_n N_Q_c_1070_n
+ Q Q PM_SKY130_FD_SC_HS__DLRTP_4%Q
x_PM_SKY130_FD_SC_HS__DLRTP_4%VGND N_VGND_M1019_d N_VGND_M1024_d N_VGND_M1026_d
+ N_VGND_M1020_d N_VGND_M1011_s N_VGND_M1015_s N_VGND_M1029_s N_VGND_c_1142_n
+ N_VGND_c_1143_n N_VGND_c_1144_n N_VGND_c_1145_n N_VGND_c_1146_n
+ N_VGND_c_1147_n N_VGND_c_1148_n N_VGND_c_1149_n N_VGND_c_1150_n
+ N_VGND_c_1151_n N_VGND_c_1152_n VGND N_VGND_c_1153_n N_VGND_c_1154_n
+ N_VGND_c_1155_n N_VGND_c_1156_n N_VGND_c_1157_n N_VGND_c_1158_n
+ N_VGND_c_1159_n N_VGND_c_1160_n N_VGND_c_1161_n N_VGND_c_1162_n
+ PM_SKY130_FD_SC_HS__DLRTP_4%VGND
x_PM_SKY130_FD_SC_HS__DLRTP_4%A_938_74# N_A_938_74#_M1000_d N_A_938_74#_M1006_d
+ N_A_938_74#_M1028_s N_A_938_74#_c_1269_n N_A_938_74#_c_1270_n
+ N_A_938_74#_c_1271_n N_A_938_74#_c_1280_n N_A_938_74#_c_1291_n
+ N_A_938_74#_c_1281_n N_A_938_74#_c_1272_n N_A_938_74#_c_1273_n
+ PM_SKY130_FD_SC_HS__DLRTP_4%A_938_74#
cc_1 VNB N_D_M1019_g 0.0375298f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.905
cc_2 VNB N_D_c_179_n 0.0247413f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.895
cc_3 VNB N_D_c_180_n 0.00883608f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.615
cc_4 VNB N_GATE_c_204_n 0.0213973f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.45
cc_5 VNB N_GATE_M1004_g 0.0323638f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.39
cc_6 VNB GATE 0.00357568f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_7 VNB N_A_240_394#_c_237_n 0.0203645f $X=-0.19 $Y=-0.245 $X2=0.407 $Y2=1.615
cc_8 VNB N_A_240_394#_M1002_g 0.0345097f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A_240_394#_c_239_n 0.0365985f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_240_394#_c_240_n 0.0129513f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_240_394#_c_241_n 0.00543282f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_240_394#_c_242_n 2.56964e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_240_394#_c_243_n 0.00636489f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_240_394#_c_244_n 0.00512304f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_240_394#_c_245_n 0.00202103f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_240_394#_c_246_n 0.0215614f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_240_394#_c_247_n 0.00182119f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_240_394#_c_248_n 0.00387937f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_240_394#_c_249_n 0.0562046f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_240_394#_c_250_n 0.00482344f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_27_126#_M1001_g 0.0367238f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_27_126#_c_387_n 0.0277721f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.615
cc_23 VNB N_A_27_126#_c_388_n 0.0229205f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.615
cc_24 VNB N_A_27_126#_c_389_n 0.00295866f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_27_126#_c_390_n 0.00965227f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_27_126#_c_391_n 0.00747638f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_27_126#_c_392_n 0.00145416f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_364_120#_c_475_n 0.00149766f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_364_120#_c_476_n 0.0163195f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_364_120#_c_477_n 0.00167324f $X=-0.19 $Y=-0.245 $X2=0.385
+ $Y2=1.615
cc_31 VNB N_A_364_120#_c_478_n 0.00331517f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_364_120#_c_479_n 0.0305134f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_364_120#_c_480_n 0.0174433f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_797_48#_c_581_n 0.0152835f $X=-0.19 $Y=-0.245 $X2=0.407 $Y2=1.615
cc_35 VNB N_A_797_48#_c_582_n 0.0304119f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.615
cc_36 VNB N_A_797_48#_c_583_n 0.00620855f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_797_48#_c_584_n 0.037999f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_797_48#_M1011_g 0.0240095f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_797_48#_M1015_g 0.020319f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_797_48#_M1023_g 0.0202914f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_797_48#_M1029_g 0.0232598f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_797_48#_c_589_n 0.00875582f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_797_48#_c_590_n 0.00496676f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_797_48#_c_591_n 0.00212473f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_A_797_48#_c_592_n 0.00227286f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_A_797_48#_c_593_n 0.00236205f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_797_48#_c_594_n 0.00356754f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_797_48#_c_595_n 0.00981913f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A_797_48#_c_596_n 0.12584f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_A_640_74#_M1000_g 0.0325439f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_A_640_74#_c_774_n 0.029019f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.615
cc_52 VNB N_A_640_74#_c_775_n 0.00984954f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_A_640_74#_M1006_g 0.0208553f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_A_640_74#_c_777_n 0.00861992f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_A_640_74#_c_778_n 0.0147763f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_A_640_74#_c_779_n 0.00534236f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_A_640_74#_c_780_n 0.00304287f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_RESET_B_c_883_n 0.0168755f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.45
cc_59 VNB N_RESET_B_c_884_n 0.0118789f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.895
cc_60 VNB N_RESET_B_c_885_n 0.0191027f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_RESET_B_c_886_n 0.012091f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.615
cc_62 VNB RESET_B 0.0041731f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_RESET_B_c_888_n 0.0516666f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_VPWR_c_947_n 0.382608f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_Q_c_1065_n 0.0018817f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_Q_c_1066_n 0.00205904f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_Q_c_1067_n 0.00308327f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_Q_c_1068_n 0.00168586f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_Q_c_1069_n 0.0118257f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_Q_c_1070_n 0.00145912f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB Q 0.0262974f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_VGND_c_1142_n 0.0193117f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_VGND_c_1143_n 0.0152056f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_VGND_c_1144_n 0.0153789f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_VGND_c_1145_n 0.00340259f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_VGND_c_1146_n 0.0187456f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_VGND_c_1147_n 0.0172414f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_VGND_c_1148_n 0.002601f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VNB N_VGND_c_1149_n 0.0120272f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_VGND_c_1150_n 0.022631f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_81 VNB N_VGND_c_1151_n 0.0367891f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_82 VNB N_VGND_c_1152_n 0.00480499f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_83 VNB N_VGND_c_1153_n 0.0394586f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_84 VNB N_VGND_c_1154_n 0.0383268f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_85 VNB N_VGND_c_1155_n 0.0169145f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_86 VNB N_VGND_c_1156_n 0.0150599f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_87 VNB N_VGND_c_1157_n 0.0285952f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_88 VNB N_VGND_c_1158_n 0.00613689f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_89 VNB N_VGND_c_1159_n 0.00601668f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_90 VNB N_VGND_c_1160_n 0.00500104f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_91 VNB N_VGND_c_1161_n 0.00604233f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_92 VNB N_VGND_c_1162_n 0.50317f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_93 VNB N_A_938_74#_c_1269_n 0.00985803f $X=-0.19 $Y=-0.245 $X2=0.385
+ $Y2=1.615
cc_94 VNB N_A_938_74#_c_1270_n 0.00451548f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_95 VNB N_A_938_74#_c_1271_n 0.00419496f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_96 VNB N_A_938_74#_c_1272_n 0.00193746f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_97 VNB N_A_938_74#_c_1273_n 0.00627934f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_98 VPB N_D_c_179_n 0.0481409f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.895
cc_99 VPB N_D_c_180_n 0.00541046f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.615
cc_100 VPB N_GATE_c_204_n 0.0423845f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.45
cc_101 VPB GATE 8.30128e-19 $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_102 VPB N_A_240_394#_c_251_n 0.0204044f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.39
cc_103 VPB N_A_240_394#_c_252_n 0.0145896f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=1.615
cc_104 VPB N_A_240_394#_c_253_n 0.0299379f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.615
cc_105 VPB N_A_240_394#_c_254_n 0.010221f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_106 VPB N_A_240_394#_c_239_n 0.0148942f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_107 VPB N_A_240_394#_c_240_n 0.00813043f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_108 VPB N_A_240_394#_c_257_n 0.00909847f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_109 VPB N_A_240_394#_c_242_n 0.00368783f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_110 VPB N_A_240_394#_c_247_n 7.67686e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_111 VPB N_A_240_394#_c_249_n 0.00968701f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_112 VPB N_A_27_126#_c_387_n 0.0278773f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.615
cc_113 VPB N_A_27_126#_c_391_n 0.00577071f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_114 VPB N_A_27_126#_c_395_n 0.00894256f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_115 VPB N_A_27_126#_c_396_n 0.00111793f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_116 VPB N_A_27_126#_c_397_n 0.0431134f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_117 VPB N_A_364_120#_c_481_n 0.065333f $X=-0.19 $Y=1.66 $X2=0.407 $Y2=1.615
cc_118 VPB N_A_364_120#_c_475_n 0.00243696f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_119 VPB N_A_364_120#_c_478_n 0.00224784f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_120 VPB N_A_364_120#_c_484_n 0.00615053f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_121 VPB N_A_364_120#_c_485_n 0.00202743f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_122 VPB N_A_364_120#_c_486_n 0.00131657f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_123 VPB N_A_364_120#_c_487_n 0.00180638f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_124 VPB N_A_797_48#_c_597_n 0.0552879f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_125 VPB N_A_797_48#_c_584_n 0.0280057f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_126 VPB N_A_797_48#_c_599_n 0.0172689f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_127 VPB N_A_797_48#_c_600_n 0.0156157f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_128 VPB N_A_797_48#_c_601_n 0.0156499f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_129 VPB N_A_797_48#_c_602_n 0.0170534f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_130 VPB N_A_797_48#_c_603_n 0.0119988f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_131 VPB N_A_797_48#_c_604_n 3.39932e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_132 VPB N_A_797_48#_c_590_n 0.00528369f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_133 VPB N_A_797_48#_c_606_n 0.00474574f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_134 VPB N_A_797_48#_c_592_n 8.84457e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_135 VPB N_A_797_48#_c_594_n 0.003521f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_136 VPB N_A_797_48#_c_595_n 0.00296695f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_137 VPB N_A_797_48#_c_596_n 0.0277913f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_138 VPB N_A_640_74#_c_774_n 0.0305205f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.615
cc_139 VPB N_A_640_74#_c_777_n 6.56313e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_140 VPB N_A_640_74#_c_783_n 0.0205584f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_141 VPB N_A_640_74#_c_779_n 3.14364e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_142 VPB N_A_640_74#_c_785_n 0.0300083f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_143 VPB N_A_640_74#_c_786_n 0.00540289f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_144 VPB N_A_640_74#_c_780_n 4.66164e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_145 VPB N_A_640_74#_c_788_n 0.00292687f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_146 VPB N_RESET_B_c_884_n 6.84519e-19 $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.895
cc_147 VPB N_RESET_B_c_890_n 0.0206524f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.39
cc_148 VPB N_RESET_B_c_886_n 7.01837e-19 $X=-0.19 $Y=1.66 $X2=0.24 $Y2=1.615
cc_149 VPB N_RESET_B_c_892_n 0.0214833f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_150 VPB N_VPWR_c_948_n 0.0204129f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_151 VPB N_VPWR_c_949_n 0.0127171f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_152 VPB N_VPWR_c_950_n 0.0202868f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_153 VPB N_VPWR_c_951_n 0.0303394f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_154 VPB N_VPWR_c_952_n 0.016486f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_155 VPB N_VPWR_c_953_n 0.00517393f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_156 VPB N_VPWR_c_954_n 0.0147428f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_157 VPB N_VPWR_c_955_n 0.0439511f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_158 VPB N_VPWR_c_956_n 0.0208961f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_159 VPB N_VPWR_c_957_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_160 VPB N_VPWR_c_958_n 0.0208961f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_161 VPB N_VPWR_c_959_n 0.00614127f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_162 VPB N_VPWR_c_960_n 0.0175706f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_163 VPB N_VPWR_c_961_n 0.00614127f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_164 VPB N_VPWR_c_962_n 0.0430552f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_165 VPB N_VPWR_c_963_n 0.0420502f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_166 VPB N_VPWR_c_964_n 0.0185368f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_167 VPB N_VPWR_c_965_n 0.027231f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_168 VPB N_VPWR_c_966_n 0.00615173f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_169 VPB N_VPWR_c_967_n 0.0105653f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_170 VPB N_VPWR_c_947_n 0.123582f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_171 VPB N_Q_c_1072_n 0.00216998f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_172 VPB N_Q_c_1073_n 0.00229638f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_173 VPB N_Q_c_1074_n 0.00193406f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_174 VPB N_Q_c_1075_n 0.00326964f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_175 VPB N_Q_c_1076_n 0.0128296f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_176 VPB N_Q_c_1077_n 0.0020352f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_177 VPB Q 0.00747008f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_178 N_D_c_179_n N_GATE_c_204_n 0.0306386f $X=0.505 $Y=1.895 $X2=-0.19
+ $Y2=-0.245
cc_179 N_D_M1019_g N_GATE_M1004_g 0.013513f $X=0.495 $Y=0.905 $X2=0 $Y2=0
cc_180 N_D_M1019_g N_A_240_394#_c_246_n 8.79535e-19 $X=0.495 $Y=0.905 $X2=0
+ $Y2=0
cc_181 N_D_M1019_g N_A_27_126#_c_388_n 0.0103282f $X=0.495 $Y=0.905 $X2=0 $Y2=0
cc_182 N_D_M1019_g N_A_27_126#_c_389_n 0.0122469f $X=0.495 $Y=0.905 $X2=0 $Y2=0
cc_183 N_D_c_179_n N_A_27_126#_c_389_n 7.44236e-19 $X=0.505 $Y=1.895 $X2=0 $Y2=0
cc_184 N_D_c_180_n N_A_27_126#_c_389_n 0.00496499f $X=0.385 $Y=1.615 $X2=0 $Y2=0
cc_185 N_D_M1019_g N_A_27_126#_c_390_n 0.00418246f $X=0.495 $Y=0.905 $X2=0 $Y2=0
cc_186 N_D_c_179_n N_A_27_126#_c_390_n 0.00465635f $X=0.505 $Y=1.895 $X2=0 $Y2=0
cc_187 N_D_c_180_n N_A_27_126#_c_390_n 0.0272332f $X=0.385 $Y=1.615 $X2=0 $Y2=0
cc_188 N_D_M1019_g N_A_27_126#_c_391_n 0.00421485f $X=0.495 $Y=0.905 $X2=0 $Y2=0
cc_189 N_D_c_179_n N_A_27_126#_c_391_n 0.00726158f $X=0.505 $Y=1.895 $X2=0 $Y2=0
cc_190 N_D_c_180_n N_A_27_126#_c_391_n 0.0250891f $X=0.385 $Y=1.615 $X2=0 $Y2=0
cc_191 N_D_c_179_n N_A_27_126#_c_397_n 0.0377902f $X=0.505 $Y=1.895 $X2=0 $Y2=0
cc_192 N_D_c_180_n N_A_27_126#_c_397_n 0.0328357f $X=0.385 $Y=1.615 $X2=0 $Y2=0
cc_193 N_D_c_179_n N_VPWR_c_948_n 0.0043785f $X=0.505 $Y=1.895 $X2=0 $Y2=0
cc_194 N_D_c_179_n N_VPWR_c_965_n 0.00463088f $X=0.505 $Y=1.895 $X2=0 $Y2=0
cc_195 N_D_c_179_n N_VPWR_c_947_n 0.00499434f $X=0.505 $Y=1.895 $X2=0 $Y2=0
cc_196 N_D_M1019_g N_VGND_c_1142_n 0.00655179f $X=0.495 $Y=0.905 $X2=0 $Y2=0
cc_197 N_D_M1019_g N_VGND_c_1157_n 0.00397467f $X=0.495 $Y=0.905 $X2=0 $Y2=0
cc_198 N_D_M1019_g N_VGND_c_1162_n 0.00468052f $X=0.495 $Y=0.905 $X2=0 $Y2=0
cc_199 N_GATE_c_204_n N_A_240_394#_c_239_n 0.0173832f $X=1.125 $Y=1.895 $X2=0
+ $Y2=0
cc_200 GATE N_A_240_394#_c_239_n 3.1363e-19 $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_201 N_GATE_c_204_n N_A_240_394#_c_257_n 0.00674487f $X=1.125 $Y=1.895 $X2=0
+ $Y2=0
cc_202 GATE N_A_240_394#_c_257_n 0.00803258f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_203 N_GATE_M1004_g N_A_240_394#_c_241_n 0.00566034f $X=1.19 $Y=0.81 $X2=0
+ $Y2=0
cc_204 N_GATE_c_204_n N_A_240_394#_c_242_n 0.00366002f $X=1.125 $Y=1.895 $X2=0
+ $Y2=0
cc_205 N_GATE_c_204_n N_A_240_394#_c_246_n 0.00185341f $X=1.125 $Y=1.895 $X2=0
+ $Y2=0
cc_206 N_GATE_M1004_g N_A_240_394#_c_246_n 0.0142314f $X=1.19 $Y=0.81 $X2=0
+ $Y2=0
cc_207 GATE N_A_240_394#_c_246_n 0.00293385f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_208 N_GATE_c_204_n N_A_240_394#_c_247_n 0.00220635f $X=1.125 $Y=1.895 $X2=0
+ $Y2=0
cc_209 GATE N_A_240_394#_c_247_n 0.026282f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_210 N_GATE_M1004_g N_A_27_126#_c_388_n 7.88473e-19 $X=1.19 $Y=0.81 $X2=0
+ $Y2=0
cc_211 N_GATE_M1004_g N_A_27_126#_c_389_n 0.00195644f $X=1.19 $Y=0.81 $X2=0
+ $Y2=0
cc_212 N_GATE_c_204_n N_A_27_126#_c_391_n 0.00460466f $X=1.125 $Y=1.895 $X2=0
+ $Y2=0
cc_213 N_GATE_M1004_g N_A_27_126#_c_391_n 0.00178944f $X=1.19 $Y=0.81 $X2=0
+ $Y2=0
cc_214 GATE N_A_27_126#_c_391_n 0.0243916f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_215 N_GATE_c_204_n N_A_27_126#_c_395_n 0.0163239f $X=1.125 $Y=1.895 $X2=0
+ $Y2=0
cc_216 GATE N_A_27_126#_c_395_n 0.00378022f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_217 N_GATE_c_204_n N_A_27_126#_c_397_n 0.00822393f $X=1.125 $Y=1.895 $X2=0
+ $Y2=0
cc_218 N_GATE_c_204_n N_VPWR_c_948_n 0.00663705f $X=1.125 $Y=1.895 $X2=0 $Y2=0
cc_219 N_GATE_c_204_n N_VPWR_c_962_n 0.00475172f $X=1.125 $Y=1.895 $X2=0 $Y2=0
cc_220 N_GATE_c_204_n N_VPWR_c_947_n 0.00499434f $X=1.125 $Y=1.895 $X2=0 $Y2=0
cc_221 N_GATE_c_204_n N_VGND_c_1142_n 2.80107e-19 $X=1.125 $Y=1.895 $X2=0 $Y2=0
cc_222 N_GATE_M1004_g N_VGND_c_1142_n 0.0107555f $X=1.19 $Y=0.81 $X2=0 $Y2=0
cc_223 N_GATE_M1004_g N_VGND_c_1153_n 0.00504315f $X=1.19 $Y=0.81 $X2=0 $Y2=0
cc_224 N_GATE_M1004_g N_VGND_c_1162_n 0.00523671f $X=1.19 $Y=0.81 $X2=0 $Y2=0
cc_225 N_A_240_394#_c_237_n N_A_27_126#_M1001_g 0.0287084f $X=2.205 $Y=1.45
+ $X2=0 $Y2=0
cc_226 N_A_240_394#_c_243_n N_A_27_126#_M1001_g 0.0112826f $X=2.835 $Y=0.855
+ $X2=0 $Y2=0
cc_227 N_A_240_394#_c_245_n N_A_27_126#_M1001_g 0.00113528f $X=3.005 $Y=0.34
+ $X2=0 $Y2=0
cc_228 N_A_240_394#_c_251_n N_A_27_126#_c_387_n 0.0230391f $X=2.19 $Y=1.885
+ $X2=0 $Y2=0
cc_229 N_A_240_394#_c_252_n N_A_27_126#_c_387_n 0.0547507f $X=3.125 $Y=1.885
+ $X2=0 $Y2=0
cc_230 N_A_240_394#_c_254_n N_A_27_126#_c_387_n 0.0119319f $X=3.215 $Y=1.765
+ $X2=0 $Y2=0
cc_231 N_A_240_394#_c_240_n N_A_27_126#_c_387_n 0.0232067f $X=2.19 $Y=1.667
+ $X2=0 $Y2=0
cc_232 N_A_240_394#_c_241_n N_A_27_126#_c_389_n 0.00274328f $X=1.545 $Y=1.45
+ $X2=0 $Y2=0
cc_233 N_A_240_394#_c_246_n N_A_27_126#_c_389_n 0.00404324f $X=1.405 $Y=0.585
+ $X2=0 $Y2=0
cc_234 N_A_240_394#_c_241_n N_A_27_126#_c_391_n 0.00522563f $X=1.545 $Y=1.45
+ $X2=0 $Y2=0
cc_235 N_A_240_394#_c_242_n N_A_27_126#_c_391_n 0.00520786f $X=1.545 $Y=1.95
+ $X2=0 $Y2=0
cc_236 N_A_240_394#_M1007_d N_A_27_126#_c_395_n 0.0102693f $X=1.2 $Y=1.97 $X2=0
+ $Y2=0
cc_237 N_A_240_394#_c_251_n N_A_27_126#_c_395_n 0.0149669f $X=2.19 $Y=1.885
+ $X2=0 $Y2=0
cc_238 N_A_240_394#_c_239_n N_A_27_126#_c_395_n 0.00321241f $X=2.1 $Y=1.615
+ $X2=0 $Y2=0
cc_239 N_A_240_394#_c_257_n N_A_27_126#_c_395_n 0.0297023f $X=1.46 $Y=2.075
+ $X2=0 $Y2=0
cc_240 N_A_240_394#_c_247_n N_A_27_126#_c_395_n 0.00500743f $X=1.735 $Y=1.615
+ $X2=0 $Y2=0
cc_241 N_A_240_394#_c_251_n N_A_27_126#_c_396_n 0.00561239f $X=2.19 $Y=1.885
+ $X2=0 $Y2=0
cc_242 N_A_240_394#_c_252_n N_A_27_126#_c_396_n 2.76464e-19 $X=3.125 $Y=1.885
+ $X2=0 $Y2=0
cc_243 N_A_240_394#_c_240_n N_A_27_126#_c_396_n 5.87186e-19 $X=2.19 $Y=1.667
+ $X2=0 $Y2=0
cc_244 N_A_240_394#_c_257_n N_A_27_126#_c_397_n 0.012627f $X=1.46 $Y=2.075 $X2=0
+ $Y2=0
cc_245 N_A_240_394#_c_240_n N_A_27_126#_c_392_n 0.00136035f $X=2.19 $Y=1.667
+ $X2=0 $Y2=0
cc_246 N_A_240_394#_c_243_n N_A_364_120#_M1024_s 0.00837187f $X=2.835 $Y=0.855
+ $X2=-0.19 $Y2=-0.245
cc_247 N_A_240_394#_c_252_n N_A_364_120#_c_481_n 0.0221802f $X=3.125 $Y=1.885
+ $X2=0 $Y2=0
cc_248 N_A_240_394#_c_253_n N_A_364_120#_c_481_n 0.0133755f $X=3.625 $Y=1.765
+ $X2=0 $Y2=0
cc_249 N_A_240_394#_c_249_n N_A_364_120#_c_481_n 0.00376644f $X=3.985 $Y=1.39
+ $X2=0 $Y2=0
cc_250 N_A_240_394#_c_251_n N_A_364_120#_c_475_n 0.00400504f $X=2.19 $Y=1.885
+ $X2=0 $Y2=0
cc_251 N_A_240_394#_c_237_n N_A_364_120#_c_475_n 0.00616191f $X=2.205 $Y=1.45
+ $X2=0 $Y2=0
cc_252 N_A_240_394#_c_239_n N_A_364_120#_c_475_n 0.00637978f $X=2.1 $Y=1.615
+ $X2=0 $Y2=0
cc_253 N_A_240_394#_c_240_n N_A_364_120#_c_475_n 0.0113743f $X=2.19 $Y=1.667
+ $X2=0 $Y2=0
cc_254 N_A_240_394#_c_257_n N_A_364_120#_c_475_n 0.00176069f $X=1.46 $Y=2.075
+ $X2=0 $Y2=0
cc_255 N_A_240_394#_c_241_n N_A_364_120#_c_475_n 0.00654383f $X=1.545 $Y=1.45
+ $X2=0 $Y2=0
cc_256 N_A_240_394#_c_242_n N_A_364_120#_c_475_n 0.00661438f $X=1.545 $Y=1.95
+ $X2=0 $Y2=0
cc_257 N_A_240_394#_c_247_n N_A_364_120#_c_475_n 0.0240999f $X=1.735 $Y=1.615
+ $X2=0 $Y2=0
cc_258 N_A_240_394#_c_237_n N_A_364_120#_c_476_n 0.00526154f $X=2.205 $Y=1.45
+ $X2=0 $Y2=0
cc_259 N_A_240_394#_c_254_n N_A_364_120#_c_476_n 0.00132929f $X=3.215 $Y=1.765
+ $X2=0 $Y2=0
cc_260 N_A_240_394#_M1002_g N_A_364_120#_c_476_n 3.56739e-19 $X=3.7 $Y=0.58
+ $X2=0 $Y2=0
cc_261 N_A_240_394#_c_243_n N_A_364_120#_c_476_n 0.0131302f $X=2.835 $Y=0.855
+ $X2=0 $Y2=0
cc_262 N_A_240_394#_c_237_n N_A_364_120#_c_477_n 0.00355682f $X=2.205 $Y=1.45
+ $X2=0 $Y2=0
cc_263 N_A_240_394#_c_239_n N_A_364_120#_c_477_n 0.00894632f $X=2.1 $Y=1.615
+ $X2=0 $Y2=0
cc_264 N_A_240_394#_c_243_n N_A_364_120#_c_477_n 0.062109f $X=2.835 $Y=0.855
+ $X2=0 $Y2=0
cc_265 N_A_240_394#_c_246_n N_A_364_120#_c_477_n 0.0146026f $X=1.405 $Y=0.585
+ $X2=0 $Y2=0
cc_266 N_A_240_394#_c_247_n N_A_364_120#_c_477_n 0.00741013f $X=1.735 $Y=1.615
+ $X2=0 $Y2=0
cc_267 N_A_240_394#_c_252_n N_A_364_120#_c_478_n 0.00182659f $X=3.125 $Y=1.885
+ $X2=0 $Y2=0
cc_268 N_A_240_394#_c_254_n N_A_364_120#_c_478_n 0.00617016f $X=3.215 $Y=1.765
+ $X2=0 $Y2=0
cc_269 N_A_240_394#_c_249_n N_A_364_120#_c_478_n 0.00115307f $X=3.985 $Y=1.39
+ $X2=0 $Y2=0
cc_270 N_A_240_394#_c_252_n N_A_364_120#_c_484_n 0.0131227f $X=3.125 $Y=1.885
+ $X2=0 $Y2=0
cc_271 N_A_240_394#_c_252_n N_A_364_120#_c_486_n 5.05727e-19 $X=3.125 $Y=1.885
+ $X2=0 $Y2=0
cc_272 N_A_240_394#_c_251_n N_A_364_120#_c_487_n 0.00542873f $X=2.19 $Y=1.885
+ $X2=0 $Y2=0
cc_273 N_A_240_394#_c_239_n N_A_364_120#_c_487_n 0.00792532f $X=2.1 $Y=1.615
+ $X2=0 $Y2=0
cc_274 N_A_240_394#_c_257_n N_A_364_120#_c_487_n 0.0156346f $X=1.46 $Y=2.075
+ $X2=0 $Y2=0
cc_275 N_A_240_394#_c_247_n N_A_364_120#_c_487_n 0.00571739f $X=1.735 $Y=1.615
+ $X2=0 $Y2=0
cc_276 N_A_240_394#_c_252_n N_A_364_120#_c_518_n 0.00713047f $X=3.125 $Y=1.885
+ $X2=0 $Y2=0
cc_277 N_A_240_394#_c_254_n N_A_364_120#_c_479_n 0.0177015f $X=3.215 $Y=1.765
+ $X2=0 $Y2=0
cc_278 N_A_240_394#_M1002_g N_A_364_120#_c_479_n 0.0155829f $X=3.7 $Y=0.58 $X2=0
+ $Y2=0
cc_279 N_A_240_394#_M1002_g N_A_364_120#_c_480_n 0.0171818f $X=3.7 $Y=0.58 $X2=0
+ $Y2=0
cc_280 N_A_240_394#_c_244_n N_A_364_120#_c_480_n 0.0130565f $X=3.85 $Y=0.34
+ $X2=0 $Y2=0
cc_281 N_A_240_394#_M1002_g N_A_797_48#_c_581_n 0.0463045f $X=3.7 $Y=0.58 $X2=0
+ $Y2=0
cc_282 N_A_240_394#_c_244_n N_A_797_48#_c_581_n 0.00364564f $X=3.85 $Y=0.34
+ $X2=0 $Y2=0
cc_283 N_A_240_394#_c_250_n N_A_797_48#_c_581_n 0.00792101f $X=4 $Y=1.225 $X2=0
+ $Y2=0
cc_284 N_A_240_394#_c_248_n N_A_797_48#_c_583_n 9.77689e-19 $X=3.985 $Y=1.39
+ $X2=0 $Y2=0
cc_285 N_A_240_394#_c_249_n N_A_797_48#_c_583_n 0.0108375f $X=3.985 $Y=1.39
+ $X2=0 $Y2=0
cc_286 N_A_240_394#_c_250_n N_A_797_48#_c_583_n 0.00540005f $X=4 $Y=1.225 $X2=0
+ $Y2=0
cc_287 N_A_240_394#_M1002_g N_A_797_48#_c_584_n 0.00252594f $X=3.7 $Y=0.58 $X2=0
+ $Y2=0
cc_288 N_A_240_394#_c_248_n N_A_797_48#_c_584_n 0.00163189f $X=3.985 $Y=1.39
+ $X2=0 $Y2=0
cc_289 N_A_240_394#_c_249_n N_A_797_48#_c_584_n 0.0268484f $X=3.985 $Y=1.39
+ $X2=0 $Y2=0
cc_290 N_A_240_394#_c_250_n N_A_797_48#_c_584_n 0.00384494f $X=4 $Y=1.225 $X2=0
+ $Y2=0
cc_291 N_A_240_394#_c_244_n N_A_640_74#_M1027_d 0.00342046f $X=3.85 $Y=0.34
+ $X2=-0.19 $Y2=-0.245
cc_292 N_A_240_394#_M1002_g N_A_640_74#_c_790_n 0.0100375f $X=3.7 $Y=0.58 $X2=0
+ $Y2=0
cc_293 N_A_240_394#_c_244_n N_A_640_74#_c_790_n 0.0280773f $X=3.85 $Y=0.34 $X2=0
+ $Y2=0
cc_294 N_A_240_394#_c_250_n N_A_640_74#_c_790_n 0.0255025f $X=4 $Y=1.225 $X2=0
+ $Y2=0
cc_295 N_A_240_394#_c_253_n N_A_640_74#_c_779_n 0.00416099f $X=3.625 $Y=1.765
+ $X2=0 $Y2=0
cc_296 N_A_240_394#_M1002_g N_A_640_74#_c_779_n 0.0061534f $X=3.7 $Y=0.58 $X2=0
+ $Y2=0
cc_297 N_A_240_394#_c_249_n N_A_640_74#_c_779_n 0.0155912f $X=3.985 $Y=1.39
+ $X2=0 $Y2=0
cc_298 N_A_240_394#_c_250_n N_A_640_74#_c_779_n 0.044736f $X=4 $Y=1.225 $X2=0
+ $Y2=0
cc_299 N_A_240_394#_c_248_n N_A_640_74#_c_785_n 0.0232488f $X=3.985 $Y=1.39
+ $X2=0 $Y2=0
cc_300 N_A_240_394#_c_249_n N_A_640_74#_c_785_n 0.0111488f $X=3.985 $Y=1.39
+ $X2=0 $Y2=0
cc_301 N_A_240_394#_c_253_n N_A_640_74#_c_786_n 0.0158225f $X=3.625 $Y=1.765
+ $X2=0 $Y2=0
cc_302 N_A_240_394#_c_254_n N_A_640_74#_c_786_n 0.00103999f $X=3.215 $Y=1.765
+ $X2=0 $Y2=0
cc_303 N_A_240_394#_c_249_n N_A_640_74#_c_786_n 9.23073e-19 $X=3.985 $Y=1.39
+ $X2=0 $Y2=0
cc_304 N_A_240_394#_c_248_n N_A_640_74#_c_780_n 0.00558489f $X=3.985 $Y=1.39
+ $X2=0 $Y2=0
cc_305 N_A_240_394#_c_252_n N_A_640_74#_c_803_n 0.0038846f $X=3.125 $Y=1.885
+ $X2=0 $Y2=0
cc_306 N_A_240_394#_c_253_n N_A_640_74#_c_803_n 0.00139529f $X=3.625 $Y=1.765
+ $X2=0 $Y2=0
cc_307 N_A_240_394#_c_252_n N_A_640_74#_c_788_n 0.00613848f $X=3.125 $Y=1.885
+ $X2=0 $Y2=0
cc_308 N_A_240_394#_c_253_n N_A_640_74#_c_788_n 0.00151884f $X=3.625 $Y=1.765
+ $X2=0 $Y2=0
cc_309 N_A_240_394#_c_251_n N_VPWR_c_949_n 0.00616258f $X=2.19 $Y=1.885 $X2=0
+ $Y2=0
cc_310 N_A_240_394#_c_252_n N_VPWR_c_949_n 2.75324e-19 $X=3.125 $Y=1.885 $X2=0
+ $Y2=0
cc_311 N_A_240_394#_c_251_n N_VPWR_c_962_n 0.00469064f $X=2.19 $Y=1.885 $X2=0
+ $Y2=0
cc_312 N_A_240_394#_c_252_n N_VPWR_c_963_n 0.00278271f $X=3.125 $Y=1.885 $X2=0
+ $Y2=0
cc_313 N_A_240_394#_c_251_n N_VPWR_c_947_n 0.0049649f $X=2.19 $Y=1.885 $X2=0
+ $Y2=0
cc_314 N_A_240_394#_c_252_n N_VPWR_c_947_n 0.00354129f $X=3.125 $Y=1.885 $X2=0
+ $Y2=0
cc_315 N_A_240_394#_c_243_n N_VGND_M1024_d 0.0052357f $X=2.835 $Y=0.855 $X2=0
+ $Y2=0
cc_316 N_A_240_394#_c_246_n N_VGND_c_1142_n 0.0324324f $X=1.405 $Y=0.585 $X2=0
+ $Y2=0
cc_317 N_A_240_394#_c_237_n N_VGND_c_1143_n 0.0036648f $X=2.205 $Y=1.45 $X2=0
+ $Y2=0
cc_318 N_A_240_394#_c_243_n N_VGND_c_1143_n 0.0212609f $X=2.835 $Y=0.855 $X2=0
+ $Y2=0
cc_319 N_A_240_394#_c_245_n N_VGND_c_1143_n 0.0117237f $X=3.005 $Y=0.34 $X2=0
+ $Y2=0
cc_320 N_A_240_394#_c_244_n N_VGND_c_1144_n 0.011728f $X=3.85 $Y=0.34 $X2=0
+ $Y2=0
cc_321 N_A_240_394#_c_250_n N_VGND_c_1144_n 0.0137718f $X=4 $Y=1.225 $X2=0 $Y2=0
cc_322 N_A_240_394#_M1002_g N_VGND_c_1151_n 0.00278271f $X=3.7 $Y=0.58 $X2=0
+ $Y2=0
cc_323 N_A_240_394#_c_244_n N_VGND_c_1151_n 0.0655656f $X=3.85 $Y=0.34 $X2=0
+ $Y2=0
cc_324 N_A_240_394#_c_245_n N_VGND_c_1151_n 0.0121935f $X=3.005 $Y=0.34 $X2=0
+ $Y2=0
cc_325 N_A_240_394#_c_237_n N_VGND_c_1153_n 0.00428744f $X=2.205 $Y=1.45 $X2=0
+ $Y2=0
cc_326 N_A_240_394#_c_246_n N_VGND_c_1153_n 0.0134308f $X=1.405 $Y=0.585 $X2=0
+ $Y2=0
cc_327 N_A_240_394#_c_237_n N_VGND_c_1162_n 0.00476395f $X=2.205 $Y=1.45 $X2=0
+ $Y2=0
cc_328 N_A_240_394#_M1002_g N_VGND_c_1162_n 0.00354117f $X=3.7 $Y=0.58 $X2=0
+ $Y2=0
cc_329 N_A_240_394#_c_243_n N_VGND_c_1162_n 0.0319198f $X=2.835 $Y=0.855 $X2=0
+ $Y2=0
cc_330 N_A_240_394#_c_244_n N_VGND_c_1162_n 0.036846f $X=3.85 $Y=0.34 $X2=0
+ $Y2=0
cc_331 N_A_240_394#_c_245_n N_VGND_c_1162_n 0.00661049f $X=3.005 $Y=0.34 $X2=0
+ $Y2=0
cc_332 N_A_240_394#_c_246_n N_VGND_c_1162_n 0.0136871f $X=1.405 $Y=0.585 $X2=0
+ $Y2=0
cc_333 N_A_240_394#_c_243_n A_559_74# 0.00171183f $X=2.835 $Y=0.855 $X2=-0.19
+ $Y2=-0.245
cc_334 N_A_240_394#_c_382_p A_559_74# 3.28781e-19 $X=2.92 $Y=0.77 $X2=-0.19
+ $Y2=-0.245
cc_335 N_A_240_394#_c_244_n A_755_74# 6.48644e-19 $X=3.85 $Y=0.34 $X2=-0.19
+ $Y2=-0.245
cc_336 N_A_240_394#_c_250_n A_755_74# 0.00344737f $X=4 $Y=1.225 $X2=-0.19
+ $Y2=-0.245
cc_337 N_A_240_394#_c_250_n N_A_938_74#_c_1269_n 0.00603064f $X=4 $Y=1.225 $X2=0
+ $Y2=0
cc_338 N_A_27_126#_c_395_n N_A_364_120#_M1016_s 0.00796132f $X=2.495 $Y=2.455
+ $X2=0 $Y2=0
cc_339 N_A_27_126#_M1001_g N_A_364_120#_c_475_n 0.00104046f $X=2.72 $Y=0.69
+ $X2=0 $Y2=0
cc_340 N_A_27_126#_c_387_n N_A_364_120#_c_475_n 0.00131739f $X=2.735 $Y=1.885
+ $X2=0 $Y2=0
cc_341 N_A_27_126#_c_392_n N_A_364_120#_c_475_n 0.028364f $X=2.66 $Y=1.635 $X2=0
+ $Y2=0
cc_342 N_A_27_126#_M1001_g N_A_364_120#_c_476_n 0.0153961f $X=2.72 $Y=0.69 $X2=0
+ $Y2=0
cc_343 N_A_27_126#_c_387_n N_A_364_120#_c_476_n 0.00220216f $X=2.735 $Y=1.885
+ $X2=0 $Y2=0
cc_344 N_A_27_126#_c_392_n N_A_364_120#_c_476_n 0.0200999f $X=2.66 $Y=1.635
+ $X2=0 $Y2=0
cc_345 N_A_27_126#_c_387_n N_A_364_120#_c_478_n 0.006947f $X=2.735 $Y=1.885
+ $X2=0 $Y2=0
cc_346 N_A_27_126#_c_396_n N_A_364_120#_c_478_n 0.0081106f $X=2.58 $Y=2.37 $X2=0
+ $Y2=0
cc_347 N_A_27_126#_c_392_n N_A_364_120#_c_478_n 0.0245577f $X=2.66 $Y=1.635
+ $X2=0 $Y2=0
cc_348 N_A_27_126#_c_387_n N_A_364_120#_c_485_n 0.00113586f $X=2.735 $Y=1.885
+ $X2=0 $Y2=0
cc_349 N_A_27_126#_c_395_n N_A_364_120#_c_487_n 0.0273154f $X=2.495 $Y=2.455
+ $X2=0 $Y2=0
cc_350 N_A_27_126#_c_396_n N_A_364_120#_c_487_n 0.00987581f $X=2.58 $Y=2.37
+ $X2=0 $Y2=0
cc_351 N_A_27_126#_M1001_g N_A_364_120#_c_479_n 0.0172227f $X=2.72 $Y=0.69 $X2=0
+ $Y2=0
cc_352 N_A_27_126#_M1001_g N_A_364_120#_c_480_n 0.0397761f $X=2.72 $Y=0.69 $X2=0
+ $Y2=0
cc_353 N_A_27_126#_c_395_n N_VPWR_M1009_d 0.00691116f $X=2.495 $Y=2.455
+ $X2=-0.19 $Y2=-0.245
cc_354 N_A_27_126#_c_397_n N_VPWR_M1009_d 0.0105582f $X=0.28 $Y=2.115 $X2=-0.19
+ $Y2=-0.245
cc_355 N_A_27_126#_c_395_n N_VPWR_M1016_d 0.00997037f $X=2.495 $Y=2.455 $X2=0
+ $Y2=0
cc_356 N_A_27_126#_c_396_n N_VPWR_M1016_d 0.00445296f $X=2.58 $Y=2.37 $X2=0
+ $Y2=0
cc_357 N_A_27_126#_c_395_n N_VPWR_c_948_n 0.00981701f $X=2.495 $Y=2.455 $X2=0
+ $Y2=0
cc_358 N_A_27_126#_c_397_n N_VPWR_c_948_n 0.0260068f $X=0.28 $Y=2.115 $X2=0
+ $Y2=0
cc_359 N_A_27_126#_c_387_n N_VPWR_c_949_n 0.00613608f $X=2.735 $Y=1.885 $X2=0
+ $Y2=0
cc_360 N_A_27_126#_c_395_n N_VPWR_c_949_n 0.0223222f $X=2.495 $Y=2.455 $X2=0
+ $Y2=0
cc_361 N_A_27_126#_c_387_n N_VPWR_c_963_n 0.00444681f $X=2.735 $Y=1.885 $X2=0
+ $Y2=0
cc_362 N_A_27_126#_c_397_n N_VPWR_c_965_n 0.00908884f $X=0.28 $Y=2.115 $X2=0
+ $Y2=0
cc_363 N_A_27_126#_c_387_n N_VPWR_c_947_n 0.00877228f $X=2.735 $Y=1.885 $X2=0
+ $Y2=0
cc_364 N_A_27_126#_c_395_n N_VPWR_c_947_n 0.0496159f $X=2.495 $Y=2.455 $X2=0
+ $Y2=0
cc_365 N_A_27_126#_c_397_n N_VPWR_c_947_n 0.019667f $X=0.28 $Y=2.115 $X2=0 $Y2=0
cc_366 N_A_27_126#_c_389_n N_VGND_M1019_d 0.0052407f $X=0.685 $Y=1.195 $X2=-0.19
+ $Y2=-0.245
cc_367 N_A_27_126#_c_388_n N_VGND_c_1142_n 0.019979f $X=0.28 $Y=0.905 $X2=0
+ $Y2=0
cc_368 N_A_27_126#_c_389_n N_VGND_c_1142_n 0.0153275f $X=0.685 $Y=1.195 $X2=0
+ $Y2=0
cc_369 N_A_27_126#_M1001_g N_VGND_c_1143_n 0.00688998f $X=2.72 $Y=0.69 $X2=0
+ $Y2=0
cc_370 N_A_27_126#_M1001_g N_VGND_c_1151_n 0.00398535f $X=2.72 $Y=0.69 $X2=0
+ $Y2=0
cc_371 N_A_27_126#_c_388_n N_VGND_c_1157_n 0.00693787f $X=0.28 $Y=0.905 $X2=0
+ $Y2=0
cc_372 N_A_27_126#_M1001_g N_VGND_c_1162_n 0.00383716f $X=2.72 $Y=0.69 $X2=0
+ $Y2=0
cc_373 N_A_27_126#_c_388_n N_VGND_c_1162_n 0.0101027f $X=0.28 $Y=0.905 $X2=0
+ $Y2=0
cc_374 N_A_364_120#_c_481_n N_A_797_48#_c_597_n 0.0352503f $X=3.66 $Y=2.465
+ $X2=0 $Y2=0
cc_375 N_A_364_120#_c_484_n N_A_797_48#_c_597_n 0.001726f $X=3.655 $Y=2.99 $X2=0
+ $Y2=0
cc_376 N_A_364_120#_c_486_n N_A_797_48#_c_597_n 0.00722594f $X=3.82 $Y=2.215
+ $X2=0 $Y2=0
cc_377 N_A_364_120#_c_481_n N_A_797_48#_c_603_n 0.00125622f $X=3.66 $Y=2.465
+ $X2=0 $Y2=0
cc_378 N_A_364_120#_c_486_n N_A_797_48#_c_603_n 0.0282952f $X=3.82 $Y=2.215
+ $X2=0 $Y2=0
cc_379 N_A_364_120#_c_484_n N_A_640_74#_M1008_d 0.00471713f $X=3.655 $Y=2.99
+ $X2=0 $Y2=0
cc_380 N_A_364_120#_c_476_n N_A_640_74#_c_790_n 0.0103344f $X=2.955 $Y=1.195
+ $X2=0 $Y2=0
cc_381 N_A_364_120#_c_479_n N_A_640_74#_c_790_n 0.00186128f $X=3.2 $Y=1.285
+ $X2=0 $Y2=0
cc_382 N_A_364_120#_c_480_n N_A_640_74#_c_790_n 0.00398872f $X=3.2 $Y=1.12 $X2=0
+ $Y2=0
cc_383 N_A_364_120#_c_476_n N_A_640_74#_c_779_n 0.025899f $X=2.955 $Y=1.195
+ $X2=0 $Y2=0
cc_384 N_A_364_120#_c_478_n N_A_640_74#_c_779_n 0.0114796f $X=3.04 $Y=1.97 $X2=0
+ $Y2=0
cc_385 N_A_364_120#_c_479_n N_A_640_74#_c_779_n 0.00205802f $X=3.2 $Y=1.285
+ $X2=0 $Y2=0
cc_386 N_A_364_120#_c_480_n N_A_640_74#_c_779_n 0.00319937f $X=3.2 $Y=1.12 $X2=0
+ $Y2=0
cc_387 N_A_364_120#_c_481_n N_A_640_74#_c_786_n 0.00442567f $X=3.66 $Y=2.465
+ $X2=0 $Y2=0
cc_388 N_A_364_120#_c_476_n N_A_640_74#_c_786_n 0.00215189f $X=2.955 $Y=1.195
+ $X2=0 $Y2=0
cc_389 N_A_364_120#_c_478_n N_A_640_74#_c_786_n 0.0130063f $X=3.04 $Y=1.97 $X2=0
+ $Y2=0
cc_390 N_A_364_120#_c_486_n N_A_640_74#_c_786_n 0.0261741f $X=3.82 $Y=2.215
+ $X2=0 $Y2=0
cc_391 N_A_364_120#_c_479_n N_A_640_74#_c_786_n 2.22933e-19 $X=3.2 $Y=1.285
+ $X2=0 $Y2=0
cc_392 N_A_364_120#_c_481_n N_A_640_74#_c_803_n 0.0021223f $X=3.66 $Y=2.465
+ $X2=0 $Y2=0
cc_393 N_A_364_120#_c_484_n N_A_640_74#_c_803_n 0.0165122f $X=3.655 $Y=2.99
+ $X2=0 $Y2=0
cc_394 N_A_364_120#_c_481_n N_A_640_74#_c_788_n 0.00385009f $X=3.66 $Y=2.465
+ $X2=0 $Y2=0
cc_395 N_A_364_120#_c_478_n N_A_640_74#_c_788_n 0.00535066f $X=3.04 $Y=1.97
+ $X2=0 $Y2=0
cc_396 N_A_364_120#_c_486_n N_A_640_74#_c_788_n 0.046187f $X=3.82 $Y=2.215 $X2=0
+ $Y2=0
cc_397 N_A_364_120#_c_518_n N_A_640_74#_c_788_n 0.0123107f $X=3.04 $Y=2.055
+ $X2=0 $Y2=0
cc_398 N_A_364_120#_c_485_n N_VPWR_c_949_n 0.0112232f $X=3.015 $Y=2.99 $X2=0
+ $Y2=0
cc_399 N_A_364_120#_c_481_n N_VPWR_c_950_n 4.07984e-19 $X=3.66 $Y=2.465 $X2=0
+ $Y2=0
cc_400 N_A_364_120#_c_484_n N_VPWR_c_950_n 0.00839268f $X=3.655 $Y=2.99 $X2=0
+ $Y2=0
cc_401 N_A_364_120#_c_486_n N_VPWR_c_950_n 0.0115445f $X=3.82 $Y=2.215 $X2=0
+ $Y2=0
cc_402 N_A_364_120#_c_481_n N_VPWR_c_963_n 0.00278193f $X=3.66 $Y=2.465 $X2=0
+ $Y2=0
cc_403 N_A_364_120#_c_484_n N_VPWR_c_963_n 0.0638747f $X=3.655 $Y=2.99 $X2=0
+ $Y2=0
cc_404 N_A_364_120#_c_485_n N_VPWR_c_963_n 0.0121867f $X=3.015 $Y=2.99 $X2=0
+ $Y2=0
cc_405 N_A_364_120#_c_481_n N_VPWR_c_947_n 0.00356044f $X=3.66 $Y=2.465 $X2=0
+ $Y2=0
cc_406 N_A_364_120#_c_484_n N_VPWR_c_947_n 0.0355129f $X=3.655 $Y=2.99 $X2=0
+ $Y2=0
cc_407 N_A_364_120#_c_485_n N_VPWR_c_947_n 0.00660921f $X=3.015 $Y=2.99 $X2=0
+ $Y2=0
cc_408 N_A_364_120#_c_572_p A_562_392# 0.00327032f $X=2.93 $Y=2.905 $X2=-0.19
+ $Y2=-0.245
cc_409 N_A_364_120#_c_478_n A_562_392# 2.12418e-19 $X=3.04 $Y=1.97 $X2=-0.19
+ $Y2=-0.245
cc_410 N_A_364_120#_c_518_n A_562_392# 0.00387782f $X=3.04 $Y=2.055 $X2=-0.19
+ $Y2=-0.245
cc_411 N_A_364_120#_c_484_n A_747_508# 8.83155e-19 $X=3.655 $Y=2.99 $X2=-0.19
+ $Y2=-0.245
cc_412 N_A_364_120#_c_486_n A_747_508# 0.00570902f $X=3.82 $Y=2.215 $X2=-0.19
+ $Y2=-0.245
cc_413 N_A_364_120#_c_476_n N_VGND_M1024_d 0.0084682f $X=2.955 $Y=1.195 $X2=0
+ $Y2=0
cc_414 N_A_364_120#_c_480_n N_VGND_c_1143_n 2.69111e-19 $X=3.2 $Y=1.12 $X2=0
+ $Y2=0
cc_415 N_A_364_120#_c_480_n N_VGND_c_1151_n 0.00278271f $X=3.2 $Y=1.12 $X2=0
+ $Y2=0
cc_416 N_A_364_120#_c_480_n N_VGND_c_1162_n 0.00354575f $X=3.2 $Y=1.12 $X2=0
+ $Y2=0
cc_417 N_A_797_48#_c_582_n N_A_640_74#_M1000_g 0.0107002f $X=4.36 $Y=0.94 $X2=0
+ $Y2=0
cc_418 N_A_797_48#_c_589_n N_A_640_74#_M1000_g 0.00800438f $X=5.275 $Y=1.62
+ $X2=0 $Y2=0
cc_419 N_A_797_48#_c_597_n N_A_640_74#_c_774_n 0.0151176f $X=4.285 $Y=2.465
+ $X2=0 $Y2=0
cc_420 N_A_797_48#_c_584_n N_A_640_74#_c_774_n 0.0304384f $X=4.435 $Y=2.05 $X2=0
+ $Y2=0
cc_421 N_A_797_48#_c_603_n N_A_640_74#_c_774_n 0.037179f $X=5.11 $Y=2.272 $X2=0
+ $Y2=0
cc_422 N_A_797_48#_c_589_n N_A_640_74#_c_774_n 9.59198e-19 $X=5.275 $Y=1.62
+ $X2=0 $Y2=0
cc_423 N_A_797_48#_c_604_n N_A_640_74#_c_774_n 0.00411748f $X=5.275 $Y=1.965
+ $X2=0 $Y2=0
cc_424 N_A_797_48#_c_592_n N_A_640_74#_c_774_n 0.00144296f $X=5.315 $Y=1.705
+ $X2=0 $Y2=0
cc_425 N_A_797_48#_c_589_n N_A_640_74#_c_775_n 0.0117026f $X=5.275 $Y=1.62 $X2=0
+ $Y2=0
cc_426 N_A_797_48#_c_589_n N_A_640_74#_M1006_g 0.00548896f $X=5.275 $Y=1.62
+ $X2=0 $Y2=0
cc_427 N_A_797_48#_c_589_n N_A_640_74#_c_777_n 0.00286293f $X=5.275 $Y=1.62
+ $X2=0 $Y2=0
cc_428 N_A_797_48#_c_590_n N_A_640_74#_c_777_n 0.00706648f $X=6.11 $Y=1.705
+ $X2=0 $Y2=0
cc_429 N_A_797_48#_c_592_n N_A_640_74#_c_777_n 0.00218178f $X=5.315 $Y=1.705
+ $X2=0 $Y2=0
cc_430 N_A_797_48#_c_603_n N_A_640_74#_c_783_n 0.00882052f $X=5.11 $Y=2.272
+ $X2=0 $Y2=0
cc_431 N_A_797_48#_c_604_n N_A_640_74#_c_783_n 0.00472301f $X=5.275 $Y=1.965
+ $X2=0 $Y2=0
cc_432 N_A_797_48#_c_590_n N_A_640_74#_c_783_n 0.00918933f $X=6.11 $Y=1.705
+ $X2=0 $Y2=0
cc_433 N_A_797_48#_c_592_n N_A_640_74#_c_783_n 0.00168501f $X=5.315 $Y=1.705
+ $X2=0 $Y2=0
cc_434 N_A_797_48#_c_581_n N_A_640_74#_c_790_n 2.75457e-19 $X=4.06 $Y=0.865
+ $X2=0 $Y2=0
cc_435 N_A_797_48#_c_584_n N_A_640_74#_c_779_n 8.2402e-19 $X=4.435 $Y=2.05 $X2=0
+ $Y2=0
cc_436 N_A_797_48#_c_597_n N_A_640_74#_c_785_n 0.0047245f $X=4.285 $Y=2.465
+ $X2=0 $Y2=0
cc_437 N_A_797_48#_c_584_n N_A_640_74#_c_785_n 0.0173533f $X=4.435 $Y=2.05 $X2=0
+ $Y2=0
cc_438 N_A_797_48#_c_603_n N_A_640_74#_c_785_n 0.0608084f $X=5.11 $Y=2.272 $X2=0
+ $Y2=0
cc_439 N_A_797_48#_c_604_n N_A_640_74#_c_785_n 0.00851136f $X=5.275 $Y=1.965
+ $X2=0 $Y2=0
cc_440 N_A_797_48#_c_592_n N_A_640_74#_c_785_n 0.00575192f $X=5.315 $Y=1.705
+ $X2=0 $Y2=0
cc_441 N_A_797_48#_c_584_n N_A_640_74#_c_780_n 0.00267497f $X=4.435 $Y=2.05
+ $X2=0 $Y2=0
cc_442 N_A_797_48#_c_589_n N_A_640_74#_c_780_n 0.019545f $X=5.275 $Y=1.62 $X2=0
+ $Y2=0
cc_443 N_A_797_48#_c_592_n N_A_640_74#_c_780_n 0.00875914f $X=5.315 $Y=1.705
+ $X2=0 $Y2=0
cc_444 N_A_797_48#_c_589_n N_RESET_B_c_884_n 2.03747e-19 $X=5.275 $Y=1.62 $X2=0
+ $Y2=0
cc_445 N_A_797_48#_c_590_n N_RESET_B_c_884_n 0.0047603f $X=6.11 $Y=1.705 $X2=0
+ $Y2=0
cc_446 N_A_797_48#_c_604_n N_RESET_B_c_890_n 5.41384e-19 $X=5.275 $Y=1.965 $X2=0
+ $Y2=0
cc_447 N_A_797_48#_c_590_n N_RESET_B_c_890_n 0.0115103f $X=6.11 $Y=1.705 $X2=0
+ $Y2=0
cc_448 N_A_797_48#_c_606_n N_RESET_B_c_890_n 0.00541891f $X=6.275 $Y=1.985 $X2=0
+ $Y2=0
cc_449 N_A_797_48#_c_593_n N_RESET_B_c_886_n 0.00130753f $X=6.275 $Y=1.705 $X2=0
+ $Y2=0
cc_450 N_A_797_48#_c_594_n N_RESET_B_c_886_n 0.00346963f $X=6.765 $Y=1.545 $X2=0
+ $Y2=0
cc_451 N_A_797_48#_c_599_n N_RESET_B_c_892_n 0.0134013f $X=7.035 $Y=1.765 $X2=0
+ $Y2=0
cc_452 N_A_797_48#_c_606_n N_RESET_B_c_892_n 0.0139459f $X=6.275 $Y=1.985 $X2=0
+ $Y2=0
cc_453 N_A_797_48#_c_593_n N_RESET_B_c_892_n 0.00220783f $X=6.275 $Y=1.705 $X2=0
+ $Y2=0
cc_454 N_A_797_48#_c_594_n N_RESET_B_c_892_n 0.00915018f $X=6.765 $Y=1.545 $X2=0
+ $Y2=0
cc_455 N_A_797_48#_M1011_g RESET_B 0.00299663f $X=7.335 $Y=0.74 $X2=0 $Y2=0
cc_456 N_A_797_48#_c_589_n RESET_B 0.0107502f $X=5.275 $Y=1.62 $X2=0 $Y2=0
cc_457 N_A_797_48#_c_590_n RESET_B 0.016199f $X=6.11 $Y=1.705 $X2=0 $Y2=0
cc_458 N_A_797_48#_c_593_n RESET_B 0.0276979f $X=6.275 $Y=1.705 $X2=0 $Y2=0
cc_459 N_A_797_48#_c_594_n RESET_B 0.0110744f $X=6.765 $Y=1.545 $X2=0 $Y2=0
cc_460 N_A_797_48#_c_595_n RESET_B 0.0139089f $X=6.935 $Y=1.545 $X2=0 $Y2=0
cc_461 N_A_797_48#_c_596_n RESET_B 4.10407e-19 $X=8.505 $Y=1.532 $X2=0 $Y2=0
cc_462 N_A_797_48#_M1011_g N_RESET_B_c_888_n 0.00215545f $X=7.335 $Y=0.74 $X2=0
+ $Y2=0
cc_463 N_A_797_48#_c_589_n N_RESET_B_c_888_n 3.11476e-19 $X=5.275 $Y=1.62 $X2=0
+ $Y2=0
cc_464 N_A_797_48#_c_590_n N_RESET_B_c_888_n 0.00206683f $X=6.11 $Y=1.705 $X2=0
+ $Y2=0
cc_465 N_A_797_48#_c_593_n N_RESET_B_c_888_n 0.00381358f $X=6.275 $Y=1.705 $X2=0
+ $Y2=0
cc_466 N_A_797_48#_c_595_n N_RESET_B_c_888_n 0.00545341f $X=6.935 $Y=1.545 $X2=0
+ $Y2=0
cc_467 N_A_797_48#_c_596_n N_RESET_B_c_888_n 0.0143445f $X=8.505 $Y=1.532 $X2=0
+ $Y2=0
cc_468 N_A_797_48#_c_603_n N_VPWR_M1003_d 0.00629892f $X=5.11 $Y=2.272 $X2=0
+ $Y2=0
cc_469 N_A_797_48#_c_597_n N_VPWR_c_950_n 0.0170985f $X=4.285 $Y=2.465 $X2=0
+ $Y2=0
cc_470 N_A_797_48#_c_603_n N_VPWR_c_950_n 0.048649f $X=5.11 $Y=2.272 $X2=0 $Y2=0
cc_471 N_A_797_48#_c_604_n N_VPWR_c_951_n 0.028357f $X=5.275 $Y=1.965 $X2=0
+ $Y2=0
cc_472 N_A_797_48#_c_590_n N_VPWR_c_951_n 0.0234881f $X=6.11 $Y=1.705 $X2=0
+ $Y2=0
cc_473 N_A_797_48#_c_606_n N_VPWR_c_951_n 0.028557f $X=6.275 $Y=1.985 $X2=0
+ $Y2=0
cc_474 N_A_797_48#_c_599_n N_VPWR_c_952_n 0.015653f $X=7.035 $Y=1.765 $X2=0
+ $Y2=0
cc_475 N_A_797_48#_c_600_n N_VPWR_c_952_n 6.73991e-19 $X=7.485 $Y=1.765 $X2=0
+ $Y2=0
cc_476 N_A_797_48#_c_606_n N_VPWR_c_952_n 0.0497671f $X=6.275 $Y=1.985 $X2=0
+ $Y2=0
cc_477 N_A_797_48#_c_591_n N_VPWR_c_952_n 0.00119971f $X=8.43 $Y=1.465 $X2=0
+ $Y2=0
cc_478 N_A_797_48#_c_594_n N_VPWR_c_952_n 0.023541f $X=6.765 $Y=1.545 $X2=0
+ $Y2=0
cc_479 N_A_797_48#_c_600_n N_VPWR_c_953_n 0.00621531f $X=7.485 $Y=1.765 $X2=0
+ $Y2=0
cc_480 N_A_797_48#_c_601_n N_VPWR_c_953_n 0.0146474f $X=7.985 $Y=1.765 $X2=0
+ $Y2=0
cc_481 N_A_797_48#_c_602_n N_VPWR_c_953_n 5.23608e-19 $X=8.505 $Y=1.765 $X2=0
+ $Y2=0
cc_482 N_A_797_48#_c_602_n N_VPWR_c_955_n 0.00787188f $X=8.505 $Y=1.765 $X2=0
+ $Y2=0
cc_483 N_A_797_48#_c_603_n N_VPWR_c_956_n 0.00663854f $X=5.11 $Y=2.272 $X2=0
+ $Y2=0
cc_484 N_A_797_48#_c_606_n N_VPWR_c_958_n 0.0066794f $X=6.275 $Y=1.985 $X2=0
+ $Y2=0
cc_485 N_A_797_48#_c_599_n N_VPWR_c_960_n 0.00413917f $X=7.035 $Y=1.765 $X2=0
+ $Y2=0
cc_486 N_A_797_48#_c_600_n N_VPWR_c_960_n 0.00445602f $X=7.485 $Y=1.765 $X2=0
+ $Y2=0
cc_487 N_A_797_48#_c_597_n N_VPWR_c_963_n 0.00413917f $X=4.285 $Y=2.465 $X2=0
+ $Y2=0
cc_488 N_A_797_48#_c_601_n N_VPWR_c_964_n 0.00413917f $X=7.985 $Y=1.765 $X2=0
+ $Y2=0
cc_489 N_A_797_48#_c_602_n N_VPWR_c_964_n 0.00461464f $X=8.505 $Y=1.765 $X2=0
+ $Y2=0
cc_490 N_A_797_48#_c_597_n N_VPWR_c_947_n 0.00418196f $X=4.285 $Y=2.465 $X2=0
+ $Y2=0
cc_491 N_A_797_48#_c_599_n N_VPWR_c_947_n 0.00817726f $X=7.035 $Y=1.765 $X2=0
+ $Y2=0
cc_492 N_A_797_48#_c_600_n N_VPWR_c_947_n 0.00857378f $X=7.485 $Y=1.765 $X2=0
+ $Y2=0
cc_493 N_A_797_48#_c_601_n N_VPWR_c_947_n 0.0081836f $X=7.985 $Y=1.765 $X2=0
+ $Y2=0
cc_494 N_A_797_48#_c_602_n N_VPWR_c_947_n 0.0091227f $X=8.505 $Y=1.765 $X2=0
+ $Y2=0
cc_495 N_A_797_48#_c_603_n N_VPWR_c_947_n 0.0236112f $X=5.11 $Y=2.272 $X2=0
+ $Y2=0
cc_496 N_A_797_48#_c_606_n N_VPWR_c_947_n 0.00997343f $X=6.275 $Y=1.985 $X2=0
+ $Y2=0
cc_497 N_A_797_48#_c_599_n N_Q_c_1072_n 0.00378511f $X=7.035 $Y=1.765 $X2=0
+ $Y2=0
cc_498 N_A_797_48#_c_600_n N_Q_c_1072_n 0.0120819f $X=7.485 $Y=1.765 $X2=0 $Y2=0
cc_499 N_A_797_48#_c_601_n N_Q_c_1072_n 5.64826e-19 $X=7.985 $Y=1.765 $X2=0
+ $Y2=0
cc_500 N_A_797_48#_M1011_g N_Q_c_1065_n 0.00326509f $X=7.335 $Y=0.74 $X2=0 $Y2=0
cc_501 N_A_797_48#_c_591_n N_Q_c_1065_n 0.0218166f $X=8.43 $Y=1.465 $X2=0 $Y2=0
cc_502 N_A_797_48#_c_596_n N_Q_c_1065_n 0.00259093f $X=8.505 $Y=1.532 $X2=0
+ $Y2=0
cc_503 N_A_797_48#_M1011_g N_Q_c_1066_n 0.00615025f $X=7.335 $Y=0.74 $X2=0 $Y2=0
cc_504 N_A_797_48#_M1015_g N_Q_c_1066_n 2.27367e-19 $X=7.765 $Y=0.74 $X2=0 $Y2=0
cc_505 N_A_797_48#_c_600_n N_Q_c_1073_n 0.0122806f $X=7.485 $Y=1.765 $X2=0 $Y2=0
cc_506 N_A_797_48#_c_601_n N_Q_c_1073_n 0.0155315f $X=7.985 $Y=1.765 $X2=0 $Y2=0
cc_507 N_A_797_48#_c_591_n N_Q_c_1073_n 0.0492159f $X=8.43 $Y=1.465 $X2=0 $Y2=0
cc_508 N_A_797_48#_c_596_n N_Q_c_1073_n 0.0102128f $X=8.505 $Y=1.532 $X2=0 $Y2=0
cc_509 N_A_797_48#_c_599_n N_Q_c_1074_n 0.00455961f $X=7.035 $Y=1.765 $X2=0
+ $Y2=0
cc_510 N_A_797_48#_c_600_n N_Q_c_1074_n 8.24772e-19 $X=7.485 $Y=1.765 $X2=0
+ $Y2=0
cc_511 N_A_797_48#_c_591_n N_Q_c_1074_n 0.0210155f $X=8.43 $Y=1.465 $X2=0 $Y2=0
cc_512 N_A_797_48#_c_596_n N_Q_c_1074_n 0.00613849f $X=8.505 $Y=1.532 $X2=0
+ $Y2=0
cc_513 N_A_797_48#_M1015_g N_Q_c_1067_n 0.0146497f $X=7.765 $Y=0.74 $X2=0 $Y2=0
cc_514 N_A_797_48#_M1023_g N_Q_c_1067_n 0.0146497f $X=8.195 $Y=0.74 $X2=0 $Y2=0
cc_515 N_A_797_48#_c_591_n N_Q_c_1067_n 0.0506171f $X=8.43 $Y=1.465 $X2=0 $Y2=0
cc_516 N_A_797_48#_c_596_n N_Q_c_1067_n 0.00265643f $X=8.505 $Y=1.532 $X2=0
+ $Y2=0
cc_517 N_A_797_48#_c_601_n N_Q_c_1075_n 0.0056973f $X=7.985 $Y=1.765 $X2=0 $Y2=0
cc_518 N_A_797_48#_c_602_n N_Q_c_1075_n 4.83874e-19 $X=8.505 $Y=1.765 $X2=0
+ $Y2=0
cc_519 N_A_797_48#_M1023_g N_Q_c_1068_n 2.26494e-19 $X=8.195 $Y=0.74 $X2=0 $Y2=0
cc_520 N_A_797_48#_M1029_g N_Q_c_1068_n 2.26494e-19 $X=8.625 $Y=0.74 $X2=0 $Y2=0
cc_521 N_A_797_48#_c_602_n N_Q_c_1076_n 0.0152094f $X=8.505 $Y=1.765 $X2=0 $Y2=0
cc_522 N_A_797_48#_c_591_n N_Q_c_1076_n 0.0121772f $X=8.43 $Y=1.465 $X2=0 $Y2=0
cc_523 N_A_797_48#_c_596_n N_Q_c_1076_n 0.00324158f $X=8.505 $Y=1.532 $X2=0
+ $Y2=0
cc_524 N_A_797_48#_M1029_g N_Q_c_1069_n 0.0176989f $X=8.625 $Y=0.74 $X2=0 $Y2=0
cc_525 N_A_797_48#_c_591_n N_Q_c_1069_n 0.00675171f $X=8.43 $Y=1.465 $X2=0 $Y2=0
cc_526 N_A_797_48#_c_591_n N_Q_c_1077_n 0.0278299f $X=8.43 $Y=1.465 $X2=0 $Y2=0
cc_527 N_A_797_48#_c_596_n N_Q_c_1077_n 0.00879386f $X=8.505 $Y=1.532 $X2=0
+ $Y2=0
cc_528 N_A_797_48#_c_591_n N_Q_c_1070_n 0.0160251f $X=8.43 $Y=1.465 $X2=0 $Y2=0
cc_529 N_A_797_48#_c_596_n N_Q_c_1070_n 0.00247261f $X=8.505 $Y=1.532 $X2=0
+ $Y2=0
cc_530 N_A_797_48#_c_602_n Q 0.00118721f $X=8.505 $Y=1.765 $X2=0 $Y2=0
cc_531 N_A_797_48#_M1029_g Q 0.0112421f $X=8.625 $Y=0.74 $X2=0 $Y2=0
cc_532 N_A_797_48#_c_591_n Q 0.0267934f $X=8.43 $Y=1.465 $X2=0 $Y2=0
cc_533 N_A_797_48#_c_596_n Q 0.00620365f $X=8.505 $Y=1.532 $X2=0 $Y2=0
cc_534 N_A_797_48#_c_581_n N_VGND_c_1144_n 0.00413902f $X=4.06 $Y=0.865 $X2=0
+ $Y2=0
cc_535 N_A_797_48#_c_582_n N_VGND_c_1144_n 0.0121899f $X=4.36 $Y=0.94 $X2=0
+ $Y2=0
cc_536 N_A_797_48#_M1011_g N_VGND_c_1147_n 0.00486281f $X=7.335 $Y=0.74 $X2=0
+ $Y2=0
cc_537 N_A_797_48#_c_591_n N_VGND_c_1147_n 0.021758f $X=8.43 $Y=1.465 $X2=0
+ $Y2=0
cc_538 N_A_797_48#_c_596_n N_VGND_c_1147_n 0.00663321f $X=8.505 $Y=1.532 $X2=0
+ $Y2=0
cc_539 N_A_797_48#_M1011_g N_VGND_c_1148_n 4.8057e-19 $X=7.335 $Y=0.74 $X2=0
+ $Y2=0
cc_540 N_A_797_48#_M1015_g N_VGND_c_1148_n 0.00811288f $X=7.765 $Y=0.74 $X2=0
+ $Y2=0
cc_541 N_A_797_48#_M1023_g N_VGND_c_1148_n 0.00797557f $X=8.195 $Y=0.74 $X2=0
+ $Y2=0
cc_542 N_A_797_48#_M1029_g N_VGND_c_1148_n 4.67172e-19 $X=8.625 $Y=0.74 $X2=0
+ $Y2=0
cc_543 N_A_797_48#_M1023_g N_VGND_c_1150_n 4.67172e-19 $X=8.195 $Y=0.74 $X2=0
+ $Y2=0
cc_544 N_A_797_48#_M1029_g N_VGND_c_1150_n 0.00908683f $X=8.625 $Y=0.74 $X2=0
+ $Y2=0
cc_545 N_A_797_48#_c_581_n N_VGND_c_1151_n 0.00418685f $X=4.06 $Y=0.865 $X2=0
+ $Y2=0
cc_546 N_A_797_48#_M1011_g N_VGND_c_1155_n 0.00434596f $X=7.335 $Y=0.74 $X2=0
+ $Y2=0
cc_547 N_A_797_48#_M1015_g N_VGND_c_1155_n 0.00383152f $X=7.765 $Y=0.74 $X2=0
+ $Y2=0
cc_548 N_A_797_48#_M1023_g N_VGND_c_1156_n 0.00383152f $X=8.195 $Y=0.74 $X2=0
+ $Y2=0
cc_549 N_A_797_48#_M1029_g N_VGND_c_1156_n 0.00383152f $X=8.625 $Y=0.74 $X2=0
+ $Y2=0
cc_550 N_A_797_48#_c_581_n N_VGND_c_1162_n 0.00783021f $X=4.06 $Y=0.865 $X2=0
+ $Y2=0
cc_551 N_A_797_48#_c_582_n N_VGND_c_1162_n 0.00290734f $X=4.36 $Y=0.94 $X2=0
+ $Y2=0
cc_552 N_A_797_48#_M1011_g N_VGND_c_1162_n 0.00825326f $X=7.335 $Y=0.74 $X2=0
+ $Y2=0
cc_553 N_A_797_48#_M1015_g N_VGND_c_1162_n 0.0075754f $X=7.765 $Y=0.74 $X2=0
+ $Y2=0
cc_554 N_A_797_48#_M1023_g N_VGND_c_1162_n 0.0075754f $X=8.195 $Y=0.74 $X2=0
+ $Y2=0
cc_555 N_A_797_48#_M1029_g N_VGND_c_1162_n 0.0075754f $X=8.625 $Y=0.74 $X2=0
+ $Y2=0
cc_556 N_A_797_48#_c_581_n N_A_938_74#_c_1269_n 0.00148506f $X=4.06 $Y=0.865
+ $X2=0 $Y2=0
cc_557 N_A_797_48#_c_582_n N_A_938_74#_c_1269_n 0.00248848f $X=4.36 $Y=0.94
+ $X2=0 $Y2=0
cc_558 N_A_797_48#_c_589_n N_A_938_74#_c_1269_n 0.00541431f $X=5.275 $Y=1.62
+ $X2=0 $Y2=0
cc_559 N_A_797_48#_M1000_s N_A_938_74#_c_1270_n 0.00181776f $X=5.125 $Y=0.37
+ $X2=0 $Y2=0
cc_560 N_A_797_48#_c_769_p N_A_938_74#_c_1270_n 0.0130519f $X=5.265 $Y=0.785
+ $X2=0 $Y2=0
cc_561 N_A_797_48#_c_590_n N_A_938_74#_c_1280_n 0.00637007f $X=6.11 $Y=1.705
+ $X2=0 $Y2=0
cc_562 N_A_797_48#_c_590_n N_A_938_74#_c_1281_n 0.00191168f $X=6.11 $Y=1.705
+ $X2=0 $Y2=0
cc_563 N_A_797_48#_c_594_n N_A_938_74#_c_1272_n 0.00395242f $X=6.765 $Y=1.545
+ $X2=0 $Y2=0
cc_564 N_A_640_74#_M1006_g N_RESET_B_c_883_n 0.014182f $X=5.485 $Y=0.69
+ $X2=-0.19 $Y2=-0.245
cc_565 N_A_640_74#_c_778_n N_RESET_B_c_884_n 0.00640412f $X=5.5 $Y=1.425 $X2=0
+ $Y2=0
cc_566 N_A_640_74#_c_777_n N_RESET_B_c_890_n 0.00640412f $X=5.5 $Y=1.675 $X2=0
+ $Y2=0
cc_567 N_A_640_74#_c_783_n N_RESET_B_c_890_n 0.0189663f $X=5.5 $Y=1.765 $X2=0
+ $Y2=0
cc_568 N_A_640_74#_M1006_g RESET_B 2.70034e-19 $X=5.485 $Y=0.69 $X2=0 $Y2=0
cc_569 N_A_640_74#_c_778_n RESET_B 9.68654e-19 $X=5.5 $Y=1.425 $X2=0 $Y2=0
cc_570 N_A_640_74#_c_778_n N_RESET_B_c_888_n 0.0139072f $X=5.5 $Y=1.425 $X2=0
+ $Y2=0
cc_571 N_A_640_74#_c_785_n N_VPWR_M1003_d 0.00239978f $X=4.72 $Y=1.81 $X2=0
+ $Y2=0
cc_572 N_A_640_74#_c_774_n N_VPWR_c_950_n 0.00425767f $X=5.05 $Y=1.765 $X2=0
+ $Y2=0
cc_573 N_A_640_74#_c_783_n N_VPWR_c_951_n 0.00716215f $X=5.5 $Y=1.765 $X2=0
+ $Y2=0
cc_574 N_A_640_74#_c_774_n N_VPWR_c_956_n 0.00393873f $X=5.05 $Y=1.765 $X2=0
+ $Y2=0
cc_575 N_A_640_74#_c_783_n N_VPWR_c_956_n 0.00393873f $X=5.5 $Y=1.765 $X2=0
+ $Y2=0
cc_576 N_A_640_74#_c_774_n N_VPWR_c_947_n 0.00462577f $X=5.05 $Y=1.765 $X2=0
+ $Y2=0
cc_577 N_A_640_74#_c_783_n N_VPWR_c_947_n 0.00462577f $X=5.5 $Y=1.765 $X2=0
+ $Y2=0
cc_578 N_A_640_74#_M1000_g N_VGND_c_1144_n 0.0019888f $X=5.05 $Y=0.69 $X2=0
+ $Y2=0
cc_579 N_A_640_74#_M1006_g N_VGND_c_1145_n 3.45328e-19 $X=5.485 $Y=0.69 $X2=0
+ $Y2=0
cc_580 N_A_640_74#_M1000_g N_VGND_c_1154_n 0.00281867f $X=5.05 $Y=0.69 $X2=0
+ $Y2=0
cc_581 N_A_640_74#_M1006_g N_VGND_c_1154_n 0.00281867f $X=5.485 $Y=0.69 $X2=0
+ $Y2=0
cc_582 N_A_640_74#_M1000_g N_VGND_c_1162_n 0.00359088f $X=5.05 $Y=0.69 $X2=0
+ $Y2=0
cc_583 N_A_640_74#_M1006_g N_VGND_c_1162_n 0.00354187f $X=5.485 $Y=0.69 $X2=0
+ $Y2=0
cc_584 N_A_640_74#_M1000_g N_A_938_74#_c_1269_n 0.0079864f $X=5.05 $Y=0.69 $X2=0
+ $Y2=0
cc_585 N_A_640_74#_c_774_n N_A_938_74#_c_1269_n 0.00185769f $X=5.05 $Y=1.765
+ $X2=0 $Y2=0
cc_586 N_A_640_74#_M1006_g N_A_938_74#_c_1269_n 5.58328e-19 $X=5.485 $Y=0.69
+ $X2=0 $Y2=0
cc_587 N_A_640_74#_c_780_n N_A_938_74#_c_1269_n 0.0150779f $X=4.885 $Y=1.515
+ $X2=0 $Y2=0
cc_588 N_A_640_74#_M1000_g N_A_938_74#_c_1270_n 0.0102214f $X=5.05 $Y=0.69 $X2=0
+ $Y2=0
cc_589 N_A_640_74#_M1006_g N_A_938_74#_c_1270_n 0.0116265f $X=5.485 $Y=0.69
+ $X2=0 $Y2=0
cc_590 N_A_640_74#_M1000_g N_A_938_74#_c_1271_n 0.00234788f $X=5.05 $Y=0.69
+ $X2=0 $Y2=0
cc_591 N_A_640_74#_M1006_g N_A_938_74#_c_1280_n 0.00258785f $X=5.485 $Y=0.69
+ $X2=0 $Y2=0
cc_592 N_A_640_74#_M1000_g N_A_938_74#_c_1291_n 4.80353e-19 $X=5.05 $Y=0.69
+ $X2=0 $Y2=0
cc_593 N_A_640_74#_M1006_g N_A_938_74#_c_1291_n 0.00449095f $X=5.485 $Y=0.69
+ $X2=0 $Y2=0
cc_594 N_RESET_B_c_890_n N_VPWR_c_951_n 0.0121096f $X=6 $Y=1.765 $X2=0 $Y2=0
cc_595 N_RESET_B_c_892_n N_VPWR_c_951_n 7.62576e-19 $X=6.5 $Y=1.765 $X2=0 $Y2=0
cc_596 N_RESET_B_c_892_n N_VPWR_c_952_n 0.00979494f $X=6.5 $Y=1.765 $X2=0 $Y2=0
cc_597 N_RESET_B_c_890_n N_VPWR_c_958_n 0.00361294f $X=6 $Y=1.765 $X2=0 $Y2=0
cc_598 N_RESET_B_c_892_n N_VPWR_c_958_n 0.00393873f $X=6.5 $Y=1.765 $X2=0 $Y2=0
cc_599 N_RESET_B_c_890_n N_VPWR_c_947_n 0.00419404f $X=6 $Y=1.765 $X2=0 $Y2=0
cc_600 N_RESET_B_c_892_n N_VPWR_c_947_n 0.00462577f $X=6.5 $Y=1.765 $X2=0 $Y2=0
cc_601 N_RESET_B_c_883_n N_VGND_c_1145_n 0.00642841f $X=5.915 $Y=1.12 $X2=0
+ $Y2=0
cc_602 N_RESET_B_c_885_n N_VGND_c_1145_n 0.00738466f $X=6.345 $Y=1.12 $X2=0
+ $Y2=0
cc_603 N_RESET_B_c_885_n N_VGND_c_1146_n 0.00383152f $X=6.345 $Y=1.12 $X2=0
+ $Y2=0
cc_604 N_RESET_B_c_885_n N_VGND_c_1147_n 0.00579698f $X=6.345 $Y=1.12 $X2=0
+ $Y2=0
cc_605 RESET_B N_VGND_c_1147_n 4.66402e-19 $X=6.395 $Y=1.21 $X2=0 $Y2=0
cc_606 N_RESET_B_c_883_n N_VGND_c_1154_n 0.00383152f $X=5.915 $Y=1.12 $X2=0
+ $Y2=0
cc_607 N_RESET_B_c_883_n N_VGND_c_1162_n 0.00369368f $X=5.915 $Y=1.12 $X2=0
+ $Y2=0
cc_608 N_RESET_B_c_885_n N_VGND_c_1162_n 0.00374269f $X=6.345 $Y=1.12 $X2=0
+ $Y2=0
cc_609 N_RESET_B_c_883_n N_A_938_74#_c_1270_n 7.41618e-19 $X=5.915 $Y=1.12 $X2=0
+ $Y2=0
cc_610 N_RESET_B_c_883_n N_A_938_74#_c_1281_n 0.0102338f $X=5.915 $Y=1.12 $X2=0
+ $Y2=0
cc_611 N_RESET_B_c_885_n N_A_938_74#_c_1281_n 0.00969758f $X=6.345 $Y=1.12 $X2=0
+ $Y2=0
cc_612 RESET_B N_A_938_74#_c_1281_n 0.0365275f $X=6.395 $Y=1.21 $X2=0 $Y2=0
cc_613 N_RESET_B_c_888_n N_A_938_74#_c_1281_n 0.00263297f $X=6.5 $Y=1.285 $X2=0
+ $Y2=0
cc_614 RESET_B N_A_938_74#_c_1272_n 0.0101265f $X=6.395 $Y=1.21 $X2=0 $Y2=0
cc_615 N_RESET_B_c_888_n N_A_938_74#_c_1272_n 0.00334602f $X=6.5 $Y=1.285 $X2=0
+ $Y2=0
cc_616 N_RESET_B_c_885_n N_A_938_74#_c_1273_n 5.59302e-19 $X=6.345 $Y=1.12 $X2=0
+ $Y2=0
cc_617 N_VPWR_c_952_n N_Q_c_1072_n 0.067717f $X=6.81 $Y=2.045 $X2=0 $Y2=0
cc_618 N_VPWR_c_953_n N_Q_c_1072_n 0.0309964f $X=7.76 $Y=2.225 $X2=0 $Y2=0
cc_619 N_VPWR_c_960_n N_Q_c_1072_n 0.0110241f $X=7.595 $Y=3.33 $X2=0 $Y2=0
cc_620 N_VPWR_c_947_n N_Q_c_1072_n 0.00909194f $X=8.88 $Y=3.33 $X2=0 $Y2=0
cc_621 N_VPWR_M1012_s N_Q_c_1073_n 0.00250873f $X=7.56 $Y=1.84 $X2=0 $Y2=0
cc_622 N_VPWR_c_953_n N_Q_c_1073_n 0.0202249f $X=7.76 $Y=2.225 $X2=0 $Y2=0
cc_623 N_VPWR_c_952_n N_Q_c_1074_n 7.28337e-19 $X=6.81 $Y=2.045 $X2=0 $Y2=0
cc_624 N_VPWR_c_953_n N_Q_c_1075_n 0.0323093f $X=7.76 $Y=2.225 $X2=0 $Y2=0
cc_625 N_VPWR_c_955_n N_Q_c_1075_n 0.00158095f $X=8.76 $Y=2.225 $X2=0 $Y2=0
cc_626 N_VPWR_c_964_n N_Q_c_1075_n 0.0146357f $X=8.595 $Y=3.33 $X2=0 $Y2=0
cc_627 N_VPWR_c_947_n N_Q_c_1075_n 0.0121141f $X=8.88 $Y=3.33 $X2=0 $Y2=0
cc_628 N_VPWR_M1014_s N_Q_c_1076_n 0.00393524f $X=8.58 $Y=1.84 $X2=0 $Y2=0
cc_629 N_VPWR_c_955_n N_Q_c_1076_n 0.0247803f $X=8.76 $Y=2.225 $X2=0 $Y2=0
cc_630 N_Q_c_1067_n N_VGND_M1015_s 0.00178571f $X=8.315 $Y=1.005 $X2=0 $Y2=0
cc_631 N_Q_c_1069_n N_VGND_M1029_s 0.00384658f $X=8.765 $Y=1.005 $X2=0 $Y2=0
cc_632 N_Q_c_1065_n N_VGND_c_1147_n 0.0112967f $X=7.515 $Y=0.88 $X2=0 $Y2=0
cc_633 N_Q_c_1066_n N_VGND_c_1147_n 0.0187552f $X=7.55 $Y=0.53 $X2=0 $Y2=0
cc_634 N_Q_c_1066_n N_VGND_c_1148_n 0.0131057f $X=7.55 $Y=0.53 $X2=0 $Y2=0
cc_635 N_Q_c_1067_n N_VGND_c_1148_n 0.0175375f $X=8.315 $Y=1.005 $X2=0 $Y2=0
cc_636 N_Q_c_1068_n N_VGND_c_1148_n 0.0130983f $X=8.41 $Y=0.53 $X2=0 $Y2=0
cc_637 N_Q_c_1068_n N_VGND_c_1150_n 0.0130983f $X=8.41 $Y=0.53 $X2=0 $Y2=0
cc_638 N_Q_c_1069_n N_VGND_c_1150_n 0.0232381f $X=8.765 $Y=1.005 $X2=0 $Y2=0
cc_639 N_Q_c_1066_n N_VGND_c_1155_n 0.0107879f $X=7.55 $Y=0.53 $X2=0 $Y2=0
cc_640 N_Q_c_1068_n N_VGND_c_1156_n 0.00791198f $X=8.41 $Y=0.53 $X2=0 $Y2=0
cc_641 N_Q_c_1066_n N_VGND_c_1162_n 0.00932577f $X=7.55 $Y=0.53 $X2=0 $Y2=0
cc_642 N_Q_c_1068_n N_VGND_c_1162_n 0.00688042f $X=8.41 $Y=0.53 $X2=0 $Y2=0
cc_643 N_VGND_c_1144_n N_A_938_74#_c_1269_n 0.0237374f $X=4.275 $Y=0.58 $X2=0
+ $Y2=0
cc_644 N_VGND_c_1145_n N_A_938_74#_c_1270_n 0.0101043f $X=6.13 $Y=0.515 $X2=0
+ $Y2=0
cc_645 N_VGND_c_1154_n N_A_938_74#_c_1270_n 0.0444371f $X=5.965 $Y=0 $X2=0 $Y2=0
cc_646 N_VGND_c_1162_n N_A_938_74#_c_1270_n 0.0281303f $X=8.88 $Y=0 $X2=0 $Y2=0
cc_647 N_VGND_c_1144_n N_A_938_74#_c_1271_n 0.011925f $X=4.275 $Y=0.58 $X2=0
+ $Y2=0
cc_648 N_VGND_c_1154_n N_A_938_74#_c_1271_n 0.0203379f $X=5.965 $Y=0 $X2=0 $Y2=0
cc_649 N_VGND_c_1162_n N_A_938_74#_c_1271_n 0.0125576f $X=8.88 $Y=0 $X2=0 $Y2=0
cc_650 N_VGND_M1020_d N_A_938_74#_c_1281_n 0.0032758f $X=5.99 $Y=0.37 $X2=0
+ $Y2=0
cc_651 N_VGND_c_1145_n N_A_938_74#_c_1281_n 0.0166614f $X=6.13 $Y=0.515 $X2=0
+ $Y2=0
cc_652 N_VGND_c_1162_n N_A_938_74#_c_1281_n 0.0122318f $X=8.88 $Y=0 $X2=0 $Y2=0
cc_653 N_VGND_c_1147_n N_A_938_74#_c_1272_n 0.0126613f $X=7.12 $Y=0.53 $X2=0
+ $Y2=0
cc_654 N_VGND_c_1145_n N_A_938_74#_c_1273_n 0.0105313f $X=6.13 $Y=0.515 $X2=0
+ $Y2=0
cc_655 N_VGND_c_1146_n N_A_938_74#_c_1273_n 0.0116481f $X=6.955 $Y=0 $X2=0 $Y2=0
cc_656 N_VGND_c_1147_n N_A_938_74#_c_1273_n 0.0276046f $X=7.12 $Y=0.53 $X2=0
+ $Y2=0
cc_657 N_VGND_c_1162_n N_A_938_74#_c_1273_n 0.00951991f $X=8.88 $Y=0 $X2=0 $Y2=0
