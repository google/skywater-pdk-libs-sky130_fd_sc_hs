* File: sky130_fd_sc_hs__sdfrbp_2.pex.spice
* Created: Thu Aug 27 21:08:27 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HS__SDFRBP_2%A_27_79# 1 2 9 11 13 14 17 20 23 27 30 34
+ 37 38
c83 30 0 1.3813e-19 $X=2.275 $Y=2.405
r84 34 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.44
+ $Y=1.995 $X2=2.44 $Y2=1.995
r85 32 34 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=2.44 $Y=2.32
+ $X2=2.44 $Y2=1.995
r86 31 38 2.76166 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.445 $Y=2.405
+ $X2=0.28 $Y2=2.405
r87 30 32 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.275 $Y=2.405
+ $X2=2.44 $Y2=2.32
r88 30 31 119.39 $w=1.68e-07 $l=1.83e-06 $layer=LI1_cond $X=2.275 $Y=2.405
+ $X2=0.445 $Y2=2.405
r89 27 28 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.23
+ $Y=1.415 $X2=1.23 $Y2=1.415
r90 25 37 0.221902 $w=3.3e-07 $l=1.25e-07 $layer=LI1_cond $X=0.365 $Y=1.415
+ $X2=0.24 $Y2=1.415
r91 25 27 30.208 $w=3.28e-07 $l=8.65e-07 $layer=LI1_cond $X=0.365 $Y=1.415
+ $X2=1.23 $Y2=1.415
r92 21 38 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.28 $Y=2.49 $X2=0.28
+ $Y2=2.405
r93 21 23 5.5876 $w=3.28e-07 $l=1.6e-07 $layer=LI1_cond $X=0.28 $Y=2.49 $X2=0.28
+ $Y2=2.65
r94 20 38 3.70735 $w=2.5e-07 $l=1.18427e-07 $layer=LI1_cond $X=0.2 $Y=2.32
+ $X2=0.28 $Y2=2.405
r95 19 37 7.38875 $w=2.1e-07 $l=1.83916e-07 $layer=LI1_cond $X=0.2 $Y=1.58
+ $X2=0.24 $Y2=1.415
r96 19 20 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=0.2 $Y=1.58 $X2=0.2
+ $Y2=2.32
r97 15 37 7.38875 $w=2.1e-07 $l=1.65e-07 $layer=LI1_cond $X=0.24 $Y=1.25
+ $X2=0.24 $Y2=1.415
r98 15 17 29.733 $w=2.48e-07 $l=6.45e-07 $layer=LI1_cond $X=0.24 $Y=1.25
+ $X2=0.24 $Y2=0.605
r99 14 28 29.7264 $w=3.3e-07 $l=1.7e-07 $layer=POLY_cond $X=1.4 $Y=1.415
+ $X2=1.23 $Y2=1.415
r100 11 35 50.023 $w=3.78e-07 $l=3.06186e-07 $layer=POLY_cond $X=2.615 $Y=2.245
+ $X2=2.49 $Y2=1.995
r101 11 13 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=2.615 $Y=2.245
+ $X2=2.615 $Y2=2.64
r102 7 14 32.1775 $w=3.3e-07 $l=1.98997e-07 $layer=POLY_cond $X=1.475 $Y=1.25
+ $X2=1.4 $Y2=1.415
r103 7 9 330.734 $w=1.5e-07 $l=6.45e-07 $layer=POLY_cond $X=1.475 $Y=1.25
+ $X2=1.475 $Y2=0.605
r104 2 23 600 $w=1.7e-07 $l=3.95917e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.32 $X2=0.28 $Y2=2.65
r105 1 17 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.395 $X2=0.28 $Y2=0.605
.ends

.subckt PM_SKY130_FD_SC_HS__SDFRBP_2%SCE 2 3 5 6 8 9 11 14 18 23 24 26 27 29 30
+ 31 36 46
r86 41 42 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.385
+ $Y=1.985 $X2=1.385 $Y2=1.985
r87 36 41 12.5952 $w=3.3e-07 $l=1.11041e-07 $layer=POLY_cond $X=1.37 $Y=1.985
+ $X2=1.46 $Y2=2.032
r88 36 38 116.283 $w=3.3e-07 $l=6.65e-07 $layer=POLY_cond $X=1.37 $Y=1.985
+ $X2=0.705 $Y2=1.985
r89 31 46 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.71 $Y=1.985
+ $X2=1.625 $Y2=1.985
r90 31 46 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=1.61 $Y=1.985
+ $X2=1.625 $Y2=1.985
r91 31 42 7.85757 $w=3.28e-07 $l=2.25e-07 $layer=LI1_cond $X=1.61 $Y=1.985
+ $X2=1.385 $Y2=1.985
r92 30 42 6.46067 $w=3.28e-07 $l=1.85e-07 $layer=LI1_cond $X=1.2 $Y=1.985
+ $X2=1.385 $Y2=1.985
r93 29 30 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=0.705 $Y=1.985
+ $X2=1.2 $Y2=1.985
r94 29 38 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=0.705
+ $Y=1.985 $X2=0.705 $Y2=1.985
r95 27 44 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.57 $Y=1.455
+ $X2=2.57 $Y2=1.29
r96 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.57
+ $Y=1.455 $X2=2.57 $Y2=1.455
r97 24 26 34.3517 $w=2.58e-07 $l=7.75e-07 $layer=LI1_cond $X=1.795 $Y=1.49
+ $X2=2.57 $Y2=1.49
r98 23 31 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.71 $Y=1.82
+ $X2=1.71 $Y2=1.985
r99 22 24 7.21222 $w=2.6e-07 $l=1.67183e-07 $layer=LI1_cond $X=1.71 $Y=1.62
+ $X2=1.795 $Y2=1.49
r100 22 23 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=1.71 $Y=1.62 $X2=1.71
+ $Y2=1.82
r101 21 38 19.2347 $w=3.3e-07 $l=1.1e-07 $layer=POLY_cond $X=0.595 $Y=1.985
+ $X2=0.705 $Y2=1.985
r102 16 18 43.5851 $w=1.5e-07 $l=8.5e-08 $layer=POLY_cond $X=0.41 $Y=0.965
+ $X2=0.495 $Y2=0.965
r103 14 44 351.245 $w=1.5e-07 $l=6.85e-07 $layer=POLY_cond $X=2.66 $Y=0.605
+ $X2=2.66 $Y2=1.29
r104 9 41 19.5823 $w=1.5e-07 $l=2.13e-07 $layer=POLY_cond $X=1.46 $Y=2.245
+ $X2=1.46 $Y2=2.032
r105 9 11 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=1.46 $Y=2.245
+ $X2=1.46 $Y2=2.64
r106 6 21 64.077 $w=2.08e-07 $l=2.79285e-07 $layer=POLY_cond $X=0.505 $Y=2.245
+ $X2=0.465 $Y2=1.985
r107 6 8 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=0.505 $Y=2.245
+ $X2=0.505 $Y2=2.64
r108 3 18 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.495 $Y=0.89
+ $X2=0.495 $Y2=0.965
r109 3 5 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=0.495 $Y=0.89
+ $X2=0.495 $Y2=0.605
r110 2 21 42.0626 $w=2.08e-07 $l=1.90526e-07 $layer=POLY_cond $X=0.41 $Y=1.82
+ $X2=0.465 $Y2=1.985
r111 1 16 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.41 $Y=1.04
+ $X2=0.41 $Y2=0.965
r112 1 2 399.957 $w=1.5e-07 $l=7.8e-07 $layer=POLY_cond $X=0.41 $Y=1.04 $X2=0.41
+ $Y2=1.82
.ends

.subckt PM_SKY130_FD_SC_HS__SDFRBP_2%D 3 5 6 8 9 12 13 14
r47 12 15 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.925 $Y=1.09
+ $X2=1.925 $Y2=1.255
r48 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.925 $Y=1.09
+ $X2=1.925 $Y2=0.925
r49 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.925
+ $Y=1.09 $X2=1.925 $Y2=1.09
r50 9 13 7.43022 $w=3.78e-07 $l=2.45e-07 $layer=LI1_cond $X=1.68 $Y=1 $X2=1.925
+ $Y2=1
r51 6 8 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=1.88 $Y=2.245
+ $X2=1.88 $Y2=2.64
r52 5 6 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=1.88 $Y=2.155 $X2=1.88
+ $Y2=2.245
r53 5 15 349.839 $w=1.8e-07 $l=9e-07 $layer=POLY_cond $X=1.88 $Y=2.155 $X2=1.88
+ $Y2=1.255
r54 3 14 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.865 $Y=0.605
+ $X2=1.865 $Y2=0.925
.ends

.subckt PM_SKY130_FD_SC_HS__SDFRBP_2%SCD 1 3 6 10 11 12 16
c44 11 0 1.2788e-19 $X=3.12 $Y=1.665
c45 1 0 2.38726e-19 $X=3.035 $Y=2.245
r46 11 12 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=3.11 $Y=1.605
+ $X2=3.11 $Y2=2.035
r47 11 16 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.11
+ $Y=1.605 $X2=3.11 $Y2=1.605
r48 10 16 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=3.11 $Y=1.945
+ $X2=3.11 $Y2=1.605
r49 9 16 41.8716 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.11 $Y=1.44
+ $X2=3.11 $Y2=1.605
r50 6 9 428.16 $w=1.5e-07 $l=8.35e-07 $layer=POLY_cond $X=3.05 $Y=0.605 $X2=3.05
+ $Y2=1.44
r51 1 10 55.1908 $w=2.62e-07 $l=3.3541e-07 $layer=POLY_cond $X=3.035 $Y=2.245
+ $X2=3.11 $Y2=1.945
r52 1 3 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=3.035 $Y=2.245
+ $X2=3.035 $Y2=2.64
.ends

.subckt PM_SKY130_FD_SC_HS__SDFRBP_2%RESET_B 3 5 7 8 10 11 12 13 15 17 20 23 24
+ 26 29 31 32 33 34 42 45 48 50 53 64
c190 64 0 1.25229e-19 $X=10.8 $Y=2.035
c191 45 0 1.2788e-19 $X=3.605 $Y=2.032
r192 55 64 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.945
+ $Y=1.985 $X2=10.945 $Y2=1.985
r193 52 53 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.825
+ $Y=1.96 $X2=7.825 $Y2=1.96
r194 50 52 14.7051 $w=2.95e-07 $l=9e-08 $layer=POLY_cond $X=7.735 $Y=2.002
+ $X2=7.825 $Y2=2.002
r195 47 48 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.95
+ $Y=1.985 $X2=3.95 $Y2=1.985
r196 45 47 46.4497 $w=3.58e-07 $l=3.45e-07 $layer=POLY_cond $X=3.605 $Y=2.032
+ $X2=3.95 $Y2=2.032
r197 44 45 2.01955 $w=3.58e-07 $l=1.5e-08 $layer=POLY_cond $X=3.59 $Y=2.032
+ $X2=3.605 $Y2=2.032
r198 42 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.8 $Y=2.035
+ $X2=10.8 $Y2=2.035
r199 40 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=2.035
+ $X2=7.92 $Y2=2.035
r200 36 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=2.035
+ $X2=4.08 $Y2=2.035
r201 34 40 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=8.065 $Y=2.035
+ $X2=7.92 $Y2=2.035
r202 33 42 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=10.655 $Y=2.035
+ $X2=10.8 $Y2=2.035
r203 33 34 3.20544 $w=1.4e-07 $l=2.59e-06 $layer=MET1_cond $X=10.655 $Y=2.035
+ $X2=8.065 $Y2=2.035
r204 32 36 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.225 $Y=2.035
+ $X2=4.08 $Y2=2.035
r205 31 40 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=7.775 $Y=2.035
+ $X2=7.92 $Y2=2.035
r206 31 32 4.39356 $w=1.4e-07 $l=3.55e-06 $layer=MET1_cond $X=7.775 $Y=2.035
+ $X2=4.225 $Y2=2.035
r207 27 29 71.7872 $w=1.5e-07 $l=1.4e-07 $layer=POLY_cond $X=10.715 $Y=1.55
+ $X2=10.855 $Y2=1.55
r208 24 55 60.4771 $w=2.87e-07 $l=3.23612e-07 $layer=POLY_cond $X=11.005 $Y=2.28
+ $X2=10.945 $Y2=1.985
r209 24 26 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=11.005 $Y=2.28
+ $X2=11.005 $Y2=2.565
r210 23 55 38.6443 $w=2.87e-07 $l=2.05122e-07 $layer=POLY_cond $X=10.855 $Y=1.82
+ $X2=10.945 $Y2=1.985
r211 22 29 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=10.855 $Y=1.625
+ $X2=10.855 $Y2=1.55
r212 22 23 99.9894 $w=1.5e-07 $l=1.95e-07 $layer=POLY_cond $X=10.855 $Y=1.625
+ $X2=10.855 $Y2=1.82
r213 18 27 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=10.715 $Y=1.475
+ $X2=10.715 $Y2=1.55
r214 18 20 458.926 $w=1.5e-07 $l=8.95e-07 $layer=POLY_cond $X=10.715 $Y=1.475
+ $X2=10.715 $Y2=0.58
r215 17 50 18.5736 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=7.735 $Y=1.795
+ $X2=7.735 $Y2=2.002
r216 16 17 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=7.735 $Y=1.235
+ $X2=7.735 $Y2=1.795
r217 13 50 34.3119 $w=2.95e-07 $l=2.96277e-07 $layer=POLY_cond $X=7.525 $Y=2.21
+ $X2=7.735 $Y2=2.002
r218 13 15 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=7.525 $Y=2.21
+ $X2=7.525 $Y2=2.495
r219 11 16 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=7.66 $Y=1.16
+ $X2=7.735 $Y2=1.235
r220 11 12 135.883 $w=1.5e-07 $l=2.65e-07 $layer=POLY_cond $X=7.66 $Y=1.16
+ $X2=7.395 $Y2=1.16
r221 8 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=7.32 $Y=1.085
+ $X2=7.395 $Y2=1.16
r222 8 10 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=7.32 $Y=1.085
+ $X2=7.32 $Y2=0.8
r223 5 45 23.1716 $w=1.5e-07 $l=2.13e-07 $layer=POLY_cond $X=3.605 $Y=2.245
+ $X2=3.605 $Y2=2.032
r224 5 7 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=3.605 $Y=2.245
+ $X2=3.605 $Y2=2.64
r225 1 44 23.1716 $w=1.5e-07 $l=2.12e-07 $layer=POLY_cond $X=3.59 $Y=1.82
+ $X2=3.59 $Y2=2.032
r226 1 3 623.011 $w=1.5e-07 $l=1.215e-06 $layer=POLY_cond $X=3.59 $Y=1.82
+ $X2=3.59 $Y2=0.605
.ends

.subckt PM_SKY130_FD_SC_HS__SDFRBP_2%CLK 1 3 4 6 8 9
c52 1 0 1.25894e-19 $X=4.62 $Y=1.22
r53 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.07
+ $Y=1.385 $X2=4.07 $Y2=1.385
r54 9 13 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=4.07 $Y=1.295 $X2=4.07
+ $Y2=1.385
r55 8 12 83.0591 $w=3.3e-07 $l=4.75e-07 $layer=POLY_cond $X=4.545 $Y=1.385
+ $X2=4.07 $Y2=1.385
r56 4 8 100.419 $w=1.86e-07 $l=3.82492e-07 $layer=POLY_cond $X=4.645 $Y=1.765
+ $X2=4.64 $Y2=1.385
r57 4 6 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=4.645 $Y=1.765
+ $X2=4.645 $Y2=2.4
r58 1 8 44.7042 $w=1.86e-07 $l=1.74714e-07 $layer=POLY_cond $X=4.62 $Y=1.22
+ $X2=4.64 $Y2=1.385
r59 1 3 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=4.62 $Y=1.22 $X2=4.62
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HS__SDFRBP_2%A_1025_74# 1 2 8 9 11 12 16 18 20 21 22 23
+ 25 29 30 31 33 34 36 39 42 43 44 46 51 56 63 64 67 69 71
c204 64 0 3.17494e-19 $X=9.475 $Y=1.07
c205 63 0 2.9567e-20 $X=9.475 $Y=1.07
c206 51 0 1.25894e-19 $X=5.56 $Y=1.075
c207 39 0 2.30857e-19 $X=8.155 $Y=0.665
c208 33 0 5.66018e-20 $X=5.56 $Y=1.5
c209 16 0 6.36741e-20 $X=6.54 $Y=0.8
r210 67 69 5.06676 $w=4.43e-07 $l=1.65e-07 $layer=LI1_cond $X=9.532 $Y=2.03
+ $X2=9.532 $Y2=1.865
r211 67 68 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.615
+ $Y=2.03 $X2=9.615 $Y2=2.03
r212 64 77 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=9.475 $Y=1.07
+ $X2=9.475 $Y2=1.16
r213 63 64 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.475
+ $Y=1.07 $X2=9.475 $Y2=1.07
r214 60 63 10.1275 $w=3.28e-07 $l=2.9e-07 $layer=LI1_cond $X=9.185 $Y=1.07
+ $X2=9.475 $Y2=1.07
r215 56 58 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=7.085 $Y=0.395
+ $X2=7.085 $Y2=0.665
r216 47 63 0.716491 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=9.475 $Y=1.235
+ $X2=9.475 $Y2=1.07
r217 47 69 22.0012 $w=3.28e-07 $l=6.3e-07 $layer=LI1_cond $X=9.475 $Y=1.235
+ $X2=9.475 $Y2=1.865
r218 46 60 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.185 $Y=0.905
+ $X2=9.185 $Y2=1.07
r219 45 46 31.3155 $w=1.68e-07 $l=4.8e-07 $layer=LI1_cond $X=9.185 $Y=0.425
+ $X2=9.185 $Y2=0.905
r220 43 45 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.1 $Y=0.34
+ $X2=9.185 $Y2=0.425
r221 43 44 50.5615 $w=1.68e-07 $l=7.75e-07 $layer=LI1_cond $X=9.1 $Y=0.34
+ $X2=8.325 $Y2=0.34
r222 41 44 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.24 $Y=0.425
+ $X2=8.325 $Y2=0.34
r223 41 42 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=8.24 $Y=0.425
+ $X2=8.24 $Y2=0.58
r224 40 58 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.17 $Y=0.665
+ $X2=7.085 $Y2=0.665
r225 39 42 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.155 $Y=0.665
+ $X2=8.24 $Y2=0.58
r226 39 40 64.262 $w=1.68e-07 $l=9.85e-07 $layer=LI1_cond $X=8.155 $Y=0.665
+ $X2=7.17 $Y2=0.665
r227 37 74 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.045 $Y=1.665
+ $X2=6.045 $Y2=1.83
r228 37 71 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=6.045 $Y=1.665
+ $X2=6.045 $Y2=1.575
r229 36 37 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.045
+ $Y=1.665 $X2=6.045 $Y2=1.665
r230 34 55 12.2 $w=3.3e-07 $l=4.35603e-07 $layer=LI1_cond $X=5.645 $Y=1.665
+ $X2=5.4 $Y2=1.995
r231 34 36 13.969 $w=3.28e-07 $l=4e-07 $layer=LI1_cond $X=5.645 $Y=1.665
+ $X2=6.045 $Y2=1.665
r232 33 34 8.95823 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=5.56 $Y=1.5
+ $X2=5.645 $Y2=1.665
r233 32 51 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.56 $Y=1.16
+ $X2=5.56 $Y2=1.075
r234 32 33 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=5.56 $Y=1.16
+ $X2=5.56 $Y2=1.5
r235 30 56 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7 $Y=0.395
+ $X2=7.085 $Y2=0.395
r236 30 31 102.428 $w=1.68e-07 $l=1.57e-06 $layer=LI1_cond $X=7 $Y=0.395
+ $X2=5.43 $Y2=0.395
r237 27 51 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=5.265 $Y=1.075
+ $X2=5.56 $Y2=1.075
r238 27 29 16.5882 $w=3.28e-07 $l=4.75e-07 $layer=LI1_cond $X=5.265 $Y=0.99
+ $X2=5.265 $Y2=0.515
r239 26 31 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=5.265 $Y=0.48
+ $X2=5.43 $Y2=0.395
r240 26 29 1.22229 $w=3.28e-07 $l=3.5e-08 $layer=LI1_cond $X=5.265 $Y=0.48
+ $X2=5.265 $Y2=0.515
r241 23 68 51.8789 $w=3.07e-07 $l=2.87228e-07 $layer=POLY_cond $X=9.7 $Y=2.28
+ $X2=9.62 $Y2=2.03
r242 23 25 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=9.7 $Y=2.28 $X2=9.7
+ $Y2=2.565
r243 21 77 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.31 $Y=1.16
+ $X2=9.475 $Y2=1.16
r244 21 22 184.596 $w=1.5e-07 $l=3.6e-07 $layer=POLY_cond $X=9.31 $Y=1.16
+ $X2=8.95 $Y2=1.16
r245 18 22 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=8.875 $Y=1.085
+ $X2=8.95 $Y2=1.16
r246 18 20 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=8.875 $Y=1.085
+ $X2=8.875 $Y2=0.69
r247 14 16 358.936 $w=1.5e-07 $l=7e-07 $layer=POLY_cond $X=6.54 $Y=1.5 $X2=6.54
+ $Y2=0.8
r248 13 71 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.21 $Y=1.575
+ $X2=6.045 $Y2=1.575
r249 12 14 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=6.465 $Y=1.575
+ $X2=6.54 $Y2=1.5
r250 12 13 130.755 $w=1.5e-07 $l=2.55e-07 $layer=POLY_cond $X=6.465 $Y=1.575
+ $X2=6.21 $Y2=1.575
r251 9 11 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=6.1 $Y=2.21 $X2=6.1
+ $Y2=2.495
r252 8 9 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=6.1 $Y=2.12 $X2=6.1
+ $Y2=2.21
r253 8 74 112.726 $w=1.8e-07 $l=2.9e-07 $layer=POLY_cond $X=6.1 $Y=2.12 $X2=6.1
+ $Y2=1.83
r254 2 55 600 $w=1.7e-07 $l=2.17428e-07 $layer=licon1_PDIFF $count=1 $X=5.17
+ $Y=1.84 $X2=5.32 $Y2=1.995
r255 1 29 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=5.125
+ $Y=0.37 $X2=5.265 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__SDFRBP_2%A_1370_289# 1 2 8 11 13 15 18 19 22 23 25
+ 33 34 36
c97 34 0 1.87681e-19 $X=8.845 $Y=0.842
c98 22 0 6.36741e-20 $X=7.21 $Y=1.005
c99 19 0 8.03528e-20 $X=7.105 $Y=1.61
c100 11 0 1.82451e-19 $X=6.93 $Y=0.8
r101 37 39 1.74861 $w=3.3e-07 $l=1e-08 $layer=POLY_cond $X=6.93 $Y=1.61 $X2=6.94
+ $Y2=1.61
r102 32 34 4.47019 $w=4.93e-07 $l=1.85e-07 $layer=LI1_cond $X=8.66 $Y=0.842
+ $X2=8.845 $Y2=0.842
r103 32 33 9.48656 $w=4.93e-07 $l=1.65e-07 $layer=LI1_cond $X=8.66 $Y=0.842
+ $X2=8.495 $Y2=0.842
r104 29 34 7.09362 $w=1.7e-07 $l=2.48e-07 $layer=LI1_cond $X=8.845 $Y=1.09
+ $X2=8.845 $Y2=0.842
r105 29 36 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=8.845 $Y=1.09
+ $X2=8.845 $Y2=1.745
r106 25 27 27.0228 $w=2.88e-07 $l=6.8e-07 $layer=LI1_cond $X=8.785 $Y=1.91
+ $X2=8.785 $Y2=2.59
r107 23 36 7.71909 $w=2.88e-07 $l=1.45e-07 $layer=LI1_cond $X=8.785 $Y=1.89
+ $X2=8.785 $Y2=1.745
r108 23 25 0.794788 $w=2.88e-07 $l=2e-08 $layer=LI1_cond $X=8.785 $Y=1.89
+ $X2=8.785 $Y2=1.91
r109 22 33 83.8342 $w=1.68e-07 $l=1.285e-06 $layer=LI1_cond $X=7.21 $Y=1.005
+ $X2=8.495 $Y2=1.005
r110 19 39 28.8521 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=7.105 $Y=1.61
+ $X2=6.94 $Y2=1.61
r111 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.105
+ $Y=1.61 $X2=7.105 $Y2=1.61
r112 16 22 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=7.105 $Y=1.09
+ $X2=7.21 $Y2=1.005
r113 16 18 27.4632 $w=2.08e-07 $l=5.2e-07 $layer=LI1_cond $X=7.105 $Y=1.09
+ $X2=7.105 $Y2=1.61
r114 13 15 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=6.94 $Y=2.21
+ $X2=6.94 $Y2=2.495
r115 9 37 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.93 $Y=1.445
+ $X2=6.93 $Y2=1.61
r116 9 11 330.734 $w=1.5e-07 $l=6.45e-07 $layer=POLY_cond $X=6.93 $Y=1.445
+ $X2=6.93 $Y2=0.8
r117 8 13 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=6.94 $Y=2.12 $X2=6.94
+ $Y2=2.21
r118 7 39 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=6.94 $Y=1.775
+ $X2=6.94 $Y2=1.61
r119 7 8 134.105 $w=1.8e-07 $l=3.45e-07 $layer=POLY_cond $X=6.94 $Y=1.775
+ $X2=6.94 $Y2=2.12
r120 2 27 400 $w=1.7e-07 $l=9.26971e-07 $layer=licon1_PDIFF $count=1 $X=8.575
+ $Y=1.735 $X2=8.725 $Y2=2.59
r121 2 25 400 $w=1.7e-07 $l=2.38485e-07 $layer=licon1_PDIFF $count=1 $X=8.575
+ $Y=1.735 $X2=8.725 $Y2=1.91
r122 1 32 182 $w=1.7e-07 $l=5.05173e-07 $layer=licon1_NDIFF $count=1 $X=8.52
+ $Y=0.37 $X2=8.66 $Y2=0.81
.ends

.subckt PM_SKY130_FD_SC_HS__SDFRBP_2%A_1223_118# 1 2 3 12 14 16 17 22 23 24 26
+ 27 29
c104 29 0 1.03439e-19 $X=8.425 $Y=1.41
c105 12 0 2.9567e-20 $X=8.445 $Y=0.69
r106 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.425
+ $Y=1.41 $X2=8.425 $Y2=1.41
r107 27 29 32.0123 $w=3.13e-07 $l=8.75e-07 $layer=LI1_cond $X=7.55 $Y=1.417
+ $X2=8.425 $Y2=1.417
r108 26 37 10.3482 $w=3.36e-07 $l=3.72552e-07 $layer=LI1_cond $X=7.465 $Y=2.32
+ $X2=7.75 $Y2=2.522
r109 25 27 7.64049 $w=3.15e-07 $l=1.95944e-07 $layer=LI1_cond $X=7.465 $Y=1.575
+ $X2=7.55 $Y2=1.417
r110 25 26 48.6043 $w=1.68e-07 $l=7.45e-07 $layer=LI1_cond $X=7.465 $Y=1.575
+ $X2=7.465 $Y2=2.32
r111 23 26 6.05874 $w=3.36e-07 $l=1.41244e-07 $layer=LI1_cond $X=7.38 $Y=2.425
+ $X2=7.465 $Y2=2.32
r112 23 24 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=7.38 $Y=2.425
+ $X2=6.83 $Y2=2.425
r113 22 24 6.00066 $w=3.3e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.745 $Y=2.34
+ $X2=6.83 $Y2=2.425
r114 22 33 15.5273 $w=3.3e-07 $l=5.06991e-07 $layer=LI1_cond $X=6.745 $Y=2.34
+ $X2=6.325 $Y2=2.532
r115 21 22 90.6845 $w=1.68e-07 $l=1.39e-06 $layer=LI1_cond $X=6.745 $Y=0.95
+ $X2=6.745 $Y2=2.34
r116 17 21 7.51767 $w=3e-07 $l=1.8775e-07 $layer=LI1_cond $X=6.66 $Y=0.8
+ $X2=6.745 $Y2=0.95
r117 17 19 12.8689 $w=2.98e-07 $l=3.35e-07 $layer=LI1_cond $X=6.66 $Y=0.8
+ $X2=6.325 $Y2=0.8
r118 14 30 52.2586 $w=2.99e-07 $l=2.85044e-07 $layer=POLY_cond $X=8.5 $Y=1.66
+ $X2=8.425 $Y2=1.41
r119 14 16 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=8.5 $Y=1.66
+ $X2=8.5 $Y2=2.235
r120 10 30 38.5562 $w=2.99e-07 $l=1.74714e-07 $layer=POLY_cond $X=8.445 $Y=1.245
+ $X2=8.425 $Y2=1.41
r121 10 12 284.585 $w=1.5e-07 $l=5.55e-07 $layer=POLY_cond $X=8.445 $Y=1.245
+ $X2=8.445 $Y2=0.69
r122 3 37 600 $w=1.7e-07 $l=3.00791e-07 $layer=licon1_PDIFF $count=1 $X=7.6
+ $Y=2.285 $X2=7.75 $Y2=2.52
r123 2 33 600 $w=1.7e-07 $l=3.11087e-07 $layer=licon1_PDIFF $count=1 $X=6.175
+ $Y=2.285 $X2=6.325 $Y2=2.53
r124 1 19 182 $w=1.7e-07 $l=2.96985e-07 $layer=licon1_NDIFF $count=1 $X=6.115
+ $Y=0.59 $X2=6.325 $Y2=0.8
.ends

.subckt PM_SKY130_FD_SC_HS__SDFRBP_2%A_852_74# 1 2 9 11 13 14 17 18 20 21 22 24
+ 25 26 27 29 30 32 33 37 38 39 42 44 48 51 54 56 57 60 61 62 68 70
c194 61 0 1.55498e-19 $X=4.407 $Y=1.01
c195 39 0 1.3138e-19 $X=9.04 $Y=1.55
c196 38 0 1.34905e-19 $X=9.85 $Y=1.55
c197 17 0 5.24149e-20 $X=5.595 $Y=3.075
c198 11 0 5.66018e-20 $X=5.095 $Y=1.765
c199 9 0 3.89357e-20 $X=5.05 $Y=0.74
r200 71 73 14.8055 $w=2.93e-07 $l=9e-08 $layer=POLY_cond $X=5.14 $Y=1.495
+ $X2=5.14 $Y2=1.405
r201 70 71 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.14
+ $Y=1.495 $X2=5.14 $Y2=1.495
r202 67 70 8.3814 $w=3.28e-07 $l=2.4e-07 $layer=LI1_cond $X=4.9 $Y=1.495
+ $X2=5.14 $Y2=1.495
r203 67 68 5.66838 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=4.9 $Y=1.495
+ $X2=4.815 $Y2=1.495
r204 62 65 4.37928 $w=2.48e-07 $l=9.5e-08 $layer=LI1_cond $X=4.46 $Y=1.905
+ $X2=4.46 $Y2=2
r205 59 67 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.9 $Y=1.66 $X2=4.9
+ $Y2=1.495
r206 59 60 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=4.9 $Y=1.66 $X2=4.9
+ $Y2=1.82
r207 58 62 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.585 $Y=1.905
+ $X2=4.46 $Y2=1.905
r208 57 60 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.815 $Y=1.905
+ $X2=4.9 $Y2=1.82
r209 57 58 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=4.815 $Y=1.905
+ $X2=4.585 $Y2=1.905
r210 56 68 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=4.575 $Y=1.415
+ $X2=4.815 $Y2=1.415
r211 54 56 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.49 $Y=1.33
+ $X2=4.575 $Y2=1.415
r212 54 61 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=4.49 $Y=1.33
+ $X2=4.49 $Y2=1.01
r213 49 61 8.53494 $w=3.33e-07 $l=1.67e-07 $layer=LI1_cond $X=4.407 $Y=0.843
+ $X2=4.407 $Y2=1.01
r214 49 51 11.2836 $w=3.33e-07 $l=3.28e-07 $layer=LI1_cond $X=4.407 $Y=0.843
+ $X2=4.407 $Y2=0.515
r215 46 47 31.303 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=5.58 $Y=1.405
+ $X2=5.58 $Y2=1.48
r216 44 46 85.5161 $w=1.8e-07 $l=2.2e-07 $layer=POLY_cond $X=5.58 $Y=1.185
+ $X2=5.58 $Y2=1.405
r217 40 42 458.926 $w=1.5e-07 $l=8.95e-07 $layer=POLY_cond $X=9.925 $Y=1.475
+ $X2=9.925 $Y2=0.58
r218 38 40 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=9.85 $Y=1.55
+ $X2=9.925 $Y2=1.475
r219 38 39 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=9.85 $Y=1.55
+ $X2=9.04 $Y2=1.55
r220 35 37 294.84 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=8.95 $Y=2.81
+ $X2=8.95 $Y2=2.235
r221 34 39 26.9307 $w=1.5e-07 $l=1.48324e-07 $layer=POLY_cond $X=8.95 $Y=1.66
+ $X2=9.04 $Y2=1.55
r222 34 37 294.84 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=8.95 $Y=1.66
+ $X2=8.95 $Y2=2.235
r223 32 35 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=8.95 $Y=2.9 $X2=8.95
+ $Y2=2.81
r224 32 33 68.0242 $w=1.8e-07 $l=1.75e-07 $layer=POLY_cond $X=8.95 $Y=2.9
+ $X2=8.95 $Y2=3.075
r225 31 48 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=6.64 $Y=3.15 $X2=6.55
+ $Y2=3.15
r226 30 33 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=8.86 $Y=3.15
+ $X2=8.95 $Y2=3.075
r227 30 31 1138.34 $w=1.5e-07 $l=2.22e-06 $layer=POLY_cond $X=8.86 $Y=3.15
+ $X2=6.64 $Y2=3.15
r228 27 29 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=6.55 $Y=2.78
+ $X2=6.55 $Y2=2.495
r229 26 48 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=6.55 $Y=3.075
+ $X2=6.55 $Y2=3.15
r230 25 27 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=6.55 $Y=2.87 $X2=6.55
+ $Y2=2.78
r231 25 26 79.6855 $w=1.8e-07 $l=2.05e-07 $layer=POLY_cond $X=6.55 $Y=2.87
+ $X2=6.55 $Y2=3.075
r232 22 24 99.6133 $w=1.5e-07 $l=3.1e-07 $layer=POLY_cond $X=6.04 $Y=1.11
+ $X2=6.04 $Y2=0.8
r233 20 48 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=6.46 $Y=3.15 $X2=6.55
+ $Y2=3.15
r234 20 21 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=6.46 $Y=3.15
+ $X2=5.67 $Y2=3.15
r235 19 44 7.1379 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=5.67 $Y=1.185 $X2=5.58
+ $Y2=1.185
r236 18 22 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.965 $Y=1.185
+ $X2=6.04 $Y2=1.11
r237 18 19 151.266 $w=1.5e-07 $l=2.95e-07 $layer=POLY_cond $X=5.965 $Y=1.185
+ $X2=5.67 $Y2=1.185
r238 17 21 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.595 $Y=3.075
+ $X2=5.67 $Y2=3.15
r239 17 47 817.862 $w=1.5e-07 $l=1.595e-06 $layer=POLY_cond $X=5.595 $Y=3.075
+ $X2=5.595 $Y2=1.48
r240 15 73 18.414 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.305 $Y=1.405
+ $X2=5.14 $Y2=1.405
r241 14 46 7.1379 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=5.49 $Y=1.405 $X2=5.58
+ $Y2=1.405
r242 14 15 94.8617 $w=1.5e-07 $l=1.85e-07 $layer=POLY_cond $X=5.49 $Y=1.405
+ $X2=5.305 $Y2=1.405
r243 11 71 55.8646 $w=2.93e-07 $l=2.91633e-07 $layer=POLY_cond $X=5.095 $Y=1.765
+ $X2=5.14 $Y2=1.495
r244 11 13 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=5.095 $Y=1.765
+ $X2=5.095 $Y2=2.4
r245 7 73 23.7861 $w=2.93e-07 $l=1.21861e-07 $layer=POLY_cond $X=5.05 $Y=1.33
+ $X2=5.14 $Y2=1.405
r246 7 9 302.532 $w=1.5e-07 $l=5.9e-07 $layer=POLY_cond $X=5.05 $Y=1.33 $X2=5.05
+ $Y2=0.74
r247 2 65 600 $w=1.7e-07 $l=2.20907e-07 $layer=licon1_PDIFF $count=1 $X=4.275
+ $Y=1.84 $X2=4.42 $Y2=2
r248 1 51 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=4.26
+ $Y=0.37 $X2=4.405 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__SDFRBP_2%A_2006_373# 1 2 7 9 12 17 19 20 21 22 25 27
+ 28 30 31 37
c110 21 0 3.10546e-20 $X=11.065 $Y=2.405
c111 20 0 1.34905e-19 $X=10.545 $Y=1.565
c112 12 0 1.25229e-19 $X=10.285 $Y=0.58
r113 36 37 22.2151 $w=3.58e-07 $l=1.65e-07 $layer=POLY_cond $X=10.12 $Y=2.072
+ $X2=10.285 $Y2=2.072
r114 31 34 5.5876 $w=3.28e-07 $l=1.6e-07 $layer=LI1_cond $X=11.23 $Y=2.405
+ $X2=11.23 $Y2=2.565
r115 29 30 39.4706 $w=1.68e-07 $l=6.05e-07 $layer=LI1_cond $X=11.775 $Y=0.875
+ $X2=11.775 $Y2=1.48
r116 27 29 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=11.69 $Y=0.79
+ $X2=11.775 $Y2=0.875
r117 27 28 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=11.69 $Y=0.79
+ $X2=11.455 $Y2=0.79
r118 23 28 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=11.29 $Y=0.705
+ $X2=11.455 $Y2=0.79
r119 23 25 4.36531 $w=3.28e-07 $l=1.25e-07 $layer=LI1_cond $X=11.29 $Y=0.705
+ $X2=11.29 $Y2=0.58
r120 21 31 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.065 $Y=2.405
+ $X2=11.23 $Y2=2.405
r121 21 22 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=11.065 $Y=2.405
+ $X2=10.545 $Y2=2.405
r122 19 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=11.69 $Y=1.565
+ $X2=11.775 $Y2=1.48
r123 19 20 74.7005 $w=1.68e-07 $l=1.145e-06 $layer=LI1_cond $X=11.69 $Y=1.565
+ $X2=10.545 $Y2=1.565
r124 18 37 16.1564 $w=3.58e-07 $l=1.2e-07 $layer=POLY_cond $X=10.405 $Y=2.072
+ $X2=10.285 $Y2=2.072
r125 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.405
+ $Y=2.03 $X2=10.405 $Y2=2.03
r126 15 22 7.36005 $w=1.7e-07 $l=1.77482e-07 $layer=LI1_cond $X=10.405 $Y=2.32
+ $X2=10.545 $Y2=2.405
r127 15 17 11.936 $w=2.78e-07 $l=2.9e-07 $layer=LI1_cond $X=10.405 $Y=2.32
+ $X2=10.405 $Y2=2.03
r128 14 20 7.36005 $w=1.7e-07 $l=1.77482e-07 $layer=LI1_cond $X=10.405 $Y=1.65
+ $X2=10.545 $Y2=1.565
r129 14 17 15.6403 $w=2.78e-07 $l=3.8e-07 $layer=LI1_cond $X=10.405 $Y=1.65
+ $X2=10.405 $Y2=2.03
r130 10 37 23.1716 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=10.285 $Y=1.865
+ $X2=10.285 $Y2=2.072
r131 10 12 658.904 $w=1.5e-07 $l=1.285e-06 $layer=POLY_cond $X=10.285 $Y=1.865
+ $X2=10.285 $Y2=0.58
r132 7 36 23.1716 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=10.12 $Y=2.28
+ $X2=10.12 $Y2=2.072
r133 7 9 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=10.12 $Y=2.28
+ $X2=10.12 $Y2=2.565
r134 2 34 600 $w=1.7e-07 $l=2.74955e-07 $layer=licon1_PDIFF $count=1 $X=11.08
+ $Y=2.355 $X2=11.23 $Y2=2.565
r135 1 25 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=11.15
+ $Y=0.37 $X2=11.29 $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_HS__SDFRBP_2%A_1790_74# 1 2 9 11 12 13 15 16 18 20 23 25
+ 27 30 32 33 34 36 39 47 51 56 58 61 64
c151 58 0 1.03069e-19 $X=10.01 $Y=2.365
c152 56 0 1.57754e-19 $X=10.01 $Y=1.045
c153 13 0 3.10546e-20 $X=11.455 $Y=2.28
c154 12 0 7.64129e-20 $X=11.455 $Y=2.19
r155 61 62 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=11.355
+ $Y=1.175 $X2=11.355 $Y2=1.175
r156 59 64 0.195364 $w=2.65e-07 $l=8.5e-08 $layer=LI1_cond $X=10.095 $Y=1.177
+ $X2=10.01 $Y2=1.177
r157 59 61 54.7954 $w=2.63e-07 $l=1.26e-06 $layer=LI1_cond $X=10.095 $Y=1.177
+ $X2=11.355 $Y2=1.177
r158 57 64 7.34436 $w=1.7e-07 $l=1.33e-07 $layer=LI1_cond $X=10.01 $Y=1.31
+ $X2=10.01 $Y2=1.177
r159 57 58 68.8289 $w=1.68e-07 $l=1.055e-06 $layer=LI1_cond $X=10.01 $Y=1.31
+ $X2=10.01 $Y2=2.365
r160 56 64 7.34436 $w=1.7e-07 $l=1.32e-07 $layer=LI1_cond $X=10.01 $Y=1.045
+ $X2=10.01 $Y2=1.177
r161 55 56 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=10.01 $Y=0.735
+ $X2=10.01 $Y2=1.045
r162 51 55 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=9.925 $Y=0.57
+ $X2=10.01 $Y2=0.735
r163 51 53 9.42908 $w=3.28e-07 $l=2.7e-07 $layer=LI1_cond $X=9.925 $Y=0.57
+ $X2=9.655 $Y2=0.57
r164 47 58 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=9.925 $Y=2.53
+ $X2=10.01 $Y2=2.365
r165 47 49 19.382 $w=3.28e-07 $l=5.55e-07 $layer=LI1_cond $X=9.925 $Y=2.53
+ $X2=9.37 $Y2=2.53
r166 43 44 9.38961 $w=3.85e-07 $l=7.5e-08 $layer=POLY_cond $X=12.44 $Y=1.51
+ $X2=12.515 $Y2=1.51
r167 42 43 44.4442 $w=3.85e-07 $l=3.55e-07 $layer=POLY_cond $X=12.085 $Y=1.51
+ $X2=12.44 $Y2=1.51
r168 41 42 11.8935 $w=3.85e-07 $l=9.5e-08 $layer=POLY_cond $X=11.99 $Y=1.51
+ $X2=12.085 $Y2=1.51
r169 37 46 24.9301 $w=1.5e-07 $l=2.55e-07 $layer=POLY_cond $X=12.99 $Y=1.255
+ $X2=12.99 $Y2=1.51
r170 37 39 289.713 $w=1.5e-07 $l=5.65e-07 $layer=POLY_cond $X=12.99 $Y=1.255
+ $X2=12.99 $Y2=0.69
r171 34 36 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=12.945 $Y=1.885
+ $X2=12.945 $Y2=2.46
r172 33 34 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=12.945 $Y=1.795
+ $X2=12.945 $Y2=1.885
r173 32 46 5.63377 $w=3.85e-07 $l=4.5e-08 $layer=POLY_cond $X=12.945 $Y=1.51
+ $X2=12.99 $Y2=1.51
r174 32 44 53.8338 $w=3.85e-07 $l=4.3e-07 $layer=POLY_cond $X=12.945 $Y=1.51
+ $X2=12.515 $Y2=1.51
r175 32 33 81.629 $w=1.8e-07 $l=2.1e-07 $layer=POLY_cond $X=12.945 $Y=1.585
+ $X2=12.945 $Y2=1.795
r176 28 44 24.9301 $w=1.5e-07 $l=2.55e-07 $layer=POLY_cond $X=12.515 $Y=1.255
+ $X2=12.515 $Y2=1.51
r177 28 30 264.074 $w=1.5e-07 $l=5.15e-07 $layer=POLY_cond $X=12.515 $Y=1.255
+ $X2=12.515 $Y2=0.74
r178 25 43 24.9301 $w=1.5e-07 $l=2.55e-07 $layer=POLY_cond $X=12.44 $Y=1.765
+ $X2=12.44 $Y2=1.51
r179 25 27 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=12.44 $Y=1.765
+ $X2=12.44 $Y2=2.4
r180 21 42 24.9301 $w=1.5e-07 $l=2.55e-07 $layer=POLY_cond $X=12.085 $Y=1.255
+ $X2=12.085 $Y2=1.51
r181 21 23 264.074 $w=1.5e-07 $l=5.15e-07 $layer=POLY_cond $X=12.085 $Y=1.255
+ $X2=12.085 $Y2=0.74
r182 18 41 24.9301 $w=1.5e-07 $l=2.55e-07 $layer=POLY_cond $X=11.99 $Y=1.765
+ $X2=11.99 $Y2=1.51
r183 18 20 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=11.99 $Y=1.765
+ $X2=11.99 $Y2=2.4
r184 17 62 36.297 $w=3.28e-07 $l=3.76776e-07 $layer=POLY_cond $X=11.545 $Y=1.422
+ $X2=11.272 $Y2=1.175
r185 16 41 12.2091 $w=3.85e-07 $l=1.2657e-07 $layer=POLY_cond $X=11.9 $Y=1.422
+ $X2=11.99 $Y2=1.51
r186 16 17 61.1493 $w=3.35e-07 $l=3.55e-07 $layer=POLY_cond $X=11.9 $Y=1.422
+ $X2=11.545 $Y2=1.422
r187 13 15 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=11.455 $Y=2.28
+ $X2=11.455 $Y2=2.565
r188 12 13 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=11.455 $Y=2.19
+ $X2=11.455 $Y2=2.28
r189 11 17 34.4294 $w=3.28e-07 $l=2.08192e-07 $layer=POLY_cond $X=11.455 $Y=1.59
+ $X2=11.545 $Y2=1.422
r190 11 12 233.226 $w=1.8e-07 $l=6e-07 $layer=POLY_cond $X=11.455 $Y=1.59
+ $X2=11.455 $Y2=2.19
r191 7 62 38.5876 $w=3.28e-07 $l=2.67047e-07 $layer=POLY_cond $X=11.075 $Y=1.01
+ $X2=11.272 $Y2=1.175
r192 7 9 220.489 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=11.075 $Y=1.01
+ $X2=11.075 $Y2=0.58
r193 2 49 600 $w=1.7e-07 $l=9.51998e-07 $layer=licon1_PDIFF $count=1 $X=9.025
+ $Y=1.735 $X2=9.37 $Y2=2.53
r194 1 53 182 $w=1.7e-07 $l=7.98765e-07 $layer=licon1_NDIFF $count=1 $X=8.95
+ $Y=0.37 $X2=9.655 $Y2=0.57
.ends

.subckt PM_SKY130_FD_SC_HS__SDFRBP_2%A_2604_392# 1 2 7 9 12 14 16 19 21 24 28 32
+ 38 41
r51 38 39 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=13.8
+ $Y=1.465 $X2=13.8 $Y2=1.465
r52 36 41 0.499868 $w=3.3e-07 $l=1.3e-07 $layer=LI1_cond $X=13.325 $Y=1.465
+ $X2=13.195 $Y2=1.465
r53 36 38 16.5882 $w=3.28e-07 $l=4.75e-07 $layer=LI1_cond $X=13.325 $Y=1.465
+ $X2=13.8 $Y2=1.465
r54 32 34 31.4706 $w=2.58e-07 $l=7.1e-07 $layer=LI1_cond $X=13.195 $Y=2.105
+ $X2=13.195 $Y2=2.815
r55 30 41 6.26932 $w=2.6e-07 $l=1.65e-07 $layer=LI1_cond $X=13.195 $Y=1.63
+ $X2=13.195 $Y2=1.465
r56 30 32 21.0542 $w=2.58e-07 $l=4.75e-07 $layer=LI1_cond $X=13.195 $Y=1.63
+ $X2=13.195 $Y2=2.105
r57 26 41 6.26932 $w=2.6e-07 $l=1.65e-07 $layer=LI1_cond $X=13.195 $Y=1.3
+ $X2=13.195 $Y2=1.465
r58 26 28 34.7949 $w=2.58e-07 $l=7.85e-07 $layer=LI1_cond $X=13.195 $Y=1.3
+ $X2=13.195 $Y2=0.515
r59 24 25 1.77641 $w=4.07e-07 $l=1.5e-08 $layer=POLY_cond $X=14.385 $Y=1.532
+ $X2=14.4 $Y2=1.532
r60 23 24 49.1474 $w=4.07e-07 $l=4.15e-07 $layer=POLY_cond $X=13.97 $Y=1.532
+ $X2=14.385 $Y2=1.532
r61 22 23 4.14496 $w=4.07e-07 $l=3.5e-08 $layer=POLY_cond $X=13.935 $Y=1.532
+ $X2=13.97 $Y2=1.532
r62 21 39 7.86876 $w=3.3e-07 $l=4.5e-08 $layer=POLY_cond $X=13.845 $Y=1.465
+ $X2=13.8 $Y2=1.465
r63 21 22 12.5251 $w=4.07e-07 $l=1.1887e-07 $layer=POLY_cond $X=13.845 $Y=1.465
+ $X2=13.935 $Y2=1.532
r64 17 25 26.2866 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=14.4 $Y=1.3
+ $X2=14.4 $Y2=1.532
r65 17 19 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=14.4 $Y=1.3 $X2=14.4
+ $Y2=0.74
r66 14 24 26.2866 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=14.385 $Y=1.765
+ $X2=14.385 $Y2=1.532
r67 14 16 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=14.385 $Y=1.765
+ $X2=14.385 $Y2=2.4
r68 10 23 26.2866 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=13.97 $Y=1.3
+ $X2=13.97 $Y2=1.532
r69 10 12 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=13.97 $Y=1.3
+ $X2=13.97 $Y2=0.74
r70 7 22 26.2866 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=13.935 $Y=1.765
+ $X2=13.935 $Y2=1.532
r71 7 9 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=13.935 $Y=1.765
+ $X2=13.935 $Y2=2.4
r72 2 34 400 $w=1.7e-07 $l=9.26971e-07 $layer=licon1_PDIFF $count=1 $X=13.02
+ $Y=1.96 $X2=13.17 $Y2=2.815
r73 2 32 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=13.02
+ $Y=1.96 $X2=13.17 $Y2=2.105
r74 1 28 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=13.065
+ $Y=0.37 $X2=13.205 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__SDFRBP_2%VPWR 1 2 3 4 5 6 7 8 9 10 33 37 41 45 49 53
+ 59 65 69 71 76 77 79 80 81 88 106 110 115 120 125 133 136 138 141 144 151 154
+ 157 161
r182 160 161 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=14.64 $Y=3.33
+ $X2=14.64 $Y2=3.33
r183 157 158 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.68 $Y=3.33
+ $X2=13.68 $Y2=3.33
r184 154 155 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.72 $Y=3.33
+ $X2=12.72 $Y2=3.33
r185 151 152 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.76 $Y=3.33
+ $X2=11.76 $Y2=3.33
r186 142 148 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=8.4 $Y=3.33
+ $X2=10.32 $Y2=3.33
r187 141 142 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=8.4 $Y=3.33
+ $X2=8.4 $Y2=3.33
r188 138 139 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r189 135 136 10.7086 $w=6.83e-07 $l=1.65e-07 $layer=LI1_cond $X=1.235 $Y=3.072
+ $X2=1.4 $Y2=3.072
r190 131 135 0.611135 $w=6.83e-07 $l=3.5e-08 $layer=LI1_cond $X=1.2 $Y=3.072
+ $X2=1.235 $Y2=3.072
r191 131 133 18.0422 $w=6.83e-07 $l=5.85e-07 $layer=LI1_cond $X=1.2 $Y=3.072
+ $X2=0.615 $Y2=3.072
r192 131 132 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r193 129 161 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=14.16 $Y=3.33
+ $X2=14.64 $Y2=3.33
r194 129 158 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=14.16 $Y=3.33
+ $X2=13.68 $Y2=3.33
r195 128 129 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=14.16 $Y=3.33
+ $X2=14.16 $Y2=3.33
r196 126 157 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=13.875 $Y=3.33
+ $X2=13.71 $Y2=3.33
r197 126 128 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=13.875 $Y=3.33
+ $X2=14.16 $Y2=3.33
r198 125 160 4.29523 $w=1.7e-07 $l=1.92e-07 $layer=LI1_cond $X=14.495 $Y=3.33
+ $X2=14.687 $Y2=3.33
r199 125 128 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=14.495 $Y=3.33
+ $X2=14.16 $Y2=3.33
r200 124 158 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=13.2 $Y=3.33
+ $X2=13.68 $Y2=3.33
r201 124 155 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=13.2 $Y=3.33
+ $X2=12.72 $Y2=3.33
r202 123 124 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.2 $Y=3.33
+ $X2=13.2 $Y2=3.33
r203 121 154 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=12.83 $Y=3.33
+ $X2=12.685 $Y2=3.33
r204 121 123 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=12.83 $Y=3.33
+ $X2=13.2 $Y2=3.33
r205 120 157 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=13.545 $Y=3.33
+ $X2=13.71 $Y2=3.33
r206 120 123 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=13.545 $Y=3.33
+ $X2=13.2 $Y2=3.33
r207 119 155 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.24 $Y=3.33
+ $X2=12.72 $Y2=3.33
r208 119 152 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.24 $Y=3.33
+ $X2=11.76 $Y2=3.33
r209 118 119 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.24 $Y=3.33
+ $X2=12.24 $Y2=3.33
r210 116 151 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=11.85 $Y=3.33
+ $X2=11.725 $Y2=3.33
r211 116 118 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=11.85 $Y=3.33
+ $X2=12.24 $Y2=3.33
r212 115 154 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=12.54 $Y=3.33
+ $X2=12.685 $Y2=3.33
r213 115 118 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=12.54 $Y=3.33
+ $X2=12.24 $Y2=3.33
r214 114 152 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.28 $Y=3.33
+ $X2=11.76 $Y2=3.33
r215 114 148 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=11.28 $Y=3.33
+ $X2=10.32 $Y2=3.33
r216 113 114 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=11.28 $Y=3.33
+ $X2=11.28 $Y2=3.33
r217 111 113 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=10.86 $Y=3.33
+ $X2=11.28 $Y2=3.33
r218 110 151 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=11.6 $Y=3.33
+ $X2=11.725 $Y2=3.33
r219 110 113 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=11.6 $Y=3.33
+ $X2=11.28 $Y2=3.33
r220 109 142 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=3.33
+ $X2=8.4 $Y2=3.33
r221 108 109 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r222 106 141 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.19 $Y=3.33
+ $X2=8.315 $Y2=3.33
r223 106 108 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=8.19 $Y=3.33
+ $X2=7.92 $Y2=3.33
r224 104 105 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r225 102 105 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=6.96 $Y2=3.33
r226 101 104 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=5.04 $Y=3.33
+ $X2=6.96 $Y2=3.33
r227 101 102 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r228 99 102 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=5.04 $Y2=3.33
r229 98 99 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r230 96 99 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.56 $Y2=3.33
r231 96 139 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=3.12 $Y2=3.33
r232 95 98 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=3.6 $Y=3.33 $X2=4.56
+ $Y2=3.33
r233 95 96 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r234 93 138 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.445 $Y=3.33
+ $X2=3.28 $Y2=3.33
r235 93 95 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=3.445 $Y=3.33
+ $X2=3.6 $Y2=3.33
r236 92 139 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=3.12 $Y2=3.33
r237 92 132 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r238 91 136 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=1.68 $Y=3.33
+ $X2=1.4 $Y2=3.33
r239 91 92 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r240 88 138 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.115 $Y=3.33
+ $X2=3.28 $Y2=3.33
r241 88 91 93.6203 $w=1.68e-07 $l=1.435e-06 $layer=LI1_cond $X=3.115 $Y=3.33
+ $X2=1.68 $Y2=3.33
r242 86 132 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=1.2 $Y2=3.33
r243 85 133 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=0.24 $Y=3.33
+ $X2=0.615 $Y2=3.33
r244 85 86 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r245 81 109 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=7.92 $Y2=3.33
r246 81 105 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=6.96 $Y2=3.33
r247 79 104 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=7.07 $Y=3.33
+ $X2=6.96 $Y2=3.33
r248 79 80 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.07 $Y=3.33
+ $X2=7.195 $Y2=3.33
r249 78 108 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=7.32 $Y=3.33
+ $X2=7.92 $Y2=3.33
r250 78 80 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.32 $Y=3.33
+ $X2=7.195 $Y2=3.33
r251 76 98 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=4.705 $Y=3.33
+ $X2=4.56 $Y2=3.33
r252 76 77 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.705 $Y=3.33
+ $X2=4.87 $Y2=3.33
r253 75 101 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=5.035 $Y=3.33
+ $X2=5.04 $Y2=3.33
r254 75 77 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.035 $Y=3.33
+ $X2=4.87 $Y2=3.33
r255 71 74 34.1617 $w=2.78e-07 $l=8.3e-07 $layer=LI1_cond $X=14.635 $Y=1.985
+ $X2=14.635 $Y2=2.815
r256 69 160 3.06482 $w=2.8e-07 $l=1.07912e-07 $layer=LI1_cond $X=14.635 $Y=3.245
+ $X2=14.687 $Y2=3.33
r257 69 74 17.6982 $w=2.78e-07 $l=4.3e-07 $layer=LI1_cond $X=14.635 $Y=3.245
+ $X2=14.635 $Y2=2.815
r258 65 68 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=13.71 $Y=1.985
+ $X2=13.71 $Y2=2.815
r259 63 157 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=13.71 $Y=3.245
+ $X2=13.71 $Y2=3.33
r260 63 68 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=13.71 $Y=3.245
+ $X2=13.71 $Y2=2.815
r261 59 62 29.0098 $w=2.88e-07 $l=7.3e-07 $layer=LI1_cond $X=12.685 $Y=2.085
+ $X2=12.685 $Y2=2.815
r262 57 154 0.489042 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=12.685 $Y=3.245
+ $X2=12.685 $Y2=3.33
r263 57 62 17.0879 $w=2.88e-07 $l=4.3e-07 $layer=LI1_cond $X=12.685 $Y=3.245
+ $X2=12.685 $Y2=2.815
r264 53 56 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=11.725 $Y=1.985
+ $X2=11.725 $Y2=2.815
r265 51 151 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=11.725 $Y=3.245
+ $X2=11.725 $Y2=3.33
r266 51 56 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=11.725 $Y=3.245
+ $X2=11.725 $Y2=2.815
r267 50 141 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.44 $Y=3.33
+ $X2=8.315 $Y2=3.33
r268 49 111 8.26286 $w=1.7e-07 $l=2.98e-07 $layer=LI1_cond $X=10.562 $Y=3.33
+ $X2=10.86 $Y2=3.33
r269 49 148 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=10.32 $Y=3.33
+ $X2=10.32 $Y2=3.33
r270 49 144 10.1516 $w=5.93e-07 $l=5.05e-07 $layer=LI1_cond $X=10.562 $Y=3.33
+ $X2=10.562 $Y2=2.825
r271 49 50 119.064 $w=1.68e-07 $l=1.825e-06 $layer=LI1_cond $X=10.265 $Y=3.33
+ $X2=8.44 $Y2=3.33
r272 45 48 31.3464 $w=2.48e-07 $l=6.8e-07 $layer=LI1_cond $X=8.315 $Y=1.91
+ $X2=8.315 $Y2=2.59
r273 43 141 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=8.315 $Y=3.245
+ $X2=8.315 $Y2=3.33
r274 43 48 30.194 $w=2.48e-07 $l=6.55e-07 $layer=LI1_cond $X=8.315 $Y=3.245
+ $X2=8.315 $Y2=2.59
r275 39 80 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=7.195 $Y=3.245
+ $X2=7.195 $Y2=3.33
r276 39 41 18.4391 $w=2.48e-07 $l=4e-07 $layer=LI1_cond $X=7.195 $Y=3.245
+ $X2=7.195 $Y2=2.845
r277 35 77 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.87 $Y=3.245
+ $X2=4.87 $Y2=3.33
r278 35 37 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=4.87 $Y=3.245
+ $X2=4.87 $Y2=2.795
r279 31 138 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.28 $Y=3.245
+ $X2=3.28 $Y2=3.33
r280 31 33 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=3.28 $Y=3.245
+ $X2=3.28 $Y2=2.78
r281 10 74 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=14.46
+ $Y=1.84 $X2=14.61 $Y2=2.815
r282 10 71 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=14.46
+ $Y=1.84 $X2=14.61 $Y2=1.985
r283 9 68 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=13.565
+ $Y=1.84 $X2=13.71 $Y2=2.815
r284 9 65 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=13.565
+ $Y=1.84 $X2=13.71 $Y2=1.985
r285 8 62 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=12.515
+ $Y=1.84 $X2=12.665 $Y2=2.815
r286 8 59 400 $w=1.7e-07 $l=3.11087e-07 $layer=licon1_PDIFF $count=1 $X=12.515
+ $Y=1.84 $X2=12.665 $Y2=2.085
r287 7 56 600 $w=1.7e-07 $l=5.6542e-07 $layer=licon1_PDIFF $count=1 $X=11.53
+ $Y=2.355 $X2=11.765 $Y2=2.815
r288 7 53 300 $w=1.7e-07 $l=4.73128e-07 $layer=licon1_PDIFF $count=2 $X=11.53
+ $Y=2.355 $X2=11.765 $Y2=1.985
r289 6 144 600 $w=1.7e-07 $l=6.26458e-07 $layer=licon1_PDIFF $count=1 $X=10.195
+ $Y=2.355 $X2=10.56 $Y2=2.825
r290 5 48 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=8.15
+ $Y=1.735 $X2=8.275 $Y2=2.59
r291 5 45 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=8.15
+ $Y=1.735 $X2=8.275 $Y2=1.91
r292 4 41 600 $w=1.7e-07 $l=6.60908e-07 $layer=licon1_PDIFF $count=1 $X=7.015
+ $Y=2.285 $X2=7.235 $Y2=2.845
r293 3 37 600 $w=1.7e-07 $l=1.02727e-06 $layer=licon1_PDIFF $count=1 $X=4.72
+ $Y=1.84 $X2=4.87 $Y2=2.795
r294 2 33 600 $w=1.7e-07 $l=5.38331e-07 $layer=licon1_PDIFF $count=1 $X=3.11
+ $Y=2.32 $X2=3.28 $Y2=2.78
r295 1 135 300 $w=1.7e-07 $l=8.679e-07 $layer=licon1_PDIFF $count=2 $X=0.58
+ $Y=2.32 $X2=1.235 $Y2=2.815
.ends

.subckt PM_SKY130_FD_SC_HS__SDFRBP_2%A_388_79# 1 2 3 4 5 16 22 24 25 27 28 29 31
+ 32 35 36 40 41 42 43 44 46 50 54
c155 46 0 5.24149e-20 $X=6.405 $Y=2
c156 44 0 3.46724e-20 $X=5.99 $Y=1.205
c157 40 0 4.26327e-21 $X=5.905 $Y=1.12
c158 36 0 1.00595e-19 $X=3.995 $Y=2.435
c159 24 0 1.55498e-19 $X=3.445 $Y=1.09
r160 45 46 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=6.405 $Y=1.29
+ $X2=6.405 $Y2=2
r161 43 45 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.32 $Y=1.205
+ $X2=6.405 $Y2=1.29
r162 43 44 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=6.32 $Y=1.205
+ $X2=5.99 $Y2=1.205
r163 41 46 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.32 $Y=2.085
+ $X2=6.405 $Y2=2
r164 41 42 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=6.32 $Y=2.085
+ $X2=5.985 $Y2=2.085
r165 40 44 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.905 $Y=1.12
+ $X2=5.99 $Y2=1.205
r166 39 50 0.716491 $w=1.7e-07 $l=1.18427e-07 $layer=LI1_cond $X=5.905 $Y=0.82
+ $X2=5.825 $Y2=0.735
r167 39 40 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=5.905 $Y=0.82
+ $X2=5.905 $Y2=1.12
r168 37 42 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.9 $Y=2.17
+ $X2=5.985 $Y2=2.085
r169 37 54 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=5.9 $Y=2.17 $X2=5.9
+ $Y2=2.33
r170 35 56 3.77163 $w=2.73e-07 $l=9e-08 $layer=LI1_cond $X=5.847 $Y=2.435
+ $X2=5.847 $Y2=2.525
r171 35 54 6.06982 $w=2.73e-07 $l=1.05e-07 $layer=LI1_cond $X=5.847 $Y=2.435
+ $X2=5.847 $Y2=2.33
r172 35 36 111.888 $w=1.68e-07 $l=1.715e-06 $layer=LI1_cond $X=5.71 $Y=2.435
+ $X2=3.995 $Y2=2.435
r173 32 36 12.363 $w=1.9e-07 $l=1.97358e-07 $layer=LI1_cond $X=3.805 $Y=2.42
+ $X2=3.995 $Y2=2.435
r174 32 47 17.6579 $w=1.9e-07 $l=2.75e-07 $layer=LI1_cond $X=3.805 $Y=2.42
+ $X2=3.53 $Y2=2.42
r175 32 34 4.17368 $w=3.8e-07 $l=1.3e-07 $layer=LI1_cond $X=3.805 $Y=2.52
+ $X2=3.805 $Y2=2.65
r176 31 47 1.386 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=3.53 $Y=2.32 $X2=3.53
+ $Y2=2.42
r177 30 31 74.7005 $w=1.68e-07 $l=1.145e-06 $layer=LI1_cond $X=3.53 $Y=1.175
+ $X2=3.53 $Y2=2.32
r178 28 47 5.62091 $w=1.9e-07 $l=9.21954e-08 $layer=LI1_cond $X=3.445 $Y=2.405
+ $X2=3.53 $Y2=2.42
r179 28 29 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=3.445 $Y=2.405
+ $X2=2.945 $Y2=2.405
r180 26 29 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.86 $Y=2.49
+ $X2=2.945 $Y2=2.405
r181 26 27 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=2.86 $Y=2.49
+ $X2=2.86 $Y2=2.66
r182 24 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.445 $Y=1.09
+ $X2=3.53 $Y2=1.175
r183 24 25 54.4759 $w=1.68e-07 $l=8.35e-07 $layer=LI1_cond $X=3.445 $Y=1.09
+ $X2=2.61 $Y2=1.09
r184 20 25 7.93686 $w=1.7e-07 $l=2.13307e-07 $layer=LI1_cond $X=2.435 $Y=1.005
+ $X2=2.61 $Y2=1.09
r185 20 22 10.7013 $w=3.48e-07 $l=3.25e-07 $layer=LI1_cond $X=2.435 $Y=1.005
+ $X2=2.435 $Y2=0.68
r186 16 27 7.14316 $w=2.5e-07 $l=1.62019e-07 $layer=LI1_cond $X=2.775 $Y=2.785
+ $X2=2.86 $Y2=2.66
r187 16 18 24.4318 $w=2.48e-07 $l=5.3e-07 $layer=LI1_cond $X=2.775 $Y=2.785
+ $X2=2.245 $Y2=2.785
r188 5 56 600 $w=1.7e-07 $l=2.97993e-07 $layer=licon1_PDIFF $count=1 $X=5.745
+ $Y=2.285 $X2=5.875 $Y2=2.525
r189 4 34 600 $w=1.7e-07 $l=3.97995e-07 $layer=licon1_PDIFF $count=1 $X=3.68
+ $Y=2.32 $X2=3.83 $Y2=2.65
r190 3 18 600 $w=1.7e-07 $l=5.51249e-07 $layer=licon1_PDIFF $count=1 $X=1.955
+ $Y=2.32 $X2=2.245 $Y2=2.745
r191 2 50 182 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=1 $X=5.68
+ $Y=0.59 $X2=5.825 $Y2=0.735
r192 1 22 182 $w=1.7e-07 $l=6.21369e-07 $layer=licon1_NDIFF $count=1 $X=1.94
+ $Y=0.395 $X2=2.435 $Y2=0.68
.ends

.subckt PM_SKY130_FD_SC_HS__SDFRBP_2%Q_N 1 2 7 8 9 16 30
r28 30 31 0.96397 $w=4.33e-07 $l=1e-08 $layer=LI1_cond $X=12.247 $Y=0.925
+ $X2=12.247 $Y2=0.915
r29 25 27 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=12.195 $Y=1.985
+ $X2=12.195 $Y2=2.815
r30 9 25 11.1752 $w=3.28e-07 $l=3.2e-07 $layer=LI1_cond $X=12.195 $Y=1.665
+ $X2=12.195 $Y2=1.985
r31 8 9 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=12.195 $Y=1.295
+ $X2=12.195 $Y2=1.665
r32 8 33 7.33373 $w=3.28e-07 $l=2.1e-07 $layer=LI1_cond $X=12.195 $Y=1.295
+ $X2=12.195 $Y2=1.085
r33 7 33 3.95767 $w=4.33e-07 $l=1.23e-07 $layer=LI1_cond $X=12.247 $Y=0.962
+ $X2=12.247 $Y2=1.085
r34 7 30 0.980239 $w=4.33e-07 $l=3.7e-08 $layer=LI1_cond $X=12.247 $Y=0.962
+ $X2=12.247 $Y2=0.925
r35 7 31 1.32706 $w=3.28e-07 $l=3.8e-08 $layer=LI1_cond $X=12.3 $Y=0.877
+ $X2=12.3 $Y2=0.915
r36 7 16 12.642 $w=3.28e-07 $l=3.62e-07 $layer=LI1_cond $X=12.3 $Y=0.877
+ $X2=12.3 $Y2=0.515
r37 2 27 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=12.065
+ $Y=1.84 $X2=12.215 $Y2=2.815
r38 2 25 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=12.065
+ $Y=1.84 $X2=12.215 $Y2=1.985
r39 1 16 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=12.16
+ $Y=0.37 $X2=12.3 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__SDFRBP_2%Q 1 2 7 10
r16 7 16 35.427 $w=2.68e-07 $l=8.3e-07 $layer=LI1_cond $X=14.19 $Y=1.985
+ $X2=14.19 $Y2=2.815
r17 7 10 62.7441 $w=2.68e-07 $l=1.47e-06 $layer=LI1_cond $X=14.19 $Y=1.985
+ $X2=14.19 $Y2=0.515
r18 2 16 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=14.01
+ $Y=1.84 $X2=14.16 $Y2=2.815
r19 2 7 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=14.01
+ $Y=1.84 $X2=14.16 $Y2=1.985
r20 1 10 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=14.045
+ $Y=0.37 $X2=14.185 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__SDFRBP_2%VGND 1 2 3 4 5 6 7 8 9 30 34 38 42 46 50 52
+ 56 58 60 63 64 66 67 69 70 71 73 99 103 108 114 118 122 124 127 130 134
c157 134 0 3.19474e-20 $X=14.64 $Y=0
r158 133 134 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=14.64 $Y=0
+ $X2=14.64 $Y2=0
r159 130 131 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=13.68 $Y=0
+ $X2=13.68 $Y2=0
r160 128 131 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=12.72 $Y=0
+ $X2=13.68 $Y2=0
r161 127 128 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.72 $Y=0
+ $X2=12.72 $Y2=0
r162 124 125 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.76 $Y=0
+ $X2=11.76 $Y2=0
r163 120 122 7.07024 $w=4.93e-07 $l=6.5e-08 $layer=LI1_cond $X=7.92 $Y=0.162
+ $X2=7.985 $Y2=0.162
r164 120 121 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=7.92 $Y=0
+ $X2=7.92 $Y2=0
r165 117 120 4.95346 $w=4.93e-07 $l=2.05e-07 $layer=LI1_cond $X=7.715 $Y=0.162
+ $X2=7.92 $Y2=0.162
r166 117 118 11.9029 $w=4.93e-07 $l=2.65e-07 $layer=LI1_cond $X=7.715 $Y=0.162
+ $X2=7.45 $Y2=0.162
r167 114 115 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0
+ $X2=0.72 $Y2=0
r168 112 134 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=14.16 $Y=0
+ $X2=14.64 $Y2=0
r169 112 131 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=14.16 $Y=0
+ $X2=13.68 $Y2=0
r170 111 112 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=14.16 $Y=0
+ $X2=14.16 $Y2=0
r171 109 130 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=13.84 $Y=0
+ $X2=13.755 $Y2=0
r172 109 111 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=13.84 $Y=0
+ $X2=14.16 $Y2=0
r173 108 133 4.34417 $w=1.7e-07 $l=1.92e-07 $layer=LI1_cond $X=14.495 $Y=0
+ $X2=14.687 $Y2=0
r174 108 111 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=14.495 $Y=0
+ $X2=14.16 $Y2=0
r175 107 128 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.24 $Y=0
+ $X2=12.72 $Y2=0
r176 107 125 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.24 $Y=0
+ $X2=11.76 $Y2=0
r177 106 107 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.24 $Y=0
+ $X2=12.24 $Y2=0
r178 104 124 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=11.895 $Y=0
+ $X2=11.77 $Y2=0
r179 104 106 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=11.895 $Y=0
+ $X2=12.24 $Y2=0
r180 103 127 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=12.635 $Y=0
+ $X2=12.765 $Y2=0
r181 103 106 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=12.635 $Y=0
+ $X2=12.24 $Y2=0
r182 102 125 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.28 $Y=0
+ $X2=11.76 $Y2=0
r183 101 102 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=11.28 $Y=0
+ $X2=11.28 $Y2=0
r184 99 124 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=11.645 $Y=0
+ $X2=11.77 $Y2=0
r185 99 101 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=11.645 $Y=0
+ $X2=11.28 $Y2=0
r186 98 102 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=10.32 $Y=0
+ $X2=11.28 $Y2=0
r187 98 121 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=10.32 $Y=0
+ $X2=7.92 $Y2=0
r188 97 122 152.337 $w=1.68e-07 $l=2.335e-06 $layer=LI1_cond $X=10.32 $Y=0
+ $X2=7.985 $Y2=0
r189 97 98 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=10.32 $Y=0
+ $X2=10.32 $Y2=0
r190 93 118 0.652406 $w=1.68e-07 $l=1e-08 $layer=LI1_cond $X=7.44 $Y=0 $X2=7.45
+ $Y2=0
r191 90 93 156.578 $w=1.68e-07 $l=2.4e-06 $layer=LI1_cond $X=5.04 $Y=0 $X2=7.44
+ $Y2=0
r192 90 91 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r193 87 91 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=5.04
+ $Y2=0
r194 86 87 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r195 84 87 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.56
+ $Y2=0
r196 83 84 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r197 81 84 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=1.2 $Y=0 $X2=3.6
+ $Y2=0
r198 81 115 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r199 80 83 156.578 $w=1.68e-07 $l=2.4e-06 $layer=LI1_cond $X=1.2 $Y=0 $X2=3.6
+ $Y2=0
r200 80 81 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r201 78 114 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.875 $Y=0
+ $X2=0.71 $Y2=0
r202 78 80 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.875 $Y=0 $X2=1.2
+ $Y2=0
r203 76 115 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0
+ $X2=0.72 $Y2=0
r204 75 76 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r205 73 114 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.545 $Y=0
+ $X2=0.71 $Y2=0
r206 73 75 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.545 $Y=0
+ $X2=0.24 $Y2=0
r207 71 121 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=0
+ $X2=7.92 $Y2=0
r208 71 91 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=7.44 $Y=0 $X2=5.04
+ $Y2=0
r209 71 93 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=7.44 $Y=0 $X2=7.44
+ $Y2=0
r210 69 97 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=10.335 $Y=0
+ $X2=10.32 $Y2=0
r211 69 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.335 $Y=0
+ $X2=10.5 $Y2=0
r212 68 101 40.123 $w=1.68e-07 $l=6.15e-07 $layer=LI1_cond $X=10.665 $Y=0
+ $X2=11.28 $Y2=0
r213 68 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.665 $Y=0
+ $X2=10.5 $Y2=0
r214 66 86 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=4.75 $Y=0 $X2=4.56
+ $Y2=0
r215 66 67 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.75 $Y=0 $X2=4.835
+ $Y2=0
r216 65 90 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=4.92 $Y=0 $X2=5.04
+ $Y2=0
r217 65 67 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.92 $Y=0 $X2=4.835
+ $Y2=0
r218 63 83 2.60963 $w=1.68e-07 $l=4e-08 $layer=LI1_cond $X=3.64 $Y=0 $X2=3.6
+ $Y2=0
r219 63 64 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.64 $Y=0 $X2=3.805
+ $Y2=0
r220 62 86 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=3.97 $Y=0 $X2=4.56
+ $Y2=0
r221 62 64 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.97 $Y=0 $X2=3.805
+ $Y2=0
r222 58 133 3.0545 $w=2.85e-07 $l=1.07121e-07 $layer=LI1_cond $X=14.637 $Y=0.085
+ $X2=14.687 $Y2=0
r223 58 60 17.3877 $w=2.83e-07 $l=4.3e-07 $layer=LI1_cond $X=14.637 $Y=0.085
+ $X2=14.637 $Y2=0.515
r224 54 130 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=13.755 $Y=0.085
+ $X2=13.755 $Y2=0
r225 54 56 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=13.755 $Y=0.085
+ $X2=13.755 $Y2=0.515
r226 53 127 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=12.895 $Y=0
+ $X2=12.765 $Y2=0
r227 52 130 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=13.67 $Y=0
+ $X2=13.755 $Y2=0
r228 52 53 50.5615 $w=1.68e-07 $l=7.75e-07 $layer=LI1_cond $X=13.67 $Y=0
+ $X2=12.895 $Y2=0
r229 48 127 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=12.765 $Y=0.085
+ $X2=12.765 $Y2=0
r230 48 50 20.3894 $w=2.58e-07 $l=4.6e-07 $layer=LI1_cond $X=12.765 $Y=0.085
+ $X2=12.765 $Y2=0.545
r231 44 124 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=11.77 $Y=0.085
+ $X2=11.77 $Y2=0
r232 44 46 13.1378 $w=2.48e-07 $l=2.85e-07 $layer=LI1_cond $X=11.77 $Y=0.085
+ $X2=11.77 $Y2=0.37
r233 40 70 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=10.5 $Y=0.085
+ $X2=10.5 $Y2=0
r234 40 42 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=10.5 $Y=0.085
+ $X2=10.5 $Y2=0.58
r235 36 67 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.835 $Y=0.085
+ $X2=4.835 $Y2=0
r236 36 38 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=4.835 $Y=0.085
+ $X2=4.835 $Y2=0.515
r237 32 64 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.805 $Y=0.085
+ $X2=3.805 $Y2=0
r238 32 34 18.1597 $w=3.28e-07 $l=5.2e-07 $layer=LI1_cond $X=3.805 $Y=0.085
+ $X2=3.805 $Y2=0.605
r239 28 114 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.71 $Y=0.085
+ $X2=0.71 $Y2=0
r240 28 30 18.1597 $w=3.28e-07 $l=5.2e-07 $layer=LI1_cond $X=0.71 $Y=0.085
+ $X2=0.71 $Y2=0.605
r241 9 60 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=14.475
+ $Y=0.37 $X2=14.615 $Y2=0.515
r242 8 56 91 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_NDIFF $count=2 $X=13.6
+ $Y=0.37 $X2=13.755 $Y2=0.515
r243 7 50 91 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_NDIFF $count=2 $X=12.59
+ $Y=0.37 $X2=12.73 $Y2=0.545
r244 6 46 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=11.685
+ $Y=0.225 $X2=11.81 $Y2=0.37
r245 5 42 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=10.36
+ $Y=0.37 $X2=10.5 $Y2=0.58
r246 4 117 182 $w=1.7e-07 $l=4.32666e-07 $layer=licon1_NDIFF $count=1 $X=7.395
+ $Y=0.59 $X2=7.715 $Y2=0.325
r247 3 38 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=4.695
+ $Y=0.37 $X2=4.835 $Y2=0.515
r248 2 34 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=3.665
+ $Y=0.395 $X2=3.805 $Y2=0.605
r249 1 30 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.395 $X2=0.71 $Y2=0.605
.ends

.subckt PM_SKY130_FD_SC_HS__SDFRBP_2%noxref_25 1 2 9 11 12 15
r35 13 15 6.28605 $w=3.28e-07 $l=1.8e-07 $layer=LI1_cond $X=3.265 $Y=0.425
+ $X2=3.265 $Y2=0.605
r36 11 13 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.1 $Y=0.34
+ $X2=3.265 $Y2=0.425
r37 11 12 114.497 $w=1.68e-07 $l=1.755e-06 $layer=LI1_cond $X=3.1 $Y=0.34
+ $X2=1.345 $Y2=0.34
r38 7 12 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.22 $Y=0.425
+ $X2=1.345 $Y2=0.34
r39 7 9 8.29759 $w=2.48e-07 $l=1.8e-07 $layer=LI1_cond $X=1.22 $Y=0.425 $X2=1.22
+ $Y2=0.605
r40 2 15 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=3.125
+ $Y=0.395 $X2=3.265 $Y2=0.605
r41 1 9 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=1.115
+ $Y=0.395 $X2=1.26 $Y2=0.605
.ends

