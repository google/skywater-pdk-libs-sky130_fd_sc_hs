* File: sky130_fd_sc_hs__sdfstp_1.pxi.spice
* Created: Thu Aug 27 21:09:27 2020
* 
x_PM_SKY130_FD_SC_HS__SDFSTP_1%SCE N_SCE_c_302_n N_SCE_c_303_n N_SCE_M1025_g
+ N_SCE_M1021_g N_SCE_c_304_n N_SCE_c_305_n N_SCE_c_306_n N_SCE_M1024_g
+ N_SCE_M1004_g N_SCE_c_296_n N_SCE_c_308_n N_SCE_c_297_n N_SCE_c_298_n
+ N_SCE_c_299_n SCE N_SCE_c_301_n PM_SKY130_FD_SC_HS__SDFSTP_1%SCE
x_PM_SKY130_FD_SC_HS__SDFSTP_1%A_27_464# N_A_27_464#_M1021_s N_A_27_464#_M1025_s
+ N_A_27_464#_M1002_g N_A_27_464#_c_389_n N_A_27_464#_M1020_g
+ N_A_27_464#_c_383_n N_A_27_464#_c_384_n N_A_27_464#_c_401_n
+ N_A_27_464#_c_385_n N_A_27_464#_c_391_n N_A_27_464#_c_386_n
+ N_A_27_464#_c_392_n N_A_27_464#_c_387_n N_A_27_464#_c_388_n
+ PM_SKY130_FD_SC_HS__SDFSTP_1%A_27_464#
x_PM_SKY130_FD_SC_HS__SDFSTP_1%D N_D_c_466_n N_D_M1031_g N_D_M1026_g D
+ N_D_c_468_n PM_SKY130_FD_SC_HS__SDFSTP_1%D
x_PM_SKY130_FD_SC_HS__SDFSTP_1%SCD N_SCD_c_501_n N_SCD_M1003_g N_SCD_c_505_n
+ N_SCD_M1028_g N_SCD_c_506_n SCD SCD SCD N_SCD_c_503_n N_SCD_c_504_n
+ PM_SKY130_FD_SC_HS__SDFSTP_1%SCD
x_PM_SKY130_FD_SC_HS__SDFSTP_1%CLK N_CLK_c_546_n N_CLK_M1005_g N_CLK_c_547_n
+ N_CLK_M1032_g CLK PM_SKY130_FD_SC_HS__SDFSTP_1%CLK
x_PM_SKY130_FD_SC_HS__SDFSTP_1%A_800_74# N_A_800_74#_M1015_d N_A_800_74#_M1037_d
+ N_A_800_74#_c_580_n N_A_800_74#_M1014_g N_A_800_74#_M1011_g
+ N_A_800_74#_c_582_n N_A_800_74#_M1001_g N_A_800_74#_c_583_n
+ N_A_800_74#_c_597_n N_A_800_74#_M1009_g N_A_800_74#_c_584_n
+ N_A_800_74#_c_713_p N_A_800_74#_c_585_n N_A_800_74#_c_586_n
+ N_A_800_74#_c_598_n N_A_800_74#_c_599_n N_A_800_74#_c_587_n
+ N_A_800_74#_c_588_n N_A_800_74#_c_601_n N_A_800_74#_c_602_n
+ N_A_800_74#_c_619_p N_A_800_74#_c_603_n N_A_800_74#_c_604_n
+ N_A_800_74#_c_605_n N_A_800_74#_c_606_n N_A_800_74#_c_607_n
+ N_A_800_74#_c_608_n N_A_800_74#_c_646_p N_A_800_74#_c_589_n
+ N_A_800_74#_c_610_n N_A_800_74#_c_590_n N_A_800_74#_c_611_n
+ N_A_800_74#_c_809_p N_A_800_74#_c_591_n N_A_800_74#_c_592_n
+ N_A_800_74#_c_593_n N_A_800_74#_c_594_n PM_SKY130_FD_SC_HS__SDFSTP_1%A_800_74#
x_PM_SKY130_FD_SC_HS__SDFSTP_1%A_1198_55# N_A_1198_55#_M1023_s
+ N_A_1198_55#_M1033_d N_A_1198_55#_c_832_n N_A_1198_55#_M1008_g
+ N_A_1198_55#_c_838_n N_A_1198_55#_M1039_g N_A_1198_55#_c_833_n
+ N_A_1198_55#_c_840_n N_A_1198_55#_c_834_n N_A_1198_55#_c_841_n
+ N_A_1198_55#_c_842_n N_A_1198_55#_c_835_n N_A_1198_55#_c_836_n
+ N_A_1198_55#_c_837_n PM_SKY130_FD_SC_HS__SDFSTP_1%A_1198_55#
x_PM_SKY130_FD_SC_HS__SDFSTP_1%A_998_81# N_A_998_81#_M1013_d N_A_998_81#_M1014_d
+ N_A_998_81#_c_941_n N_A_998_81#_c_942_n N_A_998_81#_M1033_g
+ N_A_998_81#_c_925_n N_A_998_81#_M1023_g N_A_998_81#_c_943_n
+ N_A_998_81#_M1027_g N_A_998_81#_c_926_n N_A_998_81#_M1000_g
+ N_A_998_81#_c_927_n N_A_998_81#_c_928_n N_A_998_81#_c_929_n
+ N_A_998_81#_c_930_n N_A_998_81#_c_931_n N_A_998_81#_c_932_n
+ N_A_998_81#_c_933_n N_A_998_81#_c_934_n N_A_998_81#_c_945_n
+ N_A_998_81#_c_935_n N_A_998_81#_c_936_n N_A_998_81#_c_937_n
+ N_A_998_81#_c_938_n N_A_998_81#_c_939_n N_A_998_81#_c_940_n
+ PM_SKY130_FD_SC_HS__SDFSTP_1%A_998_81#
x_PM_SKY130_FD_SC_HS__SDFSTP_1%SET_B N_SET_B_c_1103_n N_SET_B_c_1104_n
+ N_SET_B_M1030_g N_SET_B_M1012_g N_SET_B_M1017_g N_SET_B_c_1105_n
+ N_SET_B_c_1106_n N_SET_B_M1036_g N_SET_B_c_1096_n N_SET_B_c_1108_n
+ N_SET_B_c_1097_n N_SET_B_c_1110_n SET_B N_SET_B_c_1099_n N_SET_B_c_1100_n
+ N_SET_B_c_1101_n N_SET_B_c_1102_n PM_SKY130_FD_SC_HS__SDFSTP_1%SET_B
x_PM_SKY130_FD_SC_HS__SDFSTP_1%A_599_74# N_A_599_74#_M1005_s N_A_599_74#_M1032_s
+ N_A_599_74#_M1015_g N_A_599_74#_c_1246_n N_A_599_74#_M1037_g
+ N_A_599_74#_c_1234_n N_A_599_74#_c_1235_n N_A_599_74#_c_1248_n
+ N_A_599_74#_c_1249_n N_A_599_74#_c_1236_n N_A_599_74#_c_1237_n
+ N_A_599_74#_c_1250_n N_A_599_74#_c_1251_n N_A_599_74#_M1013_g
+ N_A_599_74#_c_1252_n N_A_599_74#_c_1253_n N_A_599_74#_c_1254_n
+ N_A_599_74#_M1019_g N_A_599_74#_c_1255_n N_A_599_74#_M1035_g
+ N_A_599_74#_c_1240_n N_A_599_74#_c_1241_n N_A_599_74#_M1022_g
+ N_A_599_74#_c_1258_n N_A_599_74#_c_1259_n N_A_599_74#_c_1260_n
+ N_A_599_74#_c_1261_n N_A_599_74#_c_1242_n N_A_599_74#_c_1243_n
+ N_A_599_74#_c_1263_n N_A_599_74#_c_1264_n N_A_599_74#_c_1244_n
+ N_A_599_74#_c_1245_n PM_SKY130_FD_SC_HS__SDFSTP_1%A_599_74#
x_PM_SKY130_FD_SC_HS__SDFSTP_1%A_1958_48# N_A_1958_48#_M1038_d
+ N_A_1958_48#_M1016_s N_A_1958_48#_c_1423_n N_A_1958_48#_M1007_g
+ N_A_1958_48#_c_1424_n N_A_1958_48#_c_1433_n N_A_1958_48#_M1029_g
+ N_A_1958_48#_c_1434_n N_A_1958_48#_c_1425_n N_A_1958_48#_c_1426_n
+ N_A_1958_48#_c_1435_n N_A_1958_48#_c_1427_n N_A_1958_48#_c_1428_n
+ N_A_1958_48#_c_1429_n N_A_1958_48#_c_1430_n N_A_1958_48#_c_1437_n
+ N_A_1958_48#_c_1431_n PM_SKY130_FD_SC_HS__SDFSTP_1%A_1958_48#
x_PM_SKY130_FD_SC_HS__SDFSTP_1%A_1764_74# N_A_1764_74#_M1001_d
+ N_A_1764_74#_M1009_d N_A_1764_74#_M1036_d N_A_1764_74#_M1038_g
+ N_A_1764_74#_c_1528_n N_A_1764_74#_c_1529_n N_A_1764_74#_c_1530_n
+ N_A_1764_74#_M1016_g N_A_1764_74#_c_1531_n N_A_1764_74#_M1010_g
+ N_A_1764_74#_c_1533_n N_A_1764_74#_M1034_g N_A_1764_74#_c_1521_n
+ N_A_1764_74#_c_1535_n N_A_1764_74#_c_1536_n N_A_1764_74#_c_1537_n
+ N_A_1764_74#_c_1538_n N_A_1764_74#_c_1522_n N_A_1764_74#_c_1523_n
+ N_A_1764_74#_c_1540_n N_A_1764_74#_c_1541_n N_A_1764_74#_c_1542_n
+ N_A_1764_74#_c_1543_n N_A_1764_74#_c_1524_n N_A_1764_74#_c_1525_n
+ N_A_1764_74#_c_1545_n N_A_1764_74#_c_1526_n N_A_1764_74#_c_1527_n
+ N_A_1764_74#_c_1547_n N_A_1764_74#_c_1548_n
+ PM_SKY130_FD_SC_HS__SDFSTP_1%A_1764_74#
x_PM_SKY130_FD_SC_HS__SDFSTP_1%A_2395_94# N_A_2395_94#_M1010_s
+ N_A_2395_94#_M1034_s N_A_2395_94#_c_1674_n N_A_2395_94#_M1018_g
+ N_A_2395_94#_c_1675_n N_A_2395_94#_M1006_g N_A_2395_94#_c_1676_n
+ N_A_2395_94#_c_1682_n N_A_2395_94#_c_1677_n N_A_2395_94#_c_1678_n
+ N_A_2395_94#_c_1689_n N_A_2395_94#_c_1679_n N_A_2395_94#_c_1680_n
+ PM_SKY130_FD_SC_HS__SDFSTP_1%A_2395_94#
x_PM_SKY130_FD_SC_HS__SDFSTP_1%VPWR N_VPWR_M1025_d N_VPWR_M1028_d N_VPWR_M1032_d
+ N_VPWR_M1039_d N_VPWR_M1030_d N_VPWR_M1029_d N_VPWR_M1016_d N_VPWR_M1034_d
+ N_VPWR_c_1735_n N_VPWR_c_1736_n N_VPWR_c_1737_n N_VPWR_c_1738_n
+ N_VPWR_c_1739_n N_VPWR_c_1740_n N_VPWR_c_1741_n N_VPWR_c_1742_n
+ N_VPWR_c_1743_n N_VPWR_c_1744_n N_VPWR_c_1745_n N_VPWR_c_1746_n
+ N_VPWR_c_1747_n N_VPWR_c_1748_n N_VPWR_c_1749_n N_VPWR_c_1750_n
+ N_VPWR_c_1751_n VPWR N_VPWR_c_1752_n N_VPWR_c_1753_n N_VPWR_c_1754_n
+ N_VPWR_c_1755_n N_VPWR_c_1734_n N_VPWR_c_1757_n N_VPWR_c_1758_n
+ N_VPWR_c_1759_n N_VPWR_c_1760_n PM_SKY130_FD_SC_HS__SDFSTP_1%VPWR
x_PM_SKY130_FD_SC_HS__SDFSTP_1%A_289_464# N_A_289_464#_M1026_d
+ N_A_289_464#_M1013_s N_A_289_464#_M1031_d N_A_289_464#_M1014_s
+ N_A_289_464#_c_1907_n N_A_289_464#_c_1896_n N_A_289_464#_c_1897_n
+ N_A_289_464#_c_1898_n N_A_289_464#_c_1899_n N_A_289_464#_c_1903_n
+ N_A_289_464#_c_1900_n N_A_289_464#_c_1928_n N_A_289_464#_c_1981_n
+ N_A_289_464#_c_1901_n N_A_289_464#_c_1905_n N_A_289_464#_c_1906_n
+ PM_SKY130_FD_SC_HS__SDFSTP_1%A_289_464#
x_PM_SKY130_FD_SC_HS__SDFSTP_1%A_1610_341# N_A_1610_341#_M1027_d
+ N_A_1610_341#_M1022_d N_A_1610_341#_c_2026_n N_A_1610_341#_c_2027_n
+ N_A_1610_341#_c_2028_n N_A_1610_341#_c_2029_n
+ PM_SKY130_FD_SC_HS__SDFSTP_1%A_1610_341#
x_PM_SKY130_FD_SC_HS__SDFSTP_1%A_1721_374# N_A_1721_374#_M1009_s
+ N_A_1721_374#_M1029_s N_A_1721_374#_c_2070_n N_A_1721_374#_c_2071_n
+ N_A_1721_374#_c_2072_n PM_SKY130_FD_SC_HS__SDFSTP_1%A_1721_374#
x_PM_SKY130_FD_SC_HS__SDFSTP_1%Q N_Q_M1018_d N_Q_M1006_d Q Q Q Q Q Q Q
+ N_Q_c_2102_n PM_SKY130_FD_SC_HS__SDFSTP_1%Q
x_PM_SKY130_FD_SC_HS__SDFSTP_1%VGND N_VGND_M1021_d N_VGND_M1003_d N_VGND_M1005_d
+ N_VGND_M1008_d N_VGND_M1012_d N_VGND_M1017_d N_VGND_M1010_d N_VGND_c_2117_n
+ N_VGND_c_2118_n N_VGND_c_2119_n N_VGND_c_2120_n N_VGND_c_2121_n
+ N_VGND_c_2122_n N_VGND_c_2123_n N_VGND_c_2124_n N_VGND_c_2125_n
+ N_VGND_c_2126_n N_VGND_c_2127_n N_VGND_c_2128_n N_VGND_c_2129_n
+ N_VGND_c_2130_n N_VGND_c_2131_n VGND N_VGND_c_2132_n N_VGND_c_2133_n
+ N_VGND_c_2134_n N_VGND_c_2135_n N_VGND_c_2136_n N_VGND_c_2137_n
+ N_VGND_c_2138_n PM_SKY130_FD_SC_HS__SDFSTP_1%VGND
cc_1 VNB N_SCE_M1021_g 0.0463948f $X=-0.19 $Y=-0.245 $X2=0.575 $Y2=0.58
cc_2 VNB N_SCE_M1004_g 0.0346073f $X=-0.19 $Y=-0.245 $X2=1.935 $Y2=0.58
cc_3 VNB N_SCE_c_296_n 0.018605f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=1.8
cc_4 VNB N_SCE_c_297_n 0.0283175f $X=-0.19 $Y=-0.245 $X2=1.79 $Y2=1.525
cc_5 VNB N_SCE_c_298_n 0.00282835f $X=-0.19 $Y=-0.245 $X2=1.955 $Y2=1.425
cc_6 VNB N_SCE_c_299_n 0.0310386f $X=-0.19 $Y=-0.245 $X2=1.955 $Y2=1.425
cc_7 VNB SCE 0.00942657f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_8 VNB N_SCE_c_301_n 0.0192919f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=1.445
cc_9 VNB N_A_27_464#_M1002_g 0.0207302f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_27_464#_c_383_n 0.0297558f $X=-0.19 $Y=-0.245 $X2=0.95 $Y2=2.64
cc_11 VNB N_A_27_464#_c_384_n 0.0257186f $X=-0.19 $Y=-0.245 $X2=1.935 $Y2=0.58
cc_12 VNB N_A_27_464#_c_385_n 0.00560691f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=1.875
cc_13 VNB N_A_27_464#_c_386_n 0.0135551f $X=-0.19 $Y=-0.245 $X2=1.917 $Y2=1.525
cc_14 VNB N_A_27_464#_c_387_n 0.00566304f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_27_464#_c_388_n 0.0352197f $X=-0.19 $Y=-0.245 $X2=1.955 $Y2=1.425
cc_16 VNB N_D_M1026_g 0.0617671f $X=-0.19 $Y=-0.245 $X2=0.575 $Y2=1.28
cc_17 VNB N_SCD_c_501_n 0.0179466f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=1.95
cc_18 VNB SCD 0.00602448f $X=-0.19 $Y=-0.245 $X2=0.575 $Y2=0.58
cc_19 VNB N_SCD_c_503_n 0.0560964f $X=-0.19 $Y=-0.245 $X2=0.95 $Y2=2.245
cc_20 VNB N_SCD_c_504_n 0.0258121f $X=-0.19 $Y=-0.245 $X2=0.95 $Y2=2.64
cc_21 VNB N_CLK_c_546_n 0.0206756f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=1.95
cc_22 VNB N_CLK_c_547_n 0.0400053f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=2.64
cc_23 VNB CLK 0.00813745f $X=-0.19 $Y=-0.245 $X2=0.575 $Y2=0.58
cc_24 VNB N_A_800_74#_c_580_n 0.028217f $X=-0.19 $Y=-0.245 $X2=0.575 $Y2=0.58
cc_25 VNB N_A_800_74#_M1011_g 0.0601441f $X=-0.19 $Y=-0.245 $X2=0.95 $Y2=2.245
cc_26 VNB N_A_800_74#_c_582_n 0.0196751f $X=-0.19 $Y=-0.245 $X2=0.95 $Y2=2.64
cc_27 VNB N_A_800_74#_c_583_n 0.0135603f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_800_74#_c_584_n 0.00205227f $X=-0.19 $Y=-0.245 $X2=0.835 $Y2=1.525
cc_29 VNB N_A_800_74#_c_585_n 0.017153f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_800_74#_c_586_n 0.00182933f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_31 VNB N_A_800_74#_c_587_n 0.0039887f $X=-0.19 $Y=-0.245 $X2=1.955 $Y2=1.425
cc_32 VNB N_A_800_74#_c_588_n 0.00215354f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.525
cc_33 VNB N_A_800_74#_c_589_n 0.00546133f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_800_74#_c_590_n 0.00648542f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_800_74#_c_591_n 0.00801137f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_800_74#_c_592_n 0.0065757f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_800_74#_c_593_n 0.00487818f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_800_74#_c_594_n 0.0353129f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_1198_55#_c_832_n 0.0182748f $X=-0.19 $Y=-0.245 $X2=0.575 $Y2=0.58
cc_40 VNB N_A_1198_55#_c_833_n 0.0223302f $X=-0.19 $Y=-0.245 $X2=0.95 $Y2=2.245
cc_41 VNB N_A_1198_55#_c_834_n 0.0055764f $X=-0.19 $Y=-0.245 $X2=1.935 $Y2=1.26
cc_42 VNB N_A_1198_55#_c_835_n 0.00460268f $X=-0.19 $Y=-0.245 $X2=1.955
+ $Y2=1.425
cc_43 VNB N_A_1198_55#_c_836_n 0.00955618f $X=-0.19 $Y=-0.245 $X2=0.515
+ $Y2=1.445
cc_44 VNB N_A_1198_55#_c_837_n 0.0479272f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.525
cc_45 VNB N_A_998_81#_c_925_n 0.0170678f $X=-0.19 $Y=-0.245 $X2=0.95 $Y2=2.245
cc_46 VNB N_A_998_81#_c_926_n 0.0217435f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_998_81#_c_927_n 0.022046f $X=-0.19 $Y=-0.245 $X2=1.79 $Y2=1.525
cc_48 VNB N_A_998_81#_c_928_n 0.00719981f $X=-0.19 $Y=-0.245 $X2=1.917 $Y2=1.525
cc_49 VNB N_A_998_81#_c_929_n 0.0083873f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_50 VNB N_A_998_81#_c_930_n 0.0123286f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_A_998_81#_c_931_n 0.00884798f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=1.445
cc_52 VNB N_A_998_81#_c_932_n 0.00141219f $X=-0.19 $Y=-0.245 $X2=1.955 $Y2=1.26
cc_53 VNB N_A_998_81#_c_933_n 0.00204548f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.445
cc_54 VNB N_A_998_81#_c_934_n 0.0620238f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.525
cc_55 VNB N_A_998_81#_c_935_n 0.00292199f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_A_998_81#_c_936_n 0.012354f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_A_998_81#_c_937_n 0.0050355f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_A_998_81#_c_938_n 0.0148924f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_A_998_81#_c_939_n 0.0184439f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_A_998_81#_c_940_n 0.0136403f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_SET_B_M1012_g 0.0395334f $X=-0.19 $Y=-0.245 $X2=0.575 $Y2=0.58
cc_62 VNB N_SET_B_M1017_g 0.0486142f $X=-0.19 $Y=-0.245 $X2=0.95 $Y2=1.95
cc_63 VNB N_SET_B_c_1096_n 0.00663708f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=1.445
cc_64 VNB N_SET_B_c_1097_n 0.0198309f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=1.8
cc_65 VNB SET_B 9.43259e-19 $X=-0.19 $Y=-0.245 $X2=1.955 $Y2=1.425
cc_66 VNB N_SET_B_c_1099_n 0.0142941f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_SET_B_c_1100_n 0.0151291f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=1.445
cc_68 VNB N_SET_B_c_1101_n 7.89065e-19 $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=1.445
cc_69 VNB N_SET_B_c_1102_n 0.00492784f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.665
cc_70 VNB N_A_599_74#_M1015_g 0.0277354f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_A_599_74#_c_1234_n 0.0104075f $X=-0.19 $Y=-0.245 $X2=0.95 $Y2=2.64
cc_72 VNB N_A_599_74#_c_1235_n 0.0397652f $X=-0.19 $Y=-0.245 $X2=0.95 $Y2=2.64
cc_73 VNB N_A_599_74#_c_1236_n 0.029759f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_A_599_74#_c_1237_n 0.010303f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=1.445
cc_75 VNB N_A_599_74#_M1013_g 0.0272008f $X=-0.19 $Y=-0.245 $X2=0.835 $Y2=1.525
cc_76 VNB N_A_599_74#_M1035_g 0.0519158f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=1.445
cc_77 VNB N_A_599_74#_c_1240_n 0.00967691f $X=-0.19 $Y=-0.245 $X2=1.955 $Y2=1.26
cc_78 VNB N_A_599_74#_c_1241_n 0.0105053f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VNB N_A_599_74#_c_1242_n 0.00794834f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_A_599_74#_c_1243_n 0.0115249f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_81 VNB N_A_599_74#_c_1244_n 0.00127679f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_82 VNB N_A_599_74#_c_1245_n 0.00217364f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_83 VNB N_A_1958_48#_c_1423_n 0.0214478f $X=-0.19 $Y=-0.245 $X2=0.575 $Y2=0.58
cc_84 VNB N_A_1958_48#_c_1424_n 0.0235266f $X=-0.19 $Y=-0.245 $X2=0.68 $Y2=1.875
cc_85 VNB N_A_1958_48#_c_1425_n 0.027047f $X=-0.19 $Y=-0.245 $X2=1.935 $Y2=0.58
cc_86 VNB N_A_1958_48#_c_1426_n 0.0174244f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=1.8
cc_87 VNB N_A_1958_48#_c_1427_n 0.00290066f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_88 VNB N_A_1958_48#_c_1428_n 0.0011848f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_89 VNB N_A_1958_48#_c_1429_n 0.0200994f $X=-0.19 $Y=-0.245 $X2=0.515
+ $Y2=1.445
cc_90 VNB N_A_1958_48#_c_1430_n 0.0124734f $X=-0.19 $Y=-0.245 $X2=0.515
+ $Y2=1.445
cc_91 VNB N_A_1958_48#_c_1431_n 0.0801756f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.445
cc_92 VNB N_A_1764_74#_M1038_g 0.0553638f $X=-0.19 $Y=-0.245 $X2=0.95 $Y2=1.95
cc_93 VNB N_A_1764_74#_M1010_g 0.0492609f $X=-0.19 $Y=-0.245 $X2=1.79 $Y2=1.525
cc_94 VNB N_A_1764_74#_c_1521_n 0.00802345f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_95 VNB N_A_1764_74#_c_1522_n 0.0131473f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.665
cc_96 VNB N_A_1764_74#_c_1523_n 0.00641707f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_97 VNB N_A_1764_74#_c_1524_n 0.0039198f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_98 VNB N_A_1764_74#_c_1525_n 0.0167777f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_99 VNB N_A_1764_74#_c_1526_n 0.00690449f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_100 VNB N_A_1764_74#_c_1527_n 0.00132259f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_101 VNB N_A_2395_94#_c_1674_n 0.0225183f $X=-0.19 $Y=-0.245 $X2=0.575
+ $Y2=0.58
cc_102 VNB N_A_2395_94#_c_1675_n 0.0516645f $X=-0.19 $Y=-0.245 $X2=0.86
+ $Y2=1.875
cc_103 VNB N_A_2395_94#_c_1676_n 0.00171495f $X=-0.19 $Y=-0.245 $X2=1.935
+ $Y2=0.58
cc_104 VNB N_A_2395_94#_c_1677_n 0.0069597f $X=-0.19 $Y=-0.245 $X2=1.917
+ $Y2=1.425
cc_105 VNB N_A_2395_94#_c_1678_n 0.00372599f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_106 VNB N_A_2395_94#_c_1679_n 0.00535858f $X=-0.19 $Y=-0.245 $X2=0.515
+ $Y2=1.445
cc_107 VNB N_A_2395_94#_c_1680_n 0.0017163f $X=-0.19 $Y=-0.245 $X2=0.515
+ $Y2=1.445
cc_108 VNB N_VPWR_c_1734_n 0.581632f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_109 VNB N_A_289_464#_c_1896_n 0.00240191f $X=-0.19 $Y=-0.245 $X2=1.935
+ $Y2=0.58
cc_110 VNB N_A_289_464#_c_1897_n 0.0125962f $X=-0.19 $Y=-0.245 $X2=0.515
+ $Y2=1.445
cc_111 VNB N_A_289_464#_c_1898_n 0.00305822f $X=-0.19 $Y=-0.245 $X2=0.515
+ $Y2=1.28
cc_112 VNB N_A_289_464#_c_1899_n 0.00445618f $X=-0.19 $Y=-0.245 $X2=0.515
+ $Y2=1.875
cc_113 VNB N_A_289_464#_c_1900_n 0.00786979f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_114 VNB N_A_289_464#_c_1901_n 0.00308811f $X=-0.19 $Y=-0.245 $X2=0.63
+ $Y2=1.445
cc_115 VNB Q 0.0093606f $X=-0.19 $Y=-0.245 $X2=0.575 $Y2=0.58
cc_116 VNB Q 0.0310914f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_117 VNB N_Q_c_2102_n 0.0243787f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=1.8
cc_118 VNB N_VGND_c_2117_n 0.0098156f $X=-0.19 $Y=-0.245 $X2=0.835 $Y2=1.525
cc_119 VNB N_VGND_c_2118_n 0.0108557f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_120 VNB N_VGND_c_2119_n 0.00929157f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_121 VNB N_VGND_c_2120_n 0.0176331f $X=-0.19 $Y=-0.245 $X2=1.955 $Y2=1.425
cc_122 VNB N_VGND_c_2121_n 0.0187613f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.525
cc_123 VNB N_VGND_c_2122_n 0.00925226f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_124 VNB N_VGND_c_2123_n 0.0135044f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_125 VNB N_VGND_c_2124_n 0.0401758f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_126 VNB N_VGND_c_2125_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_127 VNB N_VGND_c_2126_n 0.0599553f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_128 VNB N_VGND_c_2127_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_129 VNB N_VGND_c_2128_n 0.0753746f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_130 VNB N_VGND_c_2129_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_131 VNB N_VGND_c_2130_n 0.0479194f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_132 VNB N_VGND_c_2131_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_133 VNB N_VGND_c_2132_n 0.021877f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_134 VNB N_VGND_c_2133_n 0.0304154f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_135 VNB N_VGND_c_2134_n 0.0213543f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_136 VNB N_VGND_c_2135_n 0.802468f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_137 VNB N_VGND_c_2136_n 0.0271854f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_138 VNB N_VGND_c_2137_n 0.00634377f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_139 VNB N_VGND_c_2138_n 0.01616f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_140 VPB N_SCE_c_302_n 0.0118202f $X=-0.19 $Y=1.66 $X2=0.5 $Y2=2.155
cc_141 VPB N_SCE_c_303_n 0.0257096f $X=-0.19 $Y=1.66 $X2=0.5 $Y2=2.245
cc_142 VPB N_SCE_c_304_n 0.0208388f $X=-0.19 $Y=1.66 $X2=0.86 $Y2=1.875
cc_143 VPB N_SCE_c_305_n 0.010552f $X=-0.19 $Y=1.66 $X2=0.95 $Y2=2.155
cc_144 VPB N_SCE_c_306_n 0.02065f $X=-0.19 $Y=1.66 $X2=0.95 $Y2=2.245
cc_145 VPB N_SCE_c_296_n 0.0120846f $X=-0.19 $Y=1.66 $X2=0.515 $Y2=1.8
cc_146 VPB N_SCE_c_308_n 0.0108158f $X=-0.19 $Y=1.66 $X2=0.515 $Y2=1.875
cc_147 VPB SCE 0.00331308f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_148 VPB N_A_27_464#_c_389_n 0.0538563f $X=-0.19 $Y=1.66 $X2=0.68 $Y2=1.875
cc_149 VPB N_A_27_464#_c_384_n 0.0305746f $X=-0.19 $Y=1.66 $X2=1.935 $Y2=0.58
cc_150 VPB N_A_27_464#_c_391_n 0.00358649f $X=-0.19 $Y=1.66 $X2=1.955 $Y2=1.425
cc_151 VPB N_A_27_464#_c_392_n 0.033598f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_152 VPB N_D_c_466_n 0.0508621f $X=-0.19 $Y=1.66 $X2=0.5 $Y2=1.95
cc_153 VPB N_D_M1026_g 0.0120832f $X=-0.19 $Y=1.66 $X2=0.575 $Y2=1.28
cc_154 VPB N_D_c_468_n 0.00809561f $X=-0.19 $Y=1.66 $X2=0.95 $Y2=1.95
cc_155 VPB N_SCD_c_505_n 0.0180284f $X=-0.19 $Y=1.66 $X2=0.5 $Y2=2.64
cc_156 VPB N_SCD_c_506_n 0.032947f $X=-0.19 $Y=1.66 $X2=0.575 $Y2=0.58
cc_157 VPB SCD 0.00307097f $X=-0.19 $Y=1.66 $X2=0.575 $Y2=0.58
cc_158 VPB N_SCD_c_504_n 0.033944f $X=-0.19 $Y=1.66 $X2=0.95 $Y2=2.64
cc_159 VPB N_CLK_c_547_n 0.0247386f $X=-0.19 $Y=1.66 $X2=0.5 $Y2=2.64
cc_160 VPB N_A_800_74#_c_580_n 0.0623157f $X=-0.19 $Y=1.66 $X2=0.575 $Y2=0.58
cc_161 VPB N_A_800_74#_c_583_n 0.00307434f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_162 VPB N_A_800_74#_c_597_n 0.026261f $X=-0.19 $Y=1.66 $X2=0.515 $Y2=1.445
cc_163 VPB N_A_800_74#_c_598_n 0.0224469f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_164 VPB N_A_800_74#_c_599_n 0.00255231f $X=-0.19 $Y=1.66 $X2=0.515 $Y2=1.445
cc_165 VPB N_A_800_74#_c_587_n 0.0017748f $X=-0.19 $Y=1.66 $X2=1.955 $Y2=1.425
cc_166 VPB N_A_800_74#_c_601_n 0.0060661f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_167 VPB N_A_800_74#_c_602_n 0.00353126f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_168 VPB N_A_800_74#_c_603_n 0.0022219f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_169 VPB N_A_800_74#_c_604_n 0.0147183f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_170 VPB N_A_800_74#_c_605_n 0.00268313f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_171 VPB N_A_800_74#_c_606_n 0.00377515f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_172 VPB N_A_800_74#_c_607_n 0.00653425f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_173 VPB N_A_800_74#_c_608_n 5.45154e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_174 VPB N_A_800_74#_c_589_n 0.012091f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_175 VPB N_A_800_74#_c_610_n 0.00121771f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_176 VPB N_A_800_74#_c_611_n 0.0050852f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_177 VPB N_A_800_74#_c_591_n 0.0038037f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_178 VPB N_A_800_74#_c_592_n 0.0121093f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_179 VPB N_A_800_74#_c_593_n 0.0269856f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_180 VPB N_A_1198_55#_c_838_n 0.0583161f $X=-0.19 $Y=1.66 $X2=0.86 $Y2=1.875
cc_181 VPB N_A_1198_55#_c_833_n 0.00572465f $X=-0.19 $Y=1.66 $X2=0.95 $Y2=2.245
cc_182 VPB N_A_1198_55#_c_840_n 0.0157022f $X=-0.19 $Y=1.66 $X2=0.95 $Y2=2.64
cc_183 VPB N_A_1198_55#_c_841_n 0.00322755f $X=-0.19 $Y=1.66 $X2=0.515 $Y2=1.445
cc_184 VPB N_A_1198_55#_c_842_n 0.00344228f $X=-0.19 $Y=1.66 $X2=0.515 $Y2=1.875
cc_185 VPB N_A_998_81#_c_941_n 0.0161802f $X=-0.19 $Y=1.66 $X2=0.575 $Y2=0.58
cc_186 VPB N_A_998_81#_c_942_n 0.0209182f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_187 VPB N_A_998_81#_c_943_n 0.0155009f $X=-0.19 $Y=1.66 $X2=1.935 $Y2=1.26
cc_188 VPB N_A_998_81#_c_934_n 0.00800624f $X=-0.19 $Y=1.66 $X2=0.63 $Y2=1.525
cc_189 VPB N_A_998_81#_c_945_n 0.00447893f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_190 VPB N_A_998_81#_c_935_n 0.00889936f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_191 VPB N_A_998_81#_c_937_n 9.66089e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_192 VPB N_A_998_81#_c_938_n 0.0163809f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_193 VPB N_SET_B_c_1103_n 0.017663f $X=-0.19 $Y=1.66 $X2=0.5 $Y2=2.155
cc_194 VPB N_SET_B_c_1104_n 0.0204031f $X=-0.19 $Y=1.66 $X2=0.5 $Y2=2.245
cc_195 VPB N_SET_B_c_1105_n 0.0206116f $X=-0.19 $Y=1.66 $X2=0.95 $Y2=2.64
cc_196 VPB N_SET_B_c_1106_n 0.0270358f $X=-0.19 $Y=1.66 $X2=0.95 $Y2=2.64
cc_197 VPB N_SET_B_c_1096_n 0.0130413f $X=-0.19 $Y=1.66 $X2=0.515 $Y2=1.445
cc_198 VPB N_SET_B_c_1108_n 0.0135089f $X=-0.19 $Y=1.66 $X2=0.515 $Y2=1.28
cc_199 VPB N_SET_B_c_1097_n 0.00532363f $X=-0.19 $Y=1.66 $X2=0.515 $Y2=1.8
cc_200 VPB N_SET_B_c_1110_n 0.00135275f $X=-0.19 $Y=1.66 $X2=0.515 $Y2=1.875
cc_201 VPB SET_B 7.51643e-19 $X=-0.19 $Y=1.66 $X2=1.955 $Y2=1.425
cc_202 VPB N_SET_B_c_1100_n 0.0217114f $X=-0.19 $Y=1.66 $X2=0.515 $Y2=1.445
cc_203 VPB N_SET_B_c_1101_n 0.00305913f $X=-0.19 $Y=1.66 $X2=0.515 $Y2=1.445
cc_204 VPB N_SET_B_c_1102_n 0.0058464f $X=-0.19 $Y=1.66 $X2=0.63 $Y2=1.665
cc_205 VPB N_A_599_74#_c_1246_n 0.0150929f $X=-0.19 $Y=1.66 $X2=0.68 $Y2=1.875
cc_206 VPB N_A_599_74#_c_1235_n 0.0172467f $X=-0.19 $Y=1.66 $X2=0.95 $Y2=2.64
cc_207 VPB N_A_599_74#_c_1248_n 0.0304814f $X=-0.19 $Y=1.66 $X2=1.935 $Y2=1.26
cc_208 VPB N_A_599_74#_c_1249_n 0.036817f $X=-0.19 $Y=1.66 $X2=1.935 $Y2=0.58
cc_209 VPB N_A_599_74#_c_1250_n 0.0561446f $X=-0.19 $Y=1.66 $X2=0.515 $Y2=1.28
cc_210 VPB N_A_599_74#_c_1251_n 0.0124073f $X=-0.19 $Y=1.66 $X2=0.515 $Y2=1.8
cc_211 VPB N_A_599_74#_c_1252_n 0.00764189f $X=-0.19 $Y=1.66 $X2=1.955 $Y2=1.425
cc_212 VPB N_A_599_74#_c_1253_n 0.0159949f $X=-0.19 $Y=1.66 $X2=1.955 $Y2=1.425
cc_213 VPB N_A_599_74#_c_1254_n 0.0142625f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_214 VPB N_A_599_74#_c_1255_n 0.281038f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_215 VPB N_A_599_74#_c_1241_n 0.00226299f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_216 VPB N_A_599_74#_M1022_g 0.0103322f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_217 VPB N_A_599_74#_c_1258_n 0.0142113f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_218 VPB N_A_599_74#_c_1259_n 0.0089867f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_219 VPB N_A_599_74#_c_1260_n 0.00735577f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_220 VPB N_A_599_74#_c_1261_n 0.0250273f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_221 VPB N_A_599_74#_c_1243_n 0.00353072f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_222 VPB N_A_599_74#_c_1263_n 0.0127604f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_223 VPB N_A_599_74#_c_1264_n 0.00529758f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_224 VPB N_A_599_74#_c_1244_n 0.00154997f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_225 VPB N_A_1958_48#_c_1424_n 0.0362527f $X=-0.19 $Y=1.66 $X2=0.68 $Y2=1.875
cc_226 VPB N_A_1958_48#_c_1433_n 0.0183538f $X=-0.19 $Y=1.66 $X2=0.95 $Y2=1.95
cc_227 VPB N_A_1958_48#_c_1434_n 0.0191211f $X=-0.19 $Y=1.66 $X2=0.95 $Y2=2.64
cc_228 VPB N_A_1958_48#_c_1435_n 0.00821621f $X=-0.19 $Y=1.66 $X2=1.917
+ $Y2=1.425
cc_229 VPB N_A_1958_48#_c_1430_n 0.00438907f $X=-0.19 $Y=1.66 $X2=0.515
+ $Y2=1.445
cc_230 VPB N_A_1958_48#_c_1437_n 0.00424424f $X=-0.19 $Y=1.66 $X2=0.515
+ $Y2=1.445
cc_231 VPB N_A_1764_74#_c_1528_n 0.01924f $X=-0.19 $Y=1.66 $X2=0.95 $Y2=2.245
cc_232 VPB N_A_1764_74#_c_1529_n 0.0214817f $X=-0.19 $Y=1.66 $X2=0.95 $Y2=2.64
cc_233 VPB N_A_1764_74#_c_1530_n 0.0358602f $X=-0.19 $Y=1.66 $X2=0.95 $Y2=2.64
cc_234 VPB N_A_1764_74#_c_1531_n 0.0571373f $X=-0.19 $Y=1.66 $X2=0.515 $Y2=1.445
cc_235 VPB N_A_1764_74#_M1010_g 0.00921161f $X=-0.19 $Y=1.66 $X2=1.79 $Y2=1.525
cc_236 VPB N_A_1764_74#_c_1533_n 0.0172244f $X=-0.19 $Y=1.66 $X2=1.917 $Y2=1.425
cc_237 VPB N_A_1764_74#_c_1521_n 0.00913166f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_238 VPB N_A_1764_74#_c_1535_n 0.0173434f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_239 VPB N_A_1764_74#_c_1536_n 0.0142511f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_240 VPB N_A_1764_74#_c_1537_n 0.0164481f $X=-0.19 $Y=1.66 $X2=0.515 $Y2=1.445
cc_241 VPB N_A_1764_74#_c_1538_n 0.00182726f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_242 VPB N_A_1764_74#_c_1523_n 0.0122696f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_243 VPB N_A_1764_74#_c_1540_n 0.0095607f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_244 VPB N_A_1764_74#_c_1541_n 0.0112967f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_245 VPB N_A_1764_74#_c_1542_n 0.00342968f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_246 VPB N_A_1764_74#_c_1543_n 0.00935552f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_247 VPB N_A_1764_74#_c_1524_n 0.00103751f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_248 VPB N_A_1764_74#_c_1545_n 0.00340406f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_249 VPB N_A_1764_74#_c_1527_n 0.00151413f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_250 VPB N_A_1764_74#_c_1547_n 0.00910443f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_251 VPB N_A_1764_74#_c_1548_n 0.0087065f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_252 VPB N_A_2395_94#_c_1675_n 0.0288043f $X=-0.19 $Y=1.66 $X2=0.86 $Y2=1.875
cc_253 VPB N_A_2395_94#_c_1682_n 0.0147073f $X=-0.19 $Y=1.66 $X2=0.515 $Y2=1.8
cc_254 VPB N_A_2395_94#_c_1680_n 0.00317993f $X=-0.19 $Y=1.66 $X2=0.515
+ $Y2=1.445
cc_255 VPB N_VPWR_c_1735_n 0.00396467f $X=-0.19 $Y=1.66 $X2=1.917 $Y2=1.425
cc_256 VPB N_VPWR_c_1736_n 0.0108081f $X=-0.19 $Y=1.66 $X2=1.917 $Y2=1.525
cc_257 VPB N_VPWR_c_1737_n 0.0193021f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_258 VPB N_VPWR_c_1738_n 0.00396467f $X=-0.19 $Y=1.66 $X2=0.515 $Y2=1.445
cc_259 VPB N_VPWR_c_1739_n 0.00505111f $X=-0.19 $Y=1.66 $X2=0.63 $Y2=1.445
cc_260 VPB N_VPWR_c_1740_n 0.00825927f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_261 VPB N_VPWR_c_1741_n 0.00770537f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_262 VPB N_VPWR_c_1742_n 0.01631f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_263 VPB N_VPWR_c_1743_n 0.0113828f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_264 VPB N_VPWR_c_1744_n 0.0565312f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_265 VPB N_VPWR_c_1745_n 0.00330333f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_266 VPB N_VPWR_c_1746_n 0.0278712f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_267 VPB N_VPWR_c_1747_n 0.00330333f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_268 VPB N_VPWR_c_1748_n 0.066491f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_269 VPB N_VPWR_c_1749_n 0.00324402f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_270 VPB N_VPWR_c_1750_n 0.0349132f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_271 VPB N_VPWR_c_1751_n 0.0047828f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_272 VPB N_VPWR_c_1752_n 0.0176729f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_273 VPB N_VPWR_c_1753_n 0.0458344f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_274 VPB N_VPWR_c_1754_n 0.0204452f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_275 VPB N_VPWR_c_1755_n 0.0178682f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_276 VPB N_VPWR_c_1734_n 0.117281f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_277 VPB N_VPWR_c_1757_n 0.00601644f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_278 VPB N_VPWR_c_1758_n 0.00631651f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_279 VPB N_VPWR_c_1759_n 0.00601644f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_280 VPB N_VPWR_c_1760_n 0.00614589f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_281 VPB N_A_289_464#_c_1899_n 0.00530771f $X=-0.19 $Y=1.66 $X2=0.515
+ $Y2=1.875
cc_282 VPB N_A_289_464#_c_1903_n 0.0108447f $X=-0.19 $Y=1.66 $X2=1.79 $Y2=1.525
cc_283 VPB N_A_289_464#_c_1900_n 0.00433549f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_284 VPB N_A_289_464#_c_1905_n 0.0020854f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_285 VPB N_A_289_464#_c_1906_n 0.0121761f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_286 VPB N_A_1610_341#_c_2026_n 0.00642798f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_287 VPB N_A_1610_341#_c_2027_n 0.0178686f $X=-0.19 $Y=1.66 $X2=0.68 $Y2=1.875
cc_288 VPB N_A_1610_341#_c_2028_n 0.00933115f $X=-0.19 $Y=1.66 $X2=0.95 $Y2=1.95
cc_289 VPB N_A_1610_341#_c_2029_n 0.00340035f $X=-0.19 $Y=1.66 $X2=0.95 $Y2=2.64
cc_290 VPB N_A_1721_374#_c_2070_n 0.0286811f $X=-0.19 $Y=1.66 $X2=0.575 $Y2=0.58
cc_291 VPB N_A_1721_374#_c_2071_n 0.00439198f $X=-0.19 $Y=1.66 $X2=0.68
+ $Y2=1.875
cc_292 VPB N_A_1721_374#_c_2072_n 0.0120766f $X=-0.19 $Y=1.66 $X2=0.95 $Y2=2.245
cc_293 VPB Q 0.0545272f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_294 N_SCE_M1021_g N_A_27_464#_M1002_g 0.0127562f $X=0.575 $Y=0.58 $X2=0 $Y2=0
cc_295 N_SCE_c_298_n N_A_27_464#_c_389_n 9.21434e-19 $X=1.955 $Y=1.425 $X2=0
+ $Y2=0
cc_296 N_SCE_c_299_n N_A_27_464#_c_389_n 0.0191888f $X=1.955 $Y=1.425 $X2=0
+ $Y2=0
cc_297 N_SCE_M1021_g N_A_27_464#_c_383_n 0.0123462f $X=0.575 $Y=0.58 $X2=0 $Y2=0
cc_298 N_SCE_c_302_n N_A_27_464#_c_384_n 0.0104444f $X=0.5 $Y=2.155 $X2=0 $Y2=0
cc_299 N_SCE_M1021_g N_A_27_464#_c_384_n 0.00267154f $X=0.575 $Y=0.58 $X2=0
+ $Y2=0
cc_300 SCE N_A_27_464#_c_384_n 0.0514619f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_301 N_SCE_c_301_n N_A_27_464#_c_384_n 0.0169652f $X=0.515 $Y=1.445 $X2=0
+ $Y2=0
cc_302 N_SCE_c_303_n N_A_27_464#_c_401_n 0.0109094f $X=0.5 $Y=2.245 $X2=0 $Y2=0
cc_303 N_SCE_c_304_n N_A_27_464#_c_401_n 5.37693e-19 $X=0.86 $Y=1.875 $X2=0
+ $Y2=0
cc_304 N_SCE_c_306_n N_A_27_464#_c_401_n 0.0160194f $X=0.95 $Y=2.245 $X2=0 $Y2=0
cc_305 N_SCE_c_308_n N_A_27_464#_c_401_n 0.00105942f $X=0.515 $Y=1.875 $X2=0
+ $Y2=0
cc_306 SCE N_A_27_464#_c_401_n 0.0155689f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_307 N_SCE_M1021_g N_A_27_464#_c_385_n 0.0108485f $X=0.575 $Y=0.58 $X2=0 $Y2=0
cc_308 N_SCE_c_304_n N_A_27_464#_c_385_n 5.08606e-19 $X=0.86 $Y=1.875 $X2=0
+ $Y2=0
cc_309 N_SCE_c_297_n N_A_27_464#_c_385_n 0.00259318f $X=1.79 $Y=1.525 $X2=0
+ $Y2=0
cc_310 SCE N_A_27_464#_c_385_n 0.0199325f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_311 N_SCE_c_301_n N_A_27_464#_c_385_n 2.0866e-19 $X=0.515 $Y=1.445 $X2=0
+ $Y2=0
cc_312 N_SCE_c_298_n N_A_27_464#_c_391_n 0.0175876f $X=1.955 $Y=1.425 $X2=0
+ $Y2=0
cc_313 N_SCE_c_299_n N_A_27_464#_c_391_n 3.072e-19 $X=1.955 $Y=1.425 $X2=0 $Y2=0
cc_314 N_SCE_M1021_g N_A_27_464#_c_386_n 0.00444475f $X=0.575 $Y=0.58 $X2=0
+ $Y2=0
cc_315 SCE N_A_27_464#_c_386_n 0.00879333f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_316 N_SCE_c_301_n N_A_27_464#_c_386_n 0.00419179f $X=0.515 $Y=1.445 $X2=0
+ $Y2=0
cc_317 N_SCE_c_303_n N_A_27_464#_c_392_n 0.00597294f $X=0.5 $Y=2.245 $X2=0 $Y2=0
cc_318 N_SCE_c_308_n N_A_27_464#_c_392_n 3.93953e-19 $X=0.515 $Y=1.875 $X2=0
+ $Y2=0
cc_319 N_SCE_M1021_g N_A_27_464#_c_387_n 8.8179e-19 $X=0.575 $Y=0.58 $X2=0 $Y2=0
cc_320 N_SCE_c_297_n N_A_27_464#_c_387_n 0.0247729f $X=1.79 $Y=1.525 $X2=0 $Y2=0
cc_321 N_SCE_c_298_n N_A_27_464#_c_387_n 2.71085e-19 $X=1.955 $Y=1.425 $X2=0
+ $Y2=0
cc_322 N_SCE_M1021_g N_A_27_464#_c_388_n 0.0179354f $X=0.575 $Y=0.58 $X2=0 $Y2=0
cc_323 N_SCE_c_304_n N_A_27_464#_c_388_n 0.00261864f $X=0.86 $Y=1.875 $X2=0
+ $Y2=0
cc_324 N_SCE_c_297_n N_A_27_464#_c_388_n 0.00182006f $X=1.79 $Y=1.525 $X2=0
+ $Y2=0
cc_325 N_SCE_c_304_n N_D_c_466_n 0.0202955f $X=0.86 $Y=1.875 $X2=-0.19
+ $Y2=-0.245
cc_326 N_SCE_c_305_n N_D_c_466_n 0.00567408f $X=0.95 $Y=2.155 $X2=-0.19
+ $Y2=-0.245
cc_327 N_SCE_c_306_n N_D_c_466_n 0.0400037f $X=0.95 $Y=2.245 $X2=-0.19
+ $Y2=-0.245
cc_328 N_SCE_c_297_n N_D_c_466_n 0.00445723f $X=1.79 $Y=1.525 $X2=-0.19
+ $Y2=-0.245
cc_329 N_SCE_c_304_n N_D_M1026_g 7.44858e-19 $X=0.86 $Y=1.875 $X2=0 $Y2=0
cc_330 N_SCE_M1004_g N_D_M1026_g 0.0288701f $X=1.935 $Y=0.58 $X2=0 $Y2=0
cc_331 N_SCE_c_297_n N_D_M1026_g 0.0164371f $X=1.79 $Y=1.525 $X2=0 $Y2=0
cc_332 N_SCE_c_298_n N_D_M1026_g 0.00136336f $X=1.955 $Y=1.425 $X2=0 $Y2=0
cc_333 N_SCE_c_299_n N_D_M1026_g 0.0212203f $X=1.955 $Y=1.425 $X2=0 $Y2=0
cc_334 SCE N_D_M1026_g 0.00474552f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_335 N_SCE_c_304_n N_D_c_468_n 0.00702109f $X=0.86 $Y=1.875 $X2=0 $Y2=0
cc_336 N_SCE_c_297_n N_D_c_468_n 0.0318724f $X=1.79 $Y=1.525 $X2=0 $Y2=0
cc_337 SCE N_D_c_468_n 0.00808759f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_338 N_SCE_M1004_g N_SCD_c_501_n 0.0399302f $X=1.935 $Y=0.58 $X2=-0.19
+ $Y2=-0.245
cc_339 N_SCE_M1004_g N_SCD_c_503_n 0.00748008f $X=1.935 $Y=0.58 $X2=0 $Y2=0
cc_340 N_SCE_c_298_n N_SCD_c_503_n 2.84458e-19 $X=1.955 $Y=1.425 $X2=0 $Y2=0
cc_341 N_SCE_c_299_n N_SCD_c_503_n 0.0172124f $X=1.955 $Y=1.425 $X2=0 $Y2=0
cc_342 N_SCE_c_303_n N_VPWR_c_1735_n 0.0101271f $X=0.5 $Y=2.245 $X2=0 $Y2=0
cc_343 N_SCE_c_306_n N_VPWR_c_1735_n 0.00946621f $X=0.95 $Y=2.245 $X2=0 $Y2=0
cc_344 N_SCE_c_303_n N_VPWR_c_1752_n 0.00413917f $X=0.5 $Y=2.245 $X2=0 $Y2=0
cc_345 N_SCE_c_306_n N_VPWR_c_1753_n 0.00413917f $X=0.95 $Y=2.245 $X2=0 $Y2=0
cc_346 N_SCE_c_303_n N_VPWR_c_1734_n 0.00417983f $X=0.5 $Y=2.245 $X2=0 $Y2=0
cc_347 N_SCE_c_306_n N_VPWR_c_1734_n 0.00414311f $X=0.95 $Y=2.245 $X2=0 $Y2=0
cc_348 N_SCE_c_306_n N_A_289_464#_c_1907_n 7.12872e-19 $X=0.95 $Y=2.245 $X2=0
+ $Y2=0
cc_349 N_SCE_M1004_g N_A_289_464#_c_1896_n 0.0119647f $X=1.935 $Y=0.58 $X2=0
+ $Y2=0
cc_350 N_SCE_M1004_g N_A_289_464#_c_1897_n 0.0111068f $X=1.935 $Y=0.58 $X2=0
+ $Y2=0
cc_351 N_SCE_c_298_n N_A_289_464#_c_1897_n 0.0115612f $X=1.955 $Y=1.425 $X2=0
+ $Y2=0
cc_352 N_SCE_c_299_n N_A_289_464#_c_1897_n 0.00309472f $X=1.955 $Y=1.425 $X2=0
+ $Y2=0
cc_353 N_SCE_M1004_g N_A_289_464#_c_1898_n 0.00274486f $X=1.935 $Y=0.58 $X2=0
+ $Y2=0
cc_354 N_SCE_c_297_n N_A_289_464#_c_1898_n 0.0118057f $X=1.79 $Y=1.525 $X2=0
+ $Y2=0
cc_355 N_SCE_c_298_n N_A_289_464#_c_1898_n 0.00788548f $X=1.955 $Y=1.425 $X2=0
+ $Y2=0
cc_356 N_SCE_c_299_n N_A_289_464#_c_1898_n 5.46117e-19 $X=1.955 $Y=1.425 $X2=0
+ $Y2=0
cc_357 N_SCE_M1004_g N_A_289_464#_c_1899_n 0.00346458f $X=1.935 $Y=0.58 $X2=0
+ $Y2=0
cc_358 N_SCE_c_298_n N_A_289_464#_c_1899_n 0.0258733f $X=1.955 $Y=1.425 $X2=0
+ $Y2=0
cc_359 N_SCE_c_299_n N_A_289_464#_c_1899_n 0.00217771f $X=1.955 $Y=1.425 $X2=0
+ $Y2=0
cc_360 N_SCE_M1021_g N_VGND_c_2117_n 0.00560918f $X=0.575 $Y=0.58 $X2=0 $Y2=0
cc_361 N_SCE_M1004_g N_VGND_c_2118_n 0.00169331f $X=1.935 $Y=0.58 $X2=0 $Y2=0
cc_362 N_SCE_M1004_g N_VGND_c_2124_n 0.00434272f $X=1.935 $Y=0.58 $X2=0 $Y2=0
cc_363 N_SCE_M1021_g N_VGND_c_2135_n 0.00824991f $X=0.575 $Y=0.58 $X2=0 $Y2=0
cc_364 N_SCE_M1004_g N_VGND_c_2135_n 0.00821077f $X=1.935 $Y=0.58 $X2=0 $Y2=0
cc_365 N_SCE_M1021_g N_VGND_c_2136_n 0.00434272f $X=0.575 $Y=0.58 $X2=0 $Y2=0
cc_366 N_A_27_464#_c_389_n N_D_c_466_n 0.0433856f $X=2 $Y=2.245 $X2=-0.19
+ $Y2=-0.245
cc_367 N_A_27_464#_c_401_n N_D_c_466_n 0.0156036f $X=1.79 $Y=2.405 $X2=-0.19
+ $Y2=-0.245
cc_368 N_A_27_464#_c_391_n N_D_c_466_n 0.00361884f $X=1.955 $Y=1.995 $X2=-0.19
+ $Y2=-0.245
cc_369 N_A_27_464#_M1002_g N_D_M1026_g 0.0355306f $X=1.115 $Y=0.58 $X2=0 $Y2=0
cc_370 N_A_27_464#_c_387_n N_D_M1026_g 0.00167343f $X=1.055 $Y=1.025 $X2=0 $Y2=0
cc_371 N_A_27_464#_c_388_n N_D_M1026_g 0.0203659f $X=1.055 $Y=1.105 $X2=0 $Y2=0
cc_372 N_A_27_464#_c_389_n N_D_c_468_n 0.00111062f $X=2 $Y=2.245 $X2=0 $Y2=0
cc_373 N_A_27_464#_c_401_n N_D_c_468_n 0.0327247f $X=1.79 $Y=2.405 $X2=0 $Y2=0
cc_374 N_A_27_464#_c_391_n N_D_c_468_n 0.020556f $X=1.955 $Y=1.995 $X2=0 $Y2=0
cc_375 N_A_27_464#_c_389_n N_SCD_c_505_n 0.0380188f $X=2 $Y=2.245 $X2=0 $Y2=0
cc_376 N_A_27_464#_c_389_n N_SCD_c_506_n 0.0141771f $X=2 $Y=2.245 $X2=0 $Y2=0
cc_377 N_A_27_464#_c_391_n N_SCD_c_506_n 2.23507e-19 $X=1.955 $Y=1.995 $X2=0
+ $Y2=0
cc_378 N_A_27_464#_c_389_n N_SCD_c_504_n 0.00885359f $X=2 $Y=2.245 $X2=0 $Y2=0
cc_379 N_A_27_464#_c_401_n N_VPWR_M1025_d 0.00455834f $X=1.79 $Y=2.405 $X2=-0.19
+ $Y2=-0.245
cc_380 N_A_27_464#_c_401_n N_VPWR_c_1735_n 0.0168032f $X=1.79 $Y=2.405 $X2=0
+ $Y2=0
cc_381 N_A_27_464#_c_392_n N_VPWR_c_1735_n 0.021643f $X=0.275 $Y=2.465 $X2=0
+ $Y2=0
cc_382 N_A_27_464#_c_392_n N_VPWR_c_1752_n 0.0121815f $X=0.275 $Y=2.465 $X2=0
+ $Y2=0
cc_383 N_A_27_464#_c_389_n N_VPWR_c_1753_n 0.00300876f $X=2 $Y=2.245 $X2=0 $Y2=0
cc_384 N_A_27_464#_c_389_n N_VPWR_c_1734_n 0.00370184f $X=2 $Y=2.245 $X2=0 $Y2=0
cc_385 N_A_27_464#_c_401_n N_VPWR_c_1734_n 0.0242263f $X=1.79 $Y=2.405 $X2=0
+ $Y2=0
cc_386 N_A_27_464#_c_392_n N_VPWR_c_1734_n 0.0100828f $X=0.275 $Y=2.465 $X2=0
+ $Y2=0
cc_387 N_A_27_464#_c_401_n A_205_464# 0.00476675f $X=1.79 $Y=2.405 $X2=-0.19
+ $Y2=-0.245
cc_388 N_A_27_464#_c_401_n N_A_289_464#_M1031_d 0.0134049f $X=1.79 $Y=2.405
+ $X2=0 $Y2=0
cc_389 N_A_27_464#_c_389_n N_A_289_464#_c_1907_n 0.0148646f $X=2 $Y=2.245 $X2=0
+ $Y2=0
cc_390 N_A_27_464#_c_401_n N_A_289_464#_c_1907_n 0.0374179f $X=1.79 $Y=2.405
+ $X2=0 $Y2=0
cc_391 N_A_27_464#_M1002_g N_A_289_464#_c_1896_n 0.00195271f $X=1.115 $Y=0.58
+ $X2=0 $Y2=0
cc_392 N_A_27_464#_c_387_n N_A_289_464#_c_1898_n 0.00693658f $X=1.055 $Y=1.025
+ $X2=0 $Y2=0
cc_393 N_A_27_464#_c_388_n N_A_289_464#_c_1898_n 4.32194e-19 $X=1.055 $Y=1.105
+ $X2=0 $Y2=0
cc_394 N_A_27_464#_c_389_n N_A_289_464#_c_1899_n 0.00764248f $X=2 $Y=2.245 $X2=0
+ $Y2=0
cc_395 N_A_27_464#_c_401_n N_A_289_464#_c_1899_n 0.0133253f $X=1.79 $Y=2.405
+ $X2=0 $Y2=0
cc_396 N_A_27_464#_c_391_n N_A_289_464#_c_1899_n 0.0360394f $X=1.955 $Y=1.995
+ $X2=0 $Y2=0
cc_397 N_A_27_464#_c_389_n N_A_289_464#_c_1928_n 2.73782e-19 $X=2 $Y=2.245 $X2=0
+ $Y2=0
cc_398 N_A_27_464#_M1002_g N_VGND_c_2117_n 0.00366419f $X=1.115 $Y=0.58 $X2=0
+ $Y2=0
cc_399 N_A_27_464#_c_383_n N_VGND_c_2117_n 0.0172589f $X=0.36 $Y=0.58 $X2=0
+ $Y2=0
cc_400 N_A_27_464#_c_385_n N_VGND_c_2117_n 0.0155481f $X=0.89 $Y=1.025 $X2=0
+ $Y2=0
cc_401 N_A_27_464#_c_387_n N_VGND_c_2117_n 0.00919007f $X=1.055 $Y=1.025 $X2=0
+ $Y2=0
cc_402 N_A_27_464#_c_388_n N_VGND_c_2117_n 9.28411e-19 $X=1.055 $Y=1.105 $X2=0
+ $Y2=0
cc_403 N_A_27_464#_M1002_g N_VGND_c_2124_n 0.00461464f $X=1.115 $Y=0.58 $X2=0
+ $Y2=0
cc_404 N_A_27_464#_M1002_g N_VGND_c_2135_n 0.00908175f $X=1.115 $Y=0.58 $X2=0
+ $Y2=0
cc_405 N_A_27_464#_c_383_n N_VGND_c_2135_n 0.016061f $X=0.36 $Y=0.58 $X2=0 $Y2=0
cc_406 N_A_27_464#_c_383_n N_VGND_c_2136_n 0.0194722f $X=0.36 $Y=0.58 $X2=0
+ $Y2=0
cc_407 N_D_c_466_n N_VPWR_c_1735_n 0.0016042f $X=1.37 $Y=2.245 $X2=0 $Y2=0
cc_408 N_D_c_466_n N_VPWR_c_1753_n 0.00445405f $X=1.37 $Y=2.245 $X2=0 $Y2=0
cc_409 N_D_c_466_n N_VPWR_c_1734_n 0.00456649f $X=1.37 $Y=2.245 $X2=0 $Y2=0
cc_410 N_D_c_466_n N_A_289_464#_c_1907_n 0.00888514f $X=1.37 $Y=2.245 $X2=0
+ $Y2=0
cc_411 N_D_M1026_g N_A_289_464#_c_1896_n 0.0122205f $X=1.505 $Y=0.58 $X2=0 $Y2=0
cc_412 N_D_M1026_g N_A_289_464#_c_1898_n 0.00495141f $X=1.505 $Y=0.58 $X2=0
+ $Y2=0
cc_413 N_D_M1026_g N_A_289_464#_c_1899_n 0.00446889f $X=1.505 $Y=0.58 $X2=0
+ $Y2=0
cc_414 N_D_c_468_n N_A_289_464#_c_1899_n 2.55684e-19 $X=1.415 $Y=1.985 $X2=0
+ $Y2=0
cc_415 N_D_M1026_g N_VGND_c_2124_n 0.00434272f $X=1.505 $Y=0.58 $X2=0 $Y2=0
cc_416 N_D_M1026_g N_VGND_c_2135_n 0.00821077f $X=1.505 $Y=0.58 $X2=0 $Y2=0
cc_417 N_SCD_c_503_n N_CLK_c_546_n 0.00160779f $X=2.602 $Y=1.382 $X2=-0.19
+ $Y2=-0.245
cc_418 N_SCD_c_503_n N_CLK_c_547_n 0.00716655f $X=2.602 $Y=1.382 $X2=0 $Y2=0
cc_419 N_SCD_c_504_n N_CLK_c_547_n 0.00657478f $X=2.68 $Y=1.985 $X2=0 $Y2=0
cc_420 N_SCD_c_501_n N_A_599_74#_c_1242_n 0.00370057f $X=2.325 $Y=0.87 $X2=0
+ $Y2=0
cc_421 SCD N_A_599_74#_c_1243_n 0.0499674f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_422 N_SCD_c_503_n N_A_599_74#_c_1243_n 0.00678132f $X=2.602 $Y=1.382 $X2=0
+ $Y2=0
cc_423 SCD N_A_599_74#_c_1264_n 0.0206534f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_424 N_SCD_c_504_n N_A_599_74#_c_1264_n 0.00305239f $X=2.68 $Y=1.985 $X2=0
+ $Y2=0
cc_425 N_SCD_c_503_n N_A_599_74#_c_1245_n 0.0052344f $X=2.602 $Y=1.382 $X2=0
+ $Y2=0
cc_426 N_SCD_c_505_n N_VPWR_c_1736_n 0.00917915f $X=2.42 $Y=2.245 $X2=0 $Y2=0
cc_427 N_SCD_c_505_n N_VPWR_c_1753_n 0.00323217f $X=2.42 $Y=2.245 $X2=0 $Y2=0
cc_428 N_SCD_c_505_n N_VPWR_c_1734_n 0.00411202f $X=2.42 $Y=2.245 $X2=0 $Y2=0
cc_429 N_SCD_c_505_n N_A_289_464#_c_1907_n 2.90607e-19 $X=2.42 $Y=2.245 $X2=0
+ $Y2=0
cc_430 N_SCD_c_501_n N_A_289_464#_c_1896_n 0.00198339f $X=2.325 $Y=0.87 $X2=0
+ $Y2=0
cc_431 N_SCD_c_503_n N_A_289_464#_c_1897_n 0.0160259f $X=2.602 $Y=1.382 $X2=0
+ $Y2=0
cc_432 N_SCD_c_505_n N_A_289_464#_c_1899_n 0.0117162f $X=2.42 $Y=2.245 $X2=0
+ $Y2=0
cc_433 N_SCD_c_506_n N_A_289_464#_c_1899_n 0.00924272f $X=2.602 $Y=2 $X2=0 $Y2=0
cc_434 SCD N_A_289_464#_c_1899_n 0.0704084f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_435 N_SCD_c_503_n N_A_289_464#_c_1899_n 0.00713563f $X=2.602 $Y=1.382 $X2=0
+ $Y2=0
cc_436 N_SCD_c_504_n N_A_289_464#_c_1899_n 0.0163108f $X=2.68 $Y=1.985 $X2=0
+ $Y2=0
cc_437 N_SCD_c_505_n N_A_289_464#_c_1903_n 0.0136435f $X=2.42 $Y=2.245 $X2=0
+ $Y2=0
cc_438 N_SCD_c_506_n N_A_289_464#_c_1903_n 0.00389725f $X=2.602 $Y=2 $X2=0 $Y2=0
cc_439 SCD N_A_289_464#_c_1903_n 0.0114021f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_440 N_SCD_c_505_n N_A_289_464#_c_1928_n 0.012524f $X=2.42 $Y=2.245 $X2=0
+ $Y2=0
cc_441 N_SCD_c_501_n N_VGND_c_2118_n 0.0127161f $X=2.325 $Y=0.87 $X2=0 $Y2=0
cc_442 SCD N_VGND_c_2118_n 0.00683314f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_443 N_SCD_c_503_n N_VGND_c_2118_n 0.00696599f $X=2.602 $Y=1.382 $X2=0 $Y2=0
cc_444 N_SCD_c_501_n N_VGND_c_2124_n 0.00383152f $X=2.325 $Y=0.87 $X2=0 $Y2=0
cc_445 N_SCD_c_501_n N_VGND_c_2135_n 0.0075725f $X=2.325 $Y=0.87 $X2=0 $Y2=0
cc_446 N_CLK_c_546_n N_A_800_74#_c_584_n 6.66341e-19 $X=3.355 $Y=1.22 $X2=0
+ $Y2=0
cc_447 N_CLK_c_546_n N_A_599_74#_M1015_g 0.0209385f $X=3.355 $Y=1.22 $X2=0 $Y2=0
cc_448 N_CLK_c_547_n N_A_599_74#_M1015_g 0.0143265f $X=3.515 $Y=1.765 $X2=0
+ $Y2=0
cc_449 CLK N_A_599_74#_M1015_g 0.00542511f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_450 N_CLK_c_547_n N_A_599_74#_c_1246_n 0.0403776f $X=3.515 $Y=1.765 $X2=0
+ $Y2=0
cc_451 N_CLK_c_547_n N_A_599_74#_c_1235_n 0.0133518f $X=3.515 $Y=1.765 $X2=0
+ $Y2=0
cc_452 CLK N_A_599_74#_c_1235_n 3.59763e-19 $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_453 N_CLK_c_546_n N_A_599_74#_c_1242_n 0.00571692f $X=3.355 $Y=1.22 $X2=0
+ $Y2=0
cc_454 N_CLK_c_546_n N_A_599_74#_c_1243_n 0.00514607f $X=3.355 $Y=1.22 $X2=0
+ $Y2=0
cc_455 N_CLK_c_547_n N_A_599_74#_c_1243_n 0.00840616f $X=3.515 $Y=1.765 $X2=0
+ $Y2=0
cc_456 CLK N_A_599_74#_c_1243_n 0.0281662f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_457 N_CLK_c_547_n N_A_599_74#_c_1263_n 0.0167884f $X=3.515 $Y=1.765 $X2=0
+ $Y2=0
cc_458 CLK N_A_599_74#_c_1263_n 0.021989f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_459 N_CLK_c_547_n N_A_599_74#_c_1244_n 0.00266154f $X=3.515 $Y=1.765 $X2=0
+ $Y2=0
cc_460 CLK N_A_599_74#_c_1244_n 0.0160701f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_461 N_CLK_c_546_n N_A_599_74#_c_1245_n 0.00282765f $X=3.355 $Y=1.22 $X2=0
+ $Y2=0
cc_462 N_CLK_c_547_n N_VPWR_c_1736_n 0.00646829f $X=3.515 $Y=1.765 $X2=0 $Y2=0
cc_463 N_CLK_c_547_n N_VPWR_c_1737_n 0.00413917f $X=3.515 $Y=1.765 $X2=0 $Y2=0
cc_464 N_CLK_c_547_n N_VPWR_c_1738_n 0.0211242f $X=3.515 $Y=1.765 $X2=0 $Y2=0
cc_465 N_CLK_c_547_n N_VPWR_c_1734_n 0.00822528f $X=3.515 $Y=1.765 $X2=0 $Y2=0
cc_466 N_CLK_c_547_n N_A_289_464#_c_1905_n 0.0151682f $X=3.515 $Y=1.765 $X2=0
+ $Y2=0
cc_467 N_CLK_c_546_n N_VGND_c_2118_n 0.00341885f $X=3.355 $Y=1.22 $X2=0 $Y2=0
cc_468 N_CLK_c_546_n N_VGND_c_2119_n 0.0072585f $X=3.355 $Y=1.22 $X2=0 $Y2=0
cc_469 N_CLK_c_547_n N_VGND_c_2119_n 8.76711e-19 $X=3.515 $Y=1.765 $X2=0 $Y2=0
cc_470 CLK N_VGND_c_2119_n 0.0203996f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_471 N_CLK_c_546_n N_VGND_c_2132_n 0.00434272f $X=3.355 $Y=1.22 $X2=0 $Y2=0
cc_472 N_CLK_c_546_n N_VGND_c_2135_n 0.00826311f $X=3.355 $Y=1.22 $X2=0 $Y2=0
cc_473 N_A_800_74#_M1011_g N_A_1198_55#_c_832_n 0.0416609f $X=5.675 $Y=0.615
+ $X2=0 $Y2=0
cc_474 N_A_800_74#_c_601_n N_A_1198_55#_c_838_n 0.00866774f $X=5.76 $Y=2.345
+ $X2=0 $Y2=0
cc_475 N_A_800_74#_c_602_n N_A_1198_55#_c_838_n 0.00501742f $X=5.76 $Y=2.895
+ $X2=0 $Y2=0
cc_476 N_A_800_74#_c_619_p N_A_1198_55#_c_838_n 0.0124844f $X=6.645 $Y=2.43
+ $X2=0 $Y2=0
cc_477 N_A_800_74#_c_603_n N_A_1198_55#_c_838_n 0.00288342f $X=6.73 $Y=2.895
+ $X2=0 $Y2=0
cc_478 N_A_800_74#_c_611_n N_A_1198_55#_c_838_n 8.96868e-19 $X=5.615 $Y=1.78
+ $X2=0 $Y2=0
cc_479 N_A_800_74#_c_593_n N_A_1198_55#_c_838_n 0.00939204f $X=5.675 $Y=1.78
+ $X2=0 $Y2=0
cc_480 N_A_800_74#_c_611_n N_A_1198_55#_c_833_n 4.71005e-19 $X=5.615 $Y=1.78
+ $X2=0 $Y2=0
cc_481 N_A_800_74#_c_593_n N_A_1198_55#_c_833_n 0.00312148f $X=5.675 $Y=1.78
+ $X2=0 $Y2=0
cc_482 N_A_800_74#_c_619_p N_A_1198_55#_c_840_n 0.03315f $X=6.645 $Y=2.43 $X2=0
+ $Y2=0
cc_483 N_A_800_74#_c_606_n N_A_1198_55#_c_840_n 0.00278944f $X=7.41 $Y=2.895
+ $X2=0 $Y2=0
cc_484 N_A_800_74#_c_608_n N_A_1198_55#_c_840_n 0.0119127f $X=7.495 $Y=2.055
+ $X2=0 $Y2=0
cc_485 N_A_800_74#_c_619_p N_A_1198_55#_c_841_n 0.0133617f $X=6.645 $Y=2.43
+ $X2=0 $Y2=0
cc_486 N_A_800_74#_c_603_n N_A_1198_55#_c_841_n 0.0147353f $X=6.73 $Y=2.895
+ $X2=0 $Y2=0
cc_487 N_A_800_74#_c_604_n N_A_1198_55#_c_841_n 0.0133613f $X=7.325 $Y=2.98
+ $X2=0 $Y2=0
cc_488 N_A_800_74#_c_606_n N_A_1198_55#_c_841_n 0.0387111f $X=7.41 $Y=2.895
+ $X2=0 $Y2=0
cc_489 N_A_800_74#_c_601_n N_A_1198_55#_c_842_n 0.0172478f $X=5.76 $Y=2.345
+ $X2=0 $Y2=0
cc_490 N_A_800_74#_c_619_p N_A_1198_55#_c_842_n 0.0229228f $X=6.645 $Y=2.43
+ $X2=0 $Y2=0
cc_491 N_A_800_74#_c_611_n N_A_1198_55#_c_842_n 0.011929f $X=5.615 $Y=1.78 $X2=0
+ $Y2=0
cc_492 N_A_800_74#_M1011_g N_A_1198_55#_c_835_n 0.00182235f $X=5.675 $Y=0.615
+ $X2=0 $Y2=0
cc_493 N_A_800_74#_M1011_g N_A_1198_55#_c_837_n 0.00961436f $X=5.675 $Y=0.615
+ $X2=0 $Y2=0
cc_494 N_A_800_74#_c_585_n N_A_998_81#_M1013_d 2.28826e-19 $X=5.035 $Y=0.34
+ $X2=-0.19 $Y2=-0.245
cc_495 N_A_800_74#_c_588_n N_A_998_81#_M1013_d 0.00542902f $X=5.12 $Y=0.935
+ $X2=-0.19 $Y2=-0.245
cc_496 N_A_800_74#_c_608_n N_A_998_81#_c_941_n 2.72515e-19 $X=7.495 $Y=2.055
+ $X2=0 $Y2=0
cc_497 N_A_800_74#_c_619_p N_A_998_81#_c_942_n 0.00665945f $X=6.645 $Y=2.43
+ $X2=0 $Y2=0
cc_498 N_A_800_74#_c_603_n N_A_998_81#_c_942_n 0.00933479f $X=6.73 $Y=2.895
+ $X2=0 $Y2=0
cc_499 N_A_800_74#_c_604_n N_A_998_81#_c_942_n 0.00220266f $X=7.325 $Y=2.98
+ $X2=0 $Y2=0
cc_500 N_A_800_74#_c_606_n N_A_998_81#_c_942_n 5.13915e-19 $X=7.41 $Y=2.895
+ $X2=0 $Y2=0
cc_501 N_A_800_74#_c_606_n N_A_998_81#_c_943_n 0.00223878f $X=7.41 $Y=2.895
+ $X2=0 $Y2=0
cc_502 N_A_800_74#_c_607_n N_A_998_81#_c_943_n 0.00687625f $X=7.775 $Y=2.055
+ $X2=0 $Y2=0
cc_503 N_A_800_74#_c_646_p N_A_998_81#_c_943_n 0.00992602f $X=7.86 $Y=1.97 $X2=0
+ $Y2=0
cc_504 N_A_800_74#_c_589_n N_A_998_81#_c_943_n 0.00859808f $X=8.67 $Y=1.665
+ $X2=0 $Y2=0
cc_505 N_A_800_74#_c_610_n N_A_998_81#_c_943_n 0.00156287f $X=7.945 $Y=1.665
+ $X2=0 $Y2=0
cc_506 N_A_800_74#_c_582_n N_A_998_81#_c_926_n 0.0316178f $X=8.745 $Y=1.12 $X2=0
+ $Y2=0
cc_507 N_A_800_74#_M1011_g N_A_998_81#_c_928_n 0.0240557f $X=5.675 $Y=0.615
+ $X2=0 $Y2=0
cc_508 N_A_800_74#_c_585_n N_A_998_81#_c_928_n 0.00340526f $X=5.035 $Y=0.34
+ $X2=0 $Y2=0
cc_509 N_A_800_74#_c_587_n N_A_998_81#_c_928_n 0.00785173f $X=4.905 $Y=1.565
+ $X2=0 $Y2=0
cc_510 N_A_800_74#_c_588_n N_A_998_81#_c_928_n 0.0384131f $X=5.12 $Y=0.935 $X2=0
+ $Y2=0
cc_511 N_A_800_74#_c_590_n N_A_998_81#_c_928_n 0.0140238f $X=5.12 $Y=1.02 $X2=0
+ $Y2=0
cc_512 N_A_800_74#_M1011_g N_A_998_81#_c_929_n 0.0110534f $X=5.675 $Y=0.615
+ $X2=0 $Y2=0
cc_513 N_A_800_74#_c_611_n N_A_998_81#_c_929_n 0.00581005f $X=5.615 $Y=1.78
+ $X2=0 $Y2=0
cc_514 N_A_800_74#_c_593_n N_A_998_81#_c_929_n 7.26027e-19 $X=5.675 $Y=1.78
+ $X2=0 $Y2=0
cc_515 N_A_800_74#_c_580_n N_A_998_81#_c_930_n 5.55528e-19 $X=5.065 $Y=2.21
+ $X2=0 $Y2=0
cc_516 N_A_800_74#_M1011_g N_A_998_81#_c_930_n 0.00418906f $X=5.675 $Y=0.615
+ $X2=0 $Y2=0
cc_517 N_A_800_74#_c_587_n N_A_998_81#_c_930_n 0.0142704f $X=4.905 $Y=1.565
+ $X2=0 $Y2=0
cc_518 N_A_800_74#_c_590_n N_A_998_81#_c_930_n 0.00225903f $X=5.12 $Y=1.02 $X2=0
+ $Y2=0
cc_519 N_A_800_74#_c_611_n N_A_998_81#_c_930_n 0.0159608f $X=5.615 $Y=1.78 $X2=0
+ $Y2=0
cc_520 N_A_800_74#_c_592_n N_A_998_81#_c_930_n 0.00635901f $X=5.45 $Y=1.78 $X2=0
+ $Y2=0
cc_521 N_A_800_74#_c_610_n N_A_998_81#_c_932_n 0.0125464f $X=7.945 $Y=1.665
+ $X2=0 $Y2=0
cc_522 N_A_800_74#_c_589_n N_A_998_81#_c_933_n 0.0323341f $X=8.67 $Y=1.665 $X2=0
+ $Y2=0
cc_523 N_A_800_74#_c_591_n N_A_998_81#_c_933_n 0.0174856f $X=8.835 $Y=1.285
+ $X2=0 $Y2=0
cc_524 N_A_800_74#_c_594_n N_A_998_81#_c_933_n 3.65e-19 $X=8.945 $Y=1.285 $X2=0
+ $Y2=0
cc_525 N_A_800_74#_c_607_n N_A_998_81#_c_934_n 2.57581e-19 $X=7.775 $Y=2.055
+ $X2=0 $Y2=0
cc_526 N_A_800_74#_c_589_n N_A_998_81#_c_934_n 0.0128095f $X=8.67 $Y=1.665 $X2=0
+ $Y2=0
cc_527 N_A_800_74#_c_610_n N_A_998_81#_c_934_n 0.00456332f $X=7.945 $Y=1.665
+ $X2=0 $Y2=0
cc_528 N_A_800_74#_c_591_n N_A_998_81#_c_934_n 0.00357473f $X=8.835 $Y=1.285
+ $X2=0 $Y2=0
cc_529 N_A_800_74#_c_594_n N_A_998_81#_c_934_n 0.0316178f $X=8.945 $Y=1.285
+ $X2=0 $Y2=0
cc_530 N_A_800_74#_c_598_n N_A_998_81#_c_945_n 0.0254316f $X=5.675 $Y=2.98 $X2=0
+ $Y2=0
cc_531 N_A_800_74#_c_601_n N_A_998_81#_c_945_n 0.00371663f $X=5.76 $Y=2.345
+ $X2=0 $Y2=0
cc_532 N_A_800_74#_c_602_n N_A_998_81#_c_945_n 0.00859454f $X=5.76 $Y=2.895
+ $X2=0 $Y2=0
cc_533 N_A_800_74#_c_592_n N_A_998_81#_c_945_n 0.00286705f $X=5.45 $Y=1.78 $X2=0
+ $Y2=0
cc_534 N_A_800_74#_c_593_n N_A_998_81#_c_945_n 0.00151223f $X=5.675 $Y=1.78
+ $X2=0 $Y2=0
cc_535 N_A_800_74#_c_580_n N_A_998_81#_c_935_n 0.013507f $X=5.065 $Y=2.21 $X2=0
+ $Y2=0
cc_536 N_A_800_74#_M1011_g N_A_998_81#_c_935_n 0.00172059f $X=5.675 $Y=0.615
+ $X2=0 $Y2=0
cc_537 N_A_800_74#_c_587_n N_A_998_81#_c_935_n 0.0449923f $X=4.905 $Y=1.565
+ $X2=0 $Y2=0
cc_538 N_A_800_74#_c_601_n N_A_998_81#_c_935_n 0.0151612f $X=5.76 $Y=2.345 $X2=0
+ $Y2=0
cc_539 N_A_800_74#_c_611_n N_A_998_81#_c_935_n 0.0239806f $X=5.615 $Y=1.78 $X2=0
+ $Y2=0
cc_540 N_A_800_74#_c_592_n N_A_998_81#_c_935_n 0.0122968f $X=5.45 $Y=1.78 $X2=0
+ $Y2=0
cc_541 N_A_800_74#_c_593_n N_A_998_81#_c_935_n 0.00130548f $X=5.675 $Y=1.78
+ $X2=0 $Y2=0
cc_542 N_A_800_74#_M1011_g N_A_998_81#_c_936_n 0.00214522f $X=5.675 $Y=0.615
+ $X2=0 $Y2=0
cc_543 N_A_800_74#_c_607_n N_A_998_81#_c_939_n 0.00248073f $X=7.775 $Y=2.055
+ $X2=0 $Y2=0
cc_544 N_A_800_74#_c_608_n N_SET_B_c_1103_n 0.00584181f $X=7.495 $Y=2.055 $X2=0
+ $Y2=0
cc_545 N_A_800_74#_c_646_p N_SET_B_c_1103_n 0.00237034f $X=7.86 $Y=1.97 $X2=0
+ $Y2=0
cc_546 N_A_800_74#_c_603_n N_SET_B_c_1104_n 4.2076e-19 $X=6.73 $Y=2.895 $X2=0
+ $Y2=0
cc_547 N_A_800_74#_c_604_n N_SET_B_c_1104_n 0.00294494f $X=7.325 $Y=2.98 $X2=0
+ $Y2=0
cc_548 N_A_800_74#_c_606_n N_SET_B_c_1104_n 0.0175183f $X=7.41 $Y=2.895 $X2=0
+ $Y2=0
cc_549 N_A_800_74#_c_608_n N_SET_B_c_1104_n 6.26731e-19 $X=7.495 $Y=2.055 $X2=0
+ $Y2=0
cc_550 N_A_800_74#_c_583_n N_SET_B_c_1097_n 0.00530545f $X=8.945 $Y=1.705 $X2=0
+ $Y2=0
cc_551 N_A_800_74#_c_597_n N_SET_B_c_1097_n 0.0034234f $X=8.945 $Y=1.795 $X2=0
+ $Y2=0
cc_552 N_A_800_74#_c_607_n N_SET_B_c_1097_n 0.00541562f $X=7.775 $Y=2.055 $X2=0
+ $Y2=0
cc_553 N_A_800_74#_c_589_n N_SET_B_c_1097_n 0.0418279f $X=8.67 $Y=1.665 $X2=0
+ $Y2=0
cc_554 N_A_800_74#_c_610_n N_SET_B_c_1097_n 0.0103963f $X=7.945 $Y=1.665 $X2=0
+ $Y2=0
cc_555 N_A_800_74#_c_591_n N_SET_B_c_1097_n 0.0189741f $X=8.835 $Y=1.285 $X2=0
+ $Y2=0
cc_556 N_A_800_74#_c_607_n N_SET_B_c_1110_n 0.00140564f $X=7.775 $Y=2.055 $X2=0
+ $Y2=0
cc_557 N_A_800_74#_c_608_n N_SET_B_c_1110_n 0.00134863f $X=7.495 $Y=2.055 $X2=0
+ $Y2=0
cc_558 N_A_800_74#_c_646_p N_SET_B_c_1110_n 8.58547e-19 $X=7.86 $Y=1.97 $X2=0
+ $Y2=0
cc_559 N_A_800_74#_c_610_n N_SET_B_c_1110_n 8.95816e-19 $X=7.945 $Y=1.665 $X2=0
+ $Y2=0
cc_560 N_A_800_74#_c_607_n N_SET_B_c_1100_n 6.84012e-19 $X=7.775 $Y=2.055 $X2=0
+ $Y2=0
cc_561 N_A_800_74#_c_608_n N_SET_B_c_1100_n 0.00312373f $X=7.495 $Y=2.055 $X2=0
+ $Y2=0
cc_562 N_A_800_74#_c_646_p N_SET_B_c_1100_n 8.92125e-19 $X=7.86 $Y=1.97 $X2=0
+ $Y2=0
cc_563 N_A_800_74#_c_610_n N_SET_B_c_1100_n 5.42773e-19 $X=7.945 $Y=1.665 $X2=0
+ $Y2=0
cc_564 N_A_800_74#_c_607_n N_SET_B_c_1101_n 0.00412744f $X=7.775 $Y=2.055 $X2=0
+ $Y2=0
cc_565 N_A_800_74#_c_608_n N_SET_B_c_1101_n 0.0124557f $X=7.495 $Y=2.055 $X2=0
+ $Y2=0
cc_566 N_A_800_74#_c_646_p N_SET_B_c_1101_n 0.00274736f $X=7.86 $Y=1.97 $X2=0
+ $Y2=0
cc_567 N_A_800_74#_c_610_n N_SET_B_c_1101_n 0.00966396f $X=7.945 $Y=1.665 $X2=0
+ $Y2=0
cc_568 N_A_800_74#_c_584_n N_A_599_74#_M1015_g 0.0101255f $X=4.14 $Y=0.515 $X2=0
+ $Y2=0
cc_569 N_A_800_74#_c_586_n N_A_599_74#_M1015_g 0.0046413f $X=4.225 $Y=0.34 $X2=0
+ $Y2=0
cc_570 N_A_800_74#_c_713_p N_A_599_74#_c_1246_n 0.00102022f $X=4.19 $Y=2.78
+ $X2=0 $Y2=0
cc_571 N_A_800_74#_c_599_n N_A_599_74#_c_1246_n 0.00137141f $X=4.275 $Y=2.98
+ $X2=0 $Y2=0
cc_572 N_A_800_74#_c_587_n N_A_599_74#_c_1234_n 0.00121065f $X=4.905 $Y=1.565
+ $X2=0 $Y2=0
cc_573 N_A_800_74#_c_580_n N_A_599_74#_c_1235_n 0.042661f $X=5.065 $Y=2.21 $X2=0
+ $Y2=0
cc_574 N_A_800_74#_c_584_n N_A_599_74#_c_1235_n 0.00137178f $X=4.14 $Y=0.515
+ $X2=0 $Y2=0
cc_575 N_A_800_74#_c_587_n N_A_599_74#_c_1235_n 6.61103e-19 $X=4.905 $Y=1.565
+ $X2=0 $Y2=0
cc_576 N_A_800_74#_c_580_n N_A_599_74#_c_1248_n 0.00516838f $X=5.065 $Y=2.21
+ $X2=0 $Y2=0
cc_577 N_A_800_74#_c_713_p N_A_599_74#_c_1249_n 0.00414441f $X=4.19 $Y=2.78
+ $X2=0 $Y2=0
cc_578 N_A_800_74#_c_598_n N_A_599_74#_c_1249_n 0.0122491f $X=5.675 $Y=2.98
+ $X2=0 $Y2=0
cc_579 N_A_800_74#_c_580_n N_A_599_74#_c_1236_n 0.016576f $X=5.065 $Y=2.21 $X2=0
+ $Y2=0
cc_580 N_A_800_74#_c_587_n N_A_599_74#_c_1236_n 0.00606086f $X=4.905 $Y=1.565
+ $X2=0 $Y2=0
cc_581 N_A_800_74#_c_590_n N_A_599_74#_c_1236_n 0.0045459f $X=5.12 $Y=1.02 $X2=0
+ $Y2=0
cc_582 N_A_800_74#_c_584_n N_A_599_74#_c_1237_n 8.3837e-19 $X=4.14 $Y=0.515
+ $X2=0 $Y2=0
cc_583 N_A_800_74#_c_585_n N_A_599_74#_c_1237_n 0.00171731f $X=5.035 $Y=0.34
+ $X2=0 $Y2=0
cc_584 N_A_800_74#_c_580_n N_A_599_74#_c_1250_n 0.00737233f $X=5.065 $Y=2.21
+ $X2=0 $Y2=0
cc_585 N_A_800_74#_c_598_n N_A_599_74#_c_1250_n 0.0133502f $X=5.675 $Y=2.98
+ $X2=0 $Y2=0
cc_586 N_A_800_74#_M1011_g N_A_599_74#_M1013_g 0.00870034f $X=5.675 $Y=0.615
+ $X2=0 $Y2=0
cc_587 N_A_800_74#_c_584_n N_A_599_74#_M1013_g 0.00267053f $X=4.14 $Y=0.515
+ $X2=0 $Y2=0
cc_588 N_A_800_74#_c_585_n N_A_599_74#_M1013_g 0.0133546f $X=5.035 $Y=0.34 $X2=0
+ $Y2=0
cc_589 N_A_800_74#_c_588_n N_A_599_74#_M1013_g 0.00484065f $X=5.12 $Y=0.935
+ $X2=0 $Y2=0
cc_590 N_A_800_74#_c_590_n N_A_599_74#_M1013_g 0.00787712f $X=5.12 $Y=1.02 $X2=0
+ $Y2=0
cc_591 N_A_800_74#_c_580_n N_A_599_74#_c_1252_n 0.00215536f $X=5.065 $Y=2.21
+ $X2=0 $Y2=0
cc_592 N_A_800_74#_c_602_n N_A_599_74#_c_1252_n 0.00386835f $X=5.76 $Y=2.895
+ $X2=0 $Y2=0
cc_593 N_A_800_74#_c_598_n N_A_599_74#_c_1253_n 0.0185011f $X=5.675 $Y=2.98
+ $X2=0 $Y2=0
cc_594 N_A_800_74#_c_580_n N_A_599_74#_c_1254_n 0.011853f $X=5.065 $Y=2.21 $X2=0
+ $Y2=0
cc_595 N_A_800_74#_c_601_n N_A_599_74#_c_1254_n 0.00166632f $X=5.76 $Y=2.345
+ $X2=0 $Y2=0
cc_596 N_A_800_74#_c_602_n N_A_599_74#_c_1254_n 0.00261594f $X=5.76 $Y=2.895
+ $X2=0 $Y2=0
cc_597 N_A_800_74#_c_611_n N_A_599_74#_c_1254_n 9.63591e-19 $X=5.615 $Y=1.78
+ $X2=0 $Y2=0
cc_598 N_A_800_74#_c_593_n N_A_599_74#_c_1254_n 0.0102932f $X=5.675 $Y=1.78
+ $X2=0 $Y2=0
cc_599 N_A_800_74#_c_597_n N_A_599_74#_c_1255_n 0.00158277f $X=8.945 $Y=1.795
+ $X2=0 $Y2=0
cc_600 N_A_800_74#_c_598_n N_A_599_74#_c_1255_n 0.00463142f $X=5.675 $Y=2.98
+ $X2=0 $Y2=0
cc_601 N_A_800_74#_c_619_p N_A_599_74#_c_1255_n 0.00914224f $X=6.645 $Y=2.43
+ $X2=0 $Y2=0
cc_602 N_A_800_74#_c_604_n N_A_599_74#_c_1255_n 0.0124701f $X=7.325 $Y=2.98
+ $X2=0 $Y2=0
cc_603 N_A_800_74#_c_605_n N_A_599_74#_c_1255_n 0.00297952f $X=6.815 $Y=2.98
+ $X2=0 $Y2=0
cc_604 N_A_800_74#_c_582_n N_A_599_74#_M1035_g 0.0129467f $X=8.745 $Y=1.12 $X2=0
+ $Y2=0
cc_605 N_A_800_74#_c_594_n N_A_599_74#_M1035_g 0.00627896f $X=8.945 $Y=1.285
+ $X2=0 $Y2=0
cc_606 N_A_800_74#_c_583_n N_A_599_74#_c_1240_n 0.00627896f $X=8.945 $Y=1.705
+ $X2=0 $Y2=0
cc_607 N_A_800_74#_c_597_n N_A_599_74#_c_1241_n 0.00627896f $X=8.945 $Y=1.795
+ $X2=0 $Y2=0
cc_608 N_A_800_74#_c_597_n N_A_599_74#_M1022_g 0.0111261f $X=8.945 $Y=1.795
+ $X2=0 $Y2=0
cc_609 N_A_800_74#_c_580_n N_A_599_74#_c_1258_n 0.0113248f $X=5.065 $Y=2.21
+ $X2=0 $Y2=0
cc_610 N_A_800_74#_c_598_n N_A_599_74#_c_1258_n 0.00150742f $X=5.675 $Y=2.98
+ $X2=0 $Y2=0
cc_611 N_A_800_74#_M1037_d N_A_599_74#_c_1263_n 0.0035556f $X=4.04 $Y=1.84 $X2=0
+ $Y2=0
cc_612 N_A_800_74#_c_584_n N_A_599_74#_c_1244_n 0.0174263f $X=4.14 $Y=0.515
+ $X2=0 $Y2=0
cc_613 N_A_800_74#_c_597_n N_A_1764_74#_c_1538_n 0.0106055f $X=8.945 $Y=1.795
+ $X2=0 $Y2=0
cc_614 N_A_800_74#_c_582_n N_A_1764_74#_c_1522_n 0.00236787f $X=8.745 $Y=1.12
+ $X2=0 $Y2=0
cc_615 N_A_800_74#_c_591_n N_A_1764_74#_c_1522_n 0.0278927f $X=8.835 $Y=1.285
+ $X2=0 $Y2=0
cc_616 N_A_800_74#_c_594_n N_A_1764_74#_c_1522_n 0.00362269f $X=8.945 $Y=1.285
+ $X2=0 $Y2=0
cc_617 N_A_800_74#_c_582_n N_A_1764_74#_c_1526_n 0.0212902f $X=8.745 $Y=1.12
+ $X2=0 $Y2=0
cc_618 N_A_800_74#_c_591_n N_A_1764_74#_c_1526_n 0.0136985f $X=8.835 $Y=1.285
+ $X2=0 $Y2=0
cc_619 N_A_800_74#_c_594_n N_A_1764_74#_c_1526_n 0.00283805f $X=8.945 $Y=1.285
+ $X2=0 $Y2=0
cc_620 N_A_800_74#_c_583_n N_A_1764_74#_c_1527_n 0.00247309f $X=8.945 $Y=1.705
+ $X2=0 $Y2=0
cc_621 N_A_800_74#_c_591_n N_A_1764_74#_c_1527_n 0.00692424f $X=8.835 $Y=1.285
+ $X2=0 $Y2=0
cc_622 N_A_800_74#_c_619_p N_VPWR_M1039_d 0.0106053f $X=6.645 $Y=2.43 $X2=0
+ $Y2=0
cc_623 N_A_800_74#_c_603_n N_VPWR_M1039_d 0.00276934f $X=6.73 $Y=2.895 $X2=0
+ $Y2=0
cc_624 N_A_800_74#_c_606_n N_VPWR_M1030_d 0.00402165f $X=7.41 $Y=2.895 $X2=0
+ $Y2=0
cc_625 N_A_800_74#_c_607_n N_VPWR_M1030_d 0.00615897f $X=7.775 $Y=2.055 $X2=0
+ $Y2=0
cc_626 N_A_800_74#_c_646_p N_VPWR_M1030_d 0.0027465f $X=7.86 $Y=1.97 $X2=0 $Y2=0
cc_627 N_A_800_74#_c_610_n N_VPWR_M1030_d 3.16266e-19 $X=7.945 $Y=1.665 $X2=0
+ $Y2=0
cc_628 N_A_800_74#_c_713_p N_VPWR_c_1738_n 0.0204859f $X=4.19 $Y=2.78 $X2=0
+ $Y2=0
cc_629 N_A_800_74#_c_599_n N_VPWR_c_1738_n 0.0125705f $X=4.275 $Y=2.98 $X2=0
+ $Y2=0
cc_630 N_A_800_74#_c_598_n N_VPWR_c_1739_n 0.0084381f $X=5.675 $Y=2.98 $X2=0
+ $Y2=0
cc_631 N_A_800_74#_c_602_n N_VPWR_c_1739_n 0.00923416f $X=5.76 $Y=2.895 $X2=0
+ $Y2=0
cc_632 N_A_800_74#_c_619_p N_VPWR_c_1739_n 0.0196908f $X=6.645 $Y=2.43 $X2=0
+ $Y2=0
cc_633 N_A_800_74#_c_603_n N_VPWR_c_1739_n 0.0159221f $X=6.73 $Y=2.895 $X2=0
+ $Y2=0
cc_634 N_A_800_74#_c_605_n N_VPWR_c_1739_n 0.0146017f $X=6.815 $Y=2.98 $X2=0
+ $Y2=0
cc_635 N_A_800_74#_c_604_n N_VPWR_c_1740_n 0.0147459f $X=7.325 $Y=2.98 $X2=0
+ $Y2=0
cc_636 N_A_800_74#_c_606_n N_VPWR_c_1740_n 0.0442428f $X=7.41 $Y=2.895 $X2=0
+ $Y2=0
cc_637 N_A_800_74#_c_607_n N_VPWR_c_1740_n 0.0155942f $X=7.775 $Y=2.055 $X2=0
+ $Y2=0
cc_638 N_A_800_74#_c_598_n N_VPWR_c_1744_n 0.0953299f $X=5.675 $Y=2.98 $X2=0
+ $Y2=0
cc_639 N_A_800_74#_c_599_n N_VPWR_c_1744_n 0.0111798f $X=4.275 $Y=2.98 $X2=0
+ $Y2=0
cc_640 N_A_800_74#_c_604_n N_VPWR_c_1746_n 0.0423147f $X=7.325 $Y=2.98 $X2=0
+ $Y2=0
cc_641 N_A_800_74#_c_605_n N_VPWR_c_1746_n 0.0115071f $X=6.815 $Y=2.98 $X2=0
+ $Y2=0
cc_642 N_A_800_74#_c_598_n N_VPWR_c_1734_n 0.053125f $X=5.675 $Y=2.98 $X2=0
+ $Y2=0
cc_643 N_A_800_74#_c_599_n N_VPWR_c_1734_n 0.0065196f $X=4.275 $Y=2.98 $X2=0
+ $Y2=0
cc_644 N_A_800_74#_c_619_p N_VPWR_c_1734_n 0.0176797f $X=6.645 $Y=2.43 $X2=0
+ $Y2=0
cc_645 N_A_800_74#_c_604_n N_VPWR_c_1734_n 0.0229174f $X=7.325 $Y=2.98 $X2=0
+ $Y2=0
cc_646 N_A_800_74#_c_605_n N_VPWR_c_1734_n 0.00591013f $X=6.815 $Y=2.98 $X2=0
+ $Y2=0
cc_647 N_A_800_74#_c_585_n N_A_289_464#_M1013_s 0.0023403f $X=5.035 $Y=0.34
+ $X2=0 $Y2=0
cc_648 N_A_800_74#_c_580_n N_A_289_464#_c_1900_n 0.00542355f $X=5.065 $Y=2.21
+ $X2=0 $Y2=0
cc_649 N_A_800_74#_c_584_n N_A_289_464#_c_1900_n 0.0227634f $X=4.14 $Y=0.515
+ $X2=0 $Y2=0
cc_650 N_A_800_74#_c_587_n N_A_289_464#_c_1900_n 0.0708417f $X=4.905 $Y=1.565
+ $X2=0 $Y2=0
cc_651 N_A_800_74#_c_588_n N_A_289_464#_c_1900_n 0.00550965f $X=5.12 $Y=0.935
+ $X2=0 $Y2=0
cc_652 N_A_800_74#_c_590_n N_A_289_464#_c_1900_n 0.0131283f $X=5.12 $Y=1.02
+ $X2=0 $Y2=0
cc_653 N_A_800_74#_c_584_n N_A_289_464#_c_1901_n 0.0114406f $X=4.14 $Y=0.515
+ $X2=0 $Y2=0
cc_654 N_A_800_74#_c_585_n N_A_289_464#_c_1901_n 0.0249427f $X=5.035 $Y=0.34
+ $X2=0 $Y2=0
cc_655 N_A_800_74#_c_590_n N_A_289_464#_c_1901_n 0.0037314f $X=5.12 $Y=1.02
+ $X2=0 $Y2=0
cc_656 N_A_800_74#_M1037_d N_A_289_464#_c_1905_n 0.00520944f $X=4.04 $Y=1.84
+ $X2=0 $Y2=0
cc_657 N_A_800_74#_c_713_p N_A_289_464#_c_1905_n 0.0132996f $X=4.19 $Y=2.78
+ $X2=0 $Y2=0
cc_658 N_A_800_74#_c_598_n N_A_289_464#_c_1905_n 0.00578449f $X=5.675 $Y=2.98
+ $X2=0 $Y2=0
cc_659 N_A_800_74#_c_580_n N_A_289_464#_c_1906_n 0.01044f $X=5.065 $Y=2.21 $X2=0
+ $Y2=0
cc_660 N_A_800_74#_c_713_p N_A_289_464#_c_1906_n 0.0117768f $X=4.19 $Y=2.78
+ $X2=0 $Y2=0
cc_661 N_A_800_74#_c_598_n N_A_289_464#_c_1906_n 0.0417738f $X=5.675 $Y=2.98
+ $X2=0 $Y2=0
cc_662 N_A_800_74#_c_587_n N_A_289_464#_c_1906_n 0.0187789f $X=4.905 $Y=1.565
+ $X2=0 $Y2=0
cc_663 N_A_800_74#_c_601_n A_1128_457# 0.00109788f $X=5.76 $Y=2.345 $X2=-0.19
+ $Y2=-0.245
cc_664 N_A_800_74#_c_602_n A_1128_457# 0.00353079f $X=5.76 $Y=2.895 $X2=-0.19
+ $Y2=-0.245
cc_665 N_A_800_74#_c_619_p A_1128_457# 0.00474497f $X=6.645 $Y=2.43 $X2=-0.19
+ $Y2=-0.245
cc_666 N_A_800_74#_c_809_p A_1128_457# 0.00120442f $X=5.76 $Y=2.43 $X2=-0.19
+ $Y2=-0.245
cc_667 N_A_800_74#_c_589_n N_A_1610_341#_M1027_d 0.0028906f $X=8.67 $Y=1.665
+ $X2=-0.19 $Y2=-0.245
cc_668 N_A_800_74#_c_597_n N_A_1610_341#_c_2026_n 0.0108373f $X=8.945 $Y=1.795
+ $X2=0 $Y2=0
cc_669 N_A_800_74#_c_606_n N_A_1610_341#_c_2026_n 0.00499483f $X=7.41 $Y=2.895
+ $X2=0 $Y2=0
cc_670 N_A_800_74#_c_607_n N_A_1610_341#_c_2026_n 0.0136304f $X=7.775 $Y=2.055
+ $X2=0 $Y2=0
cc_671 N_A_800_74#_c_646_p N_A_1610_341#_c_2026_n 0.00358428f $X=7.86 $Y=1.97
+ $X2=0 $Y2=0
cc_672 N_A_800_74#_c_589_n N_A_1610_341#_c_2026_n 0.0182299f $X=8.67 $Y=1.665
+ $X2=0 $Y2=0
cc_673 N_A_800_74#_c_597_n N_A_1610_341#_c_2027_n 0.0100302f $X=8.945 $Y=1.795
+ $X2=0 $Y2=0
cc_674 N_A_800_74#_c_589_n N_A_1610_341#_c_2027_n 0.00759599f $X=8.67 $Y=1.665
+ $X2=0 $Y2=0
cc_675 N_A_800_74#_c_591_n N_A_1610_341#_c_2027_n 0.00473873f $X=8.835 $Y=1.285
+ $X2=0 $Y2=0
cc_676 N_A_800_74#_c_597_n N_A_1610_341#_c_2029_n 8.15798e-19 $X=8.945 $Y=1.795
+ $X2=0 $Y2=0
cc_677 N_A_800_74#_c_597_n N_A_1721_374#_c_2070_n 3.50003e-19 $X=8.945 $Y=1.795
+ $X2=0 $Y2=0
cc_678 N_A_800_74#_c_586_n N_VGND_c_2119_n 0.011924f $X=4.225 $Y=0.34 $X2=0
+ $Y2=0
cc_679 N_A_800_74#_M1011_g N_VGND_c_2120_n 0.00140857f $X=5.675 $Y=0.615 $X2=0
+ $Y2=0
cc_680 N_A_800_74#_c_582_n N_VGND_c_2121_n 0.00221822f $X=8.745 $Y=1.12 $X2=0
+ $Y2=0
cc_681 N_A_800_74#_M1011_g N_VGND_c_2126_n 0.00527282f $X=5.675 $Y=0.615 $X2=0
+ $Y2=0
cc_682 N_A_800_74#_c_585_n N_VGND_c_2126_n 0.0643073f $X=5.035 $Y=0.34 $X2=0
+ $Y2=0
cc_683 N_A_800_74#_c_586_n N_VGND_c_2126_n 0.0178338f $X=4.225 $Y=0.34 $X2=0
+ $Y2=0
cc_684 N_A_800_74#_c_582_n N_VGND_c_2128_n 0.00434272f $X=8.745 $Y=1.12 $X2=0
+ $Y2=0
cc_685 N_A_800_74#_M1011_g N_VGND_c_2135_n 0.00534666f $X=5.675 $Y=0.615 $X2=0
+ $Y2=0
cc_686 N_A_800_74#_c_582_n N_VGND_c_2135_n 0.00823237f $X=8.745 $Y=1.12 $X2=0
+ $Y2=0
cc_687 N_A_800_74#_c_585_n N_VGND_c_2135_n 0.0370554f $X=5.035 $Y=0.34 $X2=0
+ $Y2=0
cc_688 N_A_800_74#_c_586_n N_VGND_c_2135_n 0.00960503f $X=4.225 $Y=0.34 $X2=0
+ $Y2=0
cc_689 N_A_1198_55#_c_838_n N_A_998_81#_c_941_n 0.00959585f $X=6.08 $Y=2.21
+ $X2=0 $Y2=0
cc_690 N_A_1198_55#_c_840_n N_A_998_81#_c_941_n 0.00717704f $X=6.985 $Y=2.09
+ $X2=0 $Y2=0
cc_691 N_A_1198_55#_c_842_n N_A_998_81#_c_941_n 0.00108968f $X=6.18 $Y=1.96
+ $X2=0 $Y2=0
cc_692 N_A_1198_55#_c_838_n N_A_998_81#_c_942_n 0.0120433f $X=6.08 $Y=2.21 $X2=0
+ $Y2=0
cc_693 N_A_1198_55#_c_840_n N_A_998_81#_c_942_n 0.00719911f $X=6.985 $Y=2.09
+ $X2=0 $Y2=0
cc_694 N_A_1198_55#_c_841_n N_A_998_81#_c_942_n 0.0048688f $X=7.07 $Y=2.495
+ $X2=0 $Y2=0
cc_695 N_A_1198_55#_c_835_n N_A_998_81#_c_925_n 3.06001e-19 $X=6.36 $Y=0.945
+ $X2=0 $Y2=0
cc_696 N_A_1198_55#_c_836_n N_A_998_81#_c_925_n 0.00935872f $X=6.84 $Y=0.8 $X2=0
+ $Y2=0
cc_697 N_A_1198_55#_c_837_n N_A_998_81#_c_925_n 0.00332378f $X=6.27 $Y=1.1 $X2=0
+ $Y2=0
cc_698 N_A_1198_55#_c_835_n N_A_998_81#_c_927_n 7.71548e-19 $X=6.36 $Y=0.945
+ $X2=0 $Y2=0
cc_699 N_A_1198_55#_c_836_n N_A_998_81#_c_927_n 0.00631535f $X=6.84 $Y=0.8 $X2=0
+ $Y2=0
cc_700 N_A_1198_55#_c_837_n N_A_998_81#_c_927_n 0.0108004f $X=6.27 $Y=1.1 $X2=0
+ $Y2=0
cc_701 N_A_1198_55#_c_832_n N_A_998_81#_c_928_n 0.00248725f $X=6.065 $Y=0.935
+ $X2=0 $Y2=0
cc_702 N_A_1198_55#_c_835_n N_A_998_81#_c_928_n 0.0102689f $X=6.36 $Y=0.945
+ $X2=0 $Y2=0
cc_703 N_A_1198_55#_c_837_n N_A_998_81#_c_928_n 3.63752e-19 $X=6.27 $Y=1.1 $X2=0
+ $Y2=0
cc_704 N_A_1198_55#_c_838_n N_A_998_81#_c_931_n 5.27518e-19 $X=6.08 $Y=2.21
+ $X2=0 $Y2=0
cc_705 N_A_1198_55#_c_833_n N_A_998_81#_c_931_n 0.0115491f $X=6.27 $Y=1.795
+ $X2=0 $Y2=0
cc_706 N_A_1198_55#_c_840_n N_A_998_81#_c_931_n 0.0125408f $X=6.985 $Y=2.09
+ $X2=0 $Y2=0
cc_707 N_A_1198_55#_c_834_n N_A_998_81#_c_931_n 0.00685084f $X=6.675 $Y=0.945
+ $X2=0 $Y2=0
cc_708 N_A_1198_55#_c_842_n N_A_998_81#_c_931_n 0.0186632f $X=6.18 $Y=1.96 $X2=0
+ $Y2=0
cc_709 N_A_1198_55#_c_835_n N_A_998_81#_c_931_n 0.0178707f $X=6.36 $Y=0.945
+ $X2=0 $Y2=0
cc_710 N_A_1198_55#_c_837_n N_A_998_81#_c_931_n 0.00471412f $X=6.27 $Y=1.1 $X2=0
+ $Y2=0
cc_711 N_A_1198_55#_c_838_n N_A_998_81#_c_936_n 0.00100091f $X=6.08 $Y=2.21
+ $X2=0 $Y2=0
cc_712 N_A_1198_55#_c_833_n N_A_998_81#_c_936_n 0.00229733f $X=6.27 $Y=1.795
+ $X2=0 $Y2=0
cc_713 N_A_1198_55#_c_842_n N_A_998_81#_c_936_n 0.00393284f $X=6.18 $Y=1.96
+ $X2=0 $Y2=0
cc_714 N_A_1198_55#_c_837_n N_A_998_81#_c_936_n 0.00235485f $X=6.27 $Y=1.1 $X2=0
+ $Y2=0
cc_715 N_A_1198_55#_c_833_n N_A_998_81#_c_937_n 0.00314281f $X=6.27 $Y=1.795
+ $X2=0 $Y2=0
cc_716 N_A_1198_55#_c_840_n N_A_998_81#_c_937_n 0.0218193f $X=6.985 $Y=2.09
+ $X2=0 $Y2=0
cc_717 N_A_1198_55#_c_834_n N_A_998_81#_c_937_n 0.00201556f $X=6.675 $Y=0.945
+ $X2=0 $Y2=0
cc_718 N_A_1198_55#_c_842_n N_A_998_81#_c_937_n 0.0018598f $X=6.18 $Y=1.96 $X2=0
+ $Y2=0
cc_719 N_A_1198_55#_c_835_n N_A_998_81#_c_937_n 0.0049682f $X=6.36 $Y=0.945
+ $X2=0 $Y2=0
cc_720 N_A_1198_55#_c_836_n N_A_998_81#_c_937_n 0.0225526f $X=6.84 $Y=0.8 $X2=0
+ $Y2=0
cc_721 N_A_1198_55#_c_837_n N_A_998_81#_c_937_n 4.13851e-19 $X=6.27 $Y=1.1 $X2=0
+ $Y2=0
cc_722 N_A_1198_55#_c_833_n N_A_998_81#_c_938_n 0.0172093f $X=6.27 $Y=1.795
+ $X2=0 $Y2=0
cc_723 N_A_1198_55#_c_840_n N_A_998_81#_c_938_n 0.00188537f $X=6.985 $Y=2.09
+ $X2=0 $Y2=0
cc_724 N_A_1198_55#_c_834_n N_A_998_81#_c_938_n 3.17845e-19 $X=6.675 $Y=0.945
+ $X2=0 $Y2=0
cc_725 N_A_1198_55#_c_836_n N_A_998_81#_c_938_n 3.09804e-19 $X=6.84 $Y=0.8 $X2=0
+ $Y2=0
cc_726 N_A_1198_55#_c_840_n N_A_998_81#_c_939_n 0.00689216f $X=6.985 $Y=2.09
+ $X2=0 $Y2=0
cc_727 N_A_1198_55#_c_836_n N_A_998_81#_c_939_n 0.00528032f $X=6.84 $Y=0.8 $X2=0
+ $Y2=0
cc_728 N_A_1198_55#_c_833_n N_A_998_81#_c_940_n 0.00599859f $X=6.27 $Y=1.795
+ $X2=0 $Y2=0
cc_729 N_A_1198_55#_c_840_n N_SET_B_c_1103_n 0.00145788f $X=6.985 $Y=2.09 $X2=0
+ $Y2=0
cc_730 N_A_1198_55#_c_841_n N_SET_B_c_1104_n 0.00225137f $X=7.07 $Y=2.495 $X2=0
+ $Y2=0
cc_731 N_A_1198_55#_c_836_n N_SET_B_M1012_g 0.00147235f $X=6.84 $Y=0.8 $X2=0
+ $Y2=0
cc_732 N_A_1198_55#_c_840_n N_SET_B_c_1100_n 2.42105e-19 $X=6.985 $Y=2.09 $X2=0
+ $Y2=0
cc_733 N_A_1198_55#_c_840_n N_SET_B_c_1101_n 7.24365e-19 $X=6.985 $Y=2.09 $X2=0
+ $Y2=0
cc_734 N_A_1198_55#_c_838_n N_A_599_74#_c_1252_n 0.00142457f $X=6.08 $Y=2.21
+ $X2=0 $Y2=0
cc_735 N_A_1198_55#_c_838_n N_A_599_74#_c_1254_n 0.0156838f $X=6.08 $Y=2.21
+ $X2=0 $Y2=0
cc_736 N_A_1198_55#_c_838_n N_A_599_74#_c_1255_n 0.0085954f $X=6.08 $Y=2.21
+ $X2=0 $Y2=0
cc_737 N_A_1198_55#_c_838_n N_VPWR_c_1739_n 0.00202668f $X=6.08 $Y=2.21 $X2=0
+ $Y2=0
cc_738 N_A_1198_55#_c_838_n N_VPWR_c_1734_n 9.49986e-19 $X=6.08 $Y=2.21 $X2=0
+ $Y2=0
cc_739 N_A_1198_55#_c_832_n N_VGND_c_2120_n 0.0112257f $X=6.065 $Y=0.935 $X2=0
+ $Y2=0
cc_740 N_A_1198_55#_c_835_n N_VGND_c_2120_n 0.0175896f $X=6.36 $Y=0.945 $X2=0
+ $Y2=0
cc_741 N_A_1198_55#_c_836_n N_VGND_c_2120_n 0.00809021f $X=6.84 $Y=0.8 $X2=0
+ $Y2=0
cc_742 N_A_1198_55#_c_837_n N_VGND_c_2120_n 0.00418202f $X=6.27 $Y=1.1 $X2=0
+ $Y2=0
cc_743 N_A_1198_55#_c_836_n N_VGND_c_2121_n 0.0133548f $X=6.84 $Y=0.8 $X2=0
+ $Y2=0
cc_744 N_A_1198_55#_c_832_n N_VGND_c_2126_n 0.0045897f $X=6.065 $Y=0.935 $X2=0
+ $Y2=0
cc_745 N_A_1198_55#_c_836_n N_VGND_c_2133_n 0.00737755f $X=6.84 $Y=0.8 $X2=0
+ $Y2=0
cc_746 N_A_1198_55#_c_832_n N_VGND_c_2135_n 0.0044912f $X=6.065 $Y=0.935 $X2=0
+ $Y2=0
cc_747 N_A_1198_55#_c_834_n N_VGND_c_2135_n 0.00662207f $X=6.675 $Y=0.945 $X2=0
+ $Y2=0
cc_748 N_A_1198_55#_c_835_n N_VGND_c_2135_n 0.00197194f $X=6.36 $Y=0.945 $X2=0
+ $Y2=0
cc_749 N_A_1198_55#_c_836_n N_VGND_c_2135_n 0.0102344f $X=6.84 $Y=0.8 $X2=0
+ $Y2=0
cc_750 N_A_998_81#_c_941_n N_SET_B_c_1103_n 0.00773715f $X=6.815 $Y=2.12 $X2=0
+ $Y2=0
cc_751 N_A_998_81#_c_943_n N_SET_B_c_1103_n 0.00671011f $X=7.975 $Y=1.63 $X2=0
+ $Y2=0
cc_752 N_A_998_81#_c_942_n N_SET_B_c_1104_n 0.0147605f $X=6.815 $Y=2.21 $X2=0
+ $Y2=0
cc_753 N_A_998_81#_c_943_n N_SET_B_c_1104_n 0.00740895f $X=7.975 $Y=1.63 $X2=0
+ $Y2=0
cc_754 N_A_998_81#_c_925_n N_SET_B_M1012_g 0.0407573f $X=7.055 $Y=1.09 $X2=0
+ $Y2=0
cc_755 N_A_998_81#_c_932_n N_SET_B_M1012_g 7.58155e-19 $X=7.905 $Y=1.265 $X2=0
+ $Y2=0
cc_756 N_A_998_81#_c_934_n N_SET_B_M1012_g 0.0246954f $X=8.265 $Y=1.285 $X2=0
+ $Y2=0
cc_757 N_A_998_81#_c_937_n N_SET_B_M1012_g 0.00209379f $X=6.792 $Y=1.285 $X2=0
+ $Y2=0
cc_758 N_A_998_81#_c_939_n N_SET_B_M1012_g 0.013397f $X=7.76 $Y=1.265 $X2=0
+ $Y2=0
cc_759 N_A_998_81#_c_940_n N_SET_B_M1012_g 0.00511507f $X=6.77 $Y=1.505 $X2=0
+ $Y2=0
cc_760 N_A_998_81#_c_932_n N_SET_B_c_1097_n 0.00523122f $X=7.905 $Y=1.265 $X2=0
+ $Y2=0
cc_761 N_A_998_81#_c_934_n N_SET_B_c_1097_n 3.67435e-19 $X=8.265 $Y=1.285 $X2=0
+ $Y2=0
cc_762 N_A_998_81#_c_939_n N_SET_B_c_1097_n 0.00505085f $X=7.76 $Y=1.265 $X2=0
+ $Y2=0
cc_763 N_A_998_81#_c_934_n N_SET_B_c_1110_n 4.35473e-19 $X=8.265 $Y=1.285 $X2=0
+ $Y2=0
cc_764 N_A_998_81#_c_937_n N_SET_B_c_1110_n 0.00114135f $X=6.792 $Y=1.285 $X2=0
+ $Y2=0
cc_765 N_A_998_81#_c_939_n N_SET_B_c_1110_n 0.00285173f $X=7.76 $Y=1.265 $X2=0
+ $Y2=0
cc_766 N_A_998_81#_c_943_n N_SET_B_c_1100_n 0.00608765f $X=7.975 $Y=1.63 $X2=0
+ $Y2=0
cc_767 N_A_998_81#_c_937_n N_SET_B_c_1100_n 0.00139743f $X=6.792 $Y=1.285 $X2=0
+ $Y2=0
cc_768 N_A_998_81#_c_938_n N_SET_B_c_1100_n 0.0211517f $X=6.77 $Y=1.67 $X2=0
+ $Y2=0
cc_769 N_A_998_81#_c_939_n N_SET_B_c_1100_n 0.00613036f $X=7.76 $Y=1.265 $X2=0
+ $Y2=0
cc_770 N_A_998_81#_c_940_n N_SET_B_c_1100_n 0.00130643f $X=6.77 $Y=1.505 $X2=0
+ $Y2=0
cc_771 N_A_998_81#_c_943_n N_SET_B_c_1101_n 3.98831e-19 $X=7.975 $Y=1.63 $X2=0
+ $Y2=0
cc_772 N_A_998_81#_c_934_n N_SET_B_c_1101_n 7.4972e-19 $X=8.265 $Y=1.285 $X2=0
+ $Y2=0
cc_773 N_A_998_81#_c_937_n N_SET_B_c_1101_n 0.0152931f $X=6.792 $Y=1.285 $X2=0
+ $Y2=0
cc_774 N_A_998_81#_c_938_n N_SET_B_c_1101_n 8.99015e-19 $X=6.77 $Y=1.67 $X2=0
+ $Y2=0
cc_775 N_A_998_81#_c_939_n N_SET_B_c_1101_n 0.0281284f $X=7.76 $Y=1.265 $X2=0
+ $Y2=0
cc_776 N_A_998_81#_c_928_n N_A_599_74#_c_1236_n 3.52825e-19 $X=5.46 $Y=0.615
+ $X2=0 $Y2=0
cc_777 N_A_998_81#_c_928_n N_A_599_74#_M1013_g 0.00136003f $X=5.46 $Y=0.615
+ $X2=0 $Y2=0
cc_778 N_A_998_81#_c_945_n N_A_599_74#_c_1252_n 4.209e-19 $X=5.34 $Y=2.495 $X2=0
+ $Y2=0
cc_779 N_A_998_81#_c_945_n N_A_599_74#_c_1254_n 0.00563224f $X=5.34 $Y=2.495
+ $X2=0 $Y2=0
cc_780 N_A_998_81#_c_935_n N_A_599_74#_c_1254_n 9.16728e-19 $X=5.34 $Y=2.265
+ $X2=0 $Y2=0
cc_781 N_A_998_81#_c_942_n N_A_599_74#_c_1255_n 0.00739034f $X=6.815 $Y=2.21
+ $X2=0 $Y2=0
cc_782 N_A_998_81#_c_943_n N_A_599_74#_c_1255_n 0.00900015f $X=7.975 $Y=1.63
+ $X2=0 $Y2=0
cc_783 N_A_998_81#_c_926_n N_A_1764_74#_c_1526_n 0.00166343f $X=8.355 $Y=1.12
+ $X2=0 $Y2=0
cc_784 N_A_998_81#_c_942_n N_VPWR_c_1739_n 4.93046e-19 $X=6.815 $Y=2.21 $X2=0
+ $Y2=0
cc_785 N_A_998_81#_c_943_n N_VPWR_c_1740_n 0.00910757f $X=7.975 $Y=1.63 $X2=0
+ $Y2=0
cc_786 N_A_998_81#_c_943_n N_VPWR_c_1734_n 8.6132e-19 $X=7.975 $Y=1.63 $X2=0
+ $Y2=0
cc_787 N_A_998_81#_c_935_n N_A_289_464#_c_1900_n 0.00554858f $X=5.34 $Y=2.265
+ $X2=0 $Y2=0
cc_788 N_A_998_81#_c_935_n N_A_289_464#_c_1906_n 0.0223757f $X=5.34 $Y=2.265
+ $X2=0 $Y2=0
cc_789 N_A_998_81#_c_943_n N_A_1610_341#_c_2026_n 0.00362997f $X=7.975 $Y=1.63
+ $X2=0 $Y2=0
cc_790 N_A_998_81#_c_943_n N_A_1610_341#_c_2028_n 0.00211568f $X=7.975 $Y=1.63
+ $X2=0 $Y2=0
cc_791 N_A_998_81#_c_943_n N_A_1721_374#_c_2072_n 0.00181692f $X=7.975 $Y=1.63
+ $X2=0 $Y2=0
cc_792 N_A_998_81#_c_925_n N_VGND_c_2120_n 0.00307153f $X=7.055 $Y=1.09 $X2=0
+ $Y2=0
cc_793 N_A_998_81#_c_928_n N_VGND_c_2120_n 0.00946137f $X=5.46 $Y=0.615 $X2=0
+ $Y2=0
cc_794 N_A_998_81#_c_925_n N_VGND_c_2121_n 0.00169427f $X=7.055 $Y=1.09 $X2=0
+ $Y2=0
cc_795 N_A_998_81#_c_926_n N_VGND_c_2121_n 0.0158476f $X=8.355 $Y=1.12 $X2=0
+ $Y2=0
cc_796 N_A_998_81#_c_932_n N_VGND_c_2121_n 0.0400007f $X=7.905 $Y=1.265 $X2=0
+ $Y2=0
cc_797 N_A_998_81#_c_934_n N_VGND_c_2121_n 0.0125225f $X=8.265 $Y=1.285 $X2=0
+ $Y2=0
cc_798 N_A_998_81#_c_939_n N_VGND_c_2121_n 0.0158592f $X=7.76 $Y=1.265 $X2=0
+ $Y2=0
cc_799 N_A_998_81#_c_928_n N_VGND_c_2126_n 0.00963155f $X=5.46 $Y=0.615 $X2=0
+ $Y2=0
cc_800 N_A_998_81#_c_926_n N_VGND_c_2128_n 0.00383152f $X=8.355 $Y=1.12 $X2=0
+ $Y2=0
cc_801 N_A_998_81#_c_925_n N_VGND_c_2133_n 0.00417655f $X=7.055 $Y=1.09 $X2=0
+ $Y2=0
cc_802 N_A_998_81#_c_925_n N_VGND_c_2135_n 0.00479212f $X=7.055 $Y=1.09 $X2=0
+ $Y2=0
cc_803 N_A_998_81#_c_926_n N_VGND_c_2135_n 0.0075725f $X=8.355 $Y=1.12 $X2=0
+ $Y2=0
cc_804 N_A_998_81#_c_928_n N_VGND_c_2135_n 0.00894247f $X=5.46 $Y=0.615 $X2=0
+ $Y2=0
cc_805 N_SET_B_c_1104_n N_A_599_74#_c_1255_n 0.00738456f $X=7.295 $Y=2.21 $X2=0
+ $Y2=0
cc_806 N_SET_B_c_1097_n N_A_599_74#_c_1241_n 0.00829212f $X=10.655 $Y=1.665
+ $X2=0 $Y2=0
cc_807 N_SET_B_c_1105_n N_A_1958_48#_c_1424_n 0.00770846f $X=10.94 $Y=2.375
+ $X2=0 $Y2=0
cc_808 N_SET_B_c_1096_n N_A_1958_48#_c_1424_n 0.0320032f $X=10.865 $Y=1.885
+ $X2=0 $Y2=0
cc_809 N_SET_B_c_1097_n N_A_1958_48#_c_1424_n 0.00672379f $X=10.655 $Y=1.665
+ $X2=0 $Y2=0
cc_810 SET_B N_A_1958_48#_c_1424_n 0.00132361f $X=10.715 $Y=1.58 $X2=0 $Y2=0
cc_811 N_SET_B_c_1102_n N_A_1958_48#_c_1424_n 0.00797244f $X=10.8 $Y=1.665 $X2=0
+ $Y2=0
cc_812 N_SET_B_c_1106_n N_A_1958_48#_c_1433_n 0.00867398f $X=10.94 $Y=2.465
+ $X2=0 $Y2=0
cc_813 N_SET_B_c_1105_n N_A_1958_48#_c_1434_n 0.0084548f $X=10.94 $Y=2.375 $X2=0
+ $Y2=0
cc_814 N_SET_B_M1017_g N_A_1958_48#_c_1425_n 0.0172945f $X=10.775 $Y=0.58 $X2=0
+ $Y2=0
cc_815 N_SET_B_c_1097_n N_A_1958_48#_c_1425_n 0.0073669f $X=10.655 $Y=1.665
+ $X2=0 $Y2=0
cc_816 SET_B N_A_1958_48#_c_1425_n 0.00254262f $X=10.715 $Y=1.58 $X2=0 $Y2=0
cc_817 N_SET_B_c_1099_n N_A_1958_48#_c_1425_n 0.00477338f $X=10.865 $Y=1.545
+ $X2=0 $Y2=0
cc_818 N_SET_B_c_1102_n N_A_1958_48#_c_1425_n 0.0263263f $X=10.8 $Y=1.665 $X2=0
+ $Y2=0
cc_819 N_SET_B_M1017_g N_A_1958_48#_c_1426_n 9.3065e-19 $X=10.775 $Y=0.58 $X2=0
+ $Y2=0
cc_820 N_SET_B_c_1106_n N_A_1958_48#_c_1435_n 0.00141534f $X=10.94 $Y=2.465
+ $X2=0 $Y2=0
cc_821 N_SET_B_c_1097_n N_A_1958_48#_c_1427_n 0.0189182f $X=10.655 $Y=1.665
+ $X2=0 $Y2=0
cc_822 N_SET_B_M1017_g N_A_1958_48#_c_1428_n 6.3608e-19 $X=10.775 $Y=0.58 $X2=0
+ $Y2=0
cc_823 N_SET_B_c_1105_n N_A_1958_48#_c_1437_n 4.53641e-19 $X=10.94 $Y=2.375
+ $X2=0 $Y2=0
cc_824 N_SET_B_M1017_g N_A_1958_48#_c_1431_n 0.0320032f $X=10.775 $Y=0.58 $X2=0
+ $Y2=0
cc_825 N_SET_B_c_1097_n N_A_1958_48#_c_1431_n 0.0127068f $X=10.655 $Y=1.665
+ $X2=0 $Y2=0
cc_826 N_SET_B_M1017_g N_A_1764_74#_M1038_g 0.0248374f $X=10.775 $Y=0.58 $X2=0
+ $Y2=0
cc_827 N_SET_B_c_1108_n N_A_1764_74#_c_1529_n 0.0122682f $X=10.865 $Y=2.05 $X2=0
+ $Y2=0
cc_828 N_SET_B_c_1096_n N_A_1764_74#_c_1521_n 0.0122682f $X=10.865 $Y=1.885
+ $X2=0 $Y2=0
cc_829 N_SET_B_c_1097_n N_A_1764_74#_c_1522_n 0.0102706f $X=10.655 $Y=1.665
+ $X2=0 $Y2=0
cc_830 N_SET_B_c_1097_n N_A_1764_74#_c_1523_n 0.0469026f $X=10.655 $Y=1.665
+ $X2=0 $Y2=0
cc_831 SET_B N_A_1764_74#_c_1523_n 0.00117398f $X=10.715 $Y=1.58 $X2=0 $Y2=0
cc_832 N_SET_B_c_1102_n N_A_1764_74#_c_1523_n 0.00473775f $X=10.8 $Y=1.665 $X2=0
+ $Y2=0
cc_833 N_SET_B_c_1102_n N_A_1764_74#_c_1540_n 0.0104575f $X=10.8 $Y=1.665 $X2=0
+ $Y2=0
cc_834 N_SET_B_c_1105_n N_A_1764_74#_c_1541_n 0.00616862f $X=10.94 $Y=2.375
+ $X2=0 $Y2=0
cc_835 N_SET_B_c_1106_n N_A_1764_74#_c_1541_n 0.00684393f $X=10.94 $Y=2.465
+ $X2=0 $Y2=0
cc_836 N_SET_B_c_1108_n N_A_1764_74#_c_1541_n 0.00395407f $X=10.865 $Y=2.05
+ $X2=0 $Y2=0
cc_837 N_SET_B_c_1097_n N_A_1764_74#_c_1541_n 0.0130314f $X=10.655 $Y=1.665
+ $X2=0 $Y2=0
cc_838 SET_B N_A_1764_74#_c_1541_n 0.00216871f $X=10.715 $Y=1.58 $X2=0 $Y2=0
cc_839 N_SET_B_c_1102_n N_A_1764_74#_c_1541_n 0.0236725f $X=10.8 $Y=1.665 $X2=0
+ $Y2=0
cc_840 N_SET_B_c_1106_n N_A_1764_74#_c_1543_n 0.0120075f $X=10.94 $Y=2.465 $X2=0
+ $Y2=0
cc_841 SET_B N_A_1764_74#_c_1524_n 0.00146379f $X=10.715 $Y=1.58 $X2=0 $Y2=0
cc_842 N_SET_B_c_1099_n N_A_1764_74#_c_1524_n 0.00116472f $X=10.865 $Y=1.545
+ $X2=0 $Y2=0
cc_843 N_SET_B_c_1102_n N_A_1764_74#_c_1524_n 0.0524781f $X=10.8 $Y=1.665 $X2=0
+ $Y2=0
cc_844 N_SET_B_c_1099_n N_A_1764_74#_c_1525_n 0.0122682f $X=10.865 $Y=1.545
+ $X2=0 $Y2=0
cc_845 N_SET_B_c_1102_n N_A_1764_74#_c_1525_n 7.37528e-19 $X=10.8 $Y=1.665 $X2=0
+ $Y2=0
cc_846 N_SET_B_c_1105_n N_A_1764_74#_c_1545_n 0.00295726f $X=10.94 $Y=2.375
+ $X2=0 $Y2=0
cc_847 N_SET_B_c_1097_n N_A_1764_74#_c_1527_n 0.0119743f $X=10.655 $Y=1.665
+ $X2=0 $Y2=0
cc_848 N_SET_B_c_1105_n N_A_1764_74#_c_1547_n 0.00406017f $X=10.94 $Y=2.375
+ $X2=0 $Y2=0
cc_849 N_SET_B_c_1106_n N_A_1764_74#_c_1547_n 3.53113e-19 $X=10.94 $Y=2.465
+ $X2=0 $Y2=0
cc_850 N_SET_B_c_1102_n N_A_1764_74#_c_1547_n 0.00252403f $X=10.8 $Y=1.665 $X2=0
+ $Y2=0
cc_851 N_SET_B_c_1096_n N_A_1764_74#_c_1548_n 0.00116472f $X=10.865 $Y=1.885
+ $X2=0 $Y2=0
cc_852 N_SET_B_c_1108_n N_A_1764_74#_c_1548_n 0.00295726f $X=10.865 $Y=2.05
+ $X2=0 $Y2=0
cc_853 N_SET_B_c_1097_n N_VPWR_M1030_d 0.00121062f $X=10.655 $Y=1.665 $X2=0
+ $Y2=0
cc_854 N_SET_B_c_1104_n N_VPWR_c_1740_n 0.0015589f $X=7.295 $Y=2.21 $X2=0 $Y2=0
cc_855 N_SET_B_c_1097_n N_VPWR_c_1740_n 5.40074e-19 $X=10.655 $Y=1.665 $X2=0
+ $Y2=0
cc_856 N_SET_B_c_1106_n N_VPWR_c_1741_n 0.00408025f $X=10.94 $Y=2.465 $X2=0
+ $Y2=0
cc_857 N_SET_B_c_1106_n N_VPWR_c_1750_n 0.00445602f $X=10.94 $Y=2.465 $X2=0
+ $Y2=0
cc_858 N_SET_B_c_1106_n N_VPWR_c_1734_n 0.00900303f $X=10.94 $Y=2.465 $X2=0
+ $Y2=0
cc_859 N_SET_B_c_1097_n N_A_1610_341#_c_2026_n 0.00207987f $X=10.655 $Y=1.665
+ $X2=0 $Y2=0
cc_860 N_SET_B_c_1097_n N_A_1610_341#_c_2027_n 0.011428f $X=10.655 $Y=1.665
+ $X2=0 $Y2=0
cc_861 N_SET_B_c_1097_n N_A_1610_341#_c_2029_n 0.00246007f $X=10.655 $Y=1.665
+ $X2=0 $Y2=0
cc_862 N_SET_B_M1012_g N_VGND_c_2121_n 0.0167388f $X=7.445 $Y=0.8 $X2=0 $Y2=0
cc_863 N_SET_B_M1017_g N_VGND_c_2122_n 0.0278489f $X=10.775 $Y=0.58 $X2=0 $Y2=0
cc_864 N_SET_B_M1017_g N_VGND_c_2128_n 0.00383152f $X=10.775 $Y=0.58 $X2=0 $Y2=0
cc_865 N_SET_B_M1012_g N_VGND_c_2133_n 0.00245125f $X=7.445 $Y=0.8 $X2=0 $Y2=0
cc_866 N_SET_B_M1012_g N_VGND_c_2135_n 0.00274748f $X=7.445 $Y=0.8 $X2=0 $Y2=0
cc_867 N_SET_B_M1017_g N_VGND_c_2135_n 0.00762539f $X=10.775 $Y=0.58 $X2=0 $Y2=0
cc_868 N_A_599_74#_M1035_g N_A_1958_48#_c_1423_n 0.0579151f $X=9.475 $Y=0.58
+ $X2=0 $Y2=0
cc_869 N_A_599_74#_c_1240_n N_A_1958_48#_c_1424_n 0.00623099f $X=9.497 $Y=1.507
+ $X2=0 $Y2=0
cc_870 N_A_599_74#_M1035_g N_A_1958_48#_c_1427_n 0.00117669f $X=9.475 $Y=0.58
+ $X2=0 $Y2=0
cc_871 N_A_599_74#_M1022_g N_A_1764_74#_c_1538_n 0.00478202f $X=9.505 $Y=2.37
+ $X2=0 $Y2=0
cc_872 N_A_599_74#_c_1240_n N_A_1764_74#_c_1522_n 0.0115551f $X=9.497 $Y=1.507
+ $X2=0 $Y2=0
cc_873 N_A_599_74#_c_1241_n N_A_1764_74#_c_1523_n 0.00842342f $X=9.497 $Y=1.698
+ $X2=0 $Y2=0
cc_874 N_A_599_74#_c_1260_n N_A_1764_74#_c_1523_n 0.00891585f $X=9.497 $Y=1.795
+ $X2=0 $Y2=0
cc_875 N_A_599_74#_M1022_g N_A_1764_74#_c_1540_n 0.00368179f $X=9.505 $Y=2.37
+ $X2=0 $Y2=0
cc_876 N_A_599_74#_M1022_g N_A_1764_74#_c_1542_n 4.29783e-19 $X=9.505 $Y=2.37
+ $X2=0 $Y2=0
cc_877 N_A_599_74#_M1035_g N_A_1764_74#_c_1526_n 0.0115551f $X=9.475 $Y=0.58
+ $X2=0 $Y2=0
cc_878 N_A_599_74#_c_1263_n N_VPWR_M1032_d 0.00200574f $X=3.885 $Y=1.945 $X2=0
+ $Y2=0
cc_879 N_A_599_74#_c_1246_n N_VPWR_c_1738_n 0.00766026f $X=3.965 $Y=1.765 $X2=0
+ $Y2=0
cc_880 N_A_599_74#_c_1249_n N_VPWR_c_1738_n 2.85455e-19 $X=4.545 $Y=3.075 $X2=0
+ $Y2=0
cc_881 N_A_599_74#_c_1251_n N_VPWR_c_1738_n 0.00209543f $X=4.62 $Y=3.15 $X2=0
+ $Y2=0
cc_882 N_A_599_74#_c_1253_n N_VPWR_c_1739_n 0.00115529f $X=5.565 $Y=3.075 $X2=0
+ $Y2=0
cc_883 N_A_599_74#_c_1255_n N_VPWR_c_1739_n 0.0209548f $X=9.415 $Y=3.15 $X2=0
+ $Y2=0
cc_884 N_A_599_74#_c_1255_n N_VPWR_c_1740_n 0.0214344f $X=9.415 $Y=3.15 $X2=0
+ $Y2=0
cc_885 N_A_599_74#_c_1246_n N_VPWR_c_1744_n 0.00413917f $X=3.965 $Y=1.765 $X2=0
+ $Y2=0
cc_886 N_A_599_74#_c_1251_n N_VPWR_c_1744_n 0.0430697f $X=4.62 $Y=3.15 $X2=0
+ $Y2=0
cc_887 N_A_599_74#_c_1255_n N_VPWR_c_1746_n 0.0291914f $X=9.415 $Y=3.15 $X2=0
+ $Y2=0
cc_888 N_A_599_74#_c_1255_n N_VPWR_c_1748_n 0.0418256f $X=9.415 $Y=3.15 $X2=0
+ $Y2=0
cc_889 N_A_599_74#_c_1246_n N_VPWR_c_1734_n 0.00818839f $X=3.965 $Y=1.765 $X2=0
+ $Y2=0
cc_890 N_A_599_74#_c_1250_n N_VPWR_c_1734_n 0.0201381f $X=5.475 $Y=3.15 $X2=0
+ $Y2=0
cc_891 N_A_599_74#_c_1251_n N_VPWR_c_1734_n 0.00600709f $X=4.62 $Y=3.15 $X2=0
+ $Y2=0
cc_892 N_A_599_74#_c_1255_n N_VPWR_c_1734_n 0.0901069f $X=9.415 $Y=3.15 $X2=0
+ $Y2=0
cc_893 N_A_599_74#_c_1259_n N_VPWR_c_1734_n 0.00441804f $X=5.565 $Y=3.15 $X2=0
+ $Y2=0
cc_894 N_A_599_74#_c_1261_n N_VPWR_c_1734_n 0.00674811f $X=9.505 $Y=3.15 $X2=0
+ $Y2=0
cc_895 N_A_599_74#_c_1245_n N_A_289_464#_c_1897_n 0.00538292f $X=3.14 $Y=1.01
+ $X2=0 $Y2=0
cc_896 N_A_599_74#_c_1243_n N_A_289_464#_c_1899_n 0.00138544f $X=3.06 $Y=1.82
+ $X2=0 $Y2=0
cc_897 N_A_599_74#_M1032_s N_A_289_464#_c_1903_n 0.00435898f $X=3.145 $Y=1.84
+ $X2=0 $Y2=0
cc_898 N_A_599_74#_c_1263_n N_A_289_464#_c_1903_n 0.00343748f $X=3.885 $Y=1.945
+ $X2=0 $Y2=0
cc_899 N_A_599_74#_c_1264_n N_A_289_464#_c_1903_n 0.00759792f $X=3.145 $Y=1.945
+ $X2=0 $Y2=0
cc_900 N_A_599_74#_M1015_g N_A_289_464#_c_1900_n 0.00165105f $X=3.925 $Y=0.74
+ $X2=0 $Y2=0
cc_901 N_A_599_74#_c_1246_n N_A_289_464#_c_1900_n 0.00118962f $X=3.965 $Y=1.765
+ $X2=0 $Y2=0
cc_902 N_A_599_74#_c_1234_n N_A_289_464#_c_1900_n 0.00614702f $X=4.455 $Y=1.35
+ $X2=0 $Y2=0
cc_903 N_A_599_74#_c_1235_n N_A_289_464#_c_1900_n 0.00986722f $X=4.455 $Y=1.68
+ $X2=0 $Y2=0
cc_904 N_A_599_74#_c_1248_n N_A_289_464#_c_1900_n 0.0132241f $X=4.455 $Y=2.31
+ $X2=0 $Y2=0
cc_905 N_A_599_74#_c_1236_n N_A_289_464#_c_1900_n 0.00684609f $X=4.84 $Y=1.115
+ $X2=0 $Y2=0
cc_906 N_A_599_74#_c_1237_n N_A_289_464#_c_1900_n 0.00443795f $X=4.53 $Y=1.115
+ $X2=0 $Y2=0
cc_907 N_A_599_74#_M1013_g N_A_289_464#_c_1900_n 0.00316996f $X=4.915 $Y=0.615
+ $X2=0 $Y2=0
cc_908 N_A_599_74#_c_1258_n N_A_289_464#_c_1900_n 6.48894e-19 $X=4.545 $Y=2.385
+ $X2=0 $Y2=0
cc_909 N_A_599_74#_c_1263_n N_A_289_464#_c_1900_n 0.0156781f $X=3.885 $Y=1.945
+ $X2=0 $Y2=0
cc_910 N_A_599_74#_c_1244_n N_A_289_464#_c_1900_n 0.0268895f $X=4.05 $Y=1.515
+ $X2=0 $Y2=0
cc_911 N_A_599_74#_M1032_s N_A_289_464#_c_1981_n 0.0153888f $X=3.145 $Y=1.84
+ $X2=0 $Y2=0
cc_912 N_A_599_74#_c_1263_n N_A_289_464#_c_1981_n 0.0118235f $X=3.885 $Y=1.945
+ $X2=0 $Y2=0
cc_913 N_A_599_74#_M1015_g N_A_289_464#_c_1901_n 4.83415e-19 $X=3.925 $Y=0.74
+ $X2=0 $Y2=0
cc_914 N_A_599_74#_c_1236_n N_A_289_464#_c_1901_n 0.00520089f $X=4.84 $Y=1.115
+ $X2=0 $Y2=0
cc_915 N_A_599_74#_c_1237_n N_A_289_464#_c_1901_n 6.03498e-19 $X=4.53 $Y=1.115
+ $X2=0 $Y2=0
cc_916 N_A_599_74#_M1013_g N_A_289_464#_c_1901_n 0.0024395f $X=4.915 $Y=0.615
+ $X2=0 $Y2=0
cc_917 N_A_599_74#_c_1246_n N_A_289_464#_c_1905_n 0.0150499f $X=3.965 $Y=1.765
+ $X2=0 $Y2=0
cc_918 N_A_599_74#_c_1235_n N_A_289_464#_c_1905_n 0.00482991f $X=4.455 $Y=1.68
+ $X2=0 $Y2=0
cc_919 N_A_599_74#_c_1248_n N_A_289_464#_c_1905_n 0.00419091f $X=4.455 $Y=2.31
+ $X2=0 $Y2=0
cc_920 N_A_599_74#_c_1258_n N_A_289_464#_c_1905_n 0.00289641f $X=4.545 $Y=2.385
+ $X2=0 $Y2=0
cc_921 N_A_599_74#_c_1263_n N_A_289_464#_c_1905_n 0.0454795f $X=3.885 $Y=1.945
+ $X2=0 $Y2=0
cc_922 N_A_599_74#_c_1246_n N_A_289_464#_c_1906_n 0.00304778f $X=3.965 $Y=1.765
+ $X2=0 $Y2=0
cc_923 N_A_599_74#_c_1248_n N_A_289_464#_c_1906_n 0.0019469f $X=4.455 $Y=2.31
+ $X2=0 $Y2=0
cc_924 N_A_599_74#_c_1249_n N_A_289_464#_c_1906_n 0.0114214f $X=4.545 $Y=3.075
+ $X2=0 $Y2=0
cc_925 N_A_599_74#_c_1258_n N_A_289_464#_c_1906_n 0.00738559f $X=4.545 $Y=2.385
+ $X2=0 $Y2=0
cc_926 N_A_599_74#_c_1255_n N_A_1610_341#_c_2027_n 0.00597285f $X=9.415 $Y=3.15
+ $X2=0 $Y2=0
cc_927 N_A_599_74#_M1022_g N_A_1610_341#_c_2027_n 0.0200802f $X=9.505 $Y=2.37
+ $X2=0 $Y2=0
cc_928 N_A_599_74#_c_1255_n N_A_1610_341#_c_2028_n 0.00496234f $X=9.415 $Y=3.15
+ $X2=0 $Y2=0
cc_929 N_A_599_74#_M1022_g N_A_1610_341#_c_2029_n 0.00633949f $X=9.505 $Y=2.37
+ $X2=0 $Y2=0
cc_930 N_A_599_74#_c_1255_n N_A_1721_374#_c_2070_n 0.010569f $X=9.415 $Y=3.15
+ $X2=0 $Y2=0
cc_931 N_A_599_74#_M1022_g N_A_1721_374#_c_2070_n 0.00655f $X=9.505 $Y=2.37
+ $X2=0 $Y2=0
cc_932 N_A_599_74#_c_1261_n N_A_1721_374#_c_2070_n 0.0102073f $X=9.505 $Y=3.15
+ $X2=0 $Y2=0
cc_933 N_A_599_74#_M1022_g N_A_1721_374#_c_2071_n 0.0040068f $X=9.505 $Y=2.37
+ $X2=0 $Y2=0
cc_934 N_A_599_74#_c_1255_n N_A_1721_374#_c_2072_n 0.00743665f $X=9.415 $Y=3.15
+ $X2=0 $Y2=0
cc_935 N_A_599_74#_M1022_g N_A_1721_374#_c_2072_n 0.00523797f $X=9.505 $Y=2.37
+ $X2=0 $Y2=0
cc_936 N_A_599_74#_c_1261_n N_A_1721_374#_c_2072_n 2.9957e-19 $X=9.505 $Y=3.15
+ $X2=0 $Y2=0
cc_937 N_A_599_74#_c_1242_n N_VGND_c_2118_n 0.0241477f $X=3.14 $Y=0.515 $X2=0
+ $Y2=0
cc_938 N_A_599_74#_M1015_g N_VGND_c_2119_n 0.00537119f $X=3.925 $Y=0.74 $X2=0
+ $Y2=0
cc_939 N_A_599_74#_c_1242_n N_VGND_c_2119_n 0.0255177f $X=3.14 $Y=0.515 $X2=0
+ $Y2=0
cc_940 N_A_599_74#_M1015_g N_VGND_c_2126_n 0.00430908f $X=3.925 $Y=0.74 $X2=0
+ $Y2=0
cc_941 N_A_599_74#_M1013_g N_VGND_c_2126_n 9.15902e-19 $X=4.915 $Y=0.615 $X2=0
+ $Y2=0
cc_942 N_A_599_74#_M1035_g N_VGND_c_2128_n 0.00461464f $X=9.475 $Y=0.58 $X2=0
+ $Y2=0
cc_943 N_A_599_74#_c_1242_n N_VGND_c_2132_n 0.0145488f $X=3.14 $Y=0.515 $X2=0
+ $Y2=0
cc_944 N_A_599_74#_M1015_g N_VGND_c_2135_n 0.00821709f $X=3.925 $Y=0.74 $X2=0
+ $Y2=0
cc_945 N_A_599_74#_M1035_g N_VGND_c_2135_n 0.00911286f $X=9.475 $Y=0.58 $X2=0
+ $Y2=0
cc_946 N_A_599_74#_c_1242_n N_VGND_c_2135_n 0.0119924f $X=3.14 $Y=0.515 $X2=0
+ $Y2=0
cc_947 N_A_1958_48#_c_1425_n N_A_1764_74#_M1038_g 0.0136598f $X=11.395 $Y=1.095
+ $X2=0 $Y2=0
cc_948 N_A_1958_48#_c_1426_n N_A_1764_74#_M1038_g 0.0142424f $X=11.56 $Y=0.58
+ $X2=0 $Y2=0
cc_949 N_A_1958_48#_c_1429_n N_A_1764_74#_M1038_g 0.00601154f $X=11.395 $Y=0.98
+ $X2=0 $Y2=0
cc_950 N_A_1958_48#_c_1430_n N_A_1764_74#_M1038_g 0.00337861f $X=11.74 $Y=2.22
+ $X2=0 $Y2=0
cc_951 N_A_1958_48#_c_1429_n N_A_1764_74#_c_1528_n 0.00226477f $X=11.395 $Y=0.98
+ $X2=0 $Y2=0
cc_952 N_A_1958_48#_c_1430_n N_A_1764_74#_c_1528_n 0.0103432f $X=11.74 $Y=2.22
+ $X2=0 $Y2=0
cc_953 N_A_1958_48#_c_1437_n N_A_1764_74#_c_1529_n 0.00830212f $X=11.74 $Y=2.39
+ $X2=0 $Y2=0
cc_954 N_A_1958_48#_c_1435_n N_A_1764_74#_c_1530_n 0.0127504f $X=11.705 $Y=2.75
+ $X2=0 $Y2=0
cc_955 N_A_1958_48#_c_1437_n N_A_1764_74#_c_1530_n 0.00858249f $X=11.74 $Y=2.39
+ $X2=0 $Y2=0
cc_956 N_A_1958_48#_c_1430_n N_A_1764_74#_c_1535_n 0.00713398f $X=11.74 $Y=2.22
+ $X2=0 $Y2=0
cc_957 N_A_1958_48#_c_1437_n N_A_1764_74#_c_1535_n 0.0030711f $X=11.74 $Y=2.39
+ $X2=0 $Y2=0
cc_958 N_A_1958_48#_c_1430_n N_A_1764_74#_c_1536_n 0.00940162f $X=11.74 $Y=2.22
+ $X2=0 $Y2=0
cc_959 N_A_1958_48#_c_1427_n N_A_1764_74#_c_1522_n 0.0131299f $X=10.295 $Y=1.145
+ $X2=0 $Y2=0
cc_960 N_A_1958_48#_c_1424_n N_A_1764_74#_c_1523_n 0.00251996f $X=10.385 $Y=2.29
+ $X2=0 $Y2=0
cc_961 N_A_1958_48#_c_1427_n N_A_1764_74#_c_1523_n 0.015616f $X=10.295 $Y=1.145
+ $X2=0 $Y2=0
cc_962 N_A_1958_48#_c_1431_n N_A_1764_74#_c_1523_n 0.00961424f $X=10.385
+ $Y=1.087 $X2=0 $Y2=0
cc_963 N_A_1958_48#_c_1424_n N_A_1764_74#_c_1540_n 0.0128818f $X=10.385 $Y=2.29
+ $X2=0 $Y2=0
cc_964 N_A_1958_48#_c_1424_n N_A_1764_74#_c_1541_n 0.00655896f $X=10.385 $Y=2.29
+ $X2=0 $Y2=0
cc_965 N_A_1958_48#_c_1434_n N_A_1764_74#_c_1541_n 0.0148569f $X=10.385 $Y=2.377
+ $X2=0 $Y2=0
cc_966 N_A_1958_48#_c_1433_n N_A_1764_74#_c_1543_n 5.72855e-19 $X=10.49 $Y=2.465
+ $X2=0 $Y2=0
cc_967 N_A_1958_48#_c_1434_n N_A_1764_74#_c_1543_n 3.64083e-19 $X=10.385
+ $Y=2.377 $X2=0 $Y2=0
cc_968 N_A_1958_48#_c_1435_n N_A_1764_74#_c_1543_n 0.0494732f $X=11.705 $Y=2.75
+ $X2=0 $Y2=0
cc_969 N_A_1958_48#_c_1425_n N_A_1764_74#_c_1524_n 0.0156367f $X=11.395 $Y=1.095
+ $X2=0 $Y2=0
cc_970 N_A_1958_48#_c_1429_n N_A_1764_74#_c_1524_n 0.0180555f $X=11.395 $Y=0.98
+ $X2=0 $Y2=0
cc_971 N_A_1958_48#_c_1430_n N_A_1764_74#_c_1524_n 0.0500166f $X=11.74 $Y=2.22
+ $X2=0 $Y2=0
cc_972 N_A_1958_48#_c_1429_n N_A_1764_74#_c_1525_n 0.00140137f $X=11.395 $Y=0.98
+ $X2=0 $Y2=0
cc_973 N_A_1958_48#_c_1430_n N_A_1764_74#_c_1525_n 0.00915197f $X=11.74 $Y=2.22
+ $X2=0 $Y2=0
cc_974 N_A_1958_48#_c_1430_n N_A_1764_74#_c_1545_n 0.00498176f $X=11.74 $Y=2.22
+ $X2=0 $Y2=0
cc_975 N_A_1958_48#_c_1437_n N_A_1764_74#_c_1547_n 0.015248f $X=11.74 $Y=2.39
+ $X2=0 $Y2=0
cc_976 N_A_1958_48#_c_1437_n N_A_1764_74#_c_1548_n 0.00516543f $X=11.74 $Y=2.39
+ $X2=0 $Y2=0
cc_977 N_A_1958_48#_c_1429_n N_A_2395_94#_c_1676_n 0.00592413f $X=11.395 $Y=0.98
+ $X2=0 $Y2=0
cc_978 N_A_1958_48#_c_1430_n N_A_2395_94#_c_1676_n 3.18868e-19 $X=11.74 $Y=2.22
+ $X2=0 $Y2=0
cc_979 N_A_1958_48#_c_1435_n N_A_2395_94#_c_1682_n 0.00477139f $X=11.705 $Y=2.75
+ $X2=0 $Y2=0
cc_980 N_A_1958_48#_c_1437_n N_A_2395_94#_c_1682_n 0.0124192f $X=11.74 $Y=2.39
+ $X2=0 $Y2=0
cc_981 N_A_1958_48#_c_1426_n N_A_2395_94#_c_1678_n 0.0275804f $X=11.56 $Y=0.58
+ $X2=0 $Y2=0
cc_982 N_A_1958_48#_c_1426_n N_A_2395_94#_c_1689_n 0.00365017f $X=11.56 $Y=0.58
+ $X2=0 $Y2=0
cc_983 N_A_1958_48#_c_1429_n N_A_2395_94#_c_1689_n 8.41437e-19 $X=11.395 $Y=0.98
+ $X2=0 $Y2=0
cc_984 N_A_1958_48#_c_1430_n N_A_2395_94#_c_1679_n 0.0118548f $X=11.74 $Y=2.22
+ $X2=0 $Y2=0
cc_985 N_A_1958_48#_c_1430_n N_A_2395_94#_c_1680_n 0.0124192f $X=11.74 $Y=2.22
+ $X2=0 $Y2=0
cc_986 N_A_1958_48#_c_1433_n N_VPWR_c_1741_n 0.00253053f $X=10.49 $Y=2.465 $X2=0
+ $Y2=0
cc_987 N_A_1958_48#_c_1435_n N_VPWR_c_1742_n 0.028191f $X=11.705 $Y=2.75 $X2=0
+ $Y2=0
cc_988 N_A_1958_48#_c_1433_n N_VPWR_c_1748_n 0.0044313f $X=10.49 $Y=2.465 $X2=0
+ $Y2=0
cc_989 N_A_1958_48#_c_1435_n N_VPWR_c_1750_n 0.0145938f $X=11.705 $Y=2.75 $X2=0
+ $Y2=0
cc_990 N_A_1958_48#_c_1433_n N_VPWR_c_1734_n 0.00858246f $X=10.49 $Y=2.465 $X2=0
+ $Y2=0
cc_991 N_A_1958_48#_c_1434_n N_VPWR_c_1734_n 3.07368e-19 $X=10.385 $Y=2.377
+ $X2=0 $Y2=0
cc_992 N_A_1958_48#_c_1435_n N_VPWR_c_1734_n 0.0120466f $X=11.705 $Y=2.75 $X2=0
+ $Y2=0
cc_993 N_A_1958_48#_c_1433_n N_A_1610_341#_c_2027_n 0.00289959f $X=10.49
+ $Y=2.465 $X2=0 $Y2=0
cc_994 N_A_1958_48#_c_1434_n N_A_1610_341#_c_2027_n 0.00261194f $X=10.385
+ $Y=2.377 $X2=0 $Y2=0
cc_995 N_A_1958_48#_c_1424_n N_A_1610_341#_c_2029_n 9.84231e-19 $X=10.385
+ $Y=2.29 $X2=0 $Y2=0
cc_996 N_A_1958_48#_c_1433_n N_A_1721_374#_c_2070_n 0.00455905f $X=10.49
+ $Y=2.465 $X2=0 $Y2=0
cc_997 N_A_1958_48#_c_1433_n N_A_1721_374#_c_2071_n 0.00399792f $X=10.49
+ $Y=2.465 $X2=0 $Y2=0
cc_998 N_A_1958_48#_c_1434_n N_A_1721_374#_c_2071_n 0.00244865f $X=10.385
+ $Y=2.377 $X2=0 $Y2=0
cc_999 N_A_1958_48#_c_1425_n N_VGND_c_2122_n 0.028083f $X=11.395 $Y=1.095 $X2=0
+ $Y2=0
cc_1000 N_A_1958_48#_c_1426_n N_VGND_c_2122_n 0.027728f $X=11.56 $Y=0.58 $X2=0
+ $Y2=0
cc_1001 N_A_1958_48#_c_1423_n N_VGND_c_2128_n 0.00461464f $X=9.865 $Y=0.865
+ $X2=0 $Y2=0
cc_1002 N_A_1958_48#_c_1426_n N_VGND_c_2130_n 0.0165719f $X=11.56 $Y=0.58 $X2=0
+ $Y2=0
cc_1003 N_A_1958_48#_c_1423_n N_VGND_c_2135_n 0.00914027f $X=9.865 $Y=0.865
+ $X2=0 $Y2=0
cc_1004 N_A_1958_48#_c_1426_n N_VGND_c_2135_n 0.0136604f $X=11.56 $Y=0.58 $X2=0
+ $Y2=0
cc_1005 N_A_1958_48#_c_1431_n N_VGND_c_2135_n 0.0124312f $X=10.385 $Y=1.087
+ $X2=0 $Y2=0
cc_1006 N_A_1764_74#_M1010_g N_A_2395_94#_c_1674_n 0.0179677f $X=12.75 $Y=0.79
+ $X2=0 $Y2=0
cc_1007 N_A_1764_74#_M1010_g N_A_2395_94#_c_1675_n 0.0240619f $X=12.75 $Y=0.79
+ $X2=0 $Y2=0
cc_1008 N_A_1764_74#_c_1533_n N_A_2395_94#_c_1675_n 0.0173812f $X=12.92 $Y=1.94
+ $X2=0 $Y2=0
cc_1009 N_A_1764_74#_c_1537_n N_A_2395_94#_c_1675_n 0.0058249f $X=12.92 $Y=1.865
+ $X2=0 $Y2=0
cc_1010 N_A_1764_74#_M1010_g N_A_2395_94#_c_1676_n 0.00704048f $X=12.75 $Y=0.79
+ $X2=0 $Y2=0
cc_1011 N_A_1764_74#_c_1530_n N_A_2395_94#_c_1682_n 0.00503702f $X=11.93
+ $Y=2.465 $X2=0 $Y2=0
cc_1012 N_A_1764_74#_c_1533_n N_A_2395_94#_c_1682_n 0.0128442f $X=12.92 $Y=1.94
+ $X2=0 $Y2=0
cc_1013 N_A_1764_74#_c_1535_n N_A_2395_94#_c_1682_n 0.00300593f $X=11.93 $Y=2.29
+ $X2=0 $Y2=0
cc_1014 N_A_1764_74#_c_1537_n N_A_2395_94#_c_1682_n 0.0020013f $X=12.92 $Y=1.865
+ $X2=0 $Y2=0
cc_1015 N_A_1764_74#_M1010_g N_A_2395_94#_c_1677_n 0.0157388f $X=12.75 $Y=0.79
+ $X2=0 $Y2=0
cc_1016 N_A_1764_74#_c_1537_n N_A_2395_94#_c_1677_n 0.00705322f $X=12.92
+ $Y=1.865 $X2=0 $Y2=0
cc_1017 N_A_1764_74#_M1038_g N_A_2395_94#_c_1678_n 7.60313e-19 $X=11.345 $Y=0.58
+ $X2=0 $Y2=0
cc_1018 N_A_1764_74#_M1010_g N_A_2395_94#_c_1689_n 0.00791034f $X=12.75 $Y=0.79
+ $X2=0 $Y2=0
cc_1019 N_A_1764_74#_M1010_g N_A_2395_94#_c_1679_n 0.0064711f $X=12.75 $Y=0.79
+ $X2=0 $Y2=0
cc_1020 N_A_1764_74#_c_1531_n N_A_2395_94#_c_1680_n 0.0109169f $X=12.675
+ $Y=1.865 $X2=0 $Y2=0
cc_1021 N_A_1764_74#_M1010_g N_A_2395_94#_c_1680_n 0.00895062f $X=12.75 $Y=0.79
+ $X2=0 $Y2=0
cc_1022 N_A_1764_74#_c_1533_n N_A_2395_94#_c_1680_n 0.00189951f $X=12.92 $Y=1.94
+ $X2=0 $Y2=0
cc_1023 N_A_1764_74#_c_1536_n N_A_2395_94#_c_1680_n 0.00300593f $X=11.945
+ $Y=1.92 $X2=0 $Y2=0
cc_1024 N_A_1764_74#_c_1537_n N_A_2395_94#_c_1680_n 0.00383457f $X=12.92
+ $Y=1.865 $X2=0 $Y2=0
cc_1025 N_A_1764_74#_c_1541_n N_VPWR_c_1741_n 0.0138919f $X=11 $Y=2.305 $X2=0
+ $Y2=0
cc_1026 N_A_1764_74#_c_1543_n N_VPWR_c_1741_n 0.0276292f $X=11.165 $Y=2.75 $X2=0
+ $Y2=0
cc_1027 N_A_1764_74#_c_1530_n N_VPWR_c_1742_n 0.00649842f $X=11.93 $Y=2.465
+ $X2=0 $Y2=0
cc_1028 N_A_1764_74#_c_1531_n N_VPWR_c_1742_n 0.00538998f $X=12.675 $Y=1.865
+ $X2=0 $Y2=0
cc_1029 N_A_1764_74#_c_1533_n N_VPWR_c_1742_n 0.00324414f $X=12.92 $Y=1.94 $X2=0
+ $Y2=0
cc_1030 N_A_1764_74#_c_1533_n N_VPWR_c_1743_n 0.00803512f $X=12.92 $Y=1.94 $X2=0
+ $Y2=0
cc_1031 N_A_1764_74#_c_1530_n N_VPWR_c_1750_n 0.00445602f $X=11.93 $Y=2.465
+ $X2=0 $Y2=0
cc_1032 N_A_1764_74#_c_1543_n N_VPWR_c_1750_n 0.0163786f $X=11.165 $Y=2.75 $X2=0
+ $Y2=0
cc_1033 N_A_1764_74#_c_1533_n N_VPWR_c_1754_n 0.00491343f $X=12.92 $Y=1.94 $X2=0
+ $Y2=0
cc_1034 N_A_1764_74#_c_1530_n N_VPWR_c_1734_n 0.00904625f $X=11.93 $Y=2.465
+ $X2=0 $Y2=0
cc_1035 N_A_1764_74#_c_1533_n N_VPWR_c_1734_n 0.00512916f $X=12.92 $Y=1.94 $X2=0
+ $Y2=0
cc_1036 N_A_1764_74#_c_1543_n N_VPWR_c_1734_n 0.0135239f $X=11.165 $Y=2.75 $X2=0
+ $Y2=0
cc_1037 N_A_1764_74#_M1009_d N_A_1610_341#_c_2027_n 0.0054832f $X=9.02 $Y=1.87
+ $X2=0 $Y2=0
cc_1038 N_A_1764_74#_c_1538_n N_A_1610_341#_c_2027_n 0.0217217f $X=9.275
+ $Y=2.015 $X2=0 $Y2=0
cc_1039 N_A_1764_74#_c_1523_n N_A_1610_341#_c_2027_n 0.00386096f $X=10.065
+ $Y=1.705 $X2=0 $Y2=0
cc_1040 N_A_1764_74#_c_1542_n N_A_1610_341#_c_2027_n 0.00374779f $X=10.235
+ $Y=2.305 $X2=0 $Y2=0
cc_1041 N_A_1764_74#_c_1538_n N_A_1610_341#_c_2029_n 0.0148589f $X=9.275
+ $Y=2.015 $X2=0 $Y2=0
cc_1042 N_A_1764_74#_c_1523_n N_A_1610_341#_c_2029_n 0.0224145f $X=10.065
+ $Y=1.705 $X2=0 $Y2=0
cc_1043 N_A_1764_74#_c_1540_n N_A_1610_341#_c_2029_n 0.0205759f $X=10.15 $Y=2.22
+ $X2=0 $Y2=0
cc_1044 N_A_1764_74#_c_1542_n N_A_1610_341#_c_2029_n 0.0114578f $X=10.235
+ $Y=2.305 $X2=0 $Y2=0
cc_1045 N_A_1764_74#_c_1542_n N_A_1721_374#_c_2070_n 0.00135116f $X=10.235
+ $Y=2.305 $X2=0 $Y2=0
cc_1046 N_A_1764_74#_c_1541_n N_A_1721_374#_c_2071_n 0.0127126f $X=11 $Y=2.305
+ $X2=0 $Y2=0
cc_1047 N_A_1764_74#_c_1542_n N_A_1721_374#_c_2071_n 0.0121231f $X=10.235
+ $Y=2.305 $X2=0 $Y2=0
cc_1048 N_A_1764_74#_c_1526_n N_VGND_c_2121_n 0.0206027f $X=9.07 $Y=0.515 $X2=0
+ $Y2=0
cc_1049 N_A_1764_74#_M1038_g N_VGND_c_2122_n 0.00713799f $X=11.345 $Y=0.58 $X2=0
+ $Y2=0
cc_1050 N_A_1764_74#_M1010_g N_VGND_c_2123_n 0.00726265f $X=12.75 $Y=0.79 $X2=0
+ $Y2=0
cc_1051 N_A_1764_74#_c_1526_n N_VGND_c_2128_n 0.0250915f $X=9.07 $Y=0.515 $X2=0
+ $Y2=0
cc_1052 N_A_1764_74#_M1038_g N_VGND_c_2130_n 0.00434272f $X=11.345 $Y=0.58 $X2=0
+ $Y2=0
cc_1053 N_A_1764_74#_M1010_g N_VGND_c_2130_n 0.00486038f $X=12.75 $Y=0.79 $X2=0
+ $Y2=0
cc_1054 N_A_1764_74#_M1038_g N_VGND_c_2135_n 0.00827521f $X=11.345 $Y=0.58 $X2=0
+ $Y2=0
cc_1055 N_A_1764_74#_M1010_g N_VGND_c_2135_n 0.00514438f $X=12.75 $Y=0.79 $X2=0
+ $Y2=0
cc_1056 N_A_1764_74#_c_1526_n N_VGND_c_2135_n 0.0207918f $X=9.07 $Y=0.515 $X2=0
+ $Y2=0
cc_1057 N_A_2395_94#_c_1682_n N_VPWR_c_1742_n 0.022154f $X=12.695 $Y=2.16 $X2=0
+ $Y2=0
cc_1058 N_A_2395_94#_c_1675_n N_VPWR_c_1743_n 0.0257364f $X=13.425 $Y=1.765
+ $X2=0 $Y2=0
cc_1059 N_A_2395_94#_c_1682_n N_VPWR_c_1743_n 0.0345631f $X=12.695 $Y=2.16 $X2=0
+ $Y2=0
cc_1060 N_A_2395_94#_c_1677_n N_VPWR_c_1743_n 0.0118229f $X=13.23 $Y=1.385 $X2=0
+ $Y2=0
cc_1061 N_A_2395_94#_c_1682_n N_VPWR_c_1754_n 0.0102252f $X=12.695 $Y=2.16 $X2=0
+ $Y2=0
cc_1062 N_A_2395_94#_c_1675_n N_VPWR_c_1755_n 0.00429299f $X=13.425 $Y=1.765
+ $X2=0 $Y2=0
cc_1063 N_A_2395_94#_c_1675_n N_VPWR_c_1734_n 0.00851182f $X=13.425 $Y=1.765
+ $X2=0 $Y2=0
cc_1064 N_A_2395_94#_c_1682_n N_VPWR_c_1734_n 0.0113067f $X=12.695 $Y=2.16 $X2=0
+ $Y2=0
cc_1065 N_A_2395_94#_c_1674_n Q 0.0029127f $X=13.33 $Y=1.22 $X2=0 $Y2=0
cc_1066 N_A_2395_94#_c_1675_n Q 0.00391287f $X=13.425 $Y=1.765 $X2=0 $Y2=0
cc_1067 N_A_2395_94#_c_1677_n Q 0.00112015f $X=13.23 $Y=1.385 $X2=0 $Y2=0
cc_1068 N_A_2395_94#_c_1674_n Q 0.00561171f $X=13.33 $Y=1.22 $X2=0 $Y2=0
cc_1069 N_A_2395_94#_c_1675_n Q 0.0292597f $X=13.425 $Y=1.765 $X2=0 $Y2=0
cc_1070 N_A_2395_94#_c_1677_n Q 0.0269563f $X=13.23 $Y=1.385 $X2=0 $Y2=0
cc_1071 N_A_2395_94#_c_1674_n N_Q_c_2102_n 0.00562579f $X=13.33 $Y=1.22 $X2=0
+ $Y2=0
cc_1072 N_A_2395_94#_c_1674_n N_VGND_c_2123_n 0.00890609f $X=13.33 $Y=1.22 $X2=0
+ $Y2=0
cc_1073 N_A_2395_94#_c_1675_n N_VGND_c_2123_n 0.00332106f $X=13.425 $Y=1.765
+ $X2=0 $Y2=0
cc_1074 N_A_2395_94#_c_1677_n N_VGND_c_2123_n 0.0273042f $X=13.23 $Y=1.385 $X2=0
+ $Y2=0
cc_1075 N_A_2395_94#_c_1678_n N_VGND_c_2130_n 0.0165214f $X=12.37 $Y=0.772 $X2=0
+ $Y2=0
cc_1076 N_A_2395_94#_c_1674_n N_VGND_c_2134_n 0.00434272f $X=13.33 $Y=1.22 $X2=0
+ $Y2=0
cc_1077 N_A_2395_94#_c_1674_n N_VGND_c_2135_n 0.00829f $X=13.33 $Y=1.22 $X2=0
+ $Y2=0
cc_1078 N_A_2395_94#_c_1678_n N_VGND_c_2135_n 0.0235982f $X=12.37 $Y=0.772 $X2=0
+ $Y2=0
cc_1079 N_VPWR_c_1735_n N_A_289_464#_c_1907_n 0.00764771f $X=0.725 $Y=2.78 $X2=0
+ $Y2=0
cc_1080 N_VPWR_c_1753_n N_A_289_464#_c_1907_n 0.0221221f $X=2.565 $Y=3.33 $X2=0
+ $Y2=0
cc_1081 N_VPWR_c_1734_n N_A_289_464#_c_1907_n 0.0259323f $X=13.68 $Y=3.33 $X2=0
+ $Y2=0
cc_1082 N_VPWR_M1028_d N_A_289_464#_c_1903_n 0.00992545f $X=2.495 $Y=2.32 $X2=0
+ $Y2=0
cc_1083 N_VPWR_c_1736_n N_A_289_464#_c_1903_n 0.0253286f $X=2.73 $Y=2.995 $X2=0
+ $Y2=0
cc_1084 N_VPWR_c_1737_n N_A_289_464#_c_1903_n 0.00567825f $X=3.575 $Y=3.33 $X2=0
+ $Y2=0
cc_1085 N_VPWR_c_1753_n N_A_289_464#_c_1903_n 0.00236889f $X=2.565 $Y=3.33 $X2=0
+ $Y2=0
cc_1086 N_VPWR_c_1734_n N_A_289_464#_c_1903_n 0.0153638f $X=13.68 $Y=3.33 $X2=0
+ $Y2=0
cc_1087 N_VPWR_c_1736_n N_A_289_464#_c_1928_n 0.0056644f $X=2.73 $Y=2.995 $X2=0
+ $Y2=0
cc_1088 N_VPWR_c_1753_n N_A_289_464#_c_1928_n 0.00470407f $X=2.565 $Y=3.33 $X2=0
+ $Y2=0
cc_1089 N_VPWR_c_1734_n N_A_289_464#_c_1928_n 0.00574301f $X=13.68 $Y=3.33 $X2=0
+ $Y2=0
cc_1090 N_VPWR_c_1737_n N_A_289_464#_c_1981_n 0.00272847f $X=3.575 $Y=3.33 $X2=0
+ $Y2=0
cc_1091 N_VPWR_c_1734_n N_A_289_464#_c_1981_n 0.00485809f $X=13.68 $Y=3.33 $X2=0
+ $Y2=0
cc_1092 N_VPWR_M1032_d N_A_289_464#_c_1905_n 0.00395925f $X=3.59 $Y=1.84 $X2=0
+ $Y2=0
cc_1093 N_VPWR_c_1738_n N_A_289_464#_c_1905_n 0.0172656f $X=3.74 $Y=2.78 $X2=0
+ $Y2=0
cc_1094 N_VPWR_c_1740_n N_A_1610_341#_c_2026_n 0.00259305f $X=7.75 $Y=2.515
+ $X2=0 $Y2=0
cc_1095 N_VPWR_c_1734_n N_A_1610_341#_c_2027_n 0.00775297f $X=13.68 $Y=3.33
+ $X2=0 $Y2=0
cc_1096 N_VPWR_c_1740_n N_A_1610_341#_c_2028_n 0.0257014f $X=7.75 $Y=2.515 $X2=0
+ $Y2=0
cc_1097 N_VPWR_c_1748_n N_A_1610_341#_c_2028_n 0.00538584f $X=10.63 $Y=3.33
+ $X2=0 $Y2=0
cc_1098 N_VPWR_c_1734_n N_A_1610_341#_c_2028_n 0.00676831f $X=13.68 $Y=3.33
+ $X2=0 $Y2=0
cc_1099 N_VPWR_c_1741_n N_A_1721_374#_c_2070_n 0.0119328f $X=10.715 $Y=2.77
+ $X2=0 $Y2=0
cc_1100 N_VPWR_c_1748_n N_A_1721_374#_c_2070_n 0.0988914f $X=10.63 $Y=3.33 $X2=0
+ $Y2=0
cc_1101 N_VPWR_c_1734_n N_A_1721_374#_c_2070_n 0.0543782f $X=13.68 $Y=3.33 $X2=0
+ $Y2=0
cc_1102 N_VPWR_c_1741_n N_A_1721_374#_c_2071_n 0.0224393f $X=10.715 $Y=2.77
+ $X2=0 $Y2=0
cc_1103 N_VPWR_c_1740_n N_A_1721_374#_c_2072_n 0.0105193f $X=7.75 $Y=2.515 $X2=0
+ $Y2=0
cc_1104 N_VPWR_c_1748_n N_A_1721_374#_c_2072_n 0.0214714f $X=10.63 $Y=3.33 $X2=0
+ $Y2=0
cc_1105 N_VPWR_c_1734_n N_A_1721_374#_c_2072_n 0.0110721f $X=13.68 $Y=3.33 $X2=0
+ $Y2=0
cc_1106 N_VPWR_c_1743_n Q 0.0648352f $X=13.195 $Y=2.16 $X2=0 $Y2=0
cc_1107 N_VPWR_c_1755_n Q 0.011066f $X=13.68 $Y=3.33 $X2=0 $Y2=0
cc_1108 N_VPWR_c_1734_n Q 0.00915947f $X=13.68 $Y=3.33 $X2=0 $Y2=0
cc_1109 N_A_289_464#_c_1907_n A_415_464# 0.00499203f $X=2.215 $Y=2.785 $X2=-0.19
+ $Y2=-0.245
cc_1110 N_A_289_464#_c_1899_n A_415_464# 0.00139793f $X=2.3 $Y=2.49 $X2=-0.19
+ $Y2=-0.245
cc_1111 N_A_289_464#_c_1928_n A_415_464# 0.00350847f $X=2.3 $Y=2.575 $X2=-0.19
+ $Y2=-0.245
cc_1112 N_A_289_464#_c_1896_n N_VGND_c_2117_n 0.00656395f $X=1.72 $Y=0.58 $X2=0
+ $Y2=0
cc_1113 N_A_289_464#_c_1896_n N_VGND_c_2118_n 0.0126723f $X=1.72 $Y=0.58 $X2=0
+ $Y2=0
cc_1114 N_A_289_464#_c_1897_n N_VGND_c_2118_n 7.61858e-19 $X=2.215 $Y=1.005
+ $X2=0 $Y2=0
cc_1115 N_A_289_464#_c_1896_n N_VGND_c_2124_n 0.0144922f $X=1.72 $Y=0.58 $X2=0
+ $Y2=0
cc_1116 N_A_289_464#_c_1896_n N_VGND_c_2135_n 0.0118826f $X=1.72 $Y=0.58 $X2=0
+ $Y2=0
cc_1117 N_A_1610_341#_c_2027_n N_A_1721_374#_M1009_s 0.00507898f $X=9.565
+ $Y=2.435 $X2=-0.19 $Y2=1.66
cc_1118 N_A_1610_341#_c_2027_n N_A_1721_374#_c_2070_n 0.0436761f $X=9.565
+ $Y=2.435 $X2=0 $Y2=0
cc_1119 N_A_1610_341#_c_2027_n N_A_1721_374#_c_2071_n 0.0128284f $X=9.565
+ $Y=2.435 $X2=0 $Y2=0
cc_1120 N_A_1610_341#_c_2027_n N_A_1721_374#_c_2072_n 0.0266315f $X=9.565
+ $Y=2.435 $X2=0 $Y2=0
cc_1121 N_A_1610_341#_c_2028_n N_A_1721_374#_c_2072_n 0.00239231f $X=8.365
+ $Y=2.435 $X2=0 $Y2=0
cc_1122 N_Q_c_2102_n N_VGND_c_2123_n 0.0281509f $X=13.545 $Y=0.515 $X2=0 $Y2=0
cc_1123 N_Q_c_2102_n N_VGND_c_2134_n 0.0192663f $X=13.545 $Y=0.515 $X2=0 $Y2=0
cc_1124 N_Q_c_2102_n N_VGND_c_2135_n 0.0158831f $X=13.545 $Y=0.515 $X2=0 $Y2=0
