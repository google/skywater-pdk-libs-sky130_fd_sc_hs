* NGSPICE file created from sky130_fd_sc_hs__sdfbbn_1.ext - technology: sky130A

.subckt sky130_fd_sc_hs__sdfbbn_1 CLK_N D RESET_B SCD SCE SET_B VGND VNB VPB VPWR
+ Q Q_N
M1000 a_305_119# D a_197_119# VNB nlowvt w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=3.129e+11p ps=3.17e+06u
M1001 a_197_119# a_867_82# a_1159_497# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.176e+11p ps=1.4e+06u
M1002 VGND RESET_B a_1579_258# VNB nlowvt w=420000u l=150000u
+  ad=2.11888e+12p pd=1.742e+07u as=1.197e+11p ps=1.41e+06u
M1003 a_977_243# a_1159_497# a_1434_78# VNB nlowvt w=550000u l=150000u
+  ad=2.09e+11p pd=1.86e+06u as=5.1045e+11p ps=4.25e+06u
M1004 a_119_119# SCD VGND VNB nlowvt w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=0p ps=0u
M1005 Q_N a_2133_410# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1006 Q_N a_2133_410# VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=3.304e+11p pd=2.83e+06u as=3.0812e+12p ps=2.468e+07u
M1007 a_2392_74# SET_B VGND VNB nlowvt w=740000u l=150000u
+  ad=4.947e+11p pd=4.37e+06u as=0p ps=0u
M1008 a_2133_410# a_1954_119# a_2509_392# VPB pshort w=1e+06u l=150000u
+  ad=5.9e+11p pd=5.18e+06u as=2.7e+11p ps=2.54e+06u
M1009 VPWR RESET_B a_1579_258# VPB pshort w=640000u l=150000u
+  ad=0p pd=0u as=3.625e+11p ps=3.71e+06u
M1010 VGND a_2133_410# a_2164_119# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.638e+11p ps=1.62e+06u
M1011 a_1081_497# a_977_243# VPWR VPB pshort w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=0p ps=0u
M1012 a_1903_424# a_977_243# VPWR VPB pshort w=840000u l=150000u
+  ad=2.016e+11p pd=2.16e+06u as=0p ps=0u
M1013 a_353_93# SCE VPWR VPB pshort w=640000u l=150000u
+  ad=1.888e+11p pd=1.87e+06u as=0p ps=0u
M1014 a_212_464# SCE VPWR VPB pshort w=640000u l=150000u
+  ad=1.728e+11p pd=1.82e+06u as=0p ps=0u
M1015 VGND CLK_N a_662_82# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1016 a_867_82# a_662_82# VGND VNB nlowvt w=740000u l=150000u
+  ad=3.219e+11p pd=2.35e+06u as=0p ps=0u
M1017 a_1159_497# a_662_82# a_1151_119# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=8.82e+10p ps=1.26e+06u
M1018 a_353_93# SCE VGND VNB nlowvt w=420000u l=150000u
+  ad=1.197e+11p pd=1.41e+06u as=0p ps=0u
M1019 VGND a_2133_410# a_3078_384# VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=1.5675e+11p ps=1.67e+06u
M1020 VPWR SCD a_27_464# VPB pshort w=640000u l=150000u
+  ad=0p pd=0u as=3.744e+11p ps=3.73e+06u
M1021 a_1151_119# a_977_243# VGND VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 VPWR a_1579_258# a_1528_424# VPB pshort w=840000u l=150000u
+  ad=0p pd=0u as=2.268e+11p ps=2.22e+06u
M1023 a_197_119# D a_212_464# VPB pshort w=640000u l=150000u
+  ad=4.128e+11p pd=3.85e+06u as=0p ps=0u
M1024 VPWR a_2133_410# a_2088_508# VPB pshort w=420000u l=150000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1025 VGND SET_B a_1434_78# VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 a_977_243# SET_B VPWR VPB pshort w=840000u l=150000u
+  ad=6.342e+11p pd=4.87e+06u as=0p ps=0u
M1027 a_1954_119# a_662_82# a_1876_119# VNB nlowvt w=550000u l=150000u
+  ad=4.807e+11p pd=2.9e+06u as=1.32e+11p ps=1.58e+06u
M1028 VPWR a_2133_410# a_3078_384# VPB pshort w=840000u l=150000u
+  ad=0p pd=0u as=2.478e+11p ps=2.27e+06u
M1029 a_27_464# a_353_93# a_197_119# VPB pshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1030 a_1159_497# a_867_82# a_1081_497# VPB pshort w=420000u l=150000u
+  ad=2.266e+11p pd=2.05e+06u as=0p ps=0u
M1031 a_197_119# a_662_82# a_1159_497# VPB pshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1032 a_2392_74# a_1954_119# a_2133_410# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.812e+11p ps=2.24e+06u
M1033 a_197_119# SCE a_119_119# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1034 VGND a_353_93# a_305_119# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1035 a_2509_392# a_1579_258# VPWR VPB pshort w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1036 Q a_3078_384# VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=3.304e+11p pd=2.83e+06u as=0p ps=0u
M1037 Q a_3078_384# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1038 a_2133_410# a_1579_258# a_2392_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1039 a_2164_119# a_867_82# a_1954_119# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1040 VPWR CLK_N a_662_82# VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=3.304e+11p ps=2.83e+06u
M1041 a_2088_508# a_662_82# a_1954_119# VPB pshort w=420000u l=150000u
+  ad=0p pd=0u as=2.856e+11p ps=2.45e+06u
M1042 VPWR SET_B a_2133_410# VPB pshort w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1043 a_1876_119# a_977_243# VGND VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1044 a_1954_119# a_867_82# a_1903_424# VPB pshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1045 a_867_82# a_662_82# VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=3.304e+11p pd=2.83e+06u as=0p ps=0u
M1046 a_1528_424# a_1159_497# a_977_243# VPB pshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1047 a_1434_78# a_1579_258# a_977_243# VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

