* File: sky130_fd_sc_hs__nor3b_4.pxi.spice
* Created: Thu Aug 27 20:54:32 2020
* 
x_PM_SKY130_FD_SC_HS__NOR3B_4%B N_B_M1003_g N_B_c_118_n N_B_M1010_g N_B_M1008_g
+ N_B_c_119_n N_B_M1012_g N_B_c_120_n N_B_M1014_g N_B_M1024_g N_B_c_121_n
+ N_B_M1016_g N_B_M1026_g B B B B N_B_c_117_n PM_SKY130_FD_SC_HS__NOR3B_4%B
x_PM_SKY130_FD_SC_HS__NOR3B_4%A_468_264# N_A_468_264#_M1006_d
+ N_A_468_264#_M1004_d N_A_468_264#_c_203_n N_A_468_264#_M1018_g
+ N_A_468_264#_M1000_g N_A_468_264#_c_204_n N_A_468_264#_M1020_g
+ N_A_468_264#_M1001_g N_A_468_264#_c_205_n N_A_468_264#_M1023_g
+ N_A_468_264#_M1009_g N_A_468_264#_c_206_n N_A_468_264#_M1025_g
+ N_A_468_264#_M1013_g N_A_468_264#_c_198_n N_A_468_264#_c_208_n
+ N_A_468_264#_c_209_n N_A_468_264#_c_210_n N_A_468_264#_c_199_n
+ N_A_468_264#_c_200_n N_A_468_264#_c_233_p N_A_468_264#_c_201_n
+ N_A_468_264#_c_202_n PM_SKY130_FD_SC_HS__NOR3B_4%A_468_264#
x_PM_SKY130_FD_SC_HS__NOR3B_4%A N_A_c_343_n N_A_M1002_g N_A_c_350_n N_A_M1007_g
+ N_A_c_344_n N_A_M1011_g N_A_c_351_n N_A_M1017_g N_A_c_345_n N_A_M1015_g
+ N_A_c_352_n N_A_M1019_g N_A_c_346_n N_A_M1022_g N_A_c_353_n N_A_M1021_g A
+ N_A_c_348_n N_A_c_349_n PM_SKY130_FD_SC_HS__NOR3B_4%A
x_PM_SKY130_FD_SC_HS__NOR3B_4%C_N N_C_N_c_432_n N_C_N_M1006_g N_C_N_c_435_n
+ N_C_N_M1004_g N_C_N_c_436_n N_C_N_M1005_g C_N N_C_N_c_434_n
+ PM_SKY130_FD_SC_HS__NOR3B_4%C_N
x_PM_SKY130_FD_SC_HS__NOR3B_4%A_27_368# N_A_27_368#_M1010_d N_A_27_368#_M1012_d
+ N_A_27_368#_M1016_d N_A_27_368#_M1020_s N_A_27_368#_M1025_s
+ N_A_27_368#_c_470_n N_A_27_368#_c_471_n N_A_27_368#_c_472_n
+ N_A_27_368#_c_500_p N_A_27_368#_c_473_n N_A_27_368#_c_485_n
+ N_A_27_368#_c_474_n N_A_27_368#_c_475_n N_A_27_368#_c_489_n
+ N_A_27_368#_c_491_n N_A_27_368#_c_476_n PM_SKY130_FD_SC_HS__NOR3B_4%A_27_368#
x_PM_SKY130_FD_SC_HS__NOR3B_4%A_126_368# N_A_126_368#_M1010_s
+ N_A_126_368#_M1014_s N_A_126_368#_M1007_d N_A_126_368#_M1019_d
+ N_A_126_368#_c_539_n N_A_126_368#_c_536_n N_A_126_368#_c_537_n
+ N_A_126_368#_c_561_n N_A_126_368#_c_562_n N_A_126_368#_c_538_n
+ N_A_126_368#_c_544_n N_A_126_368#_c_549_n N_A_126_368#_c_563_n
+ PM_SKY130_FD_SC_HS__NOR3B_4%A_126_368#
x_PM_SKY130_FD_SC_HS__NOR3B_4%Y N_Y_M1003_s N_Y_M1024_s N_Y_M1000_s N_Y_M1009_s
+ N_Y_M1002_d N_Y_M1015_d N_Y_M1018_d N_Y_M1023_d N_Y_c_604_n N_Y_c_605_n
+ N_Y_c_606_n N_Y_c_607_n N_Y_c_630_n N_Y_c_618_n N_Y_c_608_n N_Y_c_609_n
+ N_Y_c_610_n N_Y_c_663_n N_Y_c_611_n N_Y_c_685_n N_Y_c_612_n N_Y_c_613_n
+ N_Y_c_614_n N_Y_c_615_n N_Y_c_616_n N_Y_c_693_n Y
+ PM_SKY130_FD_SC_HS__NOR3B_4%Y
x_PM_SKY130_FD_SC_HS__NOR3B_4%VPWR N_VPWR_M1007_s N_VPWR_M1017_s N_VPWR_M1021_s
+ N_VPWR_M1005_s N_VPWR_c_743_n N_VPWR_c_744_n N_VPWR_c_745_n N_VPWR_c_746_n
+ N_VPWR_c_747_n VPWR N_VPWR_c_748_n N_VPWR_c_749_n N_VPWR_c_750_n
+ N_VPWR_c_751_n N_VPWR_c_752_n N_VPWR_c_753_n N_VPWR_c_754_n N_VPWR_c_742_n
+ PM_SKY130_FD_SC_HS__NOR3B_4%VPWR
x_PM_SKY130_FD_SC_HS__NOR3B_4%VGND N_VGND_M1003_d N_VGND_M1008_d N_VGND_M1026_d
+ N_VGND_M1001_d N_VGND_M1013_d N_VGND_M1011_s N_VGND_M1022_s N_VGND_c_836_n
+ N_VGND_c_837_n N_VGND_c_838_n N_VGND_c_839_n N_VGND_c_840_n N_VGND_c_841_n
+ N_VGND_c_842_n N_VGND_c_843_n N_VGND_c_844_n N_VGND_c_845_n N_VGND_c_846_n
+ N_VGND_c_847_n VGND N_VGND_c_848_n N_VGND_c_849_n N_VGND_c_850_n
+ N_VGND_c_851_n N_VGND_c_852_n N_VGND_c_853_n N_VGND_c_854_n N_VGND_c_855_n
+ N_VGND_c_856_n N_VGND_c_857_n PM_SKY130_FD_SC_HS__NOR3B_4%VGND
cc_1 VNB N_B_M1003_g 0.030989f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=0.74
cc_2 VNB N_B_M1008_g 0.0252957f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=0.74
cc_3 VNB N_B_M1024_g 0.0248983f $X=-0.19 $Y=-0.245 $X2=1.565 $Y2=0.74
cc_4 VNB N_B_M1026_g 0.023399f $X=-0.19 $Y=-0.245 $X2=1.995 $Y2=0.74
cc_5 VNB B 0.018482f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=1.58
cc_6 VNB N_B_c_117_n 0.0768894f $X=-0.19 $Y=-0.245 $X2=1.98 $Y2=1.557
cc_7 VNB N_A_468_264#_M1000_g 0.0222712f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=1.765
cc_8 VNB N_A_468_264#_M1001_g 0.0220929f $X=-0.19 $Y=-0.245 $X2=1.565 $Y2=0.74
cc_9 VNB N_A_468_264#_M1009_g 0.0226931f $X=-0.19 $Y=-0.245 $X2=1.995 $Y2=0.74
cc_10 VNB N_A_468_264#_M1013_g 0.0241345f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_468_264#_c_198_n 0.00717215f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_468_264#_c_199_n 0.0289376f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_468_264#_c_200_n 0.031855f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.565
cc_14 VNB N_A_468_264#_c_201_n 0.00697138f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_468_264#_c_202_n 0.104613f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_c_343_n 0.0185806f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=1.35
cc_17 VNB N_A_c_344_n 0.0191883f $X=-0.19 $Y=-0.245 $X2=0.555 $Y2=2.4
cc_18 VNB N_A_c_345_n 0.0198403f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=2.4
cc_19 VNB N_A_c_346_n 0.0179355f $X=-0.19 $Y=-0.245 $X2=1.565 $Y2=0.74
cc_20 VNB A 0.00598605f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_c_348_n 0.138284f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=1.557
cc_22 VNB N_A_c_349_n 0.00358389f $X=-0.19 $Y=-0.245 $X2=1.65 $Y2=1.557
cc_23 VNB N_C_N_c_432_n 0.0236108f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=1.35
cc_24 VNB C_N 0.00374395f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=0.74
cc_25 VNB N_C_N_c_434_n 0.0735994f $X=-0.19 $Y=-0.245 $X2=1.455 $Y2=1.765
cc_26 VNB N_Y_c_604_n 0.00280814f $X=-0.19 $Y=-0.245 $X2=1.995 $Y2=0.74
cc_27 VNB N_Y_c_605_n 0.00273768f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_28 VNB N_Y_c_606_n 0.00239855f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_Y_c_607_n 0.00224624f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_Y_c_608_n 0.00178908f $X=-0.19 $Y=-0.245 $X2=1.565 $Y2=1.557
cc_31 VNB N_Y_c_609_n 0.00317099f $X=-0.19 $Y=-0.245 $X2=1.65 $Y2=1.515
cc_32 VNB N_Y_c_610_n 0.00240191f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.565
cc_33 VNB N_Y_c_611_n 0.00240319f $X=-0.19 $Y=-0.245 $X2=1.2 $Y2=1.565
cc_34 VNB N_Y_c_612_n 0.0028001f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_Y_c_613_n 0.00323083f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_Y_c_614_n 0.00554939f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_Y_c_615_n 0.00127131f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_Y_c_616_n 0.00230427f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB Y 0.00464838f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_VPWR_c_742_n 0.322901f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_836_n 0.0122168f $X=-0.19 $Y=-0.245 $X2=1.98 $Y2=1.765
cc_42 VNB N_VGND_c_837_n 0.0454867f $X=-0.19 $Y=-0.245 $X2=1.98 $Y2=2.4
cc_43 VNB N_VGND_c_838_n 0.00830803f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_839_n 0.0186948f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_45 VNB N_VGND_c_840_n 0.00498656f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_VGND_c_841_n 0.00498656f $X=-0.19 $Y=-0.245 $X2=0.555 $Y2=1.557
cc_47 VNB N_VGND_c_842_n 0.00830803f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=1.557
cc_48 VNB N_VGND_c_843_n 0.0186948f $X=-0.19 $Y=-0.245 $X2=1.455 $Y2=1.557
cc_49 VNB N_VGND_c_844_n 0.00967485f $X=-0.19 $Y=-0.245 $X2=1.65 $Y2=1.515
cc_50 VNB N_VGND_c_845_n 0.00586131f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_VGND_c_846_n 0.0185368f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.565
cc_52 VNB N_VGND_c_847_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_VGND_c_848_n 0.018682f $X=-0.19 $Y=-0.245 $X2=1.65 $Y2=1.565
cc_54 VNB N_VGND_c_849_n 0.0151736f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_VGND_c_850_n 0.0186948f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_VGND_c_851_n 0.0342743f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_VGND_c_852_n 0.412273f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_VGND_c_853_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_VGND_c_854_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_VGND_c_855_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_VGND_c_856_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_VGND_c_857_n 0.00884799f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VPB N_B_c_118_n 0.0186669f $X=-0.19 $Y=1.66 $X2=0.555 $Y2=1.765
cc_64 VPB N_B_c_119_n 0.014664f $X=-0.19 $Y=1.66 $X2=1.005 $Y2=1.765
cc_65 VPB N_B_c_120_n 0.0152196f $X=-0.19 $Y=1.66 $X2=1.455 $Y2=1.765
cc_66 VPB N_B_c_121_n 0.0150144f $X=-0.19 $Y=1.66 $X2=1.98 $Y2=1.765
cc_67 VPB B 0.0188074f $X=-0.19 $Y=1.66 $X2=1.595 $Y2=1.58
cc_68 VPB N_B_c_117_n 0.0504594f $X=-0.19 $Y=1.66 $X2=1.98 $Y2=1.557
cc_69 VPB N_A_468_264#_c_203_n 0.0151318f $X=-0.19 $Y=1.66 $X2=0.555 $Y2=2.4
cc_70 VPB N_A_468_264#_c_204_n 0.0155385f $X=-0.19 $Y=1.66 $X2=1.005 $Y2=2.4
cc_71 VPB N_A_468_264#_c_205_n 0.0155643f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_72 VPB N_A_468_264#_c_206_n 0.0173429f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_73 VPB N_A_468_264#_c_198_n 0.00416751f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_74 VPB N_A_468_264#_c_208_n 0.0202079f $X=-0.19 $Y=1.66 $X2=1.005 $Y2=1.557
cc_75 VPB N_A_468_264#_c_209_n 0.00350815f $X=-0.19 $Y=1.66 $X2=1.98 $Y2=1.557
cc_76 VPB N_A_468_264#_c_210_n 0.0121029f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=1.565
cc_77 VPB N_A_468_264#_c_200_n 0.00283905f $X=-0.19 $Y=1.66 $X2=0.63 $Y2=1.565
cc_78 VPB N_A_468_264#_c_202_n 0.0260456f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_79 VPB N_A_c_350_n 0.0173759f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_80 VPB N_A_c_351_n 0.0144397f $X=-0.19 $Y=1.66 $X2=0.995 $Y2=0.74
cc_81 VPB N_A_c_352_n 0.0144414f $X=-0.19 $Y=1.66 $X2=1.455 $Y2=2.4
cc_82 VPB N_A_c_353_n 0.0157487f $X=-0.19 $Y=1.66 $X2=1.98 $Y2=1.765
cc_83 VPB N_A_c_348_n 0.0263331f $X=-0.19 $Y=1.66 $X2=1.005 $Y2=1.557
cc_84 VPB N_C_N_c_435_n 0.0157152f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_85 VPB N_C_N_c_436_n 0.0170788f $X=-0.19 $Y=1.66 $X2=0.555 $Y2=2.4
cc_86 VPB N_C_N_c_434_n 0.0214551f $X=-0.19 $Y=1.66 $X2=1.455 $Y2=1.765
cc_87 VPB N_A_27_368#_c_470_n 0.0366851f $X=-0.19 $Y=1.66 $X2=1.565 $Y2=1.35
cc_88 VPB N_A_27_368#_c_471_n 0.0028338f $X=-0.19 $Y=1.66 $X2=1.98 $Y2=1.765
cc_89 VPB N_A_27_368#_c_472_n 0.0101535f $X=-0.19 $Y=1.66 $X2=1.98 $Y2=2.4
cc_90 VPB N_A_27_368#_c_473_n 0.00318897f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_91 VPB N_A_27_368#_c_474_n 0.00123754f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_92 VPB N_A_27_368#_c_475_n 0.00217207f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_93 VPB N_A_27_368#_c_476_n 0.00328928f $X=-0.19 $Y=1.66 $X2=1.565 $Y2=1.557
cc_94 VPB N_A_126_368#_c_536_n 0.0131354f $X=-0.19 $Y=1.66 $X2=1.455 $Y2=2.4
cc_95 VPB N_A_126_368#_c_537_n 0.0019689f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_96 VPB N_A_126_368#_c_538_n 0.00239564f $X=-0.19 $Y=1.66 $X2=1.995 $Y2=0.74
cc_97 VPB N_Y_c_618_n 0.00674186f $X=-0.19 $Y=1.66 $X2=0.63 $Y2=1.515
cc_98 VPB Y 0.00150537f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_99 VPB N_VPWR_c_743_n 0.0104359f $X=-0.19 $Y=1.66 $X2=1.455 $Y2=1.765
cc_100 VPB N_VPWR_c_744_n 0.0026822f $X=-0.19 $Y=1.66 $X2=1.565 $Y2=0.74
cc_101 VPB N_VPWR_c_745_n 0.0125948f $X=-0.19 $Y=1.66 $X2=1.98 $Y2=2.4
cc_102 VPB N_VPWR_c_746_n 0.0121909f $X=-0.19 $Y=1.66 $X2=1.995 $Y2=0.74
cc_103 VPB N_VPWR_c_747_n 0.0510603f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_104 VPB N_VPWR_c_748_n 0.110141f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_105 VPB N_VPWR_c_749_n 0.0164205f $X=-0.19 $Y=1.66 $X2=0.63 $Y2=1.515
cc_106 VPB N_VPWR_c_750_n 0.017373f $X=-0.19 $Y=1.66 $X2=1.65 $Y2=1.557
cc_107 VPB N_VPWR_c_751_n 0.0195748f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=1.565
cc_108 VPB N_VPWR_c_752_n 0.00614127f $X=-0.19 $Y=1.66 $X2=1.2 $Y2=1.565
cc_109 VPB N_VPWR_c_753_n 0.00601644f $X=-0.19 $Y=1.66 $X2=1.68 $Y2=1.565
cc_110 VPB N_VPWR_c_754_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_111 VPB N_VPWR_c_742_n 0.101959f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_112 N_B_c_121_n N_A_468_264#_c_203_n 0.038933f $X=1.98 $Y=1.765 $X2=0 $Y2=0
cc_113 N_B_M1026_g N_A_468_264#_M1000_g 0.0264048f $X=1.995 $Y=0.74 $X2=0 $Y2=0
cc_114 N_B_M1026_g N_A_468_264#_c_198_n 2.25772e-19 $X=1.995 $Y=0.74 $X2=0 $Y2=0
cc_115 N_B_M1026_g N_A_468_264#_c_202_n 0.0204851f $X=1.995 $Y=0.74 $X2=0 $Y2=0
cc_116 B N_A_27_368#_c_470_n 0.027274f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_117 N_B_c_118_n N_A_27_368#_c_471_n 0.0149468f $X=0.555 $Y=1.765 $X2=0 $Y2=0
cc_118 N_B_c_119_n N_A_27_368#_c_471_n 0.0128349f $X=1.005 $Y=1.765 $X2=0 $Y2=0
cc_119 N_B_c_120_n N_A_27_368#_c_473_n 0.0135069f $X=1.455 $Y=1.765 $X2=0 $Y2=0
cc_120 N_B_c_121_n N_A_27_368#_c_473_n 0.00915599f $X=1.98 $Y=1.765 $X2=0 $Y2=0
cc_121 N_B_c_120_n N_A_27_368#_c_475_n 6.61559e-19 $X=1.455 $Y=1.765 $X2=0 $Y2=0
cc_122 N_B_c_121_n N_A_27_368#_c_475_n 0.00735891f $X=1.98 $Y=1.765 $X2=0 $Y2=0
cc_123 N_B_c_119_n N_A_126_368#_c_539_n 0.0120074f $X=1.005 $Y=1.765 $X2=0 $Y2=0
cc_124 N_B_c_120_n N_A_126_368#_c_539_n 0.0127448f $X=1.455 $Y=1.765 $X2=0 $Y2=0
cc_125 B N_A_126_368#_c_539_n 0.0401171f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_126 N_B_c_117_n N_A_126_368#_c_539_n 0.001316f $X=1.98 $Y=1.557 $X2=0 $Y2=0
cc_127 N_B_c_121_n N_A_126_368#_c_536_n 0.0168026f $X=1.98 $Y=1.765 $X2=0 $Y2=0
cc_128 N_B_c_118_n N_A_126_368#_c_544_n 0.0102476f $X=0.555 $Y=1.765 $X2=0 $Y2=0
cc_129 N_B_c_119_n N_A_126_368#_c_544_n 0.0101535f $X=1.005 $Y=1.765 $X2=0 $Y2=0
cc_130 N_B_c_120_n N_A_126_368#_c_544_n 5.7282e-19 $X=1.455 $Y=1.765 $X2=0 $Y2=0
cc_131 B N_A_126_368#_c_544_n 0.0237598f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_132 N_B_c_117_n N_A_126_368#_c_544_n 0.00144338f $X=1.98 $Y=1.557 $X2=0 $Y2=0
cc_133 N_B_c_119_n N_A_126_368#_c_549_n 5.66701e-19 $X=1.005 $Y=1.765 $X2=0
+ $Y2=0
cc_134 N_B_c_120_n N_A_126_368#_c_549_n 0.0102531f $X=1.455 $Y=1.765 $X2=0 $Y2=0
cc_135 B N_A_126_368#_c_549_n 0.0229997f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_136 N_B_c_117_n N_A_126_368#_c_549_n 0.0034054f $X=1.98 $Y=1.557 $X2=0 $Y2=0
cc_137 N_B_M1003_g N_Y_c_604_n 4.71232e-19 $X=0.54 $Y=0.74 $X2=0 $Y2=0
cc_138 N_B_M1008_g N_Y_c_604_n 0.00959262f $X=0.995 $Y=0.74 $X2=0 $Y2=0
cc_139 N_B_M1024_g N_Y_c_604_n 6.3028e-19 $X=1.565 $Y=0.74 $X2=0 $Y2=0
cc_140 N_B_M1003_g N_Y_c_605_n 0.00190113f $X=0.54 $Y=0.74 $X2=0 $Y2=0
cc_141 N_B_M1008_g N_Y_c_605_n 0.0016171f $X=0.995 $Y=0.74 $X2=0 $Y2=0
cc_142 B N_Y_c_605_n 0.028235f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_143 N_B_c_117_n N_Y_c_605_n 0.00291196f $X=1.98 $Y=1.557 $X2=0 $Y2=0
cc_144 N_B_M1008_g N_Y_c_606_n 5.35648e-19 $X=0.995 $Y=0.74 $X2=0 $Y2=0
cc_145 N_B_M1024_g N_Y_c_606_n 0.00916462f $X=1.565 $Y=0.74 $X2=0 $Y2=0
cc_146 N_B_M1026_g N_Y_c_606_n 0.00924167f $X=1.995 $Y=0.74 $X2=0 $Y2=0
cc_147 N_B_c_120_n N_Y_c_630_n 3.30234e-19 $X=1.455 $Y=1.765 $X2=0 $Y2=0
cc_148 N_B_c_121_n N_Y_c_630_n 0.00698673f $X=1.98 $Y=1.765 $X2=0 $Y2=0
cc_149 N_B_M1008_g N_Y_c_613_n 0.0118691f $X=0.995 $Y=0.74 $X2=0 $Y2=0
cc_150 N_B_M1024_g N_Y_c_613_n 0.0118691f $X=1.565 $Y=0.74 $X2=0 $Y2=0
cc_151 B N_Y_c_613_n 0.0658285f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_152 N_B_c_117_n N_Y_c_613_n 0.00547601f $X=1.98 $Y=1.557 $X2=0 $Y2=0
cc_153 N_B_M1024_g N_Y_c_614_n 0.00220179f $X=1.565 $Y=0.74 $X2=0 $Y2=0
cc_154 N_B_M1026_g N_Y_c_614_n 0.0177513f $X=1.995 $Y=0.74 $X2=0 $Y2=0
cc_155 N_B_c_117_n N_Y_c_614_n 0.0024863f $X=1.98 $Y=1.557 $X2=0 $Y2=0
cc_156 N_B_M1024_g Y 8.28286e-19 $X=1.565 $Y=0.74 $X2=0 $Y2=0
cc_157 N_B_c_121_n Y 0.00135565f $X=1.98 $Y=1.765 $X2=0 $Y2=0
cc_158 N_B_M1026_g Y 0.00472643f $X=1.995 $Y=0.74 $X2=0 $Y2=0
cc_159 B Y 0.0265484f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_160 N_B_c_117_n Y 0.0109934f $X=1.98 $Y=1.557 $X2=0 $Y2=0
cc_161 N_B_c_118_n N_VPWR_c_748_n 0.00278271f $X=0.555 $Y=1.765 $X2=0 $Y2=0
cc_162 N_B_c_119_n N_VPWR_c_748_n 0.00278271f $X=1.005 $Y=1.765 $X2=0 $Y2=0
cc_163 N_B_c_120_n N_VPWR_c_748_n 0.00278271f $X=1.455 $Y=1.765 $X2=0 $Y2=0
cc_164 N_B_c_121_n N_VPWR_c_748_n 0.00279479f $X=1.98 $Y=1.765 $X2=0 $Y2=0
cc_165 N_B_c_118_n N_VPWR_c_742_n 0.00357472f $X=0.555 $Y=1.765 $X2=0 $Y2=0
cc_166 N_B_c_119_n N_VPWR_c_742_n 0.00353823f $X=1.005 $Y=1.765 $X2=0 $Y2=0
cc_167 N_B_c_120_n N_VPWR_c_742_n 0.00354498f $X=1.455 $Y=1.765 $X2=0 $Y2=0
cc_168 N_B_c_121_n N_VPWR_c_742_n 0.00353672f $X=1.98 $Y=1.765 $X2=0 $Y2=0
cc_169 N_B_M1003_g N_VGND_c_837_n 0.00549949f $X=0.54 $Y=0.74 $X2=0 $Y2=0
cc_170 B N_VGND_c_837_n 0.0239925f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_171 N_B_M1008_g N_VGND_c_838_n 0.00484409f $X=0.995 $Y=0.74 $X2=0 $Y2=0
cc_172 N_B_M1024_g N_VGND_c_838_n 0.00484409f $X=1.565 $Y=0.74 $X2=0 $Y2=0
cc_173 N_B_M1024_g N_VGND_c_839_n 0.00434272f $X=1.565 $Y=0.74 $X2=0 $Y2=0
cc_174 N_B_M1026_g N_VGND_c_839_n 0.00434272f $X=1.995 $Y=0.74 $X2=0 $Y2=0
cc_175 N_B_M1026_g N_VGND_c_840_n 0.00417204f $X=1.995 $Y=0.74 $X2=0 $Y2=0
cc_176 N_B_M1003_g N_VGND_c_848_n 0.00461464f $X=0.54 $Y=0.74 $X2=0 $Y2=0
cc_177 N_B_M1008_g N_VGND_c_848_n 0.00434272f $X=0.995 $Y=0.74 $X2=0 $Y2=0
cc_178 N_B_M1003_g N_VGND_c_852_n 0.00911596f $X=0.54 $Y=0.74 $X2=0 $Y2=0
cc_179 N_B_M1008_g N_VGND_c_852_n 0.00821539f $X=0.995 $Y=0.74 $X2=0 $Y2=0
cc_180 N_B_M1024_g N_VGND_c_852_n 0.00821294f $X=1.565 $Y=0.74 $X2=0 $Y2=0
cc_181 N_B_M1026_g N_VGND_c_852_n 0.00820772f $X=1.995 $Y=0.74 $X2=0 $Y2=0
cc_182 N_A_468_264#_M1013_g N_A_c_343_n 0.0161937f $X=3.855 $Y=0.74 $X2=-0.19
+ $Y2=-0.245
cc_183 N_A_468_264#_c_198_n N_A_c_350_n 2.77155e-19 $X=3.89 $Y=1.485 $X2=0 $Y2=0
cc_184 N_A_468_264#_c_208_n N_A_c_350_n 0.00865136f $X=6.785 $Y=1.805 $X2=0
+ $Y2=0
cc_185 N_A_468_264#_c_208_n N_A_c_351_n 0.00690449f $X=6.785 $Y=1.805 $X2=0
+ $Y2=0
cc_186 N_A_468_264#_c_208_n N_A_c_352_n 0.00690449f $X=6.785 $Y=1.805 $X2=0
+ $Y2=0
cc_187 N_A_468_264#_c_208_n N_A_c_353_n 0.0114581f $X=6.785 $Y=1.805 $X2=0 $Y2=0
cc_188 N_A_468_264#_c_209_n N_A_c_353_n 9.00694e-19 $X=6.95 $Y=1.985 $X2=0 $Y2=0
cc_189 N_A_468_264#_c_198_n N_A_c_348_n 0.00706164f $X=3.89 $Y=1.485 $X2=0 $Y2=0
cc_190 N_A_468_264#_c_208_n N_A_c_348_n 0.0357388f $X=6.785 $Y=1.805 $X2=0 $Y2=0
cc_191 N_A_468_264#_c_202_n N_A_c_348_n 0.0161937f $X=3.78 $Y=1.542 $X2=0 $Y2=0
cc_192 N_A_468_264#_M1013_g N_A_c_349_n 4.72901e-19 $X=3.855 $Y=0.74 $X2=0 $Y2=0
cc_193 N_A_468_264#_c_198_n N_A_c_349_n 0.014508f $X=3.89 $Y=1.485 $X2=0 $Y2=0
cc_194 N_A_468_264#_c_208_n N_A_c_349_n 0.160908f $X=6.785 $Y=1.805 $X2=0 $Y2=0
cc_195 N_A_468_264#_c_201_n N_C_N_c_432_n 0.0094203f $X=7.4 $Y=0.5 $X2=-0.19
+ $Y2=-0.245
cc_196 N_A_468_264#_c_208_n N_C_N_c_435_n 0.00946684f $X=6.785 $Y=1.805 $X2=0
+ $Y2=0
cc_197 N_A_468_264#_c_209_n N_C_N_c_435_n 0.0120477f $X=6.95 $Y=1.985 $X2=0
+ $Y2=0
cc_198 N_A_468_264#_c_233_p N_C_N_c_435_n 0.00109449f $X=6.92 $Y=1.805 $X2=0
+ $Y2=0
cc_199 N_A_468_264#_c_209_n N_C_N_c_436_n 8.84821e-19 $X=6.95 $Y=1.985 $X2=0
+ $Y2=0
cc_200 N_A_468_264#_c_210_n N_C_N_c_436_n 0.0113224f $X=7.395 $Y=1.805 $X2=0
+ $Y2=0
cc_201 N_A_468_264#_c_208_n C_N 0.00134249f $X=6.785 $Y=1.805 $X2=0 $Y2=0
cc_202 N_A_468_264#_c_210_n C_N 0.00279147f $X=7.395 $Y=1.805 $X2=0 $Y2=0
cc_203 N_A_468_264#_c_200_n C_N 0.0183654f $X=7.48 $Y=1.72 $X2=0 $Y2=0
cc_204 N_A_468_264#_c_233_p C_N 0.0218449f $X=6.92 $Y=1.805 $X2=0 $Y2=0
cc_205 N_A_468_264#_c_201_n C_N 0.0286132f $X=7.4 $Y=0.5 $X2=0 $Y2=0
cc_206 N_A_468_264#_c_208_n N_C_N_c_434_n 0.00914245f $X=6.785 $Y=1.805 $X2=0
+ $Y2=0
cc_207 N_A_468_264#_c_210_n N_C_N_c_434_n 0.0103356f $X=7.395 $Y=1.805 $X2=0
+ $Y2=0
cc_208 N_A_468_264#_c_200_n N_C_N_c_434_n 0.0162405f $X=7.48 $Y=1.72 $X2=0 $Y2=0
cc_209 N_A_468_264#_c_233_p N_C_N_c_434_n 0.0113514f $X=6.92 $Y=1.805 $X2=0
+ $Y2=0
cc_210 N_A_468_264#_c_201_n N_C_N_c_434_n 0.0144772f $X=7.4 $Y=0.5 $X2=0 $Y2=0
cc_211 N_A_468_264#_c_198_n N_A_27_368#_M1025_s 0.00435851f $X=3.89 $Y=1.485
+ $X2=0 $Y2=0
cc_212 N_A_468_264#_c_205_n N_A_27_368#_c_485_n 0.00871022f $X=3.33 $Y=1.765
+ $X2=0 $Y2=0
cc_213 N_A_468_264#_c_206_n N_A_27_368#_c_485_n 0.00928899f $X=3.78 $Y=1.765
+ $X2=0 $Y2=0
cc_214 N_A_468_264#_c_203_n N_A_27_368#_c_475_n 0.0083814f $X=2.43 $Y=1.765
+ $X2=0 $Y2=0
cc_215 N_A_468_264#_c_204_n N_A_27_368#_c_475_n 0.00133759f $X=2.88 $Y=1.765
+ $X2=0 $Y2=0
cc_216 N_A_468_264#_c_203_n N_A_27_368#_c_489_n 0.00925828f $X=2.43 $Y=1.765
+ $X2=0 $Y2=0
cc_217 N_A_468_264#_c_204_n N_A_27_368#_c_489_n 0.00871022f $X=2.88 $Y=1.765
+ $X2=0 $Y2=0
cc_218 N_A_468_264#_c_203_n N_A_27_368#_c_491_n 4.70346e-19 $X=2.43 $Y=1.765
+ $X2=0 $Y2=0
cc_219 N_A_468_264#_c_204_n N_A_27_368#_c_491_n 0.00339823f $X=2.88 $Y=1.765
+ $X2=0 $Y2=0
cc_220 N_A_468_264#_c_205_n N_A_27_368#_c_491_n 0.00339823f $X=3.33 $Y=1.765
+ $X2=0 $Y2=0
cc_221 N_A_468_264#_c_206_n N_A_27_368#_c_491_n 4.70346e-19 $X=3.78 $Y=1.765
+ $X2=0 $Y2=0
cc_222 N_A_468_264#_c_205_n N_A_27_368#_c_476_n 5.54287e-19 $X=3.33 $Y=1.765
+ $X2=0 $Y2=0
cc_223 N_A_468_264#_c_206_n N_A_27_368#_c_476_n 0.00385514f $X=3.78 $Y=1.765
+ $X2=0 $Y2=0
cc_224 N_A_468_264#_c_208_n N_A_126_368#_M1007_d 0.00196679f $X=6.785 $Y=1.805
+ $X2=0 $Y2=0
cc_225 N_A_468_264#_c_208_n N_A_126_368#_M1019_d 0.00197722f $X=6.785 $Y=1.805
+ $X2=0 $Y2=0
cc_226 N_A_468_264#_c_203_n N_A_126_368#_c_536_n 0.0106672f $X=2.43 $Y=1.765
+ $X2=0 $Y2=0
cc_227 N_A_468_264#_c_204_n N_A_126_368#_c_536_n 0.0107326f $X=2.88 $Y=1.765
+ $X2=0 $Y2=0
cc_228 N_A_468_264#_c_205_n N_A_126_368#_c_536_n 0.0107326f $X=3.33 $Y=1.765
+ $X2=0 $Y2=0
cc_229 N_A_468_264#_c_206_n N_A_126_368#_c_536_n 0.0144433f $X=3.78 $Y=1.765
+ $X2=0 $Y2=0
cc_230 N_A_468_264#_c_198_n N_A_126_368#_c_536_n 0.0173386f $X=3.89 $Y=1.485
+ $X2=0 $Y2=0
cc_231 N_A_468_264#_c_208_n N_A_126_368#_c_536_n 0.0234885f $X=6.785 $Y=1.805
+ $X2=0 $Y2=0
cc_232 N_A_468_264#_c_208_n N_A_126_368#_c_561_n 0.0343572f $X=6.785 $Y=1.805
+ $X2=0 $Y2=0
cc_233 N_A_468_264#_c_208_n N_A_126_368#_c_562_n 0.0162332f $X=6.785 $Y=1.805
+ $X2=0 $Y2=0
cc_234 N_A_468_264#_c_208_n N_A_126_368#_c_563_n 0.0193054f $X=6.785 $Y=1.805
+ $X2=0 $Y2=0
cc_235 N_A_468_264#_M1000_g N_Y_c_606_n 8.87957e-19 $X=2.495 $Y=0.74 $X2=0 $Y2=0
cc_236 N_A_468_264#_M1000_g N_Y_c_607_n 0.0151238f $X=2.495 $Y=0.74 $X2=0 $Y2=0
cc_237 N_A_468_264#_c_198_n N_Y_c_607_n 0.00334513f $X=3.89 $Y=1.485 $X2=0 $Y2=0
cc_238 N_A_468_264#_c_202_n N_Y_c_607_n 0.0024651f $X=3.78 $Y=1.542 $X2=0 $Y2=0
cc_239 N_A_468_264#_c_203_n N_Y_c_618_n 0.0129339f $X=2.43 $Y=1.765 $X2=0 $Y2=0
cc_240 N_A_468_264#_c_204_n N_Y_c_618_n 0.0110106f $X=2.88 $Y=1.765 $X2=0 $Y2=0
cc_241 N_A_468_264#_c_205_n N_Y_c_618_n 0.0110106f $X=3.33 $Y=1.765 $X2=0 $Y2=0
cc_242 N_A_468_264#_c_206_n N_Y_c_618_n 0.00959754f $X=3.78 $Y=1.765 $X2=0 $Y2=0
cc_243 N_A_468_264#_c_198_n N_Y_c_618_n 0.0906723f $X=3.89 $Y=1.485 $X2=0 $Y2=0
cc_244 N_A_468_264#_c_202_n N_Y_c_618_n 0.0237691f $X=3.78 $Y=1.542 $X2=0 $Y2=0
cc_245 N_A_468_264#_M1000_g N_Y_c_608_n 3.92313e-19 $X=2.495 $Y=0.74 $X2=0 $Y2=0
cc_246 N_A_468_264#_M1001_g N_Y_c_608_n 3.92313e-19 $X=2.925 $Y=0.74 $X2=0 $Y2=0
cc_247 N_A_468_264#_M1001_g N_Y_c_609_n 0.0131239f $X=2.925 $Y=0.74 $X2=0 $Y2=0
cc_248 N_A_468_264#_M1009_g N_Y_c_609_n 0.0115433f $X=3.425 $Y=0.74 $X2=0 $Y2=0
cc_249 N_A_468_264#_c_198_n N_Y_c_609_n 0.0500092f $X=3.89 $Y=1.485 $X2=0 $Y2=0
cc_250 N_A_468_264#_c_202_n N_Y_c_609_n 0.00385261f $X=3.78 $Y=1.542 $X2=0 $Y2=0
cc_251 N_A_468_264#_M1001_g N_Y_c_610_n 4.13007e-19 $X=2.925 $Y=0.74 $X2=0 $Y2=0
cc_252 N_A_468_264#_M1009_g N_Y_c_610_n 0.00721977f $X=3.425 $Y=0.74 $X2=0 $Y2=0
cc_253 N_A_468_264#_M1013_g N_Y_c_610_n 0.00834185f $X=3.855 $Y=0.74 $X2=0 $Y2=0
cc_254 N_A_468_264#_M1013_g N_Y_c_663_n 0.0120704f $X=3.855 $Y=0.74 $X2=0 $Y2=0
cc_255 N_A_468_264#_c_198_n N_Y_c_663_n 0.0202341f $X=3.89 $Y=1.485 $X2=0 $Y2=0
cc_256 N_A_468_264#_c_208_n N_Y_c_663_n 0.00575327f $X=6.785 $Y=1.805 $X2=0
+ $Y2=0
cc_257 N_A_468_264#_M1013_g N_Y_c_611_n 6.03013e-19 $X=3.855 $Y=0.74 $X2=0 $Y2=0
cc_258 N_A_468_264#_M1000_g N_Y_c_614_n 8.44859e-19 $X=2.495 $Y=0.74 $X2=0 $Y2=0
cc_259 N_A_468_264#_c_198_n N_Y_c_615_n 0.0143381f $X=3.89 $Y=1.485 $X2=0 $Y2=0
cc_260 N_A_468_264#_c_202_n N_Y_c_615_n 0.00232957f $X=3.78 $Y=1.542 $X2=0 $Y2=0
cc_261 N_A_468_264#_M1001_g N_Y_c_616_n 4.68741e-19 $X=2.925 $Y=0.74 $X2=0 $Y2=0
cc_262 N_A_468_264#_M1009_g N_Y_c_616_n 0.00330557f $X=3.425 $Y=0.74 $X2=0 $Y2=0
cc_263 N_A_468_264#_M1013_g N_Y_c_616_n 0.00342047f $X=3.855 $Y=0.74 $X2=0 $Y2=0
cc_264 N_A_468_264#_c_198_n N_Y_c_616_n 0.0276081f $X=3.89 $Y=1.485 $X2=0 $Y2=0
cc_265 N_A_468_264#_c_202_n N_Y_c_616_n 0.00232957f $X=3.78 $Y=1.542 $X2=0 $Y2=0
cc_266 N_A_468_264#_c_203_n Y 0.00133661f $X=2.43 $Y=1.765 $X2=0 $Y2=0
cc_267 N_A_468_264#_M1000_g Y 0.00326736f $X=2.495 $Y=0.74 $X2=0 $Y2=0
cc_268 N_A_468_264#_c_198_n Y 0.0172568f $X=3.89 $Y=1.485 $X2=0 $Y2=0
cc_269 N_A_468_264#_c_202_n Y 0.00640982f $X=3.78 $Y=1.542 $X2=0 $Y2=0
cc_270 N_A_468_264#_c_208_n N_VPWR_M1007_s 0.00383277f $X=6.785 $Y=1.805
+ $X2=-0.19 $Y2=-0.245
cc_271 N_A_468_264#_c_208_n N_VPWR_M1017_s 0.00198204f $X=6.785 $Y=1.805 $X2=0
+ $Y2=0
cc_272 N_A_468_264#_c_208_n N_VPWR_M1021_s 0.00391969f $X=6.785 $Y=1.805 $X2=0
+ $Y2=0
cc_273 N_A_468_264#_c_210_n N_VPWR_M1005_s 0.00286151f $X=7.395 $Y=1.805 $X2=0
+ $Y2=0
cc_274 N_A_468_264#_c_206_n N_VPWR_c_743_n 0.00411922f $X=3.78 $Y=1.765 $X2=0
+ $Y2=0
cc_275 N_A_468_264#_c_208_n N_VPWR_c_745_n 0.0249771f $X=6.785 $Y=1.805 $X2=0
+ $Y2=0
cc_276 N_A_468_264#_c_209_n N_VPWR_c_745_n 0.0424201f $X=6.95 $Y=1.985 $X2=0
+ $Y2=0
cc_277 N_A_468_264#_c_209_n N_VPWR_c_747_n 0.0236749f $X=6.95 $Y=1.985 $X2=0
+ $Y2=0
cc_278 N_A_468_264#_c_210_n N_VPWR_c_747_n 0.0234519f $X=7.395 $Y=1.805 $X2=0
+ $Y2=0
cc_279 N_A_468_264#_c_203_n N_VPWR_c_748_n 0.00317151f $X=2.43 $Y=1.765 $X2=0
+ $Y2=0
cc_280 N_A_468_264#_c_204_n N_VPWR_c_748_n 0.00318204f $X=2.88 $Y=1.765 $X2=0
+ $Y2=0
cc_281 N_A_468_264#_c_205_n N_VPWR_c_748_n 0.00318204f $X=3.33 $Y=1.765 $X2=0
+ $Y2=0
cc_282 N_A_468_264#_c_206_n N_VPWR_c_748_n 0.00319263f $X=3.78 $Y=1.765 $X2=0
+ $Y2=0
cc_283 N_A_468_264#_c_209_n N_VPWR_c_751_n 0.00545158f $X=6.95 $Y=1.985 $X2=0
+ $Y2=0
cc_284 N_A_468_264#_c_203_n N_VPWR_c_742_n 0.00395545f $X=2.43 $Y=1.765 $X2=0
+ $Y2=0
cc_285 N_A_468_264#_c_204_n N_VPWR_c_742_n 0.0039788f $X=2.88 $Y=1.765 $X2=0
+ $Y2=0
cc_286 N_A_468_264#_c_205_n N_VPWR_c_742_n 0.0039788f $X=3.33 $Y=1.765 $X2=0
+ $Y2=0
cc_287 N_A_468_264#_c_206_n N_VPWR_c_742_n 0.00401657f $X=3.78 $Y=1.765 $X2=0
+ $Y2=0
cc_288 N_A_468_264#_c_209_n N_VPWR_c_742_n 0.00814593f $X=6.95 $Y=1.985 $X2=0
+ $Y2=0
cc_289 N_A_468_264#_M1000_g N_VGND_c_840_n 0.0100169f $X=2.495 $Y=0.74 $X2=0
+ $Y2=0
cc_290 N_A_468_264#_M1001_g N_VGND_c_840_n 4.62684e-19 $X=2.925 $Y=0.74 $X2=0
+ $Y2=0
cc_291 N_A_468_264#_M1000_g N_VGND_c_841_n 4.62684e-19 $X=2.495 $Y=0.74 $X2=0
+ $Y2=0
cc_292 N_A_468_264#_M1001_g N_VGND_c_841_n 0.0100169f $X=2.925 $Y=0.74 $X2=0
+ $Y2=0
cc_293 N_A_468_264#_M1009_g N_VGND_c_841_n 0.00417204f $X=3.425 $Y=0.74 $X2=0
+ $Y2=0
cc_294 N_A_468_264#_M1013_g N_VGND_c_842_n 0.00405455f $X=3.855 $Y=0.74 $X2=0
+ $Y2=0
cc_295 N_A_468_264#_c_201_n N_VGND_c_845_n 0.0284697f $X=7.4 $Y=0.5 $X2=0 $Y2=0
cc_296 N_A_468_264#_M1000_g N_VGND_c_849_n 0.00383152f $X=2.495 $Y=0.74 $X2=0
+ $Y2=0
cc_297 N_A_468_264#_M1001_g N_VGND_c_849_n 0.00383152f $X=2.925 $Y=0.74 $X2=0
+ $Y2=0
cc_298 N_A_468_264#_M1009_g N_VGND_c_850_n 0.00434272f $X=3.425 $Y=0.74 $X2=0
+ $Y2=0
cc_299 N_A_468_264#_M1013_g N_VGND_c_850_n 0.00434272f $X=3.855 $Y=0.74 $X2=0
+ $Y2=0
cc_300 N_A_468_264#_c_199_n N_VGND_c_851_n 0.00758556f $X=7.48 $Y=1.01 $X2=0
+ $Y2=0
cc_301 N_A_468_264#_c_201_n N_VGND_c_851_n 0.0349297f $X=7.4 $Y=0.5 $X2=0 $Y2=0
cc_302 N_A_468_264#_M1000_g N_VGND_c_852_n 0.0075754f $X=2.495 $Y=0.74 $X2=0
+ $Y2=0
cc_303 N_A_468_264#_M1001_g N_VGND_c_852_n 0.0075754f $X=2.925 $Y=0.74 $X2=0
+ $Y2=0
cc_304 N_A_468_264#_M1009_g N_VGND_c_852_n 0.00820718f $X=3.425 $Y=0.74 $X2=0
+ $Y2=0
cc_305 N_A_468_264#_M1013_g N_VGND_c_852_n 0.00821312f $X=3.855 $Y=0.74 $X2=0
+ $Y2=0
cc_306 N_A_468_264#_c_199_n N_VGND_c_852_n 0.00627867f $X=7.48 $Y=1.01 $X2=0
+ $Y2=0
cc_307 N_A_468_264#_c_201_n N_VGND_c_852_n 0.0289999f $X=7.4 $Y=0.5 $X2=0 $Y2=0
cc_308 N_A_c_346_n N_C_N_c_432_n 0.0116655f $X=6.055 $Y=1.22 $X2=-0.19
+ $Y2=-0.245
cc_309 A N_C_N_c_432_n 0.00650444f $X=6.395 $Y=1.21 $X2=-0.19 $Y2=-0.245
cc_310 N_A_c_353_n N_C_N_c_435_n 0.0214491f $X=6.14 $Y=1.765 $X2=0 $Y2=0
cc_311 A C_N 0.030054f $X=6.395 $Y=1.21 $X2=0 $Y2=0
cc_312 A N_C_N_c_434_n 0.0102326f $X=6.395 $Y=1.21 $X2=0 $Y2=0
cc_313 N_A_c_348_n N_C_N_c_434_n 0.0244096f $X=6.055 $Y=1.492 $X2=0 $Y2=0
cc_314 N_A_c_350_n N_A_126_368#_c_536_n 0.0110088f $X=4.79 $Y=1.765 $X2=0 $Y2=0
cc_315 N_A_c_350_n N_A_126_368#_c_537_n 0.00471036f $X=4.79 $Y=1.765 $X2=0 $Y2=0
cc_316 N_A_c_351_n N_A_126_368#_c_561_n 0.0126853f $X=5.24 $Y=1.765 $X2=0 $Y2=0
cc_317 N_A_c_352_n N_A_126_368#_c_561_n 0.0126342f $X=5.69 $Y=1.765 $X2=0 $Y2=0
cc_318 N_A_c_353_n N_A_126_368#_c_562_n 0.00185023f $X=6.14 $Y=1.765 $X2=0 $Y2=0
cc_319 N_A_c_352_n N_A_126_368#_c_538_n 2.33402e-19 $X=5.69 $Y=1.765 $X2=0 $Y2=0
cc_320 N_A_c_353_n N_A_126_368#_c_538_n 0.00780419f $X=6.14 $Y=1.765 $X2=0 $Y2=0
cc_321 N_A_c_350_n N_A_126_368#_c_563_n 0.014276f $X=4.79 $Y=1.765 $X2=0 $Y2=0
cc_322 N_A_c_351_n N_A_126_368#_c_563_n 0.00579718f $X=5.24 $Y=1.765 $X2=0 $Y2=0
cc_323 N_A_c_343_n N_Y_c_610_n 6.03013e-19 $X=4.425 $Y=1.22 $X2=0 $Y2=0
cc_324 N_A_c_343_n N_Y_c_663_n 0.0127102f $X=4.425 $Y=1.22 $X2=0 $Y2=0
cc_325 N_A_c_349_n N_Y_c_663_n 0.00246555f $X=6.365 $Y=1.365 $X2=0 $Y2=0
cc_326 N_A_c_343_n N_Y_c_611_n 0.00834185f $X=4.425 $Y=1.22 $X2=0 $Y2=0
cc_327 N_A_c_344_n N_Y_c_611_n 0.00907544f $X=4.855 $Y=1.22 $X2=0 $Y2=0
cc_328 N_A_c_345_n N_Y_c_611_n 8.95441e-19 $X=5.555 $Y=1.22 $X2=0 $Y2=0
cc_329 N_A_c_344_n N_Y_c_685_n 0.0121454f $X=4.855 $Y=1.22 $X2=0 $Y2=0
cc_330 N_A_c_345_n N_Y_c_685_n 0.0128634f $X=5.555 $Y=1.22 $X2=0 $Y2=0
cc_331 N_A_c_348_n N_Y_c_685_n 0.0140774f $X=6.055 $Y=1.492 $X2=0 $Y2=0
cc_332 N_A_c_349_n N_Y_c_685_n 0.0783501f $X=6.365 $Y=1.365 $X2=0 $Y2=0
cc_333 N_A_c_344_n N_Y_c_612_n 8.95441e-19 $X=4.855 $Y=1.22 $X2=0 $Y2=0
cc_334 N_A_c_345_n N_Y_c_612_n 0.00908017f $X=5.555 $Y=1.22 $X2=0 $Y2=0
cc_335 N_A_c_346_n N_Y_c_612_n 0.00282572f $X=6.055 $Y=1.22 $X2=0 $Y2=0
cc_336 N_A_c_343_n N_Y_c_616_n 4.52963e-19 $X=4.425 $Y=1.22 $X2=0 $Y2=0
cc_337 N_A_c_343_n N_Y_c_693_n 7.18016e-19 $X=4.425 $Y=1.22 $X2=0 $Y2=0
cc_338 N_A_c_344_n N_Y_c_693_n 7.18016e-19 $X=4.855 $Y=1.22 $X2=0 $Y2=0
cc_339 N_A_c_348_n N_Y_c_693_n 0.00232761f $X=6.055 $Y=1.492 $X2=0 $Y2=0
cc_340 N_A_c_349_n N_Y_c_693_n 0.021954f $X=6.365 $Y=1.365 $X2=0 $Y2=0
cc_341 N_A_c_350_n N_VPWR_c_743_n 0.00942993f $X=4.79 $Y=1.765 $X2=0 $Y2=0
cc_342 N_A_c_351_n N_VPWR_c_743_n 4.21336e-19 $X=5.24 $Y=1.765 $X2=0 $Y2=0
cc_343 N_A_c_350_n N_VPWR_c_744_n 4.73012e-19 $X=4.79 $Y=1.765 $X2=0 $Y2=0
cc_344 N_A_c_351_n N_VPWR_c_744_n 0.00982773f $X=5.24 $Y=1.765 $X2=0 $Y2=0
cc_345 N_A_c_352_n N_VPWR_c_744_n 0.00963862f $X=5.69 $Y=1.765 $X2=0 $Y2=0
cc_346 N_A_c_353_n N_VPWR_c_744_n 4.7857e-19 $X=6.14 $Y=1.765 $X2=0 $Y2=0
cc_347 N_A_c_353_n N_VPWR_c_745_n 0.0113505f $X=6.14 $Y=1.765 $X2=0 $Y2=0
cc_348 N_A_c_350_n N_VPWR_c_749_n 0.00413917f $X=4.79 $Y=1.765 $X2=0 $Y2=0
cc_349 N_A_c_351_n N_VPWR_c_749_n 0.00413917f $X=5.24 $Y=1.765 $X2=0 $Y2=0
cc_350 N_A_c_352_n N_VPWR_c_750_n 0.00413917f $X=5.69 $Y=1.765 $X2=0 $Y2=0
cc_351 N_A_c_353_n N_VPWR_c_750_n 0.00445475f $X=6.14 $Y=1.765 $X2=0 $Y2=0
cc_352 N_A_c_350_n N_VPWR_c_742_n 0.00817726f $X=4.79 $Y=1.765 $X2=0 $Y2=0
cc_353 N_A_c_351_n N_VPWR_c_742_n 0.00817726f $X=5.24 $Y=1.765 $X2=0 $Y2=0
cc_354 N_A_c_352_n N_VPWR_c_742_n 0.00817726f $X=5.69 $Y=1.765 $X2=0 $Y2=0
cc_355 N_A_c_353_n N_VPWR_c_742_n 0.00861625f $X=6.14 $Y=1.765 $X2=0 $Y2=0
cc_356 N_A_c_343_n N_VGND_c_842_n 0.00405455f $X=4.425 $Y=1.22 $X2=0 $Y2=0
cc_357 N_A_c_343_n N_VGND_c_843_n 0.00434272f $X=4.425 $Y=1.22 $X2=0 $Y2=0
cc_358 N_A_c_344_n N_VGND_c_843_n 0.00434272f $X=4.855 $Y=1.22 $X2=0 $Y2=0
cc_359 N_A_c_344_n N_VGND_c_844_n 0.00460818f $X=4.855 $Y=1.22 $X2=0 $Y2=0
cc_360 N_A_c_345_n N_VGND_c_844_n 0.00460818f $X=5.555 $Y=1.22 $X2=0 $Y2=0
cc_361 N_A_c_345_n N_VGND_c_845_n 5.39035e-19 $X=5.555 $Y=1.22 $X2=0 $Y2=0
cc_362 N_A_c_346_n N_VGND_c_845_n 0.011573f $X=6.055 $Y=1.22 $X2=0 $Y2=0
cc_363 A N_VGND_c_845_n 0.00553831f $X=6.395 $Y=1.21 $X2=0 $Y2=0
cc_364 N_A_c_348_n N_VGND_c_845_n 3.80797e-19 $X=6.055 $Y=1.492 $X2=0 $Y2=0
cc_365 N_A_c_349_n N_VGND_c_845_n 0.016837f $X=6.365 $Y=1.365 $X2=0 $Y2=0
cc_366 N_A_c_345_n N_VGND_c_846_n 0.00434272f $X=5.555 $Y=1.22 $X2=0 $Y2=0
cc_367 N_A_c_346_n N_VGND_c_846_n 0.00383152f $X=6.055 $Y=1.22 $X2=0 $Y2=0
cc_368 N_A_c_343_n N_VGND_c_852_n 0.00821312f $X=4.425 $Y=1.22 $X2=0 $Y2=0
cc_369 N_A_c_344_n N_VGND_c_852_n 0.00822177f $X=4.855 $Y=1.22 $X2=0 $Y2=0
cc_370 N_A_c_345_n N_VGND_c_852_n 0.00822835f $X=5.555 $Y=1.22 $X2=0 $Y2=0
cc_371 N_A_c_346_n N_VGND_c_852_n 0.00758198f $X=6.055 $Y=1.22 $X2=0 $Y2=0
cc_372 N_C_N_c_435_n N_VPWR_c_745_n 0.00791943f $X=6.725 $Y=1.765 $X2=0 $Y2=0
cc_373 N_C_N_c_435_n N_VPWR_c_747_n 5.91896e-19 $X=6.725 $Y=1.765 $X2=0 $Y2=0
cc_374 N_C_N_c_436_n N_VPWR_c_747_n 0.0114144f $X=7.175 $Y=1.765 $X2=0 $Y2=0
cc_375 N_C_N_c_435_n N_VPWR_c_751_n 0.00393873f $X=6.725 $Y=1.765 $X2=0 $Y2=0
cc_376 N_C_N_c_436_n N_VPWR_c_751_n 0.00361294f $X=7.175 $Y=1.765 $X2=0 $Y2=0
cc_377 N_C_N_c_435_n N_VPWR_c_742_n 0.00462577f $X=6.725 $Y=1.765 $X2=0 $Y2=0
cc_378 N_C_N_c_436_n N_VPWR_c_742_n 0.00419404f $X=7.175 $Y=1.765 $X2=0 $Y2=0
cc_379 N_C_N_c_432_n N_VGND_c_845_n 0.00661609f $X=6.555 $Y=1.22 $X2=0 $Y2=0
cc_380 N_C_N_c_432_n N_VGND_c_851_n 0.00433162f $X=6.555 $Y=1.22 $X2=0 $Y2=0
cc_381 N_C_N_c_432_n N_VGND_c_852_n 0.00822119f $X=6.555 $Y=1.22 $X2=0 $Y2=0
cc_382 N_A_27_368#_c_471_n N_A_126_368#_M1010_s 0.00197722f $X=1.145 $Y=2.99
+ $X2=-0.19 $Y2=1.66
cc_383 N_A_27_368#_c_473_n N_A_126_368#_M1014_s 0.00281931f $X=2.04 $Y=2.99
+ $X2=0 $Y2=0
cc_384 N_A_27_368#_M1012_d N_A_126_368#_c_539_n 0.00408911f $X=1.08 $Y=1.84
+ $X2=0 $Y2=0
cc_385 N_A_27_368#_c_500_p N_A_126_368#_c_539_n 0.0136682f $X=1.23 $Y=2.455
+ $X2=0 $Y2=0
cc_386 N_A_27_368#_M1016_d N_A_126_368#_c_536_n 0.00395503f $X=2.055 $Y=1.84
+ $X2=0 $Y2=0
cc_387 N_A_27_368#_M1020_s N_A_126_368#_c_536_n 0.00378973f $X=2.955 $Y=1.84
+ $X2=0 $Y2=0
cc_388 N_A_27_368#_M1025_s N_A_126_368#_c_536_n 0.00712616f $X=3.855 $Y=1.84
+ $X2=0 $Y2=0
cc_389 N_A_27_368#_c_473_n N_A_126_368#_c_536_n 0.0038303f $X=2.04 $Y=2.99 $X2=0
+ $Y2=0
cc_390 N_A_27_368#_c_475_n N_A_126_368#_c_536_n 0.0167456f $X=2.205 $Y=2.665
+ $X2=0 $Y2=0
cc_391 N_A_27_368#_c_489_n N_A_126_368#_c_536_n 0.079835f $X=2.94 $Y=2.745 $X2=0
+ $Y2=0
cc_392 N_A_27_368#_c_476_n N_A_126_368#_c_536_n 0.0207579f $X=4.005 $Y=2.665
+ $X2=0 $Y2=0
cc_393 N_A_27_368#_c_471_n N_A_126_368#_c_544_n 0.0160777f $X=1.145 $Y=2.99
+ $X2=0 $Y2=0
cc_394 N_A_27_368#_c_500_p N_A_126_368#_c_544_n 0.0289859f $X=1.23 $Y=2.455
+ $X2=0 $Y2=0
cc_395 N_A_27_368#_c_500_p N_A_126_368#_c_549_n 0.0284797f $X=1.23 $Y=2.455
+ $X2=0 $Y2=0
cc_396 N_A_27_368#_c_473_n N_A_126_368#_c_549_n 0.0201846f $X=2.04 $Y=2.99 $X2=0
+ $Y2=0
cc_397 N_A_27_368#_c_489_n N_Y_M1018_d 0.00501057f $X=2.94 $Y=2.745 $X2=0 $Y2=0
cc_398 N_A_27_368#_c_485_n N_Y_M1023_d 0.00501057f $X=3.84 $Y=2.665 $X2=0 $Y2=0
cc_399 N_A_27_368#_M1016_d N_Y_c_630_n 0.00180824f $X=2.055 $Y=1.84 $X2=0 $Y2=0
cc_400 N_A_27_368#_M1016_d N_Y_c_618_n 2.37238e-19 $X=2.055 $Y=1.84 $X2=0 $Y2=0
cc_401 N_A_27_368#_M1020_s N_Y_c_618_n 0.00200574f $X=2.955 $Y=1.84 $X2=0 $Y2=0
cc_402 N_A_27_368#_c_476_n N_VPWR_c_743_n 0.0222482f $X=4.005 $Y=2.665 $X2=0
+ $Y2=0
cc_403 N_A_27_368#_c_471_n N_VPWR_c_748_n 0.0441612f $X=1.145 $Y=2.99 $X2=0
+ $Y2=0
cc_404 N_A_27_368#_c_472_n N_VPWR_c_748_n 0.0236566f $X=0.445 $Y=2.99 $X2=0
+ $Y2=0
cc_405 N_A_27_368#_c_473_n N_VPWR_c_748_n 0.0458445f $X=2.04 $Y=2.99 $X2=0 $Y2=0
cc_406 N_A_27_368#_c_485_n N_VPWR_c_748_n 0.00999853f $X=3.84 $Y=2.665 $X2=0
+ $Y2=0
cc_407 N_A_27_368#_c_474_n N_VPWR_c_748_n 0.0121867f $X=1.23 $Y=2.99 $X2=0 $Y2=0
cc_408 N_A_27_368#_c_475_n N_VPWR_c_748_n 0.0228653f $X=2.205 $Y=2.665 $X2=0
+ $Y2=0
cc_409 N_A_27_368#_c_489_n N_VPWR_c_748_n 0.00999853f $X=2.94 $Y=2.745 $X2=0
+ $Y2=0
cc_410 N_A_27_368#_c_491_n N_VPWR_c_748_n 0.00888684f $X=3.27 $Y=2.745 $X2=0
+ $Y2=0
cc_411 N_A_27_368#_c_476_n N_VPWR_c_748_n 0.00970993f $X=4.005 $Y=2.665 $X2=0
+ $Y2=0
cc_412 N_A_27_368#_c_471_n N_VPWR_c_742_n 0.0249452f $X=1.145 $Y=2.99 $X2=0
+ $Y2=0
cc_413 N_A_27_368#_c_472_n N_VPWR_c_742_n 0.0128296f $X=0.445 $Y=2.99 $X2=0
+ $Y2=0
cc_414 N_A_27_368#_c_473_n N_VPWR_c_742_n 0.0259575f $X=2.04 $Y=2.99 $X2=0 $Y2=0
cc_415 N_A_27_368#_c_485_n N_VPWR_c_742_n 0.0156417f $X=3.84 $Y=2.665 $X2=0
+ $Y2=0
cc_416 N_A_27_368#_c_474_n N_VPWR_c_742_n 0.00660921f $X=1.23 $Y=2.99 $X2=0
+ $Y2=0
cc_417 N_A_27_368#_c_475_n N_VPWR_c_742_n 0.0125201f $X=2.205 $Y=2.665 $X2=0
+ $Y2=0
cc_418 N_A_27_368#_c_489_n N_VPWR_c_742_n 0.0156417f $X=2.94 $Y=2.745 $X2=0
+ $Y2=0
cc_419 N_A_27_368#_c_491_n N_VPWR_c_742_n 0.0111774f $X=3.27 $Y=2.745 $X2=0
+ $Y2=0
cc_420 N_A_27_368#_c_476_n N_VPWR_c_742_n 0.0112088f $X=4.005 $Y=2.665 $X2=0
+ $Y2=0
cc_421 N_A_126_368#_c_536_n N_Y_M1018_d 0.00378973f $X=4.795 $Y=2.325 $X2=0
+ $Y2=0
cc_422 N_A_126_368#_c_536_n N_Y_M1023_d 0.00378973f $X=4.795 $Y=2.325 $X2=0
+ $Y2=0
cc_423 N_A_126_368#_c_536_n N_Y_c_630_n 0.0139811f $X=4.795 $Y=2.325 $X2=0 $Y2=0
cc_424 N_A_126_368#_c_536_n N_Y_c_618_n 0.0757524f $X=4.795 $Y=2.325 $X2=0 $Y2=0
cc_425 N_A_126_368#_c_536_n N_VPWR_M1007_s 0.00685669f $X=4.795 $Y=2.325
+ $X2=-0.19 $Y2=1.66
cc_426 N_A_126_368#_c_561_n N_VPWR_M1017_s 0.00385521f $X=5.81 $Y=2.145 $X2=0
+ $Y2=0
cc_427 N_A_126_368#_c_536_n N_VPWR_c_743_n 0.0219924f $X=4.795 $Y=2.325 $X2=0
+ $Y2=0
cc_428 N_A_126_368#_c_537_n N_VPWR_c_743_n 0.0267471f $X=5.015 $Y=2.485 $X2=0
+ $Y2=0
cc_429 N_A_126_368#_c_561_n N_VPWR_c_744_n 0.0171814f $X=5.81 $Y=2.145 $X2=0
+ $Y2=0
cc_430 N_A_126_368#_c_538_n N_VPWR_c_744_n 0.0222705f $X=5.915 $Y=2.485 $X2=0
+ $Y2=0
cc_431 N_A_126_368#_c_563_n N_VPWR_c_744_n 0.038469f $X=5.015 $Y=2.145 $X2=0
+ $Y2=0
cc_432 N_A_126_368#_c_538_n N_VPWR_c_745_n 0.0288238f $X=5.915 $Y=2.485 $X2=0
+ $Y2=0
cc_433 N_A_126_368#_c_537_n N_VPWR_c_749_n 0.00780931f $X=5.015 $Y=2.485 $X2=0
+ $Y2=0
cc_434 N_A_126_368#_c_538_n N_VPWR_c_750_n 0.0124152f $X=5.915 $Y=2.485 $X2=0
+ $Y2=0
cc_435 N_A_126_368#_c_537_n N_VPWR_c_742_n 0.00624184f $X=5.015 $Y=2.485 $X2=0
+ $Y2=0
cc_436 N_A_126_368#_c_538_n N_VPWR_c_742_n 0.00989001f $X=5.915 $Y=2.485 $X2=0
+ $Y2=0
cc_437 N_Y_c_613_n N_VGND_M1008_d 0.00358162f $X=1.615 $Y=1.08 $X2=0 $Y2=0
cc_438 N_Y_c_607_n N_VGND_M1026_d 9.24827e-19 $X=2.625 $Y=1.065 $X2=0 $Y2=0
cc_439 N_Y_c_614_n N_VGND_M1026_d 0.00158118f $X=2.275 $Y=1.08 $X2=0 $Y2=0
cc_440 N_Y_c_609_n N_VGND_M1001_d 0.00250873f $X=3.475 $Y=1.065 $X2=0 $Y2=0
cc_441 N_Y_c_663_n N_VGND_M1013_d 0.00859297f $X=4.475 $Y=0.965 $X2=0 $Y2=0
cc_442 N_Y_c_685_n N_VGND_M1011_s 0.0104519f $X=5.605 $Y=0.965 $X2=0 $Y2=0
cc_443 N_Y_c_604_n N_VGND_c_837_n 0.0256697f $X=0.78 $Y=0.515 $X2=0 $Y2=0
cc_444 N_Y_c_605_n N_VGND_c_837_n 0.00630154f $X=0.945 $Y=1.095 $X2=0 $Y2=0
cc_445 N_Y_c_604_n N_VGND_c_838_n 0.0191765f $X=0.78 $Y=0.515 $X2=0 $Y2=0
cc_446 N_Y_c_606_n N_VGND_c_838_n 0.0191765f $X=1.78 $Y=0.515 $X2=0 $Y2=0
cc_447 N_Y_c_613_n N_VGND_c_838_n 0.0248957f $X=1.615 $Y=1.08 $X2=0 $Y2=0
cc_448 N_Y_c_606_n N_VGND_c_839_n 0.0144124f $X=1.78 $Y=0.515 $X2=0 $Y2=0
cc_449 N_Y_c_606_n N_VGND_c_840_n 0.0180508f $X=1.78 $Y=0.515 $X2=0 $Y2=0
cc_450 N_Y_c_608_n N_VGND_c_840_n 0.0171736f $X=2.71 $Y=0.515 $X2=0 $Y2=0
cc_451 N_Y_c_614_n N_VGND_c_840_n 0.0210834f $X=2.275 $Y=1.08 $X2=0 $Y2=0
cc_452 N_Y_c_608_n N_VGND_c_841_n 0.0171736f $X=2.71 $Y=0.515 $X2=0 $Y2=0
cc_453 N_Y_c_609_n N_VGND_c_841_n 0.0209867f $X=3.475 $Y=1.065 $X2=0 $Y2=0
cc_454 N_Y_c_610_n N_VGND_c_841_n 0.0180508f $X=3.64 $Y=0.515 $X2=0 $Y2=0
cc_455 N_Y_c_610_n N_VGND_c_842_n 0.0142986f $X=3.64 $Y=0.515 $X2=0 $Y2=0
cc_456 N_Y_c_663_n N_VGND_c_842_n 0.0248957f $X=4.475 $Y=0.965 $X2=0 $Y2=0
cc_457 N_Y_c_611_n N_VGND_c_842_n 0.0142986f $X=4.64 $Y=0.515 $X2=0 $Y2=0
cc_458 N_Y_c_611_n N_VGND_c_843_n 0.0145227f $X=4.64 $Y=0.515 $X2=0 $Y2=0
cc_459 N_Y_c_611_n N_VGND_c_844_n 0.0132136f $X=4.64 $Y=0.515 $X2=0 $Y2=0
cc_460 N_Y_c_685_n N_VGND_c_844_n 0.0314257f $X=5.605 $Y=0.965 $X2=0 $Y2=0
cc_461 N_Y_c_612_n N_VGND_c_844_n 0.0132136f $X=5.77 $Y=0.515 $X2=0 $Y2=0
cc_462 N_Y_c_612_n N_VGND_c_845_n 0.0206774f $X=5.77 $Y=0.515 $X2=0 $Y2=0
cc_463 N_Y_c_612_n N_VGND_c_846_n 0.0145947f $X=5.77 $Y=0.515 $X2=0 $Y2=0
cc_464 N_Y_c_604_n N_VGND_c_848_n 0.0145639f $X=0.78 $Y=0.515 $X2=0 $Y2=0
cc_465 N_Y_c_608_n N_VGND_c_849_n 0.00749631f $X=2.71 $Y=0.515 $X2=0 $Y2=0
cc_466 N_Y_c_610_n N_VGND_c_850_n 0.0144922f $X=3.64 $Y=0.515 $X2=0 $Y2=0
cc_467 N_Y_c_604_n N_VGND_c_852_n 0.0119984f $X=0.78 $Y=0.515 $X2=0 $Y2=0
cc_468 N_Y_c_606_n N_VGND_c_852_n 0.0118513f $X=1.78 $Y=0.515 $X2=0 $Y2=0
cc_469 N_Y_c_608_n N_VGND_c_852_n 0.0062048f $X=2.71 $Y=0.515 $X2=0 $Y2=0
cc_470 N_Y_c_610_n N_VGND_c_852_n 0.0118826f $X=3.64 $Y=0.515 $X2=0 $Y2=0
cc_471 N_Y_c_611_n N_VGND_c_852_n 0.0118946f $X=4.64 $Y=0.515 $X2=0 $Y2=0
cc_472 N_Y_c_612_n N_VGND_c_852_n 0.0120104f $X=5.77 $Y=0.515 $X2=0 $Y2=0
