* File: sky130_fd_sc_hs__o21a_4.spice
* Created: Tue Sep  1 20:14:24 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hs__o21a_4.pex.spice"
.subckt sky130_fd_sc_hs__o21a_4  VNB VPB A2 A1 B1 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* B1	B1
* A1	A1
* A2	A2
* VPB	VPB
* VNB	VNB
MM1010 N_VGND_M1010_d N_A1_M1010_g N_A_27_125#_M1010_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.1136 AS=0.1824 PD=0.995 PS=1.85 NRD=13.116 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75002.7 A=0.096 P=1.58 MULT=1
MM1005 N_A_27_125#_M1005_d N_A2_M1005_g N_VGND_M1010_d VNB NLOWVT L=0.15 W=0.64
+ AD=0.0896 AS=0.1136 PD=0.92 PS=0.995 NRD=0 NRS=0.936 M=1 R=4.26667 SA=75000.7
+ SB=75002.2 A=0.096 P=1.58 MULT=1
MM1006 N_A_27_125#_M1005_d N_A2_M1006_g N_VGND_M1006_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.0896 AS=0.1376 PD=0.92 PS=1.07 NRD=0 NRS=14.988 M=1 R=4.26667 SA=75001.1
+ SB=75001.7 A=0.096 P=1.58 MULT=1
MM1012 N_VGND_M1006_s N_A1_M1012_g N_A_27_125#_M1012_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.1376 AS=0.0896 PD=1.07 PS=0.92 NRD=13.116 NRS=0 M=1 R=4.26667 SA=75001.7
+ SB=75001.1 A=0.096 P=1.58 MULT=1
MM1009 N_A_27_125#_M1012_s N_B1_M1009_g N_A_216_387#_M1009_s VNB NLOWVT L=0.15
+ W=0.64 AD=0.0896 AS=0.0896 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75002.2 SB=75000.7 A=0.096 P=1.58 MULT=1
MM1014 N_A_27_125#_M1014_d N_B1_M1014_g N_A_216_387#_M1009_s VNB NLOWVT L=0.15
+ W=0.64 AD=0.2336 AS=0.0896 PD=2.01 PS=0.92 NRD=14.988 NRS=0 M=1 R=4.26667
+ SA=75002.6 SB=75000.3 A=0.096 P=1.58 MULT=1
MM1001 N_VGND_M1001_d N_A_216_387#_M1001_g N_X_M1001_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.1036 PD=2.05 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75001.5 A=0.111 P=1.78 MULT=1
MM1002 N_VGND_M1002_d N_A_216_387#_M1002_g N_X_M1001_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.11655 AS=0.1036 PD=1.055 PS=1.02 NRD=2.424 NRS=0 M=1 R=4.93333 SA=75000.6
+ SB=75001.1 A=0.111 P=1.78 MULT=1
MM1007 N_VGND_M1002_d N_A_216_387#_M1007_g N_X_M1007_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.11655 AS=0.1036 PD=1.055 PS=1.02 NRD=3.24 NRS=0 M=1 R=4.93333 SA=75001.1
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1008 N_VGND_M1008_d N_A_216_387#_M1008_g N_X_M1007_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.1036 PD=2.05 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.5
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1017 N_VPWR_M1017_d N_A1_M1017_g N_A_116_387#_M1017_s VPB PSHORT L=0.15 W=1
+ AD=0.295 AS=0.175 PD=2.59 PS=1.35 NRD=1.9503 NRS=11.8003 M=1 R=6.66667
+ SA=75000.2 SB=75004.4 A=0.15 P=2.3 MULT=1
MM1015 N_A_216_387#_M1015_d N_A2_M1015_g N_A_116_387#_M1017_s VPB PSHORT L=0.15
+ W=1 AD=0.15 AS=0.175 PD=1.3 PS=1.35 NRD=1.9503 NRS=1.9503 M=1 R=6.66667
+ SA=75000.7 SB=75003.9 A=0.15 P=2.3 MULT=1
MM1018 N_A_216_387#_M1015_d N_A2_M1018_g N_A_116_387#_M1018_s VPB PSHORT L=0.15
+ W=1 AD=0.15 AS=0.175 PD=1.3 PS=1.35 NRD=1.9503 NRS=11.8003 M=1 R=6.66667
+ SA=75001.2 SB=75003.5 A=0.15 P=2.3 MULT=1
MM1019 N_VPWR_M1019_d N_A1_M1019_g N_A_116_387#_M1018_s VPB PSHORT L=0.15 W=1
+ AD=0.201087 AS=0.175 PD=1.51087 PS=1.35 NRD=11.8003 NRS=1.9503 M=1 R=6.66667
+ SA=75001.7 SB=75003 A=0.15 P=2.3 MULT=1
MM1003 N_VPWR_M1019_d N_B1_M1003_g N_A_216_387#_M1003_s VPB PSHORT L=0.15 W=0.84
+ AD=0.168913 AS=0.1596 PD=1.26913 PS=1.22 NRD=11.7215 NRS=4.6886 M=1 R=5.6
+ SA=75002.2 SB=75003 A=0.126 P=1.98 MULT=1
MM1004 N_VPWR_M1004_d N_B1_M1004_g N_A_216_387#_M1003_s VPB PSHORT L=0.15 W=0.84
+ AD=0.2406 AS=0.1596 PD=1.45714 PS=1.22 NRD=28.1316 NRS=18.7544 M=1 R=5.6
+ SA=75002.7 SB=75002.4 A=0.126 P=1.98 MULT=1
MM1000 N_VPWR_M1004_d N_A_216_387#_M1000_g N_X_M1000_s VPB PSHORT L=0.15 W=1.12
+ AD=0.3208 AS=0.168 PD=1.94286 PS=1.42 NRD=31.6579 NRS=1.7533 M=1 R=7.46667
+ SA=75002.6 SB=75001.7 A=0.168 P=2.54 MULT=1
MM1011 N_VPWR_M1011_d N_A_216_387#_M1011_g N_X_M1000_s VPB PSHORT L=0.15 W=1.12
+ AD=0.224 AS=0.168 PD=1.52 PS=1.42 NRD=10.5395 NRS=1.7533 M=1 R=7.46667
+ SA=75003.1 SB=75001.3 A=0.168 P=2.54 MULT=1
MM1013 N_VPWR_M1011_d N_A_216_387#_M1013_g N_X_M1013_s VPB PSHORT L=0.15 W=1.12
+ AD=0.224 AS=0.168 PD=1.52 PS=1.42 NRD=10.5395 NRS=1.7533 M=1 R=7.46667
+ SA=75003.6 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1016 N_VPWR_M1016_d N_A_216_387#_M1016_g N_X_M1013_s VPB PSHORT L=0.15 W=1.12
+ AD=0.3864 AS=0.168 PD=2.93 PS=1.42 NRD=10.5395 NRS=1.7533 M=1 R=7.46667
+ SA=75004.1 SB=75000.3 A=0.168 P=2.54 MULT=1
DX20_noxref VNB VPB NWDIODE A=11.4204 P=16
*
.include "sky130_fd_sc_hs__o21a_4.pxi.spice"
*
.ends
*
*
