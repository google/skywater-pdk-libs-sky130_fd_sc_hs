* File: sky130_fd_sc_hs__mux2_1.pex.spice
* Created: Thu Aug 27 20:48:45 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HS__MUX2_1%S 3 5 7 8 10 13 16 17 18 19 23
c57 16 0 7.03863e-20 $X=0.505 $Y=1.557
c58 13 0 1.07726e-19 $X=1.055 $Y=0.74
r59 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.67
+ $Y=1.515 $X2=0.67 $Y2=1.515
r60 19 23 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=0.67 $Y=1.665
+ $X2=0.67 $Y2=1.515
r61 17 22 48.9612 $w=3.3e-07 $l=2.8e-07 $layer=POLY_cond $X=0.95 $Y=1.515
+ $X2=0.67 $Y2=1.515
r62 17 18 5.03009 $w=3.3e-07 $l=1.08995e-07 $layer=POLY_cond $X=0.95 $Y=1.515
+ $X2=1.04 $Y2=1.557
r63 15 22 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=0.595 $Y=1.515
+ $X2=0.67 $Y2=1.515
r64 15 16 5.03009 $w=3.3e-07 $l=1.08995e-07 $layer=POLY_cond $X=0.595 $Y=1.515
+ $X2=0.505 $Y2=1.557
r65 11 18 37.0704 $w=1.5e-07 $l=2.14369e-07 $layer=POLY_cond $X=1.055 $Y=1.35
+ $X2=1.04 $Y2=1.557
r66 11 13 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.055 $Y=1.35
+ $X2=1.055 $Y2=0.74
r67 8 18 37.0704 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=1.04 $Y=1.765
+ $X2=1.04 $Y2=1.557
r68 8 10 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=1.04 $Y=1.765
+ $X2=1.04 $Y2=2.34
r69 5 16 37.0704 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=0.505 $Y=1.765
+ $X2=0.505 $Y2=1.557
r70 5 7 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=0.505 $Y=1.765
+ $X2=0.505 $Y2=2.26
r71 1 16 37.0704 $w=1.5e-07 $l=2.11941e-07 $layer=POLY_cond $X=0.495 $Y=1.35
+ $X2=0.505 $Y2=1.557
r72 1 3 264.074 $w=1.5e-07 $l=5.15e-07 $layer=POLY_cond $X=0.495 $Y=1.35
+ $X2=0.495 $Y2=0.835
.ends

.subckt PM_SKY130_FD_SC_HS__MUX2_1%A1 3 4 6 8 9 10 13 15 17 18 23 28
c62 23 0 1.32486e-19 $X=1.51 $Y=1.22
c63 10 0 1.07726e-19 $X=1.685 $Y=0.895
r64 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.62
+ $Y=1.385 $X2=2.62 $Y2=1.385
r65 18 27 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=2.62 $Y=1.295 $X2=2.62
+ $Y2=1.385
r66 17 28 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.62 $Y=0.895 $X2=2.62
+ $Y2=0.98
r67 17 18 10.4768 $w=3.28e-07 $l=3e-07 $layer=LI1_cond $X=2.62 $Y=0.995 $X2=2.62
+ $Y2=1.295
r68 17 28 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=2.62 $Y=0.995
+ $X2=2.62 $Y2=0.98
r69 13 23 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.51 $Y=1.385
+ $X2=1.51 $Y2=1.22
r70 12 15 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=1.51 $Y=1.385 $X2=1.6
+ $Y2=1.385
r71 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.51
+ $Y=1.385 $X2=1.51 $Y2=1.385
r72 9 17 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.455 $Y=0.895
+ $X2=2.62 $Y2=0.895
r73 9 10 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=2.455 $Y=0.895
+ $X2=1.685 $Y2=0.895
r74 8 15 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.6 $Y=1.22 $X2=1.6
+ $Y2=1.385
r75 7 10 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.6 $Y=0.98
+ $X2=1.685 $Y2=0.895
r76 7 8 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=1.6 $Y=0.98 $X2=1.6
+ $Y2=1.22
r77 4 26 77.2841 $w=2.7e-07 $l=4.15812e-07 $layer=POLY_cond $X=2.545 $Y=1.765
+ $X2=2.62 $Y2=1.385
r78 4 6 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=2.545 $Y=1.765
+ $X2=2.545 $Y2=2.34
r79 3 23 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.445 $Y=0.74
+ $X2=1.445 $Y2=1.22
.ends

.subckt PM_SKY130_FD_SC_HS__MUX2_1%A0 1 3 4 6 7
c29 7 0 1.1756e-19 $X=2.16 $Y=1.295
r30 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.05
+ $Y=1.385 $X2=2.05 $Y2=1.385
r31 7 11 3.42618 $w=3.68e-07 $l=1.1e-07 $layer=LI1_cond $X=2.16 $Y=1.365
+ $X2=2.05 $Y2=1.365
r32 4 10 38.9026 $w=2.7e-07 $l=2.05122e-07 $layer=POLY_cond $X=2.14 $Y=1.22
+ $X2=2.05 $Y2=1.385
r33 4 6 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=2.14 $Y=1.22 $X2=2.14
+ $Y2=0.74
r34 1 10 77.2841 $w=2.7e-07 $l=4.01871e-07 $layer=POLY_cond $X=2.005 $Y=1.765
+ $X2=2.05 $Y2=1.385
r35 1 3 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=2.005 $Y=1.765
+ $X2=2.005 $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_HS__MUX2_1%A_27_112# 1 2 9 11 13 16 19 22 25 26 27 29 30
+ 32 36
c90 9 0 8.6251e-20 $X=3.1 $Y=0.74
r91 36 37 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.19
+ $Y=1.485 $X2=3.19 $Y2=1.485
r92 33 36 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=3.04 $Y=1.485
+ $X2=3.19 $Y2=1.485
r93 28 33 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.04 $Y=1.65
+ $X2=3.04 $Y2=1.485
r94 28 29 81.877 $w=1.68e-07 $l=1.255e-06 $layer=LI1_cond $X=3.04 $Y=1.65
+ $X2=3.04 $Y2=2.905
r95 26 29 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.955 $Y=2.99
+ $X2=3.04 $Y2=2.905
r96 26 27 106.668 $w=1.68e-07 $l=1.635e-06 $layer=LI1_cond $X=2.955 $Y=2.99
+ $X2=1.32 $Y2=2.99
r97 25 27 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.235 $Y=2.905
+ $X2=1.32 $Y2=2.99
r98 24 25 44.0374 $w=1.68e-07 $l=6.75e-07 $layer=LI1_cond $X=1.235 $Y=2.23
+ $X2=1.235 $Y2=2.905
r99 23 32 2.76166 $w=1.7e-07 $l=1.90526e-07 $layer=LI1_cond $X=0.445 $Y=2.145
+ $X2=0.28 $Y2=2.09
r100 22 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.15 $Y=2.145
+ $X2=1.235 $Y2=2.23
r101 22 23 45.9947 $w=1.68e-07 $l=7.05e-07 $layer=LI1_cond $X=1.15 $Y=2.145
+ $X2=0.445 $Y2=2.145
r102 19 32 3.70735 $w=2.5e-07 $l=1.75499e-07 $layer=LI1_cond $X=0.2 $Y=1.95
+ $X2=0.28 $Y2=2.09
r103 19 30 53.4973 $w=1.68e-07 $l=8.2e-07 $layer=LI1_cond $X=0.2 $Y=1.95 $X2=0.2
+ $Y2=1.13
r104 14 30 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=0.28 $Y=0.965
+ $X2=0.28 $Y2=1.13
r105 14 16 4.53993 $w=3.28e-07 $l=1.3e-07 $layer=LI1_cond $X=0.28 $Y=0.965
+ $X2=0.28 $Y2=0.835
r106 11 37 57.6553 $w=2.91e-07 $l=3.15278e-07 $layer=POLY_cond $X=3.115 $Y=1.765
+ $X2=3.19 $Y2=1.485
r107 11 13 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=3.115 $Y=1.765
+ $X2=3.115 $Y2=2.34
r108 7 37 38.6072 $w=2.91e-07 $l=2.05122e-07 $layer=POLY_cond $X=3.1 $Y=1.32
+ $X2=3.19 $Y2=1.485
r109 7 9 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=3.1 $Y=1.32 $X2=3.1
+ $Y2=0.74
r110 2 32 300 $w=1.7e-07 $l=2.83373e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.06
r111 1 16 182 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.56 $X2=0.28 $Y2=0.835
.ends

.subckt PM_SKY130_FD_SC_HS__MUX2_1%A_304_74# 1 2 7 9 12 15 17 18 19 20 21 26 29
+ 30 31 33 36 41
c102 19 0 3.72132e-20 $X=1.175 $Y=1.805
c103 15 0 3.31731e-20 $X=1.09 $Y=1.72
c104 7 0 1.16478e-19 $X=3.735 $Y=1.765
r105 41 42 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.73
+ $Y=1.465 $X2=3.73 $Y2=1.465
r106 38 41 4.1907 $w=3.28e-07 $l=1.2e-07 $layer=LI1_cond $X=3.61 $Y=1.465
+ $X2=3.73 $Y2=1.465
r107 34 36 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=1.09 $Y=0.935
+ $X2=1.26 $Y2=0.935
r108 33 38 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.61 $Y=1.3
+ $X2=3.61 $Y2=1.465
r109 32 33 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=3.61 $Y=1.15
+ $X2=3.61 $Y2=1.3
r110 30 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.525 $Y=1.065
+ $X2=3.61 $Y2=1.15
r111 30 31 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=3.525 $Y=1.065
+ $X2=3.125 $Y2=1.065
r112 29 31 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.04 $Y=0.98
+ $X2=3.125 $Y2=1.065
r113 28 29 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=3.04 $Y=0.64
+ $X2=3.04 $Y2=0.98
r114 24 26 3.31764 $w=3.28e-07 $l=9.5e-08 $layer=LI1_cond $X=2.23 $Y=1.89
+ $X2=2.23 $Y2=1.985
r115 21 23 20.5135 $w=2.48e-07 $l=4.45e-07 $layer=LI1_cond $X=1.345 $Y=0.515
+ $X2=1.79 $Y2=0.515
r116 20 28 7.14316 $w=2.5e-07 $l=1.62019e-07 $layer=LI1_cond $X=2.955 $Y=0.515
+ $X2=3.04 $Y2=0.64
r117 20 23 53.7038 $w=2.48e-07 $l=1.165e-06 $layer=LI1_cond $X=2.955 $Y=0.515
+ $X2=1.79 $Y2=0.515
r118 18 24 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.065 $Y=1.805
+ $X2=2.23 $Y2=1.89
r119 18 19 58.0642 $w=1.68e-07 $l=8.9e-07 $layer=LI1_cond $X=2.065 $Y=1.805
+ $X2=1.175 $Y2=1.805
r120 17 36 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.26 $Y=0.85
+ $X2=1.26 $Y2=0.935
r121 16 21 7.14316 $w=2.5e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.26 $Y=0.64
+ $X2=1.345 $Y2=0.515
r122 16 17 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=1.26 $Y=0.64
+ $X2=1.26 $Y2=0.85
r123 15 19 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.09 $Y=1.72
+ $X2=1.175 $Y2=1.805
r124 14 34 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.09 $Y=1.02
+ $X2=1.09 $Y2=0.935
r125 14 15 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=1.09 $Y=1.02 $X2=1.09
+ $Y2=1.72
r126 10 42 38.6549 $w=2.86e-07 $l=2.03101e-07 $layer=POLY_cond $X=3.815 $Y=1.3
+ $X2=3.73 $Y2=1.465
r127 10 12 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=3.815 $Y=1.3
+ $X2=3.815 $Y2=0.74
r128 7 42 61.4066 $w=2.86e-07 $l=3.0249e-07 $layer=POLY_cond $X=3.735 $Y=1.765
+ $X2=3.73 $Y2=1.465
r129 7 9 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.735 $Y=1.765
+ $X2=3.735 $Y2=2.4
r130 2 26 300 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=2 $X=2.08
+ $Y=1.84 $X2=2.23 $Y2=1.985
r131 1 23 182 $w=1.7e-07 $l=3.505e-07 $layer=licon1_NDIFF $count=1 $X=1.52
+ $Y=0.37 $X2=1.79 $Y2=0.555
.ends

.subckt PM_SKY130_FD_SC_HS__MUX2_1%VPWR 1 2 11 15 20 21 22 32 33 36
r41 36 37 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r42 32 33 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r43 30 33 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=4.08 $Y2=3.33
r44 29 30 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r45 27 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r46 26 29 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=1.2 $Y=3.33
+ $X2=3.12 $Y2=3.33
r47 26 27 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r48 24 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.98 $Y=3.33
+ $X2=0.815 $Y2=3.33
r49 24 26 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=0.98 $Y=3.33 $X2=1.2
+ $Y2=3.33
r50 22 30 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=3.12 $Y2=3.33
r51 22 27 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.2 $Y2=3.33
r52 20 29 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=3.295 $Y=3.33
+ $X2=3.12 $Y2=3.33
r53 20 21 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.295 $Y=3.33
+ $X2=3.46 $Y2=3.33
r54 19 32 29.6845 $w=1.68e-07 $l=4.55e-07 $layer=LI1_cond $X=3.625 $Y=3.33
+ $X2=4.08 $Y2=3.33
r55 19 21 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.625 $Y=3.33
+ $X2=3.46 $Y2=3.33
r56 15 18 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=3.46 $Y=1.985
+ $X2=3.46 $Y2=2.815
r57 13 21 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.46 $Y=3.245
+ $X2=3.46 $Y2=3.33
r58 13 18 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=3.46 $Y=3.245
+ $X2=3.46 $Y2=2.815
r59 9 36 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.815 $Y=3.245
+ $X2=0.815 $Y2=3.33
r60 9 11 25.668 $w=3.28e-07 $l=7.35e-07 $layer=LI1_cond $X=0.815 $Y=3.245
+ $X2=0.815 $Y2=2.51
r61 2 18 600 $w=1.7e-07 $l=1.10176e-06 $layer=licon1_PDIFF $count=1 $X=3.19
+ $Y=1.84 $X2=3.46 $Y2=2.815
r62 2 15 300 $w=1.7e-07 $l=3.34739e-07 $layer=licon1_PDIFF $count=2 $X=3.19
+ $Y=1.84 $X2=3.46 $Y2=1.985
r63 1 11 600 $w=1.7e-07 $l=7.78685e-07 $layer=licon1_PDIFF $count=1 $X=0.58
+ $Y=1.84 $X2=0.815 $Y2=2.51
.ends

.subckt PM_SKY130_FD_SC_HS__MUX2_1%X 1 2 9 13 14 15 16 31 32 35
c24 13 0 2.02729e-19 $X=4.05 $Y=1.13
r25 31 32 8.83531 $w=4.38e-07 $l=1.65e-07 $layer=LI1_cond $X=4.015 $Y=1.985
+ $X2=4.015 $Y2=1.82
r26 21 35 0.130959 $w=4.38e-07 $l=5e-09 $layer=LI1_cond $X=4.015 $Y=2.04
+ $X2=4.015 $Y2=2.035
r27 16 28 1.04768 $w=4.38e-07 $l=4e-08 $layer=LI1_cond $X=4.015 $Y=2.775
+ $X2=4.015 $Y2=2.815
r28 15 16 9.691 $w=4.38e-07 $l=3.7e-07 $layer=LI1_cond $X=4.015 $Y=2.405
+ $X2=4.015 $Y2=2.775
r29 14 35 1.04768 $w=4.38e-07 $l=4e-08 $layer=LI1_cond $X=4.015 $Y=1.995
+ $X2=4.015 $Y2=2.035
r30 14 31 0.261919 $w=4.38e-07 $l=1e-08 $layer=LI1_cond $X=4.015 $Y=1.995
+ $X2=4.015 $Y2=1.985
r31 14 15 8.51236 $w=4.38e-07 $l=3.25e-07 $layer=LI1_cond $X=4.015 $Y=2.08
+ $X2=4.015 $Y2=2.405
r32 14 21 1.04768 $w=4.38e-07 $l=4e-08 $layer=LI1_cond $X=4.015 $Y=2.08
+ $X2=4.015 $Y2=2.04
r33 13 32 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=4.15 $Y=1.13 $X2=4.15
+ $Y2=1.82
r34 7 13 9.16175 $w=3.68e-07 $l=1.85e-07 $layer=LI1_cond $X=4.05 $Y=0.945
+ $X2=4.05 $Y2=1.13
r35 7 9 13.3933 $w=3.68e-07 $l=4.3e-07 $layer=LI1_cond $X=4.05 $Y=0.945 $X2=4.05
+ $Y2=0.515
r36 2 31 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=3.81
+ $Y=1.84 $X2=3.96 $Y2=1.985
r37 2 28 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=3.81
+ $Y=1.84 $X2=3.96 $Y2=2.815
r38 1 9 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.89
+ $Y=0.37 $X2=4.03 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__MUX2_1%VGND 1 2 8 11 15 18 21 22 23 25 38 39 42
c51 18 0 1.49261e-20 $X=0.815 $Y=0.515
r52 42 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r53 38 39 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r54 36 39 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=4.08
+ $Y2=0
r55 35 36 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r56 33 43 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r57 32 35 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=1.2 $Y=0 $X2=3.12
+ $Y2=0
r58 32 33 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r59 30 42 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.005 $Y=0 $X2=0.815
+ $Y2=0
r60 30 32 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=1.005 $Y=0 $X2=1.2
+ $Y2=0
r61 28 43 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r62 27 28 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r63 25 42 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.625 $Y=0 $X2=0.815
+ $Y2=0
r64 25 27 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=0.625 $Y=0 $X2=0.24
+ $Y2=0
r65 23 36 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=3.12
+ $Y2=0
r66 23 33 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.2
+ $Y2=0
r67 21 35 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=3.295 $Y=0 $X2=3.12
+ $Y2=0
r68 21 22 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.295 $Y=0 $X2=3.46
+ $Y2=0
r69 20 38 29.6845 $w=1.68e-07 $l=4.55e-07 $layer=LI1_cond $X=3.625 $Y=0 $X2=4.08
+ $Y2=0
r70 20 22 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.625 $Y=0 $X2=3.46
+ $Y2=0
r71 18 19 7.29301 $w=3.78e-07 $l=1.65e-07 $layer=LI1_cond $X=0.815 $Y=0.515
+ $X2=0.815 $Y2=0.68
r72 13 22 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.46 $Y=0.085
+ $X2=3.46 $Y2=0
r73 13 15 19.5566 $w=3.28e-07 $l=5.6e-07 $layer=LI1_cond $X=3.46 $Y=0.085
+ $X2=3.46 $Y2=0.645
r74 11 19 15.0519 $w=2.08e-07 $l=2.85e-07 $layer=LI1_cond $X=0.73 $Y=0.965
+ $X2=0.73 $Y2=0.68
r75 8 18 0.758186 $w=3.78e-07 $l=2.5e-08 $layer=LI1_cond $X=0.815 $Y=0.49
+ $X2=0.815 $Y2=0.515
r76 7 42 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=0.815 $Y=0.085
+ $X2=0.815 $Y2=0
r77 7 8 12.2826 $w=3.78e-07 $l=4.05e-07 $layer=LI1_cond $X=0.815 $Y=0.085
+ $X2=0.815 $Y2=0.49
r78 2 15 182 $w=1.7e-07 $l=3.995e-07 $layer=licon1_NDIFF $count=1 $X=3.175
+ $Y=0.37 $X2=3.46 $Y2=0.645
r79 1 18 182 $w=1.7e-07 $l=2.66552e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.56 $X2=0.815 $Y2=0.515
r80 1 11 182 $w=1.7e-07 $l=4.76235e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.56 $X2=0.725 $Y2=0.965
.ends

