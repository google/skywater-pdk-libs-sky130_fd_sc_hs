* File: sky130_fd_sc_hs__clkdlyinv3sd2_1.pex.spice
* Created: Tue Sep  1 19:58:05 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HS__CLKDLYINV3SD2_1%A 3 6 7 9 10 11 15
r37 15 18 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.57 $Y=1.355
+ $X2=0.57 $Y2=1.52
r38 15 17 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.57 $Y=1.355
+ $X2=0.57 $Y2=1.19
r39 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.57
+ $Y=1.355 $X2=0.57 $Y2=1.355
r40 11 16 5.88547 $w=6.28e-07 $l=3.1e-07 $layer=LI1_cond $X=0.415 $Y=1.665
+ $X2=0.415 $Y2=1.355
r41 10 16 1.13912 $w=6.28e-07 $l=6e-08 $layer=LI1_cond $X=0.415 $Y=1.295
+ $X2=0.415 $Y2=1.355
r42 7 9 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.495 $Y=1.765
+ $X2=0.495 $Y2=2.4
r43 6 7 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=0.495 $Y=1.675 $X2=0.495
+ $Y2=1.765
r44 6 18 60.25 $w=1.8e-07 $l=1.55e-07 $layer=POLY_cond $X=0.495 $Y=1.675
+ $X2=0.495 $Y2=1.52
r45 3 17 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=0.48 $Y=0.58 $X2=0.48
+ $Y2=1.19
.ends

.subckt PM_SKY130_FD_SC_HS__CLKDLYINV3SD2_1%A_28_74# 1 2 9 13 17 19 21 23 25 26
+ 30 31
r62 31 36 59.3793 $w=5e-07 $l=4.3e-07 $layer=POLY_cond $X=1.195 $Y=1.295
+ $X2=1.195 $Y2=1.725
r63 31 35 40.7881 $w=5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.195 $Y=1.295
+ $X2=1.195 $Y2=1.13
r64 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.14
+ $Y=1.295 $X2=1.14 $Y2=1.295
r65 28 30 25.668 $w=3.28e-07 $l=7.35e-07 $layer=LI1_cond $X=1.14 $Y=2.03
+ $X2=1.14 $Y2=1.295
r66 27 30 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=1.14 $Y=1.02
+ $X2=1.14 $Y2=1.295
r67 25 27 7.36389 $w=2e-07 $l=2.09105e-07 $layer=LI1_cond $X=0.975 $Y=0.92
+ $X2=1.14 $Y2=1.02
r68 25 26 31.3318 $w=1.98e-07 $l=5.65e-07 $layer=LI1_cond $X=0.975 $Y=0.92
+ $X2=0.41 $Y2=0.92
r69 24 33 4.75367 $w=1.75e-07 $l=1.53e-07 $layer=LI1_cond $X=0.4 $Y=2.117
+ $X2=0.247 $Y2=2.117
r70 23 28 7.68689 $w=1.75e-07 $l=2.03912e-07 $layer=LI1_cond $X=0.975 $Y=2.117
+ $X2=1.14 $Y2=2.03
r71 23 24 36.4416 $w=1.73e-07 $l=5.75e-07 $layer=LI1_cond $X=0.975 $Y=2.117
+ $X2=0.4 $Y2=2.117
r72 19 33 2.73414 $w=3.05e-07 $l=8.8e-08 $layer=LI1_cond $X=0.247 $Y=2.205
+ $X2=0.247 $Y2=2.117
r73 19 21 13.4137 $w=3.03e-07 $l=3.55e-07 $layer=LI1_cond $X=0.247 $Y=2.205
+ $X2=0.247 $Y2=2.56
r74 15 26 7.26812 $w=2e-07 $l=2.01901e-07 $layer=LI1_cond $X=0.252 $Y=0.82
+ $X2=0.41 $Y2=0.92
r75 15 17 8.78052 $w=3.13e-07 $l=2.4e-07 $layer=LI1_cond $X=0.252 $Y=0.82
+ $X2=0.252 $Y2=0.58
r76 13 35 213.79 $w=1.8e-07 $l=5.5e-07 $layer=POLY_cond $X=1.35 $Y=0.58 $X2=1.35
+ $Y2=1.13
r77 9 36 182.613 $w=2.5e-07 $l=7.35e-07 $layer=POLY_cond $X=1.32 $Y=2.46
+ $X2=1.32 $Y2=1.725
r78 2 33 600 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_PDIFF $count=1 $X=0.14
+ $Y=1.84 $X2=0.265 $Y2=2.115
r79 2 21 600 $w=1.7e-07 $l=7.8e-07 $layer=licon1_PDIFF $count=1 $X=0.14 $Y=1.84
+ $X2=0.265 $Y2=2.56
r80 1 17 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.14
+ $Y=0.37 $X2=0.265 $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_HS__CLKDLYINV3SD2_1%A_288_74# 1 2 9 11 13 16 21 24 28 31
r41 28 29 6.17723 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=1.58 $Y=2.815
+ $X2=1.58 $Y2=2.65
r42 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.275
+ $Y=1.46 $X2=2.275 $Y2=1.46
r43 22 31 0.466467 $w=3.3e-07 $l=1.35e-07 $layer=LI1_cond $X=1.745 $Y=1.46
+ $X2=1.61 $Y2=1.46
r44 22 24 18.5089 $w=3.28e-07 $l=5.3e-07 $layer=LI1_cond $X=1.745 $Y=1.46
+ $X2=2.275 $Y2=1.46
r45 21 29 23.2623 $w=2.68e-07 $l=5.45e-07 $layer=LI1_cond $X=1.61 $Y=2.105
+ $X2=1.61 $Y2=2.65
r46 18 31 6.31733 $w=2.57e-07 $l=1.65e-07 $layer=LI1_cond $X=1.61 $Y=1.625
+ $X2=1.61 $Y2=1.46
r47 18 21 20.4879 $w=2.68e-07 $l=4.8e-07 $layer=LI1_cond $X=1.61 $Y=1.625
+ $X2=1.61 $Y2=2.105
r48 14 31 6.31733 $w=2.57e-07 $l=1.71377e-07 $layer=LI1_cond $X=1.597 $Y=1.295
+ $X2=1.61 $Y2=1.46
r49 14 16 33.6325 $w=2.43e-07 $l=7.15e-07 $layer=LI1_cond $X=1.597 $Y=1.295
+ $X2=1.597 $Y2=0.58
r50 11 25 62.3432 $w=2.85e-07 $l=3.29052e-07 $layer=POLY_cond $X=2.325 $Y=1.765
+ $X2=2.275 $Y2=1.46
r51 11 13 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.325 $Y=1.765
+ $X2=2.325 $Y2=2.4
r52 7 25 38.666 $w=2.85e-07 $l=1.83916e-07 $layer=POLY_cond $X=2.315 $Y=1.295
+ $X2=2.275 $Y2=1.46
r53 7 9 366.628 $w=1.5e-07 $l=7.15e-07 $layer=POLY_cond $X=2.315 $Y=1.295
+ $X2=2.315 $Y2=0.58
r54 2 28 600 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=1.445
+ $Y=1.96 $X2=1.58 $Y2=2.815
r55 2 21 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=1.445
+ $Y=1.96 $X2=1.58 $Y2=2.105
r56 1 16 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.44
+ $Y=0.37 $X2=1.58 $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_HS__CLKDLYINV3SD2_1%VPWR 1 2 9 13 17 19 24 31 32 35 38
+ 46
r33 39 46 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.92 $Y2=3.33
r34 38 39 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r35 35 36 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r36 32 39 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=2.16 $Y2=3.33
r37 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r38 29 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.265 $Y=3.33
+ $X2=2.1 $Y2=3.33
r39 29 31 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=2.265 $Y=3.33
+ $X2=2.64 $Y2=3.33
r40 28 46 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.92 $Y2=3.33
r41 27 28 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r42 25 35 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.905 $Y=3.33
+ $X2=0.74 $Y2=3.33
r43 25 27 50.5615 $w=1.68e-07 $l=7.75e-07 $layer=LI1_cond $X=0.905 $Y=3.33
+ $X2=1.68 $Y2=3.33
r44 24 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.935 $Y=3.33
+ $X2=2.1 $Y2=3.33
r45 24 27 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=1.935 $Y=3.33
+ $X2=1.68 $Y2=3.33
r46 22 36 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r47 21 22 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r48 19 35 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.575 $Y=3.33
+ $X2=0.74 $Y2=3.33
r49 19 21 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=0.575 $Y=3.33
+ $X2=0.24 $Y2=3.33
r50 17 28 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.44 $Y=3.33
+ $X2=1.68 $Y2=3.33
r51 17 36 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.44 $Y=3.33
+ $X2=0.72 $Y2=3.33
r52 13 16 28.8111 $w=3.28e-07 $l=8.25e-07 $layer=LI1_cond $X=2.1 $Y=1.985
+ $X2=2.1 $Y2=2.81
r53 11 38 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.1 $Y=3.245 $X2=2.1
+ $Y2=3.33
r54 11 16 15.1913 $w=3.28e-07 $l=4.35e-07 $layer=LI1_cond $X=2.1 $Y=3.245
+ $X2=2.1 $Y2=2.81
r55 7 35 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.74 $Y=3.245 $X2=0.74
+ $Y2=3.33
r56 7 9 27.2396 $w=3.28e-07 $l=7.8e-07 $layer=LI1_cond $X=0.74 $Y=3.245 $X2=0.74
+ $Y2=2.465
r57 2 16 400 $w=1.7e-07 $l=1.03061e-06 $layer=licon1_PDIFF $count=1 $X=1.975
+ $Y=1.84 $X2=2.1 $Y2=2.81
r58 2 13 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=1.975
+ $Y=1.84 $X2=2.1 $Y2=1.985
r59 1 9 300 $w=1.7e-07 $l=7.04894e-07 $layer=licon1_PDIFF $count=2 $X=0.57
+ $Y=1.84 $X2=0.74 $Y2=2.465
.ends

.subckt PM_SKY130_FD_SC_HS__CLKDLYINV3SD2_1%Y 1 2 7 8 9 10 11 12 13 32
r16 44 45 6.10729 $w=3.58e-07 $l=1.65e-07 $layer=LI1_cond $X=2.615 $Y=0.59
+ $X2=2.615 $Y2=0.755
r17 30 32 1.28049 $w=3.58e-07 $l=4e-08 $layer=LI1_cond $X=2.615 $Y=1.995
+ $X2=2.615 $Y2=2.035
r18 13 47 6.52326 $w=2.63e-07 $l=1.5e-07 $layer=LI1_cond $X=2.662 $Y=1.665
+ $X2=2.662 $Y2=1.815
r19 11 12 11.8446 $w=3.58e-07 $l=3.7e-07 $layer=LI1_cond $X=2.615 $Y=2.405
+ $X2=2.615 $Y2=2.775
r20 10 30 0.736283 $w=3.58e-07 $l=2.3e-08 $layer=LI1_cond $X=2.615 $Y=1.972
+ $X2=2.615 $Y2=1.995
r21 10 47 5.85119 $w=3.58e-07 $l=1.57e-07 $layer=LI1_cond $X=2.615 $Y=1.972
+ $X2=2.615 $Y2=1.815
r22 10 11 11.1403 $w=3.58e-07 $l=3.48e-07 $layer=LI1_cond $X=2.615 $Y=2.057
+ $X2=2.615 $Y2=2.405
r23 10 32 0.704271 $w=3.58e-07 $l=2.2e-08 $layer=LI1_cond $X=2.615 $Y=2.057
+ $X2=2.615 $Y2=2.035
r24 9 13 16.0907 $w=2.63e-07 $l=3.7e-07 $layer=LI1_cond $X=2.662 $Y=1.295
+ $X2=2.662 $Y2=1.665
r25 8 9 16.0907 $w=2.63e-07 $l=3.7e-07 $layer=LI1_cond $X=2.662 $Y=0.925
+ $X2=2.662 $Y2=1.295
r26 8 45 7.39303 $w=2.63e-07 $l=1.7e-07 $layer=LI1_cond $X=2.662 $Y=0.925
+ $X2=2.662 $Y2=0.755
r27 7 44 1.12043 $w=3.58e-07 $l=3.5e-08 $layer=LI1_cond $X=2.615 $Y=0.555
+ $X2=2.615 $Y2=0.59
r28 2 10 400 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_PDIFF $count=1 $X=2.4
+ $Y=1.84 $X2=2.555 $Y2=1.985
r29 2 12 400 $w=1.7e-07 $l=1.04463e-06 $layer=licon1_PDIFF $count=1 $X=2.4
+ $Y=1.84 $X2=2.555 $Y2=2.81
r30 1 44 182 $w=1.7e-07 $l=2.81425e-07 $layer=licon1_NDIFF $count=1 $X=2.39
+ $Y=0.37 $X2=2.53 $Y2=0.59
.ends

.subckt PM_SKY130_FD_SC_HS__CLKDLYINV3SD2_1%VGND 1 2 9 13 15 17 22 29 30 33 36
+ 44
r32 37 44 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.92
+ $Y2=0
r33 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r34 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r35 30 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=2.16
+ $Y2=0
r36 29 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r37 27 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.265 $Y=0 $X2=2.1
+ $Y2=0
r38 27 29 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=2.265 $Y=0 $X2=2.64
+ $Y2=0
r39 26 44 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.92
+ $Y2=0
r40 25 26 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r41 23 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.915 $Y=0 $X2=0.75
+ $Y2=0
r42 23 25 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=0.915 $Y=0 $X2=1.68
+ $Y2=0
r43 22 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.935 $Y=0 $X2=2.1
+ $Y2=0
r44 22 25 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=1.935 $Y=0 $X2=1.68
+ $Y2=0
r45 20 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r46 19 20 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r47 17 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.585 $Y=0 $X2=0.75
+ $Y2=0
r48 17 19 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.585 $Y=0 $X2=0.24
+ $Y2=0
r49 15 26 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.44 $Y=0 $X2=1.68
+ $Y2=0
r50 15 34 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.44 $Y=0 $X2=0.72
+ $Y2=0
r51 11 36 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.1 $Y=0.085 $X2=2.1
+ $Y2=0
r52 11 13 17.4613 $w=3.28e-07 $l=5e-07 $layer=LI1_cond $X=2.1 $Y=0.085 $X2=2.1
+ $Y2=0.585
r53 7 33 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.75 $Y=0.085 $X2=0.75
+ $Y2=0
r54 7 9 16.7628 $w=3.28e-07 $l=4.8e-07 $layer=LI1_cond $X=0.75 $Y=0.085 $X2=0.75
+ $Y2=0.565
r55 2 13 182 $w=1.7e-07 $l=2.7037e-07 $layer=licon1_NDIFF $count=1 $X=1.975
+ $Y=0.37 $X2=2.1 $Y2=0.585
r56 1 9 182 $w=1.7e-07 $l=2.75772e-07 $layer=licon1_NDIFF $count=1 $X=0.555
+ $Y=0.37 $X2=0.75 $Y2=0.565
.ends

