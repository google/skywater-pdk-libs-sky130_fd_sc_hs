* File: sky130_fd_sc_hs__o41a_2.spice
* Created: Tue Sep  1 20:19:16 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hs__o41a_2.pex.spice"
.subckt sky130_fd_sc_hs__o41a_2  VNB VPB A1 A2 A3 A4 B1 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* B1	B1
* A4	A4
* A3	A3
* A2	A2
* A1	A1
* VPB	VPB
* VNB	VNB
MM1011 N_VGND_M1011_d N_A1_M1011_g N_A_27_74#_M1011_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1554 AS=0.2109 PD=1.16 PS=2.05 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75002.5 A=0.111 P=1.78 MULT=1
MM1013 N_A_27_74#_M1013_d N_A2_M1013_g N_VGND_M1011_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1554 PD=1.02 PS=1.16 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75000.8
+ SB=75001.9 A=0.111 P=1.78 MULT=1
MM1006 N_VGND_M1006_d N_A3_M1006_g N_A_27_74#_M1013_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.21645 AS=0.1036 PD=1.325 PS=1.02 NRD=25.944 NRS=0 M=1 R=4.93333
+ SA=75001.2 SB=75001.5 A=0.111 P=1.78 MULT=1
MM1004 N_A_27_74#_M1004_d N_A4_M1004_g N_VGND_M1006_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.10915 AS=0.21645 PD=1.035 PS=1.325 NRD=2.424 NRS=23.508 M=1 R=4.93333
+ SA=75001.9 SB=75000.7 A=0.111 P=1.78 MULT=1
MM1009 N_A_428_368#_M1009_d N_B1_M1009_g N_A_27_74#_M1004_d VNB NLOWVT L=0.15
+ W=0.74 AD=0.2627 AS=0.10915 PD=2.19 PS=1.035 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75002.4 SB=75000.3 A=0.111 P=1.78 MULT=1
MM1005 N_X_M1005_d N_A_428_368#_M1005_g N_VGND_M1005_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.2627 PD=1.02 PS=2.19 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.3
+ SB=75000.7 A=0.111 P=1.78 MULT=1
MM1008 N_X_M1005_d N_A_428_368#_M1008_g N_VGND_M1008_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.2627 PD=1.02 PS=2.19 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.7
+ SB=75000.3 A=0.111 P=1.78 MULT=1
MM1007 A_116_368# N_A1_M1007_g N_VPWR_M1007_s VPB PSHORT L=0.15 W=1.12 AD=0.1512
+ AS=0.3304 PD=1.39 PS=2.83 NRD=14.0658 NRS=1.7533 M=1 R=7.46667 SA=75000.2
+ SB=75003.8 A=0.168 P=2.54 MULT=1
MM1001 A_200_368# N_A2_M1001_g A_116_368# VPB PSHORT L=0.15 W=1.12 AD=0.2352
+ AS=0.1512 PD=1.54 PS=1.39 NRD=27.2451 NRS=14.0658 M=1 R=7.46667 SA=75000.6
+ SB=75003.4 A=0.168 P=2.54 MULT=1
MM1012 A_314_368# N_A3_M1012_g A_200_368# VPB PSHORT L=0.15 W=1.12 AD=0.2352
+ AS=0.2352 PD=1.54 PS=1.54 NRD=27.2451 NRS=27.2451 M=1 R=7.46667 SA=75001.2
+ SB=75002.8 A=0.168 P=2.54 MULT=1
MM1010 N_A_428_368#_M1010_d N_A4_M1010_g A_314_368# VPB PSHORT L=0.15 W=1.12
+ AD=0.240589 AS=0.2352 PD=1.62717 PS=1.54 NRD=1.7533 NRS=27.2451 M=1 R=7.46667
+ SA=75001.8 SB=75002.2 A=0.168 P=2.54 MULT=1
MM1000 N_VPWR_M1000_d N_B1_M1000_g N_A_428_368#_M1010_d VPB PSHORT L=0.15 W=1
+ AD=0.515 AS=0.214811 PD=2.0566 PS=1.45283 NRD=1.9503 NRS=25.9252 M=1 R=6.66667
+ SA=75002.3 SB=75001.9 A=0.15 P=2.3 MULT=1
MM1002 N_X_M1002_d N_A_428_368#_M1002_g N_VPWR_M1000_d VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.5768 PD=1.42 PS=2.3034 NRD=1.7533 NRS=2.6201 M=1 R=7.46667
+ SA=75003.2 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1003 N_X_M1002_d N_A_428_368#_M1003_g N_VPWR_M1003_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.3304 PD=1.42 PS=2.83 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75003.6 SB=75000.2 A=0.168 P=2.54 MULT=1
DX14_noxref VNB VPB NWDIODE A=9.6348 P=14.08
*
.include "sky130_fd_sc_hs__o41a_2.pxi.spice"
*
.ends
*
*
