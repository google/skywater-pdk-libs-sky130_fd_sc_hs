* File: sky130_fd_sc_hs__inv_2.spice
* Created: Tue Sep  1 20:06:59 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hs__inv_2.pex.spice"
.subckt sky130_fd_sc_hs__inv_2  VNB VPB A VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A	A
* VPB	VPB
* VNB	VNB
MM1002 N_Y_M1002_d N_A_M1002_g N_VGND_M1002_s VNB NLOWVT L=0.15 W=0.74 AD=0.1036
+ AS=0.2109 PD=1.02 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2 SB=75000.6
+ A=0.111 P=1.78 MULT=1
MM1003 N_Y_M1002_d N_A_M1003_g N_VGND_M1003_s VNB NLOWVT L=0.15 W=0.74 AD=0.1036
+ AS=0.2109 PD=1.02 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.6 SB=75000.2
+ A=0.111 P=1.78 MULT=1
MM1000 N_Y_M1000_d N_A_M1000_g N_VPWR_M1000_s VPB PSHORT L=0.15 W=1.12 AD=0.168
+ AS=0.3192 PD=1.42 PS=2.81 NRD=1.7533 NRS=1.7533 M=1 R=7.46667 SA=75000.2
+ SB=75000.7 A=0.168 P=2.54 MULT=1
MM1001 N_Y_M1000_d N_A_M1001_g N_VPWR_M1001_s VPB PSHORT L=0.15 W=1.12 AD=0.168
+ AS=0.3192 PD=1.42 PS=2.81 NRD=1.7533 NRS=1.7533 M=1 R=7.46667 SA=75000.7
+ SB=75000.2 A=0.168 P=2.54 MULT=1
DX4_noxref VNB VPB NWDIODE A=3.3852 P=7.36
*
.include "sky130_fd_sc_hs__inv_2.pxi.spice"
*
.ends
*
*
