* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hs__sdfrtp_1 CLK D RESET_B SCD SCE VGND VNB VPB VPWR Q
X0 a_1233_118# a_1034_368# a_1319_118# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X1 a_1972_74# a_1997_272# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X2 a_225_81# a_27_88# a_312_81# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X3 a_225_81# RESET_B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X4 a_1367_92# a_1034_368# a_1745_74# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X5 VPWR SCE a_216_464# VPB sky130_fd_pr__pfet_01v8 w=640000u l=150000u
X6 a_855_368# CLK VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X7 a_1367_92# a_855_368# a_1745_74# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=150000u
X8 a_1745_74# a_855_368# a_1972_74# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X9 a_300_464# a_27_88# a_538_464# VPB sky130_fd_pr__pfet_01v8 w=640000u l=150000u
X10 VPWR a_1745_74# a_2399_424# VPB sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X11 VGND a_2399_424# Q VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X12 a_1343_461# a_1367_92# VPWR VPB sky130_fd_pr__pfet_01v8 w=420000u l=150000u
X13 VPWR RESET_B a_1997_272# VPB sky130_fd_pr__pfet_01v8 w=420000u l=150000u
X14 a_1397_118# RESET_B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X15 a_545_81# SCD a_225_81# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X16 a_538_464# SCD VPWR VPB sky130_fd_pr__pfet_01v8 w=640000u l=150000u
X17 VGND a_1745_74# a_2399_424# VNB sky130_fd_pr__nfet_01v8_lvt w=550000u l=150000u
X18 a_300_464# a_855_368# a_1233_118# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X19 a_1233_118# a_855_368# a_1343_461# VPB sky130_fd_pr__pfet_01v8 w=420000u l=150000u
X20 VGND a_855_368# a_1034_368# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X21 VPWR a_1233_118# a_1367_92# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=150000u
X22 a_1319_118# a_1367_92# a_1397_118# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X23 VGND RESET_B a_2135_74# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X24 a_300_464# SCE a_545_81# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X25 a_855_368# CLK VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X26 a_2135_74# a_1745_74# a_1997_272# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X27 a_300_464# a_1034_368# a_1233_118# VPB sky130_fd_pr__pfet_01v8 w=420000u l=150000u
X28 a_1993_508# a_1997_272# VPWR VPB sky130_fd_pr__pfet_01v8 w=420000u l=150000u
X29 a_216_464# D a_300_464# VPB sky130_fd_pr__pfet_01v8 w=640000u l=150000u
X30 VPWR a_855_368# a_1034_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X31 a_1997_272# a_1745_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=420000u l=150000u
X32 a_27_88# SCE VPWR VPB sky130_fd_pr__pfet_01v8 w=640000u l=150000u
X33 a_1745_74# a_1034_368# a_1993_508# VPB sky130_fd_pr__pfet_01v8 w=420000u l=150000u
X34 VGND a_1233_118# a_1367_92# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X35 VPWR RESET_B a_1233_118# VPB sky130_fd_pr__pfet_01v8 w=420000u l=150000u
X36 a_27_88# SCE VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X37 VPWR a_2399_424# Q VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X38 VPWR RESET_B a_300_464# VPB sky130_fd_pr__pfet_01v8 w=640000u l=150000u
X39 a_312_81# D a_300_464# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
.ends
