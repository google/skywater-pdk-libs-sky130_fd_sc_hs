* NGSPICE file created from sky130_fd_sc_hs__xnor3_2.ext - technology: sky130A

.subckt sky130_fd_sc_hs__xnor3_2 A B C VGND VNB VPB VPWR X
M1000 VPWR C a_1027_48# VPB pshort w=640000u l=150000u
+  ad=1.6338e+12p pd=1.205e+07u as=1.856e+11p ps=1.86e+06u
M1001 a_83_247# a_397_21# a_332_373# VNB nlowvt w=640000u l=150000u
+  ad=5.925e+11p pd=4.86e+06u as=4.512e+11p ps=3.97e+06u
M1002 VPWR B a_397_21# VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=3.248e+11p ps=2.82e+06u
M1003 a_332_373# B a_27_373# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=3.886e+11p ps=3.85e+06u
M1004 a_83_247# A VPWR VPB pshort w=1e+06u l=150000u
+  ad=7.498e+11p pd=5.67e+06u as=0p ps=0u
M1005 a_27_373# a_397_21# a_329_81# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=4.22e+11p ps=4.25e+06u
M1006 a_83_247# a_397_21# a_329_81# VPB pshort w=840000u l=150000u
+  ad=0p pd=0u as=5.522e+11p ps=4.72e+06u
M1007 X a_1057_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.072e+11p pd=2.04e+06u as=1.54235e+12p ps=1.041e+07u
M1008 a_83_247# A VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_332_373# B a_83_247# VPB pshort w=840000u l=150000u
+  ad=5.92e+11p pd=4.86e+06u as=0p ps=0u
M1010 VGND a_83_247# a_27_373# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VGND C a_1027_48# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.197e+11p ps=1.41e+06u
M1012 X a_1057_74# VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=3.36e+11p pd=2.84e+06u as=0p ps=0u
M1013 a_1057_74# a_1027_48# a_332_373# VPB pshort w=840000u l=150000u
+  ad=4.2765e+11p pd=2.87e+06u as=0p ps=0u
M1014 a_329_81# C a_1057_74# VPB pshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VPWR a_1057_74# X VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VGND B a_397_21# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1017 VGND a_1057_74# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_27_373# a_397_21# a_332_373# VPB pshort w=640000u l=150000u
+  ad=4.998e+11p pd=4.51e+06u as=0p ps=0u
M1019 a_329_81# B a_83_247# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_332_373# C a_1057_74# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=2.24e+11p ps=1.98e+06u
M1021 a_329_81# B a_27_373# VPB pshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 VPWR a_83_247# a_27_373# VPB pshort w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_1057_74# a_1027_48# a_329_81# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

