* File: sky130_fd_sc_hs__a31oi_1.pex.spice
* Created: Thu Aug 27 20:29:31 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HS__A31OI_1%A3 1 3 4 6 8 9
r25 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.29
+ $Y=1.385 $X2=0.29 $Y2=1.385
r26 9 13 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=0.29 $Y=1.295 $X2=0.29
+ $Y2=1.385
r27 8 12 39.3438 $w=3.3e-07 $l=2.25e-07 $layer=POLY_cond $X=0.515 $Y=1.385
+ $X2=0.29 $Y2=1.385
r28 4 8 43.1139 $w=1.98e-07 $l=1.79374e-07 $layer=POLY_cond $X=0.65 $Y=1.22
+ $X2=0.62 $Y2=1.385
r29 4 6 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=0.65 $Y=1.22 $X2=0.65
+ $Y2=0.74
r30 1 8 95.4523 $w=1.98e-07 $l=3.87427e-07 $layer=POLY_cond $X=0.605 $Y=1.765
+ $X2=0.62 $Y2=1.385
r31 1 3 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.605 $Y=1.765
+ $X2=0.605 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_HS__A31OI_1%A2 1 3 4 6 7 8
c28 1 0 3.79312e-20 $X=1.04 $Y=1.22
r29 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.13
+ $Y=1.385 $X2=1.13 $Y2=1.385
r30 8 13 2.96342 $w=3.48e-07 $l=9e-08 $layer=LI1_cond $X=1.14 $Y=1.295 $X2=1.14
+ $Y2=1.385
r31 7 8 12.183 $w=3.48e-07 $l=3.7e-07 $layer=LI1_cond $X=1.14 $Y=0.925 $X2=1.14
+ $Y2=1.295
r32 4 12 77.2841 $w=2.7e-07 $l=4.15812e-07 $layer=POLY_cond $X=1.055 $Y=1.765
+ $X2=1.13 $Y2=1.385
r33 4 6 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.055 $Y=1.765
+ $X2=1.055 $Y2=2.4
r34 1 12 38.9026 $w=2.7e-07 $l=2.05122e-07 $layer=POLY_cond $X=1.04 $Y=1.22
+ $X2=1.13 $Y2=1.385
r35 1 3 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.04 $Y=1.22 $X2=1.04
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HS__A31OI_1%A1 1 3 4 6 7
c32 7 0 1.697e-19 $X=1.68 $Y=1.295
c33 1 0 1.15392e-19 $X=1.61 $Y=1.22
r34 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.7
+ $Y=1.385 $X2=1.7 $Y2=1.385
r35 7 11 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=1.7 $Y=1.295 $X2=1.7
+ $Y2=1.385
r36 4 10 77.2841 $w=2.7e-07 $l=3.82492e-07 $layer=POLY_cond $X=1.695 $Y=1.765
+ $X2=1.7 $Y2=1.385
r37 4 6 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.695 $Y=1.765
+ $X2=1.695 $Y2=2.4
r38 1 10 38.9026 $w=2.7e-07 $l=2.05122e-07 $layer=POLY_cond $X=1.61 $Y=1.22
+ $X2=1.7 $Y2=1.385
r39 1 3 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.61 $Y=1.22 $X2=1.61
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HS__A31OI_1%B1 3 4 6 8 9 10 11 15
c27 11 0 1.15392e-19 $X=2.64 $Y=1.295
c28 9 0 1.31769e-19 $X=2.195 $Y=1.22
r29 15 16 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.61
+ $Y=1.385 $X2=2.61 $Y2=1.385
r30 11 16 0.934413 $w=3.68e-07 $l=3e-08 $layer=LI1_cond $X=2.64 $Y=1.365
+ $X2=2.61 $Y2=1.365
r31 10 16 14.0162 $w=3.68e-07 $l=4.5e-07 $layer=LI1_cond $X=2.16 $Y=1.365
+ $X2=2.61 $Y2=1.365
r32 8 15 56.8299 $w=3.3e-07 $l=3.25e-07 $layer=POLY_cond $X=2.285 $Y=1.385
+ $X2=2.61 $Y2=1.385
r33 8 9 66.2869 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=2.195 $Y=1.385
+ $X2=2.195 $Y2=1.22
r34 4 8 149.859 $w=1.8e-07 $l=3.8e-07 $layer=POLY_cond $X=2.195 $Y=1.765
+ $X2=2.195 $Y2=1.385
r35 4 6 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.195 $Y=1.765
+ $X2=2.195 $Y2=2.4
r36 3 9 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=2.18 $Y=0.74 $X2=2.18
+ $Y2=1.22
.ends

.subckt PM_SKY130_FD_SC_HS__A31OI_1%VPWR 1 2 7 9 15 18 19 20 30 31
r35 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r36 30 31 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r37 28 31 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.64 $Y2=3.33
r38 27 30 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.68 $Y=3.33 $X2=2.64
+ $Y2=3.33
r39 27 28 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r40 25 35 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.24 $Y2=3.33
r41 24 25 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r42 22 34 4.70928 $w=1.7e-07 $l=2.28e-07 $layer=LI1_cond $X=0.455 $Y=3.33
+ $X2=0.227 $Y2=3.33
r43 22 24 48.6043 $w=1.68e-07 $l=7.45e-07 $layer=LI1_cond $X=0.455 $Y=3.33
+ $X2=1.2 $Y2=3.33
r44 20 28 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.44 $Y=3.33
+ $X2=1.68 $Y2=3.33
r45 20 25 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.44 $Y=3.33
+ $X2=1.2 $Y2=3.33
r46 18 24 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=1.205 $Y=3.33 $X2=1.2
+ $Y2=3.33
r47 18 19 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.205 $Y=3.33
+ $X2=1.37 $Y2=3.33
r48 17 27 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=1.535 $Y=3.33
+ $X2=1.68 $Y2=3.33
r49 17 19 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.535 $Y=3.33
+ $X2=1.37 $Y2=3.33
r50 13 19 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.37 $Y=3.245
+ $X2=1.37 $Y2=3.33
r51 13 15 26.5411 $w=3.28e-07 $l=7.6e-07 $layer=LI1_cond $X=1.37 $Y=3.245
+ $X2=1.37 $Y2=2.485
r52 9 12 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=0.29 $Y=1.985
+ $X2=0.29 $Y2=2.815
r53 7 34 3.0569 $w=3.3e-07 $l=1.12161e-07 $layer=LI1_cond $X=0.29 $Y=3.245
+ $X2=0.227 $Y2=3.33
r54 7 12 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=0.29 $Y=3.245
+ $X2=0.29 $Y2=2.815
r55 2 15 300 $w=1.7e-07 $l=7.5553e-07 $layer=licon1_PDIFF $count=2 $X=1.13
+ $Y=1.84 $X2=1.37 $Y2=2.485
r56 1 12 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=0.145
+ $Y=1.84 $X2=0.29 $Y2=2.815
r57 1 9 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.145
+ $Y=1.84 $X2=0.29 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HS__A31OI_1%A_136_368# 1 2 7 9 11 13 15
r31 13 20 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.92 $Y=2.23 $X2=1.92
+ $Y2=2.145
r32 13 15 20.7789 $w=3.28e-07 $l=5.95e-07 $layer=LI1_cond $X=1.92 $Y=2.23
+ $X2=1.92 $Y2=2.825
r33 12 18 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.995 $Y=2.145
+ $X2=0.83 $Y2=2.145
r34 11 20 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.755 $Y=2.145
+ $X2=1.92 $Y2=2.145
r35 11 12 49.5829 $w=1.68e-07 $l=7.6e-07 $layer=LI1_cond $X=1.755 $Y=2.145
+ $X2=0.995 $Y2=2.145
r36 7 18 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.83 $Y=2.23 $X2=0.83
+ $Y2=2.145
r37 7 9 20.7789 $w=3.28e-07 $l=5.95e-07 $layer=LI1_cond $X=0.83 $Y=2.23 $X2=0.83
+ $Y2=2.825
r38 2 20 400 $w=1.7e-07 $l=3.72525e-07 $layer=licon1_PDIFF $count=1 $X=1.77
+ $Y=1.84 $X2=1.92 $Y2=2.145
r39 2 15 400 $w=1.7e-07 $l=1.05734e-06 $layer=licon1_PDIFF $count=1 $X=1.77
+ $Y=1.84 $X2=1.92 $Y2=2.825
r40 1 18 400 $w=1.7e-07 $l=3.72525e-07 $layer=licon1_PDIFF $count=1 $X=0.68
+ $Y=1.84 $X2=0.83 $Y2=2.145
r41 1 9 400 $w=1.7e-07 $l=1.05734e-06 $layer=licon1_PDIFF $count=1 $X=0.68
+ $Y=1.84 $X2=0.83 $Y2=2.825
.ends

.subckt PM_SKY130_FD_SC_HS__A31OI_1%Y 1 2 8 9 10 11 12 16 18 19 20 25
r56 20 33 0.956863 $w=4.98e-07 $l=4e-08 $layer=LI1_cond $X=2.505 $Y=2.775
+ $X2=2.505 $Y2=2.815
r57 19 20 8.85098 $w=4.98e-07 $l=3.7e-07 $layer=LI1_cond $X=2.505 $Y=2.405
+ $X2=2.505 $Y2=2.775
r58 18 19 8.85098 $w=4.98e-07 $l=3.7e-07 $layer=LI1_cond $X=2.505 $Y=2.035
+ $X2=2.505 $Y2=2.405
r59 18 25 1.19608 $w=4.98e-07 $l=5e-08 $layer=LI1_cond $X=2.505 $Y=2.035
+ $X2=2.505 $Y2=1.985
r60 17 25 2.27255 $w=4.98e-07 $l=9.5e-08 $layer=LI1_cond $X=2.505 $Y=1.89
+ $X2=2.505 $Y2=1.985
r61 11 17 9.23067 $w=1.7e-07 $l=2.89396e-07 $layer=LI1_cond $X=2.255 $Y=1.805
+ $X2=2.505 $Y2=1.89
r62 11 12 95.2513 $w=1.68e-07 $l=1.46e-06 $layer=LI1_cond $X=2.255 $Y=1.805
+ $X2=0.795 $Y2=1.805
r63 9 16 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.73 $Y=0.435
+ $X2=1.895 $Y2=0.435
r64 9 10 61 $w=1.68e-07 $l=9.35e-07 $layer=LI1_cond $X=1.73 $Y=0.435 $X2=0.795
+ $Y2=0.435
r65 8 12 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.71 $Y=1.72
+ $X2=0.795 $Y2=1.805
r66 7 10 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.71 $Y=0.52
+ $X2=0.795 $Y2=0.435
r67 7 8 78.2888 $w=1.68e-07 $l=1.2e-06 $layer=LI1_cond $X=0.71 $Y=0.52 $X2=0.71
+ $Y2=1.72
r68 2 33 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=2.27
+ $Y=1.84 $X2=2.42 $Y2=2.815
r69 2 25 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=2.27
+ $Y=1.84 $X2=2.42 $Y2=1.985
r70 1 16 91 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=2 $X=1.685
+ $Y=0.37 $X2=1.895 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__A31OI_1%VGND 1 2 7 9 13 16 17 18 28 29
r31 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r32 28 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r33 26 29 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r34 25 26 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r35 23 33 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r36 22 25 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=0.72 $Y=0 $X2=2.16
+ $Y2=0
r37 22 23 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r38 20 32 4.70928 $w=1.7e-07 $l=2.28e-07 $layer=LI1_cond $X=0.455 $Y=0 $X2=0.227
+ $Y2=0
r39 20 22 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.455 $Y=0 $X2=0.72
+ $Y2=0
r40 18 26 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.44 $Y=0 $X2=2.16
+ $Y2=0
r41 18 23 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.44 $Y=0 $X2=0.72
+ $Y2=0
r42 16 25 4.56684 $w=1.68e-07 $l=7e-08 $layer=LI1_cond $X=2.23 $Y=0 $X2=2.16
+ $Y2=0
r43 16 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.23 $Y=0 $X2=2.395
+ $Y2=0
r44 15 28 5.21925 $w=1.68e-07 $l=8e-08 $layer=LI1_cond $X=2.56 $Y=0 $X2=2.64
+ $Y2=0
r45 15 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.56 $Y=0 $X2=2.395
+ $Y2=0
r46 11 17 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.395 $Y=0.085
+ $X2=2.395 $Y2=0
r47 11 13 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=2.395 $Y=0.085
+ $X2=2.395 $Y2=0.515
r48 7 32 3.0569 $w=3.3e-07 $l=1.12161e-07 $layer=LI1_cond $X=0.29 $Y=0.085
+ $X2=0.227 $Y2=0
r49 7 9 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=0.29 $Y=0.085 $X2=0.29
+ $Y2=0.515
r50 2 13 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.255
+ $Y=0.37 $X2=2.395 $Y2=0.515
r51 1 9 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.145
+ $Y=0.37 $X2=0.29 $Y2=0.515
.ends

