/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */

`ifndef SKY130_FD_SC_HS__MUX4_SYMBOL_V
`define SKY130_FD_SC_HS__MUX4_SYMBOL_V

/**
 * mux4: 4-input multiplexer.
 *
 * Verilog stub (without power pins) for graphical symbol definition
 * generation.
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none

(* blackbox *)
module sky130_fd_sc_hs__mux4 (
    //# {{data|Data Signals}}
    input  A0,
    input  A1,
    input  A2,
    input  A3,
    output X ,

    //# {{control|Control Signals}}
    input  S0,
    input  S1
);

    // Voltage supply signals
    supply1 VPWR;
    supply0 VGND;

endmodule

`default_nettype wire
`endif  // SKY130_FD_SC_HS__MUX4_SYMBOL_V
