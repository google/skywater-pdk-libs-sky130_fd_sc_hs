# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_hs__o21ba_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hs__o21ba_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.840000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.261000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.405000 1.180000 3.735000 1.550000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.261000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.720000 1.180000 3.235000 1.550000 ;
    END
  END A2
  PIN B1_N
    ANTENNAGATEAREA  0.208500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.300000 0.455000 1.780000 ;
    END
  END B1_N
  PIN X
    ANTENNADIFFAREA  0.543200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.010000 0.350000 1.340000 1.130000 ;
        RECT 1.010000 1.130000 1.180000 1.820000 ;
        RECT 1.010000 1.820000 1.440000 2.070000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 3.840000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 3.840000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.840000 0.085000 ;
      RECT 0.000000  3.245000 3.840000 3.415000 ;
      RECT 0.105000  0.455000 0.355000 0.960000 ;
      RECT 0.105000  0.960000 0.795000 1.130000 ;
      RECT 0.115000  1.950000 0.795000 2.240000 ;
      RECT 0.115000  2.240000 2.210000 2.410000 ;
      RECT 0.115000  2.410000 0.445000 2.700000 ;
      RECT 0.535000  0.085000 0.785000 0.790000 ;
      RECT 0.625000  1.130000 0.795000 1.950000 ;
      RECT 0.650000  2.580000 0.980000 3.245000 ;
      RECT 1.350000  1.300000 1.680000 1.630000 ;
      RECT 1.510000  1.010000 2.550000 1.180000 ;
      RECT 1.510000  1.180000 1.680000 1.300000 ;
      RECT 1.520000  0.085000 1.770000 0.820000 ;
      RECT 1.565000  2.580000 2.235000 3.245000 ;
      RECT 1.890000  1.350000 2.210000 2.240000 ;
      RECT 1.980000  0.350000 2.230000 1.010000 ;
      RECT 2.380000  1.180000 2.550000 1.820000 ;
      RECT 2.380000  1.820000 2.775000 2.410000 ;
      RECT 2.410000  0.350000 2.740000 0.670000 ;
      RECT 2.410000  0.670000 3.740000 0.840000 ;
      RECT 2.445000  2.410000 2.775000 2.860000 ;
      RECT 2.910000  0.085000 3.240000 0.500000 ;
      RECT 3.405000  1.820000 3.735000 3.245000 ;
      RECT 3.410000  0.350000 3.740000 0.670000 ;
      RECT 3.410000  0.840000 3.740000 1.010000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
  END
END sky130_fd_sc_hs__o21ba_2
END LIBRARY
