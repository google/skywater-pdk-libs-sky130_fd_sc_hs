* File: sky130_fd_sc_hs__and4_1.spice
* Created: Tue Sep  1 19:55:44 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hs__and4_1.pex.spice"
.subckt sky130_fd_sc_hs__and4_1  VNB VPB A B C D VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* D	D
* C	C
* B	B
* A	A
* VPB	VPB
* VNB	VNB
MM1009 A_179_74# N_A_M1009_g N_A_96_74#_M1009_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.0768 AS=0.1696 PD=0.88 PS=1.81 NRD=12.18 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75002.1 A=0.096 P=1.58 MULT=1
MM1006 A_257_74# N_B_M1006_g A_179_74# VNB NLOWVT L=0.15 W=0.64 AD=0.0768
+ AS=0.0768 PD=0.88 PS=0.88 NRD=12.18 NRS=12.18 M=1 R=4.26667 SA=75000.6
+ SB=75001.7 A=0.096 P=1.58 MULT=1
MM1007 A_335_74# N_C_M1007_g A_257_74# VNB NLOWVT L=0.15 W=0.64 AD=0.1344
+ AS=0.0768 PD=1.06 PS=0.88 NRD=29.052 NRS=12.18 M=1 R=4.26667 SA=75001
+ SB=75001.3 A=0.096 P=1.58 MULT=1
MM1000 N_VGND_M1000_d N_D_M1000_g A_335_74# VNB NLOWVT L=0.15 W=0.64 AD=0.118446
+ AS=0.1344 PD=1.02029 PS=1.06 NRD=0 NRS=29.052 M=1 R=4.26667 SA=75001.5
+ SB=75000.7 A=0.096 P=1.58 MULT=1
MM1001 N_X_M1001_d N_A_96_74#_M1001_g N_VGND_M1000_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.136954 PD=2.05 PS=1.17971 NRD=0 NRS=12.972 M=1 R=4.93333
+ SA=75001.8 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1005 N_A_96_74#_M1005_d N_A_M1005_g N_VPWR_M1005_s VPB PSHORT L=0.15 W=0.84
+ AD=0.147 AS=0.2898 PD=1.19 PS=2.37 NRD=2.3443 NRS=14.0658 M=1 R=5.6 SA=75000.3
+ SB=75002.5 A=0.126 P=1.98 MULT=1
MM1002 N_VPWR_M1002_d N_B_M1002_g N_A_96_74#_M1005_d VPB PSHORT L=0.15 W=0.84
+ AD=0.2352 AS=0.147 PD=1.4 PS=1.19 NRD=32.8202 NRS=14.0658 M=1 R=5.6 SA=75000.8
+ SB=75002 A=0.126 P=1.98 MULT=1
MM1003 N_A_96_74#_M1003_d N_C_M1003_g N_VPWR_M1002_d VPB PSHORT L=0.15 W=0.84
+ AD=0.147 AS=0.2352 PD=1.19 PS=1.4 NRD=14.0658 NRS=32.8202 M=1 R=5.6 SA=75001.5
+ SB=75001.3 A=0.126 P=1.98 MULT=1
MM1004 N_VPWR_M1004_d N_D_M1004_g N_A_96_74#_M1003_d VPB PSHORT L=0.15 W=0.84
+ AD=0.1884 AS=0.147 PD=1.33286 PS=1.19 NRD=22.261 NRS=2.3443 M=1 R=5.6 SA=75002
+ SB=75000.8 A=0.126 P=1.98 MULT=1
MM1008 N_X_M1008_d N_A_96_74#_M1008_g N_VPWR_M1004_d VPB PSHORT L=0.15 W=1.12
+ AD=0.3304 AS=0.2512 PD=2.83 PS=1.77714 NRD=1.7533 NRS=10.5395 M=1 R=7.46667
+ SA=75002 SB=75000.2 A=0.168 P=2.54 MULT=1
DX10_noxref VNB VPB NWDIODE A=6.9564 P=11.2
*
.include "sky130_fd_sc_hs__and4_1.pxi.spice"
*
.ends
*
*
