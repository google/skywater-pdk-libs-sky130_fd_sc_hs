* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hs__xnor2_1 A B VGND VNB VPB VPWR Y
M1000 VGND A a_293_74# VNB nlowvt w=740000u l=150000u
+  ad=5.4e+11p pd=4.52e+06u as=4.107e+11p ps=4.07e+06u
M1001 a_138_385# A VPWR VPB pshort w=840000u l=150000u
+  ad=2.52e+11p pd=2.28e+06u as=1.19585e+12p ps=8.62e+06u
M1002 VPWR a_138_385# Y VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=4.704e+11p ps=3.08e+06u
M1003 Y B a_376_368# VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=3.024e+11p ps=2.78e+06u
M1004 VPWR B a_138_385# VPB pshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_138_385# B a_112_119# VNB nlowvt w=640000u l=150000u
+  ad=1.76e+11p pd=1.83e+06u as=1.344e+11p ps=1.7e+06u
M1006 Y a_138_385# a_293_74# VNB nlowvt w=740000u l=150000u
+  ad=2.294e+11p pd=2.1e+06u as=0p ps=0u
M1007 a_376_368# A VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_112_119# A VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_293_74# B VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
