* File: sky130_fd_sc_hs__dlxbp_1.spice
* Created: Tue Sep  1 20:02:51 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hs__dlxbp_1.pex.spice"
.subckt sky130_fd_sc_hs__dlxbp_1  VNB VPB D GATE VPWR Q Q_N VGND
* 
* VGND	VGND
* Q_N	Q_N
* Q	Q
* VPWR	VPWR
* GATE	GATE
* D	D
* VPB	VPB
* VNB	VNB
MM1006 N_VGND_M1006_d N_D_M1006_g N_A_27_413#_M1006_s VNB NLOWVT L=0.15 W=0.55
+ AD=0.129591 AS=0.15675 PD=0.997674 PS=1.67 NRD=18 NRS=0 M=1 R=3.66667
+ SA=75000.2 SB=75000.8 A=0.0825 P=1.4 MULT=1
MM1003 N_A_231_74#_M1003_d N_GATE_M1003_g N_VGND_M1006_d VNB NLOWVT L=0.15
+ W=0.74 AD=0.2109 AS=0.174359 PD=2.05 PS=1.34233 NRD=0 NRS=11.34 M=1 R=4.93333
+ SA=75000.7 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1017 N_VGND_M1017_d N_A_231_74#_M1017_g N_A_373_82#_M1017_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.224922 AS=0.2109 PD=1.57116 PS=2.05 NRD=40.368 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75002 A=0.111 P=1.78 MULT=1
MM1013 A_589_80# N_A_27_413#_M1013_g N_VGND_M1017_d VNB NLOWVT L=0.15 W=0.64
+ AD=0.0768 AS=0.194528 PD=0.88 PS=1.35884 NRD=12.18 NRS=21.552 M=1 R=4.26667
+ SA=75000.8 SB=75001.7 A=0.096 P=1.58 MULT=1
MM1012 N_A_664_392#_M1012_d N_A_373_82#_M1012_g A_589_80# VNB NLOWVT L=0.15
+ W=0.64 AD=0.182823 AS=0.0768 PD=1.48528 PS=0.88 NRD=29.052 NRS=12.18 M=1
+ R=4.26667 SA=75001.2 SB=75001.3 A=0.096 P=1.58 MULT=1
MM1004 A_815_124# N_A_231_74#_M1004_g N_A_664_392#_M1012_d VNB NLOWVT L=0.15
+ W=0.42 AD=0.0504 AS=0.119977 PD=0.66 PS=0.974717 NRD=18.564 NRS=44.28 M=1
+ R=2.8 SA=75002 SB=75001.2 A=0.063 P=1.14 MULT=1
MM1019 N_VGND_M1019_d N_A_863_98#_M1019_g A_815_124# VNB NLOWVT L=0.15 W=0.42
+ AD=0.106521 AS=0.0504 PD=0.847241 PS=0.66 NRD=22.848 NRS=18.564 M=1 R=2.8
+ SA=75002.4 SB=75000.8 A=0.063 P=1.14 MULT=1
MM1008 N_A_863_98#_M1008_d N_A_664_392#_M1008_g N_VGND_M1019_d VNB NLOWVT L=0.15
+ W=0.74 AD=0.2109 AS=0.187679 PD=2.05 PS=1.49276 NRD=0 NRS=11.34 M=1 R=4.93333
+ SA=75001.8 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1015 N_VGND_M1015_d N_A_863_98#_M1015_g N_Q_M1015_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.137674 AS=0.2072 PD=1.25054 PS=2.04 NRD=5.664 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75000.6 A=0.111 P=1.78 MULT=1
MM1016 N_A_1347_424#_M1016_d N_A_863_98#_M1016_g N_VGND_M1015_d VNB NLOWVT
+ L=0.15 W=0.55 AD=0.15675 AS=0.102326 PD=1.67 PS=0.929457 NRD=0 NRS=7.632 M=1
+ R=3.66667 SA=75000.7 SB=75000.2 A=0.0825 P=1.4 MULT=1
MM1009 N_Q_N_M1009_d N_A_1347_424#_M1009_g N_VGND_M1009_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.2109 AS=0.2109 PD=2.05 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1018 N_VPWR_M1018_d N_D_M1018_g N_A_27_413#_M1018_s VPB PSHORT L=0.15 W=0.84
+ AD=0.2338 AS=0.2436 PD=1.59 PS=2.26 NRD=52.3626 NRS=2.3443 M=1 R=5.6
+ SA=75000.2 SB=75000.8 A=0.126 P=1.98 MULT=1
MM1020 N_A_231_74#_M1020_d N_GATE_M1020_g N_VPWR_M1018_d VPB PSHORT L=0.15
+ W=0.84 AD=0.2478 AS=0.2338 PD=2.27 PS=1.59 NRD=2.3443 NRS=52.3626 M=1 R=5.6
+ SA=75000.8 SB=75000.2 A=0.126 P=1.98 MULT=1
MM1005 N_VPWR_M1005_d N_A_231_74#_M1005_g N_A_373_82#_M1005_s VPB PSHORT L=0.15
+ W=0.84 AD=0.222623 AS=0.2478 PD=1.4563 PS=2.27 NRD=49.25 NRS=2.3443 M=1 R=5.6
+ SA=75000.2 SB=75001.8 A=0.126 P=1.98 MULT=1
MM1007 A_586_392# N_A_27_413#_M1007_g N_VPWR_M1005_d VPB PSHORT L=0.15 W=1
+ AD=0.12 AS=0.265027 PD=1.24 PS=1.7337 NRD=12.7853 NRS=19.6803 M=1 R=6.66667
+ SA=75000.7 SB=75001.4 A=0.15 P=2.3 MULT=1
MM1000 N_A_664_392#_M1000_d N_A_231_74#_M1000_g A_586_392# VPB PSHORT L=0.15 W=1
+ AD=0.230845 AS=0.12 PD=1.94366 PS=1.24 NRD=1.9503 NRS=12.7853 M=1 R=6.66667
+ SA=75001.1 SB=75001 A=0.15 P=2.3 MULT=1
MM1010 A_770_508# N_A_373_82#_M1010_g N_A_664_392#_M1000_d VPB PSHORT L=0.15
+ W=0.42 AD=0.10605 AS=0.0969549 PD=0.925 PS=0.816338 NRD=92.6294 NRS=82.4642
+ M=1 R=2.8 SA=75001.6 SB=75001.6 A=0.063 P=1.14 MULT=1
MM1001 N_VPWR_M1001_d N_A_863_98#_M1001_g A_770_508# VPB PSHORT L=0.15 W=0.42
+ AD=0.115309 AS=0.10605 PD=0.919091 PS=0.925 NRD=53.9386 NRS=92.6294 M=1 R=2.8
+ SA=75002.2 SB=75000.9 A=0.063 P=1.14 MULT=1
MM1011 N_A_863_98#_M1011_d N_A_664_392#_M1011_g N_VPWR_M1001_d VPB PSHORT L=0.15
+ W=1.12 AD=0.3304 AS=0.307491 PD=2.83 PS=2.45091 NRD=1.7533 NRS=29.8849 M=1
+ R=7.46667 SA=75001.2 SB=75000.2 A=0.168 P=2.54 MULT=1
MM1002 N_VPWR_M1002_d N_A_863_98#_M1002_g N_Q_M1002_s VPB PSHORT L=0.15 W=1.12
+ AD=0.2128 AS=0.3304 PD=1.68571 PS=2.83 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75000.6 A=0.168 P=2.54 MULT=1
MM1021 N_A_1347_424#_M1021_d N_A_863_98#_M1021_g N_VPWR_M1002_d VPB PSHORT
+ L=0.15 W=0.84 AD=0.2436 AS=0.1596 PD=2.26 PS=1.26429 NRD=2.3443 NRS=15.2281
+ M=1 R=5.6 SA=75000.7 SB=75000.2 A=0.126 P=1.98 MULT=1
MM1014 N_Q_N_M1014_d N_A_1347_424#_M1014_g N_VPWR_M1014_s VPB PSHORT L=0.15
+ W=1.12 AD=0.3248 AS=0.3248 PD=2.82 PS=2.82 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75000.2 SB=75000.2 A=0.168 P=2.54 MULT=1
DX22_noxref VNB VPB NWDIODE A=15.8844 P=20.8
*
.include "sky130_fd_sc_hs__dlxbp_1.pxi.spice"
*
.ends
*
*
