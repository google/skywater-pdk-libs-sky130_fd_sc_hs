# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_hs__dfrtp_4
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_hs__dfrtp_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  13.44000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.000000 0.515000 2.180000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  1.207100 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 11.035000 1.800000 12.740000 1.970000 ;
        RECT 11.035000 1.970000 11.365000 2.980000 ;
        RECT 11.595000 0.365000 11.910000 0.880000 ;
        RECT 11.595000 0.880000 12.825000 1.130000 ;
        RECT 12.410000 1.610000 13.315000 1.780000 ;
        RECT 12.410000 1.780000 12.740000 1.800000 ;
        RECT 12.410000 1.970000 12.740000 2.980000 ;
        RECT 12.575000 0.350000 12.825000 0.880000 ;
        RECT 12.575000 1.130000 12.825000 1.270000 ;
        RECT 12.575000 1.270000 13.315000 1.610000 ;
    END
  END Q
  PIN RESET_B
    ANTENNAGATEAREA  0.378000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.025000 1.130000 1.285000 2.140000 ;
        RECT 5.085000 1.670000 5.635000 2.120000 ;
        RECT 8.765000 1.920000 9.140000 2.275000 ;
      LAYER mcon ;
        RECT 1.115000 1.950000 1.285000 2.120000 ;
        RECT 5.435000 1.950000 5.605000 2.120000 ;
        RECT 8.795000 1.950000 8.965000 2.120000 ;
      LAYER met1 ;
        RECT 1.055000 1.920000 1.345000 1.965000 ;
        RECT 1.055000 1.965000 9.025000 2.105000 ;
        RECT 1.055000 2.105000 1.345000 2.150000 ;
        RECT 5.375000 1.920000 5.665000 1.965000 ;
        RECT 5.375000 2.105000 5.665000 2.150000 ;
        RECT 8.735000 1.920000 9.025000 1.965000 ;
        RECT 8.735000 2.105000 9.025000 2.150000 ;
    END
  END RESET_B
  PIN CLK
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 1.795000 1.310000 2.275000 1.640000 ;
        RECT 2.045000 1.640000 2.275000 1.780000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT  0.000000 -0.085000 13.440000 0.085000 ;
        RECT  1.065000  0.085000  1.235000 0.830000 ;
        RECT  2.045000  0.085000  2.375000 0.800000 ;
        RECT  4.895000  0.085000  5.225000 0.370000 ;
        RECT  8.625000  0.085000  8.955000 0.845000 ;
        RECT 10.115000  0.085000 10.390000 1.130000 ;
        RECT 11.120000  0.085000 11.410000 1.130000 ;
        RECT 12.080000  0.085000 12.405000 0.710000 ;
        RECT 13.005000  0.085000 13.335000 1.100000 ;
      LAYER mcon ;
        RECT  0.155000 -0.085000  0.325000 0.085000 ;
        RECT  0.635000 -0.085000  0.805000 0.085000 ;
        RECT  1.115000 -0.085000  1.285000 0.085000 ;
        RECT  1.595000 -0.085000  1.765000 0.085000 ;
        RECT  2.075000 -0.085000  2.245000 0.085000 ;
        RECT  2.555000 -0.085000  2.725000 0.085000 ;
        RECT  3.035000 -0.085000  3.205000 0.085000 ;
        RECT  3.515000 -0.085000  3.685000 0.085000 ;
        RECT  3.995000 -0.085000  4.165000 0.085000 ;
        RECT  4.475000 -0.085000  4.645000 0.085000 ;
        RECT  4.955000 -0.085000  5.125000 0.085000 ;
        RECT  5.435000 -0.085000  5.605000 0.085000 ;
        RECT  5.915000 -0.085000  6.085000 0.085000 ;
        RECT  6.395000 -0.085000  6.565000 0.085000 ;
        RECT  6.875000 -0.085000  7.045000 0.085000 ;
        RECT  7.355000 -0.085000  7.525000 0.085000 ;
        RECT  7.835000 -0.085000  8.005000 0.085000 ;
        RECT  8.315000 -0.085000  8.485000 0.085000 ;
        RECT  8.795000 -0.085000  8.965000 0.085000 ;
        RECT  9.275000 -0.085000  9.445000 0.085000 ;
        RECT  9.755000 -0.085000  9.925000 0.085000 ;
        RECT 10.235000 -0.085000 10.405000 0.085000 ;
        RECT 10.715000 -0.085000 10.885000 0.085000 ;
        RECT 11.195000 -0.085000 11.365000 0.085000 ;
        RECT 11.675000 -0.085000 11.845000 0.085000 ;
        RECT 12.155000 -0.085000 12.325000 0.085000 ;
        RECT 12.635000 -0.085000 12.805000 0.085000 ;
        RECT 13.115000 -0.085000 13.285000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.245000 13.440000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT  0.000000 3.245000 13.440000 3.415000 ;
        RECT  0.110000 2.520000  0.360000 3.245000 ;
        RECT  1.090000 2.650000  1.340000 3.245000 ;
        RECT  2.005000 2.680000  2.335000 3.245000 ;
        RECT  4.400000 2.740000  4.730000 3.245000 ;
        RECT  5.830000 2.745000  6.165000 3.245000 ;
        RECT  8.580000 2.445000  8.910000 3.245000 ;
        RECT  9.650000 2.445000  9.900000 3.245000 ;
        RECT 10.535000 2.025000 10.865000 3.245000 ;
        RECT 11.535000 2.140000 12.240000 3.245000 ;
        RECT 12.910000 1.950000 13.240000 3.245000 ;
      LAYER mcon ;
        RECT  0.155000 3.245000  0.325000 3.415000 ;
        RECT  0.635000 3.245000  0.805000 3.415000 ;
        RECT  1.115000 3.245000  1.285000 3.415000 ;
        RECT  1.595000 3.245000  1.765000 3.415000 ;
        RECT  2.075000 3.245000  2.245000 3.415000 ;
        RECT  2.555000 3.245000  2.725000 3.415000 ;
        RECT  3.035000 3.245000  3.205000 3.415000 ;
        RECT  3.515000 3.245000  3.685000 3.415000 ;
        RECT  3.995000 3.245000  4.165000 3.415000 ;
        RECT  4.475000 3.245000  4.645000 3.415000 ;
        RECT  4.955000 3.245000  5.125000 3.415000 ;
        RECT  5.435000 3.245000  5.605000 3.415000 ;
        RECT  5.915000 3.245000  6.085000 3.415000 ;
        RECT  6.395000 3.245000  6.565000 3.415000 ;
        RECT  6.875000 3.245000  7.045000 3.415000 ;
        RECT  7.355000 3.245000  7.525000 3.415000 ;
        RECT  7.835000 3.245000  8.005000 3.415000 ;
        RECT  8.315000 3.245000  8.485000 3.415000 ;
        RECT  8.795000 3.245000  8.965000 3.415000 ;
        RECT  9.275000 3.245000  9.445000 3.415000 ;
        RECT  9.755000 3.245000  9.925000 3.415000 ;
        RECT 10.235000 3.245000 10.405000 3.415000 ;
        RECT 10.715000 3.245000 10.885000 3.415000 ;
        RECT 11.195000 3.245000 11.365000 3.415000 ;
        RECT 11.675000 3.245000 11.845000 3.415000 ;
        RECT 12.155000 3.245000 12.325000 3.415000 ;
        RECT 12.635000 3.245000 12.805000 3.415000 ;
        RECT 13.115000 3.245000 13.285000 3.415000 ;
      LAYER met1 ;
        RECT 0.000000 3.085000 13.440000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.165000 0.370000  0.495000 0.660000 ;
      RECT  0.165000 0.660000  0.855000 0.830000 ;
      RECT  0.560000 2.520000  0.890000 2.980000 ;
      RECT  0.685000 0.830000  0.855000 2.310000 ;
      RECT  0.685000 2.310000  1.680000 2.340000 ;
      RECT  0.685000 2.340000  3.360000 2.480000 ;
      RECT  0.685000 2.480000  0.890000 2.520000 ;
      RECT  1.455000 0.350000  1.875000 0.970000 ;
      RECT  1.455000 0.970000  2.675000 1.140000 ;
      RECT  1.455000 1.140000  1.625000 1.810000 ;
      RECT  1.455000 1.810000  1.805000 2.140000 ;
      RECT  1.510000 2.480000  3.360000 2.510000 ;
      RECT  2.445000 1.140000  2.675000 1.550000 ;
      RECT  2.455000 1.720000  3.455000 1.890000 ;
      RECT  2.455000 1.890000  2.845000 2.170000 ;
      RECT  2.545000 0.330000  4.475000 0.500000 ;
      RECT  2.545000 0.500000  3.015000 0.800000 ;
      RECT  2.845000 0.800000  3.015000 1.720000 ;
      RECT  3.030000 2.060000  3.795000 2.230000 ;
      RECT  3.030000 2.230000  3.360000 2.340000 ;
      RECT  3.030000 2.510000  3.360000 2.755000 ;
      RECT  3.185000 0.670000  3.435000 1.220000 ;
      RECT  3.185000 1.220000  3.795000 1.390000 ;
      RECT  3.190000 1.560000  3.455000 1.720000 ;
      RECT  3.560000 2.400000  5.180000 2.570000 ;
      RECT  3.560000 2.570000  3.810000 2.755000 ;
      RECT  3.605000 0.670000  3.935000 0.880000 ;
      RECT  3.605000 0.880000  4.135000 1.050000 ;
      RECT  3.625000 1.390000  3.795000 2.060000 ;
      RECT  3.965000 1.050000  4.135000 2.400000 ;
      RECT  4.305000 0.500000  4.475000 0.540000 ;
      RECT  4.305000 0.540000  5.565000 0.710000 ;
      RECT  4.305000 0.880000  6.990000 1.050000 ;
      RECT  4.305000 1.050000  4.570000 2.105000 ;
      RECT  4.745000 1.220000  5.985000 1.500000 ;
      RECT  4.745000 1.500000  4.915000 2.295000 ;
      RECT  4.745000 2.295000  5.180000 2.400000 ;
      RECT  4.915000 2.570000  5.180000 2.755000 ;
      RECT  5.395000 0.255000  8.275000 0.425000 ;
      RECT  5.395000 0.425000  5.565000 0.540000 ;
      RECT  5.395000 2.290000  5.725000 2.405000 ;
      RECT  5.395000 2.405000  6.955000 2.575000 ;
      RECT  5.735000 0.720000  6.990000 0.880000 ;
      RECT  6.155000 1.050000  6.325000 1.940000 ;
      RECT  6.155000 1.940000  6.615000 2.235000 ;
      RECT  6.495000 1.260000  6.955000 1.590000 ;
      RECT  6.785000 1.590000  6.955000 2.405000 ;
      RECT  7.125000 2.475000  8.410000 2.805000 ;
      RECT  7.160000 0.595000  7.935000 0.845000 ;
      RECT  7.160000 0.845000  7.330000 2.475000 ;
      RECT  7.545000 1.015000  8.275000 1.345000 ;
      RECT  7.740000 1.345000  8.070000 2.305000 ;
      RECT  8.105000 0.425000  8.275000 1.015000 ;
      RECT  8.240000 1.535000  9.605000 1.705000 ;
      RECT  8.240000 1.705000  8.410000 2.475000 ;
      RECT  8.445000 1.035000  9.945000 1.205000 ;
      RECT  8.445000 1.205000  8.775000 1.365000 ;
      RECT  9.080000 2.445000  9.480000 2.905000 ;
      RECT  9.310000 1.875000  9.945000 2.045000 ;
      RECT  9.310000 2.045000  9.480000 2.445000 ;
      RECT  9.345000 1.375000  9.605000 1.535000 ;
      RECT  9.500000 0.385000  9.830000 1.035000 ;
      RECT  9.775000 1.205000  9.945000 1.875000 ;
      RECT 10.115000 1.460000 12.240000 1.630000 ;
      RECT 10.115000 1.630000 10.365000 2.905000 ;
      RECT 10.560000 0.350000 10.890000 1.300000 ;
      RECT 10.560000 1.300000 12.240000 1.460000 ;
  END
END sky130_fd_sc_hs__dfrtp_4
