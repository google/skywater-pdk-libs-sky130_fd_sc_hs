* File: sky130_fd_sc_hs__bufinv_16.pex.spice
* Created: Thu Aug 27 20:35:07 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HS__BUFINV_16%A 3 5 7 8 10 13 15 17 20 22 23 24 37 38
r66 38 39 0.647849 $w=3.72e-07 $l=5e-09 $layer=POLY_cond $X=1.41 $Y=1.557
+ $X2=1.415 $Y2=1.557
r67 36 38 18.7876 $w=3.72e-07 $l=1.45e-07 $layer=POLY_cond $X=1.265 $Y=1.557
+ $X2=1.41 $Y2=1.557
r68 36 37 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.265
+ $Y=1.515 $X2=1.265 $Y2=1.515
r69 34 36 36.2796 $w=3.72e-07 $l=2.8e-07 $layer=POLY_cond $X=0.985 $Y=1.557
+ $X2=1.265 $Y2=1.557
r70 33 34 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=0.96 $Y=1.557
+ $X2=0.985 $Y2=1.557
r71 31 33 48.5887 $w=3.72e-07 $l=3.75e-07 $layer=POLY_cond $X=0.585 $Y=1.557
+ $X2=0.96 $Y2=1.557
r72 31 32 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=0.585
+ $Y=1.515 $X2=0.585 $Y2=1.515
r73 29 31 9.71774 $w=3.72e-07 $l=7.5e-08 $layer=POLY_cond $X=0.51 $Y=1.557
+ $X2=0.585 $Y2=1.557
r74 28 29 1.94355 $w=3.72e-07 $l=1.5e-08 $layer=POLY_cond $X=0.495 $Y=1.557
+ $X2=0.51 $Y2=1.557
r75 24 37 1.74206 $w=4.28e-07 $l=6.5e-08 $layer=LI1_cond $X=1.2 $Y=1.565
+ $X2=1.265 $Y2=1.565
r76 23 24 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=0.72 $Y=1.565
+ $X2=1.2 $Y2=1.565
r77 23 32 3.61813 $w=4.28e-07 $l=1.35e-07 $layer=LI1_cond $X=0.72 $Y=1.565
+ $X2=0.585 $Y2=1.565
r78 22 32 9.24634 $w=4.28e-07 $l=3.45e-07 $layer=LI1_cond $X=0.24 $Y=1.565
+ $X2=0.585 $Y2=1.565
r79 18 39 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.415 $Y=1.35
+ $X2=1.415 $Y2=1.557
r80 18 20 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.415 $Y=1.35
+ $X2=1.415 $Y2=0.74
r81 15 38 24.0971 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=1.41 $Y=1.765
+ $X2=1.41 $Y2=1.557
r82 15 17 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.41 $Y=1.765
+ $X2=1.41 $Y2=2.4
r83 11 34 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.985 $Y=1.35
+ $X2=0.985 $Y2=1.557
r84 11 13 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=0.985 $Y=1.35
+ $X2=0.985 $Y2=0.74
r85 8 33 24.0971 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=0.96 $Y=1.765
+ $X2=0.96 $Y2=1.557
r86 8 10 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.96 $Y=1.765
+ $X2=0.96 $Y2=2.4
r87 5 29 24.0971 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=0.51 $Y=1.765
+ $X2=0.51 $Y2=1.557
r88 5 7 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.51 $Y=1.765
+ $X2=0.51 $Y2=2.4
r89 1 28 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.495 $Y=1.35
+ $X2=0.495 $Y2=1.557
r90 1 3 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=0.495 $Y=1.35
+ $X2=0.495 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HS__BUFINV_16%A_27_74# 1 2 3 4 15 17 19 22 24 26 29 31
+ 33 36 38 40 43 45 47 48 49 52 55 56 58 59 62 64 66 68 69 70 74 78 80 82 85 91
+ 97 98 99
c201 38 0 1.61688e-19 $X=3.23 $Y=1.765
c202 15 0 1.71373e-19 $X=1.845 $Y=0.74
r203 112 113 5.56154 $w=3.9e-07 $l=4.5e-08 $layer=POLY_cond $X=3.635 $Y=1.532
+ $X2=3.68 $Y2=1.532
r204 109 110 11.741 $w=3.9e-07 $l=9.5e-08 $layer=POLY_cond $X=3.135 $Y=1.532
+ $X2=3.23 $Y2=1.532
r205 108 109 43.8744 $w=3.9e-07 $l=3.55e-07 $layer=POLY_cond $X=2.78 $Y=1.532
+ $X2=3.135 $Y2=1.532
r206 107 108 9.26923 $w=3.9e-07 $l=7.5e-08 $layer=POLY_cond $X=2.705 $Y=1.532
+ $X2=2.78 $Y2=1.532
r207 106 107 46.3462 $w=3.9e-07 $l=3.75e-07 $layer=POLY_cond $X=2.33 $Y=1.532
+ $X2=2.705 $Y2=1.532
r208 105 106 6.79744 $w=3.9e-07 $l=5.5e-08 $layer=POLY_cond $X=2.275 $Y=1.532
+ $X2=2.33 $Y2=1.532
r209 102 103 1.85385 $w=3.9e-07 $l=1.5e-08 $layer=POLY_cond $X=1.845 $Y=1.532
+ $X2=1.86 $Y2=1.532
r210 92 112 42.0205 $w=3.9e-07 $l=3.4e-07 $layer=POLY_cond $X=3.295 $Y=1.532
+ $X2=3.635 $Y2=1.532
r211 92 110 8.03333 $w=3.9e-07 $l=6.5e-08 $layer=POLY_cond $X=3.295 $Y=1.532
+ $X2=3.23 $Y2=1.532
r212 91 92 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=3.295
+ $Y=1.465 $X2=3.295 $Y2=1.465
r213 89 105 42.0205 $w=3.9e-07 $l=3.4e-07 $layer=POLY_cond $X=1.935 $Y=1.532
+ $X2=2.275 $Y2=1.532
r214 89 103 9.26923 $w=3.9e-07 $l=7.5e-08 $layer=POLY_cond $X=1.935 $Y=1.532
+ $X2=1.86 $Y2=1.532
r215 88 91 47.4946 $w=3.28e-07 $l=1.36e-06 $layer=LI1_cond $X=1.935 $Y=1.465
+ $X2=3.295 $Y2=1.465
r216 88 89 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=1.935
+ $Y=1.465 $X2=1.935 $Y2=1.465
r217 86 99 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=1.685 $Y=1.465
+ $X2=1.685 $Y2=1.095
r218 86 88 5.76222 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=1.77 $Y=1.465
+ $X2=1.935 $Y2=1.465
r219 84 86 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=1.685 $Y=1.63
+ $X2=1.685 $Y2=1.465
r220 84 85 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=1.685 $Y=1.63
+ $X2=1.685 $Y2=1.95
r221 83 97 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.35 $Y=2.035
+ $X2=1.185 $Y2=2.035
r222 82 85 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.6 $Y=2.035
+ $X2=1.685 $Y2=1.95
r223 82 83 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=1.6 $Y=2.035
+ $X2=1.35 $Y2=2.035
r224 81 98 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.285 $Y=1.095
+ $X2=1.2 $Y2=1.095
r225 80 99 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.6 $Y=1.095
+ $X2=1.685 $Y2=1.095
r226 80 81 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=1.6 $Y=1.095
+ $X2=1.285 $Y2=1.095
r227 76 98 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.2 $Y=1.01 $X2=1.2
+ $Y2=1.095
r228 76 78 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=1.2 $Y=1.01
+ $X2=1.2 $Y2=0.515
r229 72 97 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.185 $Y=2.12
+ $X2=1.185 $Y2=2.035
r230 72 74 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=1.185 $Y=2.12
+ $X2=1.185 $Y2=2.815
r231 71 95 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.45 $Y=2.035
+ $X2=0.285 $Y2=2.035
r232 70 97 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.02 $Y=2.035
+ $X2=1.185 $Y2=2.035
r233 70 71 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=1.02 $Y=2.035
+ $X2=0.45 $Y2=2.035
r234 68 98 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.115 $Y=1.095
+ $X2=1.2 $Y2=1.095
r235 68 69 48.9305 $w=1.68e-07 $l=7.5e-07 $layer=LI1_cond $X=1.115 $Y=1.095
+ $X2=0.365 $Y2=1.095
r236 64 95 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.285 $Y=2.12
+ $X2=0.285 $Y2=2.035
r237 64 66 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=0.285 $Y=2.12
+ $X2=0.285 $Y2=2.815
r238 60 69 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.24 $Y=1.01
+ $X2=0.365 $Y2=1.095
r239 60 62 22.8184 $w=2.48e-07 $l=4.95e-07 $layer=LI1_cond $X=0.24 $Y=1.01
+ $X2=0.24 $Y2=0.515
r240 56 58 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=4.13 $Y=1.765
+ $X2=4.13 $Y2=2.4
r241 55 56 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=4.13 $Y=1.675
+ $X2=4.13 $Y2=1.765
r242 54 59 18.8402 $w=1.65e-07 $l=8.66025e-08 $layer=POLY_cond $X=4.13 $Y=1.45
+ $X2=4.105 $Y2=1.375
r243 54 55 87.4597 $w=1.8e-07 $l=2.25e-07 $layer=POLY_cond $X=4.13 $Y=1.45
+ $X2=4.13 $Y2=1.675
r244 50 59 18.8402 $w=1.65e-07 $l=9.28709e-08 $layer=POLY_cond $X=4.065 $Y=1.3
+ $X2=4.105 $Y2=1.375
r245 50 52 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=4.065 $Y=1.3
+ $X2=4.065 $Y2=0.74
r246 49 113 30.126 $w=3.9e-07 $l=1.96924e-07 $layer=POLY_cond $X=3.77 $Y=1.375
+ $X2=3.68 $Y2=1.532
r247 48 59 6.66866 $w=1.5e-07 $l=1.15e-07 $layer=POLY_cond $X=3.99 $Y=1.375
+ $X2=4.105 $Y2=1.375
r248 48 49 112.809 $w=1.5e-07 $l=2.2e-07 $layer=POLY_cond $X=3.99 $Y=1.375
+ $X2=3.77 $Y2=1.375
r249 45 113 25.2441 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=3.68 $Y=1.765
+ $X2=3.68 $Y2=1.532
r250 45 47 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.68 $Y=1.765
+ $X2=3.68 $Y2=2.4
r251 41 112 25.2441 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=3.635 $Y=1.3
+ $X2=3.635 $Y2=1.532
r252 41 43 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=3.635 $Y=1.3
+ $X2=3.635 $Y2=0.74
r253 38 110 25.2441 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=3.23 $Y=1.765
+ $X2=3.23 $Y2=1.532
r254 38 40 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.23 $Y=1.765
+ $X2=3.23 $Y2=2.4
r255 34 109 25.2441 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=3.135 $Y=1.3
+ $X2=3.135 $Y2=1.532
r256 34 36 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=3.135 $Y=1.3
+ $X2=3.135 $Y2=0.74
r257 31 108 25.2441 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=2.78 $Y=1.765
+ $X2=2.78 $Y2=1.532
r258 31 33 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.78 $Y=1.765
+ $X2=2.78 $Y2=2.4
r259 27 107 25.2441 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=2.705 $Y=1.3
+ $X2=2.705 $Y2=1.532
r260 27 29 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=2.705 $Y=1.3
+ $X2=2.705 $Y2=0.74
r261 24 106 25.2441 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=2.33 $Y=1.765
+ $X2=2.33 $Y2=1.532
r262 24 26 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.33 $Y=1.765
+ $X2=2.33 $Y2=2.4
r263 20 105 25.2441 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=2.275 $Y=1.3
+ $X2=2.275 $Y2=1.532
r264 20 22 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=2.275 $Y=1.3
+ $X2=2.275 $Y2=0.74
r265 17 103 25.2441 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=1.86 $Y=1.765
+ $X2=1.86 $Y2=1.532
r266 17 19 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.86 $Y=1.765
+ $X2=1.86 $Y2=2.4
r267 13 102 25.2441 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=1.845 $Y=1.3
+ $X2=1.845 $Y2=1.532
r268 13 15 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=1.845 $Y=1.3
+ $X2=1.845 $Y2=0.74
r269 4 97 400 $w=1.7e-07 $l=3.4187e-07 $layer=licon1_PDIFF $count=1 $X=1.035
+ $Y=1.84 $X2=1.185 $Y2=2.115
r270 4 74 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=1.035
+ $Y=1.84 $X2=1.185 $Y2=2.815
r271 3 95 400 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_PDIFF $count=1 $X=0.14
+ $Y=1.84 $X2=0.285 $Y2=2.115
r272 3 66 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=0.14
+ $Y=1.84 $X2=0.285 $Y2=2.815
r273 2 78 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.06
+ $Y=0.37 $X2=1.2 $Y2=0.515
r274 1 62 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__BUFINV_16%A_384_74# 1 2 3 4 5 6 21 23 25 28 30 32 35
+ 37 39 42 44 46 49 51 53 56 58 60 61 63 66 70 72 74 75 77 80 82 84 87 89 91 94
+ 98 100 102 105 107 109 112 114 116 117 119 122 126 128 130 133 139 141 142 143
+ 144 147 151 155 157 161 163 165 169 170 194 203 210 217 224 231 238 245 248
c456 163 0 1.61688e-19 $X=3.905 $Y=1.97
c457 142 0 1.71373e-19 $X=2.145 $Y=1.045
r458 248 249 5.64844 $w=3.84e-07 $l=4.5e-08 $layer=POLY_cond $X=11.435 $Y=1.532
+ $X2=11.48 $Y2=1.532
r459 247 248 53.974 $w=3.84e-07 $l=4.3e-07 $layer=POLY_cond $X=11.005 $Y=1.532
+ $X2=11.435 $Y2=1.532
r460 246 247 1.88281 $w=3.84e-07 $l=1.5e-08 $layer=POLY_cond $X=10.99 $Y=1.532
+ $X2=11.005 $Y2=1.532
r461 244 246 35.1458 $w=3.84e-07 $l=2.8e-07 $layer=POLY_cond $X=10.71 $Y=1.532
+ $X2=10.99 $Y2=1.532
r462 244 245 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.71
+ $Y=1.465 $X2=10.71 $Y2=1.465
r463 242 244 22.5938 $w=3.84e-07 $l=1.8e-07 $layer=POLY_cond $X=10.53 $Y=1.532
+ $X2=10.71 $Y2=1.532
r464 241 242 3.13802 $w=3.84e-07 $l=2.5e-08 $layer=POLY_cond $X=10.505 $Y=1.532
+ $X2=10.53 $Y2=1.532
r465 240 241 53.3464 $w=3.84e-07 $l=4.25e-07 $layer=POLY_cond $X=10.08 $Y=1.532
+ $X2=10.505 $Y2=1.532
r466 239 240 0.627604 $w=3.84e-07 $l=5e-09 $layer=POLY_cond $X=10.075 $Y=1.532
+ $X2=10.08 $Y2=1.532
r467 237 239 37.0286 $w=3.84e-07 $l=2.95e-07 $layer=POLY_cond $X=9.78 $Y=1.532
+ $X2=10.075 $Y2=1.532
r468 237 238 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.78
+ $Y=1.465 $X2=9.78 $Y2=1.465
r469 235 237 25.1042 $w=3.84e-07 $l=2e-07 $layer=POLY_cond $X=9.58 $Y=1.532
+ $X2=9.78 $Y2=1.532
r470 234 235 0.627604 $w=3.84e-07 $l=5e-09 $layer=POLY_cond $X=9.575 $Y=1.532
+ $X2=9.58 $Y2=1.532
r471 233 234 53.974 $w=3.84e-07 $l=4.3e-07 $layer=POLY_cond $X=9.145 $Y=1.532
+ $X2=9.575 $Y2=1.532
r472 232 233 1.88281 $w=3.84e-07 $l=1.5e-08 $layer=POLY_cond $X=9.13 $Y=1.532
+ $X2=9.145 $Y2=1.532
r473 230 232 35.1458 $w=3.84e-07 $l=2.8e-07 $layer=POLY_cond $X=8.85 $Y=1.532
+ $X2=9.13 $Y2=1.532
r474 230 231 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.85
+ $Y=1.465 $X2=8.85 $Y2=1.465
r475 228 230 25.7318 $w=3.84e-07 $l=2.05e-07 $layer=POLY_cond $X=8.645 $Y=1.532
+ $X2=8.85 $Y2=1.532
r476 227 228 1.88281 $w=3.84e-07 $l=1.5e-08 $layer=POLY_cond $X=8.63 $Y=1.532
+ $X2=8.645 $Y2=1.532
r477 226 227 52.0911 $w=3.84e-07 $l=4.15e-07 $layer=POLY_cond $X=8.215 $Y=1.532
+ $X2=8.63 $Y2=1.532
r478 225 226 4.39323 $w=3.84e-07 $l=3.5e-08 $layer=POLY_cond $X=8.18 $Y=1.532
+ $X2=8.215 $Y2=1.532
r479 223 225 32.0078 $w=3.84e-07 $l=2.55e-07 $layer=POLY_cond $X=7.925 $Y=1.532
+ $X2=8.18 $Y2=1.532
r480 223 224 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.925
+ $Y=1.465 $X2=7.925 $Y2=1.465
r481 221 223 24.4766 $w=3.84e-07 $l=1.95e-07 $layer=POLY_cond $X=7.73 $Y=1.532
+ $X2=7.925 $Y2=1.532
r482 220 221 1.88281 $w=3.84e-07 $l=1.5e-08 $layer=POLY_cond $X=7.715 $Y=1.532
+ $X2=7.73 $Y2=1.532
r483 219 220 53.974 $w=3.84e-07 $l=4.3e-07 $layer=POLY_cond $X=7.285 $Y=1.532
+ $X2=7.715 $Y2=1.532
r484 218 219 0.627604 $w=3.84e-07 $l=5e-09 $layer=POLY_cond $X=7.28 $Y=1.532
+ $X2=7.285 $Y2=1.532
r485 216 218 34.5182 $w=3.84e-07 $l=2.75e-07 $layer=POLY_cond $X=7.005 $Y=1.532
+ $X2=7.28 $Y2=1.532
r486 216 217 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.005
+ $Y=1.465 $X2=7.005 $Y2=1.465
r487 214 216 21.9661 $w=3.84e-07 $l=1.75e-07 $layer=POLY_cond $X=6.83 $Y=1.532
+ $X2=7.005 $Y2=1.532
r488 213 214 5.64844 $w=3.84e-07 $l=4.5e-08 $layer=POLY_cond $X=6.785 $Y=1.532
+ $X2=6.83 $Y2=1.532
r489 212 213 50.8359 $w=3.84e-07 $l=4.05e-07 $layer=POLY_cond $X=6.38 $Y=1.532
+ $X2=6.785 $Y2=1.532
r490 211 212 3.13802 $w=3.84e-07 $l=2.5e-08 $layer=POLY_cond $X=6.355 $Y=1.532
+ $X2=6.38 $Y2=1.532
r491 209 211 36.401 $w=3.84e-07 $l=2.9e-07 $layer=POLY_cond $X=6.065 $Y=1.532
+ $X2=6.355 $Y2=1.532
r492 209 210 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.065
+ $Y=1.465 $X2=6.065 $Y2=1.465
r493 207 209 16.9453 $w=3.84e-07 $l=1.35e-07 $layer=POLY_cond $X=5.93 $Y=1.532
+ $X2=6.065 $Y2=1.532
r494 206 207 9.41406 $w=3.84e-07 $l=7.5e-08 $layer=POLY_cond $X=5.855 $Y=1.532
+ $X2=5.93 $Y2=1.532
r495 205 206 47.0703 $w=3.84e-07 $l=3.75e-07 $layer=POLY_cond $X=5.48 $Y=1.532
+ $X2=5.855 $Y2=1.532
r496 204 205 6.90365 $w=3.84e-07 $l=5.5e-08 $layer=POLY_cond $X=5.425 $Y=1.532
+ $X2=5.48 $Y2=1.532
r497 202 204 31.3802 $w=3.84e-07 $l=2.5e-07 $layer=POLY_cond $X=5.175 $Y=1.532
+ $X2=5.425 $Y2=1.532
r498 202 203 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.175
+ $Y=1.465 $X2=5.175 $Y2=1.465
r499 200 202 18.2005 $w=3.84e-07 $l=1.45e-07 $layer=POLY_cond $X=5.03 $Y=1.532
+ $X2=5.175 $Y2=1.532
r500 199 200 4.39323 $w=3.84e-07 $l=3.5e-08 $layer=POLY_cond $X=4.995 $Y=1.532
+ $X2=5.03 $Y2=1.532
r501 198 199 52.0911 $w=3.84e-07 $l=4.15e-07 $layer=POLY_cond $X=4.58 $Y=1.532
+ $X2=4.995 $Y2=1.532
r502 197 198 1.88281 $w=3.84e-07 $l=1.5e-08 $layer=POLY_cond $X=4.565 $Y=1.532
+ $X2=4.58 $Y2=1.532
r503 195 245 6.9845 $w=3.28e-07 $l=2e-07 $layer=LI1_cond $X=10.71 $Y=1.665
+ $X2=10.71 $Y2=1.465
r504 194 195 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.71 $Y=1.665
+ $X2=10.71 $Y2=1.665
r505 192 238 6.9845 $w=3.28e-07 $l=2e-07 $layer=LI1_cond $X=9.78 $Y=1.665
+ $X2=9.78 $Y2=1.465
r506 191 194 0.5999 $w=2.3e-07 $l=9.35e-07 $layer=MET1_cond $X=9.775 $Y=1.665
+ $X2=10.71 $Y2=1.665
r507 191 192 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.775 $Y=1.665
+ $X2=9.775 $Y2=1.665
r508 189 231 6.9845 $w=3.28e-07 $l=2e-07 $layer=LI1_cond $X=8.85 $Y=1.665
+ $X2=8.85 $Y2=1.465
r509 188 191 0.593484 $w=2.3e-07 $l=9.25e-07 $layer=MET1_cond $X=8.85 $Y=1.665
+ $X2=9.775 $Y2=1.665
r510 188 189 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.85 $Y=1.665
+ $X2=8.85 $Y2=1.665
r511 186 224 6.9845 $w=3.28e-07 $l=2e-07 $layer=LI1_cond $X=7.925 $Y=1.665
+ $X2=7.925 $Y2=1.465
r512 185 188 0.596692 $w=2.3e-07 $l=9.3e-07 $layer=MET1_cond $X=7.92 $Y=1.665
+ $X2=8.85 $Y2=1.665
r513 185 186 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=1.665
+ $X2=7.92 $Y2=1.665
r514 183 217 6.9845 $w=3.28e-07 $l=2e-07 $layer=LI1_cond $X=7.005 $Y=1.665
+ $X2=7.005 $Y2=1.465
r515 182 185 0.587068 $w=2.3e-07 $l=9.15e-07 $layer=MET1_cond $X=7.005 $Y=1.665
+ $X2=7.92 $Y2=1.665
r516 182 183 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.005 $Y=1.665
+ $X2=7.005 $Y2=1.665
r517 180 210 6.9845 $w=3.28e-07 $l=2e-07 $layer=LI1_cond $X=6.065 $Y=1.665
+ $X2=6.065 $Y2=1.465
r518 179 182 0.603108 $w=2.3e-07 $l=9.4e-07 $layer=MET1_cond $X=6.065 $Y=1.665
+ $X2=7.005 $Y2=1.665
r519 179 180 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.065 $Y=1.665
+ $X2=6.065 $Y2=1.665
r520 177 203 8.53661 $w=2.68e-07 $l=2e-07 $layer=LI1_cond $X=5.17 $Y=1.665
+ $X2=5.17 $Y2=1.465
r521 176 179 0.571028 $w=2.3e-07 $l=8.9e-07 $layer=MET1_cond $X=5.175 $Y=1.665
+ $X2=6.065 $Y2=1.665
r522 176 177 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.175 $Y=1.665
+ $X2=5.175 $Y2=1.665
r523 173 280 5.77204 $w=4.65e-07 $l=2.2e-07 $layer=LI1_cond $X=4.06 $Y=1.665
+ $X2=4.06 $Y2=1.885
r524 172 176 0.554988 $w=2.3e-07 $l=8.65e-07 $layer=MET1_cond $X=4.31 $Y=1.665
+ $X2=5.175 $Y2=1.665
r525 172 173 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.31 $Y=1.665
+ $X2=4.31 $Y2=1.665
r526 165 167 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=3.905 $Y=1.985
+ $X2=3.905 $Y2=2.815
r527 163 280 3.27514 $w=4.65e-07 $l=1.92873e-07 $layer=LI1_cond $X=3.905 $Y=1.97
+ $X2=4.06 $Y2=1.885
r528 163 165 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=3.905 $Y=1.97
+ $X2=3.905 $Y2=1.985
r529 159 161 20.5135 $w=2.48e-07 $l=4.45e-07 $layer=LI1_cond $X=3.81 $Y=0.96
+ $X2=3.81 $Y2=0.515
r530 158 170 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.17 $Y=1.885
+ $X2=3.005 $Y2=1.885
r531 157 280 6.7035 $w=1.7e-07 $l=3.2e-07 $layer=LI1_cond $X=3.74 $Y=1.885
+ $X2=4.06 $Y2=1.885
r532 157 158 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=3.74 $Y=1.885
+ $X2=3.17 $Y2=1.885
r533 156 169 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.005 $Y=1.045
+ $X2=2.88 $Y2=1.045
r534 155 173 16.2667 $w=4.65e-07 $l=7.8543e-07 $layer=LI1_cond $X=3.685 $Y=1.045
+ $X2=4.06 $Y2=1.665
r535 155 159 4.82172 $w=4.65e-07 $l=1.62019e-07 $layer=LI1_cond $X=3.685
+ $Y=1.045 $X2=3.81 $Y2=0.96
r536 155 156 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=3.685 $Y=1.045
+ $X2=3.005 $Y2=1.045
r537 151 153 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=3.005 $Y=1.985
+ $X2=3.005 $Y2=2.815
r538 149 170 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.005 $Y=1.97
+ $X2=3.005 $Y2=1.885
r539 149 151 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=3.005 $Y=1.97
+ $X2=3.005 $Y2=1.985
r540 145 169 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.88 $Y=0.96
+ $X2=2.88 $Y2=1.045
r541 145 147 20.5135 $w=2.48e-07 $l=4.45e-07 $layer=LI1_cond $X=2.88 $Y=0.96
+ $X2=2.88 $Y2=0.515
r542 143 170 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.84 $Y=1.885
+ $X2=3.005 $Y2=1.885
r543 143 144 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=2.84 $Y=1.885
+ $X2=2.27 $Y2=1.885
r544 141 169 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.755 $Y=1.045
+ $X2=2.88 $Y2=1.045
r545 141 142 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=2.755 $Y=1.045
+ $X2=2.145 $Y2=1.045
r546 137 142 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.06 $Y=0.96
+ $X2=2.145 $Y2=1.045
r547 137 139 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=2.06 $Y=0.96
+ $X2=2.06 $Y2=0.515
r548 133 135 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=2.105 $Y=1.985
+ $X2=2.105 $Y2=2.815
r549 131 144 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.105 $Y=1.97
+ $X2=2.27 $Y2=1.885
r550 131 133 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=2.105 $Y=1.97
+ $X2=2.105 $Y2=1.985
r551 128 249 24.8669 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=11.48 $Y=1.765
+ $X2=11.48 $Y2=1.532
r552 128 130 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=11.48 $Y=1.765
+ $X2=11.48 $Y2=2.4
r553 124 248 24.8669 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=11.435 $Y=1.3
+ $X2=11.435 $Y2=1.532
r554 124 126 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=11.435 $Y=1.3
+ $X2=11.435 $Y2=0.74
r555 120 247 24.8669 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=11.005 $Y=1.3
+ $X2=11.005 $Y2=1.532
r556 120 122 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=11.005 $Y=1.3
+ $X2=11.005 $Y2=0.74
r557 117 246 24.8669 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=10.99 $Y=1.765
+ $X2=10.99 $Y2=1.532
r558 117 119 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=10.99 $Y=1.765
+ $X2=10.99 $Y2=2.4
r559 114 242 24.8669 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=10.53 $Y=1.765
+ $X2=10.53 $Y2=1.532
r560 114 116 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=10.53 $Y=1.765
+ $X2=10.53 $Y2=2.4
r561 110 241 24.8669 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=10.505 $Y=1.3
+ $X2=10.505 $Y2=1.532
r562 110 112 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=10.505 $Y=1.3
+ $X2=10.505 $Y2=0.74
r563 107 240 24.8669 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=10.08 $Y=1.765
+ $X2=10.08 $Y2=1.532
r564 107 109 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=10.08 $Y=1.765
+ $X2=10.08 $Y2=2.4
r565 103 239 24.8669 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=10.075 $Y=1.3
+ $X2=10.075 $Y2=1.532
r566 103 105 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=10.075 $Y=1.3
+ $X2=10.075 $Y2=0.74
r567 100 235 24.8669 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=9.58 $Y=1.765
+ $X2=9.58 $Y2=1.532
r568 100 102 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=9.58 $Y=1.765
+ $X2=9.58 $Y2=2.4
r569 96 234 24.8669 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=9.575 $Y=1.3
+ $X2=9.575 $Y2=1.532
r570 96 98 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=9.575 $Y=1.3
+ $X2=9.575 $Y2=0.74
r571 92 233 24.8669 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=9.145 $Y=1.3
+ $X2=9.145 $Y2=1.532
r572 92 94 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=9.145 $Y=1.3
+ $X2=9.145 $Y2=0.74
r573 89 232 24.8669 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=9.13 $Y=1.765
+ $X2=9.13 $Y2=1.532
r574 89 91 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=9.13 $Y=1.765
+ $X2=9.13 $Y2=2.4
r575 85 228 24.8669 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=8.645 $Y=1.3
+ $X2=8.645 $Y2=1.532
r576 85 87 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=8.645 $Y=1.3
+ $X2=8.645 $Y2=0.74
r577 82 227 24.8669 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=8.63 $Y=1.765
+ $X2=8.63 $Y2=1.532
r578 82 84 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=8.63 $Y=1.765
+ $X2=8.63 $Y2=2.4
r579 78 226 24.8669 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=8.215 $Y=1.3
+ $X2=8.215 $Y2=1.532
r580 78 80 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=8.215 $Y=1.3
+ $X2=8.215 $Y2=0.74
r581 75 225 24.8669 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=8.18 $Y=1.765
+ $X2=8.18 $Y2=1.532
r582 75 77 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=8.18 $Y=1.765
+ $X2=8.18 $Y2=2.4
r583 72 221 24.8669 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=7.73 $Y=1.765
+ $X2=7.73 $Y2=1.532
r584 72 74 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=7.73 $Y=1.765
+ $X2=7.73 $Y2=2.4
r585 68 220 24.8669 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=7.715 $Y=1.3
+ $X2=7.715 $Y2=1.532
r586 68 70 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=7.715 $Y=1.3
+ $X2=7.715 $Y2=0.74
r587 64 219 24.8669 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=7.285 $Y=1.3
+ $X2=7.285 $Y2=1.532
r588 64 66 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=7.285 $Y=1.3
+ $X2=7.285 $Y2=0.74
r589 61 218 24.8669 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=7.28 $Y=1.765
+ $X2=7.28 $Y2=1.532
r590 61 63 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=7.28 $Y=1.765
+ $X2=7.28 $Y2=2.4
r591 58 214 24.8669 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=6.83 $Y=1.765
+ $X2=6.83 $Y2=1.532
r592 58 60 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=6.83 $Y=1.765
+ $X2=6.83 $Y2=2.4
r593 54 213 24.8669 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=6.785 $Y=1.3
+ $X2=6.785 $Y2=1.532
r594 54 56 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=6.785 $Y=1.3
+ $X2=6.785 $Y2=0.74
r595 51 212 24.8669 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=6.38 $Y=1.765
+ $X2=6.38 $Y2=1.532
r596 51 53 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=6.38 $Y=1.765
+ $X2=6.38 $Y2=2.4
r597 47 211 24.8669 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=6.355 $Y=1.3
+ $X2=6.355 $Y2=1.532
r598 47 49 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=6.355 $Y=1.3
+ $X2=6.355 $Y2=0.74
r599 44 207 24.8669 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=5.93 $Y=1.765
+ $X2=5.93 $Y2=1.532
r600 44 46 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=5.93 $Y=1.765
+ $X2=5.93 $Y2=2.4
r601 40 206 24.8669 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=5.855 $Y=1.3
+ $X2=5.855 $Y2=1.532
r602 40 42 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=5.855 $Y=1.3
+ $X2=5.855 $Y2=0.74
r603 37 205 24.8669 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=5.48 $Y=1.765
+ $X2=5.48 $Y2=1.532
r604 37 39 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=5.48 $Y=1.765
+ $X2=5.48 $Y2=2.4
r605 33 204 24.8669 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=5.425 $Y=1.3
+ $X2=5.425 $Y2=1.532
r606 33 35 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=5.425 $Y=1.3
+ $X2=5.425 $Y2=0.74
r607 30 200 24.8669 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=5.03 $Y=1.765
+ $X2=5.03 $Y2=1.532
r608 30 32 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=5.03 $Y=1.765
+ $X2=5.03 $Y2=2.4
r609 26 199 24.8669 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=4.995 $Y=1.3
+ $X2=4.995 $Y2=1.532
r610 26 28 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=4.995 $Y=1.3
+ $X2=4.995 $Y2=0.74
r611 23 198 24.8669 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=4.58 $Y=1.765
+ $X2=4.58 $Y2=1.532
r612 23 25 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=4.58 $Y=1.765
+ $X2=4.58 $Y2=2.4
r613 19 197 24.8669 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=4.565 $Y=1.3
+ $X2=4.565 $Y2=1.532
r614 19 21 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=4.565 $Y=1.3
+ $X2=4.565 $Y2=0.74
r615 6 167 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=3.755
+ $Y=1.84 $X2=3.905 $Y2=2.815
r616 6 165 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=3.755
+ $Y=1.84 $X2=3.905 $Y2=1.985
r617 5 153 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=2.855
+ $Y=1.84 $X2=3.005 $Y2=2.815
r618 5 151 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=2.855
+ $Y=1.84 $X2=3.005 $Y2=1.985
r619 4 135 400 $w=1.7e-07 $l=1.05659e-06 $layer=licon1_PDIFF $count=1 $X=1.935
+ $Y=1.84 $X2=2.105 $Y2=2.815
r620 4 133 400 $w=1.7e-07 $l=2.31409e-07 $layer=licon1_PDIFF $count=1 $X=1.935
+ $Y=1.84 $X2=2.105 $Y2=1.985
r621 3 161 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.71
+ $Y=0.37 $X2=3.85 $Y2=0.515
r622 2 147 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.78
+ $Y=0.37 $X2=2.92 $Y2=0.515
r623 1 139 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.92
+ $Y=0.37 $X2=2.06 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__BUFINV_16%VPWR 1 2 3 4 5 6 7 8 9 10 11 12 13 44 48
+ 52 56 60 66 72 78 82 86 92 98 104 108 110 115 116 118 119 121 122 124 125 127
+ 128 130 131 132 133 134 158 163 168 173 179 182 185 188 191 195
r223 194 195 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.76 $Y=3.33
+ $X2=11.76 $Y2=3.33
r224 191 192 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.8 $Y=3.33
+ $X2=10.8 $Y2=3.33
r225 188 189 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.84 $Y=3.33
+ $X2=9.84 $Y2=3.33
r226 185 186 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r227 182 183 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r228 179 180 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r229 177 195 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.28 $Y=3.33
+ $X2=11.76 $Y2=3.33
r230 177 192 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.28 $Y=3.33
+ $X2=10.8 $Y2=3.33
r231 176 177 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.28 $Y=3.33
+ $X2=11.28 $Y2=3.33
r232 174 191 6.25164 $w=1.7e-07 $l=1.08e-07 $layer=LI1_cond $X=10.885 $Y=3.33
+ $X2=10.777 $Y2=3.33
r233 174 176 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=10.885 $Y=3.33
+ $X2=11.28 $Y2=3.33
r234 173 194 3.99177 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=11.62 $Y=3.33
+ $X2=11.81 $Y2=3.33
r235 173 176 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=11.62 $Y=3.33
+ $X2=11.28 $Y2=3.33
r236 172 192 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.32 $Y=3.33
+ $X2=10.8 $Y2=3.33
r237 172 189 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.32 $Y=3.33
+ $X2=9.84 $Y2=3.33
r238 171 172 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.32 $Y=3.33
+ $X2=10.32 $Y2=3.33
r239 169 188 6.70225 $w=1.7e-07 $l=1.18e-07 $layer=LI1_cond $X=9.955 $Y=3.33
+ $X2=9.837 $Y2=3.33
r240 169 171 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=9.955 $Y=3.33
+ $X2=10.32 $Y2=3.33
r241 168 191 6.25164 $w=1.7e-07 $l=1.07e-07 $layer=LI1_cond $X=10.67 $Y=3.33
+ $X2=10.777 $Y2=3.33
r242 168 171 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=10.67 $Y=3.33
+ $X2=10.32 $Y2=3.33
r243 167 189 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.36 $Y=3.33
+ $X2=9.84 $Y2=3.33
r244 167 186 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.36 $Y=3.33
+ $X2=8.88 $Y2=3.33
r245 166 167 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.36 $Y=3.33
+ $X2=9.36 $Y2=3.33
r246 164 185 6.47928 $w=1.7e-07 $l=1.13e-07 $layer=LI1_cond $X=8.995 $Y=3.33
+ $X2=8.882 $Y2=3.33
r247 164 166 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=8.995 $Y=3.33
+ $X2=9.36 $Y2=3.33
r248 163 188 6.70225 $w=1.7e-07 $l=1.17e-07 $layer=LI1_cond $X=9.72 $Y=3.33
+ $X2=9.837 $Y2=3.33
r249 163 166 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=9.72 $Y=3.33
+ $X2=9.36 $Y2=3.33
r250 162 186 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=3.33
+ $X2=8.88 $Y2=3.33
r251 162 183 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=3.33
+ $X2=7.92 $Y2=3.33
r252 161 162 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=3.33
+ $X2=8.4 $Y2=3.33
r253 159 182 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.04 $Y=3.33
+ $X2=7.955 $Y2=3.33
r254 159 161 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=8.04 $Y=3.33
+ $X2=8.4 $Y2=3.33
r255 158 185 6.47928 $w=1.7e-07 $l=1.12e-07 $layer=LI1_cond $X=8.77 $Y=3.33
+ $X2=8.882 $Y2=3.33
r256 158 161 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=8.77 $Y=3.33
+ $X2=8.4 $Y2=3.33
r257 157 183 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=7.92 $Y2=3.33
r258 156 157 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r259 150 151 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r260 148 151 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=5.04 $Y2=3.33
r261 147 148 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r262 145 148 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=4.08 $Y2=3.33
r263 144 145 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r264 142 145 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=3.12 $Y2=3.33
r265 141 142 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r266 139 142 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.16 $Y2=3.33
r267 139 180 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r268 138 139 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r269 136 179 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.82 $Y=3.33
+ $X2=0.735 $Y2=3.33
r270 136 138 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=0.82 $Y=3.33
+ $X2=1.2 $Y2=3.33
r271 134 157 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6 $Y=3.33
+ $X2=6.96 $Y2=3.33
r272 134 151 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6 $Y=3.33
+ $X2=5.04 $Y2=3.33
r273 134 153 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r274 132 156 0.652406 $w=1.68e-07 $l=1e-08 $layer=LI1_cond $X=6.97 $Y=3.33
+ $X2=6.96 $Y2=3.33
r275 132 133 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.97 $Y=3.33
+ $X2=7.055 $Y2=3.33
r276 130 153 4.56684 $w=1.68e-07 $l=7e-08 $layer=LI1_cond $X=6.07 $Y=3.33 $X2=6
+ $Y2=3.33
r277 130 131 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.07 $Y=3.33
+ $X2=6.155 $Y2=3.33
r278 129 156 46.9733 $w=1.68e-07 $l=7.2e-07 $layer=LI1_cond $X=6.24 $Y=3.33
+ $X2=6.96 $Y2=3.33
r279 129 131 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.24 $Y=3.33
+ $X2=6.155 $Y2=3.33
r280 127 150 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=5.17 $Y=3.33
+ $X2=5.04 $Y2=3.33
r281 127 128 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.17 $Y=3.33
+ $X2=5.255 $Y2=3.33
r282 126 153 43.0588 $w=1.68e-07 $l=6.6e-07 $layer=LI1_cond $X=5.34 $Y=3.33
+ $X2=6 $Y2=3.33
r283 126 128 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.34 $Y=3.33
+ $X2=5.255 $Y2=3.33
r284 124 147 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=4.27 $Y=3.33
+ $X2=4.08 $Y2=3.33
r285 124 125 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.27 $Y=3.33
+ $X2=4.355 $Y2=3.33
r286 123 150 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=4.44 $Y=3.33
+ $X2=5.04 $Y2=3.33
r287 123 125 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.44 $Y=3.33
+ $X2=4.355 $Y2=3.33
r288 121 144 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=3.37 $Y=3.33
+ $X2=3.12 $Y2=3.33
r289 121 122 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.37 $Y=3.33
+ $X2=3.455 $Y2=3.33
r290 120 147 35.2299 $w=1.68e-07 $l=5.4e-07 $layer=LI1_cond $X=3.54 $Y=3.33
+ $X2=4.08 $Y2=3.33
r291 120 122 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.54 $Y=3.33
+ $X2=3.455 $Y2=3.33
r292 118 141 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=2.47 $Y=3.33
+ $X2=2.16 $Y2=3.33
r293 118 119 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.47 $Y=3.33
+ $X2=2.555 $Y2=3.33
r294 117 144 31.3155 $w=1.68e-07 $l=4.8e-07 $layer=LI1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r295 117 119 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.64 $Y=3.33
+ $X2=2.555 $Y2=3.33
r296 115 138 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=1.55 $Y=3.33
+ $X2=1.2 $Y2=3.33
r297 115 116 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.55 $Y=3.33
+ $X2=1.635 $Y2=3.33
r298 114 141 28.7059 $w=1.68e-07 $l=4.4e-07 $layer=LI1_cond $X=1.72 $Y=3.33
+ $X2=2.16 $Y2=3.33
r299 114 116 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.72 $Y=3.33
+ $X2=1.635 $Y2=3.33
r300 110 113 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=11.745 $Y=1.985
+ $X2=11.745 $Y2=2.815
r301 108 194 3.1514 $w=2.5e-07 $l=1.12916e-07 $layer=LI1_cond $X=11.745 $Y=3.245
+ $X2=11.81 $Y2=3.33
r302 108 113 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=11.745 $Y=3.245
+ $X2=11.745 $Y2=2.815
r303 104 107 39.1295 $w=2.13e-07 $l=7.3e-07 $layer=LI1_cond $X=10.777 $Y=2.085
+ $X2=10.777 $Y2=2.815
r304 102 191 0.512231 $w=2.15e-07 $l=8.5e-08 $layer=LI1_cond $X=10.777 $Y=3.245
+ $X2=10.777 $Y2=3.33
r305 102 107 23.0489 $w=2.13e-07 $l=4.3e-07 $layer=LI1_cond $X=10.777 $Y=3.245
+ $X2=10.777 $Y2=2.815
r306 98 101 35.7993 $w=2.33e-07 $l=7.3e-07 $layer=LI1_cond $X=9.837 $Y=2.085
+ $X2=9.837 $Y2=2.815
r307 96 188 0.207053 $w=2.35e-07 $l=8.5e-08 $layer=LI1_cond $X=9.837 $Y=3.245
+ $X2=9.837 $Y2=3.33
r308 96 101 21.0873 $w=2.33e-07 $l=4.3e-07 $layer=LI1_cond $X=9.837 $Y=3.245
+ $X2=9.837 $Y2=2.815
r309 92 95 37.3904 $w=2.23e-07 $l=7.3e-07 $layer=LI1_cond $X=8.882 $Y=2.085
+ $X2=8.882 $Y2=2.815
r310 90 185 0.355529 $w=2.25e-07 $l=8.5e-08 $layer=LI1_cond $X=8.882 $Y=3.245
+ $X2=8.882 $Y2=3.33
r311 90 95 22.0245 $w=2.23e-07 $l=4.3e-07 $layer=LI1_cond $X=8.882 $Y=3.245
+ $X2=8.882 $Y2=2.815
r312 86 89 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=7.955 $Y=2.085
+ $X2=7.955 $Y2=2.815
r313 84 182 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.955 $Y=3.245
+ $X2=7.955 $Y2=3.33
r314 84 89 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=7.955 $Y=3.245
+ $X2=7.955 $Y2=2.815
r315 83 133 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.14 $Y=3.33
+ $X2=7.055 $Y2=3.33
r316 82 182 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.87 $Y=3.33
+ $X2=7.955 $Y2=3.33
r317 82 83 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=7.87 $Y=3.33
+ $X2=7.14 $Y2=3.33
r318 78 81 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=7.055 $Y=2.085
+ $X2=7.055 $Y2=2.815
r319 76 133 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.055 $Y=3.245
+ $X2=7.055 $Y2=3.33
r320 76 81 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=7.055 $Y=3.245
+ $X2=7.055 $Y2=2.815
r321 72 75 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=6.155 $Y=2.085
+ $X2=6.155 $Y2=2.815
r322 70 131 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.155 $Y=3.245
+ $X2=6.155 $Y2=3.33
r323 70 75 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=6.155 $Y=3.245
+ $X2=6.155 $Y2=2.815
r324 66 69 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=5.255 $Y=2.085
+ $X2=5.255 $Y2=2.815
r325 64 128 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.255 $Y=3.245
+ $X2=5.255 $Y2=3.33
r326 64 69 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=5.255 $Y=3.245
+ $X2=5.255 $Y2=2.815
r327 60 63 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=4.355 $Y=2.085
+ $X2=4.355 $Y2=2.815
r328 58 125 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.355 $Y=3.245
+ $X2=4.355 $Y2=3.33
r329 58 63 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=4.355 $Y=3.245
+ $X2=4.355 $Y2=2.815
r330 54 122 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.455 $Y=3.245
+ $X2=3.455 $Y2=3.33
r331 54 56 61.3262 $w=1.68e-07 $l=9.4e-07 $layer=LI1_cond $X=3.455 $Y=3.245
+ $X2=3.455 $Y2=2.305
r332 50 119 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.555 $Y=3.245
+ $X2=2.555 $Y2=3.33
r333 50 52 61.3262 $w=1.68e-07 $l=9.4e-07 $layer=LI1_cond $X=2.555 $Y=3.245
+ $X2=2.555 $Y2=2.305
r334 46 116 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.635 $Y=3.245
+ $X2=1.635 $Y2=3.33
r335 46 48 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=1.635 $Y=3.245
+ $X2=1.635 $Y2=2.455
r336 42 179 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.735 $Y=3.245
+ $X2=0.735 $Y2=3.33
r337 42 44 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=0.735 $Y=3.245
+ $X2=0.735 $Y2=2.455
r338 13 113 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=11.555
+ $Y=1.84 $X2=11.705 $Y2=2.815
r339 13 110 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=11.555
+ $Y=1.84 $X2=11.705 $Y2=1.985
r340 12 107 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=10.605
+ $Y=1.84 $X2=10.755 $Y2=2.815
r341 12 104 400 $w=1.7e-07 $l=3.11087e-07 $layer=licon1_PDIFF $count=1 $X=10.605
+ $Y=1.84 $X2=10.755 $Y2=2.085
r342 11 101 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=9.655
+ $Y=1.84 $X2=9.805 $Y2=2.815
r343 11 98 400 $w=1.7e-07 $l=3.11087e-07 $layer=licon1_PDIFF $count=1 $X=9.655
+ $Y=1.84 $X2=9.805 $Y2=2.085
r344 10 95 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=8.705
+ $Y=1.84 $X2=8.855 $Y2=2.815
r345 10 92 400 $w=1.7e-07 $l=3.11087e-07 $layer=licon1_PDIFF $count=1 $X=8.705
+ $Y=1.84 $X2=8.855 $Y2=2.085
r346 9 89 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=7.805
+ $Y=1.84 $X2=7.955 $Y2=2.815
r347 9 86 400 $w=1.7e-07 $l=3.11087e-07 $layer=licon1_PDIFF $count=1 $X=7.805
+ $Y=1.84 $X2=7.955 $Y2=2.085
r348 8 81 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=6.905
+ $Y=1.84 $X2=7.055 $Y2=2.815
r349 8 78 400 $w=1.7e-07 $l=3.11087e-07 $layer=licon1_PDIFF $count=1 $X=6.905
+ $Y=1.84 $X2=7.055 $Y2=2.085
r350 7 75 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=6.005
+ $Y=1.84 $X2=6.155 $Y2=2.815
r351 7 72 400 $w=1.7e-07 $l=3.11087e-07 $layer=licon1_PDIFF $count=1 $X=6.005
+ $Y=1.84 $X2=6.155 $Y2=2.085
r352 6 69 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=5.105
+ $Y=1.84 $X2=5.255 $Y2=2.815
r353 6 66 400 $w=1.7e-07 $l=3.11087e-07 $layer=licon1_PDIFF $count=1 $X=5.105
+ $Y=1.84 $X2=5.255 $Y2=2.085
r354 5 63 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=4.205
+ $Y=1.84 $X2=4.355 $Y2=2.815
r355 5 60 400 $w=1.7e-07 $l=3.11087e-07 $layer=licon1_PDIFF $count=1 $X=4.205
+ $Y=1.84 $X2=4.355 $Y2=2.085
r356 4 56 300 $w=1.7e-07 $l=5.34766e-07 $layer=licon1_PDIFF $count=2 $X=3.305
+ $Y=1.84 $X2=3.455 $Y2=2.305
r357 3 52 300 $w=1.7e-07 $l=5.34766e-07 $layer=licon1_PDIFF $count=2 $X=2.405
+ $Y=1.84 $X2=2.555 $Y2=2.305
r358 2 48 300 $w=1.7e-07 $l=6.85912e-07 $layer=licon1_PDIFF $count=2 $X=1.485
+ $Y=1.84 $X2=1.635 $Y2=2.455
r359 1 44 300 $w=1.7e-07 $l=6.85912e-07 $layer=licon1_PDIFF $count=2 $X=0.585
+ $Y=1.84 $X2=0.735 $Y2=2.455
.ends

.subckt PM_SKY130_FD_SC_HS__BUFINV_16%Y 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16
+ 51 55 59 63 67 69 71 75 77 79 83 87 91 95 100 105 110 115 118 121 127 133 139
+ 145 146 151
r262 160 162 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.355 $Y=2.035
+ $X2=9.355 $Y2=2.035
r263 158 162 0.609524 $w=2.3e-07 $l=9.5e-07 $layer=MET1_cond $X=8.405 $Y=2.035
+ $X2=9.355 $Y2=2.035
r264 156 158 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.405 $Y=2.035
+ $X2=8.405 $Y2=2.035
r265 151 154 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.505 $Y=2.035
+ $X2=7.505 $Y2=2.035
r266 151 152 3.7572 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=7.505 $Y=2.005
+ $X2=7.505 $Y2=1.92
r267 145 148 27.2396 $w=3.28e-07 $l=7.8e-07 $layer=LI1_cond $X=11.255 $Y=2.035
+ $X2=11.255 $Y2=2.815
r268 145 146 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.255 $Y=2.035
+ $X2=11.255 $Y2=2.035
r269 140 146 0.609524 $w=2.3e-07 $l=9.5e-07 $layer=MET1_cond $X=10.305 $Y=2.035
+ $X2=11.255 $Y2=2.035
r270 140 162 0.609524 $w=2.3e-07 $l=9.5e-07 $layer=MET1_cond $X=10.305 $Y=2.035
+ $X2=9.355 $Y2=2.035
r271 139 142 27.2396 $w=3.28e-07 $l=7.8e-07 $layer=LI1_cond $X=10.305 $Y=2.035
+ $X2=10.305 $Y2=2.815
r272 139 140 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.305 $Y=2.035
+ $X2=10.305 $Y2=2.035
r273 134 154 0.577444 $w=2.3e-07 $l=9e-07 $layer=MET1_cond $X=6.605 $Y=2.035
+ $X2=7.505 $Y2=2.035
r274 133 136 27.2396 $w=3.28e-07 $l=7.8e-07 $layer=LI1_cond $X=6.605 $Y=2.035
+ $X2=6.605 $Y2=2.815
r275 133 134 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.605 $Y=2.035
+ $X2=6.605 $Y2=2.035
r276 128 134 0.577444 $w=2.3e-07 $l=9e-07 $layer=MET1_cond $X=5.705 $Y=2.035
+ $X2=6.605 $Y2=2.035
r277 127 130 27.2396 $w=3.28e-07 $l=7.8e-07 $layer=LI1_cond $X=5.705 $Y=2.035
+ $X2=5.705 $Y2=2.815
r278 127 128 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.705 $Y=2.035
+ $X2=5.705 $Y2=2.035
r279 122 128 0.571028 $w=2.3e-07 $l=8.9e-07 $layer=MET1_cond $X=4.815 $Y=2.035
+ $X2=5.705 $Y2=2.035
r280 121 124 27.2396 $w=3.28e-07 $l=7.8e-07 $layer=LI1_cond $X=4.805 $Y=2.035
+ $X2=4.805 $Y2=2.815
r281 121 122 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.815 $Y=2.035
+ $X2=4.815 $Y2=2.035
r282 118 158 0.240602 $w=2.3e-07 $l=3.75e-07 $layer=MET1_cond $X=8.03 $Y=2.035
+ $X2=8.405 $Y2=2.035
r283 118 154 0.336842 $w=2.3e-07 $l=5.25e-07 $layer=MET1_cond $X=8.03 $Y=2.035
+ $X2=7.505 $Y2=2.035
r284 117 145 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=11.255 $Y=2.02
+ $X2=11.255 $Y2=2.035
r285 115 117 1.23521 $w=3.63e-07 $l=3.5e-08 $layer=LI1_cond $X=11.237 $Y=1.985
+ $X2=11.237 $Y2=2.02
r286 115 116 6.28701 $w=3.63e-07 $l=1.95e-07 $layer=LI1_cond $X=11.237 $Y=1.985
+ $X2=11.237 $Y2=1.79
r287 112 139 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=10.305 $Y=2.02
+ $X2=10.305 $Y2=2.035
r288 110 112 0.501062 $w=3.43e-07 $l=1.5e-08 $layer=LI1_cond $X=10.297 $Y=2.005
+ $X2=10.297 $Y2=2.02
r289 110 111 3.73305 $w=3.43e-07 $l=8.5e-08 $layer=LI1_cond $X=10.297 $Y=2.005
+ $X2=10.297 $Y2=1.92
r290 107 133 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=6.605 $Y=2.02
+ $X2=6.605 $Y2=2.035
r291 105 107 0.545053 $w=3.48e-07 $l=1.5e-08 $layer=LI1_cond $X=6.595 $Y=2.005
+ $X2=6.595 $Y2=2.02
r292 105 106 4.0474 $w=3.48e-07 $l=8.5e-08 $layer=LI1_cond $X=6.595 $Y=2.005
+ $X2=6.595 $Y2=1.92
r293 102 127 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=5.705 $Y=2.02
+ $X2=5.705 $Y2=2.035
r294 100 102 0.581203 $w=3.58e-07 $l=1.5e-08 $layer=LI1_cond $X=5.69 $Y=2.005
+ $X2=5.69 $Y2=2.02
r295 100 101 4.57587 $w=3.58e-07 $l=8.5e-08 $layer=LI1_cond $X=5.69 $Y=2.005
+ $X2=5.69 $Y2=1.92
r296 97 121 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=4.805 $Y=2.02
+ $X2=4.805 $Y2=2.035
r297 95 97 0.561516 $w=3.53e-07 $l=1.5e-08 $layer=LI1_cond $X=4.792 $Y=2.005
+ $X2=4.792 $Y2=2.02
r298 95 96 3.78181 $w=3.53e-07 $l=8.5e-08 $layer=LI1_cond $X=4.792 $Y=2.005
+ $X2=4.792 $Y2=1.92
r299 91 116 44.5262 $w=3.28e-07 $l=1.275e-06 $layer=LI1_cond $X=11.22 $Y=0.515
+ $X2=11.22 $Y2=1.79
r300 87 111 64.7673 $w=2.48e-07 $l=1.405e-06 $layer=LI1_cond $X=10.25 $Y=0.515
+ $X2=10.25 $Y2=1.92
r301 81 160 3.13751 $w=3.28e-07 $l=8.06226e-08 $layer=LI1_cond $X=9.32 $Y=1.92
+ $X2=9.355 $Y2=1.985
r302 81 83 64.7673 $w=2.48e-07 $l=1.405e-06 $layer=LI1_cond $X=9.32 $Y=1.92
+ $X2=9.32 $Y2=0.515
r303 77 160 7.39394 $w=3.3e-07 $l=2e-07 $layer=LI1_cond $X=9.355 $Y=2.185
+ $X2=9.355 $Y2=1.985
r304 77 79 7.50834 $w=3.28e-07 $l=2.15e-07 $layer=LI1_cond $X=9.355 $Y=2.185
+ $X2=9.355 $Y2=2.4
r305 73 156 3.09497 $w=3.2e-07 $l=7.2111e-08 $layer=LI1_cond $X=8.39 $Y=1.92
+ $X2=8.405 $Y2=1.985
r306 73 75 64.7673 $w=2.48e-07 $l=1.405e-06 $layer=LI1_cond $X=8.39 $Y=1.92
+ $X2=8.39 $Y2=0.515
r307 69 156 7.39394 $w=3.3e-07 $l=2e-07 $layer=LI1_cond $X=8.405 $Y=2.185
+ $X2=8.405 $Y2=1.985
r308 69 71 7.50834 $w=3.28e-07 $l=2.15e-07 $layer=LI1_cond $X=8.405 $Y=2.185
+ $X2=8.405 $Y2=2.4
r309 65 151 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=7.505 $Y=2.085
+ $X2=7.505 $Y2=2.005
r310 65 67 25.4934 $w=3.28e-07 $l=7.3e-07 $layer=LI1_cond $X=7.505 $Y=2.085
+ $X2=7.505 $Y2=2.815
r311 63 152 66.0891 $w=2.43e-07 $l=1.405e-06 $layer=LI1_cond $X=7.462 $Y=0.515
+ $X2=7.462 $Y2=1.92
r312 59 106 68.9014 $w=2.33e-07 $l=1.405e-06 $layer=LI1_cond $X=6.537 $Y=0.515
+ $X2=6.537 $Y2=1.92
r313 55 101 75.3108 $w=2.13e-07 $l=1.405e-06 $layer=LI1_cond $X=5.617 $Y=0.515
+ $X2=5.617 $Y2=1.92
r314 51 96 64.7673 $w=2.48e-07 $l=1.405e-06 $layer=LI1_cond $X=4.74 $Y=0.515
+ $X2=4.74 $Y2=1.92
r315 16 148 400 $w=1.7e-07 $l=1.06577e-06 $layer=licon1_PDIFF $count=1 $X=11.065
+ $Y=1.84 $X2=11.255 $Y2=2.815
r316 16 115 400 $w=1.7e-07 $l=2.5229e-07 $layer=licon1_PDIFF $count=1 $X=11.065
+ $Y=1.84 $X2=11.255 $Y2=1.985
r317 15 142 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=10.155
+ $Y=1.84 $X2=10.305 $Y2=2.815
r318 15 110 400 $w=1.7e-07 $l=2.2798e-07 $layer=licon1_PDIFF $count=1 $X=10.155
+ $Y=1.84 $X2=10.305 $Y2=2.005
r319 14 160 600 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=9.205
+ $Y=1.84 $X2=9.355 $Y2=1.985
r320 14 79 300 $w=1.7e-07 $l=6.30555e-07 $layer=licon1_PDIFF $count=2 $X=9.205
+ $Y=1.84 $X2=9.355 $Y2=2.4
r321 13 156 600 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=8.255
+ $Y=1.84 $X2=8.405 $Y2=1.985
r322 13 71 300 $w=1.7e-07 $l=6.30555e-07 $layer=licon1_PDIFF $count=2 $X=8.255
+ $Y=1.84 $X2=8.405 $Y2=2.4
r323 12 151 400 $w=1.7e-07 $l=2.2798e-07 $layer=licon1_PDIFF $count=1 $X=7.355
+ $Y=1.84 $X2=7.505 $Y2=2.005
r324 12 67 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=7.355
+ $Y=1.84 $X2=7.505 $Y2=2.815
r325 11 136 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=6.455
+ $Y=1.84 $X2=6.605 $Y2=2.815
r326 11 105 400 $w=1.7e-07 $l=2.2798e-07 $layer=licon1_PDIFF $count=1 $X=6.455
+ $Y=1.84 $X2=6.605 $Y2=2.005
r327 10 130 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=5.555
+ $Y=1.84 $X2=5.705 $Y2=2.815
r328 10 100 400 $w=1.7e-07 $l=2.2798e-07 $layer=licon1_PDIFF $count=1 $X=5.555
+ $Y=1.84 $X2=5.705 $Y2=2.005
r329 9 124 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=4.655
+ $Y=1.84 $X2=4.805 $Y2=2.815
r330 9 95 400 $w=1.7e-07 $l=2.2798e-07 $layer=licon1_PDIFF $count=1 $X=4.655
+ $Y=1.84 $X2=4.805 $Y2=2.005
r331 8 91 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=11.08
+ $Y=0.37 $X2=11.22 $Y2=0.515
r332 7 87 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=10.15
+ $Y=0.37 $X2=10.29 $Y2=0.515
r333 6 83 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=9.22
+ $Y=0.37 $X2=9.36 $Y2=0.515
r334 5 75 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=8.29
+ $Y=0.37 $X2=8.43 $Y2=0.515
r335 4 63 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=7.36
+ $Y=0.37 $X2=7.5 $Y2=0.515
r336 3 59 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=6.43
+ $Y=0.37 $X2=6.57 $Y2=0.515
r337 2 55 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=5.5
+ $Y=0.37 $X2=5.64 $Y2=0.515
r338 1 51 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=4.64
+ $Y=0.37 $X2=4.78 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__BUFINV_16%VGND 1 2 3 4 5 6 7 8 9 10 11 12 13 42 46
+ 50 54 58 62 66 70 74 78 82 86 88 90 93 94 96 97 99 100 102 103 104 106 111 129
+ 133 138 143 148 153 158 164 167 170 173 176 179 182 185 189
r214 188 189 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.76 $Y=0
+ $X2=11.76 $Y2=0
r215 185 186 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.8 $Y=0
+ $X2=10.8 $Y2=0
r216 182 183 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.84 $Y=0
+ $X2=9.84 $Y2=0
r217 179 180 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=0
+ $X2=8.88 $Y2=0
r218 176 177 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=0
+ $X2=7.92 $Y2=0
r219 173 174 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=0
+ $X2=6.96 $Y2=0
r220 167 168 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0
+ $X2=1.68 $Y2=0
r221 164 165 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0
+ $X2=0.72 $Y2=0
r222 162 189 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.28 $Y=0
+ $X2=11.76 $Y2=0
r223 162 186 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.28 $Y=0
+ $X2=10.8 $Y2=0
r224 161 162 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.28 $Y=0
+ $X2=11.28 $Y2=0
r225 159 185 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.885 $Y=0
+ $X2=10.72 $Y2=0
r226 159 161 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=10.885 $Y=0
+ $X2=11.28 $Y2=0
r227 158 188 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=11.555 $Y=0
+ $X2=11.777 $Y2=0
r228 158 161 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=11.555 $Y=0
+ $X2=11.28 $Y2=0
r229 157 186 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.32 $Y=0
+ $X2=10.8 $Y2=0
r230 157 183 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.32 $Y=0
+ $X2=9.84 $Y2=0
r231 156 157 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.32 $Y=0
+ $X2=10.32 $Y2=0
r232 154 182 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.955 $Y=0
+ $X2=9.79 $Y2=0
r233 154 156 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=9.955 $Y=0
+ $X2=10.32 $Y2=0
r234 153 185 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.555 $Y=0
+ $X2=10.72 $Y2=0
r235 153 156 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=10.555 $Y=0
+ $X2=10.32 $Y2=0
r236 152 183 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.36 $Y=0
+ $X2=9.84 $Y2=0
r237 152 180 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.36 $Y=0
+ $X2=8.88 $Y2=0
r238 151 152 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.36 $Y=0
+ $X2=9.36 $Y2=0
r239 149 179 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.025 $Y=0
+ $X2=8.86 $Y2=0
r240 149 151 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=9.025 $Y=0
+ $X2=9.36 $Y2=0
r241 148 182 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.625 $Y=0
+ $X2=9.79 $Y2=0
r242 148 151 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=9.625 $Y=0
+ $X2=9.36 $Y2=0
r243 147 180 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=0
+ $X2=8.88 $Y2=0
r244 147 177 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=0
+ $X2=7.92 $Y2=0
r245 146 147 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r246 144 176 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.095 $Y=0
+ $X2=7.93 $Y2=0
r247 144 146 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=8.095 $Y=0
+ $X2=8.4 $Y2=0
r248 143 179 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.695 $Y=0
+ $X2=8.86 $Y2=0
r249 143 146 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=8.695 $Y=0
+ $X2=8.4 $Y2=0
r250 142 177 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=0
+ $X2=7.92 $Y2=0
r251 142 174 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=0
+ $X2=6.96 $Y2=0
r252 141 142 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=0
+ $X2=7.44 $Y2=0
r253 139 173 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.165 $Y=0 $X2=7
+ $Y2=0
r254 139 141 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=7.165 $Y=0
+ $X2=7.44 $Y2=0
r255 138 176 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.765 $Y=0
+ $X2=7.93 $Y2=0
r256 138 141 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=7.765 $Y=0
+ $X2=7.44 $Y2=0
r257 137 174 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=0
+ $X2=6.96 $Y2=0
r258 136 137 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=0
+ $X2=6.48 $Y2=0
r259 134 170 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.235 $Y=0
+ $X2=6.07 $Y2=0
r260 134 136 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=6.235 $Y=0
+ $X2=6.48 $Y2=0
r261 133 173 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.835 $Y=0 $X2=7
+ $Y2=0
r262 133 136 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=6.835 $Y=0
+ $X2=6.48 $Y2=0
r263 131 132 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=0
+ $X2=5.52 $Y2=0
r264 129 170 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.905 $Y=0
+ $X2=6.07 $Y2=0
r265 129 131 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=5.905 $Y=0
+ $X2=5.52 $Y2=0
r266 128 132 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=0
+ $X2=5.52 $Y2=0
r267 127 128 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.04 $Y=0
+ $X2=5.04 $Y2=0
r268 125 128 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.08 $Y=0
+ $X2=5.04 $Y2=0
r269 124 125 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=0
+ $X2=4.08 $Y2=0
r270 122 125 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=0
+ $X2=4.08 $Y2=0
r271 121 122 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=0
+ $X2=3.12 $Y2=0
r272 119 122 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0
+ $X2=3.12 $Y2=0
r273 119 168 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0
+ $X2=1.68 $Y2=0
r274 118 119 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0
+ $X2=2.16 $Y2=0
r275 116 167 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.795 $Y=0
+ $X2=1.63 $Y2=0
r276 116 118 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=1.795 $Y=0
+ $X2=2.16 $Y2=0
r277 115 168 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0
+ $X2=1.68 $Y2=0
r278 115 165 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0
+ $X2=0.72 $Y2=0
r279 114 115 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r280 112 164 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.875 $Y=0
+ $X2=0.71 $Y2=0
r281 112 114 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.875 $Y=0
+ $X2=1.2 $Y2=0
r282 111 167 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.465 $Y=0
+ $X2=1.63 $Y2=0
r283 111 114 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=1.465 $Y=0
+ $X2=1.2 $Y2=0
r284 109 165 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0
+ $X2=0.72 $Y2=0
r285 108 109 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0
+ $X2=0.24 $Y2=0
r286 106 164 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.545 $Y=0
+ $X2=0.71 $Y2=0
r287 106 108 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.545 $Y=0
+ $X2=0.24 $Y2=0
r288 104 137 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=0 $X2=6.48
+ $Y2=0
r289 104 132 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=0 $X2=5.52
+ $Y2=0
r290 104 170 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=0 $X2=6
+ $Y2=0
r291 102 127 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=5.045 $Y=0
+ $X2=5.04 $Y2=0
r292 102 103 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.045 $Y=0
+ $X2=5.17 $Y2=0
r293 101 131 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=5.295 $Y=0
+ $X2=5.52 $Y2=0
r294 101 103 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.295 $Y=0
+ $X2=5.17 $Y2=0
r295 99 124 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=4.115 $Y=0
+ $X2=4.08 $Y2=0
r296 99 100 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.115 $Y=0
+ $X2=4.28 $Y2=0
r297 98 127 38.8182 $w=1.68e-07 $l=5.95e-07 $layer=LI1_cond $X=4.445 $Y=0
+ $X2=5.04 $Y2=0
r298 98 100 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.445 $Y=0
+ $X2=4.28 $Y2=0
r299 96 121 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=3.185 $Y=0
+ $X2=3.12 $Y2=0
r300 96 97 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.185 $Y=0 $X2=3.35
+ $Y2=0
r301 95 124 36.861 $w=1.68e-07 $l=5.65e-07 $layer=LI1_cond $X=3.515 $Y=0
+ $X2=4.08 $Y2=0
r302 95 97 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.515 $Y=0 $X2=3.35
+ $Y2=0
r303 93 118 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=2.325 $Y=0
+ $X2=2.16 $Y2=0
r304 93 94 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.325 $Y=0 $X2=2.45
+ $Y2=0
r305 92 121 35.5561 $w=1.68e-07 $l=5.45e-07 $layer=LI1_cond $X=2.575 $Y=0
+ $X2=3.12 $Y2=0
r306 92 94 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.575 $Y=0 $X2=2.45
+ $Y2=0
r307 88 188 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=11.72 $Y=0.085
+ $X2=11.777 $Y2=0
r308 88 90 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=11.72 $Y=0.085
+ $X2=11.72 $Y2=0.515
r309 84 185 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=10.72 $Y=0.085
+ $X2=10.72 $Y2=0
r310 84 86 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=10.72 $Y=0.085
+ $X2=10.72 $Y2=0.515
r311 80 182 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.79 $Y=0.085
+ $X2=9.79 $Y2=0
r312 80 82 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=9.79 $Y=0.085
+ $X2=9.79 $Y2=0.515
r313 76 179 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.86 $Y=0.085
+ $X2=8.86 $Y2=0
r314 76 78 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=8.86 $Y=0.085
+ $X2=8.86 $Y2=0.515
r315 72 176 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.93 $Y=0.085
+ $X2=7.93 $Y2=0
r316 72 74 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=7.93 $Y=0.085
+ $X2=7.93 $Y2=0.515
r317 68 173 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7 $Y=0.085 $X2=7
+ $Y2=0
r318 68 70 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=7 $Y=0.085 $X2=7
+ $Y2=0.515
r319 64 170 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.07 $Y=0.085
+ $X2=6.07 $Y2=0
r320 64 66 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=6.07 $Y=0.085
+ $X2=6.07 $Y2=0.515
r321 60 103 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.17 $Y=0.085
+ $X2=5.17 $Y2=0
r322 60 62 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=5.17 $Y=0.085
+ $X2=5.17 $Y2=0.515
r323 56 100 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.28 $Y=0.085
+ $X2=4.28 $Y2=0
r324 56 58 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=4.28 $Y=0.085
+ $X2=4.28 $Y2=0.515
r325 52 97 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.35 $Y=0.085
+ $X2=3.35 $Y2=0
r326 52 54 18.8582 $w=3.28e-07 $l=5.4e-07 $layer=LI1_cond $X=3.35 $Y=0.085
+ $X2=3.35 $Y2=0.625
r327 48 94 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.45 $Y=0.085
+ $X2=2.45 $Y2=0
r328 48 50 24.8928 $w=2.48e-07 $l=5.4e-07 $layer=LI1_cond $X=2.45 $Y=0.085
+ $X2=2.45 $Y2=0.625
r329 44 167 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.63 $Y=0.085
+ $X2=1.63 $Y2=0
r330 44 46 20.6043 $w=3.28e-07 $l=5.9e-07 $layer=LI1_cond $X=1.63 $Y=0.085
+ $X2=1.63 $Y2=0.675
r331 40 164 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.71 $Y=0.085
+ $X2=0.71 $Y2=0
r332 40 42 20.6043 $w=3.28e-07 $l=5.9e-07 $layer=LI1_cond $X=0.71 $Y=0.085
+ $X2=0.71 $Y2=0.675
r333 13 90 91 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=2 $X=11.51
+ $Y=0.37 $X2=11.72 $Y2=0.515
r334 12 86 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=10.58
+ $Y=0.37 $X2=10.72 $Y2=0.515
r335 11 82 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=9.65
+ $Y=0.37 $X2=9.79 $Y2=0.515
r336 10 78 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=8.72
+ $Y=0.37 $X2=8.86 $Y2=0.515
r337 9 74 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=7.79
+ $Y=0.37 $X2=7.93 $Y2=0.515
r338 8 70 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=6.86
+ $Y=0.37 $X2=7 $Y2=0.515
r339 7 66 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=5.93
+ $Y=0.37 $X2=6.07 $Y2=0.515
r340 6 62 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=5.07
+ $Y=0.37 $X2=5.21 $Y2=0.515
r341 5 58 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=4.14
+ $Y=0.37 $X2=4.28 $Y2=0.515
r342 4 54 182 $w=1.7e-07 $l=3.17372e-07 $layer=licon1_NDIFF $count=1 $X=3.21
+ $Y=0.37 $X2=3.35 $Y2=0.625
r343 3 50 182 $w=1.7e-07 $l=3.17372e-07 $layer=licon1_NDIFF $count=1 $X=2.35
+ $Y=0.37 $X2=2.49 $Y2=0.625
r344 2 46 182 $w=1.7e-07 $l=3.68409e-07 $layer=licon1_NDIFF $count=1 $X=1.49
+ $Y=0.37 $X2=1.63 $Y2=0.675
r345 1 42 182 $w=1.7e-07 $l=3.68409e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.37 $X2=0.71 $Y2=0.675
.ends

