* File: sky130_fd_sc_hs__nor2_1.pxi.spice
* Created: Thu Aug 27 20:52:57 2020
* 
x_PM_SKY130_FD_SC_HS__NOR2_1%A N_A_c_27_n N_A_M1001_g N_A_M1003_g A N_A_c_29_n
+ PM_SKY130_FD_SC_HS__NOR2_1%A
x_PM_SKY130_FD_SC_HS__NOR2_1%B N_B_c_51_n N_B_M1000_g N_B_M1002_g B N_B_c_53_n
+ PM_SKY130_FD_SC_HS__NOR2_1%B
x_PM_SKY130_FD_SC_HS__NOR2_1%VPWR N_VPWR_M1001_s N_VPWR_c_72_n N_VPWR_c_73_n
+ VPWR N_VPWR_c_74_n N_VPWR_c_71_n PM_SKY130_FD_SC_HS__NOR2_1%VPWR
x_PM_SKY130_FD_SC_HS__NOR2_1%Y N_Y_M1003_d N_Y_M1000_d N_Y_c_88_n N_Y_c_89_n
+ N_Y_c_90_n Y Y PM_SKY130_FD_SC_HS__NOR2_1%Y
x_PM_SKY130_FD_SC_HS__NOR2_1%VGND N_VGND_M1003_s N_VGND_M1002_d N_VGND_c_114_n
+ N_VGND_c_115_n N_VGND_c_116_n N_VGND_c_117_n VGND N_VGND_c_118_n
+ N_VGND_c_119_n PM_SKY130_FD_SC_HS__NOR2_1%VGND
cc_1 VNB N_A_c_27_n 0.0591502f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.765
cc_2 VNB N_A_M1003_g 0.0271489f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=0.74
cc_3 VNB N_A_c_29_n 0.00600492f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.465
cc_4 VNB N_B_c_51_n 0.061027f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.765
cc_5 VNB N_B_M1002_g 0.028217f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=0.74
cc_6 VNB N_B_c_53_n 0.00385705f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.465
cc_7 VNB N_VPWR_c_71_n 0.0641695f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.665
cc_8 VNB N_Y_c_88_n 0.00206666f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_Y_c_89_n 0.00960735f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.465
cc_10 VNB N_Y_c_90_n 0.0022354f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.465
cc_11 VNB N_VGND_c_114_n 0.011316f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_VGND_c_115_n 0.0411496f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_VGND_c_116_n 0.0120272f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.465
cc_14 VNB N_VGND_c_117_n 0.0404679f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.465
cc_15 VNB N_VGND_c_118_n 0.0172524f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_VGND_c_119_n 0.115949f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VPB N_A_c_27_n 0.0270256f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.765
cc_18 VPB N_A_c_29_n 0.00730438f $X=-0.19 $Y=1.66 $X2=0.29 $Y2=1.465
cc_19 VPB N_B_c_51_n 0.0286509f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.765
cc_20 VPB N_B_c_53_n 0.00739755f $X=-0.19 $Y=1.66 $X2=0.29 $Y2=1.465
cc_21 VPB N_VPWR_c_72_n 0.0120106f $X=-0.19 $Y=1.66 $X2=0.515 $Y2=1.3
cc_22 VPB N_VPWR_c_73_n 0.0489132f $X=-0.19 $Y=1.66 $X2=0.515 $Y2=0.74
cc_23 VPB N_VPWR_c_74_n 0.0288332f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_24 VPB N_VPWR_c_71_n 0.0521156f $X=-0.19 $Y=1.66 $X2=0.29 $Y2=1.665
cc_25 VPB N_Y_c_89_n 0.00320283f $X=-0.19 $Y=1.66 $X2=0.29 $Y2=1.465
cc_26 VPB Y 0.0452381f $X=-0.19 $Y=1.66 $X2=0.29 $Y2=1.665
cc_27 N_A_c_27_n N_B_c_51_n 0.0783329f $X=0.505 $Y=1.765 $X2=-0.19 $Y2=-0.245
cc_28 N_A_M1003_g N_B_M1002_g 0.0144801f $X=0.515 $Y=0.74 $X2=0 $Y2=0
cc_29 N_A_c_27_n N_VPWR_c_73_n 0.0175184f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_30 N_A_c_29_n N_VPWR_c_73_n 0.0257783f $X=0.29 $Y=1.465 $X2=0 $Y2=0
cc_31 N_A_c_27_n N_VPWR_c_74_n 0.00413917f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_32 N_A_c_27_n N_VPWR_c_71_n 0.00817532f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_33 N_A_M1003_g N_Y_c_88_n 0.00809519f $X=0.515 $Y=0.74 $X2=0 $Y2=0
cc_34 N_A_c_27_n N_Y_c_89_n 0.00762011f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_35 N_A_M1003_g N_Y_c_89_n 0.00403324f $X=0.515 $Y=0.74 $X2=0 $Y2=0
cc_36 N_A_c_29_n N_Y_c_89_n 0.0331382f $X=0.29 $Y=1.465 $X2=0 $Y2=0
cc_37 N_A_c_27_n N_Y_c_90_n 2.30445e-19 $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_38 N_A_M1003_g N_Y_c_90_n 0.0027623f $X=0.515 $Y=0.74 $X2=0 $Y2=0
cc_39 N_A_c_27_n Y 0.0080758f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_40 N_A_c_27_n N_VGND_c_115_n 0.00196285f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_41 N_A_M1003_g N_VGND_c_115_n 0.00511162f $X=0.515 $Y=0.74 $X2=0 $Y2=0
cc_42 N_A_c_29_n N_VGND_c_115_n 0.0215684f $X=0.29 $Y=1.465 $X2=0 $Y2=0
cc_43 N_A_M1003_g N_VGND_c_117_n 6.14817e-19 $X=0.515 $Y=0.74 $X2=0 $Y2=0
cc_44 N_A_M1003_g N_VGND_c_118_n 0.00434272f $X=0.515 $Y=0.74 $X2=0 $Y2=0
cc_45 N_A_M1003_g N_VGND_c_119_n 0.00824106f $X=0.515 $Y=0.74 $X2=0 $Y2=0
cc_46 N_B_c_51_n N_VPWR_c_73_n 0.00152333f $X=0.925 $Y=1.765 $X2=0 $Y2=0
cc_47 N_B_c_51_n N_VPWR_c_74_n 0.00302115f $X=0.925 $Y=1.765 $X2=0 $Y2=0
cc_48 N_B_c_51_n N_VPWR_c_71_n 0.00374141f $X=0.925 $Y=1.765 $X2=0 $Y2=0
cc_49 N_B_M1002_g N_Y_c_88_n 0.00457569f $X=0.945 $Y=0.74 $X2=0 $Y2=0
cc_50 N_B_c_51_n N_Y_c_89_n 0.00565932f $X=0.925 $Y=1.765 $X2=0 $Y2=0
cc_51 N_B_c_53_n N_Y_c_89_n 0.0360321f $X=1.15 $Y=1.465 $X2=0 $Y2=0
cc_52 N_B_c_51_n Y 0.0338169f $X=0.925 $Y=1.765 $X2=0 $Y2=0
cc_53 N_B_c_53_n Y 0.0266913f $X=1.15 $Y=1.465 $X2=0 $Y2=0
cc_54 N_B_c_51_n N_VGND_c_117_n 0.00232693f $X=0.925 $Y=1.765 $X2=0 $Y2=0
cc_55 N_B_M1002_g N_VGND_c_117_n 0.0151529f $X=0.945 $Y=0.74 $X2=0 $Y2=0
cc_56 N_B_c_53_n N_VGND_c_117_n 0.0275482f $X=1.15 $Y=1.465 $X2=0 $Y2=0
cc_57 N_B_M1002_g N_VGND_c_118_n 0.00383152f $X=0.945 $Y=0.74 $X2=0 $Y2=0
cc_58 N_B_M1002_g N_VGND_c_119_n 0.00757637f $X=0.945 $Y=0.74 $X2=0 $Y2=0
cc_59 N_VPWR_c_73_n Y 0.0710044f $X=0.28 $Y=2.115 $X2=0 $Y2=0
cc_60 N_VPWR_c_74_n Y 0.0243273f $X=1.2 $Y=3.33 $X2=0 $Y2=0
cc_61 N_VPWR_c_71_n Y 0.0232642f $X=1.2 $Y=3.33 $X2=0 $Y2=0
cc_62 A_116_368# N_Y_c_89_n 0.00134547f $X=0.58 $Y=1.84 $X2=0.73 $Y2=1.95
cc_63 A_116_368# Y 0.0118291f $X=0.58 $Y=1.84 $X2=1.115 $Y2=2.69
cc_64 N_Y_c_88_n N_VGND_c_115_n 0.0282134f $X=0.73 $Y=0.515 $X2=0 $Y2=0
cc_65 N_Y_c_88_n N_VGND_c_117_n 0.0294122f $X=0.73 $Y=0.515 $X2=0 $Y2=0
cc_66 N_Y_c_88_n N_VGND_c_118_n 0.0109942f $X=0.73 $Y=0.515 $X2=0 $Y2=0
cc_67 N_Y_c_88_n N_VGND_c_119_n 0.00904371f $X=0.73 $Y=0.515 $X2=0 $Y2=0
