* File: sky130_fd_sc_hs__mux2i_2.spice
* Created: Tue Sep  1 20:07:59 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hs__mux2i_2.pex.spice"
.subckt sky130_fd_sc_hs__mux2i_2  VNB VPB A0 A1 S Y VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* Y	Y
* S	S
* A1	A1
* A0	A0
* VPB	VPB
* VNB	VNB
MM1008 N_A_115_74#_M1008_d N_A0_M1008_g N_Y_M1008_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1369 AS=0.2109 PD=1.11 PS=2.05 NRD=14.592 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75002.2 A=0.111 P=1.78 MULT=1
MM1016 N_A_115_74#_M1008_d N_A0_M1016_g N_Y_M1016_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1369 AS=0.188175 PD=1.11 PS=1.355 NRD=0 NRS=32.316 M=1 R=4.93333
+ SA=75000.7 SB=75001.7 A=0.111 P=1.78 MULT=1
MM1003 N_A_337_74#_M1003_d N_A1_M1003_g N_Y_M1016_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.270675 AS=0.188175 PD=1.505 PS=1.355 NRD=2.016 NRS=32.316 M=1 R=4.93333
+ SA=75001.3 SB=75001.1 A=0.111 P=1.78 MULT=1
MM1015 N_A_337_74#_M1003_d N_A1_M1015_g N_Y_M1015_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.270675 AS=0.2553 PD=1.505 PS=2.17 NRD=56.748 NRS=9.72 M=1 R=4.93333
+ SA=75002.2 SB=75000.3 A=0.111 P=1.78 MULT=1
MM1011 N_A_337_74#_M1011_d N_S_M1011_g N_VGND_M1011_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1221 AS=0.36 PD=1.07 PS=2.83 NRD=4.044 NRS=69.96 M=1 R=4.93333 SA=75000.3
+ SB=75002.3 A=0.111 P=1.78 MULT=1
MM1013 N_A_337_74#_M1011_d N_S_M1013_g N_VGND_M1013_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1221 AS=0.215625 PD=1.07 PS=1.505 NRD=4.044 NRS=38.328 M=1 R=4.93333
+ SA=75000.8 SB=75001.8 A=0.111 P=1.78 MULT=1
MM1002 N_VGND_M1013_s N_A_922_72#_M1002_g N_A_115_74#_M1002_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.215625 AS=0.1221 PD=1.505 PS=1.07 NRD=38.328 NRS=4.044 M=1
+ R=4.93333 SA=75001.4 SB=75001.2 A=0.111 P=1.78 MULT=1
MM1017 N_VGND_M1017_d N_A_922_72#_M1017_g N_A_115_74#_M1002_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.166607 AS=0.1221 PD=1.25478 PS=1.07 NRD=11.34 NRS=4.044 M=1
+ R=4.93333 SA=75001.9 SB=75000.7 A=0.111 P=1.78 MULT=1
MM1010 N_A_922_72#_M1010_d N_S_M1010_g N_VGND_M1017_d VNB NLOWVT L=0.15 W=0.64
+ AD=0.1824 AS=0.144093 PD=1.85 PS=1.08522 NRD=0 NRS=15.936 M=1 R=4.26667
+ SA=75002.4 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1000 N_A_118_368#_M1000_d N_A0_M1000_g N_Y_M1000_s VPB PSHORT L=0.15 W=1.12
+ AD=0.1904 AS=0.3416 PD=1.46 PS=2.85 NRD=8.7862 NRS=3.5066 M=1 R=7.46667
+ SA=75000.2 SB=75002.2 A=0.168 P=2.54 MULT=1
MM1005 N_A_118_368#_M1000_d N_A0_M1005_g N_Y_M1005_s VPB PSHORT L=0.15 W=1.12
+ AD=0.1904 AS=0.2632 PD=1.46 PS=1.59 NRD=1.7533 NRS=16.7056 M=1 R=7.46667
+ SA=75000.7 SB=75001.7 A=0.168 P=2.54 MULT=1
MM1006 N_Y_M1005_s N_A1_M1006_g N_A_340_368#_M1006_s VPB PSHORT L=0.15 W=1.12
+ AD=0.2632 AS=0.3808 PD=1.59 PS=1.8 NRD=16.7056 NRS=1.7533 M=1 R=7.46667
+ SA=75001.3 SB=75001 A=0.168 P=2.54 MULT=1
MM1007 N_Y_M1007_d N_A1_M1007_g N_A_340_368#_M1006_s VPB PSHORT L=0.15 W=1.12
+ AD=0.3304 AS=0.3808 PD=2.83 PS=1.8 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75002.2 SB=75000.2 A=0.168 P=2.54 MULT=1
MM1009 N_A_118_368#_M1009_d N_S_M1009_g N_VPWR_M1009_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.581825 PD=1.42 PS=3.6 NRD=1.7533 NRS=81.6959 M=1 R=7.46667
+ SA=75000.4 SB=75002.3 A=0.168 P=2.54 MULT=1
MM1012 N_A_118_368#_M1009_d N_S_M1012_g N_VPWR_M1012_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.3021 PD=1.42 PS=1.805 NRD=0 NRS=37.7649 M=1 R=7.46667 SA=75000.8
+ SB=75001.8 A=0.168 P=2.54 MULT=1
MM1001 N_A_340_368#_M1001_d N_A_922_72#_M1001_g N_VPWR_M1012_s VPB PSHORT L=0.15
+ W=1.12 AD=0.168 AS=0.3021 PD=1.42 PS=1.805 NRD=0 NRS=37.7649 M=1 R=7.46667
+ SA=75001.5 SB=75001.2 A=0.168 P=2.54 MULT=1
MM1004 N_A_340_368#_M1001_d N_A_922_72#_M1004_g N_VPWR_M1004_s VPB PSHORT L=0.15
+ W=1.12 AD=0.168 AS=0.251683 PD=1.42 PS=1.64302 NRD=1.7533 NRS=10.5395 M=1
+ R=7.46667 SA=75001.9 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1014 N_A_922_72#_M1014_d N_S_M1014_g N_VPWR_M1004_s VPB PSHORT L=0.15 W=1
+ AD=0.295 AS=0.224717 PD=2.59 PS=1.46698 NRD=1.9503 NRS=19.1878 M=1 R=6.66667
+ SA=75002.5 SB=75000.2 A=0.15 P=2.3 MULT=1
DX18_noxref VNB VPB NWDIODE A=12.3132 P=16.96
*
.include "sky130_fd_sc_hs__mux2i_2.pxi.spice"
*
.ends
*
*
