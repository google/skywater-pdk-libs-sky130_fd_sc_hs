* File: sky130_fd_sc_hs__o21ba_2.pxi.spice
* Created: Tue Sep  1 20:14:55 2020
* 
x_PM_SKY130_FD_SC_HS__O21BA_2%B1_N N_B1_N_M1003_g N_B1_N_c_70_n N_B1_N_M1005_g
+ B1_N N_B1_N_c_71_n PM_SKY130_FD_SC_HS__O21BA_2%B1_N
x_PM_SKY130_FD_SC_HS__O21BA_2%A_177_48# N_A_177_48#_M1011_s N_A_177_48#_M1004_d
+ N_A_177_48#_M1001_g N_A_177_48#_c_104_n N_A_177_48#_M1006_g
+ N_A_177_48#_M1009_g N_A_177_48#_c_105_n N_A_177_48#_M1008_g N_A_177_48#_c_98_n
+ N_A_177_48#_c_99_n N_A_177_48#_c_106_n N_A_177_48#_c_100_n N_A_177_48#_c_101_n
+ N_A_177_48#_c_107_n N_A_177_48#_c_102_n N_A_177_48#_c_103_n
+ PM_SKY130_FD_SC_HS__O21BA_2%A_177_48#
x_PM_SKY130_FD_SC_HS__O21BA_2%A_27_74# N_A_27_74#_M1003_s N_A_27_74#_M1005_s
+ N_A_27_74#_M1011_g N_A_27_74#_c_205_n N_A_27_74#_M1004_g N_A_27_74#_c_198_n
+ N_A_27_74#_c_199_n N_A_27_74#_c_200_n N_A_27_74#_c_201_n N_A_27_74#_c_202_n
+ N_A_27_74#_c_203_n N_A_27_74#_c_240_n N_A_27_74#_c_204_n N_A_27_74#_c_210_n
+ PM_SKY130_FD_SC_HS__O21BA_2%A_27_74#
x_PM_SKY130_FD_SC_HS__O21BA_2%A2 N_A2_c_284_n N_A2_M1002_g N_A2_c_285_n
+ N_A2_M1007_g A2 PM_SKY130_FD_SC_HS__O21BA_2%A2
x_PM_SKY130_FD_SC_HS__O21BA_2%A1 N_A1_c_316_n N_A1_M1000_g N_A1_c_317_n
+ N_A1_M1010_g A1 PM_SKY130_FD_SC_HS__O21BA_2%A1
x_PM_SKY130_FD_SC_HS__O21BA_2%VPWR N_VPWR_M1005_d N_VPWR_M1008_s N_VPWR_M1000_d
+ N_VPWR_c_339_n N_VPWR_c_340_n N_VPWR_c_341_n VPWR N_VPWR_c_342_n
+ N_VPWR_c_343_n N_VPWR_c_344_n N_VPWR_c_345_n N_VPWR_c_338_n
+ PM_SKY130_FD_SC_HS__O21BA_2%VPWR
x_PM_SKY130_FD_SC_HS__O21BA_2%X N_X_M1001_s N_X_M1006_d N_X_c_382_n N_X_c_386_n
+ X X X PM_SKY130_FD_SC_HS__O21BA_2%X
x_PM_SKY130_FD_SC_HS__O21BA_2%VGND N_VGND_M1003_d N_VGND_M1009_d N_VGND_M1002_d
+ N_VGND_c_417_n N_VGND_c_418_n N_VGND_c_419_n N_VGND_c_420_n N_VGND_c_421_n
+ VGND N_VGND_c_422_n N_VGND_c_423_n N_VGND_c_424_n N_VGND_c_425_n
+ N_VGND_c_426_n N_VGND_c_427_n PM_SKY130_FD_SC_HS__O21BA_2%VGND
x_PM_SKY130_FD_SC_HS__O21BA_2%A_487_74# N_A_487_74#_M1011_d N_A_487_74#_M1010_d
+ N_A_487_74#_c_479_n N_A_487_74#_c_473_n N_A_487_74#_c_474_n
+ PM_SKY130_FD_SC_HS__O21BA_2%A_487_74#
cc_1 VNB N_B1_N_M1003_g 0.0415411f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=0.645
cc_2 VNB N_B1_N_c_70_n 0.0599021f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.765
cc_3 VNB N_B1_N_c_71_n 0.0037649f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.465
cc_4 VNB N_A_177_48#_M1001_g 0.0234736f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_5 VNB N_A_177_48#_M1009_g 0.0223256f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_6 VNB N_A_177_48#_c_98_n 0.0164379f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_7 VNB N_A_177_48#_c_99_n 0.00911858f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_A_177_48#_c_100_n 0.00963453f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A_177_48#_c_101_n 0.00364368f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_177_48#_c_102_n 0.00360224f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_177_48#_c_103_n 0.0606756f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_27_74#_M1011_g 0.0270364f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_27_74#_c_198_n 0.0292115f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_27_74#_c_199_n 0.0111157f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.665
cc_15 VNB N_A_27_74#_c_200_n 0.0194899f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_27_74#_c_201_n 0.00436079f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_27_74#_c_202_n 0.00988676f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_27_74#_c_203_n 0.00937892f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_27_74#_c_204_n 0.00298618f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A2_c_284_n 0.0186845f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=1.3
cc_21 VNB N_A2_c_285_n 0.0400289f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB A2 0.0138799f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.26
cc_23 VNB N_A1_c_316_n 0.0673897f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=1.3
cc_24 VNB N_A1_c_317_n 0.024572f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB A1 0.00756722f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.26
cc_26 VNB N_VPWR_c_338_n 0.163682f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_X_c_382_n 0.00199855f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_28 VNB X 0.00240191f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB X 0.00419424f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.665
cc_30 VNB N_VGND_c_417_n 0.00562672f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.465
cc_31 VNB N_VGND_c_418_n 0.0136548f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_419_n 0.00790898f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_420_n 0.0174338f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_421_n 0.00461913f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_422_n 0.0207632f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_423_n 0.0310006f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_424_n 0.017961f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_425_n 0.239258f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_426_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_427_n 0.00631651f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_487_74#_c_473_n 0.00238751f $X=-0.19 $Y=-0.245 $X2=0.36 $Y2=1.465
cc_42 VNB N_A_487_74#_c_474_n 0.0284841f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.665
cc_43 VPB N_B1_N_c_70_n 0.0296259f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.765
cc_44 VPB N_B1_N_c_71_n 0.00730438f $X=-0.19 $Y=1.66 $X2=0.29 $Y2=1.465
cc_45 VPB N_A_177_48#_c_104_n 0.0169074f $X=-0.19 $Y=1.66 $X2=0.29 $Y2=1.465
cc_46 VPB N_A_177_48#_c_105_n 0.0173586f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_47 VPB N_A_177_48#_c_106_n 0.003137f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_48 VPB N_A_177_48#_c_107_n 0.00707359f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_49 VPB N_A_177_48#_c_102_n 0.00155932f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_50 VPB N_A_177_48#_c_103_n 0.0141865f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_51 VPB N_A_27_74#_c_205_n 0.015301f $X=-0.19 $Y=1.66 $X2=0.29 $Y2=1.465
cc_52 VPB N_A_27_74#_c_198_n 0.0141697f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_53 VPB N_A_27_74#_c_199_n 0.00771623f $X=-0.19 $Y=1.66 $X2=0.29 $Y2=1.665
cc_54 VPB N_A_27_74#_c_203_n 0.00312372f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_55 VPB N_A_27_74#_c_204_n 0.0027552f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_56 VPB N_A_27_74#_c_210_n 0.0348417f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_57 VPB N_A2_c_285_n 0.0230933f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_58 VPB N_A1_c_316_n 0.0290811f $X=-0.19 $Y=1.66 $X2=0.485 $Y2=1.3
cc_59 VPB N_VPWR_c_339_n 0.0165465f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_60 VPB N_VPWR_c_340_n 0.0118719f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_61 VPB N_VPWR_c_341_n 0.0617288f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_62 VPB N_VPWR_c_342_n 0.0182672f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_63 VPB N_VPWR_c_343_n 0.0351759f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_64 VPB N_VPWR_c_344_n 0.0274943f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_65 VPB N_VPWR_c_345_n 0.0273298f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_66 VPB N_VPWR_c_338_n 0.0939968f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_67 VPB N_X_c_382_n 0.00176723f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_68 VPB N_X_c_386_n 0.0023595f $X=-0.19 $Y=1.66 $X2=0.29 $Y2=1.465
cc_69 N_B1_N_M1003_g N_A_177_48#_M1001_g 0.0214791f $X=0.485 $Y=0.645 $X2=0
+ $Y2=0
cc_70 N_B1_N_c_70_n N_A_177_48#_M1001_g 0.0120528f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_71 N_B1_N_c_70_n N_A_177_48#_c_104_n 0.0234657f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_72 N_B1_N_c_70_n N_A_177_48#_c_103_n 0.00413087f $X=0.505 $Y=1.765 $X2=0
+ $Y2=0
cc_73 N_B1_N_M1003_g N_A_27_74#_c_200_n 0.00265886f $X=0.485 $Y=0.645 $X2=0
+ $Y2=0
cc_74 N_B1_N_M1003_g N_A_27_74#_c_201_n 0.0186832f $X=0.485 $Y=0.645 $X2=0 $Y2=0
cc_75 N_B1_N_c_70_n N_A_27_74#_c_201_n 0.00180385f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_76 N_B1_N_c_71_n N_A_27_74#_c_201_n 0.00749401f $X=0.29 $Y=1.465 $X2=0 $Y2=0
cc_77 N_B1_N_c_70_n N_A_27_74#_c_202_n 0.00180238f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_78 N_B1_N_c_71_n N_A_27_74#_c_202_n 0.0199042f $X=0.29 $Y=1.465 $X2=0 $Y2=0
cc_79 N_B1_N_M1003_g N_A_27_74#_c_203_n 0.00407925f $X=0.485 $Y=0.645 $X2=0
+ $Y2=0
cc_80 N_B1_N_c_70_n N_A_27_74#_c_203_n 0.00642088f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_81 N_B1_N_c_71_n N_A_27_74#_c_203_n 0.0360322f $X=0.29 $Y=1.465 $X2=0 $Y2=0
cc_82 N_B1_N_c_70_n N_A_27_74#_c_210_n 0.0323323f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_83 N_B1_N_c_71_n N_A_27_74#_c_210_n 0.026581f $X=0.29 $Y=1.465 $X2=0 $Y2=0
cc_84 N_B1_N_c_70_n N_VPWR_c_339_n 0.00418414f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_85 N_B1_N_c_70_n N_VPWR_c_344_n 0.00393265f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_86 N_B1_N_c_70_n N_VPWR_c_338_n 0.00462577f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_87 N_B1_N_M1003_g X 8.0174e-19 $X=0.485 $Y=0.645 $X2=0 $Y2=0
cc_88 N_B1_N_M1003_g N_VGND_c_417_n 0.0151909f $X=0.485 $Y=0.645 $X2=0 $Y2=0
cc_89 N_B1_N_M1003_g N_VGND_c_420_n 0.00383152f $X=0.485 $Y=0.645 $X2=0 $Y2=0
cc_90 N_B1_N_M1003_g N_VGND_c_425_n 0.00761163f $X=0.485 $Y=0.645 $X2=0 $Y2=0
cc_91 N_A_177_48#_c_99_n N_A_27_74#_M1011_g 0.00159319f $X=2.145 $Y=0.515 $X2=0
+ $Y2=0
cc_92 N_A_177_48#_c_100_n N_A_27_74#_M1011_g 0.00286806f $X=1.515 $Y=1.095 $X2=0
+ $Y2=0
cc_93 N_A_177_48#_c_101_n N_A_27_74#_M1011_g 0.0153167f $X=2.465 $Y=1.095 $X2=0
+ $Y2=0
cc_94 N_A_177_48#_c_102_n N_A_27_74#_M1011_g 0.0084954f $X=2.577 $Y=1.82 $X2=0
+ $Y2=0
cc_95 N_A_177_48#_c_103_n N_A_27_74#_M1011_g 7.05618e-19 $X=1.5 $Y=1.532 $X2=0
+ $Y2=0
cc_96 N_A_177_48#_c_106_n N_A_27_74#_c_205_n 0.0106833f $X=2.61 $Y=2.695 $X2=0
+ $Y2=0
cc_97 N_A_177_48#_c_107_n N_A_27_74#_c_205_n 0.0118395f $X=2.61 $Y=1.985 $X2=0
+ $Y2=0
cc_98 N_A_177_48#_c_102_n N_A_27_74#_c_205_n 0.0010952f $X=2.577 $Y=1.82 $X2=0
+ $Y2=0
cc_99 N_A_177_48#_c_98_n N_A_27_74#_c_198_n 0.00223955f $X=1.98 $Y=1.095 $X2=0
+ $Y2=0
cc_100 N_A_177_48#_c_100_n N_A_27_74#_c_198_n 0.00108808f $X=1.515 $Y=1.095
+ $X2=0 $Y2=0
cc_101 N_A_177_48#_c_101_n N_A_27_74#_c_198_n 0.00283481f $X=2.465 $Y=1.095
+ $X2=0 $Y2=0
cc_102 N_A_177_48#_c_103_n N_A_27_74#_c_198_n 0.0208131f $X=1.5 $Y=1.532 $X2=0
+ $Y2=0
cc_103 N_A_177_48#_c_102_n N_A_27_74#_c_199_n 0.011868f $X=2.577 $Y=1.82 $X2=0
+ $Y2=0
cc_104 N_A_177_48#_c_103_n N_A_27_74#_c_199_n 7.55131e-19 $X=1.5 $Y=1.532 $X2=0
+ $Y2=0
cc_105 N_A_177_48#_M1001_g N_A_27_74#_c_201_n 0.00150892f $X=0.96 $Y=0.74 $X2=0
+ $Y2=0
cc_106 N_A_177_48#_M1001_g N_A_27_74#_c_203_n 0.00390955f $X=0.96 $Y=0.74 $X2=0
+ $Y2=0
cc_107 N_A_177_48#_c_104_n N_A_27_74#_c_203_n 0.00131837f $X=1.05 $Y=1.765 $X2=0
+ $Y2=0
cc_108 N_A_177_48#_c_103_n N_A_27_74#_c_203_n 0.00118563f $X=1.5 $Y=1.532 $X2=0
+ $Y2=0
cc_109 N_A_177_48#_c_104_n N_A_27_74#_c_240_n 0.0166143f $X=1.05 $Y=1.765 $X2=0
+ $Y2=0
cc_110 N_A_177_48#_c_105_n N_A_27_74#_c_240_n 0.0187212f $X=1.5 $Y=1.765 $X2=0
+ $Y2=0
cc_111 N_A_177_48#_c_100_n N_A_27_74#_c_240_n 0.00561753f $X=1.515 $Y=1.095
+ $X2=0 $Y2=0
cc_112 N_A_177_48#_c_107_n N_A_27_74#_c_240_n 0.0142173f $X=2.61 $Y=1.985 $X2=0
+ $Y2=0
cc_113 N_A_177_48#_c_103_n N_A_27_74#_c_240_n 0.00178829f $X=1.5 $Y=1.532 $X2=0
+ $Y2=0
cc_114 N_A_177_48#_c_105_n N_A_27_74#_c_204_n 0.0118821f $X=1.5 $Y=1.765 $X2=0
+ $Y2=0
cc_115 N_A_177_48#_c_98_n N_A_27_74#_c_204_n 0.0253755f $X=1.98 $Y=1.095 $X2=0
+ $Y2=0
cc_116 N_A_177_48#_c_100_n N_A_27_74#_c_204_n 0.0177787f $X=1.515 $Y=1.095 $X2=0
+ $Y2=0
cc_117 N_A_177_48#_c_102_n N_A_27_74#_c_204_n 0.0669379f $X=2.577 $Y=1.82 $X2=0
+ $Y2=0
cc_118 N_A_177_48#_c_103_n N_A_27_74#_c_204_n 0.00265542f $X=1.5 $Y=1.532 $X2=0
+ $Y2=0
cc_119 N_A_177_48#_c_104_n N_A_27_74#_c_210_n 0.00646197f $X=1.05 $Y=1.765 $X2=0
+ $Y2=0
cc_120 N_A_177_48#_c_101_n N_A2_c_284_n 0.00465411f $X=2.465 $Y=1.095 $X2=-0.19
+ $Y2=-0.245
cc_121 N_A_177_48#_c_102_n N_A2_c_284_n 0.00220497f $X=2.577 $Y=1.82 $X2=-0.19
+ $Y2=-0.245
cc_122 N_A_177_48#_c_106_n N_A2_c_285_n 0.00884164f $X=2.61 $Y=2.695 $X2=0 $Y2=0
cc_123 N_A_177_48#_c_107_n N_A2_c_285_n 0.0129262f $X=2.61 $Y=1.985 $X2=0 $Y2=0
cc_124 N_A_177_48#_c_102_n N_A2_c_285_n 0.0053934f $X=2.577 $Y=1.82 $X2=0 $Y2=0
cc_125 N_A_177_48#_c_107_n A2 0.00318492f $X=2.61 $Y=1.985 $X2=0 $Y2=0
cc_126 N_A_177_48#_c_102_n A2 0.0287265f $X=2.577 $Y=1.82 $X2=0 $Y2=0
cc_127 N_A_177_48#_c_107_n N_A1_c_316_n 0.00316513f $X=2.61 $Y=1.985 $X2=-0.19
+ $Y2=-0.245
cc_128 N_A_177_48#_c_104_n N_VPWR_c_339_n 0.0117699f $X=1.05 $Y=1.765 $X2=0
+ $Y2=0
cc_129 N_A_177_48#_c_105_n N_VPWR_c_339_n 0.00148719f $X=1.5 $Y=1.765 $X2=0
+ $Y2=0
cc_130 N_A_177_48#_c_107_n N_VPWR_c_341_n 0.0264677f $X=2.61 $Y=1.985 $X2=0
+ $Y2=0
cc_131 N_A_177_48#_c_104_n N_VPWR_c_342_n 0.00444681f $X=1.05 $Y=1.765 $X2=0
+ $Y2=0
cc_132 N_A_177_48#_c_105_n N_VPWR_c_342_n 0.004307f $X=1.5 $Y=1.765 $X2=0 $Y2=0
cc_133 N_A_177_48#_c_106_n N_VPWR_c_343_n 0.00976219f $X=2.61 $Y=2.695 $X2=0
+ $Y2=0
cc_134 N_A_177_48#_c_104_n N_VPWR_c_345_n 0.00149535f $X=1.05 $Y=1.765 $X2=0
+ $Y2=0
cc_135 N_A_177_48#_c_105_n N_VPWR_c_345_n 0.0134232f $X=1.5 $Y=1.765 $X2=0 $Y2=0
cc_136 N_A_177_48#_c_106_n N_VPWR_c_345_n 0.0195791f $X=2.61 $Y=2.695 $X2=0
+ $Y2=0
cc_137 N_A_177_48#_c_104_n N_VPWR_c_338_n 0.00877716f $X=1.05 $Y=1.765 $X2=0
+ $Y2=0
cc_138 N_A_177_48#_c_105_n N_VPWR_c_338_n 0.00847721f $X=1.5 $Y=1.765 $X2=0
+ $Y2=0
cc_139 N_A_177_48#_c_106_n N_VPWR_c_338_n 0.0111764f $X=2.61 $Y=2.695 $X2=0
+ $Y2=0
cc_140 N_A_177_48#_M1001_g N_X_c_382_n 0.00395829f $X=0.96 $Y=0.74 $X2=0 $Y2=0
cc_141 N_A_177_48#_c_104_n N_X_c_382_n 0.00157573f $X=1.05 $Y=1.765 $X2=0 $Y2=0
cc_142 N_A_177_48#_M1009_g N_X_c_382_n 0.00162644f $X=1.39 $Y=0.74 $X2=0 $Y2=0
cc_143 N_A_177_48#_c_105_n N_X_c_382_n 0.00104603f $X=1.5 $Y=1.765 $X2=0 $Y2=0
cc_144 N_A_177_48#_c_100_n N_X_c_382_n 0.0323092f $X=1.515 $Y=1.095 $X2=0 $Y2=0
cc_145 N_A_177_48#_c_103_n N_X_c_382_n 0.0185548f $X=1.5 $Y=1.532 $X2=0 $Y2=0
cc_146 N_A_177_48#_c_104_n N_X_c_386_n 0.00645217f $X=1.05 $Y=1.765 $X2=0 $Y2=0
cc_147 N_A_177_48#_c_105_n N_X_c_386_n 0.00487049f $X=1.5 $Y=1.765 $X2=0 $Y2=0
cc_148 N_A_177_48#_c_100_n N_X_c_386_n 0.00637801f $X=1.515 $Y=1.095 $X2=0 $Y2=0
cc_149 N_A_177_48#_c_103_n N_X_c_386_n 0.00794145f $X=1.5 $Y=1.532 $X2=0 $Y2=0
cc_150 N_A_177_48#_M1001_g X 0.00957449f $X=0.96 $Y=0.74 $X2=0 $Y2=0
cc_151 N_A_177_48#_M1009_g X 0.00944938f $X=1.39 $Y=0.74 $X2=0 $Y2=0
cc_152 N_A_177_48#_c_99_n X 0.00535741f $X=2.145 $Y=0.515 $X2=0 $Y2=0
cc_153 N_A_177_48#_M1001_g X 0.00206898f $X=0.96 $Y=0.74 $X2=0 $Y2=0
cc_154 N_A_177_48#_M1009_g X 0.00364888f $X=1.39 $Y=0.74 $X2=0 $Y2=0
cc_155 N_A_177_48#_c_100_n X 0.00540984f $X=1.515 $Y=1.095 $X2=0 $Y2=0
cc_156 N_A_177_48#_c_103_n X 0.0018557f $X=1.5 $Y=1.532 $X2=0 $Y2=0
cc_157 N_A_177_48#_c_98_n N_VGND_M1009_d 9.80805e-19 $X=1.98 $Y=1.095 $X2=0
+ $Y2=0
cc_158 N_A_177_48#_c_100_n N_VGND_M1009_d 0.00270316f $X=1.515 $Y=1.095 $X2=0
+ $Y2=0
cc_159 N_A_177_48#_M1001_g N_VGND_c_417_n 0.00455916f $X=0.96 $Y=0.74 $X2=0
+ $Y2=0
cc_160 N_A_177_48#_M1009_g N_VGND_c_418_n 0.00631755f $X=1.39 $Y=0.74 $X2=0
+ $Y2=0
cc_161 N_A_177_48#_c_98_n N_VGND_c_418_n 0.00672294f $X=1.98 $Y=1.095 $X2=0
+ $Y2=0
cc_162 N_A_177_48#_c_99_n N_VGND_c_418_n 0.0323605f $X=2.145 $Y=0.515 $X2=0
+ $Y2=0
cc_163 N_A_177_48#_c_100_n N_VGND_c_418_n 0.0130147f $X=1.515 $Y=1.095 $X2=0
+ $Y2=0
cc_164 N_A_177_48#_c_103_n N_VGND_c_418_n 6.72525e-19 $X=1.5 $Y=1.532 $X2=0
+ $Y2=0
cc_165 N_A_177_48#_M1001_g N_VGND_c_422_n 0.00434272f $X=0.96 $Y=0.74 $X2=0
+ $Y2=0
cc_166 N_A_177_48#_M1009_g N_VGND_c_422_n 0.00434272f $X=1.39 $Y=0.74 $X2=0
+ $Y2=0
cc_167 N_A_177_48#_c_99_n N_VGND_c_423_n 0.0110419f $X=2.145 $Y=0.515 $X2=0
+ $Y2=0
cc_168 N_A_177_48#_M1001_g N_VGND_c_425_n 0.00821771f $X=0.96 $Y=0.74 $X2=0
+ $Y2=0
cc_169 N_A_177_48#_M1009_g N_VGND_c_425_n 0.00825283f $X=1.39 $Y=0.74 $X2=0
+ $Y2=0
cc_170 N_A_177_48#_c_99_n N_VGND_c_425_n 0.00915013f $X=2.145 $Y=0.515 $X2=0
+ $Y2=0
cc_171 N_A_177_48#_c_101_n N_A_487_74#_M1011_d 0.00196876f $X=2.465 $Y=1.095
+ $X2=-0.19 $Y2=-0.245
cc_172 N_A_177_48#_c_99_n N_A_487_74#_c_473_n 0.0182902f $X=2.145 $Y=0.515 $X2=0
+ $Y2=0
cc_173 N_A_177_48#_c_101_n N_A_487_74#_c_473_n 0.00637434f $X=2.465 $Y=1.095
+ $X2=0 $Y2=0
cc_174 N_A_27_74#_M1011_g N_A2_c_284_n 0.0315537f $X=2.36 $Y=0.74 $X2=-0.19
+ $Y2=-0.245
cc_175 N_A_27_74#_c_205_n N_A2_c_285_n 0.00843822f $X=2.385 $Y=1.765 $X2=0 $Y2=0
cc_176 N_A_27_74#_c_199_n N_A2_c_285_n 0.0199208f $X=2.285 $Y=1.35 $X2=0 $Y2=0
cc_177 N_A_27_74#_c_199_n A2 2.1389e-19 $X=2.285 $Y=1.35 $X2=0 $Y2=0
cc_178 N_A_27_74#_c_203_n N_VPWR_M1005_d 0.00120621f $X=0.71 $Y=1.95 $X2=-0.19
+ $Y2=-0.245
cc_179 N_A_27_74#_c_240_n N_VPWR_M1005_d 0.00526394f $X=1.89 $Y=2.325 $X2=-0.19
+ $Y2=-0.245
cc_180 N_A_27_74#_c_210_n N_VPWR_M1005_d 0.00660301f $X=0.28 $Y=2.115 $X2=-0.19
+ $Y2=-0.245
cc_181 N_A_27_74#_c_240_n N_VPWR_M1008_s 0.0206821f $X=1.89 $Y=2.325 $X2=0 $Y2=0
cc_182 N_A_27_74#_c_204_n N_VPWR_M1008_s 0.0153631f $X=2.055 $Y=1.515 $X2=0
+ $Y2=0
cc_183 N_A_27_74#_c_240_n N_VPWR_c_339_n 0.0102332f $X=1.89 $Y=2.325 $X2=0 $Y2=0
cc_184 N_A_27_74#_c_210_n N_VPWR_c_339_n 0.0210687f $X=0.28 $Y=2.115 $X2=0 $Y2=0
cc_185 N_A_27_74#_c_205_n N_VPWR_c_343_n 0.00481995f $X=2.385 $Y=1.765 $X2=0
+ $Y2=0
cc_186 N_A_27_74#_c_210_n N_VPWR_c_344_n 0.00671799f $X=0.28 $Y=2.115 $X2=0
+ $Y2=0
cc_187 N_A_27_74#_c_205_n N_VPWR_c_345_n 0.0114447f $X=2.385 $Y=1.765 $X2=0
+ $Y2=0
cc_188 N_A_27_74#_c_240_n N_VPWR_c_345_n 0.0503591f $X=1.89 $Y=2.325 $X2=0 $Y2=0
cc_189 N_A_27_74#_c_205_n N_VPWR_c_338_n 0.00508379f $X=2.385 $Y=1.765 $X2=0
+ $Y2=0
cc_190 N_A_27_74#_c_210_n N_VPWR_c_338_n 0.0100331f $X=0.28 $Y=2.115 $X2=0 $Y2=0
cc_191 N_A_27_74#_c_240_n N_X_M1006_d 0.00892559f $X=1.89 $Y=2.325 $X2=0 $Y2=0
cc_192 N_A_27_74#_c_203_n N_X_c_382_n 0.0412826f $X=0.71 $Y=1.95 $X2=0 $Y2=0
cc_193 N_A_27_74#_c_203_n N_X_c_386_n 0.00814288f $X=0.71 $Y=1.95 $X2=0 $Y2=0
cc_194 N_A_27_74#_c_240_n N_X_c_386_n 0.022884f $X=1.89 $Y=2.325 $X2=0 $Y2=0
cc_195 N_A_27_74#_c_204_n N_X_c_386_n 0.0092774f $X=2.055 $Y=1.515 $X2=0 $Y2=0
cc_196 N_A_27_74#_c_210_n N_X_c_386_n 0.00838529f $X=0.28 $Y=2.115 $X2=0 $Y2=0
cc_197 N_A_27_74#_c_200_n X 0.00264902f $X=0.27 $Y=0.645 $X2=0 $Y2=0
cc_198 N_A_27_74#_c_201_n X 0.0117316f $X=0.625 $Y=1.045 $X2=0 $Y2=0
cc_199 N_A_27_74#_c_201_n N_VGND_M1003_d 0.00400349f $X=0.625 $Y=1.045 $X2=-0.19
+ $Y2=-0.245
cc_200 N_A_27_74#_c_201_n N_VGND_c_417_n 0.0189182f $X=0.625 $Y=1.045 $X2=0
+ $Y2=0
cc_201 N_A_27_74#_M1011_g N_VGND_c_418_n 0.00342609f $X=2.36 $Y=0.74 $X2=0 $Y2=0
cc_202 N_A_27_74#_c_200_n N_VGND_c_420_n 0.00750773f $X=0.27 $Y=0.645 $X2=0
+ $Y2=0
cc_203 N_A_27_74#_M1011_g N_VGND_c_423_n 0.00434272f $X=2.36 $Y=0.74 $X2=0 $Y2=0
cc_204 N_A_27_74#_M1011_g N_VGND_c_425_n 0.00826366f $X=2.36 $Y=0.74 $X2=0 $Y2=0
cc_205 N_A_27_74#_c_200_n N_VGND_c_425_n 0.00854988f $X=0.27 $Y=0.645 $X2=0
+ $Y2=0
cc_206 N_A_27_74#_M1011_g N_A_487_74#_c_473_n 0.0070904f $X=2.36 $Y=0.74 $X2=0
+ $Y2=0
cc_207 N_A2_c_285_n N_A1_c_316_n 0.0647064f $X=2.835 $Y=1.765 $X2=-0.19
+ $Y2=-0.245
cc_208 N_A2_c_284_n N_A1_c_317_n 0.0256009f $X=2.79 $Y=1.22 $X2=0 $Y2=0
cc_209 A2 N_A1_c_317_n 0.00312957f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_210 N_A2_c_285_n A1 2.48878e-19 $X=2.835 $Y=1.765 $X2=0 $Y2=0
cc_211 A2 A1 0.0302901f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_212 N_A2_c_285_n N_VPWR_c_341_n 0.00367627f $X=2.835 $Y=1.765 $X2=0 $Y2=0
cc_213 N_A2_c_285_n N_VPWR_c_343_n 0.00481995f $X=2.835 $Y=1.765 $X2=0 $Y2=0
cc_214 N_A2_c_285_n N_VPWR_c_338_n 0.00508379f $X=2.835 $Y=1.765 $X2=0 $Y2=0
cc_215 N_A2_c_284_n N_VGND_c_419_n 0.00416106f $X=2.79 $Y=1.22 $X2=0 $Y2=0
cc_216 N_A2_c_284_n N_VGND_c_423_n 0.00324657f $X=2.79 $Y=1.22 $X2=0 $Y2=0
cc_217 N_A2_c_284_n N_VGND_c_425_n 0.00410881f $X=2.79 $Y=1.22 $X2=0 $Y2=0
cc_218 N_A2_c_284_n N_A_487_74#_c_479_n 0.0104597f $X=2.79 $Y=1.22 $X2=0 $Y2=0
cc_219 N_A2_c_285_n N_A_487_74#_c_479_n 8.52057e-19 $X=2.835 $Y=1.765 $X2=0
+ $Y2=0
cc_220 A2 N_A_487_74#_c_479_n 0.0215496f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_221 N_A2_c_284_n N_A_487_74#_c_473_n 0.00797172f $X=2.79 $Y=1.22 $X2=0 $Y2=0
cc_222 A2 N_A_487_74#_c_473_n 8.53117e-19 $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_223 N_A2_c_284_n N_A_487_74#_c_474_n 0.00142177f $X=2.79 $Y=1.22 $X2=0 $Y2=0
cc_224 N_A1_c_316_n N_VPWR_c_341_n 0.0279053f $X=3.345 $Y=1.765 $X2=0 $Y2=0
cc_225 A1 N_VPWR_c_341_n 0.0197435f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_226 N_A1_c_316_n N_VPWR_c_343_n 0.00443511f $X=3.345 $Y=1.765 $X2=0 $Y2=0
cc_227 N_A1_c_316_n N_VPWR_c_338_n 0.00460931f $X=3.345 $Y=1.765 $X2=0 $Y2=0
cc_228 N_A1_c_317_n N_VGND_c_419_n 0.00416106f $X=3.36 $Y=1.22 $X2=0 $Y2=0
cc_229 N_A1_c_317_n N_VGND_c_424_n 0.00324657f $X=3.36 $Y=1.22 $X2=0 $Y2=0
cc_230 N_A1_c_317_n N_VGND_c_425_n 0.00414389f $X=3.36 $Y=1.22 $X2=0 $Y2=0
cc_231 N_A1_c_317_n N_A_487_74#_c_479_n 0.0135231f $X=3.36 $Y=1.22 $X2=0 $Y2=0
cc_232 N_A1_c_317_n N_A_487_74#_c_473_n 6.42889e-19 $X=3.36 $Y=1.22 $X2=0 $Y2=0
cc_233 N_A1_c_316_n N_A_487_74#_c_474_n 0.00195015f $X=3.345 $Y=1.765 $X2=0
+ $Y2=0
cc_234 N_A1_c_317_n N_A_487_74#_c_474_n 0.010732f $X=3.36 $Y=1.22 $X2=0 $Y2=0
cc_235 A1 N_A_487_74#_c_474_n 0.0255896f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_236 X N_VGND_c_417_n 0.0269864f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_237 X N_VGND_c_418_n 0.0175734f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_238 X N_VGND_c_422_n 0.0144922f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_239 X N_VGND_c_425_n 0.0118826f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_240 N_VGND_M1002_d N_A_487_74#_c_479_n 0.00789873f $X=2.865 $Y=0.37 $X2=0
+ $Y2=0
cc_241 N_VGND_c_419_n N_A_487_74#_c_479_n 0.0235778f $X=3.075 $Y=0.335 $X2=0
+ $Y2=0
cc_242 N_VGND_c_423_n N_A_487_74#_c_479_n 0.00227739f $X=2.91 $Y=0 $X2=0 $Y2=0
cc_243 N_VGND_c_424_n N_A_487_74#_c_479_n 0.00227739f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_244 N_VGND_c_425_n N_A_487_74#_c_479_n 0.00966343f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_245 N_VGND_c_419_n N_A_487_74#_c_473_n 0.00641885f $X=3.075 $Y=0.335 $X2=0
+ $Y2=0
cc_246 N_VGND_c_423_n N_A_487_74#_c_473_n 0.0141563f $X=2.91 $Y=0 $X2=0 $Y2=0
cc_247 N_VGND_c_425_n N_A_487_74#_c_473_n 0.0117515f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_248 N_VGND_c_419_n N_A_487_74#_c_474_n 0.00641885f $X=3.075 $Y=0.335 $X2=0
+ $Y2=0
cc_249 N_VGND_c_424_n N_A_487_74#_c_474_n 0.0145323f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_250 N_VGND_c_425_n N_A_487_74#_c_474_n 0.0119861f $X=3.6 $Y=0 $X2=0 $Y2=0
