* File: sky130_fd_sc_hs__buf_4.pxi.spice
* Created: Tue Sep  1 19:56:54 2020
* 
x_PM_SKY130_FD_SC_HS__BUF_4%A_86_260# N_A_86_260#_M1004_d N_A_86_260#_M1003_d
+ N_A_86_260#_c_63_n N_A_86_260#_c_78_n N_A_86_260#_M1006_g N_A_86_260#_M1000_g
+ N_A_86_260#_c_65_n N_A_86_260#_c_79_n N_A_86_260#_M1007_g N_A_86_260#_M1001_g
+ N_A_86_260#_c_80_n N_A_86_260#_M1009_g N_A_86_260#_M1002_g N_A_86_260#_c_81_n
+ N_A_86_260#_M1010_g N_A_86_260#_M1008_g N_A_86_260#_c_69_n N_A_86_260#_c_70_n
+ N_A_86_260#_c_71_n N_A_86_260#_c_72_n N_A_86_260#_c_73_n N_A_86_260#_c_155_p
+ N_A_86_260#_c_83_n N_A_86_260#_c_74_n N_A_86_260#_c_75_n N_A_86_260#_c_76_n
+ PM_SKY130_FD_SC_HS__BUF_4%A_86_260#
x_PM_SKY130_FD_SC_HS__BUF_4%A N_A_c_185_n N_A_M1003_g N_A_c_186_n N_A_M1005_g
+ N_A_M1004_g A N_A_c_183_n N_A_c_184_n PM_SKY130_FD_SC_HS__BUF_4%A
x_PM_SKY130_FD_SC_HS__BUF_4%VPWR N_VPWR_M1006_s N_VPWR_M1007_s N_VPWR_M1010_s
+ N_VPWR_M1005_s N_VPWR_c_222_n N_VPWR_c_223_n N_VPWR_c_224_n N_VPWR_c_225_n
+ N_VPWR_c_226_n N_VPWR_c_227_n VPWR N_VPWR_c_228_n N_VPWR_c_229_n
+ N_VPWR_c_230_n N_VPWR_c_231_n N_VPWR_c_232_n N_VPWR_c_221_n
+ PM_SKY130_FD_SC_HS__BUF_4%VPWR
x_PM_SKY130_FD_SC_HS__BUF_4%X N_X_M1000_s N_X_M1002_s N_X_M1006_d N_X_M1009_d
+ N_X_c_275_n N_X_c_276_n N_X_c_277_n N_X_c_281_n N_X_c_282_n N_X_c_278_n
+ N_X_c_283_n N_X_c_279_n N_X_c_284_n X PM_SKY130_FD_SC_HS__BUF_4%X
x_PM_SKY130_FD_SC_HS__BUF_4%VGND N_VGND_M1000_d N_VGND_M1001_d N_VGND_M1008_d
+ N_VGND_c_340_n N_VGND_c_341_n N_VGND_c_342_n N_VGND_c_343_n VGND
+ N_VGND_c_344_n N_VGND_c_345_n N_VGND_c_346_n N_VGND_c_347_n N_VGND_c_348_n
+ PM_SKY130_FD_SC_HS__BUF_4%VGND
cc_1 VNB N_A_86_260#_c_63_n 0.0175041f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=1.675
cc_2 VNB N_A_86_260#_M1000_g 0.0265448f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=0.74
cc_3 VNB N_A_86_260#_c_65_n 0.00922324f $X=-0.19 $Y=-0.245 $X2=0.88 $Y2=1.375
cc_4 VNB N_A_86_260#_M1001_g 0.022504f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=0.74
cc_5 VNB N_A_86_260#_M1002_g 0.0225168f $X=-0.19 $Y=-0.245 $X2=1.565 $Y2=0.74
cc_6 VNB N_A_86_260#_M1008_g 0.0249635f $X=-0.19 $Y=-0.245 $X2=1.995 $Y2=0.74
cc_7 VNB N_A_86_260#_c_69_n 0.0145005f $X=-0.19 $Y=-0.245 $X2=0.535 $Y2=1.375
cc_8 VNB N_A_86_260#_c_70_n 0.00768954f $X=-0.19 $Y=-0.245 $X2=2.115 $Y2=1.465
cc_9 VNB N_A_86_260#_c_71_n 0.081977f $X=-0.19 $Y=-0.245 $X2=1.905 $Y2=1.465
cc_10 VNB N_A_86_260#_c_72_n 0.00389847f $X=-0.19 $Y=-0.245 $X2=2.2 $Y2=1.3
cc_11 VNB N_A_86_260#_c_73_n 0.00548705f $X=-0.19 $Y=-0.245 $X2=2.915 $Y2=1.045
cc_12 VNB N_A_86_260#_c_74_n 0.02581f $X=-0.19 $Y=-0.245 $X2=3.08 $Y2=0.515
cc_13 VNB N_A_86_260#_c_75_n 0.0249538f $X=-0.19 $Y=-0.245 $X2=3.16 $Y2=1.95
cc_14 VNB N_A_86_260#_c_76_n 0.0124806f $X=-0.19 $Y=-0.245 $X2=3.08 $Y2=1.045
cc_15 VNB N_A_M1004_g 0.0330952f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=1.765
cc_16 VNB N_A_c_183_n 0.00412911f $X=-0.19 $Y=-0.245 $X2=0.88 $Y2=1.375
cc_17 VNB N_A_c_184_n 0.0434583f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.375
cc_18 VNB N_VPWR_c_221_n 0.143779f $X=-0.19 $Y=-0.245 $X2=3.16 $Y2=1.95
cc_19 VNB N_X_c_275_n 0.00240191f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_X_c_276_n 0.00290742f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.375
cc_21 VNB N_X_c_277_n 0.00337286f $X=-0.19 $Y=-0.245 $X2=0.97 $Y2=1.765
cc_22 VNB N_X_c_278_n 0.00542414f $X=-0.19 $Y=-0.245 $X2=1.42 $Y2=2.4
cc_23 VNB N_X_c_279_n 0.00240191f $X=-0.19 $Y=-0.245 $X2=1.995 $Y2=0.74
cc_24 VNB N_VGND_c_340_n 0.0122168f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=2.4
cc_25 VNB N_VGND_c_341_n 0.0376574f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=1.3
cc_26 VNB N_VGND_c_342_n 0.00830803f $X=-0.19 $Y=-0.245 $X2=0.88 $Y2=1.375
cc_27 VNB N_VGND_c_343_n 0.0187266f $X=-0.19 $Y=-0.245 $X2=0.97 $Y2=1.765
cc_28 VNB N_VGND_c_344_n 0.0186948f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=0.74
cc_29 VNB N_VGND_c_345_n 0.0191816f $X=-0.19 $Y=-0.245 $X2=1.565 $Y2=0.74
cc_30 VNB N_VGND_c_346_n 0.204744f $X=-0.19 $Y=-0.245 $X2=1.565 $Y2=0.74
cc_31 VNB N_VGND_c_347_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=1.995 $Y2=0.74
cc_32 VNB N_VGND_c_348_n 0.0243944f $X=-0.19 $Y=-0.245 $X2=2.115 $Y2=1.465
cc_33 VPB N_A_86_260#_c_63_n 0.00117364f $X=-0.19 $Y=1.66 $X2=0.52 $Y2=1.675
cc_34 VPB N_A_86_260#_c_78_n 0.0274181f $X=-0.19 $Y=1.66 $X2=0.52 $Y2=1.765
cc_35 VPB N_A_86_260#_c_79_n 0.0147047f $X=-0.19 $Y=1.66 $X2=0.97 $Y2=1.765
cc_36 VPB N_A_86_260#_c_80_n 0.0147155f $X=-0.19 $Y=1.66 $X2=1.42 $Y2=1.765
cc_37 VPB N_A_86_260#_c_81_n 0.0171739f $X=-0.19 $Y=1.66 $X2=1.87 $Y2=1.765
cc_38 VPB N_A_86_260#_c_71_n 0.0198854f $X=-0.19 $Y=1.66 $X2=1.905 $Y2=1.465
cc_39 VPB N_A_86_260#_c_83_n 0.0105449f $X=-0.19 $Y=1.66 $X2=3.075 $Y2=2.075
cc_40 VPB N_A_86_260#_c_75_n 0.0122801f $X=-0.19 $Y=1.66 $X2=3.16 $Y2=1.95
cc_41 VPB N_A_c_185_n 0.0162849f $X=-0.19 $Y=1.66 $X2=2.94 $Y2=0.37
cc_42 VPB N_A_c_186_n 0.0169025f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_43 VPB N_A_c_183_n 0.00336439f $X=-0.19 $Y=1.66 $X2=0.88 $Y2=1.375
cc_44 VPB N_A_c_184_n 0.0213107f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.375
cc_45 VPB N_VPWR_c_222_n 0.0124891f $X=-0.19 $Y=1.66 $X2=0.565 $Y2=0.74
cc_46 VPB N_VPWR_c_223_n 0.0651331f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_47 VPB N_VPWR_c_224_n 0.00261791f $X=-0.19 $Y=1.66 $X2=0.995 $Y2=1.3
cc_48 VPB N_VPWR_c_225_n 0.0125404f $X=-0.19 $Y=1.66 $X2=1.42 $Y2=1.765
cc_49 VPB N_VPWR_c_226_n 0.0121909f $X=-0.19 $Y=1.66 $X2=1.565 $Y2=0.74
cc_50 VPB N_VPWR_c_227_n 0.0392892f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_51 VPB N_VPWR_c_228_n 0.0164074f $X=-0.19 $Y=1.66 $X2=1.995 $Y2=1.3
cc_52 VPB N_VPWR_c_229_n 0.0164465f $X=-0.19 $Y=1.66 $X2=2.115 $Y2=1.465
cc_53 VPB N_VPWR_c_230_n 0.0207798f $X=-0.19 $Y=1.66 $X2=1.905 $Y2=1.465
cc_54 VPB N_VPWR_c_231_n 0.00601644f $X=-0.19 $Y=1.66 $X2=2.63 $Y2=2.115
cc_55 VPB N_VPWR_c_232_n 0.00614127f $X=-0.19 $Y=1.66 $X2=3.08 $Y2=0.515
cc_56 VPB N_VPWR_c_221_n 0.0787651f $X=-0.19 $Y=1.66 $X2=3.16 $Y2=1.95
cc_57 VPB N_X_c_277_n 0.00280927f $X=-0.19 $Y=1.66 $X2=0.97 $Y2=1.765
cc_58 VPB N_X_c_281_n 0.00185483f $X=-0.19 $Y=1.66 $X2=0.995 $Y2=1.3
cc_59 VPB N_X_c_282_n 0.00446252f $X=-0.19 $Y=1.66 $X2=1.42 $Y2=1.765
cc_60 VPB N_X_c_283_n 0.00180921f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_61 VPB N_X_c_284_n 4.21926e-19 $X=-0.19 $Y=1.66 $X2=0.535 $Y2=1.375
cc_62 N_A_86_260#_c_81_n N_A_c_185_n 0.0137311f $X=1.87 $Y=1.765 $X2=-0.19
+ $Y2=-0.245
cc_63 N_A_86_260#_c_83_n N_A_c_185_n 0.00381685f $X=3.075 $Y=2.075 $X2=-0.19
+ $Y2=-0.245
cc_64 N_A_86_260#_c_83_n N_A_c_186_n 0.0176218f $X=3.075 $Y=2.075 $X2=0 $Y2=0
cc_65 N_A_86_260#_c_75_n N_A_c_186_n 0.00623977f $X=3.16 $Y=1.95 $X2=0 $Y2=0
cc_66 N_A_86_260#_M1008_g N_A_M1004_g 0.0127822f $X=1.995 $Y=0.74 $X2=0 $Y2=0
cc_67 N_A_86_260#_c_70_n N_A_M1004_g 0.00105416f $X=2.115 $Y=1.465 $X2=0 $Y2=0
cc_68 N_A_86_260#_c_72_n N_A_M1004_g 0.00275276f $X=2.2 $Y=1.3 $X2=0 $Y2=0
cc_69 N_A_86_260#_c_73_n N_A_M1004_g 0.0131472f $X=2.915 $Y=1.045 $X2=0 $Y2=0
cc_70 N_A_86_260#_c_74_n N_A_M1004_g 0.0174462f $X=3.08 $Y=0.515 $X2=0 $Y2=0
cc_71 N_A_86_260#_c_75_n N_A_M1004_g 0.00778767f $X=3.16 $Y=1.95 $X2=0 $Y2=0
cc_72 N_A_86_260#_c_76_n N_A_M1004_g 0.00204635f $X=3.08 $Y=1.045 $X2=0 $Y2=0
cc_73 N_A_86_260#_c_70_n N_A_c_183_n 0.0192045f $X=2.115 $Y=1.465 $X2=0 $Y2=0
cc_74 N_A_86_260#_c_71_n N_A_c_183_n 7.75012e-19 $X=1.905 $Y=1.465 $X2=0 $Y2=0
cc_75 N_A_86_260#_c_73_n N_A_c_183_n 0.0237625f $X=2.915 $Y=1.045 $X2=0 $Y2=0
cc_76 N_A_86_260#_c_83_n N_A_c_183_n 0.0275642f $X=3.075 $Y=2.075 $X2=0 $Y2=0
cc_77 N_A_86_260#_c_75_n N_A_c_183_n 0.0326295f $X=3.16 $Y=1.95 $X2=0 $Y2=0
cc_78 N_A_86_260#_c_70_n N_A_c_184_n 0.00188928f $X=2.115 $Y=1.465 $X2=0 $Y2=0
cc_79 N_A_86_260#_c_71_n N_A_c_184_n 0.0140442f $X=1.905 $Y=1.465 $X2=0 $Y2=0
cc_80 N_A_86_260#_c_73_n N_A_c_184_n 0.00821934f $X=2.915 $Y=1.045 $X2=0 $Y2=0
cc_81 N_A_86_260#_c_83_n N_A_c_184_n 0.0012403f $X=3.075 $Y=2.075 $X2=0 $Y2=0
cc_82 N_A_86_260#_c_75_n N_A_c_184_n 0.0101252f $X=3.16 $Y=1.95 $X2=0 $Y2=0
cc_83 N_A_86_260#_c_76_n N_A_c_184_n 2.15716e-19 $X=3.08 $Y=1.045 $X2=0 $Y2=0
cc_84 N_A_86_260#_c_83_n N_VPWR_M1005_s 0.00765411f $X=3.075 $Y=2.075 $X2=0
+ $Y2=0
cc_85 N_A_86_260#_c_75_n N_VPWR_M1005_s 0.00193837f $X=3.16 $Y=1.95 $X2=0 $Y2=0
cc_86 N_A_86_260#_c_78_n N_VPWR_c_223_n 0.0194655f $X=0.52 $Y=1.765 $X2=0 $Y2=0
cc_87 N_A_86_260#_c_79_n N_VPWR_c_223_n 6.87578e-19 $X=0.97 $Y=1.765 $X2=0 $Y2=0
cc_88 N_A_86_260#_c_78_n N_VPWR_c_224_n 5.75642e-19 $X=0.52 $Y=1.765 $X2=0 $Y2=0
cc_89 N_A_86_260#_c_79_n N_VPWR_c_224_n 0.0150018f $X=0.97 $Y=1.765 $X2=0 $Y2=0
cc_90 N_A_86_260#_c_80_n N_VPWR_c_224_n 0.0150993f $X=1.42 $Y=1.765 $X2=0 $Y2=0
cc_91 N_A_86_260#_c_81_n N_VPWR_c_224_n 5.81581e-19 $X=1.87 $Y=1.765 $X2=0 $Y2=0
cc_92 N_A_86_260#_c_80_n N_VPWR_c_225_n 6.87578e-19 $X=1.42 $Y=1.765 $X2=0 $Y2=0
cc_93 N_A_86_260#_c_81_n N_VPWR_c_225_n 0.0176941f $X=1.87 $Y=1.765 $X2=0 $Y2=0
cc_94 N_A_86_260#_c_70_n N_VPWR_c_225_n 0.02681f $X=2.115 $Y=1.465 $X2=0 $Y2=0
cc_95 N_A_86_260#_c_71_n N_VPWR_c_225_n 0.00343701f $X=1.905 $Y=1.465 $X2=0
+ $Y2=0
cc_96 N_A_86_260#_c_83_n N_VPWR_c_225_n 0.0176744f $X=3.075 $Y=2.075 $X2=0 $Y2=0
cc_97 N_A_86_260#_c_83_n N_VPWR_c_227_n 0.0236247f $X=3.075 $Y=2.075 $X2=0 $Y2=0
cc_98 N_A_86_260#_c_78_n N_VPWR_c_228_n 0.00413917f $X=0.52 $Y=1.765 $X2=0 $Y2=0
cc_99 N_A_86_260#_c_79_n N_VPWR_c_228_n 0.00413917f $X=0.97 $Y=1.765 $X2=0 $Y2=0
cc_100 N_A_86_260#_c_80_n N_VPWR_c_229_n 0.00413917f $X=1.42 $Y=1.765 $X2=0
+ $Y2=0
cc_101 N_A_86_260#_c_81_n N_VPWR_c_229_n 0.00413917f $X=1.87 $Y=1.765 $X2=0
+ $Y2=0
cc_102 N_A_86_260#_c_78_n N_VPWR_c_221_n 0.00817726f $X=0.52 $Y=1.765 $X2=0
+ $Y2=0
cc_103 N_A_86_260#_c_79_n N_VPWR_c_221_n 0.00817726f $X=0.97 $Y=1.765 $X2=0
+ $Y2=0
cc_104 N_A_86_260#_c_80_n N_VPWR_c_221_n 0.00817726f $X=1.42 $Y=1.765 $X2=0
+ $Y2=0
cc_105 N_A_86_260#_c_81_n N_VPWR_c_221_n 0.00817726f $X=1.87 $Y=1.765 $X2=0
+ $Y2=0
cc_106 N_A_86_260#_M1000_g N_X_c_275_n 0.00767507f $X=0.565 $Y=0.74 $X2=0 $Y2=0
cc_107 N_A_86_260#_M1001_g N_X_c_275_n 0.00916694f $X=0.995 $Y=0.74 $X2=0 $Y2=0
cc_108 N_A_86_260#_M1002_g N_X_c_275_n 6.18925e-19 $X=1.565 $Y=0.74 $X2=0 $Y2=0
cc_109 N_A_86_260#_M1000_g N_X_c_276_n 0.0154604f $X=0.565 $Y=0.74 $X2=0 $Y2=0
cc_110 N_A_86_260#_c_65_n N_X_c_276_n 0.00719234f $X=0.88 $Y=1.375 $X2=0 $Y2=0
cc_111 N_A_86_260#_M1001_g N_X_c_276_n 0.00546031f $X=0.995 $Y=0.74 $X2=0 $Y2=0
cc_112 N_A_86_260#_c_69_n N_X_c_276_n 0.00651236f $X=0.535 $Y=1.375 $X2=0 $Y2=0
cc_113 N_A_86_260#_c_70_n N_X_c_276_n 0.00679785f $X=2.115 $Y=1.465 $X2=0 $Y2=0
cc_114 N_A_86_260#_c_63_n N_X_c_277_n 0.00761156f $X=0.52 $Y=1.675 $X2=0 $Y2=0
cc_115 N_A_86_260#_c_78_n N_X_c_277_n 8.14381e-19 $X=0.52 $Y=1.765 $X2=0 $Y2=0
cc_116 N_A_86_260#_c_65_n N_X_c_277_n 0.00499189f $X=0.88 $Y=1.375 $X2=0 $Y2=0
cc_117 N_A_86_260#_c_79_n N_X_c_277_n 8.19586e-19 $X=0.97 $Y=1.765 $X2=0 $Y2=0
cc_118 N_A_86_260#_c_70_n N_X_c_277_n 0.014004f $X=2.115 $Y=1.465 $X2=0 $Y2=0
cc_119 N_A_86_260#_c_71_n N_X_c_277_n 0.00503443f $X=1.905 $Y=1.465 $X2=0 $Y2=0
cc_120 N_A_86_260#_c_78_n N_X_c_281_n 0.00351076f $X=0.52 $Y=1.765 $X2=0 $Y2=0
cc_121 N_A_86_260#_c_79_n N_X_c_281_n 0.00627021f $X=0.97 $Y=1.765 $X2=0 $Y2=0
cc_122 N_A_86_260#_c_79_n N_X_c_282_n 0.0152314f $X=0.97 $Y=1.765 $X2=0 $Y2=0
cc_123 N_A_86_260#_c_80_n N_X_c_282_n 0.0130213f $X=1.42 $Y=1.765 $X2=0 $Y2=0
cc_124 N_A_86_260#_c_81_n N_X_c_282_n 0.00137593f $X=1.87 $Y=1.765 $X2=0 $Y2=0
cc_125 N_A_86_260#_c_70_n N_X_c_282_n 0.0513154f $X=2.115 $Y=1.465 $X2=0 $Y2=0
cc_126 N_A_86_260#_c_71_n N_X_c_282_n 0.0143964f $X=1.905 $Y=1.465 $X2=0 $Y2=0
cc_127 N_A_86_260#_M1001_g N_X_c_278_n 0.0135268f $X=0.995 $Y=0.74 $X2=0 $Y2=0
cc_128 N_A_86_260#_M1002_g N_X_c_278_n 0.0128445f $X=1.565 $Y=0.74 $X2=0 $Y2=0
cc_129 N_A_86_260#_M1008_g N_X_c_278_n 0.00240508f $X=1.995 $Y=0.74 $X2=0 $Y2=0
cc_130 N_A_86_260#_c_70_n N_X_c_278_n 0.0687837f $X=2.115 $Y=1.465 $X2=0 $Y2=0
cc_131 N_A_86_260#_c_71_n N_X_c_278_n 0.00811464f $X=1.905 $Y=1.465 $X2=0 $Y2=0
cc_132 N_A_86_260#_c_155_p N_X_c_278_n 0.00808483f $X=2.285 $Y=1.045 $X2=0 $Y2=0
cc_133 N_A_86_260#_c_80_n N_X_c_283_n 0.00624195f $X=1.42 $Y=1.765 $X2=0 $Y2=0
cc_134 N_A_86_260#_c_81_n N_X_c_283_n 0.00348939f $X=1.87 $Y=1.765 $X2=0 $Y2=0
cc_135 N_A_86_260#_M1001_g N_X_c_279_n 6.18925e-19 $X=0.995 $Y=0.74 $X2=0 $Y2=0
cc_136 N_A_86_260#_M1002_g N_X_c_279_n 0.00916694f $X=1.565 $Y=0.74 $X2=0 $Y2=0
cc_137 N_A_86_260#_M1008_g N_X_c_279_n 0.0167949f $X=1.995 $Y=0.74 $X2=0 $Y2=0
cc_138 N_A_86_260#_c_78_n N_X_c_284_n 0.00137593f $X=0.52 $Y=1.765 $X2=0 $Y2=0
cc_139 N_A_86_260#_c_73_n N_VGND_M1008_d 0.00863822f $X=2.915 $Y=1.045 $X2=0
+ $Y2=0
cc_140 N_A_86_260#_c_155_p N_VGND_M1008_d 0.00351113f $X=2.285 $Y=1.045 $X2=0
+ $Y2=0
cc_141 N_A_86_260#_M1000_g N_VGND_c_341_n 0.0161039f $X=0.565 $Y=0.74 $X2=0
+ $Y2=0
cc_142 N_A_86_260#_c_69_n N_VGND_c_341_n 3.33459e-19 $X=0.535 $Y=1.375 $X2=0
+ $Y2=0
cc_143 N_A_86_260#_M1001_g N_VGND_c_342_n 0.00454042f $X=0.995 $Y=0.74 $X2=0
+ $Y2=0
cc_144 N_A_86_260#_M1002_g N_VGND_c_342_n 0.00454042f $X=1.565 $Y=0.74 $X2=0
+ $Y2=0
cc_145 N_A_86_260#_M1002_g N_VGND_c_343_n 0.00434272f $X=1.565 $Y=0.74 $X2=0
+ $Y2=0
cc_146 N_A_86_260#_M1008_g N_VGND_c_343_n 0.00434272f $X=1.995 $Y=0.74 $X2=0
+ $Y2=0
cc_147 N_A_86_260#_M1000_g N_VGND_c_344_n 0.00434272f $X=0.565 $Y=0.74 $X2=0
+ $Y2=0
cc_148 N_A_86_260#_M1001_g N_VGND_c_344_n 0.00434272f $X=0.995 $Y=0.74 $X2=0
+ $Y2=0
cc_149 N_A_86_260#_c_74_n N_VGND_c_345_n 0.0145639f $X=3.08 $Y=0.515 $X2=0 $Y2=0
cc_150 N_A_86_260#_M1000_g N_VGND_c_346_n 0.00823934f $X=0.565 $Y=0.74 $X2=0
+ $Y2=0
cc_151 N_A_86_260#_M1001_g N_VGND_c_346_n 0.00821294f $X=0.995 $Y=0.74 $X2=0
+ $Y2=0
cc_152 N_A_86_260#_M1002_g N_VGND_c_346_n 0.00821294f $X=1.565 $Y=0.74 $X2=0
+ $Y2=0
cc_153 N_A_86_260#_M1008_g N_VGND_c_346_n 0.00822986f $X=1.995 $Y=0.74 $X2=0
+ $Y2=0
cc_154 N_A_86_260#_c_74_n N_VGND_c_346_n 0.0119984f $X=3.08 $Y=0.515 $X2=0 $Y2=0
cc_155 N_A_86_260#_M1008_g N_VGND_c_348_n 0.00543794f $X=1.995 $Y=0.74 $X2=0
+ $Y2=0
cc_156 N_A_86_260#_c_73_n N_VGND_c_348_n 0.0251789f $X=2.915 $Y=1.045 $X2=0
+ $Y2=0
cc_157 N_A_86_260#_c_155_p N_VGND_c_348_n 0.00982229f $X=2.285 $Y=1.045 $X2=0
+ $Y2=0
cc_158 N_A_86_260#_c_74_n N_VGND_c_348_n 0.013254f $X=3.08 $Y=0.515 $X2=0 $Y2=0
cc_159 N_A_c_185_n N_VPWR_c_225_n 0.0173587f $X=2.405 $Y=1.765 $X2=0 $Y2=0
cc_160 N_A_c_185_n N_VPWR_c_227_n 0.00134042f $X=2.405 $Y=1.765 $X2=0 $Y2=0
cc_161 N_A_c_186_n N_VPWR_c_227_n 0.0114161f $X=2.855 $Y=1.765 $X2=0 $Y2=0
cc_162 N_A_c_185_n N_VPWR_c_230_n 0.00402388f $X=2.405 $Y=1.765 $X2=0 $Y2=0
cc_163 N_A_c_186_n N_VPWR_c_230_n 0.00361294f $X=2.855 $Y=1.765 $X2=0 $Y2=0
cc_164 N_A_c_185_n N_VPWR_c_221_n 0.00462577f $X=2.405 $Y=1.765 $X2=0 $Y2=0
cc_165 N_A_c_186_n N_VPWR_c_221_n 0.00419404f $X=2.855 $Y=1.765 $X2=0 $Y2=0
cc_166 N_A_M1004_g N_VGND_c_345_n 0.00434272f $X=2.865 $Y=0.74 $X2=0 $Y2=0
cc_167 N_A_M1004_g N_VGND_c_346_n 0.00826644f $X=2.865 $Y=0.74 $X2=0 $Y2=0
cc_168 N_A_M1004_g N_VGND_c_348_n 0.00703669f $X=2.865 $Y=0.74 $X2=0 $Y2=0
cc_169 N_VPWR_c_223_n N_X_c_281_n 0.0659251f $X=0.295 $Y=1.985 $X2=0 $Y2=0
cc_170 N_VPWR_c_224_n N_X_c_281_n 0.0559381f $X=1.195 $Y=2.225 $X2=0 $Y2=0
cc_171 N_VPWR_c_228_n N_X_c_281_n 0.00771942f $X=1.03 $Y=3.33 $X2=0 $Y2=0
cc_172 N_VPWR_c_221_n N_X_c_281_n 0.00638947f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_173 N_VPWR_M1007_s N_X_c_282_n 0.00197722f $X=1.045 $Y=1.84 $X2=0 $Y2=0
cc_174 N_VPWR_c_224_n N_X_c_282_n 0.0171813f $X=1.195 $Y=2.225 $X2=0 $Y2=0
cc_175 N_VPWR_c_225_n N_X_c_282_n 0.010961f $X=2.095 $Y=1.985 $X2=0 $Y2=0
cc_176 N_VPWR_c_224_n N_X_c_283_n 0.0547423f $X=1.195 $Y=2.225 $X2=0 $Y2=0
cc_177 N_VPWR_c_225_n N_X_c_283_n 0.0657834f $X=2.095 $Y=1.985 $X2=0 $Y2=0
cc_178 N_VPWR_c_229_n N_X_c_283_n 0.00749631f $X=1.93 $Y=3.33 $X2=0 $Y2=0
cc_179 N_VPWR_c_221_n N_X_c_283_n 0.0062048f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_180 N_VPWR_c_223_n N_X_c_284_n 0.010961f $X=0.295 $Y=1.985 $X2=0 $Y2=0
cc_181 N_X_c_278_n N_VGND_M1001_d 0.00374767f $X=1.615 $Y=1.045 $X2=0 $Y2=0
cc_182 N_X_c_275_n N_VGND_c_341_n 0.0236416f $X=0.78 $Y=0.515 $X2=0 $Y2=0
cc_183 N_X_c_275_n N_VGND_c_342_n 0.0173003f $X=0.78 $Y=0.515 $X2=0 $Y2=0
cc_184 N_X_c_278_n N_VGND_c_342_n 0.0248957f $X=1.615 $Y=1.045 $X2=0 $Y2=0
cc_185 N_X_c_279_n N_VGND_c_342_n 0.0173003f $X=1.78 $Y=0.515 $X2=0 $Y2=0
cc_186 N_X_c_279_n N_VGND_c_343_n 0.0144922f $X=1.78 $Y=0.515 $X2=0 $Y2=0
cc_187 N_X_c_275_n N_VGND_c_344_n 0.0144922f $X=0.78 $Y=0.515 $X2=0 $Y2=0
cc_188 N_X_c_275_n N_VGND_c_346_n 0.0118826f $X=0.78 $Y=0.515 $X2=0 $Y2=0
cc_189 N_X_c_279_n N_VGND_c_346_n 0.0118826f $X=1.78 $Y=0.515 $X2=0 $Y2=0
cc_190 N_X_c_279_n N_VGND_c_348_n 0.013254f $X=1.78 $Y=0.515 $X2=0 $Y2=0
