* File: sky130_fd_sc_hs__edfxbp_1.pex.spice
* Created: Tue Sep  1 20:04:21 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HS__EDFXBP_1%D 2 4 5 7 10 12 13 17 18 21
c44 21 0 4.29314e-20 $X=0.59 $Y=1.825
r45 21 23 40.7132 $w=3.4e-07 $l=1.65e-07 $layer=POLY_cond $X=0.585 $Y=1.825
+ $X2=0.585 $Y2=1.99
r46 21 22 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=0.59
+ $Y=1.825 $X2=0.59 $Y2=1.825
r47 17 19 46.3065 $w=3.4e-07 $l=1.65e-07 $layer=POLY_cond $X=0.585 $Y=1.145
+ $X2=0.585 $Y2=0.98
r48 17 18 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=0.59
+ $Y=1.145 $X2=0.59 $Y2=1.145
r49 13 22 4.49734 $w=4.08e-07 $l=1.6e-07 $layer=LI1_cond $X=0.63 $Y=1.665
+ $X2=0.63 $Y2=1.825
r50 12 13 10.4001 $w=4.08e-07 $l=3.7e-07 $layer=LI1_cond $X=0.63 $Y=1.295
+ $X2=0.63 $Y2=1.665
r51 12 18 4.21625 $w=4.08e-07 $l=1.5e-07 $layer=LI1_cond $X=0.63 $Y=1.295
+ $X2=0.63 $Y2=1.145
r52 10 19 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=0.65 $Y=0.58 $X2=0.65
+ $Y2=0.98
r53 5 7 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=0.505 $Y=2.465
+ $X2=0.505 $Y2=2.75
r54 4 5 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=0.505 $Y=2.375 $X2=0.505
+ $Y2=2.465
r55 4 23 149.653 $w=1.8e-07 $l=3.85e-07 $layer=POLY_cond $X=0.505 $Y=2.375
+ $X2=0.505 $Y2=1.99
r56 2 21 0.848592 $w=3.4e-07 $l=5e-09 $layer=POLY_cond $X=0.585 $Y=1.82
+ $X2=0.585 $Y2=1.825
r57 1 17 0.848592 $w=3.4e-07 $l=5e-09 $layer=POLY_cond $X=0.585 $Y=1.15
+ $X2=0.585 $Y2=1.145
r58 1 2 113.711 $w=3.4e-07 $l=6.7e-07 $layer=POLY_cond $X=0.585 $Y=1.15
+ $X2=0.585 $Y2=1.82
.ends

.subckt PM_SKY130_FD_SC_HS__EDFXBP_1%A_161_446# 1 2 7 9 12 22 23 24 25 26 27 30
+ 34 36 40 41 43
c107 40 0 1.52853e-19 $X=2.5 $Y=1.145
c108 27 0 4.29314e-20 $X=1.335 $Y=2.035
c109 7 0 1.45922e-19 $X=0.895 $Y=2.465
r110 40 41 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.5
+ $Y=1.145 $X2=2.5 $Y2=1.145
r111 38 40 28.1126 $w=3.28e-07 $l=8.05e-07 $layer=LI1_cond $X=2.5 $Y=1.95
+ $X2=2.5 $Y2=1.145
r112 37 43 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.885 $Y=2.035
+ $X2=1.8 $Y2=2.035
r113 36 38 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.335 $Y=2.035
+ $X2=2.5 $Y2=1.95
r114 36 37 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=2.335 $Y=2.035
+ $X2=1.885 $Y2=2.035
r115 32 43 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.8 $Y=2.12 $X2=1.8
+ $Y2=2.035
r116 32 34 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=1.8 $Y=2.12
+ $X2=1.8 $Y2=2.505
r117 28 30 15.311 $w=3.48e-07 $l=4.65e-07 $layer=LI1_cond $X=1.825 $Y=1.11
+ $X2=1.825 $Y2=0.645
r118 26 43 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.715 $Y=2.035
+ $X2=1.8 $Y2=2.035
r119 26 27 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=1.715 $Y=2.035
+ $X2=1.335 $Y2=2.035
r120 24 28 7.93686 $w=1.7e-07 $l=2.13307e-07 $layer=LI1_cond $X=1.65 $Y=1.195
+ $X2=1.825 $Y2=1.11
r121 24 25 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=1.65 $Y=1.195
+ $X2=1.335 $Y2=1.195
r122 22 23 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.17
+ $Y=1.615 $X2=1.17 $Y2=1.615
r123 20 27 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.17 $Y=1.95
+ $X2=1.335 $Y2=2.035
r124 20 22 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=1.17 $Y=1.95
+ $X2=1.17 $Y2=1.615
r125 19 25 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.17 $Y=1.28
+ $X2=1.335 $Y2=1.195
r126 19 22 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=1.17 $Y=1.28
+ $X2=1.17 $Y2=1.615
r127 18 41 41.8716 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.5 $Y=0.98
+ $X2=2.5 $Y2=1.145
r128 16 23 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.17 $Y=1.955
+ $X2=1.17 $Y2=1.615
r129 12 18 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=2.56 $Y=0.58 $X2=2.56
+ $Y2=0.98
r130 7 16 50.7854 $w=2.61e-07 $l=6.32732e-07 $layer=POLY_cond $X=0.895 $Y=2.465
+ $X2=1.17 $Y2=1.955
r131 7 9 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=0.895 $Y=2.465
+ $X2=0.895 $Y2=2.75
r132 2 34 600 $w=1.7e-07 $l=2.67862e-07 $layer=licon1_PDIFF $count=1 $X=1.655
+ $Y=2.3 $X2=1.8 $Y2=2.505
r133 1 30 182 $w=1.7e-07 $l=3.43875e-07 $layer=licon1_NDIFF $count=1 $X=1.67
+ $Y=0.37 $X2=1.825 $Y2=0.645
.ends

.subckt PM_SKY130_FD_SC_HS__EDFXBP_1%DE 1 3 4 5 7 8 10 12 13 15 16 19 20 22 23
+ 24 26
c86 20 0 9.62868e-20 $X=2.705 $Y=2.445
c87 16 0 2.45649e-19 $X=2.44 $Y=1.965
c88 8 0 1.52853e-19 $X=1.975 $Y=0.94
r89 29 31 37.1586 $w=4.54e-07 $l=3.5e-07 $layer=POLY_cond $X=1.845 $Y=1.615
+ $X2=1.845 $Y2=1.965
r90 26 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.74
+ $Y=1.615 $X2=1.74 $Y2=1.615
r91 24 25 50.3187 $w=1.82e-07 $l=1.9e-07 $layer=POLY_cond $X=2.515 $Y=2.337
+ $X2=2.705 $Y2=2.337
r92 20 25 7.39479 $w=1.5e-07 $l=1.08e-07 $layer=POLY_cond $X=2.705 $Y=2.445
+ $X2=2.705 $Y2=2.337
r93 20 22 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=2.705 $Y=2.445
+ $X2=2.705 $Y2=2.73
r94 19 24 7.39479 $w=1.5e-07 $l=1.07e-07 $layer=POLY_cond $X=2.515 $Y=2.23
+ $X2=2.515 $Y2=2.337
r95 18 19 97.4255 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=2.515 $Y=2.04
+ $X2=2.515 $Y2=2.23
r96 17 31 28.9869 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=2.115 $Y=1.965
+ $X2=1.845 $Y2=1.965
r97 16 18 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.44 $Y=1.965
+ $X2=2.515 $Y2=2.04
r98 16 17 166.649 $w=1.5e-07 $l=3.25e-07 $layer=POLY_cond $X=2.44 $Y=1.965
+ $X2=2.115 $Y2=1.965
r99 13 15 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=2.05 $Y=0.865
+ $X2=2.05 $Y2=0.58
r100 10 31 50.8617 $w=4.54e-07 $l=3.38231e-07 $layer=POLY_cond $X=2.025 $Y=2.225
+ $X2=1.845 $Y2=1.965
r101 10 12 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=2.025 $Y=2.225
+ $X2=2.025 $Y2=2.62
r102 9 23 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.725 $Y=0.94
+ $X2=1.65 $Y2=0.94
r103 8 13 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.975 $Y=0.94
+ $X2=2.05 $Y2=0.865
r104 8 9 128.191 $w=1.5e-07 $l=2.5e-07 $layer=POLY_cond $X=1.975 $Y=0.94
+ $X2=1.725 $Y2=0.94
r105 7 29 40.7758 $w=4.54e-07 $l=2.64953e-07 $layer=POLY_cond $X=1.65 $Y=1.45
+ $X2=1.845 $Y2=1.615
r106 6 23 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.65 $Y=1.015
+ $X2=1.65 $Y2=0.94
r107 6 7 223.053 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.65 $Y=1.015
+ $X2=1.65 $Y2=1.45
r108 4 23 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.575 $Y=0.94
+ $X2=1.65 $Y2=0.94
r109 4 5 235.872 $w=1.5e-07 $l=4.6e-07 $layer=POLY_cond $X=1.575 $Y=0.94
+ $X2=1.115 $Y2=0.94
r110 1 5 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.04 $Y=0.865
+ $X2=1.115 $Y2=0.94
r111 1 3 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=1.04 $Y=0.865 $X2=1.04
+ $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_HS__EDFXBP_1%A_575_48# 1 2 9 12 13 15 16 18 21 23 25 28
+ 32 39 41 42 44 45 47 53 54 55 61 66 67 69 71 73 81
c232 71 0 1.37757e-19 $X=3.04 $Y=1.99
c233 67 0 1.15042e-19 $X=3.04 $Y=1.145
c234 54 0 1.73187e-19 $X=12.095 $Y=1.665
c235 32 0 7.23051e-20 $X=12.155 $Y=1.922
c236 23 0 7.45843e-20 $X=13.85 $Y=1.765
r237 72 73 2.08357 $w=3.47e-07 $l=1.5e-08 $layer=POLY_cond $X=11.435 $Y=1.932
+ $X2=11.45 $Y2=1.932
r238 69 71 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.04 $Y=1.825
+ $X2=3.04 $Y2=1.99
r239 66 69 118.906 $w=3.3e-07 $l=6.8e-07 $layer=POLY_cond $X=3.04 $Y=1.145
+ $X2=3.04 $Y2=1.825
r240 66 67 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=3.04
+ $Y=1.145 $X2=3.04 $Y2=1.145
r241 62 81 40.1609 $w=3.28e-07 $l=1.15e-06 $layer=LI1_cond $X=12.32 $Y=1.665
+ $X2=12.32 $Y2=0.515
r242 61 62 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.24 $Y=1.665
+ $X2=12.24 $Y2=1.665
r243 58 67 18.1597 $w=3.28e-07 $l=5.2e-07 $layer=LI1_cond $X=3.04 $Y=1.665
+ $X2=3.04 $Y2=1.145
r244 58 69 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=3.04
+ $Y=1.825 $X2=3.04 $Y2=1.825
r245 57 58 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=1.665
+ $X2=3.12 $Y2=1.665
r246 55 57 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.265 $Y=1.665
+ $X2=3.12 $Y2=1.665
r247 54 61 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=12.095 $Y=1.665
+ $X2=12.24 $Y2=1.665
r248 54 55 10.9282 $w=1.4e-07 $l=8.83e-06 $layer=MET1_cond $X=12.095 $Y=1.665
+ $X2=3.265 $Y2=1.665
r249 51 62 2.09535 $w=3.28e-07 $l=6e-08 $layer=LI1_cond $X=12.32 $Y=1.725
+ $X2=12.32 $Y2=1.665
r250 51 53 6.62588 $w=2.9e-07 $l=1.65e-07 $layer=LI1_cond $X=12.32 $Y=1.725
+ $X2=12.155 $Y2=1.725
r251 50 81 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=12.32 $Y=0.425
+ $X2=12.32 $Y2=0.515
r252 47 48 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=13.865
+ $Y=1.485 $X2=13.865 $Y2=1.485
r253 45 47 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=13.435 $Y=1.485
+ $X2=13.865 $Y2=1.485
r254 44 45 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=13.35 $Y=1.32
+ $X2=13.435 $Y2=1.485
r255 43 44 58.3904 $w=1.68e-07 $l=8.95e-07 $layer=LI1_cond $X=13.35 $Y=0.425
+ $X2=13.35 $Y2=1.32
r256 42 50 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=12.485 $Y=0.34
+ $X2=12.32 $Y2=0.425
r257 41 43 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=13.265 $Y=0.34
+ $X2=13.35 $Y2=0.425
r258 41 42 50.8877 $w=1.68e-07 $l=7.8e-07 $layer=LI1_cond $X=13.265 $Y=0.34
+ $X2=12.485 $Y2=0.34
r259 37 53 6.62588 $w=2.9e-07 $l=5.85064e-07 $layer=LI1_cond $X=12.575 $Y=2.12
+ $X2=12.155 $Y2=1.725
r260 37 39 25.8147 $w=2.48e-07 $l=5.6e-07 $layer=LI1_cond $X=12.575 $Y=2.12
+ $X2=12.575 $Y2=2.68
r261 35 73 38.1988 $w=3.47e-07 $l=2.75e-07 $layer=POLY_cond $X=11.725 $Y=1.932
+ $X2=11.45 $Y2=1.932
r262 34 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=11.725
+ $Y=1.89 $X2=11.725 $Y2=1.89
r263 32 53 0.257366 $w=3.95e-07 $l=1.97e-07 $layer=LI1_cond $X=12.155 $Y=1.922
+ $X2=12.155 $Y2=1.725
r264 32 34 12.5456 $w=3.93e-07 $l=4.3e-07 $layer=LI1_cond $X=12.155 $Y=1.922
+ $X2=11.725 $Y2=1.922
r265 31 66 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.04 $Y=0.98
+ $X2=3.04 $Y2=1.145
r266 26 48 38.6072 $w=2.91e-07 $l=1.83916e-07 $layer=POLY_cond $X=13.905 $Y=1.32
+ $X2=13.865 $Y2=1.485
r267 26 28 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=13.905 $Y=1.32
+ $X2=13.905 $Y2=0.76
r268 23 48 57.6553 $w=2.91e-07 $l=2.87402e-07 $layer=POLY_cond $X=13.85 $Y=1.765
+ $X2=13.865 $Y2=1.485
r269 23 25 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=13.85 $Y=1.765
+ $X2=13.85 $Y2=2.4
r270 19 73 22.4223 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=11.45 $Y=1.725
+ $X2=11.45 $Y2=1.932
r271 19 21 474.309 $w=1.5e-07 $l=9.25e-07 $layer=POLY_cond $X=11.45 $Y=1.725
+ $X2=11.45 $Y2=0.8
r272 16 72 22.4223 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=11.435 $Y=2.14
+ $X2=11.435 $Y2=1.932
r273 16 18 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=11.435 $Y=2.14
+ $X2=11.435 $Y2=2.425
r274 13 15 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=3.095 $Y=2.445
+ $X2=3.095 $Y2=2.73
r275 12 13 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=3.095 $Y=2.355
+ $X2=3.095 $Y2=2.445
r276 12 71 141.879 $w=1.8e-07 $l=3.65e-07 $layer=POLY_cond $X=3.095 $Y=2.355
+ $X2=3.095 $Y2=1.99
r277 9 31 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=2.95 $Y=0.58 $X2=2.95
+ $Y2=0.98
r278 2 53 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=12.465
+ $Y=1.825 $X2=12.615 $Y2=1.97
r279 2 39 400 $w=1.7e-07 $l=9.26971e-07 $layer=licon1_PDIFF $count=1 $X=12.465
+ $Y=1.825 $X2=12.615 $Y2=2.68
r280 1 81 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=12.18
+ $Y=0.37 $X2=12.32 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__EDFXBP_1%CLK 1 3 4 6 7
r33 10 11 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.22
+ $Y=1.385 $X2=4.22 $Y2=1.385
r34 7 11 1.60667 $w=6.68e-07 $l=9e-08 $layer=LI1_cond $X=4.05 $Y=1.295 $X2=4.05
+ $Y2=1.385
r35 4 10 63.0862 $w=4.76e-07 $l=4.06571e-07 $layer=POLY_cond $X=4.105 $Y=1.765
+ $X2=4.05 $Y2=1.385
r36 4 6 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=4.105 $Y=1.765
+ $X2=4.105 $Y2=2.4
r37 1 10 41.3152 $w=4.76e-07 $l=1.81659e-07 $layer=POLY_cond $X=4.015 $Y=1.22
+ $X2=4.05 $Y2=1.385
r38 1 3 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=4.015 $Y=1.22 $X2=4.015
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HS__EDFXBP_1%A_1008_74# 1 2 7 9 10 12 13 15 17 19 20 22
+ 25 27 28 29 34 35 38 39 42 43 44 46 48 51 55 56 58 59 62 63 66 68 69 71 72 73
+ 81
c224 66 0 1.31135e-19 $X=6.72 $Y=1.18
c225 62 0 1.41465e-19 $X=6.19 $Y=2.215
c226 56 0 2.75091e-19 $X=11 $Y=1.635
c227 44 0 1.9677e-19 $X=7.81 $Y=0.34
c228 19 0 7.23051e-20 $X=10.955 $Y=2.05
c229 17 0 3.32586e-20 $X=9.395 $Y=1.26
r230 72 81 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=9.92 $Y=1.285
+ $X2=9.755 $Y2=1.285
r231 71 73 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=9.92 $Y=1.285
+ $X2=10.085 $Y2=1.285
r232 71 72 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.92
+ $Y=1.285 $X2=9.92 $Y2=1.285
r233 69 71 19.2074 $w=3.28e-07 $l=5.5e-07 $layer=LI1_cond $X=9.37 $Y=1.285
+ $X2=9.92 $Y2=1.285
r234 68 69 8.63679 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=9.2 $Y=1.207
+ $X2=9.37 $Y2=1.207
r235 66 76 21.8577 $w=3.3e-07 $l=1.25e-07 $layer=POLY_cond $X=6.72 $Y=1.18
+ $X2=6.595 $Y2=1.18
r236 65 66 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.72
+ $Y=1.18 $X2=6.72 $Y2=1.18
r237 63 65 5.9927 $w=2.48e-07 $l=1.3e-07 $layer=LI1_cond $X=6.76 $Y=1.05
+ $X2=6.76 $Y2=1.18
r238 62 75 71.6729 $w=2.69e-07 $l=4e-07 $layer=POLY_cond $X=6.19 $Y=2.257
+ $X2=6.59 $Y2=2.257
r239 61 62 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.19
+ $Y=2.215 $X2=6.19 $Y2=2.215
r240 59 61 8.7403 $w=3.35e-07 $l=2.4e-07 $layer=LI1_cond $X=6.155 $Y=1.975
+ $X2=6.155 $Y2=2.215
r241 56 85 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=11 $Y=1.635 $X2=11
+ $Y2=1.8
r242 55 56 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=11
+ $Y=1.635 $X2=11 $Y2=1.635
r243 53 55 14.7257 $w=2.68e-07 $l=3.45e-07 $layer=LI1_cond $X=10.97 $Y=1.29
+ $X2=10.97 $Y2=1.635
r244 51 53 7.28469 $w=1.7e-07 $l=1.72337e-07 $layer=LI1_cond $X=10.835 $Y=1.205
+ $X2=10.97 $Y2=1.29
r245 51 73 48.9305 $w=1.68e-07 $l=7.5e-07 $layer=LI1_cond $X=10.835 $Y=1.205
+ $X2=10.085 $Y2=1.205
r246 48 68 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=8.49 $Y=1.05
+ $X2=9.2 $Y2=1.05
r247 46 48 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.405 $Y=0.965
+ $X2=8.49 $Y2=1.05
r248 45 46 35.2299 $w=1.68e-07 $l=5.4e-07 $layer=LI1_cond $X=8.405 $Y=0.425
+ $X2=8.405 $Y2=0.965
r249 43 45 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.32 $Y=0.34
+ $X2=8.405 $Y2=0.425
r250 43 44 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=8.32 $Y=0.34
+ $X2=7.81 $Y2=0.34
r251 41 44 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.725 $Y=0.425
+ $X2=7.81 $Y2=0.34
r252 41 42 35.2299 $w=1.68e-07 $l=5.4e-07 $layer=LI1_cond $X=7.725 $Y=0.425
+ $X2=7.725 $Y2=0.965
r253 40 63 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.885 $Y=1.05
+ $X2=6.76 $Y2=1.05
r254 39 42 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.64 $Y=1.05
+ $X2=7.725 $Y2=0.965
r255 39 40 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=7.64 $Y=1.05
+ $X2=6.885 $Y2=1.05
r256 38 63 3.91831 $w=2.48e-07 $l=8.5e-08 $layer=LI1_cond $X=6.76 $Y=0.965
+ $X2=6.76 $Y2=1.05
r257 37 38 24.8928 $w=2.48e-07 $l=5.4e-07 $layer=LI1_cond $X=6.76 $Y=0.425
+ $X2=6.76 $Y2=0.965
r258 36 58 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.125 $Y=0.34
+ $X2=6.04 $Y2=0.34
r259 35 37 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=6.635 $Y=0.34
+ $X2=6.76 $Y2=0.425
r260 35 36 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=6.635 $Y=0.34
+ $X2=6.125 $Y2=0.34
r261 34 59 8.96243 $w=3.35e-07 $l=2.14942e-07 $layer=LI1_cond $X=6.04 $Y=1.81
+ $X2=6.155 $Y2=1.975
r262 33 58 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.04 $Y=0.425
+ $X2=6.04 $Y2=0.34
r263 33 34 90.3583 $w=1.68e-07 $l=1.385e-06 $layer=LI1_cond $X=6.04 $Y=0.425
+ $X2=6.04 $Y2=1.81
r264 29 59 0.808037 $w=3.3e-07 $l=2e-07 $layer=LI1_cond $X=5.955 $Y=1.975
+ $X2=6.155 $Y2=1.975
r265 29 31 8.20679 $w=3.28e-07 $l=2.35e-07 $layer=LI1_cond $X=5.955 $Y=1.975
+ $X2=5.72 $Y2=1.975
r266 27 58 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.955 $Y=0.34
+ $X2=6.04 $Y2=0.34
r267 27 28 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=5.955 $Y=0.34
+ $X2=5.345 $Y2=0.34
r268 23 28 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=5.22 $Y=0.425
+ $X2=5.345 $Y2=0.34
r269 23 25 4.14879 $w=2.48e-07 $l=9e-08 $layer=LI1_cond $X=5.22 $Y=0.425
+ $X2=5.22 $Y2=0.515
r270 20 22 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=10.955 $Y=2.14
+ $X2=10.955 $Y2=2.425
r271 19 20 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=10.955 $Y=2.05
+ $X2=10.955 $Y2=2.14
r272 19 85 97.1774 $w=1.8e-07 $l=2.5e-07 $layer=POLY_cond $X=10.955 $Y=2.05
+ $X2=10.955 $Y2=1.8
r273 17 81 184.596 $w=1.5e-07 $l=3.6e-07 $layer=POLY_cond $X=9.395 $Y=1.26
+ $X2=9.755 $Y2=1.26
r274 13 17 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=9.32 $Y=1.185
+ $X2=9.395 $Y2=1.26
r275 13 15 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=9.32 $Y=1.185
+ $X2=9.32 $Y2=0.74
r276 10 76 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.595 $Y=1.015
+ $X2=6.595 $Y2=1.18
r277 10 12 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=6.595 $Y=1.015
+ $X2=6.595 $Y2=0.695
r278 7 75 16.4183 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=6.59 $Y=2.465
+ $X2=6.59 $Y2=2.257
r279 7 9 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=6.59 $Y=2.465 $X2=6.59
+ $Y2=2.75
r280 2 31 600 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=5.57
+ $Y=1.83 $X2=5.72 $Y2=1.975
r281 1 25 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=5.04
+ $Y=0.37 $X2=5.18 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__EDFXBP_1%A_818_74# 1 2 9 11 13 15 16 20 22 25 26 28
+ 29 31 33 34 35 36 38 39 40 44 46 51 53 54 55 56 59 60 61 64 68 75 77 82 87
c220 82 0 3.39525e-20 $X=10.46 $Y=1.625
c221 77 0 1.51669e-19 $X=8.28 $Y=2.63
c222 75 0 1.41465e-19 $X=7.235 $Y=2.23
c223 34 0 1.59075e-19 $X=10.985 $Y=1.185
c224 22 0 1.37651e-20 $X=6.595 $Y=1.68
r225 87 88 33.431 $w=4.05e-07 $l=7.5e-08 $layer=POLY_cond $X=4.837 $Y=1.68
+ $X2=4.837 $Y2=1.605
r226 82 85 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=10.46 $Y=1.625
+ $X2=10.46 $Y2=1.705
r227 82 83 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.46
+ $Y=1.625 $X2=10.46 $Y2=1.625
r228 77 79 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=8.28 $Y=2.63
+ $X2=8.28 $Y2=2.84
r229 72 75 6.91466 $w=2.98e-07 $l=1.8e-07 $layer=LI1_cond $X=7.055 $Y=2.23
+ $X2=7.235 $Y2=2.23
r230 72 73 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.055
+ $Y=2.215 $X2=7.055 $Y2=2.215
r231 69 87 40.51 $w=4.05e-07 $l=2.95e-07 $layer=POLY_cond $X=4.837 $Y=1.975
+ $X2=4.837 $Y2=1.68
r232 68 69 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.8
+ $Y=1.975 $X2=4.8 $Y2=1.975
r233 66 68 5.5876 $w=3.28e-07 $l=1.6e-07 $layer=LI1_cond $X=4.64 $Y=1.975
+ $X2=4.8 $Y2=1.975
r234 60 85 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.295 $Y=1.705
+ $X2=10.46 $Y2=1.705
r235 60 61 58.0642 $w=1.68e-07 $l=8.9e-07 $layer=LI1_cond $X=10.295 $Y=1.705
+ $X2=9.405 $Y2=1.705
r236 58 61 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.32 $Y=1.79
+ $X2=9.405 $Y2=1.705
r237 58 59 62.9572 $w=1.68e-07 $l=9.65e-07 $layer=LI1_cond $X=9.32 $Y=1.79
+ $X2=9.32 $Y2=2.755
r238 57 79 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.365 $Y=2.84
+ $X2=8.28 $Y2=2.84
r239 56 59 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.235 $Y=2.84
+ $X2=9.32 $Y2=2.755
r240 56 57 56.7594 $w=1.68e-07 $l=8.7e-07 $layer=LI1_cond $X=9.235 $Y=2.84
+ $X2=8.365 $Y2=2.84
r241 54 77 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.195 $Y=2.63
+ $X2=8.28 $Y2=2.63
r242 54 55 57.0856 $w=1.68e-07 $l=8.75e-07 $layer=LI1_cond $X=8.195 $Y=2.63
+ $X2=7.32 $Y2=2.63
r243 53 55 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.235 $Y=2.545
+ $X2=7.32 $Y2=2.63
r244 52 75 4.061 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=7.235 $Y=2.38
+ $X2=7.235 $Y2=2.23
r245 52 53 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=7.235 $Y=2.38
+ $X2=7.235 $Y2=2.545
r246 51 66 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.64 $Y=1.81
+ $X2=4.64 $Y2=1.975
r247 50 64 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.64 $Y=1.01
+ $X2=4.64 $Y2=0.925
r248 50 51 52.1925 $w=1.68e-07 $l=8e-07 $layer=LI1_cond $X=4.64 $Y=1.01 $X2=4.64
+ $Y2=1.81
r249 46 66 2.96841 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=4.555 $Y=1.975
+ $X2=4.64 $Y2=1.975
r250 46 48 7.85757 $w=3.28e-07 $l=2.25e-07 $layer=LI1_cond $X=4.555 $Y=1.975
+ $X2=4.33 $Y2=1.975
r251 42 64 26.7487 $w=1.68e-07 $l=4.1e-07 $layer=LI1_cond $X=4.23 $Y=0.925
+ $X2=4.64 $Y2=0.925
r252 42 44 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=4.23 $Y=0.84
+ $X2=4.23 $Y2=0.515
r253 36 38 99.6133 $w=1.5e-07 $l=3.1e-07 $layer=POLY_cond $X=11.06 $Y=1.11
+ $X2=11.06 $Y2=0.8
r254 34 36 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=10.985 $Y=1.185
+ $X2=11.06 $Y2=1.11
r255 34 35 184.596 $w=1.5e-07 $l=3.6e-07 $layer=POLY_cond $X=10.985 $Y=1.185
+ $X2=10.625 $Y2=1.185
r256 33 83 38.5718 $w=2.96e-07 $l=2.05122e-07 $layer=POLY_cond $X=10.55 $Y=1.46
+ $X2=10.46 $Y2=1.625
r257 32 35 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=10.55 $Y=1.26
+ $X2=10.625 $Y2=1.185
r258 32 33 102.553 $w=1.5e-07 $l=2e-07 $layer=POLY_cond $X=10.55 $Y=1.26
+ $X2=10.55 $Y2=1.46
r259 29 83 54.0414 $w=2.96e-07 $l=2.95127e-07 $layer=POLY_cond $X=10.385
+ $Y=1.885 $X2=10.46 $Y2=1.625
r260 29 31 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=10.385 $Y=1.885
+ $X2=10.385 $Y2=2.46
r261 26 73 53.429 $w=2.79e-07 $l=2.57391e-07 $layer=POLY_cond $X=7.04 $Y=2.465
+ $X2=7.055 $Y2=2.215
r262 26 28 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=7.04 $Y=2.465
+ $X2=7.04 $Y2=2.75
r263 25 73 1.29086 $w=3.3e-07 $l=8.75758e-08 $layer=POLY_cond $X=7.055 $Y=2.215
+ $X2=7.055 $Y2=2.215
r264 24 25 34.9723 $w=3.3e-07 $l=2e-07 $layer=POLY_cond $X=7.055 $Y=2.015
+ $X2=7.055 $Y2=2.215
r265 23 40 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.99 $Y=1.68
+ $X2=5.915 $Y2=1.68
r266 22 24 108.771 $w=2.12e-07 $l=5.44702e-07 $layer=POLY_cond $X=6.595 $Y=1.68
+ $X2=7.055 $Y2=1.865
r267 22 23 310.223 $w=1.5e-07 $l=6.05e-07 $layer=POLY_cond $X=6.595 $Y=1.68
+ $X2=5.99 $Y2=1.68
r268 18 40 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.915 $Y=1.605
+ $X2=5.915 $Y2=1.68
r269 18 20 466.617 $w=1.5e-07 $l=9.1e-07 $layer=POLY_cond $X=5.915 $Y=1.605
+ $X2=5.915 $Y2=0.695
r270 17 39 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.57 $Y=1.68
+ $X2=5.495 $Y2=1.68
r271 16 40 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.84 $Y=1.68
+ $X2=5.915 $Y2=1.68
r272 16 17 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=5.84 $Y=1.68
+ $X2=5.57 $Y2=1.68
r273 13 39 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.495 $Y=1.755
+ $X2=5.495 $Y2=1.68
r274 13 15 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=5.495 $Y=1.755
+ $X2=5.495 $Y2=2.39
r275 12 87 26.1659 $w=1.5e-07 $l=2.03e-07 $layer=POLY_cond $X=5.04 $Y=1.68
+ $X2=4.837 $Y2=1.68
r276 11 39 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.42 $Y=1.68
+ $X2=5.495 $Y2=1.68
r277 11 12 194.851 $w=1.5e-07 $l=3.8e-07 $layer=POLY_cond $X=5.42 $Y=1.68
+ $X2=5.04 $Y2=1.68
r278 9 88 443.543 $w=1.5e-07 $l=8.65e-07 $layer=POLY_cond $X=4.965 $Y=0.74
+ $X2=4.965 $Y2=1.605
r279 2 48 600 $w=1.7e-07 $l=2.43721e-07 $layer=licon1_PDIFF $count=1 $X=4.18
+ $Y=1.84 $X2=4.33 $Y2=2.02
r280 1 44 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=4.09
+ $Y=0.37 $X2=4.23 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__EDFXBP_1%A_1419_71# 1 2 9 12 13 15 18 20 22 24 25 29
+ 31 33 38 40 41 44 46 47 50
c137 50 0 1.51669e-19 $X=8.865 $Y=2.42
c138 46 0 1.30788e-19 $X=7.535 $Y=1.437
c139 31 0 3.32586e-20 $X=8.7 $Y=1.39
c140 20 0 3.39525e-20 $X=9.89 $Y=1.81
c141 9 0 1.9677e-19 $X=7.17 $Y=0.695
r142 51 59 12.9189 $w=3.35e-07 $l=7.5e-08 $layer=POLY_cond $X=8.867 $Y=1.885
+ $X2=8.867 $Y2=1.81
r143 50 51 92.1545 $w=3.35e-07 $l=5.35e-07 $layer=POLY_cond $X=8.867 $Y=2.42
+ $X2=8.867 $Y2=1.885
r144 49 50 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=8.865
+ $Y=2.42 $X2=8.865 $Y2=2.42
r145 43 46 8.65224 $w=2.63e-07 $l=1.65e-07 $layer=LI1_cond $X=7.37 $Y=1.437
+ $X2=7.535 $Y2=1.437
r146 43 44 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.37
+ $Y=1.435 $X2=7.37 $Y2=1.435
r147 41 59 12.0576 $w=3.35e-07 $l=7e-08 $layer=POLY_cond $X=8.867 $Y=1.74
+ $X2=8.867 $Y2=1.81
r148 41 58 46.255 $w=3.35e-07 $l=1.65e-07 $layer=POLY_cond $X=8.867 $Y=1.74
+ $X2=8.867 $Y2=1.575
r149 40 41 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=8.865
+ $Y=1.74 $X2=8.865 $Y2=1.74
r150 38 49 3.2138 $w=3.3e-07 $l=2.3e-07 $layer=LI1_cond $X=8.865 $Y=2.125
+ $X2=8.865 $Y2=2.355
r151 38 40 13.4452 $w=3.28e-07 $l=3.85e-07 $layer=LI1_cond $X=8.865 $Y=2.125
+ $X2=8.865 $Y2=1.74
r152 37 40 9.25447 $w=3.28e-07 $l=2.65e-07 $layer=LI1_cond $X=8.865 $Y=1.475
+ $X2=8.865 $Y2=1.74
r153 33 49 3.77273 $w=2.5e-07 $l=2.11069e-07 $layer=LI1_cond $X=8.7 $Y=2.25
+ $X2=8.865 $Y2=2.355
r154 33 35 14.0598 $w=2.48e-07 $l=3.05e-07 $layer=LI1_cond $X=8.7 $Y=2.25
+ $X2=8.395 $Y2=2.25
r155 32 47 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.15 $Y=1.39
+ $X2=8.065 $Y2=1.39
r156 31 37 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=8.7 $Y=1.39
+ $X2=8.865 $Y2=1.475
r157 31 32 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=8.7 $Y=1.39
+ $X2=8.15 $Y2=1.39
r158 27 47 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.065 $Y=1.305
+ $X2=8.065 $Y2=1.39
r159 27 29 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=8.065 $Y=1.305
+ $X2=8.065 $Y2=0.81
r160 25 47 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.98 $Y=1.39
+ $X2=8.065 $Y2=1.39
r161 25 46 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=7.98 $Y=1.39
+ $X2=7.535 $Y2=1.39
r162 22 24 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=9.965 $Y=1.885
+ $X2=9.965 $Y2=2.46
r163 21 59 21.5811 $w=1.5e-07 $l=1.68e-07 $layer=POLY_cond $X=9.035 $Y=1.81
+ $X2=8.867 $Y2=1.81
r164 20 22 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=9.89 $Y=1.81
+ $X2=9.965 $Y2=1.885
r165 20 21 438.415 $w=1.5e-07 $l=8.55e-07 $layer=POLY_cond $X=9.89 $Y=1.81
+ $X2=9.035 $Y2=1.81
r166 18 58 428.16 $w=1.5e-07 $l=8.35e-07 $layer=POLY_cond $X=8.96 $Y=0.74
+ $X2=8.96 $Y2=1.575
r167 13 15 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=7.55 $Y=2.465
+ $X2=7.55 $Y2=2.75
r168 12 13 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=7.55 $Y=2.375
+ $X2=7.55 $Y2=2.465
r169 11 44 30.0208 $w=2.89e-07 $l=2.80936e-07 $layer=POLY_cond $X=7.55 $Y=1.625
+ $X2=7.37 $Y2=1.42
r170 11 12 291.532 $w=1.8e-07 $l=7.5e-07 $layer=POLY_cond $X=7.55 $Y=1.625
+ $X2=7.55 $Y2=2.375
r171 7 44 33.3564 $w=2.89e-07 $l=2.88141e-07 $layer=POLY_cond $X=7.17 $Y=1.215
+ $X2=7.37 $Y2=1.42
r172 7 9 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=7.17 $Y=1.215
+ $X2=7.17 $Y2=0.695
r173 2 35 600 $w=1.7e-07 $l=2.33238e-07 $layer=licon1_PDIFF $count=1 $X=8.245
+ $Y=2.12 $X2=8.395 $Y2=2.29
r174 1 29 182 $w=1.7e-07 $l=5.05173e-07 $layer=licon1_NDIFF $count=1 $X=7.925
+ $Y=0.37 $X2=8.065 $Y2=0.81
.ends

.subckt PM_SKY130_FD_SC_HS__EDFXBP_1%A_1198_97# 1 2 7 9 11 12 14 17 21 24 26 33
+ 35
r102 33 35 8.46729 $w=3.08e-07 $l=1.65e-07 $layer=LI1_cond $X=8.095 $Y=1.8
+ $X2=7.93 $Y2=1.8
r103 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.095
+ $Y=1.79 $X2=8.095 $Y2=1.79
r104 27 28 11.9654 $w=2.6e-07 $l=2.55e-07 $layer=LI1_cond $X=6.38 $Y=1.685
+ $X2=6.635 $Y2=1.685
r105 26 28 5.4494 $w=2.6e-07 $l=1.77482e-07 $layer=LI1_cond $X=6.72 $Y=1.825
+ $X2=6.635 $Y2=1.685
r106 26 35 78.9412 $w=1.68e-07 $l=1.21e-06 $layer=LI1_cond $X=6.72 $Y=1.825
+ $X2=7.93 $Y2=1.825
r107 24 31 5.95122 $w=3.69e-07 $l=2.91419e-07 $layer=LI1_cond $X=6.635 $Y=2.55
+ $X2=6.815 $Y2=2.765
r108 23 28 3.22376 $w=1.7e-07 $l=2.25e-07 $layer=LI1_cond $X=6.635 $Y=1.91
+ $X2=6.635 $Y2=1.685
r109 23 24 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=6.635 $Y=1.91
+ $X2=6.635 $Y2=2.55
r110 19 27 3.22376 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=6.38 $Y=1.515
+ $X2=6.38 $Y2=1.685
r111 19 21 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=6.38 $Y=1.515
+ $X2=6.38 $Y2=0.76
r112 15 17 79.4787 $w=1.5e-07 $l=1.55e-07 $layer=POLY_cond $X=7.85 $Y=1.16
+ $X2=8.005 $Y2=1.16
r113 12 34 53.1722 $w=2.97e-07 $l=2.90086e-07 $layer=POLY_cond $X=8.17 $Y=2.045
+ $X2=8.095 $Y2=1.79
r114 12 14 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=8.17 $Y=2.045
+ $X2=8.17 $Y2=2.54
r115 11 34 38.5662 $w=2.97e-07 $l=2.05122e-07 $layer=POLY_cond $X=8.005 $Y=1.625
+ $X2=8.095 $Y2=1.79
r116 10 17 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=8.005 $Y=1.235
+ $X2=8.005 $Y2=1.16
r117 10 11 199.979 $w=1.5e-07 $l=3.9e-07 $layer=POLY_cond $X=8.005 $Y=1.235
+ $X2=8.005 $Y2=1.625
r118 7 15 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.85 $Y=1.085
+ $X2=7.85 $Y2=1.16
r119 7 9 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=7.85 $Y=1.085
+ $X2=7.85 $Y2=0.69
r120 2 31 600 $w=1.7e-07 $l=2.90474e-07 $layer=licon1_PDIFF $count=1 $X=6.665
+ $Y=2.54 $X2=6.815 $Y2=2.765
r121 1 21 182 $w=1.7e-07 $l=5.09264e-07 $layer=licon1_NDIFF $count=1 $X=5.99
+ $Y=0.485 $X2=6.38 $Y2=0.76
.ends

.subckt PM_SKY130_FD_SC_HS__EDFXBP_1%A_1879_74# 1 2 9 11 13 14 15 16 18 20 21 23
+ 25 27 33 35 37 40 42 45 50
c129 50 0 1.03676e-19 $X=11.36 $Y=1.32
c130 27 0 1.71415e-19 $X=11.275 $Y=0.785
r131 52 53 31.2916 $w=4.39e-07 $l=2.85e-07 $layer=POLY_cond $X=12.105 $Y=1.452
+ $X2=12.39 $Y2=1.452
r132 46 52 22.508 $w=4.39e-07 $l=2.05e-07 $layer=POLY_cond $X=11.9 $Y=1.452
+ $X2=12.105 $Y2=1.452
r133 45 46 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=11.9
+ $Y=1.32 $X2=11.9 $Y2=1.32
r134 43 50 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=11.445 $Y=1.32
+ $X2=11.36 $Y2=1.32
r135 43 45 15.8897 $w=3.28e-07 $l=4.55e-07 $layer=LI1_cond $X=11.445 $Y=1.32
+ $X2=11.9 $Y2=1.32
r136 41 50 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.36 $Y=1.485
+ $X2=11.36 $Y2=1.32
r137 41 42 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=11.36 $Y=1.485
+ $X2=11.36 $Y2=1.985
r138 40 50 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.36 $Y=1.155
+ $X2=11.36 $Y2=1.32
r139 39 40 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=11.36 $Y=0.95
+ $X2=11.36 $Y2=1.155
r140 38 49 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.775 $Y=2.07
+ $X2=10.61 $Y2=2.07
r141 37 42 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=11.275 $Y=2.07
+ $X2=11.36 $Y2=1.985
r142 37 38 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=11.275 $Y=2.07
+ $X2=10.775 $Y2=2.07
r143 33 49 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=10.61 $Y=2.155
+ $X2=10.61 $Y2=2.07
r144 33 35 23.0489 $w=3.28e-07 $l=6.6e-07 $layer=LI1_cond $X=10.61 $Y=2.155
+ $X2=10.61 $Y2=2.815
r145 29 32 42.6055 $w=3.28e-07 $l=1.22e-06 $layer=LI1_cond $X=9.625 $Y=0.785
+ $X2=10.845 $Y2=0.785
r146 27 39 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=11.275 $Y=0.785
+ $X2=11.36 $Y2=0.95
r147 27 32 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=11.275 $Y=0.785
+ $X2=10.845 $Y2=0.785
r148 24 25 47.4664 $w=3.1e-07 $l=2.55e-07 $layer=POLY_cond $X=13.145 $Y=1.36
+ $X2=13.4 $Y2=1.36
r149 21 23 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=13.4 $Y=1.765
+ $X2=13.4 $Y2=2.4
r150 20 21 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=13.4 $Y=1.675
+ $X2=13.4 $Y2=1.765
r151 19 25 15.4789 $w=1.8e-07 $l=1.55e-07 $layer=POLY_cond $X=13.4 $Y=1.515
+ $X2=13.4 $Y2=1.36
r152 19 20 62.1936 $w=1.8e-07 $l=1.6e-07 $layer=POLY_cond $X=13.4 $Y=1.515
+ $X2=13.4 $Y2=1.675
r153 16 24 19.7411 $w=1.5e-07 $l=1.55e-07 $layer=POLY_cond $X=13.145 $Y=1.205
+ $X2=13.145 $Y2=1.36
r154 16 18 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=13.145 $Y=1.205
+ $X2=13.145 $Y2=0.76
r155 15 53 14.1054 $w=4.39e-07 $l=1.29399e-07 $layer=POLY_cond $X=12.48 $Y=1.36
+ $X2=12.39 $Y2=1.452
r156 14 24 13.9607 $w=3.1e-07 $l=7.5e-08 $layer=POLY_cond $X=13.07 $Y=1.36
+ $X2=13.145 $Y2=1.36
r157 14 15 109.824 $w=3.1e-07 $l=5.9e-07 $layer=POLY_cond $X=13.07 $Y=1.36
+ $X2=12.48 $Y2=1.36
r158 11 53 28.1521 $w=1.5e-07 $l=2.98e-07 $layer=POLY_cond $X=12.39 $Y=1.75
+ $X2=12.39 $Y2=1.452
r159 11 13 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=12.39 $Y=1.75
+ $X2=12.39 $Y2=2.325
r160 7 52 28.1521 $w=1.5e-07 $l=2.97e-07 $layer=POLY_cond $X=12.105 $Y=1.155
+ $X2=12.105 $Y2=1.452
r161 7 9 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=12.105 $Y=1.155
+ $X2=12.105 $Y2=0.69
r162 2 49 300 $w=1.7e-07 $l=2.2798e-07 $layer=licon1_PDIFF $count=2 $X=10.46
+ $Y=1.96 $X2=10.61 $Y2=2.125
r163 2 35 600 $w=1.7e-07 $l=9.26971e-07 $layer=licon1_PDIFF $count=1 $X=10.46
+ $Y=1.96 $X2=10.61 $Y2=2.815
r164 1 32 91 $w=1.7e-07 $l=1.64446e-06 $layer=licon1_NDIFF $count=2 $X=9.395
+ $Y=0.37 $X2=10.845 $Y2=0.785
r165 1 29 91 $w=1.7e-07 $l=5.17373e-07 $layer=licon1_NDIFF $count=2 $X=9.395
+ $Y=0.37 $X2=9.625 $Y2=0.785
.ends

.subckt PM_SKY130_FD_SC_HS__EDFXBP_1%A_27_74# 1 2 3 4 5 6 20 23 25 28 29 30 32
+ 33 34 37 40 41 44 45 47 49 52 53 55 60 62 66 68 73
c178 68 0 2.34044e-19 $X=3.35 $Y=2.385
c179 34 0 1.30607e-19 $X=2.225 $Y=2.375
c180 28 0 1.24694e-19 $X=1.46 $Y=2.905
c181 23 0 2.12276e-20 $X=0.28 $Y=2.75
r182 64 66 7.6705 $w=4.58e-07 $l=2.95e-07 $layer=LI1_cond $X=3.165 $Y=0.58
+ $X2=3.46 $Y2=0.58
r183 57 60 9.25447 $w=3.28e-07 $l=2.65e-07 $layer=LI1_cond $X=0.17 $Y=0.585
+ $X2=0.435 $Y2=0.585
r184 53 55 32.9465 $w=1.68e-07 $l=5.05e-07 $layer=LI1_cond $X=5.775 $Y=2.975
+ $X2=6.28 $Y2=2.975
r185 52 53 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.69 $Y=2.89
+ $X2=5.775 $Y2=2.975
r186 51 52 26.7487 $w=1.68e-07 $l=4.1e-07 $layer=LI1_cond $X=5.69 $Y=2.48
+ $X2=5.69 $Y2=2.89
r187 47 69 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=5.66 $Y=1.385
+ $X2=5.3 $Y2=1.385
r188 47 49 24.8928 $w=2.48e-07 $l=5.4e-07 $layer=LI1_cond $X=5.66 $Y=1.3
+ $X2=5.66 $Y2=0.76
r189 46 73 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.385 $Y=2.395
+ $X2=5.3 $Y2=2.395
r190 45 51 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.605 $Y=2.395
+ $X2=5.69 $Y2=2.48
r191 45 46 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=5.605 $Y=2.395
+ $X2=5.385 $Y2=2.395
r192 44 73 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.3 $Y=2.31 $X2=5.3
+ $Y2=2.395
r193 43 69 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.3 $Y=1.47 $X2=5.3
+ $Y2=1.385
r194 43 44 54.8021 $w=1.68e-07 $l=8.4e-07 $layer=LI1_cond $X=5.3 $Y=1.47 $X2=5.3
+ $Y2=2.31
r195 42 68 4.69131 $w=1.7e-07 $l=1.99937e-07 $layer=LI1_cond $X=3.545 $Y=2.395
+ $X2=3.35 $Y2=2.385
r196 41 73 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.215 $Y=2.395
+ $X2=5.3 $Y2=2.395
r197 41 42 108.952 $w=1.68e-07 $l=1.67e-06 $layer=LI1_cond $X=5.215 $Y=2.395
+ $X2=3.545 $Y2=2.395
r198 40 68 1.68048 $w=1.7e-07 $l=1.50167e-07 $layer=LI1_cond $X=3.46 $Y=2.29
+ $X2=3.35 $Y2=2.385
r199 39 66 6.6364 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=3.46 $Y=0.81 $X2=3.46
+ $Y2=0.58
r200 39 40 96.5562 $w=1.68e-07 $l=1.48e-06 $layer=LI1_cond $X=3.46 $Y=0.81
+ $X2=3.46 $Y2=2.29
r201 35 68 1.68048 $w=3.9e-07 $l=9.5e-08 $layer=LI1_cond $X=3.35 $Y=2.48
+ $X2=3.35 $Y2=2.385
r202 35 37 7.38745 $w=3.88e-07 $l=2.5e-07 $layer=LI1_cond $X=3.35 $Y=2.48
+ $X2=3.35 $Y2=2.73
r203 33 68 4.69131 $w=1.7e-07 $l=1.99937e-07 $layer=LI1_cond $X=3.155 $Y=2.375
+ $X2=3.35 $Y2=2.385
r204 33 34 60.6738 $w=1.68e-07 $l=9.3e-07 $layer=LI1_cond $X=3.155 $Y=2.375
+ $X2=2.225 $Y2=2.375
r205 31 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.14 $Y=2.46
+ $X2=2.225 $Y2=2.375
r206 31 32 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=2.14 $Y=2.46
+ $X2=2.14 $Y2=2.905
r207 29 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.055 $Y=2.99
+ $X2=2.14 $Y2=2.905
r208 29 30 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=2.055 $Y=2.99
+ $X2=1.545 $Y2=2.99
r209 28 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.46 $Y=2.905
+ $X2=1.545 $Y2=2.99
r210 27 28 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=1.46 $Y=2.46
+ $X2=1.46 $Y2=2.905
r211 26 62 2.98021 $w=1.7e-07 $l=1.8e-07 $layer=LI1_cond $X=0.445 $Y=2.375
+ $X2=0.265 $Y2=2.375
r212 25 27 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.375 $Y=2.375
+ $X2=1.46 $Y2=2.46
r213 25 26 60.6738 $w=1.68e-07 $l=9.3e-07 $layer=LI1_cond $X=1.375 $Y=2.375
+ $X2=0.445 $Y2=2.375
r214 21 62 3.52026 $w=2.65e-07 $l=8.5e-08 $layer=LI1_cond $X=0.265 $Y=2.46
+ $X2=0.265 $Y2=2.375
r215 21 23 9.28357 $w=3.58e-07 $l=2.9e-07 $layer=LI1_cond $X=0.265 $Y=2.46
+ $X2=0.265 $Y2=2.75
r216 20 62 3.52026 $w=2.65e-07 $l=1.30767e-07 $layer=LI1_cond $X=0.17 $Y=2.29
+ $X2=0.265 $Y2=2.375
r217 19 57 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.17 $Y=0.75
+ $X2=0.17 $Y2=0.585
r218 19 20 100.471 $w=1.68e-07 $l=1.54e-06 $layer=LI1_cond $X=0.17 $Y=0.75
+ $X2=0.17 $Y2=2.29
r219 6 55 600 $w=1.7e-07 $l=5.02295e-07 $layer=licon1_PDIFF $count=1 $X=6.135
+ $Y=2.54 $X2=6.28 $Y2=2.975
r220 5 37 600 $w=1.7e-07 $l=2.74955e-07 $layer=licon1_PDIFF $count=1 $X=3.17
+ $Y=2.52 $X2=3.32 $Y2=2.73
r221 4 23 600 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.54 $X2=0.28 $Y2=2.75
r222 3 49 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=5.575
+ $Y=0.485 $X2=5.7 $Y2=0.76
r223 2 64 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=3.025
+ $Y=0.37 $X2=3.165 $Y2=0.58
r224 1 60 182 $w=1.7e-07 $l=3.93065e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.37 $X2=0.435 $Y2=0.585
.ends

.subckt PM_SKY130_FD_SC_HS__EDFXBP_1%VPWR 1 2 3 4 5 6 7 8 27 31 35 39 43 47 53
+ 57 62 63 65 66 67 69 74 89 96 104 109 116 117 120 123 126 129 132 137
r160 137 138 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.68 $Y=3.33
+ $X2=13.68 $Y2=3.33
r161 133 135 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.24 $Y=3.33
+ $X2=11.76 $Y2=3.33
r162 132 135 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.76 $Y=3.33
+ $X2=11.76 $Y2=3.33
r163 132 133 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=12.24 $Y=3.33
+ $X2=12.24 $Y2=3.33
r164 129 130 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.84 $Y=3.33
+ $X2=9.84 $Y2=3.33
r165 126 127 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r166 123 124 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r167 120 121 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r168 117 138 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=14.16 $Y=3.33
+ $X2=13.68 $Y2=3.33
r169 116 117 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=14.16 $Y=3.33
+ $X2=14.16 $Y2=3.33
r170 114 137 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=13.79 $Y=3.33
+ $X2=13.665 $Y2=3.33
r171 114 116 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=13.79 $Y=3.33
+ $X2=14.16 $Y2=3.33
r172 113 138 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=13.2 $Y=3.33
+ $X2=13.68 $Y2=3.33
r173 113 133 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=13.2 $Y=3.33
+ $X2=12.24 $Y2=3.33
r174 112 113 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=13.2 $Y=3.33
+ $X2=13.2 $Y2=3.33
r175 110 132 14.4958 $w=1.7e-07 $l=3.93e-07 $layer=LI1_cond $X=12.28 $Y=3.33
+ $X2=11.887 $Y2=3.33
r176 110 112 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=12.28 $Y=3.33
+ $X2=13.2 $Y2=3.33
r177 109 137 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=13.54 $Y=3.33
+ $X2=13.665 $Y2=3.33
r178 109 112 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=13.54 $Y=3.33
+ $X2=13.2 $Y2=3.33
r179 108 135 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.28 $Y=3.33
+ $X2=11.76 $Y2=3.33
r180 108 130 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=11.28 $Y=3.33
+ $X2=9.84 $Y2=3.33
r181 107 108 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=11.28 $Y=3.33
+ $X2=11.28 $Y2=3.33
r182 105 129 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.905 $Y=3.33
+ $X2=9.74 $Y2=3.33
r183 105 107 89.7059 $w=1.68e-07 $l=1.375e-06 $layer=LI1_cond $X=9.905 $Y=3.33
+ $X2=11.28 $Y2=3.33
r184 104 132 14.4958 $w=1.7e-07 $l=3.92e-07 $layer=LI1_cond $X=11.495 $Y=3.33
+ $X2=11.887 $Y2=3.33
r185 104 107 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=11.495 $Y=3.33
+ $X2=11.28 $Y2=3.33
r186 103 130 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.36 $Y=3.33
+ $X2=9.84 $Y2=3.33
r187 102 103 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=9.36 $Y=3.33
+ $X2=9.36 $Y2=3.33
r188 100 103 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=8.4 $Y=3.33
+ $X2=9.36 $Y2=3.33
r189 100 127 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=3.33
+ $X2=7.92 $Y2=3.33
r190 99 102 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=8.4 $Y=3.33
+ $X2=9.36 $Y2=3.33
r191 99 100 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=8.4 $Y=3.33
+ $X2=8.4 $Y2=3.33
r192 97 126 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.025 $Y=3.33
+ $X2=7.86 $Y2=3.33
r193 97 99 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=8.025 $Y=3.33
+ $X2=8.4 $Y2=3.33
r194 96 129 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.575 $Y=3.33
+ $X2=9.74 $Y2=3.33
r195 96 102 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=9.575 $Y=3.33
+ $X2=9.36 $Y2=3.33
r196 95 127 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=7.92 $Y2=3.33
r197 94 95 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r198 91 94 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=5.52 $Y=3.33
+ $X2=7.44 $Y2=3.33
r199 91 92 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r200 89 126 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.695 $Y=3.33
+ $X2=7.86 $Y2=3.33
r201 89 94 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=7.695 $Y=3.33
+ $X2=7.44 $Y2=3.33
r202 88 92 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=5.52 $Y2=3.33
r203 87 88 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r204 85 88 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=5.04 $Y2=3.33
r205 84 87 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=4.08 $Y=3.33
+ $X2=5.04 $Y2=3.33
r206 84 85 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r207 82 85 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.08 $Y2=3.33
r208 82 124 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=2.64 $Y2=3.33
r209 81 82 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r210 79 123 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.645 $Y=3.33
+ $X2=2.52 $Y2=3.33
r211 79 81 62.3048 $w=1.68e-07 $l=9.55e-07 $layer=LI1_cond $X=2.645 $Y=3.33
+ $X2=3.6 $Y2=3.33
r212 78 124 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r213 78 121 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.2 $Y2=3.33
r214 77 78 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r215 75 120 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.205 $Y=3.33
+ $X2=1.08 $Y2=3.33
r216 75 77 62.3048 $w=1.68e-07 $l=9.55e-07 $layer=LI1_cond $X=1.205 $Y=3.33
+ $X2=2.16 $Y2=3.33
r217 74 123 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.395 $Y=3.33
+ $X2=2.52 $Y2=3.33
r218 74 77 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=2.395 $Y=3.33
+ $X2=2.16 $Y2=3.33
r219 72 121 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r220 71 72 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r221 69 120 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.955 $Y=3.33
+ $X2=1.08 $Y2=3.33
r222 69 71 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=0.955 $Y=3.33
+ $X2=0.72 $Y2=3.33
r223 67 95 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=7.2 $Y=3.33
+ $X2=7.44 $Y2=3.33
r224 67 92 0.468274 $w=4.9e-07 $l=1.68e-06 $layer=MET1_cond $X=7.2 $Y=3.33
+ $X2=5.52 $Y2=3.33
r225 65 87 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=5.105 $Y=3.33
+ $X2=5.04 $Y2=3.33
r226 65 66 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.105 $Y=3.33
+ $X2=5.27 $Y2=3.33
r227 64 91 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=5.435 $Y=3.33
+ $X2=5.52 $Y2=3.33
r228 64 66 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.435 $Y=3.33
+ $X2=5.27 $Y2=3.33
r229 62 81 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=3.715 $Y=3.33
+ $X2=3.6 $Y2=3.33
r230 62 63 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.715 $Y=3.33
+ $X2=3.88 $Y2=3.33
r231 61 84 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=4.045 $Y=3.33
+ $X2=4.08 $Y2=3.33
r232 61 63 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.045 $Y=3.33
+ $X2=3.88 $Y2=3.33
r233 57 60 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=13.665 $Y=1.985
+ $X2=13.665 $Y2=2.815
r234 55 137 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=13.665 $Y=3.245
+ $X2=13.665 $Y2=3.33
r235 55 60 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=13.665 $Y=3.245
+ $X2=13.665 $Y2=2.815
r236 51 132 3.09511 $w=7.85e-07 $l=8.5e-08 $layer=LI1_cond $X=11.887 $Y=3.245
+ $X2=11.887 $Y2=3.33
r237 51 53 11.5037 $w=7.83e-07 $l=7.55e-07 $layer=LI1_cond $X=11.887 $Y=3.245
+ $X2=11.887 $Y2=2.49
r238 47 50 24.0965 $w=3.28e-07 $l=6.9e-07 $layer=LI1_cond $X=9.74 $Y=2.125
+ $X2=9.74 $Y2=2.815
r239 45 129 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.74 $Y=3.245
+ $X2=9.74 $Y2=3.33
r240 45 50 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=9.74 $Y=3.245
+ $X2=9.74 $Y2=2.815
r241 41 126 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.86 $Y=3.245
+ $X2=7.86 $Y2=3.33
r242 41 43 6.80989 $w=3.28e-07 $l=1.95e-07 $layer=LI1_cond $X=7.86 $Y=3.245
+ $X2=7.86 $Y2=3.05
r243 37 66 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.27 $Y=3.245
+ $X2=5.27 $Y2=3.33
r244 37 39 16.5882 $w=3.28e-07 $l=4.75e-07 $layer=LI1_cond $X=5.27 $Y=3.245
+ $X2=5.27 $Y2=2.77
r245 33 63 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.88 $Y=3.245
+ $X2=3.88 $Y2=3.33
r246 33 35 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=3.88 $Y=3.245
+ $X2=3.88 $Y2=2.815
r247 29 123 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.52 $Y=3.245
+ $X2=2.52 $Y2=3.33
r248 29 31 20.744 $w=2.48e-07 $l=4.5e-07 $layer=LI1_cond $X=2.52 $Y=3.245
+ $X2=2.52 $Y2=2.795
r249 25 120 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.08 $Y=3.245
+ $X2=1.08 $Y2=3.33
r250 25 27 20.283 $w=2.48e-07 $l=4.4e-07 $layer=LI1_cond $X=1.08 $Y=3.245
+ $X2=1.08 $Y2=2.805
r251 8 60 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=13.475
+ $Y=1.84 $X2=13.625 $Y2=2.815
r252 8 57 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=13.475
+ $Y=1.84 $X2=13.625 $Y2=1.985
r253 7 53 300 $w=1.7e-07 $l=7.29657e-07 $layer=licon1_PDIFF $count=2 $X=11.51
+ $Y=2.215 $X2=12.115 $Y2=2.49
r254 6 50 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=9.595
+ $Y=1.96 $X2=9.74 $Y2=2.815
r255 6 47 400 $w=1.7e-07 $l=2.26164e-07 $layer=licon1_PDIFF $count=1 $X=9.595
+ $Y=1.96 $X2=9.74 $Y2=2.125
r256 5 43 600 $w=1.7e-07 $l=6.16401e-07 $layer=licon1_PDIFF $count=1 $X=7.625
+ $Y=2.54 $X2=7.86 $Y2=3.05
r257 4 39 600 $w=1.7e-07 $l=1.0099e-06 $layer=licon1_PDIFF $count=1 $X=5.125
+ $Y=1.83 $X2=5.27 $Y2=2.77
r258 3 35 600 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=3.735
+ $Y=1.84 $X2=3.88 $Y2=2.815
r259 2 31 600 $w=1.7e-07 $l=6.58122e-07 $layer=licon1_PDIFF $count=1 $X=2.1
+ $Y=2.3 $X2=2.48 $Y2=2.795
r260 1 27 600 $w=1.7e-07 $l=3.31625e-07 $layer=licon1_PDIFF $count=1 $X=0.97
+ $Y=2.54 $X2=1.12 $Y2=2.805
.ends

.subckt PM_SKY130_FD_SC_HS__EDFXBP_1%Q 1 2 10 13 14 15 22 32
c33 32 0 7.45843e-20 $X=13.132 $Y=1.82
r34 20 22 0.222158 $w=4.13e-07 $l=8e-09 $layer=LI1_cond $X=13.132 $Y=2.027
+ $X2=13.132 $Y2=2.035
r35 14 15 10.2748 $w=4.13e-07 $l=3.7e-07 $layer=LI1_cond $X=13.132 $Y=2.405
+ $X2=13.132 $Y2=2.775
r36 13 20 1.16633 $w=4.13e-07 $l=4.2e-08 $layer=LI1_cond $X=13.132 $Y=1.985
+ $X2=13.132 $Y2=2.027
r37 13 32 8.71334 $w=4.13e-07 $l=1.65e-07 $layer=LI1_cond $X=13.132 $Y=1.985
+ $X2=13.132 $Y2=1.82
r38 13 14 9.21954 $w=4.13e-07 $l=3.32e-07 $layer=LI1_cond $X=13.132 $Y=2.073
+ $X2=13.132 $Y2=2.405
r39 13 22 1.05525 $w=4.13e-07 $l=3.8e-08 $layer=LI1_cond $X=13.132 $Y=2.073
+ $X2=13.132 $Y2=2.035
r40 12 32 53.4973 $w=1.68e-07 $l=8.2e-07 $layer=LI1_cond $X=13.01 $Y=1 $X2=13.01
+ $Y2=1.82
r41 10 12 9.33524 $w=3.28e-07 $l=1.9e-07 $layer=LI1_cond $X=12.93 $Y=0.81
+ $X2=12.93 $Y2=1
r42 2 13 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=13.03
+ $Y=1.84 $X2=13.175 $Y2=1.985
r43 2 15 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=13.03
+ $Y=1.84 $X2=13.175 $Y2=2.815
r44 1 10 182 $w=1.7e-07 $l=4.87134e-07 $layer=licon1_NDIFF $count=1 $X=12.785
+ $Y=0.39 $X2=12.93 $Y2=0.81
.ends

.subckt PM_SKY130_FD_SC_HS__EDFXBP_1%Q_N 1 2 7 9 15 16 17 28
r20 21 28 1.44055 $w=3.58e-07 $l=4.5e-08 $layer=LI1_cond $X=14.135 $Y=0.97
+ $X2=14.135 $Y2=0.925
r21 17 30 8.35096 $w=3.58e-07 $l=1.6e-07 $layer=LI1_cond $X=14.135 $Y=0.99
+ $X2=14.135 $Y2=1.15
r22 17 21 0.640246 $w=3.58e-07 $l=2e-08 $layer=LI1_cond $X=14.135 $Y=0.99
+ $X2=14.135 $Y2=0.97
r23 17 28 0.640246 $w=3.58e-07 $l=2e-08 $layer=LI1_cond $X=14.135 $Y=0.905
+ $X2=14.135 $Y2=0.925
r24 16 17 11.8446 $w=3.58e-07 $l=3.7e-07 $layer=LI1_cond $X=14.135 $Y=0.535
+ $X2=14.135 $Y2=0.905
r25 15 30 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=14.23 $Y=1.82
+ $X2=14.23 $Y2=1.15
r26 9 11 29.4316 $w=3.23e-07 $l=8.3e-07 $layer=LI1_cond $X=14.152 $Y=1.985
+ $X2=14.152 $Y2=2.815
r27 7 15 8.35379 $w=3.23e-07 $l=1.62e-07 $layer=LI1_cond $X=14.152 $Y=1.982
+ $X2=14.152 $Y2=1.82
r28 7 9 0.106379 $w=3.23e-07 $l=3e-09 $layer=LI1_cond $X=14.152 $Y=1.982
+ $X2=14.152 $Y2=1.985
r29 2 11 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=13.925
+ $Y=1.84 $X2=14.075 $Y2=2.815
r30 2 9 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=13.925
+ $Y=1.84 $X2=14.075 $Y2=1.985
r31 1 16 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=13.98
+ $Y=0.39 $X2=14.12 $Y2=0.535
.ends

.subckt PM_SKY130_FD_SC_HS__EDFXBP_1%VGND 1 2 3 4 5 6 7 8 27 31 35 39 43 47 51
+ 55 58 59 61 62 64 65 66 68 86 93 98 103 110 111 114 117 120 123 126
r153 126 127 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=13.68 $Y=0
+ $X2=13.68 $Y2=0
r154 123 124 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.76 $Y=0
+ $X2=11.76 $Y2=0
r155 120 121 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=8.88 $Y=0
+ $X2=8.88 $Y2=0
r156 117 118 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=7.44 $Y=0
+ $X2=7.44 $Y2=0
r157 114 115 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r158 111 127 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=14.16 $Y=0
+ $X2=13.68 $Y2=0
r159 110 111 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=14.16 $Y=0
+ $X2=14.16 $Y2=0
r160 108 126 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=13.775 $Y=0
+ $X2=13.69 $Y2=0
r161 108 110 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=13.775 $Y=0
+ $X2=14.16 $Y2=0
r162 107 127 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=12.24 $Y=0
+ $X2=13.68 $Y2=0
r163 107 124 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.24 $Y=0
+ $X2=11.76 $Y2=0
r164 106 107 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=12.24 $Y=0
+ $X2=12.24 $Y2=0
r165 104 123 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.985 $Y=0
+ $X2=11.82 $Y2=0
r166 104 106 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=11.985 $Y=0
+ $X2=12.24 $Y2=0
r167 103 126 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=13.605 $Y=0
+ $X2=13.69 $Y2=0
r168 103 106 89.0535 $w=1.68e-07 $l=1.365e-06 $layer=LI1_cond $X=13.605 $Y=0
+ $X2=12.24 $Y2=0
r169 102 124 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.28 $Y=0
+ $X2=11.76 $Y2=0
r170 102 121 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=11.28 $Y=0
+ $X2=8.88 $Y2=0
r171 101 102 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=11.28 $Y=0
+ $X2=11.28 $Y2=0
r172 99 120 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.91 $Y=0
+ $X2=8.785 $Y2=0
r173 99 101 154.62 $w=1.68e-07 $l=2.37e-06 $layer=LI1_cond $X=8.91 $Y=0
+ $X2=11.28 $Y2=0
r174 98 123 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.655 $Y=0
+ $X2=11.82 $Y2=0
r175 98 101 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=11.655 $Y=0
+ $X2=11.28 $Y2=0
r176 97 121 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=0 $X2=8.88
+ $Y2=0
r177 97 118 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=8.4 $Y=0 $X2=7.44
+ $Y2=0
r178 96 97 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r179 94 117 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.47 $Y=0
+ $X2=7.345 $Y2=0
r180 94 96 60.6738 $w=1.68e-07 $l=9.3e-07 $layer=LI1_cond $X=7.47 $Y=0 $X2=8.4
+ $Y2=0
r181 93 120 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.66 $Y=0
+ $X2=8.785 $Y2=0
r182 93 96 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=8.66 $Y=0 $X2=8.4
+ $Y2=0
r183 91 92 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6.96 $Y=0
+ $X2=6.96 $Y2=0
r184 89 92 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=5.04 $Y=0
+ $X2=6.96 $Y2=0
r185 88 91 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=5.04 $Y=0 $X2=6.96
+ $Y2=0
r186 88 89 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=5.04 $Y=0
+ $X2=5.04 $Y2=0
r187 86 117 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.22 $Y=0
+ $X2=7.345 $Y2=0
r188 86 91 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=7.22 $Y=0 $X2=6.96
+ $Y2=0
r189 85 89 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=5.04
+ $Y2=0
r190 84 85 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r191 82 85 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.56
+ $Y2=0
r192 81 82 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r193 79 82 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.6
+ $Y2=0
r194 78 81 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=2.64 $Y=0 $X2=3.6
+ $Y2=0
r195 78 79 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r196 76 79 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r197 76 115 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.2
+ $Y2=0
r198 75 76 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r199 73 114 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.42 $Y=0
+ $X2=1.255 $Y2=0
r200 73 75 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=1.42 $Y=0 $X2=2.16
+ $Y2=0
r201 71 115 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r202 70 71 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r203 68 114 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.09 $Y=0
+ $X2=1.255 $Y2=0
r204 68 70 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=1.09 $Y=0 $X2=0.72
+ $Y2=0
r205 66 118 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=7.2 $Y=0
+ $X2=7.44 $Y2=0
r206 66 92 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=7.2 $Y=0 $X2=6.96
+ $Y2=0
r207 64 84 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=4.585 $Y=0 $X2=4.56
+ $Y2=0
r208 64 65 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.585 $Y=0 $X2=4.75
+ $Y2=0
r209 63 88 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=4.915 $Y=0
+ $X2=5.04 $Y2=0
r210 63 65 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.915 $Y=0 $X2=4.75
+ $Y2=0
r211 61 81 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=3.715 $Y=0 $X2=3.6
+ $Y2=0
r212 61 62 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.715 $Y=0 $X2=3.8
+ $Y2=0
r213 60 84 44.0374 $w=1.68e-07 $l=6.75e-07 $layer=LI1_cond $X=3.885 $Y=0
+ $X2=4.56 $Y2=0
r214 60 62 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.885 $Y=0 $X2=3.8
+ $Y2=0
r215 58 75 0.652406 $w=1.68e-07 $l=1e-08 $layer=LI1_cond $X=2.17 $Y=0 $X2=2.16
+ $Y2=0
r216 58 59 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.17 $Y=0 $X2=2.335
+ $Y2=0
r217 57 78 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=2.5 $Y=0 $X2=2.64
+ $Y2=0
r218 57 59 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.5 $Y=0 $X2=2.335
+ $Y2=0
r219 53 126 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=13.69 $Y=0.085
+ $X2=13.69 $Y2=0
r220 53 55 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=13.69 $Y=0.085
+ $X2=13.69 $Y2=0.535
r221 49 123 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=11.82 $Y=0.085
+ $X2=11.82 $Y2=0
r222 49 51 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=11.82 $Y=0.085
+ $X2=11.82 $Y2=0.515
r223 45 120 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=8.785 $Y=0.085
+ $X2=8.785 $Y2=0
r224 45 47 23.5098 $w=2.48e-07 $l=5.1e-07 $layer=LI1_cond $X=8.785 $Y=0.085
+ $X2=8.785 $Y2=0.595
r225 41 117 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=7.345 $Y=0.085
+ $X2=7.345 $Y2=0
r226 41 43 25.1233 $w=2.48e-07 $l=5.45e-07 $layer=LI1_cond $X=7.345 $Y=0.085
+ $X2=7.345 $Y2=0.63
r227 37 65 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.75 $Y=0.085
+ $X2=4.75 $Y2=0
r228 37 39 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=4.75 $Y=0.085
+ $X2=4.75 $Y2=0.55
r229 33 62 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.8 $Y=0.085 $X2=3.8
+ $Y2=0
r230 33 35 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=3.8 $Y=0.085
+ $X2=3.8 $Y2=0.505
r231 29 59 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.335 $Y=0.085
+ $X2=2.335 $Y2=0
r232 29 31 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=2.335 $Y=0.085
+ $X2=2.335 $Y2=0.58
r233 25 114 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.255 $Y=0.085
+ $X2=1.255 $Y2=0
r234 25 27 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=1.255 $Y=0.085
+ $X2=1.255 $Y2=0.58
r235 8 55 91 $w=1.7e-07 $l=5.37634e-07 $layer=licon1_NDIFF $count=2 $X=13.22
+ $Y=0.39 $X2=13.69 $Y2=0.535
r236 7 51 91 $w=1.7e-07 $l=3.30379e-07 $layer=licon1_NDIFF $count=2 $X=11.525
+ $Y=0.59 $X2=11.82 $Y2=0.515
r237 6 47 182 $w=1.7e-07 $l=2.88531e-07 $layer=licon1_NDIFF $count=1 $X=8.6
+ $Y=0.37 $X2=8.745 $Y2=0.595
r238 5 43 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=7.245
+ $Y=0.485 $X2=7.385 $Y2=0.63
r239 4 39 182 $w=1.7e-07 $l=2.34307e-07 $layer=licon1_NDIFF $count=1 $X=4.625
+ $Y=0.37 $X2=4.75 $Y2=0.55
r240 3 35 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=3.655
+ $Y=0.37 $X2=3.8 $Y2=0.505
r241 2 31 182 $w=1.7e-07 $l=2.96985e-07 $layer=licon1_NDIFF $count=1 $X=2.125
+ $Y=0.37 $X2=2.335 $Y2=0.58
r242 1 27 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.115
+ $Y=0.37 $X2=1.255 $Y2=0.58
.ends

