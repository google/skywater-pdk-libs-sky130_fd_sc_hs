# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_hs__a211oi_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.800000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.558000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.180000 0.480000 1.550000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.558000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.085000 1.430000 2.275000 1.780000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.447000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.005000 1.180000 3.715000 1.550000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.447000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.965000 1.180000 4.675000 1.550000 ;
    END
  END C1
  PIN Y
    ANTENNADIFFAREA  1.076000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.650000 0.635000 0.830000 1.090000 ;
        RECT 0.650000 1.090000 2.755000 1.260000 ;
        RECT 2.525000 1.260000 2.755000 1.720000 ;
        RECT 2.525000 1.720000 4.145000 1.890000 ;
        RECT 2.585000 0.840000 3.590000 1.010000 ;
        RECT 2.585000 1.010000 2.755000 1.090000 ;
        RECT 2.960000 0.330000 3.590000 0.840000 ;
        RECT 3.815000 1.890000 4.145000 2.735000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 4.800000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 4.800000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.800000 0.085000 ;
      RECT 0.000000  3.245000 4.800000 3.415000 ;
      RECT 0.105000  1.820000 0.355000 3.245000 ;
      RECT 0.150000  0.255000 1.260000 0.425000 ;
      RECT 0.150000  0.425000 0.480000 1.010000 ;
      RECT 0.555000  1.820000 0.805000 1.950000 ;
      RECT 0.555000  1.950000 2.355000 2.060000 ;
      RECT 0.555000  2.060000 3.245000 2.120000 ;
      RECT 0.555000  2.120000 0.805000 2.980000 ;
      RECT 1.005000  2.290000 1.335000 3.245000 ;
      RECT 1.010000  0.425000 1.260000 0.750000 ;
      RECT 1.010000  0.750000 2.240000 0.920000 ;
      RECT 1.440000  0.085000 1.610000 0.330000 ;
      RECT 1.440000  0.330000 1.810000 0.580000 ;
      RECT 1.535000  2.120000 3.245000 2.230000 ;
      RECT 1.535000  2.230000 1.705000 2.980000 ;
      RECT 1.905000  2.400000 2.235000 3.245000 ;
      RECT 1.990000  0.330000 2.240000 0.750000 ;
      RECT 2.460000  0.085000 2.790000 0.670000 ;
      RECT 2.465000  2.400000 2.795000 2.905000 ;
      RECT 2.465000  2.905000 4.595000 3.075000 ;
      RECT 2.965000  2.230000 3.245000 2.735000 ;
      RECT 3.445000  2.060000 3.615000 2.905000 ;
      RECT 3.760000  0.085000 4.090000 1.010000 ;
      RECT 4.345000  1.820000 4.595000 2.905000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
  END
END sky130_fd_sc_hs__a211oi_2
END LIBRARY
