* File: sky130_fd_sc_hs__clkinv_16.spice
* Created: Tue Sep  1 19:58:34 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hs__clkinv_16.pex.spice"
.subckt sky130_fd_sc_hs__clkinv_16  VNB VPB A VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A	A
* VPB	VPB
* VNB	VNB
MM1000 N_Y_M1000_d N_A_M1000_g N_VGND_M1000_s VNB NLOWVT L=0.15 W=0.42 AD=0.0588
+ AS=0.1197 PD=0.7 PS=1.41 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2 SB=75008.5 A=0.063
+ P=1.14 MULT=1
MM1001 N_Y_M1000_d N_A_M1001_g N_VGND_M1001_s VNB NLOWVT L=0.15 W=0.42 AD=0.0588
+ AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6 SB=75008.1 A=0.063
+ P=1.14 MULT=1
MM1005 N_Y_M1005_d N_A_M1005_g N_VGND_M1001_s VNB NLOWVT L=0.15 W=0.42 AD=0.0588
+ AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75001.1 SB=75007.6 A=0.063
+ P=1.14 MULT=1
MM1008 N_Y_M1005_d N_A_M1008_g N_VGND_M1008_s VNB NLOWVT L=0.15 W=0.42 AD=0.0588
+ AS=0.0735 PD=0.7 PS=0.77 NRD=0 NRS=0 M=1 R=2.8 SA=75001.5 SB=75007.2 A=0.063
+ P=1.14 MULT=1
MM1009 N_Y_M1009_d N_A_M1009_g N_VGND_M1008_s VNB NLOWVT L=0.15 W=0.42 AD=0.0588
+ AS=0.0735 PD=0.7 PS=0.77 NRD=0 NRS=19.992 M=1 R=2.8 SA=75002 SB=75006.7
+ A=0.063 P=1.14 MULT=1
MM1014 N_Y_M1009_d N_A_M1014_g N_VGND_M1014_s VNB NLOWVT L=0.15 W=0.42 AD=0.0588
+ AS=0.0735 PD=0.7 PS=0.77 NRD=0 NRS=0 M=1 R=2.8 SA=75002.4 SB=75006.3 A=0.063
+ P=1.14 MULT=1
MM1016 N_Y_M1016_d N_A_M1016_g N_VGND_M1014_s VNB NLOWVT L=0.15 W=0.42 AD=0.0588
+ AS=0.0735 PD=0.7 PS=0.77 NRD=0 NRS=19.992 M=1 R=2.8 SA=75002.9 SB=75005.8
+ A=0.063 P=1.14 MULT=1
MM1017 N_Y_M1016_d N_A_M1017_g N_VGND_M1017_s VNB NLOWVT L=0.15 W=0.42 AD=0.0588
+ AS=0.0882 PD=0.7 PS=0.84 NRD=0 NRS=19.992 M=1 R=2.8 SA=75003.4 SB=75005.4
+ A=0.063 P=1.14 MULT=1
MM1022 N_Y_M1022_d N_A_M1022_g N_VGND_M1017_s VNB NLOWVT L=0.15 W=0.42 AD=0.0588
+ AS=0.0882 PD=0.7 PS=0.84 NRD=0 NRS=19.992 M=1 R=2.8 SA=75003.9 SB=75004.8
+ A=0.063 P=1.14 MULT=1
MM1027 N_Y_M1022_d N_A_M1027_g N_VGND_M1027_s VNB NLOWVT L=0.15 W=0.42 AD=0.0588
+ AS=0.0882 PD=0.7 PS=0.84 NRD=0 NRS=19.992 M=1 R=2.8 SA=75004.4 SB=75004.4
+ A=0.063 P=1.14 MULT=1
MM1028 N_Y_M1028_d N_A_M1028_g N_VGND_M1027_s VNB NLOWVT L=0.15 W=0.42 AD=0.0588
+ AS=0.0882 PD=0.7 PS=0.84 NRD=0 NRS=19.992 M=1 R=2.8 SA=75004.9 SB=75003.8
+ A=0.063 P=1.14 MULT=1
MM1030 N_Y_M1028_d N_A_M1030_g N_VGND_M1030_s VNB NLOWVT L=0.15 W=0.42 AD=0.0588
+ AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75005.4 SB=75003.4 A=0.063
+ P=1.14 MULT=1
MM1032 N_Y_M1032_d N_A_M1032_g N_VGND_M1030_s VNB NLOWVT L=0.15 W=0.42 AD=0.0588
+ AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75005.8 SB=75002.9 A=0.063
+ P=1.14 MULT=1
MM1036 N_Y_M1032_d N_A_M1036_g N_VGND_M1036_s VNB NLOWVT L=0.15 W=0.42 AD=0.0588
+ AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75006.2 SB=75002.5 A=0.063
+ P=1.14 MULT=1
MM1037 N_Y_M1037_d N_A_M1037_g N_VGND_M1036_s VNB NLOWVT L=0.15 W=0.42 AD=0.0588
+ AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75006.6 SB=75002.1 A=0.063
+ P=1.14 MULT=1
MM1038 N_Y_M1037_d N_A_M1038_g N_VGND_M1038_s VNB NLOWVT L=0.15 W=0.42 AD=0.0588
+ AS=0.71835 PD=0.7 PS=5.57 NRD=0 NRS=19.992 M=1 R=2.8 SA=75007.1 SB=75001.6
+ A=0.063 P=1.14 MULT=1
MM1002 N_Y_M1002_d N_A_M1002_g N_VPWR_M1002_s VPB PSHORT L=0.15 W=1.12 AD=0.168
+ AS=0.3304 PD=1.42 PS=2.83 NRD=1.7533 NRS=1.7533 M=1 R=7.46667 SA=75000.2
+ SB=75010.7 A=0.168 P=2.54 MULT=1
MM1003 N_Y_M1002_d N_A_M1003_g N_VPWR_M1003_s VPB PSHORT L=0.15 W=1.12 AD=0.168
+ AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667 SA=75000.7
+ SB=75010.3 A=0.168 P=2.54 MULT=1
MM1004 N_Y_M1004_d N_A_M1004_g N_VPWR_M1003_s VPB PSHORT L=0.15 W=1.12 AD=0.168
+ AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667 SA=75001.1
+ SB=75009.8 A=0.168 P=2.54 MULT=1
MM1006 N_Y_M1004_d N_A_M1006_g N_VPWR_M1006_s VPB PSHORT L=0.15 W=1.12 AD=0.168
+ AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667 SA=75001.6
+ SB=75009.4 A=0.168 P=2.54 MULT=1
MM1007 N_Y_M1007_d N_A_M1007_g N_VPWR_M1006_s VPB PSHORT L=0.15 W=1.12 AD=0.168
+ AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667 SA=75002
+ SB=75008.9 A=0.168 P=2.54 MULT=1
MM1010 N_Y_M1007_d N_A_M1010_g N_VPWR_M1010_s VPB PSHORT L=0.15 W=1.12 AD=0.168
+ AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667 SA=75002.5
+ SB=75008.5 A=0.168 P=2.54 MULT=1
MM1011 N_Y_M1011_d N_A_M1011_g N_VPWR_M1010_s VPB PSHORT L=0.15 W=1.12 AD=0.168
+ AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667 SA=75002.9
+ SB=75008 A=0.168 P=2.54 MULT=1
MM1012 N_Y_M1011_d N_A_M1012_g N_VPWR_M1012_s VPB PSHORT L=0.15 W=1.12 AD=0.168
+ AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667 SA=75003.4
+ SB=75007.6 A=0.168 P=2.54 MULT=1
MM1013 N_Y_M1013_d N_A_M1013_g N_VPWR_M1012_s VPB PSHORT L=0.15 W=1.12 AD=0.168
+ AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667 SA=75003.8
+ SB=75007.1 A=0.168 P=2.54 MULT=1
MM1015 N_Y_M1013_d N_A_M1015_g N_VPWR_M1015_s VPB PSHORT L=0.15 W=1.12 AD=0.168
+ AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667 SA=75004.3
+ SB=75006.7 A=0.168 P=2.54 MULT=1
MM1018 N_Y_M1018_d N_A_M1018_g N_VPWR_M1015_s VPB PSHORT L=0.15 W=1.12 AD=0.168
+ AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667 SA=75004.7
+ SB=75006.2 A=0.168 P=2.54 MULT=1
MM1019 N_Y_M1018_d N_A_M1019_g N_VPWR_M1019_s VPB PSHORT L=0.15 W=1.12 AD=0.168
+ AS=0.196 PD=1.42 PS=1.47 NRD=1.7533 NRS=1.7533 M=1 R=7.46667 SA=75005.2
+ SB=75005.8 A=0.168 P=2.54 MULT=1
MM1020 N_Y_M1020_d N_A_M1020_g N_VPWR_M1019_s VPB PSHORT L=0.15 W=1.12 AD=0.168
+ AS=0.196 PD=1.42 PS=1.47 NRD=1.7533 NRS=10.5395 M=1 R=7.46667 SA=75005.7
+ SB=75005.3 A=0.168 P=2.54 MULT=1
MM1021 N_Y_M1020_d N_A_M1021_g N_VPWR_M1021_s VPB PSHORT L=0.15 W=1.12 AD=0.168
+ AS=0.196 PD=1.42 PS=1.47 NRD=1.7533 NRS=1.7533 M=1 R=7.46667 SA=75006.1
+ SB=75004.8 A=0.168 P=2.54 MULT=1
MM1023 N_Y_M1023_d N_A_M1023_g N_VPWR_M1021_s VPB PSHORT L=0.15 W=1.12 AD=0.2016
+ AS=0.196 PD=1.48 PS=1.47 NRD=7.0329 NRS=10.5395 M=1 R=7.46667 SA=75006.6
+ SB=75004.3 A=0.168 P=2.54 MULT=1
MM1024 N_Y_M1023_d N_A_M1024_g N_VPWR_M1024_s VPB PSHORT L=0.15 W=1.12 AD=0.2016
+ AS=0.168 PD=1.48 PS=1.42 NRD=7.0329 NRS=1.7533 M=1 R=7.46667 SA=75007.1
+ SB=75003.8 A=0.168 P=2.54 MULT=1
MM1025 N_Y_M1025_d N_A_M1025_g N_VPWR_M1024_s VPB PSHORT L=0.15 W=1.12 AD=0.168
+ AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667 SA=75007.6
+ SB=75003.4 A=0.168 P=2.54 MULT=1
MM1026 N_Y_M1025_d N_A_M1026_g N_VPWR_M1026_s VPB PSHORT L=0.15 W=1.12 AD=0.168
+ AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667 SA=75008
+ SB=75002.9 A=0.168 P=2.54 MULT=1
MM1029 N_Y_M1029_d N_A_M1029_g N_VPWR_M1026_s VPB PSHORT L=0.15 W=1.12 AD=0.168
+ AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667 SA=75008.5
+ SB=75002.5 A=0.168 P=2.54 MULT=1
MM1031 N_Y_M1029_d N_A_M1031_g N_VPWR_M1031_s VPB PSHORT L=0.15 W=1.12 AD=0.168
+ AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667 SA=75008.9
+ SB=75002 A=0.168 P=2.54 MULT=1
MM1033 N_Y_M1033_d N_A_M1033_g N_VPWR_M1031_s VPB PSHORT L=0.15 W=1.12 AD=0.168
+ AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667 SA=75009.4
+ SB=75001.6 A=0.168 P=2.54 MULT=1
MM1034 N_Y_M1033_d N_A_M1034_g N_VPWR_M1034_s VPB PSHORT L=0.15 W=1.12 AD=0.168
+ AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667 SA=75009.8
+ SB=75001.1 A=0.168 P=2.54 MULT=1
MM1035 N_Y_M1035_d N_A_M1035_g N_VPWR_M1034_s VPB PSHORT L=0.15 W=1.12 AD=0.168
+ AS=0.168 PD=1.42 PS=1.42 NRD=1.7533 NRS=1.7533 M=1 R=7.46667 SA=75010.3
+ SB=75000.7 A=0.168 P=2.54 MULT=1
MM1039 N_Y_M1035_d N_A_M1039_g N_VPWR_M1039_s VPB PSHORT L=0.15 W=1.12 AD=0.168
+ AS=0.3304 PD=1.42 PS=2.83 NRD=1.7533 NRS=1.7533 M=1 R=7.46667 SA=75010.7
+ SB=75000.2 A=0.168 P=2.54 MULT=1
DX40_noxref VNB VPB NWDIODE A=22.134 P=27.52
*
.include "sky130_fd_sc_hs__clkinv_16.pxi.spice"
*
.ends
*
*
