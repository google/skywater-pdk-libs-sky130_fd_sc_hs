* File: sky130_fd_sc_hs__sdlclkp_2.spice
* Created: Tue Sep  1 20:24:07 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hs__sdlclkp_2.pex.spice"
.subckt sky130_fd_sc_hs__sdlclkp_2  VNB VPB SCE GATE CLK VPWR GCLK VGND
* 
* VGND	VGND
* GCLK	GCLK
* VPWR	VPWR
* CLK	CLK
* GATE	GATE
* SCE	SCE
* VPB	VPB
* VNB	VNB
MM1013 N_A_114_112#_M1013_d N_SCE_M1013_g N_VGND_M1013_s VNB NLOWVT L=0.15
+ W=0.55 AD=0.077 AS=0.15675 PD=0.83 PS=1.67 NRD=0 NRS=0 M=1 R=3.66667
+ SA=75000.2 SB=75001.2 A=0.0825 P=1.4 MULT=1
MM1012 N_VGND_M1012_d N_GATE_M1012_g N_A_114_112#_M1013_d VNB NLOWVT L=0.15
+ W=0.55 AD=0.161184 AS=0.077 PD=1.20233 PS=0.83 NRD=51.936 NRS=0 M=1 R=3.66667
+ SA=75000.6 SB=75000.8 A=0.0825 P=1.4 MULT=1
MM1002 N_A_318_74#_M1002_d N_A_288_48#_M1002_g N_VGND_M1012_d VNB NLOWVT L=0.15
+ W=0.74 AD=0.2109 AS=0.216866 PD=2.05 PS=1.61767 NRD=0 NRS=38.604 M=1 R=4.93333
+ SA=75001 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1023 N_A_580_74#_M1023_d N_A_288_48#_M1023_g N_A_114_112#_M1023_s VNB NLOWVT
+ L=0.15 W=0.55 AD=0.110425 AS=0.33275 PD=1.04897 PS=2.31 NRD=2.172 NRS=69.816
+ M=1 R=3.66667 SA=75000.5 SB=75001.4 A=0.0825 P=1.4 MULT=1
MM1018 A_685_81# N_A_318_74#_M1018_g N_A_580_74#_M1023_d VNB NLOWVT L=0.15
+ W=0.42 AD=0.0504 AS=0.0843247 PD=0.66 PS=0.801031 NRD=18.564 NRS=24.276 M=1
+ R=2.8 SA=75001.1 SB=75001.3 A=0.063 P=1.14 MULT=1
MM1019 N_VGND_M1019_d N_A_706_317#_M1019_g A_685_81# VNB NLOWVT L=0.15 W=0.42
+ AD=0.109562 AS=0.0504 PD=0.919655 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8
+ SA=75001.4 SB=75000.9 A=0.063 P=1.14 MULT=1
MM1001 N_A_706_317#_M1001_d N_A_580_74#_M1001_g N_VGND_M1019_d VNB NLOWVT L=0.15
+ W=0.74 AD=0.2109 AS=0.193038 PD=2.05 PS=1.62034 NRD=0 NRS=40.536 M=1 R=4.93333
+ SA=75001.3 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1000 N_VGND_M1000_d N_CLK_M1000_g N_A_288_48#_M1000_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.13135 AS=0.2109 PD=1.095 PS=2.05 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75001.1 A=0.111 P=1.78 MULT=1
MM1015 A_1198_74# N_CLK_M1015_g N_VGND_M1000_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.0777 AS=0.13135 PD=0.95 PS=1.095 NRD=8.1 NRS=0.804 M=1 R=4.93333
+ SA=75000.7 SB=75000.6 A=0.111 P=1.78 MULT=1
MM1010 N_A_1195_374#_M1010_d N_A_706_317#_M1010_g A_1198_74# VNB NLOWVT L=0.15
+ W=0.74 AD=0.2035 AS=0.0777 PD=2.03 PS=0.95 NRD=0 NRS=8.1 M=1 R=4.93333
+ SA=75001.1 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1007 N_GCLK_M1007_d N_A_1195_374#_M1007_g N_VGND_M1007_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.2035 PD=1.02 PS=2.03 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75000.6 A=0.111 P=1.78 MULT=1
MM1016 N_GCLK_M1007_d N_A_1195_374#_M1016_g N_VGND_M1016_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.2035 PD=1.02 PS=2.03 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.6 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1005 A_114_424# N_SCE_M1005_g N_VPWR_M1005_s VPB PSHORT L=0.15 W=0.84
+ AD=0.1008 AS=0.2394 PD=1.08 PS=2.25 NRD=15.2281 NRS=2.3443 M=1 R=5.6
+ SA=75000.2 SB=75000.6 A=0.126 P=1.98 MULT=1
MM1022 N_A_114_112#_M1022_d N_GATE_M1022_g A_114_424# VPB PSHORT L=0.15 W=0.84
+ AD=0.2394 AS=0.1008 PD=2.25 PS=1.08 NRD=2.3443 NRS=15.2281 M=1 R=5.6
+ SA=75000.6 SB=75000.2 A=0.126 P=1.98 MULT=1
MM1020 N_A_318_74#_M1020_d N_A_288_48#_M1020_g N_VPWR_M1020_s VPB PSHORT L=0.15
+ W=0.84 AD=0.2394 AS=0.3807 PD=2.25 PS=2.98 NRD=2.3443 NRS=93.378 M=1 R=5.6
+ SA=75000.3 SB=75000.2 A=0.126 P=1.98 MULT=1
MM1008 N_A_580_74#_M1008_d N_A_318_74#_M1008_g N_A_114_112#_M1008_s VPB PSHORT
+ L=0.15 W=0.84 AD=0.1848 AS=0.2394 PD=1.62 PS=2.25 NRD=2.3443 NRS=2.3443 M=1
+ R=5.6 SA=75000.2 SB=75000.9 A=0.126 P=1.98 MULT=1
MM1021 A_708_451# N_A_288_48#_M1021_g N_A_580_74#_M1008_d VPB PSHORT L=0.15
+ W=0.42 AD=0.0504 AS=0.0924 PD=0.66 PS=0.81 NRD=30.4759 NRS=39.8531 M=1 R=2.8
+ SA=75000.7 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1011 N_VPWR_M1011_d N_A_706_317#_M1011_g A_708_451# VPB PSHORT L=0.15 W=0.42
+ AD=0.0973636 AS=0.0504 PD=0.815455 PS=0.66 NRD=42.1974 NRS=30.4759 M=1 R=2.8
+ SA=75001.1 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1014 N_A_706_317#_M1014_d N_A_580_74#_M1014_g N_VPWR_M1011_d VPB PSHORT L=0.15
+ W=1.12 AD=0.3192 AS=0.259636 PD=2.81 PS=2.17455 NRD=1.7533 NRS=1.7533 M=1
+ R=7.46667 SA=75000.7 SB=75000.2 A=0.168 P=2.54 MULT=1
MM1017 N_VPWR_M1017_d N_CLK_M1017_g N_A_288_48#_M1017_s VPB PSHORT L=0.15 W=0.84
+ AD=0.17729 AS=0.2394 PD=1.3787 PS=2.25 NRD=36.5829 NRS=2.3443 M=1 R=5.6
+ SA=75000.2 SB=75002.1 A=0.126 P=1.98 MULT=1
MM1003 N_A_1195_374#_M1003_d N_CLK_M1003_g N_VPWR_M1017_d VPB PSHORT L=0.15 W=1
+ AD=0.2575 AS=0.21106 PD=1.515 PS=1.6413 NRD=44.325 NRS=1.9503 M=1 R=6.66667
+ SA=75000.6 SB=75001.9 A=0.15 P=2.3 MULT=1
MM1004 N_VPWR_M1004_d N_A_706_317#_M1004_g N_A_1195_374#_M1003_d VPB PSHORT
+ L=0.15 W=1 AD=0.223585 AS=0.2575 PD=1.46698 PS=1.515 NRD=19.2075 NRS=1.9503
+ M=1 R=6.66667 SA=75001.3 SB=75001.3 A=0.15 P=2.3 MULT=1
MM1006 N_GCLK_M1006_d N_A_1195_374#_M1006_g N_VPWR_M1004_d VPB PSHORT L=0.15
+ W=1.12 AD=0.168 AS=0.250415 PD=1.42 PS=1.64302 NRD=1.7533 NRS=10.5395 M=1
+ R=7.46667 SA=75001.7 SB=75000.7 A=0.168 P=2.54 MULT=1
MM1009 N_GCLK_M1006_d N_A_1195_374#_M1009_g N_VPWR_M1009_s VPB PSHORT L=0.15
+ W=1.12 AD=0.168 AS=0.3304 PD=1.42 PS=2.83 NRD=1.7533 NRS=1.7533 M=1 R=7.46667
+ SA=75002.1 SB=75000.2 A=0.168 P=2.54 MULT=1
DX24_noxref VNB VPB NWDIODE A=16.0894 P=21
*
.include "sky130_fd_sc_hs__sdlclkp_2.pxi.spice"
*
.ends
*
*
