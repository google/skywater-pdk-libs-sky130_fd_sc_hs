* NGSPICE file created from sky130_fd_sc_hs__sdlclkp_2.ext - technology: sky130A

.subckt sky130_fd_sc_hs__sdlclkp_2 CLK GATE SCE VGND VNB VPB VPWR GCLK
M1000 VGND CLK a_288_48# VNB nlowvt w=740000u l=150000u
+  ad=1.5071e+12p pd=1.328e+07u as=2.109e+11p ps=2.05e+06u
M1001 a_706_317# a_580_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1002 a_318_74# a_288_48# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1003 a_1195_374# CLK VPWR VPB pshort w=1e+06u l=150000u
+  ad=5.15e+11p pd=3.03e+06u as=2.16985e+12p ps=1.718e+07u
M1004 VPWR a_706_317# a_1195_374# VPB pshort w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_114_424# SCE VPWR VPB pshort w=840000u l=150000u
+  ad=2.016e+11p pd=2.16e+06u as=0p ps=0u
M1006 GCLK a_1195_374# VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=3.36e+11p pd=2.84e+06u as=0p ps=0u
M1007 GCLK a_1195_374# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.072e+11p pd=2.04e+06u as=0p ps=0u
M1008 a_580_74# a_318_74# a_114_112# VPB pshort w=840000u l=150000u
+  ad=2.772e+11p pd=2.43e+06u as=4.788e+11p ps=4.5e+06u
M1009 VPWR a_1195_374# GCLK VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_1195_374# a_706_317# a_1198_74# VNB nlowvt w=740000u l=150000u
+  ad=2.035e+11p pd=2.03e+06u as=1.554e+11p ps=1.9e+06u
M1011 VPWR a_706_317# a_708_451# VPB pshort w=420000u l=150000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1012 VGND GATE a_114_112# VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=4.8675e+11p ps=3.97e+06u
M1013 a_114_112# SCE VGND VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_706_317# a_580_74# VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=3.192e+11p pd=2.81e+06u as=0p ps=0u
M1015 a_1198_74# CLK VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VGND a_1195_374# GCLK VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 VPWR CLK a_288_48# VPB pshort w=840000u l=150000u
+  ad=0p pd=0u as=2.394e+11p ps=2.25e+06u
M1018 a_685_81# a_318_74# a_580_74# VNB nlowvt w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=1.9475e+11p ps=1.85e+06u
M1019 VGND a_706_317# a_685_81# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_318_74# a_288_48# VPWR VPB pshort w=840000u l=150000u
+  ad=2.394e+11p pd=2.25e+06u as=0p ps=0u
M1021 a_708_451# a_288_48# a_580_74# VPB pshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_114_112# GATE a_114_424# VPB pshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_580_74# a_288_48# a_114_112# VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

