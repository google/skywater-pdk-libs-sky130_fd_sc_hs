* File: sky130_fd_sc_hs__nor3b_1.pxi.spice
* Created: Tue Sep  1 20:11:44 2020
* 
x_PM_SKY130_FD_SC_HS__NOR3B_1%C_N N_C_N_c_48_n N_C_N_M1001_g N_C_N_c_49_n
+ N_C_N_M1005_g C_N PM_SKY130_FD_SC_HS__NOR3B_1%C_N
x_PM_SKY130_FD_SC_HS__NOR3B_1%A N_A_c_75_n N_A_M1002_g N_A_M1007_g A N_A_c_77_n
+ PM_SKY130_FD_SC_HS__NOR3B_1%A
x_PM_SKY130_FD_SC_HS__NOR3B_1%B N_B_c_104_n N_B_M1004_g N_B_M1006_g B
+ N_B_c_106_n PM_SKY130_FD_SC_HS__NOR3B_1%B
x_PM_SKY130_FD_SC_HS__NOR3B_1%A_27_112# N_A_27_112#_M1005_s N_A_27_112#_M1001_s
+ N_A_27_112#_c_137_n N_A_27_112#_M1003_g N_A_27_112#_M1000_g
+ N_A_27_112#_c_148_n N_A_27_112#_c_143_n N_A_27_112#_c_139_n
+ N_A_27_112#_c_144_n N_A_27_112#_c_140_n N_A_27_112#_c_146_n
+ N_A_27_112#_c_141_n PM_SKY130_FD_SC_HS__NOR3B_1%A_27_112#
x_PM_SKY130_FD_SC_HS__NOR3B_1%VPWR N_VPWR_M1001_d N_VPWR_c_200_n N_VPWR_c_201_n
+ N_VPWR_c_202_n VPWR N_VPWR_c_203_n N_VPWR_c_199_n
+ PM_SKY130_FD_SC_HS__NOR3B_1%VPWR
x_PM_SKY130_FD_SC_HS__NOR3B_1%Y N_Y_M1007_d N_Y_M1000_d N_Y_M1003_d N_Y_c_225_n
+ N_Y_c_226_n N_Y_c_227_n N_Y_c_231_n N_Y_c_228_n Y Y N_Y_c_229_n N_Y_c_230_n
+ PM_SKY130_FD_SC_HS__NOR3B_1%Y
x_PM_SKY130_FD_SC_HS__NOR3B_1%VGND N_VGND_M1005_d N_VGND_M1006_d N_VGND_c_270_n
+ N_VGND_c_271_n N_VGND_c_272_n N_VGND_c_273_n N_VGND_c_274_n N_VGND_c_275_n
+ VGND N_VGND_c_276_n N_VGND_c_277_n PM_SKY130_FD_SC_HS__NOR3B_1%VGND
cc_1 VNB N_C_N_c_48_n 0.0411324f $X=-0.19 $Y=-0.245 $X2=0.655 $Y2=1.765
cc_2 VNB N_C_N_c_49_n 0.0224251f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=1.22
cc_3 VNB C_N 0.0104207f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_4 VNB N_A_c_75_n 0.0267844f $X=-0.19 $Y=-0.245 $X2=0.655 $Y2=1.765
cc_5 VNB N_A_M1007_g 0.0268153f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=0.835
cc_6 VNB N_A_c_77_n 0.0023516f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.365
cc_7 VNB N_B_c_104_n 0.0270077f $X=-0.19 $Y=-0.245 $X2=0.655 $Y2=1.765
cc_8 VNB N_B_M1006_g 0.026332f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=0.835
cc_9 VNB N_B_c_106_n 0.00165701f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.365
cc_10 VNB N_A_27_112#_c_137_n 0.0289667f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_11 VNB N_A_27_112#_M1000_g 0.0321102f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.365
cc_12 VNB N_A_27_112#_c_139_n 0.0138636f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_27_112#_c_140_n 0.0299402f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_27_112#_c_141_n 0.00165828f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_VPWR_c_199_n 0.123877f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_Y_c_225_n 0.00280874f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.365
cc_17 VNB N_Y_c_226_n 0.00951425f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.365
cc_18 VNB N_Y_c_227_n 0.0107024f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_Y_c_228_n 0.0227107f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_Y_c_229_n 0.0332097f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_Y_c_230_n 0.0157047f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_VGND_c_270_n 0.0162763f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.385
cc_23 VNB N_VGND_c_271_n 0.00900728f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_VGND_c_272_n 0.0263417f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_VGND_c_273_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_VGND_c_274_n 0.0186436f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_VGND_c_275_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_276_n 0.0214382f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_277_n 0.188982f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VPB N_C_N_c_48_n 0.0280237f $X=-0.19 $Y=1.66 $X2=0.655 $Y2=1.765
cc_31 VPB N_A_c_75_n 0.028441f $X=-0.19 $Y=1.66 $X2=0.655 $Y2=1.765
cc_32 VPB N_A_c_77_n 0.00286496f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=1.365
cc_33 VPB N_B_c_104_n 0.0279325f $X=-0.19 $Y=1.66 $X2=0.655 $Y2=1.765
cc_34 VPB N_B_c_106_n 0.00246919f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=1.365
cc_35 VPB N_A_27_112#_c_137_n 0.0327793f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.21
cc_36 VPB N_A_27_112#_c_143_n 0.00168917f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_37 VPB N_A_27_112#_c_144_n 0.0217384f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_38 VPB N_A_27_112#_c_140_n 0.00811534f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_39 VPB N_A_27_112#_c_146_n 0.0328014f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_40 VPB N_A_27_112#_c_141_n 0.00241918f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_41 VPB N_VPWR_c_200_n 0.0171181f $X=-0.19 $Y=1.66 $X2=0.7 $Y2=0.835
cc_42 VPB N_VPWR_c_201_n 0.0265205f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=1.385
cc_43 VPB N_VPWR_c_202_n 0.00614127f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=1.385
cc_44 VPB N_VPWR_c_203_n 0.0525134f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_45 VPB N_VPWR_c_199_n 0.0879731f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_46 VPB N_Y_c_231_n 0.0385529f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_47 VPB N_Y_c_228_n 0.0308317f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_48 N_C_N_c_48_n N_A_c_75_n 0.0418823f $X=0.655 $Y=1.765 $X2=-0.19 $Y2=-0.245
cc_49 C_N N_A_c_75_n 0.00113494f $X=0.635 $Y=1.21 $X2=-0.19 $Y2=-0.245
cc_50 N_C_N_c_49_n N_A_M1007_g 0.014565f $X=0.7 $Y=1.22 $X2=0 $Y2=0
cc_51 C_N N_A_M1007_g 0.00343954f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_52 N_C_N_c_48_n N_A_c_77_n 0.00335781f $X=0.655 $Y=1.765 $X2=0 $Y2=0
cc_53 C_N N_A_c_77_n 0.0159708f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_54 N_C_N_c_48_n N_A_27_112#_c_148_n 0.014246f $X=0.655 $Y=1.765 $X2=0 $Y2=0
cc_55 C_N N_A_27_112#_c_148_n 0.00722565f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_56 N_C_N_c_48_n N_A_27_112#_c_139_n 0.00105773f $X=0.655 $Y=1.765 $X2=0 $Y2=0
cc_57 N_C_N_c_49_n N_A_27_112#_c_139_n 0.00429074f $X=0.7 $Y=1.22 $X2=0 $Y2=0
cc_58 C_N N_A_27_112#_c_139_n 0.014413f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_59 N_C_N_c_48_n N_A_27_112#_c_144_n 0.00721244f $X=0.655 $Y=1.765 $X2=0 $Y2=0
cc_60 C_N N_A_27_112#_c_144_n 0.00890472f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_61 N_C_N_c_48_n N_A_27_112#_c_140_n 0.0105299f $X=0.655 $Y=1.765 $X2=0 $Y2=0
cc_62 N_C_N_c_49_n N_A_27_112#_c_140_n 0.00459385f $X=0.7 $Y=1.22 $X2=0 $Y2=0
cc_63 C_N N_A_27_112#_c_140_n 0.0282012f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_64 N_C_N_c_48_n N_A_27_112#_c_146_n 0.0123352f $X=0.655 $Y=1.765 $X2=0 $Y2=0
cc_65 N_C_N_c_48_n N_VPWR_c_200_n 0.0068216f $X=0.655 $Y=1.765 $X2=0 $Y2=0
cc_66 N_C_N_c_48_n N_VPWR_c_201_n 0.00393873f $X=0.655 $Y=1.765 $X2=0 $Y2=0
cc_67 N_C_N_c_48_n N_VPWR_c_199_n 0.00462577f $X=0.655 $Y=1.765 $X2=0 $Y2=0
cc_68 N_C_N_c_49_n N_VGND_c_270_n 0.00619988f $X=0.7 $Y=1.22 $X2=0 $Y2=0
cc_69 N_C_N_c_49_n N_VGND_c_272_n 0.00434489f $X=0.7 $Y=1.22 $X2=0 $Y2=0
cc_70 N_C_N_c_49_n N_VGND_c_277_n 0.00487769f $X=0.7 $Y=1.22 $X2=0 $Y2=0
cc_71 N_A_c_75_n N_B_c_104_n 0.0856124f $X=1.225 $Y=1.765 $X2=-0.19 $Y2=-0.245
cc_72 N_A_c_77_n N_B_c_104_n 0.00154866f $X=1.15 $Y=1.515 $X2=-0.19 $Y2=-0.245
cc_73 N_A_M1007_g N_B_M1006_g 0.0165331f $X=1.24 $Y=0.74 $X2=0 $Y2=0
cc_74 N_A_c_75_n N_B_c_106_n 0.00154866f $X=1.225 $Y=1.765 $X2=0 $Y2=0
cc_75 N_A_c_77_n N_B_c_106_n 0.0246243f $X=1.15 $Y=1.515 $X2=0 $Y2=0
cc_76 N_A_c_75_n N_A_27_112#_c_148_n 0.0159168f $X=1.225 $Y=1.765 $X2=0 $Y2=0
cc_77 N_A_c_77_n N_A_27_112#_c_148_n 0.0226548f $X=1.15 $Y=1.515 $X2=0 $Y2=0
cc_78 N_A_c_75_n N_A_27_112#_c_144_n 0.00135095f $X=1.225 $Y=1.765 $X2=0 $Y2=0
cc_79 N_A_c_75_n N_VPWR_c_200_n 0.0170305f $X=1.225 $Y=1.765 $X2=0 $Y2=0
cc_80 N_A_c_75_n N_VPWR_c_203_n 0.00413917f $X=1.225 $Y=1.765 $X2=0 $Y2=0
cc_81 N_A_c_75_n N_VPWR_c_199_n 0.00817532f $X=1.225 $Y=1.765 $X2=0 $Y2=0
cc_82 N_A_M1007_g N_Y_c_225_n 4.78065e-19 $X=1.24 $Y=0.74 $X2=0 $Y2=0
cc_83 N_A_M1007_g N_Y_c_227_n 0.00233828f $X=1.24 $Y=0.74 $X2=0 $Y2=0
cc_84 N_A_c_75_n N_VGND_c_270_n 0.00104209f $X=1.225 $Y=1.765 $X2=0 $Y2=0
cc_85 N_A_M1007_g N_VGND_c_270_n 0.00395387f $X=1.24 $Y=0.74 $X2=0 $Y2=0
cc_86 N_A_c_77_n N_VGND_c_270_n 0.00718896f $X=1.15 $Y=1.515 $X2=0 $Y2=0
cc_87 N_A_M1007_g N_VGND_c_274_n 0.00461464f $X=1.24 $Y=0.74 $X2=0 $Y2=0
cc_88 N_A_M1007_g N_VGND_c_277_n 0.00912669f $X=1.24 $Y=0.74 $X2=0 $Y2=0
cc_89 N_B_c_104_n N_A_27_112#_c_137_n 0.058845f $X=1.645 $Y=1.765 $X2=0 $Y2=0
cc_90 N_B_c_106_n N_A_27_112#_c_137_n 0.00188012f $X=1.72 $Y=1.515 $X2=0 $Y2=0
cc_91 N_B_M1006_g N_A_27_112#_M1000_g 0.0260254f $X=1.71 $Y=0.74 $X2=0 $Y2=0
cc_92 N_B_c_104_n N_A_27_112#_c_148_n 0.0163414f $X=1.645 $Y=1.765 $X2=0 $Y2=0
cc_93 N_B_c_106_n N_A_27_112#_c_148_n 0.0226548f $X=1.72 $Y=1.515 $X2=0 $Y2=0
cc_94 N_B_c_104_n N_A_27_112#_c_143_n 0.00145222f $X=1.645 $Y=1.765 $X2=0 $Y2=0
cc_95 N_B_c_104_n N_A_27_112#_c_141_n 0.00121489f $X=1.645 $Y=1.765 $X2=0 $Y2=0
cc_96 N_B_c_106_n N_A_27_112#_c_141_n 0.0246767f $X=1.72 $Y=1.515 $X2=0 $Y2=0
cc_97 N_B_c_104_n N_VPWR_c_200_n 0.00385876f $X=1.645 $Y=1.765 $X2=0 $Y2=0
cc_98 N_B_c_104_n N_VPWR_c_203_n 0.00461464f $X=1.645 $Y=1.765 $X2=0 $Y2=0
cc_99 N_B_c_104_n N_VPWR_c_199_n 0.00910574f $X=1.645 $Y=1.765 $X2=0 $Y2=0
cc_100 N_B_M1006_g N_Y_c_225_n 0.00963749f $X=1.71 $Y=0.74 $X2=0 $Y2=0
cc_101 N_B_c_104_n N_Y_c_226_n 6.97898e-19 $X=1.645 $Y=1.765 $X2=0 $Y2=0
cc_102 N_B_M1006_g N_Y_c_226_n 0.0117933f $X=1.71 $Y=0.74 $X2=0 $Y2=0
cc_103 N_B_c_106_n N_Y_c_226_n 0.0167639f $X=1.72 $Y=1.515 $X2=0 $Y2=0
cc_104 N_B_c_104_n N_Y_c_227_n 6.18732e-19 $X=1.645 $Y=1.765 $X2=0 $Y2=0
cc_105 N_B_M1006_g N_Y_c_227_n 0.00153788f $X=1.71 $Y=0.74 $X2=0 $Y2=0
cc_106 N_B_c_106_n N_Y_c_227_n 0.00886294f $X=1.72 $Y=1.515 $X2=0 $Y2=0
cc_107 N_B_c_104_n N_Y_c_231_n 0.00308082f $X=1.645 $Y=1.765 $X2=0 $Y2=0
cc_108 N_B_M1006_g N_Y_c_229_n 6.27049e-19 $X=1.71 $Y=0.74 $X2=0 $Y2=0
cc_109 N_B_M1006_g N_VGND_c_271_n 0.00484409f $X=1.71 $Y=0.74 $X2=0 $Y2=0
cc_110 N_B_M1006_g N_VGND_c_274_n 0.00434272f $X=1.71 $Y=0.74 $X2=0 $Y2=0
cc_111 N_B_M1006_g N_VGND_c_277_n 0.0082177f $X=1.71 $Y=0.74 $X2=0 $Y2=0
cc_112 N_A_27_112#_c_148_n N_VPWR_M1001_d 0.0130612f $X=2.125 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_113 N_A_27_112#_c_148_n N_VPWR_c_200_n 0.0219335f $X=2.125 $Y=2.035 $X2=0
+ $Y2=0
cc_114 N_A_27_112#_c_146_n N_VPWR_c_200_n 0.025186f $X=0.35 $Y=2.035 $X2=0 $Y2=0
cc_115 N_A_27_112#_c_146_n N_VPWR_c_201_n 0.00995358f $X=0.35 $Y=2.035 $X2=0
+ $Y2=0
cc_116 N_A_27_112#_c_137_n N_VPWR_c_203_n 0.00445602f $X=2.215 $Y=1.765 $X2=0
+ $Y2=0
cc_117 N_A_27_112#_c_137_n N_VPWR_c_199_n 0.00863322f $X=2.215 $Y=1.765 $X2=0
+ $Y2=0
cc_118 N_A_27_112#_c_146_n N_VPWR_c_199_n 0.0148468f $X=0.35 $Y=2.035 $X2=0
+ $Y2=0
cc_119 N_A_27_112#_c_148_n A_260_368# 0.0119045f $X=2.125 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_120 N_A_27_112#_c_148_n A_344_368# 0.0207543f $X=2.125 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_121 N_A_27_112#_M1000_g N_Y_c_225_n 6.28869e-19 $X=2.28 $Y=0.74 $X2=0 $Y2=0
cc_122 N_A_27_112#_c_137_n N_Y_c_226_n 5.50399e-19 $X=2.215 $Y=1.765 $X2=0 $Y2=0
cc_123 N_A_27_112#_M1000_g N_Y_c_226_n 0.0117933f $X=2.28 $Y=0.74 $X2=0 $Y2=0
cc_124 N_A_27_112#_c_141_n N_Y_c_226_n 0.0156476f $X=2.29 $Y=1.515 $X2=0 $Y2=0
cc_125 N_A_27_112#_c_137_n N_Y_c_231_n 0.015735f $X=2.215 $Y=1.765 $X2=0 $Y2=0
cc_126 N_A_27_112#_c_148_n N_Y_c_231_n 0.00114401f $X=2.125 $Y=2.035 $X2=0 $Y2=0
cc_127 N_A_27_112#_c_141_n N_Y_c_231_n 0.00392504f $X=2.29 $Y=1.515 $X2=0 $Y2=0
cc_128 N_A_27_112#_c_137_n N_Y_c_228_n 0.0145585f $X=2.215 $Y=1.765 $X2=0 $Y2=0
cc_129 N_A_27_112#_M1000_g N_Y_c_228_n 0.00367585f $X=2.28 $Y=0.74 $X2=0 $Y2=0
cc_130 N_A_27_112#_c_143_n N_Y_c_228_n 0.00985212f $X=2.21 $Y=1.95 $X2=0 $Y2=0
cc_131 N_A_27_112#_c_141_n N_Y_c_228_n 0.0248017f $X=2.29 $Y=1.515 $X2=0 $Y2=0
cc_132 N_A_27_112#_M1000_g N_Y_c_229_n 0.0104715f $X=2.28 $Y=0.74 $X2=0 $Y2=0
cc_133 N_A_27_112#_c_137_n N_Y_c_230_n 7.83559e-19 $X=2.215 $Y=1.765 $X2=0 $Y2=0
cc_134 N_A_27_112#_M1000_g N_Y_c_230_n 0.002266f $X=2.28 $Y=0.74 $X2=0 $Y2=0
cc_135 N_A_27_112#_c_141_n N_Y_c_230_n 0.0103958f $X=2.29 $Y=1.515 $X2=0 $Y2=0
cc_136 N_A_27_112#_M1000_g N_VGND_c_271_n 0.00622602f $X=2.28 $Y=0.74 $X2=0
+ $Y2=0
cc_137 N_A_27_112#_c_139_n N_VGND_c_272_n 0.00858362f $X=0.485 $Y=0.845 $X2=0
+ $Y2=0
cc_138 N_A_27_112#_M1000_g N_VGND_c_276_n 0.00434272f $X=2.28 $Y=0.74 $X2=0
+ $Y2=0
cc_139 N_A_27_112#_M1000_g N_VGND_c_277_n 0.00825279f $X=2.28 $Y=0.74 $X2=0
+ $Y2=0
cc_140 N_A_27_112#_c_139_n N_VGND_c_277_n 0.0154187f $X=0.485 $Y=0.845 $X2=0
+ $Y2=0
cc_141 N_VPWR_c_203_n N_Y_c_231_n 0.0230883f $X=2.64 $Y=3.33 $X2=0 $Y2=0
cc_142 N_VPWR_c_199_n N_Y_c_231_n 0.0190704f $X=2.64 $Y=3.33 $X2=0 $Y2=0
cc_143 N_Y_c_226_n N_VGND_M1006_d 0.00358162f $X=2.33 $Y=1.095 $X2=0 $Y2=0
cc_144 N_Y_c_225_n N_VGND_c_270_n 0.00158095f $X=1.495 $Y=0.515 $X2=0 $Y2=0
cc_145 N_Y_c_225_n N_VGND_c_271_n 0.0191765f $X=1.495 $Y=0.515 $X2=0 $Y2=0
cc_146 N_Y_c_226_n N_VGND_c_271_n 0.0248957f $X=2.33 $Y=1.095 $X2=0 $Y2=0
cc_147 N_Y_c_229_n N_VGND_c_271_n 0.0201667f $X=2.495 $Y=0.515 $X2=0 $Y2=0
cc_148 N_Y_c_225_n N_VGND_c_274_n 0.0145639f $X=1.495 $Y=0.515 $X2=0 $Y2=0
cc_149 N_Y_c_229_n N_VGND_c_276_n 0.0205877f $X=2.495 $Y=0.515 $X2=0 $Y2=0
cc_150 N_Y_c_225_n N_VGND_c_277_n 0.0119984f $X=1.495 $Y=0.515 $X2=0 $Y2=0
cc_151 N_Y_c_229_n N_VGND_c_277_n 0.0169844f $X=2.495 $Y=0.515 $X2=0 $Y2=0
