* File: sky130_fd_sc_hs__a222o_2.spice
* Created: Tue Sep  1 19:50:48 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hs__a222o_2.pex.spice"
.subckt sky130_fd_sc_hs__a222o_2  VNB VPB C1 C2 A1 B1 B2 A2 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A2	A2
* B2	B2
* B1	B1
* A1	A1
* C2	C2
* C1	C1
* VPB	VPB
* VNB	VNB
MM1002 A_114_82# N_C1_M1002_g N_A_27_82#_M1002_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.0768 AS=0.1824 PD=0.88 PS=1.85 NRD=12.18 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75001.8 A=0.096 P=1.58 MULT=1
MM1015 N_VGND_M1015_d N_C2_M1015_g A_114_82# VNB NLOWVT L=0.15 W=0.64
+ AD=0.192649 AS=0.0768 PD=1.25217 PS=0.88 NRD=0 NRS=12.18 M=1 R=4.26667
+ SA=75000.6 SB=75001.4 A=0.096 P=1.58 MULT=1
MM1004 N_X_M1004_d N_A_27_82#_M1004_g N_VGND_M1015_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.222751 PD=1.02 PS=1.44783 NRD=0 NRS=53.508 M=1 R=4.93333
+ SA=75001.2 SB=75000.6 A=0.111 P=1.78 MULT=1
MM1010 N_X_M1004_d N_A_27_82#_M1010_g N_VGND_M1010_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.2586 PD=1.02 PS=2.67 NRD=0 NRS=47.748 M=1 R=4.93333 SA=75001.6
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1008 N_A_27_82#_M1008_d N_A1_M1008_g N_A_557_74#_M1008_s VNB NLOWVT L=0.15
+ W=0.64 AD=0.1504 AS=0.1971 PD=1.11 PS=1.92 NRD=20.616 NRS=6.552 M=1 R=4.26667
+ SA=75000.2 SB=75001.8 A=0.096 P=1.58 MULT=1
MM1011 A_775_74# N_B1_M1011_g N_A_27_82#_M1008_d VNB NLOWVT L=0.15 W=0.64
+ AD=0.0768 AS=0.1504 PD=0.88 PS=1.11 NRD=12.18 NRS=14.988 M=1 R=4.26667
+ SA=75000.9 SB=75001.2 A=0.096 P=1.58 MULT=1
MM1012 N_VGND_M1012_d N_B2_M1012_g A_775_74# VNB NLOWVT L=0.15 W=0.64 AD=0.1344
+ AS=0.0768 PD=1.06 PS=0.88 NRD=3.744 NRS=12.18 M=1 R=4.26667 SA=75001.2
+ SB=75000.8 A=0.096 P=1.58 MULT=1
MM1000 N_A_557_74#_M1000_d N_A2_M1000_g N_VGND_M1012_d VNB NLOWVT L=0.15 W=0.64
+ AD=0.1824 AS=0.1344 PD=1.85 PS=1.06 NRD=0 NRS=22.488 M=1 R=4.26667 SA=75001.8
+ SB=75000.2 A=0.096 P=1.58 MULT=1
MM1006 N_A_116_392#_M1006_d N_C1_M1006_g N_A_27_82#_M1006_s VPB PSHORT L=0.15
+ W=1 AD=0.15 AS=0.295 PD=1.3 PS=2.59 NRD=1.9503 NRS=1.9503 M=1 R=6.66667
+ SA=75000.2 SB=75000.7 A=0.15 P=2.3 MULT=1
MM1007 N_A_27_82#_M1007_d N_C2_M1007_g N_A_116_392#_M1006_d VPB PSHORT L=0.15
+ W=1 AD=0.295 AS=0.15 PD=2.59 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=6.66667
+ SA=75000.7 SB=75000.2 A=0.15 P=2.3 MULT=1
MM1013 N_X_M1013_d N_A_27_82#_M1013_g N_VPWR_M1013_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.34065 PD=1.42 PS=3.12 NRD=1.7533 NRS=17.5724 M=1 R=7.46667
+ SA=75000.2 SB=75002.7 A=0.168 P=2.54 MULT=1
MM1014 N_X_M1013_d N_A_27_82#_M1014_g N_VPWR_M1014_s VPB PSHORT L=0.15 W=1.12
+ AD=0.168 AS=0.281585 PD=1.42 PS=1.7434 NRD=1.7533 NRS=17.5724 M=1 R=7.46667
+ SA=75000.7 SB=75002.3 A=0.168 P=2.54 MULT=1
MM1009 N_A_639_368#_M1009_d N_A1_M1009_g N_VPWR_M1014_s VPB PSHORT L=0.15 W=1
+ AD=0.28175 AS=0.251415 PD=1.685 PS=1.5566 NRD=22.655 NRS=19.6803 M=1 R=6.66667
+ SA=75001.3 SB=75001.9 A=0.15 P=2.3 MULT=1
MM1003 N_A_116_392#_M1003_d N_B1_M1003_g N_A_639_368#_M1009_d VPB PSHORT L=0.15
+ W=1 AD=0.15 AS=0.28175 PD=1.3 PS=1.685 NRD=0 NRS=44.6599 M=1 R=6.66667
+ SA=75001.9 SB=75001.2 A=0.15 P=2.3 MULT=1
MM1005 N_A_639_368#_M1005_d N_B2_M1005_g N_A_116_392#_M1003_d VPB PSHORT L=0.15
+ W=1 AD=0.2 AS=0.15 PD=1.4 PS=1.3 NRD=11.8003 NRS=1.9503 M=1 R=6.66667
+ SA=75002.4 SB=75000.8 A=0.15 P=2.3 MULT=1
MM1001 N_VPWR_M1001_d N_A2_M1001_g N_A_639_368#_M1005_d VPB PSHORT L=0.15 W=1
+ AD=0.295 AS=0.2 PD=2.59 PS=1.4 NRD=1.9503 NRS=11.8003 M=1 R=6.66667 SA=75002.9
+ SB=75000.2 A=0.15 P=2.3 MULT=1
DX16_noxref VNB VPB NWDIODE A=10.5276 P=15.04
c_655 A_775_74# 0 2.49076e-20 $X=3.875 $Y=0.37
*
.include "sky130_fd_sc_hs__a222o_2.pxi.spice"
*
.ends
*
*
