* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hs__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
M1000 Y A2 a_162_368# VPB pshort w=1.12e+06u l=150000u
+  ad=5.656e+11p pd=3.25e+06u as=3.024e+11p ps=2.78e+06u
M1001 a_27_74# A2 VGND VNB nlowvt w=740000u l=150000u
+  ad=4.181e+11p pd=4.09e+06u as=6.722e+11p ps=3.36e+06u
M1002 VPWR B1 Y VPB pshort w=1.12e+06u l=150000u
+  ad=7.952e+11p pd=5.9e+06u as=0p ps=0u
M1003 Y B1 a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=2.627e+11p pd=2.19e+06u as=0p ps=0u
M1004 VGND A1 a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_162_368# A1 VPWR VPB pshort w=1.12e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
