* File: sky130_fd_sc_hs__a211oi_4.pex.spice
* Created: Tue Sep  1 19:48:53 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HS__A211OI_4%A2 1 3 6 8 10 13 15 17 20 22 24 27 29 30 31
+ 32 33 51
c81 33 0 9.93954e-20 $X=2.16 $Y=1.665
c82 27 0 2.04552e-19 $X=2.09 $Y=0.74
c83 22 0 1.30641e-20 $X=2.085 $Y=1.765
r84 51 52 0.651351 $w=3.7e-07 $l=5e-09 $layer=POLY_cond $X=2.085 $Y=1.557
+ $X2=2.09 $Y2=1.557
r85 49 51 33.2189 $w=3.7e-07 $l=2.55e-07 $layer=POLY_cond $X=1.83 $Y=1.557
+ $X2=2.085 $Y2=1.557
r86 49 50 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.83
+ $Y=1.515 $X2=1.83 $Y2=1.515
r87 47 49 22.1459 $w=3.7e-07 $l=1.7e-07 $layer=POLY_cond $X=1.66 $Y=1.557
+ $X2=1.83 $Y2=1.557
r88 46 47 3.25676 $w=3.7e-07 $l=2.5e-08 $layer=POLY_cond $X=1.635 $Y=1.557
+ $X2=1.66 $Y2=1.557
r89 45 46 52.7595 $w=3.7e-07 $l=4.05e-07 $layer=POLY_cond $X=1.23 $Y=1.557
+ $X2=1.635 $Y2=1.557
r90 44 45 5.86216 $w=3.7e-07 $l=4.5e-08 $layer=POLY_cond $X=1.185 $Y=1.557
+ $X2=1.23 $Y2=1.557
r91 42 44 48.8514 $w=3.7e-07 $l=3.75e-07 $layer=POLY_cond $X=0.81 $Y=1.557
+ $X2=1.185 $Y2=1.557
r92 42 43 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.81
+ $Y=1.515 $X2=0.81 $Y2=1.515
r93 40 42 1.3027 $w=3.7e-07 $l=1e-08 $layer=POLY_cond $X=0.8 $Y=1.557 $X2=0.81
+ $Y2=1.557
r94 39 40 8.46757 $w=3.7e-07 $l=6.5e-08 $layer=POLY_cond $X=0.735 $Y=1.557
+ $X2=0.8 $Y2=1.557
r95 33 50 8.84433 $w=4.28e-07 $l=3.3e-07 $layer=LI1_cond $X=2.16 $Y=1.565
+ $X2=1.83 $Y2=1.565
r96 32 50 4.02015 $w=4.28e-07 $l=1.5e-07 $layer=LI1_cond $X=1.68 $Y=1.565
+ $X2=1.83 $Y2=1.565
r97 31 32 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=1.2 $Y=1.565
+ $X2=1.68 $Y2=1.565
r98 31 43 10.4524 $w=4.28e-07 $l=3.9e-07 $layer=LI1_cond $X=1.2 $Y=1.565
+ $X2=0.81 $Y2=1.565
r99 30 43 2.41209 $w=4.28e-07 $l=9e-08 $layer=LI1_cond $X=0.72 $Y=1.565 $X2=0.81
+ $Y2=1.565
r100 29 30 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=0.24 $Y=1.565
+ $X2=0.72 $Y2=1.565
r101 25 52 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.09 $Y=1.35
+ $X2=2.09 $Y2=1.557
r102 25 27 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.09 $Y=1.35
+ $X2=2.09 $Y2=0.74
r103 22 51 23.9667 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=2.085 $Y=1.765
+ $X2=2.085 $Y2=1.557
r104 22 24 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.085 $Y=1.765
+ $X2=2.085 $Y2=2.4
r105 18 47 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.66 $Y=1.35
+ $X2=1.66 $Y2=1.557
r106 18 20 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.66 $Y=1.35
+ $X2=1.66 $Y2=0.74
r107 15 46 23.9667 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=1.635 $Y=1.765
+ $X2=1.635 $Y2=1.557
r108 15 17 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.635 $Y=1.765
+ $X2=1.635 $Y2=2.4
r109 11 45 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.23 $Y=1.35
+ $X2=1.23 $Y2=1.557
r110 11 13 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.23 $Y=1.35
+ $X2=1.23 $Y2=0.74
r111 8 44 23.9667 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=1.185 $Y=1.765
+ $X2=1.185 $Y2=1.557
r112 8 10 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.185 $Y=1.765
+ $X2=1.185 $Y2=2.4
r113 4 40 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.8 $Y=1.35 $X2=0.8
+ $Y2=1.557
r114 4 6 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=0.8 $Y=1.35 $X2=0.8
+ $Y2=0.74
r115 1 39 23.9667 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=0.735 $Y=1.765
+ $X2=0.735 $Y2=1.557
r116 1 3 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.735 $Y=1.765
+ $X2=0.735 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_HS__A211OI_4%A1 3 5 7 10 12 14 17 19 21 24 26 28 29 30
+ 31 46 47
c74 46 0 1.30641e-20 $X=3.69 $Y=1.515
c75 5 0 9.93954e-20 $X=2.535 $Y=1.765
r76 47 48 9.77027 $w=3.7e-07 $l=7.5e-08 $layer=POLY_cond $X=3.81 $Y=1.557
+ $X2=3.885 $Y2=1.557
r77 45 47 15.6324 $w=3.7e-07 $l=1.2e-07 $layer=POLY_cond $X=3.69 $Y=1.557
+ $X2=3.81 $Y2=1.557
r78 45 46 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.69
+ $Y=1.515 $X2=3.69 $Y2=1.515
r79 43 45 33.2189 $w=3.7e-07 $l=2.55e-07 $layer=POLY_cond $X=3.435 $Y=1.557
+ $X2=3.69 $Y2=1.557
r80 42 43 7.16487 $w=3.7e-07 $l=5.5e-08 $layer=POLY_cond $X=3.38 $Y=1.557
+ $X2=3.435 $Y2=1.557
r81 41 42 51.4568 $w=3.7e-07 $l=3.95e-07 $layer=POLY_cond $X=2.985 $Y=1.557
+ $X2=3.38 $Y2=1.557
r82 40 41 4.55946 $w=3.7e-07 $l=3.5e-08 $layer=POLY_cond $X=2.95 $Y=1.557
+ $X2=2.985 $Y2=1.557
r83 38 40 36.4757 $w=3.7e-07 $l=2.8e-07 $layer=POLY_cond $X=2.67 $Y=1.557
+ $X2=2.95 $Y2=1.557
r84 38 39 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.67
+ $Y=1.515 $X2=2.67 $Y2=1.515
r85 36 38 17.5865 $w=3.7e-07 $l=1.35e-07 $layer=POLY_cond $X=2.535 $Y=1.557
+ $X2=2.67 $Y2=1.557
r86 35 36 1.95405 $w=3.7e-07 $l=1.5e-08 $layer=POLY_cond $X=2.52 $Y=1.557
+ $X2=2.535 $Y2=1.557
r87 31 46 2.41209 $w=4.28e-07 $l=9e-08 $layer=LI1_cond $X=3.6 $Y=1.565 $X2=3.69
+ $Y2=1.565
r88 30 31 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=3.12 $Y=1.565
+ $X2=3.6 $Y2=1.565
r89 30 39 12.0604 $w=4.28e-07 $l=4.5e-07 $layer=LI1_cond $X=3.12 $Y=1.565
+ $X2=2.67 $Y2=1.565
r90 29 39 0.80403 $w=4.28e-07 $l=3e-08 $layer=LI1_cond $X=2.64 $Y=1.565 $X2=2.67
+ $Y2=1.565
r91 26 48 23.9667 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=3.885 $Y=1.765
+ $X2=3.885 $Y2=1.557
r92 26 28 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.885 $Y=1.765
+ $X2=3.885 $Y2=2.4
r93 22 47 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.81 $Y=1.35
+ $X2=3.81 $Y2=1.557
r94 22 24 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=3.81 $Y=1.35
+ $X2=3.81 $Y2=0.74
r95 19 43 23.9667 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=3.435 $Y=1.765
+ $X2=3.435 $Y2=1.557
r96 19 21 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=3.435 $Y=1.765
+ $X2=3.435 $Y2=2.4
r97 15 42 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.38 $Y=1.35
+ $X2=3.38 $Y2=1.557
r98 15 17 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=3.38 $Y=1.35
+ $X2=3.38 $Y2=0.74
r99 12 41 23.9667 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=2.985 $Y=1.765
+ $X2=2.985 $Y2=1.557
r100 12 14 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.985 $Y=1.765
+ $X2=2.985 $Y2=2.4
r101 8 40 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.95 $Y=1.35
+ $X2=2.95 $Y2=1.557
r102 8 10 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.95 $Y=1.35
+ $X2=2.95 $Y2=0.74
r103 5 36 23.9667 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=2.535 $Y=1.765
+ $X2=2.535 $Y2=1.557
r104 5 7 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.535 $Y=1.765
+ $X2=2.535 $Y2=2.4
r105 1 35 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.52 $Y=1.35
+ $X2=2.52 $Y2=1.557
r106 1 3 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.52 $Y=1.35 $X2=2.52
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HS__A211OI_4%B1 1 3 4 6 7 9 12 16 18 20 21 22 23 24 39
c77 39 0 1.7359e-19 $X=6.19 $Y=1.532
c78 18 0 1.26549e-19 $X=6.205 $Y=1.765
r79 39 40 1.83969 $w=3.93e-07 $l=1.5e-08 $layer=POLY_cond $X=6.19 $Y=1.532
+ $X2=6.205 $Y2=1.532
r80 37 39 29.4351 $w=3.93e-07 $l=2.4e-07 $layer=POLY_cond $X=5.95 $Y=1.532
+ $X2=6.19 $Y2=1.532
r81 37 38 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.95
+ $Y=1.465 $X2=5.95 $Y2=1.465
r82 35 37 23.3028 $w=3.93e-07 $l=1.9e-07 $layer=POLY_cond $X=5.76 $Y=1.532
+ $X2=5.95 $Y2=1.532
r83 34 35 0.613232 $w=3.93e-07 $l=5e-09 $layer=POLY_cond $X=5.755 $Y=1.532
+ $X2=5.76 $Y2=1.532
r84 33 34 55.1908 $w=3.93e-07 $l=4.5e-07 $layer=POLY_cond $X=5.305 $Y=1.532
+ $X2=5.755 $Y2=1.532
r85 31 33 45.9924 $w=3.93e-07 $l=3.75e-07 $layer=POLY_cond $X=4.93 $Y=1.532
+ $X2=5.305 $Y2=1.532
r86 31 32 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.93
+ $Y=1.465 $X2=4.93 $Y2=1.465
r87 29 31 9.19847 $w=3.93e-07 $l=7.5e-08 $layer=POLY_cond $X=4.855 $Y=1.532
+ $X2=4.93 $Y2=1.532
r88 24 38 1.24592 $w=4.78e-07 $l=5e-08 $layer=LI1_cond $X=6 $Y=1.54 $X2=5.95
+ $Y2=1.54
r89 23 38 10.7149 $w=4.78e-07 $l=4.3e-07 $layer=LI1_cond $X=5.52 $Y=1.54
+ $X2=5.95 $Y2=1.54
r90 22 23 11.9608 $w=4.78e-07 $l=4.8e-07 $layer=LI1_cond $X=5.04 $Y=1.54
+ $X2=5.52 $Y2=1.54
r91 22 32 2.74101 $w=4.78e-07 $l=1.1e-07 $layer=LI1_cond $X=5.04 $Y=1.54
+ $X2=4.93 $Y2=1.54
r92 21 32 9.21977 $w=4.78e-07 $l=3.7e-07 $layer=LI1_cond $X=4.56 $Y=1.54
+ $X2=4.93 $Y2=1.54
r93 18 40 25.4309 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=6.205 $Y=1.765
+ $X2=6.205 $Y2=1.532
r94 18 20 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=6.205 $Y=1.765
+ $X2=6.205 $Y2=2.4
r95 14 39 25.4309 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=6.19 $Y=1.3
+ $X2=6.19 $Y2=1.532
r96 14 16 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=6.19 $Y=1.3 $X2=6.19
+ $Y2=0.74
r97 10 35 25.4309 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=5.76 $Y=1.3
+ $X2=5.76 $Y2=1.532
r98 10 12 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=5.76 $Y=1.3 $X2=5.76
+ $Y2=0.74
r99 7 34 25.4309 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=5.755 $Y=1.765
+ $X2=5.755 $Y2=1.532
r100 7 9 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=5.755 $Y=1.765
+ $X2=5.755 $Y2=2.4
r101 4 33 25.4309 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=5.305 $Y=1.765
+ $X2=5.305 $Y2=1.532
r102 4 6 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=5.305 $Y=1.765
+ $X2=5.305 $Y2=2.4
r103 1 29 25.4309 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=4.855 $Y=1.765
+ $X2=4.855 $Y2=1.532
r104 1 3 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=4.855 $Y=1.765
+ $X2=4.855 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_HS__A211OI_4%C1 3 5 7 10 12 14 15 17 18 20 21 22 23 37
c64 23 0 1.26549e-19 $X=7.44 $Y=1.665
r65 37 38 54.3609 $w=3.99e-07 $l=4.5e-07 $layer=POLY_cond $X=7.555 $Y=1.542
+ $X2=8.005 $Y2=1.542
r66 35 37 19.9323 $w=3.99e-07 $l=1.65e-07 $layer=POLY_cond $X=7.39 $Y=1.542
+ $X2=7.555 $Y2=1.542
r67 35 36 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=7.39
+ $Y=1.515 $X2=7.39 $Y2=1.515
r68 33 35 34.4286 $w=3.99e-07 $l=2.85e-07 $layer=POLY_cond $X=7.105 $Y=1.542
+ $X2=7.39 $Y2=1.542
r69 32 33 6.64411 $w=3.99e-07 $l=5.5e-08 $layer=POLY_cond $X=7.05 $Y=1.542
+ $X2=7.105 $Y2=1.542
r70 30 32 41.0727 $w=3.99e-07 $l=3.4e-07 $layer=POLY_cond $X=6.71 $Y=1.542
+ $X2=7.05 $Y2=1.542
r71 30 31 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=6.71
+ $Y=1.515 $X2=6.71 $Y2=1.515
r72 28 30 6.64411 $w=3.99e-07 $l=5.5e-08 $layer=POLY_cond $X=6.655 $Y=1.542
+ $X2=6.71 $Y2=1.542
r73 27 28 4.22807 $w=3.99e-07 $l=3.5e-08 $layer=POLY_cond $X=6.62 $Y=1.542
+ $X2=6.655 $Y2=1.542
r74 23 36 1.34005 $w=4.28e-07 $l=5e-08 $layer=LI1_cond $X=7.44 $Y=1.565 $X2=7.39
+ $Y2=1.565
r75 22 36 11.5244 $w=4.28e-07 $l=4.3e-07 $layer=LI1_cond $X=6.96 $Y=1.565
+ $X2=7.39 $Y2=1.565
r76 22 31 6.70025 $w=4.28e-07 $l=2.5e-07 $layer=LI1_cond $X=6.96 $Y=1.565
+ $X2=6.71 $Y2=1.565
r77 21 31 6.16423 $w=4.28e-07 $l=2.3e-07 $layer=LI1_cond $X=6.48 $Y=1.565
+ $X2=6.71 $Y2=1.565
r78 18 38 25.8008 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=8.005 $Y=1.765
+ $X2=8.005 $Y2=1.542
r79 18 20 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=8.005 $Y=1.765
+ $X2=8.005 $Y2=2.4
r80 15 37 25.8008 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=7.555 $Y=1.765
+ $X2=7.555 $Y2=1.542
r81 15 17 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=7.555 $Y=1.765
+ $X2=7.555 $Y2=2.4
r82 12 33 25.8008 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=7.105 $Y=1.765
+ $X2=7.105 $Y2=1.542
r83 12 14 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=7.105 $Y=1.765
+ $X2=7.105 $Y2=2.4
r84 8 32 25.8008 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=7.05 $Y=1.32
+ $X2=7.05 $Y2=1.542
r85 8 10 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=7.05 $Y=1.32 $X2=7.05
+ $Y2=0.74
r86 5 28 25.8008 $w=1.5e-07 $l=2.23e-07 $layer=POLY_cond $X=6.655 $Y=1.765
+ $X2=6.655 $Y2=1.542
r87 5 7 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=6.655 $Y=1.765
+ $X2=6.655 $Y2=2.4
r88 1 27 25.8008 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=6.62 $Y=1.32
+ $X2=6.62 $Y2=1.542
r89 1 3 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=6.62 $Y=1.32 $X2=6.62
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HS__A211OI_4%A_77_368# 1 2 3 4 5 6 7 22 24 26 30 32 36
+ 38 42 44 48 50 54 56 58 60 65 67 69 71 73
c99 50 0 1.7359e-19 $X=4.995 $Y=2.035
r100 58 75 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.02 $Y=2.12
+ $X2=6.02 $Y2=2.035
r101 58 60 20.744 $w=2.48e-07 $l=4.5e-07 $layer=LI1_cond $X=6.02 $Y=2.12
+ $X2=6.02 $Y2=2.57
r102 57 73 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.165 $Y=2.035
+ $X2=5.08 $Y2=2.035
r103 56 75 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.895 $Y=2.035
+ $X2=6.02 $Y2=2.035
r104 56 57 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=5.895 $Y=2.035
+ $X2=5.165 $Y2=2.035
r105 52 73 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.08 $Y=2.12
+ $X2=5.08 $Y2=2.035
r106 52 54 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=5.08 $Y=2.12
+ $X2=5.08 $Y2=2.57
r107 51 71 7.02821 $w=1.7e-07 $l=1.5411e-07 $layer=LI1_cond $X=4.275 $Y=2.035
+ $X2=4.15 $Y2=1.97
r108 50 73 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.995 $Y=2.035
+ $X2=5.08 $Y2=2.035
r109 50 51 46.9733 $w=1.68e-07 $l=7.2e-07 $layer=LI1_cond $X=4.995 $Y=2.035
+ $X2=4.275 $Y2=2.035
r110 46 71 0.00168595 $w=2.5e-07 $l=1.5e-07 $layer=LI1_cond $X=4.15 $Y=2.12
+ $X2=4.15 $Y2=1.97
r111 46 48 12.9074 $w=2.48e-07 $l=2.8e-07 $layer=LI1_cond $X=4.15 $Y=2.12
+ $X2=4.15 $Y2=2.4
r112 45 69 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.295 $Y=2.035
+ $X2=3.21 $Y2=2.035
r113 44 71 7.02821 $w=1.7e-07 $l=1.5411e-07 $layer=LI1_cond $X=4.025 $Y=2.035
+ $X2=4.15 $Y2=1.97
r114 44 45 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=4.025 $Y=2.035
+ $X2=3.295 $Y2=2.035
r115 40 69 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.21 $Y=2.12
+ $X2=3.21 $Y2=2.035
r116 40 42 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=3.21 $Y=2.12
+ $X2=3.21 $Y2=2.445
r117 39 67 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.395 $Y=2.035
+ $X2=2.31 $Y2=2.035
r118 38 69 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.125 $Y=2.035
+ $X2=3.21 $Y2=2.035
r119 38 39 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=3.125 $Y=2.035
+ $X2=2.395 $Y2=2.035
r120 34 67 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.31 $Y=2.12
+ $X2=2.31 $Y2=2.035
r121 34 36 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=2.31 $Y=2.12
+ $X2=2.31 $Y2=2.445
r122 33 65 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.495 $Y=2.035
+ $X2=1.37 $Y2=2.035
r123 32 67 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.225 $Y=2.035
+ $X2=2.31 $Y2=2.035
r124 32 33 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=2.225 $Y=2.035
+ $X2=1.495 $Y2=2.035
r125 28 65 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.37 $Y=2.12
+ $X2=1.37 $Y2=2.035
r126 28 30 14.9818 $w=2.48e-07 $l=3.25e-07 $layer=LI1_cond $X=1.37 $Y=2.12
+ $X2=1.37 $Y2=2.445
r127 27 63 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.675 $Y=2.035
+ $X2=0.51 $Y2=2.035
r128 26 65 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.245 $Y=2.035
+ $X2=1.37 $Y2=2.035
r129 26 27 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=1.245 $Y=2.035
+ $X2=0.675 $Y2=2.035
r130 22 63 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.51 $Y=2.12 $X2=0.51
+ $Y2=2.035
r131 22 24 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=0.51 $Y=2.12
+ $X2=0.51 $Y2=2.815
r132 7 75 600 $w=1.7e-07 $l=2.59374e-07 $layer=licon1_PDIFF $count=1 $X=5.83
+ $Y=1.84 $X2=5.98 $Y2=2.035
r133 7 60 600 $w=1.7e-07 $l=8.01499e-07 $layer=licon1_PDIFF $count=1 $X=5.83
+ $Y=1.84 $X2=5.98 $Y2=2.57
r134 6 73 600 $w=1.7e-07 $l=2.59374e-07 $layer=licon1_PDIFF $count=1 $X=4.93
+ $Y=1.84 $X2=5.08 $Y2=2.035
r135 6 54 600 $w=1.7e-07 $l=8.01499e-07 $layer=licon1_PDIFF $count=1 $X=4.93
+ $Y=1.84 $X2=5.08 $Y2=2.57
r136 5 71 600 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=3.96
+ $Y=1.84 $X2=4.11 $Y2=1.985
r137 5 48 300 $w=1.7e-07 $l=6.30555e-07 $layer=licon1_PDIFF $count=2 $X=3.96
+ $Y=1.84 $X2=4.11 $Y2=2.4
r138 4 69 600 $w=1.7e-07 $l=2.59374e-07 $layer=licon1_PDIFF $count=1 $X=3.06
+ $Y=1.84 $X2=3.21 $Y2=2.035
r139 4 42 300 $w=1.7e-07 $l=6.75851e-07 $layer=licon1_PDIFF $count=2 $X=3.06
+ $Y=1.84 $X2=3.21 $Y2=2.445
r140 3 67 600 $w=1.7e-07 $l=2.59374e-07 $layer=licon1_PDIFF $count=1 $X=2.16
+ $Y=1.84 $X2=2.31 $Y2=2.035
r141 3 36 300 $w=1.7e-07 $l=6.75851e-07 $layer=licon1_PDIFF $count=2 $X=2.16
+ $Y=1.84 $X2=2.31 $Y2=2.445
r142 2 65 600 $w=1.7e-07 $l=2.59374e-07 $layer=licon1_PDIFF $count=1 $X=1.26
+ $Y=1.84 $X2=1.41 $Y2=2.035
r143 2 30 300 $w=1.7e-07 $l=6.75851e-07 $layer=licon1_PDIFF $count=2 $X=1.26
+ $Y=1.84 $X2=1.41 $Y2=2.445
r144 1 63 400 $w=1.7e-07 $l=2.498e-07 $layer=licon1_PDIFF $count=1 $X=0.385
+ $Y=1.84 $X2=0.51 $Y2=2.035
r145 1 24 400 $w=1.7e-07 $l=1.03562e-06 $layer=licon1_PDIFF $count=1 $X=0.385
+ $Y=1.84 $X2=0.51 $Y2=2.815
.ends

.subckt PM_SKY130_FD_SC_HS__A211OI_4%VPWR 1 2 3 4 15 19 21 25 29 32 33 34 35 36
+ 45 55 56 59 62
r103 62 63 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r104 59 60 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r105 55 56 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=8.4 $Y=3.33
+ $X2=8.4 $Y2=3.33
r106 53 63 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=3.6 $Y2=3.33
r107 52 55 281.84 $w=1.68e-07 $l=4.32e-06 $layer=LI1_cond $X=4.08 $Y=3.33
+ $X2=8.4 $Y2=3.33
r108 52 53 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r109 50 62 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.825 $Y=3.33
+ $X2=3.66 $Y2=3.33
r110 50 52 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=3.825 $Y=3.33
+ $X2=4.08 $Y2=3.33
r111 49 63 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=3.6 $Y2=3.33
r112 49 60 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=2.64 $Y2=3.33
r113 48 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r114 46 59 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.925 $Y=3.33
+ $X2=2.76 $Y2=3.33
r115 46 48 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=2.925 $Y=3.33
+ $X2=3.12 $Y2=3.33
r116 45 62 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.495 $Y=3.33
+ $X2=3.66 $Y2=3.33
r117 45 48 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=3.495 $Y=3.33
+ $X2=3.12 $Y2=3.33
r118 44 60 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.64 $Y2=3.33
r119 43 44 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r120 40 44 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.68 $Y2=3.33
r121 39 40 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r122 36 56 1.13724 $w=4.9e-07 $l=4.08e-06 $layer=MET1_cond $X=4.32 $Y=3.33
+ $X2=8.4 $Y2=3.33
r123 36 53 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=4.32 $Y=3.33
+ $X2=4.08 $Y2=3.33
r124 34 43 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=1.695 $Y=3.33
+ $X2=1.68 $Y2=3.33
r125 34 35 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.695 $Y=3.33
+ $X2=1.86 $Y2=3.33
r126 32 39 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=0.875 $Y=3.33
+ $X2=0.72 $Y2=3.33
r127 32 33 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.875 $Y=3.33
+ $X2=0.96 $Y2=3.33
r128 31 43 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=1.045 $Y=3.33
+ $X2=1.68 $Y2=3.33
r129 31 33 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.045 $Y=3.33
+ $X2=0.96 $Y2=3.33
r130 27 62 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.66 $Y=3.245
+ $X2=3.66 $Y2=3.33
r131 27 29 29.1603 $w=3.28e-07 $l=8.35e-07 $layer=LI1_cond $X=3.66 $Y=3.245
+ $X2=3.66 $Y2=2.41
r132 23 59 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.76 $Y=3.245
+ $X2=2.76 $Y2=3.33
r133 23 25 29.1603 $w=3.28e-07 $l=8.35e-07 $layer=LI1_cond $X=2.76 $Y=3.245
+ $X2=2.76 $Y2=2.41
r134 22 35 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.025 $Y=3.33
+ $X2=1.86 $Y2=3.33
r135 21 59 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.595 $Y=3.33
+ $X2=2.76 $Y2=3.33
r136 21 22 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=2.595 $Y=3.33
+ $X2=2.025 $Y2=3.33
r137 17 35 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.86 $Y=3.245
+ $X2=1.86 $Y2=3.33
r138 17 19 29.1603 $w=3.28e-07 $l=8.35e-07 $layer=LI1_cond $X=1.86 $Y=3.245
+ $X2=1.86 $Y2=2.41
r139 13 33 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.96 $Y=3.245
+ $X2=0.96 $Y2=3.33
r140 13 15 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=0.96 $Y=3.245
+ $X2=0.96 $Y2=2.455
r141 4 29 300 $w=1.7e-07 $l=6.40625e-07 $layer=licon1_PDIFF $count=2 $X=3.51
+ $Y=1.84 $X2=3.66 $Y2=2.41
r142 3 25 300 $w=1.7e-07 $l=6.40625e-07 $layer=licon1_PDIFF $count=2 $X=2.61
+ $Y=1.84 $X2=2.76 $Y2=2.41
r143 2 19 300 $w=1.7e-07 $l=6.40625e-07 $layer=licon1_PDIFF $count=2 $X=1.71
+ $Y=1.84 $X2=1.86 $Y2=2.41
r144 1 15 300 $w=1.7e-07 $l=6.85912e-07 $layer=licon1_PDIFF $count=2 $X=0.81
+ $Y=1.84 $X2=0.96 $Y2=2.455
.ends

.subckt PM_SKY130_FD_SC_HS__A211OI_4%A_901_368# 1 2 3 4 5 18 20 21 24 26 30 34
+ 38 40 44 46 47 48
r80 42 44 21.652 $w=3.28e-07 $l=6.2e-07 $layer=LI1_cond $X=8.23 $Y=2.905
+ $X2=8.23 $Y2=2.285
r81 41 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.495 $Y=2.99
+ $X2=7.33 $Y2=2.99
r82 40 42 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=8.065 $Y=2.99
+ $X2=8.23 $Y2=2.905
r83 40 41 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=8.065 $Y=2.99
+ $X2=7.495 $Y2=2.99
r84 36 48 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.33 $Y=2.905
+ $X2=7.33 $Y2=2.99
r85 36 38 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=7.33 $Y=2.905
+ $X2=7.33 $Y2=2.455
r86 35 47 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=6.595 $Y=2.99
+ $X2=6.455 $Y2=2.99
r87 34 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.165 $Y=2.99
+ $X2=7.33 $Y2=2.99
r88 34 35 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=7.165 $Y=2.99
+ $X2=6.595 $Y2=2.99
r89 30 33 28.8111 $w=2.78e-07 $l=7e-07 $layer=LI1_cond $X=6.455 $Y=2.115
+ $X2=6.455 $Y2=2.815
r90 28 47 0.375625 $w=2.8e-07 $l=8.5e-08 $layer=LI1_cond $X=6.455 $Y=2.905
+ $X2=6.455 $Y2=2.99
r91 28 33 3.70428 $w=2.78e-07 $l=9e-08 $layer=LI1_cond $X=6.455 $Y=2.905
+ $X2=6.455 $Y2=2.815
r92 27 46 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.695 $Y=2.99
+ $X2=5.53 $Y2=2.99
r93 26 47 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=6.315 $Y=2.99
+ $X2=6.455 $Y2=2.99
r94 26 27 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=6.315 $Y=2.99
+ $X2=5.695 $Y2=2.99
r95 22 46 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.53 $Y=2.905
+ $X2=5.53 $Y2=2.99
r96 22 24 17.8105 $w=3.28e-07 $l=5.1e-07 $layer=LI1_cond $X=5.53 $Y=2.905
+ $X2=5.53 $Y2=2.395
r97 20 46 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.365 $Y=2.99
+ $X2=5.53 $Y2=2.99
r98 20 21 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=5.365 $Y=2.99
+ $X2=4.795 $Y2=2.99
r99 16 21 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.63 $Y=2.905
+ $X2=4.795 $Y2=2.99
r100 16 18 17.8105 $w=3.28e-07 $l=5.1e-07 $layer=LI1_cond $X=4.63 $Y=2.905
+ $X2=4.63 $Y2=2.395
r101 5 44 300 $w=1.7e-07 $l=5.14563e-07 $layer=licon1_PDIFF $count=2 $X=8.08
+ $Y=1.84 $X2=8.23 $Y2=2.285
r102 4 38 300 $w=1.7e-07 $l=6.85912e-07 $layer=licon1_PDIFF $count=2 $X=7.18
+ $Y=1.84 $X2=7.33 $Y2=2.455
r103 3 33 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=6.28
+ $Y=1.84 $X2=6.43 $Y2=2.815
r104 3 30 400 $w=1.7e-07 $l=3.4187e-07 $layer=licon1_PDIFF $count=1 $X=6.28
+ $Y=1.84 $X2=6.43 $Y2=2.115
r105 2 24 300 $w=1.7e-07 $l=6.2552e-07 $layer=licon1_PDIFF $count=2 $X=5.38
+ $Y=1.84 $X2=5.53 $Y2=2.395
r106 1 18 300 $w=1.7e-07 $l=6.14329e-07 $layer=licon1_PDIFF $count=2 $X=4.505
+ $Y=1.84 $X2=4.63 $Y2=2.395
.ends

.subckt PM_SKY130_FD_SC_HS__A211OI_4%Y 1 2 3 4 5 6 7 22 26 30 32 36 38 42 48 49
+ 50 52 53 54 55 56 57 58 59 60
c77 22 0 4.29123e-20 $X=3.588 $Y=0.957
r78 56 60 11.6415 $w=1.7e-07 $l=5.53e-07 $layer=LI1_cond $X=7.847 $Y=1.665
+ $X2=8.4 $Y2=1.665
r79 55 56 4.56883 $w=9.88e-07 $l=3.7e-07 $layer=LI1_cond $X=7.847 $Y=1.295
+ $X2=7.847 $Y2=1.665
r80 55 59 11.6415 $w=1.7e-07 $l=5.53e-07 $layer=LI1_cond $X=7.847 $Y=1.295
+ $X2=8.4 $Y2=1.295
r81 55 77 2.46964 $w=9.88e-07 $l=2e-07 $layer=LI1_cond $X=7.847 $Y=1.295
+ $X2=7.847 $Y2=1.095
r82 54 77 2.09919 $w=9.88e-07 $l=1.7e-07 $layer=LI1_cond $X=7.847 $Y=0.925
+ $X2=7.847 $Y2=1.095
r83 54 58 11.6415 $w=1.7e-07 $l=5.53e-07 $layer=LI1_cond $X=7.847 $Y=0.925
+ $X2=8.4 $Y2=0.925
r84 53 54 4.56883 $w=9.88e-07 $l=3.7e-07 $layer=LI1_cond $X=7.847 $Y=0.555
+ $X2=7.847 $Y2=0.925
r85 53 57 11.6415 $w=1.7e-07 $l=5.53e-07 $layer=LI1_cond $X=7.847 $Y=0.555
+ $X2=8.4 $Y2=0.555
r86 53 70 0.493927 $w=9.88e-07 $l=4e-08 $layer=LI1_cond $X=7.847 $Y=0.555
+ $X2=7.847 $Y2=0.515
r87 47 48 8.4794 $w=3.43e-07 $l=1.65e-07 $layer=LI1_cond $X=3.595 $Y=0.957
+ $X2=3.76 $Y2=0.957
r88 43 52 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.965 $Y=2.035
+ $X2=6.88 $Y2=2.035
r89 42 56 4.56883 $w=9.88e-07 $l=3.7e-07 $layer=LI1_cond $X=7.847 $Y=2.035
+ $X2=7.847 $Y2=1.665
r90 42 43 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=7.695 $Y=2.035
+ $X2=6.965 $Y2=2.035
r91 39 50 5.16603 $w=1.7e-07 $l=9.66954e-08 $layer=LI1_cond $X=6.49 $Y=1.095
+ $X2=6.405 $Y2=1.07
r92 38 77 11.6415 $w=1.7e-07 $l=6.67e-07 $layer=LI1_cond $X=7.18 $Y=1.095
+ $X2=7.847 $Y2=1.095
r93 38 39 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=7.18 $Y=1.095
+ $X2=6.49 $Y2=1.095
r94 34 50 1.34256 $w=1.7e-07 $l=1.1e-07 $layer=LI1_cond $X=6.405 $Y=0.96
+ $X2=6.405 $Y2=1.07
r95 34 36 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=6.405 $Y=0.96
+ $X2=6.405 $Y2=0.515
r96 33 49 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.63 $Y=1.045
+ $X2=5.505 $Y2=1.045
r97 32 50 5.16603 $w=1.7e-07 $l=9.66954e-08 $layer=LI1_cond $X=6.32 $Y=1.045
+ $X2=6.405 $Y2=1.07
r98 32 33 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=6.32 $Y=1.045
+ $X2=5.63 $Y2=1.045
r99 28 49 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.505 $Y=0.96
+ $X2=5.505 $Y2=1.045
r100 28 30 20.5135 $w=2.48e-07 $l=4.45e-07 $layer=LI1_cond $X=5.505 $Y=0.96
+ $X2=5.505 $Y2=0.515
r101 26 49 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.38 $Y=1.045
+ $X2=5.505 $Y2=1.045
r102 26 48 105.69 $w=1.68e-07 $l=1.62e-06 $layer=LI1_cond $X=5.38 $Y=1.045
+ $X2=3.76 $Y2=1.045
r103 22 47 0.233829 $w=3.43e-07 $l=7e-09 $layer=LI1_cond $X=3.588 $Y=0.957
+ $X2=3.595 $Y2=0.957
r104 22 24 28.4937 $w=3.43e-07 $l=8.53e-07 $layer=LI1_cond $X=3.588 $Y=0.957
+ $X2=2.735 $Y2=0.957
r105 7 42 300 $w=1.7e-07 $l=3.4187e-07 $layer=licon1_PDIFF $count=2 $X=7.63
+ $Y=1.84 $X2=7.78 $Y2=2.115
r106 6 52 300 $w=1.7e-07 $l=3.4187e-07 $layer=licon1_PDIFF $count=2 $X=6.73
+ $Y=1.84 $X2=6.88 $Y2=2.115
r107 5 70 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=7.125
+ $Y=0.37 $X2=7.265 $Y2=0.515
r108 4 36 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=6.265
+ $Y=0.37 $X2=6.405 $Y2=0.515
r109 3 30 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=5.42
+ $Y=0.37 $X2=5.545 $Y2=0.515
r110 2 47 182 $w=1.7e-07 $l=6.4622e-07 $layer=licon1_NDIFF $count=1 $X=3.455
+ $Y=0.37 $X2=3.595 $Y2=0.95
r111 1 24 182 $w=1.7e-07 $l=6.4622e-07 $layer=licon1_NDIFF $count=1 $X=2.595
+ $Y=0.37 $X2=2.735 $Y2=0.95
.ends

.subckt PM_SKY130_FD_SC_HS__A211OI_4%A_92_74# 1 2 3 4 5 18 20 21 24 26 28 36 38
c51 28 0 1.6164e-19 $X=2.305 $Y=0.615
r52 34 36 37.4 $w=2.63e-07 $l=8.6e-07 $layer=LI1_cond $X=3.165 $Y=0.482
+ $X2=4.025 $Y2=0.482
r53 32 40 2.82608 $w=2.65e-07 $l=8.5e-08 $layer=LI1_cond $X=2.39 $Y=0.482
+ $X2=2.305 $Y2=0.482
r54 32 34 33.7035 $w=2.63e-07 $l=7.75e-07 $layer=LI1_cond $X=2.39 $Y=0.482
+ $X2=3.165 $Y2=0.482
r55 29 31 2.93583 $w=1.68e-07 $l=4.5e-08 $layer=LI1_cond $X=2.305 $Y=1.01
+ $X2=2.305 $Y2=0.965
r56 28 40 4.42198 $w=1.7e-07 $l=1.33e-07 $layer=LI1_cond $X=2.305 $Y=0.615
+ $X2=2.305 $Y2=0.482
r57 28 31 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=2.305 $Y=0.615
+ $X2=2.305 $Y2=0.965
r58 27 38 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.53 $Y=1.095
+ $X2=1.445 $Y2=1.095
r59 26 29 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.22 $Y=1.095
+ $X2=2.305 $Y2=1.01
r60 26 27 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=2.22 $Y=1.095
+ $X2=1.53 $Y2=1.095
r61 22 38 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.445 $Y=1.01
+ $X2=1.445 $Y2=1.095
r62 22 24 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=1.445 $Y=1.01
+ $X2=1.445 $Y2=0.515
r63 20 38 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.36 $Y=1.095
+ $X2=1.445 $Y2=1.095
r64 20 21 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.36 $Y=1.095
+ $X2=0.67 $Y2=1.095
r65 16 21 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.545 $Y=1.01
+ $X2=0.67 $Y2=1.095
r66 16 18 22.8184 $w=2.48e-07 $l=4.95e-07 $layer=LI1_cond $X=0.545 $Y=1.01
+ $X2=0.545 $Y2=0.515
r67 5 36 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=3.885
+ $Y=0.37 $X2=4.025 $Y2=0.515
r68 4 34 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=3.025
+ $Y=0.37 $X2=3.165 $Y2=0.515
r69 3 40 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=2.165
+ $Y=0.37 $X2=2.305 $Y2=0.515
r70 3 31 182 $w=1.7e-07 $l=6.61306e-07 $layer=licon1_NDIFF $count=1 $X=2.165
+ $Y=0.37 $X2=2.305 $Y2=0.965
r71 2 24 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.305
+ $Y=0.37 $X2=1.445 $Y2=0.515
r72 1 18 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.46
+ $Y=0.37 $X2=0.585 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__A211OI_4%VGND 1 2 3 4 15 19 23 27 30 31 33 34 35 44
+ 51 58 59 62 65
r81 65 66 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.96 $Y=0 $X2=6.96
+ $Y2=0
r82 62 63 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=0 $X2=6 $Y2=0
r83 59 66 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=8.4 $Y=0 $X2=6.96
+ $Y2=0
r84 58 59 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r85 56 65 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7 $Y=0 $X2=6.835
+ $Y2=0
r86 56 58 91.3369 $w=1.68e-07 $l=1.4e-06 $layer=LI1_cond $X=7 $Y=0 $X2=8.4 $Y2=0
r87 55 66 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=0 $X2=6.96
+ $Y2=0
r88 55 63 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=0 $X2=6
+ $Y2=0
r89 54 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=0 $X2=6.48
+ $Y2=0
r90 52 62 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.14 $Y=0 $X2=5.975
+ $Y2=0
r91 52 54 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=6.14 $Y=0 $X2=6.48
+ $Y2=0
r92 51 65 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.67 $Y=0 $X2=6.835
+ $Y2=0
r93 51 54 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=6.67 $Y=0 $X2=6.48
+ $Y2=0
r94 50 63 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=6
+ $Y2=0
r95 49 50 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r96 46 49 219.209 $w=1.68e-07 $l=3.36e-06 $layer=LI1_cond $X=2.16 $Y=0 $X2=5.52
+ $Y2=0
r97 46 47 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r98 44 62 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.81 $Y=0 $X2=5.975
+ $Y2=0
r99 44 49 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=5.81 $Y=0 $X2=5.52
+ $Y2=0
r100 43 47 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r101 42 43 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r102 39 43 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r103 38 39 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r104 35 50 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=4.32 $Y=0 $X2=5.52
+ $Y2=0
r105 35 47 0.602067 $w=4.9e-07 $l=2.16e-06 $layer=MET1_cond $X=4.32 $Y=0
+ $X2=2.16 $Y2=0
r106 33 42 1.95722 $w=1.68e-07 $l=3e-08 $layer=LI1_cond $X=1.71 $Y=0 $X2=1.68
+ $Y2=0
r107 33 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.71 $Y=0 $X2=1.875
+ $Y2=0
r108 32 46 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=2.04 $Y=0 $X2=2.16
+ $Y2=0
r109 32 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.04 $Y=0 $X2=1.875
+ $Y2=0
r110 30 38 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=0.85 $Y=0 $X2=0.72
+ $Y2=0
r111 30 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.85 $Y=0 $X2=1.015
+ $Y2=0
r112 29 42 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=1.18 $Y=0 $X2=1.68
+ $Y2=0
r113 29 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.18 $Y=0 $X2=1.015
+ $Y2=0
r114 25 65 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.835 $Y=0.085
+ $X2=6.835 $Y2=0
r115 25 27 20.6043 $w=3.28e-07 $l=5.9e-07 $layer=LI1_cond $X=6.835 $Y=0.085
+ $X2=6.835 $Y2=0.675
r116 21 62 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.975 $Y=0.085
+ $X2=5.975 $Y2=0
r117 21 23 18.8582 $w=3.28e-07 $l=5.4e-07 $layer=LI1_cond $X=5.975 $Y=0.085
+ $X2=5.975 $Y2=0.625
r118 17 34 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.875 $Y=0.085
+ $X2=1.875 $Y2=0
r119 17 19 20.6043 $w=3.28e-07 $l=5.9e-07 $layer=LI1_cond $X=1.875 $Y=0.085
+ $X2=1.875 $Y2=0.675
r120 13 31 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.015 $Y=0.085
+ $X2=1.015 $Y2=0
r121 13 15 20.6043 $w=3.28e-07 $l=5.9e-07 $layer=LI1_cond $X=1.015 $Y=0.085
+ $X2=1.015 $Y2=0.675
r122 4 27 182 $w=1.7e-07 $l=3.68409e-07 $layer=licon1_NDIFF $count=1 $X=6.695
+ $Y=0.37 $X2=6.835 $Y2=0.675
r123 3 23 182 $w=1.7e-07 $l=3.17372e-07 $layer=licon1_NDIFF $count=1 $X=5.835
+ $Y=0.37 $X2=5.975 $Y2=0.625
r124 2 19 182 $w=1.7e-07 $l=3.68409e-07 $layer=licon1_NDIFF $count=1 $X=1.735
+ $Y=0.37 $X2=1.875 $Y2=0.675
r125 1 15 182 $w=1.7e-07 $l=3.68409e-07 $layer=licon1_NDIFF $count=1 $X=0.875
+ $Y=0.37 $X2=1.015 $Y2=0.675
.ends

