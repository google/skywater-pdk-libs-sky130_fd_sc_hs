* File: sky130_fd_sc_hs__o21ai_2.pxi.spice
* Created: Tue Sep  1 20:14:36 2020
* 
x_PM_SKY130_FD_SC_HS__O21AI_2%A1 N_A1_M1009_g N_A1_c_63_n N_A1_M1002_g
+ N_A1_M1010_g N_A1_c_65_n N_A1_M1005_g N_A1_c_66_n N_A1_c_74_p N_A1_c_96_p A1
+ N_A1_c_67_n PM_SKY130_FD_SC_HS__O21AI_2%A1
x_PM_SKY130_FD_SC_HS__O21AI_2%A2 N_A2_c_140_n N_A2_M1003_g N_A2_M1001_g
+ N_A2_M1011_g N_A2_c_141_n N_A2_M1004_g A2 N_A2_c_138_n N_A2_c_139_n
+ PM_SKY130_FD_SC_HS__O21AI_2%A2
x_PM_SKY130_FD_SC_HS__O21AI_2%B1 N_B1_M1000_g N_B1_c_194_n N_B1_M1006_g
+ N_B1_c_195_n N_B1_c_196_n N_B1_M1008_g N_B1_c_197_n N_B1_M1007_g B1
+ PM_SKY130_FD_SC_HS__O21AI_2%B1
x_PM_SKY130_FD_SC_HS__O21AI_2%VPWR N_VPWR_M1002_d N_VPWR_M1005_d N_VPWR_M1008_s
+ N_VPWR_c_240_n N_VPWR_c_241_n N_VPWR_c_242_n N_VPWR_c_243_n N_VPWR_c_244_n
+ VPWR N_VPWR_c_245_n N_VPWR_c_246_n N_VPWR_c_247_n N_VPWR_c_239_n
+ PM_SKY130_FD_SC_HS__O21AI_2%VPWR
x_PM_SKY130_FD_SC_HS__O21AI_2%A_116_368# N_A_116_368#_M1002_s
+ N_A_116_368#_M1004_s N_A_116_368#_c_294_n N_A_116_368#_c_288_n
+ N_A_116_368#_c_289_n N_A_116_368#_c_290_n
+ PM_SKY130_FD_SC_HS__O21AI_2%A_116_368#
x_PM_SKY130_FD_SC_HS__O21AI_2%Y N_Y_M1000_d N_Y_M1003_d N_Y_M1006_d N_Y_c_325_n
+ N_Y_c_360_p N_Y_c_327_n N_Y_c_319_n Y Y Y Y N_Y_c_320_n
+ PM_SKY130_FD_SC_HS__O21AI_2%Y
x_PM_SKY130_FD_SC_HS__O21AI_2%A_27_74# N_A_27_74#_M1009_d N_A_27_74#_M1001_d
+ N_A_27_74#_M1010_d N_A_27_74#_M1007_s N_A_27_74#_c_361_n N_A_27_74#_c_362_n
+ N_A_27_74#_c_363_n N_A_27_74#_c_364_n N_A_27_74#_c_365_n N_A_27_74#_c_366_n
+ N_A_27_74#_c_367_n N_A_27_74#_c_368_n N_A_27_74#_c_369_n
+ PM_SKY130_FD_SC_HS__O21AI_2%A_27_74#
x_PM_SKY130_FD_SC_HS__O21AI_2%VGND N_VGND_M1009_s N_VGND_M1011_s N_VGND_c_421_n
+ N_VGND_c_422_n VGND N_VGND_c_423_n N_VGND_c_424_n N_VGND_c_425_n
+ N_VGND_c_426_n N_VGND_c_427_n N_VGND_c_428_n PM_SKY130_FD_SC_HS__O21AI_2%VGND
cc_1 VNB N_A1_M1009_g 0.0340607f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_2 VNB N_A1_c_63_n 0.0374247f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.765
cc_3 VNB N_A1_M1010_g 0.0246779f $X=-0.19 $Y=-0.245 $X2=1.925 $Y2=0.74
cc_4 VNB N_A1_c_65_n 0.0248396f $X=-0.19 $Y=-0.245 $X2=1.955 $Y2=1.765
cc_5 VNB N_A1_c_66_n 0.00166865f $X=-0.19 $Y=-0.245 $X2=0.43 $Y2=1.515
cc_6 VNB N_A1_c_67_n 0.00562447f $X=-0.19 $Y=-0.245 $X2=1.92 $Y2=1.515
cc_7 VNB N_A2_M1001_g 0.0239739f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_8 VNB N_A2_M1011_g 0.0245225f $X=-0.19 $Y=-0.245 $X2=1.925 $Y2=0.74
cc_9 VNB N_A2_c_138_n 0.00175883f $X=-0.19 $Y=-0.245 $X2=0.595 $Y2=2.035
cc_10 VNB N_A2_c_139_n 0.040003f $X=-0.19 $Y=-0.245 $X2=2.015 $Y2=1.95
cc_11 VNB N_B1_M1000_g 0.0262343f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_12 VNB N_B1_c_194_n 0.011794f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.765
cc_13 VNB N_B1_c_195_n 0.0186258f $X=-0.19 $Y=-0.245 $X2=1.925 $Y2=1.35
cc_14 VNB N_B1_c_196_n 0.0619018f $X=-0.19 $Y=-0.245 $X2=1.925 $Y2=0.74
cc_15 VNB N_B1_c_197_n 0.0233164f $X=-0.19 $Y=-0.245 $X2=1.955 $Y2=2.4
cc_16 VNB B1 0.00877571f $X=-0.19 $Y=-0.245 $X2=0.43 $Y2=1.515
cc_17 VNB N_VPWR_c_239_n 0.143779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_Y_c_319_n 0.00235393f $X=-0.19 $Y=-0.245 $X2=2.075 $Y2=1.58
cc_19 VNB N_Y_c_320_n 0.00472487f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_27_74#_c_361_n 0.0277086f $X=-0.19 $Y=-0.245 $X2=0.43 $Y2=1.95
cc_21 VNB N_A_27_74#_c_362_n 0.00973995f $X=-0.19 $Y=-0.245 $X2=0.43 $Y2=1.515
cc_22 VNB N_A_27_74#_c_363_n 0.0143688f $X=-0.19 $Y=-0.245 $X2=0.43 $Y2=1.515
cc_23 VNB N_A_27_74#_c_364_n 0.00220643f $X=-0.19 $Y=-0.245 $X2=0.595 $Y2=2.035
cc_24 VNB N_A_27_74#_c_365_n 0.0124022f $X=-0.19 $Y=-0.245 $X2=2.075 $Y2=1.58
cc_25 VNB N_A_27_74#_c_366_n 0.00232545f $X=-0.19 $Y=-0.245 $X2=0.43 $Y2=1.515
cc_26 VNB N_A_27_74#_c_367_n 0.00279725f $X=-0.19 $Y=-0.245 $X2=1.92 $Y2=1.515
cc_27 VNB N_A_27_74#_c_368_n 0.00187632f $X=-0.19 $Y=-0.245 $X2=2.015 $Y2=1.665
cc_28 VNB N_A_27_74#_c_369_n 0.0287634f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_421_n 0.00578139f $X=-0.19 $Y=-0.245 $X2=1.925 $Y2=0.74
cc_30 VNB N_VGND_c_422_n 0.00557884f $X=-0.19 $Y=-0.245 $X2=1.955 $Y2=2.4
cc_31 VNB N_VGND_c_423_n 0.0191515f $X=-0.19 $Y=-0.245 $X2=0.43 $Y2=1.515
cc_32 VNB N_VGND_c_424_n 0.0169342f $X=-0.19 $Y=-0.245 $X2=2.015 $Y2=1.95
cc_33 VNB N_VGND_c_425_n 0.0399491f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_426_n 0.207539f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_427_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_428_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VPB N_A1_c_63_n 0.0289996f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.765
cc_38 VPB N_A1_c_65_n 0.0255169f $X=-0.19 $Y=1.66 $X2=1.955 $Y2=1.765
cc_39 VPB N_A1_c_66_n 0.00674617f $X=-0.19 $Y=1.66 $X2=0.43 $Y2=1.515
cc_40 VPB N_A1_c_67_n 0.00264206f $X=-0.19 $Y=1.66 $X2=1.92 $Y2=1.515
cc_41 VPB N_A2_c_140_n 0.0151474f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.35
cc_42 VPB N_A2_c_141_n 0.0155885f $X=-0.19 $Y=1.66 $X2=1.955 $Y2=1.765
cc_43 VPB N_A2_c_138_n 0.00430556f $X=-0.19 $Y=1.66 $X2=0.595 $Y2=2.035
cc_44 VPB N_A2_c_139_n 0.0221376f $X=-0.19 $Y=1.66 $X2=2.015 $Y2=1.95
cc_45 VPB N_B1_c_194_n 0.0218396f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.765
cc_46 VPB N_B1_c_196_n 0.0276353f $X=-0.19 $Y=1.66 $X2=1.925 $Y2=0.74
cc_47 VPB N_VPWR_c_240_n 0.0106521f $X=-0.19 $Y=1.66 $X2=1.925 $Y2=0.74
cc_48 VPB N_VPWR_c_241_n 0.0373712f $X=-0.19 $Y=1.66 $X2=1.955 $Y2=1.765
cc_49 VPB N_VPWR_c_242_n 0.00481327f $X=-0.19 $Y=1.66 $X2=0.43 $Y2=1.515
cc_50 VPB N_VPWR_c_243_n 0.0106521f $X=-0.19 $Y=1.66 $X2=0.43 $Y2=1.515
cc_51 VPB N_VPWR_c_244_n 0.055977f $X=-0.19 $Y=1.66 $X2=1.755 $Y2=2.035
cc_52 VPB N_VPWR_c_245_n 0.0419554f $X=-0.19 $Y=1.66 $X2=1.92 $Y2=1.515
cc_53 VPB N_VPWR_c_246_n 0.0183691f $X=-0.19 $Y=1.66 $X2=2.015 $Y2=1.665
cc_54 VPB N_VPWR_c_247_n 0.00460249f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_55 VPB N_VPWR_c_239_n 0.0637314f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_56 VPB N_A_116_368#_c_288_n 0.00297669f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_57 VPB N_A_116_368#_c_289_n 0.0021839f $X=-0.19 $Y=1.66 $X2=1.955 $Y2=1.765
cc_58 VPB N_A_116_368#_c_290_n 0.00248006f $X=-0.19 $Y=1.66 $X2=1.955 $Y2=2.4
cc_59 VPB Y 6.90925e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_60 VPB Y 0.0023458f $X=-0.19 $Y=1.66 $X2=0.43 $Y2=1.515
cc_61 VPB N_Y_c_320_n 0.00258439f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_62 N_A1_c_63_n N_A2_c_140_n 0.0261308f $X=0.505 $Y=1.765 $X2=-0.19 $Y2=-0.245
cc_63 N_A1_c_66_n N_A2_c_140_n 0.00159252f $X=0.43 $Y=1.515 $X2=-0.19 $Y2=-0.245
cc_64 N_A1_c_74_p N_A2_c_140_n 0.0151016f $X=1.755 $Y=2.035 $X2=-0.19 $Y2=-0.245
cc_65 N_A1_M1009_g N_A2_M1001_g 0.0292811f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_66 N_A1_M1010_g N_A2_M1011_g 0.0256098f $X=1.925 $Y=0.74 $X2=0 $Y2=0
cc_67 N_A1_c_65_n N_A2_c_141_n 0.0387077f $X=1.955 $Y=1.765 $X2=0 $Y2=0
cc_68 N_A1_c_74_p N_A2_c_141_n 0.0116004f $X=1.755 $Y=2.035 $X2=0 $Y2=0
cc_69 N_A1_c_67_n N_A2_c_141_n 0.00429709f $X=1.92 $Y=1.515 $X2=0 $Y2=0
cc_70 N_A1_c_63_n N_A2_c_138_n 0.00185053f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_71 N_A1_c_65_n N_A2_c_138_n 0.00125098f $X=1.955 $Y=1.765 $X2=0 $Y2=0
cc_72 N_A1_c_66_n N_A2_c_138_n 0.0255979f $X=0.43 $Y=1.515 $X2=0 $Y2=0
cc_73 N_A1_c_74_p N_A2_c_138_n 0.0461579f $X=1.755 $Y=2.035 $X2=0 $Y2=0
cc_74 N_A1_c_67_n N_A2_c_138_n 0.0271976f $X=1.92 $Y=1.515 $X2=0 $Y2=0
cc_75 N_A1_c_63_n N_A2_c_139_n 0.0209265f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_76 N_A1_c_65_n N_A2_c_139_n 0.022834f $X=1.955 $Y=1.765 $X2=0 $Y2=0
cc_77 N_A1_c_66_n N_A2_c_139_n 0.00152602f $X=0.43 $Y=1.515 $X2=0 $Y2=0
cc_78 N_A1_c_74_p N_A2_c_139_n 0.00157644f $X=1.755 $Y=2.035 $X2=0 $Y2=0
cc_79 N_A1_c_67_n N_A2_c_139_n 0.00198112f $X=1.92 $Y=1.515 $X2=0 $Y2=0
cc_80 N_A1_M1010_g N_B1_M1000_g 0.0156839f $X=1.925 $Y=0.74 $X2=0 $Y2=0
cc_81 N_A1_c_65_n N_B1_M1000_g 0.00921114f $X=1.955 $Y=1.765 $X2=0 $Y2=0
cc_82 N_A1_c_67_n N_B1_M1000_g 0.00173955f $X=1.92 $Y=1.515 $X2=0 $Y2=0
cc_83 N_A1_c_65_n N_B1_c_194_n 0.0510023f $X=1.955 $Y=1.765 $X2=0 $Y2=0
cc_84 N_A1_c_67_n N_B1_c_194_n 0.00358933f $X=1.92 $Y=1.515 $X2=0 $Y2=0
cc_85 N_A1_c_66_n N_VPWR_M1002_d 0.00450592f $X=0.43 $Y=1.515 $X2=-0.19
+ $Y2=-0.245
cc_86 N_A1_c_96_p N_VPWR_M1002_d 0.00915927f $X=0.595 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_87 N_A1_c_74_p N_VPWR_M1005_d 0.0026248f $X=1.755 $Y=2.035 $X2=0 $Y2=0
cc_88 N_A1_c_67_n N_VPWR_M1005_d 2.48634e-19 $X=1.92 $Y=1.515 $X2=0 $Y2=0
cc_89 N_A1_c_63_n N_VPWR_c_241_n 0.00577175f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_90 N_A1_c_96_p N_VPWR_c_241_n 0.00888093f $X=0.595 $Y=2.035 $X2=0 $Y2=0
cc_91 N_A1_c_65_n N_VPWR_c_242_n 0.00239895f $X=1.955 $Y=1.765 $X2=0 $Y2=0
cc_92 N_A1_c_63_n N_VPWR_c_245_n 0.0044313f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_93 N_A1_c_65_n N_VPWR_c_245_n 0.00444353f $X=1.955 $Y=1.765 $X2=0 $Y2=0
cc_94 N_A1_c_63_n N_VPWR_c_239_n 0.00856939f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_95 N_A1_c_65_n N_VPWR_c_239_n 0.00857665f $X=1.955 $Y=1.765 $X2=0 $Y2=0
cc_96 N_A1_c_74_p N_A_116_368#_M1002_s 0.00907415f $X=1.755 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_97 N_A1_c_74_p N_A_116_368#_M1004_s 0.00889481f $X=1.755 $Y=2.035 $X2=0 $Y2=0
cc_98 N_A1_c_67_n N_A_116_368#_M1004_s 0.00150594f $X=1.92 $Y=1.515 $X2=0 $Y2=0
cc_99 N_A1_c_63_n N_A_116_368#_c_294_n 0.00678385f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_100 N_A1_c_74_p N_A_116_368#_c_294_n 0.016157f $X=1.755 $Y=2.035 $X2=0 $Y2=0
cc_101 N_A1_c_96_p N_A_116_368#_c_294_n 0.00114279f $X=0.595 $Y=2.035 $X2=0
+ $Y2=0
cc_102 N_A1_c_63_n N_A_116_368#_c_289_n 0.00332677f $X=0.505 $Y=1.765 $X2=0
+ $Y2=0
cc_103 N_A1_c_65_n N_A_116_368#_c_290_n 0.00615477f $X=1.955 $Y=1.765 $X2=0
+ $Y2=0
cc_104 N_A1_c_74_p N_Y_M1003_d 0.00455513f $X=1.755 $Y=2.035 $X2=0 $Y2=0
cc_105 N_A1_c_65_n N_Y_c_325_n 0.0150988f $X=1.955 $Y=1.765 $X2=0 $Y2=0
cc_106 N_A1_c_74_p N_Y_c_325_n 0.0533629f $X=1.755 $Y=2.035 $X2=0 $Y2=0
cc_107 N_A1_c_65_n N_Y_c_327_n 8.24416e-19 $X=1.955 $Y=1.765 $X2=0 $Y2=0
cc_108 N_A1_c_74_p N_Y_c_327_n 0.0195846f $X=1.755 $Y=2.035 $X2=0 $Y2=0
cc_109 N_A1_c_67_n N_Y_c_320_n 0.0301739f $X=1.92 $Y=1.515 $X2=0 $Y2=0
cc_110 N_A1_M1009_g N_A_27_74#_c_361_n 0.0101985f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_111 N_A1_M1009_g N_A_27_74#_c_362_n 0.0114775f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_112 N_A1_c_66_n N_A_27_74#_c_362_n 0.0114058f $X=0.43 $Y=1.515 $X2=0 $Y2=0
cc_113 N_A1_M1009_g N_A_27_74#_c_363_n 0.00214612f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_114 N_A1_c_63_n N_A_27_74#_c_363_n 0.00121873f $X=0.505 $Y=1.765 $X2=0 $Y2=0
cc_115 N_A1_c_66_n N_A_27_74#_c_363_n 0.0158461f $X=0.43 $Y=1.515 $X2=0 $Y2=0
cc_116 N_A1_M1010_g N_A_27_74#_c_364_n 9.34885e-19 $X=1.925 $Y=0.74 $X2=0 $Y2=0
cc_117 N_A1_M1010_g N_A_27_74#_c_365_n 0.0133221f $X=1.925 $Y=0.74 $X2=0 $Y2=0
cc_118 N_A1_c_65_n N_A_27_74#_c_365_n 0.00128239f $X=1.955 $Y=1.765 $X2=0 $Y2=0
cc_119 N_A1_c_67_n N_A_27_74#_c_365_n 0.0436794f $X=1.92 $Y=1.515 $X2=0 $Y2=0
cc_120 N_A1_M1009_g N_VGND_c_421_n 0.00565822f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_121 N_A1_M1010_g N_VGND_c_422_n 0.0106192f $X=1.925 $Y=0.74 $X2=0 $Y2=0
cc_122 N_A1_M1009_g N_VGND_c_423_n 0.00434272f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_123 N_A1_M1010_g N_VGND_c_425_n 0.00383152f $X=1.925 $Y=0.74 $X2=0 $Y2=0
cc_124 N_A1_M1009_g N_VGND_c_426_n 0.00824429f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_125 N_A1_M1010_g N_VGND_c_426_n 0.00758041f $X=1.925 $Y=0.74 $X2=0 $Y2=0
cc_126 N_A2_c_140_n N_VPWR_c_245_n 0.00278257f $X=0.955 $Y=1.765 $X2=0 $Y2=0
cc_127 N_A2_c_141_n N_VPWR_c_245_n 0.00278271f $X=1.455 $Y=1.765 $X2=0 $Y2=0
cc_128 N_A2_c_140_n N_VPWR_c_239_n 0.00354366f $X=0.955 $Y=1.765 $X2=0 $Y2=0
cc_129 N_A2_c_141_n N_VPWR_c_239_n 0.00354798f $X=1.455 $Y=1.765 $X2=0 $Y2=0
cc_130 N_A2_c_140_n N_A_116_368#_c_294_n 0.0076826f $X=0.955 $Y=1.765 $X2=0
+ $Y2=0
cc_131 N_A2_c_141_n N_A_116_368#_c_294_n 6.5039e-19 $X=1.455 $Y=1.765 $X2=0
+ $Y2=0
cc_132 N_A2_c_140_n N_A_116_368#_c_288_n 0.011054f $X=0.955 $Y=1.765 $X2=0 $Y2=0
cc_133 N_A2_c_141_n N_A_116_368#_c_288_n 0.00978708f $X=1.455 $Y=1.765 $X2=0
+ $Y2=0
cc_134 N_A2_c_140_n N_A_116_368#_c_289_n 0.00171731f $X=0.955 $Y=1.765 $X2=0
+ $Y2=0
cc_135 N_A2_c_141_n N_A_116_368#_c_290_n 5.05939e-19 $X=1.455 $Y=1.765 $X2=0
+ $Y2=0
cc_136 N_A2_c_141_n N_Y_c_325_n 0.00996205f $X=1.455 $Y=1.765 $X2=0 $Y2=0
cc_137 N_A2_c_141_n N_Y_c_327_n 0.00596455f $X=1.455 $Y=1.765 $X2=0 $Y2=0
cc_138 N_A2_M1001_g N_A_27_74#_c_361_n 9.46832e-19 $X=0.995 $Y=0.74 $X2=0 $Y2=0
cc_139 N_A2_M1001_g N_A_27_74#_c_362_n 0.0134647f $X=0.995 $Y=0.74 $X2=0 $Y2=0
cc_140 N_A2_c_138_n N_A_27_74#_c_362_n 0.0209068f $X=1.35 $Y=1.515 $X2=0 $Y2=0
cc_141 N_A2_c_139_n N_A_27_74#_c_362_n 5.17477e-19 $X=1.44 $Y=1.557 $X2=0 $Y2=0
cc_142 N_A2_M1001_g N_A_27_74#_c_364_n 4.13268e-19 $X=0.995 $Y=0.74 $X2=0 $Y2=0
cc_143 N_A2_M1011_g N_A_27_74#_c_364_n 0.00837823f $X=1.44 $Y=0.74 $X2=0 $Y2=0
cc_144 N_A2_M1011_g N_A_27_74#_c_365_n 0.0124938f $X=1.44 $Y=0.74 $X2=0 $Y2=0
cc_145 N_A2_c_138_n N_A_27_74#_c_365_n 0.0101599f $X=1.35 $Y=1.515 $X2=0 $Y2=0
cc_146 N_A2_c_139_n N_A_27_74#_c_365_n 9.98122e-19 $X=1.44 $Y=1.557 $X2=0 $Y2=0
cc_147 N_A2_M1011_g N_A_27_74#_c_368_n 0.00115653f $X=1.44 $Y=0.74 $X2=0 $Y2=0
cc_148 N_A2_c_138_n N_A_27_74#_c_368_n 0.0215332f $X=1.35 $Y=1.515 $X2=0 $Y2=0
cc_149 N_A2_c_139_n N_A_27_74#_c_368_n 9.10195e-19 $X=1.44 $Y=1.557 $X2=0 $Y2=0
cc_150 N_A2_M1001_g N_VGND_c_421_n 0.0106183f $X=0.995 $Y=0.74 $X2=0 $Y2=0
cc_151 N_A2_M1011_g N_VGND_c_421_n 5.10607e-19 $X=1.44 $Y=0.74 $X2=0 $Y2=0
cc_152 N_A2_M1011_g N_VGND_c_422_n 0.00233634f $X=1.44 $Y=0.74 $X2=0 $Y2=0
cc_153 N_A2_M1001_g N_VGND_c_424_n 0.00383152f $X=0.995 $Y=0.74 $X2=0 $Y2=0
cc_154 N_A2_M1011_g N_VGND_c_424_n 0.00451267f $X=1.44 $Y=0.74 $X2=0 $Y2=0
cc_155 N_A2_M1001_g N_VGND_c_426_n 0.00757689f $X=0.995 $Y=0.74 $X2=0 $Y2=0
cc_156 N_A2_M1011_g N_VGND_c_426_n 0.00875489f $X=1.44 $Y=0.74 $X2=0 $Y2=0
cc_157 N_B1_c_194_n N_VPWR_c_242_n 0.00716461f $X=2.405 $Y=1.765 $X2=0 $Y2=0
cc_158 N_B1_c_196_n N_VPWR_c_242_n 4.42881e-19 $X=2.855 $Y=1.765 $X2=0 $Y2=0
cc_159 N_B1_c_196_n N_VPWR_c_244_n 0.010561f $X=2.855 $Y=1.765 $X2=0 $Y2=0
cc_160 B1 N_VPWR_c_244_n 0.0143742f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_161 N_B1_c_194_n N_VPWR_c_246_n 0.00413917f $X=2.405 $Y=1.765 $X2=0 $Y2=0
cc_162 N_B1_c_196_n N_VPWR_c_246_n 0.00445602f $X=2.855 $Y=1.765 $X2=0 $Y2=0
cc_163 N_B1_c_194_n N_VPWR_c_239_n 0.00817726f $X=2.405 $Y=1.765 $X2=0 $Y2=0
cc_164 N_B1_c_196_n N_VPWR_c_239_n 0.00861084f $X=2.855 $Y=1.765 $X2=0 $Y2=0
cc_165 N_B1_c_194_n N_Y_c_325_n 0.0169719f $X=2.405 $Y=1.765 $X2=0 $Y2=0
cc_166 N_B1_M1000_g N_Y_c_319_n 3.52947e-19 $X=2.4 $Y=0.74 $X2=0 $Y2=0
cc_167 N_B1_c_197_n N_Y_c_319_n 0.00177298f $X=2.865 $Y=1.22 $X2=0 $Y2=0
cc_168 N_B1_c_195_n Y 0.00137454f $X=2.765 $Y=1.492 $X2=0 $Y2=0
cc_169 N_B1_c_196_n Y 0.00319333f $X=2.855 $Y=1.765 $X2=0 $Y2=0
cc_170 N_B1_c_194_n Y 2.68607e-19 $X=2.405 $Y=1.765 $X2=0 $Y2=0
cc_171 N_B1_c_196_n Y 0.00799488f $X=2.855 $Y=1.765 $X2=0 $Y2=0
cc_172 N_B1_c_196_n Y 0.00383175f $X=2.855 $Y=1.765 $X2=0 $Y2=0
cc_173 N_B1_M1000_g N_Y_c_320_n 0.00491952f $X=2.4 $Y=0.74 $X2=0 $Y2=0
cc_174 N_B1_c_194_n N_Y_c_320_n 0.00208883f $X=2.405 $Y=1.765 $X2=0 $Y2=0
cc_175 N_B1_c_195_n N_Y_c_320_n 0.021036f $X=2.765 $Y=1.492 $X2=0 $Y2=0
cc_176 N_B1_c_196_n N_Y_c_320_n 0.00699998f $X=2.855 $Y=1.765 $X2=0 $Y2=0
cc_177 B1 N_Y_c_320_n 0.0275294f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_178 N_B1_M1000_g N_A_27_74#_c_365_n 7.03414e-19 $X=2.4 $Y=0.74 $X2=0 $Y2=0
cc_179 N_B1_M1000_g N_A_27_74#_c_367_n 0.0128435f $X=2.4 $Y=0.74 $X2=0 $Y2=0
cc_180 N_B1_c_197_n N_A_27_74#_c_367_n 0.0107617f $X=2.865 $Y=1.22 $X2=0 $Y2=0
cc_181 N_B1_M1000_g N_A_27_74#_c_369_n 6.09607e-19 $X=2.4 $Y=0.74 $X2=0 $Y2=0
cc_182 N_B1_c_196_n N_A_27_74#_c_369_n 0.00191466f $X=2.855 $Y=1.765 $X2=0 $Y2=0
cc_183 N_B1_c_197_n N_A_27_74#_c_369_n 0.00847698f $X=2.865 $Y=1.22 $X2=0 $Y2=0
cc_184 B1 N_A_27_74#_c_369_n 0.0251165f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_185 N_B1_M1000_g N_VGND_c_422_n 5.93944e-19 $X=2.4 $Y=0.74 $X2=0 $Y2=0
cc_186 N_B1_M1000_g N_VGND_c_425_n 0.00291649f $X=2.4 $Y=0.74 $X2=0 $Y2=0
cc_187 N_B1_c_197_n N_VGND_c_425_n 0.00291626f $X=2.865 $Y=1.22 $X2=0 $Y2=0
cc_188 N_B1_M1000_g N_VGND_c_426_n 0.00359962f $X=2.4 $Y=0.74 $X2=0 $Y2=0
cc_189 N_B1_c_197_n N_VGND_c_426_n 0.00363101f $X=2.865 $Y=1.22 $X2=0 $Y2=0
cc_190 N_VPWR_c_241_n N_A_116_368#_c_294_n 0.0412035f $X=0.28 $Y=2.455 $X2=0
+ $Y2=0
cc_191 N_VPWR_c_245_n N_A_116_368#_c_288_n 0.0423044f $X=2.095 $Y=3.33 $X2=0
+ $Y2=0
cc_192 N_VPWR_c_239_n N_A_116_368#_c_288_n 0.0238902f $X=3.12 $Y=3.33 $X2=0
+ $Y2=0
cc_193 N_VPWR_c_241_n N_A_116_368#_c_289_n 0.012272f $X=0.28 $Y=2.455 $X2=0
+ $Y2=0
cc_194 N_VPWR_c_245_n N_A_116_368#_c_289_n 0.0235512f $X=2.095 $Y=3.33 $X2=0
+ $Y2=0
cc_195 N_VPWR_c_239_n N_A_116_368#_c_289_n 0.0126924f $X=3.12 $Y=3.33 $X2=0
+ $Y2=0
cc_196 N_VPWR_c_242_n N_A_116_368#_c_290_n 0.0300075f $X=2.18 $Y=2.805 $X2=0
+ $Y2=0
cc_197 N_VPWR_c_245_n N_A_116_368#_c_290_n 0.0227333f $X=2.095 $Y=3.33 $X2=0
+ $Y2=0
cc_198 N_VPWR_c_239_n N_A_116_368#_c_290_n 0.0125508f $X=3.12 $Y=3.33 $X2=0
+ $Y2=0
cc_199 N_VPWR_M1005_d N_Y_c_325_n 0.00420216f $X=2.03 $Y=1.84 $X2=0 $Y2=0
cc_200 N_VPWR_c_242_n N_Y_c_325_n 0.0154248f $X=2.18 $Y=2.805 $X2=0 $Y2=0
cc_201 N_VPWR_c_244_n Y 0.0310109f $X=3.08 $Y=1.985 $X2=0 $Y2=0
cc_202 N_VPWR_c_242_n Y 0.0127584f $X=2.18 $Y=2.805 $X2=0 $Y2=0
cc_203 N_VPWR_c_244_n Y 0.0464479f $X=3.08 $Y=1.985 $X2=0 $Y2=0
cc_204 N_VPWR_c_246_n Y 0.0119166f $X=2.995 $Y=3.33 $X2=0 $Y2=0
cc_205 N_VPWR_c_239_n Y 0.00983061f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_206 N_A_116_368#_c_288_n N_Y_M1003_d 0.00250873f $X=1.565 $Y=2.99 $X2=0 $Y2=0
cc_207 N_A_116_368#_M1004_s N_Y_c_325_n 0.00495191f $X=1.53 $Y=1.84 $X2=0 $Y2=0
cc_208 N_A_116_368#_c_288_n N_Y_c_325_n 0.00419805f $X=1.565 $Y=2.99 $X2=0 $Y2=0
cc_209 N_A_116_368#_c_290_n N_Y_c_325_n 0.0195451f $X=1.73 $Y=2.805 $X2=0 $Y2=0
cc_210 N_A_116_368#_c_288_n N_Y_c_327_n 0.0183575f $X=1.565 $Y=2.99 $X2=0 $Y2=0
cc_211 N_Y_c_319_n N_A_27_74#_c_365_n 0.00427071f $X=2.605 $Y=1.13 $X2=0 $Y2=0
cc_212 N_Y_c_320_n N_A_27_74#_c_365_n 0.00353683f $X=2.66 $Y=1.82 $X2=0 $Y2=0
cc_213 N_Y_M1000_d N_A_27_74#_c_367_n 0.00226551f $X=2.475 $Y=0.37 $X2=0 $Y2=0
cc_214 N_Y_c_360_p N_A_27_74#_c_367_n 0.0138835f $X=2.645 $Y=0.88 $X2=0 $Y2=0
cc_215 N_A_27_74#_c_362_n N_VGND_M1009_s 0.00256964f $X=1.125 $Y=1.095 $X2=-0.19
+ $Y2=-0.245
cc_216 N_A_27_74#_c_365_n N_VGND_M1011_s 0.00240632f $X=2.055 $Y=1.095 $X2=0
+ $Y2=0
cc_217 N_A_27_74#_c_361_n N_VGND_c_421_n 0.0188012f $X=0.28 $Y=0.515 $X2=0 $Y2=0
cc_218 N_A_27_74#_c_362_n N_VGND_c_421_n 0.0201026f $X=1.125 $Y=1.095 $X2=0
+ $Y2=0
cc_219 N_A_27_74#_c_364_n N_VGND_c_421_n 0.0179318f $X=1.21 $Y=0.515 $X2=0 $Y2=0
cc_220 N_A_27_74#_c_364_n N_VGND_c_422_n 0.018051f $X=1.21 $Y=0.515 $X2=0 $Y2=0
cc_221 N_A_27_74#_c_365_n N_VGND_c_422_n 0.0189333f $X=2.055 $Y=1.095 $X2=0
+ $Y2=0
cc_222 N_A_27_74#_c_366_n N_VGND_c_422_n 0.00697079f $X=2.18 $Y=0.52 $X2=0 $Y2=0
cc_223 N_A_27_74#_c_361_n N_VGND_c_423_n 0.0145639f $X=0.28 $Y=0.515 $X2=0 $Y2=0
cc_224 N_A_27_74#_c_364_n N_VGND_c_424_n 0.0110391f $X=1.21 $Y=0.515 $X2=0 $Y2=0
cc_225 N_A_27_74#_c_366_n N_VGND_c_425_n 0.0111552f $X=2.18 $Y=0.52 $X2=0 $Y2=0
cc_226 N_A_27_74#_c_367_n N_VGND_c_425_n 0.0239026f $X=2.915 $Y=0.435 $X2=0
+ $Y2=0
cc_227 N_A_27_74#_c_369_n N_VGND_c_425_n 0.0146186f $X=3.08 $Y=0.515 $X2=0 $Y2=0
cc_228 N_A_27_74#_c_361_n N_VGND_c_426_n 0.0119984f $X=0.28 $Y=0.515 $X2=0 $Y2=0
cc_229 N_A_27_74#_c_364_n N_VGND_c_426_n 0.00911606f $X=1.21 $Y=0.515 $X2=0
+ $Y2=0
cc_230 N_A_27_74#_c_366_n N_VGND_c_426_n 0.00923333f $X=2.18 $Y=0.52 $X2=0 $Y2=0
cc_231 N_A_27_74#_c_367_n N_VGND_c_426_n 0.02025f $X=2.915 $Y=0.435 $X2=0 $Y2=0
cc_232 N_A_27_74#_c_369_n N_VGND_c_426_n 0.0120551f $X=3.08 $Y=0.515 $X2=0 $Y2=0
