* File: sky130_fd_sc_hs__mux2_1.spice
* Created: Thu Aug 27 20:48:45 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hs__mux2_1.pex.spice"
.subckt sky130_fd_sc_hs__mux2_1  VNB VPB S A1 A0 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A0	A0
* A1	A1
* S	S
* VPB	VPB
* VNB	VNB
MM1003 N_VGND_M1003_d N_S_M1003_g N_A_27_112#_M1003_s VNB NLOWVT L=0.15 W=0.55
+ AD=0.123281 AS=0.15675 PD=0.98062 PS=1.67 NRD=13.632 NRS=0 M=1 R=3.66667
+ SA=75000.2 SB=75003.5 A=0.0825 P=1.4 MULT=1
MM1006 A_226_74# N_S_M1006_g N_VGND_M1003_d VNB NLOWVT L=0.15 W=0.74 AD=0.0888
+ AS=0.165869 PD=0.98 PS=1.31938 NRD=10.536 NRS=11.34 M=1 R=4.93333 SA=75000.6
+ SB=75003 A=0.111 P=1.78 MULT=1
MM1004 N_A_304_74#_M1004_d N_A1_M1004_g A_226_74# VNB NLOWVT L=0.15 W=0.74
+ AD=0.20165 AS=0.0888 PD=1.285 PS=0.98 NRD=21.072 NRS=10.536 M=1 R=4.93333
+ SA=75001 SB=75002.6 A=0.111 P=1.78 MULT=1
MM1001 A_443_74# N_A0_M1001_g N_A_304_74#_M1004_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.2997 AS=0.20165 PD=1.55 PS=1.285 NRD=56.748 NRS=21.888 M=1 R=4.93333
+ SA=75001.7 SB=75001.9 A=0.111 P=1.78 MULT=1
MM1008 N_VGND_M1008_d N_A_27_112#_M1008_g A_443_74# VNB NLOWVT L=0.15 W=0.74
+ AD=0.20905 AS=0.2997 PD=1.305 PS=1.55 NRD=23.508 NRS=56.748 M=1 R=4.93333
+ SA=75002.7 SB=75000.9 A=0.111 P=1.78 MULT=1
MM1009 N_X_M1009_d N_A_304_74#_M1009_g N_VGND_M1008_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.20905 PD=2.05 PS=1.305 NRD=0 NRS=22.692 M=1 R=4.93333
+ SA=75003.4 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1005 N_VPWR_M1005_d N_S_M1005_g N_A_27_112#_M1005_s VPB PSHORT L=0.15 W=0.84
+ AD=0.169187 AS=0.2478 PD=1.26457 PS=2.27 NRD=22.261 NRS=2.3443 M=1 R=5.6
+ SA=75000.2 SB=75003.4 A=0.126 P=1.98 MULT=1
MM1000 A_223_368# N_S_M1000_g N_VPWR_M1005_d VPB PSHORT L=0.15 W=1 AD=0.4075
+ AS=0.201413 PD=1.815 PS=1.50543 NRD=69.4228 NRS=1.9503 M=1 R=6.66667
+ SA=75000.7 SB=75002.9 A=0.15 P=2.3 MULT=1
MM1002 N_A_304_74#_M1002_d N_A0_M1002_g A_223_368# VPB PSHORT L=0.15 W=1
+ AD=0.195 AS=0.4075 PD=1.39 PS=1.815 NRD=1.9503 NRS=69.4228 M=1 R=6.66667
+ SA=75001.6 SB=75001.9 A=0.15 P=2.3 MULT=1
MM1011 A_524_368# N_A1_M1011_g N_A_304_74#_M1002_d VPB PSHORT L=0.15 W=1 AD=0.21
+ AS=0.195 PD=1.42 PS=1.39 NRD=30.5153 NRS=19.7 M=1 R=6.66667 SA=75002.2
+ SB=75001.4 A=0.15 P=2.3 MULT=1
MM1007 N_VPWR_M1007_d N_A_27_112#_M1007_g A_524_368# VPB PSHORT L=0.15 W=1
+ AD=0.241226 AS=0.21 PD=1.5 PS=1.42 NRD=25.9252 NRS=30.5153 M=1 R=6.66667
+ SA=75002.7 SB=75000.8 A=0.15 P=2.3 MULT=1
MM1010 N_X_M1010_d N_A_304_74#_M1010_g N_VPWR_M1007_d VPB PSHORT L=0.15 W=1.12
+ AD=0.3304 AS=0.270174 PD=2.83 PS=1.68 NRD=1.7533 NRS=10.5395 M=1 R=7.46667
+ SA=75003 SB=75000.2 A=0.168 P=2.54 MULT=1
DX12_noxref VNB VPB NWDIODE A=8.742 P=13.12
*
.include "sky130_fd_sc_hs__mux2_1.pxi.spice"
*
.ends
*
*
