* File: sky130_fd_sc_hs__mux2_4.spice
* Created: Thu Aug 27 20:49:00 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hs__mux2_4.pex.spice"
.subckt sky130_fd_sc_hs__mux2_4  VNB VPB S A0 A1 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A1	A1
* A0	A0
* S	S
* VPB	VPB
* VNB	VNB
MM1003 N_VGND_M1003_d N_S_M1003_g N_A_27_368#_M1003_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.136255 AS=0.1824 PD=1.07594 PS=1.85 NRD=13.116 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75004.4 A=0.096 P=1.58 MULT=1
MM1009 N_X_M1009_d N_A_193_241#_M1009_g N_VGND_M1003_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.1184 AS=0.157545 PD=1.06 PS=1.24406 NRD=6.48 NRS=11.34 M=1 R=4.93333
+ SA=75000.7 SB=75003.5 A=0.111 P=1.78 MULT=1
MM1014 N_X_M1009_d N_A_193_241#_M1014_g N_VGND_M1014_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1184 AS=0.1628 PD=1.06 PS=1.18 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75001.2
+ SB=75003.1 A=0.111 P=1.78 MULT=1
MM1021 N_X_M1021_d N_A_193_241#_M1021_g N_VGND_M1014_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1628 PD=1.02 PS=1.18 NRD=0 NRS=14.592 M=1 R=4.93333 SA=75001.8
+ SB=75002.5 A=0.111 P=1.78 MULT=1
MM1023 N_X_M1021_d N_A_193_241#_M1023_g N_VGND_M1023_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.249804 PD=1.02 PS=1.56043 NRD=0 NRS=27.156 M=1 R=4.93333
+ SA=75002.2 SB=75002.1 A=0.111 P=1.78 MULT=1
MM1001 N_A_709_119#_M1001_d N_S_M1001_g N_VGND_M1023_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.112 AS=0.216046 PD=0.99 PS=1.34957 NRD=0 NRS=73.116 M=1 R=4.26667
+ SA=75002.6 SB=75001.9 A=0.096 P=1.58 MULT=1
MM1024 N_A_709_119#_M1001_d N_S_M1024_g N_VGND_M1024_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.112 AS=0.1568 PD=0.99 PS=1.13 NRD=13.116 NRS=13.116 M=1 R=4.26667
+ SA=75003.1 SB=75001.4 A=0.096 P=1.58 MULT=1
MM1005 N_A_937_119#_M1005_d N_A_27_368#_M1005_g N_VGND_M1024_s VNB NLOWVT L=0.15
+ W=0.64 AD=0.0896 AS=0.1568 PD=0.92 PS=1.13 NRD=0 NRS=26.244 M=1 R=4.26667
+ SA=75003.7 SB=75000.8 A=0.096 P=1.58 MULT=1
MM1010 N_A_937_119#_M1005_d N_A_27_368#_M1010_g N_VGND_M1010_s VNB NLOWVT L=0.15
+ W=0.64 AD=0.0896 AS=0.3692 PD=0.92 PS=2.64 NRD=0 NRS=97.848 M=1 R=4.26667
+ SA=75004.2 SB=75000.4 A=0.096 P=1.58 MULT=1
MM1017 N_A_937_119#_M1017_d N_A0_M1017_g N_A_193_241#_M1017_s VNB NLOWVT L=0.15
+ W=0.64 AD=0.096 AS=0.4992 PD=0.94 PS=2.84 NRD=0 NRS=13.116 M=1 R=4.26667
+ SA=75000.7 SB=75001.6 A=0.096 P=1.58 MULT=1
MM1022 N_A_937_119#_M1017_d N_A0_M1022_g N_A_193_241#_M1022_s VNB NLOWVT L=0.15
+ W=0.64 AD=0.096 AS=0.1056 PD=0.94 PS=0.97 NRD=3.744 NRS=9.372 M=1 R=4.26667
+ SA=75001.2 SB=75001.2 A=0.096 P=1.58 MULT=1
MM1015 N_A_193_241#_M1022_s N_A1_M1015_g N_A_709_119#_M1015_s VNB NLOWVT L=0.15
+ W=0.64 AD=0.1056 AS=0.0992 PD=0.97 PS=0.95 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75001.6 SB=75000.7 A=0.096 P=1.58 MULT=1
MM1025 N_A_193_241#_M1025_d N_A1_M1025_g N_A_709_119#_M1015_s VNB NLOWVT L=0.15
+ W=0.64 AD=0.2112 AS=0.0992 PD=1.94 PS=0.95 NRD=7.488 NRS=5.616 M=1 R=4.26667
+ SA=75002.1 SB=75000.3 A=0.096 P=1.58 MULT=1
MM1016 N_VPWR_M1016_d N_S_M1016_g N_A_27_368#_M1016_s VPB PSHORT L=0.15 W=1
+ AD=0.206226 AS=0.295 PD=1.43396 PS=2.59 NRD=20.6653 NRS=1.9503 M=1 R=6.66667
+ SA=75000.2 SB=75004.6 A=0.15 P=2.3 MULT=1
MM1006 N_VPWR_M1016_d N_A_193_241#_M1006_g N_X_M1006_s VPB PSHORT L=0.15 W=1.12
+ AD=0.230974 AS=0.29075 PD=1.60604 PS=1.78 NRD=0 NRS=35.9722 M=1 R=7.46667
+ SA=75000.7 SB=75004.1 A=0.168 P=2.54 MULT=1
MM1011 N_VPWR_M1011_d N_A_193_241#_M1011_g N_X_M1006_s VPB PSHORT L=0.15 W=1.12
+ AD=0.290025 AS=0.29075 PD=1.775 PS=1.78 NRD=17.5724 NRS=17.5724 M=1 R=7.46667
+ SA=75001.3 SB=75003.4 A=0.168 P=2.54 MULT=1
MM1012 N_VPWR_M1011_d N_A_193_241#_M1012_g N_X_M1012_s VPB PSHORT L=0.15 W=1.12
+ AD=0.290025 AS=0.275525 PD=1.775 PS=1.675 NRD=35.854 NRS=3.94 M=1 R=7.46667
+ SA=75002 SB=75002.8 A=0.168 P=2.54 MULT=1
MM1013 N_VPWR_M1013_d N_A_193_241#_M1013_g N_X_M1012_s VPB PSHORT L=0.15 W=1.12
+ AD=0.293749 AS=0.275525 PD=1.87547 PS=1.675 NRD=36.445 NRS=3.94 M=1 R=7.46667
+ SA=75002.6 SB=75002.2 A=0.168 P=2.54 MULT=1
MM1002 N_A_722_391#_M1002_d N_S_M1002_g N_VPWR_M1013_d VPB PSHORT L=0.15 W=1
+ AD=0.15 AS=0.262276 PD=1.3 PS=1.67453 NRD=0 NRS=40.8184 M=1 R=6.66667
+ SA=75003.2 SB=75001.8 A=0.15 P=2.3 MULT=1
MM1007 N_A_722_391#_M1002_d N_S_M1007_g N_VPWR_M1007_s VPB PSHORT L=0.15 W=1
+ AD=0.15 AS=0.25385 PD=1.3 PS=1.6 NRD=1.9503 NRS=19.6803 M=1 R=6.66667
+ SA=75003.6 SB=75001.4 A=0.15 P=2.3 MULT=1
MM1000 N_VPWR_M1007_s N_A_27_368#_M1000_g N_A_936_391#_M1000_s VPB PSHORT L=0.15
+ W=1 AD=0.25385 AS=0.15 PD=1.6 PS=1.3 NRD=19.6803 NRS=1.9503 M=1 R=6.66667
+ SA=75004.3 SB=75000.8 A=0.15 P=2.3 MULT=1
MM1020 N_VPWR_M1020_d N_A_27_368#_M1020_g N_A_936_391#_M1000_s VPB PSHORT L=0.15
+ W=1 AD=0.4177 AS=0.15 PD=3.02 PS=1.3 NRD=19.6803 NRS=1.9503 M=1 R=6.66667
+ SA=75004.7 SB=75000.3 A=0.15 P=2.3 MULT=1
MM1004 N_A_722_391#_M1004_d N_A0_M1004_g N_A_193_241#_M1004_s VPB PSHORT L=0.15
+ W=1 AD=0.15 AS=0.33 PD=1.3 PS=2.66 NRD=1.9503 NRS=5.8903 M=1 R=6.66667
+ SA=75000.3 SB=75001.6 A=0.15 P=2.3 MULT=1
MM1008 N_A_722_391#_M1004_d N_A0_M1008_g N_A_193_241#_M1008_s VPB PSHORT L=0.15
+ W=1 AD=0.15 AS=0.155 PD=1.3 PS=1.31 NRD=1.9503 NRS=2.9353 M=1 R=6.66667
+ SA=75000.7 SB=75001.2 A=0.15 P=2.3 MULT=1
MM1018 N_A_936_391#_M1018_d N_A1_M1018_g N_A_193_241#_M1008_s VPB PSHORT L=0.15
+ W=1 AD=0.15 AS=0.155 PD=1.3 PS=1.31 NRD=1.9503 NRS=2.9353 M=1 R=6.66667
+ SA=75001.2 SB=75000.7 A=0.15 P=2.3 MULT=1
MM1019 N_A_936_391#_M1018_d N_A1_M1019_g N_A_193_241#_M1019_s VPB PSHORT L=0.15
+ W=1 AD=0.15 AS=0.345 PD=1.3 PS=2.69 NRD=1.9503 NRS=11.8003 M=1 R=6.66667
+ SA=75001.6 SB=75000.3 A=0.15 P=2.3 MULT=1
DX26_noxref VNB VPB NWDIODE A=17.0422 P=22.14
*
.include "sky130_fd_sc_hs__mux2_4.pxi.spice"
*
.ends
*
*
