* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hs__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
X0 a_817_138# a_837_359# a_895_138# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X1 a_696_457# a_306_74# a_786_457# VPB sky130_fd_pr__pfet_01v8 w=420000u l=150000u
X2 a_1271_74# a_490_362# a_1478_493# VPB sky130_fd_pr__pfet_01v8 w=420000u l=150000u
X3 a_30_78# a_306_74# a_696_457# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X4 a_1481_81# a_1525_212# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X5 a_306_74# CLK VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X6 VGND a_1271_74# a_1921_409# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X7 VPWR D a_30_78# VPB sky130_fd_pr__pfet_01v8 w=420000u l=150000u
X8 a_306_74# CLK VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X9 a_696_457# a_490_362# a_817_138# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X10 a_1525_212# a_1271_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=420000u l=150000u
X11 VGND a_696_457# a_837_359# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X12 Q a_1921_409# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X13 a_30_78# a_490_362# a_696_457# VPB sky130_fd_pr__pfet_01v8 w=420000u l=150000u
X14 VPWR RESET_B a_696_457# VPB sky130_fd_pr__pfet_01v8 w=420000u l=150000u
X15 Q a_1921_409# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X16 a_895_138# RESET_B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X17 VGND a_1921_409# Q VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X18 VPWR a_696_457# a_837_359# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=150000u
X19 VGND a_306_74# a_490_362# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X20 a_1271_74# a_306_74# a_1481_81# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X21 a_786_457# a_837_359# VPWR VPB sky130_fd_pr__pfet_01v8 w=420000u l=150000u
X22 a_1478_493# a_1525_212# VPWR VPB sky130_fd_pr__pfet_01v8 w=420000u l=150000u
X23 a_837_359# a_306_74# a_1271_74# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=150000u
X24 a_117_78# RESET_B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X25 VPWR a_1271_74# a_1921_409# VPB sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X26 a_1663_81# a_1271_74# a_1525_212# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X27 VPWR a_306_74# a_490_362# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X28 a_30_78# D a_117_78# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X29 a_837_359# a_490_362# a_1271_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X30 VGND RESET_B a_1663_81# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X31 VPWR RESET_B a_1525_212# VPB sky130_fd_pr__pfet_01v8 w=420000u l=150000u
X32 VPWR a_1921_409# Q VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X33 a_30_78# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8 w=420000u l=150000u
.ends
