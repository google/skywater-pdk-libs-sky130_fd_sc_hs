# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_hs__or4b_1
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_hs__or4b_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.320000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.232500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.995000 1.350000 3.325000 1.780000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.232500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.455000 1.180000 2.785000 1.780000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.232500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.885000 1.045000 2.275000 1.780000 ;
    END
  END C
  PIN D_N
    ANTENNAGATEAREA  0.208500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.450000 0.570000 1.780000 ;
    END
  END D_N
  PIN X
    ANTENNADIFFAREA  0.541300 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.835000 0.350000 4.235000 1.130000 ;
        RECT 3.835000 1.820000 4.235000 2.980000 ;
        RECT 4.065000 1.130000 4.235000 1.820000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 4.320000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 4.320000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.320000 0.085000 ;
      RECT 0.000000  3.245000 4.320000 3.415000 ;
      RECT 0.115000  0.350000 0.445000 1.110000 ;
      RECT 0.115000  1.110000 0.980000 1.280000 ;
      RECT 0.120000  1.950000 0.980000 2.120000 ;
      RECT 0.120000  2.120000 0.450000 2.980000 ;
      RECT 0.615000  0.085000 0.945000 0.940000 ;
      RECT 0.620000  2.290000 0.950000 3.245000 ;
      RECT 0.810000  1.280000 0.980000 1.580000 ;
      RECT 0.810000  1.580000 1.140000 1.910000 ;
      RECT 0.810000  1.910000 0.980000 1.950000 ;
      RECT 1.115000  0.545000 2.090000 0.875000 ;
      RECT 1.315000  0.875000 1.645000 1.950000 ;
      RECT 1.315000  1.950000 3.665000 2.120000 ;
      RECT 1.315000  2.120000 1.645000 2.860000 ;
      RECT 2.260000  0.085000 2.590000 0.875000 ;
      RECT 2.760000  0.350000 3.125000 0.940000 ;
      RECT 2.955000  0.940000 3.125000 1.010000 ;
      RECT 2.955000  1.010000 3.665000 1.180000 ;
      RECT 3.295000  0.085000 3.625000 0.840000 ;
      RECT 3.335000  2.290000 3.665000 3.245000 ;
      RECT 3.495000  1.180000 3.665000 1.300000 ;
      RECT 3.495000  1.300000 3.895000 1.630000 ;
      RECT 3.495000  1.630000 3.665000 1.950000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
  END
END sky130_fd_sc_hs__or4b_1
