* File: sky130_fd_sc_hs__o22a_1.pex.spice
* Created: Thu Aug 27 21:00:00 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HS__O22A_1%A_83_260# 1 2 9 11 13 15 16 21 24 26 30 34 35
+ 40
c78 35 0 1.80886e-19 $X=2.26 $Y=1.202
c79 30 0 4.2886e-20 $X=0.93 $Y=1.465
c80 21 0 1.97013e-19 $X=2.26 $Y=1.97
c81 11 0 1.53455e-19 $X=0.505 $Y=1.765
r82 37 40 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=2.26 $Y=2.055 $X2=2.56
+ $Y2=2.055
r83 33 35 9.669 $w=1.93e-07 $l=1.7e-07 $layer=LI1_cond $X=2.09 $Y=1.202 $X2=2.26
+ $Y2=1.202
r84 33 34 10.7338 $w=1.93e-07 $l=1.85e-07 $layer=LI1_cond $X=2.09 $Y=1.202
+ $X2=1.905 $Y2=1.202
r85 24 40 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=2.56 $Y=2.815
+ $X2=2.56 $Y2=2.14
r86 21 37 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.26 $Y=1.97
+ $X2=2.26 $Y2=2.055
r87 20 35 1.54022 $w=1.7e-07 $l=9.8e-08 $layer=LI1_cond $X=2.26 $Y=1.3 $X2=2.26
+ $Y2=1.202
r88 20 21 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.26 $Y=1.3 $X2=2.26
+ $Y2=1.97
r89 19 26 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.095 $Y=1.215
+ $X2=1.01 $Y2=1.215
r90 19 34 52.8449 $w=1.68e-07 $l=8.1e-07 $layer=LI1_cond $X=1.095 $Y=1.215
+ $X2=1.905 $Y2=1.215
r91 16 30 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.93
+ $Y=1.465 $X2=0.93 $Y2=1.465
r92 16 26 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=1.01 $Y=1.465
+ $X2=1.01 $Y2=1.215
r93 14 30 58.5785 $w=3.3e-07 $l=3.35e-07 $layer=POLY_cond $X=0.595 $Y=1.465
+ $X2=0.93 $Y2=1.465
r94 14 15 5.03009 $w=3.3e-07 $l=1.1887e-07 $layer=POLY_cond $X=0.595 $Y=1.465
+ $X2=0.505 $Y2=1.532
r95 11 15 37.0704 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=0.505 $Y=1.765
+ $X2=0.505 $Y2=1.532
r96 11 13 204.047 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.505 $Y=1.765
+ $X2=0.505 $Y2=2.4
r97 7 15 37.0704 $w=1.5e-07 $l=2.36947e-07 $layer=POLY_cond $X=0.495 $Y=1.3
+ $X2=0.505 $Y2=1.532
r98 7 9 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=0.495 $Y=1.3 $X2=0.495
+ $Y2=0.74
r99 2 40 400 $w=1.7e-07 $l=2.38485e-07 $layer=licon1_PDIFF $count=1 $X=2.41
+ $Y=1.96 $X2=2.56 $Y2=2.135
r100 2 24 400 $w=1.7e-07 $l=9.26971e-07 $layer=licon1_PDIFF $count=1 $X=2.41
+ $Y=1.96 $X2=2.56 $Y2=2.815
r101 1 33 182 $w=1.7e-07 $l=5.69408e-07 $layer=licon1_NDIFF $count=1 $X=1.93
+ $Y=0.695 $X2=2.09 $Y2=1.19
.ends

.subckt PM_SKY130_FD_SC_HS__O22A_1%B1 1 5 7 9 10 14
r38 10 14 0.535558 $w=6.68e-07 $l=3e-08 $layer=LI1_cond $X=1.67 $Y=1.665
+ $X2=1.67 $Y2=1.635
r39 7 9 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=1.915 $Y=1.885
+ $X2=1.915 $Y2=2.46
r40 3 5 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=1.855 $Y=1.47
+ $X2=1.855 $Y2=1.015
r41 1 7 60.5037 $w=2.15e-07 $l=2.61247e-07 $layer=POLY_cond $X=1.892 $Y=1.635
+ $X2=1.915 $Y2=1.885
r42 1 14 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.84
+ $Y=1.635 $X2=1.84 $Y2=1.635
r43 1 3 41.4478 $w=2.15e-07 $l=1.82565e-07 $layer=POLY_cond $X=1.892 $Y=1.635
+ $X2=1.855 $Y2=1.47
.ends

.subckt PM_SKY130_FD_SC_HS__O22A_1%B2 1 2 6 7 9 13 14 16 24
c48 24 0 4.2886e-20 $X=1.305 $Y=0.462
c49 13 0 6.69395e-20 $X=2.305 $Y=0.42
r50 16 24 3.43205 $w=4.13e-07 $l=1.05e-07 $layer=LI1_cond $X=1.2 $Y=0.462
+ $X2=1.305 $Y2=0.462
r51 14 20 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.305 $Y=0.42
+ $X2=2.305 $Y2=0.585
r52 13 24 34.9225 $w=3.28e-07 $l=1e-06 $layer=LI1_cond $X=2.305 $Y=0.42
+ $X2=1.305 $Y2=0.42
r53 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.305
+ $Y=0.42 $X2=2.305 $Y2=0.42
r54 7 9 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=2.335 $Y=1.885
+ $X2=2.335 $Y2=2.46
r55 6 10 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=2.325 $Y=1.015
+ $X2=2.325 $Y2=1.41
r56 6 20 220.489 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=2.325 $Y=1.015
+ $X2=2.325 $Y2=0.585
r57 2 7 36.0588 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=2.335 $Y=1.795 $X2=2.335
+ $Y2=1.885
r58 1 10 36.5962 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=2.335 $Y=1.5 $X2=2.335
+ $Y2=1.41
r59 1 2 114.669 $w=1.8e-07 $l=2.95e-07 $layer=POLY_cond $X=2.335 $Y=1.5
+ $X2=2.335 $Y2=1.795
.ends

.subckt PM_SKY130_FD_SC_HS__O22A_1%A2 3 5 7 8 12
c37 3 0 2.47825e-19 $X=2.755 $Y=1.015
r38 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.83
+ $Y=1.635 $X2=2.83 $Y2=1.635
r39 8 12 6.63528 $w=3.28e-07 $l=1.9e-07 $layer=LI1_cond $X=2.64 $Y=1.635
+ $X2=2.83 $Y2=1.635
r40 5 11 52.2586 $w=2.99e-07 $l=2.7157e-07 $layer=POLY_cond $X=2.785 $Y=1.885
+ $X2=2.83 $Y2=1.635
r41 5 7 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=2.785 $Y=1.885
+ $X2=2.785 $Y2=2.46
r42 1 11 38.5562 $w=2.99e-07 $l=1.98997e-07 $layer=POLY_cond $X=2.755 $Y=1.47
+ $X2=2.83 $Y2=1.635
r43 1 3 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=2.755 $Y=1.47
+ $X2=2.755 $Y2=1.015
.ends

.subckt PM_SKY130_FD_SC_HS__O22A_1%A1 1 3 6 8
r24 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.4
+ $Y=1.635 $X2=3.4 $Y2=1.635
r25 8 12 6.9845 $w=3.28e-07 $l=2e-07 $layer=LI1_cond $X=3.6 $Y=1.635 $X2=3.4
+ $Y2=1.635
r26 4 11 38.5562 $w=2.99e-07 $l=1.90526e-07 $layer=POLY_cond $X=3.345 $Y=1.47
+ $X2=3.4 $Y2=1.635
r27 4 6 256.383 $w=1.5e-07 $l=5e-07 $layer=POLY_cond $X=3.345 $Y=1.47 $X2=3.345
+ $Y2=0.97
r28 1 11 52.2586 $w=2.99e-07 $l=2.85044e-07 $layer=POLY_cond $X=3.325 $Y=1.885
+ $X2=3.4 $Y2=1.635
r29 1 3 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=3.325 $Y=1.885
+ $X2=3.325 $Y2=2.46
.ends

.subckt PM_SKY130_FD_SC_HS__O22A_1%X 1 2 9 13 14 15 16 23 32
c21 32 0 1.53455e-19 $X=0.265 $Y=1.82
r22 21 23 1.12043 $w=3.58e-07 $l=3.5e-08 $layer=LI1_cond $X=0.265 $Y=2 $X2=0.265
+ $Y2=2.035
r23 15 16 11.8446 $w=3.58e-07 $l=3.7e-07 $layer=LI1_cond $X=0.265 $Y=2.405
+ $X2=0.265 $Y2=2.775
r24 14 21 0.800308 $w=3.58e-07 $l=2.5e-08 $layer=LI1_cond $X=0.265 $Y=1.975
+ $X2=0.265 $Y2=2
r25 14 32 8.1909 $w=3.58e-07 $l=1.55e-07 $layer=LI1_cond $X=0.265 $Y=1.975
+ $X2=0.265 $Y2=1.82
r26 14 15 11.0442 $w=3.58e-07 $l=3.45e-07 $layer=LI1_cond $X=0.265 $Y=2.06
+ $X2=0.265 $Y2=2.405
r27 14 23 0.800308 $w=3.58e-07 $l=2.5e-08 $layer=LI1_cond $X=0.265 $Y=2.06
+ $X2=0.265 $Y2=2.035
r28 13 32 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=0.17 $Y=1.13 $X2=0.17
+ $Y2=1.82
r29 7 13 7.52792 $w=2.78e-07 $l=1.4e-07 $layer=LI1_cond $X=0.225 $Y=0.99
+ $X2=0.225 $Y2=1.13
r30 7 9 19.5504 $w=2.78e-07 $l=4.75e-07 $layer=LI1_cond $X=0.225 $Y=0.99
+ $X2=0.225 $Y2=0.515
r31 2 14 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=1.985
r32 2 16 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.815
r33 1 9 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__O22A_1%VPWR 1 2 9 16 18 22 24 29 38 44
r38 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r39 39 41 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=0.72 $Y2=3.33
r40 38 41 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r41 38 39 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r42 36 44 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=3.6 $Y2=3.33
r43 35 36 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r44 33 36 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=3.12 $Y2=3.33
r45 32 35 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=2.16 $Y=3.33 $X2=3.12
+ $Y2=3.33
r46 32 33 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r47 30 38 17.8809 $w=1.7e-07 $l=6.18e-07 $layer=LI1_cond $X=1.85 $Y=3.33
+ $X2=1.232 $Y2=3.33
r48 30 32 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=1.85 $Y=3.33
+ $X2=2.16 $Y2=3.33
r49 29 43 4.71369 $w=1.7e-07 $l=2.27e-07 $layer=LI1_cond $X=3.385 $Y=3.33
+ $X2=3.612 $Y2=3.33
r50 29 35 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=3.385 $Y=3.33
+ $X2=3.12 $Y2=3.33
r51 27 41 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r52 26 27 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r53 24 38 17.8809 $w=1.7e-07 $l=6.17e-07 $layer=LI1_cond $X=0.615 $Y=3.33
+ $X2=1.232 $Y2=3.33
r54 24 26 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=0.615 $Y=3.33
+ $X2=0.24 $Y2=3.33
r55 22 33 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=2.16 $Y2=3.33
r56 22 39 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=1.68 $Y2=3.33
r57 18 21 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=3.55 $Y=2.135
+ $X2=3.55 $Y2=2.815
r58 16 43 3.05248 $w=3.3e-07 $l=1.11781e-07 $layer=LI1_cond $X=3.55 $Y=3.245
+ $X2=3.612 $Y2=3.33
r59 16 21 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=3.55 $Y=3.245
+ $X2=3.55 $Y2=2.815
r60 12 15 3.3587 $w=1.233e-06 $l=3.4e-07 $layer=LI1_cond $X=1.232 $Y=2.49
+ $X2=1.232 $Y2=2.83
r61 9 12 3.3587 $w=1.233e-06 $l=3.4e-07 $layer=LI1_cond $X=1.232 $Y=2.15
+ $X2=1.232 $Y2=2.49
r62 7 38 3.84952 $w=1.235e-06 $l=8.5e-08 $layer=LI1_cond $X=1.232 $Y=3.245
+ $X2=1.232 $Y2=3.33
r63 7 15 4.0996 $w=1.233e-06 $l=4.15e-07 $layer=LI1_cond $X=1.232 $Y=3.245
+ $X2=1.232 $Y2=2.83
r64 2 21 400 $w=1.7e-07 $l=9.26971e-07 $layer=licon1_PDIFF $count=1 $X=3.4
+ $Y=1.96 $X2=3.55 $Y2=2.815
r65 2 18 400 $w=1.7e-07 $l=2.38485e-07 $layer=licon1_PDIFF $count=1 $X=3.4
+ $Y=1.96 $X2=3.55 $Y2=2.135
r66 1 15 266.667 $w=1.7e-07 $l=1.27615e-06 $layer=licon1_PDIFF $count=2 $X=0.58
+ $Y=1.84 $X2=1.235 $Y2=2.83
r67 1 12 266.667 $w=1.7e-07 $l=1.39258e-06 $layer=licon1_PDIFF $count=2 $X=0.58
+ $Y=1.84 $X2=1.685 $Y2=2.49
r68 1 12 266.667 $w=1.7e-07 $l=7.2336e-07 $layer=licon1_PDIFF $count=2 $X=0.58
+ $Y=1.84 $X2=0.735 $Y2=2.49
r69 1 9 266.667 $w=1.7e-07 $l=7.95031e-07 $layer=licon1_PDIFF $count=2 $X=0.58
+ $Y=1.84 $X2=1.235 $Y2=2.15
.ends

.subckt PM_SKY130_FD_SC_HS__O22A_1%VGND 1 2 9 13 15 17 22 32 33 36 39
r40 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r41 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r42 33 40 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=3.12
+ $Y2=0
r43 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r44 30 39 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=3.225 $Y=0 $X2=3.055
+ $Y2=0
r45 30 32 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=3.225 $Y=0 $X2=3.6
+ $Y2=0
r46 29 40 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r47 28 29 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r48 26 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r49 25 28 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.2 $Y=0 $X2=2.64
+ $Y2=0
r50 25 26 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r51 23 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.875 $Y=0 $X2=0.71
+ $Y2=0
r52 23 25 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.875 $Y=0 $X2=1.2
+ $Y2=0
r53 22 39 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=2.885 $Y=0 $X2=3.055
+ $Y2=0
r54 22 28 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=2.885 $Y=0 $X2=2.64
+ $Y2=0
r55 20 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r56 19 20 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r57 17 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.545 $Y=0 $X2=0.71
+ $Y2=0
r58 17 19 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.545 $Y=0 $X2=0.24
+ $Y2=0
r59 15 29 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=2.64
+ $Y2=0
r60 15 26 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=1.2
+ $Y2=0
r61 11 39 0.987631 $w=3.4e-07 $l=8.5e-08 $layer=LI1_cond $X=3.055 $Y=0.085
+ $X2=3.055 $Y2=0
r62 11 13 24.0657 $w=3.38e-07 $l=7.1e-07 $layer=LI1_cond $X=3.055 $Y=0.085
+ $X2=3.055 $Y2=0.795
r63 7 36 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.71 $Y=0.085 $X2=0.71
+ $Y2=0
r64 7 9 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=0.71 $Y=0.085 $X2=0.71
+ $Y2=0.515
r65 2 13 182 $w=1.7e-07 $l=2.70416e-07 $layer=licon1_NDIFF $count=1 $X=2.83
+ $Y=0.695 $X2=3.055 $Y2=0.795
r66 1 9 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=0.57
+ $Y=0.37 $X2=0.71 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HS__O22A_1%A_299_139# 1 2 3 10 14 15 16 17 20
r39 18 20 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=3.56 $Y=1.13
+ $X2=3.56 $Y2=0.795
r40 16 18 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.395 $Y=1.215
+ $X2=3.56 $Y2=1.13
r41 16 17 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=3.395 $Y=1.215
+ $X2=2.705 $Y2=1.215
r42 15 17 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.62 $Y=1.13
+ $X2=2.705 $Y2=1.215
r43 14 23 3.50935 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=2.62 $Y=0.935 $X2=2.62
+ $Y2=0.845
r44 14 15 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=2.62 $Y=0.935
+ $X2=2.62 $Y2=1.13
r45 10 23 3.31438 $w=1.8e-07 $l=8.5e-08 $layer=LI1_cond $X=2.535 $Y=0.845
+ $X2=2.62 $Y2=0.845
r46 10 12 55.1465 $w=1.78e-07 $l=8.95e-07 $layer=LI1_cond $X=2.535 $Y=0.845
+ $X2=1.64 $Y2=0.845
r47 3 20 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.42
+ $Y=0.65 $X2=3.56 $Y2=0.795
r48 2 23 182 $w=1.7e-07 $l=2.08567e-07 $layer=licon1_NDIFF $count=1 $X=2.4
+ $Y=0.695 $X2=2.54 $Y2=0.845
r49 1 12 182 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_NDIFF $count=1 $X=1.495
+ $Y=0.695 $X2=1.64 $Y2=0.845
.ends

