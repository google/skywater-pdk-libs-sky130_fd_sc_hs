* File: sky130_fd_sc_hs__o22a_4.pxi.spice
* Created: Thu Aug 27 21:00:16 2020
* 
x_PM_SKY130_FD_SC_HS__O22A_4%A2 N_A2_c_119_n N_A2_M1010_g N_A2_M1018_g
+ N_A2_c_116_n N_A2_M1019_g N_A2_c_120_n N_A2_M1011_g A2 N_A2_c_117_n
+ N_A2_c_118_n PM_SKY130_FD_SC_HS__O22A_4%A2
x_PM_SKY130_FD_SC_HS__O22A_4%A1 N_A1_c_172_n N_A1_c_173_n N_A1_M1020_g
+ N_A1_c_181_n N_A1_M1008_g N_A1_c_175_n N_A1_c_176_n N_A1_c_177_n N_A1_M1009_g
+ N_A1_M1021_g A1 PM_SKY130_FD_SC_HS__O22A_4%A1
x_PM_SKY130_FD_SC_HS__O22A_4%B2 N_B2_M1013_g N_B2_c_243_n N_B2_M1005_g
+ N_B2_c_240_n N_B2_M1017_g N_B2_c_244_n N_B2_M1006_g B2 B2 N_B2_c_241_n
+ N_B2_c_242_n PM_SKY130_FD_SC_HS__O22A_4%B2
x_PM_SKY130_FD_SC_HS__O22A_4%B1 N_B1_M1001_g N_B1_c_299_n N_B1_c_300_n
+ N_B1_c_308_n N_B1_M1002_g N_B1_c_301_n N_B1_M1023_g N_B1_c_303_n N_B1_c_310_n
+ N_B1_M1003_g N_B1_c_304_n B1 N_B1_c_306_n PM_SKY130_FD_SC_HS__O22A_4%B1
x_PM_SKY130_FD_SC_HS__O22A_4%A_206_392# N_A_206_392#_M1001_s
+ N_A_206_392#_M1017_d N_A_206_392#_M1010_d N_A_206_392#_M1005_d
+ N_A_206_392#_c_390_n N_A_206_392#_M1000_g N_A_206_392#_M1004_g
+ N_A_206_392#_c_391_n N_A_206_392#_M1012_g N_A_206_392#_M1007_g
+ N_A_206_392#_c_392_n N_A_206_392#_M1014_g N_A_206_392#_M1016_g
+ N_A_206_392#_c_393_n N_A_206_392#_M1015_g N_A_206_392#_M1022_g
+ N_A_206_392#_c_394_n N_A_206_392#_c_395_n N_A_206_392#_c_396_n
+ N_A_206_392#_c_383_n N_A_206_392#_c_384_n N_A_206_392#_c_385_n
+ N_A_206_392#_c_386_n N_A_206_392#_c_482_p N_A_206_392#_c_398_n
+ N_A_206_392#_c_399_n N_A_206_392#_c_411_n N_A_206_392#_c_387_n
+ N_A_206_392#_c_388_n N_A_206_392#_c_389_n
+ PM_SKY130_FD_SC_HS__O22A_4%A_206_392#
x_PM_SKY130_FD_SC_HS__O22A_4%VPWR N_VPWR_M1008_d N_VPWR_M1009_d N_VPWR_M1003_s
+ N_VPWR_M1012_d N_VPWR_M1015_d N_VPWR_c_556_n N_VPWR_c_557_n N_VPWR_c_558_n
+ N_VPWR_c_559_n N_VPWR_c_560_n N_VPWR_c_561_n N_VPWR_c_562_n N_VPWR_c_563_n
+ N_VPWR_c_564_n N_VPWR_c_565_n N_VPWR_c_566_n VPWR N_VPWR_c_567_n
+ N_VPWR_c_568_n N_VPWR_c_569_n N_VPWR_c_555_n PM_SKY130_FD_SC_HS__O22A_4%VPWR
x_PM_SKY130_FD_SC_HS__O22A_4%A_116_392# N_A_116_392#_M1008_s
+ N_A_116_392#_M1011_s N_A_116_392#_c_636_n N_A_116_392#_c_637_n
+ N_A_116_392#_c_638_n N_A_116_392#_c_649_n
+ PM_SKY130_FD_SC_HS__O22A_4%A_116_392#
x_PM_SKY130_FD_SC_HS__O22A_4%A_516_392# N_A_516_392#_M1002_d
+ N_A_516_392#_M1006_s N_A_516_392#_c_665_n N_A_516_392#_c_663_n
+ N_A_516_392#_c_664_n N_A_516_392#_c_673_n
+ PM_SKY130_FD_SC_HS__O22A_4%A_516_392#
x_PM_SKY130_FD_SC_HS__O22A_4%X N_X_M1004_s N_X_M1016_s N_X_M1000_s N_X_M1014_s
+ N_X_c_697_n N_X_c_694_n N_X_c_702_n N_X_c_688_n N_X_c_689_n N_X_c_690_n
+ N_X_c_695_n N_X_c_691_n N_X_c_692_n N_X_c_696_n N_X_c_730_n X
+ PM_SKY130_FD_SC_HS__O22A_4%X
x_PM_SKY130_FD_SC_HS__O22A_4%A_27_136# N_A_27_136#_M1020_d N_A_27_136#_M1018_d
+ N_A_27_136#_M1021_d N_A_27_136#_M1013_s N_A_27_136#_M1023_d
+ N_A_27_136#_c_758_n N_A_27_136#_c_763_n N_A_27_136#_c_759_n
+ N_A_27_136#_c_760_n N_A_27_136#_c_769_n N_A_27_136#_c_772_n
+ N_A_27_136#_c_782_n N_A_27_136#_c_761_n N_A_27_136#_c_784_n
+ PM_SKY130_FD_SC_HS__O22A_4%A_27_136#
x_PM_SKY130_FD_SC_HS__O22A_4%VGND N_VGND_M1020_s N_VGND_M1019_s N_VGND_M1004_d
+ N_VGND_M1007_d N_VGND_M1022_d N_VGND_c_820_n N_VGND_c_821_n N_VGND_c_822_n
+ N_VGND_c_823_n N_VGND_c_824_n N_VGND_c_825_n VGND N_VGND_c_826_n
+ N_VGND_c_827_n N_VGND_c_828_n N_VGND_c_829_n N_VGND_c_830_n N_VGND_c_831_n
+ N_VGND_c_832_n N_VGND_c_833_n N_VGND_c_834_n N_VGND_c_835_n
+ PM_SKY130_FD_SC_HS__O22A_4%VGND
cc_1 VNB N_A2_M1018_g 0.0160698f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=1
cc_2 VNB N_A2_c_116_n 0.0140801f $X=-0.19 $Y=-0.245 $X2=1.425 $Y2=1.395
cc_3 VNB N_A2_c_117_n 0.00161204f $X=-0.19 $Y=-0.245 $X2=1.35 $Y2=1.615
cc_4 VNB N_A2_c_118_n 0.0330027f $X=-0.19 $Y=-0.245 $X2=1.425 $Y2=1.64
cc_5 VNB N_A1_c_172_n 0.00204037f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=2.46
cc_6 VNB N_A1_c_173_n 0.0209762f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=1.45
cc_7 VNB N_A1_M1020_g 0.0365474f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=1
cc_8 VNB N_A1_c_175_n 0.102022f $X=-0.19 $Y=-0.245 $X2=1.425 $Y2=1
cc_9 VNB N_A1_c_176_n 0.0139749f $X=-0.19 $Y=-0.245 $X2=1.455 $Y2=1.885
cc_10 VNB N_A1_c_177_n 0.0172835f $X=-0.19 $Y=-0.245 $X2=1.455 $Y2=2.46
cc_11 VNB N_A1_M1021_g 0.0286707f $X=-0.19 $Y=-0.245 $X2=1.35 $Y2=1.64
cc_12 VNB A1 0.0040904f $X=-0.19 $Y=-0.245 $X2=1.35 $Y2=1.615
cc_13 VNB N_B2_M1013_g 0.0170753f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=2.46
cc_14 VNB N_B2_c_240_n 0.0139501f $X=-0.19 $Y=-0.245 $X2=1.425 $Y2=1.395
cc_15 VNB N_B2_c_241_n 0.00223017f $X=-0.19 $Y=-0.245 $X2=1.455 $Y2=1.64
cc_16 VNB N_B2_c_242_n 0.0312223f $X=-0.19 $Y=-0.245 $X2=1.18 $Y2=1.615
cc_17 VNB N_B1_M1001_g 0.0105364f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=1.45
cc_18 VNB N_B1_c_299_n 0.00571253f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=1
cc_19 VNB N_B1_c_300_n 0.00838574f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=1
cc_20 VNB N_B1_c_301_n 0.0945597f $X=-0.19 $Y=-0.245 $X2=1.425 $Y2=1
cc_21 VNB N_B1_M1023_g 0.0365291f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_B1_c_303_n 0.00577572f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=1.64
cc_23 VNB N_B1_c_304_n 0.0147434f $X=-0.19 $Y=-0.245 $X2=1.18 $Y2=1.615
cc_24 VNB B1 0.0199191f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_B1_c_306_n 0.0426747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_206_392#_M1004_g 0.0255061f $X=-0.19 $Y=-0.245 $X2=1.35 $Y2=1.64
cc_27 VNB N_A_206_392#_M1007_g 0.0224691f $X=-0.19 $Y=-0.245 $X2=1.18 $Y2=1.665
cc_28 VNB N_A_206_392#_M1016_g 0.0224203f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_206_392#_M1022_g 0.0283548f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_206_392#_c_383_n 0.00814028f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_206_392#_c_384_n 0.0042854f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_206_392#_c_385_n 0.00205537f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_206_392#_c_386_n 0.00727975f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_206_392#_c_387_n 0.00290147f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_206_392#_c_388_n 0.00222088f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_206_392#_c_389_n 0.109886f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_VPWR_c_555_n 0.283096f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_X_c_688_n 0.00206666f $X=-0.19 $Y=-0.245 $X2=1.425 $Y2=1.64
cc_39 VNB N_X_c_689_n 0.00357067f $X=-0.19 $Y=-0.245 $X2=1.18 $Y2=1.615
cc_40 VNB N_X_c_690_n 0.00178779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_X_c_691_n 0.00192086f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_X_c_692_n 0.00278817f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB X 0.0183882f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_27_136#_c_758_n 0.0212786f $X=-0.19 $Y=-0.245 $X2=1.35 $Y2=1.64
cc_45 VNB N_A_27_136#_c_759_n 0.0155989f $X=-0.19 $Y=-0.245 $X2=1.425 $Y2=1.64
cc_46 VNB N_A_27_136#_c_760_n 0.00218255f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_27_136#_c_761_n 0.00474714f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_VGND_c_820_n 0.00936742f $X=-0.19 $Y=-0.245 $X2=1.35 $Y2=1.64
cc_49 VNB N_VGND_c_821_n 0.010435f $X=-0.19 $Y=-0.245 $X2=1.455 $Y2=1.64
cc_50 VNB N_VGND_c_822_n 0.0119348f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_VGND_c_823_n 0.00262088f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_VGND_c_824_n 0.0120318f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_VGND_c_825_n 0.0340824f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_VGND_c_826_n 0.0196398f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_VGND_c_827_n 0.0166097f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_VGND_c_828_n 0.069427f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_VGND_c_829_n 0.0172524f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_VGND_c_830_n 0.0152155f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_VGND_c_831_n 0.00506589f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_VGND_c_832_n 0.00506589f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_VGND_c_833_n 0.00632082f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_VGND_c_834_n 0.00604233f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_VGND_c_835_n 0.352068f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VPB N_A2_c_119_n 0.0152201f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=1.885
cc_65 VPB N_A2_c_120_n 0.0155314f $X=-0.19 $Y=1.66 $X2=1.455 $Y2=1.885
cc_66 VPB N_A2_c_117_n 0.00369885f $X=-0.19 $Y=1.66 $X2=1.35 $Y2=1.615
cc_67 VPB N_A2_c_118_n 0.0373936f $X=-0.19 $Y=1.66 $X2=1.425 $Y2=1.64
cc_68 VPB N_A1_c_172_n 0.0114052f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=2.46
cc_69 VPB N_A1_c_181_n 0.0263421f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_70 VPB N_A1_c_177_n 0.034755f $X=-0.19 $Y=1.66 $X2=1.455 $Y2=2.46
cc_71 VPB A1 0.0027167f $X=-0.19 $Y=1.66 $X2=1.35 $Y2=1.615
cc_72 VPB N_B2_c_243_n 0.0151407f $X=-0.19 $Y=1.66 $X2=0.995 $Y2=1
cc_73 VPB N_B2_c_244_n 0.015481f $X=-0.19 $Y=1.66 $X2=1.455 $Y2=1.885
cc_74 VPB N_B2_c_241_n 0.00223017f $X=-0.19 $Y=1.66 $X2=1.455 $Y2=1.64
cc_75 VPB N_B2_c_242_n 0.0353646f $X=-0.19 $Y=1.66 $X2=1.18 $Y2=1.615
cc_76 VPB N_B1_c_300_n 0.00660151f $X=-0.19 $Y=1.66 $X2=0.995 $Y2=1
cc_77 VPB N_B1_c_308_n 0.0224027f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_78 VPB N_B1_c_303_n 0.00808091f $X=-0.19 $Y=1.66 $X2=0.995 $Y2=1.64
cc_79 VPB N_B1_c_310_n 0.0235105f $X=-0.19 $Y=1.66 $X2=1.35 $Y2=1.64
cc_80 VPB N_A_206_392#_c_390_n 0.0169254f $X=-0.19 $Y=1.66 $X2=1.455 $Y2=2.46
cc_81 VPB N_A_206_392#_c_391_n 0.0176723f $X=-0.19 $Y=1.66 $X2=1.35 $Y2=1.615
cc_82 VPB N_A_206_392#_c_392_n 0.0173658f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_83 VPB N_A_206_392#_c_393_n 0.0174177f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_84 VPB N_A_206_392#_c_394_n 0.0124298f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_85 VPB N_A_206_392#_c_395_n 0.00241927f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_86 VPB N_A_206_392#_c_396_n 0.00478819f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_87 VPB N_A_206_392#_c_384_n 0.00509758f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_88 VPB N_A_206_392#_c_398_n 0.00198056f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_89 VPB N_A_206_392#_c_399_n 0.00193086f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_90 VPB N_A_206_392#_c_389_n 0.0606446f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_91 VPB N_VPWR_c_556_n 0.0106521f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=1.64
cc_92 VPB N_VPWR_c_557_n 0.0538358f $X=-0.19 $Y=1.66 $X2=1.35 $Y2=1.64
cc_93 VPB N_VPWR_c_558_n 0.00886797f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_94 VPB N_VPWR_c_559_n 0.0104602f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_95 VPB N_VPWR_c_560_n 0.00993726f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_96 VPB N_VPWR_c_561_n 0.0121909f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_97 VPB N_VPWR_c_562_n 0.061496f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_98 VPB N_VPWR_c_563_n 0.0411572f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_99 VPB N_VPWR_c_564_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_100 VPB N_VPWR_c_565_n 0.021877f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_101 VPB N_VPWR_c_566_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_102 VPB N_VPWR_c_567_n 0.0409981f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_103 VPB N_VPWR_c_568_n 0.0210814f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_104 VPB N_VPWR_c_569_n 0.00631418f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_105 VPB N_VPWR_c_555_n 0.0846214f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_106 VPB N_A_116_392#_c_636_n 0.00470716f $X=-0.19 $Y=1.66 $X2=1.425 $Y2=1
cc_107 VPB N_A_116_392#_c_637_n 0.00502722f $X=-0.19 $Y=1.66 $X2=1.455 $Y2=2.46
cc_108 VPB N_A_116_392#_c_638_n 0.0021839f $X=-0.19 $Y=1.66 $X2=1.115 $Y2=1.58
cc_109 VPB N_A_516_392#_c_663_n 0.00502722f $X=-0.19 $Y=1.66 $X2=1.455 $Y2=1.885
cc_110 VPB N_A_516_392#_c_664_n 0.0021839f $X=-0.19 $Y=1.66 $X2=1.455 $Y2=2.46
cc_111 VPB N_X_c_694_n 0.00290214f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_112 VPB N_X_c_695_n 0.00257348f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_113 VPB N_X_c_696_n 0.00150441f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_114 N_A2_c_118_n N_A1_c_172_n 0.00563966f $X=1.425 $Y=1.64 $X2=0 $Y2=0
cc_115 N_A2_c_117_n N_A1_c_173_n 0.00211029f $X=1.35 $Y=1.615 $X2=0 $Y2=0
cc_116 N_A2_c_118_n N_A1_c_173_n 0.0185231f $X=1.425 $Y=1.64 $X2=0 $Y2=0
cc_117 N_A2_M1018_g N_A1_M1020_g 0.023421f $X=0.995 $Y=1 $X2=0 $Y2=0
cc_118 N_A2_c_119_n N_A1_c_181_n 0.00882862f $X=0.955 $Y=1.885 $X2=0 $Y2=0
cc_119 N_A2_M1018_g N_A1_c_175_n 0.00902846f $X=0.995 $Y=1 $X2=0 $Y2=0
cc_120 N_A2_c_116_n N_A1_c_175_n 0.00904974f $X=1.425 $Y=1.395 $X2=0 $Y2=0
cc_121 N_A2_c_120_n N_A1_c_177_n 0.0271482f $X=1.455 $Y=1.885 $X2=0 $Y2=0
cc_122 N_A2_c_117_n N_A1_c_177_n 4.05682e-19 $X=1.35 $Y=1.615 $X2=0 $Y2=0
cc_123 N_A2_c_118_n N_A1_c_177_n 0.0182639f $X=1.425 $Y=1.64 $X2=0 $Y2=0
cc_124 N_A2_c_116_n N_A1_M1021_g 0.0181273f $X=1.425 $Y=1.395 $X2=0 $Y2=0
cc_125 N_A2_c_118_n N_A1_M1021_g 0.00214132f $X=1.425 $Y=1.64 $X2=0 $Y2=0
cc_126 N_A2_c_117_n A1 0.015639f $X=1.35 $Y=1.615 $X2=0 $Y2=0
cc_127 N_A2_c_118_n A1 0.00152916f $X=1.425 $Y=1.64 $X2=0 $Y2=0
cc_128 N_A2_c_120_n N_A_206_392#_c_394_n 0.0123597f $X=1.455 $Y=1.885 $X2=0
+ $Y2=0
cc_129 N_A2_c_117_n N_A_206_392#_c_394_n 0.00850855f $X=1.35 $Y=1.615 $X2=0
+ $Y2=0
cc_130 N_A2_c_118_n N_A_206_392#_c_394_n 4.58792e-19 $X=1.425 $Y=1.64 $X2=0
+ $Y2=0
cc_131 N_A2_c_119_n N_A_206_392#_c_398_n 9.42736e-19 $X=0.955 $Y=1.885 $X2=0
+ $Y2=0
cc_132 N_A2_c_120_n N_A_206_392#_c_398_n 0.0089121f $X=1.455 $Y=1.885 $X2=0
+ $Y2=0
cc_133 N_A2_c_117_n N_A_206_392#_c_398_n 0.0278981f $X=1.35 $Y=1.615 $X2=0 $Y2=0
cc_134 N_A2_c_118_n N_A_206_392#_c_398_n 0.0028188f $X=1.425 $Y=1.64 $X2=0 $Y2=0
cc_135 N_A2_c_119_n N_VPWR_c_567_n 0.00278257f $X=0.955 $Y=1.885 $X2=0 $Y2=0
cc_136 N_A2_c_120_n N_VPWR_c_567_n 0.00278271f $X=1.455 $Y=1.885 $X2=0 $Y2=0
cc_137 N_A2_c_119_n N_VPWR_c_555_n 0.00354366f $X=0.955 $Y=1.885 $X2=0 $Y2=0
cc_138 N_A2_c_120_n N_VPWR_c_555_n 0.00354798f $X=1.455 $Y=1.885 $X2=0 $Y2=0
cc_139 N_A2_c_119_n N_A_116_392#_c_636_n 0.0110453f $X=0.955 $Y=1.885 $X2=0
+ $Y2=0
cc_140 N_A2_c_120_n N_A_116_392#_c_636_n 6.68308e-19 $X=1.455 $Y=1.885 $X2=0
+ $Y2=0
cc_141 N_A2_c_117_n N_A_116_392#_c_636_n 0.00400453f $X=1.35 $Y=1.615 $X2=0
+ $Y2=0
cc_142 N_A2_c_118_n N_A_116_392#_c_636_n 5.69468e-19 $X=1.425 $Y=1.64 $X2=0
+ $Y2=0
cc_143 N_A2_c_119_n N_A_116_392#_c_637_n 0.0111147f $X=0.955 $Y=1.885 $X2=0
+ $Y2=0
cc_144 N_A2_c_120_n N_A_116_392#_c_637_n 0.0140663f $X=1.455 $Y=1.885 $X2=0
+ $Y2=0
cc_145 N_A2_c_119_n N_A_116_392#_c_638_n 0.00171731f $X=0.955 $Y=1.885 $X2=0
+ $Y2=0
cc_146 N_A2_M1018_g N_A_27_136#_c_758_n 6.53685e-19 $X=0.995 $Y=1 $X2=0 $Y2=0
cc_147 N_A2_M1018_g N_A_27_136#_c_763_n 0.0137182f $X=0.995 $Y=1 $X2=0 $Y2=0
cc_148 N_A2_c_117_n N_A_27_136#_c_763_n 0.0162559f $X=1.35 $Y=1.615 $X2=0 $Y2=0
cc_149 N_A2_c_118_n N_A_27_136#_c_763_n 3.93021e-19 $X=1.425 $Y=1.64 $X2=0 $Y2=0
cc_150 N_A2_M1018_g N_A_27_136#_c_759_n 2.84014e-19 $X=0.995 $Y=1 $X2=0 $Y2=0
cc_151 N_A2_M1018_g N_A_27_136#_c_760_n 5.44783e-19 $X=0.995 $Y=1 $X2=0 $Y2=0
cc_152 N_A2_c_116_n N_A_27_136#_c_760_n 0.00769338f $X=1.425 $Y=1.395 $X2=0
+ $Y2=0
cc_153 N_A2_c_116_n N_A_27_136#_c_769_n 0.00211405f $X=1.425 $Y=1.395 $X2=0
+ $Y2=0
cc_154 N_A2_c_117_n N_A_27_136#_c_769_n 0.0179043f $X=1.35 $Y=1.615 $X2=0 $Y2=0
cc_155 N_A2_c_118_n N_A_27_136#_c_769_n 7.81311e-19 $X=1.425 $Y=1.64 $X2=0 $Y2=0
cc_156 N_A2_c_116_n N_A_27_136#_c_772_n 0.0113587f $X=1.425 $Y=1.395 $X2=0 $Y2=0
cc_157 N_A2_c_117_n N_A_27_136#_c_772_n 0.00946756f $X=1.35 $Y=1.615 $X2=0 $Y2=0
cc_158 N_A2_M1018_g N_VGND_c_820_n 0.00707853f $X=0.995 $Y=1 $X2=0 $Y2=0
cc_159 N_A2_c_116_n N_VGND_c_820_n 4.68906e-19 $X=1.425 $Y=1.395 $X2=0 $Y2=0
cc_160 N_A2_c_116_n N_VGND_c_821_n 0.00335184f $X=1.425 $Y=1.395 $X2=0 $Y2=0
cc_161 N_A2_M1018_g N_VGND_c_835_n 7.45466e-19 $X=0.995 $Y=1 $X2=0 $Y2=0
cc_162 N_A2_c_116_n N_VGND_c_835_n 8.87459e-19 $X=1.425 $Y=1.395 $X2=0 $Y2=0
cc_163 N_A1_c_177_n N_B2_c_241_n 2.98498e-19 $X=1.955 $Y=1.885 $X2=0 $Y2=0
cc_164 A1 N_B2_c_241_n 0.0210577f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_165 N_A1_M1021_g N_B1_M1001_g 0.0205874f $X=1.965 $Y=1 $X2=0 $Y2=0
cc_166 N_A1_c_177_n N_B1_c_299_n 0.0165839f $X=1.955 $Y=1.885 $X2=0 $Y2=0
cc_167 A1 N_B1_c_299_n 0.00239116f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_168 N_A1_c_177_n N_B1_c_300_n 0.00424127f $X=1.955 $Y=1.885 $X2=0 $Y2=0
cc_169 N_A1_c_177_n N_B1_c_308_n 0.0297442f $X=1.955 $Y=1.885 $X2=0 $Y2=0
cc_170 N_A1_c_175_n B1 0.00359425f $X=1.89 $Y=0.235 $X2=0 $Y2=0
cc_171 N_A1_c_175_n N_B1_c_306_n 0.0217819f $X=1.89 $Y=0.235 $X2=0 $Y2=0
cc_172 N_A1_c_177_n N_A_206_392#_c_394_n 0.0197409f $X=1.955 $Y=1.885 $X2=0
+ $Y2=0
cc_173 A1 N_A_206_392#_c_394_n 0.0321683f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_174 N_A1_c_177_n N_A_206_392#_c_398_n 7.18055e-19 $X=1.955 $Y=1.885 $X2=0
+ $Y2=0
cc_175 N_A1_M1021_g N_A_206_392#_c_411_n 3.26818e-19 $X=1.965 $Y=1 $X2=0 $Y2=0
cc_176 N_A1_c_181_n N_VPWR_c_557_n 0.00721488f $X=0.505 $Y=1.885 $X2=0 $Y2=0
cc_177 N_A1_c_177_n N_VPWR_c_558_n 0.00546951f $X=1.955 $Y=1.885 $X2=0 $Y2=0
cc_178 N_A1_c_181_n N_VPWR_c_567_n 0.0044313f $X=0.505 $Y=1.885 $X2=0 $Y2=0
cc_179 N_A1_c_177_n N_VPWR_c_567_n 0.0044313f $X=1.955 $Y=1.885 $X2=0 $Y2=0
cc_180 N_A1_c_181_n N_VPWR_c_555_n 0.00856939f $X=0.505 $Y=1.885 $X2=0 $Y2=0
cc_181 N_A1_c_177_n N_VPWR_c_555_n 0.00854111f $X=1.955 $Y=1.885 $X2=0 $Y2=0
cc_182 N_A1_c_181_n N_A_116_392#_c_636_n 0.0111335f $X=0.505 $Y=1.885 $X2=0
+ $Y2=0
cc_183 N_A1_c_177_n N_A_116_392#_c_637_n 0.00331203f $X=1.955 $Y=1.885 $X2=0
+ $Y2=0
cc_184 N_A1_c_181_n N_A_116_392#_c_638_n 0.00332677f $X=0.505 $Y=1.885 $X2=0
+ $Y2=0
cc_185 N_A1_c_177_n N_A_116_392#_c_649_n 0.00608374f $X=1.955 $Y=1.885 $X2=0
+ $Y2=0
cc_186 N_A1_M1020_g N_A_27_136#_c_758_n 0.0070629f $X=0.495 $Y=1 $X2=0 $Y2=0
cc_187 N_A1_M1020_g N_A_27_136#_c_763_n 0.0150928f $X=0.495 $Y=1 $X2=0 $Y2=0
cc_188 N_A1_c_173_n N_A_27_136#_c_759_n 2.6096e-19 $X=0.495 $Y=1.395 $X2=0 $Y2=0
cc_189 N_A1_M1020_g N_A_27_136#_c_759_n 0.00315149f $X=0.495 $Y=1 $X2=0 $Y2=0
cc_190 N_A1_c_175_n N_A_27_136#_c_760_n 0.00458512f $X=1.89 $Y=0.235 $X2=0 $Y2=0
cc_191 N_A1_M1021_g N_A_27_136#_c_760_n 3.645e-19 $X=1.965 $Y=1 $X2=0 $Y2=0
cc_192 N_A1_M1021_g N_A_27_136#_c_772_n 0.0138807f $X=1.965 $Y=1 $X2=0 $Y2=0
cc_193 A1 N_A_27_136#_c_772_n 0.0290809f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_194 N_A1_c_177_n N_A_27_136#_c_782_n 0.00295011f $X=1.955 $Y=1.885 $X2=0
+ $Y2=0
cc_195 N_A1_M1020_g N_VGND_c_820_n 0.0148276f $X=0.495 $Y=1 $X2=0 $Y2=0
cc_196 N_A1_c_175_n N_VGND_c_820_n 0.0251128f $X=1.89 $Y=0.235 $X2=0 $Y2=0
cc_197 N_A1_c_175_n N_VGND_c_821_n 0.0226067f $X=1.89 $Y=0.235 $X2=0 $Y2=0
cc_198 N_A1_M1021_g N_VGND_c_821_n 0.00705239f $X=1.965 $Y=1 $X2=0 $Y2=0
cc_199 N_A1_c_176_n N_VGND_c_826_n 0.00663676f $X=0.57 $Y=0.235 $X2=0 $Y2=0
cc_200 N_A1_c_175_n N_VGND_c_827_n 0.0167629f $X=1.89 $Y=0.235 $X2=0 $Y2=0
cc_201 N_A1_c_175_n N_VGND_c_828_n 0.00580908f $X=1.89 $Y=0.235 $X2=0 $Y2=0
cc_202 N_A1_c_175_n N_VGND_c_835_n 0.0334926f $X=1.89 $Y=0.235 $X2=0 $Y2=0
cc_203 N_A1_c_176_n N_VGND_c_835_n 0.00954248f $X=0.57 $Y=0.235 $X2=0 $Y2=0
cc_204 N_B2_M1013_g N_B1_M1001_g 0.022149f $X=2.925 $Y=1 $X2=0 $Y2=0
cc_205 N_B2_M1013_g N_B1_c_299_n 0.00305567f $X=2.925 $Y=1 $X2=0 $Y2=0
cc_206 N_B2_c_241_n N_B1_c_299_n 0.00164403f $X=3.34 $Y=1.615 $X2=0 $Y2=0
cc_207 N_B2_c_242_n N_B1_c_299_n 0.0181632f $X=3.43 $Y=1.64 $X2=0 $Y2=0
cc_208 N_B2_c_241_n N_B1_c_300_n 0.00851467f $X=3.34 $Y=1.615 $X2=0 $Y2=0
cc_209 N_B2_c_242_n N_B1_c_300_n 0.00563966f $X=3.43 $Y=1.64 $X2=0 $Y2=0
cc_210 N_B2_c_243_n N_B1_c_308_n 0.0215037f $X=2.955 $Y=1.885 $X2=0 $Y2=0
cc_211 N_B2_M1013_g N_B1_c_301_n 0.00852312f $X=2.925 $Y=1 $X2=0 $Y2=0
cc_212 N_B2_c_240_n N_B1_c_301_n 0.00850324f $X=3.43 $Y=1.395 $X2=0 $Y2=0
cc_213 N_B2_c_240_n N_B1_M1023_g 0.0238464f $X=3.43 $Y=1.395 $X2=0 $Y2=0
cc_214 N_B2_c_242_n N_B1_c_303_n 0.0114955f $X=3.43 $Y=1.64 $X2=0 $Y2=0
cc_215 N_B2_c_244_n N_B1_c_310_n 0.0246307f $X=3.455 $Y=1.885 $X2=0 $Y2=0
cc_216 N_B2_c_241_n N_B1_c_304_n 3.97735e-19 $X=3.34 $Y=1.615 $X2=0 $Y2=0
cc_217 N_B2_c_242_n N_B1_c_304_n 0.0090932f $X=3.43 $Y=1.64 $X2=0 $Y2=0
cc_218 N_B2_M1013_g N_B1_c_306_n 0.00100933f $X=2.925 $Y=1 $X2=0 $Y2=0
cc_219 N_B2_c_243_n N_A_206_392#_c_394_n 0.0151078f $X=2.955 $Y=1.885 $X2=0
+ $Y2=0
cc_220 N_B2_c_241_n N_A_206_392#_c_394_n 0.0407699f $X=3.34 $Y=1.615 $X2=0 $Y2=0
cc_221 N_B2_c_242_n N_A_206_392#_c_394_n 0.00215124f $X=3.43 $Y=1.64 $X2=0 $Y2=0
cc_222 N_B2_c_244_n N_A_206_392#_c_395_n 0.0122431f $X=3.455 $Y=1.885 $X2=0
+ $Y2=0
cc_223 N_B2_c_241_n N_A_206_392#_c_395_n 0.00782149f $X=3.34 $Y=1.615 $X2=0
+ $Y2=0
cc_224 N_B2_c_242_n N_A_206_392#_c_395_n 5.02084e-19 $X=3.43 $Y=1.64 $X2=0 $Y2=0
cc_225 N_B2_c_244_n N_A_206_392#_c_396_n 0.00141334f $X=3.455 $Y=1.885 $X2=0
+ $Y2=0
cc_226 N_B2_c_241_n N_A_206_392#_c_396_n 0.00787349f $X=3.34 $Y=1.615 $X2=0
+ $Y2=0
cc_227 N_B2_c_242_n N_A_206_392#_c_396_n 0.00317596f $X=3.43 $Y=1.64 $X2=0 $Y2=0
cc_228 N_B2_c_241_n N_A_206_392#_c_385_n 0.0151554f $X=3.34 $Y=1.615 $X2=0 $Y2=0
cc_229 N_B2_c_242_n N_A_206_392#_c_385_n 0.00149989f $X=3.43 $Y=1.64 $X2=0 $Y2=0
cc_230 N_B2_c_244_n N_A_206_392#_c_399_n 0.00893175f $X=3.455 $Y=1.885 $X2=0
+ $Y2=0
cc_231 N_B2_c_241_n N_A_206_392#_c_399_n 0.0277622f $X=3.34 $Y=1.615 $X2=0 $Y2=0
cc_232 N_B2_c_242_n N_A_206_392#_c_399_n 0.0079453f $X=3.43 $Y=1.64 $X2=0 $Y2=0
cc_233 N_B2_M1013_g N_A_206_392#_c_411_n 0.00977946f $X=2.925 $Y=1 $X2=0 $Y2=0
cc_234 N_B2_c_240_n N_A_206_392#_c_411_n 0.00856975f $X=3.43 $Y=1.395 $X2=0
+ $Y2=0
cc_235 N_B2_M1013_g N_A_206_392#_c_387_n 3.73061e-19 $X=2.925 $Y=1 $X2=0 $Y2=0
cc_236 N_B2_c_240_n N_A_206_392#_c_387_n 0.00285677f $X=3.43 $Y=1.395 $X2=0
+ $Y2=0
cc_237 N_B2_c_243_n N_VPWR_c_563_n 0.00278257f $X=2.955 $Y=1.885 $X2=0 $Y2=0
cc_238 N_B2_c_244_n N_VPWR_c_563_n 0.00278271f $X=3.455 $Y=1.885 $X2=0 $Y2=0
cc_239 N_B2_c_243_n N_VPWR_c_555_n 0.00354366f $X=2.955 $Y=1.885 $X2=0 $Y2=0
cc_240 N_B2_c_244_n N_VPWR_c_555_n 0.00354798f $X=3.455 $Y=1.885 $X2=0 $Y2=0
cc_241 N_B2_c_243_n N_A_516_392#_c_665_n 0.00769091f $X=2.955 $Y=1.885 $X2=0
+ $Y2=0
cc_242 N_B2_c_244_n N_A_516_392#_c_665_n 5.85804e-19 $X=3.455 $Y=1.885 $X2=0
+ $Y2=0
cc_243 N_B2_c_243_n N_A_516_392#_c_663_n 0.0111147f $X=2.955 $Y=1.885 $X2=0
+ $Y2=0
cc_244 N_B2_c_244_n N_A_516_392#_c_663_n 0.0140663f $X=3.455 $Y=1.885 $X2=0
+ $Y2=0
cc_245 N_B2_c_243_n N_A_516_392#_c_664_n 0.00171731f $X=2.955 $Y=1.885 $X2=0
+ $Y2=0
cc_246 N_B2_c_240_n N_A_27_136#_c_761_n 2.88213e-19 $X=3.43 $Y=1.395 $X2=0 $Y2=0
cc_247 N_B2_M1013_g N_A_27_136#_c_784_n 0.00896296f $X=2.925 $Y=1 $X2=0 $Y2=0
cc_248 N_B2_c_240_n N_A_27_136#_c_784_n 0.00893001f $X=3.43 $Y=1.395 $X2=0 $Y2=0
cc_249 N_B2_c_241_n N_A_27_136#_c_784_n 0.0646255f $X=3.34 $Y=1.615 $X2=0 $Y2=0
cc_250 N_B2_c_242_n N_A_27_136#_c_784_n 0.00393357f $X=3.43 $Y=1.64 $X2=0 $Y2=0
cc_251 N_B2_M1013_g N_VGND_c_835_n 8.87459e-19 $X=2.925 $Y=1 $X2=0 $Y2=0
cc_252 N_B2_c_240_n N_VGND_c_835_n 8.87459e-19 $X=3.43 $Y=1.395 $X2=0 $Y2=0
cc_253 N_B1_c_303_n N_A_206_392#_c_390_n 0.00310411f $X=3.955 $Y=1.795 $X2=0
+ $Y2=0
cc_254 N_B1_c_310_n N_A_206_392#_c_390_n 0.013969f $X=3.955 $Y=1.885 $X2=0 $Y2=0
cc_255 N_B1_c_308_n N_A_206_392#_c_394_n 0.0176709f $X=2.505 $Y=1.885 $X2=0
+ $Y2=0
cc_256 N_B1_c_310_n N_A_206_392#_c_395_n 9.58769e-19 $X=3.955 $Y=1.885 $X2=0
+ $Y2=0
cc_257 N_B1_c_303_n N_A_206_392#_c_396_n 0.00468492f $X=3.955 $Y=1.795 $X2=0
+ $Y2=0
cc_258 N_B1_c_310_n N_A_206_392#_c_396_n 6.07706e-19 $X=3.955 $Y=1.885 $X2=0
+ $Y2=0
cc_259 N_B1_M1023_g N_A_206_392#_c_383_n 0.010793f $X=3.86 $Y=1 $X2=0 $Y2=0
cc_260 N_B1_c_303_n N_A_206_392#_c_384_n 0.0127143f $X=3.955 $Y=1.795 $X2=0
+ $Y2=0
cc_261 N_B1_c_304_n N_A_206_392#_c_384_n 0.00373309f $X=3.915 $Y=1.545 $X2=0
+ $Y2=0
cc_262 N_B1_c_304_n N_A_206_392#_c_385_n 0.00279055f $X=3.915 $Y=1.545 $X2=0
+ $Y2=0
cc_263 N_B1_M1023_g N_A_206_392#_c_386_n 0.00347845f $X=3.86 $Y=1 $X2=0 $Y2=0
cc_264 N_B1_c_310_n N_A_206_392#_c_399_n 7.18055e-19 $X=3.955 $Y=1.885 $X2=0
+ $Y2=0
cc_265 N_B1_M1001_g N_A_206_392#_c_411_n 0.00327726f $X=2.49 $Y=1 $X2=0 $Y2=0
cc_266 N_B1_c_301_n N_A_206_392#_c_411_n 0.00872661f $X=3.785 $Y=0.235 $X2=0
+ $Y2=0
cc_267 B1 N_A_206_392#_c_411_n 0.00304187f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_268 N_B1_c_301_n N_A_206_392#_c_387_n 0.00368783f $X=3.785 $Y=0.235 $X2=0
+ $Y2=0
cc_269 N_B1_M1023_g N_A_206_392#_c_387_n 0.00541004f $X=3.86 $Y=1 $X2=0 $Y2=0
cc_270 N_B1_M1023_g N_A_206_392#_c_388_n 2.39625e-19 $X=3.86 $Y=1 $X2=0 $Y2=0
cc_271 N_B1_c_304_n N_A_206_392#_c_388_n 7.14715e-19 $X=3.915 $Y=1.545 $X2=0
+ $Y2=0
cc_272 N_B1_M1023_g N_A_206_392#_c_389_n 9.06986e-19 $X=3.86 $Y=1 $X2=0 $Y2=0
cc_273 N_B1_c_304_n N_A_206_392#_c_389_n 0.0118639f $X=3.915 $Y=1.545 $X2=0
+ $Y2=0
cc_274 N_B1_c_308_n N_VPWR_c_558_n 0.00546951f $X=2.505 $Y=1.885 $X2=0 $Y2=0
cc_275 N_B1_c_310_n N_VPWR_c_559_n 0.0151574f $X=3.955 $Y=1.885 $X2=0 $Y2=0
cc_276 N_B1_c_308_n N_VPWR_c_563_n 0.0044313f $X=2.505 $Y=1.885 $X2=0 $Y2=0
cc_277 N_B1_c_310_n N_VPWR_c_563_n 0.0044313f $X=3.955 $Y=1.885 $X2=0 $Y2=0
cc_278 N_B1_c_308_n N_VPWR_c_555_n 0.0085368f $X=2.505 $Y=1.885 $X2=0 $Y2=0
cc_279 N_B1_c_310_n N_VPWR_c_555_n 0.00854895f $X=3.955 $Y=1.885 $X2=0 $Y2=0
cc_280 N_B1_c_308_n N_A_516_392#_c_665_n 0.00608374f $X=2.505 $Y=1.885 $X2=0
+ $Y2=0
cc_281 N_B1_c_310_n N_A_516_392#_c_663_n 0.00345428f $X=3.955 $Y=1.885 $X2=0
+ $Y2=0
cc_282 N_B1_c_308_n N_A_516_392#_c_664_n 0.00313312f $X=2.505 $Y=1.885 $X2=0
+ $Y2=0
cc_283 N_B1_c_310_n N_A_516_392#_c_673_n 0.00679059f $X=3.955 $Y=1.885 $X2=0
+ $Y2=0
cc_284 B1 N_A_27_136#_c_782_n 0.021796f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_285 N_B1_c_306_n N_A_27_136#_c_782_n 6.11396e-19 $X=2.445 $Y=0.235 $X2=0
+ $Y2=0
cc_286 N_B1_M1023_g N_A_27_136#_c_761_n 0.00255763f $X=3.86 $Y=1 $X2=0 $Y2=0
cc_287 N_B1_c_304_n N_A_27_136#_c_761_n 0.00331306f $X=3.915 $Y=1.545 $X2=0
+ $Y2=0
cc_288 N_B1_M1001_g N_A_27_136#_c_784_n 0.0148964f $X=2.49 $Y=1 $X2=0 $Y2=0
cc_289 N_B1_M1023_g N_A_27_136#_c_784_n 0.00809366f $X=3.86 $Y=1 $X2=0 $Y2=0
cc_290 B1 N_A_27_136#_c_784_n 0.00434556f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_291 B1 N_VGND_c_821_n 0.0353558f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_292 N_B1_c_306_n N_VGND_c_821_n 7.523e-19 $X=2.445 $Y=0.235 $X2=0 $Y2=0
cc_293 N_B1_c_301_n N_VGND_c_822_n 0.0101887f $X=3.785 $Y=0.235 $X2=0 $Y2=0
cc_294 B1 N_VGND_c_828_n 0.0375355f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_295 N_B1_c_306_n N_VGND_c_828_n 0.0380973f $X=2.445 $Y=0.235 $X2=0 $Y2=0
cc_296 N_B1_c_301_n N_VGND_c_835_n 0.0397068f $X=3.785 $Y=0.235 $X2=0 $Y2=0
cc_297 B1 N_VGND_c_835_n 0.0201025f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_298 N_B1_c_306_n N_VGND_c_835_n 0.00857772f $X=2.445 $Y=0.235 $X2=0 $Y2=0
cc_299 N_A_206_392#_c_394_n N_VPWR_M1009_d 0.00339226f $X=3.065 $Y=2.035 $X2=0
+ $Y2=0
cc_300 N_A_206_392#_c_394_n N_VPWR_c_558_n 0.0232685f $X=3.065 $Y=2.035 $X2=0
+ $Y2=0
cc_301 N_A_206_392#_c_390_n N_VPWR_c_559_n 0.0036738f $X=4.505 $Y=1.765 $X2=0
+ $Y2=0
cc_302 N_A_206_392#_c_395_n N_VPWR_c_559_n 0.00540156f $X=3.675 $Y=2.035 $X2=0
+ $Y2=0
cc_303 N_A_206_392#_c_396_n N_VPWR_c_559_n 0.00593922f $X=3.76 $Y=1.95 $X2=0
+ $Y2=0
cc_304 N_A_206_392#_c_384_n N_VPWR_c_559_n 0.0240754f $X=4.415 $Y=1.595 $X2=0
+ $Y2=0
cc_305 N_A_206_392#_c_391_n N_VPWR_c_560_n 0.0114743f $X=4.99 $Y=1.765 $X2=0
+ $Y2=0
cc_306 N_A_206_392#_c_392_n N_VPWR_c_560_n 0.0117072f $X=5.715 $Y=1.765 $X2=0
+ $Y2=0
cc_307 N_A_206_392#_c_393_n N_VPWR_c_562_n 0.0275367f $X=6.165 $Y=1.765 $X2=0
+ $Y2=0
cc_308 N_A_206_392#_c_389_n N_VPWR_c_562_n 4.87993e-19 $X=6.165 $Y=1.557 $X2=0
+ $Y2=0
cc_309 N_A_206_392#_c_390_n N_VPWR_c_565_n 0.00460063f $X=4.505 $Y=1.765 $X2=0
+ $Y2=0
cc_310 N_A_206_392#_c_391_n N_VPWR_c_565_n 0.00445602f $X=4.99 $Y=1.765 $X2=0
+ $Y2=0
cc_311 N_A_206_392#_c_392_n N_VPWR_c_568_n 0.00445602f $X=5.715 $Y=1.765 $X2=0
+ $Y2=0
cc_312 N_A_206_392#_c_393_n N_VPWR_c_568_n 0.00445602f $X=6.165 $Y=1.765 $X2=0
+ $Y2=0
cc_313 N_A_206_392#_c_390_n N_VPWR_c_555_n 0.0090873f $X=4.505 $Y=1.765 $X2=0
+ $Y2=0
cc_314 N_A_206_392#_c_391_n N_VPWR_c_555_n 0.00860744f $X=4.99 $Y=1.765 $X2=0
+ $Y2=0
cc_315 N_A_206_392#_c_392_n N_VPWR_c_555_n 0.00860417f $X=5.715 $Y=1.765 $X2=0
+ $Y2=0
cc_316 N_A_206_392#_c_393_n N_VPWR_c_555_n 0.00860566f $X=6.165 $Y=1.765 $X2=0
+ $Y2=0
cc_317 N_A_206_392#_c_394_n N_A_116_392#_M1011_s 0.00250873f $X=3.065 $Y=2.035
+ $X2=0 $Y2=0
cc_318 N_A_206_392#_c_398_n N_A_116_392#_c_636_n 0.00682867f $X=1.23 $Y=2.115
+ $X2=0 $Y2=0
cc_319 N_A_206_392#_M1010_d N_A_116_392#_c_637_n 0.00250873f $X=1.03 $Y=1.96
+ $X2=0 $Y2=0
cc_320 N_A_206_392#_c_398_n N_A_116_392#_c_637_n 0.018923f $X=1.23 $Y=2.115
+ $X2=0 $Y2=0
cc_321 N_A_206_392#_c_394_n N_A_116_392#_c_649_n 0.0202249f $X=3.065 $Y=2.035
+ $X2=0 $Y2=0
cc_322 N_A_206_392#_c_394_n N_A_516_392#_M1002_d 0.00197722f $X=3.065 $Y=2.035
+ $X2=-0.19 $Y2=-0.245
cc_323 N_A_206_392#_c_395_n N_A_516_392#_M1006_s 0.0034954f $X=3.675 $Y=2.035
+ $X2=0 $Y2=0
cc_324 N_A_206_392#_c_394_n N_A_516_392#_c_665_n 0.0171814f $X=3.065 $Y=2.035
+ $X2=0 $Y2=0
cc_325 N_A_206_392#_M1005_d N_A_516_392#_c_663_n 0.00250873f $X=3.03 $Y=1.96
+ $X2=0 $Y2=0
cc_326 N_A_206_392#_c_399_n N_A_516_392#_c_663_n 0.018923f $X=3.23 $Y=2.115
+ $X2=0 $Y2=0
cc_327 N_A_206_392#_c_395_n N_A_516_392#_c_673_n 0.0203604f $X=3.675 $Y=2.035
+ $X2=0 $Y2=0
cc_328 N_A_206_392#_c_384_n N_A_516_392#_c_673_n 8.25517e-19 $X=4.415 $Y=1.595
+ $X2=0 $Y2=0
cc_329 N_A_206_392#_c_391_n N_X_c_697_n 4.27055e-19 $X=4.99 $Y=1.765 $X2=0 $Y2=0
cc_330 N_A_206_392#_c_482_p N_X_c_697_n 0.0229494f $X=5.6 $Y=1.515 $X2=0 $Y2=0
cc_331 N_A_206_392#_c_389_n N_X_c_697_n 0.00692546f $X=6.165 $Y=1.557 $X2=0
+ $Y2=0
cc_332 N_A_206_392#_c_390_n N_X_c_694_n 2.77814e-19 $X=4.505 $Y=1.765 $X2=0
+ $Y2=0
cc_333 N_A_206_392#_c_391_n N_X_c_694_n 0.017719f $X=4.99 $Y=1.765 $X2=0 $Y2=0
cc_334 N_A_206_392#_c_391_n N_X_c_702_n 0.013143f $X=4.99 $Y=1.765 $X2=0 $Y2=0
cc_335 N_A_206_392#_c_392_n N_X_c_702_n 0.0132756f $X=5.715 $Y=1.765 $X2=0 $Y2=0
cc_336 N_A_206_392#_c_482_p N_X_c_702_n 0.05685f $X=5.6 $Y=1.515 $X2=0 $Y2=0
cc_337 N_A_206_392#_c_389_n N_X_c_702_n 0.0133942f $X=6.165 $Y=1.557 $X2=0 $Y2=0
cc_338 N_A_206_392#_M1004_g N_X_c_688_n 0.014854f $X=4.93 $Y=0.74 $X2=0 $Y2=0
cc_339 N_A_206_392#_M1007_g N_X_c_688_n 3.97481e-19 $X=5.36 $Y=0.74 $X2=0 $Y2=0
cc_340 N_A_206_392#_c_383_n N_X_c_688_n 0.00719656f $X=4.415 $Y=0.835 $X2=0
+ $Y2=0
cc_341 N_A_206_392#_c_386_n N_X_c_688_n 0.00335992f $X=4.5 $Y=1.35 $X2=0 $Y2=0
cc_342 N_A_206_392#_M1007_g N_X_c_689_n 0.0130932f $X=5.36 $Y=0.74 $X2=0 $Y2=0
cc_343 N_A_206_392#_M1016_g N_X_c_689_n 0.0142578f $X=5.79 $Y=0.74 $X2=0 $Y2=0
cc_344 N_A_206_392#_c_482_p N_X_c_689_n 0.0394261f $X=5.6 $Y=1.515 $X2=0 $Y2=0
cc_345 N_A_206_392#_c_389_n N_X_c_689_n 0.00224206f $X=6.165 $Y=1.557 $X2=0
+ $Y2=0
cc_346 N_A_206_392#_M1004_g N_X_c_690_n 0.00398706f $X=4.93 $Y=0.74 $X2=0 $Y2=0
cc_347 N_A_206_392#_c_386_n N_X_c_690_n 0.00704875f $X=4.5 $Y=1.35 $X2=0 $Y2=0
cc_348 N_A_206_392#_c_482_p N_X_c_690_n 0.0209731f $X=5.6 $Y=1.515 $X2=0 $Y2=0
cc_349 N_A_206_392#_c_389_n N_X_c_690_n 0.00232957f $X=6.165 $Y=1.557 $X2=0
+ $Y2=0
cc_350 N_A_206_392#_c_392_n N_X_c_695_n 0.0172378f $X=5.715 $Y=1.765 $X2=0 $Y2=0
cc_351 N_A_206_392#_c_393_n N_X_c_695_n 0.0101903f $X=6.165 $Y=1.765 $X2=0 $Y2=0
cc_352 N_A_206_392#_M1016_g N_X_c_691_n 3.93409e-19 $X=5.79 $Y=0.74 $X2=0 $Y2=0
cc_353 N_A_206_392#_M1022_g N_X_c_691_n 4.02936e-19 $X=6.22 $Y=0.74 $X2=0 $Y2=0
cc_354 N_A_206_392#_M1016_g N_X_c_692_n 0.00518759f $X=5.79 $Y=0.74 $X2=0 $Y2=0
cc_355 N_A_206_392#_M1022_g N_X_c_692_n 0.00222852f $X=6.22 $Y=0.74 $X2=0 $Y2=0
cc_356 N_A_206_392#_c_482_p N_X_c_692_n 0.00498327f $X=5.6 $Y=1.515 $X2=0 $Y2=0
cc_357 N_A_206_392#_c_389_n N_X_c_692_n 0.00425872f $X=6.165 $Y=1.557 $X2=0
+ $Y2=0
cc_358 N_A_206_392#_c_392_n N_X_c_696_n 0.00177248f $X=5.715 $Y=1.765 $X2=0
+ $Y2=0
cc_359 N_A_206_392#_c_393_n N_X_c_696_n 0.00300856f $X=6.165 $Y=1.765 $X2=0
+ $Y2=0
cc_360 N_A_206_392#_c_482_p N_X_c_696_n 0.0204571f $X=5.6 $Y=1.515 $X2=0 $Y2=0
cc_361 N_A_206_392#_c_389_n N_X_c_696_n 0.0280382f $X=6.165 $Y=1.557 $X2=0 $Y2=0
cc_362 N_A_206_392#_c_392_n N_X_c_730_n 6.21797e-19 $X=5.715 $Y=1.765 $X2=0
+ $Y2=0
cc_363 N_A_206_392#_c_393_n N_X_c_730_n 0.00170116f $X=6.165 $Y=1.765 $X2=0
+ $Y2=0
cc_364 N_A_206_392#_c_389_n N_X_c_730_n 0.00401853f $X=6.165 $Y=1.557 $X2=0
+ $Y2=0
cc_365 N_A_206_392#_M1022_g X 0.013491f $X=6.22 $Y=0.74 $X2=0 $Y2=0
cc_366 N_A_206_392#_c_389_n X 0.0100839f $X=6.165 $Y=1.557 $X2=0 $Y2=0
cc_367 N_A_206_392#_c_411_n N_A_27_136#_M1013_s 0.00612404f $X=3.48 $Y=0.79
+ $X2=0 $Y2=0
cc_368 N_A_206_392#_c_383_n N_A_27_136#_M1023_d 0.00781687f $X=4.415 $Y=0.835
+ $X2=0 $Y2=0
cc_369 N_A_206_392#_c_394_n N_A_27_136#_c_772_n 0.0139844f $X=3.065 $Y=2.035
+ $X2=0 $Y2=0
cc_370 N_A_206_392#_c_384_n N_A_27_136#_c_761_n 0.0249888f $X=4.415 $Y=1.595
+ $X2=0 $Y2=0
cc_371 N_A_206_392#_c_386_n N_A_27_136#_c_761_n 0.0202415f $X=4.5 $Y=1.35 $X2=0
+ $Y2=0
cc_372 N_A_206_392#_c_387_n N_A_27_136#_c_761_n 0.0467438f $X=3.81 $Y=0.79 $X2=0
+ $Y2=0
cc_373 N_A_206_392#_M1001_s N_A_27_136#_c_784_n 0.00365692f $X=2.565 $Y=0.68
+ $X2=0 $Y2=0
cc_374 N_A_206_392#_M1017_d N_A_27_136#_c_784_n 0.00481535f $X=3.505 $Y=0.68
+ $X2=0 $Y2=0
cc_375 N_A_206_392#_c_395_n N_A_27_136#_c_784_n 0.00382984f $X=3.675 $Y=2.035
+ $X2=0 $Y2=0
cc_376 N_A_206_392#_c_384_n N_A_27_136#_c_784_n 0.00343635f $X=4.415 $Y=1.595
+ $X2=0 $Y2=0
cc_377 N_A_206_392#_c_385_n N_A_27_136#_c_784_n 0.0092339f $X=3.845 $Y=1.595
+ $X2=0 $Y2=0
cc_378 N_A_206_392#_c_411_n N_A_27_136#_c_784_n 0.0467438f $X=3.48 $Y=0.79 $X2=0
+ $Y2=0
cc_379 N_A_206_392#_c_383_n N_VGND_M1004_d 0.0041238f $X=4.415 $Y=0.835 $X2=0
+ $Y2=0
cc_380 N_A_206_392#_c_386_n N_VGND_M1004_d 0.00332348f $X=4.5 $Y=1.35 $X2=0
+ $Y2=0
cc_381 N_A_206_392#_M1004_g N_VGND_c_822_n 0.00760845f $X=4.93 $Y=0.74 $X2=0
+ $Y2=0
cc_382 N_A_206_392#_c_383_n N_VGND_c_822_n 0.00997876f $X=4.415 $Y=0.835 $X2=0
+ $Y2=0
cc_383 N_A_206_392#_M1004_g N_VGND_c_823_n 5.04273e-19 $X=4.93 $Y=0.74 $X2=0
+ $Y2=0
cc_384 N_A_206_392#_M1007_g N_VGND_c_823_n 0.00974296f $X=5.36 $Y=0.74 $X2=0
+ $Y2=0
cc_385 N_A_206_392#_M1016_g N_VGND_c_823_n 0.00961487f $X=5.79 $Y=0.74 $X2=0
+ $Y2=0
cc_386 N_A_206_392#_M1022_g N_VGND_c_823_n 4.57434e-19 $X=6.22 $Y=0.74 $X2=0
+ $Y2=0
cc_387 N_A_206_392#_M1016_g N_VGND_c_825_n 5.07085e-19 $X=5.79 $Y=0.74 $X2=0
+ $Y2=0
cc_388 N_A_206_392#_M1022_g N_VGND_c_825_n 0.0119952f $X=6.22 $Y=0.74 $X2=0
+ $Y2=0
cc_389 N_A_206_392#_c_383_n N_VGND_c_828_n 0.00883251f $X=4.415 $Y=0.835 $X2=0
+ $Y2=0
cc_390 N_A_206_392#_c_411_n N_VGND_c_828_n 0.010721f $X=3.48 $Y=0.79 $X2=0 $Y2=0
cc_391 N_A_206_392#_c_387_n N_VGND_c_828_n 0.00578134f $X=3.81 $Y=0.79 $X2=0
+ $Y2=0
cc_392 N_A_206_392#_M1004_g N_VGND_c_829_n 0.00434272f $X=4.93 $Y=0.74 $X2=0
+ $Y2=0
cc_393 N_A_206_392#_M1007_g N_VGND_c_829_n 0.00383152f $X=5.36 $Y=0.74 $X2=0
+ $Y2=0
cc_394 N_A_206_392#_M1016_g N_VGND_c_830_n 0.00383152f $X=5.79 $Y=0.74 $X2=0
+ $Y2=0
cc_395 N_A_206_392#_M1022_g N_VGND_c_830_n 0.00398535f $X=6.22 $Y=0.74 $X2=0
+ $Y2=0
cc_396 N_A_206_392#_M1004_g N_VGND_c_835_n 0.00825283f $X=4.93 $Y=0.74 $X2=0
+ $Y2=0
cc_397 N_A_206_392#_M1007_g N_VGND_c_835_n 0.0075754f $X=5.36 $Y=0.74 $X2=0
+ $Y2=0
cc_398 N_A_206_392#_M1016_g N_VGND_c_835_n 0.0075754f $X=5.79 $Y=0.74 $X2=0
+ $Y2=0
cc_399 N_A_206_392#_M1022_g N_VGND_c_835_n 0.00787535f $X=6.22 $Y=0.74 $X2=0
+ $Y2=0
cc_400 N_A_206_392#_c_383_n N_VGND_c_835_n 0.0172305f $X=4.415 $Y=0.835 $X2=0
+ $Y2=0
cc_401 N_A_206_392#_c_411_n N_VGND_c_835_n 0.0193611f $X=3.48 $Y=0.79 $X2=0
+ $Y2=0
cc_402 N_A_206_392#_c_387_n N_VGND_c_835_n 0.00804027f $X=3.81 $Y=0.79 $X2=0
+ $Y2=0
cc_403 N_VPWR_c_557_n N_A_116_392#_c_636_n 0.0640156f $X=0.28 $Y=2.105 $X2=0
+ $Y2=0
cc_404 N_VPWR_c_558_n N_A_116_392#_c_637_n 0.0119239f $X=2.23 $Y=2.455 $X2=0
+ $Y2=0
cc_405 N_VPWR_c_567_n N_A_116_392#_c_637_n 0.0658792f $X=2.065 $Y=3.33 $X2=0
+ $Y2=0
cc_406 N_VPWR_c_555_n N_A_116_392#_c_637_n 0.0366471f $X=6.48 $Y=3.33 $X2=0
+ $Y2=0
cc_407 N_VPWR_c_557_n N_A_116_392#_c_638_n 0.012272f $X=0.28 $Y=2.105 $X2=0
+ $Y2=0
cc_408 N_VPWR_c_567_n N_A_116_392#_c_638_n 0.0235512f $X=2.065 $Y=3.33 $X2=0
+ $Y2=0
cc_409 N_VPWR_c_555_n N_A_116_392#_c_638_n 0.0126924f $X=6.48 $Y=3.33 $X2=0
+ $Y2=0
cc_410 N_VPWR_c_559_n N_A_516_392#_c_663_n 0.0122955f $X=4.265 $Y=2.015 $X2=0
+ $Y2=0
cc_411 N_VPWR_c_563_n N_A_516_392#_c_663_n 0.0658792f $X=4.1 $Y=3.33 $X2=0 $Y2=0
cc_412 N_VPWR_c_555_n N_A_516_392#_c_663_n 0.0366471f $X=6.48 $Y=3.33 $X2=0
+ $Y2=0
cc_413 N_VPWR_c_558_n N_A_516_392#_c_664_n 0.0119239f $X=2.23 $Y=2.455 $X2=0
+ $Y2=0
cc_414 N_VPWR_c_563_n N_A_516_392#_c_664_n 0.0235512f $X=4.1 $Y=3.33 $X2=0 $Y2=0
cc_415 N_VPWR_c_555_n N_A_516_392#_c_664_n 0.0126924f $X=6.48 $Y=3.33 $X2=0
+ $Y2=0
cc_416 N_VPWR_c_559_n N_A_516_392#_c_673_n 0.0413021f $X=4.265 $Y=2.015 $X2=0
+ $Y2=0
cc_417 N_VPWR_c_559_n N_X_c_694_n 0.0398566f $X=4.265 $Y=2.015 $X2=0 $Y2=0
cc_418 N_VPWR_c_560_n N_X_c_694_n 0.0430465f $X=5.365 $Y=2.355 $X2=0 $Y2=0
cc_419 N_VPWR_c_565_n N_X_c_694_n 0.0145938f $X=5.2 $Y=3.33 $X2=0 $Y2=0
cc_420 N_VPWR_c_555_n N_X_c_694_n 0.0120466f $X=6.48 $Y=3.33 $X2=0 $Y2=0
cc_421 N_VPWR_M1012_d N_X_c_702_n 0.0143236f $X=5.065 $Y=1.84 $X2=0 $Y2=0
cc_422 N_VPWR_c_560_n N_X_c_702_n 0.0266856f $X=5.365 $Y=2.355 $X2=0 $Y2=0
cc_423 N_VPWR_c_560_n N_X_c_695_n 0.0463616f $X=5.365 $Y=2.355 $X2=0 $Y2=0
cc_424 N_VPWR_c_562_n N_X_c_695_n 0.0367744f $X=6.44 $Y=1.985 $X2=0 $Y2=0
cc_425 N_VPWR_c_568_n N_X_c_695_n 0.014552f $X=6.275 $Y=3.33 $X2=0 $Y2=0
cc_426 N_VPWR_c_555_n N_X_c_695_n 0.0119791f $X=6.48 $Y=3.33 $X2=0 $Y2=0
cc_427 N_VPWR_c_562_n N_X_c_696_n 0.00177331f $X=6.44 $Y=1.985 $X2=0 $Y2=0
cc_428 N_VPWR_c_562_n X 0.0148615f $X=6.44 $Y=1.985 $X2=0 $Y2=0
cc_429 N_VPWR_c_557_n N_A_27_136#_c_759_n 0.0096123f $X=0.28 $Y=2.105 $X2=0
+ $Y2=0
cc_430 N_A_116_392#_c_636_n N_A_27_136#_c_763_n 0.00780496f $X=0.73 $Y=2.115
+ $X2=0 $Y2=0
cc_431 N_X_c_689_n N_VGND_M1007_d 0.00197509f $X=5.92 $Y=1.095 $X2=0 $Y2=0
cc_432 N_X_c_688_n N_VGND_c_822_n 0.00865936f $X=5.145 $Y=0.515 $X2=0 $Y2=0
cc_433 N_X_c_688_n N_VGND_c_823_n 0.0164981f $X=5.145 $Y=0.515 $X2=0 $Y2=0
cc_434 N_X_c_689_n N_VGND_c_823_n 0.0140541f $X=5.92 $Y=1.095 $X2=0 $Y2=0
cc_435 N_X_c_691_n N_VGND_c_823_n 0.0164656f $X=6.005 $Y=0.515 $X2=0 $Y2=0
cc_436 N_X_c_691_n N_VGND_c_825_n 0.0254889f $X=6.005 $Y=0.515 $X2=0 $Y2=0
cc_437 X N_VGND_c_825_n 0.0242353f $X=6.395 $Y=1.21 $X2=0 $Y2=0
cc_438 N_X_c_688_n N_VGND_c_829_n 0.0109942f $X=5.145 $Y=0.515 $X2=0 $Y2=0
cc_439 N_X_c_691_n N_VGND_c_830_n 0.00816563f $X=6.005 $Y=0.515 $X2=0 $Y2=0
cc_440 N_X_c_688_n N_VGND_c_835_n 0.00904371f $X=5.145 $Y=0.515 $X2=0 $Y2=0
cc_441 N_X_c_691_n N_VGND_c_835_n 0.0067588f $X=6.005 $Y=0.515 $X2=0 $Y2=0
cc_442 N_A_27_136#_c_763_n N_VGND_M1020_s 0.00726894f $X=1.125 $Y=1.195
+ $X2=-0.19 $Y2=-0.245
cc_443 N_A_27_136#_c_772_n N_VGND_M1019_s 0.00902368f $X=2.045 $Y=1.06 $X2=0
+ $Y2=0
cc_444 N_A_27_136#_c_758_n N_VGND_c_820_n 0.0112968f $X=0.28 $Y=0.825 $X2=0
+ $Y2=0
cc_445 N_A_27_136#_c_763_n N_VGND_c_820_n 0.0209867f $X=1.125 $Y=1.195 $X2=0
+ $Y2=0
cc_446 N_A_27_136#_c_760_n N_VGND_c_820_n 0.0107635f $X=1.21 $Y=0.97 $X2=0 $Y2=0
cc_447 N_A_27_136#_c_760_n N_VGND_c_821_n 0.0108591f $X=1.21 $Y=0.97 $X2=0 $Y2=0
cc_448 N_A_27_136#_c_772_n N_VGND_c_821_n 0.022455f $X=2.045 $Y=1.06 $X2=0 $Y2=0
cc_449 N_A_27_136#_c_758_n N_VGND_c_826_n 0.00625741f $X=0.28 $Y=0.825 $X2=0
+ $Y2=0
cc_450 N_A_27_136#_c_760_n N_VGND_c_827_n 0.0046738f $X=1.21 $Y=0.97 $X2=0 $Y2=0
cc_451 N_A_27_136#_c_758_n N_VGND_c_835_n 0.00964803f $X=0.28 $Y=0.825 $X2=0
+ $Y2=0
cc_452 N_A_27_136#_c_760_n N_VGND_c_835_n 0.00635481f $X=1.21 $Y=0.97 $X2=0
+ $Y2=0
